`define BIT_SIZE 31 
`define EXP_SIZE 7
`define MANT_SIZE 22
`define BIAS 127
`define EXP_SHIFT 4
