
module fpu ( clk, rmode, fpu_op, opa, opb, out, inf, snan, qnan, ine, overflow, 
        underflow, zero, div_by_zero );
  input [1:0] rmode;
  input [2:0] fpu_op;
  input [63:0] opa;
  input [63:0] opb;
  output [63:0] out;
  input clk;
  output inf, snan, qnan, ine, overflow, underflow, zero, div_by_zero;
  wire   inf_d, ind_d, snan_d, opa_nan, opb_nan, opa_00, opb_00, opa_inf,
         opb_inf, opa_dn, opb_dn, sign_fasu, nan_sign_d, result_zero_sign_d,
         sign_fasu_r, sign_mul, sign_exe, inf_mul, sign_mul_r, sign_exe_r,
         exp_ovf_r_0_, N256, N257, N258, N259, N260, N261, N262, N263, N264,
         N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337,
         N340, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374,
         N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385,
         N386, N387, N388, N389, N390, N391, N392, N393, N394, N395, N396,
         N501, N502, N503, N504, N505, N506, N507, N508, N509, N510, N511,
         N512, N513, N514, N515, N516, N517, N518, N519, N520, N521, N522,
         N523, N524, N525, N526, N527, N528, N529, N530, N531, N532, N533,
         N534, N535, N536, N537, N538, N539, N540, N541, N542, N543, N544,
         N545, N546, N547, N548, N549, N550, N551, N552, N553, N554, N555,
         N556, N557, N710, N711, N712, N713, N714, N715, N716, N717, N718,
         N719, N720, N721, N722, N723, N724, N725, N726, N727, N728, N729,
         N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740,
         N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751,
         N752, N753, N754, N755, N756, N757, N758, N759, N760, N761, N762,
         N763, N764, N765, N766, N767, N768, N769, opas_r1, opas_r2, sign,
         N789, fasu_op_r1, N793, N794, N795, N796, N797, N798, N799, N800,
         N801, N802, N803, N804, N805, N806, N807, N808, N809, N810, N811,
         N812, N813, N814, N815, N816, N817, N818, N819, N820, N821, N822,
         N823, N824, N825, N826, N827, N828, N829, N830, N831, N832, N833,
         N834, N835, N836, N837, N838, N839, N840, N841, N842, N843, N844,
         N845, N846, N847, N848, N849, N850, N851, N852, N853, N854, N855,
         N875, N889, N899, N902, N904, N906, N911, N912, opa_nan_r, N913, N923,
         u0_N17, u0_N16, u0_fractb_00, u0_fracta_00, u0_expb_00, u0_expa_00,
         u0_N11, u0_N10, u0_N7, u0_N6, u0_snan_r_b, u0_N5, u0_qnan_r_b,
         u0_snan_r_a, u0_N4, u0_qnan_r_a, u0_infb_f_r, u0_infa_f_r, u0_expb_ff,
         u0_expa_ff, u1_N232, u1_N229, u1_fracta_eq_fractb, u1_N220,
         u1_fracta_lt_fractb, u1_N219, u1_N218, u1_add_r, u1_signb_r,
         u1_signa_r, u1_sign_d, u1_fractb_lt_fracta, u1_adj_op_out_sft_0_,
         u1_adj_op_out_sft_1_, u1_adj_op_out_sft_2_, u1_adj_op_out_sft_3_,
         u1_adj_op_out_sft_4_, u1_adj_op_out_sft_5_, u1_adj_op_out_sft_6_,
         u1_adj_op_out_sft_7_, u1_adj_op_out_sft_8_, u1_adj_op_out_sft_9_,
         u1_adj_op_out_sft_10_, u1_adj_op_out_sft_11_, u1_adj_op_out_sft_12_,
         u1_adj_op_out_sft_13_, u1_adj_op_out_sft_14_, u1_adj_op_out_sft_15_,
         u1_adj_op_out_sft_16_, u1_adj_op_out_sft_17_, u1_adj_op_out_sft_18_,
         u1_adj_op_out_sft_19_, u1_adj_op_out_sft_20_, u1_adj_op_out_sft_21_,
         u1_adj_op_out_sft_22_, u1_adj_op_out_sft_23_, u1_adj_op_out_sft_24_,
         u1_adj_op_out_sft_25_, u1_adj_op_out_sft_26_, u1_adj_op_out_sft_27_,
         u1_adj_op_out_sft_28_, u1_adj_op_out_sft_29_, u1_adj_op_out_sft_30_,
         u1_adj_op_out_sft_31_, u1_adj_op_out_sft_32_, u1_adj_op_out_sft_33_,
         u1_adj_op_out_sft_34_, u1_adj_op_out_sft_35_, u1_adj_op_out_sft_36_,
         u1_adj_op_out_sft_37_, u1_adj_op_out_sft_38_, u1_adj_op_out_sft_39_,
         u1_adj_op_out_sft_40_, u1_adj_op_out_sft_41_, u1_adj_op_out_sft_42_,
         u1_adj_op_out_sft_43_, u1_adj_op_out_sft_44_, u1_adj_op_out_sft_45_,
         u1_adj_op_out_sft_46_, u1_adj_op_out_sft_47_, u1_adj_op_out_sft_48_,
         u1_adj_op_out_sft_49_, u1_adj_op_out_sft_50_, u1_adj_op_out_sft_51_,
         u1_adj_op_out_sft_52_, u1_adj_op_out_sft_53_, u1_adj_op_out_sft_54_,
         u1_adj_op_out_sft_55_, u1_adj_op_0_, u1_adj_op_3_, u1_adj_op_10_,
         u1_adj_op_11_, u1_adj_op_15_, u1_adj_op_16_, u1_adj_op_17_,
         u1_adj_op_20_, u1_adj_op_21_, u1_adj_op_22_, u1_adj_op_27_,
         u1_adj_op_28_, u1_adj_op_32_, u1_adj_op_36_, u1_adj_op_37_,
         u1_adj_op_38_, u1_adj_op_42_, u1_adj_op_44_, u1_adj_op_51_, u1_N62,
         u1_N61, u1_N60, u1_N59, u1_N58, u1_N57, u1_N56, u1_N55, u1_N54,
         u1_N53, u1_N52, u1_N46, u1_exp_large_0_, u1_exp_large_1_,
         u1_exp_large_2_, u1_exp_large_3_, u1_exp_large_4_, u1_exp_large_5_,
         u1_exp_large_6_, u1_exp_large_7_, u1_exp_large_10_, u2_N157, u2_N121,
         u2_sign_d, u2_N114, u2_exp_ovf_d_0_, u2_exp_ovf_d_1_, u2_N86, u2_N85,
         u2_N84, u2_N83, u2_N82, u2_N81, u2_N80, u2_N79, u2_N78, u2_N77,
         u2_N76, u2_N64, u2_N63, u2_N62, u2_N61, u2_N60, u2_N59, u2_N58,
         u2_N57, u2_N56, u2_N55, u2_N54, u2_exp_tmp4_0_, u2_exp_tmp4_1_,
         u2_exp_tmp4_2_, u2_exp_tmp4_3_, u2_exp_tmp4_4_, u2_exp_tmp4_5_,
         u2_exp_tmp4_6_, u2_exp_tmp4_7_, u2_exp_tmp4_8_, u2_exp_tmp4_9_,
         u2_exp_tmp4_10_, u2_exp_tmp3_0_, u2_exp_tmp3_1_, u2_exp_tmp3_2_,
         u2_exp_tmp3_3_, u2_exp_tmp3_4_, u2_exp_tmp3_5_, u2_exp_tmp3_6_,
         u2_exp_tmp3_7_, u2_exp_tmp3_8_, u2_exp_tmp3_9_, u2_exp_tmp3_10_,
         u2_N29, u2_N28, u2_N27, u2_N26, u2_N25, u2_N24, u2_N23, u2_N22,
         u2_N21, u2_N20, u2_N19, u2_N18, u2_N17, u2_N16, u2_N15, u2_N14,
         u2_N13, u2_N12, u2_N11, u2_N10, u2_N9, u2_N8, u2_N7, u2_N6, u3_N116,
         u3_N115, u3_N114, u3_N113, u3_N112, u3_N111, u3_N110, u3_N109,
         u3_N108, u3_N107, u3_N106, u3_N105, u3_N104, u3_N103, u3_N102,
         u3_N101, u3_N100, u3_N99, u3_N98, u3_N97, u3_N96, u3_N95, u3_N94,
         u3_N93, u3_N92, u3_N91, u3_N90, u3_N89, u3_N88, u3_N87, u3_N86,
         u3_N85, u3_N84, u3_N83, u3_N82, u3_N81, u3_N80, u3_N79, u3_N78,
         u3_N77, u3_N76, u3_N75, u3_N74, u3_N73, u3_N72, u3_N71, u3_N70,
         u3_N69, u3_N68, u3_N67, u3_N66, u3_N65, u3_N64, u3_N63, u3_N62,
         u3_N61, u3_N60, u3_N59, u3_N58, u3_N57, u3_N56, u3_N55, u3_N54,
         u3_N53, u3_N52, u3_N51, u3_N50, u3_N49, u3_N48, u3_N47, u3_N46,
         u3_N45, u3_N44, u3_N43, u3_N42, u3_N41, u3_N40, u3_N39, u3_N38,
         u3_N37, u3_N36, u3_N35, u3_N34, u3_N33, u3_N32, u3_N31, u3_N30,
         u3_N29, u3_N28, u3_N27, u3_N26, u3_N25, u3_N24, u3_N23, u3_N22,
         u3_N21, u3_N20, u3_N19, u3_N18, u3_N17, u3_N16, u3_N15, u3_N14,
         u3_N13, u3_N12, u3_N11, u3_N10, u3_N9, u3_N8, u3_N7, u3_N6, u3_N5,
         u3_N4, u3_N3, u5_N105, u5_N104, u5_N103, u5_N102, u5_N101, u5_N100,
         u5_N99, u5_N98, u5_N97, u5_N96, u5_N95, u5_N94, u5_N93, u5_N92,
         u5_N91, u5_N90, u5_N89, u5_N88, u5_N87, u5_N86, u5_N85, u5_N84,
         u5_N83, u5_N82, u5_N81, u5_N80, u5_N79, u5_N78, u5_N77, u5_N76,
         u5_N75, u5_N74, u5_N73, u5_N72, u5_N71, u5_N70, u5_N69, u5_N68,
         u5_N67, u5_N66, u5_N65, u5_N64, u5_N63, u5_N62, u5_N61, u5_N60,
         u5_N59, u5_N58, u5_N57, u5_N56, u5_N55, u5_N54, u5_N53, u5_N52,
         u5_N51, u5_N50, u5_N49, u5_N48, u5_N47, u5_N46, u5_N45, u5_N44,
         u5_N43, u5_N42, u5_N41, u5_N40, u5_N39, u5_N38, u5_N37, u5_N36,
         u5_N35, u5_N34, u5_N33, u5_N32, u5_N31, u5_N30, u5_N29, u5_N28,
         u5_N27, u5_N26, u5_N25, u5_N24, u5_N23, u5_N22, u5_N21, u5_N20,
         u5_N19, u5_N18, u5_N17, u5_N16, u5_N15, u5_N14, u5_N13, u5_N12,
         u5_N11, u5_N10, u5_N9, u5_N8, u5_N7, u5_N6, u5_N5, u5_N4, u5_N3,
         u5_N2, u5_N1, u5_N0, u6_N107, u6_N106, u6_N105, u6_N104, u6_N103,
         u6_N102, u6_N101, u6_N100, u6_N99, u6_N98, u6_N97, u6_N96, u6_N95,
         u6_N94, u6_N93, u6_N92, u6_N91, u6_N90, u6_N89, u6_N88, u6_N87,
         u6_N86, u6_N85, u6_N84, u6_N83, u6_N82, u6_N81, u6_N80, u6_N79,
         u6_N78, u6_N77, u6_N76, u6_N75, u6_N74, u6_N73, u6_N72, u6_N71,
         u6_N70, u6_N69, u6_N68, u6_N67, u6_N66, u6_N65, u6_N64, u6_N63,
         u6_N62, u6_N61, u6_N60, u6_N59, u6_N58, u6_N57, u6_N56, u6_N55,
         u6_N52, u6_N51, u6_N50, u6_N49, u6_N48, u6_N46, u6_N45, u6_N43,
         u6_N40, u6_N39, u6_N37, u6_N36, u6_N35, u6_N33, u6_N32, u6_N31,
         u6_N30, u6_N29, u6_N27, u6_N26, u6_N25, u6_N24, u6_N23, u6_N22,
         u6_N21, u6_N20, u6_N19, u6_N18, u6_N17, u6_N16, u6_N15, u6_N14,
         u6_N13, u6_N12, u6_N11, u6_N10, u6_N9, u6_N8, u6_N7, u6_N6, u6_N5,
         u6_N4, u6_N3, u6_N2, u6_N1, u6_N0, u4_N6917, u4_N6916, u4_N6463,
         u4_N6462, u4_N6461, u4_N6460, u4_N6459, u4_N6457, u4_N6456, u4_N6455,
         u4_N6454, u4_N6280, u4_div_exp2_0_, u4_div_exp2_1_, u4_div_exp2_2_,
         u4_div_exp2_3_, u4_div_exp2_4_, u4_div_exp2_5_, u4_div_exp2_6_,
         u4_div_exp2_7_, u4_div_exp2_8_, u4_div_exp2_9_, u4_div_exp2_10_,
         u4_div_exp1_0_, u4_div_exp1_1_, u4_div_exp1_2_, u4_div_exp1_3_,
         u4_div_exp1_4_, u4_div_exp1_5_, u4_div_exp1_6_, u4_div_exp1_7_,
         u4_div_exp1_8_, u4_div_exp1_9_, u4_div_exp1_10_, u4_fi_ldz_2a_2_,
         u4_fi_ldz_2a_4_, u4_fi_ldz_2a_5_, u4_fi_ldz_2a_6_, u4_ldz_all_0_,
         u4_ldz_all_1_, u4_ldz_all_2_, u4_ldz_all_3_, u4_ldz_all_4_,
         u4_ldz_all_5_, u4_ldz_all_6_, u4_exp_f2i_1_108_, u4_exp_out1_1_,
         u4_exp_out_pl1_0_, u4_exp_out_pl1_1_, u4_exp_out_pl1_2_,
         u4_exp_out_pl1_3_, u4_exp_out_pl1_4_, u4_exp_out_pl1_5_,
         u4_exp_out_pl1_6_, u4_exp_out_pl1_7_, u4_exp_out_pl1_8_,
         u4_exp_out_pl1_9_, u4_exp_out_pl1_10_, u4_fi_ldz_mi1_1_,
         u4_fi_ldz_mi1_3_, u4_fi_ldz_mi1_4_, u4_fi_ldz_mi1_5_,
         u4_fi_ldz_mi1_6_, u4_N6119, u4_N6118, u4_N6117, u4_N6116, u4_N6115,
         u4_N6114, u4_N6113, u4_N6112, u4_N6111, u4_N6110, u4_N6109, u4_N6108,
         u4_N6107, u4_N6106, u4_N6105, u4_N6104, u4_N6103, u4_N6102, u4_N6101,
         u4_N6100, u4_N6099, u4_N6098, u4_N6097, u4_N6096, u4_N6095, u4_N6094,
         u4_N6093, u4_N6092, u4_N6091, u4_N6090, u4_N6089, u4_N6088, u4_N6087,
         u4_N6086, u4_N6085, u4_N6084, u4_N6083, u4_N6082, u4_N6081, u4_N6080,
         u4_N6079, u4_N6078, u4_N6077, u4_N6076, u4_N6075, u4_N6074, u4_N6073,
         u4_N6072, u4_N6071, u4_N6070, u4_N6069, u4_N6068, u4_N6067, u4_N6066,
         u4_N6065, u4_N6064, u4_N6063, u4_N6062, u4_N6061, u4_N6060, u4_N6059,
         u4_N6058, u4_N6057, u4_N6056, u4_N6055, u4_N6054, u4_N6053, u4_N6052,
         u4_N6051, u4_N6050, u4_N6049, u4_N6048, u4_N6047, u4_N6046, u4_N6045,
         u4_N6044, u4_N6043, u4_N6042, u4_N6041, u4_N6040, u4_N6039, u4_N6038,
         u4_N6037, u4_N6036, u4_N6035, u4_N6034, u4_N6033, u4_N6032, u4_N6031,
         u4_N6030, u4_N6029, u4_N6028, u4_N6027, u4_N6026, u4_N6025, u4_N6024,
         u4_N6023, u4_N6022, u4_N6021, u4_N6020, u4_N6019, u4_N6018, u4_N6017,
         u4_N6016, u4_N6015, u4_N6014, u4_N6011, u4_N6010, u4_N6009, u4_N6008,
         u4_N6007, u4_N6006, u4_N6005, u4_N6004, u4_N6003, u4_N6002, u4_N6001,
         u4_N6000, u4_N5999, u4_N5998, u4_N5997, u4_N5996, u4_N5995, u4_N5994,
         u4_N5993, u4_N5992, u4_N5991, u4_N5990, u4_N5989, u4_N5988, u4_N5987,
         u4_N5986, u4_N5985, u4_N5984, u4_N5983, u4_N5982, u4_N5981, u4_N5980,
         u4_N5979, u4_N5978, u4_N5977, u4_N5976, u4_N5975, u4_N5974, u4_N5973,
         u4_N5972, u4_N5971, u4_N5970, u4_N5969, u4_N5968, u4_N5967, u4_N5966,
         u4_N5965, u4_N5964, u4_N5963, u4_N5962, u4_N5961, u4_N5960, u4_N5959,
         u4_N5958, u4_N5957, u4_N5956, u4_N5955, u4_N5954, u4_N5953, u4_N5952,
         u4_N5951, u4_N5950, u4_N5949, u4_N5948, u4_N5947, u4_N5946, u4_N5945,
         u4_N5944, u4_N5943, u4_N5942, u4_N5941, u4_N5940, u4_N5939, u4_N5938,
         u4_N5937, u4_N5936, u4_N5935, u4_N5934, u4_N5933, u4_N5932, u4_N5931,
         u4_N5930, u4_N5929, u4_N5928, u4_N5927, u4_N5926, u4_N5925, u4_N5924,
         u4_N5923, u4_N5922, u4_N5921, u4_N5920, u4_N5919, u4_N5918, u4_N5917,
         u4_N5916, u4_N5915, u4_N5914, u4_N5913, u4_N5912, u4_N5911, u4_N5910,
         u4_N5909, u4_N5908, u4_N5907, u4_N5906, u4_N5904, u4_exp_in_pl1_0_,
         u4_exp_in_pl1_1_, u4_exp_in_pl1_2_, u4_exp_in_pl1_3_,
         u4_exp_in_pl1_4_, u4_exp_in_pl1_5_, u4_exp_in_pl1_6_,
         u4_exp_in_pl1_7_, u4_exp_in_pl1_8_, u4_exp_in_pl1_9_,
         u4_exp_in_pl1_10_, u4_exp_in_pl1_11_, u4_f2i_shft_2_, u4_f2i_shft_3_,
         u4_f2i_shft_6_, u4_f2i_shft_7_, u4_f2i_shft_8_, u4_f2i_shft_9_,
         u4_f2i_shft_10_, u4_exp_in_mi1_1_, u4_exp_in_mi1_2_, u4_exp_in_mi1_3_,
         u4_exp_in_mi1_4_, u4_exp_in_mi1_6_, u4_exp_in_mi1_7_,
         u4_exp_in_mi1_8_, u4_exp_in_mi1_9_, u4_exp_in_mi1_10_,
         u4_exp_in_mi1_11_, u4_fract_out_pl1_0_, u4_fract_out_pl1_1_,
         u4_fract_out_pl1_2_, u4_fract_out_pl1_3_, u4_fract_out_pl1_4_,
         u4_fract_out_pl1_5_, u4_fract_out_pl1_6_, u4_fract_out_pl1_7_,
         u4_fract_out_pl1_8_, u4_fract_out_pl1_9_, u4_fract_out_pl1_10_,
         u4_fract_out_pl1_11_, u4_fract_out_pl1_12_, u4_fract_out_pl1_13_,
         u4_fract_out_pl1_14_, u4_fract_out_pl1_15_, u4_fract_out_pl1_16_,
         u4_fract_out_pl1_17_, u4_fract_out_pl1_18_, u4_fract_out_pl1_19_,
         u4_fract_out_pl1_20_, u4_fract_out_pl1_21_, u4_fract_out_pl1_22_,
         u4_fract_out_pl1_23_, u4_fract_out_pl1_24_, u4_fract_out_pl1_25_,
         u4_fract_out_pl1_26_, u4_fract_out_pl1_27_, u4_fract_out_pl1_28_,
         u4_fract_out_pl1_29_, u4_fract_out_pl1_30_, u4_fract_out_pl1_31_,
         u4_fract_out_pl1_32_, u4_fract_out_pl1_33_, u4_fract_out_pl1_34_,
         u4_fract_out_pl1_35_, u4_fract_out_pl1_36_, u4_fract_out_pl1_37_,
         u4_fract_out_pl1_38_, u4_fract_out_pl1_39_, u4_fract_out_pl1_40_,
         u4_fract_out_pl1_41_, u4_fract_out_pl1_42_, u4_fract_out_pl1_43_,
         u4_fract_out_pl1_44_, u4_fract_out_pl1_45_, u4_fract_out_pl1_46_,
         u4_fract_out_pl1_47_, u4_fract_out_pl1_48_, u4_fract_out_pl1_49_,
         u4_fract_out_pl1_50_, u4_fract_out_pl1_51_, u4_fract_out_pl1_52_,
         u4_exp_next_mi_0_, u4_exp_next_mi_1_, u4_exp_next_mi_2_,
         u4_exp_next_mi_3_, u4_exp_next_mi_4_, u4_exp_next_mi_5_,
         u4_exp_next_mi_6_, u4_exp_next_mi_7_, u4_exp_next_mi_8_,
         u4_exp_next_mi_9_, u4_exp_next_mi_10_, u4_exp_next_mi_11_,
         u4_fract_out_0_, u4_fract_out_1_, u4_fract_out_2_, u4_fract_out_3_,
         u4_fract_out_4_, u4_fract_out_5_, u4_fract_out_6_, u4_fract_out_7_,
         u4_fract_out_8_, u4_fract_out_9_, u4_fract_out_10_, u4_fract_out_11_,
         u4_fract_out_12_, u4_fract_out_13_, u4_fract_out_14_,
         u4_fract_out_15_, u4_fract_out_16_, u4_fract_out_17_,
         u4_fract_out_18_, u4_fract_out_19_, u4_fract_out_20_,
         u4_fract_out_21_, u4_fract_out_22_, u4_fract_out_23_,
         u4_fract_out_24_, u4_fract_out_25_, u4_fract_out_26_,
         u4_fract_out_27_, u4_fract_out_28_, u4_fract_out_29_,
         u4_fract_out_30_, u4_fract_out_31_, u4_fract_out_32_,
         u4_fract_out_33_, u4_fract_out_34_, u4_fract_out_35_,
         u4_fract_out_36_, u4_fract_out_37_, u4_fract_out_38_,
         u4_fract_out_39_, u4_fract_out_40_, u4_fract_out_41_,
         u4_fract_out_42_, u4_fract_out_43_, u4_fract_out_44_,
         u4_fract_out_45_, u4_fract_out_46_, u4_fract_out_47_,
         u4_fract_out_48_, u4_fract_out_49_, u4_fract_out_50_,
         u4_fract_out_51_, u4_exp_out_0_, u4_exp_out_1_, u4_exp_out_2_,
         u4_exp_out_3_, u4_exp_out_4_, u4_exp_out_5_, u4_exp_out_6_,
         u4_exp_out_7_, u4_exp_out_8_, u4_exp_out_9_, u4_exp_out_10_,
         u4_fi_ldz_1_, u4_fi_ldz_2_, u4_fi_ldz_3_, u4_fi_ldz_4_, u4_fi_ldz_5_,
         n2399, n2402, n2404, n2408, n2409, n2412, n2415, n2417, n2419, n2421,
         n2442, n2476, n2477, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3074, n3078,
         n3081, n3096, n3097, n3098, n3100, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3203, n3293, n3294, n3295, n3296, n3341, n3355,
         n3356, n3357, n3358, n3359, n3360, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3378, n3381, n3382, n3385, n3626, n3629, n3636,
         n3638, n3641, n3644, n3650, n3652, n3654, n3662, n3664, n3666, n3675,
         n3677, n3679, n3687, n3689, n3691, n3699, n3702, n3709, n3712, n3715,
         n3717, n3720, n3724, n3727, n3731, n3865, n3888, n3897, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, u4_ldz_dif_9_, u4_ldz_dif_8_, u4_ldz_dif_7_,
         u4_ldz_dif_6_, u4_ldz_dif_5_, u4_ldz_dif_4_, u4_ldz_dif_3_,
         u4_ldz_dif_2_, u4_ldz_dif_1_, u4_ldz_dif_10_, u4_ldz_dif_0_, net33546,
         net33547, net33548, net33549, net33550, net33551, net33552, net33554,
         net33558, net33559, net33561, net33562, net33563, net33564, net33565,
         net33566, net33568, net33569, net33572, net33573, net33575, net33577,
         net33578, net33579, net33581, net33583, net33584, net33585, net33586,
         net33587, net33625, net33641, net33642, net33647, net33648, net34242,
         net34243, net34244, net43686, net44696, net44706, net44770, net44903,
         net45055, net45067, net45071, net57229, net57230, net57232, net57240,
         net57241, net57252, net57260, net57265, net57268, net57276, net57281,
         net57282, net57285, net58419, net58420, net58421, net58422, net58423,
         net58424, net58425, net58427, net58429, net58431, net58433, net58434,
         net58437, net58438, net58440, net58472, net58474, net58475, net58476,
         net58477, net58478, net58479, net58480, net58481, net58482, net58483,
         net58484, net58485, net58486, net58487, net58488, net58489, net58490,
         net58491, net58493, net58494, net58495, net58506, net58517, net58523,
         net58524, net58525, net58526, net58533, net58535, net58537, net58540,
         net58544, net58547, net58550, net58579, net58580, net58581, net58583,
         net58584, net58585, net58586, net58587, net58589, net58590, net58591,
         net58592, net58609, net58613, net58615, net58617, net58623, net58624,
         net58628, net58629, net58631, net58634, net58636, net58638, net58641,
         net58643, net58644, net58645, net58646, net58648, net58649, net58650,
         net58653, net58655, net58658, net58662, net58664, net58666, net58673,
         net58674, net58676, net58681, net58682, net58687, net58688, net58700,
         net58701, net58706, net58707, net58711, net58714, net58716, net58718,
         net58719, net58728, net58733, net58735, net58741, net58743, net58750,
         net58752, net58759, net58762, net58767, net58769, net58771, net58772,
         net58773, net58774, net58775, net58780, net58781, net58783, net58787,
         net58789, net58790, net58792, net58793, net58795, net58799, net58800,
         net58801, net58802, net58803, net58808, net58820, net58825, net58826,
         net58827, net58835, net58886, net58925, net58932, net58935, net58936,
         net58937, net58938, net58939, net58941, net58947, net58951, net58952,
         net58953, net58956, net58957, net58974, net58975, net58976, net58980,
         net58981, net58982, net58983, net58985, net58986, net58987, net58988,
         net58997, net58998, net59008, net59010, net59012, net59013, net59014,
         net59017, net59019, net59020, net59024, net59026, net59027, net59028,
         net59030, net59032, net59054, net59057, net59064, net59070, net59072,
         net59078, net59079, net59081, net59083, net59084, net59087, net59088,
         net59091, net59093, net59097, net59099, net59100, net59107, net59110,
         net59111, net59117, net59120, net59142, net59143, net59144, net59146,
         net59153, net59154, net59155, net59159, net59166, net59169, net59171,
         net59183, net59184, net59189, net59192, net59193, net59195, net59200,
         net59201, net59207, net59208, net59209, net59210, net59212, net59214,
         net59215, net59216, net59217, net59218, net59219, net59224, net59225,
         net59226, net59228, net59231, net59260, net59270, net59275, net59283,
         net59295, net59296, net59309, net59323, net59324, net59328, net59333,
         net59338, net59341, net59347, net59349, net59355, net59356, net59423,
         net59424, net59427, net59430, net59433, net59435, net59442, net59443,
         net59504, net59505, net59506, net59517, net59519, net59531, net59540,
         net59541, net59543, net59551, net59553, net59555, net59563, net59565,
         net59568, net59578, net59579, net59582, net59588, net59589, net59592,
         net59593, net59594, net59600, net59626, net59632, net59635, net59642,
         net59644, net59645, net59651, net59670, net59674, net59678, net59679,
         net59693, net59694, net59695, net59696, net59697, net59698, net59699,
         net59700, net59701, net59717, net59719, net59721, net59722, net59723,
         net59724, net59726, net59731, net59765, net59768, net59785, net59792,
         net59799, net59812, net59826, net59835, net59849, net59850, net59851,
         net59863, net59865, net59868, net59869, net59886, net59888, net59891,
         net59892, net59901, net59910, net59911, net59914, net59917, net59920,
         net59921, net59922, net59923, net59927, net59939, net59941, net59946,
         net59950, net59951, net59952, net59954, net59955, net59956, net59957,
         net59958, net59959, net59962, net59965, net59966, net59974, net59975,
         net59976, net59980, net59982, net59984, net59986, net59988, net59990,
         net59991, net59993, net60002, net60004, net60007, net60008, net60011,
         net60020, net60022, net60026, net60028, net60032, net60038, net60040,
         net60044, net60047, net60048, net60049, net60050, net60051, net60054,
         net60055, net60056, net60057, net60058, net60060, net60062, net60065,
         net60073, net60077, net60078, net60081, net60082, net60084, net60085,
         net60088, net60089, net60090, net60092, net60094, net60095, net60096,
         net60097, net60105, net60107, net60110, net60112, net60113, net60114,
         net60117, net60147, net60150, net60151, net60152, net60153, net60157,
         net60158, net60173, net60174, net60176, net60177, net60178, net60180,
         net60182, net60183, net60185, net60186, net60189, net60190, net60197,
         net60199, net60202, net60204, net60208, net60215, net60219, net60220,
         net60221, net60223, net60230, net60231, net60232, net60237, net60273,
         net60275, net60276, net60279, net60281, net60283, net60284, net60285,
         net60288, net60289, net60290, net60291, net60292, net60293, net60295,
         net60300, net60301, net60302, net60303, net60306, net60308, net60310,
         net60311, net60312, net60314, net60316, net60317, net60318, net60322,
         net60329, net60330, net60340, net60346, net60460, net60461, net60462,
         net60509, net60510, net60536, net60537, net60548, net60549, net60587,
         net60588, net60599, net60600, net60606, net60607, net60610, net60646,
         net60647, net60649, net60652, net60653, net63089, net63085, net63083,
         net63079, net63217, net63293, net63291, net63289, net63287, net63333,
         net63331, net63329, net63327, net63325, net63323, net63321, net63319,
         net63317, net63347, net63343, net63341, net63339, net63335, net63513,
         net63511, net63509, net63507, net63503, net63529, net63527, net63523,
         net63537, net63555, net63553, net63551, net63547, net63545, net63543,
         net63541, net63575, net63573, net63571, net63569, net63567, net63565,
         net63561, net63559, net63587, net63585, net63583, net63579, net63577,
         net66835, net66839, net66851, net66863, net66871, net66870, net66875,
         net66897, net66896, net66895, net66914, net66912, net66911, net66910,
         net66907, net66906, net66905, net66904, net66930, net66929, net66928,
         net87237, net87917, net96080, net58729, net60005, net59999, net59998,
         net59997, net59996, net59995, net59269, net59268, net59267, net59265,
         net59262, net59198, net59124, net60196, net58768, net58426, net58637,
         net58528, net58428, net60345, net60344, net59322, net59339, net59007,
         net58996, net58995, net58993, net58991, net58656, net60286, net60135,
         net58966, net60236, net60235, net60146, net60145, net60144, net60142,
         net60139, net60137, net60136, net60106, net59945, net59307, net59306,
         net59590, net60201, net60192, net59041, net59040, net59039, net58657,
         net60349, net60348, net60159, net59331, net59953, net59591, net58926,
         net59345, net59343, net59311, net58963, net58633, net58630, net60132,
         net60130, net60129, net60128, net60121, net60120, net60119, net59981,
         net66850, net59122, net59121, net59114, net59113, net60611, net59462,
         net59461, net59460, net59448, net59255, net59912, net60324, net60353,
         net60352, net60325, net60131, net59715, net59709, net59708, net59707,
         net59706, net59705, net59704, net59703, net59426, net59243, net59310,
         net59241, net63517, net60193, net58962, net58961, net58958, net58950,
         net58635, net59476, net59475, net59459, net59421, net59352, net59344,
         net59222, net59221, net58779, net58778, net58776, net59315, net59220,
         net60206, net59326, net58846, net58492, net59085, net59082, net59076,
         net59074, net59073, net58990, net58972, net58971, net58970, net58969,
         net58968, net59480, net59479, net59477, net59047, net59046, net59045,
         net59038, net59354, net59353, net59351, net59350, net59342, net59118,
         net58984, net60200, net60194, net60093, net60650, net59669, net59668,
         net59667, net59666, net59566, net58652, net58651, fract_denorm_105_,
         net59278, net60282, net60191, net66927, net60697, net60134, net60133,
         net59840, net59488, net59487, net59478, net59071, net59069, net59068,
         net59053, net59050, net59049, net59048, net59044, net59021, net59009,
         net58994, net59129, net59128, net59127, net59126, net59123, net59031,
         net58973, net59576, net59573, net63221, net60354, net60304, net60111,
         net60006, net59961, net59429, net59428, net60168, net60167, net60164,
         net60163, net60162, net60101, net60100, net60099, net60098, net60086,
         net60053, net59994, net59913, net59449, net59447, n3935, n3934, n3933,
         n3932, n3931, n3930, n3929, n3928, n3927, n3926, n3925, n3924, n3923,
         n3922, n3921, n3920, net60205, net60184, net59973, net59330, net63351,
         net63349, net59503, net59348, net58642, net44995, n3704, net60287,
         net60187, net60072, net59329, net59305, net59261, net59259, net59258,
         net58777, net60696, net60207, net59340, net59337, net59336, net59335,
         net59334, net59332, net59327, net59325, net59321, net59318, net59312,
         net58955, net58948, net59233, net59230, net59132, net59125, net59101,
         net59029, net57231, net59664, net59662, net59641, net59574, net58817,
         net58816, net58818, net58810, net58809, net58805, net58804, net63589,
         net58960, net58959, net58836, net58530, net58529, net58471, net58430,
         net58821, net58791, net66894, net63521, net63515, net60694, net60468,
         net60305, net60155, net60154, net59919, net59918, net58443, net59149,
         net59148, net59145, net59112, net59239, net59237, net59236, net59235,
         net59234, net59194, net59191, net59170, net59161, net63295, net63093,
         net60695, net59042, net59034, net59033, net58989, net58964, net58632,
         net58848, net58847, net58833, net58832, net58831, net58830, net58829,
         net58828, net58823, net58812, net58616, net58610, net58593, net58546,
         net58432, u4_N6458, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4764, n4765, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4790, n4791, n4792, n4793, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4835,
         n4836, n4837, n4838, n4839, n4840, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, u4_sub_473_n14, u4_sub_473_n13, u4_sub_473_n12, u4_sub_473_n11,
         u4_sub_473_n10, u4_sub_473_n9, u4_sub_473_n8, u4_sub_473_n7,
         u4_sub_473_n6, u4_sub_473_n5, u4_sub_473_n4, u4_sub_473_n3,
         u4_sub_473_n2, u4_sub_473_n1, u4_sub_473_carry_1_,
         u4_sub_473_carry_2_, u4_sub_473_carry_3_, u4_sub_473_carry_4_,
         u4_sub_473_carry_5_, u4_sub_473_carry_6_, u4_sub_473_carry_7_,
         u4_sub_473_carry_8_, u4_sub_473_carry_9_, u4_sub_473_carry_10_,
         u4_sub_472_n14, u4_sub_472_n13, u4_sub_472_n12, u4_sub_472_n11,
         u4_sub_472_n10, u4_sub_472_n9, u4_sub_472_n8, u4_sub_472_n7,
         u4_sub_472_n6, u4_sub_472_n5, u4_sub_472_n4, u4_sub_472_n3,
         u4_sub_472_n2, u4_sub_472_n1, u4_sub_472_carry_1_,
         u4_sub_472_carry_2_, u4_sub_472_carry_3_, u4_sub_472_carry_4_,
         u4_sub_472_carry_5_, u4_sub_472_carry_6_, u4_sub_472_carry_7_,
         u4_sub_472_carry_8_, u4_sub_472_carry_9_, u4_sub_472_carry_10_,
         u4_srl_453_n911, u4_srl_453_n910, u4_srl_453_n909, u4_srl_453_n908,
         u4_srl_453_n907, u4_srl_453_n906, u4_srl_453_n905, u4_srl_453_n904,
         u4_srl_453_n903, u4_srl_453_n902, u4_srl_453_n901, u4_srl_453_n900,
         u4_srl_453_n899, u4_srl_453_n898, u4_srl_453_n897, u4_srl_453_n896,
         u4_srl_453_n895, u4_srl_453_n894, u4_srl_453_n893, u4_srl_453_n892,
         u4_srl_453_n891, u4_srl_453_n890, u4_srl_453_n889, u4_srl_453_n888,
         u4_srl_453_n887, u4_srl_453_n886, u4_srl_453_n885, u4_srl_453_n884,
         u4_srl_453_n883, u4_srl_453_n882, u4_srl_453_n881, u4_srl_453_n880,
         u4_srl_453_n879, u4_srl_453_n878, u4_srl_453_n877, u4_srl_453_n876,
         u4_srl_453_n875, u4_srl_453_n874, u4_srl_453_n873, u4_srl_453_n872,
         u4_srl_453_n871, u4_srl_453_n870, u4_srl_453_n869, u4_srl_453_n868,
         u4_srl_453_n867, u4_srl_453_n866, u4_srl_453_n865, u4_srl_453_n864,
         u4_srl_453_n863, u4_srl_453_n862, u4_srl_453_n861, u4_srl_453_n860,
         u4_srl_453_n859, u4_srl_453_n858, u4_srl_453_n857, u4_srl_453_n856,
         u4_srl_453_n855, u4_srl_453_n854, u4_srl_453_n853, u4_srl_453_n852,
         u4_srl_453_n851, u4_srl_453_n850, u4_srl_453_n849, u4_srl_453_n848,
         u4_srl_453_n847, u4_srl_453_n846, u4_srl_453_n845, u4_srl_453_n844,
         u4_srl_453_n843, u4_srl_453_n842, u4_srl_453_n841, u4_srl_453_n840,
         u4_srl_453_n839, u4_srl_453_n838, u4_srl_453_n837, u4_srl_453_n836,
         u4_srl_453_n835, u4_srl_453_n834, u4_srl_453_n833, u4_srl_453_n832,
         u4_srl_453_n831, u4_srl_453_n830, u4_srl_453_n829, u4_srl_453_n828,
         u4_srl_453_n827, u4_srl_453_n826, u4_srl_453_n825, u4_srl_453_n824,
         u4_srl_453_n823, u4_srl_453_n822, u4_srl_453_n821, u4_srl_453_n820,
         u4_srl_453_n819, u4_srl_453_n818, u4_srl_453_n817, u4_srl_453_n816,
         u4_srl_453_n815, u4_srl_453_n814, u4_srl_453_n813, u4_srl_453_n812,
         u4_srl_453_n811, u4_srl_453_n810, u4_srl_453_n809, u4_srl_453_n808,
         u4_srl_453_n807, u4_srl_453_n806, u4_srl_453_n805, u4_srl_453_n804,
         u4_srl_453_n803, u4_srl_453_n802, u4_srl_453_n801, u4_srl_453_n800,
         u4_srl_453_n799, u4_srl_453_n798, u4_srl_453_n797, u4_srl_453_n796,
         u4_srl_453_n795, u4_srl_453_n794, u4_srl_453_n793, u4_srl_453_n792,
         u4_srl_453_n791, u4_srl_453_n790, u4_srl_453_n789, u4_srl_453_n788,
         u4_srl_453_n787, u4_srl_453_n786, u4_srl_453_n785, u4_srl_453_n784,
         u4_srl_453_n783, u4_srl_453_n782, u4_srl_453_n781, u4_srl_453_n780,
         u4_srl_453_n779, u4_srl_453_n778, u4_srl_453_n777, u4_srl_453_n776,
         u4_srl_453_n775, u4_srl_453_n774, u4_srl_453_n773, u4_srl_453_n772,
         u4_srl_453_n771, u4_srl_453_n770, u4_srl_453_n769, u4_srl_453_n768,
         u4_srl_453_n767, u4_srl_453_n766, u4_srl_453_n765, u4_srl_453_n764,
         u4_srl_453_n763, u4_srl_453_n762, u4_srl_453_n761, u4_srl_453_n760,
         u4_srl_453_n759, u4_srl_453_n758, u4_srl_453_n757, u4_srl_453_n756,
         u4_srl_453_n755, u4_srl_453_n754, u4_srl_453_n753, u4_srl_453_n752,
         u4_srl_453_n751, u4_srl_453_n750, u4_srl_453_n749, u4_srl_453_n748,
         u4_srl_453_n747, u4_srl_453_n746, u4_srl_453_n745, u4_srl_453_n744,
         u4_srl_453_n743, u4_srl_453_n742, u4_srl_453_n741, u4_srl_453_n740,
         u4_srl_453_n739, u4_srl_453_n738, u4_srl_453_n737, u4_srl_453_n736,
         u4_srl_453_n735, u4_srl_453_n734, u4_srl_453_n733, u4_srl_453_n732,
         u4_srl_453_n731, u4_srl_453_n730, u4_srl_453_n729, u4_srl_453_n728,
         u4_srl_453_n727, u4_srl_453_n726, u4_srl_453_n725, u4_srl_453_n724,
         u4_srl_453_n723, u4_srl_453_n722, u4_srl_453_n721, u4_srl_453_n720,
         u4_srl_453_n719, u4_srl_453_n718, u4_srl_453_n717, u4_srl_453_n716,
         u4_srl_453_n715, u4_srl_453_n714, u4_srl_453_n713, u4_srl_453_n712,
         u4_srl_453_n711, u4_srl_453_n710, u4_srl_453_n709, u4_srl_453_n708,
         u4_srl_453_n707, u4_srl_453_n706, u4_srl_453_n705, u4_srl_453_n704,
         u4_srl_453_n703, u4_srl_453_n702, u4_srl_453_n701, u4_srl_453_n700,
         u4_srl_453_n699, u4_srl_453_n698, u4_srl_453_n697, u4_srl_453_n696,
         u4_srl_453_n695, u4_srl_453_n694, u4_srl_453_n693, u4_srl_453_n692,
         u4_srl_453_n691, u4_srl_453_n690, u4_srl_453_n689, u4_srl_453_n688,
         u4_srl_453_n687, u4_srl_453_n686, u4_srl_453_n685, u4_srl_453_n684,
         u4_srl_453_n683, u4_srl_453_n682, u4_srl_453_n681, u4_srl_453_n680,
         u4_srl_453_n679, u4_srl_453_n678, u4_srl_453_n677, u4_srl_453_n676,
         u4_srl_453_n675, u4_srl_453_n674, u4_srl_453_n673, u4_srl_453_n672,
         u4_srl_453_n671, u4_srl_453_n670, u4_srl_453_n669, u4_srl_453_n668,
         u4_srl_453_n667, u4_srl_453_n666, u4_srl_453_n665, u4_srl_453_n664,
         u4_srl_453_n663, u4_srl_453_n662, u4_srl_453_n661, u4_srl_453_n660,
         u4_srl_453_n659, u4_srl_453_n658, u4_srl_453_n657, u4_srl_453_n656,
         u4_srl_453_n655, u4_srl_453_n654, u4_srl_453_n653, u4_srl_453_n652,
         u4_srl_453_n651, u4_srl_453_n650, u4_srl_453_n649, u4_srl_453_n648,
         u4_srl_453_n647, u4_srl_453_n646, u4_srl_453_n645, u4_srl_453_n644,
         u4_srl_453_n643, u4_srl_453_n642, u4_srl_453_n641, u4_srl_453_n640,
         u4_srl_453_n639, u4_srl_453_n638, u4_srl_453_n637, u4_srl_453_n636,
         u4_srl_453_n635, u4_srl_453_n634, u4_srl_453_n633, u4_srl_453_n632,
         u4_srl_453_n631, u4_srl_453_n630, u4_srl_453_n629, u4_srl_453_n628,
         u4_srl_453_n627, u4_srl_453_n626, u4_srl_453_n625, u4_srl_453_n624,
         u4_srl_453_n623, u4_srl_453_n622, u4_srl_453_n621, u4_srl_453_n620,
         u4_srl_453_n619, u4_srl_453_n618, u4_srl_453_n617, u4_srl_453_n616,
         u4_srl_453_n615, u4_srl_453_n614, u4_srl_453_n613, u4_srl_453_n612,
         u4_srl_453_n611, u4_srl_453_n610, u4_srl_453_n609, u4_srl_453_n608,
         u4_srl_453_n607, u4_srl_453_n606, u4_srl_453_n605, u4_srl_453_n604,
         u4_srl_453_n603, u4_srl_453_n602, u4_srl_453_n601, u4_srl_453_n600,
         u4_srl_453_n599, u4_srl_453_n598, u4_srl_453_n597, u4_srl_453_n596,
         u4_srl_453_n595, u4_srl_453_n594, u4_srl_453_n593, u4_srl_453_n592,
         u4_srl_453_n591, u4_srl_453_n590, u4_srl_453_n589, u4_srl_453_n588,
         u4_srl_453_n587, u4_srl_453_n586, u4_srl_453_n585, u4_srl_453_n584,
         u4_srl_453_n583, u4_srl_453_n582, u4_srl_453_n581, u4_srl_453_n580,
         u4_srl_453_n579, u4_srl_453_n578, u4_srl_453_n577, u4_srl_453_n576,
         u4_srl_453_n575, u4_srl_453_n574, u4_srl_453_n573, u4_srl_453_n572,
         u4_srl_453_n571, u4_srl_453_n570, u4_srl_453_n569, u4_srl_453_n568,
         u4_srl_453_n567, u4_srl_453_n566, u4_srl_453_n565, u4_srl_453_n564,
         u4_srl_453_n563, u4_srl_453_n562, u4_srl_453_n561, u4_srl_453_n560,
         u4_srl_453_n559, u4_srl_453_n558, u4_srl_453_n557, u4_srl_453_n556,
         u4_srl_453_n555, u4_srl_453_n554, u4_srl_453_n553, u4_srl_453_n552,
         u4_srl_453_n551, u4_srl_453_n550, u4_srl_453_n549, u4_srl_453_n548,
         u4_srl_453_n547, u4_srl_453_n546, u4_srl_453_n545, u4_srl_453_n544,
         u4_srl_453_n543, u4_srl_453_n542, u4_srl_453_n541, u4_srl_453_n540,
         u4_srl_453_n539, u4_srl_453_n538, u4_srl_453_n537, u4_srl_453_n536,
         u4_srl_453_n535, u4_srl_453_n534, u4_srl_453_n533, u4_srl_453_n532,
         u4_srl_453_n531, u4_srl_453_n530, u4_srl_453_n529, u4_srl_453_n528,
         u4_srl_453_n527, u4_srl_453_n526, u4_srl_453_n525, u4_srl_453_n524,
         u4_srl_453_n523, u4_srl_453_n522, u4_srl_453_n521, u4_srl_453_n520,
         u4_srl_453_n519, u4_srl_453_n518, u4_srl_453_n517, u4_srl_453_n516,
         u4_srl_453_n515, u4_srl_453_n514, u4_srl_453_n513, u4_srl_453_n512,
         u4_srl_453_n511, u4_srl_453_n510, u4_srl_453_n509, u4_srl_453_n508,
         u4_srl_453_n507, u4_srl_453_n506, u4_srl_453_n505, u4_srl_453_n504,
         u4_srl_453_n503, u4_srl_453_n502, u4_srl_453_n501, u4_srl_453_n500,
         u4_srl_453_n499, u4_srl_453_n498, u4_srl_453_n497, u4_srl_453_n496,
         u4_srl_453_n495, u4_srl_453_n494, u4_srl_453_n493, u4_srl_453_n492,
         u4_srl_453_n491, u4_srl_453_n490, u4_srl_453_n489, u4_srl_453_n488,
         u4_srl_453_n487, u4_srl_453_n486, u4_srl_453_n485, u4_srl_453_n484,
         u4_srl_453_n483, u4_srl_453_n482, u4_srl_453_n481, u4_srl_453_n480,
         u4_srl_453_n479, u4_srl_453_n478, u4_srl_453_n477, u4_srl_453_n476,
         u4_srl_453_n475, u4_srl_453_n474, u4_srl_453_n473, u4_srl_453_n472,
         u4_srl_453_n471, u4_srl_453_n470, u4_srl_453_n469, u4_srl_453_n468,
         u4_srl_453_n467, u4_srl_453_n466, u4_srl_453_n465, u4_srl_453_n464,
         u4_srl_453_n463, u4_srl_453_n462, u4_srl_453_n461, u4_srl_453_n460,
         u4_srl_453_n459, u4_srl_453_n458, u4_srl_453_n457, u4_srl_453_n456,
         u4_srl_453_n455, u4_srl_453_n454, u4_srl_453_n453, u4_srl_453_n452,
         u4_srl_453_n451, u4_srl_453_n450, u4_srl_453_n449, u4_srl_453_n448,
         u4_srl_453_n447, u4_srl_453_n446, u4_srl_453_n445, u4_srl_453_n444,
         u4_srl_453_n443, u4_srl_453_n442, u4_srl_453_n441, u4_srl_453_n440,
         u4_srl_453_n439, u4_srl_453_n438, u4_srl_453_n437, u4_srl_453_n436,
         u4_srl_453_n435, u4_srl_453_n434, u4_srl_453_n433, u4_srl_453_n432,
         u4_srl_453_n431, u4_srl_453_n430, u4_srl_453_n429, u4_srl_453_n428,
         u4_srl_453_n427, u4_srl_453_n426, u4_srl_453_n425, u4_srl_453_n424,
         u4_srl_453_n423, u4_srl_453_n422, u4_srl_453_n421, u4_srl_453_n420,
         u4_srl_453_n419, u4_srl_453_n418, u4_srl_453_n417, u4_srl_453_n416,
         u4_srl_453_n415, u4_srl_453_n414, u4_srl_453_n413, u4_srl_453_n412,
         u4_srl_453_n411, u4_srl_453_n410, u4_srl_453_n409, u4_srl_453_n408,
         u4_srl_453_n407, u4_srl_453_n406, u4_srl_453_n405, u4_srl_453_n404,
         u4_srl_453_n403, u4_srl_453_n402, u4_srl_453_n401, u4_srl_453_n400,
         u4_srl_453_n399, u4_srl_453_n398, u4_srl_453_n397, u4_srl_453_n396,
         u4_srl_453_n395, u4_srl_453_n394, u4_srl_453_n393, u4_srl_453_n392,
         u4_srl_453_n391, u4_srl_453_n390, u4_srl_453_n389, u4_srl_453_n388,
         u4_srl_453_n387, u4_srl_453_n386, u4_srl_453_n385, u4_srl_453_n384,
         u4_srl_453_n383, u4_srl_453_n382, u4_srl_453_n381, u4_srl_453_n380,
         u4_srl_453_n379, u4_srl_453_n378, u4_srl_453_n377, u4_srl_453_n376,
         u4_srl_453_n375, u4_srl_453_n374, u4_srl_453_n373, u4_srl_453_n372,
         u4_srl_453_n371, u4_srl_453_n370, u4_srl_453_n369, u4_srl_453_n368,
         u4_srl_453_n367, u4_srl_453_n366, u4_srl_453_n365, u4_srl_453_n364,
         u4_srl_453_n363, u4_srl_453_n362, u4_srl_453_n361, u4_srl_453_n360,
         u4_srl_453_n359, u4_srl_453_n358, u4_srl_453_n357, u4_srl_453_n356,
         u4_srl_453_n355, u4_srl_453_n354, u4_srl_453_n353, u4_srl_453_n352,
         u4_srl_453_n351, u4_srl_453_n350, u4_srl_453_n349, u4_srl_453_n348,
         u4_srl_453_n347, u4_srl_453_n346, u4_srl_453_n345, u4_srl_453_n344,
         u4_srl_453_n343, u4_srl_453_n342, u4_srl_453_n341, u4_srl_453_n340,
         u4_srl_453_n339, u4_srl_453_n338, u4_srl_453_n337, u4_srl_453_n336,
         u4_srl_453_n335, u4_srl_453_n334, u4_srl_453_n333, u4_srl_453_n332,
         u4_srl_453_n331, u4_srl_453_n330, u4_srl_453_n329, u4_srl_453_n328,
         u4_srl_453_n327, u4_srl_453_n326, u4_srl_453_n325, u4_srl_453_n324,
         u4_srl_453_n323, u4_srl_453_n322, u4_srl_453_n321, u4_srl_453_n320,
         u4_srl_453_n319, u4_srl_453_n318, u4_srl_453_n317, u4_srl_453_n316,
         u4_srl_453_n315, u4_srl_453_n314, u4_srl_453_n313, u4_srl_453_n312,
         u4_srl_453_n311, u4_srl_453_n310, u4_srl_453_n309, u4_srl_453_n308,
         u4_srl_453_n307, u4_srl_453_n306, u4_srl_453_n305, u4_srl_453_n304,
         u4_srl_453_n303, u4_srl_453_n302, u4_srl_453_n301, u4_srl_453_n300,
         u4_srl_453_n299, u4_srl_453_n298, u4_srl_453_n297, u4_srl_453_n296,
         u4_srl_453_n295, u4_srl_453_n294, u4_srl_453_n293, u4_srl_453_n292,
         u4_srl_453_n291, u4_srl_453_n290, u4_srl_453_n289, u4_srl_453_n288,
         u4_srl_453_n287, u4_srl_453_n286, u4_srl_453_n285, u4_srl_453_n284,
         u4_srl_453_n283, u4_srl_453_n282, u4_srl_453_n281, u4_srl_453_n280,
         u4_srl_453_n279, u4_srl_453_n278, u4_srl_453_n277, u4_srl_453_n276,
         u4_srl_453_n275, u4_srl_453_n274, u4_srl_453_n273, u4_srl_453_n272,
         u4_srl_453_n271, u4_srl_453_n270, u4_srl_453_n269, u4_srl_453_n268,
         u4_srl_453_n267, u4_srl_453_n266, u4_srl_453_n265, u4_srl_453_n264,
         u4_srl_453_n263, u4_srl_453_n262, u4_srl_453_n261, u4_srl_453_n260,
         u4_srl_453_n259, u4_srl_453_n258, u4_srl_453_n257, u4_srl_453_n256,
         u4_srl_453_n255, u4_srl_453_n254, u4_srl_453_n253, u4_srl_453_n252,
         u4_srl_453_n251, u4_srl_453_n250, u4_srl_453_n249, u4_srl_453_n248,
         u4_srl_453_n247, u4_srl_453_n246, u4_srl_453_n245, u4_srl_453_n244,
         u4_srl_453_n243, u4_srl_453_n242, u4_srl_453_n241, u4_srl_453_n240,
         u4_srl_453_n239, u4_srl_453_n238, u4_srl_453_n237, u4_srl_453_n236,
         u4_srl_453_n235, u4_srl_453_n234, u4_srl_453_n233, u4_srl_453_n232,
         u4_srl_453_n231, u4_srl_453_n230, u4_srl_453_n229, u4_srl_453_n228,
         u4_srl_453_n227, u4_srl_453_n226, u4_srl_453_n225, u4_srl_453_n224,
         u4_srl_453_n223, u4_srl_453_n222, u4_srl_453_n221, u4_srl_453_n220,
         u4_srl_453_n219, u4_srl_453_n218, u4_srl_453_n217, u4_srl_453_n216,
         u4_srl_453_n215, u4_srl_453_n214, u4_srl_453_n213, u4_srl_453_n212,
         u4_srl_453_n211, u4_srl_453_n210, u4_srl_453_n209, u4_srl_453_n208,
         u4_srl_453_n207, u4_srl_453_n206, u4_srl_453_n205, u4_srl_453_n204,
         u4_srl_453_n203, u4_srl_453_n202, u4_srl_453_n201, u4_srl_453_n200,
         u4_srl_453_n199, u4_srl_453_n198, u4_srl_453_n197, u4_srl_453_n196,
         u4_srl_453_n195, u4_srl_453_n194, u4_srl_453_n193, u4_srl_453_n192,
         u4_srl_453_n191, u4_srl_453_n190, u4_srl_453_n189, u4_srl_453_n188,
         u4_srl_453_n187, u4_srl_453_n186, u4_srl_453_n185, u4_srl_453_n184,
         u4_srl_453_n183, u4_srl_453_n182, u4_srl_453_n181, u4_srl_453_n180,
         u4_srl_453_n179, u4_srl_453_n178, u4_srl_453_n177, u4_srl_453_n176,
         u4_srl_453_n175, u4_srl_453_n174, u4_srl_453_n173, u4_srl_453_n172,
         u4_srl_453_n171, u4_srl_453_n170, u4_srl_453_n169, u4_srl_453_n168,
         u4_srl_453_n167, u4_srl_453_n166, u4_srl_453_n165, u4_srl_453_n164,
         u4_srl_453_n163, u4_srl_453_n162, u4_srl_453_n161, u4_srl_453_n160,
         u4_srl_453_n159, u4_srl_453_n158, u4_srl_453_n157, u4_srl_453_n156,
         u4_srl_453_n155, u4_srl_453_n154, u4_srl_453_n153, u4_srl_453_n152,
         u4_srl_453_n151, u4_srl_453_n150, u4_srl_453_n149, u4_srl_453_n148,
         u4_srl_453_n147, u4_srl_453_n146, u4_srl_453_n145, u4_srl_453_n144,
         u4_srl_453_n143, u4_srl_453_n142, u4_srl_453_n141, u4_srl_453_n140,
         u4_srl_453_n139, u4_srl_453_n138, u4_srl_453_n137, u4_srl_453_n136,
         u4_srl_453_n135, u4_srl_453_n134, u4_srl_453_n133, u4_srl_453_n132,
         u4_srl_453_n131, u4_srl_453_n130, u4_srl_453_n129, u4_srl_453_n128,
         u4_srl_453_n127, u4_srl_453_n126, u4_srl_453_n125, u4_srl_453_n124,
         u4_srl_453_n123, u4_srl_453_n122, u4_srl_453_n121, u4_srl_453_n120,
         u4_srl_453_n119, u4_srl_453_n118, u4_srl_453_n117, u4_srl_453_n116,
         u4_srl_453_n115, u4_srl_453_n114, u4_srl_453_n113, u4_srl_453_n112,
         u4_srl_453_n111, u4_srl_453_n110, u4_srl_453_n109, u4_srl_453_n108,
         u4_srl_453_n107, u4_srl_453_n106, u4_srl_453_n105, u4_srl_453_n104,
         u4_srl_453_n103, u4_srl_453_n102, u4_srl_453_n101, u4_srl_453_n100,
         u4_srl_453_n99, u4_srl_453_n98, u4_srl_453_n97, u4_srl_453_n96,
         u4_srl_453_n95, u4_srl_453_n94, u4_srl_453_n93, u4_srl_453_n92,
         u4_srl_453_n91, u4_srl_453_n90, u4_srl_453_n89, u4_srl_453_n88,
         u4_srl_453_n87, u4_srl_453_n86, u4_srl_453_n85, u4_srl_453_n84,
         u4_srl_453_n83, u4_srl_453_n82, u4_srl_453_n81, u4_srl_453_n80,
         u4_srl_453_n79, u4_srl_453_n78, u4_srl_453_n77, u4_srl_453_n76,
         u4_srl_453_n75, u4_srl_453_n74, u4_srl_453_n73, u4_srl_453_n72,
         u4_srl_453_n71, u4_srl_453_n70, u4_srl_453_n69, u4_srl_453_n68,
         u4_srl_453_n67, u4_srl_453_n66, u4_srl_453_n65, u4_srl_453_n64,
         u4_srl_453_n63, u4_srl_453_n62, u4_srl_453_n61, u4_srl_453_n60,
         u4_srl_453_n59, u4_srl_453_n58, u4_srl_453_n57, u4_srl_453_n56,
         u4_srl_453_n55, u4_srl_453_n54, u4_srl_453_n53, u4_srl_453_n52,
         u4_srl_453_n51, u4_srl_453_n50, u4_srl_453_n49, u4_srl_453_n48,
         u4_srl_453_n47, u4_srl_453_n46, u4_srl_453_n45, u4_srl_453_n44,
         u4_srl_453_n43, u4_srl_453_n42, u4_srl_453_n41, u4_srl_453_n40,
         u4_srl_453_n39, u4_srl_453_n38, u4_srl_453_n37, u4_srl_453_n36,
         u4_srl_453_n35, u4_srl_453_n34, u4_srl_453_n33, u4_srl_453_n32,
         u4_srl_453_n31, u4_srl_453_n30, u4_srl_453_n29, u4_srl_453_n28,
         u4_srl_453_n27, u4_srl_453_n26, u4_srl_453_n25, u4_srl_453_n24,
         u4_srl_453_n23, u4_srl_453_n22, u4_srl_453_n21, u4_srl_453_n20,
         u4_srl_453_n19, u4_srl_453_n18, u4_srl_453_n17, u4_srl_453_n16,
         u4_srl_453_n15, u4_srl_453_n14, u4_srl_453_n13, u4_srl_453_n12,
         u4_srl_453_n11, u4_srl_453_n10, u4_srl_453_n9, u4_srl_453_n8,
         u4_srl_453_n7, u4_srl_453_n6, u4_srl_453_n5, u4_srl_453_n4,
         u4_srl_453_n3, u4_srl_453_n2, u4_srl_453_n1, u4_sll_482_n59,
         u4_sll_482_n58, u4_sll_482_n57, u4_sll_482_n56, u4_sll_482_n55,
         u4_sll_482_n54, u4_sll_482_n53, u4_sll_482_n52, u4_sll_482_n51,
         u4_sll_482_n50, u4_sll_482_n49, u4_sll_482_n48, u4_sll_482_n47,
         u4_sll_482_n46, u4_sll_482_n45, u4_sll_482_n44, u4_sll_482_n43,
         u4_sll_482_n42, u4_sll_482_n41, u4_sll_482_n40, u4_sll_482_n39,
         u4_sll_482_n38, u4_sll_482_n37, u4_sll_482_n36, u4_sll_482_n35,
         u4_sll_482_n34, u4_sll_482_n33, u4_sll_482_n32, u4_sll_482_n31,
         u4_sll_482_n30, u4_sll_482_n29, u4_sll_482_n28, u4_sll_482_n27,
         u4_sll_482_n26, u4_sll_482_n25, u4_sll_482_n24, u4_sll_482_n23,
         u4_sll_482_n22, u4_sll_482_n21, u4_sll_482_n20, u4_sll_482_n19,
         u4_sll_482_n18, u4_sll_482_n17, u4_sll_482_n16, u4_sll_482_n15,
         u4_sll_482_n14, u4_sll_482_n13, u4_sll_482_n12, u4_sll_482_n11,
         u4_sll_482_n10, u4_sll_482_n9, u4_sll_482_n8, u4_sll_482_n7,
         u4_sll_482_n6, u4_sll_482_n5, u4_sll_482_n4, u4_sll_482_n3,
         u4_sll_482_n2, u4_sll_482_n1, u4_sll_482_ML_int_7__108_,
         u4_sll_482_ML_int_6__44_, u4_sll_482_ML_int_6__108_,
         u4_sll_482_ML_int_5__12_, u4_sll_482_ML_int_5__44_,
         u4_sll_482_ML_int_5__76_, u4_sll_482_ML_int_5__108_,
         u4_sll_482_ML_int_4__12_, u4_sll_482_ML_int_4__28_,
         u4_sll_482_ML_int_4__44_, u4_sll_482_ML_int_4__60_,
         u4_sll_482_ML_int_4__76_, u4_sll_482_ML_int_4__92_,
         u4_sll_482_ML_int_4__108_, u4_sll_482_ML_int_3__4_,
         u4_sll_482_ML_int_3__12_, u4_sll_482_ML_int_3__20_,
         u4_sll_482_ML_int_3__28_, u4_sll_482_ML_int_3__36_,
         u4_sll_482_ML_int_3__44_, u4_sll_482_ML_int_3__52_,
         u4_sll_482_ML_int_3__60_, u4_sll_482_ML_int_3__68_,
         u4_sll_482_ML_int_3__76_, u4_sll_482_ML_int_3__84_,
         u4_sll_482_ML_int_3__92_, u4_sll_482_ML_int_3__100_,
         u4_sll_482_ML_int_3__108_, u4_sll_482_ML_int_2__4_,
         u4_sll_482_ML_int_2__8_, u4_sll_482_ML_int_2__12_,
         u4_sll_482_ML_int_2__16_, u4_sll_482_ML_int_2__20_,
         u4_sll_482_ML_int_2__24_, u4_sll_482_ML_int_2__28_,
         u4_sll_482_ML_int_2__32_, u4_sll_482_ML_int_2__36_,
         u4_sll_482_ML_int_2__40_, u4_sll_482_ML_int_2__44_,
         u4_sll_482_ML_int_2__48_, u4_sll_482_ML_int_2__52_,
         u4_sll_482_ML_int_2__56_, u4_sll_482_ML_int_2__60_,
         u4_sll_482_ML_int_2__64_, u4_sll_482_ML_int_2__68_,
         u4_sll_482_ML_int_2__72_, u4_sll_482_ML_int_2__76_,
         u4_sll_482_ML_int_2__80_, u4_sll_482_ML_int_2__84_,
         u4_sll_482_ML_int_2__88_, u4_sll_482_ML_int_2__92_,
         u4_sll_482_ML_int_2__96_, u4_sll_482_ML_int_2__100_,
         u4_sll_482_ML_int_2__104_, u4_sll_482_ML_int_2__108_,
         u4_sll_482_ML_int_1__0_, u4_sll_482_ML_int_1__2_,
         u4_sll_482_ML_int_1__4_, u4_sll_482_ML_int_1__6_,
         u4_sll_482_ML_int_1__8_, u4_sll_482_ML_int_1__10_,
         u4_sll_482_ML_int_1__12_, u4_sll_482_ML_int_1__14_,
         u4_sll_482_ML_int_1__16_, u4_sll_482_ML_int_1__18_,
         u4_sll_482_ML_int_1__20_, u4_sll_482_ML_int_1__22_,
         u4_sll_482_ML_int_1__24_, u4_sll_482_ML_int_1__26_,
         u4_sll_482_ML_int_1__28_, u4_sll_482_ML_int_1__30_,
         u4_sll_482_ML_int_1__32_, u4_sll_482_ML_int_1__34_,
         u4_sll_482_ML_int_1__36_, u4_sll_482_ML_int_1__38_,
         u4_sll_482_ML_int_1__40_, u4_sll_482_ML_int_1__42_,
         u4_sll_482_ML_int_1__44_, u4_sll_482_ML_int_1__46_,
         u4_sll_482_ML_int_1__48_, u4_sll_482_ML_int_1__50_,
         u4_sll_482_ML_int_1__52_, u4_sll_482_ML_int_1__54_,
         u4_sll_482_ML_int_1__56_, u4_sll_482_ML_int_1__58_,
         u4_sll_482_ML_int_1__60_, u4_sll_482_ML_int_1__62_,
         u4_sll_482_ML_int_1__64_, u4_sll_482_ML_int_1__66_,
         u4_sll_482_ML_int_1__68_, u4_sll_482_ML_int_1__70_,
         u4_sll_482_ML_int_1__72_, u4_sll_482_ML_int_1__74_,
         u4_sll_482_ML_int_1__76_, u4_sll_482_ML_int_1__78_,
         u4_sll_482_ML_int_1__80_, u4_sll_482_ML_int_1__82_,
         u4_sll_482_ML_int_1__84_, u4_sll_482_ML_int_1__86_,
         u4_sll_482_ML_int_1__88_, u4_sll_482_ML_int_1__90_,
         u4_sll_482_ML_int_1__92_, u4_sll_482_ML_int_1__94_,
         u4_sll_482_ML_int_1__96_, u4_sll_482_ML_int_1__98_,
         u4_sll_482_ML_int_1__100_, u4_sll_482_ML_int_1__102_,
         u4_sll_482_ML_int_1__104_, u4_sll_482_ML_int_1__106_,
         u4_sll_482_ML_int_1__108_, u4_sll_482_temp_int_SH_0_,
         u4_sll_482_temp_int_SH_2_, u4_sll_482_temp_int_SH_3_, u4_add_489_n2,
         u4_add_489__UDW__88324_net67898, u4_add_489_carry_1_,
         u4_add_489_carry_2_, u4_add_489_carry_3_, u4_add_489_carry_4_,
         u4_add_489_carry_5_, u4_add_489__UDW__88324_net67896,
         u4_add_489__UDW__88319_net67884, u4_add_494_n7, u4_add_494_n6,
         u4_add_494_n3, u4_add_494_carry_2_, u4_add_494_carry_3_,
         u4_add_494_carry_4_, u4_add_494_carry_5_, u4_add_494_carry_6_,
         u4_add_494_carry_7_, u4_add_494_carry_8_, u4_add_494_carry_9_,
         u4_add_494_carry_10_, u3_sub_63_n59, u3_sub_63_n58, u3_sub_63_n57,
         u3_sub_63_n56, u3_sub_63_n55, u3_sub_63_n54, u3_sub_63_n53,
         u3_sub_63_n52, u3_sub_63_n51, u3_sub_63_n50, u3_sub_63_n49,
         u3_sub_63_n48, u3_sub_63_n47, u3_sub_63_n46, u3_sub_63_n45,
         u3_sub_63_n44, u3_sub_63_n43, u3_sub_63_n42, u3_sub_63_n41,
         u3_sub_63_n40, u3_sub_63_n39, u3_sub_63_n38, u3_sub_63_n37,
         u3_sub_63_n36, u3_sub_63_n35, u3_sub_63_n34, u3_sub_63_n33,
         u3_sub_63_n32, u3_sub_63_n31, u3_sub_63_n30, u3_sub_63_n29,
         u3_sub_63_n28, u3_sub_63_n27, u3_sub_63_n26, u3_sub_63_n25,
         u3_sub_63_n24, u3_sub_63_n23, u3_sub_63_n22, u3_sub_63_n21,
         u3_sub_63_n20, u3_sub_63_n19, u3_sub_63_n18, u3_sub_63_n17,
         u3_sub_63_n16, u3_sub_63_n15, u3_sub_63_n14, u3_sub_63_n13,
         u3_sub_63_n12, u3_sub_63_n11, u3_sub_63_n10, u3_sub_63_n9,
         u3_sub_63_n8, u3_sub_63_n7, u3_sub_63_n6, u3_sub_63_n5, u3_sub_63_n4,
         u3_sub_63_n2, u3_sub_63_n1, u3_add_63_n2, u2_add_115_n2,
         u2_sub_115_n14, u2_sub_115_n13, u2_sub_115_n12, u2_sub_115_n11,
         u2_sub_115_n10, u2_sub_115_n9, u2_sub_115_n8, u2_sub_115_n7,
         u2_sub_115_n6, u2_sub_115_n5, u2_sub_115_n4, u2_sub_115_n2,
         u2_sub_115_n1, u1_srl_151_n375, u1_srl_151_n374, u1_srl_151_n373,
         u1_srl_151_n372, u1_srl_151_n371, u1_srl_151_n370, u1_srl_151_n369,
         u1_srl_151_n368, u1_srl_151_n367, u1_srl_151_n366, u1_srl_151_n365,
         u1_srl_151_n364, u1_srl_151_n363, u1_srl_151_n362, u1_srl_151_n361,
         u1_srl_151_n360, u1_srl_151_n359, u1_srl_151_n358, u1_srl_151_n357,
         u1_srl_151_n356, u1_srl_151_n355, u1_srl_151_n354, u1_srl_151_n353,
         u1_srl_151_n352, u1_srl_151_n351, u1_srl_151_n350, u1_srl_151_n349,
         u1_srl_151_n348, u1_srl_151_n347, u1_srl_151_n346, u1_srl_151_n345,
         u1_srl_151_n344, u1_srl_151_n343, u1_srl_151_n342, u1_srl_151_n341,
         u1_srl_151_n340, u1_srl_151_n339, u1_srl_151_n338, u1_srl_151_n337,
         u1_srl_151_n336, u1_srl_151_n335, u1_srl_151_n334, u1_srl_151_n333,
         u1_srl_151_n332, u1_srl_151_n331, u1_srl_151_n330, u1_srl_151_n329,
         u1_srl_151_n328, u1_srl_151_n327, u1_srl_151_n326, u1_srl_151_n325,
         u1_srl_151_n324, u1_srl_151_n323, u1_srl_151_n322, u1_srl_151_n321,
         u1_srl_151_n320, u1_srl_151_n319, u1_srl_151_n318, u1_srl_151_n317,
         u1_srl_151_n316, u1_srl_151_n315, u1_srl_151_n314, u1_srl_151_n313,
         u1_srl_151_n312, u1_srl_151_n311, u1_srl_151_n310, u1_srl_151_n309,
         u1_srl_151_n308, u1_srl_151_n307, u1_srl_151_n306, u1_srl_151_n305,
         u1_srl_151_n304, u1_srl_151_n303, u1_srl_151_n302, u1_srl_151_n301,
         u1_srl_151_n300, u1_srl_151_n299, u1_srl_151_n298, u1_srl_151_n297,
         u1_srl_151_n296, u1_srl_151_n295, u1_srl_151_n294, u1_srl_151_n293,
         u1_srl_151_n292, u1_srl_151_n291, u1_srl_151_n290, u1_srl_151_n289,
         u1_srl_151_n288, u1_srl_151_n287, u1_srl_151_n286, u1_srl_151_n285,
         u1_srl_151_n284, u1_srl_151_n283, u1_srl_151_n282, u1_srl_151_n281,
         u1_srl_151_n280, u1_srl_151_n279, u1_srl_151_n278, u1_srl_151_n277,
         u1_srl_151_n276, u1_srl_151_n275, u1_srl_151_n274, u1_srl_151_n273,
         u1_srl_151_n272, u1_srl_151_n271, u1_srl_151_n270, u1_srl_151_n269,
         u1_srl_151_n268, u1_srl_151_n267, u1_srl_151_n266, u1_srl_151_n265,
         u1_srl_151_n264, u1_srl_151_n263, u1_srl_151_n262, u1_srl_151_n261,
         u1_srl_151_n260, u1_srl_151_n259, u1_srl_151_n258, u1_srl_151_n257,
         u1_srl_151_n256, u1_srl_151_n255, u1_srl_151_n254, u1_srl_151_n253,
         u1_srl_151_n252, u1_srl_151_n251, u1_srl_151_n250, u1_srl_151_n249,
         u1_srl_151_n248, u1_srl_151_n247, u1_srl_151_n246, u1_srl_151_n245,
         u1_srl_151_n244, u1_srl_151_n243, u1_srl_151_n242, u1_srl_151_n241,
         u1_srl_151_n240, u1_srl_151_n239, u1_srl_151_n238, u1_srl_151_n237,
         u1_srl_151_n236, u1_srl_151_n235, u1_srl_151_n234, u1_srl_151_n233,
         u1_srl_151_n232, u1_srl_151_n231, u1_srl_151_n230, u1_srl_151_n229,
         u1_srl_151_n228, u1_srl_151_n227, u1_srl_151_n226, u1_srl_151_n225,
         u1_srl_151_n224, u1_srl_151_n223, u1_srl_151_n222, u1_srl_151_n221,
         u1_srl_151_n220, u1_srl_151_n219, u1_srl_151_n218, u1_srl_151_n217,
         u1_srl_151_n216, u1_srl_151_n215, u1_srl_151_n214, u1_srl_151_n213,
         u1_srl_151_n212, u1_srl_151_n211, u1_srl_151_n210, u1_srl_151_n209,
         u1_srl_151_n208, u1_srl_151_n207, u1_srl_151_n206, u1_srl_151_n205,
         u1_srl_151_n204, u1_srl_151_n203, u1_srl_151_n202, u1_srl_151_n201,
         u1_srl_151_n200, u1_srl_151_n199, u1_srl_151_n198, u1_srl_151_n197,
         u1_srl_151_n196, u1_srl_151_n195, u1_srl_151_n194, u1_srl_151_n193,
         u1_srl_151_n192, u1_srl_151_n191, u1_srl_151_n190, u1_srl_151_n189,
         u1_srl_151_n188, u1_srl_151_n187, u1_srl_151_n186, u1_srl_151_n185,
         u1_srl_151_n184, u1_srl_151_n183, u1_srl_151_n182, u1_srl_151_n181,
         u1_srl_151_n180, u1_srl_151_n179, u1_srl_151_n178, u1_srl_151_n177,
         u1_srl_151_n176, u1_srl_151_n175, u1_srl_151_n174, u1_srl_151_n173,
         u1_srl_151_n172, u1_srl_151_n171, u1_srl_151_n170, u1_srl_151_n169,
         u1_srl_151_n168, u1_srl_151_n167, u1_srl_151_n166, u1_srl_151_n165,
         u1_srl_151_n164, u1_srl_151_n163, u1_srl_151_n162, u1_srl_151_n161,
         u1_srl_151_n160, u1_srl_151_n159, u1_srl_151_n158, u1_srl_151_n157,
         u1_srl_151_n156, u1_srl_151_n155, u1_srl_151_n154, u1_srl_151_n153,
         u1_srl_151_n152, u1_srl_151_n151, u1_srl_151_n150, u1_srl_151_n149,
         u1_srl_151_n148, u1_srl_151_n147, u1_srl_151_n146, u1_srl_151_n145,
         u1_srl_151_n144, u1_srl_151_n143, u1_srl_151_n142, u1_srl_151_n141,
         u1_srl_151_n140, u1_srl_151_n139, u1_srl_151_n138, u1_srl_151_n137,
         u1_srl_151_n136, u1_srl_151_n135, u1_srl_151_n134, u1_srl_151_n133,
         u1_srl_151_n132, u1_srl_151_n131, u1_srl_151_n130, u1_srl_151_n129,
         u1_srl_151_n128, u1_srl_151_n127, u1_srl_151_n126, u1_srl_151_n125,
         u1_srl_151_n124, u1_srl_151_n123, u1_srl_151_n122, u1_srl_151_n121,
         u1_srl_151_n120, u1_srl_151_n119, u1_srl_151_n118, u1_srl_151_n117,
         u1_srl_151_n116, u1_srl_151_n115, u1_srl_151_n114, u1_srl_151_n113,
         u1_srl_151_n112, u1_srl_151_n111, u1_srl_151_n110, u1_srl_151_n109,
         u1_srl_151_n108, u1_srl_151_n107, u1_srl_151_n106, u1_srl_151_n105,
         u1_srl_151_n104, u1_srl_151_n103, u1_srl_151_n102, u1_srl_151_n101,
         u1_srl_151_n100, u1_srl_151_n99, u1_srl_151_n98, u1_srl_151_n97,
         u1_srl_151_n96, u1_srl_151_n95, u1_srl_151_n94, u1_srl_151_n93,
         u1_srl_151_n92, u1_srl_151_n91, u1_srl_151_n90, u1_srl_151_n89,
         u1_srl_151_n88, u1_srl_151_n87, u1_srl_151_n86, u1_srl_151_n85,
         u1_srl_151_n84, u1_srl_151_n83, u1_srl_151_n82, u1_srl_151_n81,
         u1_srl_151_n80, u1_srl_151_n79, u1_srl_151_n78, u1_srl_151_n77,
         u1_srl_151_n76, u1_srl_151_n75, u1_srl_151_n74, u1_srl_151_n73,
         u1_srl_151_n72, u1_srl_151_n71, u1_srl_151_n70, u1_srl_151_n69,
         u1_srl_151_n68, u1_srl_151_n67, u1_srl_151_n66, u1_srl_151_n65,
         u1_srl_151_n64, u1_srl_151_n63, u1_srl_151_n62, u1_srl_151_n61,
         u1_srl_151_n60, u1_srl_151_n59, u1_srl_151_n58, u1_srl_151_n57,
         u1_srl_151_n56, u1_srl_151_n55, u1_srl_151_n54, u1_srl_151_n53,
         u1_srl_151_n52, u1_srl_151_n51, u1_srl_151_n50, u1_srl_151_n49,
         u1_srl_151_n48, u1_srl_151_n47, u1_srl_151_n46, u1_srl_151_n45,
         u1_srl_151_n44, u1_srl_151_n43, u1_srl_151_n42, u1_srl_151_n41,
         u1_srl_151_n40, u1_srl_151_n39, u1_srl_151_n38, u1_srl_151_n37,
         u1_srl_151_n36, u1_srl_151_n35, u1_srl_151_n34, u1_srl_151_n33,
         u1_srl_151_n32, u1_srl_151_n31, u1_srl_151_n30, u1_srl_151_n29,
         u1_srl_151_n28, u1_srl_151_n27, u1_srl_151_n26, u1_srl_151_n25,
         u1_srl_151_n24, u1_srl_151_n23, u1_srl_151_n22, u1_srl_151_n21,
         u1_srl_151_n20, u1_srl_151_n19, u1_srl_151_n18, u1_srl_151_n17,
         u1_srl_151_n16, u1_srl_151_n15, u1_srl_151_n14, u1_srl_151_n13,
         u1_srl_151_n12, u1_srl_151_n11, u1_srl_151_n10, u1_srl_151_n9,
         u1_srl_151_n8, u1_srl_151_n7, u1_srl_151_n6, u1_srl_151_n5,
         u1_srl_151_n4, u1_srl_151_n3, u1_srl_151_n2, u1_srl_151_n1,
         sub_1_root_u1_sub_133_aco_n12, sub_1_root_u1_sub_133_aco_n11,
         sub_1_root_u1_sub_133_aco_n10, sub_1_root_u1_sub_133_aco_n9,
         sub_1_root_u1_sub_133_aco_n8, sub_1_root_u1_sub_133_aco_n7,
         sub_1_root_u1_sub_133_aco_n6, sub_1_root_u1_sub_133_aco_n5,
         sub_1_root_u1_sub_133_aco_n4, sub_1_root_u1_sub_133_aco_n3,
         sub_1_root_u1_sub_133_aco_n2, sub_1_root_u1_sub_133_aco_n1,
         sub_436_3_n171, sub_436_3_n170, sub_436_3_n169, sub_436_3_n168,
         sub_436_3_n167, sub_436_3_n166, sub_436_3_n165, sub_436_3_n164,
         sub_436_3_n163, sub_436_3_n162, sub_436_3_n161, sub_436_3_n160,
         sub_436_3_n159, sub_436_3_n158, sub_436_3_n157, sub_436_3_n156,
         sub_436_3_n155, sub_436_3_n154, sub_436_3_n153, sub_436_3_n152,
         sub_436_3_n151, sub_436_3_n150, sub_436_3_n149, sub_436_3_n148,
         sub_436_3_n147, sub_436_3_n146, sub_436_3_n145, sub_436_3_n144,
         sub_436_3_n143, sub_436_3_n142, sub_436_3_n141, sub_436_3_n140,
         sub_436_3_n139, sub_436_3_n138, sub_436_3_n137, sub_436_3_n136,
         sub_436_3_n135, sub_436_3_n134, sub_436_3_n133, sub_436_3_n132,
         sub_436_3_n131, sub_436_3_n130, sub_436_3_n129, sub_436_3_n128,
         sub_436_3_n127, sub_436_3_n126, sub_436_3_n125, sub_436_3_n124,
         sub_436_3_n123, sub_436_3_n122, sub_436_3_n121, sub_436_3_n120,
         sub_436_3_n119, sub_436_3_n118, sub_436_3_n117, sub_436_3_n116,
         sub_436_3_n115, sub_436_3_n114, sub_436_3_n113, sub_436_3_n112,
         sub_436_3_n111, sub_436_3_n110, sub_436_3_n109, sub_436_3_n108,
         sub_436_3_n107, sub_436_3_n106, sub_436_3_n105, sub_436_3_n104,
         sub_436_3_n103, sub_436_3_n102, sub_436_3_n101, sub_436_3_n100,
         sub_436_3_n99, sub_436_3_n98, sub_436_3_n97, sub_436_3_n96,
         sub_436_3_n95, sub_436_3_n94, sub_436_3_n93, sub_436_3_n92,
         sub_436_3_n91, sub_436_3_n90, sub_436_3_n89, sub_436_3_n88,
         sub_436_3_n87, sub_436_3_n86, sub_436_3_n85, sub_436_3_n84,
         sub_436_3_n83, sub_436_3_n82, sub_436_3_n81, sub_436_3_n80,
         sub_436_3_n79, sub_436_3_n78, sub_436_3_n77, sub_436_3_n76,
         sub_436_3_n75, sub_436_3_n74, sub_436_3_n73, sub_436_3_n72,
         sub_436_3_n71, sub_436_3_n70, sub_436_3_n69, sub_436_3_n68,
         sub_436_3_n67, sub_436_3_n66, sub_436_3_n65, sub_436_3_n64,
         sub_436_3_n63, sub_436_3_n62, sub_436_3_n61, sub_436_3_n60,
         sub_436_3_n59, sub_436_3_n58, sub_436_3_n57, sub_436_3_n56,
         sub_436_3_n55, sub_436_3_n54, sub_436_3_n53, sub_436_3_n52,
         sub_436_3_n51, sub_436_3_n50, sub_436_3_n49, sub_436_3_n48,
         sub_436_3_n47, sub_436_3_n46, sub_436_3_n45, sub_436_3_n44,
         sub_436_3_n43, sub_436_3_n42, sub_436_3_n41, sub_436_3_n40,
         sub_436_3_n39, sub_436_3_n38, sub_436_3_n37, sub_436_3_n36,
         sub_436_3_n35, sub_436_3_n34, sub_436_3_n33, sub_436_3_n32,
         sub_436_3_n31, sub_436_3_n30, sub_436_3_n29, sub_436_3_n28,
         sub_436_3_n27, sub_436_3_n26, sub_436_3_carry_50_,
         sub_436_3_carry_51_, sub_436_3_carry_52_, sub_436_3_carry_53_,
         sub_436_3_carry_54_, sub_436_3_carry_55_, sub_436_3_carry_56_,
         sub_436_3_carry_57_, sub_436_3_carry_58_, sub_436_3_carry_59_,
         sub_436_3_carry_60_, sub_436_3_carry_61_, sub_436_3_carry_62_,
         sub_436_3_carry_63_, sub_436_3_carry_64_, sub_436_3_carry_65_,
         sub_436_3_carry_66_, sub_436_3_carry_67_, sub_436_3_carry_68_,
         sub_436_3_carry_69_, sub_436_3_carry_70_, sub_436_3_carry_71_,
         sub_436_3_carry_72_, sub_436_3_carry_73_, sub_436_3_carry_74_,
         sub_436_3_carry_75_, sub_436_3_carry_76_, sub_436_3_carry_77_,
         sub_436_3_carry_78_, sub_436_3_carry_79_, sub_436_3_carry_80_,
         sub_436_3_carry_81_, sub_436_3_carry_82_, sub_436_3_carry_83_,
         sub_436_3_carry_84_, sub_436_3_carry_85_, sub_436_3_carry_86_,
         sub_436_3_carry_87_, sub_436_3_carry_88_, sub_436_3_carry_89_,
         sub_436_3_carry_90_, sub_436_3_carry_91_, sub_436_3_carry_92_,
         sub_436_3_carry_93_, sub_436_3_carry_94_, sub_436_3_carry_95_,
         sub_436_3_carry_96_, sub_436_3_carry_97_, sub_436_3_carry_98_,
         sub_436_3_carry_99_, sub_436_3_carry_100_, sub_436_3_carry_101_,
         sub_436_3_carry_102_, sub_436_3_carry_103_, sub_436_3_carry_104_,
         sub_436_3_carry_105_, sub_436_b0_n157, sub_436_b0_n156,
         sub_436_b0_n155, sub_436_b0_n154, sub_436_b0_n153, sub_436_b0_n152,
         sub_436_b0_n151, sub_436_b0_n150, sub_436_b0_n149, sub_436_b0_n148,
         sub_436_b0_n147, sub_436_b0_n146, sub_436_b0_n145, sub_436_b0_n144,
         sub_436_b0_n143, sub_436_b0_n142, sub_436_b0_n141, sub_436_b0_n140,
         sub_436_b0_n139, sub_436_b0_n138, sub_436_b0_n137, sub_436_b0_n136,
         sub_436_b0_n135, sub_436_b0_n134, sub_436_b0_n133, sub_436_b0_n132,
         sub_436_b0_n131, sub_436_b0_n130, sub_436_b0_n129, sub_436_b0_n128,
         sub_436_b0_n127, sub_436_b0_n126, sub_436_b0_n125, sub_436_b0_n124,
         sub_436_b0_n123, sub_436_b0_n122, sub_436_b0_n121, sub_436_b0_n120,
         sub_436_b0_n119, sub_436_b0_n118, sub_436_b0_n117, sub_436_b0_n116,
         sub_436_b0_n115, sub_436_b0_n114, sub_436_b0_n113, sub_436_b0_n112,
         sub_436_b0_n111, sub_436_b0_n110, sub_436_b0_n109, sub_436_b0_n108,
         sub_436_b0_n107, sub_436_b0_n106, sub_436_b0_n105, sub_436_b0_n104,
         sub_436_b0_n103, sub_436_b0_n102, sub_436_b0_n101, sub_436_b0_n100,
         sub_436_b0_n99, sub_436_b0_n98, sub_436_b0_n97, sub_436_b0_n96,
         sub_436_b0_n95, sub_436_b0_n94, sub_436_b0_n93, sub_436_b0_n92,
         sub_436_b0_n91, sub_436_b0_n90, sub_436_b0_n89, sub_436_b0_n88,
         sub_436_b0_n87, sub_436_b0_n86, sub_436_b0_n85, sub_436_b0_n84,
         sub_436_b0_n83, sub_436_b0_n82, sub_436_b0_n81, sub_436_b0_n80,
         sub_436_b0_n79, sub_436_b0_n78, sub_436_b0_n77, sub_436_b0_n76,
         sub_436_b0_n75, sub_436_b0_n74, sub_436_b0_n73, sub_436_b0_n72,
         sub_436_b0_n71, sub_436_b0_n70, sub_436_b0_n69, sub_436_b0_n68,
         sub_436_b0_n67, sub_436_b0_n66, sub_436_b0_n65, sub_436_b0_n64,
         sub_436_b0_n63, sub_436_b0_n62, sub_436_b0_n61, sub_436_b0_n60,
         sub_436_b0_n59, sub_436_b0_n58, sub_436_b0_n57, sub_436_b0_n56,
         sub_436_b0_n55, sub_436_b0_n54, sub_436_b0_n53, sub_436_b0_n52,
         sub_436_b0_n51, sub_436_b0_n50, sub_436_b0_n49, sub_436_b0_n48,
         sub_436_b0_n47, sub_436_b0_n46, sub_436_b0_n45, sub_436_b0_n44,
         sub_436_b0_n43, sub_436_b0_n42, sub_436_b0_n41, sub_436_b0_n40,
         sub_436_b0_n39, sub_436_b0_n38, sub_436_b0_n37, sub_436_b0_n36,
         sub_436_b0_n35, sub_436_b0_n34, sub_436_b0_n33, sub_436_b0_n32,
         sub_436_b0_n31, sub_436_b0_carry_2_, sub_436_b0_carry_3_,
         sub_436_b0_carry_4_, sub_436_b0_carry_5_, sub_436_b0_carry_6_,
         sub_436_b0_carry_7_, sub_436_b0_carry_8_, sub_436_b0_carry_9_,
         sub_436_b0_carry_10_, sub_436_b0_carry_11_, sub_436_b0_carry_12_,
         sub_436_b0_carry_13_, sub_436_b0_carry_14_, sub_436_b0_carry_15_,
         sub_436_b0_carry_16_, sub_436_b0_carry_17_, sub_436_b0_carry_18_,
         sub_436_b0_carry_19_, sub_436_b0_carry_20_, sub_436_b0_carry_21_,
         sub_436_b0_carry_22_, sub_436_b0_carry_23_, sub_436_b0_carry_24_,
         sub_436_b0_carry_25_, sub_436_b0_carry_26_, sub_436_b0_carry_27_,
         sub_436_b0_carry_28_, sub_436_b0_carry_29_, sub_436_b0_carry_30_,
         sub_436_b0_carry_31_, sub_436_b0_carry_32_, sub_436_b0_carry_33_,
         sub_436_b0_carry_34_, sub_436_b0_carry_35_, sub_436_b0_carry_36_,
         sub_436_b0_carry_37_, sub_436_b0_carry_38_, sub_436_b0_carry_39_,
         sub_436_b0_carry_40_, sub_436_b0_carry_41_, sub_436_b0_carry_42_,
         sub_436_b0_carry_43_, sub_436_b0_carry_44_, sub_436_b0_carry_45_,
         sub_436_b0_carry_46_, sub_436_b0_carry_47_, sub_436_b0_carry_48_,
         sub_436_b0_carry_49_, sub_436_b0_carry_50_, sub_436_b0_carry_51_,
         sub_436_b0_carry_52_, sll_386_n41, sll_386_n40, sll_386_n39,
         sll_386_n38, sll_386_n37, sll_386_n36, sll_386_n35, sll_386_n34,
         sll_386_n33, sll_386_n32, sll_386_n31, sll_386_n30, sll_386_n29,
         sll_386_n28, sll_386_n27, sll_386_n26, sll_386_n25, sll_386_n24,
         sll_386_n23, sll_386_n22, sll_386_n21, sll_386_n20, sll_386_n19,
         sll_386_n18, sll_386_n17, sll_386_n16, sll_386_n15, sll_386_n14,
         sll_386_n13, sll_386_n12, sll_386_n11, sll_386_n10, sll_386_n9,
         sll_386_n8, sll_386_n7, sll_386_n6, sll_386_n5, sll_386_n4,
         sll_386_n3, sll_386_n2, sll_386_n1, sll_386_ML_int_4__8_,
         sll_386_ML_int_4__9_, sll_386_ML_int_4__10_, sll_386_ML_int_4__11_,
         sll_386_ML_int_4__12_, sll_386_ML_int_4__13_, sll_386_ML_int_4__14_,
         sll_386_ML_int_4__15_, sll_386_ML_int_4__16_, sll_386_ML_int_4__17_,
         sll_386_ML_int_4__18_, sll_386_ML_int_4__19_, sll_386_ML_int_4__20_,
         sll_386_ML_int_4__21_, sll_386_ML_int_4__22_, sll_386_ML_int_4__23_,
         sll_386_ML_int_4__24_, sll_386_ML_int_4__25_, sll_386_ML_int_4__26_,
         sll_386_ML_int_4__27_, sll_386_ML_int_4__28_, sll_386_ML_int_4__29_,
         sll_386_ML_int_4__30_, sll_386_ML_int_4__31_, sll_386_ML_int_4__32_,
         sll_386_ML_int_4__33_, sll_386_ML_int_4__34_, sll_386_ML_int_4__35_,
         sll_386_ML_int_4__36_, sll_386_ML_int_4__37_, sll_386_ML_int_4__38_,
         sll_386_ML_int_4__39_, sll_386_ML_int_4__40_, sll_386_ML_int_4__41_,
         sll_386_ML_int_4__42_, sll_386_ML_int_4__43_, sll_386_ML_int_4__44_,
         sll_386_ML_int_4__45_, sll_386_ML_int_4__46_, sll_386_ML_int_4__47_,
         sll_386_ML_int_4__48_, sll_386_ML_int_4__49_, sll_386_ML_int_4__50_,
         sll_386_ML_int_4__51_, sll_386_ML_int_4__52_, sll_386_ML_int_3__0_,
         sll_386_ML_int_3__1_, sll_386_ML_int_3__2_, sll_386_ML_int_3__3_,
         sll_386_ML_int_3__4_, sll_386_ML_int_3__5_, sll_386_ML_int_3__6_,
         sll_386_ML_int_3__7_, sll_386_ML_int_3__8_, sll_386_ML_int_3__9_,
         sll_386_ML_int_3__10_, sll_386_ML_int_3__11_, sll_386_ML_int_3__12_,
         sll_386_ML_int_3__13_, sll_386_ML_int_3__14_, sll_386_ML_int_3__15_,
         sll_386_ML_int_3__16_, sll_386_ML_int_3__17_, sll_386_ML_int_3__18_,
         sll_386_ML_int_3__19_, sll_386_ML_int_3__20_, sll_386_ML_int_3__21_,
         sll_386_ML_int_3__22_, sll_386_ML_int_3__23_, sll_386_ML_int_3__24_,
         sll_386_ML_int_3__25_, sll_386_ML_int_3__26_, sll_386_ML_int_3__27_,
         sll_386_ML_int_3__28_, sll_386_ML_int_3__29_, sll_386_ML_int_3__30_,
         sll_386_ML_int_3__31_, sll_386_ML_int_3__32_, sll_386_ML_int_3__33_,
         sll_386_ML_int_3__34_, sll_386_ML_int_3__35_, sll_386_ML_int_3__36_,
         sll_386_ML_int_3__37_, sll_386_ML_int_3__38_, sll_386_ML_int_3__39_,
         sll_386_ML_int_3__40_, sll_386_ML_int_3__41_, sll_386_ML_int_3__42_,
         sll_386_ML_int_3__43_, sll_386_ML_int_3__44_, sll_386_ML_int_3__45_,
         sll_386_ML_int_3__46_, sll_386_ML_int_3__47_, sll_386_ML_int_3__48_,
         sll_386_ML_int_3__49_, sll_386_ML_int_3__50_, sll_386_ML_int_3__51_,
         sll_386_ML_int_3__52_, sll_386_ML_int_2__0_, sll_386_ML_int_2__1_,
         sll_386_ML_int_2__2_, sll_386_ML_int_2__3_, sll_386_ML_int_2__4_,
         sll_386_ML_int_2__5_, sll_386_ML_int_2__6_, sll_386_ML_int_2__7_,
         sll_386_ML_int_2__8_, sll_386_ML_int_2__9_, sll_386_ML_int_2__10_,
         sll_386_ML_int_2__11_, sll_386_ML_int_2__12_, sll_386_ML_int_2__13_,
         sll_386_ML_int_2__14_, sll_386_ML_int_2__15_, sll_386_ML_int_2__16_,
         sll_386_ML_int_2__17_, sll_386_ML_int_2__18_, sll_386_ML_int_2__19_,
         sll_386_ML_int_2__20_, sll_386_ML_int_2__21_, sll_386_ML_int_2__22_,
         sll_386_ML_int_2__23_, sll_386_ML_int_2__24_, sll_386_ML_int_2__25_,
         sll_386_ML_int_2__26_, sll_386_ML_int_2__27_, sll_386_ML_int_2__28_,
         sll_386_ML_int_2__29_, sll_386_ML_int_2__30_, sll_386_ML_int_2__31_,
         sll_386_ML_int_2__32_, sll_386_ML_int_2__33_, sll_386_ML_int_2__34_,
         sll_386_ML_int_2__35_, sll_386_ML_int_2__36_, sll_386_ML_int_2__37_,
         sll_386_ML_int_2__38_, sll_386_ML_int_2__39_, sll_386_ML_int_2__40_,
         sll_386_ML_int_2__41_, sll_386_ML_int_2__42_, sll_386_ML_int_2__43_,
         sll_386_ML_int_2__44_, sll_386_ML_int_2__45_, sll_386_ML_int_2__46_,
         sll_386_ML_int_2__47_, sll_386_ML_int_2__48_, sll_386_ML_int_2__49_,
         sll_386_ML_int_2__50_, sll_386_ML_int_2__51_, sll_386_ML_int_2__52_,
         sll_386_ML_int_1__0_, sll_386_ML_int_1__1_, sll_386_ML_int_1__2_,
         sll_386_ML_int_1__3_, sll_386_ML_int_1__4_, sll_386_ML_int_1__5_,
         sll_386_ML_int_1__6_, sll_386_ML_int_1__7_, sll_386_ML_int_1__8_,
         sll_386_ML_int_1__9_, sll_386_ML_int_1__10_, sll_386_ML_int_1__11_,
         sll_386_ML_int_1__12_, sll_386_ML_int_1__13_, sll_386_ML_int_1__14_,
         sll_386_ML_int_1__15_, sll_386_ML_int_1__16_, sll_386_ML_int_1__17_,
         sll_386_ML_int_1__18_, sll_386_ML_int_1__19_, sll_386_ML_int_1__20_,
         sll_386_ML_int_1__21_, sll_386_ML_int_1__22_, sll_386_ML_int_1__23_,
         sll_386_ML_int_1__24_, sll_386_ML_int_1__25_, sll_386_ML_int_1__26_,
         sll_386_ML_int_1__27_, sll_386_ML_int_1__28_, sll_386_ML_int_1__29_,
         sll_386_ML_int_1__30_, sll_386_ML_int_1__31_, sll_386_ML_int_1__32_,
         sll_386_ML_int_1__33_, sll_386_ML_int_1__34_, sll_386_ML_int_1__35_,
         sll_386_ML_int_1__36_, sll_386_ML_int_1__37_, sll_386_ML_int_1__38_,
         sll_386_ML_int_1__39_, sll_386_ML_int_1__40_, sll_386_ML_int_1__41_,
         sll_386_ML_int_1__42_, sll_386_ML_int_1__43_, sll_386_ML_int_1__44_,
         sll_386_ML_int_1__45_, sll_386_ML_int_1__46_, sll_386_ML_int_1__47_,
         sll_386_ML_int_1__48_, sll_386_ML_int_1__49_, sll_386_ML_int_1__50_,
         sll_386_ML_int_1__51_, sll_386_ML_int_1__52_, r471_n178, r471_n177,
         r471_n176, r471_n175, r471_n174, r471_n173, r471_n172, r471_n171,
         r471_n170, r471_n169, r471_n168, r471_n167, r471_n166, r471_n165,
         r471_n164, r471_n163, r471_n162, r471_n161, r471_n160, r471_n159,
         r471_n158, r471_n157, r471_n156, r471_n155, r471_n154, r471_n153,
         r471_n152, r471_n151, r471_n150, r471_n149, r471_n148, r471_n147,
         r471_n146, r471_n145, r471_n144, r471_n143, r471_n142, r471_n141,
         r471_n140, r471_n139, r471_n138, r471_n137, r471_n136, r471_n135,
         r471_n134, r471_n133, r471_n132, r471_n131, r471_n130, r471_n129,
         r471_n128, r471_n127, r471_n126, r471_n125, r471_n124, r471_n123,
         r471_n122, r471_n121, r471_n120, r471_n119, r471_n118, r471_n117,
         r471_n116, r471_n115, r471_n114, r471_n113, r471_n112, r471_n111,
         r471_n110, r471_n109, r471_n108, r471_n107, r471_n106, r471_n105,
         r471_n104, r471_n103, r471_n102, r471_n101, r471_n100, r471_n99,
         r471_n98, r471_n97, r471_n96, r471_n95, r471_n94, r471_n93, r471_n92,
         r471_n91, r471_n90, r471_n89, r471_n88, r471_n87, r471_n86, r471_n85,
         r471_n84, r471_n83, r471_n82, r471_n81, r471_n80, r471_n79, r471_n78,
         r471_n77, r471_n76, r471_n75, r471_n74, r471_n73, r471_n72, r471_n71,
         r471_n70, r471_n69, r471_n68, r471_n67, r471_n66, r471_n65, r471_n64,
         r471_n63, r471_n62, r471_n61, r471_n60, r471_n59, r471_n58, r471_n57,
         r471_n56, r471_n55, r471_n54, r471_n53, r471_n52, r471_n51, r471_n50,
         r471_n49, r471_n48, r471_n47, r471_n46, r471_n45, r471_n44, r471_n43,
         r471_n42, r471_n41, r471_n40, r471_n39, r471_n38, r471_n37, r471_n36,
         r471_n35, r471_n34, r471_n33, r471_n32, r471_n31, r471_n30, r471_n29,
         r471_n28, r471_n27, r471_n26, r471_n25, r471_n24, r471_n23, r471_n22,
         r471_n21, r471_n20, r471_n19, r471_n18, r471_n17, r471_n16, r471_n15,
         r471_n14, r471_n13, r471_n12, r471_n11, r471_n10, r471_n9, r471_n8,
         r471_n7, r471_n6, r471_n5, r471_n4, r471_n3, r471_n2, r471_n1,
         add_0_root_sub_0_root_u4_add_497_n7,
         add_0_root_sub_0_root_u4_add_497_n6,
         add_0_root_sub_0_root_u4_add_497_n5,
         add_0_root_sub_0_root_u4_add_497_n1,
         add_0_root_sub_0_root_u4_add_497_carry_2_,
         add_0_root_sub_0_root_u4_add_497_carry_3_,
         add_0_root_sub_0_root_u4_add_497_carry_4_,
         add_0_root_sub_0_root_u4_add_497_carry_5_,
         add_0_root_sub_0_root_u4_add_497_carry_6_,
         add_0_root_sub_0_root_u4_add_497_carry_7_,
         add_0_root_sub_0_root_u4_add_497_carry_8_,
         add_0_root_sub_0_root_u4_add_497_carry_9_,
         add_0_root_sub_0_root_u4_add_497_carry_10_, u5_mult_82_n7022,
         u5_mult_82_n7021, u5_mult_82_n7020, u5_mult_82_n7019,
         u5_mult_82_n7018, u5_mult_82_n7017, u5_mult_82_n7016,
         u5_mult_82_n7015, u5_mult_82_n7014, u5_mult_82_n7013,
         u5_mult_82_n7012, u5_mult_82_n7011, u5_mult_82_n7010,
         u5_mult_82_n7009, u5_mult_82_n7008, u5_mult_82_n7007,
         u5_mult_82_n7006, u5_mult_82_n7005, u5_mult_82_n7004,
         u5_mult_82_n7003, u5_mult_82_n7002, u5_mult_82_n7001,
         u5_mult_82_n7000, u5_mult_82_n6999, u5_mult_82_n6998,
         u5_mult_82_n6997, u5_mult_82_n6996, u5_mult_82_n6995,
         u5_mult_82_n6994, u5_mult_82_n6993, u5_mult_82_n6992,
         u5_mult_82_n6991, u5_mult_82_n6990, u5_mult_82_n6989,
         u5_mult_82_n6988, u5_mult_82_n6987, u5_mult_82_n6986,
         u5_mult_82_n6985, u5_mult_82_n6984, u5_mult_82_n6983,
         u5_mult_82_n6982, u5_mult_82_n6981, u5_mult_82_n6980,
         u5_mult_82_n6979, u5_mult_82_n6978, u5_mult_82_n6977,
         u5_mult_82_n6976, u5_mult_82_n6975, u5_mult_82_n6974,
         u5_mult_82_n6973, u5_mult_82_n6972, u5_mult_82_n6971,
         u5_mult_82_n6970, u5_mult_82_n6969, u5_mult_82_n6968,
         u5_mult_82_n6967, u5_mult_82_n6966, u5_mult_82_n6965,
         u5_mult_82_n6964, u5_mult_82_n6963, u5_mult_82_n6962,
         u5_mult_82_n6961, u5_mult_82_n6960, u5_mult_82_n6959,
         u5_mult_82_n6958, u5_mult_82_n6957, u5_mult_82_n6956,
         u5_mult_82_n6955, u5_mult_82_n6954, u5_mult_82_n6953,
         u5_mult_82_n6952, u5_mult_82_n6951, u5_mult_82_n6950,
         u5_mult_82_n6949, u5_mult_82_n6948, u5_mult_82_n6947,
         u5_mult_82_n6946, u5_mult_82_n6945, u5_mult_82_n6944,
         u5_mult_82_n6943, u5_mult_82_n6942, u5_mult_82_n6941,
         u5_mult_82_n6940, u5_mult_82_n6939, u5_mult_82_n6938,
         u5_mult_82_n6937, u5_mult_82_n6936, u5_mult_82_n6935,
         u5_mult_82_n6934, u5_mult_82_n6933, u5_mult_82_n6932,
         u5_mult_82_n6931, u5_mult_82_n6930, u5_mult_82_n6929,
         u5_mult_82_n6928, u5_mult_82_n6927, u5_mult_82_n6926,
         u5_mult_82_n6925, u5_mult_82_n6924, u5_mult_82_n6923,
         u5_mult_82_n6922, u5_mult_82_n6921, u5_mult_82_n6920,
         u5_mult_82_n6919, u5_mult_82_n6918, u5_mult_82_n6917,
         u5_mult_82_n6916, u5_mult_82_n6915, u5_mult_82_n6914,
         u5_mult_82_n6913, u5_mult_82_n6912, u5_mult_82_n6911,
         u5_mult_82_n6910, u5_mult_82_n6909, u5_mult_82_n6908,
         u5_mult_82_n6907, u5_mult_82_n6906, u5_mult_82_n6905,
         u5_mult_82_n6904, u5_mult_82_n6903, u5_mult_82_n6902,
         u5_mult_82_n6901, u5_mult_82_n6900, u5_mult_82_n6899,
         u5_mult_82_n6898, u5_mult_82_n6897, u5_mult_82_n6896,
         u5_mult_82_n6895, u5_mult_82_n6894, u5_mult_82_n6893,
         u5_mult_82_n6892, u5_mult_82_n6891, u5_mult_82_n6890,
         u5_mult_82_n6889, u5_mult_82_n6888, u5_mult_82_n6887,
         u5_mult_82_n6886, u5_mult_82_n6885, u5_mult_82_n6884,
         u5_mult_82_n6883, u5_mult_82_n6882, u5_mult_82_n6881,
         u5_mult_82_n6880, u5_mult_82_n6879, u5_mult_82_n6878,
         u5_mult_82_n6877, u5_mult_82_n6876, u5_mult_82_n6875,
         u5_mult_82_n6874, u5_mult_82_n6873, u5_mult_82_n6872,
         u5_mult_82_n6871, u5_mult_82_n6870, u5_mult_82_n6869,
         u5_mult_82_n6868, u5_mult_82_n6867, u5_mult_82_n6866,
         u5_mult_82_n6865, u5_mult_82_n6864, u5_mult_82_n6863,
         u5_mult_82_n6862, u5_mult_82_n6861, u5_mult_82_n6860,
         u5_mult_82_n6859, u5_mult_82_n6858, u5_mult_82_n6857,
         u5_mult_82_n6856, u5_mult_82_n6855, u5_mult_82_n6854,
         u5_mult_82_n6853, u5_mult_82_n6852, u5_mult_82_n6851,
         u5_mult_82_n6850, u5_mult_82_n6849, u5_mult_82_n6848,
         u5_mult_82_n6847, u5_mult_82_n6846, u5_mult_82_n6845,
         u5_mult_82_n6844, u5_mult_82_n6843, u5_mult_82_n6842,
         u5_mult_82_n6841, u5_mult_82_n6840, u5_mult_82_n6839,
         u5_mult_82_n6838, u5_mult_82_n6837, u5_mult_82_n6836,
         u5_mult_82_n6835, u5_mult_82_n6834, u5_mult_82_n6833,
         u5_mult_82_n6832, u5_mult_82_n6831, u5_mult_82_n6830,
         u5_mult_82_n6829, u5_mult_82_n6828, u5_mult_82_n6827,
         u5_mult_82_n6826, u5_mult_82_n6825, u5_mult_82_n6824,
         u5_mult_82_n6823, u5_mult_82_n6822, u5_mult_82_n6821,
         u5_mult_82_n6820, u5_mult_82_n6819, u5_mult_82_n6818,
         u5_mult_82_n6817, u5_mult_82_n6816, u5_mult_82_n6815,
         u5_mult_82_n6814, u5_mult_82_n6813, u5_mult_82_n6812,
         u5_mult_82_n6811, u5_mult_82_n6810, u5_mult_82_n6809,
         u5_mult_82_n6808, u5_mult_82_n6807, u5_mult_82_n6806,
         u5_mult_82_n6805, u5_mult_82_n6804, u5_mult_82_n6803,
         u5_mult_82_n6802, u5_mult_82_n6801, u5_mult_82_n6800,
         u5_mult_82_n6799, u5_mult_82_n6798, u5_mult_82_n6797,
         u5_mult_82_n6796, u5_mult_82_n6795, u5_mult_82_n6794,
         u5_mult_82_n6793, u5_mult_82_n6792, u5_mult_82_n6791,
         u5_mult_82_n6790, u5_mult_82_n6789, u5_mult_82_n6788,
         u5_mult_82_n6787, u5_mult_82_n6786, u5_mult_82_n6785,
         u5_mult_82_n6784, u5_mult_82_n6783, u5_mult_82_n6782,
         u5_mult_82_n6781, u5_mult_82_n6780, u5_mult_82_n6779,
         u5_mult_82_n6778, u5_mult_82_n6777, u5_mult_82_n6776,
         u5_mult_82_n6775, u5_mult_82_n6774, u5_mult_82_n6773,
         u5_mult_82_n6772, u5_mult_82_n6771, u5_mult_82_n6770,
         u5_mult_82_n6769, u5_mult_82_n6768, u5_mult_82_n6767,
         u5_mult_82_n6766, u5_mult_82_n6765, u5_mult_82_n6764,
         u5_mult_82_n6763, u5_mult_82_n6762, u5_mult_82_n6761,
         u5_mult_82_n6760, u5_mult_82_n6759, u5_mult_82_n6758,
         u5_mult_82_n6757, u5_mult_82_n6756, u5_mult_82_n6755,
         u5_mult_82_n6754, u5_mult_82_n6753, u5_mult_82_n6752,
         u5_mult_82_n6751, u5_mult_82_n6750, u5_mult_82_n6749,
         u5_mult_82_n6748, u5_mult_82_n6747, u5_mult_82_n6746,
         u5_mult_82_n6745, u5_mult_82_n6744, u5_mult_82_n6743,
         u5_mult_82_n6742, u5_mult_82_n6741, u5_mult_82_n6740,
         u5_mult_82_n6739, u5_mult_82_n6738, u5_mult_82_n6737,
         u5_mult_82_n6736, u5_mult_82_n6735, u5_mult_82_n6734,
         u5_mult_82_n6733, u5_mult_82_n6732, u5_mult_82_n6731,
         u5_mult_82_n6730, u5_mult_82_n6729, u5_mult_82_n6728,
         u5_mult_82_n6727, u5_mult_82_n6726, u5_mult_82_n6725,
         u5_mult_82_n6724, u5_mult_82_n6723, u5_mult_82_n6722,
         u5_mult_82_n6721, u5_mult_82_n6720, u5_mult_82_n6719,
         u5_mult_82_n6718, u5_mult_82_n6717, u5_mult_82_n6716,
         u5_mult_82_n6715, u5_mult_82_n6714, u5_mult_82_n6713,
         u5_mult_82_n6712, u5_mult_82_n6711, u5_mult_82_n6710,
         u5_mult_82_n6709, u5_mult_82_n6708, u5_mult_82_n6707,
         u5_mult_82_n6706, u5_mult_82_n6705, u5_mult_82_n6704,
         u5_mult_82_n6703, u5_mult_82_n6702, u5_mult_82_n6701,
         u5_mult_82_n6700, u5_mult_82_n6699, u5_mult_82_n6698,
         u5_mult_82_n6697, u5_mult_82_n6696, u5_mult_82_n6695,
         u5_mult_82_n6694, u5_mult_82_n6693, u5_mult_82_n6692,
         u5_mult_82_n6691, u5_mult_82_n6690, u5_mult_82_n6689,
         u5_mult_82_n6688, u5_mult_82_n6687, u5_mult_82_n6686,
         u5_mult_82_n6685, u5_mult_82_n6684, u5_mult_82_n6683,
         u5_mult_82_n6682, u5_mult_82_n6681, u5_mult_82_n6680,
         u5_mult_82_n6679, u5_mult_82_n6678, u5_mult_82_n6677,
         u5_mult_82_n6676, u5_mult_82_n6675, u5_mult_82_n6674,
         u5_mult_82_n6673, u5_mult_82_n6672, u5_mult_82_n6671,
         u5_mult_82_n6670, u5_mult_82_n6669, u5_mult_82_n6668,
         u5_mult_82_n6667, u5_mult_82_n6666, u5_mult_82_n6665,
         u5_mult_82_n6664, u5_mult_82_n6663, u5_mult_82_n6662,
         u5_mult_82_n6661, u5_mult_82_n6660, u5_mult_82_n6659,
         u5_mult_82_n6658, u5_mult_82_n6657, u5_mult_82_n6656,
         u5_mult_82_n6655, u5_mult_82_n6654, u5_mult_82_n6653,
         u5_mult_82_n6652, u5_mult_82_n6651, u5_mult_82_n6650,
         u5_mult_82_n6649, u5_mult_82_n6648, u5_mult_82_n6647,
         u5_mult_82_n6646, u5_mult_82_n6645, u5_mult_82_n6644,
         u5_mult_82_n6643, u5_mult_82_n6642, u5_mult_82_n6641,
         u5_mult_82_n6640, u5_mult_82_n6639, u5_mult_82_n6638,
         u5_mult_82_n6637, u5_mult_82_n6636, u5_mult_82_n6635,
         u5_mult_82_n6634, u5_mult_82_n6633, u5_mult_82_n6632,
         u5_mult_82_n6631, u5_mult_82_n6630, u5_mult_82_n6629,
         u5_mult_82_n6628, u5_mult_82_n6627, u5_mult_82_n6626,
         u5_mult_82_n6625, u5_mult_82_n6624, u5_mult_82_n6623,
         u5_mult_82_n6622, u5_mult_82_n6621, u5_mult_82_n6620,
         u5_mult_82_n6619, u5_mult_82_n6618, u5_mult_82_n6617,
         u5_mult_82_n6616, u5_mult_82_n6615, u5_mult_82_n6614,
         u5_mult_82_n6613, u5_mult_82_n6612, u5_mult_82_n6611,
         u5_mult_82_n6610, u5_mult_82_n6609, u5_mult_82_n6608,
         u5_mult_82_n6607, u5_mult_82_n6606, u5_mult_82_n6605,
         u5_mult_82_n6604, u5_mult_82_n6603, u5_mult_82_n6602,
         u5_mult_82_n6601, u5_mult_82_n6600, u5_mult_82_n6599,
         u5_mult_82_n6598, u5_mult_82_n6597, u5_mult_82_n6596,
         u5_mult_82_n6595, u5_mult_82_n6594, u5_mult_82_n6593,
         u5_mult_82_n6592, u5_mult_82_n6591, u5_mult_82_n6590,
         u5_mult_82_n6589, u5_mult_82_n6588, u5_mult_82_n6587,
         u5_mult_82_n6586, u5_mult_82_n6585, u5_mult_82_n6584,
         u5_mult_82_n6583, u5_mult_82_n6582, u5_mult_82_n6581,
         u5_mult_82_n6580, u5_mult_82_n6579, u5_mult_82_n6578,
         u5_mult_82_n6577, u5_mult_82_n6576, u5_mult_82_n6575,
         u5_mult_82_n6574, u5_mult_82_n6573, u5_mult_82_n6572,
         u5_mult_82_n6571, u5_mult_82_n6570, u5_mult_82_n6569,
         u5_mult_82_n6568, u5_mult_82_n6567, u5_mult_82_n6566,
         u5_mult_82_n6565, u5_mult_82_n6564, u5_mult_82_n6563,
         u5_mult_82_n6562, u5_mult_82_n6561, u5_mult_82_n6560,
         u5_mult_82_n6559, u5_mult_82_n6558, u5_mult_82_n6557,
         u5_mult_82_n6556, u5_mult_82_n6555, u5_mult_82_n6554,
         u5_mult_82_n6553, u5_mult_82_n6552, u5_mult_82_n6551,
         u5_mult_82_n6550, u5_mult_82_n6549, u5_mult_82_n6548,
         u5_mult_82_n6547, u5_mult_82_n6546, u5_mult_82_n6545,
         u5_mult_82_n6544, u5_mult_82_n6543, u5_mult_82_n6542,
         u5_mult_82_n6541, u5_mult_82_n6540, u5_mult_82_n6539,
         u5_mult_82_n6538, u5_mult_82_n6537, u5_mult_82_n6536,
         u5_mult_82_n6535, u5_mult_82_n6534, u5_mult_82_n6533,
         u5_mult_82_n6532, u5_mult_82_n6531, u5_mult_82_n6530,
         u5_mult_82_n6529, u5_mult_82_n6528, u5_mult_82_n6527,
         u5_mult_82_n6526, u5_mult_82_n6525, u5_mult_82_n6524,
         u5_mult_82_n6523, u5_mult_82_n6522, u5_mult_82_n6521,
         u5_mult_82_n6520, u5_mult_82_n6519, u5_mult_82_n6518,
         u5_mult_82_n6517, u5_mult_82_n6516, u5_mult_82_n6515,
         u5_mult_82_n6514, u5_mult_82_n6513, u5_mult_82_n6512,
         u5_mult_82_n6511, u5_mult_82_n6510, u5_mult_82_n6509,
         u5_mult_82_n6508, u5_mult_82_n6507, u5_mult_82_n6506,
         u5_mult_82_n6505, u5_mult_82_n6504, u5_mult_82_n6503,
         u5_mult_82_n6502, u5_mult_82_n6501, u5_mult_82_n6500,
         u5_mult_82_n6499, u5_mult_82_n6498, u5_mult_82_n6497,
         u5_mult_82_n6496, u5_mult_82_n6495, u5_mult_82_n6494,
         u5_mult_82_n6493, u5_mult_82_n6492, u5_mult_82_n6491,
         u5_mult_82_n6490, u5_mult_82_n6489, u5_mult_82_n6488,
         u5_mult_82_n6487, u5_mult_82_n6486, u5_mult_82_n6485,
         u5_mult_82_n6484, u5_mult_82_n6483, u5_mult_82_n6482,
         u5_mult_82_n6481, u5_mult_82_n6480, u5_mult_82_n6479,
         u5_mult_82_n6478, u5_mult_82_n6477, u5_mult_82_n6476,
         u5_mult_82_n6475, u5_mult_82_n6474, u5_mult_82_n6473,
         u5_mult_82_n6472, u5_mult_82_n6471, u5_mult_82_n6470,
         u5_mult_82_n6469, u5_mult_82_n6468, u5_mult_82_n6467,
         u5_mult_82_n6466, u5_mult_82_n6465, u5_mult_82_n6464,
         u5_mult_82_n6463, u5_mult_82_n6462, u5_mult_82_n6461,
         u5_mult_82_n6460, u5_mult_82_n6459, u5_mult_82_n6458,
         u5_mult_82_n6457, u5_mult_82_n6456, u5_mult_82_n6455,
         u5_mult_82_n6454, u5_mult_82_n6453, u5_mult_82_n6452,
         u5_mult_82_n6451, u5_mult_82_n6450, u5_mult_82_n6449,
         u5_mult_82_n6448, u5_mult_82_n6447, u5_mult_82_n6446,
         u5_mult_82_n6445, u5_mult_82_n6444, u5_mult_82_n6443,
         u5_mult_82_n6442, u5_mult_82_n6441, u5_mult_82_n6440,
         u5_mult_82_n6439, u5_mult_82_n6438, u5_mult_82_n6437,
         u5_mult_82_n6436, u5_mult_82_n6435, u5_mult_82_n6434,
         u5_mult_82_n6433, u5_mult_82_n6432, u5_mult_82_n6431,
         u5_mult_82_n6430, u5_mult_82_n6429, u5_mult_82_n6428,
         u5_mult_82_n6427, u5_mult_82_n6426, u5_mult_82_n6425,
         u5_mult_82_n6424, u5_mult_82_n6423, u5_mult_82_n6422,
         u5_mult_82_n6421, u5_mult_82_n6420, u5_mult_82_n6419,
         u5_mult_82_n6418, u5_mult_82_n6417, u5_mult_82_n6416,
         u5_mult_82_n6415, u5_mult_82_n6414, u5_mult_82_n6413,
         u5_mult_82_n6412, u5_mult_82_n6411, u5_mult_82_n6410,
         u5_mult_82_n6409, u5_mult_82_n6408, u5_mult_82_n6407,
         u5_mult_82_n6406, u5_mult_82_n6405, u5_mult_82_n6404,
         u5_mult_82_n6403, u5_mult_82_n6402, u5_mult_82_n6401,
         u5_mult_82_n6400, u5_mult_82_n6399, u5_mult_82_n6398,
         u5_mult_82_n6397, u5_mult_82_n6396, u5_mult_82_n6395,
         u5_mult_82_n6394, u5_mult_82_n6393, u5_mult_82_n6392,
         u5_mult_82_n6391, u5_mult_82_n6390, u5_mult_82_n6389,
         u5_mult_82_n6388, u5_mult_82_n6387, u5_mult_82_n6386,
         u5_mult_82_n6385, u5_mult_82_n6384, u5_mult_82_n6383,
         u5_mult_82_n6382, u5_mult_82_n6381, u5_mult_82_n6380,
         u5_mult_82_n6379, u5_mult_82_n6378, u5_mult_82_n6377,
         u5_mult_82_n6376, u5_mult_82_n6375, u5_mult_82_n6374,
         u5_mult_82_n6373, u5_mult_82_n6372, u5_mult_82_n6371,
         u5_mult_82_n6370, u5_mult_82_n6369, u5_mult_82_n6368,
         u5_mult_82_n6367, u5_mult_82_n6366, u5_mult_82_n6365,
         u5_mult_82_n6364, u5_mult_82_n6363, u5_mult_82_n6362,
         u5_mult_82_n6361, u5_mult_82_n6360, u5_mult_82_n6359,
         u5_mult_82_n6358, u5_mult_82_n6357, u5_mult_82_n6356,
         u5_mult_82_n6355, u5_mult_82_n6354, u5_mult_82_n6353,
         u5_mult_82_n6352, u5_mult_82_n6351, u5_mult_82_n6350,
         u5_mult_82_n6349, u5_mult_82_n6348, u5_mult_82_n6347,
         u5_mult_82_n6346, u5_mult_82_n6345, u5_mult_82_n6344,
         u5_mult_82_n6343, u5_mult_82_n6342, u5_mult_82_n6341,
         u5_mult_82_n6340, u5_mult_82_n6339, u5_mult_82_n6338,
         u5_mult_82_n6337, u5_mult_82_n6336, u5_mult_82_n6335,
         u5_mult_82_n6334, u5_mult_82_n6333, u5_mult_82_n6332,
         u5_mult_82_n6331, u5_mult_82_n6330, u5_mult_82_n6329,
         u5_mult_82_n6328, u5_mult_82_n6327, u5_mult_82_n6326,
         u5_mult_82_n6325, u5_mult_82_n6324, u5_mult_82_n6323,
         u5_mult_82_n6322, u5_mult_82_n6321, u5_mult_82_n6320,
         u5_mult_82_n6319, u5_mult_82_n6318, u5_mult_82_n6317,
         u5_mult_82_n6316, u5_mult_82_n6315, u5_mult_82_n6314,
         u5_mult_82_n6313, u5_mult_82_n6312, u5_mult_82_n6311,
         u5_mult_82_n6310, u5_mult_82_n6309, u5_mult_82_n6308,
         u5_mult_82_n6307, u5_mult_82_n6306, u5_mult_82_n6305,
         u5_mult_82_n6304, u5_mult_82_n6303, u5_mult_82_n6302,
         u5_mult_82_n6301, u5_mult_82_n6300, u5_mult_82_n6299,
         u5_mult_82_n6298, u5_mult_82_n6297, u5_mult_82_n6296,
         u5_mult_82_n6295, u5_mult_82_n6294, u5_mult_82_n6293,
         u5_mult_82_n6292, u5_mult_82_n6291, u5_mult_82_n6290,
         u5_mult_82_n6289, u5_mult_82_n6288, u5_mult_82_n6287,
         u5_mult_82_n6286, u5_mult_82_n6285, u5_mult_82_n6284,
         u5_mult_82_n6283, u5_mult_82_n6282, u5_mult_82_n6281,
         u5_mult_82_n6280, u5_mult_82_n6279, u5_mult_82_n6278,
         u5_mult_82_n6277, u5_mult_82_n6276, u5_mult_82_n6275,
         u5_mult_82_n6274, u5_mult_82_n6273, u5_mult_82_n6272,
         u5_mult_82_n6271, u5_mult_82_n6270, u5_mult_82_n6269,
         u5_mult_82_n6268, u5_mult_82_n6267, u5_mult_82_n6266,
         u5_mult_82_n6265, u5_mult_82_n6264, u5_mult_82_n6263,
         u5_mult_82_n6262, u5_mult_82_n6261, u5_mult_82_n6260,
         u5_mult_82_n6259, u5_mult_82_n6258, u5_mult_82_n6257,
         u5_mult_82_n6256, u5_mult_82_n6255, u5_mult_82_n6254,
         u5_mult_82_n6253, u5_mult_82_n6252, u5_mult_82_n6251,
         u5_mult_82_n6250, u5_mult_82_n6249, u5_mult_82_n6248,
         u5_mult_82_n6247, u5_mult_82_n6246, u5_mult_82_n6245,
         u5_mult_82_n6244, u5_mult_82_n6243, u5_mult_82_n6242,
         u5_mult_82_n6241, u5_mult_82_n6240, u5_mult_82_n6239,
         u5_mult_82_n6238, u5_mult_82_n6237, u5_mult_82_n6236,
         u5_mult_82_n6235, u5_mult_82_n6234, u5_mult_82_n6233,
         u5_mult_82_n6232, u5_mult_82_n6231, u5_mult_82_n6230,
         u5_mult_82_n6229, u5_mult_82_n6228, u5_mult_82_n6227,
         u5_mult_82_n6226, u5_mult_82_n6225, u5_mult_82_n6224,
         u5_mult_82_n6223, u5_mult_82_n6222, u5_mult_82_n6221,
         u5_mult_82_n6220, u5_mult_82_n6219, u5_mult_82_n6218,
         u5_mult_82_n6217, u5_mult_82_n6216, u5_mult_82_n6215,
         u5_mult_82_n6214, u5_mult_82_n6213, u5_mult_82_n6212,
         u5_mult_82_n6211, u5_mult_82_n6210, u5_mult_82_n6209,
         u5_mult_82_n6208, u5_mult_82_n6207, u5_mult_82_n6206,
         u5_mult_82_n6205, u5_mult_82_n6204, u5_mult_82_n6203,
         u5_mult_82_n6202, u5_mult_82_n6201, u5_mult_82_n6200,
         u5_mult_82_n6199, u5_mult_82_n6198, u5_mult_82_n6197,
         u5_mult_82_n6196, u5_mult_82_n6195, u5_mult_82_n6194,
         u5_mult_82_n6193, u5_mult_82_n6192, u5_mult_82_n6191,
         u5_mult_82_n6190, u5_mult_82_n6189, u5_mult_82_n6188,
         u5_mult_82_n6187, u5_mult_82_n6186, u5_mult_82_n6185,
         u5_mult_82_n6184, u5_mult_82_n6183, u5_mult_82_n6182,
         u5_mult_82_n6181, u5_mult_82_n6180, u5_mult_82_n6179,
         u5_mult_82_n6178, u5_mult_82_n6177, u5_mult_82_n6176,
         u5_mult_82_n6175, u5_mult_82_n6174, u5_mult_82_n6173,
         u5_mult_82_n6172, u5_mult_82_n6171, u5_mult_82_n6170,
         u5_mult_82_n6169, u5_mult_82_n6168, u5_mult_82_n6167,
         u5_mult_82_n6166, u5_mult_82_n6165, u5_mult_82_n6164,
         u5_mult_82_n6163, u5_mult_82_n6162, u5_mult_82_n6161,
         u5_mult_82_n6160, u5_mult_82_n6159, u5_mult_82_n6158,
         u5_mult_82_n6157, u5_mult_82_n6156, u5_mult_82_n6155,
         u5_mult_82_n6154, u5_mult_82_n6153, u5_mult_82_n6152,
         u5_mult_82_n6151, u5_mult_82_n6150, u5_mult_82_n6149,
         u5_mult_82_n6148, u5_mult_82_n6147, u5_mult_82_n6146,
         u5_mult_82_n6145, u5_mult_82_n6144, u5_mult_82_n6143,
         u5_mult_82_n6142, u5_mult_82_n6141, u5_mult_82_n6140,
         u5_mult_82_n6139, u5_mult_82_n6138, u5_mult_82_n6137,
         u5_mult_82_n6136, u5_mult_82_n6135, u5_mult_82_n6134,
         u5_mult_82_n6133, u5_mult_82_n6132, u5_mult_82_n6131,
         u5_mult_82_n6130, u5_mult_82_n6129, u5_mult_82_n6128,
         u5_mult_82_n6127, u5_mult_82_n6126, u5_mult_82_n6125,
         u5_mult_82_n6124, u5_mult_82_n6123, u5_mult_82_n6122,
         u5_mult_82_n6121, u5_mult_82_n6120, u5_mult_82_n6119,
         u5_mult_82_n6118, u5_mult_82_n6117, u5_mult_82_n6116,
         u5_mult_82_n6115, u5_mult_82_n6114, u5_mult_82_n6113,
         u5_mult_82_n6112, u5_mult_82_n6111, u5_mult_82_n6110,
         u5_mult_82_n6109, u5_mult_82_n6108, u5_mult_82_n6107,
         u5_mult_82_n6106, u5_mult_82_n6105, u5_mult_82_n6104,
         u5_mult_82_n6103, u5_mult_82_n6102, u5_mult_82_n6101,
         u5_mult_82_n6100, u5_mult_82_n6099, u5_mult_82_n6098,
         u5_mult_82_n6097, u5_mult_82_n6096, u5_mult_82_n6095,
         u5_mult_82_n6094, u5_mult_82_n6093, u5_mult_82_n6092,
         u5_mult_82_n6091, u5_mult_82_n6090, u5_mult_82_n6089,
         u5_mult_82_n6088, u5_mult_82_n6087, u5_mult_82_n6086,
         u5_mult_82_n6085, u5_mult_82_n6084, u5_mult_82_n6083,
         u5_mult_82_n6082, u5_mult_82_n6081, u5_mult_82_n6080,
         u5_mult_82_n6079, u5_mult_82_n6078, u5_mult_82_n6077,
         u5_mult_82_n6076, u5_mult_82_n6075, u5_mult_82_n6074,
         u5_mult_82_n6073, u5_mult_82_n6072, u5_mult_82_n6071,
         u5_mult_82_n6070, u5_mult_82_n6069, u5_mult_82_n6068,
         u5_mult_82_n6067, u5_mult_82_n6066, u5_mult_82_n6065,
         u5_mult_82_n6064, u5_mult_82_n6063, u5_mult_82_n6062,
         u5_mult_82_n6061, u5_mult_82_n6060, u5_mult_82_n6059,
         u5_mult_82_n6058, u5_mult_82_n6057, u5_mult_82_n6056,
         u5_mult_82_n6055, u5_mult_82_n6054, u5_mult_82_n6053,
         u5_mult_82_n6052, u5_mult_82_n6051, u5_mult_82_n6050,
         u5_mult_82_n6049, u5_mult_82_n6048, u5_mult_82_n6047,
         u5_mult_82_n6046, u5_mult_82_n6045, u5_mult_82_n6044,
         u5_mult_82_n6043, u5_mult_82_n6042, u5_mult_82_n6041,
         u5_mult_82_n6040, u5_mult_82_n6039, u5_mult_82_n6038,
         u5_mult_82_n6037, u5_mult_82_n6036, u5_mult_82_n6035,
         u5_mult_82_n6034, u5_mult_82_n6033, u5_mult_82_n6032,
         u5_mult_82_n6031, u5_mult_82_n6030, u5_mult_82_n6029,
         u5_mult_82_n6028, u5_mult_82_n6027, u5_mult_82_n6026,
         u5_mult_82_n6025, u5_mult_82_n6024, u5_mult_82_n6023,
         u5_mult_82_n6022, u5_mult_82_n6021, u5_mult_82_n6020,
         u5_mult_82_n6019, u5_mult_82_n6018, u5_mult_82_n6017,
         u5_mult_82_n6016, u5_mult_82_n6015, u5_mult_82_n6014,
         u5_mult_82_n6013, u5_mult_82_n6012, u5_mult_82_n6011,
         u5_mult_82_n6010, u5_mult_82_n6009, u5_mult_82_n6008,
         u5_mult_82_n6007, u5_mult_82_n6006, u5_mult_82_n6005,
         u5_mult_82_n6004, u5_mult_82_n6003, u5_mult_82_n6002,
         u5_mult_82_n6001, u5_mult_82_n6000, u5_mult_82_n5999,
         u5_mult_82_n5998, u5_mult_82_n5997, u5_mult_82_n5996,
         u5_mult_82_n5995, u5_mult_82_n5994, u5_mult_82_n5993,
         u5_mult_82_n5992, u5_mult_82_n5991, u5_mult_82_n5990,
         u5_mult_82_n5989, u5_mult_82_n5988, u5_mult_82_n5987,
         u5_mult_82_n5986, u5_mult_82_n5985, u5_mult_82_n5984,
         u5_mult_82_n5983, u5_mult_82_n5982, u5_mult_82_n5981,
         u5_mult_82_n5980, u5_mult_82_n5979, u5_mult_82_n5978,
         u5_mult_82_n5977, u5_mult_82_n5976, u5_mult_82_n5975,
         u5_mult_82_n5974, u5_mult_82_n5973, u5_mult_82_n5972,
         u5_mult_82_n5971, u5_mult_82_n5970, u5_mult_82_n5969,
         u5_mult_82_n5968, u5_mult_82_n5967, u5_mult_82_n5966,
         u5_mult_82_n5965, u5_mult_82_n5964, u5_mult_82_n5963,
         u5_mult_82_n5962, u5_mult_82_n5961, u5_mult_82_n5960,
         u5_mult_82_n5959, u5_mult_82_n5958, u5_mult_82_n5957,
         u5_mult_82_n5956, u5_mult_82_n5955, u5_mult_82_n5954,
         u5_mult_82_n5953, u5_mult_82_n5952, u5_mult_82_n5951,
         u5_mult_82_n5950, u5_mult_82_n5949, u5_mult_82_n5948,
         u5_mult_82_n5947, u5_mult_82_n5946, u5_mult_82_n5945,
         u5_mult_82_n5944, u5_mult_82_n5943, u5_mult_82_n5942,
         u5_mult_82_n5941, u5_mult_82_n5940, u5_mult_82_n5939,
         u5_mult_82_n5938, u5_mult_82_n5937, u5_mult_82_n5936,
         u5_mult_82_n5935, u5_mult_82_n5934, u5_mult_82_n5933,
         u5_mult_82_n5932, u5_mult_82_n5931, u5_mult_82_n5930,
         u5_mult_82_n5929, u5_mult_82_n5928, u5_mult_82_n5927,
         u5_mult_82_n5926, u5_mult_82_n5925, u5_mult_82_n5924,
         u5_mult_82_n5923, u5_mult_82_n5922, u5_mult_82_n5921,
         u5_mult_82_n5920, u5_mult_82_n5919, u5_mult_82_n5918,
         u5_mult_82_n5917, u5_mult_82_n5916, u5_mult_82_n5915,
         u5_mult_82_n5914, u5_mult_82_n5913, u5_mult_82_n5912,
         u5_mult_82_n5911, u5_mult_82_n5910, u5_mult_82_n5909,
         u5_mult_82_n5908, u5_mult_82_n5907, u5_mult_82_n5906,
         u5_mult_82_n5905, u5_mult_82_n5904, u5_mult_82_n5903,
         u5_mult_82_n5902, u5_mult_82_n5901, u5_mult_82_n5900,
         u5_mult_82_n5899, u5_mult_82_n5898, u5_mult_82_n5897,
         u5_mult_82_n5896, u5_mult_82_n5895, u5_mult_82_n5894,
         u5_mult_82_n5893, u5_mult_82_n5892, u5_mult_82_n5891,
         u5_mult_82_n5890, u5_mult_82_n5889, u5_mult_82_n5888,
         u5_mult_82_n5887, u5_mult_82_n5886, u5_mult_82_n5885,
         u5_mult_82_n5884, u5_mult_82_n5883, u5_mult_82_n5882,
         u5_mult_82_n5881, u5_mult_82_n5880, u5_mult_82_n5879,
         u5_mult_82_n5878, u5_mult_82_n5877, u5_mult_82_n5876,
         u5_mult_82_n5875, u5_mult_82_n5874, u5_mult_82_n5873,
         u5_mult_82_n5872, u5_mult_82_n5871, u5_mult_82_n5870,
         u5_mult_82_n5869, u5_mult_82_n5868, u5_mult_82_n5867,
         u5_mult_82_n5866, u5_mult_82_n5865, u5_mult_82_n5864,
         u5_mult_82_n5863, u5_mult_82_n5862, u5_mult_82_n5861,
         u5_mult_82_n5860, u5_mult_82_n5859, u5_mult_82_n5858,
         u5_mult_82_n5857, u5_mult_82_n5856, u5_mult_82_n5855,
         u5_mult_82_n5854, u5_mult_82_n5853, u5_mult_82_n5852,
         u5_mult_82_n5851, u5_mult_82_n5850, u5_mult_82_n5849,
         u5_mult_82_n5848, u5_mult_82_n5847, u5_mult_82_n5846,
         u5_mult_82_n5845, u5_mult_82_n5844, u5_mult_82_n5843,
         u5_mult_82_n5842, u5_mult_82_n5841, u5_mult_82_n5840,
         u5_mult_82_n5839, u5_mult_82_n5838, u5_mult_82_n5837,
         u5_mult_82_n5836, u5_mult_82_n5835, u5_mult_82_n5834,
         u5_mult_82_n5833, u5_mult_82_n5832, u5_mult_82_n5831,
         u5_mult_82_n5830, u5_mult_82_n5829, u5_mult_82_n5828,
         u5_mult_82_n5827, u5_mult_82_n5826, u5_mult_82_n5825,
         u5_mult_82_n5824, u5_mult_82_n5823, u5_mult_82_n5822,
         u5_mult_82_n5821, u5_mult_82_n5820, u5_mult_82_n5819,
         u5_mult_82_n5818, u5_mult_82_n5817, u5_mult_82_n5816,
         u5_mult_82_n5815, u5_mult_82_n5814, u5_mult_82_n5813,
         u5_mult_82_n5812, u5_mult_82_n5811, u5_mult_82_n5810,
         u5_mult_82_n5809, u5_mult_82_n5808, u5_mult_82_n5807,
         u5_mult_82_n5806, u5_mult_82_n5805, u5_mult_82_n5804,
         u5_mult_82_n5803, u5_mult_82_n5802, u5_mult_82_n5801,
         u5_mult_82_n5800, u5_mult_82_n5799, u5_mult_82_n5798,
         u5_mult_82_n5797, u5_mult_82_n5796, u5_mult_82_n5795,
         u5_mult_82_n5794, u5_mult_82_n5793, u5_mult_82_n5792,
         u5_mult_82_n5791, u5_mult_82_n5790, u5_mult_82_n5789,
         u5_mult_82_n5788, u5_mult_82_n5787, u5_mult_82_n5786,
         u5_mult_82_n5785, u5_mult_82_n5784, u5_mult_82_n5783,
         u5_mult_82_n5782, u5_mult_82_n5781, u5_mult_82_n5780,
         u5_mult_82_n5779, u5_mult_82_n5778, u5_mult_82_n5777,
         u5_mult_82_n5776, u5_mult_82_n5775, u5_mult_82_n5774,
         u5_mult_82_n5773, u5_mult_82_n5772, u5_mult_82_n5771,
         u5_mult_82_n5770, u5_mult_82_n5769, u5_mult_82_n5768,
         u5_mult_82_n5767, u5_mult_82_n5766, u5_mult_82_n5765,
         u5_mult_82_n5764, u5_mult_82_n5763, u5_mult_82_n5762,
         u5_mult_82_n5761, u5_mult_82_n5760, u5_mult_82_n5759,
         u5_mult_82_n5758, u5_mult_82_n5757, u5_mult_82_n5756,
         u5_mult_82_n5755, u5_mult_82_n5754, u5_mult_82_n5753,
         u5_mult_82_n5752, u5_mult_82_n5751, u5_mult_82_n5750,
         u5_mult_82_n5749, u5_mult_82_n5748, u5_mult_82_n5747,
         u5_mult_82_n5746, u5_mult_82_n5745, u5_mult_82_n5744,
         u5_mult_82_n5743, u5_mult_82_n5742, u5_mult_82_n5741,
         u5_mult_82_n5740, u5_mult_82_n5739, u5_mult_82_n5738,
         u5_mult_82_n5737, u5_mult_82_n5736, u5_mult_82_n5735,
         u5_mult_82_n5734, u5_mult_82_n5733, u5_mult_82_n5732,
         u5_mult_82_n5731, u5_mult_82_n5730, u5_mult_82_n5729,
         u5_mult_82_n5728, u5_mult_82_n5727, u5_mult_82_n5726,
         u5_mult_82_n5725, u5_mult_82_n5724, u5_mult_82_n5723,
         u5_mult_82_n5722, u5_mult_82_n5721, u5_mult_82_n5720,
         u5_mult_82_n5719, u5_mult_82_n5718, u5_mult_82_n5717,
         u5_mult_82_n5716, u5_mult_82_n5715, u5_mult_82_n5714,
         u5_mult_82_n5713, u5_mult_82_n5712, u5_mult_82_n5711,
         u5_mult_82_n5710, u5_mult_82_n5709, u5_mult_82_n5708,
         u5_mult_82_n5707, u5_mult_82_n5706, u5_mult_82_n5705,
         u5_mult_82_n5704, u5_mult_82_n5703, u5_mult_82_n5702,
         u5_mult_82_n5701, u5_mult_82_n5700, u5_mult_82_n5699,
         u5_mult_82_n5698, u5_mult_82_n5697, u5_mult_82_n5696,
         u5_mult_82_n5695, u5_mult_82_n5694, u5_mult_82_n5693,
         u5_mult_82_n5692, u5_mult_82_n5691, u5_mult_82_n5690,
         u5_mult_82_n5689, u5_mult_82_n5688, u5_mult_82_n5687,
         u5_mult_82_n5686, u5_mult_82_n5685, u5_mult_82_n5684,
         u5_mult_82_n5683, u5_mult_82_n5682, u5_mult_82_n5681,
         u5_mult_82_n5680, u5_mult_82_n5679, u5_mult_82_n5678,
         u5_mult_82_n5677, u5_mult_82_n5676, u5_mult_82_n5675,
         u5_mult_82_n5674, u5_mult_82_n5673, u5_mult_82_n5672,
         u5_mult_82_n5671, u5_mult_82_n5670, u5_mult_82_n5669,
         u5_mult_82_n5668, u5_mult_82_n5667, u5_mult_82_n5666,
         u5_mult_82_n5665, u5_mult_82_n5664, u5_mult_82_n5663,
         u5_mult_82_n5662, u5_mult_82_n5661, u5_mult_82_n5660,
         u5_mult_82_n5659, u5_mult_82_n5658, u5_mult_82_n5657,
         u5_mult_82_n5656, u5_mult_82_n5655, u5_mult_82_n5654,
         u5_mult_82_n5653, u5_mult_82_n5652, u5_mult_82_n5651,
         u5_mult_82_n5650, u5_mult_82_n5649, u5_mult_82_n5648,
         u5_mult_82_n5647, u5_mult_82_n5646, u5_mult_82_n5645,
         u5_mult_82_n5644, u5_mult_82_n5643, u5_mult_82_n5642,
         u5_mult_82_n5641, u5_mult_82_n5640, u5_mult_82_n5639,
         u5_mult_82_n5638, u5_mult_82_n5637, u5_mult_82_n5636,
         u5_mult_82_n5635, u5_mult_82_n5634, u5_mult_82_n5633,
         u5_mult_82_n5632, u5_mult_82_n5631, u5_mult_82_n5630,
         u5_mult_82_n5629, u5_mult_82_n5628, u5_mult_82_n5627,
         u5_mult_82_n5626, u5_mult_82_n5625, u5_mult_82_n5624,
         u5_mult_82_n5623, u5_mult_82_n5622, u5_mult_82_n5621,
         u5_mult_82_n5620, u5_mult_82_n5619, u5_mult_82_n5618,
         u5_mult_82_n5617, u5_mult_82_n5616, u5_mult_82_n5615,
         u5_mult_82_n5614, u5_mult_82_n5613, u5_mult_82_n5612,
         u5_mult_82_n5611, u5_mult_82_n5610, u5_mult_82_n5609,
         u5_mult_82_n5608, u5_mult_82_n5607, u5_mult_82_n5606,
         u5_mult_82_n5605, u5_mult_82_n5604, u5_mult_82_n5603,
         u5_mult_82_n5602, u5_mult_82_n5601, u5_mult_82_n5600,
         u5_mult_82_n5599, u5_mult_82_n5598, u5_mult_82_n5597,
         u5_mult_82_n5596, u5_mult_82_n5595, u5_mult_82_n5594,
         u5_mult_82_n5593, u5_mult_82_n5592, u5_mult_82_n5591,
         u5_mult_82_n5590, u5_mult_82_n5589, u5_mult_82_n5588,
         u5_mult_82_n5587, u5_mult_82_n5586, u5_mult_82_n5585,
         u5_mult_82_n5584, u5_mult_82_n5583, u5_mult_82_n5582,
         u5_mult_82_n5581, u5_mult_82_n5580, u5_mult_82_n5579,
         u5_mult_82_n5578, u5_mult_82_n5577, u5_mult_82_n5576,
         u5_mult_82_n5575, u5_mult_82_n5574, u5_mult_82_n5573,
         u5_mult_82_n5572, u5_mult_82_n5571, u5_mult_82_n5570,
         u5_mult_82_n5569, u5_mult_82_n5568, u5_mult_82_n5567,
         u5_mult_82_n5566, u5_mult_82_n5565, u5_mult_82_n5564,
         u5_mult_82_n5563, u5_mult_82_n5562, u5_mult_82_n5561,
         u5_mult_82_n5560, u5_mult_82_n5559, u5_mult_82_n5558,
         u5_mult_82_n5557, u5_mult_82_n5556, u5_mult_82_n5555,
         u5_mult_82_n5554, u5_mult_82_n5553, u5_mult_82_n5552,
         u5_mult_82_n5551, u5_mult_82_n5550, u5_mult_82_n5549,
         u5_mult_82_n5548, u5_mult_82_n5547, u5_mult_82_n5546,
         u5_mult_82_n5545, u5_mult_82_n5544, u5_mult_82_n5543,
         u5_mult_82_n5542, u5_mult_82_n5541, u5_mult_82_n5540,
         u5_mult_82_n5539, u5_mult_82_n5538, u5_mult_82_n5537,
         u5_mult_82_n5536, u5_mult_82_n5535, u5_mult_82_n5534,
         u5_mult_82_n5533, u5_mult_82_n5532, u5_mult_82_n5531,
         u5_mult_82_n5530, u5_mult_82_n5529, u5_mult_82_n5528,
         u5_mult_82_n5527, u5_mult_82_n5526, u5_mult_82_n5525,
         u5_mult_82_n5524, u5_mult_82_n5523, u5_mult_82_n5522,
         u5_mult_82_n5521, u5_mult_82_n5520, u5_mult_82_n5519,
         u5_mult_82_n5518, u5_mult_82_n5517, u5_mult_82_n5516,
         u5_mult_82_n5515, u5_mult_82_n5514, u5_mult_82_n5513,
         u5_mult_82_n5512, u5_mult_82_n5511, u5_mult_82_n5510,
         u5_mult_82_n5509, u5_mult_82_n5508, u5_mult_82_n5507,
         u5_mult_82_n5506, u5_mult_82_n5505, u5_mult_82_n5504,
         u5_mult_82_n5503, u5_mult_82_n5502, u5_mult_82_n5501,
         u5_mult_82_n5500, u5_mult_82_n5499, u5_mult_82_n5498,
         u5_mult_82_n5497, u5_mult_82_n5496, u5_mult_82_n5495,
         u5_mult_82_n5494, u5_mult_82_n5493, u5_mult_82_n5492,
         u5_mult_82_n5491, u5_mult_82_n5490, u5_mult_82_n5489,
         u5_mult_82_n5488, u5_mult_82_n5487, u5_mult_82_n5486,
         u5_mult_82_n5485, u5_mult_82_n5484, u5_mult_82_n5483,
         u5_mult_82_n5482, u5_mult_82_n5481, u5_mult_82_n5480,
         u5_mult_82_n5479, u5_mult_82_n5478, u5_mult_82_n5477,
         u5_mult_82_n5476, u5_mult_82_n5475, u5_mult_82_n5474,
         u5_mult_82_n5473, u5_mult_82_n5472, u5_mult_82_n5471,
         u5_mult_82_n5470, u5_mult_82_n5469, u5_mult_82_n5468,
         u5_mult_82_n5467, u5_mult_82_n5466, u5_mult_82_n5465,
         u5_mult_82_n5464, u5_mult_82_n5463, u5_mult_82_n5462,
         u5_mult_82_n5461, u5_mult_82_n5460, u5_mult_82_n5459,
         u5_mult_82_n5458, u5_mult_82_n5457, u5_mult_82_n5456,
         u5_mult_82_n5455, u5_mult_82_n5454, u5_mult_82_n5453,
         u5_mult_82_n5452, u5_mult_82_n5451, u5_mult_82_n5450,
         u5_mult_82_n5449, u5_mult_82_n5448, u5_mult_82_n5447,
         u5_mult_82_n5446, u5_mult_82_n5445, u5_mult_82_n5444,
         u5_mult_82_n5443, u5_mult_82_n5442, u5_mult_82_n5441,
         u5_mult_82_n5440, u5_mult_82_n5439, u5_mult_82_n5438,
         u5_mult_82_n5437, u5_mult_82_n5436, u5_mult_82_n5435,
         u5_mult_82_n5434, u5_mult_82_n5433, u5_mult_82_n5432,
         u5_mult_82_n5431, u5_mult_82_n5430, u5_mult_82_n5429,
         u5_mult_82_n5428, u5_mult_82_n5427, u5_mult_82_n5426,
         u5_mult_82_n5425, u5_mult_82_n5424, u5_mult_82_n5423,
         u5_mult_82_n5422, u5_mult_82_n5421, u5_mult_82_n5420,
         u5_mult_82_n5419, u5_mult_82_n5418, u5_mult_82_n5417,
         u5_mult_82_n5416, u5_mult_82_n5415, u5_mult_82_n5414,
         u5_mult_82_n5413, u5_mult_82_n5412, u5_mult_82_n5411,
         u5_mult_82_n5410, u5_mult_82_n5409, u5_mult_82_n5408,
         u5_mult_82_n5407, u5_mult_82_n5406, u5_mult_82_n5405,
         u5_mult_82_n5404, u5_mult_82_n5403, u5_mult_82_n5402,
         u5_mult_82_n5401, u5_mult_82_n5400, u5_mult_82_n5399,
         u5_mult_82_n5398, u5_mult_82_n5397, u5_mult_82_n5396,
         u5_mult_82_n5395, u5_mult_82_n5394, u5_mult_82_n5393,
         u5_mult_82_n5392, u5_mult_82_n5391, u5_mult_82_n5390,
         u5_mult_82_n5389, u5_mult_82_n5388, u5_mult_82_n5387,
         u5_mult_82_n5386, u5_mult_82_n5385, u5_mult_82_n5384,
         u5_mult_82_n5383, u5_mult_82_n5382, u5_mult_82_n5381,
         u5_mult_82_n5380, u5_mult_82_n5379, u5_mult_82_n5378,
         u5_mult_82_n5377, u5_mult_82_n5376, u5_mult_82_n5375,
         u5_mult_82_n5374, u5_mult_82_n5373, u5_mult_82_n5372,
         u5_mult_82_n5371, u5_mult_82_n5370, u5_mult_82_n5369,
         u5_mult_82_n5368, u5_mult_82_n5367, u5_mult_82_n5366,
         u5_mult_82_n5365, u5_mult_82_n5364, u5_mult_82_n5363,
         u5_mult_82_n5362, u5_mult_82_n5361, u5_mult_82_n5360,
         u5_mult_82_n5359, u5_mult_82_n5358, u5_mult_82_n5357,
         u5_mult_82_n5356, u5_mult_82_n5355, u5_mult_82_n5354,
         u5_mult_82_n5353, u5_mult_82_n5352, u5_mult_82_n5351,
         u5_mult_82_n5350, u5_mult_82_n5349, u5_mult_82_n5348,
         u5_mult_82_n5347, u5_mult_82_n5346, u5_mult_82_n5345,
         u5_mult_82_n5344, u5_mult_82_n5343, u5_mult_82_n5342,
         u5_mult_82_n5341, u5_mult_82_n5340, u5_mult_82_n5339,
         u5_mult_82_n5338, u5_mult_82_n5337, u5_mult_82_n5336,
         u5_mult_82_n5335, u5_mult_82_n5334, u5_mult_82_n5333,
         u5_mult_82_n5332, u5_mult_82_n5331, u5_mult_82_n5330,
         u5_mult_82_n5329, u5_mult_82_n5328, u5_mult_82_n5327,
         u5_mult_82_n5326, u5_mult_82_n5325, u5_mult_82_n5324,
         u5_mult_82_n5323, u5_mult_82_n5322, u5_mult_82_n5321,
         u5_mult_82_n5320, u5_mult_82_n5319, u5_mult_82_n5318,
         u5_mult_82_n5317, u5_mult_82_n5316, u5_mult_82_n5315,
         u5_mult_82_n5314, u5_mult_82_n5313, u5_mult_82_n5312,
         u5_mult_82_n5311, u5_mult_82_n5310, u5_mult_82_n5309,
         u5_mult_82_n5308, u5_mult_82_n5307, u5_mult_82_n5306,
         u5_mult_82_n5305, u5_mult_82_n5304, u5_mult_82_n5303,
         u5_mult_82_n5302, u5_mult_82_n5301, u5_mult_82_n5300,
         u5_mult_82_n5299, u5_mult_82_n5298, u5_mult_82_n5297,
         u5_mult_82_n5296, u5_mult_82_n5295, u5_mult_82_n5294,
         u5_mult_82_n5293, u5_mult_82_n5292, u5_mult_82_n5291,
         u5_mult_82_n5290, u5_mult_82_n5289, u5_mult_82_n5288,
         u5_mult_82_n5287, u5_mult_82_n5286, u5_mult_82_n5285,
         u5_mult_82_n5284, u5_mult_82_n5283, u5_mult_82_n5282,
         u5_mult_82_n5281, u5_mult_82_n5280, u5_mult_82_n5279,
         u5_mult_82_n5278, u5_mult_82_n5277, u5_mult_82_n5276,
         u5_mult_82_n5275, u5_mult_82_n5274, u5_mult_82_n5273,
         u5_mult_82_n5272, u5_mult_82_n5271, u5_mult_82_n5270,
         u5_mult_82_n5269, u5_mult_82_n5268, u5_mult_82_n5267,
         u5_mult_82_n5266, u5_mult_82_n5265, u5_mult_82_n5264,
         u5_mult_82_n5263, u5_mult_82_n5262, u5_mult_82_n5261,
         u5_mult_82_n5260, u5_mult_82_n5259, u5_mult_82_n5258,
         u5_mult_82_n5257, u5_mult_82_n5256, u5_mult_82_n5255,
         u5_mult_82_n5254, u5_mult_82_n5253, u5_mult_82_n5252,
         u5_mult_82_n5251, u5_mult_82_n5250, u5_mult_82_n5249,
         u5_mult_82_n5248, u5_mult_82_n5247, u5_mult_82_n5246,
         u5_mult_82_n5245, u5_mult_82_n5244, u5_mult_82_n5243,
         u5_mult_82_n5242, u5_mult_82_n5241, u5_mult_82_n5240,
         u5_mult_82_n5239, u5_mult_82_n5238, u5_mult_82_n5237,
         u5_mult_82_n5236, u5_mult_82_n5235, u5_mult_82_n5234,
         u5_mult_82_n5233, u5_mult_82_n5232, u5_mult_82_n5231,
         u5_mult_82_n5230, u5_mult_82_n5229, u5_mult_82_n5228,
         u5_mult_82_n5227, u5_mult_82_n5226, u5_mult_82_n5225,
         u5_mult_82_n5224, u5_mult_82_n5223, u5_mult_82_n5222,
         u5_mult_82_n5221, u5_mult_82_n5220, u5_mult_82_n5219,
         u5_mult_82_n5218, u5_mult_82_n5217, u5_mult_82_n5216,
         u5_mult_82_n5215, u5_mult_82_n5214, u5_mult_82_n5213,
         u5_mult_82_n5212, u5_mult_82_n5211, u5_mult_82_n5210,
         u5_mult_82_n5209, u5_mult_82_n5208, u5_mult_82_n5207,
         u5_mult_82_n5206, u5_mult_82_n5205, u5_mult_82_n5204,
         u5_mult_82_n5203, u5_mult_82_n5202, u5_mult_82_n5201,
         u5_mult_82_n5200, u5_mult_82_n5199, u5_mult_82_n5198,
         u5_mult_82_n5197, u5_mult_82_n5196, u5_mult_82_n5195,
         u5_mult_82_n5194, u5_mult_82_n5193, u5_mult_82_n5192,
         u5_mult_82_n5191, u5_mult_82_n5190, u5_mult_82_n5189,
         u5_mult_82_n5188, u5_mult_82_n5187, u5_mult_82_n5186,
         u5_mult_82_n5185, u5_mult_82_n5184, u5_mult_82_n5183,
         u5_mult_82_n5182, u5_mult_82_n5181, u5_mult_82_n5180,
         u5_mult_82_n5179, u5_mult_82_n5178, u5_mult_82_n5177,
         u5_mult_82_n5176, u5_mult_82_n5175, u5_mult_82_n5174,
         u5_mult_82_n5173, u5_mult_82_n5172, u5_mult_82_n5171,
         u5_mult_82_n5170, u5_mult_82_n5169, u5_mult_82_n5168,
         u5_mult_82_n5167, u5_mult_82_n5166, u5_mult_82_n5165,
         u5_mult_82_n5164, u5_mult_82_n5163, u5_mult_82_n5162,
         u5_mult_82_n5161, u5_mult_82_n5160, u5_mult_82_n5159,
         u5_mult_82_n5158, u5_mult_82_n5157, u5_mult_82_n5156,
         u5_mult_82_n5155, u5_mult_82_n5154, u5_mult_82_n5153,
         u5_mult_82_n5152, u5_mult_82_n5151, u5_mult_82_n5150,
         u5_mult_82_n5149, u5_mult_82_n5148, u5_mult_82_n5147,
         u5_mult_82_n5146, u5_mult_82_n5145, u5_mult_82_n5144,
         u5_mult_82_n5143, u5_mult_82_n5142, u5_mult_82_n5141,
         u5_mult_82_n5140, u5_mult_82_n5139, u5_mult_82_n5138,
         u5_mult_82_n5137, u5_mult_82_n5136, u5_mult_82_n5135,
         u5_mult_82_n5134, u5_mult_82_n5133, u5_mult_82_n5132,
         u5_mult_82_n5131, u5_mult_82_n5130, u5_mult_82_n5129,
         u5_mult_82_n5128, u5_mult_82_n5127, u5_mult_82_n5126,
         u5_mult_82_n5125, u5_mult_82_n5124, u5_mult_82_n5123,
         u5_mult_82_n5122, u5_mult_82_n5121, u5_mult_82_n5120,
         u5_mult_82_n5119, u5_mult_82_n5118, u5_mult_82_n5117,
         u5_mult_82_n5116, u5_mult_82_n5115, u5_mult_82_n5114,
         u5_mult_82_n5113, u5_mult_82_n5112, u5_mult_82_n5111,
         u5_mult_82_n5110, u5_mult_82_n5109, u5_mult_82_n5108,
         u5_mult_82_n5107, u5_mult_82_n5106, u5_mult_82_n5105,
         u5_mult_82_n5104, u5_mult_82_n5103, u5_mult_82_n5102,
         u5_mult_82_n5101, u5_mult_82_n5100, u5_mult_82_n5099,
         u5_mult_82_n5098, u5_mult_82_n5097, u5_mult_82_n5096,
         u5_mult_82_n5095, u5_mult_82_n5094, u5_mult_82_n5093,
         u5_mult_82_n5092, u5_mult_82_n5091, u5_mult_82_n5090,
         u5_mult_82_n5089, u5_mult_82_n5088, u5_mult_82_n5087,
         u5_mult_82_n5086, u5_mult_82_n5085, u5_mult_82_n5084,
         u5_mult_82_n5083, u5_mult_82_n5082, u5_mult_82_n5081,
         u5_mult_82_n5080, u5_mult_82_n5079, u5_mult_82_n5078,
         u5_mult_82_n5077, u5_mult_82_n5076, u5_mult_82_n5075,
         u5_mult_82_n5074, u5_mult_82_n5073, u5_mult_82_n5072,
         u5_mult_82_n5071, u5_mult_82_n5070, u5_mult_82_n5069,
         u5_mult_82_n5068, u5_mult_82_n5067, u5_mult_82_n5066,
         u5_mult_82_n5065, u5_mult_82_n5064, u5_mult_82_n5063,
         u5_mult_82_n5062, u5_mult_82_n5061, u5_mult_82_n5060,
         u5_mult_82_n5059, u5_mult_82_n5058, u5_mult_82_n5057,
         u5_mult_82_n5056, u5_mult_82_n5055, u5_mult_82_n5054,
         u5_mult_82_n5053, u5_mult_82_n5052, u5_mult_82_n5051,
         u5_mult_82_n5050, u5_mult_82_n5049, u5_mult_82_n5048,
         u5_mult_82_n5047, u5_mult_82_n5046, u5_mult_82_n5045,
         u5_mult_82_n5044, u5_mult_82_n5043, u5_mult_82_n5042,
         u5_mult_82_n5041, u5_mult_82_n5040, u5_mult_82_n5039,
         u5_mult_82_n5038, u5_mult_82_n5037, u5_mult_82_n5036,
         u5_mult_82_n5035, u5_mult_82_n5034, u5_mult_82_n5033,
         u5_mult_82_n5032, u5_mult_82_n5031, u5_mult_82_n5030,
         u5_mult_82_n5029, u5_mult_82_n5028, u5_mult_82_n5027,
         u5_mult_82_n5026, u5_mult_82_n5025, u5_mult_82_n5024,
         u5_mult_82_n5023, u5_mult_82_n5022, u5_mult_82_n5021,
         u5_mult_82_n5020, u5_mult_82_n5019, u5_mult_82_n5018,
         u5_mult_82_n5017, u5_mult_82_n5016, u5_mult_82_n5015,
         u5_mult_82_n5014, u5_mult_82_n5013, u5_mult_82_n5012,
         u5_mult_82_n5011, u5_mult_82_n5010, u5_mult_82_n5009,
         u5_mult_82_n5008, u5_mult_82_n5007, u5_mult_82_n5006,
         u5_mult_82_n5005, u5_mult_82_n5004, u5_mult_82_n5003,
         u5_mult_82_n5002, u5_mult_82_n5001, u5_mult_82_n5000,
         u5_mult_82_n4999, u5_mult_82_n4998, u5_mult_82_n4997,
         u5_mult_82_n4996, u5_mult_82_n4995, u5_mult_82_n4994,
         u5_mult_82_n4993, u5_mult_82_n4992, u5_mult_82_n4991,
         u5_mult_82_n4990, u5_mult_82_n4989, u5_mult_82_n4988,
         u5_mult_82_n4987, u5_mult_82_n4986, u5_mult_82_n4985,
         u5_mult_82_n4984, u5_mult_82_n4983, u5_mult_82_n4982,
         u5_mult_82_n4981, u5_mult_82_n4980, u5_mult_82_n4979,
         u5_mult_82_n4978, u5_mult_82_n4977, u5_mult_82_n4976,
         u5_mult_82_n4975, u5_mult_82_n4974, u5_mult_82_n4973,
         u5_mult_82_n4972, u5_mult_82_n4971, u5_mult_82_n4970,
         u5_mult_82_n4969, u5_mult_82_n4968, u5_mult_82_n4967,
         u5_mult_82_n4966, u5_mult_82_n4965, u5_mult_82_n4964,
         u5_mult_82_n4963, u5_mult_82_n4962, u5_mult_82_n4961,
         u5_mult_82_n4960, u5_mult_82_n4959, u5_mult_82_n4958,
         u5_mult_82_n4957, u5_mult_82_n4956, u5_mult_82_n4955,
         u5_mult_82_n4954, u5_mult_82_n4953, u5_mult_82_n4952,
         u5_mult_82_n4951, u5_mult_82_n4950, u5_mult_82_n4949,
         u5_mult_82_n4948, u5_mult_82_n4947, u5_mult_82_n4946,
         u5_mult_82_n4945, u5_mult_82_n4944, u5_mult_82_n4943,
         u5_mult_82_n4942, u5_mult_82_n4941, u5_mult_82_n4940,
         u5_mult_82_n4939, u5_mult_82_n4938, u5_mult_82_n4937,
         u5_mult_82_n4936, u5_mult_82_n4935, u5_mult_82_n4934,
         u5_mult_82_n4933, u5_mult_82_n4932, u5_mult_82_n4931,
         u5_mult_82_n4930, u5_mult_82_n4929, u5_mult_82_n4928,
         u5_mult_82_n4927, u5_mult_82_n4926, u5_mult_82_n4925,
         u5_mult_82_n4924, u5_mult_82_n4923, u5_mult_82_n4922,
         u5_mult_82_n4921, u5_mult_82_n4920, u5_mult_82_n4919,
         u5_mult_82_n4918, u5_mult_82_n4917, u5_mult_82_n4916,
         u5_mult_82_n4915, u5_mult_82_n4914, u5_mult_82_n4913,
         u5_mult_82_n4912, u5_mult_82_n4911, u5_mult_82_n4910,
         u5_mult_82_n4909, u5_mult_82_n4908, u5_mult_82_n4907,
         u5_mult_82_n4906, u5_mult_82_n4905, u5_mult_82_n4904,
         u5_mult_82_n4903, u5_mult_82_n4902, u5_mult_82_n4901,
         u5_mult_82_n4900, u5_mult_82_n4899, u5_mult_82_n4898,
         u5_mult_82_n4897, u5_mult_82_n4896, u5_mult_82_n4895,
         u5_mult_82_n4894, u5_mult_82_n4893, u5_mult_82_n4892,
         u5_mult_82_n4891, u5_mult_82_n4890, u5_mult_82_n4889,
         u5_mult_82_n4888, u5_mult_82_n4887, u5_mult_82_n4886,
         u5_mult_82_n4885, u5_mult_82_n4884, u5_mult_82_n4883,
         u5_mult_82_n4882, u5_mult_82_n4881, u5_mult_82_n4880,
         u5_mult_82_n4879, u5_mult_82_n4878, u5_mult_82_n4877,
         u5_mult_82_n4876, u5_mult_82_n4875, u5_mult_82_n4874,
         u5_mult_82_n4873, u5_mult_82_n4872, u5_mult_82_n4871,
         u5_mult_82_n4870, u5_mult_82_n4869, u5_mult_82_n4868,
         u5_mult_82_n4867, u5_mult_82_n4866, u5_mult_82_n4865,
         u5_mult_82_n4864, u5_mult_82_n4863, u5_mult_82_n4862,
         u5_mult_82_n4861, u5_mult_82_n4860, u5_mult_82_n4859,
         u5_mult_82_n4858, u5_mult_82_n4857, u5_mult_82_n4856,
         u5_mult_82_n4855, u5_mult_82_n4854, u5_mult_82_n4853,
         u5_mult_82_n4852, u5_mult_82_n4851, u5_mult_82_n4850,
         u5_mult_82_n4849, u5_mult_82_n4848, u5_mult_82_n4847,
         u5_mult_82_n4846, u5_mult_82_n4845, u5_mult_82_n4844,
         u5_mult_82_n4843, u5_mult_82_n4842, u5_mult_82_n4841,
         u5_mult_82_n4840, u5_mult_82_n4839, u5_mult_82_n4838,
         u5_mult_82_n4837, u5_mult_82_n4836, u5_mult_82_n4835,
         u5_mult_82_n4834, u5_mult_82_n4833, u5_mult_82_n4832,
         u5_mult_82_n4831, u5_mult_82_n4830, u5_mult_82_n4829,
         u5_mult_82_n4828, u5_mult_82_n4827, u5_mult_82_n4826,
         u5_mult_82_n4825, u5_mult_82_n4824, u5_mult_82_n4823,
         u5_mult_82_n4822, u5_mult_82_n4821, u5_mult_82_n4820,
         u5_mult_82_n4819, u5_mult_82_n4818, u5_mult_82_n4817,
         u5_mult_82_n4816, u5_mult_82_n4815, u5_mult_82_n4814,
         u5_mult_82_n4813, u5_mult_82_n4812, u5_mult_82_n4811,
         u5_mult_82_n4810, u5_mult_82_n4809, u5_mult_82_n4808,
         u5_mult_82_n4807, u5_mult_82_n4806, u5_mult_82_n4805,
         u5_mult_82_n4804, u5_mult_82_n4803, u5_mult_82_n4802,
         u5_mult_82_n4801, u5_mult_82_n4800, u5_mult_82_n4799,
         u5_mult_82_n4798, u5_mult_82_n4797, u5_mult_82_n4796,
         u5_mult_82_n4795, u5_mult_82_n4794, u5_mult_82_n4793,
         u5_mult_82_n4792, u5_mult_82_n4791, u5_mult_82_n4790,
         u5_mult_82_n4789, u5_mult_82_n4788, u5_mult_82_n4787,
         u5_mult_82_n4786, u5_mult_82_n4785, u5_mult_82_n4784,
         u5_mult_82_n4783, u5_mult_82_n4782, u5_mult_82_n4781,
         u5_mult_82_n4780, u5_mult_82_n4779, u5_mult_82_n4778,
         u5_mult_82_n4777, u5_mult_82_n4776, u5_mult_82_n4775,
         u5_mult_82_n4774, u5_mult_82_n4773, u5_mult_82_n4772,
         u5_mult_82_n4771, u5_mult_82_n4770, u5_mult_82_n4769,
         u5_mult_82_n4768, u5_mult_82_n4767, u5_mult_82_n4766,
         u5_mult_82_n4765, u5_mult_82_n4764, u5_mult_82_n4763,
         u5_mult_82_n4762, u5_mult_82_n4761, u5_mult_82_n4760,
         u5_mult_82_n4759, u5_mult_82_n4758, u5_mult_82_n4757,
         u5_mult_82_n4756, u5_mult_82_n4755, u5_mult_82_n4754,
         u5_mult_82_n4753, u5_mult_82_n4752, u5_mult_82_n4751,
         u5_mult_82_n4750, u5_mult_82_n4749, u5_mult_82_n4748,
         u5_mult_82_n4747, u5_mult_82_n4746, u5_mult_82_n4745,
         u5_mult_82_n4744, u5_mult_82_n4743, u5_mult_82_n4742,
         u5_mult_82_n4741, u5_mult_82_n4740, u5_mult_82_n4739,
         u5_mult_82_n4738, u5_mult_82_n4737, u5_mult_82_n4736,
         u5_mult_82_n4735, u5_mult_82_n4734, u5_mult_82_n4733,
         u5_mult_82_n4732, u5_mult_82_n4731, u5_mult_82_n4730,
         u5_mult_82_n4729, u5_mult_82_n4728, u5_mult_82_n4727,
         u5_mult_82_n4726, u5_mult_82_n4725, u5_mult_82_n4724,
         u5_mult_82_n4723, u5_mult_82_n4722, u5_mult_82_n4721,
         u5_mult_82_n4720, u5_mult_82_n4719, u5_mult_82_n4718,
         u5_mult_82_n4717, u5_mult_82_n4716, u5_mult_82_n4715,
         u5_mult_82_n4714, u5_mult_82_n4713, u5_mult_82_n4712,
         u5_mult_82_n4711, u5_mult_82_n4710, u5_mult_82_n4709,
         u5_mult_82_n4708, u5_mult_82_n4707, u5_mult_82_n4706,
         u5_mult_82_n4705, u5_mult_82_n4704, u5_mult_82_n4703,
         u5_mult_82_n4702, u5_mult_82_n4701, u5_mult_82_n4700,
         u5_mult_82_n4699, u5_mult_82_n4698, u5_mult_82_n4697,
         u5_mult_82_n4696, u5_mult_82_n4695, u5_mult_82_n4694,
         u5_mult_82_n4693, u5_mult_82_n4692, u5_mult_82_n4691,
         u5_mult_82_n4690, u5_mult_82_n4689, u5_mult_82_n4688,
         u5_mult_82_n4687, u5_mult_82_n4686, u5_mult_82_n4685,
         u5_mult_82_n4684, u5_mult_82_n4683, u5_mult_82_n4682,
         u5_mult_82_n4681, u5_mult_82_n4680, u5_mult_82_n4679,
         u5_mult_82_n4678, u5_mult_82_n4677, u5_mult_82_n4676,
         u5_mult_82_n4675, u5_mult_82_n4674, u5_mult_82_n4673,
         u5_mult_82_n4672, u5_mult_82_n4671, u5_mult_82_n4670,
         u5_mult_82_n4669, u5_mult_82_n4668, u5_mult_82_n4667,
         u5_mult_82_n4666, u5_mult_82_n4665, u5_mult_82_n4664,
         u5_mult_82_n4663, u5_mult_82_n4662, u5_mult_82_n4661,
         u5_mult_82_n4660, u5_mult_82_n4659, u5_mult_82_n4658,
         u5_mult_82_n4657, u5_mult_82_n4656, u5_mult_82_n4655,
         u5_mult_82_n4654, u5_mult_82_n4653, u5_mult_82_n4652,
         u5_mult_82_n4651, u5_mult_82_n4650, u5_mult_82_n4649,
         u5_mult_82_n4648, u5_mult_82_n4647, u5_mult_82_n4646,
         u5_mult_82_n4645, u5_mult_82_n4644, u5_mult_82_n4643,
         u5_mult_82_n4642, u5_mult_82_n4641, u5_mult_82_n4640,
         u5_mult_82_n4639, u5_mult_82_n4638, u5_mult_82_n4637,
         u5_mult_82_n4636, u5_mult_82_n4635, u5_mult_82_n4634,
         u5_mult_82_n4633, u5_mult_82_n4632, u5_mult_82_n4631,
         u5_mult_82_n4630, u5_mult_82_n4629, u5_mult_82_n4628,
         u5_mult_82_n4627, u5_mult_82_n4626, u5_mult_82_n4625,
         u5_mult_82_n4624, u5_mult_82_n4623, u5_mult_82_n4622,
         u5_mult_82_n4621, u5_mult_82_n4620, u5_mult_82_n4619,
         u5_mult_82_n4618, u5_mult_82_n4617, u5_mult_82_n4616,
         u5_mult_82_n4615, u5_mult_82_n4614, u5_mult_82_n4613,
         u5_mult_82_n4612, u5_mult_82_n4611, u5_mult_82_n4610,
         u5_mult_82_n4609, u5_mult_82_n4608, u5_mult_82_n4607,
         u5_mult_82_n4606, u5_mult_82_n4605, u5_mult_82_n4604,
         u5_mult_82_n4603, u5_mult_82_n4602, u5_mult_82_n4601,
         u5_mult_82_n4600, u5_mult_82_n4599, u5_mult_82_n4598,
         u5_mult_82_n4597, u5_mult_82_n4596, u5_mult_82_n4595,
         u5_mult_82_n4594, u5_mult_82_n4593, u5_mult_82_n4592,
         u5_mult_82_n4591, u5_mult_82_n4590, u5_mult_82_n4589,
         u5_mult_82_n4588, u5_mult_82_n4587, u5_mult_82_n4586,
         u5_mult_82_n4585, u5_mult_82_n4584, u5_mult_82_n4583,
         u5_mult_82_n4582, u5_mult_82_n4581, u5_mult_82_n4580,
         u5_mult_82_n4579, u5_mult_82_n4578, u5_mult_82_n4577,
         u5_mult_82_n4576, u5_mult_82_n4575, u5_mult_82_n4574,
         u5_mult_82_n4573, u5_mult_82_n4572, u5_mult_82_n4571,
         u5_mult_82_n4570, u5_mult_82_n4569, u5_mult_82_n4568,
         u5_mult_82_n4567, u5_mult_82_n4566, u5_mult_82_n4565,
         u5_mult_82_n4564, u5_mult_82_n4563, u5_mult_82_n4562,
         u5_mult_82_n4561, u5_mult_82_n4560, u5_mult_82_n4559,
         u5_mult_82_n4558, u5_mult_82_n4557, u5_mult_82_n4556,
         u5_mult_82_n4555, u5_mult_82_n4554, u5_mult_82_n4553,
         u5_mult_82_n4552, u5_mult_82_n4551, u5_mult_82_n4550,
         u5_mult_82_n4549, u5_mult_82_n4548, u5_mult_82_n4547,
         u5_mult_82_n4546, u5_mult_82_n4545, u5_mult_82_n4544,
         u5_mult_82_n4543, u5_mult_82_n4542, u5_mult_82_n4541,
         u5_mult_82_n4540, u5_mult_82_n4539, u5_mult_82_n4538,
         u5_mult_82_n4537, u5_mult_82_n4536, u5_mult_82_n4535,
         u5_mult_82_n4534, u5_mult_82_n4533, u5_mult_82_n4532,
         u5_mult_82_n4531, u5_mult_82_n4530, u5_mult_82_n4529,
         u5_mult_82_n4528, u5_mult_82_n4527, u5_mult_82_n4526,
         u5_mult_82_n4525, u5_mult_82_n4524, u5_mult_82_n4523,
         u5_mult_82_n4522, u5_mult_82_n4521, u5_mult_82_n4520,
         u5_mult_82_n4519, u5_mult_82_n4518, u5_mult_82_n4517,
         u5_mult_82_n4516, u5_mult_82_n4515, u5_mult_82_n4514,
         u5_mult_82_n4513, u5_mult_82_n4512, u5_mult_82_n4511,
         u5_mult_82_n4510, u5_mult_82_n4509, u5_mult_82_n4508,
         u5_mult_82_n4507, u5_mult_82_n4506, u5_mult_82_n4505,
         u5_mult_82_n4504, u5_mult_82_n4503, u5_mult_82_n4502,
         u5_mult_82_n4501, u5_mult_82_n4500, u5_mult_82_n4499,
         u5_mult_82_n4498, u5_mult_82_n4497, u5_mult_82_n4496,
         u5_mult_82_n4495, u5_mult_82_n4494, u5_mult_82_n4493,
         u5_mult_82_n4492, u5_mult_82_n4491, u5_mult_82_n4490,
         u5_mult_82_n4489, u5_mult_82_n4488, u5_mult_82_n4487,
         u5_mult_82_n4486, u5_mult_82_n4485, u5_mult_82_n4484,
         u5_mult_82_n4483, u5_mult_82_n4482, u5_mult_82_n4481,
         u5_mult_82_n4480, u5_mult_82_n4479, u5_mult_82_n4478,
         u5_mult_82_n4477, u5_mult_82_n4476, u5_mult_82_n4475,
         u5_mult_82_n4474, u5_mult_82_n4473, u5_mult_82_n4472,
         u5_mult_82_n4471, u5_mult_82_n4470, u5_mult_82_n4469,
         u5_mult_82_n4468, u5_mult_82_n4467, u5_mult_82_n4466,
         u5_mult_82_n4465, u5_mult_82_n4464, u5_mult_82_n4463,
         u5_mult_82_n4462, u5_mult_82_n4461, u5_mult_82_n4460,
         u5_mult_82_n4459, u5_mult_82_n4458, u5_mult_82_n4457,
         u5_mult_82_n4456, u5_mult_82_n4455, u5_mult_82_n4454,
         u5_mult_82_n4453, u5_mult_82_n4452, u5_mult_82_n4451,
         u5_mult_82_n4450, u5_mult_82_n4449, u5_mult_82_n4448,
         u5_mult_82_n4447, u5_mult_82_n4446, u5_mult_82_n4445,
         u5_mult_82_n4444, u5_mult_82_n4443, u5_mult_82_n4442,
         u5_mult_82_n4441, u5_mult_82_n4440, u5_mult_82_n4439,
         u5_mult_82_n4438, u5_mult_82_n4437, u5_mult_82_n4436,
         u5_mult_82_n4435, u5_mult_82_n4434, u5_mult_82_n4433,
         u5_mult_82_n4432, u5_mult_82_n4431, u5_mult_82_n4430,
         u5_mult_82_n4429, u5_mult_82_n4428, u5_mult_82_n4427,
         u5_mult_82_n4426, u5_mult_82_n4425, u5_mult_82_n4424,
         u5_mult_82_n4423, u5_mult_82_n4422, u5_mult_82_n4421,
         u5_mult_82_n4420, u5_mult_82_n4419, u5_mult_82_n4418,
         u5_mult_82_n4417, u5_mult_82_n4416, u5_mult_82_n4415,
         u5_mult_82_n4414, u5_mult_82_n4413, u5_mult_82_n4412,
         u5_mult_82_n4411, u5_mult_82_n4410, u5_mult_82_n4409,
         u5_mult_82_n4408, u5_mult_82_n4407, u5_mult_82_n4406,
         u5_mult_82_n4405, u5_mult_82_n4404, u5_mult_82_n4403,
         u5_mult_82_n4402, u5_mult_82_n4401, u5_mult_82_n4400,
         u5_mult_82_n4399, u5_mult_82_n4398, u5_mult_82_n4397,
         u5_mult_82_n4396, u5_mult_82_n4395, u5_mult_82_n4394,
         u5_mult_82_n4393, u5_mult_82_n4392, u5_mult_82_n4391,
         u5_mult_82_n4390, u5_mult_82_n4389, u5_mult_82_n4388,
         u5_mult_82_n4387, u5_mult_82_n4386, u5_mult_82_n4385,
         u5_mult_82_n4384, u5_mult_82_n4383, u5_mult_82_n4382,
         u5_mult_82_n4381, u5_mult_82_n4380, u5_mult_82_n4379,
         u5_mult_82_n4378, u5_mult_82_n4377, u5_mult_82_n4376,
         u5_mult_82_n4375, u5_mult_82_n4374, u5_mult_82_n4373,
         u5_mult_82_n4372, u5_mult_82_n4371, u5_mult_82_n4370,
         u5_mult_82_n4369, u5_mult_82_n4368, u5_mult_82_n4367,
         u5_mult_82_n4366, u5_mult_82_n4365, u5_mult_82_n4364,
         u5_mult_82_n4363, u5_mult_82_n4362, u5_mult_82_n4361,
         u5_mult_82_n4360, u5_mult_82_n4359, u5_mult_82_n4358,
         u5_mult_82_n4357, u5_mult_82_n4356, u5_mult_82_n4355,
         u5_mult_82_n4354, u5_mult_82_n4353, u5_mult_82_n4352,
         u5_mult_82_n4351, u5_mult_82_n4350, u5_mult_82_n4349,
         u5_mult_82_n4348, u5_mult_82_n4347, u5_mult_82_n4346,
         u5_mult_82_n4345, u5_mult_82_n4344, u5_mult_82_n4343,
         u5_mult_82_n4342, u5_mult_82_n4341, u5_mult_82_n4340,
         u5_mult_82_n4339, u5_mult_82_n4338, u5_mult_82_n4337,
         u5_mult_82_n4336, u5_mult_82_n4335, u5_mult_82_n4334,
         u5_mult_82_n4333, u5_mult_82_n4332, u5_mult_82_n4331,
         u5_mult_82_n4330, u5_mult_82_n4329, u5_mult_82_n4328,
         u5_mult_82_n4327, u5_mult_82_n4326, u5_mult_82_n4325,
         u5_mult_82_n4324, u5_mult_82_n4323, u5_mult_82_n4322,
         u5_mult_82_n4321, u5_mult_82_n4320, u5_mult_82_n4319,
         u5_mult_82_n4318, u5_mult_82_n4317, u5_mult_82_n4316,
         u5_mult_82_n4315, u5_mult_82_n4314, u5_mult_82_n4313,
         u5_mult_82_n4312, u5_mult_82_n4311, u5_mult_82_n4310,
         u5_mult_82_n4309, u5_mult_82_n4308, u5_mult_82_n4307,
         u5_mult_82_n4306, u5_mult_82_n4305, u5_mult_82_n4304,
         u5_mult_82_n4303, u5_mult_82_n4302, u5_mult_82_n4301,
         u5_mult_82_n4300, u5_mult_82_n4299, u5_mult_82_n4298,
         u5_mult_82_n4297, u5_mult_82_n4296, u5_mult_82_n4295,
         u5_mult_82_n4294, u5_mult_82_n4293, u5_mult_82_n4292,
         u5_mult_82_n4291, u5_mult_82_n4290, u5_mult_82_n4289,
         u5_mult_82_n4288, u5_mult_82_n4287, u5_mult_82_n4286,
         u5_mult_82_n4285, u5_mult_82_n4284, u5_mult_82_n4283,
         u5_mult_82_n4282, u5_mult_82_n4281, u5_mult_82_n4280,
         u5_mult_82_n4279, u5_mult_82_n4278, u5_mult_82_n4277,
         u5_mult_82_n4276, u5_mult_82_n4275, u5_mult_82_n4274,
         u5_mult_82_n4273, u5_mult_82_n4272, u5_mult_82_n4271,
         u5_mult_82_n4270, u5_mult_82_n4269, u5_mult_82_n4268,
         u5_mult_82_n4267, u5_mult_82_n4266, u5_mult_82_n4265,
         u5_mult_82_n4264, u5_mult_82_n4263, u5_mult_82_n4262,
         u5_mult_82_n4261, u5_mult_82_n4260, u5_mult_82_n4259,
         u5_mult_82_n4258, u5_mult_82_n4257, u5_mult_82_n4256,
         u5_mult_82_n4255, u5_mult_82_n4254, u5_mult_82_n4253,
         u5_mult_82_n4252, u5_mult_82_n4251, u5_mult_82_n4250,
         u5_mult_82_n4249, u5_mult_82_n4248, u5_mult_82_n4247,
         u5_mult_82_n4246, u5_mult_82_n4245, u5_mult_82_n4244,
         u5_mult_82_n4243, u5_mult_82_n4242, u5_mult_82_n4241,
         u5_mult_82_n4240, u5_mult_82_n4239, u5_mult_82_n4238,
         u5_mult_82_n4237, u5_mult_82_n4236, u5_mult_82_n4235,
         u5_mult_82_n4234, u5_mult_82_n4233, u5_mult_82_n4232,
         u5_mult_82_n4231, u5_mult_82_n4230, u5_mult_82_n4229,
         u5_mult_82_n4228, u5_mult_82_n4227, u5_mult_82_n4226,
         u5_mult_82_n4225, u5_mult_82_n4224, u5_mult_82_n4223,
         u5_mult_82_n4222, u5_mult_82_n4221, u5_mult_82_n4220,
         u5_mult_82_n4219, u5_mult_82_n4218, u5_mult_82_n4217,
         u5_mult_82_n4216, u5_mult_82_n4215, u5_mult_82_n4214,
         u5_mult_82_n4213, u5_mult_82_n4212, u5_mult_82_n4211,
         u5_mult_82_n4210, u5_mult_82_n4209, u5_mult_82_n4208,
         u5_mult_82_n4207, u5_mult_82_n4206, u5_mult_82_n4205,
         u5_mult_82_n4204, u5_mult_82_n4203, u5_mult_82_n4202,
         u5_mult_82_n4201, u5_mult_82_n4200, u5_mult_82_n4199,
         u5_mult_82_n4198, u5_mult_82_n4197, u5_mult_82_n4196,
         u5_mult_82_n4195, u5_mult_82_n4194, u5_mult_82_n4193,
         u5_mult_82_n4192, u5_mult_82_n4191, u5_mult_82_n4190,
         u5_mult_82_n4189, u5_mult_82_n4188, u5_mult_82_n4187,
         u5_mult_82_n4186, u5_mult_82_n4185, u5_mult_82_n4184,
         u5_mult_82_n4183, u5_mult_82_n4182, u5_mult_82_n4181,
         u5_mult_82_n4180, u5_mult_82_n4179, u5_mult_82_n4178,
         u5_mult_82_n4177, u5_mult_82_n4176, u5_mult_82_n4175,
         u5_mult_82_n4174, u5_mult_82_n4173, u5_mult_82_n4172,
         u5_mult_82_n4171, u5_mult_82_n4170, u5_mult_82_n4169,
         u5_mult_82_n4168, u5_mult_82_n4167, u5_mult_82_n4166,
         u5_mult_82_n4165, u5_mult_82_n4164, u5_mult_82_n4163,
         u5_mult_82_n4162, u5_mult_82_n4161, u5_mult_82_n4160,
         u5_mult_82_n4159, u5_mult_82_n4158, u5_mult_82_n4157,
         u5_mult_82_n4156, u5_mult_82_n4155, u5_mult_82_n4154,
         u5_mult_82_n4153, u5_mult_82_n4152, u5_mult_82_n4151,
         u5_mult_82_n4150, u5_mult_82_n4149, u5_mult_82_n4148,
         u5_mult_82_n4147, u5_mult_82_n4146, u5_mult_82_n4145,
         u5_mult_82_n4144, u5_mult_82_n4143, u5_mult_82_n4142,
         u5_mult_82_n4141, u5_mult_82_n4140, u5_mult_82_n4139,
         u5_mult_82_n4138, u5_mult_82_n4137, u5_mult_82_n4136,
         u5_mult_82_n4135, u5_mult_82_n4134, u5_mult_82_n4133,
         u5_mult_82_n4132, u5_mult_82_n4131, u5_mult_82_n4130,
         u5_mult_82_n4129, u5_mult_82_n4128, u5_mult_82_n4127,
         u5_mult_82_n4126, u5_mult_82_n4125, u5_mult_82_n4124,
         u5_mult_82_n4123, u5_mult_82_n4122, u5_mult_82_n4121,
         u5_mult_82_n4120, u5_mult_82_n4119, u5_mult_82_n4118,
         u5_mult_82_n4117, u5_mult_82_n4116, u5_mult_82_n4115,
         u5_mult_82_n4114, u5_mult_82_n4113, u5_mult_82_n4112,
         u5_mult_82_n4111, u5_mult_82_n4110, u5_mult_82_n4109,
         u5_mult_82_n4108, u5_mult_82_n4107, u5_mult_82_n4106,
         u5_mult_82_n4105, u5_mult_82_n4104, u5_mult_82_n4103,
         u5_mult_82_n4102, u5_mult_82_n4101, u5_mult_82_n4100,
         u5_mult_82_n4099, u5_mult_82_n4098, u5_mult_82_n4097,
         u5_mult_82_n4096, u5_mult_82_n4095, u5_mult_82_n4094,
         u5_mult_82_n4093, u5_mult_82_n4092, u5_mult_82_n4091,
         u5_mult_82_n4090, u5_mult_82_n4089, u5_mult_82_n4088,
         u5_mult_82_n4087, u5_mult_82_n4086, u5_mult_82_n4085,
         u5_mult_82_n4084, u5_mult_82_n4083, u5_mult_82_n4082,
         u5_mult_82_n4081, u5_mult_82_n4080, u5_mult_82_n4079,
         u5_mult_82_n4078, u5_mult_82_n4077, u5_mult_82_n4076,
         u5_mult_82_n4075, u5_mult_82_n4074, u5_mult_82_n4073,
         u5_mult_82_n4072, u5_mult_82_n4071, u5_mult_82_n4070,
         u5_mult_82_n4069, u5_mult_82_n4068, u5_mult_82_n4067,
         u5_mult_82_n4066, u5_mult_82_n4065, u5_mult_82_n4064,
         u5_mult_82_n4063, u5_mult_82_n4062, u5_mult_82_n4061,
         u5_mult_82_n4060, u5_mult_82_n4059, u5_mult_82_n4058,
         u5_mult_82_n4057, u5_mult_82_n4056, u5_mult_82_n4055,
         u5_mult_82_n4054, u5_mult_82_n4053, u5_mult_82_n4052,
         u5_mult_82_n4051, u5_mult_82_n4050, u5_mult_82_n4049,
         u5_mult_82_n4048, u5_mult_82_n4047, u5_mult_82_n4046,
         u5_mult_82_n4045, u5_mult_82_n4044, u5_mult_82_n4043,
         u5_mult_82_n4042, u5_mult_82_n4041, u5_mult_82_n4040,
         u5_mult_82_n4039, u5_mult_82_n4038, u5_mult_82_n4037,
         u5_mult_82_n4036, u5_mult_82_n4035, u5_mult_82_n4034,
         u5_mult_82_n4033, u5_mult_82_n4032, u5_mult_82_n4031,
         u5_mult_82_n4030, u5_mult_82_n4029, u5_mult_82_n4028,
         u5_mult_82_n4027, u5_mult_82_n4026, u5_mult_82_n4025,
         u5_mult_82_n4024, u5_mult_82_n4023, u5_mult_82_n4022,
         u5_mult_82_n4021, u5_mult_82_n4020, u5_mult_82_n4019,
         u5_mult_82_n4018, u5_mult_82_n4017, u5_mult_82_n4016,
         u5_mult_82_n4015, u5_mult_82_n4014, u5_mult_82_n4013,
         u5_mult_82_n4012, u5_mult_82_n4011, u5_mult_82_n4010,
         u5_mult_82_n4009, u5_mult_82_n4008, u5_mult_82_n4007,
         u5_mult_82_n4006, u5_mult_82_n4005, u5_mult_82_n4004,
         u5_mult_82_n4003, u5_mult_82_n4002, u5_mult_82_n4001,
         u5_mult_82_n4000, u5_mult_82_n3999, u5_mult_82_n3998,
         u5_mult_82_n3997, u5_mult_82_n3996, u5_mult_82_n3995,
         u5_mult_82_n3994, u5_mult_82_n3993, u5_mult_82_n3992,
         u5_mult_82_n3991, u5_mult_82_n3990, u5_mult_82_n3989,
         u5_mult_82_n3988, u5_mult_82_n3987, u5_mult_82_n3986,
         u5_mult_82_n3985, u5_mult_82_n3984, u5_mult_82_n3983,
         u5_mult_82_n3982, u5_mult_82_n3981, u5_mult_82_n3980,
         u5_mult_82_n3979, u5_mult_82_n3978, u5_mult_82_n3977,
         u5_mult_82_n3976, u5_mult_82_n3975, u5_mult_82_n3974,
         u5_mult_82_n3973, u5_mult_82_n3972, u5_mult_82_n3971,
         u5_mult_82_n3970, u5_mult_82_n3969, u5_mult_82_n3968,
         u5_mult_82_n3967, u5_mult_82_n3966, u5_mult_82_n3965,
         u5_mult_82_n3964, u5_mult_82_n3963, u5_mult_82_n3962,
         u5_mult_82_n3961, u5_mult_82_n3960, u5_mult_82_n3959,
         u5_mult_82_n3958, u5_mult_82_n3957, u5_mult_82_n3956,
         u5_mult_82_n3955, u5_mult_82_n3954, u5_mult_82_n3953,
         u5_mult_82_n3952, u5_mult_82_n3951, u5_mult_82_n3950,
         u5_mult_82_n3949, u5_mult_82_n3948, u5_mult_82_n3947,
         u5_mult_82_n3946, u5_mult_82_n3945, u5_mult_82_n3944,
         u5_mult_82_n3943, u5_mult_82_n3942, u5_mult_82_n3941,
         u5_mult_82_n3940, u5_mult_82_n3939, u5_mult_82_n3938,
         u5_mult_82_n3937, u5_mult_82_n3936, u5_mult_82_n3935,
         u5_mult_82_n3934, u5_mult_82_n3933, u5_mult_82_n3932,
         u5_mult_82_n3931, u5_mult_82_n3930, u5_mult_82_n3929,
         u5_mult_82_n3928, u5_mult_82_n3927, u5_mult_82_n3926,
         u5_mult_82_n3925, u5_mult_82_n3924, u5_mult_82_n3923,
         u5_mult_82_n3922, u5_mult_82_n3921, u5_mult_82_n3920,
         u5_mult_82_n3919, u5_mult_82_n3918, u5_mult_82_n3917,
         u5_mult_82_n3916, u5_mult_82_n3915, u5_mult_82_n3914,
         u5_mult_82_n3913, u5_mult_82_n3912, u5_mult_82_n3911,
         u5_mult_82_n3910, u5_mult_82_n3909, u5_mult_82_n3908,
         u5_mult_82_n3907, u5_mult_82_n3906, u5_mult_82_n3905,
         u5_mult_82_n3904, u5_mult_82_n3903, u5_mult_82_n3902,
         u5_mult_82_n3901, u5_mult_82_n3900, u5_mult_82_n3899,
         u5_mult_82_n3898, u5_mult_82_n3897, u5_mult_82_n3896,
         u5_mult_82_n3895, u5_mult_82_n3894, u5_mult_82_n3893,
         u5_mult_82_n3892, u5_mult_82_n3891, u5_mult_82_n3890,
         u5_mult_82_n3889, u5_mult_82_n3888, u5_mult_82_n3887,
         u5_mult_82_n3886, u5_mult_82_n3885, u5_mult_82_n3884,
         u5_mult_82_n3883, u5_mult_82_n3882, u5_mult_82_n3881,
         u5_mult_82_n3880, u5_mult_82_n3879, u5_mult_82_n3878,
         u5_mult_82_n3877, u5_mult_82_n3876, u5_mult_82_n3875,
         u5_mult_82_n3874, u5_mult_82_n3873, u5_mult_82_n3872,
         u5_mult_82_n3871, u5_mult_82_n3870, u5_mult_82_n3869,
         u5_mult_82_n3868, u5_mult_82_n3867, u5_mult_82_n3866,
         u5_mult_82_n3865, u5_mult_82_n3864, u5_mult_82_n3863,
         u5_mult_82_n3862, u5_mult_82_n3861, u5_mult_82_n3860,
         u5_mult_82_n3859, u5_mult_82_n3858, u5_mult_82_n3857,
         u5_mult_82_n3856, u5_mult_82_n3855, u5_mult_82_n3854,
         u5_mult_82_n3853, u5_mult_82_n3852, u5_mult_82_n3851,
         u5_mult_82_n3850, u5_mult_82_n3849, u5_mult_82_n3848,
         u5_mult_82_n3847, u5_mult_82_n3846, u5_mult_82_n3845,
         u5_mult_82_n3844, u5_mult_82_n3843, u5_mult_82_n3842,
         u5_mult_82_n3841, u5_mult_82_n3840, u5_mult_82_n3839,
         u5_mult_82_n3838, u5_mult_82_n3837, u5_mult_82_n3836,
         u5_mult_82_n3835, u5_mult_82_n3834, u5_mult_82_n3833,
         u5_mult_82_n3832, u5_mult_82_n3831, u5_mult_82_n3830,
         u5_mult_82_n3829, u5_mult_82_n3828, u5_mult_82_n3827,
         u5_mult_82_n3826, u5_mult_82_n3825, u5_mult_82_n3824,
         u5_mult_82_n3823, u5_mult_82_n3822, u5_mult_82_n3821,
         u5_mult_82_n3820, u5_mult_82_n3819, u5_mult_82_n3818,
         u5_mult_82_n3817, u5_mult_82_n3816, u5_mult_82_n3815,
         u5_mult_82_n3814, u5_mult_82_n3813, u5_mult_82_n3812,
         u5_mult_82_n3811, u5_mult_82_n3810, u5_mult_82_n3809,
         u5_mult_82_n3808, u5_mult_82_n3807, u5_mult_82_n3806,
         u5_mult_82_n3805, u5_mult_82_n3804, u5_mult_82_n3803,
         u5_mult_82_n3802, u5_mult_82_n3801, u5_mult_82_n3800,
         u5_mult_82_n3799, u5_mult_82_n3798, u5_mult_82_n3797,
         u5_mult_82_n3796, u5_mult_82_n3795, u5_mult_82_n3794,
         u5_mult_82_n3793, u5_mult_82_n3792, u5_mult_82_n3791,
         u5_mult_82_n3790, u5_mult_82_n3789, u5_mult_82_n3788,
         u5_mult_82_n3787, u5_mult_82_n3786, u5_mult_82_n3785,
         u5_mult_82_n3784, u5_mult_82_n3783, u5_mult_82_n3782,
         u5_mult_82_n3781, u5_mult_82_n3780, u5_mult_82_n3779,
         u5_mult_82_n3778, u5_mult_82_n3777, u5_mult_82_n3776,
         u5_mult_82_n3775, u5_mult_82_n3774, u5_mult_82_n3773,
         u5_mult_82_n3772, u5_mult_82_n3771, u5_mult_82_n3770,
         u5_mult_82_n3769, u5_mult_82_n3768, u5_mult_82_n3767,
         u5_mult_82_n3766, u5_mult_82_n3765, u5_mult_82_n3764,
         u5_mult_82_n3763, u5_mult_82_n3762, u5_mult_82_n3761,
         u5_mult_82_n3760, u5_mult_82_n3759, u5_mult_82_n3758,
         u5_mult_82_n3757, u5_mult_82_n3756, u5_mult_82_n3755,
         u5_mult_82_n3754, u5_mult_82_n3753, u5_mult_82_n3752,
         u5_mult_82_n3751, u5_mult_82_n3750, u5_mult_82_n3749,
         u5_mult_82_n3748, u5_mult_82_n3747, u5_mult_82_n3746,
         u5_mult_82_n3745, u5_mult_82_n3744, u5_mult_82_n3743,
         u5_mult_82_n3742, u5_mult_82_n3741, u5_mult_82_n3740,
         u5_mult_82_n3739, u5_mult_82_n3738, u5_mult_82_n3737,
         u5_mult_82_n3736, u5_mult_82_n3735, u5_mult_82_n3734,
         u5_mult_82_n3733, u5_mult_82_n3732, u5_mult_82_n3731,
         u5_mult_82_n3730, u5_mult_82_n3729, u5_mult_82_n3728,
         u5_mult_82_n3727, u5_mult_82_n3726, u5_mult_82_n3725,
         u5_mult_82_n3724, u5_mult_82_n3723, u5_mult_82_n3722,
         u5_mult_82_n3721, u5_mult_82_n3720, u5_mult_82_n3719,
         u5_mult_82_n3718, u5_mult_82_n3717, u5_mult_82_n3716,
         u5_mult_82_n3715, u5_mult_82_n3714, u5_mult_82_n3713,
         u5_mult_82_n3712, u5_mult_82_n3711, u5_mult_82_n3710,
         u5_mult_82_n3709, u5_mult_82_n3708, u5_mult_82_n3707,
         u5_mult_82_n3706, u5_mult_82_n3705, u5_mult_82_n3704,
         u5_mult_82_n3703, u5_mult_82_n3702, u5_mult_82_n3701,
         u5_mult_82_n3700, u5_mult_82_n3699, u5_mult_82_n3698,
         u5_mult_82_n3697, u5_mult_82_n3696, u5_mult_82_n3695,
         u5_mult_82_n3694, u5_mult_82_n3693, u5_mult_82_n3692,
         u5_mult_82_n3691, u5_mult_82_n3690, u5_mult_82_n3689,
         u5_mult_82_n3688, u5_mult_82_n3687, u5_mult_82_n3686,
         u5_mult_82_n3685, u5_mult_82_n3684, u5_mult_82_n3683,
         u5_mult_82_n3682, u5_mult_82_n3681, u5_mult_82_n3680,
         u5_mult_82_n3679, u5_mult_82_n3678, u5_mult_82_n3677,
         u5_mult_82_n3676, u5_mult_82_n3675, u5_mult_82_n3674,
         u5_mult_82_n3673, u5_mult_82_n3672, u5_mult_82_n3671,
         u5_mult_82_n3670, u5_mult_82_n3669, u5_mult_82_n3668,
         u5_mult_82_n3667, u5_mult_82_n3666, u5_mult_82_n3665,
         u5_mult_82_n3664, u5_mult_82_n3663, u5_mult_82_n3662,
         u5_mult_82_n3661, u5_mult_82_n3660, u5_mult_82_n3659,
         u5_mult_82_n3658, u5_mult_82_n3657, u5_mult_82_n3656,
         u5_mult_82_n3655, u5_mult_82_n3654, u5_mult_82_n3653,
         u5_mult_82_n3652, u5_mult_82_n3651, u5_mult_82_n3650,
         u5_mult_82_n3649, u5_mult_82_n3648, u5_mult_82_n3647,
         u5_mult_82_n3646, u5_mult_82_n3645, u5_mult_82_n3644,
         u5_mult_82_n3643, u5_mult_82_n3642, u5_mult_82_n3641,
         u5_mult_82_n3640, u5_mult_82_n3639, u5_mult_82_n3638,
         u5_mult_82_n3637, u5_mult_82_n3636, u5_mult_82_n3635,
         u5_mult_82_n3634, u5_mult_82_n3633, u5_mult_82_n3632,
         u5_mult_82_n3631, u5_mult_82_n3630, u5_mult_82_n3629,
         u5_mult_82_n3628, u5_mult_82_n3627, u5_mult_82_n3626,
         u5_mult_82_n3625, u5_mult_82_n3624, u5_mult_82_n3623,
         u5_mult_82_n3622, u5_mult_82_n3621, u5_mult_82_n3620,
         u5_mult_82_n3619, u5_mult_82_n3618, u5_mult_82_n3617,
         u5_mult_82_n3616, u5_mult_82_n3615, u5_mult_82_n3614,
         u5_mult_82_n3613, u5_mult_82_n3612, u5_mult_82_n3611,
         u5_mult_82_n3610, u5_mult_82_n3609, u5_mult_82_n3608,
         u5_mult_82_n3607, u5_mult_82_n3606, u5_mult_82_n3605,
         u5_mult_82_n3604, u5_mult_82_n3603, u5_mult_82_n3602,
         u5_mult_82_n3601, u5_mult_82_n3600, u5_mult_82_n3599,
         u5_mult_82_n3598, u5_mult_82_n3597, u5_mult_82_n3596,
         u5_mult_82_n3595, u5_mult_82_n3594, u5_mult_82_n3593,
         u5_mult_82_n3592, u5_mult_82_n3591, u5_mult_82_n3590,
         u5_mult_82_n3589, u5_mult_82_n3588, u5_mult_82_n3587,
         u5_mult_82_n3586, u5_mult_82_n3585, u5_mult_82_n3584,
         u5_mult_82_n3583, u5_mult_82_n3582, u5_mult_82_n3581,
         u5_mult_82_n3580, u5_mult_82_n3579, u5_mult_82_n3578,
         u5_mult_82_n3577, u5_mult_82_n3576, u5_mult_82_n3575,
         u5_mult_82_n3574, u5_mult_82_n3573, u5_mult_82_n3572,
         u5_mult_82_n3571, u5_mult_82_n3570, u5_mult_82_n3569,
         u5_mult_82_n3568, u5_mult_82_n3567, u5_mult_82_n3566,
         u5_mult_82_n3565, u5_mult_82_n3564, u5_mult_82_n3563,
         u5_mult_82_n3562, u5_mult_82_n3561, u5_mult_82_n3560,
         u5_mult_82_n3559, u5_mult_82_n3558, u5_mult_82_n3557,
         u5_mult_82_n3556, u5_mult_82_n3555, u5_mult_82_n3554,
         u5_mult_82_n3553, u5_mult_82_n3552, u5_mult_82_n3551,
         u5_mult_82_n3550, u5_mult_82_n3549, u5_mult_82_n3548,
         u5_mult_82_n3547, u5_mult_82_n3546, u5_mult_82_n3545,
         u5_mult_82_n3544, u5_mult_82_n3543, u5_mult_82_n3542,
         u5_mult_82_n3541, u5_mult_82_n3540, u5_mult_82_n3539,
         u5_mult_82_n3538, u5_mult_82_n3537, u5_mult_82_n3536,
         u5_mult_82_n3535, u5_mult_82_n3534, u5_mult_82_n3533,
         u5_mult_82_n3532, u5_mult_82_n3531, u5_mult_82_n3530,
         u5_mult_82_n3529, u5_mult_82_n3528, u5_mult_82_n3527,
         u5_mult_82_n3526, u5_mult_82_n3525, u5_mult_82_n3524,
         u5_mult_82_n3523, u5_mult_82_n3522, u5_mult_82_n3521,
         u5_mult_82_n3520, u5_mult_82_n3519, u5_mult_82_n3518,
         u5_mult_82_n3517, u5_mult_82_n3516, u5_mult_82_n3515,
         u5_mult_82_n3514, u5_mult_82_n3513, u5_mult_82_n3512,
         u5_mult_82_n3511, u5_mult_82_n3510, u5_mult_82_n3509,
         u5_mult_82_n3508, u5_mult_82_n3507, u5_mult_82_n3506,
         u5_mult_82_n3505, u5_mult_82_n3504, u5_mult_82_n3503,
         u5_mult_82_n3502, u5_mult_82_n3501, u5_mult_82_n3500,
         u5_mult_82_n3499, u5_mult_82_n3498, u5_mult_82_n3497,
         u5_mult_82_n3496, u5_mult_82_n3495, u5_mult_82_n3494,
         u5_mult_82_n3493, u5_mult_82_n3492, u5_mult_82_n3491,
         u5_mult_82_n3490, u5_mult_82_n3489, u5_mult_82_n3488,
         u5_mult_82_n3487, u5_mult_82_n3486, u5_mult_82_n3485,
         u5_mult_82_n3484, u5_mult_82_n3483, u5_mult_82_n3482,
         u5_mult_82_n3481, u5_mult_82_n3480, u5_mult_82_n3479,
         u5_mult_82_n3478, u5_mult_82_n3477, u5_mult_82_n3476,
         u5_mult_82_n3475, u5_mult_82_n3474, u5_mult_82_n3473,
         u5_mult_82_n3472, u5_mult_82_n3471, u5_mult_82_n3470,
         u5_mult_82_n3469, u5_mult_82_n3468, u5_mult_82_n3467,
         u5_mult_82_n3466, u5_mult_82_n3465, u5_mult_82_n3464,
         u5_mult_82_n3463, u5_mult_82_n3462, u5_mult_82_n3461,
         u5_mult_82_n3460, u5_mult_82_n3459, u5_mult_82_n3458,
         u5_mult_82_n3457, u5_mult_82_n3456, u5_mult_82_n3455,
         u5_mult_82_n3454, u5_mult_82_n3453, u5_mult_82_n3452,
         u5_mult_82_n3451, u5_mult_82_n3450, u5_mult_82_n3449,
         u5_mult_82_n3448, u5_mult_82_n3447, u5_mult_82_n3446,
         u5_mult_82_n3445, u5_mult_82_n3444, u5_mult_82_n3443,
         u5_mult_82_n3442, u5_mult_82_n3441, u5_mult_82_n3440,
         u5_mult_82_n3439, u5_mult_82_n3438, u5_mult_82_n3437,
         u5_mult_82_n3436, u5_mult_82_n3435, u5_mult_82_n3434,
         u5_mult_82_n3433, u5_mult_82_n3432, u5_mult_82_n3431,
         u5_mult_82_n3430, u5_mult_82_n3429, u5_mult_82_n3428,
         u5_mult_82_n3427, u5_mult_82_n3426, u5_mult_82_n3425,
         u5_mult_82_n3424, u5_mult_82_n3423, u5_mult_82_n3422,
         u5_mult_82_n3421, u5_mult_82_n3420, u5_mult_82_n3419,
         u5_mult_82_n3418, u5_mult_82_n3417, u5_mult_82_n3416,
         u5_mult_82_n3415, u5_mult_82_n3414, u5_mult_82_n3413,
         u5_mult_82_n3412, u5_mult_82_n3411, u5_mult_82_n3410,
         u5_mult_82_n3409, u5_mult_82_n3408, u5_mult_82_n3407,
         u5_mult_82_n3406, u5_mult_82_n3405, u5_mult_82_n3404,
         u5_mult_82_n3403, u5_mult_82_n3402, u5_mult_82_n3401,
         u5_mult_82_n3400, u5_mult_82_n3399, u5_mult_82_n3398,
         u5_mult_82_n3397, u5_mult_82_n3396, u5_mult_82_n3395,
         u5_mult_82_n3394, u5_mult_82_n3393, u5_mult_82_n3392,
         u5_mult_82_n3391, u5_mult_82_n3390, u5_mult_82_n3389,
         u5_mult_82_n3388, u5_mult_82_n3387, u5_mult_82_n3386,
         u5_mult_82_n3385, u5_mult_82_n3384, u5_mult_82_n3383,
         u5_mult_82_n3382, u5_mult_82_n3381, u5_mult_82_n3380,
         u5_mult_82_n3379, u5_mult_82_n3378, u5_mult_82_n3377,
         u5_mult_82_n3376, u5_mult_82_n3375, u5_mult_82_n3374,
         u5_mult_82_n3373, u5_mult_82_n3372, u5_mult_82_n3371,
         u5_mult_82_n3370, u5_mult_82_n3369, u5_mult_82_n3368,
         u5_mult_82_n3367, u5_mult_82_n3366, u5_mult_82_n3365,
         u5_mult_82_n3364, u5_mult_82_n3363, u5_mult_82_n3362,
         u5_mult_82_n3361, u5_mult_82_n3360, u5_mult_82_n3359,
         u5_mult_82_n3358, u5_mult_82_n3357, u5_mult_82_n3356,
         u5_mult_82_n3355, u5_mult_82_n3354, u5_mult_82_n3353,
         u5_mult_82_n3352, u5_mult_82_n3351, u5_mult_82_n3350,
         u5_mult_82_n3349, u5_mult_82_n3348, u5_mult_82_n3347,
         u5_mult_82_n3346, u5_mult_82_n3345, u5_mult_82_n3344,
         u5_mult_82_n3343, u5_mult_82_n3342, u5_mult_82_n3341,
         u5_mult_82_n3340, u5_mult_82_n3339, u5_mult_82_n3338,
         u5_mult_82_n3337, u5_mult_82_n3336, u5_mult_82_n3335,
         u5_mult_82_n3334, u5_mult_82_n3333, u5_mult_82_n3332,
         u5_mult_82_n3331, u5_mult_82_n3330, u5_mult_82_n3329,
         u5_mult_82_n3328, u5_mult_82_n3327, u5_mult_82_n3326,
         u5_mult_82_n3325, u5_mult_82_n3324, u5_mult_82_n3323,
         u5_mult_82_n3322, u5_mult_82_n3321, u5_mult_82_n3320,
         u5_mult_82_n3319, u5_mult_82_n3318, u5_mult_82_n3317,
         u5_mult_82_n3316, u5_mult_82_n3315, u5_mult_82_n3314,
         u5_mult_82_n3313, u5_mult_82_n3312, u5_mult_82_n3311,
         u5_mult_82_n3310, u5_mult_82_n3309, u5_mult_82_n3308,
         u5_mult_82_n3307, u5_mult_82_n3306, u5_mult_82_n3305,
         u5_mult_82_n3304, u5_mult_82_n3303, u5_mult_82_n3302,
         u5_mult_82_n3301, u5_mult_82_n3300, u5_mult_82_n3299,
         u5_mult_82_n3298, u5_mult_82_n3297, u5_mult_82_n3296,
         u5_mult_82_n3295, u5_mult_82_n3294, u5_mult_82_n3293,
         u5_mult_82_n3292, u5_mult_82_n3291, u5_mult_82_n3290,
         u5_mult_82_n3289, u5_mult_82_n3288, u5_mult_82_n3287,
         u5_mult_82_n3286, u5_mult_82_n3285, u5_mult_82_n3284,
         u5_mult_82_n3283, u5_mult_82_n3282, u5_mult_82_n3281,
         u5_mult_82_n3280, u5_mult_82_n3279, u5_mult_82_n3278,
         u5_mult_82_n3277, u5_mult_82_n3276, u5_mult_82_n3275,
         u5_mult_82_n3274, u5_mult_82_n3273, u5_mult_82_n3272,
         u5_mult_82_n3271, u5_mult_82_n3270, u5_mult_82_n3269,
         u5_mult_82_n3268, u5_mult_82_n3267, u5_mult_82_n3266,
         u5_mult_82_n3265, u5_mult_82_n3264, u5_mult_82_n3263,
         u5_mult_82_n3262, u5_mult_82_n3261, u5_mult_82_n3260,
         u5_mult_82_n3259, u5_mult_82_n3258, u5_mult_82_n3257,
         u5_mult_82_n3256, u5_mult_82_n3255, u5_mult_82_n3254,
         u5_mult_82_n3253, u5_mult_82_n3252, u5_mult_82_n3251,
         u5_mult_82_n3250, u5_mult_82_n3249, u5_mult_82_n3248,
         u5_mult_82_n3247, u5_mult_82_n3246, u5_mult_82_n3245,
         u5_mult_82_n3244, u5_mult_82_n3243, u5_mult_82_n3242,
         u5_mult_82_n3241, u5_mult_82_n3240, u5_mult_82_n3239,
         u5_mult_82_n3238, u5_mult_82_n3237, u5_mult_82_n3236,
         u5_mult_82_n3235, u5_mult_82_n3234, u5_mult_82_n3233,
         u5_mult_82_n3232, u5_mult_82_n3231, u5_mult_82_n3230,
         u5_mult_82_n3229, u5_mult_82_n3228, u5_mult_82_n3227,
         u5_mult_82_n3226, u5_mult_82_n3225, u5_mult_82_n3224,
         u5_mult_82_n3223, u5_mult_82_n3222, u5_mult_82_n3221,
         u5_mult_82_n3220, u5_mult_82_n3219, u5_mult_82_n3218,
         u5_mult_82_n3217, u5_mult_82_n3216, u5_mult_82_n3215,
         u5_mult_82_n3214, u5_mult_82_n3213, u5_mult_82_n3212,
         u5_mult_82_n3211, u5_mult_82_n3210, u5_mult_82_n3209,
         u5_mult_82_n3208, u5_mult_82_n3207, u5_mult_82_n3206,
         u5_mult_82_n3205, u5_mult_82_n3204, u5_mult_82_n3203,
         u5_mult_82_n3202, u5_mult_82_n3201, u5_mult_82_n3200,
         u5_mult_82_n3199, u5_mult_82_n3198, u5_mult_82_n3197,
         u5_mult_82_n3196, u5_mult_82_n3195, u5_mult_82_n3194,
         u5_mult_82_n3193, u5_mult_82_n3192, u5_mult_82_n3191,
         u5_mult_82_n3190, u5_mult_82_n3189, u5_mult_82_n3188,
         u5_mult_82_n3187, u5_mult_82_n3186, u5_mult_82_n3185,
         u5_mult_82_n3184, u5_mult_82_n3183, u5_mult_82_n3182,
         u5_mult_82_n3181, u5_mult_82_n3180, u5_mult_82_n3179,
         u5_mult_82_n3178, u5_mult_82_n3177, u5_mult_82_n3176,
         u5_mult_82_n3175, u5_mult_82_n3174, u5_mult_82_n3173,
         u5_mult_82_n3172, u5_mult_82_n3171, u5_mult_82_n3170,
         u5_mult_82_n3169, u5_mult_82_n3168, u5_mult_82_n3167,
         u5_mult_82_n3166, u5_mult_82_n3165, u5_mult_82_n3164,
         u5_mult_82_n3163, u5_mult_82_n3162, u5_mult_82_n3161,
         u5_mult_82_n3160, u5_mult_82_n3159, u5_mult_82_n3158,
         u5_mult_82_n3157, u5_mult_82_n3156, u5_mult_82_n3155,
         u5_mult_82_n3154, u5_mult_82_n3153, u5_mult_82_n3152,
         u5_mult_82_n3151, u5_mult_82_n3150, u5_mult_82_n3149,
         u5_mult_82_n3148, u5_mult_82_n3147, u5_mult_82_n3146,
         u5_mult_82_n3145, u5_mult_82_n3144, u5_mult_82_n3143,
         u5_mult_82_n3142, u5_mult_82_n3141, u5_mult_82_n3140,
         u5_mult_82_n3139, u5_mult_82_n3138, u5_mult_82_n3137,
         u5_mult_82_n3136, u5_mult_82_n3135, u5_mult_82_n3134,
         u5_mult_82_n3133, u5_mult_82_n3132, u5_mult_82_n3131,
         u5_mult_82_n3130, u5_mult_82_n3129, u5_mult_82_n3128,
         u5_mult_82_n3127, u5_mult_82_n3126, u5_mult_82_n3125,
         u5_mult_82_n3124, u5_mult_82_n3123, u5_mult_82_n3122,
         u5_mult_82_n3121, u5_mult_82_n3120, u5_mult_82_n3119,
         u5_mult_82_n3118, u5_mult_82_n3117, u5_mult_82_n3116,
         u5_mult_82_n3115, u5_mult_82_n3114, u5_mult_82_n3113,
         u5_mult_82_n3112, u5_mult_82_n3111, u5_mult_82_n3110,
         u5_mult_82_n3109, u5_mult_82_n3108, u5_mult_82_n3107,
         u5_mult_82_n3106, u5_mult_82_n3105, u5_mult_82_n3104,
         u5_mult_82_n3103, u5_mult_82_n3102, u5_mult_82_n3101,
         u5_mult_82_n3100, u5_mult_82_n3099, u5_mult_82_n3098,
         u5_mult_82_n3097, u5_mult_82_n3096, u5_mult_82_n3095,
         u5_mult_82_n3094, u5_mult_82_n3093, u5_mult_82_n3092,
         u5_mult_82_n3091, u5_mult_82_n3090, u5_mult_82_n3089,
         u5_mult_82_n3088, u5_mult_82_n3087, u5_mult_82_n3086,
         u5_mult_82_n3085, u5_mult_82_n3084, u5_mult_82_n3083,
         u5_mult_82_n3082, u5_mult_82_n3081, u5_mult_82_n3080,
         u5_mult_82_n3079, u5_mult_82_n3078, u5_mult_82_n3077,
         u5_mult_82_n3076, u5_mult_82_n3075, u5_mult_82_n3074,
         u5_mult_82_n3073, u5_mult_82_n3072, u5_mult_82_n3071,
         u5_mult_82_n3070, u5_mult_82_n3069, u5_mult_82_n3068,
         u5_mult_82_n3067, u5_mult_82_n3066, u5_mult_82_n3065,
         u5_mult_82_n3064, u5_mult_82_n3063, u5_mult_82_n3062,
         u5_mult_82_n3061, u5_mult_82_n3060, u5_mult_82_n3059,
         u5_mult_82_n3058, u5_mult_82_n3057, u5_mult_82_n3056,
         u5_mult_82_n3055, u5_mult_82_n3054, u5_mult_82_n3053,
         u5_mult_82_n3052, u5_mult_82_n3051, u5_mult_82_n3050,
         u5_mult_82_n3049, u5_mult_82_n3048, u5_mult_82_n3047,
         u5_mult_82_n3046, u5_mult_82_n3045, u5_mult_82_n3044,
         u5_mult_82_n3043, u5_mult_82_n3042, u5_mult_82_n3041,
         u5_mult_82_n3040, u5_mult_82_n3039, u5_mult_82_n3038,
         u5_mult_82_n3037, u5_mult_82_n3036, u5_mult_82_n3035,
         u5_mult_82_n3034, u5_mult_82_n3033, u5_mult_82_n3032,
         u5_mult_82_n3031, u5_mult_82_n3030, u5_mult_82_n3029,
         u5_mult_82_n3028, u5_mult_82_n3027, u5_mult_82_n3026,
         u5_mult_82_n3025, u5_mult_82_n3024, u5_mult_82_n3023,
         u5_mult_82_n3022, u5_mult_82_n3021, u5_mult_82_n3020,
         u5_mult_82_n3019, u5_mult_82_n3018, u5_mult_82_n3017,
         u5_mult_82_n3016, u5_mult_82_n3015, u5_mult_82_n3014,
         u5_mult_82_n3013, u5_mult_82_n3012, u5_mult_82_n3011,
         u5_mult_82_n3010, u5_mult_82_n3009, u5_mult_82_n3008,
         u5_mult_82_n3007, u5_mult_82_n3006, u5_mult_82_n3005,
         u5_mult_82_n3004, u5_mult_82_n3003, u5_mult_82_n3002,
         u5_mult_82_n3001, u5_mult_82_n3000, u5_mult_82_n2999,
         u5_mult_82_n2998, u5_mult_82_n2997, u5_mult_82_n2996,
         u5_mult_82_n2995, u5_mult_82_n2994, u5_mult_82_n2993,
         u5_mult_82_n2992, u5_mult_82_n2991, u5_mult_82_n2990,
         u5_mult_82_n2989, u5_mult_82_n2988, u5_mult_82_n2987,
         u5_mult_82_n2986, u5_mult_82_n2985, u5_mult_82_n2984,
         u5_mult_82_n2983, u5_mult_82_n2982, u5_mult_82_n2981,
         u5_mult_82_n2980, u5_mult_82_n2979, u5_mult_82_n2978,
         u5_mult_82_n2977, u5_mult_82_n2976, u5_mult_82_n2975,
         u5_mult_82_n2974, u5_mult_82_n2973, u5_mult_82_n2972,
         u5_mult_82_n2971, u5_mult_82_n2970, u5_mult_82_n2969,
         u5_mult_82_n2968, u5_mult_82_n2967, u5_mult_82_n2966,
         u5_mult_82_n2965, u5_mult_82_n2964, u5_mult_82_n2963,
         u5_mult_82_n2962, u5_mult_82_n2961, u5_mult_82_n2960,
         u5_mult_82_n2959, u5_mult_82_n2958, u5_mult_82_n2957,
         u5_mult_82_n2956, u5_mult_82_n2955, u5_mult_82_n2954,
         u5_mult_82_n2953, u5_mult_82_n2952, u5_mult_82_n2951,
         u5_mult_82_n2950, u5_mult_82_n2949, u5_mult_82_n2948,
         u5_mult_82_n2947, u5_mult_82_n2946, u5_mult_82_n2945,
         u5_mult_82_n2944, u5_mult_82_n2943, u5_mult_82_n2942,
         u5_mult_82_n2941, u5_mult_82_n2940, u5_mult_82_n2939,
         u5_mult_82_n2938, u5_mult_82_n2937, u5_mult_82_n2936,
         u5_mult_82_n2935, u5_mult_82_n2934, u5_mult_82_n2933,
         u5_mult_82_n2932, u5_mult_82_n2931, u5_mult_82_n2930,
         u5_mult_82_n2929, u5_mult_82_n2928, u5_mult_82_n2927,
         u5_mult_82_n2926, u5_mult_82_n2925, u5_mult_82_n2924,
         u5_mult_82_n2923, u5_mult_82_n2922, u5_mult_82_n2921,
         u5_mult_82_n2920, u5_mult_82_n2919, u5_mult_82_n2918,
         u5_mult_82_n2917, u5_mult_82_n2916, u5_mult_82_n2915,
         u5_mult_82_n2914, u5_mult_82_n2913, u5_mult_82_n2912,
         u5_mult_82_n2911, u5_mult_82_n2910, u5_mult_82_n2909,
         u5_mult_82_n2908, u5_mult_82_n2907, u5_mult_82_n2906,
         u5_mult_82_n2905, u5_mult_82_n2904, u5_mult_82_n2903,
         u5_mult_82_n2902, u5_mult_82_n2901, u5_mult_82_n2900,
         u5_mult_82_n2899, u5_mult_82_n2898, u5_mult_82_n2897,
         u5_mult_82_n2896, u5_mult_82_n2895, u5_mult_82_n2894,
         u5_mult_82_n2893, u5_mult_82_n2892, u5_mult_82_n2891,
         u5_mult_82_n2890, u5_mult_82_n2889, u5_mult_82_n2888,
         u5_mult_82_n2887, u5_mult_82_n2886, u5_mult_82_n2885,
         u5_mult_82_n2884, u5_mult_82_n2883, u5_mult_82_n2882,
         u5_mult_82_n2881, u5_mult_82_n2880, u5_mult_82_n2879,
         u5_mult_82_n2878, u5_mult_82_n2877, u5_mult_82_n2876,
         u5_mult_82_n2875, u5_mult_82_n2874, u5_mult_82_n2873,
         u5_mult_82_n2872, u5_mult_82_n2871, u5_mult_82_n2870,
         u5_mult_82_n2869, u5_mult_82_n2868, u5_mult_82_n2867,
         u5_mult_82_n2866, u5_mult_82_n2865, u5_mult_82_n2864,
         u5_mult_82_n2863, u5_mult_82_n2862, u5_mult_82_n2861,
         u5_mult_82_n2860, u5_mult_82_n2859, u5_mult_82_n2858,
         u5_mult_82_n2857, u5_mult_82_n2856, u5_mult_82_n2855,
         u5_mult_82_n2854, u5_mult_82_n2853, u5_mult_82_n2852,
         u5_mult_82_n2851, u5_mult_82_n2850, u5_mult_82_n2849,
         u5_mult_82_n2848, u5_mult_82_n2847, u5_mult_82_n2846,
         u5_mult_82_n2845, u5_mult_82_n2844, u5_mult_82_n2843,
         u5_mult_82_n2842, u5_mult_82_n2841, u5_mult_82_n2840,
         u5_mult_82_n2839, u5_mult_82_n2838, u5_mult_82_n2837,
         u5_mult_82_n2836, u5_mult_82_n2835, u5_mult_82_n2834,
         u5_mult_82_n2833, u5_mult_82_n2832, u5_mult_82_n2831,
         u5_mult_82_n2830, u5_mult_82_n2829, u5_mult_82_n2828,
         u5_mult_82_n2827, u5_mult_82_n2826, u5_mult_82_n2825,
         u5_mult_82_n2824, u5_mult_82_n2823, u5_mult_82_n2822,
         u5_mult_82_n2821, u5_mult_82_n2820, u5_mult_82_n2819,
         u5_mult_82_n2818, u5_mult_82_n2817, u5_mult_82_n2816,
         u5_mult_82_n2815, u5_mult_82_n2814, u5_mult_82_n2813,
         u5_mult_82_n2812, u5_mult_82_n2811, u5_mult_82_n2810,
         u5_mult_82_n2809, u5_mult_82_n2808, u5_mult_82_n2807,
         u5_mult_82_n2806, u5_mult_82_n2805, u5_mult_82_n2804,
         u5_mult_82_n2803, u5_mult_82_n2802, u5_mult_82_n2801,
         u5_mult_82_n2800, u5_mult_82_n2799, u5_mult_82_n2798,
         u5_mult_82_n2797, u5_mult_82_n2796, u5_mult_82_n2795,
         u5_mult_82_n2794, u5_mult_82_n2793, u5_mult_82_n2792,
         u5_mult_82_n2791, u5_mult_82_n2790, u5_mult_82_n2789,
         u5_mult_82_n2788, u5_mult_82_n2787, u5_mult_82_n2786,
         u5_mult_82_n2785, u5_mult_82_n2784, u5_mult_82_n2783,
         u5_mult_82_n2782, u5_mult_82_n2781, u5_mult_82_n2780,
         u5_mult_82_n2779, u5_mult_82_n2778, u5_mult_82_n2777,
         u5_mult_82_n2776, u5_mult_82_n2775, u5_mult_82_n2774,
         u5_mult_82_n2773, u5_mult_82_n2772, u5_mult_82_n2771,
         u5_mult_82_n2770, u5_mult_82_n2769, u5_mult_82_n2768,
         u5_mult_82_n2767, u5_mult_82_n2766, u5_mult_82_n2765,
         u5_mult_82_n2764, u5_mult_82_n2763, u5_mult_82_n2762,
         u5_mult_82_n2761, u5_mult_82_n2760, u5_mult_82_n2759,
         u5_mult_82_n2758, u5_mult_82_n2757, u5_mult_82_n2756,
         u5_mult_82_n2755, u5_mult_82_n2754, u5_mult_82_n2753,
         u5_mult_82_n2752, u5_mult_82_n2751, u5_mult_82_n2750,
         u5_mult_82_n2749, u5_mult_82_n2748, u5_mult_82_n2747,
         u5_mult_82_n2746, u5_mult_82_n2745, u5_mult_82_n2744,
         u5_mult_82_n2743, u5_mult_82_n2742, u5_mult_82_n2741,
         u5_mult_82_n2740, u5_mult_82_n2739, u5_mult_82_n2738,
         u5_mult_82_n2737, u5_mult_82_n2736, u5_mult_82_n2735,
         u5_mult_82_n2734, u5_mult_82_n2733, u5_mult_82_n2732,
         u5_mult_82_n2731, u5_mult_82_n2730, u5_mult_82_n2729,
         u5_mult_82_n2728, u5_mult_82_n2727, u5_mult_82_n2726,
         u5_mult_82_n2725, u5_mult_82_n2724, u5_mult_82_n2723,
         u5_mult_82_n2722, u5_mult_82_n2721, u5_mult_82_n2720,
         u5_mult_82_n2719, u5_mult_82_n2718, u5_mult_82_n2717,
         u5_mult_82_n2716, u5_mult_82_n2715, u5_mult_82_n2714,
         u5_mult_82_n2713, u5_mult_82_n2712, u5_mult_82_n2711,
         u5_mult_82_n2710, u5_mult_82_n2709, u5_mult_82_n2708,
         u5_mult_82_n2707, u5_mult_82_n2706, u5_mult_82_n2705,
         u5_mult_82_n2704, u5_mult_82_n2703, u5_mult_82_n2702,
         u5_mult_82_n2701, u5_mult_82_n2700, u5_mult_82_n2699,
         u5_mult_82_n2698, u5_mult_82_n2697, u5_mult_82_n2696,
         u5_mult_82_n2695, u5_mult_82_n2694, u5_mult_82_n2693,
         u5_mult_82_n2692, u5_mult_82_n2691, u5_mult_82_n2690,
         u5_mult_82_n2689, u5_mult_82_n2688, u5_mult_82_n2687,
         u5_mult_82_n2686, u5_mult_82_n2685, u5_mult_82_n2684,
         u5_mult_82_n2683, u5_mult_82_n2682, u5_mult_82_n2681,
         u5_mult_82_n2680, u5_mult_82_n2679, u5_mult_82_n2678,
         u5_mult_82_n2677, u5_mult_82_n2676, u5_mult_82_n2675,
         u5_mult_82_n2674, u5_mult_82_n2673, u5_mult_82_n2672,
         u5_mult_82_n2671, u5_mult_82_n2670, u5_mult_82_n2669,
         u5_mult_82_n2668, u5_mult_82_n2667, u5_mult_82_n2666,
         u5_mult_82_n2665, u5_mult_82_n2664, u5_mult_82_n2663,
         u5_mult_82_n2662, u5_mult_82_n2661, u5_mult_82_n2660,
         u5_mult_82_n2659, u5_mult_82_n2658, u5_mult_82_n2657,
         u5_mult_82_n2656, u5_mult_82_n2655, u5_mult_82_n2654,
         u5_mult_82_n2653, u5_mult_82_n2652, u5_mult_82_n2651,
         u5_mult_82_n2650, u5_mult_82_n2649, u5_mult_82_n2648,
         u5_mult_82_n2647, u5_mult_82_n2646, u5_mult_82_n2645,
         u5_mult_82_n2644, u5_mult_82_n2643, u5_mult_82_n2642,
         u5_mult_82_n2641, u5_mult_82_n2640, u5_mult_82_n2639,
         u5_mult_82_n2638, u5_mult_82_n2637, u5_mult_82_n2636,
         u5_mult_82_n2635, u5_mult_82_n2634, u5_mult_82_n2633,
         u5_mult_82_n2632, u5_mult_82_n2631, u5_mult_82_n2630,
         u5_mult_82_n2629, u5_mult_82_n2628, u5_mult_82_n2627,
         u5_mult_82_n2626, u5_mult_82_n2625, u5_mult_82_n2624,
         u5_mult_82_n2623, u5_mult_82_n2622, u5_mult_82_n2621,
         u5_mult_82_n2620, u5_mult_82_n2619, u5_mult_82_n2618,
         u5_mult_82_n2617, u5_mult_82_n2616, u5_mult_82_n2615,
         u5_mult_82_n2614, u5_mult_82_n2613, u5_mult_82_n2612,
         u5_mult_82_n2611, u5_mult_82_n2610, u5_mult_82_n2609,
         u5_mult_82_n2608, u5_mult_82_n2607, u5_mult_82_n2606,
         u5_mult_82_n2605, u5_mult_82_n2604, u5_mult_82_n2603,
         u5_mult_82_n2602, u5_mult_82_n2601, u5_mult_82_n2600,
         u5_mult_82_n2599, u5_mult_82_n2598, u5_mult_82_n2597,
         u5_mult_82_n2596, u5_mult_82_n2595, u5_mult_82_n2594,
         u5_mult_82_n2593, u5_mult_82_n2592, u5_mult_82_n2591,
         u5_mult_82_n2590, u5_mult_82_n2589, u5_mult_82_n2588,
         u5_mult_82_n2587, u5_mult_82_n2586, u5_mult_82_n2585,
         u5_mult_82_n2584, u5_mult_82_n2583, u5_mult_82_n2582,
         u5_mult_82_n2581, u5_mult_82_n2580, u5_mult_82_n2579,
         u5_mult_82_n2578, u5_mult_82_n2577, u5_mult_82_n2576,
         u5_mult_82_n2575, u5_mult_82_n2574, u5_mult_82_n2573,
         u5_mult_82_n2572, u5_mult_82_n2571, u5_mult_82_n2570,
         u5_mult_82_n2569, u5_mult_82_n2568, u5_mult_82_n2567,
         u5_mult_82_n2566, u5_mult_82_n2565, u5_mult_82_n2564,
         u5_mult_82_n2563, u5_mult_82_n2562, u5_mult_82_n2561,
         u5_mult_82_n2560, u5_mult_82_n2559, u5_mult_82_n2558,
         u5_mult_82_n2557, u5_mult_82_n2556, u5_mult_82_n2555,
         u5_mult_82_n2554, u5_mult_82_n2553, u5_mult_82_n2552,
         u5_mult_82_n2551, u5_mult_82_n2550, u5_mult_82_n2549,
         u5_mult_82_n2548, u5_mult_82_n2547, u5_mult_82_n2546,
         u5_mult_82_n2545, u5_mult_82_n2544, u5_mult_82_n2543,
         u5_mult_82_n2542, u5_mult_82_n2541, u5_mult_82_n2540,
         u5_mult_82_n2539, u5_mult_82_n2538, u5_mult_82_n2537,
         u5_mult_82_n2536, u5_mult_82_n2535, u5_mult_82_n2534,
         u5_mult_82_n2533, u5_mult_82_n2532, u5_mult_82_n2531,
         u5_mult_82_n2530, u5_mult_82_n2529, u5_mult_82_n2528,
         u5_mult_82_n2527, u5_mult_82_n2526, u5_mult_82_n2525,
         u5_mult_82_n2524, u5_mult_82_n2523, u5_mult_82_n2522,
         u5_mult_82_n2521, u5_mult_82_n2520, u5_mult_82_n2519,
         u5_mult_82_n2518, u5_mult_82_n2517, u5_mult_82_n2516,
         u5_mult_82_n2515, u5_mult_82_n2514, u5_mult_82_n2513,
         u5_mult_82_n2512, u5_mult_82_n2511, u5_mult_82_n2510,
         u5_mult_82_n2509, u5_mult_82_n2508, u5_mult_82_n2507,
         u5_mult_82_n2506, u5_mult_82_n2505, u5_mult_82_n2504,
         u5_mult_82_n2503, u5_mult_82_n2502, u5_mult_82_n2501,
         u5_mult_82_n2500, u5_mult_82_n2499, u5_mult_82_n2498,
         u5_mult_82_n2497, u5_mult_82_n2496, u5_mult_82_n2495,
         u5_mult_82_n2494, u5_mult_82_n2493, u5_mult_82_n2492,
         u5_mult_82_n2491, u5_mult_82_n2490, u5_mult_82_n2489,
         u5_mult_82_n2488, u5_mult_82_n2487, u5_mult_82_n2486,
         u5_mult_82_n2485, u5_mult_82_n2484, u5_mult_82_n2483,
         u5_mult_82_n2482, u5_mult_82_n2481, u5_mult_82_n2480,
         u5_mult_82_n2479, u5_mult_82_n2478, u5_mult_82_n2477,
         u5_mult_82_n2476, u5_mult_82_n2475, u5_mult_82_n2474,
         u5_mult_82_n2473, u5_mult_82_n2472, u5_mult_82_n2471,
         u5_mult_82_n2470, u5_mult_82_n2469, u5_mult_82_n2468,
         u5_mult_82_n2467, u5_mult_82_n2466, u5_mult_82_n2465,
         u5_mult_82_n2464, u5_mult_82_n2463, u5_mult_82_n2462,
         u5_mult_82_n2461, u5_mult_82_n2460, u5_mult_82_n2459,
         u5_mult_82_n2458, u5_mult_82_n2457, u5_mult_82_n2456,
         u5_mult_82_n2455, u5_mult_82_n2454, u5_mult_82_n2453,
         u5_mult_82_n2452, u5_mult_82_n2451, u5_mult_82_n2450,
         u5_mult_82_n2449, u5_mult_82_n2448, u5_mult_82_n2447,
         u5_mult_82_n2446, u5_mult_82_n2445, u5_mult_82_n2444,
         u5_mult_82_n2443, u5_mult_82_n2442, u5_mult_82_n2441,
         u5_mult_82_n2440, u5_mult_82_n2439, u5_mult_82_n2438,
         u5_mult_82_n2437, u5_mult_82_n2436, u5_mult_82_n2435,
         u5_mult_82_n2434, u5_mult_82_n2433, u5_mult_82_n2432,
         u5_mult_82_n2431, u5_mult_82_n2430, u5_mult_82_n2429,
         u5_mult_82_n2428, u5_mult_82_n2427, u5_mult_82_n2426,
         u5_mult_82_n2425, u5_mult_82_n2424, u5_mult_82_n2423,
         u5_mult_82_n2422, u5_mult_82_n2421, u5_mult_82_n2420,
         u5_mult_82_n2419, u5_mult_82_n2418, u5_mult_82_n2417,
         u5_mult_82_n2416, u5_mult_82_n2415, u5_mult_82_n2414,
         u5_mult_82_n2413, u5_mult_82_n2412, u5_mult_82_n2411,
         u5_mult_82_n2410, u5_mult_82_n2409, u5_mult_82_n2408,
         u5_mult_82_n2407, u5_mult_82_n2406, u5_mult_82_n2405,
         u5_mult_82_n2404, u5_mult_82_n2403, u5_mult_82_n2402,
         u5_mult_82_n2401, u5_mult_82_n2400, u5_mult_82_n2399,
         u5_mult_82_n2398, u5_mult_82_n2397, u5_mult_82_n2396,
         u5_mult_82_n2395, u5_mult_82_n2394, u5_mult_82_n2393,
         u5_mult_82_n2392, u5_mult_82_n2391, u5_mult_82_n2390,
         u5_mult_82_n2389, u5_mult_82_n2388, u5_mult_82_n2387,
         u5_mult_82_n2386, u5_mult_82_n2385, u5_mult_82_n2384,
         u5_mult_82_n2383, u5_mult_82_n2382, u5_mult_82_n2381,
         u5_mult_82_n2380, u5_mult_82_n2379, u5_mult_82_n2378,
         u5_mult_82_n2377, u5_mult_82_n2376, u5_mult_82_n2375,
         u5_mult_82_n2374, u5_mult_82_n2373, u5_mult_82_n2372,
         u5_mult_82_n2371, u5_mult_82_n2370, u5_mult_82_n2369,
         u5_mult_82_n2368, u5_mult_82_n2367, u5_mult_82_n2366,
         u5_mult_82_n2365, u5_mult_82_n2364, u5_mult_82_n2363,
         u5_mult_82_n2362, u5_mult_82_n2361, u5_mult_82_n2360,
         u5_mult_82_n2359, u5_mult_82_n2358, u5_mult_82_n2357,
         u5_mult_82_n2356, u5_mult_82_n2355, u5_mult_82_n2354,
         u5_mult_82_n2353, u5_mult_82_n2352, u5_mult_82_n2351,
         u5_mult_82_n2350, u5_mult_82_n2349, u5_mult_82_n2348,
         u5_mult_82_n2347, u5_mult_82_n2346, u5_mult_82_n2345,
         u5_mult_82_n2344, u5_mult_82_n2343, u5_mult_82_n2342,
         u5_mult_82_n2341, u5_mult_82_n2340, u5_mult_82_n2339,
         u5_mult_82_n2338, u5_mult_82_n2337, u5_mult_82_n2336,
         u5_mult_82_n2335, u5_mult_82_n2334, u5_mult_82_n2333,
         u5_mult_82_n2332, u5_mult_82_n2331, u5_mult_82_n2330,
         u5_mult_82_n2329, u5_mult_82_n2328, u5_mult_82_n2327,
         u5_mult_82_n2326, u5_mult_82_n2325, u5_mult_82_n2324,
         u5_mult_82_n2323, u5_mult_82_n2322, u5_mult_82_n2321,
         u5_mult_82_n2320, u5_mult_82_n2319, u5_mult_82_n2318,
         u5_mult_82_n2317, u5_mult_82_n2316, u5_mult_82_n2315,
         u5_mult_82_n2314, u5_mult_82_n2313, u5_mult_82_n2312,
         u5_mult_82_n2311, u5_mult_82_n2310, u5_mult_82_n2309,
         u5_mult_82_n2308, u5_mult_82_n2307, u5_mult_82_n2306,
         u5_mult_82_n2305, u5_mult_82_n2304, u5_mult_82_n2303,
         u5_mult_82_n2302, u5_mult_82_n2301, u5_mult_82_n2300,
         u5_mult_82_n2299, u5_mult_82_n2298, u5_mult_82_n2297,
         u5_mult_82_n2296, u5_mult_82_n2295, u5_mult_82_n2294,
         u5_mult_82_n2293, u5_mult_82_n2292, u5_mult_82_n2291,
         u5_mult_82_n2290, u5_mult_82_n2289, u5_mult_82_n2288,
         u5_mult_82_n2287, u5_mult_82_n2286, u5_mult_82_n2285,
         u5_mult_82_n2284, u5_mult_82_n2283, u5_mult_82_n2282,
         u5_mult_82_n2281, u5_mult_82_n2280, u5_mult_82_n2279,
         u5_mult_82_n2278, u5_mult_82_n2277, u5_mult_82_n2276,
         u5_mult_82_n2275, u5_mult_82_n2274, u5_mult_82_n2273,
         u5_mult_82_n2272, u5_mult_82_n2271, u5_mult_82_n2270,
         u5_mult_82_n2269, u5_mult_82_n2268, u5_mult_82_n2267,
         u5_mult_82_n2266, u5_mult_82_n2265, u5_mult_82_n2264,
         u5_mult_82_n2263, u5_mult_82_n2262, u5_mult_82_n2261,
         u5_mult_82_n2260, u5_mult_82_n2259, u5_mult_82_n2258,
         u5_mult_82_n2257, u5_mult_82_n2256, u5_mult_82_n2255,
         u5_mult_82_n2254, u5_mult_82_n2253, u5_mult_82_n2252,
         u5_mult_82_n2251, u5_mult_82_n2250, u5_mult_82_n2249,
         u5_mult_82_n2248, u5_mult_82_n2247, u5_mult_82_n2246,
         u5_mult_82_n2245, u5_mult_82_n2244, u5_mult_82_n2243,
         u5_mult_82_n2242, u5_mult_82_n2241, u5_mult_82_n2240,
         u5_mult_82_n2239, u5_mult_82_n2238, u5_mult_82_n2237,
         u5_mult_82_n2236, u5_mult_82_n2235, u5_mult_82_n2234,
         u5_mult_82_n2233, u5_mult_82_n2232, u5_mult_82_n2231,
         u5_mult_82_n2230, u5_mult_82_n2229, u5_mult_82_n2228,
         u5_mult_82_n2227, u5_mult_82_n2226, u5_mult_82_n2225,
         u5_mult_82_n2224, u5_mult_82_n2223, u5_mult_82_n2222,
         u5_mult_82_n2221, u5_mult_82_n2220, u5_mult_82_n2219,
         u5_mult_82_n2218, u5_mult_82_n2217, u5_mult_82_n2216,
         u5_mult_82_n2215, u5_mult_82_n2214, u5_mult_82_n2213,
         u5_mult_82_n2212, u5_mult_82_n2211, u5_mult_82_n2210,
         u5_mult_82_n2209, u5_mult_82_n2208, u5_mult_82_n2207,
         u5_mult_82_n2206, u5_mult_82_n2205, u5_mult_82_n2204,
         u5_mult_82_n2203, u5_mult_82_n2202, u5_mult_82_n2201,
         u5_mult_82_n2200, u5_mult_82_n2199, u5_mult_82_n2198,
         u5_mult_82_n2197, u5_mult_82_n2196, u5_mult_82_n2195,
         u5_mult_82_n2194, u5_mult_82_n2193, u5_mult_82_n2192,
         u5_mult_82_n2191, u5_mult_82_n2190, u5_mult_82_n2189,
         u5_mult_82_n2188, u5_mult_82_n2187, u5_mult_82_n2186,
         u5_mult_82_n2185, u5_mult_82_n2184, u5_mult_82_n2183,
         u5_mult_82_n2182, u5_mult_82_n2181, u5_mult_82_n2180,
         u5_mult_82_n2179, u5_mult_82_n2178, u5_mult_82_n2177,
         u5_mult_82_n2176, u5_mult_82_n2175, u5_mult_82_n2174,
         u5_mult_82_n2173, u5_mult_82_n2172, u5_mult_82_n2171,
         u5_mult_82_n2170, u5_mult_82_n2169, u5_mult_82_n2168,
         u5_mult_82_n2167, u5_mult_82_n2166, u5_mult_82_n2165,
         u5_mult_82_n2164, u5_mult_82_n2163, u5_mult_82_n2162,
         u5_mult_82_n2161, u5_mult_82_n2160, u5_mult_82_n2159,
         u5_mult_82_n2158, u5_mult_82_n2157, u5_mult_82_n2156,
         u5_mult_82_n2155, u5_mult_82_n2154, u5_mult_82_n2153,
         u5_mult_82_n2152, u5_mult_82_n2151, u5_mult_82_n2150,
         u5_mult_82_n2149, u5_mult_82_n2148, u5_mult_82_n2147,
         u5_mult_82_n2146, u5_mult_82_n2145, u5_mult_82_n2144,
         u5_mult_82_n2143, u5_mult_82_n2142, u5_mult_82_n2141,
         u5_mult_82_n2140, u5_mult_82_n2139, u5_mult_82_n2138,
         u5_mult_82_n2137, u5_mult_82_n2136, u5_mult_82_n2135,
         u5_mult_82_n2134, u5_mult_82_n2133, u5_mult_82_n2132,
         u5_mult_82_n2131, u5_mult_82_n2130, u5_mult_82_n2129,
         u5_mult_82_n2128, u5_mult_82_n2127, u5_mult_82_n2126,
         u5_mult_82_n2125, u5_mult_82_n2124, u5_mult_82_n2123,
         u5_mult_82_n2122, u5_mult_82_n2121, u5_mult_82_n2120,
         u5_mult_82_n2119, u5_mult_82_n2118, u5_mult_82_n2117,
         u5_mult_82_n2116, u5_mult_82_n2115, u5_mult_82_n2114,
         u5_mult_82_n2113, u5_mult_82_n2112, u5_mult_82_n2111,
         u5_mult_82_n2110, u5_mult_82_n2109, u5_mult_82_n2108,
         u5_mult_82_n2107, u5_mult_82_n2106, u5_mult_82_n2105,
         u5_mult_82_n2104, u5_mult_82_n2103, u5_mult_82_n2102,
         u5_mult_82_n2101, u5_mult_82_n2100, u5_mult_82_n2099,
         u5_mult_82_n2098, u5_mult_82_n2097, u5_mult_82_n2096,
         u5_mult_82_n2095, u5_mult_82_n2094, u5_mult_82_n2093,
         u5_mult_82_n2092, u5_mult_82_n2091, u5_mult_82_n2090,
         u5_mult_82_n2089, u5_mult_82_n2088, u5_mult_82_n2087,
         u5_mult_82_n2086, u5_mult_82_n2085, u5_mult_82_n2084,
         u5_mult_82_n2083, u5_mult_82_n2082, u5_mult_82_n2081,
         u5_mult_82_n2080, u5_mult_82_n2079, u5_mult_82_n2078,
         u5_mult_82_n2077, u5_mult_82_n2076, u5_mult_82_n2075,
         u5_mult_82_n2074, u5_mult_82_n2073, u5_mult_82_n2072,
         u5_mult_82_n2071, u5_mult_82_n2070, u5_mult_82_n2069,
         u5_mult_82_n2068, u5_mult_82_n2067, u5_mult_82_n2066,
         u5_mult_82_n2065, u5_mult_82_n2064, u5_mult_82_n2063,
         u5_mult_82_n2062, u5_mult_82_n2061, u5_mult_82_n2060,
         u5_mult_82_n2059, u5_mult_82_n2058, u5_mult_82_n2057,
         u5_mult_82_n2056, u5_mult_82_n2055, u5_mult_82_n2054,
         u5_mult_82_n2053, u5_mult_82_n2052, u5_mult_82_n2051,
         u5_mult_82_n2050, u5_mult_82_n2049, u5_mult_82_n2048,
         u5_mult_82_n2047, u5_mult_82_n2046, u5_mult_82_n2045,
         u5_mult_82_n2044, u5_mult_82_n2043, u5_mult_82_n2042,
         u5_mult_82_n2041, u5_mult_82_n2040, u5_mult_82_n2039,
         u5_mult_82_n2038, u5_mult_82_n2037, u5_mult_82_n2036,
         u5_mult_82_n2035, u5_mult_82_n2034, u5_mult_82_n2033,
         u5_mult_82_n2032, u5_mult_82_n2031, u5_mult_82_n2030,
         u5_mult_82_n2029, u5_mult_82_n2028, u5_mult_82_n2027,
         u5_mult_82_n2026, u5_mult_82_n2025, u5_mult_82_n2024,
         u5_mult_82_n2023, u5_mult_82_n2022, u5_mult_82_n2021,
         u5_mult_82_n2020, u5_mult_82_n2019, u5_mult_82_n2018,
         u5_mult_82_n2017, u5_mult_82_n2016, u5_mult_82_n2015,
         u5_mult_82_n2014, u5_mult_82_n2013, u5_mult_82_n2012,
         u5_mult_82_n2011, u5_mult_82_n2010, u5_mult_82_n2009,
         u5_mult_82_n2008, u5_mult_82_n2007, u5_mult_82_n2006,
         u5_mult_82_n2005, u5_mult_82_n2004, u5_mult_82_n2003,
         u5_mult_82_n2002, u5_mult_82_n2001, u5_mult_82_n2000,
         u5_mult_82_n1999, u5_mult_82_n1998, u5_mult_82_n1997,
         u5_mult_82_n1996, u5_mult_82_n1995, u5_mult_82_n1994,
         u5_mult_82_n1993, u5_mult_82_n1992, u5_mult_82_n1991,
         u5_mult_82_n1990, u5_mult_82_n1989, u5_mult_82_n1988,
         u5_mult_82_n1987, u5_mult_82_n1986, u5_mult_82_n1985,
         u5_mult_82_n1984, u5_mult_82_n1983, u5_mult_82_n1982,
         u5_mult_82_n1981, u5_mult_82_n1980, u5_mult_82_n1979,
         u5_mult_82_n1978, u5_mult_82_n1977, u5_mult_82_n1976,
         u5_mult_82_n1975, u5_mult_82_n1974, u5_mult_82_n1973,
         u5_mult_82_n1972, u5_mult_82_n1971, u5_mult_82_n1970,
         u5_mult_82_n1969, u5_mult_82_n1968, u5_mult_82_n1967,
         u5_mult_82_n1966, u5_mult_82_n1965, u5_mult_82_n1964,
         u5_mult_82_n1963, u5_mult_82_n1962, u5_mult_82_n1961,
         u5_mult_82_n1960, u5_mult_82_n1959, u5_mult_82_n1958,
         u5_mult_82_n1957, u5_mult_82_n1956, u5_mult_82_n1955,
         u5_mult_82_n1954, u5_mult_82_n1953, u5_mult_82_n1952,
         u5_mult_82_n1951, u5_mult_82_n1950, u5_mult_82_n1949,
         u5_mult_82_n1948, u5_mult_82_n1947, u5_mult_82_n1946,
         u5_mult_82_n1945, u5_mult_82_n1944, u5_mult_82_n1943,
         u5_mult_82_n1942, u5_mult_82_n1941, u5_mult_82_n1940,
         u5_mult_82_n1939, u5_mult_82_n1938, u5_mult_82_n1937,
         u5_mult_82_n1936, u5_mult_82_n1935, u5_mult_82_n1934,
         u5_mult_82_n1933, u5_mult_82_n1932, u5_mult_82_n1931,
         u5_mult_82_n1930, u5_mult_82_n1929, u5_mult_82_n1928,
         u5_mult_82_n1927, u5_mult_82_n1926, u5_mult_82_n1925,
         u5_mult_82_n1924, u5_mult_82_n1923, u5_mult_82_n1922,
         u5_mult_82_n1921, u5_mult_82_n1920, u5_mult_82_n1919,
         u5_mult_82_n1918, u5_mult_82_n1917, u5_mult_82_n1916,
         u5_mult_82_n1915, u5_mult_82_n1914, u5_mult_82_n1913,
         u5_mult_82_n1912, u5_mult_82_n1911, u5_mult_82_n1910,
         u5_mult_82_n1909, u5_mult_82_n1908, u5_mult_82_n1907,
         u5_mult_82_n1906, u5_mult_82_n1905, u5_mult_82_n1904,
         u5_mult_82_n1903, u5_mult_82_n1902, u5_mult_82_n1901,
         u5_mult_82_n1900, u5_mult_82_n1899, u5_mult_82_n1898,
         u5_mult_82_n1897, u5_mult_82_n1896, u5_mult_82_n1895,
         u5_mult_82_n1894, u5_mult_82_n1893, u5_mult_82_n1892,
         u5_mult_82_n1891, u5_mult_82_n1890, u5_mult_82_n1889,
         u5_mult_82_n1888, u5_mult_82_n1887, u5_mult_82_n1886,
         u5_mult_82_n1885, u5_mult_82_n1884, u5_mult_82_n1883,
         u5_mult_82_n1882, u5_mult_82_n1881, u5_mult_82_n1880,
         u5_mult_82_n1879, u5_mult_82_n1878, u5_mult_82_n1877,
         u5_mult_82_n1876, u5_mult_82_n1875, u5_mult_82_n1874,
         u5_mult_82_n1873, u5_mult_82_n1872, u5_mult_82_n1871,
         u5_mult_82_n1870, u5_mult_82_n1869, u5_mult_82_n1868,
         u5_mult_82_n1867, u5_mult_82_n1866, u5_mult_82_n1865,
         u5_mult_82_n1864, u5_mult_82_n1863, u5_mult_82_n1862,
         u5_mult_82_n1861, u5_mult_82_n1860, u5_mult_82_n1859,
         u5_mult_82_n1858, u5_mult_82_n1857, u5_mult_82_n1856,
         u5_mult_82_n1855, u5_mult_82_n1854, u5_mult_82_n1853,
         u5_mult_82_n1852, u5_mult_82_n1851, u5_mult_82_n1850,
         u5_mult_82_n1849, u5_mult_82_n1848, u5_mult_82_n1847,
         u5_mult_82_n1846, u5_mult_82_n1845, u5_mult_82_n1844,
         u5_mult_82_n1843, u5_mult_82_n1842, u5_mult_82_n1841,
         u5_mult_82_n1840, u5_mult_82_n1839, u5_mult_82_n1838,
         u5_mult_82_n1837, u5_mult_82_n1836, u5_mult_82_n1835,
         u5_mult_82_n1834, u5_mult_82_n1833, u5_mult_82_n1832,
         u5_mult_82_n1831, u5_mult_82_n1830, u5_mult_82_n1829,
         u5_mult_82_n1828, u5_mult_82_n1827, u5_mult_82_n1826,
         u5_mult_82_n1825, u5_mult_82_n1824, u5_mult_82_n1823,
         u5_mult_82_n1822, u5_mult_82_n1821, u5_mult_82_n1820,
         u5_mult_82_n1819, u5_mult_82_n1818, u5_mult_82_n1817,
         u5_mult_82_n1816, u5_mult_82_n1815, u5_mult_82_n1814,
         u5_mult_82_n1813, u5_mult_82_n1812, u5_mult_82_n1811,
         u5_mult_82_n1810, u5_mult_82_n1809, u5_mult_82_n1808,
         u5_mult_82_n1807, u5_mult_82_n1806, u5_mult_82_n1805,
         u5_mult_82_n1804, u5_mult_82_n1803, u5_mult_82_n1802,
         u5_mult_82_n1801, u5_mult_82_n1800, u5_mult_82_n1799,
         u5_mult_82_n1798, u5_mult_82_n1797, u5_mult_82_n1796,
         u5_mult_82_n1795, u5_mult_82_n1794, u5_mult_82_n1793,
         u5_mult_82_n1792, u5_mult_82_n1791, u5_mult_82_n1790,
         u5_mult_82_n1789, u5_mult_82_n1788, u5_mult_82_n1787,
         u5_mult_82_n1786, u5_mult_82_n1785, u5_mult_82_n1784,
         u5_mult_82_n1783, u5_mult_82_n1782, u5_mult_82_n1781,
         u5_mult_82_n1780, u5_mult_82_n1779, u5_mult_82_n1778,
         u5_mult_82_n1777, u5_mult_82_n1776, u5_mult_82_n1775,
         u5_mult_82_n1774, u5_mult_82_n1773, u5_mult_82_n1772,
         u5_mult_82_n1771, u5_mult_82_n1770, u5_mult_82_n1769,
         u5_mult_82_n1768, u5_mult_82_n1767, u5_mult_82_n1766,
         u5_mult_82_n1765, u5_mult_82_n1764, u5_mult_82_n1763,
         u5_mult_82_n1762, u5_mult_82_n1761, u5_mult_82_n1760,
         u5_mult_82_n1759, u5_mult_82_n1758, u5_mult_82_n1757,
         u5_mult_82_n1756, u5_mult_82_n1755, u5_mult_82_n1754,
         u5_mult_82_n1753, u5_mult_82_n1752, u5_mult_82_n1751,
         u5_mult_82_n1750, u5_mult_82_n1749, u5_mult_82_n1748,
         u5_mult_82_n1747, u5_mult_82_n1746, u5_mult_82_n1745,
         u5_mult_82_n1744, u5_mult_82_n1743, u5_mult_82_n1742,
         u5_mult_82_n1741, u5_mult_82_n1740, u5_mult_82_n1739,
         u5_mult_82_n1738, u5_mult_82_n1737, u5_mult_82_n1736,
         u5_mult_82_n1735, u5_mult_82_n1734, u5_mult_82_n1733,
         u5_mult_82_n1732, u5_mult_82_n1731, u5_mult_82_n1730,
         u5_mult_82_n1729, u5_mult_82_n1728, u5_mult_82_n1727,
         u5_mult_82_n1726, u5_mult_82_n1725, u5_mult_82_n1724,
         u5_mult_82_n1723, u5_mult_82_n1722, u5_mult_82_n1721,
         u5_mult_82_n1720, u5_mult_82_n1719, u5_mult_82_n1718,
         u5_mult_82_n1717, u5_mult_82_n1716, u5_mult_82_n1715,
         u5_mult_82_n1714, u5_mult_82_n1713, u5_mult_82_n1712,
         u5_mult_82_n1711, u5_mult_82_n1710, u5_mult_82_n1709,
         u5_mult_82_n1708, u5_mult_82_n1707, u5_mult_82_n1706,
         u5_mult_82_n1705, u5_mult_82_n1704, u5_mult_82_n1703,
         u5_mult_82_n1702, u5_mult_82_n1701, u5_mult_82_n1700,
         u5_mult_82_n1699, u5_mult_82_n1698, u5_mult_82_n1697,
         u5_mult_82_n1696, u5_mult_82_n1695, u5_mult_82_n1694,
         u5_mult_82_n1693, u5_mult_82_n1692, u5_mult_82_n1691,
         u5_mult_82_n1690, u5_mult_82_n1689, u5_mult_82_n1688,
         u5_mult_82_n1687, u5_mult_82_n1686, u5_mult_82_n1685,
         u5_mult_82_n1684, u5_mult_82_n1683, u5_mult_82_n1682,
         u5_mult_82_n1681, u5_mult_82_n1680, u5_mult_82_n1679,
         u5_mult_82_n1678, u5_mult_82_n1677, u5_mult_82_n1676,
         u5_mult_82_n1675, u5_mult_82_n1674, u5_mult_82_n1673,
         u5_mult_82_n1672, u5_mult_82_n1671, u5_mult_82_n1670,
         u5_mult_82_n1669, u5_mult_82_n1668, u5_mult_82_n1667,
         u5_mult_82_n1666, u5_mult_82_n1665, u5_mult_82_n1664,
         u5_mult_82_n1663, u5_mult_82_n1662, u5_mult_82_n1661,
         u5_mult_82_n1660, u5_mult_82_n1659, u5_mult_82_n1658,
         u5_mult_82_n1657, u5_mult_82_n1656, u5_mult_82_n1655,
         u5_mult_82_n1654, u5_mult_82_n1653, u5_mult_82_n1652,
         u5_mult_82_n1651, u5_mult_82_n1650, u5_mult_82_n1649,
         u5_mult_82_n1648, u5_mult_82_n1647, u5_mult_82_n1646,
         u5_mult_82_n1645, u5_mult_82_n1644, u5_mult_82_n1643,
         u5_mult_82_n1642, u5_mult_82_n1641, u5_mult_82_n1640,
         u5_mult_82_n1639, u5_mult_82_n1638, u5_mult_82_n1637,
         u5_mult_82_n1636, u5_mult_82_n1635, u5_mult_82_n1634,
         u5_mult_82_n1633, u5_mult_82_n1632, u5_mult_82_n1631,
         u5_mult_82_n1630, u5_mult_82_n1629, u5_mult_82_n1628,
         u5_mult_82_n1627, u5_mult_82_n1626, u5_mult_82_n1625,
         u5_mult_82_n1624, u5_mult_82_n1623, u5_mult_82_n1622,
         u5_mult_82_n1621, u5_mult_82_n1620, u5_mult_82_n1619,
         u5_mult_82_n1618, u5_mult_82_n1617, u5_mult_82_n1616,
         u5_mult_82_n1615, u5_mult_82_n1614, u5_mult_82_n1613,
         u5_mult_82_n1612, u5_mult_82_n1611, u5_mult_82_n1610,
         u5_mult_82_n1609, u5_mult_82_n1608, u5_mult_82_n1607,
         u5_mult_82_n1606, u5_mult_82_n1605, u5_mult_82_n1604,
         u5_mult_82_n1603, u5_mult_82_n1602, u5_mult_82_n1601,
         u5_mult_82_n1600, u5_mult_82_n1599, u5_mult_82_n1598,
         u5_mult_82_n1597, u5_mult_82_n1596, u5_mult_82_n1595,
         u5_mult_82_n1594, u5_mult_82_n1593, u5_mult_82_n1592,
         u5_mult_82_n1591, u5_mult_82_n1590, u5_mult_82_n1589,
         u5_mult_82_n1588, u5_mult_82_n1587, u5_mult_82_n1586,
         u5_mult_82_n1585, u5_mult_82_n1584, u5_mult_82_n1583,
         u5_mult_82_n1582, u5_mult_82_n1581, u5_mult_82_n1580,
         u5_mult_82_n1579, u5_mult_82_n1578, u5_mult_82_n1577,
         u5_mult_82_n1576, u5_mult_82_n1575, u5_mult_82_n1574,
         u5_mult_82_n1573, u5_mult_82_n1572, u5_mult_82_n1571,
         u5_mult_82_n1570, u5_mult_82_n1569, u5_mult_82_n1568,
         u5_mult_82_n1567, u5_mult_82_n1566, u5_mult_82_n1565,
         u5_mult_82_n1564, u5_mult_82_n1563, u5_mult_82_n1562,
         u5_mult_82_n1561, u5_mult_82_n1560, u5_mult_82_n1559,
         u5_mult_82_n1558, u5_mult_82_n1557, u5_mult_82_n1556,
         u5_mult_82_n1555, u5_mult_82_n1554, u5_mult_82_n1553,
         u5_mult_82_n1552, u5_mult_82_n1551, u5_mult_82_n1550,
         u5_mult_82_n1549, u5_mult_82_n1548, u5_mult_82_n1547,
         u5_mult_82_n1546, u5_mult_82_n1545, u5_mult_82_n1544,
         u5_mult_82_n1543, u5_mult_82_n1542, u5_mult_82_n1541,
         u5_mult_82_n1540, u5_mult_82_n1539, u5_mult_82_n1538,
         u5_mult_82_n1537, u5_mult_82_n1536, u5_mult_82_n1535,
         u5_mult_82_n1534, u5_mult_82_n1533, u5_mult_82_n1532,
         u5_mult_82_n1531, u5_mult_82_n1530, u5_mult_82_n1529,
         u5_mult_82_n1528, u5_mult_82_n1527, u5_mult_82_n1526,
         u5_mult_82_n1525, u5_mult_82_n1524, u5_mult_82_n1523,
         u5_mult_82_n1522, u5_mult_82_n1521, u5_mult_82_n1520,
         u5_mult_82_n1519, u5_mult_82_n1518, u5_mult_82_n1517,
         u5_mult_82_n1516, u5_mult_82_n1515, u5_mult_82_n1514,
         u5_mult_82_n1513, u5_mult_82_n1512, u5_mult_82_n1511,
         u5_mult_82_n1510, u5_mult_82_n1509, u5_mult_82_n1508,
         u5_mult_82_n1507, u5_mult_82_n1506, u5_mult_82_n1505,
         u5_mult_82_n1504, u5_mult_82_n1503, u5_mult_82_n1502,
         u5_mult_82_n1501, u5_mult_82_n1500, u5_mult_82_n1499,
         u5_mult_82_n1498, u5_mult_82_n1497, u5_mult_82_n1496,
         u5_mult_82_n1495, u5_mult_82_n1494, u5_mult_82_n1493,
         u5_mult_82_n1492, u5_mult_82_n1491, u5_mult_82_n1490,
         u5_mult_82_n1489, u5_mult_82_n1488, u5_mult_82_n1487,
         u5_mult_82_n1486, u5_mult_82_n1485, u5_mult_82_n1484,
         u5_mult_82_n1483, u5_mult_82_n1482, u5_mult_82_n1481,
         u5_mult_82_n1480, u5_mult_82_n1479, u5_mult_82_n1478,
         u5_mult_82_n1477, u5_mult_82_n1476, u5_mult_82_n1475,
         u5_mult_82_n1474, u5_mult_82_n1473, u5_mult_82_n1472,
         u5_mult_82_n1471, u5_mult_82_n1470, u5_mult_82_n1469,
         u5_mult_82_n1468, u5_mult_82_n1467, u5_mult_82_n1466,
         u5_mult_82_n1465, u5_mult_82_n1464, u5_mult_82_n1463,
         u5_mult_82_n1462, u5_mult_82_n1461, u5_mult_82_n1460,
         u5_mult_82_n1459, u5_mult_82_n1458, u5_mult_82_n1457,
         u5_mult_82_n1456, u5_mult_82_n1455, u5_mult_82_n1454,
         u5_mult_82_n1453, u5_mult_82_n1452, u5_mult_82_n1451,
         u5_mult_82_n1450, u5_mult_82_n1449, u5_mult_82_n1448,
         u5_mult_82_n1447, u5_mult_82_n1446, u5_mult_82_n1445,
         u5_mult_82_n1444, u5_mult_82_n1443, u5_mult_82_n1442,
         u5_mult_82_n1441, u5_mult_82_n1440, u5_mult_82_n1439,
         u5_mult_82_n1438, u5_mult_82_n1437, u5_mult_82_n1436,
         u5_mult_82_n1435, u5_mult_82_n1434, u5_mult_82_n1433,
         u5_mult_82_n1432, u5_mult_82_n1431, u5_mult_82_n1430,
         u5_mult_82_n1429, u5_mult_82_n1428, u5_mult_82_n1427,
         u5_mult_82_n1426, u5_mult_82_n1425, u5_mult_82_n1424,
         u5_mult_82_n1423, u5_mult_82_n1422, u5_mult_82_n1421,
         u5_mult_82_n1420, u5_mult_82_n1419, u5_mult_82_n1418,
         u5_mult_82_n1417, u5_mult_82_n1416, u5_mult_82_n1415,
         u5_mult_82_n1414, u5_mult_82_n1413, u5_mult_82_n1412,
         u5_mult_82_n1411, u5_mult_82_n1410, u5_mult_82_n1409,
         u5_mult_82_n1408, u5_mult_82_n1407, u5_mult_82_n1406,
         u5_mult_82_n1405, u5_mult_82_n1404, u5_mult_82_n1403,
         u5_mult_82_n1402, u5_mult_82_n1401, u5_mult_82_n1400,
         u5_mult_82_n1399, u5_mult_82_n1398, u5_mult_82_n1397,
         u5_mult_82_n1396, u5_mult_82_n1395, u5_mult_82_n1394,
         u5_mult_82_n1393, u5_mult_82_n1392, u5_mult_82_n1391,
         u5_mult_82_n1390, u5_mult_82_n1389, u5_mult_82_n1388,
         u5_mult_82_n1387, u5_mult_82_n1386, u5_mult_82_n1385,
         u5_mult_82_n1384, u5_mult_82_n1383, u5_mult_82_n1382,
         u5_mult_82_n1381, u5_mult_82_n1380, u5_mult_82_n1379,
         u5_mult_82_n1378, u5_mult_82_n1377, u5_mult_82_n1376,
         u5_mult_82_n1375, u5_mult_82_n1374, u5_mult_82_n1373,
         u5_mult_82_n1372, u5_mult_82_n1371, u5_mult_82_n1370,
         u5_mult_82_n1369, u5_mult_82_n1368, u5_mult_82_n1367,
         u5_mult_82_n1366, u5_mult_82_n1365, u5_mult_82_n1364,
         u5_mult_82_n1363, u5_mult_82_n1362, u5_mult_82_n1361,
         u5_mult_82_n1360, u5_mult_82_n1359, u5_mult_82_n1358,
         u5_mult_82_n1357, u5_mult_82_n1356, u5_mult_82_n1355,
         u5_mult_82_n1354, u5_mult_82_n1353, u5_mult_82_n1352,
         u5_mult_82_n1351, u5_mult_82_n1350, u5_mult_82_n1349,
         u5_mult_82_n1348, u5_mult_82_n1347, u5_mult_82_n1346,
         u5_mult_82_n1345, u5_mult_82_n1344, u5_mult_82_n1343,
         u5_mult_82_n1342, u5_mult_82_n1341, u5_mult_82_n1340,
         u5_mult_82_n1339, u5_mult_82_n1338, u5_mult_82_n1337,
         u5_mult_82_n1336, u5_mult_82_n1335, u5_mult_82_n1334,
         u5_mult_82_n1333, u5_mult_82_n1332, u5_mult_82_n1331,
         u5_mult_82_n1330, u5_mult_82_n1329, u5_mult_82_n1328,
         u5_mult_82_n1327, u5_mult_82_n1326, u5_mult_82_n1325,
         u5_mult_82_n1324, u5_mult_82_n1323, u5_mult_82_n1322,
         u5_mult_82_n1321, u5_mult_82_n1320, u5_mult_82_n1319,
         u5_mult_82_n1318, u5_mult_82_n1317, u5_mult_82_n1316,
         u5_mult_82_n1315, u5_mult_82_n1314, u5_mult_82_n1313,
         u5_mult_82_n1312, u5_mult_82_n1311, u5_mult_82_n1310,
         u5_mult_82_n1309, u5_mult_82_n1308, u5_mult_82_n1307,
         u5_mult_82_n1306, u5_mult_82_n1305, u5_mult_82_n1304,
         u5_mult_82_n1303, u5_mult_82_n1302, u5_mult_82_n1301,
         u5_mult_82_n1300, u5_mult_82_n1299, u5_mult_82_n1298,
         u5_mult_82_n1297, u5_mult_82_n1296, u5_mult_82_n1295,
         u5_mult_82_n1294, u5_mult_82_n1293, u5_mult_82_n1292,
         u5_mult_82_n1291, u5_mult_82_n1290, u5_mult_82_n1289,
         u5_mult_82_n1288, u5_mult_82_n1287, u5_mult_82_n1286,
         u5_mult_82_n1285, u5_mult_82_n1284, u5_mult_82_n1283,
         u5_mult_82_n1282, u5_mult_82_n1281, u5_mult_82_n1280,
         u5_mult_82_n1279, u5_mult_82_n1278, u5_mult_82_n1277,
         u5_mult_82_n1276, u5_mult_82_n1275, u5_mult_82_n1274,
         u5_mult_82_n1273, u5_mult_82_n1272, u5_mult_82_n1271,
         u5_mult_82_n1270, u5_mult_82_n1269, u5_mult_82_n1268,
         u5_mult_82_n1267, u5_mult_82_n1266, u5_mult_82_n1265,
         u5_mult_82_n1264, u5_mult_82_n1263, u5_mult_82_n1262,
         u5_mult_82_n1261, u5_mult_82_n1260, u5_mult_82_n1259,
         u5_mult_82_n1258, u5_mult_82_n1257, u5_mult_82_n1256,
         u5_mult_82_n1255, u5_mult_82_n1254, u5_mult_82_n1253,
         u5_mult_82_n1252, u5_mult_82_n1251, u5_mult_82_n1250,
         u5_mult_82_n1249, u5_mult_82_n1248, u5_mult_82_n1247,
         u5_mult_82_n1246, u5_mult_82_n1245, u5_mult_82_n1244,
         u5_mult_82_n1243, u5_mult_82_n1242, u5_mult_82_n1241,
         u5_mult_82_n1240, u5_mult_82_n1239, u5_mult_82_n1238,
         u5_mult_82_n1237, u5_mult_82_n1236, u5_mult_82_n1235,
         u5_mult_82_n1234, u5_mult_82_n1233, u5_mult_82_n1232,
         u5_mult_82_n1231, u5_mult_82_n1230, u5_mult_82_n1229,
         u5_mult_82_n1228, u5_mult_82_n1227, u5_mult_82_n1226,
         u5_mult_82_n1225, u5_mult_82_n1224, u5_mult_82_n1223,
         u5_mult_82_n1222, u5_mult_82_n1221, u5_mult_82_n1220,
         u5_mult_82_n1219, u5_mult_82_n1218, u5_mult_82_n1217,
         u5_mult_82_n1216, u5_mult_82_n1215, u5_mult_82_n1214,
         u5_mult_82_n1213, u5_mult_82_n1212, u5_mult_82_n1211,
         u5_mult_82_n1210, u5_mult_82_n1209, u5_mult_82_n1208,
         u5_mult_82_n1207, u5_mult_82_n1206, u5_mult_82_n1205,
         u5_mult_82_n1204, u5_mult_82_n1203, u5_mult_82_n1202,
         u5_mult_82_n1201, u5_mult_82_n1200, u5_mult_82_n1199,
         u5_mult_82_n1198, u5_mult_82_n1197, u5_mult_82_n1196,
         u5_mult_82_n1195, u5_mult_82_n1194, u5_mult_82_n1193,
         u5_mult_82_n1192, u5_mult_82_n1191, u5_mult_82_n1190,
         u5_mult_82_n1189, u5_mult_82_n1188, u5_mult_82_n1187,
         u5_mult_82_n1186, u5_mult_82_n1185, u5_mult_82_n1184,
         u5_mult_82_n1183, u5_mult_82_n1182, u5_mult_82_n1181,
         u5_mult_82_n1180, u5_mult_82_n1179, u5_mult_82_n1178,
         u5_mult_82_n1177, u5_mult_82_n1176, u5_mult_82_n1175,
         u5_mult_82_n1174, u5_mult_82_n1173, u5_mult_82_n1172,
         u5_mult_82_n1171, u5_mult_82_n1170, u5_mult_82_n1169,
         u5_mult_82_n1168, u5_mult_82_n1167, u5_mult_82_n1166,
         u5_mult_82_n1165, u5_mult_82_n1164, u5_mult_82_n1163,
         u5_mult_82_n1162, u5_mult_82_n1161, u5_mult_82_n1160,
         u5_mult_82_n1159, u5_mult_82_n1158, u5_mult_82_n1157,
         u5_mult_82_n1156, u5_mult_82_n1155, u5_mult_82_n1154,
         u5_mult_82_n1153, u5_mult_82_n1152, u5_mult_82_n1151,
         u5_mult_82_n1150, u5_mult_82_n1149, u5_mult_82_n1148,
         u5_mult_82_n1147, u5_mult_82_n1146, u5_mult_82_n1145,
         u5_mult_82_n1144, u5_mult_82_n1143, u5_mult_82_n1142,
         u5_mult_82_n1141, u5_mult_82_n1140, u5_mult_82_n1139,
         u5_mult_82_n1138, u5_mult_82_n1137, u5_mult_82_n1136,
         u5_mult_82_n1135, u5_mult_82_n1134, u5_mult_82_n1133,
         u5_mult_82_n1132, u5_mult_82_n1131, u5_mult_82_n1130,
         u5_mult_82_n1129, u5_mult_82_n1128, u5_mult_82_n1127,
         u5_mult_82_n1126, u5_mult_82_n1125, u5_mult_82_n1124,
         u5_mult_82_n1123, u5_mult_82_n1122, u5_mult_82_n1121,
         u5_mult_82_n1120, u5_mult_82_n1119, u5_mult_82_n1118,
         u5_mult_82_n1117, u5_mult_82_n1116, u5_mult_82_n1115,
         u5_mult_82_n1114, u5_mult_82_n1113, u5_mult_82_n1112,
         u5_mult_82_n1111, u5_mult_82_n1110, u5_mult_82_n1109,
         u5_mult_82_n1108, u5_mult_82_n1107, u5_mult_82_n1106,
         u5_mult_82_n1105, u5_mult_82_n1104, u5_mult_82_n1103,
         u5_mult_82_n1102, u5_mult_82_n1101, u5_mult_82_n1100,
         u5_mult_82_n1099, u5_mult_82_n1098, u5_mult_82_n1097,
         u5_mult_82_n1096, u5_mult_82_n1095, u5_mult_82_n1094,
         u5_mult_82_n1093, u5_mult_82_n1092, u5_mult_82_n1091,
         u5_mult_82_n1090, u5_mult_82_n1089, u5_mult_82_n1088,
         u5_mult_82_n1087, u5_mult_82_n1086, u5_mult_82_n1085,
         u5_mult_82_n1084, u5_mult_82_n1083, u5_mult_82_n1082,
         u5_mult_82_n1081, u5_mult_82_n1080, u5_mult_82_n1079,
         u5_mult_82_n1078, u5_mult_82_n1077, u5_mult_82_n1076,
         u5_mult_82_n1075, u5_mult_82_n1074, u5_mult_82_n1073,
         u5_mult_82_n1072, u5_mult_82_n1071, u5_mult_82_n1070,
         u5_mult_82_n1069, u5_mult_82_n1068, u5_mult_82_n1067,
         u5_mult_82_n1066, u5_mult_82_n1065, u5_mult_82_n1064,
         u5_mult_82_n1063, u5_mult_82_n1062, u5_mult_82_n1061,
         u5_mult_82_n1060, u5_mult_82_n1059, u5_mult_82_n1058,
         u5_mult_82_n1057, u5_mult_82_n1056, u5_mult_82_n1055,
         u5_mult_82_n1054, u5_mult_82_n1053, u5_mult_82_n1052,
         u5_mult_82_n1051, u5_mult_82_n1050, u5_mult_82_n1049,
         u5_mult_82_n1048, u5_mult_82_n1047, u5_mult_82_n1046,
         u5_mult_82_n1045, u5_mult_82_n1044, u5_mult_82_n1043,
         u5_mult_82_n1042, u5_mult_82_n1041, u5_mult_82_n1040,
         u5_mult_82_n1039, u5_mult_82_n1038, u5_mult_82_n1037,
         u5_mult_82_n1036, u5_mult_82_n1035, u5_mult_82_n1034,
         u5_mult_82_n1033, u5_mult_82_n1032, u5_mult_82_n1031,
         u5_mult_82_n1030, u5_mult_82_n1029, u5_mult_82_n1028,
         u5_mult_82_n1027, u5_mult_82_n1026, u5_mult_82_n1025,
         u5_mult_82_n1024, u5_mult_82_n1023, u5_mult_82_n1022,
         u5_mult_82_n1021, u5_mult_82_n1020, u5_mult_82_n1019,
         u5_mult_82_n1018, u5_mult_82_n1017, u5_mult_82_n1016,
         u5_mult_82_n1015, u5_mult_82_n1014, u5_mult_82_n1013,
         u5_mult_82_n1012, u5_mult_82_n1011, u5_mult_82_n1010,
         u5_mult_82_n1009, u5_mult_82_n1008, u5_mult_82_n1007,
         u5_mult_82_n1006, u5_mult_82_n1005, u5_mult_82_n1004,
         u5_mult_82_n1003, u5_mult_82_n1002, u5_mult_82_n1001,
         u5_mult_82_n1000, u5_mult_82_n999, u5_mult_82_n998, u5_mult_82_n997,
         u5_mult_82_n996, u5_mult_82_n995, u5_mult_82_n994, u5_mult_82_n993,
         u5_mult_82_n992, u5_mult_82_n991, u5_mult_82_n990, u5_mult_82_n989,
         u5_mult_82_n988, u5_mult_82_n987, u5_mult_82_n986, u5_mult_82_n985,
         u5_mult_82_n984, u5_mult_82_n983, u5_mult_82_n982, u5_mult_82_n981,
         u5_mult_82_n980, u5_mult_82_n979, u5_mult_82_n978, u5_mult_82_n977,
         u5_mult_82_n976, u5_mult_82_n975, u5_mult_82_n974, u5_mult_82_n973,
         u5_mult_82_n972, u5_mult_82_n971, u5_mult_82_n970, u5_mult_82_n969,
         u5_mult_82_n968, u5_mult_82_n967, u5_mult_82_n966, u5_mult_82_n965,
         u5_mult_82_n964, u5_mult_82_n963, u5_mult_82_n962, u5_mult_82_n961,
         u5_mult_82_n960, u5_mult_82_n959, u5_mult_82_n958, u5_mult_82_n957,
         u5_mult_82_n956, u5_mult_82_n955, u5_mult_82_n954, u5_mult_82_n953,
         u5_mult_82_n952, u5_mult_82_n951, u5_mult_82_n950, u5_mult_82_n949,
         u5_mult_82_n948, u5_mult_82_n947, u5_mult_82_n946, u5_mult_82_n945,
         u5_mult_82_n944, u5_mult_82_n943, u5_mult_82_n942, u5_mult_82_n941,
         u5_mult_82_n940, u5_mult_82_n939, u5_mult_82_n938, u5_mult_82_n937,
         u5_mult_82_n936, u5_mult_82_n935, u5_mult_82_n934, u5_mult_82_n933,
         u5_mult_82_n932, u5_mult_82_n931, u5_mult_82_n930, u5_mult_82_n929,
         u5_mult_82_n928, u5_mult_82_n927, u5_mult_82_n926, u5_mult_82_n925,
         u5_mult_82_n924, u5_mult_82_n923, u5_mult_82_n922, u5_mult_82_n921,
         u5_mult_82_n920, u5_mult_82_n919, u5_mult_82_n918, u5_mult_82_n917,
         u5_mult_82_n916, u5_mult_82_n915, u5_mult_82_n914, u5_mult_82_n913,
         u5_mult_82_n912, u5_mult_82_n911, u5_mult_82_n910, u5_mult_82_n909,
         u5_mult_82_n908, u5_mult_82_n907, u5_mult_82_n906, u5_mult_82_n905,
         u5_mult_82_n904, u5_mult_82_n903, u5_mult_82_n902, u5_mult_82_n901,
         u5_mult_82_n900, u5_mult_82_n899, u5_mult_82_n898, u5_mult_82_n897,
         u5_mult_82_n896, u5_mult_82_n895, u5_mult_82_n894, u5_mult_82_n893,
         u5_mult_82_n892, u5_mult_82_n891, u5_mult_82_n890, u5_mult_82_n889,
         u5_mult_82_n888, u5_mult_82_n887, u5_mult_82_n886, u5_mult_82_n885,
         u5_mult_82_n884, u5_mult_82_n883, u5_mult_82_n882, u5_mult_82_n881,
         u5_mult_82_n880, u5_mult_82_n879, u5_mult_82_n878, u5_mult_82_n877,
         u5_mult_82_n876, u5_mult_82_n875, u5_mult_82_n874, u5_mult_82_n873,
         u5_mult_82_n872, u5_mult_82_n871, u5_mult_82_n870, u5_mult_82_n869,
         u5_mult_82_n868, u5_mult_82_n867, u5_mult_82_n866, u5_mult_82_n865,
         u5_mult_82_n864, u5_mult_82_n863, u5_mult_82_n862, u5_mult_82_n861,
         u5_mult_82_n860, u5_mult_82_n859, u5_mult_82_n858, u5_mult_82_n857,
         u5_mult_82_n856, u5_mult_82_n855, u5_mult_82_n854, u5_mult_82_n853,
         u5_mult_82_n852, u5_mult_82_n851, u5_mult_82_n850, u5_mult_82_n849,
         u5_mult_82_n848, u5_mult_82_n847, u5_mult_82_n846, u5_mult_82_n845,
         u5_mult_82_n844, u5_mult_82_n843, u5_mult_82_n842, u5_mult_82_n841,
         u5_mult_82_n840, u5_mult_82_n839, u5_mult_82_n838, u5_mult_82_n837,
         u5_mult_82_n836, u5_mult_82_n835, u5_mult_82_n834, u5_mult_82_n833,
         u5_mult_82_n832, u5_mult_82_n831, u5_mult_82_n830, u5_mult_82_n829,
         u5_mult_82_n828, u5_mult_82_n827, u5_mult_82_n826, u5_mult_82_n825,
         u5_mult_82_n824, u5_mult_82_n823, u5_mult_82_n822, u5_mult_82_n821,
         u5_mult_82_n820, u5_mult_82_n819, u5_mult_82_n818, u5_mult_82_n817,
         u5_mult_82_n816, u5_mult_82_n815, u5_mult_82_n814, u5_mult_82_n813,
         u5_mult_82_n812, u5_mult_82_n811, u5_mult_82_n810, u5_mult_82_n809,
         u5_mult_82_n808, u5_mult_82_n807, u5_mult_82_n806, u5_mult_82_n805,
         u5_mult_82_n804, u5_mult_82_n803, u5_mult_82_n802, u5_mult_82_n801,
         u5_mult_82_n800, u5_mult_82_n799, u5_mult_82_n798, u5_mult_82_n797,
         u5_mult_82_n796, u5_mult_82_n795, u5_mult_82_n794, u5_mult_82_n793,
         u5_mult_82_n792, u5_mult_82_n791, u5_mult_82_n790, u5_mult_82_n789,
         u5_mult_82_n788, u5_mult_82_n787, u5_mult_82_n786, u5_mult_82_n785,
         u5_mult_82_n784, u5_mult_82_n783, u5_mult_82_n782, u5_mult_82_n781,
         u5_mult_82_n780, u5_mult_82_n779, u5_mult_82_n778, u5_mult_82_n777,
         u5_mult_82_n776, u5_mult_82_n775, u5_mult_82_n774, u5_mult_82_n773,
         u5_mult_82_n772, u5_mult_82_n771, u5_mult_82_n770, u5_mult_82_n769,
         u5_mult_82_n768, u5_mult_82_n767, u5_mult_82_n766, u5_mult_82_n765,
         u5_mult_82_n764, u5_mult_82_n763, u5_mult_82_n762, u5_mult_82_n761,
         u5_mult_82_n760, u5_mult_82_n759, u5_mult_82_n758, u5_mult_82_n757,
         u5_mult_82_n756, u5_mult_82_n755, u5_mult_82_n754, u5_mult_82_n753,
         u5_mult_82_n752, u5_mult_82_n751, u5_mult_82_n750, u5_mult_82_n749,
         u5_mult_82_n748, u5_mult_82_n747, u5_mult_82_n746, u5_mult_82_n745,
         u5_mult_82_n744, u5_mult_82_n743, u5_mult_82_n742, u5_mult_82_n741,
         u5_mult_82_n740, u5_mult_82_n739, u5_mult_82_n738, u5_mult_82_n737,
         u5_mult_82_n736, u5_mult_82_n735, u5_mult_82_n734, u5_mult_82_n733,
         u5_mult_82_n732, u5_mult_82_n731, u5_mult_82_n730, u5_mult_82_n729,
         u5_mult_82_n728, u5_mult_82_n727, u5_mult_82_n726, u5_mult_82_n725,
         u5_mult_82_n724, u5_mult_82_n723, u5_mult_82_n722, u5_mult_82_n721,
         u5_mult_82_n720, u5_mult_82_n719, u5_mult_82_n718, u5_mult_82_n717,
         u5_mult_82_n716, u5_mult_82_n715, u5_mult_82_n714, u5_mult_82_n713,
         u5_mult_82_n712, u5_mult_82_n711, u5_mult_82_n710, u5_mult_82_n709,
         u5_mult_82_n708, u5_mult_82_n707, u5_mult_82_n706, u5_mult_82_n705,
         u5_mult_82_n704, u5_mult_82_n703, u5_mult_82_n702, u5_mult_82_n701,
         u5_mult_82_n700, u5_mult_82_n699, u5_mult_82_n698, u5_mult_82_n697,
         u5_mult_82_n696, u5_mult_82_n695, u5_mult_82_n694, u5_mult_82_n693,
         u5_mult_82_n692, u5_mult_82_n691, u5_mult_82_n690, u5_mult_82_n689,
         u5_mult_82_n688, u5_mult_82_n687, u5_mult_82_n686, u5_mult_82_n685,
         u5_mult_82_n684, u5_mult_82_n683, u5_mult_82_n682, u5_mult_82_n681,
         u5_mult_82_n680, u5_mult_82_n679, u5_mult_82_n678, u5_mult_82_n677,
         u5_mult_82_n676, u5_mult_82_n675, u5_mult_82_n674, u5_mult_82_n673,
         u5_mult_82_n672, u5_mult_82_n671, u5_mult_82_n670, u5_mult_82_n669,
         u5_mult_82_n668, u5_mult_82_n667, u5_mult_82_n666, u5_mult_82_n665,
         u5_mult_82_n664, u5_mult_82_n663, u5_mult_82_n662, u5_mult_82_n661,
         u5_mult_82_n660, u5_mult_82_n659, u5_mult_82_n658, u5_mult_82_n657,
         u5_mult_82_n656, u5_mult_82_n655, u5_mult_82_n654, u5_mult_82_n653,
         u5_mult_82_n652, u5_mult_82_n651, u5_mult_82_n650, u5_mult_82_n649,
         u5_mult_82_n648, u5_mult_82_n647, u5_mult_82_n646, u5_mult_82_n645,
         u5_mult_82_n644, u5_mult_82_n643, u5_mult_82_n642, u5_mult_82_n641,
         u5_mult_82_n640, u5_mult_82_n639, u5_mult_82_n638, u5_mult_82_n637,
         u5_mult_82_n636, u5_mult_82_n635, u5_mult_82_n634, u5_mult_82_n633,
         u5_mult_82_n632, u5_mult_82_n631, u5_mult_82_n630, u5_mult_82_n629,
         u5_mult_82_n627, u5_mult_82_n626, u5_mult_82_n624, u5_mult_82_n623,
         u5_mult_82_n622, u5_mult_82_n621, u5_mult_82_n620, u5_mult_82_n619,
         u5_mult_82_n618, u5_mult_82_n617, u5_mult_82_n616, u5_mult_82_n615,
         u5_mult_82_n614, u5_mult_82_n613, u5_mult_82_n612, u5_mult_82_n611,
         u5_mult_82_n610, u5_mult_82_n609, u5_mult_82_n608, u5_mult_82_n607,
         u5_mult_82_n606, u5_mult_82_n605, u5_mult_82_n604, u5_mult_82_n603,
         u5_mult_82_n602, u5_mult_82_n601, u5_mult_82_n600, u5_mult_82_n599,
         u5_mult_82_n598, u5_mult_82_n597, u5_mult_82_n596, u5_mult_82_n595,
         u5_mult_82_n594, u5_mult_82_n593, u5_mult_82_n592, u5_mult_82_n591,
         u5_mult_82_n590, u5_mult_82_n589, u5_mult_82_n588, u5_mult_82_n587,
         u5_mult_82_n586, u5_mult_82_n585, u5_mult_82_n584, u5_mult_82_n583,
         u5_mult_82_n582, u5_mult_82_n581, u5_mult_82_n580, u5_mult_82_n579,
         u5_mult_82_n578, u5_mult_82_n577, u5_mult_82_n576, u5_mult_82_n575,
         u5_mult_82_n574, u5_mult_82_n573, u5_mult_82_n572, u5_mult_82_n571,
         u5_mult_82_n570, u5_mult_82_n569, u5_mult_82_n568, u5_mult_82_n567,
         u5_mult_82_n566, u5_mult_82_n565, u5_mult_82_n564, u5_mult_82_n563,
         u5_mult_82_n562, u5_mult_82_n561, u5_mult_82_n560, u5_mult_82_n559,
         u5_mult_82_n558, u5_mult_82_n557, u5_mult_82_n556, u5_mult_82_n555,
         u5_mult_82_n554, u5_mult_82_n553, u5_mult_82_n552, u5_mult_82_n551,
         u5_mult_82_n550, u5_mult_82_n549, u5_mult_82_n548, u5_mult_82_n547,
         u5_mult_82_n546, u5_mult_82_n545, u5_mult_82_n544, u5_mult_82_n543,
         u5_mult_82_n542, u5_mult_82_n541, u5_mult_82_n540, u5_mult_82_n539,
         u5_mult_82_n538, u5_mult_82_n537, u5_mult_82_n536, u5_mult_82_n535,
         u5_mult_82_n534, u5_mult_82_n533, u5_mult_82_n532, u5_mult_82_n531,
         u5_mult_82_n530, u5_mult_82_n529, u5_mult_82_n528, u5_mult_82_n527,
         u5_mult_82_n526, u5_mult_82_n525, u5_mult_82_n524, u5_mult_82_n523,
         u5_mult_82_n522, u5_mult_82_n521, u5_mult_82_n520, u5_mult_82_n519,
         u5_mult_82_n518, u5_mult_82_n517, u5_mult_82_n516, u5_mult_82_n515,
         u5_mult_82_n514, u5_mult_82_n513, u5_mult_82_n512, u5_mult_82_n511,
         u5_mult_82_n510, u5_mult_82_n509, u5_mult_82_n508, u5_mult_82_n507,
         u5_mult_82_n506, u5_mult_82_n505, u5_mult_82_n504, u5_mult_82_n503,
         u5_mult_82_n502, u5_mult_82_n501, u5_mult_82_n500, u5_mult_82_n499,
         u5_mult_82_n498, u5_mult_82_n497, u5_mult_82_n496, u5_mult_82_n495,
         u5_mult_82_n494, u5_mult_82_n493, u5_mult_82_n492, u5_mult_82_n491,
         u5_mult_82_n490, u5_mult_82_n489, u5_mult_82_n488, u5_mult_82_n487,
         u5_mult_82_n486, u5_mult_82_n485, u5_mult_82_n484, u5_mult_82_n483,
         u5_mult_82_n482, u5_mult_82_n481, u5_mult_82_n480, u5_mult_82_n479,
         u5_mult_82_n478, u5_mult_82_n477, u5_mult_82_n476, u5_mult_82_n475,
         u5_mult_82_n474, u5_mult_82_n473, u5_mult_82_n472, u5_mult_82_n471,
         u5_mult_82_n470, u5_mult_82_n469, u5_mult_82_n468, u5_mult_82_n467,
         u5_mult_82_n466, u5_mult_82_n465, u5_mult_82_n464, u5_mult_82_n463,
         u5_mult_82_n462, u5_mult_82_n461, u5_mult_82_n460, u5_mult_82_n459,
         u5_mult_82_n458, u5_mult_82_n457, u5_mult_82_n456, u5_mult_82_n455,
         u5_mult_82_n454, u5_mult_82_n453, u5_mult_82_n452, u5_mult_82_n451,
         u5_mult_82_n450, u5_mult_82_n449, u5_mult_82_n448, u5_mult_82_n447,
         u5_mult_82_n446, u5_mult_82_n445, u5_mult_82_n444, u5_mult_82_n443,
         u5_mult_82_n442, u5_mult_82_n441, u5_mult_82_n440, u5_mult_82_n439,
         u5_mult_82_n438, u5_mult_82_n437, u5_mult_82_n436, u5_mult_82_n435,
         u5_mult_82_n434, u5_mult_82_n433, u5_mult_82_n432, u5_mult_82_n431,
         u5_mult_82_n430, u5_mult_82_n429, u5_mult_82_n428, u5_mult_82_n427,
         u5_mult_82_n426, u5_mult_82_n425, u5_mult_82_n424, u5_mult_82_n423,
         u5_mult_82_n422, u5_mult_82_n421, u5_mult_82_n420, u5_mult_82_n419,
         u5_mult_82_n418, u5_mult_82_n417, u5_mult_82_n416, u5_mult_82_n415,
         u5_mult_82_n414, u5_mult_82_n413, u5_mult_82_n412, u5_mult_82_n411,
         u5_mult_82_n410, u5_mult_82_n409, u5_mult_82_n408, u5_mult_82_n407,
         u5_mult_82_n406, u5_mult_82_n405, u5_mult_82_n404, u5_mult_82_n403,
         u5_mult_82_n402, u5_mult_82_n401, u5_mult_82_n400, u5_mult_82_n399,
         u5_mult_82_n398, u5_mult_82_n397, u5_mult_82_n396, u5_mult_82_n395,
         u5_mult_82_n394, u5_mult_82_n393, u5_mult_82_n392, u5_mult_82_n391,
         u5_mult_82_n390, u5_mult_82_n389, u5_mult_82_n388, u5_mult_82_n387,
         u5_mult_82_n386, u5_mult_82_n385, u5_mult_82_n384, u5_mult_82_n383,
         u5_mult_82_n382, u5_mult_82_n381, u5_mult_82_n380, u5_mult_82_n379,
         u5_mult_82_n378, u5_mult_82_n377, u5_mult_82_n376, u5_mult_82_n375,
         u5_mult_82_n374, u5_mult_82_n373, u5_mult_82_n372, u5_mult_82_n371,
         u5_mult_82_n370, u5_mult_82_n369, u5_mult_82_n368, u5_mult_82_n367,
         u5_mult_82_n366, u5_mult_82_n365, u5_mult_82_n364, u5_mult_82_n363,
         u5_mult_82_n362, u5_mult_82_n361, u5_mult_82_n360, u5_mult_82_n359,
         u5_mult_82_n358, u5_mult_82_n357, u5_mult_82_n356, u5_mult_82_n355,
         u5_mult_82_n354, u5_mult_82_n353, u5_mult_82_n352, u5_mult_82_n351,
         u5_mult_82_n350, u5_mult_82_n349, u5_mult_82_n348, u5_mult_82_n347,
         u5_mult_82_n346, u5_mult_82_n345, u5_mult_82_n344, u5_mult_82_n343,
         u5_mult_82_n342, u5_mult_82_n341, u5_mult_82_n340, u5_mult_82_n339,
         u5_mult_82_n338, u5_mult_82_n337, u5_mult_82_n336, u5_mult_82_n335,
         u5_mult_82_n334, u5_mult_82_n333, u5_mult_82_n332, u5_mult_82_n331,
         u5_mult_82_n330, u5_mult_82_n329, u5_mult_82_n328, u5_mult_82_n327,
         u5_mult_82_n326, u5_mult_82_n325, u5_mult_82_n324, u5_mult_82_n323,
         u5_mult_82_n322, u5_mult_82_n321, u5_mult_82_n320, u5_mult_82_n319,
         u5_mult_82_n318, u5_mult_82_n317, u5_mult_82_n316, u5_mult_82_n315,
         u5_mult_82_n314, u5_mult_82_n313, u5_mult_82_n312, u5_mult_82_n311,
         u5_mult_82_n310, u5_mult_82_n309, u5_mult_82_n308, u5_mult_82_n307,
         u5_mult_82_n306, u5_mult_82_n305, u5_mult_82_n304, u5_mult_82_n303,
         u5_mult_82_n302, u5_mult_82_n301, u5_mult_82_n300, u5_mult_82_n299,
         u5_mult_82_n298, u5_mult_82_n297, u5_mult_82_n296, u5_mult_82_n295,
         u5_mult_82_n294, u5_mult_82_n293, u5_mult_82_n292, u5_mult_82_n291,
         u5_mult_82_n290, u5_mult_82_n289, u5_mult_82_n288, u5_mult_82_n287,
         u5_mult_82_n286, u5_mult_82_n285, u5_mult_82_n284, u5_mult_82_n283,
         u5_mult_82_n282, u5_mult_82_n281, u5_mult_82_n280, u5_mult_82_n279,
         u5_mult_82_n278, u5_mult_82_n277, u5_mult_82_n276, u5_mult_82_n275,
         u5_mult_82_n274, u5_mult_82_n273, u5_mult_82_n272, u5_mult_82_n271,
         u5_mult_82_n270, u5_mult_82_n269, u5_mult_82_n268, u5_mult_82_n267,
         u5_mult_82_n266, u5_mult_82_n265, u5_mult_82_n264, u5_mult_82_n263,
         u5_mult_82_n262, u5_mult_82_n261, u5_mult_82_n260, u5_mult_82_n259,
         u5_mult_82_n258, u5_mult_82_n257, u5_mult_82_n256, u5_mult_82_n255,
         u5_mult_82_n254, u5_mult_82_n253, u5_mult_82_n252, u5_mult_82_n251,
         u5_mult_82_n250, u5_mult_82_n249, u5_mult_82_n248, u5_mult_82_n247,
         u5_mult_82_n246, u5_mult_82_n245, u5_mult_82_n244, u5_mult_82_n243,
         u5_mult_82_n242, u5_mult_82_n241, u5_mult_82_n240, u5_mult_82_n239,
         u5_mult_82_n238, u5_mult_82_n237, u5_mult_82_n236, u5_mult_82_n235,
         u5_mult_82_n234, u5_mult_82_n233, u5_mult_82_n232, u5_mult_82_n231,
         u5_mult_82_n230, u5_mult_82_n229, u5_mult_82_n228, u5_mult_82_n227,
         u5_mult_82_n226, u5_mult_82_n225, u5_mult_82_n224, u5_mult_82_n223,
         u5_mult_82_n222, u5_mult_82_n221, u5_mult_82_n220, u5_mult_82_n219,
         u5_mult_82_n218, u5_mult_82_n217, u5_mult_82_n216, u5_mult_82_n215,
         u5_mult_82_n214, u5_mult_82_n213, u5_mult_82_n212, u5_mult_82_n211,
         u5_mult_82_n210, u5_mult_82_n209, u5_mult_82_n208, u5_mult_82_n207,
         u5_mult_82_n206, u5_mult_82_n205, u5_mult_82_n204, u5_mult_82_n203,
         u5_mult_82_n202, u5_mult_82_n201, u5_mult_82_n200, u5_mult_82_n199,
         u5_mult_82_n198, u5_mult_82_n197, u5_mult_82_n196, u5_mult_82_n195,
         u5_mult_82_n194, u5_mult_82_n193, u5_mult_82_n192, u5_mult_82_n191,
         u5_mult_82_n190, u5_mult_82_n189, u5_mult_82_n188, u5_mult_82_n187,
         u5_mult_82_n186, u5_mult_82_n185, u5_mult_82_n184, u5_mult_82_n183,
         u5_mult_82_n182, u5_mult_82_n181, u5_mult_82_n180, u5_mult_82_n179,
         u5_mult_82_n178, u5_mult_82_n177, u5_mult_82_n176, u5_mult_82_n175,
         u5_mult_82_n174, u5_mult_82_n173, u5_mult_82_n172, u5_mult_82_n171,
         u5_mult_82_n170, u5_mult_82_n169, u5_mult_82_n168, u5_mult_82_n167,
         u5_mult_82_n166, u5_mult_82_n165, u5_mult_82_n164, u5_mult_82_n163,
         u5_mult_82_n162, u5_mult_82_n161, u5_mult_82_n160, u5_mult_82_n159,
         u5_mult_82_n158, u5_mult_82_n157, u5_mult_82_n156, u5_mult_82_n155,
         u5_mult_82_n154, u5_mult_82_n153, u5_mult_82_n152, u5_mult_82_n151,
         u5_mult_82_n150, u5_mult_82_n149, u5_mult_82_n148, u5_mult_82_n147,
         u5_mult_82_n146, u5_mult_82_n145, u5_mult_82_n144, u5_mult_82_n143,
         u5_mult_82_n142, u5_mult_82_n141, u5_mult_82_n140, u5_mult_82_n139,
         u5_mult_82_n138, u5_mult_82_n137, u5_mult_82_n136, u5_mult_82_n135,
         u5_mult_82_n134, u5_mult_82_n133, u5_mult_82_n132, u5_mult_82_n131,
         u5_mult_82_n130, u5_mult_82_n129, u5_mult_82_n128, u5_mult_82_n127,
         u5_mult_82_n126, u5_mult_82_n125, u5_mult_82_n124, u5_mult_82_n123,
         u5_mult_82_n122, u5_mult_82_n121, u5_mult_82_n120, u5_mult_82_n119,
         u5_mult_82_n118, u5_mult_82_n117, u5_mult_82_n116, u5_mult_82_n115,
         u5_mult_82_n114, u5_mult_82_n113, u5_mult_82_n112, u5_mult_82_n111,
         u5_mult_82_n110, u5_mult_82_n109, u5_mult_82_n108, u5_mult_82_n107,
         u5_mult_82_n106, u5_mult_82_n105, u5_mult_82_n104, u5_mult_82_n103,
         u5_mult_82_n102, u5_mult_82_n101, u5_mult_82_n100, u5_mult_82_n99,
         u5_mult_82_n98, u5_mult_82_n97, u5_mult_82_n96, u5_mult_82_n95,
         u5_mult_82_n94, u5_mult_82_n93, u5_mult_82_n92, u5_mult_82_n91,
         u5_mult_82_n90, u5_mult_82_n89, u5_mult_82_n88, u5_mult_82_n87,
         u5_mult_82_n86, u5_mult_82_n85, u5_mult_82_n84, u5_mult_82_n83,
         u5_mult_82_n82, u5_mult_82_n81, u5_mult_82_n80, u5_mult_82_n79,
         u5_mult_82_n78, u5_mult_82_n77, u5_mult_82_n76, u5_mult_82_n75,
         u5_mult_82_n74, u5_mult_82_n73, u5_mult_82_n72, u5_mult_82_n71,
         u5_mult_82_n70, u5_mult_82_n69, u5_mult_82_n68, u5_mult_82_n67,
         u5_mult_82_n66, u5_mult_82_n65, u5_mult_82_n64, u5_mult_82_n63,
         u5_mult_82_n62, u5_mult_82_n61, u5_mult_82_n60, u5_mult_82_n59,
         u5_mult_82_n58, u5_mult_82_n57, u5_mult_82_n56, u5_mult_82_n55,
         u5_mult_82_n54, u5_mult_82_n53, u5_mult_82_n52, u5_mult_82_n51,
         u5_mult_82_n50, u5_mult_82_n49, u5_mult_82_n48, u5_mult_82_n47,
         u5_mult_82_n46, u5_mult_82_n45, u5_mult_82_n44, u5_mult_82_n43,
         u5_mult_82_n42, u5_mult_82_n41, u5_mult_82_n40, u5_mult_82_n39,
         u5_mult_82_n38, u5_mult_82_n37, u5_mult_82_n36, u5_mult_82_n35,
         u5_mult_82_n34, u5_mult_82_n33, u5_mult_82_n32, u5_mult_82_n31,
         u5_mult_82_n30, u5_mult_82_n29, u5_mult_82_n28, u5_mult_82_n27,
         u5_mult_82_n26, u5_mult_82_n25, u5_mult_82_n24, u5_mult_82_n23,
         u5_mult_82_n22, u5_mult_82_n21, u5_mult_82_n20, u5_mult_82_n19,
         u5_mult_82_n18, u5_mult_82_n17, u5_mult_82_n16, u5_mult_82_n15,
         u5_mult_82_n14, u5_mult_82_n13, u5_mult_82_n12, u5_mult_82_n11,
         u5_mult_82_n10, u5_mult_82_n9, u5_mult_82_n8, u5_mult_82_n7,
         u5_mult_82_n6, u5_mult_82_n5, u5_mult_82_n4, u5_mult_82_n3,
         u5_mult_82__UDW__88988_net69760, u5_mult_82_CARRYB_1__36_,
         u5_mult_82_CARRYB_2__36_, u5_mult_82_CARRYB_3__35_,
         u5_mult_82_SUMB_2__36_, u5_mult_82_SUMB_3__35_, u5_mult_82_ab_0__37_,
         u5_mult_82_CARRYB_49__6_, u5_mult_82_CARRYB_50__6_,
         u5_mult_82_SUMB_49__7_, u5_mult_82_ab_50__6_, u5_mult_82_net57179,
         u5_mult_82_net78900, u5_mult_82_net78901, u5_mult_82_net84846,
         u5_mult_82_CARRYB_39__12_, u5_mult_82_CARRYB_40__12_,
         u5_mult_82_SUMB_39__13_, u5_mult_82_ab_40__12_, u5_mult_82_net64495,
         u5_mult_82_net82471, u5_mult_82_net82472, u5_mult_82_net85894,
         u5_mult_82_CARRYB_44__9_, u5_mult_82_CARRYB_45__9_,
         u5_mult_82_SUMB_44__10_, u5_mult_82_ab_45__9_, u5_mult_82_net79320,
         u5_mult_82_net79321, u5_mult_82_net83142, u5_mult_82_CARRYB_50__5_,
         u5_mult_82_CARRYB_51__4_, u5_mult_82_CARRYB_51__5_,
         u5_mult_82_CARRYB_52__4_, u5_mult_82_SUMB_49__6_,
         u5_mult_82_SUMB_50__5_, u5_mult_82_SUMB_50__6_,
         u5_mult_82_SUMB_51__5_, u5_mult_82_SUMB_51__6_,
         u5_mult_82_SUMB_52__5_, u5_mult_82_ab_50__5_, u5_mult_82_net78789,
         u5_mult_82_net80802, u5_mult_82_net86159, u5_mult_82_net87687,
         u5_mult_82_net87846, u5_mult_82_net87847, u5_mult_82_CARRYB_4__34_,
         u5_mult_82_CARRYB_5__34_, u5_mult_82_SUMB_3__36_,
         u5_mult_82_SUMB_4__35_, u5_mult_82_SUMB_5__34_, u5_mult_82_ab_5__34_,
         u5_mult_82_net57160, u5_mult_82_net80613, u5_mult_82_net83295,
         u5_mult_82_net83296, u5_mult_82_net85316, u5_mult_82_net85323,
         u5_mult_82_CARRYB_6__34_, u5_mult_82_SUMB_5__35_,
         u5_mult_82_SUMB_6__34_, u5_mult_82_CARRYB_25__22_,
         u5_mult_82_CARRYB_26__21_, u5_mult_82_CARRYB_27__20_,
         u5_mult_82_CARRYB_28__20_, u5_mult_82_CARRYB_29__19_,
         u5_mult_82_CARRYB_30__18_, u5_mult_82_SUMB_24__23_,
         u5_mult_82_SUMB_25__22_, u5_mult_82_SUMB_26__21_,
         u5_mult_82_SUMB_27__20_, u5_mult_82_SUMB_28__20_,
         u5_mult_82_SUMB_29__19_, u5_mult_82_CARRYB_16__28_,
         u5_mult_82_CARRYB_18__26_, u5_mult_82_CARRYB_19__26_,
         u5_mult_82_SUMB_15__29_, u5_mult_82_SUMB_16__28_,
         u5_mult_82_SUMB_17__27_, u5_mult_82_SUMB_18__26_,
         u5_mult_82_SUMB_18__27_, u5_mult_82_SUMB_19__26_,
         u5_mult_82_SUMB_20__25_, u5_mult_82_CARRYB_41__11_,
         u5_mult_82_SUMB_41__12_, u5_mult_82_SUMB_42__11_,
         u5_mult_82_ab_42__11_, u5_mult_82_net83870, u5_mult_82_net86284,
         u5_mult_82_CARRYB_41__13_, u5_mult_82_CARRYB_42__12_,
         u5_mult_82_CARRYB_43__11_, u5_mult_82_SUMB_40__14_,
         u5_mult_82_SUMB_41__13_, u5_mult_82_SUMB_42__12_,
         u5_mult_82_SUMB_43__11_, u5_mult_82_ab_41__13_,
         u5_mult_82_CARRYB_10__32_, u5_mult_82_CARRYB_11__31_,
         u5_mult_82_CARRYB_12__30_, u5_mult_82_CARRYB_13__29_,
         u5_mult_82_CARRYB_14__28_, u5_mult_82_CARRYB_15__27_,
         u5_mult_82_CARRYB_6__35_, u5_mult_82_CARRYB_7__34_,
         u5_mult_82_CARRYB_8__33_, u5_mult_82_CARRYB_9__32_,
         u5_mult_82_CARRYB_9__33_, u5_mult_82_SUMB_10__32_,
         u5_mult_82_SUMB_10__33_, u5_mult_82_SUMB_11__31_,
         u5_mult_82_SUMB_11__32_, u5_mult_82_SUMB_12__30_,
         u5_mult_82_SUMB_12__31_, u5_mult_82_SUMB_13__29_,
         u5_mult_82_SUMB_14__28_, u5_mult_82_SUMB_15__27_,
         u5_mult_82_SUMB_6__35_, u5_mult_82_SUMB_7__34_,
         u5_mult_82_SUMB_8__33_, u5_mult_82_SUMB_8__34_,
         u5_mult_82_SUMB_9__33_, u5_mult_82_CARRYB_34__16_,
         u5_mult_82_CARRYB_35__15_, u5_mult_82_CARRYB_36__14_,
         u5_mult_82_SUMB_33__17_, u5_mult_82_SUMB_34__16_,
         u5_mult_82_SUMB_35__15_, u5_mult_82_SUMB_36__14_,
         u5_mult_82_SUMB_36__15_, u5_mult_82_SUMB_37__14_,
         u5_mult_82_ab_34__16_, u5_mult_82_net79082, u5_mult_82_net81198,
         u5_mult_82_net81421, u5_mult_82_net81422, u5_mult_82_net83710,
         u5_mult_82_CARRYB_46__8_, u5_mult_82_CARRYB_47__8_,
         u5_mult_82_CARRYB_48__7_, u5_mult_82_SUMB_46__9_,
         u5_mult_82_SUMB_47__8_, u5_mult_82_SUMB_48__8_, u5_mult_82_ab_47__8_,
         u5_mult_82_net81824, u5_mult_82_CARRYB_22__23_,
         u5_mult_82_CARRYB_23__23_, u5_mult_82_SUMB_22__24_,
         u5_mult_82_SUMB_23__23_, u5_mult_82_ab_23__23_,
         u5_mult_82_SUMB_50__7_, u5_mult_82_ab_51__6_,
         u5_mult_82_CARRYB_37__14_, u5_mult_82_CARRYB_38__14_,
         u5_mult_82_SUMB_37__15_, u5_mult_82_SUMB_38__14_,
         u5_mult_82_ab_38__14_, u5_mult_82_net79087, u5_mult_82_net79088,
         u5_mult_82_net79089, u5_mult_82_CARRYB_5__35_, u5_mult_82_SUMB_5__36_,
         u5_mult_82_ab_6__35_, u5_mult_82_SUMB_29__20_,
         u5_mult_82_SUMB_30__19_, u5_mult_82_SUMB_31__18_, u5_mult_82_net79209,
         u5_mult_82_net82042, u5_mult_82_net86279, u5_mult_82_net86280,
         u5_mult_82_net86281, u5_mult_82_net87269, u5_mult_82_ab_43__10_,
         u5_mult_82_net78856, u5_mult_82_net78857, u5_mult_82_SUMB_40__13_,
         u5_mult_82_ab_41__12_, u5_mult_82_net64497, u5_mult_82_net64499,
         u5_mult_82_net64569, u5_mult_82_net64571, u5_mult_82_net65521,
         u5_mult_82_net65525, u5_mult_82_ab_25__22_, u5_mult_82_net88595,
         u5_mult_82_net88132, u5_mult_82_net88030, u5_mult_82_net87436,
         u5_mult_82_net87435, u5_mult_82_net87429, u5_mult_82_net87430,
         u5_mult_82_net87325, u5_mult_82_net86976, u5_mult_82_net86966,
         u5_mult_82_net86863, u5_mult_82_net86784, u5_mult_82_net86785,
         u5_mult_82_net86288, u5_mult_82_net86289, u5_mult_82_net86290,
         u5_mult_82_net86084, u5_mult_82_net86085, u5_mult_82_net85540,
         u5_mult_82_net85541, u5_mult_82_net85371, u5_mult_82_net85372,
         u5_mult_82_net85373, u5_mult_82_net84888, u5_mult_82_net84890,
         u5_mult_82_net84845, u5_mult_82_net84599, u5_mult_82_net84601,
         u5_mult_82_net84580, u5_mult_82_net84453, u5_mult_82_net84440,
         u5_mult_82_net84441, u5_mult_82_net84443, u5_mult_82_net84193,
         u5_mult_82_net84194, u5_mult_82_net84199, u5_mult_82_net83655,
         u5_mult_82_net83288, u5_mult_82_net83289, u5_mult_82_net83290,
         u5_mult_82_net83292, u5_mult_82_net83293, u5_mult_82_net83273,
         u5_mult_82_net83274, u5_mult_82_net83139, u5_mult_82_net83047,
         u5_mult_82_net82990, u5_mult_82_net82676, u5_mult_82_net82678,
         u5_mult_82_net82468, u5_mult_82_net82469, u5_mult_82_net82039,
         u5_mult_82_net82040, u5_mult_82_net82046, u5_mult_82_net82047,
         u5_mult_82_net82048, u5_mult_82_net82055, u5_mult_82_net82056,
         u5_mult_82_net81962, u5_mult_82_net81825, u5_mult_82_net81827,
         u5_mult_82_net81828, u5_mult_82_net81829, u5_mult_82_net81830,
         u5_mult_82_net81531, u5_mult_82_net81534, u5_mult_82_net81536,
         u5_mult_82_net81427, u5_mult_82_net81428, u5_mult_82_net81335,
         u5_mult_82_net80793, u5_mult_82_net80795, u5_mult_82_net80797,
         u5_mult_82_net80806, u5_mult_82_net80807, u5_mult_82_net80808,
         u5_mult_82_net80786, u5_mult_82_net80645, u5_mult_82_net80647,
         u5_mult_82_net80614, u5_mult_82_net80616, u5_mult_82_net80618,
         u5_mult_82_net80619, u5_mult_82_net80535, u5_mult_82_net80537,
         u5_mult_82_net80542, u5_mult_82_net80543, u5_mult_82_net80364,
         u5_mult_82_net80252, u5_mult_82_net80254, u5_mult_82_net80255,
         u5_mult_82_net80183, u5_mult_82_net80185, u5_mult_82_net80187,
         u5_mult_82_net80188, u5_mult_82_net80190, u5_mult_82_net80099,
         u5_mult_82_net79785, u5_mult_82_net79786, u5_mult_82_net79780,
         u5_mult_82_net79444, u5_mult_82_net79446, u5_mult_82_net79317,
         u5_mult_82_net79318, u5_mult_82_net79263, u5_mult_82_net79208,
         u5_mult_82_net79210, u5_mult_82_net79212, u5_mult_82_net79213,
         u5_mult_82_net79214, u5_mult_82_net79215, u5_mult_82_net79084,
         u5_mult_82_net79086, u5_mult_82_net78954, u5_mult_82_net78850,
         u5_mult_82_net78851, u5_mult_82_net78852, u5_mult_82_net78853,
         u5_mult_82_net78790, u5_mult_82_net78791, u5_mult_82_net78792,
         u5_mult_82__UDW__89408_net70938, u5_mult_82__UDW__88983_net69746,
         u5_mult_82_net66121, u5_mult_82_net66107, u5_mult_82_net66109,
         u5_mult_82_net66111, u5_mult_82_net66087, u5_mult_82_net66089,
         u5_mult_82_net66091, u5_mult_82_net66093, u5_mult_82_net66097,
         u5_mult_82_net66033, u5_mult_82_net66035, u5_mult_82_net66037,
         u5_mult_82_net66039, u5_mult_82_net66041, u5_mult_82_net66043,
         u5_mult_82_net66017, u5_mult_82_net66019, u5_mult_82_net66021,
         u5_mult_82_net66023, u5_mult_82_net66025, u5_mult_82_net65711,
         u5_mult_82_net65713, u5_mult_82_net65717, u5_mult_82_net65721,
         u5_mult_82_net65675, u5_mult_82_net65677, u5_mult_82_net65679,
         u5_mult_82_net65681, u5_mult_82_net65685, u5_mult_82_net65513,
         u5_mult_82_net65515, u5_mult_82_net65517, u5_mult_82_net65519,
         u5_mult_82_net65523, u5_mult_82_net65441, u5_mult_82_net65443,
         u5_mult_82_net65445, u5_mult_82_net65447, u5_mult_82_net65451,
         u5_mult_82_net65403, u5_mult_82_net65405, u5_mult_82_net65407,
         u5_mult_82_net65409, u5_mult_82_net65411, u5_mult_82_net65385,
         u5_mult_82_net65387, u5_mult_82_net65389, u5_mult_82_net65391,
         u5_mult_82_net65393, u5_mult_82_net65369, u5_mult_82_net65371,
         u5_mult_82_net65373, u5_mult_82_net65375, u5_mult_82_net65379,
         u5_mult_82_net65349, u5_mult_82_net65351, u5_mult_82_net65353,
         u5_mult_82_net65355, u5_mult_82_net65361, u5_mult_82_net65313,
         u5_mult_82_net65315, u5_mult_82_net65319, u5_mult_82_net65321,
         u5_mult_82_net65293, u5_mult_82_net65277, u5_mult_82_net65279,
         u5_mult_82_net65283, u5_mult_82_net65285, u5_mult_82_net65287,
         u5_mult_82_net65223, u5_mult_82_net65225, u5_mult_82_net65229,
         u5_mult_82_net65189, u5_mult_82_net65191, u5_mult_82_net65193,
         u5_mult_82_net65197, u5_mult_82_net64957, u5_mult_82_net64959,
         u5_mult_82_net64961, u5_mult_82_net64949, u5_mult_82_net64935,
         u5_mult_82_net64937, u5_mult_82_net64939, u5_mult_82_net64941,
         u5_mult_82_net64943, u5_mult_82_net64945, u5_mult_82_net64947,
         u5_mult_82_net64921, u5_mult_82_net64923, u5_mult_82_net64913,
         u5_mult_82_net64915, u5_mult_82_net64899, u5_mult_82_net64901,
         u5_mult_82_net64903, u5_mult_82_net64905, u5_mult_82_net64911,
         u5_mult_82_net64881, u5_mult_82_net64883, u5_mult_82_net64885,
         u5_mult_82_net64887, u5_mult_82_net64893, u5_mult_82_net64683,
         u5_mult_82_net64685, u5_mult_82_net64687, u5_mult_82_net64689,
         u5_mult_82_net64695, u5_mult_82_net64665, u5_mult_82_net64667,
         u5_mult_82_net64669, u5_mult_82_net64671, u5_mult_82_net64673,
         u5_mult_82_net64677, u5_mult_82_net64559, u5_mult_82_net64561,
         u5_mult_82_net64563, u5_mult_82_net64565, u5_mult_82_net64567,
         u5_mult_82_net64535, u5_mult_82_net64523, u5_mult_82_net64525,
         u5_mult_82_net64527, u5_mult_82_net64531, u5_mult_82_net64533,
         u5_mult_82_net64517, u5_mult_82_net64505, u5_mult_82_net64507,
         u5_mult_82_net64509, u5_mult_82_net64511, u5_mult_82_net64513,
         u5_mult_82_net64515, u5_mult_82_net64487, u5_mult_82_net64489,
         u5_mult_82_net64491, u5_mult_82_net64469, u5_mult_82_net64471,
         u5_mult_82_net64473, u5_mult_82_net64475, u5_mult_82_net64477,
         u5_mult_82_net64451, u5_mult_82_net64453, u5_mult_82_net64455,
         u5_mult_82_net64459, u5_mult_82_net64433, u5_mult_82_net64435,
         u5_mult_82_net64437, u5_mult_82_net64441, u5_mult_82_net64427,
         u5_mult_82_net64415, u5_mult_82_net64417, u5_mult_82_net64419,
         u5_mult_82_net64423, u5_mult_82_net64425, u5_mult_82_net64379,
         u5_mult_82_net64381, u5_mult_82_net64383, u5_mult_82_net64385,
         u5_mult_82_net64387, u5_mult_82_net64373, u5_mult_82_net64361,
         u5_mult_82_net64363, u5_mult_82_net64365, u5_mult_82_net64367,
         u5_mult_82_net64369, u5_mult_82_net64371, u5_mult_82_net64217,
         u5_mult_82_net64219, u5_mult_82_net64223, u5_mult_82_net64225,
         u5_mult_82_net57182, u5_mult_82_net57161, u5_mult_82_SUMB_43__18_,
         u5_mult_82_SUMB_43__19_, u5_mult_82_SUMB_43__20_,
         u5_mult_82_SUMB_43__21_, u5_mult_82_SUMB_43__22_,
         u5_mult_82_SUMB_43__23_, u5_mult_82_SUMB_43__24_,
         u5_mult_82_SUMB_43__25_, u5_mult_82_SUMB_43__26_,
         u5_mult_82_SUMB_43__27_, u5_mult_82_SUMB_43__28_,
         u5_mult_82_SUMB_43__29_, u5_mult_82_SUMB_43__30_,
         u5_mult_82_SUMB_43__31_, u5_mult_82_SUMB_43__32_,
         u5_mult_82_SUMB_43__33_, u5_mult_82_SUMB_43__34_,
         u5_mult_82_SUMB_43__35_, u5_mult_82_SUMB_43__36_,
         u5_mult_82_SUMB_43__37_, u5_mult_82_SUMB_43__38_,
         u5_mult_82_SUMB_43__39_, u5_mult_82_SUMB_43__40_,
         u5_mult_82_SUMB_43__41_, u5_mult_82_SUMB_43__42_,
         u5_mult_82_SUMB_43__43_, u5_mult_82_SUMB_43__44_,
         u5_mult_82_SUMB_43__45_, u5_mult_82_SUMB_43__46_,
         u5_mult_82_SUMB_43__47_, u5_mult_82_SUMB_43__48_,
         u5_mult_82_SUMB_43__49_, u5_mult_82_SUMB_43__50_,
         u5_mult_82_SUMB_43__51_, u5_mult_82_SUMB_44__1_,
         u5_mult_82_SUMB_44__2_, u5_mult_82_SUMB_44__3_,
         u5_mult_82_SUMB_44__4_, u5_mult_82_SUMB_44__5_,
         u5_mult_82_SUMB_44__6_, u5_mult_82_SUMB_44__7_,
         u5_mult_82_SUMB_44__8_, u5_mult_82_SUMB_44__9_,
         u5_mult_82_SUMB_44__11_, u5_mult_82_SUMB_44__12_,
         u5_mult_82_SUMB_44__13_, u5_mult_82_SUMB_44__14_,
         u5_mult_82_SUMB_44__15_, u5_mult_82_SUMB_44__16_,
         u5_mult_82_SUMB_44__17_, u5_mult_82_SUMB_44__18_,
         u5_mult_82_SUMB_44__19_, u5_mult_82_SUMB_44__20_,
         u5_mult_82_SUMB_44__21_, u5_mult_82_SUMB_44__22_,
         u5_mult_82_SUMB_44__23_, u5_mult_82_SUMB_44__24_,
         u5_mult_82_SUMB_44__25_, u5_mult_82_SUMB_44__26_,
         u5_mult_82_SUMB_44__27_, u5_mult_82_SUMB_44__28_,
         u5_mult_82_SUMB_44__29_, u5_mult_82_SUMB_44__30_,
         u5_mult_82_SUMB_44__31_, u5_mult_82_SUMB_44__32_,
         u5_mult_82_SUMB_44__33_, u5_mult_82_SUMB_44__34_,
         u5_mult_82_SUMB_44__35_, u5_mult_82_SUMB_44__36_,
         u5_mult_82_SUMB_44__37_, u5_mult_82_SUMB_44__38_,
         u5_mult_82_SUMB_44__39_, u5_mult_82_SUMB_44__40_,
         u5_mult_82_SUMB_44__41_, u5_mult_82_SUMB_44__42_,
         u5_mult_82_SUMB_44__43_, u5_mult_82_SUMB_44__44_,
         u5_mult_82_SUMB_44__45_, u5_mult_82_SUMB_44__46_,
         u5_mult_82_SUMB_44__47_, u5_mult_82_SUMB_44__48_,
         u5_mult_82_SUMB_44__49_, u5_mult_82_SUMB_44__50_,
         u5_mult_82_SUMB_44__51_, u5_mult_82_SUMB_45__1_,
         u5_mult_82_SUMB_45__2_, u5_mult_82_SUMB_45__3_,
         u5_mult_82_SUMB_45__4_, u5_mult_82_SUMB_45__5_,
         u5_mult_82_SUMB_45__6_, u5_mult_82_SUMB_45__7_,
         u5_mult_82_SUMB_45__8_, u5_mult_82_SUMB_45__9_,
         u5_mult_82_SUMB_45__10_, u5_mult_82_SUMB_45__11_,
         u5_mult_82_SUMB_45__12_, u5_mult_82_SUMB_45__13_,
         u5_mult_82_SUMB_45__14_, u5_mult_82_SUMB_45__15_,
         u5_mult_82_SUMB_45__16_, u5_mult_82_SUMB_45__17_,
         u5_mult_82_SUMB_45__18_, u5_mult_82_SUMB_45__19_,
         u5_mult_82_SUMB_45__20_, u5_mult_82_SUMB_45__21_,
         u5_mult_82_SUMB_45__22_, u5_mult_82_SUMB_45__23_,
         u5_mult_82_SUMB_45__24_, u5_mult_82_SUMB_45__25_,
         u5_mult_82_SUMB_45__26_, u5_mult_82_SUMB_45__27_,
         u5_mult_82_SUMB_45__28_, u5_mult_82_SUMB_45__29_,
         u5_mult_82_SUMB_45__30_, u5_mult_82_SUMB_45__31_,
         u5_mult_82_SUMB_45__32_, u5_mult_82_SUMB_45__33_,
         u5_mult_82_SUMB_45__34_, u5_mult_82_SUMB_45__35_,
         u5_mult_82_SUMB_45__36_, u5_mult_82_SUMB_45__37_,
         u5_mult_82_SUMB_45__38_, u5_mult_82_SUMB_45__39_,
         u5_mult_82_SUMB_45__40_, u5_mult_82_SUMB_45__41_,
         u5_mult_82_SUMB_45__42_, u5_mult_82_SUMB_45__43_,
         u5_mult_82_SUMB_45__44_, u5_mult_82_SUMB_45__45_,
         u5_mult_82_SUMB_45__46_, u5_mult_82_SUMB_45__47_,
         u5_mult_82_SUMB_45__48_, u5_mult_82_SUMB_45__49_,
         u5_mult_82_SUMB_45__50_, u5_mult_82_SUMB_45__51_,
         u5_mult_82_SUMB_46__1_, u5_mult_82_SUMB_46__2_,
         u5_mult_82_SUMB_46__3_, u5_mult_82_SUMB_46__4_,
         u5_mult_82_SUMB_46__5_, u5_mult_82_SUMB_46__6_,
         u5_mult_82_SUMB_46__7_, u5_mult_82_SUMB_46__8_,
         u5_mult_82_SUMB_46__10_, u5_mult_82_SUMB_46__11_,
         u5_mult_82_SUMB_46__12_, u5_mult_82_SUMB_46__13_,
         u5_mult_82_SUMB_46__14_, u5_mult_82_SUMB_46__15_,
         u5_mult_82_SUMB_46__16_, u5_mult_82_SUMB_46__17_,
         u5_mult_82_SUMB_46__18_, u5_mult_82_SUMB_46__19_,
         u5_mult_82_SUMB_46__20_, u5_mult_82_SUMB_46__21_,
         u5_mult_82_SUMB_46__22_, u5_mult_82_SUMB_46__23_,
         u5_mult_82_SUMB_46__24_, u5_mult_82_SUMB_46__25_,
         u5_mult_82_SUMB_46__26_, u5_mult_82_SUMB_46__27_,
         u5_mult_82_SUMB_46__28_, u5_mult_82_SUMB_46__29_,
         u5_mult_82_SUMB_46__30_, u5_mult_82_SUMB_46__31_,
         u5_mult_82_SUMB_46__32_, u5_mult_82_SUMB_46__33_,
         u5_mult_82_SUMB_46__34_, u5_mult_82_SUMB_46__35_,
         u5_mult_82_SUMB_46__36_, u5_mult_82_SUMB_46__37_,
         u5_mult_82_SUMB_46__38_, u5_mult_82_SUMB_46__39_,
         u5_mult_82_SUMB_46__40_, u5_mult_82_SUMB_46__41_,
         u5_mult_82_SUMB_46__42_, u5_mult_82_SUMB_46__43_,
         u5_mult_82_SUMB_46__44_, u5_mult_82_SUMB_46__45_,
         u5_mult_82_SUMB_46__46_, u5_mult_82_SUMB_46__47_,
         u5_mult_82_SUMB_46__48_, u5_mult_82_SUMB_46__49_,
         u5_mult_82_SUMB_46__50_, u5_mult_82_SUMB_46__51_,
         u5_mult_82_SUMB_47__1_, u5_mult_82_SUMB_47__2_,
         u5_mult_82_SUMB_47__3_, u5_mult_82_SUMB_47__4_,
         u5_mult_82_SUMB_47__5_, u5_mult_82_SUMB_47__6_,
         u5_mult_82_SUMB_47__7_, u5_mult_82_SUMB_47__9_,
         u5_mult_82_SUMB_47__10_, u5_mult_82_SUMB_47__11_,
         u5_mult_82_SUMB_47__12_, u5_mult_82_SUMB_47__13_,
         u5_mult_82_SUMB_47__14_, u5_mult_82_SUMB_47__15_,
         u5_mult_82_SUMB_47__16_, u5_mult_82_SUMB_47__17_,
         u5_mult_82_SUMB_47__18_, u5_mult_82_SUMB_47__19_,
         u5_mult_82_SUMB_47__20_, u5_mult_82_SUMB_47__21_,
         u5_mult_82_SUMB_47__22_, u5_mult_82_SUMB_47__23_,
         u5_mult_82_SUMB_47__24_, u5_mult_82_SUMB_47__25_,
         u5_mult_82_SUMB_47__26_, u5_mult_82_SUMB_47__27_,
         u5_mult_82_SUMB_47__28_, u5_mult_82_SUMB_47__29_,
         u5_mult_82_SUMB_47__30_, u5_mult_82_SUMB_47__31_,
         u5_mult_82_SUMB_47__32_, u5_mult_82_SUMB_47__33_,
         u5_mult_82_SUMB_47__34_, u5_mult_82_SUMB_47__35_,
         u5_mult_82_SUMB_47__37_, u5_mult_82_SUMB_47__38_,
         u5_mult_82_SUMB_47__39_, u5_mult_82_SUMB_47__40_,
         u5_mult_82_SUMB_47__41_, u5_mult_82_SUMB_47__42_,
         u5_mult_82_SUMB_47__43_, u5_mult_82_SUMB_47__44_,
         u5_mult_82_SUMB_47__45_, u5_mult_82_SUMB_47__46_,
         u5_mult_82_SUMB_47__47_, u5_mult_82_SUMB_47__48_,
         u5_mult_82_SUMB_47__49_, u5_mult_82_SUMB_47__50_,
         u5_mult_82_SUMB_47__51_, u5_mult_82_SUMB_48__1_,
         u5_mult_82_SUMB_48__2_, u5_mult_82_SUMB_48__3_,
         u5_mult_82_SUMB_48__4_, u5_mult_82_SUMB_48__5_,
         u5_mult_82_SUMB_48__6_, u5_mult_82_SUMB_48__7_,
         u5_mult_82_SUMB_48__9_, u5_mult_82_SUMB_48__10_,
         u5_mult_82_SUMB_48__11_, u5_mult_82_SUMB_48__12_,
         u5_mult_82_SUMB_48__13_, u5_mult_82_SUMB_48__14_,
         u5_mult_82_SUMB_48__16_, u5_mult_82_SUMB_48__17_,
         u5_mult_82_SUMB_48__18_, u5_mult_82_SUMB_48__19_,
         u5_mult_82_SUMB_48__20_, u5_mult_82_SUMB_48__21_,
         u5_mult_82_SUMB_48__22_, u5_mult_82_SUMB_48__23_,
         u5_mult_82_SUMB_48__24_, u5_mult_82_SUMB_48__25_,
         u5_mult_82_SUMB_48__26_, u5_mult_82_SUMB_48__27_,
         u5_mult_82_SUMB_48__28_, u5_mult_82_SUMB_48__29_,
         u5_mult_82_SUMB_48__30_, u5_mult_82_SUMB_48__31_,
         u5_mult_82_SUMB_48__32_, u5_mult_82_SUMB_48__33_,
         u5_mult_82_SUMB_48__34_, u5_mult_82_SUMB_48__35_,
         u5_mult_82_SUMB_48__36_, u5_mult_82_SUMB_48__37_,
         u5_mult_82_SUMB_48__38_, u5_mult_82_SUMB_48__39_,
         u5_mult_82_SUMB_48__40_, u5_mult_82_SUMB_48__41_,
         u5_mult_82_SUMB_48__42_, u5_mult_82_SUMB_48__43_,
         u5_mult_82_SUMB_48__44_, u5_mult_82_SUMB_48__45_,
         u5_mult_82_SUMB_48__46_, u5_mult_82_SUMB_48__47_,
         u5_mult_82_SUMB_48__48_, u5_mult_82_SUMB_48__49_,
         u5_mult_82_SUMB_48__50_, u5_mult_82_SUMB_48__51_,
         u5_mult_82_SUMB_49__1_, u5_mult_82_SUMB_49__2_,
         u5_mult_82_SUMB_49__3_, u5_mult_82_SUMB_49__4_,
         u5_mult_82_SUMB_49__5_, u5_mult_82_SUMB_49__8_,
         u5_mult_82_SUMB_49__9_, u5_mult_82_SUMB_49__10_,
         u5_mult_82_SUMB_49__11_, u5_mult_82_SUMB_49__12_,
         u5_mult_82_SUMB_49__13_, u5_mult_82_SUMB_49__14_,
         u5_mult_82_SUMB_49__15_, u5_mult_82_SUMB_49__16_,
         u5_mult_82_SUMB_49__17_, u5_mult_82_SUMB_49__18_,
         u5_mult_82_SUMB_49__19_, u5_mult_82_SUMB_49__20_,
         u5_mult_82_SUMB_49__21_, u5_mult_82_SUMB_49__22_,
         u5_mult_82_SUMB_49__23_, u5_mult_82_SUMB_49__24_,
         u5_mult_82_SUMB_49__25_, u5_mult_82_SUMB_49__26_,
         u5_mult_82_SUMB_49__27_, u5_mult_82_SUMB_49__28_,
         u5_mult_82_SUMB_49__29_, u5_mult_82_SUMB_49__30_,
         u5_mult_82_SUMB_49__31_, u5_mult_82_SUMB_49__32_,
         u5_mult_82_SUMB_49__33_, u5_mult_82_SUMB_49__34_,
         u5_mult_82_SUMB_49__35_, u5_mult_82_SUMB_49__36_,
         u5_mult_82_SUMB_49__37_, u5_mult_82_SUMB_49__38_,
         u5_mult_82_SUMB_49__39_, u5_mult_82_SUMB_49__40_,
         u5_mult_82_SUMB_49__41_, u5_mult_82_SUMB_49__42_,
         u5_mult_82_SUMB_49__43_, u5_mult_82_SUMB_49__44_,
         u5_mult_82_SUMB_49__45_, u5_mult_82_SUMB_49__46_,
         u5_mult_82_SUMB_49__47_, u5_mult_82_SUMB_49__48_,
         u5_mult_82_SUMB_49__49_, u5_mult_82_SUMB_49__50_,
         u5_mult_82_SUMB_49__51_, u5_mult_82_SUMB_50__1_,
         u5_mult_82_SUMB_50__2_, u5_mult_82_SUMB_50__3_,
         u5_mult_82_SUMB_50__4_, u5_mult_82_SUMB_50__8_,
         u5_mult_82_SUMB_50__9_, u5_mult_82_SUMB_50__10_,
         u5_mult_82_SUMB_50__11_, u5_mult_82_SUMB_50__12_,
         u5_mult_82_SUMB_50__13_, u5_mult_82_SUMB_50__14_,
         u5_mult_82_SUMB_50__15_, u5_mult_82_SUMB_50__16_,
         u5_mult_82_SUMB_50__17_, u5_mult_82_SUMB_50__18_,
         u5_mult_82_SUMB_50__19_, u5_mult_82_SUMB_50__20_,
         u5_mult_82_SUMB_50__21_, u5_mult_82_SUMB_50__22_,
         u5_mult_82_SUMB_50__23_, u5_mult_82_SUMB_50__24_,
         u5_mult_82_SUMB_50__25_, u5_mult_82_SUMB_50__26_,
         u5_mult_82_SUMB_50__27_, u5_mult_82_SUMB_50__28_,
         u5_mult_82_SUMB_50__29_, u5_mult_82_SUMB_50__30_,
         u5_mult_82_SUMB_50__31_, u5_mult_82_SUMB_50__32_,
         u5_mult_82_SUMB_50__33_, u5_mult_82_SUMB_50__34_,
         u5_mult_82_SUMB_50__35_, u5_mult_82_SUMB_50__36_,
         u5_mult_82_SUMB_50__37_, u5_mult_82_SUMB_50__38_,
         u5_mult_82_SUMB_50__39_, u5_mult_82_SUMB_50__40_,
         u5_mult_82_SUMB_50__41_, u5_mult_82_SUMB_50__42_,
         u5_mult_82_SUMB_50__43_, u5_mult_82_SUMB_50__44_,
         u5_mult_82_SUMB_50__45_, u5_mult_82_SUMB_50__46_,
         u5_mult_82_SUMB_50__47_, u5_mult_82_SUMB_50__48_,
         u5_mult_82_SUMB_50__49_, u5_mult_82_SUMB_50__50_,
         u5_mult_82_SUMB_50__51_, u5_mult_82_SUMB_51__1_,
         u5_mult_82_SUMB_51__2_, u5_mult_82_SUMB_51__3_,
         u5_mult_82_SUMB_51__4_, u5_mult_82_SUMB_51__7_,
         u5_mult_82_SUMB_51__8_, u5_mult_82_SUMB_51__9_,
         u5_mult_82_SUMB_51__10_, u5_mult_82_SUMB_51__11_,
         u5_mult_82_SUMB_51__12_, u5_mult_82_SUMB_51__13_,
         u5_mult_82_SUMB_51__14_, u5_mult_82_SUMB_51__15_,
         u5_mult_82_SUMB_51__16_, u5_mult_82_SUMB_51__17_,
         u5_mult_82_SUMB_51__18_, u5_mult_82_SUMB_51__19_,
         u5_mult_82_SUMB_51__20_, u5_mult_82_SUMB_51__21_,
         u5_mult_82_SUMB_51__22_, u5_mult_82_SUMB_51__23_,
         u5_mult_82_SUMB_51__24_, u5_mult_82_SUMB_51__25_,
         u5_mult_82_SUMB_51__26_, u5_mult_82_SUMB_51__27_,
         u5_mult_82_SUMB_51__28_, u5_mult_82_SUMB_51__29_,
         u5_mult_82_SUMB_51__30_, u5_mult_82_SUMB_51__31_,
         u5_mult_82_SUMB_51__32_, u5_mult_82_SUMB_51__33_,
         u5_mult_82_SUMB_51__34_, u5_mult_82_SUMB_51__35_,
         u5_mult_82_SUMB_51__36_, u5_mult_82_SUMB_51__37_,
         u5_mult_82_SUMB_51__38_, u5_mult_82_SUMB_51__39_,
         u5_mult_82_SUMB_51__40_, u5_mult_82_SUMB_51__41_,
         u5_mult_82_SUMB_51__42_, u5_mult_82_SUMB_51__43_,
         u5_mult_82_SUMB_51__44_, u5_mult_82_SUMB_51__45_,
         u5_mult_82_SUMB_51__46_, u5_mult_82_SUMB_51__47_,
         u5_mult_82_SUMB_51__48_, u5_mult_82_SUMB_51__49_,
         u5_mult_82_SUMB_51__50_, u5_mult_82_SUMB_51__51_,
         u5_mult_82_SUMB_52__1_, u5_mult_82_SUMB_52__2_,
         u5_mult_82_SUMB_52__3_, u5_mult_82_SUMB_52__4_,
         u5_mult_82_SUMB_52__6_, u5_mult_82_SUMB_52__7_,
         u5_mult_82_SUMB_52__8_, u5_mult_82_SUMB_52__9_,
         u5_mult_82_SUMB_52__10_, u5_mult_82_SUMB_52__11_,
         u5_mult_82_SUMB_52__12_, u5_mult_82_SUMB_52__13_,
         u5_mult_82_SUMB_52__14_, u5_mult_82_SUMB_52__15_,
         u5_mult_82_SUMB_52__16_, u5_mult_82_SUMB_52__17_,
         u5_mult_82_SUMB_52__18_, u5_mult_82_SUMB_52__19_,
         u5_mult_82_SUMB_52__20_, u5_mult_82_SUMB_52__21_,
         u5_mult_82_SUMB_52__22_, u5_mult_82_SUMB_52__23_,
         u5_mult_82_SUMB_52__24_, u5_mult_82_SUMB_52__25_,
         u5_mult_82_SUMB_52__26_, u5_mult_82_SUMB_52__27_,
         u5_mult_82_SUMB_52__28_, u5_mult_82_SUMB_52__29_,
         u5_mult_82_SUMB_52__30_, u5_mult_82_SUMB_52__31_,
         u5_mult_82_SUMB_52__32_, u5_mult_82_SUMB_52__33_,
         u5_mult_82_SUMB_52__34_, u5_mult_82_SUMB_52__35_,
         u5_mult_82_SUMB_52__36_, u5_mult_82_SUMB_52__37_,
         u5_mult_82_SUMB_52__38_, u5_mult_82_SUMB_52__39_,
         u5_mult_82_SUMB_52__40_, u5_mult_82_SUMB_52__41_,
         u5_mult_82_SUMB_52__42_, u5_mult_82_SUMB_52__43_,
         u5_mult_82_SUMB_52__44_, u5_mult_82_SUMB_52__45_,
         u5_mult_82_SUMB_52__46_, u5_mult_82_SUMB_52__47_,
         u5_mult_82_SUMB_52__48_, u5_mult_82_SUMB_52__49_,
         u5_mult_82_SUMB_52__50_, u5_mult_82_SUMB_52__51_,
         u5_mult_82_CARRYB_43__18_, u5_mult_82_CARRYB_43__19_,
         u5_mult_82_CARRYB_43__20_, u5_mult_82_CARRYB_43__21_,
         u5_mult_82_CARRYB_43__22_, u5_mult_82_CARRYB_43__23_,
         u5_mult_82_CARRYB_43__24_, u5_mult_82_CARRYB_43__25_,
         u5_mult_82_CARRYB_43__26_, u5_mult_82_CARRYB_43__27_,
         u5_mult_82_CARRYB_43__28_, u5_mult_82_CARRYB_43__29_,
         u5_mult_82_CARRYB_43__30_, u5_mult_82_CARRYB_43__31_,
         u5_mult_82_CARRYB_43__32_, u5_mult_82_CARRYB_43__33_,
         u5_mult_82_CARRYB_43__34_, u5_mult_82_CARRYB_43__35_,
         u5_mult_82_CARRYB_43__36_, u5_mult_82_CARRYB_43__37_,
         u5_mult_82_CARRYB_43__38_, u5_mult_82_CARRYB_43__39_,
         u5_mult_82_CARRYB_43__40_, u5_mult_82_CARRYB_43__41_,
         u5_mult_82_CARRYB_43__42_, u5_mult_82_CARRYB_43__43_,
         u5_mult_82_CARRYB_43__44_, u5_mult_82_CARRYB_43__45_,
         u5_mult_82_CARRYB_43__46_, u5_mult_82_CARRYB_43__47_,
         u5_mult_82_CARRYB_43__48_, u5_mult_82_CARRYB_43__49_,
         u5_mult_82_CARRYB_43__50_, u5_mult_82_CARRYB_43__51_,
         u5_mult_82_CARRYB_44__0_, u5_mult_82_CARRYB_44__1_,
         u5_mult_82_CARRYB_44__2_, u5_mult_82_CARRYB_44__3_,
         u5_mult_82_CARRYB_44__4_, u5_mult_82_CARRYB_44__5_,
         u5_mult_82_CARRYB_44__6_, u5_mult_82_CARRYB_44__7_,
         u5_mult_82_CARRYB_44__8_, u5_mult_82_CARRYB_44__10_,
         u5_mult_82_CARRYB_44__11_, u5_mult_82_CARRYB_44__12_,
         u5_mult_82_CARRYB_44__13_, u5_mult_82_CARRYB_44__14_,
         u5_mult_82_CARRYB_44__15_, u5_mult_82_CARRYB_44__16_,
         u5_mult_82_CARRYB_44__17_, u5_mult_82_CARRYB_44__18_,
         u5_mult_82_CARRYB_44__19_, u5_mult_82_CARRYB_44__20_,
         u5_mult_82_CARRYB_44__21_, u5_mult_82_CARRYB_44__22_,
         u5_mult_82_CARRYB_44__23_, u5_mult_82_CARRYB_44__24_,
         u5_mult_82_CARRYB_44__25_, u5_mult_82_CARRYB_44__26_,
         u5_mult_82_CARRYB_44__27_, u5_mult_82_CARRYB_44__28_,
         u5_mult_82_CARRYB_44__29_, u5_mult_82_CARRYB_44__30_,
         u5_mult_82_CARRYB_44__31_, u5_mult_82_CARRYB_44__32_,
         u5_mult_82_CARRYB_44__33_, u5_mult_82_CARRYB_44__34_,
         u5_mult_82_CARRYB_44__35_, u5_mult_82_CARRYB_44__36_,
         u5_mult_82_CARRYB_44__37_, u5_mult_82_CARRYB_44__38_,
         u5_mult_82_CARRYB_44__39_, u5_mult_82_CARRYB_44__40_,
         u5_mult_82_CARRYB_44__41_, u5_mult_82_CARRYB_44__42_,
         u5_mult_82_CARRYB_44__43_, u5_mult_82_CARRYB_44__44_,
         u5_mult_82_CARRYB_44__45_, u5_mult_82_CARRYB_44__46_,
         u5_mult_82_CARRYB_44__47_, u5_mult_82_CARRYB_44__48_,
         u5_mult_82_CARRYB_44__49_, u5_mult_82_CARRYB_44__50_,
         u5_mult_82_CARRYB_44__51_, u5_mult_82_CARRYB_45__0_,
         u5_mult_82_CARRYB_45__1_, u5_mult_82_CARRYB_45__2_,
         u5_mult_82_CARRYB_45__3_, u5_mult_82_CARRYB_45__4_,
         u5_mult_82_CARRYB_45__5_, u5_mult_82_CARRYB_45__6_,
         u5_mult_82_CARRYB_45__7_, u5_mult_82_CARRYB_45__8_,
         u5_mult_82_CARRYB_45__10_, u5_mult_82_CARRYB_45__11_,
         u5_mult_82_CARRYB_45__12_, u5_mult_82_CARRYB_45__13_,
         u5_mult_82_CARRYB_45__14_, u5_mult_82_CARRYB_45__15_,
         u5_mult_82_CARRYB_45__16_, u5_mult_82_CARRYB_45__17_,
         u5_mult_82_CARRYB_45__18_, u5_mult_82_CARRYB_45__19_,
         u5_mult_82_CARRYB_45__20_, u5_mult_82_CARRYB_45__21_,
         u5_mult_82_CARRYB_45__22_, u5_mult_82_CARRYB_45__23_,
         u5_mult_82_CARRYB_45__24_, u5_mult_82_CARRYB_45__25_,
         u5_mult_82_CARRYB_45__26_, u5_mult_82_CARRYB_45__27_,
         u5_mult_82_CARRYB_45__28_, u5_mult_82_CARRYB_45__29_,
         u5_mult_82_CARRYB_45__30_, u5_mult_82_CARRYB_45__31_,
         u5_mult_82_CARRYB_45__32_, u5_mult_82_CARRYB_45__33_,
         u5_mult_82_CARRYB_45__34_, u5_mult_82_CARRYB_45__35_,
         u5_mult_82_CARRYB_45__36_, u5_mult_82_CARRYB_45__37_,
         u5_mult_82_CARRYB_45__38_, u5_mult_82_CARRYB_45__39_,
         u5_mult_82_CARRYB_45__40_, u5_mult_82_CARRYB_45__41_,
         u5_mult_82_CARRYB_45__42_, u5_mult_82_CARRYB_45__43_,
         u5_mult_82_CARRYB_45__44_, u5_mult_82_CARRYB_45__45_,
         u5_mult_82_CARRYB_45__46_, u5_mult_82_CARRYB_45__47_,
         u5_mult_82_CARRYB_45__48_, u5_mult_82_CARRYB_45__49_,
         u5_mult_82_CARRYB_45__50_, u5_mult_82_CARRYB_45__51_,
         u5_mult_82_CARRYB_46__0_, u5_mult_82_CARRYB_46__1_,
         u5_mult_82_CARRYB_46__2_, u5_mult_82_CARRYB_46__3_,
         u5_mult_82_CARRYB_46__4_, u5_mult_82_CARRYB_46__5_,
         u5_mult_82_CARRYB_46__6_, u5_mult_82_CARRYB_46__7_,
         u5_mult_82_CARRYB_46__9_, u5_mult_82_CARRYB_46__10_,
         u5_mult_82_CARRYB_46__11_, u5_mult_82_CARRYB_46__12_,
         u5_mult_82_CARRYB_46__13_, u5_mult_82_CARRYB_46__14_,
         u5_mult_82_CARRYB_46__15_, u5_mult_82_CARRYB_46__16_,
         u5_mult_82_CARRYB_46__17_, u5_mult_82_CARRYB_46__18_,
         u5_mult_82_CARRYB_46__19_, u5_mult_82_CARRYB_46__20_,
         u5_mult_82_CARRYB_46__21_, u5_mult_82_CARRYB_46__22_,
         u5_mult_82_CARRYB_46__23_, u5_mult_82_CARRYB_46__24_,
         u5_mult_82_CARRYB_46__25_, u5_mult_82_CARRYB_46__26_,
         u5_mult_82_CARRYB_46__27_, u5_mult_82_CARRYB_46__28_,
         u5_mult_82_CARRYB_46__29_, u5_mult_82_CARRYB_46__30_,
         u5_mult_82_CARRYB_46__31_, u5_mult_82_CARRYB_46__32_,
         u5_mult_82_CARRYB_46__33_, u5_mult_82_CARRYB_46__34_,
         u5_mult_82_CARRYB_46__35_, u5_mult_82_CARRYB_46__36_,
         u5_mult_82_CARRYB_46__37_, u5_mult_82_CARRYB_46__38_,
         u5_mult_82_CARRYB_46__39_, u5_mult_82_CARRYB_46__40_,
         u5_mult_82_CARRYB_46__41_, u5_mult_82_CARRYB_46__42_,
         u5_mult_82_CARRYB_46__43_, u5_mult_82_CARRYB_46__44_,
         u5_mult_82_CARRYB_46__45_, u5_mult_82_CARRYB_46__46_,
         u5_mult_82_CARRYB_46__47_, u5_mult_82_CARRYB_46__48_,
         u5_mult_82_CARRYB_46__49_, u5_mult_82_CARRYB_46__50_,
         u5_mult_82_CARRYB_46__51_, u5_mult_82_CARRYB_47__0_,
         u5_mult_82_CARRYB_47__1_, u5_mult_82_CARRYB_47__2_,
         u5_mult_82_CARRYB_47__3_, u5_mult_82_CARRYB_47__4_,
         u5_mult_82_CARRYB_47__5_, u5_mult_82_CARRYB_47__6_,
         u5_mult_82_CARRYB_47__7_, u5_mult_82_CARRYB_47__9_,
         u5_mult_82_CARRYB_47__10_, u5_mult_82_CARRYB_47__11_,
         u5_mult_82_CARRYB_47__12_, u5_mult_82_CARRYB_47__13_,
         u5_mult_82_CARRYB_47__14_, u5_mult_82_CARRYB_47__15_,
         u5_mult_82_CARRYB_47__16_, u5_mult_82_CARRYB_47__17_,
         u5_mult_82_CARRYB_47__18_, u5_mult_82_CARRYB_47__19_,
         u5_mult_82_CARRYB_47__20_, u5_mult_82_CARRYB_47__21_,
         u5_mult_82_CARRYB_47__22_, u5_mult_82_CARRYB_47__23_,
         u5_mult_82_CARRYB_47__24_, u5_mult_82_CARRYB_47__25_,
         u5_mult_82_CARRYB_47__26_, u5_mult_82_CARRYB_47__27_,
         u5_mult_82_CARRYB_47__28_, u5_mult_82_CARRYB_47__29_,
         u5_mult_82_CARRYB_47__30_, u5_mult_82_CARRYB_47__31_,
         u5_mult_82_CARRYB_47__32_, u5_mult_82_CARRYB_47__33_,
         u5_mult_82_CARRYB_47__34_, u5_mult_82_CARRYB_47__35_,
         u5_mult_82_CARRYB_47__36_, u5_mult_82_CARRYB_47__37_,
         u5_mult_82_CARRYB_47__38_, u5_mult_82_CARRYB_47__39_,
         u5_mult_82_CARRYB_47__40_, u5_mult_82_CARRYB_47__41_,
         u5_mult_82_CARRYB_47__42_, u5_mult_82_CARRYB_47__43_,
         u5_mult_82_CARRYB_47__44_, u5_mult_82_CARRYB_47__45_,
         u5_mult_82_CARRYB_47__46_, u5_mult_82_CARRYB_47__47_,
         u5_mult_82_CARRYB_47__48_, u5_mult_82_CARRYB_47__49_,
         u5_mult_82_CARRYB_47__50_, u5_mult_82_CARRYB_47__51_,
         u5_mult_82_CARRYB_48__0_, u5_mult_82_CARRYB_48__1_,
         u5_mult_82_CARRYB_48__2_, u5_mult_82_CARRYB_48__3_,
         u5_mult_82_CARRYB_48__4_, u5_mult_82_CARRYB_48__5_,
         u5_mult_82_CARRYB_48__6_, u5_mult_82_CARRYB_48__8_,
         u5_mult_82_CARRYB_48__9_, u5_mult_82_CARRYB_48__10_,
         u5_mult_82_CARRYB_48__11_, u5_mult_82_CARRYB_48__12_,
         u5_mult_82_CARRYB_48__13_, u5_mult_82_CARRYB_48__14_,
         u5_mult_82_CARRYB_48__15_, u5_mult_82_CARRYB_48__16_,
         u5_mult_82_CARRYB_48__17_, u5_mult_82_CARRYB_48__18_,
         u5_mult_82_CARRYB_48__19_, u5_mult_82_CARRYB_48__20_,
         u5_mult_82_CARRYB_48__21_, u5_mult_82_CARRYB_48__22_,
         u5_mult_82_CARRYB_48__23_, u5_mult_82_CARRYB_48__24_,
         u5_mult_82_CARRYB_48__25_, u5_mult_82_CARRYB_48__26_,
         u5_mult_82_CARRYB_48__27_, u5_mult_82_CARRYB_48__28_,
         u5_mult_82_CARRYB_48__29_, u5_mult_82_CARRYB_48__30_,
         u5_mult_82_CARRYB_48__31_, u5_mult_82_CARRYB_48__32_,
         u5_mult_82_CARRYB_48__33_, u5_mult_82_CARRYB_48__34_,
         u5_mult_82_CARRYB_48__35_, u5_mult_82_CARRYB_48__36_,
         u5_mult_82_CARRYB_48__37_, u5_mult_82_CARRYB_48__38_,
         u5_mult_82_CARRYB_48__39_, u5_mult_82_CARRYB_48__40_,
         u5_mult_82_CARRYB_48__41_, u5_mult_82_CARRYB_48__42_,
         u5_mult_82_CARRYB_48__43_, u5_mult_82_CARRYB_48__44_,
         u5_mult_82_CARRYB_48__45_, u5_mult_82_CARRYB_48__46_,
         u5_mult_82_CARRYB_48__47_, u5_mult_82_CARRYB_48__48_,
         u5_mult_82_CARRYB_48__49_, u5_mult_82_CARRYB_48__50_,
         u5_mult_82_CARRYB_48__51_, u5_mult_82_CARRYB_49__0_,
         u5_mult_82_CARRYB_49__1_, u5_mult_82_CARRYB_49__2_,
         u5_mult_82_CARRYB_49__3_, u5_mult_82_CARRYB_49__4_,
         u5_mult_82_CARRYB_49__5_, u5_mult_82_CARRYB_49__7_,
         u5_mult_82_CARRYB_49__8_, u5_mult_82_CARRYB_49__9_,
         u5_mult_82_CARRYB_49__10_, u5_mult_82_CARRYB_49__11_,
         u5_mult_82_CARRYB_49__12_, u5_mult_82_CARRYB_49__14_,
         u5_mult_82_CARRYB_49__15_, u5_mult_82_CARRYB_49__16_,
         u5_mult_82_CARRYB_49__17_, u5_mult_82_CARRYB_49__18_,
         u5_mult_82_CARRYB_49__19_, u5_mult_82_CARRYB_49__20_,
         u5_mult_82_CARRYB_49__21_, u5_mult_82_CARRYB_49__22_,
         u5_mult_82_CARRYB_49__23_, u5_mult_82_CARRYB_49__24_,
         u5_mult_82_CARRYB_49__25_, u5_mult_82_CARRYB_49__26_,
         u5_mult_82_CARRYB_49__27_, u5_mult_82_CARRYB_49__28_,
         u5_mult_82_CARRYB_49__29_, u5_mult_82_CARRYB_49__30_,
         u5_mult_82_CARRYB_49__31_, u5_mult_82_CARRYB_49__32_,
         u5_mult_82_CARRYB_49__33_, u5_mult_82_CARRYB_49__34_,
         u5_mult_82_CARRYB_49__35_, u5_mult_82_CARRYB_49__36_,
         u5_mult_82_CARRYB_49__37_, u5_mult_82_CARRYB_49__38_,
         u5_mult_82_CARRYB_49__39_, u5_mult_82_CARRYB_49__40_,
         u5_mult_82_CARRYB_49__41_, u5_mult_82_CARRYB_49__42_,
         u5_mult_82_CARRYB_49__43_, u5_mult_82_CARRYB_49__44_,
         u5_mult_82_CARRYB_49__45_, u5_mult_82_CARRYB_49__46_,
         u5_mult_82_CARRYB_49__47_, u5_mult_82_CARRYB_49__48_,
         u5_mult_82_CARRYB_49__49_, u5_mult_82_CARRYB_49__50_,
         u5_mult_82_CARRYB_49__51_, u5_mult_82_CARRYB_50__0_,
         u5_mult_82_CARRYB_50__1_, u5_mult_82_CARRYB_50__2_,
         u5_mult_82_CARRYB_50__3_, u5_mult_82_CARRYB_50__4_,
         u5_mult_82_CARRYB_50__7_, u5_mult_82_CARRYB_50__8_,
         u5_mult_82_CARRYB_50__9_, u5_mult_82_CARRYB_50__10_,
         u5_mult_82_CARRYB_50__11_, u5_mult_82_CARRYB_50__12_,
         u5_mult_82_CARRYB_50__13_, u5_mult_82_CARRYB_50__14_,
         u5_mult_82_CARRYB_50__15_, u5_mult_82_CARRYB_50__16_,
         u5_mult_82_CARRYB_50__17_, u5_mult_82_CARRYB_50__18_,
         u5_mult_82_CARRYB_50__19_, u5_mult_82_CARRYB_50__20_,
         u5_mult_82_CARRYB_50__21_, u5_mult_82_CARRYB_50__22_,
         u5_mult_82_CARRYB_50__23_, u5_mult_82_CARRYB_50__24_,
         u5_mult_82_CARRYB_50__25_, u5_mult_82_CARRYB_50__26_,
         u5_mult_82_CARRYB_50__27_, u5_mult_82_CARRYB_50__28_,
         u5_mult_82_CARRYB_50__29_, u5_mult_82_CARRYB_50__30_,
         u5_mult_82_CARRYB_50__31_, u5_mult_82_CARRYB_50__32_,
         u5_mult_82_CARRYB_50__33_, u5_mult_82_CARRYB_50__34_,
         u5_mult_82_CARRYB_50__35_, u5_mult_82_CARRYB_50__36_,
         u5_mult_82_CARRYB_50__37_, u5_mult_82_CARRYB_50__38_,
         u5_mult_82_CARRYB_50__39_, u5_mult_82_CARRYB_50__40_,
         u5_mult_82_CARRYB_50__41_, u5_mult_82_CARRYB_50__42_,
         u5_mult_82_CARRYB_50__43_, u5_mult_82_CARRYB_50__44_,
         u5_mult_82_CARRYB_50__45_, u5_mult_82_CARRYB_50__46_,
         u5_mult_82_CARRYB_50__47_, u5_mult_82_CARRYB_50__48_,
         u5_mult_82_CARRYB_50__49_, u5_mult_82_CARRYB_50__50_,
         u5_mult_82_CARRYB_50__51_, u5_mult_82_CARRYB_51__0_,
         u5_mult_82_CARRYB_51__1_, u5_mult_82_CARRYB_51__2_,
         u5_mult_82_CARRYB_51__3_, u5_mult_82_CARRYB_51__6_,
         u5_mult_82_CARRYB_51__7_, u5_mult_82_CARRYB_51__8_,
         u5_mult_82_CARRYB_51__9_, u5_mult_82_CARRYB_51__10_,
         u5_mult_82_CARRYB_51__11_, u5_mult_82_CARRYB_51__12_,
         u5_mult_82_CARRYB_51__13_, u5_mult_82_CARRYB_51__14_,
         u5_mult_82_CARRYB_51__15_, u5_mult_82_CARRYB_51__16_,
         u5_mult_82_CARRYB_51__17_, u5_mult_82_CARRYB_51__18_,
         u5_mult_82_CARRYB_51__19_, u5_mult_82_CARRYB_51__20_,
         u5_mult_82_CARRYB_51__21_, u5_mult_82_CARRYB_51__22_,
         u5_mult_82_CARRYB_51__23_, u5_mult_82_CARRYB_51__24_,
         u5_mult_82_CARRYB_51__25_, u5_mult_82_CARRYB_51__26_,
         u5_mult_82_CARRYB_51__27_, u5_mult_82_CARRYB_51__28_,
         u5_mult_82_CARRYB_51__29_, u5_mult_82_CARRYB_51__30_,
         u5_mult_82_CARRYB_51__31_, u5_mult_82_CARRYB_51__32_,
         u5_mult_82_CARRYB_51__33_, u5_mult_82_CARRYB_51__34_,
         u5_mult_82_CARRYB_51__35_, u5_mult_82_CARRYB_51__36_,
         u5_mult_82_CARRYB_51__37_, u5_mult_82_CARRYB_51__38_,
         u5_mult_82_CARRYB_51__39_, u5_mult_82_CARRYB_51__40_,
         u5_mult_82_CARRYB_51__41_, u5_mult_82_CARRYB_51__42_,
         u5_mult_82_CARRYB_51__43_, u5_mult_82_CARRYB_51__44_,
         u5_mult_82_CARRYB_51__45_, u5_mult_82_CARRYB_51__46_,
         u5_mult_82_CARRYB_51__47_, u5_mult_82_CARRYB_51__48_,
         u5_mult_82_CARRYB_51__49_, u5_mult_82_CARRYB_51__50_,
         u5_mult_82_CARRYB_51__51_, u5_mult_82_CARRYB_52__0_,
         u5_mult_82_CARRYB_52__1_, u5_mult_82_CARRYB_52__2_,
         u5_mult_82_CARRYB_52__3_, u5_mult_82_CARRYB_52__5_,
         u5_mult_82_CARRYB_52__6_, u5_mult_82_CARRYB_52__7_,
         u5_mult_82_CARRYB_52__8_, u5_mult_82_CARRYB_52__9_,
         u5_mult_82_CARRYB_52__10_, u5_mult_82_CARRYB_52__11_,
         u5_mult_82_CARRYB_52__12_, u5_mult_82_CARRYB_52__13_,
         u5_mult_82_CARRYB_52__14_, u5_mult_82_CARRYB_52__15_,
         u5_mult_82_CARRYB_52__16_, u5_mult_82_CARRYB_52__17_,
         u5_mult_82_CARRYB_52__18_, u5_mult_82_CARRYB_52__19_,
         u5_mult_82_CARRYB_52__20_, u5_mult_82_CARRYB_52__21_,
         u5_mult_82_CARRYB_52__22_, u5_mult_82_CARRYB_52__23_,
         u5_mult_82_CARRYB_52__24_, u5_mult_82_CARRYB_52__25_,
         u5_mult_82_CARRYB_52__26_, u5_mult_82_CARRYB_52__27_,
         u5_mult_82_CARRYB_52__28_, u5_mult_82_CARRYB_52__29_,
         u5_mult_82_CARRYB_52__30_, u5_mult_82_CARRYB_52__31_,
         u5_mult_82_CARRYB_52__32_, u5_mult_82_CARRYB_52__33_,
         u5_mult_82_CARRYB_52__34_, u5_mult_82_CARRYB_52__35_,
         u5_mult_82_CARRYB_52__36_, u5_mult_82_CARRYB_52__37_,
         u5_mult_82_CARRYB_52__38_, u5_mult_82_CARRYB_52__39_,
         u5_mult_82_CARRYB_52__40_, u5_mult_82_CARRYB_52__41_,
         u5_mult_82_CARRYB_52__42_, u5_mult_82_CARRYB_52__43_,
         u5_mult_82_CARRYB_52__44_, u5_mult_82_CARRYB_52__45_,
         u5_mult_82_CARRYB_52__46_, u5_mult_82_CARRYB_52__47_,
         u5_mult_82_CARRYB_52__48_, u5_mult_82_CARRYB_52__49_,
         u5_mult_82_CARRYB_52__50_, u5_mult_82_CARRYB_52__51_,
         u5_mult_82_SUMB_33__36_, u5_mult_82_SUMB_33__37_,
         u5_mult_82_SUMB_33__38_, u5_mult_82_SUMB_33__39_,
         u5_mult_82_SUMB_33__40_, u5_mult_82_SUMB_33__41_,
         u5_mult_82_SUMB_33__42_, u5_mult_82_SUMB_33__43_,
         u5_mult_82_SUMB_33__44_, u5_mult_82_SUMB_33__45_,
         u5_mult_82_SUMB_33__46_, u5_mult_82_SUMB_33__47_,
         u5_mult_82_SUMB_33__48_, u5_mult_82_SUMB_33__49_,
         u5_mult_82_SUMB_33__50_, u5_mult_82_SUMB_33__51_,
         u5_mult_82_SUMB_34__1_, u5_mult_82_SUMB_34__2_,
         u5_mult_82_SUMB_34__3_, u5_mult_82_SUMB_34__4_,
         u5_mult_82_SUMB_34__5_, u5_mult_82_SUMB_34__6_,
         u5_mult_82_SUMB_34__7_, u5_mult_82_SUMB_34__8_,
         u5_mult_82_SUMB_34__9_, u5_mult_82_SUMB_34__10_,
         u5_mult_82_SUMB_34__11_, u5_mult_82_SUMB_34__12_,
         u5_mult_82_SUMB_34__13_, u5_mult_82_SUMB_34__14_,
         u5_mult_82_SUMB_34__15_, u5_mult_82_SUMB_34__17_,
         u5_mult_82_SUMB_34__18_, u5_mult_82_SUMB_34__19_,
         u5_mult_82_SUMB_34__20_, u5_mult_82_SUMB_34__21_,
         u5_mult_82_SUMB_34__22_, u5_mult_82_SUMB_34__23_,
         u5_mult_82_SUMB_34__24_, u5_mult_82_SUMB_34__25_,
         u5_mult_82_SUMB_34__26_, u5_mult_82_SUMB_34__27_,
         u5_mult_82_SUMB_34__28_, u5_mult_82_SUMB_34__29_,
         u5_mult_82_SUMB_34__30_, u5_mult_82_SUMB_34__31_,
         u5_mult_82_SUMB_34__32_, u5_mult_82_SUMB_34__33_,
         u5_mult_82_SUMB_34__34_, u5_mult_82_SUMB_34__35_,
         u5_mult_82_SUMB_34__36_, u5_mult_82_SUMB_34__37_,
         u5_mult_82_SUMB_34__38_, u5_mult_82_SUMB_34__39_,
         u5_mult_82_SUMB_34__40_, u5_mult_82_SUMB_34__41_,
         u5_mult_82_SUMB_34__42_, u5_mult_82_SUMB_34__43_,
         u5_mult_82_SUMB_34__44_, u5_mult_82_SUMB_34__45_,
         u5_mult_82_SUMB_34__46_, u5_mult_82_SUMB_34__47_,
         u5_mult_82_SUMB_34__48_, u5_mult_82_SUMB_34__49_,
         u5_mult_82_SUMB_34__50_, u5_mult_82_SUMB_34__51_,
         u5_mult_82_SUMB_35__1_, u5_mult_82_SUMB_35__2_,
         u5_mult_82_SUMB_35__3_, u5_mult_82_SUMB_35__4_,
         u5_mult_82_SUMB_35__5_, u5_mult_82_SUMB_35__6_,
         u5_mult_82_SUMB_35__7_, u5_mult_82_SUMB_35__8_,
         u5_mult_82_SUMB_35__9_, u5_mult_82_SUMB_35__10_,
         u5_mult_82_SUMB_35__11_, u5_mult_82_SUMB_35__12_,
         u5_mult_82_SUMB_35__13_, u5_mult_82_SUMB_35__14_,
         u5_mult_82_SUMB_35__17_, u5_mult_82_SUMB_35__18_,
         u5_mult_82_SUMB_35__19_, u5_mult_82_SUMB_35__20_,
         u5_mult_82_SUMB_35__21_, u5_mult_82_SUMB_35__22_,
         u5_mult_82_SUMB_35__23_, u5_mult_82_SUMB_35__24_,
         u5_mult_82_SUMB_35__25_, u5_mult_82_SUMB_35__26_,
         u5_mult_82_SUMB_35__27_, u5_mult_82_SUMB_35__28_,
         u5_mult_82_SUMB_35__29_, u5_mult_82_SUMB_35__30_,
         u5_mult_82_SUMB_35__31_, u5_mult_82_SUMB_35__32_,
         u5_mult_82_SUMB_35__33_, u5_mult_82_SUMB_35__34_,
         u5_mult_82_SUMB_35__35_, u5_mult_82_SUMB_35__36_,
         u5_mult_82_SUMB_35__37_, u5_mult_82_SUMB_35__38_,
         u5_mult_82_SUMB_35__39_, u5_mult_82_SUMB_35__40_,
         u5_mult_82_SUMB_35__41_, u5_mult_82_SUMB_35__42_,
         u5_mult_82_SUMB_35__43_, u5_mult_82_SUMB_35__44_,
         u5_mult_82_SUMB_35__45_, u5_mult_82_SUMB_35__46_,
         u5_mult_82_SUMB_35__47_, u5_mult_82_SUMB_35__48_,
         u5_mult_82_SUMB_35__49_, u5_mult_82_SUMB_35__50_,
         u5_mult_82_SUMB_35__51_, u5_mult_82_SUMB_36__1_,
         u5_mult_82_SUMB_36__2_, u5_mult_82_SUMB_36__3_,
         u5_mult_82_SUMB_36__4_, u5_mult_82_SUMB_36__5_,
         u5_mult_82_SUMB_36__6_, u5_mult_82_SUMB_36__7_,
         u5_mult_82_SUMB_36__8_, u5_mult_82_SUMB_36__9_,
         u5_mult_82_SUMB_36__10_, u5_mult_82_SUMB_36__11_,
         u5_mult_82_SUMB_36__12_, u5_mult_82_SUMB_36__13_,
         u5_mult_82_SUMB_36__16_, u5_mult_82_SUMB_36__17_,
         u5_mult_82_SUMB_36__18_, u5_mult_82_SUMB_36__19_,
         u5_mult_82_SUMB_36__20_, u5_mult_82_SUMB_36__21_,
         u5_mult_82_SUMB_36__22_, u5_mult_82_SUMB_36__23_,
         u5_mult_82_SUMB_36__24_, u5_mult_82_SUMB_36__25_,
         u5_mult_82_SUMB_36__26_, u5_mult_82_SUMB_36__27_,
         u5_mult_82_SUMB_36__28_, u5_mult_82_SUMB_36__29_,
         u5_mult_82_SUMB_36__30_, u5_mult_82_SUMB_36__31_,
         u5_mult_82_SUMB_36__32_, u5_mult_82_SUMB_36__33_,
         u5_mult_82_SUMB_36__34_, u5_mult_82_SUMB_36__35_,
         u5_mult_82_SUMB_36__36_, u5_mult_82_SUMB_36__37_,
         u5_mult_82_SUMB_36__38_, u5_mult_82_SUMB_36__39_,
         u5_mult_82_SUMB_36__40_, u5_mult_82_SUMB_36__41_,
         u5_mult_82_SUMB_36__42_, u5_mult_82_SUMB_36__43_,
         u5_mult_82_SUMB_36__44_, u5_mult_82_SUMB_36__45_,
         u5_mult_82_SUMB_36__46_, u5_mult_82_SUMB_36__47_,
         u5_mult_82_SUMB_36__48_, u5_mult_82_SUMB_36__49_,
         u5_mult_82_SUMB_36__50_, u5_mult_82_SUMB_36__51_,
         u5_mult_82_SUMB_37__1_, u5_mult_82_SUMB_37__2_,
         u5_mult_82_SUMB_37__3_, u5_mult_82_SUMB_37__4_,
         u5_mult_82_SUMB_37__5_, u5_mult_82_SUMB_37__6_,
         u5_mult_82_SUMB_37__7_, u5_mult_82_SUMB_37__8_,
         u5_mult_82_SUMB_37__9_, u5_mult_82_SUMB_37__10_,
         u5_mult_82_SUMB_37__11_, u5_mult_82_SUMB_37__12_,
         u5_mult_82_SUMB_37__13_, u5_mult_82_SUMB_37__16_,
         u5_mult_82_SUMB_37__17_, u5_mult_82_SUMB_37__18_,
         u5_mult_82_SUMB_37__19_, u5_mult_82_SUMB_37__20_,
         u5_mult_82_SUMB_37__21_, u5_mult_82_SUMB_37__22_,
         u5_mult_82_SUMB_37__23_, u5_mult_82_SUMB_37__24_,
         u5_mult_82_SUMB_37__25_, u5_mult_82_SUMB_37__26_,
         u5_mult_82_SUMB_37__27_, u5_mult_82_SUMB_37__28_,
         u5_mult_82_SUMB_37__29_, u5_mult_82_SUMB_37__30_,
         u5_mult_82_SUMB_37__31_, u5_mult_82_SUMB_37__32_,
         u5_mult_82_SUMB_37__33_, u5_mult_82_SUMB_37__34_,
         u5_mult_82_SUMB_37__35_, u5_mult_82_SUMB_37__36_,
         u5_mult_82_SUMB_37__37_, u5_mult_82_SUMB_37__38_,
         u5_mult_82_SUMB_37__39_, u5_mult_82_SUMB_37__40_,
         u5_mult_82_SUMB_37__41_, u5_mult_82_SUMB_37__42_,
         u5_mult_82_SUMB_37__43_, u5_mult_82_SUMB_37__44_,
         u5_mult_82_SUMB_37__45_, u5_mult_82_SUMB_37__46_,
         u5_mult_82_SUMB_37__47_, u5_mult_82_SUMB_37__48_,
         u5_mult_82_SUMB_37__49_, u5_mult_82_SUMB_37__50_,
         u5_mult_82_SUMB_37__51_, u5_mult_82_SUMB_38__1_,
         u5_mult_82_SUMB_38__2_, u5_mult_82_SUMB_38__3_,
         u5_mult_82_SUMB_38__4_, u5_mult_82_SUMB_38__5_,
         u5_mult_82_SUMB_38__6_, u5_mult_82_SUMB_38__7_,
         u5_mult_82_SUMB_38__8_, u5_mult_82_SUMB_38__9_,
         u5_mult_82_SUMB_38__10_, u5_mult_82_SUMB_38__11_,
         u5_mult_82_SUMB_38__12_, u5_mult_82_SUMB_38__13_,
         u5_mult_82_SUMB_38__15_, u5_mult_82_SUMB_38__16_,
         u5_mult_82_SUMB_38__17_, u5_mult_82_SUMB_38__18_,
         u5_mult_82_SUMB_38__19_, u5_mult_82_SUMB_38__20_,
         u5_mult_82_SUMB_38__21_, u5_mult_82_SUMB_38__22_,
         u5_mult_82_SUMB_38__23_, u5_mult_82_SUMB_38__24_,
         u5_mult_82_SUMB_38__25_, u5_mult_82_SUMB_38__26_,
         u5_mult_82_SUMB_38__27_, u5_mult_82_SUMB_38__28_,
         u5_mult_82_SUMB_38__29_, u5_mult_82_SUMB_38__30_,
         u5_mult_82_SUMB_38__31_, u5_mult_82_SUMB_38__32_,
         u5_mult_82_SUMB_38__33_, u5_mult_82_SUMB_38__34_,
         u5_mult_82_SUMB_38__35_, u5_mult_82_SUMB_38__36_,
         u5_mult_82_SUMB_38__37_, u5_mult_82_SUMB_38__38_,
         u5_mult_82_SUMB_38__39_, u5_mult_82_SUMB_38__40_,
         u5_mult_82_SUMB_38__41_, u5_mult_82_SUMB_38__42_,
         u5_mult_82_SUMB_38__43_, u5_mult_82_SUMB_38__44_,
         u5_mult_82_SUMB_38__45_, u5_mult_82_SUMB_38__46_,
         u5_mult_82_SUMB_38__47_, u5_mult_82_SUMB_38__48_,
         u5_mult_82_SUMB_38__49_, u5_mult_82_SUMB_38__50_,
         u5_mult_82_SUMB_38__51_, u5_mult_82_SUMB_39__1_,
         u5_mult_82_SUMB_39__2_, u5_mult_82_SUMB_39__3_,
         u5_mult_82_SUMB_39__4_, u5_mult_82_SUMB_39__5_,
         u5_mult_82_SUMB_39__6_, u5_mult_82_SUMB_39__7_,
         u5_mult_82_SUMB_39__8_, u5_mult_82_SUMB_39__9_,
         u5_mult_82_SUMB_39__10_, u5_mult_82_SUMB_39__11_,
         u5_mult_82_SUMB_39__12_, u5_mult_82_SUMB_39__14_,
         u5_mult_82_SUMB_39__15_, u5_mult_82_SUMB_39__16_,
         u5_mult_82_SUMB_39__17_, u5_mult_82_SUMB_39__18_,
         u5_mult_82_SUMB_39__19_, u5_mult_82_SUMB_39__20_,
         u5_mult_82_SUMB_39__21_, u5_mult_82_SUMB_39__22_,
         u5_mult_82_SUMB_39__23_, u5_mult_82_SUMB_39__24_,
         u5_mult_82_SUMB_39__25_, u5_mult_82_SUMB_39__26_,
         u5_mult_82_SUMB_39__27_, u5_mult_82_SUMB_39__28_,
         u5_mult_82_SUMB_39__29_, u5_mult_82_SUMB_39__30_,
         u5_mult_82_SUMB_39__31_, u5_mult_82_SUMB_39__32_,
         u5_mult_82_SUMB_39__33_, u5_mult_82_SUMB_39__34_,
         u5_mult_82_SUMB_39__35_, u5_mult_82_SUMB_39__36_,
         u5_mult_82_SUMB_39__37_, u5_mult_82_SUMB_39__38_,
         u5_mult_82_SUMB_39__39_, u5_mult_82_SUMB_39__40_,
         u5_mult_82_SUMB_39__41_, u5_mult_82_SUMB_39__42_,
         u5_mult_82_SUMB_39__43_, u5_mult_82_SUMB_39__44_,
         u5_mult_82_SUMB_39__45_, u5_mult_82_SUMB_39__46_,
         u5_mult_82_SUMB_39__47_, u5_mult_82_SUMB_39__48_,
         u5_mult_82_SUMB_39__49_, u5_mult_82_SUMB_39__50_,
         u5_mult_82_SUMB_39__51_, u5_mult_82_SUMB_40__1_,
         u5_mult_82_SUMB_40__2_, u5_mult_82_SUMB_40__3_,
         u5_mult_82_SUMB_40__4_, u5_mult_82_SUMB_40__5_,
         u5_mult_82_SUMB_40__6_, u5_mult_82_SUMB_40__7_,
         u5_mult_82_SUMB_40__8_, u5_mult_82_SUMB_40__9_,
         u5_mult_82_SUMB_40__10_, u5_mult_82_SUMB_40__11_,
         u5_mult_82_SUMB_40__12_, u5_mult_82_SUMB_40__15_,
         u5_mult_82_SUMB_40__16_, u5_mult_82_SUMB_40__17_,
         u5_mult_82_SUMB_40__18_, u5_mult_82_SUMB_40__19_,
         u5_mult_82_SUMB_40__20_, u5_mult_82_SUMB_40__21_,
         u5_mult_82_SUMB_40__22_, u5_mult_82_SUMB_40__23_,
         u5_mult_82_SUMB_40__24_, u5_mult_82_SUMB_40__25_,
         u5_mult_82_SUMB_40__26_, u5_mult_82_SUMB_40__27_,
         u5_mult_82_SUMB_40__28_, u5_mult_82_SUMB_40__29_,
         u5_mult_82_SUMB_40__30_, u5_mult_82_SUMB_40__31_,
         u5_mult_82_SUMB_40__32_, u5_mult_82_SUMB_40__33_,
         u5_mult_82_SUMB_40__34_, u5_mult_82_SUMB_40__35_,
         u5_mult_82_SUMB_40__36_, u5_mult_82_SUMB_40__37_,
         u5_mult_82_SUMB_40__38_, u5_mult_82_SUMB_40__39_,
         u5_mult_82_SUMB_40__40_, u5_mult_82_SUMB_40__41_,
         u5_mult_82_SUMB_40__42_, u5_mult_82_SUMB_40__43_,
         u5_mult_82_SUMB_40__44_, u5_mult_82_SUMB_40__45_,
         u5_mult_82_SUMB_40__46_, u5_mult_82_SUMB_40__47_,
         u5_mult_82_SUMB_40__48_, u5_mult_82_SUMB_40__49_,
         u5_mult_82_SUMB_40__50_, u5_mult_82_SUMB_40__51_,
         u5_mult_82_SUMB_41__1_, u5_mult_82_SUMB_41__2_,
         u5_mult_82_SUMB_41__3_, u5_mult_82_SUMB_41__4_,
         u5_mult_82_SUMB_41__5_, u5_mult_82_SUMB_41__6_,
         u5_mult_82_SUMB_41__7_, u5_mult_82_SUMB_41__8_,
         u5_mult_82_SUMB_41__9_, u5_mult_82_SUMB_41__10_,
         u5_mult_82_SUMB_41__11_, u5_mult_82_SUMB_41__14_,
         u5_mult_82_SUMB_41__15_, u5_mult_82_SUMB_41__16_,
         u5_mult_82_SUMB_41__17_, u5_mult_82_SUMB_41__18_,
         u5_mult_82_SUMB_41__19_, u5_mult_82_SUMB_41__20_,
         u5_mult_82_SUMB_41__21_, u5_mult_82_SUMB_41__22_,
         u5_mult_82_SUMB_41__23_, u5_mult_82_SUMB_41__24_,
         u5_mult_82_SUMB_41__25_, u5_mult_82_SUMB_41__26_,
         u5_mult_82_SUMB_41__27_, u5_mult_82_SUMB_41__28_,
         u5_mult_82_SUMB_41__29_, u5_mult_82_SUMB_41__30_,
         u5_mult_82_SUMB_41__31_, u5_mult_82_SUMB_41__32_,
         u5_mult_82_SUMB_41__33_, u5_mult_82_SUMB_41__34_,
         u5_mult_82_SUMB_41__35_, u5_mult_82_SUMB_41__36_,
         u5_mult_82_SUMB_41__37_, u5_mult_82_SUMB_41__38_,
         u5_mult_82_SUMB_41__39_, u5_mult_82_SUMB_41__40_,
         u5_mult_82_SUMB_41__41_, u5_mult_82_SUMB_41__42_,
         u5_mult_82_SUMB_41__43_, u5_mult_82_SUMB_41__44_,
         u5_mult_82_SUMB_41__45_, u5_mult_82_SUMB_41__46_,
         u5_mult_82_SUMB_41__47_, u5_mult_82_SUMB_41__48_,
         u5_mult_82_SUMB_41__49_, u5_mult_82_SUMB_41__50_,
         u5_mult_82_SUMB_41__51_, u5_mult_82_SUMB_42__1_,
         u5_mult_82_SUMB_42__2_, u5_mult_82_SUMB_42__3_,
         u5_mult_82_SUMB_42__4_, u5_mult_82_SUMB_42__5_,
         u5_mult_82_SUMB_42__6_, u5_mult_82_SUMB_42__7_,
         u5_mult_82_SUMB_42__8_, u5_mult_82_SUMB_42__9_,
         u5_mult_82_SUMB_42__10_, u5_mult_82_SUMB_42__13_,
         u5_mult_82_SUMB_42__14_, u5_mult_82_SUMB_42__15_,
         u5_mult_82_SUMB_42__16_, u5_mult_82_SUMB_42__17_,
         u5_mult_82_SUMB_42__19_, u5_mult_82_SUMB_42__20_,
         u5_mult_82_SUMB_42__21_, u5_mult_82_SUMB_42__22_,
         u5_mult_82_SUMB_42__23_, u5_mult_82_SUMB_42__24_,
         u5_mult_82_SUMB_42__25_, u5_mult_82_SUMB_42__26_,
         u5_mult_82_SUMB_42__27_, u5_mult_82_SUMB_42__28_,
         u5_mult_82_SUMB_42__29_, u5_mult_82_SUMB_42__30_,
         u5_mult_82_SUMB_42__31_, u5_mult_82_SUMB_42__32_,
         u5_mult_82_SUMB_42__33_, u5_mult_82_SUMB_42__34_,
         u5_mult_82_SUMB_42__35_, u5_mult_82_SUMB_42__36_,
         u5_mult_82_SUMB_42__37_, u5_mult_82_SUMB_42__38_,
         u5_mult_82_SUMB_42__39_, u5_mult_82_SUMB_42__40_,
         u5_mult_82_SUMB_42__41_, u5_mult_82_SUMB_42__42_,
         u5_mult_82_SUMB_42__43_, u5_mult_82_SUMB_42__44_,
         u5_mult_82_SUMB_42__45_, u5_mult_82_SUMB_42__46_,
         u5_mult_82_SUMB_42__47_, u5_mult_82_SUMB_42__48_,
         u5_mult_82_SUMB_42__49_, u5_mult_82_SUMB_42__50_,
         u5_mult_82_SUMB_42__51_, u5_mult_82_SUMB_43__1_,
         u5_mult_82_SUMB_43__2_, u5_mult_82_SUMB_43__3_,
         u5_mult_82_SUMB_43__4_, u5_mult_82_SUMB_43__5_,
         u5_mult_82_SUMB_43__6_, u5_mult_82_SUMB_43__7_,
         u5_mult_82_SUMB_43__8_, u5_mult_82_SUMB_43__9_,
         u5_mult_82_SUMB_43__10_, u5_mult_82_SUMB_43__12_,
         u5_mult_82_SUMB_43__13_, u5_mult_82_SUMB_43__14_,
         u5_mult_82_SUMB_43__15_, u5_mult_82_SUMB_43__16_,
         u5_mult_82_SUMB_43__17_, u5_mult_82_CARRYB_33__36_,
         u5_mult_82_CARRYB_33__37_, u5_mult_82_CARRYB_33__38_,
         u5_mult_82_CARRYB_33__39_, u5_mult_82_CARRYB_33__40_,
         u5_mult_82_CARRYB_33__41_, u5_mult_82_CARRYB_33__42_,
         u5_mult_82_CARRYB_33__43_, u5_mult_82_CARRYB_33__44_,
         u5_mult_82_CARRYB_33__45_, u5_mult_82_CARRYB_33__46_,
         u5_mult_82_CARRYB_33__47_, u5_mult_82_CARRYB_33__48_,
         u5_mult_82_CARRYB_33__49_, u5_mult_82_CARRYB_33__50_,
         u5_mult_82_CARRYB_33__51_, u5_mult_82_CARRYB_34__0_,
         u5_mult_82_CARRYB_34__1_, u5_mult_82_CARRYB_34__2_,
         u5_mult_82_CARRYB_34__3_, u5_mult_82_CARRYB_34__4_,
         u5_mult_82_CARRYB_34__5_, u5_mult_82_CARRYB_34__6_,
         u5_mult_82_CARRYB_34__7_, u5_mult_82_CARRYB_34__8_,
         u5_mult_82_CARRYB_34__9_, u5_mult_82_CARRYB_34__10_,
         u5_mult_82_CARRYB_34__11_, u5_mult_82_CARRYB_34__12_,
         u5_mult_82_CARRYB_34__13_, u5_mult_82_CARRYB_34__14_,
         u5_mult_82_CARRYB_34__15_, u5_mult_82_CARRYB_34__17_,
         u5_mult_82_CARRYB_34__18_, u5_mult_82_CARRYB_34__19_,
         u5_mult_82_CARRYB_34__20_, u5_mult_82_CARRYB_34__21_,
         u5_mult_82_CARRYB_34__22_, u5_mult_82_CARRYB_34__23_,
         u5_mult_82_CARRYB_34__24_, u5_mult_82_CARRYB_34__25_,
         u5_mult_82_CARRYB_34__26_, u5_mult_82_CARRYB_34__27_,
         u5_mult_82_CARRYB_34__28_, u5_mult_82_CARRYB_34__29_,
         u5_mult_82_CARRYB_34__30_, u5_mult_82_CARRYB_34__31_,
         u5_mult_82_CARRYB_34__32_, u5_mult_82_CARRYB_34__33_,
         u5_mult_82_CARRYB_34__34_, u5_mult_82_CARRYB_34__35_,
         u5_mult_82_CARRYB_34__36_, u5_mult_82_CARRYB_34__37_,
         u5_mult_82_CARRYB_34__38_, u5_mult_82_CARRYB_34__39_,
         u5_mult_82_CARRYB_34__40_, u5_mult_82_CARRYB_34__41_,
         u5_mult_82_CARRYB_34__42_, u5_mult_82_CARRYB_34__43_,
         u5_mult_82_CARRYB_34__44_, u5_mult_82_CARRYB_34__45_,
         u5_mult_82_CARRYB_34__46_, u5_mult_82_CARRYB_34__47_,
         u5_mult_82_CARRYB_34__48_, u5_mult_82_CARRYB_34__49_,
         u5_mult_82_CARRYB_34__50_, u5_mult_82_CARRYB_34__51_,
         u5_mult_82_CARRYB_35__0_, u5_mult_82_CARRYB_35__1_,
         u5_mult_82_CARRYB_35__2_, u5_mult_82_CARRYB_35__3_,
         u5_mult_82_CARRYB_35__4_, u5_mult_82_CARRYB_35__5_,
         u5_mult_82_CARRYB_35__6_, u5_mult_82_CARRYB_35__7_,
         u5_mult_82_CARRYB_35__8_, u5_mult_82_CARRYB_35__9_,
         u5_mult_82_CARRYB_35__10_, u5_mult_82_CARRYB_35__11_,
         u5_mult_82_CARRYB_35__12_, u5_mult_82_CARRYB_35__13_,
         u5_mult_82_CARRYB_35__14_, u5_mult_82_CARRYB_35__16_,
         u5_mult_82_CARRYB_35__17_, u5_mult_82_CARRYB_35__18_,
         u5_mult_82_CARRYB_35__19_, u5_mult_82_CARRYB_35__20_,
         u5_mult_82_CARRYB_35__21_, u5_mult_82_CARRYB_35__22_,
         u5_mult_82_CARRYB_35__23_, u5_mult_82_CARRYB_35__24_,
         u5_mult_82_CARRYB_35__25_, u5_mult_82_CARRYB_35__26_,
         u5_mult_82_CARRYB_35__27_, u5_mult_82_CARRYB_35__28_,
         u5_mult_82_CARRYB_35__29_, u5_mult_82_CARRYB_35__30_,
         u5_mult_82_CARRYB_35__31_, u5_mult_82_CARRYB_35__32_,
         u5_mult_82_CARRYB_35__33_, u5_mult_82_CARRYB_35__34_,
         u5_mult_82_CARRYB_35__35_, u5_mult_82_CARRYB_35__36_,
         u5_mult_82_CARRYB_35__37_, u5_mult_82_CARRYB_35__38_,
         u5_mult_82_CARRYB_35__39_, u5_mult_82_CARRYB_35__40_,
         u5_mult_82_CARRYB_35__41_, u5_mult_82_CARRYB_35__42_,
         u5_mult_82_CARRYB_35__43_, u5_mult_82_CARRYB_35__44_,
         u5_mult_82_CARRYB_35__45_, u5_mult_82_CARRYB_35__46_,
         u5_mult_82_CARRYB_35__47_, u5_mult_82_CARRYB_35__48_,
         u5_mult_82_CARRYB_35__49_, u5_mult_82_CARRYB_35__50_,
         u5_mult_82_CARRYB_35__51_, u5_mult_82_CARRYB_36__0_,
         u5_mult_82_CARRYB_36__1_, u5_mult_82_CARRYB_36__2_,
         u5_mult_82_CARRYB_36__3_, u5_mult_82_CARRYB_36__4_,
         u5_mult_82_CARRYB_36__5_, u5_mult_82_CARRYB_36__6_,
         u5_mult_82_CARRYB_36__7_, u5_mult_82_CARRYB_36__8_,
         u5_mult_82_CARRYB_36__9_, u5_mult_82_CARRYB_36__10_,
         u5_mult_82_CARRYB_36__11_, u5_mult_82_CARRYB_36__12_,
         u5_mult_82_CARRYB_36__13_, u5_mult_82_CARRYB_36__15_,
         u5_mult_82_CARRYB_36__16_, u5_mult_82_CARRYB_36__17_,
         u5_mult_82_CARRYB_36__18_, u5_mult_82_CARRYB_36__19_,
         u5_mult_82_CARRYB_36__20_, u5_mult_82_CARRYB_36__21_,
         u5_mult_82_CARRYB_36__22_, u5_mult_82_CARRYB_36__23_,
         u5_mult_82_CARRYB_36__24_, u5_mult_82_CARRYB_36__25_,
         u5_mult_82_CARRYB_36__26_, u5_mult_82_CARRYB_36__27_,
         u5_mult_82_CARRYB_36__28_, u5_mult_82_CARRYB_36__29_,
         u5_mult_82_CARRYB_36__30_, u5_mult_82_CARRYB_36__31_,
         u5_mult_82_CARRYB_36__32_, u5_mult_82_CARRYB_36__33_,
         u5_mult_82_CARRYB_36__34_, u5_mult_82_CARRYB_36__35_,
         u5_mult_82_CARRYB_36__36_, u5_mult_82_CARRYB_36__37_,
         u5_mult_82_CARRYB_36__38_, u5_mult_82_CARRYB_36__39_,
         u5_mult_82_CARRYB_36__40_, u5_mult_82_CARRYB_36__41_,
         u5_mult_82_CARRYB_36__42_, u5_mult_82_CARRYB_36__43_,
         u5_mult_82_CARRYB_36__44_, u5_mult_82_CARRYB_36__45_,
         u5_mult_82_CARRYB_36__46_, u5_mult_82_CARRYB_36__47_,
         u5_mult_82_CARRYB_36__48_, u5_mult_82_CARRYB_36__49_,
         u5_mult_82_CARRYB_36__50_, u5_mult_82_CARRYB_36__51_,
         u5_mult_82_CARRYB_37__0_, u5_mult_82_CARRYB_37__1_,
         u5_mult_82_CARRYB_37__2_, u5_mult_82_CARRYB_37__3_,
         u5_mult_82_CARRYB_37__4_, u5_mult_82_CARRYB_37__5_,
         u5_mult_82_CARRYB_37__6_, u5_mult_82_CARRYB_37__7_,
         u5_mult_82_CARRYB_37__8_, u5_mult_82_CARRYB_37__9_,
         u5_mult_82_CARRYB_37__10_, u5_mult_82_CARRYB_37__11_,
         u5_mult_82_CARRYB_37__12_, u5_mult_82_CARRYB_37__13_,
         u5_mult_82_CARRYB_37__15_, u5_mult_82_CARRYB_37__16_,
         u5_mult_82_CARRYB_37__17_, u5_mult_82_CARRYB_37__18_,
         u5_mult_82_CARRYB_37__19_, u5_mult_82_CARRYB_37__20_,
         u5_mult_82_CARRYB_37__21_, u5_mult_82_CARRYB_37__22_,
         u5_mult_82_CARRYB_37__23_, u5_mult_82_CARRYB_37__24_,
         u5_mult_82_CARRYB_37__25_, u5_mult_82_CARRYB_37__26_,
         u5_mult_82_CARRYB_37__27_, u5_mult_82_CARRYB_37__28_,
         u5_mult_82_CARRYB_37__29_, u5_mult_82_CARRYB_37__30_,
         u5_mult_82_CARRYB_37__31_, u5_mult_82_CARRYB_37__32_,
         u5_mult_82_CARRYB_37__33_, u5_mult_82_CARRYB_37__34_,
         u5_mult_82_CARRYB_37__35_, u5_mult_82_CARRYB_37__36_,
         u5_mult_82_CARRYB_37__37_, u5_mult_82_CARRYB_37__38_,
         u5_mult_82_CARRYB_37__39_, u5_mult_82_CARRYB_37__40_,
         u5_mult_82_CARRYB_37__41_, u5_mult_82_CARRYB_37__42_,
         u5_mult_82_CARRYB_37__43_, u5_mult_82_CARRYB_37__44_,
         u5_mult_82_CARRYB_37__45_, u5_mult_82_CARRYB_37__46_,
         u5_mult_82_CARRYB_37__47_, u5_mult_82_CARRYB_37__48_,
         u5_mult_82_CARRYB_37__49_, u5_mult_82_CARRYB_37__50_,
         u5_mult_82_CARRYB_37__51_, u5_mult_82_CARRYB_38__0_,
         u5_mult_82_CARRYB_38__1_, u5_mult_82_CARRYB_38__2_,
         u5_mult_82_CARRYB_38__3_, u5_mult_82_CARRYB_38__4_,
         u5_mult_82_CARRYB_38__5_, u5_mult_82_CARRYB_38__6_,
         u5_mult_82_CARRYB_38__7_, u5_mult_82_CARRYB_38__8_,
         u5_mult_82_CARRYB_38__9_, u5_mult_82_CARRYB_38__10_,
         u5_mult_82_CARRYB_38__11_, u5_mult_82_CARRYB_38__12_,
         u5_mult_82_CARRYB_38__13_, u5_mult_82_CARRYB_38__15_,
         u5_mult_82_CARRYB_38__16_, u5_mult_82_CARRYB_38__17_,
         u5_mult_82_CARRYB_38__18_, u5_mult_82_CARRYB_38__19_,
         u5_mult_82_CARRYB_38__20_, u5_mult_82_CARRYB_38__21_,
         u5_mult_82_CARRYB_38__22_, u5_mult_82_CARRYB_38__23_,
         u5_mult_82_CARRYB_38__24_, u5_mult_82_CARRYB_38__25_,
         u5_mult_82_CARRYB_38__26_, u5_mult_82_CARRYB_38__27_,
         u5_mult_82_CARRYB_38__28_, u5_mult_82_CARRYB_38__29_,
         u5_mult_82_CARRYB_38__30_, u5_mult_82_CARRYB_38__31_,
         u5_mult_82_CARRYB_38__32_, u5_mult_82_CARRYB_38__33_,
         u5_mult_82_CARRYB_38__34_, u5_mult_82_CARRYB_38__35_,
         u5_mult_82_CARRYB_38__36_, u5_mult_82_CARRYB_38__37_,
         u5_mult_82_CARRYB_38__38_, u5_mult_82_CARRYB_38__39_,
         u5_mult_82_CARRYB_38__40_, u5_mult_82_CARRYB_38__41_,
         u5_mult_82_CARRYB_38__42_, u5_mult_82_CARRYB_38__43_,
         u5_mult_82_CARRYB_38__44_, u5_mult_82_CARRYB_38__45_,
         u5_mult_82_CARRYB_38__46_, u5_mult_82_CARRYB_38__47_,
         u5_mult_82_CARRYB_38__48_, u5_mult_82_CARRYB_38__49_,
         u5_mult_82_CARRYB_38__50_, u5_mult_82_CARRYB_38__51_,
         u5_mult_82_CARRYB_39__0_, u5_mult_82_CARRYB_39__1_,
         u5_mult_82_CARRYB_39__2_, u5_mult_82_CARRYB_39__3_,
         u5_mult_82_CARRYB_39__4_, u5_mult_82_CARRYB_39__5_,
         u5_mult_82_CARRYB_39__6_, u5_mult_82_CARRYB_39__7_,
         u5_mult_82_CARRYB_39__8_, u5_mult_82_CARRYB_39__9_,
         u5_mult_82_CARRYB_39__10_, u5_mult_82_CARRYB_39__11_,
         u5_mult_82_CARRYB_39__13_, u5_mult_82_CARRYB_39__14_,
         u5_mult_82_CARRYB_39__15_, u5_mult_82_CARRYB_39__16_,
         u5_mult_82_CARRYB_39__17_, u5_mult_82_CARRYB_39__18_,
         u5_mult_82_CARRYB_39__19_, u5_mult_82_CARRYB_39__20_,
         u5_mult_82_CARRYB_39__21_, u5_mult_82_CARRYB_39__22_,
         u5_mult_82_CARRYB_39__23_, u5_mult_82_CARRYB_39__24_,
         u5_mult_82_CARRYB_39__25_, u5_mult_82_CARRYB_39__26_,
         u5_mult_82_CARRYB_39__27_, u5_mult_82_CARRYB_39__28_,
         u5_mult_82_CARRYB_39__29_, u5_mult_82_CARRYB_39__30_,
         u5_mult_82_CARRYB_39__31_, u5_mult_82_CARRYB_39__32_,
         u5_mult_82_CARRYB_39__33_, u5_mult_82_CARRYB_39__34_,
         u5_mult_82_CARRYB_39__35_, u5_mult_82_CARRYB_39__36_,
         u5_mult_82_CARRYB_39__37_, u5_mult_82_CARRYB_39__38_,
         u5_mult_82_CARRYB_39__39_, u5_mult_82_CARRYB_39__40_,
         u5_mult_82_CARRYB_39__41_, u5_mult_82_CARRYB_39__42_,
         u5_mult_82_CARRYB_39__43_, u5_mult_82_CARRYB_39__44_,
         u5_mult_82_CARRYB_39__45_, u5_mult_82_CARRYB_39__46_,
         u5_mult_82_CARRYB_39__47_, u5_mult_82_CARRYB_39__48_,
         u5_mult_82_CARRYB_39__49_, u5_mult_82_CARRYB_39__50_,
         u5_mult_82_CARRYB_39__51_, u5_mult_82_CARRYB_40__0_,
         u5_mult_82_CARRYB_40__1_, u5_mult_82_CARRYB_40__2_,
         u5_mult_82_CARRYB_40__3_, u5_mult_82_CARRYB_40__4_,
         u5_mult_82_CARRYB_40__5_, u5_mult_82_CARRYB_40__6_,
         u5_mult_82_CARRYB_40__7_, u5_mult_82_CARRYB_40__8_,
         u5_mult_82_CARRYB_40__9_, u5_mult_82_CARRYB_40__10_,
         u5_mult_82_CARRYB_40__11_, u5_mult_82_CARRYB_40__13_,
         u5_mult_82_CARRYB_40__14_, u5_mult_82_CARRYB_40__15_,
         u5_mult_82_CARRYB_40__16_, u5_mult_82_CARRYB_40__17_,
         u5_mult_82_CARRYB_40__18_, u5_mult_82_CARRYB_40__19_,
         u5_mult_82_CARRYB_40__20_, u5_mult_82_CARRYB_40__21_,
         u5_mult_82_CARRYB_40__22_, u5_mult_82_CARRYB_40__23_,
         u5_mult_82_CARRYB_40__24_, u5_mult_82_CARRYB_40__25_,
         u5_mult_82_CARRYB_40__26_, u5_mult_82_CARRYB_40__27_,
         u5_mult_82_CARRYB_40__28_, u5_mult_82_CARRYB_40__29_,
         u5_mult_82_CARRYB_40__30_, u5_mult_82_CARRYB_40__31_,
         u5_mult_82_CARRYB_40__32_, u5_mult_82_CARRYB_40__33_,
         u5_mult_82_CARRYB_40__34_, u5_mult_82_CARRYB_40__35_,
         u5_mult_82_CARRYB_40__36_, u5_mult_82_CARRYB_40__37_,
         u5_mult_82_CARRYB_40__38_, u5_mult_82_CARRYB_40__39_,
         u5_mult_82_CARRYB_40__40_, u5_mult_82_CARRYB_40__41_,
         u5_mult_82_CARRYB_40__42_, u5_mult_82_CARRYB_40__43_,
         u5_mult_82_CARRYB_40__44_, u5_mult_82_CARRYB_40__45_,
         u5_mult_82_CARRYB_40__46_, u5_mult_82_CARRYB_40__47_,
         u5_mult_82_CARRYB_40__48_, u5_mult_82_CARRYB_40__49_,
         u5_mult_82_CARRYB_40__50_, u5_mult_82_CARRYB_40__51_,
         u5_mult_82_CARRYB_41__0_, u5_mult_82_CARRYB_41__1_,
         u5_mult_82_CARRYB_41__2_, u5_mult_82_CARRYB_41__3_,
         u5_mult_82_CARRYB_41__4_, u5_mult_82_CARRYB_41__5_,
         u5_mult_82_CARRYB_41__6_, u5_mult_82_CARRYB_41__7_,
         u5_mult_82_CARRYB_41__8_, u5_mult_82_CARRYB_41__9_,
         u5_mult_82_CARRYB_41__10_, u5_mult_82_CARRYB_41__12_,
         u5_mult_82_CARRYB_41__14_, u5_mult_82_CARRYB_41__15_,
         u5_mult_82_CARRYB_41__16_, u5_mult_82_CARRYB_41__17_,
         u5_mult_82_CARRYB_41__18_, u5_mult_82_CARRYB_41__19_,
         u5_mult_82_CARRYB_41__20_, u5_mult_82_CARRYB_41__21_,
         u5_mult_82_CARRYB_41__22_, u5_mult_82_CARRYB_41__23_,
         u5_mult_82_CARRYB_41__24_, u5_mult_82_CARRYB_41__25_,
         u5_mult_82_CARRYB_41__26_, u5_mult_82_CARRYB_41__27_,
         u5_mult_82_CARRYB_41__28_, u5_mult_82_CARRYB_41__29_,
         u5_mult_82_CARRYB_41__30_, u5_mult_82_CARRYB_41__31_,
         u5_mult_82_CARRYB_41__32_, u5_mult_82_CARRYB_41__33_,
         u5_mult_82_CARRYB_41__34_, u5_mult_82_CARRYB_41__35_,
         u5_mult_82_CARRYB_41__36_, u5_mult_82_CARRYB_41__37_,
         u5_mult_82_CARRYB_41__38_, u5_mult_82_CARRYB_41__39_,
         u5_mult_82_CARRYB_41__40_, u5_mult_82_CARRYB_41__41_,
         u5_mult_82_CARRYB_41__42_, u5_mult_82_CARRYB_41__43_,
         u5_mult_82_CARRYB_41__44_, u5_mult_82_CARRYB_41__45_,
         u5_mult_82_CARRYB_41__46_, u5_mult_82_CARRYB_41__47_,
         u5_mult_82_CARRYB_41__48_, u5_mult_82_CARRYB_41__49_,
         u5_mult_82_CARRYB_41__50_, u5_mult_82_CARRYB_41__51_,
         u5_mult_82_CARRYB_42__0_, u5_mult_82_CARRYB_42__1_,
         u5_mult_82_CARRYB_42__2_, u5_mult_82_CARRYB_42__3_,
         u5_mult_82_CARRYB_42__4_, u5_mult_82_CARRYB_42__5_,
         u5_mult_82_CARRYB_42__6_, u5_mult_82_CARRYB_42__7_,
         u5_mult_82_CARRYB_42__8_, u5_mult_82_CARRYB_42__9_,
         u5_mult_82_CARRYB_42__10_, u5_mult_82_CARRYB_42__11_,
         u5_mult_82_CARRYB_42__13_, u5_mult_82_CARRYB_42__14_,
         u5_mult_82_CARRYB_42__15_, u5_mult_82_CARRYB_42__16_,
         u5_mult_82_CARRYB_42__17_, u5_mult_82_CARRYB_42__18_,
         u5_mult_82_CARRYB_42__19_, u5_mult_82_CARRYB_42__20_,
         u5_mult_82_CARRYB_42__21_, u5_mult_82_CARRYB_42__22_,
         u5_mult_82_CARRYB_42__23_, u5_mult_82_CARRYB_42__24_,
         u5_mult_82_CARRYB_42__25_, u5_mult_82_CARRYB_42__26_,
         u5_mult_82_CARRYB_42__27_, u5_mult_82_CARRYB_42__28_,
         u5_mult_82_CARRYB_42__29_, u5_mult_82_CARRYB_42__30_,
         u5_mult_82_CARRYB_42__31_, u5_mult_82_CARRYB_42__32_,
         u5_mult_82_CARRYB_42__33_, u5_mult_82_CARRYB_42__34_,
         u5_mult_82_CARRYB_42__35_, u5_mult_82_CARRYB_42__36_,
         u5_mult_82_CARRYB_42__37_, u5_mult_82_CARRYB_42__38_,
         u5_mult_82_CARRYB_42__39_, u5_mult_82_CARRYB_42__40_,
         u5_mult_82_CARRYB_42__41_, u5_mult_82_CARRYB_42__42_,
         u5_mult_82_CARRYB_42__43_, u5_mult_82_CARRYB_42__44_,
         u5_mult_82_CARRYB_42__45_, u5_mult_82_CARRYB_42__46_,
         u5_mult_82_CARRYB_42__47_, u5_mult_82_CARRYB_42__48_,
         u5_mult_82_CARRYB_42__49_, u5_mult_82_CARRYB_42__50_,
         u5_mult_82_CARRYB_42__51_, u5_mult_82_CARRYB_43__0_,
         u5_mult_82_CARRYB_43__1_, u5_mult_82_CARRYB_43__2_,
         u5_mult_82_CARRYB_43__3_, u5_mult_82_CARRYB_43__4_,
         u5_mult_82_CARRYB_43__5_, u5_mult_82_CARRYB_43__6_,
         u5_mult_82_CARRYB_43__7_, u5_mult_82_CARRYB_43__8_,
         u5_mult_82_CARRYB_43__9_, u5_mult_82_CARRYB_43__10_,
         u5_mult_82_CARRYB_43__12_, u5_mult_82_CARRYB_43__13_,
         u5_mult_82_CARRYB_43__14_, u5_mult_82_CARRYB_43__15_,
         u5_mult_82_CARRYB_43__16_, u5_mult_82_CARRYB_43__17_,
         u5_mult_82_SUMB_24__1_, u5_mult_82_SUMB_24__2_,
         u5_mult_82_SUMB_24__3_, u5_mult_82_SUMB_24__4_,
         u5_mult_82_SUMB_24__5_, u5_mult_82_SUMB_24__6_,
         u5_mult_82_SUMB_24__7_, u5_mult_82_SUMB_24__8_,
         u5_mult_82_SUMB_24__9_, u5_mult_82_SUMB_24__10_,
         u5_mult_82_SUMB_24__11_, u5_mult_82_SUMB_24__12_,
         u5_mult_82_SUMB_24__13_, u5_mult_82_SUMB_24__14_,
         u5_mult_82_SUMB_24__15_, u5_mult_82_SUMB_24__16_,
         u5_mult_82_SUMB_24__17_, u5_mult_82_SUMB_24__18_,
         u5_mult_82_SUMB_24__19_, u5_mult_82_SUMB_24__20_,
         u5_mult_82_SUMB_24__21_, u5_mult_82_SUMB_24__22_,
         u5_mult_82_SUMB_24__24_, u5_mult_82_SUMB_24__25_,
         u5_mult_82_SUMB_24__26_, u5_mult_82_SUMB_24__27_,
         u5_mult_82_SUMB_24__28_, u5_mult_82_SUMB_24__29_,
         u5_mult_82_SUMB_24__30_, u5_mult_82_SUMB_24__31_,
         u5_mult_82_SUMB_24__32_, u5_mult_82_SUMB_24__33_,
         u5_mult_82_SUMB_24__34_, u5_mult_82_SUMB_24__35_,
         u5_mult_82_SUMB_24__36_, u5_mult_82_SUMB_24__37_,
         u5_mult_82_SUMB_24__38_, u5_mult_82_SUMB_24__39_,
         u5_mult_82_SUMB_24__40_, u5_mult_82_SUMB_24__41_,
         u5_mult_82_SUMB_24__42_, u5_mult_82_SUMB_24__43_,
         u5_mult_82_SUMB_24__44_, u5_mult_82_SUMB_24__45_,
         u5_mult_82_SUMB_24__46_, u5_mult_82_SUMB_24__47_,
         u5_mult_82_SUMB_24__48_, u5_mult_82_SUMB_24__49_,
         u5_mult_82_SUMB_24__50_, u5_mult_82_SUMB_24__51_,
         u5_mult_82_SUMB_25__1_, u5_mult_82_SUMB_25__2_,
         u5_mult_82_SUMB_25__3_, u5_mult_82_SUMB_25__4_,
         u5_mult_82_SUMB_25__5_, u5_mult_82_SUMB_25__6_,
         u5_mult_82_SUMB_25__7_, u5_mult_82_SUMB_25__8_,
         u5_mult_82_SUMB_25__9_, u5_mult_82_SUMB_25__10_,
         u5_mult_82_SUMB_25__11_, u5_mult_82_SUMB_25__12_,
         u5_mult_82_SUMB_25__13_, u5_mult_82_SUMB_25__14_,
         u5_mult_82_SUMB_25__15_, u5_mult_82_SUMB_25__16_,
         u5_mult_82_SUMB_25__17_, u5_mult_82_SUMB_25__18_,
         u5_mult_82_SUMB_25__19_, u5_mult_82_SUMB_25__20_,
         u5_mult_82_SUMB_25__21_, u5_mult_82_SUMB_25__23_,
         u5_mult_82_SUMB_25__24_, u5_mult_82_SUMB_25__25_,
         u5_mult_82_SUMB_25__26_, u5_mult_82_SUMB_25__27_,
         u5_mult_82_SUMB_25__28_, u5_mult_82_SUMB_25__29_,
         u5_mult_82_SUMB_25__30_, u5_mult_82_SUMB_25__31_,
         u5_mult_82_SUMB_25__32_, u5_mult_82_SUMB_25__33_,
         u5_mult_82_SUMB_25__34_, u5_mult_82_SUMB_25__35_,
         u5_mult_82_SUMB_25__36_, u5_mult_82_SUMB_25__37_,
         u5_mult_82_SUMB_25__38_, u5_mult_82_SUMB_25__39_,
         u5_mult_82_SUMB_25__40_, u5_mult_82_SUMB_25__41_,
         u5_mult_82_SUMB_25__42_, u5_mult_82_SUMB_25__43_,
         u5_mult_82_SUMB_25__44_, u5_mult_82_SUMB_25__45_,
         u5_mult_82_SUMB_25__46_, u5_mult_82_SUMB_25__47_,
         u5_mult_82_SUMB_25__48_, u5_mult_82_SUMB_25__49_,
         u5_mult_82_SUMB_25__50_, u5_mult_82_SUMB_25__51_,
         u5_mult_82_SUMB_26__1_, u5_mult_82_SUMB_26__2_,
         u5_mult_82_SUMB_26__3_, u5_mult_82_SUMB_26__4_,
         u5_mult_82_SUMB_26__5_, u5_mult_82_SUMB_26__6_,
         u5_mult_82_SUMB_26__7_, u5_mult_82_SUMB_26__8_,
         u5_mult_82_SUMB_26__9_, u5_mult_82_SUMB_26__10_,
         u5_mult_82_SUMB_26__11_, u5_mult_82_SUMB_26__12_,
         u5_mult_82_SUMB_26__13_, u5_mult_82_SUMB_26__14_,
         u5_mult_82_SUMB_26__15_, u5_mult_82_SUMB_26__16_,
         u5_mult_82_SUMB_26__17_, u5_mult_82_SUMB_26__18_,
         u5_mult_82_SUMB_26__19_, u5_mult_82_SUMB_26__20_,
         u5_mult_82_SUMB_26__22_, u5_mult_82_SUMB_26__23_,
         u5_mult_82_SUMB_26__24_, u5_mult_82_SUMB_26__25_,
         u5_mult_82_SUMB_26__26_, u5_mult_82_SUMB_26__27_,
         u5_mult_82_SUMB_26__28_, u5_mult_82_SUMB_26__29_,
         u5_mult_82_SUMB_26__30_, u5_mult_82_SUMB_26__31_,
         u5_mult_82_SUMB_26__32_, u5_mult_82_SUMB_26__33_,
         u5_mult_82_SUMB_26__34_, u5_mult_82_SUMB_26__35_,
         u5_mult_82_SUMB_26__36_, u5_mult_82_SUMB_26__37_,
         u5_mult_82_SUMB_26__38_, u5_mult_82_SUMB_26__39_,
         u5_mult_82_SUMB_26__40_, u5_mult_82_SUMB_26__41_,
         u5_mult_82_SUMB_26__42_, u5_mult_82_SUMB_26__43_,
         u5_mult_82_SUMB_26__44_, u5_mult_82_SUMB_26__45_,
         u5_mult_82_SUMB_26__46_, u5_mult_82_SUMB_26__47_,
         u5_mult_82_SUMB_26__48_, u5_mult_82_SUMB_26__49_,
         u5_mult_82_SUMB_26__50_, u5_mult_82_SUMB_26__51_,
         u5_mult_82_SUMB_27__1_, u5_mult_82_SUMB_27__2_,
         u5_mult_82_SUMB_27__3_, u5_mult_82_SUMB_27__4_,
         u5_mult_82_SUMB_27__5_, u5_mult_82_SUMB_27__6_,
         u5_mult_82_SUMB_27__7_, u5_mult_82_SUMB_27__8_,
         u5_mult_82_SUMB_27__9_, u5_mult_82_SUMB_27__10_,
         u5_mult_82_SUMB_27__11_, u5_mult_82_SUMB_27__12_,
         u5_mult_82_SUMB_27__13_, u5_mult_82_SUMB_27__14_,
         u5_mult_82_SUMB_27__15_, u5_mult_82_SUMB_27__16_,
         u5_mult_82_SUMB_27__17_, u5_mult_82_SUMB_27__18_,
         u5_mult_82_SUMB_27__19_, u5_mult_82_SUMB_27__21_,
         u5_mult_82_SUMB_27__22_, u5_mult_82_SUMB_27__23_,
         u5_mult_82_SUMB_27__24_, u5_mult_82_SUMB_27__25_,
         u5_mult_82_SUMB_27__26_, u5_mult_82_SUMB_27__27_,
         u5_mult_82_SUMB_27__28_, u5_mult_82_SUMB_27__29_,
         u5_mult_82_SUMB_27__30_, u5_mult_82_SUMB_27__31_,
         u5_mult_82_SUMB_27__32_, u5_mult_82_SUMB_27__33_,
         u5_mult_82_SUMB_27__34_, u5_mult_82_SUMB_27__35_,
         u5_mult_82_SUMB_27__36_, u5_mult_82_SUMB_27__37_,
         u5_mult_82_SUMB_27__38_, u5_mult_82_SUMB_27__39_,
         u5_mult_82_SUMB_27__40_, u5_mult_82_SUMB_27__41_,
         u5_mult_82_SUMB_27__42_, u5_mult_82_SUMB_27__43_,
         u5_mult_82_SUMB_27__44_, u5_mult_82_SUMB_27__45_,
         u5_mult_82_SUMB_27__46_, u5_mult_82_SUMB_27__47_,
         u5_mult_82_SUMB_27__48_, u5_mult_82_SUMB_27__49_,
         u5_mult_82_SUMB_27__50_, u5_mult_82_SUMB_27__51_,
         u5_mult_82_SUMB_28__1_, u5_mult_82_SUMB_28__2_,
         u5_mult_82_SUMB_28__3_, u5_mult_82_SUMB_28__4_,
         u5_mult_82_SUMB_28__5_, u5_mult_82_SUMB_28__6_,
         u5_mult_82_SUMB_28__7_, u5_mult_82_SUMB_28__8_,
         u5_mult_82_SUMB_28__9_, u5_mult_82_SUMB_28__10_,
         u5_mult_82_SUMB_28__11_, u5_mult_82_SUMB_28__12_,
         u5_mult_82_SUMB_28__13_, u5_mult_82_SUMB_28__14_,
         u5_mult_82_SUMB_28__15_, u5_mult_82_SUMB_28__16_,
         u5_mult_82_SUMB_28__17_, u5_mult_82_SUMB_28__18_,
         u5_mult_82_SUMB_28__19_, u5_mult_82_SUMB_28__21_,
         u5_mult_82_SUMB_28__22_, u5_mult_82_SUMB_28__23_,
         u5_mult_82_SUMB_28__24_, u5_mult_82_SUMB_28__25_,
         u5_mult_82_SUMB_28__26_, u5_mult_82_SUMB_28__27_,
         u5_mult_82_SUMB_28__28_, u5_mult_82_SUMB_28__29_,
         u5_mult_82_SUMB_28__30_, u5_mult_82_SUMB_28__31_,
         u5_mult_82_SUMB_28__32_, u5_mult_82_SUMB_28__33_,
         u5_mult_82_SUMB_28__34_, u5_mult_82_SUMB_28__35_,
         u5_mult_82_SUMB_28__36_, u5_mult_82_SUMB_28__37_,
         u5_mult_82_SUMB_28__38_, u5_mult_82_SUMB_28__39_,
         u5_mult_82_SUMB_28__41_, u5_mult_82_SUMB_28__42_,
         u5_mult_82_SUMB_28__43_, u5_mult_82_SUMB_28__44_,
         u5_mult_82_SUMB_28__45_, u5_mult_82_SUMB_28__46_,
         u5_mult_82_SUMB_28__47_, u5_mult_82_SUMB_28__48_,
         u5_mult_82_SUMB_28__49_, u5_mult_82_SUMB_28__50_,
         u5_mult_82_SUMB_28__51_, u5_mult_82_SUMB_29__1_,
         u5_mult_82_SUMB_29__2_, u5_mult_82_SUMB_29__3_,
         u5_mult_82_SUMB_29__4_, u5_mult_82_SUMB_29__5_,
         u5_mult_82_SUMB_29__6_, u5_mult_82_SUMB_29__7_,
         u5_mult_82_SUMB_29__8_, u5_mult_82_SUMB_29__9_,
         u5_mult_82_SUMB_29__10_, u5_mult_82_SUMB_29__11_,
         u5_mult_82_SUMB_29__12_, u5_mult_82_SUMB_29__13_,
         u5_mult_82_SUMB_29__14_, u5_mult_82_SUMB_29__15_,
         u5_mult_82_SUMB_29__16_, u5_mult_82_SUMB_29__17_,
         u5_mult_82_SUMB_29__18_, u5_mult_82_SUMB_29__21_,
         u5_mult_82_SUMB_29__22_, u5_mult_82_SUMB_29__23_,
         u5_mult_82_SUMB_29__24_, u5_mult_82_SUMB_29__25_,
         u5_mult_82_SUMB_29__26_, u5_mult_82_SUMB_29__27_,
         u5_mult_82_SUMB_29__28_, u5_mult_82_SUMB_29__29_,
         u5_mult_82_SUMB_29__30_, u5_mult_82_SUMB_29__31_,
         u5_mult_82_SUMB_29__32_, u5_mult_82_SUMB_29__33_,
         u5_mult_82_SUMB_29__34_, u5_mult_82_SUMB_29__35_,
         u5_mult_82_SUMB_29__36_, u5_mult_82_SUMB_29__37_,
         u5_mult_82_SUMB_29__38_, u5_mult_82_SUMB_29__39_,
         u5_mult_82_SUMB_29__40_, u5_mult_82_SUMB_29__41_,
         u5_mult_82_SUMB_29__42_, u5_mult_82_SUMB_29__43_,
         u5_mult_82_SUMB_29__44_, u5_mult_82_SUMB_29__45_,
         u5_mult_82_SUMB_29__46_, u5_mult_82_SUMB_29__47_,
         u5_mult_82_SUMB_29__48_, u5_mult_82_SUMB_29__49_,
         u5_mult_82_SUMB_29__50_, u5_mult_82_SUMB_29__51_,
         u5_mult_82_SUMB_30__1_, u5_mult_82_SUMB_30__2_,
         u5_mult_82_SUMB_30__3_, u5_mult_82_SUMB_30__4_,
         u5_mult_82_SUMB_30__5_, u5_mult_82_SUMB_30__6_,
         u5_mult_82_SUMB_30__7_, u5_mult_82_SUMB_30__8_,
         u5_mult_82_SUMB_30__9_, u5_mult_82_SUMB_30__10_,
         u5_mult_82_SUMB_30__11_, u5_mult_82_SUMB_30__12_,
         u5_mult_82_SUMB_30__13_, u5_mult_82_SUMB_30__14_,
         u5_mult_82_SUMB_30__15_, u5_mult_82_SUMB_30__16_,
         u5_mult_82_SUMB_30__17_, u5_mult_82_SUMB_30__18_,
         u5_mult_82_SUMB_30__20_, u5_mult_82_SUMB_30__21_,
         u5_mult_82_SUMB_30__22_, u5_mult_82_SUMB_30__23_,
         u5_mult_82_SUMB_30__24_, u5_mult_82_SUMB_30__25_,
         u5_mult_82_SUMB_30__26_, u5_mult_82_SUMB_30__27_,
         u5_mult_82_SUMB_30__28_, u5_mult_82_SUMB_30__29_,
         u5_mult_82_SUMB_30__30_, u5_mult_82_SUMB_30__31_,
         u5_mult_82_SUMB_30__32_, u5_mult_82_SUMB_30__33_,
         u5_mult_82_SUMB_30__34_, u5_mult_82_SUMB_30__35_,
         u5_mult_82_SUMB_30__36_, u5_mult_82_SUMB_30__37_,
         u5_mult_82_SUMB_30__38_, u5_mult_82_SUMB_30__39_,
         u5_mult_82_SUMB_30__40_, u5_mult_82_SUMB_30__41_,
         u5_mult_82_SUMB_30__42_, u5_mult_82_SUMB_30__43_,
         u5_mult_82_SUMB_30__44_, u5_mult_82_SUMB_30__45_,
         u5_mult_82_SUMB_30__46_, u5_mult_82_SUMB_30__47_,
         u5_mult_82_SUMB_30__48_, u5_mult_82_SUMB_30__49_,
         u5_mult_82_SUMB_30__50_, u5_mult_82_SUMB_30__51_,
         u5_mult_82_SUMB_31__1_, u5_mult_82_SUMB_31__2_,
         u5_mult_82_SUMB_31__3_, u5_mult_82_SUMB_31__4_,
         u5_mult_82_SUMB_31__5_, u5_mult_82_SUMB_31__6_,
         u5_mult_82_SUMB_31__7_, u5_mult_82_SUMB_31__8_,
         u5_mult_82_SUMB_31__9_, u5_mult_82_SUMB_31__10_,
         u5_mult_82_SUMB_31__11_, u5_mult_82_SUMB_31__12_,
         u5_mult_82_SUMB_31__13_, u5_mult_82_SUMB_31__14_,
         u5_mult_82_SUMB_31__15_, u5_mult_82_SUMB_31__16_,
         u5_mult_82_SUMB_31__17_, u5_mult_82_SUMB_31__19_,
         u5_mult_82_SUMB_31__20_, u5_mult_82_SUMB_31__21_,
         u5_mult_82_SUMB_31__22_, u5_mult_82_SUMB_31__23_,
         u5_mult_82_SUMB_31__24_, u5_mult_82_SUMB_31__25_,
         u5_mult_82_SUMB_31__26_, u5_mult_82_SUMB_31__27_,
         u5_mult_82_SUMB_31__28_, u5_mult_82_SUMB_31__29_,
         u5_mult_82_SUMB_31__30_, u5_mult_82_SUMB_31__31_,
         u5_mult_82_SUMB_31__32_, u5_mult_82_SUMB_31__33_,
         u5_mult_82_SUMB_31__34_, u5_mult_82_SUMB_31__35_,
         u5_mult_82_SUMB_31__36_, u5_mult_82_SUMB_31__37_,
         u5_mult_82_SUMB_31__38_, u5_mult_82_SUMB_31__39_,
         u5_mult_82_SUMB_31__40_, u5_mult_82_SUMB_31__41_,
         u5_mult_82_SUMB_31__42_, u5_mult_82_SUMB_31__43_,
         u5_mult_82_SUMB_31__44_, u5_mult_82_SUMB_31__45_,
         u5_mult_82_SUMB_31__46_, u5_mult_82_SUMB_31__47_,
         u5_mult_82_SUMB_31__48_, u5_mult_82_SUMB_31__49_,
         u5_mult_82_SUMB_31__50_, u5_mult_82_SUMB_31__51_,
         u5_mult_82_SUMB_32__1_, u5_mult_82_SUMB_32__2_,
         u5_mult_82_SUMB_32__3_, u5_mult_82_SUMB_32__4_,
         u5_mult_82_SUMB_32__5_, u5_mult_82_SUMB_32__6_,
         u5_mult_82_SUMB_32__7_, u5_mult_82_SUMB_32__8_,
         u5_mult_82_SUMB_32__9_, u5_mult_82_SUMB_32__10_,
         u5_mult_82_SUMB_32__11_, u5_mult_82_SUMB_32__12_,
         u5_mult_82_SUMB_32__13_, u5_mult_82_SUMB_32__14_,
         u5_mult_82_SUMB_32__15_, u5_mult_82_SUMB_32__16_,
         u5_mult_82_SUMB_32__17_, u5_mult_82_SUMB_32__18_,
         u5_mult_82_SUMB_32__19_, u5_mult_82_SUMB_32__20_,
         u5_mult_82_SUMB_32__21_, u5_mult_82_SUMB_32__22_,
         u5_mult_82_SUMB_32__23_, u5_mult_82_SUMB_32__24_,
         u5_mult_82_SUMB_32__25_, u5_mult_82_SUMB_32__26_,
         u5_mult_82_SUMB_32__27_, u5_mult_82_SUMB_32__28_,
         u5_mult_82_SUMB_32__29_, u5_mult_82_SUMB_32__30_,
         u5_mult_82_SUMB_32__31_, u5_mult_82_SUMB_32__32_,
         u5_mult_82_SUMB_32__33_, u5_mult_82_SUMB_32__34_,
         u5_mult_82_SUMB_32__35_, u5_mult_82_SUMB_32__36_,
         u5_mult_82_SUMB_32__37_, u5_mult_82_SUMB_32__38_,
         u5_mult_82_SUMB_32__39_, u5_mult_82_SUMB_32__40_,
         u5_mult_82_SUMB_32__41_, u5_mult_82_SUMB_32__42_,
         u5_mult_82_SUMB_32__43_, u5_mult_82_SUMB_32__44_,
         u5_mult_82_SUMB_32__45_, u5_mult_82_SUMB_32__46_,
         u5_mult_82_SUMB_32__47_, u5_mult_82_SUMB_32__48_,
         u5_mult_82_SUMB_32__49_, u5_mult_82_SUMB_32__50_,
         u5_mult_82_SUMB_32__51_, u5_mult_82_SUMB_33__1_,
         u5_mult_82_SUMB_33__2_, u5_mult_82_SUMB_33__3_,
         u5_mult_82_SUMB_33__4_, u5_mult_82_SUMB_33__5_,
         u5_mult_82_SUMB_33__6_, u5_mult_82_SUMB_33__7_,
         u5_mult_82_SUMB_33__8_, u5_mult_82_SUMB_33__9_,
         u5_mult_82_SUMB_33__10_, u5_mult_82_SUMB_33__11_,
         u5_mult_82_SUMB_33__12_, u5_mult_82_SUMB_33__13_,
         u5_mult_82_SUMB_33__14_, u5_mult_82_SUMB_33__15_,
         u5_mult_82_SUMB_33__16_, u5_mult_82_SUMB_33__18_,
         u5_mult_82_SUMB_33__19_, u5_mult_82_SUMB_33__20_,
         u5_mult_82_SUMB_33__21_, u5_mult_82_SUMB_33__22_,
         u5_mult_82_SUMB_33__23_, u5_mult_82_SUMB_33__24_,
         u5_mult_82_SUMB_33__25_, u5_mult_82_SUMB_33__26_,
         u5_mult_82_SUMB_33__27_, u5_mult_82_SUMB_33__28_,
         u5_mult_82_SUMB_33__29_, u5_mult_82_SUMB_33__30_,
         u5_mult_82_SUMB_33__32_, u5_mult_82_SUMB_33__33_,
         u5_mult_82_SUMB_33__34_, u5_mult_82_SUMB_33__35_,
         u5_mult_82_CARRYB_24__1_, u5_mult_82_CARRYB_24__2_,
         u5_mult_82_CARRYB_24__3_, u5_mult_82_CARRYB_24__4_,
         u5_mult_82_CARRYB_24__5_, u5_mult_82_CARRYB_24__6_,
         u5_mult_82_CARRYB_24__7_, u5_mult_82_CARRYB_24__8_,
         u5_mult_82_CARRYB_24__9_, u5_mult_82_CARRYB_24__10_,
         u5_mult_82_CARRYB_24__11_, u5_mult_82_CARRYB_24__12_,
         u5_mult_82_CARRYB_24__13_, u5_mult_82_CARRYB_24__14_,
         u5_mult_82_CARRYB_24__15_, u5_mult_82_CARRYB_24__16_,
         u5_mult_82_CARRYB_24__17_, u5_mult_82_CARRYB_24__18_,
         u5_mult_82_CARRYB_24__19_, u5_mult_82_CARRYB_24__20_,
         u5_mult_82_CARRYB_24__21_, u5_mult_82_CARRYB_24__22_,
         u5_mult_82_CARRYB_24__23_, u5_mult_82_CARRYB_24__24_,
         u5_mult_82_CARRYB_24__25_, u5_mult_82_CARRYB_24__26_,
         u5_mult_82_CARRYB_24__27_, u5_mult_82_CARRYB_24__28_,
         u5_mult_82_CARRYB_24__29_, u5_mult_82_CARRYB_24__30_,
         u5_mult_82_CARRYB_24__31_, u5_mult_82_CARRYB_24__32_,
         u5_mult_82_CARRYB_24__33_, u5_mult_82_CARRYB_24__34_,
         u5_mult_82_CARRYB_24__35_, u5_mult_82_CARRYB_24__36_,
         u5_mult_82_CARRYB_24__37_, u5_mult_82_CARRYB_24__38_,
         u5_mult_82_CARRYB_24__39_, u5_mult_82_CARRYB_24__40_,
         u5_mult_82_CARRYB_24__41_, u5_mult_82_CARRYB_24__42_,
         u5_mult_82_CARRYB_24__43_, u5_mult_82_CARRYB_24__44_,
         u5_mult_82_CARRYB_24__45_, u5_mult_82_CARRYB_24__46_,
         u5_mult_82_CARRYB_24__47_, u5_mult_82_CARRYB_24__48_,
         u5_mult_82_CARRYB_24__49_, u5_mult_82_CARRYB_24__50_,
         u5_mult_82_CARRYB_24__51_, u5_mult_82_CARRYB_25__0_,
         u5_mult_82_CARRYB_25__1_, u5_mult_82_CARRYB_25__2_,
         u5_mult_82_CARRYB_25__3_, u5_mult_82_CARRYB_25__4_,
         u5_mult_82_CARRYB_25__5_, u5_mult_82_CARRYB_25__6_,
         u5_mult_82_CARRYB_25__7_, u5_mult_82_CARRYB_25__8_,
         u5_mult_82_CARRYB_25__9_, u5_mult_82_CARRYB_25__10_,
         u5_mult_82_CARRYB_25__11_, u5_mult_82_CARRYB_25__12_,
         u5_mult_82_CARRYB_25__13_, u5_mult_82_CARRYB_25__14_,
         u5_mult_82_CARRYB_25__15_, u5_mult_82_CARRYB_25__16_,
         u5_mult_82_CARRYB_25__17_, u5_mult_82_CARRYB_25__18_,
         u5_mult_82_CARRYB_25__19_, u5_mult_82_CARRYB_25__20_,
         u5_mult_82_CARRYB_25__21_, u5_mult_82_CARRYB_25__23_,
         u5_mult_82_CARRYB_25__24_, u5_mult_82_CARRYB_25__25_,
         u5_mult_82_CARRYB_25__26_, u5_mult_82_CARRYB_25__27_,
         u5_mult_82_CARRYB_25__28_, u5_mult_82_CARRYB_25__29_,
         u5_mult_82_CARRYB_25__30_, u5_mult_82_CARRYB_25__31_,
         u5_mult_82_CARRYB_25__32_, u5_mult_82_CARRYB_25__34_,
         u5_mult_82_CARRYB_25__35_, u5_mult_82_CARRYB_25__36_,
         u5_mult_82_CARRYB_25__37_, u5_mult_82_CARRYB_25__38_,
         u5_mult_82_CARRYB_25__39_, u5_mult_82_CARRYB_25__41_,
         u5_mult_82_CARRYB_25__42_, u5_mult_82_CARRYB_25__43_,
         u5_mult_82_CARRYB_25__44_, u5_mult_82_CARRYB_25__45_,
         u5_mult_82_CARRYB_25__46_, u5_mult_82_CARRYB_25__47_,
         u5_mult_82_CARRYB_25__48_, u5_mult_82_CARRYB_25__49_,
         u5_mult_82_CARRYB_25__50_, u5_mult_82_CARRYB_25__51_,
         u5_mult_82_CARRYB_26__0_, u5_mult_82_CARRYB_26__1_,
         u5_mult_82_CARRYB_26__2_, u5_mult_82_CARRYB_26__3_,
         u5_mult_82_CARRYB_26__4_, u5_mult_82_CARRYB_26__5_,
         u5_mult_82_CARRYB_26__6_, u5_mult_82_CARRYB_26__7_,
         u5_mult_82_CARRYB_26__8_, u5_mult_82_CARRYB_26__9_,
         u5_mult_82_CARRYB_26__10_, u5_mult_82_CARRYB_26__11_,
         u5_mult_82_CARRYB_26__12_, u5_mult_82_CARRYB_26__13_,
         u5_mult_82_CARRYB_26__14_, u5_mult_82_CARRYB_26__15_,
         u5_mult_82_CARRYB_26__16_, u5_mult_82_CARRYB_26__17_,
         u5_mult_82_CARRYB_26__18_, u5_mult_82_CARRYB_26__19_,
         u5_mult_82_CARRYB_26__20_, u5_mult_82_CARRYB_26__22_,
         u5_mult_82_CARRYB_26__23_, u5_mult_82_CARRYB_26__24_,
         u5_mult_82_CARRYB_26__25_, u5_mult_82_CARRYB_26__26_,
         u5_mult_82_CARRYB_26__27_, u5_mult_82_CARRYB_26__28_,
         u5_mult_82_CARRYB_26__29_, u5_mult_82_CARRYB_26__30_,
         u5_mult_82_CARRYB_26__31_, u5_mult_82_CARRYB_26__32_,
         u5_mult_82_CARRYB_26__33_, u5_mult_82_CARRYB_26__34_,
         u5_mult_82_CARRYB_26__35_, u5_mult_82_CARRYB_26__36_,
         u5_mult_82_CARRYB_26__37_, u5_mult_82_CARRYB_26__38_,
         u5_mult_82_CARRYB_26__39_, u5_mult_82_CARRYB_26__40_,
         u5_mult_82_CARRYB_26__41_, u5_mult_82_CARRYB_26__42_,
         u5_mult_82_CARRYB_26__43_, u5_mult_82_CARRYB_26__44_,
         u5_mult_82_CARRYB_26__45_, u5_mult_82_CARRYB_26__46_,
         u5_mult_82_CARRYB_26__47_, u5_mult_82_CARRYB_26__48_,
         u5_mult_82_CARRYB_26__49_, u5_mult_82_CARRYB_26__50_,
         u5_mult_82_CARRYB_26__51_, u5_mult_82_CARRYB_27__0_,
         u5_mult_82_CARRYB_27__1_, u5_mult_82_CARRYB_27__2_,
         u5_mult_82_CARRYB_27__3_, u5_mult_82_CARRYB_27__4_,
         u5_mult_82_CARRYB_27__5_, u5_mult_82_CARRYB_27__6_,
         u5_mult_82_CARRYB_27__7_, u5_mult_82_CARRYB_27__8_,
         u5_mult_82_CARRYB_27__9_, u5_mult_82_CARRYB_27__10_,
         u5_mult_82_CARRYB_27__11_, u5_mult_82_CARRYB_27__12_,
         u5_mult_82_CARRYB_27__13_, u5_mult_82_CARRYB_27__14_,
         u5_mult_82_CARRYB_27__15_, u5_mult_82_CARRYB_27__16_,
         u5_mult_82_CARRYB_27__17_, u5_mult_82_CARRYB_27__18_,
         u5_mult_82_CARRYB_27__19_, u5_mult_82_CARRYB_27__21_,
         u5_mult_82_CARRYB_27__22_, u5_mult_82_CARRYB_27__23_,
         u5_mult_82_CARRYB_27__24_, u5_mult_82_CARRYB_27__25_,
         u5_mult_82_CARRYB_27__26_, u5_mult_82_CARRYB_27__27_,
         u5_mult_82_CARRYB_27__28_, u5_mult_82_CARRYB_27__29_,
         u5_mult_82_CARRYB_27__30_, u5_mult_82_CARRYB_27__31_,
         u5_mult_82_CARRYB_27__32_, u5_mult_82_CARRYB_27__33_,
         u5_mult_82_CARRYB_27__34_, u5_mult_82_CARRYB_27__35_,
         u5_mult_82_CARRYB_27__36_, u5_mult_82_CARRYB_27__37_,
         u5_mult_82_CARRYB_27__38_, u5_mult_82_CARRYB_27__39_,
         u5_mult_82_CARRYB_27__40_, u5_mult_82_CARRYB_27__41_,
         u5_mult_82_CARRYB_27__42_, u5_mult_82_CARRYB_27__43_,
         u5_mult_82_CARRYB_27__44_, u5_mult_82_CARRYB_27__45_,
         u5_mult_82_CARRYB_27__46_, u5_mult_82_CARRYB_27__47_,
         u5_mult_82_CARRYB_27__48_, u5_mult_82_CARRYB_27__49_,
         u5_mult_82_CARRYB_27__50_, u5_mult_82_CARRYB_27__51_,
         u5_mult_82_CARRYB_28__0_, u5_mult_82_CARRYB_28__1_,
         u5_mult_82_CARRYB_28__2_, u5_mult_82_CARRYB_28__3_,
         u5_mult_82_CARRYB_28__4_, u5_mult_82_CARRYB_28__5_,
         u5_mult_82_CARRYB_28__6_, u5_mult_82_CARRYB_28__7_,
         u5_mult_82_CARRYB_28__8_, u5_mult_82_CARRYB_28__9_,
         u5_mult_82_CARRYB_28__10_, u5_mult_82_CARRYB_28__11_,
         u5_mult_82_CARRYB_28__12_, u5_mult_82_CARRYB_28__13_,
         u5_mult_82_CARRYB_28__14_, u5_mult_82_CARRYB_28__15_,
         u5_mult_82_CARRYB_28__16_, u5_mult_82_CARRYB_28__17_,
         u5_mult_82_CARRYB_28__18_, u5_mult_82_CARRYB_28__19_,
         u5_mult_82_CARRYB_28__21_, u5_mult_82_CARRYB_28__22_,
         u5_mult_82_CARRYB_28__23_, u5_mult_82_CARRYB_28__24_,
         u5_mult_82_CARRYB_28__25_, u5_mult_82_CARRYB_28__26_,
         u5_mult_82_CARRYB_28__27_, u5_mult_82_CARRYB_28__28_,
         u5_mult_82_CARRYB_28__29_, u5_mult_82_CARRYB_28__30_,
         u5_mult_82_CARRYB_28__31_, u5_mult_82_CARRYB_28__32_,
         u5_mult_82_CARRYB_28__33_, u5_mult_82_CARRYB_28__34_,
         u5_mult_82_CARRYB_28__35_, u5_mult_82_CARRYB_28__36_,
         u5_mult_82_CARRYB_28__37_, u5_mult_82_CARRYB_28__38_,
         u5_mult_82_CARRYB_28__39_, u5_mult_82_CARRYB_28__40_,
         u5_mult_82_CARRYB_28__41_, u5_mult_82_CARRYB_28__42_,
         u5_mult_82_CARRYB_28__43_, u5_mult_82_CARRYB_28__44_,
         u5_mult_82_CARRYB_28__45_, u5_mult_82_CARRYB_28__46_,
         u5_mult_82_CARRYB_28__47_, u5_mult_82_CARRYB_28__48_,
         u5_mult_82_CARRYB_28__49_, u5_mult_82_CARRYB_28__50_,
         u5_mult_82_CARRYB_28__51_, u5_mult_82_CARRYB_29__0_,
         u5_mult_82_CARRYB_29__1_, u5_mult_82_CARRYB_29__2_,
         u5_mult_82_CARRYB_29__3_, u5_mult_82_CARRYB_29__4_,
         u5_mult_82_CARRYB_29__5_, u5_mult_82_CARRYB_29__6_,
         u5_mult_82_CARRYB_29__7_, u5_mult_82_CARRYB_29__8_,
         u5_mult_82_CARRYB_29__9_, u5_mult_82_CARRYB_29__10_,
         u5_mult_82_CARRYB_29__11_, u5_mult_82_CARRYB_29__12_,
         u5_mult_82_CARRYB_29__13_, u5_mult_82_CARRYB_29__14_,
         u5_mult_82_CARRYB_29__15_, u5_mult_82_CARRYB_29__16_,
         u5_mult_82_CARRYB_29__17_, u5_mult_82_CARRYB_29__18_,
         u5_mult_82_CARRYB_29__20_, u5_mult_82_CARRYB_29__21_,
         u5_mult_82_CARRYB_29__22_, u5_mult_82_CARRYB_29__23_,
         u5_mult_82_CARRYB_29__24_, u5_mult_82_CARRYB_29__25_,
         u5_mult_82_CARRYB_29__26_, u5_mult_82_CARRYB_29__27_,
         u5_mult_82_CARRYB_29__28_, u5_mult_82_CARRYB_29__29_,
         u5_mult_82_CARRYB_29__30_, u5_mult_82_CARRYB_29__31_,
         u5_mult_82_CARRYB_29__32_, u5_mult_82_CARRYB_29__33_,
         u5_mult_82_CARRYB_29__34_, u5_mult_82_CARRYB_29__35_,
         u5_mult_82_CARRYB_29__36_, u5_mult_82_CARRYB_29__37_,
         u5_mult_82_CARRYB_29__38_, u5_mult_82_CARRYB_29__39_,
         u5_mult_82_CARRYB_29__40_, u5_mult_82_CARRYB_29__41_,
         u5_mult_82_CARRYB_29__42_, u5_mult_82_CARRYB_29__43_,
         u5_mult_82_CARRYB_29__44_, u5_mult_82_CARRYB_29__45_,
         u5_mult_82_CARRYB_29__46_, u5_mult_82_CARRYB_29__47_,
         u5_mult_82_CARRYB_29__48_, u5_mult_82_CARRYB_29__49_,
         u5_mult_82_CARRYB_29__50_, u5_mult_82_CARRYB_29__51_,
         u5_mult_82_CARRYB_30__0_, u5_mult_82_CARRYB_30__1_,
         u5_mult_82_CARRYB_30__2_, u5_mult_82_CARRYB_30__3_,
         u5_mult_82_CARRYB_30__4_, u5_mult_82_CARRYB_30__5_,
         u5_mult_82_CARRYB_30__6_, u5_mult_82_CARRYB_30__7_,
         u5_mult_82_CARRYB_30__8_, u5_mult_82_CARRYB_30__9_,
         u5_mult_82_CARRYB_30__10_, u5_mult_82_CARRYB_30__11_,
         u5_mult_82_CARRYB_30__12_, u5_mult_82_CARRYB_30__13_,
         u5_mult_82_CARRYB_30__14_, u5_mult_82_CARRYB_30__15_,
         u5_mult_82_CARRYB_30__16_, u5_mult_82_CARRYB_30__17_,
         u5_mult_82_CARRYB_30__19_, u5_mult_82_CARRYB_30__20_,
         u5_mult_82_CARRYB_30__21_, u5_mult_82_CARRYB_30__22_,
         u5_mult_82_CARRYB_30__23_, u5_mult_82_CARRYB_30__24_,
         u5_mult_82_CARRYB_30__25_, u5_mult_82_CARRYB_30__26_,
         u5_mult_82_CARRYB_30__27_, u5_mult_82_CARRYB_30__28_,
         u5_mult_82_CARRYB_30__29_, u5_mult_82_CARRYB_30__30_,
         u5_mult_82_CARRYB_30__31_, u5_mult_82_CARRYB_30__32_,
         u5_mult_82_CARRYB_30__33_, u5_mult_82_CARRYB_30__34_,
         u5_mult_82_CARRYB_30__35_, u5_mult_82_CARRYB_30__36_,
         u5_mult_82_CARRYB_30__37_, u5_mult_82_CARRYB_30__38_,
         u5_mult_82_CARRYB_30__39_, u5_mult_82_CARRYB_30__40_,
         u5_mult_82_CARRYB_30__41_, u5_mult_82_CARRYB_30__42_,
         u5_mult_82_CARRYB_30__43_, u5_mult_82_CARRYB_30__44_,
         u5_mult_82_CARRYB_30__45_, u5_mult_82_CARRYB_30__46_,
         u5_mult_82_CARRYB_30__47_, u5_mult_82_CARRYB_30__48_,
         u5_mult_82_CARRYB_30__49_, u5_mult_82_CARRYB_30__50_,
         u5_mult_82_CARRYB_30__51_, u5_mult_82_CARRYB_31__0_,
         u5_mult_82_CARRYB_31__1_, u5_mult_82_CARRYB_31__2_,
         u5_mult_82_CARRYB_31__3_, u5_mult_82_CARRYB_31__4_,
         u5_mult_82_CARRYB_31__5_, u5_mult_82_CARRYB_31__6_,
         u5_mult_82_CARRYB_31__7_, u5_mult_82_CARRYB_31__8_,
         u5_mult_82_CARRYB_31__9_, u5_mult_82_CARRYB_31__10_,
         u5_mult_82_CARRYB_31__11_, u5_mult_82_CARRYB_31__12_,
         u5_mult_82_CARRYB_31__13_, u5_mult_82_CARRYB_31__14_,
         u5_mult_82_CARRYB_31__15_, u5_mult_82_CARRYB_31__16_,
         u5_mult_82_CARRYB_31__17_, u5_mult_82_CARRYB_31__18_,
         u5_mult_82_CARRYB_31__19_, u5_mult_82_CARRYB_31__20_,
         u5_mult_82_CARRYB_31__21_, u5_mult_82_CARRYB_31__22_,
         u5_mult_82_CARRYB_31__23_, u5_mult_82_CARRYB_31__24_,
         u5_mult_82_CARRYB_31__25_, u5_mult_82_CARRYB_31__26_,
         u5_mult_82_CARRYB_31__27_, u5_mult_82_CARRYB_31__28_,
         u5_mult_82_CARRYB_31__29_, u5_mult_82_CARRYB_31__30_,
         u5_mult_82_CARRYB_31__31_, u5_mult_82_CARRYB_31__32_,
         u5_mult_82_CARRYB_31__33_, u5_mult_82_CARRYB_31__34_,
         u5_mult_82_CARRYB_31__35_, u5_mult_82_CARRYB_31__36_,
         u5_mult_82_CARRYB_31__37_, u5_mult_82_CARRYB_31__38_,
         u5_mult_82_CARRYB_31__39_, u5_mult_82_CARRYB_31__40_,
         u5_mult_82_CARRYB_31__41_, u5_mult_82_CARRYB_31__42_,
         u5_mult_82_CARRYB_31__43_, u5_mult_82_CARRYB_31__44_,
         u5_mult_82_CARRYB_31__45_, u5_mult_82_CARRYB_31__46_,
         u5_mult_82_CARRYB_31__47_, u5_mult_82_CARRYB_31__48_,
         u5_mult_82_CARRYB_31__49_, u5_mult_82_CARRYB_31__50_,
         u5_mult_82_CARRYB_31__51_, u5_mult_82_CARRYB_32__0_,
         u5_mult_82_CARRYB_32__1_, u5_mult_82_CARRYB_32__2_,
         u5_mult_82_CARRYB_32__3_, u5_mult_82_CARRYB_32__4_,
         u5_mult_82_CARRYB_32__5_, u5_mult_82_CARRYB_32__6_,
         u5_mult_82_CARRYB_32__7_, u5_mult_82_CARRYB_32__8_,
         u5_mult_82_CARRYB_32__9_, u5_mult_82_CARRYB_32__10_,
         u5_mult_82_CARRYB_32__11_, u5_mult_82_CARRYB_32__12_,
         u5_mult_82_CARRYB_32__13_, u5_mult_82_CARRYB_32__14_,
         u5_mult_82_CARRYB_32__15_, u5_mult_82_CARRYB_32__16_,
         u5_mult_82_CARRYB_32__17_, u5_mult_82_CARRYB_32__18_,
         u5_mult_82_CARRYB_32__19_, u5_mult_82_CARRYB_32__20_,
         u5_mult_82_CARRYB_32__21_, u5_mult_82_CARRYB_32__22_,
         u5_mult_82_CARRYB_32__23_, u5_mult_82_CARRYB_32__24_,
         u5_mult_82_CARRYB_32__25_, u5_mult_82_CARRYB_32__26_,
         u5_mult_82_CARRYB_32__27_, u5_mult_82_CARRYB_32__28_,
         u5_mult_82_CARRYB_32__29_, u5_mult_82_CARRYB_32__30_,
         u5_mult_82_CARRYB_32__31_, u5_mult_82_CARRYB_32__32_,
         u5_mult_82_CARRYB_32__33_, u5_mult_82_CARRYB_32__34_,
         u5_mult_82_CARRYB_32__35_, u5_mult_82_CARRYB_32__36_,
         u5_mult_82_CARRYB_32__37_, u5_mult_82_CARRYB_32__38_,
         u5_mult_82_CARRYB_32__39_, u5_mult_82_CARRYB_32__40_,
         u5_mult_82_CARRYB_32__41_, u5_mult_82_CARRYB_32__42_,
         u5_mult_82_CARRYB_32__43_, u5_mult_82_CARRYB_32__44_,
         u5_mult_82_CARRYB_32__45_, u5_mult_82_CARRYB_32__46_,
         u5_mult_82_CARRYB_32__47_, u5_mult_82_CARRYB_32__48_,
         u5_mult_82_CARRYB_32__49_, u5_mult_82_CARRYB_32__50_,
         u5_mult_82_CARRYB_32__51_, u5_mult_82_CARRYB_33__0_,
         u5_mult_82_CARRYB_33__1_, u5_mult_82_CARRYB_33__2_,
         u5_mult_82_CARRYB_33__3_, u5_mult_82_CARRYB_33__4_,
         u5_mult_82_CARRYB_33__5_, u5_mult_82_CARRYB_33__6_,
         u5_mult_82_CARRYB_33__7_, u5_mult_82_CARRYB_33__8_,
         u5_mult_82_CARRYB_33__9_, u5_mult_82_CARRYB_33__10_,
         u5_mult_82_CARRYB_33__11_, u5_mult_82_CARRYB_33__12_,
         u5_mult_82_CARRYB_33__13_, u5_mult_82_CARRYB_33__14_,
         u5_mult_82_CARRYB_33__15_, u5_mult_82_CARRYB_33__16_,
         u5_mult_82_CARRYB_33__17_, u5_mult_82_CARRYB_33__18_,
         u5_mult_82_CARRYB_33__19_, u5_mult_82_CARRYB_33__20_,
         u5_mult_82_CARRYB_33__21_, u5_mult_82_CARRYB_33__22_,
         u5_mult_82_CARRYB_33__23_, u5_mult_82_CARRYB_33__24_,
         u5_mult_82_CARRYB_33__25_, u5_mult_82_CARRYB_33__26_,
         u5_mult_82_CARRYB_33__27_, u5_mult_82_CARRYB_33__28_,
         u5_mult_82_CARRYB_33__29_, u5_mult_82_CARRYB_33__30_,
         u5_mult_82_CARRYB_33__31_, u5_mult_82_CARRYB_33__32_,
         u5_mult_82_CARRYB_33__33_, u5_mult_82_CARRYB_33__34_,
         u5_mult_82_CARRYB_33__35_, u5_mult_82_SUMB_14__19_,
         u5_mult_82_SUMB_14__20_, u5_mult_82_SUMB_14__21_,
         u5_mult_82_SUMB_14__22_, u5_mult_82_SUMB_14__23_,
         u5_mult_82_SUMB_14__24_, u5_mult_82_SUMB_14__25_,
         u5_mult_82_SUMB_14__26_, u5_mult_82_SUMB_14__27_,
         u5_mult_82_SUMB_14__29_, u5_mult_82_SUMB_14__30_,
         u5_mult_82_SUMB_14__31_, u5_mult_82_SUMB_14__32_,
         u5_mult_82_SUMB_14__33_, u5_mult_82_SUMB_14__34_,
         u5_mult_82_SUMB_14__35_, u5_mult_82_SUMB_14__36_,
         u5_mult_82_SUMB_14__37_, u5_mult_82_SUMB_14__38_,
         u5_mult_82_SUMB_14__39_, u5_mult_82_SUMB_14__40_,
         u5_mult_82_SUMB_14__41_, u5_mult_82_SUMB_14__42_,
         u5_mult_82_SUMB_14__43_, u5_mult_82_SUMB_14__44_,
         u5_mult_82_SUMB_14__45_, u5_mult_82_SUMB_14__46_,
         u5_mult_82_SUMB_14__47_, u5_mult_82_SUMB_14__48_,
         u5_mult_82_SUMB_14__49_, u5_mult_82_SUMB_14__50_,
         u5_mult_82_SUMB_14__51_, u5_mult_82_SUMB_15__1_,
         u5_mult_82_SUMB_15__2_, u5_mult_82_SUMB_15__3_,
         u5_mult_82_SUMB_15__4_, u5_mult_82_SUMB_15__5_,
         u5_mult_82_SUMB_15__6_, u5_mult_82_SUMB_15__7_,
         u5_mult_82_SUMB_15__8_, u5_mult_82_SUMB_15__9_,
         u5_mult_82_SUMB_15__10_, u5_mult_82_SUMB_15__11_,
         u5_mult_82_SUMB_15__12_, u5_mult_82_SUMB_15__13_,
         u5_mult_82_SUMB_15__14_, u5_mult_82_SUMB_15__15_,
         u5_mult_82_SUMB_15__16_, u5_mult_82_SUMB_15__17_,
         u5_mult_82_SUMB_15__18_, u5_mult_82_SUMB_15__19_,
         u5_mult_82_SUMB_15__20_, u5_mult_82_SUMB_15__21_,
         u5_mult_82_SUMB_15__22_, u5_mult_82_SUMB_15__23_,
         u5_mult_82_SUMB_15__24_, u5_mult_82_SUMB_15__25_,
         u5_mult_82_SUMB_15__26_, u5_mult_82_SUMB_15__28_,
         u5_mult_82_SUMB_15__30_, u5_mult_82_SUMB_15__31_,
         u5_mult_82_SUMB_15__32_, u5_mult_82_SUMB_15__33_,
         u5_mult_82_SUMB_15__34_, u5_mult_82_SUMB_15__35_,
         u5_mult_82_SUMB_15__36_, u5_mult_82_SUMB_15__38_,
         u5_mult_82_SUMB_15__39_, u5_mult_82_SUMB_15__40_,
         u5_mult_82_SUMB_15__41_, u5_mult_82_SUMB_15__42_,
         u5_mult_82_SUMB_15__43_, u5_mult_82_SUMB_15__44_,
         u5_mult_82_SUMB_15__45_, u5_mult_82_SUMB_15__46_,
         u5_mult_82_SUMB_15__47_, u5_mult_82_SUMB_15__48_,
         u5_mult_82_SUMB_15__49_, u5_mult_82_SUMB_15__50_,
         u5_mult_82_SUMB_15__51_, u5_mult_82_SUMB_16__1_,
         u5_mult_82_SUMB_16__2_, u5_mult_82_SUMB_16__3_,
         u5_mult_82_SUMB_16__4_, u5_mult_82_SUMB_16__5_,
         u5_mult_82_SUMB_16__6_, u5_mult_82_SUMB_16__7_,
         u5_mult_82_SUMB_16__8_, u5_mult_82_SUMB_16__9_,
         u5_mult_82_SUMB_16__10_, u5_mult_82_SUMB_16__11_,
         u5_mult_82_SUMB_16__12_, u5_mult_82_SUMB_16__13_,
         u5_mult_82_SUMB_16__14_, u5_mult_82_SUMB_16__15_,
         u5_mult_82_SUMB_16__16_, u5_mult_82_SUMB_16__17_,
         u5_mult_82_SUMB_16__18_, u5_mult_82_SUMB_16__19_,
         u5_mult_82_SUMB_16__20_, u5_mult_82_SUMB_16__21_,
         u5_mult_82_SUMB_16__22_, u5_mult_82_SUMB_16__23_,
         u5_mult_82_SUMB_16__24_, u5_mult_82_SUMB_16__25_,
         u5_mult_82_SUMB_16__26_, u5_mult_82_SUMB_16__27_,
         u5_mult_82_SUMB_16__29_, u5_mult_82_SUMB_16__30_,
         u5_mult_82_SUMB_16__31_, u5_mult_82_SUMB_16__32_,
         u5_mult_82_SUMB_16__33_, u5_mult_82_SUMB_16__34_,
         u5_mult_82_SUMB_16__35_, u5_mult_82_SUMB_16__36_,
         u5_mult_82_SUMB_16__37_, u5_mult_82_SUMB_16__38_,
         u5_mult_82_SUMB_16__39_, u5_mult_82_SUMB_16__40_,
         u5_mult_82_SUMB_16__41_, u5_mult_82_SUMB_16__42_,
         u5_mult_82_SUMB_16__43_, u5_mult_82_SUMB_16__44_,
         u5_mult_82_SUMB_16__45_, u5_mult_82_SUMB_16__46_,
         u5_mult_82_SUMB_16__47_, u5_mult_82_SUMB_16__48_,
         u5_mult_82_SUMB_16__49_, u5_mult_82_SUMB_16__50_,
         u5_mult_82_SUMB_16__51_, u5_mult_82_SUMB_17__1_,
         u5_mult_82_SUMB_17__2_, u5_mult_82_SUMB_17__3_,
         u5_mult_82_SUMB_17__4_, u5_mult_82_SUMB_17__5_,
         u5_mult_82_SUMB_17__6_, u5_mult_82_SUMB_17__7_,
         u5_mult_82_SUMB_17__8_, u5_mult_82_SUMB_17__9_,
         u5_mult_82_SUMB_17__10_, u5_mult_82_SUMB_17__11_,
         u5_mult_82_SUMB_17__12_, u5_mult_82_SUMB_17__13_,
         u5_mult_82_SUMB_17__14_, u5_mult_82_SUMB_17__15_,
         u5_mult_82_SUMB_17__16_, u5_mult_82_SUMB_17__17_,
         u5_mult_82_SUMB_17__18_, u5_mult_82_SUMB_17__19_,
         u5_mult_82_SUMB_17__20_, u5_mult_82_SUMB_17__21_,
         u5_mult_82_SUMB_17__22_, u5_mult_82_SUMB_17__23_,
         u5_mult_82_SUMB_17__24_, u5_mult_82_SUMB_17__25_,
         u5_mult_82_SUMB_17__26_, u5_mult_82_SUMB_17__28_,
         u5_mult_82_SUMB_17__29_, u5_mult_82_SUMB_17__30_,
         u5_mult_82_SUMB_17__31_, u5_mult_82_SUMB_17__32_,
         u5_mult_82_SUMB_17__33_, u5_mult_82_SUMB_17__34_,
         u5_mult_82_SUMB_17__35_, u5_mult_82_SUMB_17__36_,
         u5_mult_82_SUMB_17__37_, u5_mult_82_SUMB_17__38_,
         u5_mult_82_SUMB_17__39_, u5_mult_82_SUMB_17__40_,
         u5_mult_82_SUMB_17__41_, u5_mult_82_SUMB_17__42_,
         u5_mult_82_SUMB_17__43_, u5_mult_82_SUMB_17__44_,
         u5_mult_82_SUMB_17__45_, u5_mult_82_SUMB_17__46_,
         u5_mult_82_SUMB_17__47_, u5_mult_82_SUMB_17__48_,
         u5_mult_82_SUMB_17__49_, u5_mult_82_SUMB_17__50_,
         u5_mult_82_SUMB_17__51_, u5_mult_82_SUMB_18__1_,
         u5_mult_82_SUMB_18__2_, u5_mult_82_SUMB_18__3_,
         u5_mult_82_SUMB_18__4_, u5_mult_82_SUMB_18__5_,
         u5_mult_82_SUMB_18__6_, u5_mult_82_SUMB_18__7_,
         u5_mult_82_SUMB_18__8_, u5_mult_82_SUMB_18__9_,
         u5_mult_82_SUMB_18__10_, u5_mult_82_SUMB_18__11_,
         u5_mult_82_SUMB_18__12_, u5_mult_82_SUMB_18__13_,
         u5_mult_82_SUMB_18__14_, u5_mult_82_SUMB_18__15_,
         u5_mult_82_SUMB_18__16_, u5_mult_82_SUMB_18__17_,
         u5_mult_82_SUMB_18__18_, u5_mult_82_SUMB_18__19_,
         u5_mult_82_SUMB_18__20_, u5_mult_82_SUMB_18__21_,
         u5_mult_82_SUMB_18__22_, u5_mult_82_SUMB_18__23_,
         u5_mult_82_SUMB_18__24_, u5_mult_82_SUMB_18__25_,
         u5_mult_82_SUMB_18__28_, u5_mult_82_SUMB_18__29_,
         u5_mult_82_SUMB_18__30_, u5_mult_82_SUMB_18__31_,
         u5_mult_82_SUMB_18__32_, u5_mult_82_SUMB_18__33_,
         u5_mult_82_SUMB_18__34_, u5_mult_82_SUMB_18__35_,
         u5_mult_82_SUMB_18__36_, u5_mult_82_SUMB_18__37_,
         u5_mult_82_SUMB_18__38_, u5_mult_82_SUMB_18__39_,
         u5_mult_82_SUMB_18__40_, u5_mult_82_SUMB_18__41_,
         u5_mult_82_SUMB_18__42_, u5_mult_82_SUMB_18__43_,
         u5_mult_82_SUMB_18__44_, u5_mult_82_SUMB_18__45_,
         u5_mult_82_SUMB_18__46_, u5_mult_82_SUMB_18__47_,
         u5_mult_82_SUMB_18__48_, u5_mult_82_SUMB_18__49_,
         u5_mult_82_SUMB_18__50_, u5_mult_82_SUMB_18__51_,
         u5_mult_82_SUMB_19__1_, u5_mult_82_SUMB_19__2_,
         u5_mult_82_SUMB_19__3_, u5_mult_82_SUMB_19__4_,
         u5_mult_82_SUMB_19__5_, u5_mult_82_SUMB_19__6_,
         u5_mult_82_SUMB_19__7_, u5_mult_82_SUMB_19__8_,
         u5_mult_82_SUMB_19__9_, u5_mult_82_SUMB_19__10_,
         u5_mult_82_SUMB_19__11_, u5_mult_82_SUMB_19__12_,
         u5_mult_82_SUMB_19__13_, u5_mult_82_SUMB_19__14_,
         u5_mult_82_SUMB_19__15_, u5_mult_82_SUMB_19__16_,
         u5_mult_82_SUMB_19__17_, u5_mult_82_SUMB_19__18_,
         u5_mult_82_SUMB_19__19_, u5_mult_82_SUMB_19__20_,
         u5_mult_82_SUMB_19__21_, u5_mult_82_SUMB_19__22_,
         u5_mult_82_SUMB_19__23_, u5_mult_82_SUMB_19__24_,
         u5_mult_82_SUMB_19__25_, u5_mult_82_SUMB_19__27_,
         u5_mult_82_SUMB_19__28_, u5_mult_82_SUMB_19__29_,
         u5_mult_82_SUMB_19__30_, u5_mult_82_SUMB_19__31_,
         u5_mult_82_SUMB_19__32_, u5_mult_82_SUMB_19__33_,
         u5_mult_82_SUMB_19__34_, u5_mult_82_SUMB_19__35_,
         u5_mult_82_SUMB_19__36_, u5_mult_82_SUMB_19__37_,
         u5_mult_82_SUMB_19__38_, u5_mult_82_SUMB_19__39_,
         u5_mult_82_SUMB_19__40_, u5_mult_82_SUMB_19__41_,
         u5_mult_82_SUMB_19__42_, u5_mult_82_SUMB_19__43_,
         u5_mult_82_SUMB_19__44_, u5_mult_82_SUMB_19__45_,
         u5_mult_82_SUMB_19__46_, u5_mult_82_SUMB_19__47_,
         u5_mult_82_SUMB_19__48_, u5_mult_82_SUMB_19__49_,
         u5_mult_82_SUMB_19__50_, u5_mult_82_SUMB_19__51_,
         u5_mult_82_SUMB_20__1_, u5_mult_82_SUMB_20__2_,
         u5_mult_82_SUMB_20__3_, u5_mult_82_SUMB_20__4_,
         u5_mult_82_SUMB_20__5_, u5_mult_82_SUMB_20__6_,
         u5_mult_82_SUMB_20__7_, u5_mult_82_SUMB_20__8_,
         u5_mult_82_SUMB_20__9_, u5_mult_82_SUMB_20__10_,
         u5_mult_82_SUMB_20__11_, u5_mult_82_SUMB_20__12_,
         u5_mult_82_SUMB_20__13_, u5_mult_82_SUMB_20__14_,
         u5_mult_82_SUMB_20__15_, u5_mult_82_SUMB_20__16_,
         u5_mult_82_SUMB_20__17_, u5_mult_82_SUMB_20__18_,
         u5_mult_82_SUMB_20__19_, u5_mult_82_SUMB_20__20_,
         u5_mult_82_SUMB_20__21_, u5_mult_82_SUMB_20__22_,
         u5_mult_82_SUMB_20__23_, u5_mult_82_SUMB_20__24_,
         u5_mult_82_SUMB_20__26_, u5_mult_82_SUMB_20__27_,
         u5_mult_82_SUMB_20__28_, u5_mult_82_SUMB_20__29_,
         u5_mult_82_SUMB_20__30_, u5_mult_82_SUMB_20__31_,
         u5_mult_82_SUMB_20__32_, u5_mult_82_SUMB_20__33_,
         u5_mult_82_SUMB_20__34_, u5_mult_82_SUMB_20__35_,
         u5_mult_82_SUMB_20__36_, u5_mult_82_SUMB_20__37_,
         u5_mult_82_SUMB_20__38_, u5_mult_82_SUMB_20__39_,
         u5_mult_82_SUMB_20__40_, u5_mult_82_SUMB_20__41_,
         u5_mult_82_SUMB_20__42_, u5_mult_82_SUMB_20__43_,
         u5_mult_82_SUMB_20__44_, u5_mult_82_SUMB_20__45_,
         u5_mult_82_SUMB_20__46_, u5_mult_82_SUMB_20__47_,
         u5_mult_82_SUMB_20__48_, u5_mult_82_SUMB_20__49_,
         u5_mult_82_SUMB_20__50_, u5_mult_82_SUMB_20__51_,
         u5_mult_82_SUMB_21__1_, u5_mult_82_SUMB_21__2_,
         u5_mult_82_SUMB_21__3_, u5_mult_82_SUMB_21__4_,
         u5_mult_82_SUMB_21__5_, u5_mult_82_SUMB_21__6_,
         u5_mult_82_SUMB_21__7_, u5_mult_82_SUMB_21__8_,
         u5_mult_82_SUMB_21__9_, u5_mult_82_SUMB_21__10_,
         u5_mult_82_SUMB_21__11_, u5_mult_82_SUMB_21__12_,
         u5_mult_82_SUMB_21__13_, u5_mult_82_SUMB_21__14_,
         u5_mult_82_SUMB_21__15_, u5_mult_82_SUMB_21__16_,
         u5_mult_82_SUMB_21__17_, u5_mult_82_SUMB_21__18_,
         u5_mult_82_SUMB_21__19_, u5_mult_82_SUMB_21__20_,
         u5_mult_82_SUMB_21__21_, u5_mult_82_SUMB_21__22_,
         u5_mult_82_SUMB_21__23_, u5_mult_82_SUMB_21__24_,
         u5_mult_82_SUMB_21__25_, u5_mult_82_SUMB_21__26_,
         u5_mult_82_SUMB_21__27_, u5_mult_82_SUMB_21__28_,
         u5_mult_82_SUMB_21__29_, u5_mult_82_SUMB_21__30_,
         u5_mult_82_SUMB_21__31_, u5_mult_82_SUMB_21__32_,
         u5_mult_82_SUMB_21__33_, u5_mult_82_SUMB_21__34_,
         u5_mult_82_SUMB_21__35_, u5_mult_82_SUMB_21__36_,
         u5_mult_82_SUMB_21__37_, u5_mult_82_SUMB_21__38_,
         u5_mult_82_SUMB_21__39_, u5_mult_82_SUMB_21__40_,
         u5_mult_82_SUMB_21__41_, u5_mult_82_SUMB_21__42_,
         u5_mult_82_SUMB_21__43_, u5_mult_82_SUMB_21__44_,
         u5_mult_82_SUMB_21__45_, u5_mult_82_SUMB_21__46_,
         u5_mult_82_SUMB_21__47_, u5_mult_82_SUMB_21__48_,
         u5_mult_82_SUMB_21__49_, u5_mult_82_SUMB_21__50_,
         u5_mult_82_SUMB_21__51_, u5_mult_82_SUMB_22__1_,
         u5_mult_82_SUMB_22__2_, u5_mult_82_SUMB_22__3_,
         u5_mult_82_SUMB_22__4_, u5_mult_82_SUMB_22__5_,
         u5_mult_82_SUMB_22__6_, u5_mult_82_SUMB_22__7_,
         u5_mult_82_SUMB_22__8_, u5_mult_82_SUMB_22__9_,
         u5_mult_82_SUMB_22__10_, u5_mult_82_SUMB_22__11_,
         u5_mult_82_SUMB_22__12_, u5_mult_82_SUMB_22__13_,
         u5_mult_82_SUMB_22__14_, u5_mult_82_SUMB_22__15_,
         u5_mult_82_SUMB_22__16_, u5_mult_82_SUMB_22__17_,
         u5_mult_82_SUMB_22__18_, u5_mult_82_SUMB_22__19_,
         u5_mult_82_SUMB_22__20_, u5_mult_82_SUMB_22__21_,
         u5_mult_82_SUMB_22__22_, u5_mult_82_SUMB_22__23_,
         u5_mult_82_SUMB_22__25_, u5_mult_82_SUMB_22__26_,
         u5_mult_82_SUMB_22__27_, u5_mult_82_SUMB_22__28_,
         u5_mult_82_SUMB_22__29_, u5_mult_82_SUMB_22__30_,
         u5_mult_82_SUMB_22__31_, u5_mult_82_SUMB_22__32_,
         u5_mult_82_SUMB_22__33_, u5_mult_82_SUMB_22__34_,
         u5_mult_82_SUMB_22__35_, u5_mult_82_SUMB_22__36_,
         u5_mult_82_SUMB_22__37_, u5_mult_82_SUMB_22__38_,
         u5_mult_82_SUMB_22__39_, u5_mult_82_SUMB_22__40_,
         u5_mult_82_SUMB_22__41_, u5_mult_82_SUMB_22__42_,
         u5_mult_82_SUMB_22__43_, u5_mult_82_SUMB_22__44_,
         u5_mult_82_SUMB_22__45_, u5_mult_82_SUMB_22__46_,
         u5_mult_82_SUMB_22__47_, u5_mult_82_SUMB_22__48_,
         u5_mult_82_SUMB_22__49_, u5_mult_82_SUMB_22__50_,
         u5_mult_82_SUMB_22__51_, u5_mult_82_SUMB_23__1_,
         u5_mult_82_SUMB_23__2_, u5_mult_82_SUMB_23__3_,
         u5_mult_82_SUMB_23__4_, u5_mult_82_SUMB_23__5_,
         u5_mult_82_SUMB_23__6_, u5_mult_82_SUMB_23__7_,
         u5_mult_82_SUMB_23__8_, u5_mult_82_SUMB_23__9_,
         u5_mult_82_SUMB_23__10_, u5_mult_82_SUMB_23__11_,
         u5_mult_82_SUMB_23__12_, u5_mult_82_SUMB_23__13_,
         u5_mult_82_SUMB_23__14_, u5_mult_82_SUMB_23__15_,
         u5_mult_82_SUMB_23__16_, u5_mult_82_SUMB_23__17_,
         u5_mult_82_SUMB_23__18_, u5_mult_82_SUMB_23__19_,
         u5_mult_82_SUMB_23__20_, u5_mult_82_SUMB_23__21_,
         u5_mult_82_SUMB_23__22_, u5_mult_82_SUMB_23__24_,
         u5_mult_82_SUMB_23__25_, u5_mult_82_SUMB_23__26_,
         u5_mult_82_SUMB_23__27_, u5_mult_82_SUMB_23__28_,
         u5_mult_82_SUMB_23__29_, u5_mult_82_SUMB_23__30_,
         u5_mult_82_SUMB_23__31_, u5_mult_82_SUMB_23__32_,
         u5_mult_82_SUMB_23__33_, u5_mult_82_SUMB_23__34_,
         u5_mult_82_SUMB_23__35_, u5_mult_82_SUMB_23__36_,
         u5_mult_82_SUMB_23__37_, u5_mult_82_SUMB_23__38_,
         u5_mult_82_SUMB_23__39_, u5_mult_82_SUMB_23__40_,
         u5_mult_82_SUMB_23__41_, u5_mult_82_SUMB_23__42_,
         u5_mult_82_SUMB_23__43_, u5_mult_82_SUMB_23__44_,
         u5_mult_82_SUMB_23__45_, u5_mult_82_SUMB_23__46_,
         u5_mult_82_SUMB_23__47_, u5_mult_82_SUMB_23__48_,
         u5_mult_82_SUMB_23__49_, u5_mult_82_SUMB_23__50_,
         u5_mult_82_SUMB_23__51_, u5_mult_82_CARRYB_14__19_,
         u5_mult_82_CARRYB_14__20_, u5_mult_82_CARRYB_14__21_,
         u5_mult_82_CARRYB_14__22_, u5_mult_82_CARRYB_14__23_,
         u5_mult_82_CARRYB_14__24_, u5_mult_82_CARRYB_14__25_,
         u5_mult_82_CARRYB_14__26_, u5_mult_82_CARRYB_14__27_,
         u5_mult_82_CARRYB_14__29_, u5_mult_82_CARRYB_14__30_,
         u5_mult_82_CARRYB_14__31_, u5_mult_82_CARRYB_14__32_,
         u5_mult_82_CARRYB_14__33_, u5_mult_82_CARRYB_14__34_,
         u5_mult_82_CARRYB_14__35_, u5_mult_82_CARRYB_14__36_,
         u5_mult_82_CARRYB_14__37_, u5_mult_82_CARRYB_14__38_,
         u5_mult_82_CARRYB_14__39_, u5_mult_82_CARRYB_14__40_,
         u5_mult_82_CARRYB_14__41_, u5_mult_82_CARRYB_14__42_,
         u5_mult_82_CARRYB_14__43_, u5_mult_82_CARRYB_14__44_,
         u5_mult_82_CARRYB_14__45_, u5_mult_82_CARRYB_14__46_,
         u5_mult_82_CARRYB_14__47_, u5_mult_82_CARRYB_14__48_,
         u5_mult_82_CARRYB_14__49_, u5_mult_82_CARRYB_14__50_,
         u5_mult_82_CARRYB_14__51_, u5_mult_82_CARRYB_15__0_,
         u5_mult_82_CARRYB_15__1_, u5_mult_82_CARRYB_15__2_,
         u5_mult_82_CARRYB_15__3_, u5_mult_82_CARRYB_15__4_,
         u5_mult_82_CARRYB_15__5_, u5_mult_82_CARRYB_15__6_,
         u5_mult_82_CARRYB_15__7_, u5_mult_82_CARRYB_15__8_,
         u5_mult_82_CARRYB_15__9_, u5_mult_82_CARRYB_15__10_,
         u5_mult_82_CARRYB_15__11_, u5_mult_82_CARRYB_15__12_,
         u5_mult_82_CARRYB_15__13_, u5_mult_82_CARRYB_15__14_,
         u5_mult_82_CARRYB_15__15_, u5_mult_82_CARRYB_15__16_,
         u5_mult_82_CARRYB_15__17_, u5_mult_82_CARRYB_15__18_,
         u5_mult_82_CARRYB_15__19_, u5_mult_82_CARRYB_15__20_,
         u5_mult_82_CARRYB_15__21_, u5_mult_82_CARRYB_15__22_,
         u5_mult_82_CARRYB_15__23_, u5_mult_82_CARRYB_15__24_,
         u5_mult_82_CARRYB_15__25_, u5_mult_82_CARRYB_15__26_,
         u5_mult_82_CARRYB_15__28_, u5_mult_82_CARRYB_15__29_,
         u5_mult_82_CARRYB_15__30_, u5_mult_82_CARRYB_15__31_,
         u5_mult_82_CARRYB_15__32_, u5_mult_82_CARRYB_15__33_,
         u5_mult_82_CARRYB_15__34_, u5_mult_82_CARRYB_15__35_,
         u5_mult_82_CARRYB_15__36_, u5_mult_82_CARRYB_15__37_,
         u5_mult_82_CARRYB_15__38_, u5_mult_82_CARRYB_15__39_,
         u5_mult_82_CARRYB_15__40_, u5_mult_82_CARRYB_15__41_,
         u5_mult_82_CARRYB_15__42_, u5_mult_82_CARRYB_15__43_,
         u5_mult_82_CARRYB_15__44_, u5_mult_82_CARRYB_15__45_,
         u5_mult_82_CARRYB_15__46_, u5_mult_82_CARRYB_15__47_,
         u5_mult_82_CARRYB_15__48_, u5_mult_82_CARRYB_15__49_,
         u5_mult_82_CARRYB_15__50_, u5_mult_82_CARRYB_15__51_,
         u5_mult_82_CARRYB_16__0_, u5_mult_82_CARRYB_16__1_,
         u5_mult_82_CARRYB_16__2_, u5_mult_82_CARRYB_16__3_,
         u5_mult_82_CARRYB_16__4_, u5_mult_82_CARRYB_16__5_,
         u5_mult_82_CARRYB_16__6_, u5_mult_82_CARRYB_16__7_,
         u5_mult_82_CARRYB_16__8_, u5_mult_82_CARRYB_16__9_,
         u5_mult_82_CARRYB_16__10_, u5_mult_82_CARRYB_16__11_,
         u5_mult_82_CARRYB_16__12_, u5_mult_82_CARRYB_16__13_,
         u5_mult_82_CARRYB_16__14_, u5_mult_82_CARRYB_16__15_,
         u5_mult_82_CARRYB_16__16_, u5_mult_82_CARRYB_16__17_,
         u5_mult_82_CARRYB_16__18_, u5_mult_82_CARRYB_16__19_,
         u5_mult_82_CARRYB_16__20_, u5_mult_82_CARRYB_16__21_,
         u5_mult_82_CARRYB_16__22_, u5_mult_82_CARRYB_16__23_,
         u5_mult_82_CARRYB_16__24_, u5_mult_82_CARRYB_16__25_,
         u5_mult_82_CARRYB_16__26_, u5_mult_82_CARRYB_16__27_,
         u5_mult_82_CARRYB_16__29_, u5_mult_82_CARRYB_16__30_,
         u5_mult_82_CARRYB_16__31_, u5_mult_82_CARRYB_16__32_,
         u5_mult_82_CARRYB_16__33_, u5_mult_82_CARRYB_16__34_,
         u5_mult_82_CARRYB_16__35_, u5_mult_82_CARRYB_16__36_,
         u5_mult_82_CARRYB_16__37_, u5_mult_82_CARRYB_16__38_,
         u5_mult_82_CARRYB_16__39_, u5_mult_82_CARRYB_16__40_,
         u5_mult_82_CARRYB_16__41_, u5_mult_82_CARRYB_16__42_,
         u5_mult_82_CARRYB_16__43_, u5_mult_82_CARRYB_16__44_,
         u5_mult_82_CARRYB_16__45_, u5_mult_82_CARRYB_16__46_,
         u5_mult_82_CARRYB_16__47_, u5_mult_82_CARRYB_16__48_,
         u5_mult_82_CARRYB_16__49_, u5_mult_82_CARRYB_16__50_,
         u5_mult_82_CARRYB_16__51_, u5_mult_82_CARRYB_17__0_,
         u5_mult_82_CARRYB_17__1_, u5_mult_82_CARRYB_17__2_,
         u5_mult_82_CARRYB_17__3_, u5_mult_82_CARRYB_17__4_,
         u5_mult_82_CARRYB_17__5_, u5_mult_82_CARRYB_17__6_,
         u5_mult_82_CARRYB_17__7_, u5_mult_82_CARRYB_17__8_,
         u5_mult_82_CARRYB_17__9_, u5_mult_82_CARRYB_17__10_,
         u5_mult_82_CARRYB_17__11_, u5_mult_82_CARRYB_17__12_,
         u5_mult_82_CARRYB_17__13_, u5_mult_82_CARRYB_17__14_,
         u5_mult_82_CARRYB_17__15_, u5_mult_82_CARRYB_17__16_,
         u5_mult_82_CARRYB_17__17_, u5_mult_82_CARRYB_17__18_,
         u5_mult_82_CARRYB_17__19_, u5_mult_82_CARRYB_17__20_,
         u5_mult_82_CARRYB_17__21_, u5_mult_82_CARRYB_17__22_,
         u5_mult_82_CARRYB_17__23_, u5_mult_82_CARRYB_17__24_,
         u5_mult_82_CARRYB_17__25_, u5_mult_82_CARRYB_17__26_,
         u5_mult_82_CARRYB_17__27_, u5_mult_82_CARRYB_17__28_,
         u5_mult_82_CARRYB_17__29_, u5_mult_82_CARRYB_17__30_,
         u5_mult_82_CARRYB_17__31_, u5_mult_82_CARRYB_17__32_,
         u5_mult_82_CARRYB_17__33_, u5_mult_82_CARRYB_17__34_,
         u5_mult_82_CARRYB_17__35_, u5_mult_82_CARRYB_17__36_,
         u5_mult_82_CARRYB_17__37_, u5_mult_82_CARRYB_17__38_,
         u5_mult_82_CARRYB_17__39_, u5_mult_82_CARRYB_17__40_,
         u5_mult_82_CARRYB_17__41_, u5_mult_82_CARRYB_17__42_,
         u5_mult_82_CARRYB_17__43_, u5_mult_82_CARRYB_17__44_,
         u5_mult_82_CARRYB_17__45_, u5_mult_82_CARRYB_17__46_,
         u5_mult_82_CARRYB_17__47_, u5_mult_82_CARRYB_17__48_,
         u5_mult_82_CARRYB_17__49_, u5_mult_82_CARRYB_17__50_,
         u5_mult_82_CARRYB_17__51_, u5_mult_82_CARRYB_18__0_,
         u5_mult_82_CARRYB_18__1_, u5_mult_82_CARRYB_18__2_,
         u5_mult_82_CARRYB_18__3_, u5_mult_82_CARRYB_18__4_,
         u5_mult_82_CARRYB_18__5_, u5_mult_82_CARRYB_18__6_,
         u5_mult_82_CARRYB_18__7_, u5_mult_82_CARRYB_18__8_,
         u5_mult_82_CARRYB_18__9_, u5_mult_82_CARRYB_18__10_,
         u5_mult_82_CARRYB_18__11_, u5_mult_82_CARRYB_18__12_,
         u5_mult_82_CARRYB_18__13_, u5_mult_82_CARRYB_18__14_,
         u5_mult_82_CARRYB_18__15_, u5_mult_82_CARRYB_18__16_,
         u5_mult_82_CARRYB_18__17_, u5_mult_82_CARRYB_18__18_,
         u5_mult_82_CARRYB_18__19_, u5_mult_82_CARRYB_18__20_,
         u5_mult_82_CARRYB_18__21_, u5_mult_82_CARRYB_18__22_,
         u5_mult_82_CARRYB_18__23_, u5_mult_82_CARRYB_18__24_,
         u5_mult_82_CARRYB_18__25_, u5_mult_82_CARRYB_18__27_,
         u5_mult_82_CARRYB_18__28_, u5_mult_82_CARRYB_18__29_,
         u5_mult_82_CARRYB_18__30_, u5_mult_82_CARRYB_18__31_,
         u5_mult_82_CARRYB_18__32_, u5_mult_82_CARRYB_18__33_,
         u5_mult_82_CARRYB_18__34_, u5_mult_82_CARRYB_18__35_,
         u5_mult_82_CARRYB_18__36_, u5_mult_82_CARRYB_18__37_,
         u5_mult_82_CARRYB_18__38_, u5_mult_82_CARRYB_18__39_,
         u5_mult_82_CARRYB_18__40_, u5_mult_82_CARRYB_18__41_,
         u5_mult_82_CARRYB_18__42_, u5_mult_82_CARRYB_18__43_,
         u5_mult_82_CARRYB_18__44_, u5_mult_82_CARRYB_18__45_,
         u5_mult_82_CARRYB_18__46_, u5_mult_82_CARRYB_18__47_,
         u5_mult_82_CARRYB_18__48_, u5_mult_82_CARRYB_18__49_,
         u5_mult_82_CARRYB_18__50_, u5_mult_82_CARRYB_18__51_,
         u5_mult_82_CARRYB_19__0_, u5_mult_82_CARRYB_19__1_,
         u5_mult_82_CARRYB_19__2_, u5_mult_82_CARRYB_19__3_,
         u5_mult_82_CARRYB_19__4_, u5_mult_82_CARRYB_19__5_,
         u5_mult_82_CARRYB_19__6_, u5_mult_82_CARRYB_19__7_,
         u5_mult_82_CARRYB_19__8_, u5_mult_82_CARRYB_19__9_,
         u5_mult_82_CARRYB_19__10_, u5_mult_82_CARRYB_19__11_,
         u5_mult_82_CARRYB_19__12_, u5_mult_82_CARRYB_19__13_,
         u5_mult_82_CARRYB_19__14_, u5_mult_82_CARRYB_19__15_,
         u5_mult_82_CARRYB_19__16_, u5_mult_82_CARRYB_19__17_,
         u5_mult_82_CARRYB_19__18_, u5_mult_82_CARRYB_19__19_,
         u5_mult_82_CARRYB_19__20_, u5_mult_82_CARRYB_19__21_,
         u5_mult_82_CARRYB_19__22_, u5_mult_82_CARRYB_19__23_,
         u5_mult_82_CARRYB_19__24_, u5_mult_82_CARRYB_19__25_,
         u5_mult_82_CARRYB_19__27_, u5_mult_82_CARRYB_19__28_,
         u5_mult_82_CARRYB_19__29_, u5_mult_82_CARRYB_19__30_,
         u5_mult_82_CARRYB_19__31_, u5_mult_82_CARRYB_19__32_,
         u5_mult_82_CARRYB_19__33_, u5_mult_82_CARRYB_19__34_,
         u5_mult_82_CARRYB_19__35_, u5_mult_82_CARRYB_19__36_,
         u5_mult_82_CARRYB_19__37_, u5_mult_82_CARRYB_19__38_,
         u5_mult_82_CARRYB_19__39_, u5_mult_82_CARRYB_19__40_,
         u5_mult_82_CARRYB_19__41_, u5_mult_82_CARRYB_19__42_,
         u5_mult_82_CARRYB_19__43_, u5_mult_82_CARRYB_19__44_,
         u5_mult_82_CARRYB_19__45_, u5_mult_82_CARRYB_19__46_,
         u5_mult_82_CARRYB_19__47_, u5_mult_82_CARRYB_19__48_,
         u5_mult_82_CARRYB_19__49_, u5_mult_82_CARRYB_19__50_,
         u5_mult_82_CARRYB_19__51_, u5_mult_82_CARRYB_20__0_,
         u5_mult_82_CARRYB_20__1_, u5_mult_82_CARRYB_20__2_,
         u5_mult_82_CARRYB_20__3_, u5_mult_82_CARRYB_20__4_,
         u5_mult_82_CARRYB_20__5_, u5_mult_82_CARRYB_20__6_,
         u5_mult_82_CARRYB_20__7_, u5_mult_82_CARRYB_20__8_,
         u5_mult_82_CARRYB_20__9_, u5_mult_82_CARRYB_20__10_,
         u5_mult_82_CARRYB_20__11_, u5_mult_82_CARRYB_20__12_,
         u5_mult_82_CARRYB_20__13_, u5_mult_82_CARRYB_20__14_,
         u5_mult_82_CARRYB_20__15_, u5_mult_82_CARRYB_20__16_,
         u5_mult_82_CARRYB_20__17_, u5_mult_82_CARRYB_20__18_,
         u5_mult_82_CARRYB_20__19_, u5_mult_82_CARRYB_20__20_,
         u5_mult_82_CARRYB_20__21_, u5_mult_82_CARRYB_20__22_,
         u5_mult_82_CARRYB_20__23_, u5_mult_82_CARRYB_20__24_,
         u5_mult_82_CARRYB_20__25_, u5_mult_82_CARRYB_20__26_,
         u5_mult_82_CARRYB_20__27_, u5_mult_82_CARRYB_20__28_,
         u5_mult_82_CARRYB_20__29_, u5_mult_82_CARRYB_20__30_,
         u5_mult_82_CARRYB_20__31_, u5_mult_82_CARRYB_20__32_,
         u5_mult_82_CARRYB_20__33_, u5_mult_82_CARRYB_20__34_,
         u5_mult_82_CARRYB_20__35_, u5_mult_82_CARRYB_20__36_,
         u5_mult_82_CARRYB_20__37_, u5_mult_82_CARRYB_20__38_,
         u5_mult_82_CARRYB_20__39_, u5_mult_82_CARRYB_20__40_,
         u5_mult_82_CARRYB_20__41_, u5_mult_82_CARRYB_20__42_,
         u5_mult_82_CARRYB_20__43_, u5_mult_82_CARRYB_20__44_,
         u5_mult_82_CARRYB_20__45_, u5_mult_82_CARRYB_20__46_,
         u5_mult_82_CARRYB_20__47_, u5_mult_82_CARRYB_20__48_,
         u5_mult_82_CARRYB_20__49_, u5_mult_82_CARRYB_20__50_,
         u5_mult_82_CARRYB_20__51_, u5_mult_82_CARRYB_21__0_,
         u5_mult_82_CARRYB_21__1_, u5_mult_82_CARRYB_21__2_,
         u5_mult_82_CARRYB_21__3_, u5_mult_82_CARRYB_21__4_,
         u5_mult_82_CARRYB_21__5_, u5_mult_82_CARRYB_21__6_,
         u5_mult_82_CARRYB_21__7_, u5_mult_82_CARRYB_21__8_,
         u5_mult_82_CARRYB_21__9_, u5_mult_82_CARRYB_21__10_,
         u5_mult_82_CARRYB_21__11_, u5_mult_82_CARRYB_21__12_,
         u5_mult_82_CARRYB_21__13_, u5_mult_82_CARRYB_21__14_,
         u5_mult_82_CARRYB_21__15_, u5_mult_82_CARRYB_21__16_,
         u5_mult_82_CARRYB_21__17_, u5_mult_82_CARRYB_21__18_,
         u5_mult_82_CARRYB_21__19_, u5_mult_82_CARRYB_21__20_,
         u5_mult_82_CARRYB_21__21_, u5_mult_82_CARRYB_21__22_,
         u5_mult_82_CARRYB_21__23_, u5_mult_82_CARRYB_21__24_,
         u5_mult_82_CARRYB_21__25_, u5_mult_82_CARRYB_21__26_,
         u5_mult_82_CARRYB_21__27_, u5_mult_82_CARRYB_21__28_,
         u5_mult_82_CARRYB_21__29_, u5_mult_82_CARRYB_21__30_,
         u5_mult_82_CARRYB_21__31_, u5_mult_82_CARRYB_21__32_,
         u5_mult_82_CARRYB_21__33_, u5_mult_82_CARRYB_21__34_,
         u5_mult_82_CARRYB_21__35_, u5_mult_82_CARRYB_21__36_,
         u5_mult_82_CARRYB_21__37_, u5_mult_82_CARRYB_21__38_,
         u5_mult_82_CARRYB_21__39_, u5_mult_82_CARRYB_21__40_,
         u5_mult_82_CARRYB_21__41_, u5_mult_82_CARRYB_21__42_,
         u5_mult_82_CARRYB_21__43_, u5_mult_82_CARRYB_21__44_,
         u5_mult_82_CARRYB_21__45_, u5_mult_82_CARRYB_21__46_,
         u5_mult_82_CARRYB_21__47_, u5_mult_82_CARRYB_21__48_,
         u5_mult_82_CARRYB_21__49_, u5_mult_82_CARRYB_21__50_,
         u5_mult_82_CARRYB_21__51_, u5_mult_82_CARRYB_22__0_,
         u5_mult_82_CARRYB_22__1_, u5_mult_82_CARRYB_22__2_,
         u5_mult_82_CARRYB_22__3_, u5_mult_82_CARRYB_22__4_,
         u5_mult_82_CARRYB_22__5_, u5_mult_82_CARRYB_22__6_,
         u5_mult_82_CARRYB_22__7_, u5_mult_82_CARRYB_22__8_,
         u5_mult_82_CARRYB_22__9_, u5_mult_82_CARRYB_22__10_,
         u5_mult_82_CARRYB_22__11_, u5_mult_82_CARRYB_22__12_,
         u5_mult_82_CARRYB_22__13_, u5_mult_82_CARRYB_22__14_,
         u5_mult_82_CARRYB_22__15_, u5_mult_82_CARRYB_22__16_,
         u5_mult_82_CARRYB_22__17_, u5_mult_82_CARRYB_22__18_,
         u5_mult_82_CARRYB_22__19_, u5_mult_82_CARRYB_22__20_,
         u5_mult_82_CARRYB_22__21_, u5_mult_82_CARRYB_22__22_,
         u5_mult_82_CARRYB_22__24_, u5_mult_82_CARRYB_22__25_,
         u5_mult_82_CARRYB_22__26_, u5_mult_82_CARRYB_22__27_,
         u5_mult_82_CARRYB_22__28_, u5_mult_82_CARRYB_22__29_,
         u5_mult_82_CARRYB_22__30_, u5_mult_82_CARRYB_22__31_,
         u5_mult_82_CARRYB_22__32_, u5_mult_82_CARRYB_22__33_,
         u5_mult_82_CARRYB_22__34_, u5_mult_82_CARRYB_22__35_,
         u5_mult_82_CARRYB_22__36_, u5_mult_82_CARRYB_22__37_,
         u5_mult_82_CARRYB_22__38_, u5_mult_82_CARRYB_22__39_,
         u5_mult_82_CARRYB_22__40_, u5_mult_82_CARRYB_22__41_,
         u5_mult_82_CARRYB_22__42_, u5_mult_82_CARRYB_22__43_,
         u5_mult_82_CARRYB_22__44_, u5_mult_82_CARRYB_22__45_,
         u5_mult_82_CARRYB_22__46_, u5_mult_82_CARRYB_22__47_,
         u5_mult_82_CARRYB_22__48_, u5_mult_82_CARRYB_22__49_,
         u5_mult_82_CARRYB_22__50_, u5_mult_82_CARRYB_22__51_,
         u5_mult_82_CARRYB_23__0_, u5_mult_82_CARRYB_23__1_,
         u5_mult_82_CARRYB_23__2_, u5_mult_82_CARRYB_23__3_,
         u5_mult_82_CARRYB_23__4_, u5_mult_82_CARRYB_23__5_,
         u5_mult_82_CARRYB_23__6_, u5_mult_82_CARRYB_23__7_,
         u5_mult_82_CARRYB_23__8_, u5_mult_82_CARRYB_23__9_,
         u5_mult_82_CARRYB_23__10_, u5_mult_82_CARRYB_23__11_,
         u5_mult_82_CARRYB_23__12_, u5_mult_82_CARRYB_23__13_,
         u5_mult_82_CARRYB_23__14_, u5_mult_82_CARRYB_23__15_,
         u5_mult_82_CARRYB_23__16_, u5_mult_82_CARRYB_23__17_,
         u5_mult_82_CARRYB_23__18_, u5_mult_82_CARRYB_23__19_,
         u5_mult_82_CARRYB_23__20_, u5_mult_82_CARRYB_23__21_,
         u5_mult_82_CARRYB_23__22_, u5_mult_82_CARRYB_23__24_,
         u5_mult_82_CARRYB_23__25_, u5_mult_82_CARRYB_23__26_,
         u5_mult_82_CARRYB_23__27_, u5_mult_82_CARRYB_23__28_,
         u5_mult_82_CARRYB_23__29_, u5_mult_82_CARRYB_23__30_,
         u5_mult_82_CARRYB_23__31_, u5_mult_82_CARRYB_23__32_,
         u5_mult_82_CARRYB_23__33_, u5_mult_82_CARRYB_23__34_,
         u5_mult_82_CARRYB_23__35_, u5_mult_82_CARRYB_23__36_,
         u5_mult_82_CARRYB_23__37_, u5_mult_82_CARRYB_23__38_,
         u5_mult_82_CARRYB_23__39_, u5_mult_82_CARRYB_23__40_,
         u5_mult_82_CARRYB_23__41_, u5_mult_82_CARRYB_23__42_,
         u5_mult_82_CARRYB_23__43_, u5_mult_82_CARRYB_23__44_,
         u5_mult_82_CARRYB_23__45_, u5_mult_82_CARRYB_23__46_,
         u5_mult_82_CARRYB_23__47_, u5_mult_82_CARRYB_23__48_,
         u5_mult_82_CARRYB_23__49_, u5_mult_82_CARRYB_23__50_,
         u5_mult_82_CARRYB_23__51_, u5_mult_82_CARRYB_24__0_,
         u5_mult_82_SUMB_4__37_, u5_mult_82_SUMB_4__38_,
         u5_mult_82_SUMB_4__39_, u5_mult_82_SUMB_4__40_,
         u5_mult_82_SUMB_4__41_, u5_mult_82_SUMB_4__42_,
         u5_mult_82_SUMB_4__43_, u5_mult_82_SUMB_4__44_,
         u5_mult_82_SUMB_4__45_, u5_mult_82_SUMB_4__46_,
         u5_mult_82_SUMB_4__47_, u5_mult_82_SUMB_4__48_,
         u5_mult_82_SUMB_4__49_, u5_mult_82_SUMB_4__50_,
         u5_mult_82_SUMB_4__51_, u5_mult_82_SUMB_5__1_, u5_mult_82_SUMB_5__2_,
         u5_mult_82_SUMB_5__3_, u5_mult_82_SUMB_5__4_, u5_mult_82_SUMB_5__5_,
         u5_mult_82_SUMB_5__6_, u5_mult_82_SUMB_5__7_, u5_mult_82_SUMB_5__8_,
         u5_mult_82_SUMB_5__9_, u5_mult_82_SUMB_5__10_, u5_mult_82_SUMB_5__11_,
         u5_mult_82_SUMB_5__12_, u5_mult_82_SUMB_5__13_,
         u5_mult_82_SUMB_5__14_, u5_mult_82_SUMB_5__15_,
         u5_mult_82_SUMB_5__16_, u5_mult_82_SUMB_5__17_,
         u5_mult_82_SUMB_5__18_, u5_mult_82_SUMB_5__19_,
         u5_mult_82_SUMB_5__20_, u5_mult_82_SUMB_5__21_,
         u5_mult_82_SUMB_5__22_, u5_mult_82_SUMB_5__23_,
         u5_mult_82_SUMB_5__24_, u5_mult_82_SUMB_5__25_,
         u5_mult_82_SUMB_5__26_, u5_mult_82_SUMB_5__27_,
         u5_mult_82_SUMB_5__28_, u5_mult_82_SUMB_5__29_,
         u5_mult_82_SUMB_5__30_, u5_mult_82_SUMB_5__31_,
         u5_mult_82_SUMB_5__32_, u5_mult_82_SUMB_5__33_,
         u5_mult_82_SUMB_5__37_, u5_mult_82_SUMB_5__38_,
         u5_mult_82_SUMB_5__39_, u5_mult_82_SUMB_5__40_,
         u5_mult_82_SUMB_5__41_, u5_mult_82_SUMB_5__42_,
         u5_mult_82_SUMB_5__43_, u5_mult_82_SUMB_5__44_,
         u5_mult_82_SUMB_5__45_, u5_mult_82_SUMB_5__46_,
         u5_mult_82_SUMB_5__47_, u5_mult_82_SUMB_5__48_,
         u5_mult_82_SUMB_5__49_, u5_mult_82_SUMB_5__50_,
         u5_mult_82_SUMB_5__51_, u5_mult_82_SUMB_6__1_, u5_mult_82_SUMB_6__2_,
         u5_mult_82_SUMB_6__3_, u5_mult_82_SUMB_6__4_, u5_mult_82_SUMB_6__5_,
         u5_mult_82_SUMB_6__6_, u5_mult_82_SUMB_6__7_, u5_mult_82_SUMB_6__8_,
         u5_mult_82_SUMB_6__9_, u5_mult_82_SUMB_6__10_, u5_mult_82_SUMB_6__11_,
         u5_mult_82_SUMB_6__12_, u5_mult_82_SUMB_6__13_,
         u5_mult_82_SUMB_6__14_, u5_mult_82_SUMB_6__15_,
         u5_mult_82_SUMB_6__16_, u5_mult_82_SUMB_6__17_,
         u5_mult_82_SUMB_6__18_, u5_mult_82_SUMB_6__19_,
         u5_mult_82_SUMB_6__20_, u5_mult_82_SUMB_6__21_,
         u5_mult_82_SUMB_6__22_, u5_mult_82_SUMB_6__23_,
         u5_mult_82_SUMB_6__24_, u5_mult_82_SUMB_6__25_,
         u5_mult_82_SUMB_6__26_, u5_mult_82_SUMB_6__27_,
         u5_mult_82_SUMB_6__28_, u5_mult_82_SUMB_6__29_,
         u5_mult_82_SUMB_6__30_, u5_mult_82_SUMB_6__31_,
         u5_mult_82_SUMB_6__32_, u5_mult_82_SUMB_6__33_,
         u5_mult_82_SUMB_6__36_, u5_mult_82_SUMB_6__37_,
         u5_mult_82_SUMB_6__38_, u5_mult_82_SUMB_6__39_,
         u5_mult_82_SUMB_6__40_, u5_mult_82_SUMB_6__41_,
         u5_mult_82_SUMB_6__42_, u5_mult_82_SUMB_6__43_,
         u5_mult_82_SUMB_6__44_, u5_mult_82_SUMB_6__45_,
         u5_mult_82_SUMB_6__46_, u5_mult_82_SUMB_6__47_,
         u5_mult_82_SUMB_6__48_, u5_mult_82_SUMB_6__49_,
         u5_mult_82_SUMB_6__50_, u5_mult_82_SUMB_6__51_, u5_mult_82_SUMB_7__1_,
         u5_mult_82_SUMB_7__2_, u5_mult_82_SUMB_7__3_, u5_mult_82_SUMB_7__4_,
         u5_mult_82_SUMB_7__5_, u5_mult_82_SUMB_7__6_, u5_mult_82_SUMB_7__7_,
         u5_mult_82_SUMB_7__8_, u5_mult_82_SUMB_7__9_, u5_mult_82_SUMB_7__10_,
         u5_mult_82_SUMB_7__11_, u5_mult_82_SUMB_7__12_,
         u5_mult_82_SUMB_7__13_, u5_mult_82_SUMB_7__14_,
         u5_mult_82_SUMB_7__15_, u5_mult_82_SUMB_7__16_,
         u5_mult_82_SUMB_7__17_, u5_mult_82_SUMB_7__18_,
         u5_mult_82_SUMB_7__19_, u5_mult_82_SUMB_7__20_,
         u5_mult_82_SUMB_7__21_, u5_mult_82_SUMB_7__22_,
         u5_mult_82_SUMB_7__23_, u5_mult_82_SUMB_7__24_,
         u5_mult_82_SUMB_7__25_, u5_mult_82_SUMB_7__26_,
         u5_mult_82_SUMB_7__27_, u5_mult_82_SUMB_7__28_,
         u5_mult_82_SUMB_7__29_, u5_mult_82_SUMB_7__30_,
         u5_mult_82_SUMB_7__31_, u5_mult_82_SUMB_7__32_,
         u5_mult_82_SUMB_7__33_, u5_mult_82_SUMB_7__35_,
         u5_mult_82_SUMB_7__36_, u5_mult_82_SUMB_7__37_,
         u5_mult_82_SUMB_7__38_, u5_mult_82_SUMB_7__39_,
         u5_mult_82_SUMB_7__40_, u5_mult_82_SUMB_7__41_,
         u5_mult_82_SUMB_7__42_, u5_mult_82_SUMB_7__43_,
         u5_mult_82_SUMB_7__44_, u5_mult_82_SUMB_7__45_,
         u5_mult_82_SUMB_7__46_, u5_mult_82_SUMB_7__47_,
         u5_mult_82_SUMB_7__48_, u5_mult_82_SUMB_7__49_,
         u5_mult_82_SUMB_7__50_, u5_mult_82_SUMB_7__51_, u5_mult_82_SUMB_8__1_,
         u5_mult_82_SUMB_8__2_, u5_mult_82_SUMB_8__3_, u5_mult_82_SUMB_8__4_,
         u5_mult_82_SUMB_8__5_, u5_mult_82_SUMB_8__6_, u5_mult_82_SUMB_8__7_,
         u5_mult_82_SUMB_8__8_, u5_mult_82_SUMB_8__9_, u5_mult_82_SUMB_8__10_,
         u5_mult_82_SUMB_8__11_, u5_mult_82_SUMB_8__12_,
         u5_mult_82_SUMB_8__13_, u5_mult_82_SUMB_8__14_,
         u5_mult_82_SUMB_8__15_, u5_mult_82_SUMB_8__16_,
         u5_mult_82_SUMB_8__17_, u5_mult_82_SUMB_8__18_,
         u5_mult_82_SUMB_8__19_, u5_mult_82_SUMB_8__20_,
         u5_mult_82_SUMB_8__21_, u5_mult_82_SUMB_8__22_,
         u5_mult_82_SUMB_8__23_, u5_mult_82_SUMB_8__24_,
         u5_mult_82_SUMB_8__25_, u5_mult_82_SUMB_8__26_,
         u5_mult_82_SUMB_8__27_, u5_mult_82_SUMB_8__28_,
         u5_mult_82_SUMB_8__29_, u5_mult_82_SUMB_8__30_,
         u5_mult_82_SUMB_8__31_, u5_mult_82_SUMB_8__32_,
         u5_mult_82_SUMB_8__35_, u5_mult_82_SUMB_8__36_,
         u5_mult_82_SUMB_8__37_, u5_mult_82_SUMB_8__38_,
         u5_mult_82_SUMB_8__39_, u5_mult_82_SUMB_8__40_,
         u5_mult_82_SUMB_8__41_, u5_mult_82_SUMB_8__42_,
         u5_mult_82_SUMB_8__43_, u5_mult_82_SUMB_8__44_,
         u5_mult_82_SUMB_8__45_, u5_mult_82_SUMB_8__46_,
         u5_mult_82_SUMB_8__47_, u5_mult_82_SUMB_8__48_,
         u5_mult_82_SUMB_8__49_, u5_mult_82_SUMB_8__50_,
         u5_mult_82_SUMB_8__51_, u5_mult_82_SUMB_9__1_, u5_mult_82_SUMB_9__2_,
         u5_mult_82_SUMB_9__3_, u5_mult_82_SUMB_9__4_, u5_mult_82_SUMB_9__5_,
         u5_mult_82_SUMB_9__6_, u5_mult_82_SUMB_9__7_, u5_mult_82_SUMB_9__8_,
         u5_mult_82_SUMB_9__9_, u5_mult_82_SUMB_9__10_, u5_mult_82_SUMB_9__11_,
         u5_mult_82_SUMB_9__12_, u5_mult_82_SUMB_9__13_,
         u5_mult_82_SUMB_9__14_, u5_mult_82_SUMB_9__15_,
         u5_mult_82_SUMB_9__16_, u5_mult_82_SUMB_9__17_,
         u5_mult_82_SUMB_9__18_, u5_mult_82_SUMB_9__19_,
         u5_mult_82_SUMB_9__20_, u5_mult_82_SUMB_9__21_,
         u5_mult_82_SUMB_9__22_, u5_mult_82_SUMB_9__23_,
         u5_mult_82_SUMB_9__24_, u5_mult_82_SUMB_9__25_,
         u5_mult_82_SUMB_9__26_, u5_mult_82_SUMB_9__27_,
         u5_mult_82_SUMB_9__28_, u5_mult_82_SUMB_9__29_,
         u5_mult_82_SUMB_9__30_, u5_mult_82_SUMB_9__31_,
         u5_mult_82_SUMB_9__32_, u5_mult_82_SUMB_9__34_,
         u5_mult_82_SUMB_9__35_, u5_mult_82_SUMB_9__36_,
         u5_mult_82_SUMB_9__37_, u5_mult_82_SUMB_9__38_,
         u5_mult_82_SUMB_9__39_, u5_mult_82_SUMB_9__40_,
         u5_mult_82_SUMB_9__41_, u5_mult_82_SUMB_9__42_,
         u5_mult_82_SUMB_9__43_, u5_mult_82_SUMB_9__44_,
         u5_mult_82_SUMB_9__45_, u5_mult_82_SUMB_9__46_,
         u5_mult_82_SUMB_9__47_, u5_mult_82_SUMB_9__48_,
         u5_mult_82_SUMB_9__49_, u5_mult_82_SUMB_9__50_,
         u5_mult_82_SUMB_9__51_, u5_mult_82_SUMB_10__1_,
         u5_mult_82_SUMB_10__2_, u5_mult_82_SUMB_10__3_,
         u5_mult_82_SUMB_10__4_, u5_mult_82_SUMB_10__5_,
         u5_mult_82_SUMB_10__6_, u5_mult_82_SUMB_10__7_,
         u5_mult_82_SUMB_10__8_, u5_mult_82_SUMB_10__9_,
         u5_mult_82_SUMB_10__10_, u5_mult_82_SUMB_10__11_,
         u5_mult_82_SUMB_10__12_, u5_mult_82_SUMB_10__13_,
         u5_mult_82_SUMB_10__14_, u5_mult_82_SUMB_10__15_,
         u5_mult_82_SUMB_10__16_, u5_mult_82_SUMB_10__17_,
         u5_mult_82_SUMB_10__18_, u5_mult_82_SUMB_10__19_,
         u5_mult_82_SUMB_10__20_, u5_mult_82_SUMB_10__21_,
         u5_mult_82_SUMB_10__22_, u5_mult_82_SUMB_10__23_,
         u5_mult_82_SUMB_10__24_, u5_mult_82_SUMB_10__25_,
         u5_mult_82_SUMB_10__26_, u5_mult_82_SUMB_10__27_,
         u5_mult_82_SUMB_10__28_, u5_mult_82_SUMB_10__29_,
         u5_mult_82_SUMB_10__30_, u5_mult_82_SUMB_10__31_,
         u5_mult_82_SUMB_10__34_, u5_mult_82_SUMB_10__35_,
         u5_mult_82_SUMB_10__36_, u5_mult_82_SUMB_10__37_,
         u5_mult_82_SUMB_10__38_, u5_mult_82_SUMB_10__39_,
         u5_mult_82_SUMB_10__40_, u5_mult_82_SUMB_10__41_,
         u5_mult_82_SUMB_10__42_, u5_mult_82_SUMB_10__43_,
         u5_mult_82_SUMB_10__44_, u5_mult_82_SUMB_10__45_,
         u5_mult_82_SUMB_10__46_, u5_mult_82_SUMB_10__47_,
         u5_mult_82_SUMB_10__48_, u5_mult_82_SUMB_10__49_,
         u5_mult_82_SUMB_10__50_, u5_mult_82_SUMB_10__51_,
         u5_mult_82_SUMB_11__1_, u5_mult_82_SUMB_11__2_,
         u5_mult_82_SUMB_11__3_, u5_mult_82_SUMB_11__4_,
         u5_mult_82_SUMB_11__5_, u5_mult_82_SUMB_11__6_,
         u5_mult_82_SUMB_11__7_, u5_mult_82_SUMB_11__8_,
         u5_mult_82_SUMB_11__9_, u5_mult_82_SUMB_11__10_,
         u5_mult_82_SUMB_11__11_, u5_mult_82_SUMB_11__12_,
         u5_mult_82_SUMB_11__13_, u5_mult_82_SUMB_11__14_,
         u5_mult_82_SUMB_11__15_, u5_mult_82_SUMB_11__16_,
         u5_mult_82_SUMB_11__17_, u5_mult_82_SUMB_11__18_,
         u5_mult_82_SUMB_11__19_, u5_mult_82_SUMB_11__20_,
         u5_mult_82_SUMB_11__21_, u5_mult_82_SUMB_11__22_,
         u5_mult_82_SUMB_11__23_, u5_mult_82_SUMB_11__24_,
         u5_mult_82_SUMB_11__25_, u5_mult_82_SUMB_11__26_,
         u5_mult_82_SUMB_11__27_, u5_mult_82_SUMB_11__28_,
         u5_mult_82_SUMB_11__29_, u5_mult_82_SUMB_11__30_,
         u5_mult_82_SUMB_11__33_, u5_mult_82_SUMB_11__34_,
         u5_mult_82_SUMB_11__35_, u5_mult_82_SUMB_11__36_,
         u5_mult_82_SUMB_11__37_, u5_mult_82_SUMB_11__38_,
         u5_mult_82_SUMB_11__39_, u5_mult_82_SUMB_11__40_,
         u5_mult_82_SUMB_11__41_, u5_mult_82_SUMB_11__42_,
         u5_mult_82_SUMB_11__44_, u5_mult_82_SUMB_11__45_,
         u5_mult_82_SUMB_11__46_, u5_mult_82_SUMB_11__47_,
         u5_mult_82_SUMB_11__48_, u5_mult_82_SUMB_11__49_,
         u5_mult_82_SUMB_11__50_, u5_mult_82_SUMB_11__51_,
         u5_mult_82_SUMB_12__1_, u5_mult_82_SUMB_12__2_,
         u5_mult_82_SUMB_12__3_, u5_mult_82_SUMB_12__4_,
         u5_mult_82_SUMB_12__5_, u5_mult_82_SUMB_12__6_,
         u5_mult_82_SUMB_12__7_, u5_mult_82_SUMB_12__8_,
         u5_mult_82_SUMB_12__9_, u5_mult_82_SUMB_12__10_,
         u5_mult_82_SUMB_12__11_, u5_mult_82_SUMB_12__12_,
         u5_mult_82_SUMB_12__13_, u5_mult_82_SUMB_12__14_,
         u5_mult_82_SUMB_12__15_, u5_mult_82_SUMB_12__16_,
         u5_mult_82_SUMB_12__17_, u5_mult_82_SUMB_12__18_,
         u5_mult_82_SUMB_12__19_, u5_mult_82_SUMB_12__20_,
         u5_mult_82_SUMB_12__21_, u5_mult_82_SUMB_12__22_,
         u5_mult_82_SUMB_12__23_, u5_mult_82_SUMB_12__24_,
         u5_mult_82_SUMB_12__25_, u5_mult_82_SUMB_12__26_,
         u5_mult_82_SUMB_12__27_, u5_mult_82_SUMB_12__28_,
         u5_mult_82_SUMB_12__29_, u5_mult_82_SUMB_12__32_,
         u5_mult_82_SUMB_12__33_, u5_mult_82_SUMB_12__34_,
         u5_mult_82_SUMB_12__35_, u5_mult_82_SUMB_12__36_,
         u5_mult_82_SUMB_12__37_, u5_mult_82_SUMB_12__38_,
         u5_mult_82_SUMB_12__39_, u5_mult_82_SUMB_12__40_,
         u5_mult_82_SUMB_12__41_, u5_mult_82_SUMB_12__42_,
         u5_mult_82_SUMB_12__43_, u5_mult_82_SUMB_12__44_,
         u5_mult_82_SUMB_12__45_, u5_mult_82_SUMB_12__46_,
         u5_mult_82_SUMB_12__47_, u5_mult_82_SUMB_12__48_,
         u5_mult_82_SUMB_12__49_, u5_mult_82_SUMB_12__50_,
         u5_mult_82_SUMB_12__51_, u5_mult_82_SUMB_13__1_,
         u5_mult_82_SUMB_13__2_, u5_mult_82_SUMB_13__3_,
         u5_mult_82_SUMB_13__4_, u5_mult_82_SUMB_13__5_,
         u5_mult_82_SUMB_13__6_, u5_mult_82_SUMB_13__7_,
         u5_mult_82_SUMB_13__8_, u5_mult_82_SUMB_13__9_,
         u5_mult_82_SUMB_13__10_, u5_mult_82_SUMB_13__11_,
         u5_mult_82_SUMB_13__12_, u5_mult_82_SUMB_13__13_,
         u5_mult_82_SUMB_13__14_, u5_mult_82_SUMB_13__15_,
         u5_mult_82_SUMB_13__16_, u5_mult_82_SUMB_13__17_,
         u5_mult_82_SUMB_13__18_, u5_mult_82_SUMB_13__19_,
         u5_mult_82_SUMB_13__20_, u5_mult_82_SUMB_13__21_,
         u5_mult_82_SUMB_13__22_, u5_mult_82_SUMB_13__23_,
         u5_mult_82_SUMB_13__24_, u5_mult_82_SUMB_13__25_,
         u5_mult_82_SUMB_13__26_, u5_mult_82_SUMB_13__27_,
         u5_mult_82_SUMB_13__28_, u5_mult_82_SUMB_13__30_,
         u5_mult_82_SUMB_13__31_, u5_mult_82_SUMB_13__32_,
         u5_mult_82_SUMB_13__33_, u5_mult_82_SUMB_13__34_,
         u5_mult_82_SUMB_13__35_, u5_mult_82_SUMB_13__36_,
         u5_mult_82_SUMB_13__37_, u5_mult_82_SUMB_13__38_,
         u5_mult_82_SUMB_13__39_, u5_mult_82_SUMB_13__40_,
         u5_mult_82_SUMB_13__41_, u5_mult_82_SUMB_13__42_,
         u5_mult_82_SUMB_13__43_, u5_mult_82_SUMB_13__44_,
         u5_mult_82_SUMB_13__45_, u5_mult_82_SUMB_13__46_,
         u5_mult_82_SUMB_13__47_, u5_mult_82_SUMB_13__48_,
         u5_mult_82_SUMB_13__49_, u5_mult_82_SUMB_13__50_,
         u5_mult_82_SUMB_13__51_, u5_mult_82_SUMB_14__1_,
         u5_mult_82_SUMB_14__2_, u5_mult_82_SUMB_14__3_,
         u5_mult_82_SUMB_14__4_, u5_mult_82_SUMB_14__5_,
         u5_mult_82_SUMB_14__6_, u5_mult_82_SUMB_14__7_,
         u5_mult_82_SUMB_14__8_, u5_mult_82_SUMB_14__9_,
         u5_mult_82_SUMB_14__10_, u5_mult_82_SUMB_14__11_,
         u5_mult_82_SUMB_14__12_, u5_mult_82_SUMB_14__13_,
         u5_mult_82_SUMB_14__14_, u5_mult_82_SUMB_14__15_,
         u5_mult_82_SUMB_14__16_, u5_mult_82_SUMB_14__17_,
         u5_mult_82_SUMB_14__18_, u5_mult_82_CARRYB_4__37_,
         u5_mult_82_CARRYB_4__38_, u5_mult_82_CARRYB_4__39_,
         u5_mult_82_CARRYB_4__40_, u5_mult_82_CARRYB_4__41_,
         u5_mult_82_CARRYB_4__42_, u5_mult_82_CARRYB_4__43_,
         u5_mult_82_CARRYB_4__44_, u5_mult_82_CARRYB_4__45_,
         u5_mult_82_CARRYB_4__46_, u5_mult_82_CARRYB_4__47_,
         u5_mult_82_CARRYB_4__48_, u5_mult_82_CARRYB_4__49_,
         u5_mult_82_CARRYB_4__50_, u5_mult_82_CARRYB_4__51_,
         u5_mult_82_CARRYB_5__0_, u5_mult_82_CARRYB_5__1_,
         u5_mult_82_CARRYB_5__2_, u5_mult_82_CARRYB_5__3_,
         u5_mult_82_CARRYB_5__4_, u5_mult_82_CARRYB_5__5_,
         u5_mult_82_CARRYB_5__6_, u5_mult_82_CARRYB_5__7_,
         u5_mult_82_CARRYB_5__8_, u5_mult_82_CARRYB_5__9_,
         u5_mult_82_CARRYB_5__10_, u5_mult_82_CARRYB_5__11_,
         u5_mult_82_CARRYB_5__12_, u5_mult_82_CARRYB_5__13_,
         u5_mult_82_CARRYB_5__14_, u5_mult_82_CARRYB_5__15_,
         u5_mult_82_CARRYB_5__16_, u5_mult_82_CARRYB_5__17_,
         u5_mult_82_CARRYB_5__18_, u5_mult_82_CARRYB_5__19_,
         u5_mult_82_CARRYB_5__20_, u5_mult_82_CARRYB_5__21_,
         u5_mult_82_CARRYB_5__22_, u5_mult_82_CARRYB_5__23_,
         u5_mult_82_CARRYB_5__24_, u5_mult_82_CARRYB_5__25_,
         u5_mult_82_CARRYB_5__26_, u5_mult_82_CARRYB_5__27_,
         u5_mult_82_CARRYB_5__28_, u5_mult_82_CARRYB_5__29_,
         u5_mult_82_CARRYB_5__30_, u5_mult_82_CARRYB_5__31_,
         u5_mult_82_CARRYB_5__32_, u5_mult_82_CARRYB_5__33_,
         u5_mult_82_CARRYB_5__36_, u5_mult_82_CARRYB_5__37_,
         u5_mult_82_CARRYB_5__38_, u5_mult_82_CARRYB_5__39_,
         u5_mult_82_CARRYB_5__40_, u5_mult_82_CARRYB_5__41_,
         u5_mult_82_CARRYB_5__42_, u5_mult_82_CARRYB_5__43_,
         u5_mult_82_CARRYB_5__44_, u5_mult_82_CARRYB_5__45_,
         u5_mult_82_CARRYB_5__46_, u5_mult_82_CARRYB_5__47_,
         u5_mult_82_CARRYB_5__48_, u5_mult_82_CARRYB_5__49_,
         u5_mult_82_CARRYB_5__50_, u5_mult_82_CARRYB_5__51_,
         u5_mult_82_CARRYB_6__0_, u5_mult_82_CARRYB_6__1_,
         u5_mult_82_CARRYB_6__2_, u5_mult_82_CARRYB_6__3_,
         u5_mult_82_CARRYB_6__4_, u5_mult_82_CARRYB_6__5_,
         u5_mult_82_CARRYB_6__6_, u5_mult_82_CARRYB_6__7_,
         u5_mult_82_CARRYB_6__8_, u5_mult_82_CARRYB_6__9_,
         u5_mult_82_CARRYB_6__10_, u5_mult_82_CARRYB_6__11_,
         u5_mult_82_CARRYB_6__12_, u5_mult_82_CARRYB_6__13_,
         u5_mult_82_CARRYB_6__14_, u5_mult_82_CARRYB_6__15_,
         u5_mult_82_CARRYB_6__16_, u5_mult_82_CARRYB_6__17_,
         u5_mult_82_CARRYB_6__18_, u5_mult_82_CARRYB_6__19_,
         u5_mult_82_CARRYB_6__20_, u5_mult_82_CARRYB_6__21_,
         u5_mult_82_CARRYB_6__22_, u5_mult_82_CARRYB_6__23_,
         u5_mult_82_CARRYB_6__24_, u5_mult_82_CARRYB_6__25_,
         u5_mult_82_CARRYB_6__26_, u5_mult_82_CARRYB_6__27_,
         u5_mult_82_CARRYB_6__28_, u5_mult_82_CARRYB_6__29_,
         u5_mult_82_CARRYB_6__30_, u5_mult_82_CARRYB_6__31_,
         u5_mult_82_CARRYB_6__32_, u5_mult_82_CARRYB_6__33_,
         u5_mult_82_CARRYB_6__36_, u5_mult_82_CARRYB_6__37_,
         u5_mult_82_CARRYB_6__38_, u5_mult_82_CARRYB_6__39_,
         u5_mult_82_CARRYB_6__40_, u5_mult_82_CARRYB_6__41_,
         u5_mult_82_CARRYB_6__42_, u5_mult_82_CARRYB_6__43_,
         u5_mult_82_CARRYB_6__44_, u5_mult_82_CARRYB_6__45_,
         u5_mult_82_CARRYB_6__46_, u5_mult_82_CARRYB_6__47_,
         u5_mult_82_CARRYB_6__48_, u5_mult_82_CARRYB_6__49_,
         u5_mult_82_CARRYB_6__50_, u5_mult_82_CARRYB_6__51_,
         u5_mult_82_CARRYB_7__0_, u5_mult_82_CARRYB_7__1_,
         u5_mult_82_CARRYB_7__2_, u5_mult_82_CARRYB_7__3_,
         u5_mult_82_CARRYB_7__4_, u5_mult_82_CARRYB_7__5_,
         u5_mult_82_CARRYB_7__6_, u5_mult_82_CARRYB_7__7_,
         u5_mult_82_CARRYB_7__8_, u5_mult_82_CARRYB_7__9_,
         u5_mult_82_CARRYB_7__10_, u5_mult_82_CARRYB_7__11_,
         u5_mult_82_CARRYB_7__12_, u5_mult_82_CARRYB_7__13_,
         u5_mult_82_CARRYB_7__14_, u5_mult_82_CARRYB_7__15_,
         u5_mult_82_CARRYB_7__16_, u5_mult_82_CARRYB_7__17_,
         u5_mult_82_CARRYB_7__18_, u5_mult_82_CARRYB_7__19_,
         u5_mult_82_CARRYB_7__20_, u5_mult_82_CARRYB_7__21_,
         u5_mult_82_CARRYB_7__22_, u5_mult_82_CARRYB_7__23_,
         u5_mult_82_CARRYB_7__24_, u5_mult_82_CARRYB_7__25_,
         u5_mult_82_CARRYB_7__26_, u5_mult_82_CARRYB_7__27_,
         u5_mult_82_CARRYB_7__28_, u5_mult_82_CARRYB_7__29_,
         u5_mult_82_CARRYB_7__30_, u5_mult_82_CARRYB_7__31_,
         u5_mult_82_CARRYB_7__32_, u5_mult_82_CARRYB_7__33_,
         u5_mult_82_CARRYB_7__35_, u5_mult_82_CARRYB_7__36_,
         u5_mult_82_CARRYB_7__37_, u5_mult_82_CARRYB_7__38_,
         u5_mult_82_CARRYB_7__39_, u5_mult_82_CARRYB_7__40_,
         u5_mult_82_CARRYB_7__41_, u5_mult_82_CARRYB_7__42_,
         u5_mult_82_CARRYB_7__43_, u5_mult_82_CARRYB_7__44_,
         u5_mult_82_CARRYB_7__45_, u5_mult_82_CARRYB_7__46_,
         u5_mult_82_CARRYB_7__47_, u5_mult_82_CARRYB_7__48_,
         u5_mult_82_CARRYB_7__49_, u5_mult_82_CARRYB_7__50_,
         u5_mult_82_CARRYB_7__51_, u5_mult_82_CARRYB_8__0_,
         u5_mult_82_CARRYB_8__1_, u5_mult_82_CARRYB_8__2_,
         u5_mult_82_CARRYB_8__3_, u5_mult_82_CARRYB_8__4_,
         u5_mult_82_CARRYB_8__5_, u5_mult_82_CARRYB_8__6_,
         u5_mult_82_CARRYB_8__7_, u5_mult_82_CARRYB_8__8_,
         u5_mult_82_CARRYB_8__9_, u5_mult_82_CARRYB_8__10_,
         u5_mult_82_CARRYB_8__11_, u5_mult_82_CARRYB_8__12_,
         u5_mult_82_CARRYB_8__13_, u5_mult_82_CARRYB_8__14_,
         u5_mult_82_CARRYB_8__15_, u5_mult_82_CARRYB_8__16_,
         u5_mult_82_CARRYB_8__17_, u5_mult_82_CARRYB_8__18_,
         u5_mult_82_CARRYB_8__19_, u5_mult_82_CARRYB_8__20_,
         u5_mult_82_CARRYB_8__21_, u5_mult_82_CARRYB_8__22_,
         u5_mult_82_CARRYB_8__23_, u5_mult_82_CARRYB_8__24_,
         u5_mult_82_CARRYB_8__25_, u5_mult_82_CARRYB_8__26_,
         u5_mult_82_CARRYB_8__27_, u5_mult_82_CARRYB_8__28_,
         u5_mult_82_CARRYB_8__29_, u5_mult_82_CARRYB_8__30_,
         u5_mult_82_CARRYB_8__31_, u5_mult_82_CARRYB_8__32_,
         u5_mult_82_CARRYB_8__34_, u5_mult_82_CARRYB_8__35_,
         u5_mult_82_CARRYB_8__36_, u5_mult_82_CARRYB_8__37_,
         u5_mult_82_CARRYB_8__38_, u5_mult_82_CARRYB_8__39_,
         u5_mult_82_CARRYB_8__40_, u5_mult_82_CARRYB_8__41_,
         u5_mult_82_CARRYB_8__42_, u5_mult_82_CARRYB_8__43_,
         u5_mult_82_CARRYB_8__44_, u5_mult_82_CARRYB_8__45_,
         u5_mult_82_CARRYB_8__46_, u5_mult_82_CARRYB_8__47_,
         u5_mult_82_CARRYB_8__48_, u5_mult_82_CARRYB_8__49_,
         u5_mult_82_CARRYB_8__50_, u5_mult_82_CARRYB_8__51_,
         u5_mult_82_CARRYB_9__0_, u5_mult_82_CARRYB_9__1_,
         u5_mult_82_CARRYB_9__2_, u5_mult_82_CARRYB_9__3_,
         u5_mult_82_CARRYB_9__4_, u5_mult_82_CARRYB_9__5_,
         u5_mult_82_CARRYB_9__6_, u5_mult_82_CARRYB_9__7_,
         u5_mult_82_CARRYB_9__8_, u5_mult_82_CARRYB_9__9_,
         u5_mult_82_CARRYB_9__10_, u5_mult_82_CARRYB_9__11_,
         u5_mult_82_CARRYB_9__12_, u5_mult_82_CARRYB_9__13_,
         u5_mult_82_CARRYB_9__14_, u5_mult_82_CARRYB_9__15_,
         u5_mult_82_CARRYB_9__16_, u5_mult_82_CARRYB_9__17_,
         u5_mult_82_CARRYB_9__18_, u5_mult_82_CARRYB_9__19_,
         u5_mult_82_CARRYB_9__20_, u5_mult_82_CARRYB_9__21_,
         u5_mult_82_CARRYB_9__22_, u5_mult_82_CARRYB_9__23_,
         u5_mult_82_CARRYB_9__24_, u5_mult_82_CARRYB_9__25_,
         u5_mult_82_CARRYB_9__26_, u5_mult_82_CARRYB_9__27_,
         u5_mult_82_CARRYB_9__28_, u5_mult_82_CARRYB_9__29_,
         u5_mult_82_CARRYB_9__30_, u5_mult_82_CARRYB_9__31_,
         u5_mult_82_CARRYB_9__34_, u5_mult_82_CARRYB_9__35_,
         u5_mult_82_CARRYB_9__36_, u5_mult_82_CARRYB_9__37_,
         u5_mult_82_CARRYB_9__38_, u5_mult_82_CARRYB_9__39_,
         u5_mult_82_CARRYB_9__40_, u5_mult_82_CARRYB_9__41_,
         u5_mult_82_CARRYB_9__42_, u5_mult_82_CARRYB_9__43_,
         u5_mult_82_CARRYB_9__44_, u5_mult_82_CARRYB_9__45_,
         u5_mult_82_CARRYB_9__46_, u5_mult_82_CARRYB_9__47_,
         u5_mult_82_CARRYB_9__48_, u5_mult_82_CARRYB_9__49_,
         u5_mult_82_CARRYB_9__50_, u5_mult_82_CARRYB_9__51_,
         u5_mult_82_CARRYB_10__0_, u5_mult_82_CARRYB_10__1_,
         u5_mult_82_CARRYB_10__2_, u5_mult_82_CARRYB_10__3_,
         u5_mult_82_CARRYB_10__4_, u5_mult_82_CARRYB_10__5_,
         u5_mult_82_CARRYB_10__6_, u5_mult_82_CARRYB_10__7_,
         u5_mult_82_CARRYB_10__8_, u5_mult_82_CARRYB_10__9_,
         u5_mult_82_CARRYB_10__10_, u5_mult_82_CARRYB_10__11_,
         u5_mult_82_CARRYB_10__12_, u5_mult_82_CARRYB_10__13_,
         u5_mult_82_CARRYB_10__14_, u5_mult_82_CARRYB_10__15_,
         u5_mult_82_CARRYB_10__16_, u5_mult_82_CARRYB_10__17_,
         u5_mult_82_CARRYB_10__18_, u5_mult_82_CARRYB_10__19_,
         u5_mult_82_CARRYB_10__20_, u5_mult_82_CARRYB_10__21_,
         u5_mult_82_CARRYB_10__22_, u5_mult_82_CARRYB_10__23_,
         u5_mult_82_CARRYB_10__24_, u5_mult_82_CARRYB_10__25_,
         u5_mult_82_CARRYB_10__26_, u5_mult_82_CARRYB_10__27_,
         u5_mult_82_CARRYB_10__28_, u5_mult_82_CARRYB_10__29_,
         u5_mult_82_CARRYB_10__30_, u5_mult_82_CARRYB_10__31_,
         u5_mult_82_CARRYB_10__33_, u5_mult_82_CARRYB_10__34_,
         u5_mult_82_CARRYB_10__35_, u5_mult_82_CARRYB_10__36_,
         u5_mult_82_CARRYB_10__37_, u5_mult_82_CARRYB_10__38_,
         u5_mult_82_CARRYB_10__39_, u5_mult_82_CARRYB_10__40_,
         u5_mult_82_CARRYB_10__41_, u5_mult_82_CARRYB_10__42_,
         u5_mult_82_CARRYB_10__43_, u5_mult_82_CARRYB_10__44_,
         u5_mult_82_CARRYB_10__45_, u5_mult_82_CARRYB_10__46_,
         u5_mult_82_CARRYB_10__47_, u5_mult_82_CARRYB_10__48_,
         u5_mult_82_CARRYB_10__49_, u5_mult_82_CARRYB_10__50_,
         u5_mult_82_CARRYB_10__51_, u5_mult_82_CARRYB_11__0_,
         u5_mult_82_CARRYB_11__1_, u5_mult_82_CARRYB_11__2_,
         u5_mult_82_CARRYB_11__3_, u5_mult_82_CARRYB_11__4_,
         u5_mult_82_CARRYB_11__5_, u5_mult_82_CARRYB_11__6_,
         u5_mult_82_CARRYB_11__7_, u5_mult_82_CARRYB_11__8_,
         u5_mult_82_CARRYB_11__9_, u5_mult_82_CARRYB_11__10_,
         u5_mult_82_CARRYB_11__11_, u5_mult_82_CARRYB_11__12_,
         u5_mult_82_CARRYB_11__13_, u5_mult_82_CARRYB_11__14_,
         u5_mult_82_CARRYB_11__15_, u5_mult_82_CARRYB_11__16_,
         u5_mult_82_CARRYB_11__17_, u5_mult_82_CARRYB_11__18_,
         u5_mult_82_CARRYB_11__19_, u5_mult_82_CARRYB_11__20_,
         u5_mult_82_CARRYB_11__21_, u5_mult_82_CARRYB_11__22_,
         u5_mult_82_CARRYB_11__23_, u5_mult_82_CARRYB_11__24_,
         u5_mult_82_CARRYB_11__25_, u5_mult_82_CARRYB_11__26_,
         u5_mult_82_CARRYB_11__27_, u5_mult_82_CARRYB_11__28_,
         u5_mult_82_CARRYB_11__29_, u5_mult_82_CARRYB_11__30_,
         u5_mult_82_CARRYB_11__32_, u5_mult_82_CARRYB_11__33_,
         u5_mult_82_CARRYB_11__34_, u5_mult_82_CARRYB_11__35_,
         u5_mult_82_CARRYB_11__36_, u5_mult_82_CARRYB_11__37_,
         u5_mult_82_CARRYB_11__38_, u5_mult_82_CARRYB_11__39_,
         u5_mult_82_CARRYB_11__40_, u5_mult_82_CARRYB_11__41_,
         u5_mult_82_CARRYB_11__42_, u5_mult_82_CARRYB_11__43_,
         u5_mult_82_CARRYB_11__44_, u5_mult_82_CARRYB_11__45_,
         u5_mult_82_CARRYB_11__46_, u5_mult_82_CARRYB_11__47_,
         u5_mult_82_CARRYB_11__48_, u5_mult_82_CARRYB_11__49_,
         u5_mult_82_CARRYB_11__50_, u5_mult_82_CARRYB_11__51_,
         u5_mult_82_CARRYB_12__0_, u5_mult_82_CARRYB_12__1_,
         u5_mult_82_CARRYB_12__2_, u5_mult_82_CARRYB_12__3_,
         u5_mult_82_CARRYB_12__4_, u5_mult_82_CARRYB_12__5_,
         u5_mult_82_CARRYB_12__6_, u5_mult_82_CARRYB_12__7_,
         u5_mult_82_CARRYB_12__8_, u5_mult_82_CARRYB_12__9_,
         u5_mult_82_CARRYB_12__10_, u5_mult_82_CARRYB_12__11_,
         u5_mult_82_CARRYB_12__12_, u5_mult_82_CARRYB_12__13_,
         u5_mult_82_CARRYB_12__14_, u5_mult_82_CARRYB_12__15_,
         u5_mult_82_CARRYB_12__16_, u5_mult_82_CARRYB_12__17_,
         u5_mult_82_CARRYB_12__18_, u5_mult_82_CARRYB_12__19_,
         u5_mult_82_CARRYB_12__20_, u5_mult_82_CARRYB_12__21_,
         u5_mult_82_CARRYB_12__22_, u5_mult_82_CARRYB_12__23_,
         u5_mult_82_CARRYB_12__24_, u5_mult_82_CARRYB_12__25_,
         u5_mult_82_CARRYB_12__26_, u5_mult_82_CARRYB_12__27_,
         u5_mult_82_CARRYB_12__28_, u5_mult_82_CARRYB_12__29_,
         u5_mult_82_CARRYB_12__31_, u5_mult_82_CARRYB_12__32_,
         u5_mult_82_CARRYB_12__33_, u5_mult_82_CARRYB_12__34_,
         u5_mult_82_CARRYB_12__35_, u5_mult_82_CARRYB_12__36_,
         u5_mult_82_CARRYB_12__37_, u5_mult_82_CARRYB_12__38_,
         u5_mult_82_CARRYB_12__39_, u5_mult_82_CARRYB_12__40_,
         u5_mult_82_CARRYB_12__41_, u5_mult_82_CARRYB_12__42_,
         u5_mult_82_CARRYB_12__43_, u5_mult_82_CARRYB_12__44_,
         u5_mult_82_CARRYB_12__45_, u5_mult_82_CARRYB_12__46_,
         u5_mult_82_CARRYB_12__47_, u5_mult_82_CARRYB_12__48_,
         u5_mult_82_CARRYB_12__49_, u5_mult_82_CARRYB_12__50_,
         u5_mult_82_CARRYB_12__51_, u5_mult_82_CARRYB_13__0_,
         u5_mult_82_CARRYB_13__1_, u5_mult_82_CARRYB_13__2_,
         u5_mult_82_CARRYB_13__3_, u5_mult_82_CARRYB_13__4_,
         u5_mult_82_CARRYB_13__5_, u5_mult_82_CARRYB_13__6_,
         u5_mult_82_CARRYB_13__7_, u5_mult_82_CARRYB_13__8_,
         u5_mult_82_CARRYB_13__9_, u5_mult_82_CARRYB_13__10_,
         u5_mult_82_CARRYB_13__11_, u5_mult_82_CARRYB_13__12_,
         u5_mult_82_CARRYB_13__13_, u5_mult_82_CARRYB_13__14_,
         u5_mult_82_CARRYB_13__15_, u5_mult_82_CARRYB_13__16_,
         u5_mult_82_CARRYB_13__17_, u5_mult_82_CARRYB_13__18_,
         u5_mult_82_CARRYB_13__19_, u5_mult_82_CARRYB_13__20_,
         u5_mult_82_CARRYB_13__21_, u5_mult_82_CARRYB_13__22_,
         u5_mult_82_CARRYB_13__23_, u5_mult_82_CARRYB_13__24_,
         u5_mult_82_CARRYB_13__25_, u5_mult_82_CARRYB_13__26_,
         u5_mult_82_CARRYB_13__27_, u5_mult_82_CARRYB_13__28_,
         u5_mult_82_CARRYB_13__30_, u5_mult_82_CARRYB_13__31_,
         u5_mult_82_CARRYB_13__32_, u5_mult_82_CARRYB_13__33_,
         u5_mult_82_CARRYB_13__34_, u5_mult_82_CARRYB_13__35_,
         u5_mult_82_CARRYB_13__36_, u5_mult_82_CARRYB_13__37_,
         u5_mult_82_CARRYB_13__38_, u5_mult_82_CARRYB_13__39_,
         u5_mult_82_CARRYB_13__40_, u5_mult_82_CARRYB_13__41_,
         u5_mult_82_CARRYB_13__42_, u5_mult_82_CARRYB_13__43_,
         u5_mult_82_CARRYB_13__44_, u5_mult_82_CARRYB_13__45_,
         u5_mult_82_CARRYB_13__46_, u5_mult_82_CARRYB_13__47_,
         u5_mult_82_CARRYB_13__48_, u5_mult_82_CARRYB_13__49_,
         u5_mult_82_CARRYB_13__50_, u5_mult_82_CARRYB_13__51_,
         u5_mult_82_CARRYB_14__0_, u5_mult_82_CARRYB_14__1_,
         u5_mult_82_CARRYB_14__2_, u5_mult_82_CARRYB_14__3_,
         u5_mult_82_CARRYB_14__4_, u5_mult_82_CARRYB_14__5_,
         u5_mult_82_CARRYB_14__6_, u5_mult_82_CARRYB_14__7_,
         u5_mult_82_CARRYB_14__8_, u5_mult_82_CARRYB_14__9_,
         u5_mult_82_CARRYB_14__10_, u5_mult_82_CARRYB_14__11_,
         u5_mult_82_CARRYB_14__12_, u5_mult_82_CARRYB_14__13_,
         u5_mult_82_CARRYB_14__14_, u5_mult_82_CARRYB_14__15_,
         u5_mult_82_CARRYB_14__16_, u5_mult_82_CARRYB_14__17_,
         u5_mult_82_CARRYB_14__18_, u5_mult_82_SUMB_1__2_,
         u5_mult_82_SUMB_1__3_, u5_mult_82_SUMB_1__5_, u5_mult_82_SUMB_1__6_,
         u5_mult_82_SUMB_1__7_, u5_mult_82_SUMB_1__8_, u5_mult_82_SUMB_1__9_,
         u5_mult_82_SUMB_1__11_, u5_mult_82_SUMB_1__12_,
         u5_mult_82_SUMB_1__13_, u5_mult_82_SUMB_1__14_,
         u5_mult_82_SUMB_1__15_, u5_mult_82_SUMB_1__16_,
         u5_mult_82_SUMB_1__17_, u5_mult_82_SUMB_1__19_,
         u5_mult_82_SUMB_1__20_, u5_mult_82_SUMB_1__22_,
         u5_mult_82_SUMB_1__23_, u5_mult_82_SUMB_1__24_,
         u5_mult_82_SUMB_1__25_, u5_mult_82_SUMB_1__26_,
         u5_mult_82_SUMB_1__27_, u5_mult_82_SUMB_1__29_,
         u5_mult_82_SUMB_1__30_, u5_mult_82_SUMB_1__31_,
         u5_mult_82_SUMB_1__33_, u5_mult_82_SUMB_1__35_,
         u5_mult_82_SUMB_1__36_, u5_mult_82_SUMB_1__38_,
         u5_mult_82_SUMB_1__40_, u5_mult_82_SUMB_1__42_,
         u5_mult_82_SUMB_1__44_, u5_mult_82_SUMB_1__45_,
         u5_mult_82_SUMB_1__46_, u5_mult_82_SUMB_1__47_,
         u5_mult_82_SUMB_1__48_, u5_mult_82_SUMB_1__49_,
         u5_mult_82_SUMB_1__50_, u5_mult_82_SUMB_1__51_, u5_mult_82_SUMB_2__1_,
         u5_mult_82_SUMB_2__2_, u5_mult_82_SUMB_2__3_, u5_mult_82_SUMB_2__4_,
         u5_mult_82_SUMB_2__5_, u5_mult_82_SUMB_2__6_, u5_mult_82_SUMB_2__7_,
         u5_mult_82_SUMB_2__8_, u5_mult_82_SUMB_2__9_, u5_mult_82_SUMB_2__10_,
         u5_mult_82_SUMB_2__11_, u5_mult_82_SUMB_2__12_,
         u5_mult_82_SUMB_2__13_, u5_mult_82_SUMB_2__14_,
         u5_mult_82_SUMB_2__15_, u5_mult_82_SUMB_2__16_,
         u5_mult_82_SUMB_2__17_, u5_mult_82_SUMB_2__18_,
         u5_mult_82_SUMB_2__19_, u5_mult_82_SUMB_2__20_,
         u5_mult_82_SUMB_2__21_, u5_mult_82_SUMB_2__22_,
         u5_mult_82_SUMB_2__23_, u5_mult_82_SUMB_2__24_,
         u5_mult_82_SUMB_2__25_, u5_mult_82_SUMB_2__26_,
         u5_mult_82_SUMB_2__27_, u5_mult_82_SUMB_2__28_,
         u5_mult_82_SUMB_2__29_, u5_mult_82_SUMB_2__30_,
         u5_mult_82_SUMB_2__31_, u5_mult_82_SUMB_2__32_,
         u5_mult_82_SUMB_2__33_, u5_mult_82_SUMB_2__34_,
         u5_mult_82_SUMB_2__35_, u5_mult_82_SUMB_2__37_,
         u5_mult_82_SUMB_2__38_, u5_mult_82_SUMB_2__39_,
         u5_mult_82_SUMB_2__40_, u5_mult_82_SUMB_2__41_,
         u5_mult_82_SUMB_2__42_, u5_mult_82_SUMB_2__43_,
         u5_mult_82_SUMB_2__44_, u5_mult_82_SUMB_2__45_,
         u5_mult_82_SUMB_2__46_, u5_mult_82_SUMB_2__47_,
         u5_mult_82_SUMB_2__48_, u5_mult_82_SUMB_2__49_,
         u5_mult_82_SUMB_2__50_, u5_mult_82_SUMB_2__51_, u5_mult_82_SUMB_3__1_,
         u5_mult_82_SUMB_3__2_, u5_mult_82_SUMB_3__3_, u5_mult_82_SUMB_3__4_,
         u5_mult_82_SUMB_3__5_, u5_mult_82_SUMB_3__6_, u5_mult_82_SUMB_3__7_,
         u5_mult_82_SUMB_3__8_, u5_mult_82_SUMB_3__9_, u5_mult_82_SUMB_3__10_,
         u5_mult_82_SUMB_3__11_, u5_mult_82_SUMB_3__12_,
         u5_mult_82_SUMB_3__13_, u5_mult_82_SUMB_3__14_,
         u5_mult_82_SUMB_3__15_, u5_mult_82_SUMB_3__16_,
         u5_mult_82_SUMB_3__17_, u5_mult_82_SUMB_3__18_,
         u5_mult_82_SUMB_3__19_, u5_mult_82_SUMB_3__20_,
         u5_mult_82_SUMB_3__21_, u5_mult_82_SUMB_3__22_,
         u5_mult_82_SUMB_3__23_, u5_mult_82_SUMB_3__24_,
         u5_mult_82_SUMB_3__25_, u5_mult_82_SUMB_3__26_,
         u5_mult_82_SUMB_3__27_, u5_mult_82_SUMB_3__28_,
         u5_mult_82_SUMB_3__29_, u5_mult_82_SUMB_3__30_,
         u5_mult_82_SUMB_3__31_, u5_mult_82_SUMB_3__32_,
         u5_mult_82_SUMB_3__33_, u5_mult_82_SUMB_3__34_,
         u5_mult_82_SUMB_3__37_, u5_mult_82_SUMB_3__38_,
         u5_mult_82_SUMB_3__39_, u5_mult_82_SUMB_3__40_,
         u5_mult_82_SUMB_3__41_, u5_mult_82_SUMB_3__42_,
         u5_mult_82_SUMB_3__43_, u5_mult_82_SUMB_3__44_,
         u5_mult_82_SUMB_3__45_, u5_mult_82_SUMB_3__46_,
         u5_mult_82_SUMB_3__47_, u5_mult_82_SUMB_3__48_,
         u5_mult_82_SUMB_3__49_, u5_mult_82_SUMB_3__50_,
         u5_mult_82_SUMB_3__51_, u5_mult_82_SUMB_4__1_, u5_mult_82_SUMB_4__2_,
         u5_mult_82_SUMB_4__3_, u5_mult_82_SUMB_4__4_, u5_mult_82_SUMB_4__5_,
         u5_mult_82_SUMB_4__6_, u5_mult_82_SUMB_4__7_, u5_mult_82_SUMB_4__8_,
         u5_mult_82_SUMB_4__9_, u5_mult_82_SUMB_4__10_, u5_mult_82_SUMB_4__11_,
         u5_mult_82_SUMB_4__12_, u5_mult_82_SUMB_4__13_,
         u5_mult_82_SUMB_4__14_, u5_mult_82_SUMB_4__15_,
         u5_mult_82_SUMB_4__16_, u5_mult_82_SUMB_4__17_,
         u5_mult_82_SUMB_4__18_, u5_mult_82_SUMB_4__19_,
         u5_mult_82_SUMB_4__20_, u5_mult_82_SUMB_4__21_,
         u5_mult_82_SUMB_4__22_, u5_mult_82_SUMB_4__23_,
         u5_mult_82_SUMB_4__24_, u5_mult_82_SUMB_4__25_,
         u5_mult_82_SUMB_4__26_, u5_mult_82_SUMB_4__27_,
         u5_mult_82_SUMB_4__28_, u5_mult_82_SUMB_4__29_,
         u5_mult_82_SUMB_4__30_, u5_mult_82_SUMB_4__31_,
         u5_mult_82_SUMB_4__32_, u5_mult_82_SUMB_4__33_,
         u5_mult_82_SUMB_4__34_, u5_mult_82_SUMB_4__36_,
         u5_mult_82_CARRYB_1__0_, u5_mult_82_CARRYB_1__2_,
         u5_mult_82_CARRYB_1__3_, u5_mult_82_CARRYB_1__5_,
         u5_mult_82_CARRYB_1__6_, u5_mult_82_CARRYB_1__7_,
         u5_mult_82_CARRYB_1__9_, u5_mult_82_CARRYB_1__11_,
         u5_mult_82_CARRYB_1__12_, u5_mult_82_CARRYB_1__13_,
         u5_mult_82_CARRYB_1__14_, u5_mult_82_CARRYB_1__16_,
         u5_mult_82_CARRYB_1__18_, u5_mult_82_CARRYB_1__19_,
         u5_mult_82_CARRYB_1__21_, u5_mult_82_CARRYB_1__23_,
         u5_mult_82_CARRYB_1__24_, u5_mult_82_CARRYB_1__25_,
         u5_mult_82_CARRYB_1__26_, u5_mult_82_CARRYB_1__27_,
         u5_mult_82_CARRYB_1__29_, u5_mult_82_CARRYB_1__30_,
         u5_mult_82_CARRYB_1__32_, u5_mult_82_CARRYB_1__34_,
         u5_mult_82_CARRYB_1__37_, u5_mult_82_CARRYB_1__41_,
         u5_mult_82_CARRYB_1__42_, u5_mult_82_CARRYB_1__43_,
         u5_mult_82_CARRYB_1__44_, u5_mult_82_CARRYB_1__45_,
         u5_mult_82_CARRYB_1__46_, u5_mult_82_CARRYB_1__47_,
         u5_mult_82_CARRYB_1__48_, u5_mult_82_CARRYB_1__49_,
         u5_mult_82_CARRYB_1__50_, u5_mult_82_CARRYB_2__0_,
         u5_mult_82_CARRYB_2__1_, u5_mult_82_CARRYB_2__2_,
         u5_mult_82_CARRYB_2__3_, u5_mult_82_CARRYB_2__4_,
         u5_mult_82_CARRYB_2__5_, u5_mult_82_CARRYB_2__6_,
         u5_mult_82_CARRYB_2__7_, u5_mult_82_CARRYB_2__8_,
         u5_mult_82_CARRYB_2__9_, u5_mult_82_CARRYB_2__10_,
         u5_mult_82_CARRYB_2__11_, u5_mult_82_CARRYB_2__12_,
         u5_mult_82_CARRYB_2__13_, u5_mult_82_CARRYB_2__14_,
         u5_mult_82_CARRYB_2__15_, u5_mult_82_CARRYB_2__16_,
         u5_mult_82_CARRYB_2__17_, u5_mult_82_CARRYB_2__18_,
         u5_mult_82_CARRYB_2__19_, u5_mult_82_CARRYB_2__20_,
         u5_mult_82_CARRYB_2__21_, u5_mult_82_CARRYB_2__22_,
         u5_mult_82_CARRYB_2__23_, u5_mult_82_CARRYB_2__24_,
         u5_mult_82_CARRYB_2__25_, u5_mult_82_CARRYB_2__26_,
         u5_mult_82_CARRYB_2__27_, u5_mult_82_CARRYB_2__28_,
         u5_mult_82_CARRYB_2__29_, u5_mult_82_CARRYB_2__30_,
         u5_mult_82_CARRYB_2__31_, u5_mult_82_CARRYB_2__32_,
         u5_mult_82_CARRYB_2__33_, u5_mult_82_CARRYB_2__34_,
         u5_mult_82_CARRYB_2__35_, u5_mult_82_CARRYB_2__37_,
         u5_mult_82_CARRYB_2__38_, u5_mult_82_CARRYB_2__39_,
         u5_mult_82_CARRYB_2__40_, u5_mult_82_CARRYB_2__41_,
         u5_mult_82_CARRYB_2__42_, u5_mult_82_CARRYB_2__43_,
         u5_mult_82_CARRYB_2__44_, u5_mult_82_CARRYB_2__45_,
         u5_mult_82_CARRYB_2__46_, u5_mult_82_CARRYB_2__47_,
         u5_mult_82_CARRYB_2__48_, u5_mult_82_CARRYB_2__49_,
         u5_mult_82_CARRYB_2__50_, u5_mult_82_CARRYB_2__51_,
         u5_mult_82_CARRYB_3__0_, u5_mult_82_CARRYB_3__1_,
         u5_mult_82_CARRYB_3__2_, u5_mult_82_CARRYB_3__3_,
         u5_mult_82_CARRYB_3__4_, u5_mult_82_CARRYB_3__5_,
         u5_mult_82_CARRYB_3__6_, u5_mult_82_CARRYB_3__7_,
         u5_mult_82_CARRYB_3__8_, u5_mult_82_CARRYB_3__9_,
         u5_mult_82_CARRYB_3__10_, u5_mult_82_CARRYB_3__11_,
         u5_mult_82_CARRYB_3__12_, u5_mult_82_CARRYB_3__13_,
         u5_mult_82_CARRYB_3__14_, u5_mult_82_CARRYB_3__15_,
         u5_mult_82_CARRYB_3__16_, u5_mult_82_CARRYB_3__17_,
         u5_mult_82_CARRYB_3__18_, u5_mult_82_CARRYB_3__19_,
         u5_mult_82_CARRYB_3__20_, u5_mult_82_CARRYB_3__21_,
         u5_mult_82_CARRYB_3__22_, u5_mult_82_CARRYB_3__23_,
         u5_mult_82_CARRYB_3__24_, u5_mult_82_CARRYB_3__25_,
         u5_mult_82_CARRYB_3__26_, u5_mult_82_CARRYB_3__27_,
         u5_mult_82_CARRYB_3__28_, u5_mult_82_CARRYB_3__29_,
         u5_mult_82_CARRYB_3__30_, u5_mult_82_CARRYB_3__31_,
         u5_mult_82_CARRYB_3__32_, u5_mult_82_CARRYB_3__33_,
         u5_mult_82_CARRYB_3__34_, u5_mult_82_CARRYB_3__36_,
         u5_mult_82_CARRYB_3__37_, u5_mult_82_CARRYB_3__38_,
         u5_mult_82_CARRYB_3__39_, u5_mult_82_CARRYB_3__40_,
         u5_mult_82_CARRYB_3__41_, u5_mult_82_CARRYB_3__42_,
         u5_mult_82_CARRYB_3__43_, u5_mult_82_CARRYB_3__44_,
         u5_mult_82_CARRYB_3__45_, u5_mult_82_CARRYB_3__46_,
         u5_mult_82_CARRYB_3__47_, u5_mult_82_CARRYB_3__48_,
         u5_mult_82_CARRYB_3__49_, u5_mult_82_CARRYB_3__50_,
         u5_mult_82_CARRYB_3__51_, u5_mult_82_CARRYB_4__0_,
         u5_mult_82_CARRYB_4__1_, u5_mult_82_CARRYB_4__2_,
         u5_mult_82_CARRYB_4__3_, u5_mult_82_CARRYB_4__4_,
         u5_mult_82_CARRYB_4__5_, u5_mult_82_CARRYB_4__6_,
         u5_mult_82_CARRYB_4__7_, u5_mult_82_CARRYB_4__8_,
         u5_mult_82_CARRYB_4__9_, u5_mult_82_CARRYB_4__10_,
         u5_mult_82_CARRYB_4__11_, u5_mult_82_CARRYB_4__12_,
         u5_mult_82_CARRYB_4__13_, u5_mult_82_CARRYB_4__14_,
         u5_mult_82_CARRYB_4__15_, u5_mult_82_CARRYB_4__16_,
         u5_mult_82_CARRYB_4__17_, u5_mult_82_CARRYB_4__18_,
         u5_mult_82_CARRYB_4__19_, u5_mult_82_CARRYB_4__20_,
         u5_mult_82_CARRYB_4__21_, u5_mult_82_CARRYB_4__22_,
         u5_mult_82_CARRYB_4__23_, u5_mult_82_CARRYB_4__24_,
         u5_mult_82_CARRYB_4__25_, u5_mult_82_CARRYB_4__26_,
         u5_mult_82_CARRYB_4__27_, u5_mult_82_CARRYB_4__28_,
         u5_mult_82_CARRYB_4__29_, u5_mult_82_CARRYB_4__30_,
         u5_mult_82_CARRYB_4__31_, u5_mult_82_CARRYB_4__32_,
         u5_mult_82_CARRYB_4__33_, u5_mult_82_CARRYB_4__35_,
         u5_mult_82_CARRYB_4__36_, u5_mult_82_ab_0__1_, u5_mult_82_ab_0__2_,
         u5_mult_82_ab_0__3_, u5_mult_82_ab_0__4_, u5_mult_82_ab_0__5_,
         u5_mult_82_ab_0__6_, u5_mult_82_ab_0__7_, u5_mult_82_ab_0__8_,
         u5_mult_82_ab_0__9_, u5_mult_82_ab_0__10_, u5_mult_82_ab_0__11_,
         u5_mult_82_ab_0__12_, u5_mult_82_ab_0__13_, u5_mult_82_ab_0__14_,
         u5_mult_82_ab_0__15_, u5_mult_82_ab_0__16_, u5_mult_82_ab_0__17_,
         u5_mult_82_ab_0__18_, u5_mult_82_ab_0__19_, u5_mult_82_ab_0__20_,
         u5_mult_82_ab_0__21_, u5_mult_82_ab_0__22_, u5_mult_82_ab_0__23_,
         u5_mult_82_ab_0__24_, u5_mult_82_ab_0__25_, u5_mult_82_ab_0__26_,
         u5_mult_82_ab_0__27_, u5_mult_82_ab_0__28_, u5_mult_82_ab_0__29_,
         u5_mult_82_ab_0__30_, u5_mult_82_ab_0__31_, u5_mult_82_ab_0__32_,
         u5_mult_82_ab_0__33_, u5_mult_82_ab_0__34_, u5_mult_82_ab_0__35_,
         u5_mult_82_ab_0__36_, u5_mult_82_ab_0__39_, u5_mult_82_ab_0__40_,
         u5_mult_82_ab_0__41_, u5_mult_82_ab_0__42_, u5_mult_82_ab_0__43_,
         u5_mult_82_ab_0__44_, u5_mult_82_ab_0__45_, u5_mult_82_ab_0__46_,
         u5_mult_82_ab_0__47_, u5_mult_82_ab_0__48_, u5_mult_82_ab_0__49_,
         u5_mult_82_ab_0__50_, u5_mult_82_ab_0__51_, u5_mult_82_ab_1__0_,
         u5_mult_82_ab_1__1_, u5_mult_82_ab_1__2_, u5_mult_82_ab_1__3_,
         u5_mult_82_ab_1__4_, u5_mult_82_ab_1__5_, u5_mult_82_ab_1__6_,
         u5_mult_82_ab_1__7_, u5_mult_82_ab_1__8_, u5_mult_82_ab_1__9_,
         u5_mult_82_ab_1__10_, u5_mult_82_ab_1__11_, u5_mult_82_ab_1__12_,
         u5_mult_82_ab_1__13_, u5_mult_82_ab_1__14_, u5_mult_82_ab_1__15_,
         u5_mult_82_ab_1__16_, u5_mult_82_ab_1__17_, u5_mult_82_ab_1__18_,
         u5_mult_82_ab_1__19_, u5_mult_82_ab_1__20_, u5_mult_82_ab_1__21_,
         u5_mult_82_ab_1__22_, u5_mult_82_ab_1__23_, u5_mult_82_ab_1__24_,
         u5_mult_82_ab_1__25_, u5_mult_82_ab_1__26_, u5_mult_82_ab_1__27_,
         u5_mult_82_ab_1__28_, u5_mult_82_ab_1__29_, u5_mult_82_ab_1__30_,
         u5_mult_82_ab_1__31_, u5_mult_82_ab_1__32_, u5_mult_82_ab_1__33_,
         u5_mult_82_ab_1__34_, u5_mult_82_ab_1__36_, u5_mult_82_ab_1__38_,
         u5_mult_82_ab_1__41_, u5_mult_82_ab_1__42_, u5_mult_82_ab_1__43_,
         u5_mult_82_ab_1__44_, u5_mult_82_ab_1__45_, u5_mult_82_ab_1__46_,
         u5_mult_82_ab_1__47_, u5_mult_82_ab_1__48_, u5_mult_82_ab_1__49_,
         u5_mult_82_ab_1__50_, u5_mult_82_ab_1__51_, u5_mult_82_ab_1__52_,
         u5_mult_82_ab_2__0_, u5_mult_82_ab_2__1_, u5_mult_82_ab_2__2_,
         u5_mult_82_ab_2__3_, u5_mult_82_ab_2__4_, u5_mult_82_ab_2__5_,
         u5_mult_82_ab_2__6_, u5_mult_82_ab_2__7_, u5_mult_82_ab_2__8_,
         u5_mult_82_ab_2__9_, u5_mult_82_ab_2__10_, u5_mult_82_ab_2__11_,
         u5_mult_82_ab_2__12_, u5_mult_82_ab_2__13_, u5_mult_82_ab_2__14_,
         u5_mult_82_ab_2__15_, u5_mult_82_ab_2__16_, u5_mult_82_ab_2__17_,
         u5_mult_82_ab_2__18_, u5_mult_82_ab_2__19_, u5_mult_82_ab_2__20_,
         u5_mult_82_ab_2__21_, u5_mult_82_ab_2__22_, u5_mult_82_ab_2__23_,
         u5_mult_82_ab_2__24_, u5_mult_82_ab_2__25_, u5_mult_82_ab_2__26_,
         u5_mult_82_ab_2__27_, u5_mult_82_ab_2__28_, u5_mult_82_ab_2__29_,
         u5_mult_82_ab_2__30_, u5_mult_82_ab_2__31_, u5_mult_82_ab_2__32_,
         u5_mult_82_ab_2__33_, u5_mult_82_ab_2__34_, u5_mult_82_ab_2__35_,
         u5_mult_82_ab_2__37_, u5_mult_82_ab_2__38_, u5_mult_82_ab_2__39_,
         u5_mult_82_ab_2__40_, u5_mult_82_ab_2__41_, u5_mult_82_ab_2__42_,
         u5_mult_82_ab_2__43_, u5_mult_82_ab_2__44_, u5_mult_82_ab_2__45_,
         u5_mult_82_ab_2__46_, u5_mult_82_ab_2__47_, u5_mult_82_ab_2__48_,
         u5_mult_82_ab_2__49_, u5_mult_82_ab_2__50_, u5_mult_82_ab_2__51_,
         u5_mult_82_ab_2__52_, u5_mult_82_ab_3__0_, u5_mult_82_ab_3__1_,
         u5_mult_82_ab_3__2_, u5_mult_82_ab_3__3_, u5_mult_82_ab_3__4_,
         u5_mult_82_ab_3__5_, u5_mult_82_ab_3__6_, u5_mult_82_ab_3__7_,
         u5_mult_82_ab_3__8_, u5_mult_82_ab_3__9_, u5_mult_82_ab_3__10_,
         u5_mult_82_ab_3__11_, u5_mult_82_ab_3__12_, u5_mult_82_ab_3__13_,
         u5_mult_82_ab_3__14_, u5_mult_82_ab_3__15_, u5_mult_82_ab_3__16_,
         u5_mult_82_ab_3__17_, u5_mult_82_ab_3__18_, u5_mult_82_ab_3__19_,
         u5_mult_82_ab_3__20_, u5_mult_82_ab_3__21_, u5_mult_82_ab_3__22_,
         u5_mult_82_ab_3__23_, u5_mult_82_ab_3__24_, u5_mult_82_ab_3__25_,
         u5_mult_82_ab_3__26_, u5_mult_82_ab_3__27_, u5_mult_82_ab_3__28_,
         u5_mult_82_ab_3__29_, u5_mult_82_ab_3__30_, u5_mult_82_ab_3__31_,
         u5_mult_82_ab_3__32_, u5_mult_82_ab_3__33_, u5_mult_82_ab_3__34_,
         u5_mult_82_ab_3__35_, u5_mult_82_ab_3__36_, u5_mult_82_ab_3__37_,
         u5_mult_82_ab_3__38_, u5_mult_82_ab_3__39_, u5_mult_82_ab_3__40_,
         u5_mult_82_ab_3__41_, u5_mult_82_ab_3__42_, u5_mult_82_ab_3__43_,
         u5_mult_82_ab_3__44_, u5_mult_82_ab_3__45_, u5_mult_82_ab_3__46_,
         u5_mult_82_ab_3__47_, u5_mult_82_ab_3__48_, u5_mult_82_ab_3__49_,
         u5_mult_82_ab_3__50_, u5_mult_82_ab_3__51_, u5_mult_82_ab_3__52_,
         u5_mult_82_ab_4__0_, u5_mult_82_ab_4__1_, u5_mult_82_ab_4__2_,
         u5_mult_82_ab_4__3_, u5_mult_82_ab_4__4_, u5_mult_82_ab_4__5_,
         u5_mult_82_ab_4__6_, u5_mult_82_ab_4__7_, u5_mult_82_ab_4__8_,
         u5_mult_82_ab_4__9_, u5_mult_82_ab_4__10_, u5_mult_82_ab_4__11_,
         u5_mult_82_ab_4__12_, u5_mult_82_ab_4__13_, u5_mult_82_ab_4__14_,
         u5_mult_82_ab_4__15_, u5_mult_82_ab_4__16_, u5_mult_82_ab_4__17_,
         u5_mult_82_ab_4__18_, u5_mult_82_ab_4__19_, u5_mult_82_ab_4__20_,
         u5_mult_82_ab_4__21_, u5_mult_82_ab_4__22_, u5_mult_82_ab_4__23_,
         u5_mult_82_ab_4__24_, u5_mult_82_ab_4__25_, u5_mult_82_ab_4__26_,
         u5_mult_82_ab_4__27_, u5_mult_82_ab_4__28_, u5_mult_82_ab_4__29_,
         u5_mult_82_ab_4__30_, u5_mult_82_ab_4__31_, u5_mult_82_ab_4__32_,
         u5_mult_82_ab_4__33_, u5_mult_82_ab_4__34_, u5_mult_82_ab_4__35_,
         u5_mult_82_ab_4__36_, u5_mult_82_ab_4__37_, u5_mult_82_ab_4__38_,
         u5_mult_82_ab_4__39_, u5_mult_82_ab_4__40_, u5_mult_82_ab_4__41_,
         u5_mult_82_ab_4__42_, u5_mult_82_ab_4__43_, u5_mult_82_ab_4__44_,
         u5_mult_82_ab_4__45_, u5_mult_82_ab_4__46_, u5_mult_82_ab_4__47_,
         u5_mult_82_ab_4__48_, u5_mult_82_ab_4__49_, u5_mult_82_ab_4__50_,
         u5_mult_82_ab_4__51_, u5_mult_82_ab_4__52_, u5_mult_82_ab_5__0_,
         u5_mult_82_ab_5__1_, u5_mult_82_ab_5__2_, u5_mult_82_ab_5__3_,
         u5_mult_82_ab_5__4_, u5_mult_82_ab_5__5_, u5_mult_82_ab_5__6_,
         u5_mult_82_ab_5__7_, u5_mult_82_ab_5__8_, u5_mult_82_ab_5__9_,
         u5_mult_82_ab_5__10_, u5_mult_82_ab_5__11_, u5_mult_82_ab_5__12_,
         u5_mult_82_ab_5__13_, u5_mult_82_ab_5__14_, u5_mult_82_ab_5__15_,
         u5_mult_82_ab_5__16_, u5_mult_82_ab_5__17_, u5_mult_82_ab_5__18_,
         u5_mult_82_ab_5__19_, u5_mult_82_ab_5__20_, u5_mult_82_ab_5__21_,
         u5_mult_82_ab_5__22_, u5_mult_82_ab_5__23_, u5_mult_82_ab_5__24_,
         u5_mult_82_ab_5__25_, u5_mult_82_ab_5__26_, u5_mult_82_ab_5__27_,
         u5_mult_82_ab_5__28_, u5_mult_82_ab_5__29_, u5_mult_82_ab_5__30_,
         u5_mult_82_ab_5__31_, u5_mult_82_ab_5__32_, u5_mult_82_ab_5__33_,
         u5_mult_82_ab_5__35_, u5_mult_82_ab_5__36_, u5_mult_82_ab_5__37_,
         u5_mult_82_ab_5__38_, u5_mult_82_ab_5__39_, u5_mult_82_ab_5__40_,
         u5_mult_82_ab_5__41_, u5_mult_82_ab_5__42_, u5_mult_82_ab_5__43_,
         u5_mult_82_ab_5__44_, u5_mult_82_ab_5__45_, u5_mult_82_ab_5__46_,
         u5_mult_82_ab_5__47_, u5_mult_82_ab_5__48_, u5_mult_82_ab_5__49_,
         u5_mult_82_ab_5__50_, u5_mult_82_ab_5__51_, u5_mult_82_ab_5__52_,
         u5_mult_82_ab_6__0_, u5_mult_82_ab_6__1_, u5_mult_82_ab_6__2_,
         u5_mult_82_ab_6__3_, u5_mult_82_ab_6__4_, u5_mult_82_ab_6__5_,
         u5_mult_82_ab_6__6_, u5_mult_82_ab_6__7_, u5_mult_82_ab_6__8_,
         u5_mult_82_ab_6__9_, u5_mult_82_ab_6__10_, u5_mult_82_ab_6__11_,
         u5_mult_82_ab_6__12_, u5_mult_82_ab_6__13_, u5_mult_82_ab_6__14_,
         u5_mult_82_ab_6__15_, u5_mult_82_ab_6__16_, u5_mult_82_ab_6__17_,
         u5_mult_82_ab_6__18_, u5_mult_82_ab_6__19_, u5_mult_82_ab_6__20_,
         u5_mult_82_ab_6__21_, u5_mult_82_ab_6__22_, u5_mult_82_ab_6__23_,
         u5_mult_82_ab_6__24_, u5_mult_82_ab_6__25_, u5_mult_82_ab_6__26_,
         u5_mult_82_ab_6__27_, u5_mult_82_ab_6__28_, u5_mult_82_ab_6__29_,
         u5_mult_82_ab_6__30_, u5_mult_82_ab_6__31_, u5_mult_82_ab_6__32_,
         u5_mult_82_ab_6__33_, u5_mult_82_ab_6__34_, u5_mult_82_ab_6__36_,
         u5_mult_82_ab_6__37_, u5_mult_82_ab_6__38_, u5_mult_82_ab_6__39_,
         u5_mult_82_ab_6__40_, u5_mult_82_ab_6__41_, u5_mult_82_ab_6__42_,
         u5_mult_82_ab_6__43_, u5_mult_82_ab_6__44_, u5_mult_82_ab_6__45_,
         u5_mult_82_ab_6__46_, u5_mult_82_ab_6__47_, u5_mult_82_ab_6__48_,
         u5_mult_82_ab_6__49_, u5_mult_82_ab_6__50_, u5_mult_82_ab_6__51_,
         u5_mult_82_ab_6__52_, u5_mult_82_ab_7__0_, u5_mult_82_ab_7__1_,
         u5_mult_82_ab_7__2_, u5_mult_82_ab_7__3_, u5_mult_82_ab_7__4_,
         u5_mult_82_ab_7__5_, u5_mult_82_ab_7__6_, u5_mult_82_ab_7__7_,
         u5_mult_82_ab_7__8_, u5_mult_82_ab_7__9_, u5_mult_82_ab_7__10_,
         u5_mult_82_ab_7__11_, u5_mult_82_ab_7__12_, u5_mult_82_ab_7__13_,
         u5_mult_82_ab_7__14_, u5_mult_82_ab_7__15_, u5_mult_82_ab_7__16_,
         u5_mult_82_ab_7__17_, u5_mult_82_ab_7__18_, u5_mult_82_ab_7__19_,
         u5_mult_82_ab_7__20_, u5_mult_82_ab_7__21_, u5_mult_82_ab_7__22_,
         u5_mult_82_ab_7__23_, u5_mult_82_ab_7__24_, u5_mult_82_ab_7__25_,
         u5_mult_82_ab_7__26_, u5_mult_82_ab_7__27_, u5_mult_82_ab_7__28_,
         u5_mult_82_ab_7__29_, u5_mult_82_ab_7__30_, u5_mult_82_ab_7__31_,
         u5_mult_82_ab_7__32_, u5_mult_82_ab_7__33_, u5_mult_82_ab_7__34_,
         u5_mult_82_ab_7__35_, u5_mult_82_ab_7__36_, u5_mult_82_ab_7__37_,
         u5_mult_82_ab_7__38_, u5_mult_82_ab_7__39_, u5_mult_82_ab_7__40_,
         u5_mult_82_ab_7__41_, u5_mult_82_ab_7__42_, u5_mult_82_ab_7__43_,
         u5_mult_82_ab_7__44_, u5_mult_82_ab_7__45_, u5_mult_82_ab_7__46_,
         u5_mult_82_ab_7__47_, u5_mult_82_ab_7__48_, u5_mult_82_ab_7__49_,
         u5_mult_82_ab_7__50_, u5_mult_82_ab_7__51_, u5_mult_82_ab_7__52_,
         u5_mult_82_ab_8__0_, u5_mult_82_ab_8__1_, u5_mult_82_ab_8__2_,
         u5_mult_82_ab_8__3_, u5_mult_82_ab_8__4_, u5_mult_82_ab_8__5_,
         u5_mult_82_ab_8__6_, u5_mult_82_ab_8__7_, u5_mult_82_ab_8__8_,
         u5_mult_82_ab_8__9_, u5_mult_82_ab_8__10_, u5_mult_82_ab_8__11_,
         u5_mult_82_ab_8__12_, u5_mult_82_ab_8__13_, u5_mult_82_ab_8__14_,
         u5_mult_82_ab_8__15_, u5_mult_82_ab_8__16_, u5_mult_82_ab_8__17_,
         u5_mult_82_ab_8__18_, u5_mult_82_ab_8__19_, u5_mult_82_ab_8__20_,
         u5_mult_82_ab_8__21_, u5_mult_82_ab_8__22_, u5_mult_82_ab_8__23_,
         u5_mult_82_ab_8__24_, u5_mult_82_ab_8__25_, u5_mult_82_ab_8__26_,
         u5_mult_82_ab_8__27_, u5_mult_82_ab_8__28_, u5_mult_82_ab_8__29_,
         u5_mult_82_ab_8__30_, u5_mult_82_ab_8__31_, u5_mult_82_ab_8__32_,
         u5_mult_82_ab_8__33_, u5_mult_82_ab_8__34_, u5_mult_82_ab_8__35_,
         u5_mult_82_ab_8__36_, u5_mult_82_ab_8__37_, u5_mult_82_ab_8__38_,
         u5_mult_82_ab_8__39_, u5_mult_82_ab_8__40_, u5_mult_82_ab_8__41_,
         u5_mult_82_ab_8__42_, u5_mult_82_ab_8__43_, u5_mult_82_ab_8__44_,
         u5_mult_82_ab_8__45_, u5_mult_82_ab_8__46_, u5_mult_82_ab_8__47_,
         u5_mult_82_ab_8__48_, u5_mult_82_ab_8__49_, u5_mult_82_ab_8__50_,
         u5_mult_82_ab_8__51_, u5_mult_82_ab_8__52_, u5_mult_82_ab_9__0_,
         u5_mult_82_ab_9__1_, u5_mult_82_ab_9__2_, u5_mult_82_ab_9__3_,
         u5_mult_82_ab_9__4_, u5_mult_82_ab_9__5_, u5_mult_82_ab_9__6_,
         u5_mult_82_ab_9__7_, u5_mult_82_ab_9__8_, u5_mult_82_ab_9__9_,
         u5_mult_82_ab_9__10_, u5_mult_82_ab_9__11_, u5_mult_82_ab_9__12_,
         u5_mult_82_ab_9__13_, u5_mult_82_ab_9__14_, u5_mult_82_ab_9__15_,
         u5_mult_82_ab_9__16_, u5_mult_82_ab_9__17_, u5_mult_82_ab_9__18_,
         u5_mult_82_ab_9__19_, u5_mult_82_ab_9__20_, u5_mult_82_ab_9__21_,
         u5_mult_82_ab_9__22_, u5_mult_82_ab_9__23_, u5_mult_82_ab_9__24_,
         u5_mult_82_ab_9__25_, u5_mult_82_ab_9__26_, u5_mult_82_ab_9__27_,
         u5_mult_82_ab_9__28_, u5_mult_82_ab_9__29_, u5_mult_82_ab_9__30_,
         u5_mult_82_ab_9__31_, u5_mult_82_ab_9__32_, u5_mult_82_ab_9__33_,
         u5_mult_82_ab_9__34_, u5_mult_82_ab_9__35_, u5_mult_82_ab_9__36_,
         u5_mult_82_ab_9__37_, u5_mult_82_ab_9__38_, u5_mult_82_ab_9__39_,
         u5_mult_82_ab_9__40_, u5_mult_82_ab_9__41_, u5_mult_82_ab_9__42_,
         u5_mult_82_ab_9__43_, u5_mult_82_ab_9__44_, u5_mult_82_ab_9__45_,
         u5_mult_82_ab_9__46_, u5_mult_82_ab_9__47_, u5_mult_82_ab_9__48_,
         u5_mult_82_ab_9__49_, u5_mult_82_ab_9__50_, u5_mult_82_ab_9__51_,
         u5_mult_82_ab_9__52_, u5_mult_82_ab_10__0_, u5_mult_82_ab_10__1_,
         u5_mult_82_ab_10__2_, u5_mult_82_ab_10__3_, u5_mult_82_ab_10__4_,
         u5_mult_82_ab_10__5_, u5_mult_82_ab_10__6_, u5_mult_82_ab_10__7_,
         u5_mult_82_ab_10__8_, u5_mult_82_ab_10__9_, u5_mult_82_ab_10__10_,
         u5_mult_82_ab_10__11_, u5_mult_82_ab_10__12_, u5_mult_82_ab_10__13_,
         u5_mult_82_ab_10__14_, u5_mult_82_ab_10__15_, u5_mult_82_ab_10__16_,
         u5_mult_82_ab_10__17_, u5_mult_82_ab_10__18_, u5_mult_82_ab_10__19_,
         u5_mult_82_ab_10__20_, u5_mult_82_ab_10__21_, u5_mult_82_ab_10__22_,
         u5_mult_82_ab_10__23_, u5_mult_82_ab_10__24_, u5_mult_82_ab_10__25_,
         u5_mult_82_ab_10__26_, u5_mult_82_ab_10__27_, u5_mult_82_ab_10__28_,
         u5_mult_82_ab_10__29_, u5_mult_82_ab_10__30_, u5_mult_82_ab_10__31_,
         u5_mult_82_ab_10__32_, u5_mult_82_ab_10__33_, u5_mult_82_ab_10__34_,
         u5_mult_82_ab_10__35_, u5_mult_82_ab_10__36_, u5_mult_82_ab_10__37_,
         u5_mult_82_ab_10__38_, u5_mult_82_ab_10__39_, u5_mult_82_ab_10__40_,
         u5_mult_82_ab_10__41_, u5_mult_82_ab_10__42_, u5_mult_82_ab_10__43_,
         u5_mult_82_ab_10__44_, u5_mult_82_ab_10__45_, u5_mult_82_ab_10__46_,
         u5_mult_82_ab_10__47_, u5_mult_82_ab_10__48_, u5_mult_82_ab_10__49_,
         u5_mult_82_ab_10__50_, u5_mult_82_ab_10__51_, u5_mult_82_ab_10__52_,
         u5_mult_82_ab_11__0_, u5_mult_82_ab_11__1_, u5_mult_82_ab_11__2_,
         u5_mult_82_ab_11__3_, u5_mult_82_ab_11__4_, u5_mult_82_ab_11__5_,
         u5_mult_82_ab_11__6_, u5_mult_82_ab_11__7_, u5_mult_82_ab_11__8_,
         u5_mult_82_ab_11__9_, u5_mult_82_ab_11__10_, u5_mult_82_ab_11__11_,
         u5_mult_82_ab_11__12_, u5_mult_82_ab_11__13_, u5_mult_82_ab_11__14_,
         u5_mult_82_ab_11__15_, u5_mult_82_ab_11__16_, u5_mult_82_ab_11__17_,
         u5_mult_82_ab_11__18_, u5_mult_82_ab_11__19_, u5_mult_82_ab_11__20_,
         u5_mult_82_ab_11__21_, u5_mult_82_ab_11__22_, u5_mult_82_ab_11__23_,
         u5_mult_82_ab_11__24_, u5_mult_82_ab_11__25_, u5_mult_82_ab_11__26_,
         u5_mult_82_ab_11__27_, u5_mult_82_ab_11__28_, u5_mult_82_ab_11__29_,
         u5_mult_82_ab_11__30_, u5_mult_82_ab_11__31_, u5_mult_82_ab_11__32_,
         u5_mult_82_ab_11__33_, u5_mult_82_ab_11__34_, u5_mult_82_ab_11__35_,
         u5_mult_82_ab_11__36_, u5_mult_82_ab_11__37_, u5_mult_82_ab_11__38_,
         u5_mult_82_ab_11__39_, u5_mult_82_ab_11__40_, u5_mult_82_ab_11__41_,
         u5_mult_82_ab_11__42_, u5_mult_82_ab_11__43_, u5_mult_82_ab_11__44_,
         u5_mult_82_ab_11__45_, u5_mult_82_ab_11__46_, u5_mult_82_ab_11__47_,
         u5_mult_82_ab_11__48_, u5_mult_82_ab_11__49_, u5_mult_82_ab_11__50_,
         u5_mult_82_ab_11__51_, u5_mult_82_ab_11__52_, u5_mult_82_ab_12__0_,
         u5_mult_82_ab_12__1_, u5_mult_82_ab_12__2_, u5_mult_82_ab_12__3_,
         u5_mult_82_ab_12__4_, u5_mult_82_ab_12__5_, u5_mult_82_ab_12__6_,
         u5_mult_82_ab_12__7_, u5_mult_82_ab_12__8_, u5_mult_82_ab_12__9_,
         u5_mult_82_ab_12__10_, u5_mult_82_ab_12__11_, u5_mult_82_ab_12__12_,
         u5_mult_82_ab_12__13_, u5_mult_82_ab_12__14_, u5_mult_82_ab_12__15_,
         u5_mult_82_ab_12__16_, u5_mult_82_ab_12__17_, u5_mult_82_ab_12__18_,
         u5_mult_82_ab_12__19_, u5_mult_82_ab_12__20_, u5_mult_82_ab_12__21_,
         u5_mult_82_ab_12__22_, u5_mult_82_ab_12__23_, u5_mult_82_ab_12__24_,
         u5_mult_82_ab_12__25_, u5_mult_82_ab_12__26_, u5_mult_82_ab_12__27_,
         u5_mult_82_ab_12__28_, u5_mult_82_ab_12__29_, u5_mult_82_ab_12__30_,
         u5_mult_82_ab_12__31_, u5_mult_82_ab_12__32_, u5_mult_82_ab_12__33_,
         u5_mult_82_ab_12__34_, u5_mult_82_ab_12__35_, u5_mult_82_ab_12__36_,
         u5_mult_82_ab_12__37_, u5_mult_82_ab_12__38_, u5_mult_82_ab_12__39_,
         u5_mult_82_ab_12__40_, u5_mult_82_ab_12__41_, u5_mult_82_ab_12__42_,
         u5_mult_82_ab_12__43_, u5_mult_82_ab_12__44_, u5_mult_82_ab_12__45_,
         u5_mult_82_ab_12__46_, u5_mult_82_ab_12__47_, u5_mult_82_ab_12__48_,
         u5_mult_82_ab_12__49_, u5_mult_82_ab_12__50_, u5_mult_82_ab_12__51_,
         u5_mult_82_ab_12__52_, u5_mult_82_ab_13__0_, u5_mult_82_ab_13__1_,
         u5_mult_82_ab_13__2_, u5_mult_82_ab_13__3_, u5_mult_82_ab_13__4_,
         u5_mult_82_ab_13__5_, u5_mult_82_ab_13__6_, u5_mult_82_ab_13__7_,
         u5_mult_82_ab_13__8_, u5_mult_82_ab_13__9_, u5_mult_82_ab_13__10_,
         u5_mult_82_ab_13__11_, u5_mult_82_ab_13__12_, u5_mult_82_ab_13__13_,
         u5_mult_82_ab_13__14_, u5_mult_82_ab_13__15_, u5_mult_82_ab_13__16_,
         u5_mult_82_ab_13__17_, u5_mult_82_ab_13__18_, u5_mult_82_ab_13__19_,
         u5_mult_82_ab_13__20_, u5_mult_82_ab_13__21_, u5_mult_82_ab_13__22_,
         u5_mult_82_ab_13__23_, u5_mult_82_ab_13__24_, u5_mult_82_ab_13__25_,
         u5_mult_82_ab_13__26_, u5_mult_82_ab_13__27_, u5_mult_82_ab_13__28_,
         u5_mult_82_ab_13__29_, u5_mult_82_ab_13__30_, u5_mult_82_ab_13__31_,
         u5_mult_82_ab_13__32_, u5_mult_82_ab_13__33_, u5_mult_82_ab_13__34_,
         u5_mult_82_ab_13__35_, u5_mult_82_ab_13__36_, u5_mult_82_ab_13__37_,
         u5_mult_82_ab_13__38_, u5_mult_82_ab_13__39_, u5_mult_82_ab_13__40_,
         u5_mult_82_ab_13__41_, u5_mult_82_ab_13__42_, u5_mult_82_ab_13__43_,
         u5_mult_82_ab_13__44_, u5_mult_82_ab_13__45_, u5_mult_82_ab_13__46_,
         u5_mult_82_ab_13__47_, u5_mult_82_ab_13__48_, u5_mult_82_ab_13__49_,
         u5_mult_82_ab_13__50_, u5_mult_82_ab_13__51_, u5_mult_82_ab_13__52_,
         u5_mult_82_ab_14__0_, u5_mult_82_ab_14__1_, u5_mult_82_ab_14__2_,
         u5_mult_82_ab_14__3_, u5_mult_82_ab_14__4_, u5_mult_82_ab_14__5_,
         u5_mult_82_ab_14__6_, u5_mult_82_ab_14__7_, u5_mult_82_ab_14__8_,
         u5_mult_82_ab_14__9_, u5_mult_82_ab_14__10_, u5_mult_82_ab_14__11_,
         u5_mult_82_ab_14__12_, u5_mult_82_ab_14__13_, u5_mult_82_ab_14__14_,
         u5_mult_82_ab_14__15_, u5_mult_82_ab_14__16_, u5_mult_82_ab_14__17_,
         u5_mult_82_ab_14__18_, u5_mult_82_ab_14__19_, u5_mult_82_ab_14__20_,
         u5_mult_82_ab_14__21_, u5_mult_82_ab_14__22_, u5_mult_82_ab_14__23_,
         u5_mult_82_ab_14__24_, u5_mult_82_ab_14__25_, u5_mult_82_ab_14__26_,
         u5_mult_82_ab_14__27_, u5_mult_82_ab_14__28_, u5_mult_82_ab_14__29_,
         u5_mult_82_ab_14__30_, u5_mult_82_ab_14__31_, u5_mult_82_ab_14__32_,
         u5_mult_82_ab_14__33_, u5_mult_82_ab_14__34_, u5_mult_82_ab_14__35_,
         u5_mult_82_ab_14__36_, u5_mult_82_ab_14__37_, u5_mult_82_ab_14__38_,
         u5_mult_82_ab_14__39_, u5_mult_82_ab_14__40_, u5_mult_82_ab_14__41_,
         u5_mult_82_ab_14__42_, u5_mult_82_ab_14__43_, u5_mult_82_ab_14__44_,
         u5_mult_82_ab_14__45_, u5_mult_82_ab_14__46_, u5_mult_82_ab_14__47_,
         u5_mult_82_ab_14__48_, u5_mult_82_ab_14__49_, u5_mult_82_ab_14__50_,
         u5_mult_82_ab_14__51_, u5_mult_82_ab_14__52_, u5_mult_82_ab_15__0_,
         u5_mult_82_ab_15__1_, u5_mult_82_ab_15__2_, u5_mult_82_ab_15__3_,
         u5_mult_82_ab_15__4_, u5_mult_82_ab_15__5_, u5_mult_82_ab_15__6_,
         u5_mult_82_ab_15__7_, u5_mult_82_ab_15__8_, u5_mult_82_ab_15__9_,
         u5_mult_82_ab_15__10_, u5_mult_82_ab_15__11_, u5_mult_82_ab_15__12_,
         u5_mult_82_ab_15__13_, u5_mult_82_ab_15__14_, u5_mult_82_ab_15__15_,
         u5_mult_82_ab_15__16_, u5_mult_82_ab_15__17_, u5_mult_82_ab_15__18_,
         u5_mult_82_ab_15__19_, u5_mult_82_ab_15__20_, u5_mult_82_ab_15__21_,
         u5_mult_82_ab_15__22_, u5_mult_82_ab_15__23_, u5_mult_82_ab_15__24_,
         u5_mult_82_ab_15__25_, u5_mult_82_ab_15__26_, u5_mult_82_ab_15__27_,
         u5_mult_82_ab_15__28_, u5_mult_82_ab_15__29_, u5_mult_82_ab_15__30_,
         u5_mult_82_ab_15__31_, u5_mult_82_ab_15__32_, u5_mult_82_ab_15__33_,
         u5_mult_82_ab_15__34_, u5_mult_82_ab_15__35_, u5_mult_82_ab_15__36_,
         u5_mult_82_ab_15__37_, u5_mult_82_ab_15__38_, u5_mult_82_ab_15__39_,
         u5_mult_82_ab_15__40_, u5_mult_82_ab_15__41_, u5_mult_82_ab_15__42_,
         u5_mult_82_ab_15__43_, u5_mult_82_ab_15__44_, u5_mult_82_ab_15__45_,
         u5_mult_82_ab_15__46_, u5_mult_82_ab_15__47_, u5_mult_82_ab_15__48_,
         u5_mult_82_ab_15__49_, u5_mult_82_ab_15__50_, u5_mult_82_ab_15__51_,
         u5_mult_82_ab_15__52_, u5_mult_82_ab_16__0_, u5_mult_82_ab_16__1_,
         u5_mult_82_ab_16__2_, u5_mult_82_ab_16__3_, u5_mult_82_ab_16__4_,
         u5_mult_82_ab_16__5_, u5_mult_82_ab_16__6_, u5_mult_82_ab_16__7_,
         u5_mult_82_ab_16__8_, u5_mult_82_ab_16__9_, u5_mult_82_ab_16__10_,
         u5_mult_82_ab_16__11_, u5_mult_82_ab_16__12_, u5_mult_82_ab_16__13_,
         u5_mult_82_ab_16__14_, u5_mult_82_ab_16__15_, u5_mult_82_ab_16__16_,
         u5_mult_82_ab_16__17_, u5_mult_82_ab_16__18_, u5_mult_82_ab_16__19_,
         u5_mult_82_ab_16__20_, u5_mult_82_ab_16__21_, u5_mult_82_ab_16__22_,
         u5_mult_82_ab_16__23_, u5_mult_82_ab_16__24_, u5_mult_82_ab_16__25_,
         u5_mult_82_ab_16__26_, u5_mult_82_ab_16__27_, u5_mult_82_ab_16__28_,
         u5_mult_82_ab_16__29_, u5_mult_82_ab_16__30_, u5_mult_82_ab_16__31_,
         u5_mult_82_ab_16__32_, u5_mult_82_ab_16__33_, u5_mult_82_ab_16__34_,
         u5_mult_82_ab_16__35_, u5_mult_82_ab_16__36_, u5_mult_82_ab_16__37_,
         u5_mult_82_ab_16__38_, u5_mult_82_ab_16__39_, u5_mult_82_ab_16__40_,
         u5_mult_82_ab_16__41_, u5_mult_82_ab_16__42_, u5_mult_82_ab_16__43_,
         u5_mult_82_ab_16__44_, u5_mult_82_ab_16__45_, u5_mult_82_ab_16__46_,
         u5_mult_82_ab_16__47_, u5_mult_82_ab_16__48_, u5_mult_82_ab_16__49_,
         u5_mult_82_ab_16__50_, u5_mult_82_ab_16__51_, u5_mult_82_ab_16__52_,
         u5_mult_82_ab_17__0_, u5_mult_82_ab_17__1_, u5_mult_82_ab_17__2_,
         u5_mult_82_ab_17__3_, u5_mult_82_ab_17__4_, u5_mult_82_ab_17__5_,
         u5_mult_82_ab_17__6_, u5_mult_82_ab_17__7_, u5_mult_82_ab_17__8_,
         u5_mult_82_ab_17__9_, u5_mult_82_ab_17__10_, u5_mult_82_ab_17__11_,
         u5_mult_82_ab_17__12_, u5_mult_82_ab_17__13_, u5_mult_82_ab_17__14_,
         u5_mult_82_ab_17__15_, u5_mult_82_ab_17__16_, u5_mult_82_ab_17__17_,
         u5_mult_82_ab_17__18_, u5_mult_82_ab_17__19_, u5_mult_82_ab_17__20_,
         u5_mult_82_ab_17__21_, u5_mult_82_ab_17__22_, u5_mult_82_ab_17__23_,
         u5_mult_82_ab_17__24_, u5_mult_82_ab_17__25_, u5_mult_82_ab_17__26_,
         u5_mult_82_ab_17__27_, u5_mult_82_ab_17__28_, u5_mult_82_ab_17__29_,
         u5_mult_82_ab_17__30_, u5_mult_82_ab_17__31_, u5_mult_82_ab_17__32_,
         u5_mult_82_ab_17__33_, u5_mult_82_ab_17__34_, u5_mult_82_ab_17__35_,
         u5_mult_82_ab_17__36_, u5_mult_82_ab_17__37_, u5_mult_82_ab_17__38_,
         u5_mult_82_ab_17__39_, u5_mult_82_ab_17__40_, u5_mult_82_ab_17__41_,
         u5_mult_82_ab_17__42_, u5_mult_82_ab_17__43_, u5_mult_82_ab_17__44_,
         u5_mult_82_ab_17__45_, u5_mult_82_ab_17__46_, u5_mult_82_ab_17__47_,
         u5_mult_82_ab_17__48_, u5_mult_82_ab_17__49_, u5_mult_82_ab_17__50_,
         u5_mult_82_ab_17__51_, u5_mult_82_ab_17__52_, u5_mult_82_ab_18__0_,
         u5_mult_82_ab_18__1_, u5_mult_82_ab_18__2_, u5_mult_82_ab_18__3_,
         u5_mult_82_ab_18__4_, u5_mult_82_ab_18__5_, u5_mult_82_ab_18__6_,
         u5_mult_82_ab_18__7_, u5_mult_82_ab_18__8_, u5_mult_82_ab_18__9_,
         u5_mult_82_ab_18__10_, u5_mult_82_ab_18__11_, u5_mult_82_ab_18__12_,
         u5_mult_82_ab_18__13_, u5_mult_82_ab_18__14_, u5_mult_82_ab_18__15_,
         u5_mult_82_ab_18__16_, u5_mult_82_ab_18__17_, u5_mult_82_ab_18__18_,
         u5_mult_82_ab_18__19_, u5_mult_82_ab_18__20_, u5_mult_82_ab_18__21_,
         u5_mult_82_ab_18__22_, u5_mult_82_ab_18__23_, u5_mult_82_ab_18__24_,
         u5_mult_82_ab_18__25_, u5_mult_82_ab_18__26_, u5_mult_82_ab_18__27_,
         u5_mult_82_ab_18__28_, u5_mult_82_ab_18__29_, u5_mult_82_ab_18__30_,
         u5_mult_82_ab_18__31_, u5_mult_82_ab_18__32_, u5_mult_82_ab_18__33_,
         u5_mult_82_ab_18__34_, u5_mult_82_ab_18__35_, u5_mult_82_ab_18__36_,
         u5_mult_82_ab_18__37_, u5_mult_82_ab_18__38_, u5_mult_82_ab_18__39_,
         u5_mult_82_ab_18__40_, u5_mult_82_ab_18__41_, u5_mult_82_ab_18__42_,
         u5_mult_82_ab_18__43_, u5_mult_82_ab_18__44_, u5_mult_82_ab_18__45_,
         u5_mult_82_ab_18__46_, u5_mult_82_ab_18__47_, u5_mult_82_ab_18__48_,
         u5_mult_82_ab_18__49_, u5_mult_82_ab_18__50_, u5_mult_82_ab_18__51_,
         u5_mult_82_ab_18__52_, u5_mult_82_ab_19__0_, u5_mult_82_ab_19__1_,
         u5_mult_82_ab_19__2_, u5_mult_82_ab_19__3_, u5_mult_82_ab_19__4_,
         u5_mult_82_ab_19__5_, u5_mult_82_ab_19__6_, u5_mult_82_ab_19__7_,
         u5_mult_82_ab_19__8_, u5_mult_82_ab_19__9_, u5_mult_82_ab_19__10_,
         u5_mult_82_ab_19__11_, u5_mult_82_ab_19__12_, u5_mult_82_ab_19__13_,
         u5_mult_82_ab_19__14_, u5_mult_82_ab_19__15_, u5_mult_82_ab_19__16_,
         u5_mult_82_ab_19__17_, u5_mult_82_ab_19__18_, u5_mult_82_ab_19__19_,
         u5_mult_82_ab_19__20_, u5_mult_82_ab_19__21_, u5_mult_82_ab_19__22_,
         u5_mult_82_ab_19__23_, u5_mult_82_ab_19__24_, u5_mult_82_ab_19__25_,
         u5_mult_82_ab_19__26_, u5_mult_82_ab_19__27_, u5_mult_82_ab_19__28_,
         u5_mult_82_ab_19__29_, u5_mult_82_ab_19__30_, u5_mult_82_ab_19__31_,
         u5_mult_82_ab_19__32_, u5_mult_82_ab_19__33_, u5_mult_82_ab_19__34_,
         u5_mult_82_ab_19__35_, u5_mult_82_ab_19__36_, u5_mult_82_ab_19__37_,
         u5_mult_82_ab_19__38_, u5_mult_82_ab_19__39_, u5_mult_82_ab_19__40_,
         u5_mult_82_ab_19__41_, u5_mult_82_ab_19__42_, u5_mult_82_ab_19__43_,
         u5_mult_82_ab_19__44_, u5_mult_82_ab_19__45_, u5_mult_82_ab_19__46_,
         u5_mult_82_ab_19__47_, u5_mult_82_ab_19__48_, u5_mult_82_ab_19__49_,
         u5_mult_82_ab_19__50_, u5_mult_82_ab_19__51_, u5_mult_82_ab_19__52_,
         u5_mult_82_ab_20__0_, u5_mult_82_ab_20__1_, u5_mult_82_ab_20__2_,
         u5_mult_82_ab_20__3_, u5_mult_82_ab_20__4_, u5_mult_82_ab_20__5_,
         u5_mult_82_ab_20__6_, u5_mult_82_ab_20__7_, u5_mult_82_ab_20__8_,
         u5_mult_82_ab_20__9_, u5_mult_82_ab_20__10_, u5_mult_82_ab_20__11_,
         u5_mult_82_ab_20__12_, u5_mult_82_ab_20__13_, u5_mult_82_ab_20__14_,
         u5_mult_82_ab_20__15_, u5_mult_82_ab_20__16_, u5_mult_82_ab_20__17_,
         u5_mult_82_ab_20__18_, u5_mult_82_ab_20__19_, u5_mult_82_ab_20__20_,
         u5_mult_82_ab_20__21_, u5_mult_82_ab_20__22_, u5_mult_82_ab_20__23_,
         u5_mult_82_ab_20__24_, u5_mult_82_ab_20__25_, u5_mult_82_ab_20__26_,
         u5_mult_82_ab_20__27_, u5_mult_82_ab_20__28_, u5_mult_82_ab_20__29_,
         u5_mult_82_ab_20__30_, u5_mult_82_ab_20__31_, u5_mult_82_ab_20__32_,
         u5_mult_82_ab_20__33_, u5_mult_82_ab_20__34_, u5_mult_82_ab_20__35_,
         u5_mult_82_ab_20__36_, u5_mult_82_ab_20__37_, u5_mult_82_ab_20__38_,
         u5_mult_82_ab_20__39_, u5_mult_82_ab_20__40_, u5_mult_82_ab_20__41_,
         u5_mult_82_ab_20__42_, u5_mult_82_ab_20__43_, u5_mult_82_ab_20__44_,
         u5_mult_82_ab_20__45_, u5_mult_82_ab_20__46_, u5_mult_82_ab_20__47_,
         u5_mult_82_ab_20__48_, u5_mult_82_ab_20__49_, u5_mult_82_ab_20__50_,
         u5_mult_82_ab_20__51_, u5_mult_82_ab_20__52_, u5_mult_82_ab_21__0_,
         u5_mult_82_ab_21__1_, u5_mult_82_ab_21__2_, u5_mult_82_ab_21__3_,
         u5_mult_82_ab_21__4_, u5_mult_82_ab_21__5_, u5_mult_82_ab_21__6_,
         u5_mult_82_ab_21__7_, u5_mult_82_ab_21__8_, u5_mult_82_ab_21__9_,
         u5_mult_82_ab_21__10_, u5_mult_82_ab_21__11_, u5_mult_82_ab_21__12_,
         u5_mult_82_ab_21__13_, u5_mult_82_ab_21__14_, u5_mult_82_ab_21__15_,
         u5_mult_82_ab_21__16_, u5_mult_82_ab_21__17_, u5_mult_82_ab_21__18_,
         u5_mult_82_ab_21__19_, u5_mult_82_ab_21__20_, u5_mult_82_ab_21__21_,
         u5_mult_82_ab_21__22_, u5_mult_82_ab_21__23_, u5_mult_82_ab_21__24_,
         u5_mult_82_ab_21__25_, u5_mult_82_ab_21__26_, u5_mult_82_ab_21__27_,
         u5_mult_82_ab_21__28_, u5_mult_82_ab_21__29_, u5_mult_82_ab_21__30_,
         u5_mult_82_ab_21__31_, u5_mult_82_ab_21__32_, u5_mult_82_ab_21__33_,
         u5_mult_82_ab_21__34_, u5_mult_82_ab_21__35_, u5_mult_82_ab_21__36_,
         u5_mult_82_ab_21__37_, u5_mult_82_ab_21__38_, u5_mult_82_ab_21__39_,
         u5_mult_82_ab_21__40_, u5_mult_82_ab_21__41_, u5_mult_82_ab_21__42_,
         u5_mult_82_ab_21__43_, u5_mult_82_ab_21__44_, u5_mult_82_ab_21__45_,
         u5_mult_82_ab_21__46_, u5_mult_82_ab_21__47_, u5_mult_82_ab_21__48_,
         u5_mult_82_ab_21__49_, u5_mult_82_ab_21__50_, u5_mult_82_ab_21__51_,
         u5_mult_82_ab_21__52_, u5_mult_82_ab_22__0_, u5_mult_82_ab_22__1_,
         u5_mult_82_ab_22__2_, u5_mult_82_ab_22__3_, u5_mult_82_ab_22__4_,
         u5_mult_82_ab_22__5_, u5_mult_82_ab_22__6_, u5_mult_82_ab_22__7_,
         u5_mult_82_ab_22__8_, u5_mult_82_ab_22__9_, u5_mult_82_ab_22__10_,
         u5_mult_82_ab_22__11_, u5_mult_82_ab_22__12_, u5_mult_82_ab_22__13_,
         u5_mult_82_ab_22__14_, u5_mult_82_ab_22__15_, u5_mult_82_ab_22__16_,
         u5_mult_82_ab_22__17_, u5_mult_82_ab_22__18_, u5_mult_82_ab_22__19_,
         u5_mult_82_ab_22__20_, u5_mult_82_ab_22__21_, u5_mult_82_ab_22__22_,
         u5_mult_82_ab_22__23_, u5_mult_82_ab_22__24_, u5_mult_82_ab_22__25_,
         u5_mult_82_ab_22__26_, u5_mult_82_ab_22__27_, u5_mult_82_ab_22__28_,
         u5_mult_82_ab_22__29_, u5_mult_82_ab_22__30_, u5_mult_82_ab_22__31_,
         u5_mult_82_ab_22__32_, u5_mult_82_ab_22__33_, u5_mult_82_ab_22__34_,
         u5_mult_82_ab_22__35_, u5_mult_82_ab_22__36_, u5_mult_82_ab_22__37_,
         u5_mult_82_ab_22__38_, u5_mult_82_ab_22__39_, u5_mult_82_ab_22__40_,
         u5_mult_82_ab_22__41_, u5_mult_82_ab_22__42_, u5_mult_82_ab_22__43_,
         u5_mult_82_ab_22__44_, u5_mult_82_ab_22__45_, u5_mult_82_ab_22__46_,
         u5_mult_82_ab_22__47_, u5_mult_82_ab_22__48_, u5_mult_82_ab_22__49_,
         u5_mult_82_ab_22__50_, u5_mult_82_ab_22__51_, u5_mult_82_ab_22__52_,
         u5_mult_82_ab_23__0_, u5_mult_82_ab_23__1_, u5_mult_82_ab_23__2_,
         u5_mult_82_ab_23__3_, u5_mult_82_ab_23__4_, u5_mult_82_ab_23__5_,
         u5_mult_82_ab_23__6_, u5_mult_82_ab_23__7_, u5_mult_82_ab_23__8_,
         u5_mult_82_ab_23__9_, u5_mult_82_ab_23__10_, u5_mult_82_ab_23__11_,
         u5_mult_82_ab_23__12_, u5_mult_82_ab_23__13_, u5_mult_82_ab_23__14_,
         u5_mult_82_ab_23__15_, u5_mult_82_ab_23__16_, u5_mult_82_ab_23__17_,
         u5_mult_82_ab_23__18_, u5_mult_82_ab_23__19_, u5_mult_82_ab_23__20_,
         u5_mult_82_ab_23__21_, u5_mult_82_ab_23__22_, u5_mult_82_ab_23__24_,
         u5_mult_82_ab_23__25_, u5_mult_82_ab_23__26_, u5_mult_82_ab_23__27_,
         u5_mult_82_ab_23__28_, u5_mult_82_ab_23__29_, u5_mult_82_ab_23__30_,
         u5_mult_82_ab_23__31_, u5_mult_82_ab_23__32_, u5_mult_82_ab_23__33_,
         u5_mult_82_ab_23__34_, u5_mult_82_ab_23__35_, u5_mult_82_ab_23__36_,
         u5_mult_82_ab_23__37_, u5_mult_82_ab_23__38_, u5_mult_82_ab_23__39_,
         u5_mult_82_ab_23__40_, u5_mult_82_ab_23__41_, u5_mult_82_ab_23__42_,
         u5_mult_82_ab_23__43_, u5_mult_82_ab_23__44_, u5_mult_82_ab_23__45_,
         u5_mult_82_ab_23__46_, u5_mult_82_ab_23__47_, u5_mult_82_ab_23__48_,
         u5_mult_82_ab_23__49_, u5_mult_82_ab_23__50_, u5_mult_82_ab_23__51_,
         u5_mult_82_ab_23__52_, u5_mult_82_ab_24__0_, u5_mult_82_ab_24__1_,
         u5_mult_82_ab_24__2_, u5_mult_82_ab_24__3_, u5_mult_82_ab_24__4_,
         u5_mult_82_ab_24__5_, u5_mult_82_ab_24__6_, u5_mult_82_ab_24__7_,
         u5_mult_82_ab_24__8_, u5_mult_82_ab_24__9_, u5_mult_82_ab_24__10_,
         u5_mult_82_ab_24__11_, u5_mult_82_ab_24__12_, u5_mult_82_ab_24__13_,
         u5_mult_82_ab_24__14_, u5_mult_82_ab_24__15_, u5_mult_82_ab_24__16_,
         u5_mult_82_ab_24__17_, u5_mult_82_ab_24__18_, u5_mult_82_ab_24__19_,
         u5_mult_82_ab_24__20_, u5_mult_82_ab_24__21_, u5_mult_82_ab_24__22_,
         u5_mult_82_ab_24__23_, u5_mult_82_ab_24__24_, u5_mult_82_ab_24__25_,
         u5_mult_82_ab_24__26_, u5_mult_82_ab_24__27_, u5_mult_82_ab_24__28_,
         u5_mult_82_ab_24__29_, u5_mult_82_ab_24__30_, u5_mult_82_ab_24__31_,
         u5_mult_82_ab_24__32_, u5_mult_82_ab_24__33_, u5_mult_82_ab_24__34_,
         u5_mult_82_ab_24__35_, u5_mult_82_ab_24__36_, u5_mult_82_ab_24__37_,
         u5_mult_82_ab_24__38_, u5_mult_82_ab_24__39_, u5_mult_82_ab_24__40_,
         u5_mult_82_ab_24__41_, u5_mult_82_ab_24__42_, u5_mult_82_ab_24__43_,
         u5_mult_82_ab_24__44_, u5_mult_82_ab_24__45_, u5_mult_82_ab_24__46_,
         u5_mult_82_ab_24__47_, u5_mult_82_ab_24__48_, u5_mult_82_ab_24__49_,
         u5_mult_82_ab_24__50_, u5_mult_82_ab_24__51_, u5_mult_82_ab_24__52_,
         u5_mult_82_ab_25__0_, u5_mult_82_ab_25__1_, u5_mult_82_ab_25__2_,
         u5_mult_82_ab_25__3_, u5_mult_82_ab_25__4_, u5_mult_82_ab_25__5_,
         u5_mult_82_ab_25__6_, u5_mult_82_ab_25__7_, u5_mult_82_ab_25__8_,
         u5_mult_82_ab_25__9_, u5_mult_82_ab_25__10_, u5_mult_82_ab_25__11_,
         u5_mult_82_ab_25__12_, u5_mult_82_ab_25__13_, u5_mult_82_ab_25__14_,
         u5_mult_82_ab_25__15_, u5_mult_82_ab_25__16_, u5_mult_82_ab_25__17_,
         u5_mult_82_ab_25__18_, u5_mult_82_ab_25__19_, u5_mult_82_ab_25__20_,
         u5_mult_82_ab_25__21_, u5_mult_82_ab_25__23_, u5_mult_82_ab_25__24_,
         u5_mult_82_ab_25__25_, u5_mult_82_ab_25__26_, u5_mult_82_ab_25__27_,
         u5_mult_82_ab_25__28_, u5_mult_82_ab_25__29_, u5_mult_82_ab_25__30_,
         u5_mult_82_ab_25__31_, u5_mult_82_ab_25__32_, u5_mult_82_ab_25__33_,
         u5_mult_82_ab_25__34_, u5_mult_82_ab_25__35_, u5_mult_82_ab_25__36_,
         u5_mult_82_ab_25__37_, u5_mult_82_ab_25__38_, u5_mult_82_ab_25__39_,
         u5_mult_82_ab_25__40_, u5_mult_82_ab_25__41_, u5_mult_82_ab_25__42_,
         u5_mult_82_ab_25__43_, u5_mult_82_ab_25__44_, u5_mult_82_ab_25__45_,
         u5_mult_82_ab_25__46_, u5_mult_82_ab_25__47_, u5_mult_82_ab_25__48_,
         u5_mult_82_ab_25__49_, u5_mult_82_ab_25__50_, u5_mult_82_ab_25__51_,
         u5_mult_82_ab_25__52_, u5_mult_82_ab_26__0_, u5_mult_82_ab_26__1_,
         u5_mult_82_ab_26__2_, u5_mult_82_ab_26__3_, u5_mult_82_ab_26__4_,
         u5_mult_82_ab_26__5_, u5_mult_82_ab_26__6_, u5_mult_82_ab_26__7_,
         u5_mult_82_ab_26__8_, u5_mult_82_ab_26__9_, u5_mult_82_ab_26__10_,
         u5_mult_82_ab_26__11_, u5_mult_82_ab_26__12_, u5_mult_82_ab_26__13_,
         u5_mult_82_ab_26__14_, u5_mult_82_ab_26__15_, u5_mult_82_ab_26__16_,
         u5_mult_82_ab_26__17_, u5_mult_82_ab_26__18_, u5_mult_82_ab_26__19_,
         u5_mult_82_ab_26__20_, u5_mult_82_ab_26__21_, u5_mult_82_ab_26__22_,
         u5_mult_82_ab_26__23_, u5_mult_82_ab_26__24_, u5_mult_82_ab_26__25_,
         u5_mult_82_ab_26__26_, u5_mult_82_ab_26__27_, u5_mult_82_ab_26__28_,
         u5_mult_82_ab_26__29_, u5_mult_82_ab_26__30_, u5_mult_82_ab_26__31_,
         u5_mult_82_ab_26__32_, u5_mult_82_ab_26__33_, u5_mult_82_ab_26__34_,
         u5_mult_82_ab_26__35_, u5_mult_82_ab_26__36_, u5_mult_82_ab_26__37_,
         u5_mult_82_ab_26__38_, u5_mult_82_ab_26__39_, u5_mult_82_ab_26__40_,
         u5_mult_82_ab_26__41_, u5_mult_82_ab_26__42_, u5_mult_82_ab_26__43_,
         u5_mult_82_ab_26__44_, u5_mult_82_ab_26__45_, u5_mult_82_ab_26__46_,
         u5_mult_82_ab_26__47_, u5_mult_82_ab_26__48_, u5_mult_82_ab_26__49_,
         u5_mult_82_ab_26__50_, u5_mult_82_ab_26__51_, u5_mult_82_ab_26__52_,
         u5_mult_82_ab_27__0_, u5_mult_82_ab_27__1_, u5_mult_82_ab_27__2_,
         u5_mult_82_ab_27__3_, u5_mult_82_ab_27__4_, u5_mult_82_ab_27__5_,
         u5_mult_82_ab_27__6_, u5_mult_82_ab_27__7_, u5_mult_82_ab_27__8_,
         u5_mult_82_ab_27__9_, u5_mult_82_ab_27__10_, u5_mult_82_ab_27__11_,
         u5_mult_82_ab_27__12_, u5_mult_82_ab_27__13_, u5_mult_82_ab_27__14_,
         u5_mult_82_ab_27__15_, u5_mult_82_ab_27__16_, u5_mult_82_ab_27__17_,
         u5_mult_82_ab_27__18_, u5_mult_82_ab_27__19_, u5_mult_82_ab_27__20_,
         u5_mult_82_ab_27__21_, u5_mult_82_ab_27__22_, u5_mult_82_ab_27__23_,
         u5_mult_82_ab_27__24_, u5_mult_82_ab_27__25_, u5_mult_82_ab_27__26_,
         u5_mult_82_ab_27__27_, u5_mult_82_ab_27__28_, u5_mult_82_ab_27__29_,
         u5_mult_82_ab_27__30_, u5_mult_82_ab_27__31_, u5_mult_82_ab_27__32_,
         u5_mult_82_ab_27__33_, u5_mult_82_ab_27__34_, u5_mult_82_ab_27__35_,
         u5_mult_82_ab_27__36_, u5_mult_82_ab_27__37_, u5_mult_82_ab_27__38_,
         u5_mult_82_ab_27__39_, u5_mult_82_ab_27__40_, u5_mult_82_ab_27__41_,
         u5_mult_82_ab_27__42_, u5_mult_82_ab_27__43_, u5_mult_82_ab_27__44_,
         u5_mult_82_ab_27__45_, u5_mult_82_ab_27__46_, u5_mult_82_ab_27__47_,
         u5_mult_82_ab_27__48_, u5_mult_82_ab_27__49_, u5_mult_82_ab_27__50_,
         u5_mult_82_ab_27__51_, u5_mult_82_ab_27__52_, u5_mult_82_ab_28__0_,
         u5_mult_82_ab_28__1_, u5_mult_82_ab_28__2_, u5_mult_82_ab_28__3_,
         u5_mult_82_ab_28__4_, u5_mult_82_ab_28__5_, u5_mult_82_ab_28__6_,
         u5_mult_82_ab_28__7_, u5_mult_82_ab_28__8_, u5_mult_82_ab_28__9_,
         u5_mult_82_ab_28__10_, u5_mult_82_ab_28__11_, u5_mult_82_ab_28__12_,
         u5_mult_82_ab_28__13_, u5_mult_82_ab_28__14_, u5_mult_82_ab_28__15_,
         u5_mult_82_ab_28__16_, u5_mult_82_ab_28__17_, u5_mult_82_ab_28__18_,
         u5_mult_82_ab_28__19_, u5_mult_82_ab_28__20_, u5_mult_82_ab_28__21_,
         u5_mult_82_ab_28__22_, u5_mult_82_ab_28__23_, u5_mult_82_ab_28__24_,
         u5_mult_82_ab_28__25_, u5_mult_82_ab_28__26_, u5_mult_82_ab_28__27_,
         u5_mult_82_ab_28__28_, u5_mult_82_ab_28__29_, u5_mult_82_ab_28__30_,
         u5_mult_82_ab_28__31_, u5_mult_82_ab_28__32_, u5_mult_82_ab_28__33_,
         u5_mult_82_ab_28__34_, u5_mult_82_ab_28__35_, u5_mult_82_ab_28__36_,
         u5_mult_82_ab_28__37_, u5_mult_82_ab_28__38_, u5_mult_82_ab_28__39_,
         u5_mult_82_ab_28__40_, u5_mult_82_ab_28__41_, u5_mult_82_ab_28__42_,
         u5_mult_82_ab_28__43_, u5_mult_82_ab_28__44_, u5_mult_82_ab_28__45_,
         u5_mult_82_ab_28__46_, u5_mult_82_ab_28__47_, u5_mult_82_ab_28__48_,
         u5_mult_82_ab_28__49_, u5_mult_82_ab_28__50_, u5_mult_82_ab_28__51_,
         u5_mult_82_ab_28__52_, u5_mult_82_ab_29__0_, u5_mult_82_ab_29__1_,
         u5_mult_82_ab_29__2_, u5_mult_82_ab_29__3_, u5_mult_82_ab_29__4_,
         u5_mult_82_ab_29__5_, u5_mult_82_ab_29__6_, u5_mult_82_ab_29__7_,
         u5_mult_82_ab_29__8_, u5_mult_82_ab_29__9_, u5_mult_82_ab_29__10_,
         u5_mult_82_ab_29__11_, u5_mult_82_ab_29__12_, u5_mult_82_ab_29__13_,
         u5_mult_82_ab_29__14_, u5_mult_82_ab_29__15_, u5_mult_82_ab_29__16_,
         u5_mult_82_ab_29__17_, u5_mult_82_ab_29__18_, u5_mult_82_ab_29__19_,
         u5_mult_82_ab_29__20_, u5_mult_82_ab_29__21_, u5_mult_82_ab_29__22_,
         u5_mult_82_ab_29__23_, u5_mult_82_ab_29__24_, u5_mult_82_ab_29__25_,
         u5_mult_82_ab_29__26_, u5_mult_82_ab_29__27_, u5_mult_82_ab_29__28_,
         u5_mult_82_ab_29__29_, u5_mult_82_ab_29__30_, u5_mult_82_ab_29__31_,
         u5_mult_82_ab_29__32_, u5_mult_82_ab_29__33_, u5_mult_82_ab_29__34_,
         u5_mult_82_ab_29__35_, u5_mult_82_ab_29__36_, u5_mult_82_ab_29__37_,
         u5_mult_82_ab_29__38_, u5_mult_82_ab_29__39_, u5_mult_82_ab_29__40_,
         u5_mult_82_ab_29__41_, u5_mult_82_ab_29__42_, u5_mult_82_ab_29__43_,
         u5_mult_82_ab_29__44_, u5_mult_82_ab_29__45_, u5_mult_82_ab_29__46_,
         u5_mult_82_ab_29__47_, u5_mult_82_ab_29__48_, u5_mult_82_ab_29__49_,
         u5_mult_82_ab_29__50_, u5_mult_82_ab_29__51_, u5_mult_82_ab_29__52_,
         u5_mult_82_ab_30__0_, u5_mult_82_ab_30__1_, u5_mult_82_ab_30__2_,
         u5_mult_82_ab_30__3_, u5_mult_82_ab_30__4_, u5_mult_82_ab_30__5_,
         u5_mult_82_ab_30__6_, u5_mult_82_ab_30__7_, u5_mult_82_ab_30__8_,
         u5_mult_82_ab_30__9_, u5_mult_82_ab_30__10_, u5_mult_82_ab_30__11_,
         u5_mult_82_ab_30__12_, u5_mult_82_ab_30__13_, u5_mult_82_ab_30__14_,
         u5_mult_82_ab_30__15_, u5_mult_82_ab_30__16_, u5_mult_82_ab_30__17_,
         u5_mult_82_ab_30__18_, u5_mult_82_ab_30__19_, u5_mult_82_ab_30__20_,
         u5_mult_82_ab_30__21_, u5_mult_82_ab_30__22_, u5_mult_82_ab_30__23_,
         u5_mult_82_ab_30__24_, u5_mult_82_ab_30__25_, u5_mult_82_ab_30__26_,
         u5_mult_82_ab_30__27_, u5_mult_82_ab_30__28_, u5_mult_82_ab_30__29_,
         u5_mult_82_ab_30__30_, u5_mult_82_ab_30__31_, u5_mult_82_ab_30__32_,
         u5_mult_82_ab_30__33_, u5_mult_82_ab_30__34_, u5_mult_82_ab_30__35_,
         u5_mult_82_ab_30__36_, u5_mult_82_ab_30__37_, u5_mult_82_ab_30__38_,
         u5_mult_82_ab_30__39_, u5_mult_82_ab_30__40_, u5_mult_82_ab_30__41_,
         u5_mult_82_ab_30__42_, u5_mult_82_ab_30__43_, u5_mult_82_ab_30__44_,
         u5_mult_82_ab_30__45_, u5_mult_82_ab_30__46_, u5_mult_82_ab_30__47_,
         u5_mult_82_ab_30__48_, u5_mult_82_ab_30__49_, u5_mult_82_ab_30__50_,
         u5_mult_82_ab_30__51_, u5_mult_82_ab_30__52_, u5_mult_82_ab_31__0_,
         u5_mult_82_ab_31__1_, u5_mult_82_ab_31__2_, u5_mult_82_ab_31__3_,
         u5_mult_82_ab_31__4_, u5_mult_82_ab_31__5_, u5_mult_82_ab_31__6_,
         u5_mult_82_ab_31__7_, u5_mult_82_ab_31__8_, u5_mult_82_ab_31__9_,
         u5_mult_82_ab_31__10_, u5_mult_82_ab_31__11_, u5_mult_82_ab_31__12_,
         u5_mult_82_ab_31__13_, u5_mult_82_ab_31__14_, u5_mult_82_ab_31__15_,
         u5_mult_82_ab_31__16_, u5_mult_82_ab_31__17_, u5_mult_82_ab_31__18_,
         u5_mult_82_ab_31__19_, u5_mult_82_ab_31__20_, u5_mult_82_ab_31__21_,
         u5_mult_82_ab_31__22_, u5_mult_82_ab_31__23_, u5_mult_82_ab_31__24_,
         u5_mult_82_ab_31__25_, u5_mult_82_ab_31__26_, u5_mult_82_ab_31__27_,
         u5_mult_82_ab_31__28_, u5_mult_82_ab_31__29_, u5_mult_82_ab_31__30_,
         u5_mult_82_ab_31__31_, u5_mult_82_ab_31__32_, u5_mult_82_ab_31__33_,
         u5_mult_82_ab_31__34_, u5_mult_82_ab_31__35_, u5_mult_82_ab_31__36_,
         u5_mult_82_ab_31__37_, u5_mult_82_ab_31__38_, u5_mult_82_ab_31__39_,
         u5_mult_82_ab_31__40_, u5_mult_82_ab_31__41_, u5_mult_82_ab_31__42_,
         u5_mult_82_ab_31__43_, u5_mult_82_ab_31__44_, u5_mult_82_ab_31__45_,
         u5_mult_82_ab_31__46_, u5_mult_82_ab_31__47_, u5_mult_82_ab_31__48_,
         u5_mult_82_ab_31__49_, u5_mult_82_ab_31__50_, u5_mult_82_ab_31__51_,
         u5_mult_82_ab_31__52_, u5_mult_82_ab_32__0_, u5_mult_82_ab_32__1_,
         u5_mult_82_ab_32__2_, u5_mult_82_ab_32__3_, u5_mult_82_ab_32__4_,
         u5_mult_82_ab_32__5_, u5_mult_82_ab_32__6_, u5_mult_82_ab_32__7_,
         u5_mult_82_ab_32__8_, u5_mult_82_ab_32__9_, u5_mult_82_ab_32__10_,
         u5_mult_82_ab_32__11_, u5_mult_82_ab_32__12_, u5_mult_82_ab_32__13_,
         u5_mult_82_ab_32__14_, u5_mult_82_ab_32__15_, u5_mult_82_ab_32__16_,
         u5_mult_82_ab_32__17_, u5_mult_82_ab_32__18_, u5_mult_82_ab_32__19_,
         u5_mult_82_ab_32__20_, u5_mult_82_ab_32__21_, u5_mult_82_ab_32__22_,
         u5_mult_82_ab_32__23_, u5_mult_82_ab_32__24_, u5_mult_82_ab_32__25_,
         u5_mult_82_ab_32__26_, u5_mult_82_ab_32__27_, u5_mult_82_ab_32__28_,
         u5_mult_82_ab_32__29_, u5_mult_82_ab_32__30_, u5_mult_82_ab_32__31_,
         u5_mult_82_ab_32__32_, u5_mult_82_ab_32__33_, u5_mult_82_ab_32__34_,
         u5_mult_82_ab_32__35_, u5_mult_82_ab_32__36_, u5_mult_82_ab_32__37_,
         u5_mult_82_ab_32__38_, u5_mult_82_ab_32__39_, u5_mult_82_ab_32__40_,
         u5_mult_82_ab_32__41_, u5_mult_82_ab_32__42_, u5_mult_82_ab_32__43_,
         u5_mult_82_ab_32__44_, u5_mult_82_ab_32__45_, u5_mult_82_ab_32__46_,
         u5_mult_82_ab_32__47_, u5_mult_82_ab_32__48_, u5_mult_82_ab_32__49_,
         u5_mult_82_ab_32__50_, u5_mult_82_ab_32__51_, u5_mult_82_ab_32__52_,
         u5_mult_82_ab_33__0_, u5_mult_82_ab_33__1_, u5_mult_82_ab_33__2_,
         u5_mult_82_ab_33__3_, u5_mult_82_ab_33__4_, u5_mult_82_ab_33__5_,
         u5_mult_82_ab_33__6_, u5_mult_82_ab_33__7_, u5_mult_82_ab_33__8_,
         u5_mult_82_ab_33__9_, u5_mult_82_ab_33__10_, u5_mult_82_ab_33__11_,
         u5_mult_82_ab_33__12_, u5_mult_82_ab_33__13_, u5_mult_82_ab_33__14_,
         u5_mult_82_ab_33__15_, u5_mult_82_ab_33__16_, u5_mult_82_ab_33__17_,
         u5_mult_82_ab_33__18_, u5_mult_82_ab_33__19_, u5_mult_82_ab_33__20_,
         u5_mult_82_ab_33__21_, u5_mult_82_ab_33__22_, u5_mult_82_ab_33__23_,
         u5_mult_82_ab_33__24_, u5_mult_82_ab_33__25_, u5_mult_82_ab_33__26_,
         u5_mult_82_ab_33__27_, u5_mult_82_ab_33__28_, u5_mult_82_ab_33__29_,
         u5_mult_82_ab_33__30_, u5_mult_82_ab_33__31_, u5_mult_82_ab_33__32_,
         u5_mult_82_ab_33__33_, u5_mult_82_ab_33__34_, u5_mult_82_ab_33__35_,
         u5_mult_82_ab_33__36_, u5_mult_82_ab_33__37_, u5_mult_82_ab_33__38_,
         u5_mult_82_ab_33__39_, u5_mult_82_ab_33__40_, u5_mult_82_ab_33__41_,
         u5_mult_82_ab_33__42_, u5_mult_82_ab_33__43_, u5_mult_82_ab_33__44_,
         u5_mult_82_ab_33__45_, u5_mult_82_ab_33__46_, u5_mult_82_ab_33__47_,
         u5_mult_82_ab_33__48_, u5_mult_82_ab_33__49_, u5_mult_82_ab_33__50_,
         u5_mult_82_ab_33__51_, u5_mult_82_ab_33__52_, u5_mult_82_ab_34__0_,
         u5_mult_82_ab_34__1_, u5_mult_82_ab_34__2_, u5_mult_82_ab_34__3_,
         u5_mult_82_ab_34__4_, u5_mult_82_ab_34__5_, u5_mult_82_ab_34__6_,
         u5_mult_82_ab_34__7_, u5_mult_82_ab_34__8_, u5_mult_82_ab_34__9_,
         u5_mult_82_ab_34__10_, u5_mult_82_ab_34__11_, u5_mult_82_ab_34__12_,
         u5_mult_82_ab_34__13_, u5_mult_82_ab_34__14_, u5_mult_82_ab_34__15_,
         u5_mult_82_ab_34__17_, u5_mult_82_ab_34__18_, u5_mult_82_ab_34__19_,
         u5_mult_82_ab_34__20_, u5_mult_82_ab_34__21_, u5_mult_82_ab_34__22_,
         u5_mult_82_ab_34__23_, u5_mult_82_ab_34__24_, u5_mult_82_ab_34__25_,
         u5_mult_82_ab_34__26_, u5_mult_82_ab_34__27_, u5_mult_82_ab_34__28_,
         u5_mult_82_ab_34__29_, u5_mult_82_ab_34__30_, u5_mult_82_ab_34__31_,
         u5_mult_82_ab_34__32_, u5_mult_82_ab_34__33_, u5_mult_82_ab_34__34_,
         u5_mult_82_ab_34__35_, u5_mult_82_ab_34__36_, u5_mult_82_ab_34__37_,
         u5_mult_82_ab_34__38_, u5_mult_82_ab_34__39_, u5_mult_82_ab_34__40_,
         u5_mult_82_ab_34__41_, u5_mult_82_ab_34__42_, u5_mult_82_ab_34__43_,
         u5_mult_82_ab_34__44_, u5_mult_82_ab_34__45_, u5_mult_82_ab_34__46_,
         u5_mult_82_ab_34__47_, u5_mult_82_ab_34__48_, u5_mult_82_ab_34__49_,
         u5_mult_82_ab_34__50_, u5_mult_82_ab_34__51_, u5_mult_82_ab_34__52_,
         u5_mult_82_ab_35__0_, u5_mult_82_ab_35__1_, u5_mult_82_ab_35__2_,
         u5_mult_82_ab_35__3_, u5_mult_82_ab_35__4_, u5_mult_82_ab_35__5_,
         u5_mult_82_ab_35__6_, u5_mult_82_ab_35__7_, u5_mult_82_ab_35__8_,
         u5_mult_82_ab_35__9_, u5_mult_82_ab_35__10_, u5_mult_82_ab_35__11_,
         u5_mult_82_ab_35__12_, u5_mult_82_ab_35__13_, u5_mult_82_ab_35__14_,
         u5_mult_82_ab_35__15_, u5_mult_82_ab_35__16_, u5_mult_82_ab_35__17_,
         u5_mult_82_ab_35__18_, u5_mult_82_ab_35__19_, u5_mult_82_ab_35__20_,
         u5_mult_82_ab_35__21_, u5_mult_82_ab_35__22_, u5_mult_82_ab_35__23_,
         u5_mult_82_ab_35__24_, u5_mult_82_ab_35__25_, u5_mult_82_ab_35__26_,
         u5_mult_82_ab_35__27_, u5_mult_82_ab_35__28_, u5_mult_82_ab_35__29_,
         u5_mult_82_ab_35__30_, u5_mult_82_ab_35__31_, u5_mult_82_ab_35__32_,
         u5_mult_82_ab_35__33_, u5_mult_82_ab_35__34_, u5_mult_82_ab_35__35_,
         u5_mult_82_ab_35__36_, u5_mult_82_ab_35__37_, u5_mult_82_ab_35__38_,
         u5_mult_82_ab_35__39_, u5_mult_82_ab_35__40_, u5_mult_82_ab_35__41_,
         u5_mult_82_ab_35__42_, u5_mult_82_ab_35__43_, u5_mult_82_ab_35__44_,
         u5_mult_82_ab_35__45_, u5_mult_82_ab_35__46_, u5_mult_82_ab_35__47_,
         u5_mult_82_ab_35__48_, u5_mult_82_ab_35__49_, u5_mult_82_ab_35__50_,
         u5_mult_82_ab_35__51_, u5_mult_82_ab_35__52_, u5_mult_82_ab_36__0_,
         u5_mult_82_ab_36__1_, u5_mult_82_ab_36__2_, u5_mult_82_ab_36__3_,
         u5_mult_82_ab_36__4_, u5_mult_82_ab_36__5_, u5_mult_82_ab_36__6_,
         u5_mult_82_ab_36__7_, u5_mult_82_ab_36__8_, u5_mult_82_ab_36__9_,
         u5_mult_82_ab_36__10_, u5_mult_82_ab_36__11_, u5_mult_82_ab_36__12_,
         u5_mult_82_ab_36__13_, u5_mult_82_ab_36__14_, u5_mult_82_ab_36__15_,
         u5_mult_82_ab_36__16_, u5_mult_82_ab_36__17_, u5_mult_82_ab_36__18_,
         u5_mult_82_ab_36__19_, u5_mult_82_ab_36__20_, u5_mult_82_ab_36__21_,
         u5_mult_82_ab_36__22_, u5_mult_82_ab_36__23_, u5_mult_82_ab_36__24_,
         u5_mult_82_ab_36__25_, u5_mult_82_ab_36__26_, u5_mult_82_ab_36__27_,
         u5_mult_82_ab_36__28_, u5_mult_82_ab_36__29_, u5_mult_82_ab_36__30_,
         u5_mult_82_ab_36__31_, u5_mult_82_ab_36__32_, u5_mult_82_ab_36__33_,
         u5_mult_82_ab_36__34_, u5_mult_82_ab_36__35_, u5_mult_82_ab_36__36_,
         u5_mult_82_ab_36__37_, u5_mult_82_ab_36__38_, u5_mult_82_ab_36__39_,
         u5_mult_82_ab_36__40_, u5_mult_82_ab_36__41_, u5_mult_82_ab_36__42_,
         u5_mult_82_ab_36__43_, u5_mult_82_ab_36__44_, u5_mult_82_ab_36__45_,
         u5_mult_82_ab_36__46_, u5_mult_82_ab_36__47_, u5_mult_82_ab_36__48_,
         u5_mult_82_ab_36__49_, u5_mult_82_ab_36__50_, u5_mult_82_ab_36__51_,
         u5_mult_82_ab_36__52_, u5_mult_82_ab_37__0_, u5_mult_82_ab_37__1_,
         u5_mult_82_ab_37__2_, u5_mult_82_ab_37__3_, u5_mult_82_ab_37__4_,
         u5_mult_82_ab_37__5_, u5_mult_82_ab_37__6_, u5_mult_82_ab_37__7_,
         u5_mult_82_ab_37__8_, u5_mult_82_ab_37__9_, u5_mult_82_ab_37__10_,
         u5_mult_82_ab_37__11_, u5_mult_82_ab_37__12_, u5_mult_82_ab_37__13_,
         u5_mult_82_ab_37__14_, u5_mult_82_ab_37__15_, u5_mult_82_ab_37__16_,
         u5_mult_82_ab_37__17_, u5_mult_82_ab_37__18_, u5_mult_82_ab_37__19_,
         u5_mult_82_ab_37__20_, u5_mult_82_ab_37__21_, u5_mult_82_ab_37__22_,
         u5_mult_82_ab_37__23_, u5_mult_82_ab_37__24_, u5_mult_82_ab_37__25_,
         u5_mult_82_ab_37__26_, u5_mult_82_ab_37__27_, u5_mult_82_ab_37__28_,
         u5_mult_82_ab_37__29_, u5_mult_82_ab_37__30_, u5_mult_82_ab_37__31_,
         u5_mult_82_ab_37__32_, u5_mult_82_ab_37__33_, u5_mult_82_ab_37__34_,
         u5_mult_82_ab_37__35_, u5_mult_82_ab_37__36_, u5_mult_82_ab_37__37_,
         u5_mult_82_ab_37__38_, u5_mult_82_ab_37__39_, u5_mult_82_ab_37__40_,
         u5_mult_82_ab_37__41_, u5_mult_82_ab_37__42_, u5_mult_82_ab_37__43_,
         u5_mult_82_ab_37__44_, u5_mult_82_ab_37__45_, u5_mult_82_ab_37__46_,
         u5_mult_82_ab_37__47_, u5_mult_82_ab_37__48_, u5_mult_82_ab_37__49_,
         u5_mult_82_ab_37__50_, u5_mult_82_ab_37__51_, u5_mult_82_ab_37__52_,
         u5_mult_82_ab_38__0_, u5_mult_82_ab_38__1_, u5_mult_82_ab_38__2_,
         u5_mult_82_ab_38__3_, u5_mult_82_ab_38__4_, u5_mult_82_ab_38__5_,
         u5_mult_82_ab_38__6_, u5_mult_82_ab_38__7_, u5_mult_82_ab_38__8_,
         u5_mult_82_ab_38__9_, u5_mult_82_ab_38__10_, u5_mult_82_ab_38__11_,
         u5_mult_82_ab_38__12_, u5_mult_82_ab_38__13_, u5_mult_82_ab_38__15_,
         u5_mult_82_ab_38__16_, u5_mult_82_ab_38__17_, u5_mult_82_ab_38__18_,
         u5_mult_82_ab_38__19_, u5_mult_82_ab_38__20_, u5_mult_82_ab_38__21_,
         u5_mult_82_ab_38__22_, u5_mult_82_ab_38__23_, u5_mult_82_ab_38__24_,
         u5_mult_82_ab_38__25_, u5_mult_82_ab_38__26_, u5_mult_82_ab_38__27_,
         u5_mult_82_ab_38__28_, u5_mult_82_ab_38__29_, u5_mult_82_ab_38__30_,
         u5_mult_82_ab_38__31_, u5_mult_82_ab_38__32_, u5_mult_82_ab_38__33_,
         u5_mult_82_ab_38__34_, u5_mult_82_ab_38__35_, u5_mult_82_ab_38__36_,
         u5_mult_82_ab_38__37_, u5_mult_82_ab_38__38_, u5_mult_82_ab_38__39_,
         u5_mult_82_ab_38__40_, u5_mult_82_ab_38__41_, u5_mult_82_ab_38__42_,
         u5_mult_82_ab_38__43_, u5_mult_82_ab_38__44_, u5_mult_82_ab_38__45_,
         u5_mult_82_ab_38__46_, u5_mult_82_ab_38__47_, u5_mult_82_ab_38__48_,
         u5_mult_82_ab_38__49_, u5_mult_82_ab_38__50_, u5_mult_82_ab_38__51_,
         u5_mult_82_ab_38__52_, u5_mult_82_ab_39__0_, u5_mult_82_ab_39__1_,
         u5_mult_82_ab_39__2_, u5_mult_82_ab_39__3_, u5_mult_82_ab_39__4_,
         u5_mult_82_ab_39__5_, u5_mult_82_ab_39__6_, u5_mult_82_ab_39__7_,
         u5_mult_82_ab_39__8_, u5_mult_82_ab_39__9_, u5_mult_82_ab_39__10_,
         u5_mult_82_ab_39__11_, u5_mult_82_ab_39__12_, u5_mult_82_ab_39__13_,
         u5_mult_82_ab_39__14_, u5_mult_82_ab_39__15_, u5_mult_82_ab_39__16_,
         u5_mult_82_ab_39__17_, u5_mult_82_ab_39__18_, u5_mult_82_ab_39__19_,
         u5_mult_82_ab_39__20_, u5_mult_82_ab_39__21_, u5_mult_82_ab_39__22_,
         u5_mult_82_ab_39__23_, u5_mult_82_ab_39__24_, u5_mult_82_ab_39__25_,
         u5_mult_82_ab_39__26_, u5_mult_82_ab_39__27_, u5_mult_82_ab_39__28_,
         u5_mult_82_ab_39__29_, u5_mult_82_ab_39__30_, u5_mult_82_ab_39__31_,
         u5_mult_82_ab_39__32_, u5_mult_82_ab_39__33_, u5_mult_82_ab_39__34_,
         u5_mult_82_ab_39__35_, u5_mult_82_ab_39__36_, u5_mult_82_ab_39__37_,
         u5_mult_82_ab_39__38_, u5_mult_82_ab_39__39_, u5_mult_82_ab_39__40_,
         u5_mult_82_ab_39__41_, u5_mult_82_ab_39__42_, u5_mult_82_ab_39__43_,
         u5_mult_82_ab_39__44_, u5_mult_82_ab_39__45_, u5_mult_82_ab_39__46_,
         u5_mult_82_ab_39__47_, u5_mult_82_ab_39__48_, u5_mult_82_ab_39__49_,
         u5_mult_82_ab_39__50_, u5_mult_82_ab_39__51_, u5_mult_82_ab_39__52_,
         u5_mult_82_ab_40__0_, u5_mult_82_ab_40__1_, u5_mult_82_ab_40__2_,
         u5_mult_82_ab_40__3_, u5_mult_82_ab_40__4_, u5_mult_82_ab_40__5_,
         u5_mult_82_ab_40__6_, u5_mult_82_ab_40__7_, u5_mult_82_ab_40__8_,
         u5_mult_82_ab_40__9_, u5_mult_82_ab_40__10_, u5_mult_82_ab_40__11_,
         u5_mult_82_ab_40__13_, u5_mult_82_ab_40__14_, u5_mult_82_ab_40__15_,
         u5_mult_82_ab_40__16_, u5_mult_82_ab_40__17_, u5_mult_82_ab_40__18_,
         u5_mult_82_ab_40__19_, u5_mult_82_ab_40__20_, u5_mult_82_ab_40__21_,
         u5_mult_82_ab_40__22_, u5_mult_82_ab_40__23_, u5_mult_82_ab_40__24_,
         u5_mult_82_ab_40__25_, u5_mult_82_ab_40__26_, u5_mult_82_ab_40__27_,
         u5_mult_82_ab_40__28_, u5_mult_82_ab_40__29_, u5_mult_82_ab_40__30_,
         u5_mult_82_ab_40__31_, u5_mult_82_ab_40__32_, u5_mult_82_ab_40__33_,
         u5_mult_82_ab_40__34_, u5_mult_82_ab_40__35_, u5_mult_82_ab_40__36_,
         u5_mult_82_ab_40__37_, u5_mult_82_ab_40__38_, u5_mult_82_ab_40__39_,
         u5_mult_82_ab_40__40_, u5_mult_82_ab_40__41_, u5_mult_82_ab_40__42_,
         u5_mult_82_ab_40__43_, u5_mult_82_ab_40__44_, u5_mult_82_ab_40__45_,
         u5_mult_82_ab_40__46_, u5_mult_82_ab_40__47_, u5_mult_82_ab_40__48_,
         u5_mult_82_ab_40__49_, u5_mult_82_ab_40__50_, u5_mult_82_ab_40__51_,
         u5_mult_82_ab_40__52_, u5_mult_82_ab_41__0_, u5_mult_82_ab_41__1_,
         u5_mult_82_ab_41__2_, u5_mult_82_ab_41__3_, u5_mult_82_ab_41__4_,
         u5_mult_82_ab_41__5_, u5_mult_82_ab_41__6_, u5_mult_82_ab_41__7_,
         u5_mult_82_ab_41__8_, u5_mult_82_ab_41__9_, u5_mult_82_ab_41__10_,
         u5_mult_82_ab_41__11_, u5_mult_82_ab_41__14_, u5_mult_82_ab_41__15_,
         u5_mult_82_ab_41__16_, u5_mult_82_ab_41__17_, u5_mult_82_ab_41__18_,
         u5_mult_82_ab_41__19_, u5_mult_82_ab_41__20_, u5_mult_82_ab_41__21_,
         u5_mult_82_ab_41__22_, u5_mult_82_ab_41__23_, u5_mult_82_ab_41__24_,
         u5_mult_82_ab_41__25_, u5_mult_82_ab_41__26_, u5_mult_82_ab_41__27_,
         u5_mult_82_ab_41__28_, u5_mult_82_ab_41__29_, u5_mult_82_ab_41__30_,
         u5_mult_82_ab_41__31_, u5_mult_82_ab_41__32_, u5_mult_82_ab_41__33_,
         u5_mult_82_ab_41__34_, u5_mult_82_ab_41__35_, u5_mult_82_ab_41__36_,
         u5_mult_82_ab_41__37_, u5_mult_82_ab_41__38_, u5_mult_82_ab_41__39_,
         u5_mult_82_ab_41__40_, u5_mult_82_ab_41__41_, u5_mult_82_ab_41__42_,
         u5_mult_82_ab_41__43_, u5_mult_82_ab_41__44_, u5_mult_82_ab_41__45_,
         u5_mult_82_ab_41__46_, u5_mult_82_ab_41__47_, u5_mult_82_ab_41__48_,
         u5_mult_82_ab_41__49_, u5_mult_82_ab_41__50_, u5_mult_82_ab_41__51_,
         u5_mult_82_ab_41__52_, u5_mult_82_ab_42__0_, u5_mult_82_ab_42__1_,
         u5_mult_82_ab_42__2_, u5_mult_82_ab_42__3_, u5_mult_82_ab_42__4_,
         u5_mult_82_ab_42__5_, u5_mult_82_ab_42__6_, u5_mult_82_ab_42__7_,
         u5_mult_82_ab_42__8_, u5_mult_82_ab_42__9_, u5_mult_82_ab_42__10_,
         u5_mult_82_ab_42__12_, u5_mult_82_ab_42__13_, u5_mult_82_ab_42__14_,
         u5_mult_82_ab_42__15_, u5_mult_82_ab_42__16_, u5_mult_82_ab_42__17_,
         u5_mult_82_ab_42__18_, u5_mult_82_ab_42__19_, u5_mult_82_ab_42__20_,
         u5_mult_82_ab_42__21_, u5_mult_82_ab_42__22_, u5_mult_82_ab_42__23_,
         u5_mult_82_ab_42__24_, u5_mult_82_ab_42__25_, u5_mult_82_ab_42__26_,
         u5_mult_82_ab_42__27_, u5_mult_82_ab_42__28_, u5_mult_82_ab_42__29_,
         u5_mult_82_ab_42__30_, u5_mult_82_ab_42__31_, u5_mult_82_ab_42__32_,
         u5_mult_82_ab_42__33_, u5_mult_82_ab_42__34_, u5_mult_82_ab_42__35_,
         u5_mult_82_ab_42__36_, u5_mult_82_ab_42__37_, u5_mult_82_ab_42__38_,
         u5_mult_82_ab_42__39_, u5_mult_82_ab_42__40_, u5_mult_82_ab_42__41_,
         u5_mult_82_ab_42__42_, u5_mult_82_ab_42__43_, u5_mult_82_ab_42__44_,
         u5_mult_82_ab_42__45_, u5_mult_82_ab_42__46_, u5_mult_82_ab_42__47_,
         u5_mult_82_ab_42__48_, u5_mult_82_ab_42__49_, u5_mult_82_ab_42__50_,
         u5_mult_82_ab_42__51_, u5_mult_82_ab_42__52_, u5_mult_82_ab_43__0_,
         u5_mult_82_ab_43__1_, u5_mult_82_ab_43__2_, u5_mult_82_ab_43__3_,
         u5_mult_82_ab_43__4_, u5_mult_82_ab_43__5_, u5_mult_82_ab_43__6_,
         u5_mult_82_ab_43__7_, u5_mult_82_ab_43__8_, u5_mult_82_ab_43__9_,
         u5_mult_82_ab_43__11_, u5_mult_82_ab_43__12_, u5_mult_82_ab_43__13_,
         u5_mult_82_ab_43__14_, u5_mult_82_ab_43__15_, u5_mult_82_ab_43__16_,
         u5_mult_82_ab_43__17_, u5_mult_82_ab_43__18_, u5_mult_82_ab_43__19_,
         u5_mult_82_ab_43__20_, u5_mult_82_ab_43__21_, u5_mult_82_ab_43__22_,
         u5_mult_82_ab_43__23_, u5_mult_82_ab_43__24_, u5_mult_82_ab_43__25_,
         u5_mult_82_ab_43__26_, u5_mult_82_ab_43__27_, u5_mult_82_ab_43__28_,
         u5_mult_82_ab_43__29_, u5_mult_82_ab_43__30_, u5_mult_82_ab_43__31_,
         u5_mult_82_ab_43__32_, u5_mult_82_ab_43__33_, u5_mult_82_ab_43__34_,
         u5_mult_82_ab_43__35_, u5_mult_82_ab_43__36_, u5_mult_82_ab_43__37_,
         u5_mult_82_ab_43__38_, u5_mult_82_ab_43__39_, u5_mult_82_ab_43__40_,
         u5_mult_82_ab_43__41_, u5_mult_82_ab_43__42_, u5_mult_82_ab_43__43_,
         u5_mult_82_ab_43__44_, u5_mult_82_ab_43__45_, u5_mult_82_ab_43__46_,
         u5_mult_82_ab_43__47_, u5_mult_82_ab_43__48_, u5_mult_82_ab_43__49_,
         u5_mult_82_ab_43__50_, u5_mult_82_ab_43__51_, u5_mult_82_ab_43__52_,
         u5_mult_82_ab_44__0_, u5_mult_82_ab_44__1_, u5_mult_82_ab_44__2_,
         u5_mult_82_ab_44__3_, u5_mult_82_ab_44__4_, u5_mult_82_ab_44__5_,
         u5_mult_82_ab_44__6_, u5_mult_82_ab_44__7_, u5_mult_82_ab_44__8_,
         u5_mult_82_ab_44__9_, u5_mult_82_ab_44__10_, u5_mult_82_ab_44__11_,
         u5_mult_82_ab_44__12_, u5_mult_82_ab_44__13_, u5_mult_82_ab_44__14_,
         u5_mult_82_ab_44__15_, u5_mult_82_ab_44__16_, u5_mult_82_ab_44__17_,
         u5_mult_82_ab_44__18_, u5_mult_82_ab_44__19_, u5_mult_82_ab_44__20_,
         u5_mult_82_ab_44__21_, u5_mult_82_ab_44__22_, u5_mult_82_ab_44__23_,
         u5_mult_82_ab_44__24_, u5_mult_82_ab_44__25_, u5_mult_82_ab_44__26_,
         u5_mult_82_ab_44__27_, u5_mult_82_ab_44__28_, u5_mult_82_ab_44__29_,
         u5_mult_82_ab_44__30_, u5_mult_82_ab_44__31_, u5_mult_82_ab_44__32_,
         u5_mult_82_ab_44__33_, u5_mult_82_ab_44__34_, u5_mult_82_ab_44__35_,
         u5_mult_82_ab_44__36_, u5_mult_82_ab_44__37_, u5_mult_82_ab_44__38_,
         u5_mult_82_ab_44__39_, u5_mult_82_ab_44__40_, u5_mult_82_ab_44__41_,
         u5_mult_82_ab_44__42_, u5_mult_82_ab_44__43_, u5_mult_82_ab_44__44_,
         u5_mult_82_ab_44__45_, u5_mult_82_ab_44__46_, u5_mult_82_ab_44__47_,
         u5_mult_82_ab_44__48_, u5_mult_82_ab_44__49_, u5_mult_82_ab_44__50_,
         u5_mult_82_ab_44__51_, u5_mult_82_ab_44__52_, u5_mult_82_ab_45__0_,
         u5_mult_82_ab_45__1_, u5_mult_82_ab_45__2_, u5_mult_82_ab_45__3_,
         u5_mult_82_ab_45__4_, u5_mult_82_ab_45__5_, u5_mult_82_ab_45__6_,
         u5_mult_82_ab_45__7_, u5_mult_82_ab_45__8_, u5_mult_82_ab_45__10_,
         u5_mult_82_ab_45__11_, u5_mult_82_ab_45__12_, u5_mult_82_ab_45__13_,
         u5_mult_82_ab_45__14_, u5_mult_82_ab_45__15_, u5_mult_82_ab_45__16_,
         u5_mult_82_ab_45__17_, u5_mult_82_ab_45__18_, u5_mult_82_ab_45__19_,
         u5_mult_82_ab_45__20_, u5_mult_82_ab_45__21_, u5_mult_82_ab_45__22_,
         u5_mult_82_ab_45__23_, u5_mult_82_ab_45__24_, u5_mult_82_ab_45__25_,
         u5_mult_82_ab_45__26_, u5_mult_82_ab_45__27_, u5_mult_82_ab_45__28_,
         u5_mult_82_ab_45__29_, u5_mult_82_ab_45__30_, u5_mult_82_ab_45__31_,
         u5_mult_82_ab_45__32_, u5_mult_82_ab_45__33_, u5_mult_82_ab_45__34_,
         u5_mult_82_ab_45__35_, u5_mult_82_ab_45__36_, u5_mult_82_ab_45__37_,
         u5_mult_82_ab_45__38_, u5_mult_82_ab_45__39_, u5_mult_82_ab_45__40_,
         u5_mult_82_ab_45__41_, u5_mult_82_ab_45__42_, u5_mult_82_ab_45__43_,
         u5_mult_82_ab_45__44_, u5_mult_82_ab_45__45_, u5_mult_82_ab_45__46_,
         u5_mult_82_ab_45__47_, u5_mult_82_ab_45__48_, u5_mult_82_ab_45__49_,
         u5_mult_82_ab_45__50_, u5_mult_82_ab_45__51_, u5_mult_82_ab_45__52_,
         u5_mult_82_ab_46__0_, u5_mult_82_ab_46__1_, u5_mult_82_ab_46__2_,
         u5_mult_82_ab_46__3_, u5_mult_82_ab_46__4_, u5_mult_82_ab_46__5_,
         u5_mult_82_ab_46__6_, u5_mult_82_ab_46__7_, u5_mult_82_ab_46__8_,
         u5_mult_82_ab_46__9_, u5_mult_82_ab_46__10_, u5_mult_82_ab_46__11_,
         u5_mult_82_ab_46__12_, u5_mult_82_ab_46__13_, u5_mult_82_ab_46__14_,
         u5_mult_82_ab_46__15_, u5_mult_82_ab_46__16_, u5_mult_82_ab_46__17_,
         u5_mult_82_ab_46__18_, u5_mult_82_ab_46__19_, u5_mult_82_ab_46__20_,
         u5_mult_82_ab_46__21_, u5_mult_82_ab_46__22_, u5_mult_82_ab_46__23_,
         u5_mult_82_ab_46__24_, u5_mult_82_ab_46__25_, u5_mult_82_ab_46__26_,
         u5_mult_82_ab_46__27_, u5_mult_82_ab_46__28_, u5_mult_82_ab_46__29_,
         u5_mult_82_ab_46__30_, u5_mult_82_ab_46__31_, u5_mult_82_ab_46__32_,
         u5_mult_82_ab_46__33_, u5_mult_82_ab_46__34_, u5_mult_82_ab_46__35_,
         u5_mult_82_ab_46__36_, u5_mult_82_ab_46__37_, u5_mult_82_ab_46__38_,
         u5_mult_82_ab_46__39_, u5_mult_82_ab_46__40_, u5_mult_82_ab_46__41_,
         u5_mult_82_ab_46__42_, u5_mult_82_ab_46__43_, u5_mult_82_ab_46__44_,
         u5_mult_82_ab_46__45_, u5_mult_82_ab_46__46_, u5_mult_82_ab_46__47_,
         u5_mult_82_ab_46__48_, u5_mult_82_ab_46__49_, u5_mult_82_ab_46__50_,
         u5_mult_82_ab_46__51_, u5_mult_82_ab_46__52_, u5_mult_82_ab_47__0_,
         u5_mult_82_ab_47__1_, u5_mult_82_ab_47__2_, u5_mult_82_ab_47__3_,
         u5_mult_82_ab_47__4_, u5_mult_82_ab_47__5_, u5_mult_82_ab_47__6_,
         u5_mult_82_ab_47__7_, u5_mult_82_ab_47__9_, u5_mult_82_ab_47__10_,
         u5_mult_82_ab_47__11_, u5_mult_82_ab_47__12_, u5_mult_82_ab_47__13_,
         u5_mult_82_ab_47__14_, u5_mult_82_ab_47__15_, u5_mult_82_ab_47__16_,
         u5_mult_82_ab_47__17_, u5_mult_82_ab_47__18_, u5_mult_82_ab_47__19_,
         u5_mult_82_ab_47__20_, u5_mult_82_ab_47__21_, u5_mult_82_ab_47__22_,
         u5_mult_82_ab_47__23_, u5_mult_82_ab_47__24_, u5_mult_82_ab_47__25_,
         u5_mult_82_ab_47__26_, u5_mult_82_ab_47__27_, u5_mult_82_ab_47__28_,
         u5_mult_82_ab_47__29_, u5_mult_82_ab_47__30_, u5_mult_82_ab_47__31_,
         u5_mult_82_ab_47__32_, u5_mult_82_ab_47__33_, u5_mult_82_ab_47__34_,
         u5_mult_82_ab_47__35_, u5_mult_82_ab_47__36_, u5_mult_82_ab_47__37_,
         u5_mult_82_ab_47__38_, u5_mult_82_ab_47__39_, u5_mult_82_ab_47__40_,
         u5_mult_82_ab_47__41_, u5_mult_82_ab_47__42_, u5_mult_82_ab_47__43_,
         u5_mult_82_ab_47__44_, u5_mult_82_ab_47__45_, u5_mult_82_ab_47__46_,
         u5_mult_82_ab_47__47_, u5_mult_82_ab_47__48_, u5_mult_82_ab_47__49_,
         u5_mult_82_ab_47__50_, u5_mult_82_ab_47__51_, u5_mult_82_ab_47__52_,
         u5_mult_82_ab_48__0_, u5_mult_82_ab_48__1_, u5_mult_82_ab_48__2_,
         u5_mult_82_ab_48__3_, u5_mult_82_ab_48__4_, u5_mult_82_ab_48__5_,
         u5_mult_82_ab_48__6_, u5_mult_82_ab_48__7_, u5_mult_82_ab_48__8_,
         u5_mult_82_ab_48__9_, u5_mult_82_ab_48__10_, u5_mult_82_ab_48__11_,
         u5_mult_82_ab_48__12_, u5_mult_82_ab_48__13_, u5_mult_82_ab_48__14_,
         u5_mult_82_ab_48__15_, u5_mult_82_ab_48__16_, u5_mult_82_ab_48__17_,
         u5_mult_82_ab_48__18_, u5_mult_82_ab_48__19_, u5_mult_82_ab_48__20_,
         u5_mult_82_ab_48__21_, u5_mult_82_ab_48__22_, u5_mult_82_ab_48__23_,
         u5_mult_82_ab_48__24_, u5_mult_82_ab_48__25_, u5_mult_82_ab_48__26_,
         u5_mult_82_ab_48__27_, u5_mult_82_ab_48__28_, u5_mult_82_ab_48__29_,
         u5_mult_82_ab_48__30_, u5_mult_82_ab_48__31_, u5_mult_82_ab_48__32_,
         u5_mult_82_ab_48__33_, u5_mult_82_ab_48__34_, u5_mult_82_ab_48__35_,
         u5_mult_82_ab_48__36_, u5_mult_82_ab_48__37_, u5_mult_82_ab_48__38_,
         u5_mult_82_ab_48__39_, u5_mult_82_ab_48__40_, u5_mult_82_ab_48__41_,
         u5_mult_82_ab_48__42_, u5_mult_82_ab_48__43_, u5_mult_82_ab_48__44_,
         u5_mult_82_ab_48__45_, u5_mult_82_ab_48__46_, u5_mult_82_ab_48__47_,
         u5_mult_82_ab_48__48_, u5_mult_82_ab_48__49_, u5_mult_82_ab_48__50_,
         u5_mult_82_ab_48__51_, u5_mult_82_ab_48__52_, u5_mult_82_ab_49__0_,
         u5_mult_82_ab_49__1_, u5_mult_82_ab_49__2_, u5_mult_82_ab_49__3_,
         u5_mult_82_ab_49__4_, u5_mult_82_ab_49__5_, u5_mult_82_ab_49__6_,
         u5_mult_82_ab_49__7_, u5_mult_82_ab_49__8_, u5_mult_82_ab_49__9_,
         u5_mult_82_ab_49__10_, u5_mult_82_ab_49__11_, u5_mult_82_ab_49__12_,
         u5_mult_82_ab_49__13_, u5_mult_82_ab_49__14_, u5_mult_82_ab_49__15_,
         u5_mult_82_ab_49__16_, u5_mult_82_ab_49__17_, u5_mult_82_ab_49__18_,
         u5_mult_82_ab_49__19_, u5_mult_82_ab_49__20_, u5_mult_82_ab_49__21_,
         u5_mult_82_ab_49__22_, u5_mult_82_ab_49__23_, u5_mult_82_ab_49__24_,
         u5_mult_82_ab_49__25_, u5_mult_82_ab_49__26_, u5_mult_82_ab_49__27_,
         u5_mult_82_ab_49__28_, u5_mult_82_ab_49__29_, u5_mult_82_ab_49__30_,
         u5_mult_82_ab_49__31_, u5_mult_82_ab_49__32_, u5_mult_82_ab_49__33_,
         u5_mult_82_ab_49__34_, u5_mult_82_ab_49__35_, u5_mult_82_ab_49__36_,
         u5_mult_82_ab_49__37_, u5_mult_82_ab_49__38_, u5_mult_82_ab_49__39_,
         u5_mult_82_ab_49__40_, u5_mult_82_ab_49__41_, u5_mult_82_ab_49__42_,
         u5_mult_82_ab_49__43_, u5_mult_82_ab_49__44_, u5_mult_82_ab_49__45_,
         u5_mult_82_ab_49__46_, u5_mult_82_ab_49__47_, u5_mult_82_ab_49__48_,
         u5_mult_82_ab_49__49_, u5_mult_82_ab_49__50_, u5_mult_82_ab_49__51_,
         u5_mult_82_ab_49__52_, u5_mult_82_ab_50__0_, u5_mult_82_ab_50__1_,
         u5_mult_82_ab_50__2_, u5_mult_82_ab_50__3_, u5_mult_82_ab_50__4_,
         u5_mult_82_ab_50__7_, u5_mult_82_ab_50__8_, u5_mult_82_ab_50__9_,
         u5_mult_82_ab_50__10_, u5_mult_82_ab_50__11_, u5_mult_82_ab_50__12_,
         u5_mult_82_ab_50__13_, u5_mult_82_ab_50__14_, u5_mult_82_ab_50__15_,
         u5_mult_82_ab_50__16_, u5_mult_82_ab_50__17_, u5_mult_82_ab_50__18_,
         u5_mult_82_ab_50__19_, u5_mult_82_ab_50__20_, u5_mult_82_ab_50__21_,
         u5_mult_82_ab_50__22_, u5_mult_82_ab_50__23_, u5_mult_82_ab_50__24_,
         u5_mult_82_ab_50__25_, u5_mult_82_ab_50__26_, u5_mult_82_ab_50__27_,
         u5_mult_82_ab_50__28_, u5_mult_82_ab_50__29_, u5_mult_82_ab_50__30_,
         u5_mult_82_ab_50__31_, u5_mult_82_ab_50__32_, u5_mult_82_ab_50__33_,
         u5_mult_82_ab_50__34_, u5_mult_82_ab_50__35_, u5_mult_82_ab_50__36_,
         u5_mult_82_ab_50__37_, u5_mult_82_ab_50__38_, u5_mult_82_ab_50__39_,
         u5_mult_82_ab_50__40_, u5_mult_82_ab_50__41_, u5_mult_82_ab_50__42_,
         u5_mult_82_ab_50__43_, u5_mult_82_ab_50__44_, u5_mult_82_ab_50__45_,
         u5_mult_82_ab_50__46_, u5_mult_82_ab_50__47_, u5_mult_82_ab_50__48_,
         u5_mult_82_ab_50__49_, u5_mult_82_ab_50__50_, u5_mult_82_ab_50__51_,
         u5_mult_82_ab_50__52_, u5_mult_82_ab_51__0_, u5_mult_82_ab_51__1_,
         u5_mult_82_ab_51__2_, u5_mult_82_ab_51__3_, u5_mult_82_ab_51__4_,
         u5_mult_82_ab_51__5_, u5_mult_82_ab_51__7_, u5_mult_82_ab_51__8_,
         u5_mult_82_ab_51__9_, u5_mult_82_ab_51__10_, u5_mult_82_ab_51__11_,
         u5_mult_82_ab_51__12_, u5_mult_82_ab_51__13_, u5_mult_82_ab_51__14_,
         u5_mult_82_ab_51__15_, u5_mult_82_ab_51__16_, u5_mult_82_ab_51__17_,
         u5_mult_82_ab_51__18_, u5_mult_82_ab_51__19_, u5_mult_82_ab_51__20_,
         u5_mult_82_ab_51__21_, u5_mult_82_ab_51__22_, u5_mult_82_ab_51__23_,
         u5_mult_82_ab_51__24_, u5_mult_82_ab_51__25_, u5_mult_82_ab_51__26_,
         u5_mult_82_ab_51__27_, u5_mult_82_ab_51__28_, u5_mult_82_ab_51__29_,
         u5_mult_82_ab_51__30_, u5_mult_82_ab_51__31_, u5_mult_82_ab_51__32_,
         u5_mult_82_ab_51__33_, u5_mult_82_ab_51__34_, u5_mult_82_ab_51__35_,
         u5_mult_82_ab_51__36_, u5_mult_82_ab_51__37_, u5_mult_82_ab_51__38_,
         u5_mult_82_ab_51__39_, u5_mult_82_ab_51__40_, u5_mult_82_ab_51__41_,
         u5_mult_82_ab_51__42_, u5_mult_82_ab_51__43_, u5_mult_82_ab_51__44_,
         u5_mult_82_ab_51__45_, u5_mult_82_ab_51__46_, u5_mult_82_ab_51__47_,
         u5_mult_82_ab_51__48_, u5_mult_82_ab_51__49_, u5_mult_82_ab_51__50_,
         u5_mult_82_ab_51__51_, u5_mult_82_ab_51__52_, u5_mult_82_ab_52__0_,
         u5_mult_82_ab_52__1_, u5_mult_82_ab_52__2_, u5_mult_82_ab_52__3_,
         u5_mult_82_ab_52__4_, u5_mult_82_ab_52__5_, u5_mult_82_ab_52__6_,
         u5_mult_82_ab_52__7_, u5_mult_82_ab_52__8_, u5_mult_82_ab_52__9_,
         u5_mult_82_ab_52__10_, u5_mult_82_ab_52__11_, u5_mult_82_ab_52__12_,
         u5_mult_82_ab_52__13_, u5_mult_82_ab_52__14_, u5_mult_82_ab_52__15_,
         u5_mult_82_ab_52__16_, u5_mult_82_ab_52__17_, u5_mult_82_ab_52__18_,
         u5_mult_82_ab_52__19_, u5_mult_82_ab_52__20_, u5_mult_82_ab_52__21_,
         u5_mult_82_ab_52__22_, u5_mult_82_ab_52__23_, u5_mult_82_ab_52__24_,
         u5_mult_82_ab_52__25_, u5_mult_82_ab_52__26_, u5_mult_82_ab_52__27_,
         u5_mult_82_ab_52__28_, u5_mult_82_ab_52__29_, u5_mult_82_ab_52__30_,
         u5_mult_82_ab_52__31_, u5_mult_82_ab_52__32_, u5_mult_82_ab_52__33_,
         u5_mult_82_ab_52__34_, u5_mult_82_ab_52__35_, u5_mult_82_ab_52__36_,
         u5_mult_82_ab_52__37_, u5_mult_82_ab_52__38_, u5_mult_82_ab_52__39_,
         u5_mult_82_ab_52__40_, u5_mult_82_ab_52__41_, u5_mult_82_ab_52__42_,
         u5_mult_82_ab_52__43_, u5_mult_82_ab_52__44_, u5_mult_82_ab_52__45_,
         u5_mult_82_ab_52__46_, u5_mult_82_ab_52__47_, u5_mult_82_ab_52__48_,
         u5_mult_82_ab_52__49_, u5_mult_82_ab_52__50_, u5_mult_82_ab_52__51_,
         u5_mult_82_ab_52__52_, u5_mult_82_FS_1_n743, u5_mult_82_FS_1_n742,
         u5_mult_82_FS_1_n741, u5_mult_82_FS_1_n740, u5_mult_82_FS_1_n739,
         u5_mult_82_FS_1_n738, u5_mult_82_FS_1_n737, u5_mult_82_FS_1_n736,
         u5_mult_82_FS_1_n735, u5_mult_82_FS_1_n734, u5_mult_82_FS_1_n733,
         u5_mult_82_FS_1_n732, u5_mult_82_FS_1_n731, u5_mult_82_FS_1_n730,
         u5_mult_82_FS_1_n729, u5_mult_82_FS_1_n728, u5_mult_82_FS_1_n727,
         u5_mult_82_FS_1_n726, u5_mult_82_FS_1_n725, u5_mult_82_FS_1_n724,
         u5_mult_82_FS_1_n723, u5_mult_82_FS_1_n722, u5_mult_82_FS_1_n721,
         u5_mult_82_FS_1_n720, u5_mult_82_FS_1_n719, u5_mult_82_FS_1_n718,
         u5_mult_82_FS_1_n717, u5_mult_82_FS_1_n716, u5_mult_82_FS_1_n715,
         u5_mult_82_FS_1_n714, u5_mult_82_FS_1_n713, u5_mult_82_FS_1_n712,
         u5_mult_82_FS_1_n711, u5_mult_82_FS_1_n710, u5_mult_82_FS_1_n709,
         u5_mult_82_FS_1_n708, u5_mult_82_FS_1_n707, u5_mult_82_FS_1_n706,
         u5_mult_82_FS_1_n705, u5_mult_82_FS_1_n704, u5_mult_82_FS_1_n703,
         u5_mult_82_FS_1_n702, u5_mult_82_FS_1_n701, u5_mult_82_FS_1_n700,
         u5_mult_82_FS_1_n699, u5_mult_82_FS_1_n698, u5_mult_82_FS_1_n697,
         u5_mult_82_FS_1_n696, u5_mult_82_FS_1_n695, u5_mult_82_FS_1_n694,
         u5_mult_82_FS_1_n693, u5_mult_82_FS_1_n692, u5_mult_82_FS_1_n691,
         u5_mult_82_FS_1_n690, u5_mult_82_FS_1_n689, u5_mult_82_FS_1_n688,
         u5_mult_82_FS_1_n687, u5_mult_82_FS_1_n686, u5_mult_82_FS_1_n685,
         u5_mult_82_FS_1_n684, u5_mult_82_FS_1_n683, u5_mult_82_FS_1_n682,
         u5_mult_82_FS_1_n681, u5_mult_82_FS_1_n680, u5_mult_82_FS_1_n679,
         u5_mult_82_FS_1_n678, u5_mult_82_FS_1_n677, u5_mult_82_FS_1_n676,
         u5_mult_82_FS_1_n675, u5_mult_82_FS_1_n674, u5_mult_82_FS_1_n673,
         u5_mult_82_FS_1_n672, u5_mult_82_FS_1_n671, u5_mult_82_FS_1_n670,
         u5_mult_82_FS_1_n669, u5_mult_82_FS_1_n668, u5_mult_82_FS_1_n667,
         u5_mult_82_FS_1_n666, u5_mult_82_FS_1_n665, u5_mult_82_FS_1_n664,
         u5_mult_82_FS_1_n663, u5_mult_82_FS_1_n662, u5_mult_82_FS_1_n661,
         u5_mult_82_FS_1_n660, u5_mult_82_FS_1_n659, u5_mult_82_FS_1_n658,
         u5_mult_82_FS_1_n657, u5_mult_82_FS_1_n656, u5_mult_82_FS_1_n655,
         u5_mult_82_FS_1_n654, u5_mult_82_FS_1_n653, u5_mult_82_FS_1_n652,
         u5_mult_82_FS_1_n651, u5_mult_82_FS_1_n650, u5_mult_82_FS_1_n649,
         u5_mult_82_FS_1_n648, u5_mult_82_FS_1_n647, u5_mult_82_FS_1_n646,
         u5_mult_82_FS_1_n645, u5_mult_82_FS_1_n644, u5_mult_82_FS_1_n643,
         u5_mult_82_FS_1_n642, u5_mult_82_FS_1_n641, u5_mult_82_FS_1_n640,
         u5_mult_82_FS_1_n639, u5_mult_82_FS_1_n638, u5_mult_82_FS_1_n637,
         u5_mult_82_FS_1_n636, u5_mult_82_FS_1_n635, u5_mult_82_FS_1_n634,
         u5_mult_82_FS_1_n633, u5_mult_82_FS_1_n632, u5_mult_82_FS_1_n631,
         u5_mult_82_FS_1_n630, u5_mult_82_FS_1_n629, u5_mult_82_FS_1_n628,
         u5_mult_82_FS_1_n627, u5_mult_82_FS_1_n626, u5_mult_82_FS_1_n625,
         u5_mult_82_FS_1_n624, u5_mult_82_FS_1_n623, u5_mult_82_FS_1_n622,
         u5_mult_82_FS_1_n621, u5_mult_82_FS_1_n620, u5_mult_82_FS_1_n619,
         u5_mult_82_FS_1_n618, u5_mult_82_FS_1_n617, u5_mult_82_FS_1_n616,
         u5_mult_82_FS_1_n615, u5_mult_82_FS_1_n614, u5_mult_82_FS_1_n613,
         u5_mult_82_FS_1_n612, u5_mult_82_FS_1_n611, u5_mult_82_FS_1_n610,
         u5_mult_82_FS_1_n609, u5_mult_82_FS_1_n608, u5_mult_82_FS_1_n607,
         u5_mult_82_FS_1_n606, u5_mult_82_FS_1_n605, u5_mult_82_FS_1_n604,
         u5_mult_82_FS_1_n603, u5_mult_82_FS_1_n602, u5_mult_82_FS_1_n601,
         u5_mult_82_FS_1_n600, u5_mult_82_FS_1_n599, u5_mult_82_FS_1_n598,
         u5_mult_82_FS_1_n597, u5_mult_82_FS_1_n596, u5_mult_82_FS_1_n595,
         u5_mult_82_FS_1_n594, u5_mult_82_FS_1_n593, u5_mult_82_FS_1_n592,
         u5_mult_82_FS_1_n591, u5_mult_82_FS_1_n590, u5_mult_82_FS_1_n589,
         u5_mult_82_FS_1_n588, u5_mult_82_FS_1_n587, u5_mult_82_FS_1_n586,
         u5_mult_82_FS_1_n585, u5_mult_82_FS_1_n584, u5_mult_82_FS_1_n583,
         u5_mult_82_FS_1_n582, u5_mult_82_FS_1_n581, u5_mult_82_FS_1_n580,
         u5_mult_82_FS_1_n579, u5_mult_82_FS_1_n578, u5_mult_82_FS_1_n577,
         u5_mult_82_FS_1_n576, u5_mult_82_FS_1_n575, u5_mult_82_FS_1_n574,
         u5_mult_82_FS_1_n573, u5_mult_82_FS_1_n572, u5_mult_82_FS_1_n571,
         u5_mult_82_FS_1_n570, u5_mult_82_FS_1_n569, u5_mult_82_FS_1_n568,
         u5_mult_82_FS_1_n567, u5_mult_82_FS_1_n566, u5_mult_82_FS_1_n565,
         u5_mult_82_FS_1_n564, u5_mult_82_FS_1_n563, u5_mult_82_FS_1_n562,
         u5_mult_82_FS_1_n561, u5_mult_82_FS_1_n560, u5_mult_82_FS_1_n559,
         u5_mult_82_FS_1_n558, u5_mult_82_FS_1_n557, u5_mult_82_FS_1_n556,
         u5_mult_82_FS_1_n555, u5_mult_82_FS_1_n554, u5_mult_82_FS_1_n553,
         u5_mult_82_FS_1_n552, u5_mult_82_FS_1_n551, u5_mult_82_FS_1_n550,
         u5_mult_82_FS_1_n549, u5_mult_82_FS_1_n548, u5_mult_82_FS_1_n547,
         u5_mult_82_FS_1_n546, u5_mult_82_FS_1_n545, u5_mult_82_FS_1_n544,
         u5_mult_82_FS_1_n543, u5_mult_82_FS_1_n542, u5_mult_82_FS_1_n541,
         u5_mult_82_FS_1_n540, u5_mult_82_FS_1_n539, u5_mult_82_FS_1_n538,
         u5_mult_82_FS_1_n537, u5_mult_82_FS_1_n536, u5_mult_82_FS_1_n535,
         u5_mult_82_FS_1_n534, u5_mult_82_FS_1_n533, u5_mult_82_FS_1_n532,
         u5_mult_82_FS_1_n531, u5_mult_82_FS_1_n530, u5_mult_82_FS_1_n529,
         u5_mult_82_FS_1_n528, u5_mult_82_FS_1_n527, u5_mult_82_FS_1_n526,
         u5_mult_82_FS_1_n525, u5_mult_82_FS_1_n524, u5_mult_82_FS_1_n523,
         u5_mult_82_FS_1_n522, u5_mult_82_FS_1_n521, u5_mult_82_FS_1_n520,
         u5_mult_82_FS_1_n519, u5_mult_82_FS_1_n518, u5_mult_82_FS_1_n517,
         u5_mult_82_FS_1_n516, u5_mult_82_FS_1_n515, u5_mult_82_FS_1_n514,
         u5_mult_82_FS_1_n513, u5_mult_82_FS_1_n512, u5_mult_82_FS_1_n511,
         u5_mult_82_FS_1_n510, u5_mult_82_FS_1_n509, u5_mult_82_FS_1_n508,
         u5_mult_82_FS_1_n507, u5_mult_82_FS_1_n506, u5_mult_82_FS_1_n505,
         u5_mult_82_FS_1_n504, u5_mult_82_FS_1_n503, u5_mult_82_FS_1_n502,
         u5_mult_82_FS_1_n501, u5_mult_82_FS_1_n500, u5_mult_82_FS_1_n499,
         u5_mult_82_FS_1_n498, u5_mult_82_FS_1_n497, u5_mult_82_FS_1_n496,
         u5_mult_82_FS_1_n495, u5_mult_82_FS_1_n494, u5_mult_82_FS_1_n493,
         u5_mult_82_FS_1_n492, u5_mult_82_FS_1_n491, u5_mult_82_FS_1_n490,
         u5_mult_82_FS_1_n489, u5_mult_82_FS_1_n488, u5_mult_82_FS_1_n487,
         u5_mult_82_FS_1_n486, u5_mult_82_FS_1_n485, u5_mult_82_FS_1_n484,
         u5_mult_82_FS_1_n483, u5_mult_82_FS_1_n482, u5_mult_82_FS_1_n481,
         u5_mult_82_FS_1_n480, u5_mult_82_FS_1_n479, u5_mult_82_FS_1_n478,
         u5_mult_82_FS_1_n477, u5_mult_82_FS_1_n476, u5_mult_82_FS_1_n475,
         u5_mult_82_FS_1_n474, u5_mult_82_FS_1_n473, u5_mult_82_FS_1_n472,
         u5_mult_82_FS_1_n471, u5_mult_82_FS_1_n470, u5_mult_82_FS_1_n469,
         u5_mult_82_FS_1_n468, u5_mult_82_FS_1_n467, u5_mult_82_FS_1_n466,
         u5_mult_82_FS_1_n465, u5_mult_82_FS_1_n464, u5_mult_82_FS_1_n463,
         u5_mult_82_FS_1_n462, u5_mult_82_FS_1_n461, u5_mult_82_FS_1_n460,
         u5_mult_82_FS_1_n459, u5_mult_82_FS_1_n458, u5_mult_82_FS_1_n457,
         u5_mult_82_FS_1_n456, u5_mult_82_FS_1_n455, u5_mult_82_FS_1_n454,
         u5_mult_82_FS_1_n453, u5_mult_82_FS_1_n452, u5_mult_82_FS_1_n451,
         u5_mult_82_FS_1_n450, u5_mult_82_FS_1_n449, u5_mult_82_FS_1_n448,
         u5_mult_82_FS_1_n447, u5_mult_82_FS_1_n446, u5_mult_82_FS_1_n445,
         u5_mult_82_FS_1_n444, u5_mult_82_FS_1_n443, u5_mult_82_FS_1_n442,
         u5_mult_82_FS_1_n441, u5_mult_82_FS_1_n440, u5_mult_82_FS_1_n439,
         u5_mult_82_FS_1_n438, u5_mult_82_FS_1_n437, u5_mult_82_FS_1_n436,
         u5_mult_82_FS_1_n435, u5_mult_82_FS_1_n434, u5_mult_82_FS_1_n433,
         u5_mult_82_FS_1_n432, u5_mult_82_FS_1_n431, u5_mult_82_FS_1_n430,
         u5_mult_82_FS_1_n429, u5_mult_82_FS_1_n428, u5_mult_82_FS_1_n427,
         u5_mult_82_FS_1_n426, u5_mult_82_FS_1_n425, u5_mult_82_FS_1_n424,
         u5_mult_82_FS_1_n423, u5_mult_82_FS_1_n422, u5_mult_82_FS_1_n421,
         u5_mult_82_FS_1_n420, u5_mult_82_FS_1_n419, u5_mult_82_FS_1_n418,
         u5_mult_82_FS_1_n417, u5_mult_82_FS_1_n416, u5_mult_82_FS_1_n415,
         u5_mult_82_FS_1_n414, u5_mult_82_FS_1_n413, u5_mult_82_FS_1_n412,
         u5_mult_82_FS_1_n411, u5_mult_82_FS_1_n410, u5_mult_82_FS_1_n409,
         u5_mult_82_FS_1_n408, u5_mult_82_FS_1_n407, u5_mult_82_FS_1_n406,
         u5_mult_82_FS_1_n405, u5_mult_82_FS_1_n404, u5_mult_82_FS_1_n403,
         u5_mult_82_FS_1_n402, u5_mult_82_FS_1_n401, u5_mult_82_FS_1_n400,
         u5_mult_82_FS_1_n399, u5_mult_82_FS_1_n398, u5_mult_82_FS_1_n397,
         u5_mult_82_FS_1_n396, u5_mult_82_FS_1_n395, u5_mult_82_FS_1_n394,
         u5_mult_82_FS_1_n393, u5_mult_82_FS_1_n392, u5_mult_82_FS_1_n391,
         u5_mult_82_FS_1_n390, u5_mult_82_FS_1_n389, u5_mult_82_FS_1_n388,
         u5_mult_82_FS_1_n387, u5_mult_82_FS_1_n386, u5_mult_82_FS_1_n385,
         u5_mult_82_FS_1_n384, u5_mult_82_FS_1_n383, u5_mult_82_FS_1_n382,
         u5_mult_82_FS_1_n381, u5_mult_82_FS_1_n380, u5_mult_82_FS_1_n379,
         u5_mult_82_FS_1_n378, u5_mult_82_FS_1_n377, u5_mult_82_FS_1_n376,
         u5_mult_82_FS_1_n375, u5_mult_82_FS_1_n374, u5_mult_82_FS_1_n373,
         u5_mult_82_FS_1_n372, u5_mult_82_FS_1_n371, u5_mult_82_FS_1_n370,
         u5_mult_82_FS_1_n369, u5_mult_82_FS_1_n368, u5_mult_82_FS_1_n367,
         u5_mult_82_FS_1_n366, u5_mult_82_FS_1_n365, u5_mult_82_FS_1_n364,
         u5_mult_82_FS_1_n363, u5_mult_82_FS_1_n362, u5_mult_82_FS_1_n361,
         u5_mult_82_FS_1_n360, u5_mult_82_FS_1_n359, u5_mult_82_FS_1_n358,
         u5_mult_82_FS_1_n357, u5_mult_82_FS_1_n356, u5_mult_82_FS_1_n355,
         u5_mult_82_FS_1_n354, u5_mult_82_FS_1_n353, u5_mult_82_FS_1_n352,
         u5_mult_82_FS_1_n351, u5_mult_82_FS_1_n350, u5_mult_82_FS_1_n349,
         u5_mult_82_FS_1_n348, u5_mult_82_FS_1_n347, u5_mult_82_FS_1_n346,
         u5_mult_82_FS_1_n345, u5_mult_82_FS_1_n344, u5_mult_82_FS_1_n343,
         u5_mult_82_FS_1_n342, u5_mult_82_FS_1_n341, u5_mult_82_FS_1_n340,
         u5_mult_82_FS_1_n339, u5_mult_82_FS_1_n338, u5_mult_82_FS_1_n337,
         u5_mult_82_FS_1_n336, u5_mult_82_FS_1_n335, u5_mult_82_FS_1_n334,
         u5_mult_82_FS_1_n333, u5_mult_82_FS_1_n332, u5_mult_82_FS_1_n331,
         u5_mult_82_FS_1_n330, u5_mult_82_FS_1_n329, u5_mult_82_FS_1_n328,
         u5_mult_82_FS_1_n327, u5_mult_82_FS_1_n326, u5_mult_82_FS_1_n325,
         u5_mult_82_FS_1_n324, u5_mult_82_FS_1_n323, u5_mult_82_FS_1_n322,
         u5_mult_82_FS_1_n321, u5_mult_82_FS_1_n320, u5_mult_82_FS_1_n319,
         u5_mult_82_FS_1_n318, u5_mult_82_FS_1_n317, u5_mult_82_FS_1_n316,
         u5_mult_82_FS_1_n315, u5_mult_82_FS_1_n314, u5_mult_82_FS_1_n313,
         u5_mult_82_FS_1_n312, u5_mult_82_FS_1_n311, u5_mult_82_FS_1_n310,
         u5_mult_82_FS_1_n309, u5_mult_82_FS_1_n308, u5_mult_82_FS_1_n307,
         u5_mult_82_FS_1_n306, u5_mult_82_FS_1_n305, u5_mult_82_FS_1_n304,
         u5_mult_82_FS_1_n303, u5_mult_82_FS_1_n302, u5_mult_82_FS_1_n301,
         u5_mult_82_FS_1_n300, u5_mult_82_FS_1_n299, u5_mult_82_FS_1_n298,
         u5_mult_82_FS_1_n297, u5_mult_82_FS_1_n296, u5_mult_82_FS_1_n295,
         u5_mult_82_FS_1_n294, u5_mult_82_FS_1_n293, u5_mult_82_FS_1_n292,
         u5_mult_82_FS_1_n291, u5_mult_82_FS_1_n290, u5_mult_82_FS_1_n289,
         u5_mult_82_FS_1_n288, u5_mult_82_FS_1_n287, u5_mult_82_FS_1_n286,
         u5_mult_82_FS_1_n285, u5_mult_82_FS_1_n284, u5_mult_82_FS_1_n283,
         u5_mult_82_FS_1_n282, u5_mult_82_FS_1_n281, u5_mult_82_FS_1_n280,
         u5_mult_82_FS_1_n279, u5_mult_82_FS_1_n278, u5_mult_82_FS_1_n277,
         u5_mult_82_FS_1_n276, u5_mult_82_FS_1_n275, u5_mult_82_FS_1_n274,
         u5_mult_82_FS_1_n273, u5_mult_82_FS_1_n272, u5_mult_82_FS_1_n271,
         u5_mult_82_FS_1_n270, u5_mult_82_FS_1_n269, u5_mult_82_FS_1_n268,
         u5_mult_82_FS_1_n267, u5_mult_82_FS_1_n266, u5_mult_82_FS_1_n265,
         u5_mult_82_FS_1_n264, u5_mult_82_FS_1_n263, u5_mult_82_FS_1_n262,
         u5_mult_82_FS_1_n261, u5_mult_82_FS_1_n260, u5_mult_82_FS_1_n259,
         u5_mult_82_FS_1_n258, u5_mult_82_FS_1_n257, u5_mult_82_FS_1_n256,
         u5_mult_82_FS_1_n255, u5_mult_82_FS_1_n254, u5_mult_82_FS_1_n253,
         u5_mult_82_FS_1_n252, u5_mult_82_FS_1_n251, u5_mult_82_FS_1_n250,
         u5_mult_82_FS_1_n249, u5_mult_82_FS_1_n248, u5_mult_82_FS_1_n247,
         u5_mult_82_FS_1_n246, u5_mult_82_FS_1_n245, u5_mult_82_FS_1_n244,
         u5_mult_82_FS_1_n243, u5_mult_82_FS_1_n242, u5_mult_82_FS_1_n241,
         u5_mult_82_FS_1_n240, u5_mult_82_FS_1_n239, u5_mult_82_FS_1_n238,
         u5_mult_82_FS_1_n237, u5_mult_82_FS_1_n236, u5_mult_82_FS_1_n235,
         u5_mult_82_FS_1_n234, u5_mult_82_FS_1_n233, u5_mult_82_FS_1_n232,
         u5_mult_82_FS_1_n231, u5_mult_82_FS_1_n230, u5_mult_82_FS_1_n229,
         u5_mult_82_FS_1_n228, u5_mult_82_FS_1_n227, u5_mult_82_FS_1_n226,
         u5_mult_82_FS_1_n225, u5_mult_82_FS_1_n224, u5_mult_82_FS_1_n223,
         u5_mult_82_FS_1_n222, u5_mult_82_FS_1_n221, u5_mult_82_FS_1_n220,
         u5_mult_82_FS_1_n219, u5_mult_82_FS_1_n218, u5_mult_82_FS_1_n217,
         u5_mult_82_FS_1_n216, u5_mult_82_FS_1_n215, u5_mult_82_FS_1_n214,
         u5_mult_82_FS_1_n213, u5_mult_82_FS_1_n212, u5_mult_82_FS_1_n211,
         u5_mult_82_FS_1_n210, u5_mult_82_FS_1_n209, u5_mult_82_FS_1_n208,
         u5_mult_82_FS_1_n207, u5_mult_82_FS_1_n206, u5_mult_82_FS_1_n205,
         u5_mult_82_FS_1_n204, u5_mult_82_FS_1_n203, u5_mult_82_FS_1_n202,
         u5_mult_82_FS_1_n201, u5_mult_82_FS_1_n200, u5_mult_82_FS_1_n199,
         u5_mult_82_FS_1_n198, u5_mult_82_FS_1_n197, u5_mult_82_FS_1_n196,
         u5_mult_82_FS_1_n195, u5_mult_82_FS_1_n194, u5_mult_82_FS_1_n193,
         u5_mult_82_FS_1_n192, u5_mult_82_FS_1_n191, u5_mult_82_FS_1_n190,
         u5_mult_82_FS_1_n189, u5_mult_82_FS_1_n188, u5_mult_82_FS_1_n187,
         u5_mult_82_FS_1_n186, u5_mult_82_FS_1_n185, u5_mult_82_FS_1_n184,
         u5_mult_82_FS_1_n183, u5_mult_82_FS_1_n182, u5_mult_82_FS_1_n181,
         u5_mult_82_FS_1_n180, u5_mult_82_FS_1_n179, u5_mult_82_FS_1_n178,
         u5_mult_82_FS_1_n177, u5_mult_82_FS_1_n176, u5_mult_82_FS_1_n175,
         u5_mult_82_FS_1_n174, u5_mult_82_FS_1_n173, u5_mult_82_FS_1_n172,
         u5_mult_82_FS_1_n171, u5_mult_82_FS_1_n170, u5_mult_82_FS_1_n169,
         u5_mult_82_FS_1_n168, u5_mult_82_FS_1_n167, u5_mult_82_FS_1_n166,
         u5_mult_82_FS_1_n165, u5_mult_82_FS_1_n164, u5_mult_82_FS_1_n163,
         u5_mult_82_FS_1_n162, u5_mult_82_FS_1_n161, u5_mult_82_FS_1_n160,
         u5_mult_82_FS_1_n159, u5_mult_82_FS_1_n158, u5_mult_82_FS_1_n157,
         u5_mult_82_FS_1_n156, u5_mult_82_FS_1_n155, u5_mult_82_FS_1_n154,
         u5_mult_82_FS_1_n153, u5_mult_82_FS_1_n152, u5_mult_82_FS_1_n151,
         u5_mult_82_FS_1_n150, u5_mult_82_FS_1_n149, u5_mult_82_FS_1_n148,
         u5_mult_82_FS_1_n147, u5_mult_82_FS_1_n146, u5_mult_82_FS_1_n145,
         u5_mult_82_FS_1_n144, u5_mult_82_FS_1_n143, u5_mult_82_FS_1_n142,
         u5_mult_82_FS_1_n141, u5_mult_82_FS_1_n140, u5_mult_82_FS_1_n139,
         u5_mult_82_FS_1_n138, u5_mult_82_FS_1_n137, u5_mult_82_FS_1_n136,
         u5_mult_82_FS_1_n135, u5_mult_82_FS_1_n134, u5_mult_82_FS_1_n133,
         u5_mult_82_FS_1_n132, u5_mult_82_FS_1_n131, u5_mult_82_FS_1_n130,
         u5_mult_82_FS_1_n129, u5_mult_82_FS_1_n128, u5_mult_82_FS_1_n127,
         u5_mult_82_FS_1_n126, u5_mult_82_FS_1_n125, u5_mult_82_FS_1_n124,
         u5_mult_82_FS_1_n123, u5_mult_82_FS_1_n122, u5_mult_82_FS_1_n121,
         u5_mult_82_FS_1_n120, u5_mult_82_FS_1_n119, u5_mult_82_FS_1_n118,
         u5_mult_82_FS_1_n117, u5_mult_82_FS_1_n116, u5_mult_82_FS_1_n115,
         u5_mult_82_FS_1_n114, u5_mult_82_FS_1_n113, u5_mult_82_FS_1_n112,
         u5_mult_82_FS_1_n111, u5_mult_82_FS_1_n110, u5_mult_82_FS_1_n109,
         u5_mult_82_FS_1_n108, u5_mult_82_FS_1_n107, u5_mult_82_FS_1_n106,
         u5_mult_82_FS_1_n105, u5_mult_82_FS_1_n104, u5_mult_82_FS_1_n103,
         u5_mult_82_FS_1_n102, u5_mult_82_FS_1_n101, u5_mult_82_FS_1_n100,
         u5_mult_82_FS_1_n99, u5_mult_82_FS_1_n98, u5_mult_82_FS_1_n97,
         u5_mult_82_FS_1_n96, u5_mult_82_FS_1_n95, u5_mult_82_FS_1_n94,
         u5_mult_82_FS_1_n93, u5_mult_82_FS_1_n92, u5_mult_82_FS_1_n91,
         u5_mult_82_FS_1_n90, u5_mult_82_FS_1_n89, u5_mult_82_FS_1_n88,
         u5_mult_82_FS_1_n87, u5_mult_82_FS_1_n86, u5_mult_82_FS_1_n85,
         u5_mult_82_FS_1_n84, u5_mult_82_FS_1_n83, u5_mult_82_FS_1_n82,
         u5_mult_82_FS_1_n81, u5_mult_82_FS_1_n80, u5_mult_82_FS_1_n79,
         u5_mult_82_FS_1_n78, u5_mult_82_FS_1_n77, u5_mult_82_FS_1_n76,
         u5_mult_82_FS_1_n75, u5_mult_82_FS_1_n74, u5_mult_82_FS_1_n73,
         u5_mult_82_FS_1_n72, u5_mult_82_FS_1_n71, u5_mult_82_FS_1_n70,
         u5_mult_82_FS_1_n69, u5_mult_82_FS_1_n68, u5_mult_82_FS_1_n67,
         u5_mult_82_FS_1_n66, u5_mult_82_FS_1_n65, u5_mult_82_FS_1_n64,
         u5_mult_82_FS_1_n63, u5_mult_82_FS_1_n62, u5_mult_82_FS_1_n61,
         u5_mult_82_FS_1_n60, u5_mult_82_FS_1_n59, u5_mult_82_FS_1_n58,
         u5_mult_82_FS_1_n57, u5_mult_82_FS_1_n56, u5_mult_82_FS_1_n55,
         u5_mult_82_FS_1_n54, u5_mult_82_FS_1_n53, u5_mult_82_FS_1_n52,
         u5_mult_82_FS_1_n51, u5_mult_82_FS_1_n50, u5_mult_82_FS_1_n49,
         u5_mult_82_FS_1_n48, u5_mult_82_FS_1_n47, u5_mult_82_FS_1_n46,
         u5_mult_82_FS_1_n45, u5_mult_82_FS_1_n44, u5_mult_82_FS_1_n43,
         u5_mult_82_FS_1_n42, u5_mult_82_FS_1_n41, u5_mult_82_FS_1_n40,
         u5_mult_82_FS_1_n39, u5_mult_82_FS_1_n38, u5_mult_82_FS_1_n37,
         u5_mult_82_FS_1_n36, u5_mult_82_FS_1_n35, u5_mult_82_FS_1_n34,
         u5_mult_82_FS_1_n33, u5_mult_82_FS_1_n32, u5_mult_82_FS_1_n31,
         u5_mult_82_FS_1_n30, u5_mult_82_FS_1_n29, u5_mult_82_FS_1_n28,
         u5_mult_82_FS_1_n27, u5_mult_82_FS_1_n26, u5_mult_82_FS_1_n25,
         u5_mult_82_FS_1_n24, u5_mult_82_FS_1_n23, u5_mult_82_FS_1_n22,
         u5_mult_82_FS_1_n21, u5_mult_82_FS_1_n20, u5_mult_82_FS_1_n19,
         u5_mult_82_FS_1_n18, u5_mult_82_FS_1_n17, u5_mult_82_FS_1_n16,
         u5_mult_82_FS_1_n15, u5_mult_82_FS_1_n14, u5_mult_82_FS_1_n13,
         u5_mult_82_FS_1_n12, u5_mult_82_FS_1_n11, u5_mult_82_FS_1_n10,
         u5_mult_82_FS_1_n9, u5_mult_82_FS_1_n8, u5_mult_82_FS_1_n7,
         u5_mult_82_FS_1_n6, u5_mult_82_FS_1_n5, u5_mult_82_FS_1_n4,
         u5_mult_82_FS_1_n3, u5_mult_82_FS_1_n2, u5_mult_82_FS_1_n1,
         u4_sub_470_n100, u4_sub_470_n99, u4_sub_470_n98, u4_sub_470_n97,
         u4_sub_470_n96, u4_sub_470_n95, u4_sub_470_n94, u4_sub_470_n93,
         u4_sub_470_n92, u4_sub_470_n91, u4_sub_470_n90, u4_sub_470_n89,
         u4_sub_470_n88, u4_sub_470_n87, u4_sub_470_n86, u4_sub_470_n85,
         u4_sub_470_n84, u4_sub_470_n83, u4_sub_470_n82, u4_sub_470_n81,
         u4_sub_470_n80, u4_sub_470_n79, u4_sub_470_n78, u4_sub_470_n77,
         u4_sub_470_n76, u4_sub_470_n75, u4_sub_470_n74, u4_sub_470_n73,
         u4_sub_470_n72, u4_sub_470_n71, u4_sub_470_n70, u4_sub_470_n69,
         u4_sub_470_n68, u4_sub_470_n67, u4_sub_470_n66, u4_sub_470_n65,
         u4_sub_470_n64, u4_sub_470_n63, u4_sub_470_n62, u4_sub_470_n61,
         u4_sub_470_n60, u4_sub_470_n59, u4_sub_470_n58, u4_sub_470_n57,
         u4_sub_470_n56, u4_sub_470_n55, u4_sub_470_n54, u4_sub_470_n53,
         u4_sub_470_n52, u4_sub_470_n51, u4_sub_470_n50, u4_sub_470_n49,
         u4_sub_470_n48, u4_sub_470_n47, u4_sub_470_n46, u4_sub_470_n45,
         u4_sub_470_n44, u4_sub_470_n43, u4_sub_470_n42, u4_sub_470_n41,
         u4_sub_470_n40, u4_sub_470_n39, u4_sub_470_n38, u4_sub_470_n37,
         u4_sub_470_n36, u4_sub_470_n35, u4_sub_470_n34, u4_sub_470_n33,
         u4_sub_470_n32, u4_sub_470_n31, u4_sub_470_n30, u4_sub_470_n29,
         u4_sub_470_n28, u4_sub_470_n27, u4_sub_470_n26, u4_sub_470_n25,
         u4_sub_470_n24, u4_sub_470_n23, u4_sub_470_n22, u4_sub_470_n21,
         u4_sub_470_n20, u4_sub_470_n19, u4_sub_470_n18, u4_sub_470_n17,
         u4_sub_470_n16, u4_sub_470_n15, u4_sub_470_n14, u4_sub_470_n13,
         u4_sub_470_n12, u4_sub_470_n11, u4_sub_470_n10, u4_sub_470_n9,
         u4_sub_470_n8, u4_sub_470_n7, u4_sub_470_n6, u4_sub_470_n5,
         u4_sub_470_n4, u4_sub_470_n3, u4_sub_470_n2, u4_sub_470_n1,
         u4_add_464_n23, u4_add_464_n22, u4_add_464_n21, u4_add_464_n20,
         u4_add_464_n19, u4_add_464_n18, u4_add_464_n17, u4_add_464_n16,
         u4_add_464_n15, u4_add_464_n14, u4_add_464_n13, u4_add_464_n12,
         u4_add_464_n11, u4_add_464_n10, u4_add_464_n9, u4_add_464_n8,
         u4_add_464_n7, u4_add_464_n6, u4_add_464_n5, u4_add_464_n4,
         u4_add_464_n3, u4_add_464_n2, u4_add_464_n1, u4_add_396_n173,
         u4_add_396_n172, u4_add_396_n171, u4_add_396_n170, u4_add_396_n169,
         u4_add_396_n168, u4_add_396_n167, u4_add_396_n166, u4_add_396_n165,
         u4_add_396_n164, u4_add_396_n163, u4_add_396_n162, u4_add_396_n161,
         u4_add_396_n160, u4_add_396_n159, u4_add_396_n158, u4_add_396_n157,
         u4_add_396_n156, u4_add_396_n155, u4_add_396_n154, u4_add_396_n153,
         u4_add_396_n152, u4_add_396_n151, u4_add_396_n150, u4_add_396_n149,
         u4_add_396_n148, u4_add_396_n147, u4_add_396_n146, u4_add_396_n145,
         u4_add_396_n144, u4_add_396_n143, u4_add_396_n142, u4_add_396_n141,
         u4_add_396_n140, u4_add_396_n139, u4_add_396_n138, u4_add_396_n137,
         u4_add_396_n136, u4_add_396_n135, u4_add_396_n134, u4_add_396_n133,
         u4_add_396_n132, u4_add_396_n131, u4_add_396_n130, u4_add_396_n129,
         u4_add_396_n128, u4_add_396_n127, u4_add_396_n126, u4_add_396_n125,
         u4_add_396_n124, u4_add_396_n123, u4_add_396_n122, u4_add_396_n121,
         u4_add_396_n120, u4_add_396_n119, u4_add_396_n118, u4_add_396_n117,
         u4_add_396_n116, u4_add_396_n115, u4_add_396_n114, u4_add_396_n113,
         u4_add_396_n112, u4_add_396_n111, u4_add_396_n110, u4_add_396_n109,
         u4_add_396_n108, u4_add_396_n107, u4_add_396_n106, u4_add_396_n105,
         u4_add_396_n104, u4_add_396_n103, u4_add_396_n102, u4_add_396_n101,
         u4_add_396_n100, u4_add_396_n99, u4_add_396_n98, u4_add_396_n97,
         u4_add_396_n96, u4_add_396_n95, u4_add_396_n94, u4_add_396_n93,
         u4_add_396_n92, u4_add_396_n91, u4_add_396_n90, u4_add_396_n89,
         u4_add_396_n88, u4_add_396_n87, u4_add_396_n86, u4_add_396_n85,
         u4_add_396_n84, u4_add_396_n83, u4_add_396_n82, u4_add_396_n81,
         u4_add_396_n80, u4_add_396_n79, u4_add_396_n78, u4_add_396_n77,
         u4_add_396_n76, u4_add_396_n75, u4_add_396_n74, u4_add_396_n73,
         u4_add_396_n72, u4_add_396_n71, u4_add_396_n70, u4_add_396_n69,
         u4_add_396_n68, u4_add_396_n67, u4_add_396_n66, u4_add_396_n65,
         u4_add_396_n64, u4_add_396_n63, u4_add_396_n62, u4_add_396_n61,
         u4_add_396_n60, u4_add_396_n59, u4_add_396_n58, u4_add_396_n57,
         u4_add_396_n56, u4_add_396_n55, u4_add_396_n54, u4_add_396_n53,
         u4_add_396_n52, u4_add_396_n51, u4_add_396_n50, u4_add_396_n49,
         u4_add_396_n48, u4_add_396_n47, u4_add_396_n46, u4_add_396_n45,
         u4_add_396_n44, u4_add_396_n43, u4_add_396_n42, u4_add_396_n41,
         u4_add_396_n40, u4_add_396_n39, u4_add_396_n38, u4_add_396_n37,
         u4_add_396_n36, u4_add_396_n35, u4_add_396_n34, u4_add_396_n33,
         u4_add_396_n32, u4_add_396_n31, u4_add_396_n30, u4_add_396_n29,
         u4_add_396_n28, u4_add_396_n27, u4_add_396_n26, u4_add_396_n25,
         u4_add_396_n24, u4_add_396_n23, u4_add_396_n22, u4_add_396_n21,
         u4_add_396_n20, u4_add_396_n19, u4_add_396_n18, u4_add_396_n17,
         u4_add_396_n16, u4_add_396_n15, u4_add_396_n14, u4_add_396_n13,
         u4_add_396_n12, u4_add_396_n11, u4_add_396_n10, u4_add_396_n9,
         u4_add_396_n8, u4_add_396_n7, u4_add_396_n6, u4_add_396_n5,
         u4_add_396_n4, u4_add_396_n3, u4_add_396_n1, u1_gt_239_n859,
         u1_gt_239_n858, u1_gt_239_n857, u1_gt_239_n856, u1_gt_239_n855,
         u1_gt_239_n854, u1_gt_239_n853, u1_gt_239_n852, u1_gt_239_n851,
         u1_gt_239_n850, u1_gt_239_n849, u1_gt_239_n848, u1_gt_239_n847,
         u1_gt_239_n846, u1_gt_239_n845, u1_gt_239_n844, u1_gt_239_n843,
         u1_gt_239_n842, u1_gt_239_n841, u1_gt_239_n840, u1_gt_239_n839,
         u1_gt_239_n838, u1_gt_239_n837, u1_gt_239_n836, u1_gt_239_n835,
         u1_gt_239_n834, u1_gt_239_n833, u1_gt_239_n832, u1_gt_239_n831,
         u1_gt_239_n830, u1_gt_239_n829, u1_gt_239_n828, u1_gt_239_n827,
         u1_gt_239_n826, u1_gt_239_n825, u1_gt_239_n824, u1_gt_239_n823,
         u1_gt_239_n822, u1_gt_239_n821, u1_gt_239_n820, u1_gt_239_n819,
         u1_gt_239_n818, u1_gt_239_n817, u1_gt_239_n816, u1_gt_239_n815,
         u1_gt_239_n814, u1_gt_239_n813, u1_gt_239_n812, u1_gt_239_n811,
         u1_gt_239_n810, u1_gt_239_n809, u1_gt_239_n808, u1_gt_239_n807,
         u1_gt_239_n806, u1_gt_239_n805, u1_gt_239_n804, u1_gt_239_n803,
         u1_gt_239_n802, u1_gt_239_n801, u1_gt_239_n800, u1_gt_239_n799,
         u1_gt_239_n798, u1_gt_239_n797, u1_gt_239_n796, u1_gt_239_n795,
         u1_gt_239_n794, u1_gt_239_n793, u1_gt_239_n792, u1_gt_239_n791,
         u1_gt_239_n790, u1_gt_239_n789, u1_gt_239_n788, u1_gt_239_n787,
         u1_gt_239_n786, u1_gt_239_n785, u1_gt_239_n784, u1_gt_239_n783,
         u1_gt_239_n782, u1_gt_239_n781, u1_gt_239_n780, u1_gt_239_n779,
         u1_gt_239_n778, u1_gt_239_n777, u1_gt_239_n776, u1_gt_239_n775,
         u1_gt_239_n774, u1_gt_239_n773, u1_gt_239_n772, u1_gt_239_n771,
         u1_gt_239_n770, u1_gt_239_n769, u1_gt_239_n768, u1_gt_239_n767,
         u1_gt_239_n766, u1_gt_239_n765, u1_gt_239_n764, u1_gt_239_n763,
         u1_gt_239_n762, u1_gt_239_n761, u1_gt_239_n760, u1_gt_239_n759,
         u1_gt_239_n758, u1_gt_239_n757, u1_gt_239_n756, u1_gt_239_n755,
         u1_gt_239_n754, u1_gt_239_n753, u1_gt_239_n752, u1_gt_239_n751,
         u1_gt_239_n750, u1_gt_239_n749, u1_gt_239_n748, u1_gt_239_n747,
         u1_gt_239_n746, u1_gt_239_n745, u1_gt_239_n744, u1_gt_239_n743,
         u1_gt_239_n742, u1_gt_239_n741, u1_gt_239_n740, u1_gt_239_n739,
         u1_gt_239_n738, u1_gt_239_n737, u1_gt_239_n736, u1_gt_239_n735,
         u1_gt_239_n734, u1_gt_239_n733, u1_gt_239_n732, u1_gt_239_n731,
         u1_gt_239_n730, u1_gt_239_n729, u1_gt_239_n728, u1_gt_239_n727,
         u1_gt_239_n726, u1_gt_239_n725, u1_gt_239_n724, u1_gt_239_n723,
         u1_gt_239_n722, u1_gt_239_n721, u1_gt_239_n720, u1_gt_239_n719,
         u1_gt_239_n718, u1_gt_239_n717, u1_gt_239_n716, u1_gt_239_n715,
         u1_gt_239_n714, u1_gt_239_n713, u1_gt_239_n712, u1_gt_239_n711,
         u1_gt_239_n710, u1_gt_239_n709, u1_gt_239_n708, u1_gt_239_n707,
         u1_gt_239_n706, u1_gt_239_n705, u1_gt_239_n704, u1_gt_239_n703,
         u1_gt_239_n702, u1_gt_239_n701, u1_gt_239_n700, u1_gt_239_n699,
         u1_gt_239_n698, u1_gt_239_n697, u1_gt_239_n696, u1_gt_239_n695,
         u1_gt_239_n694, u1_gt_239_n693, u1_gt_239_n692, u1_gt_239_n691,
         u1_gt_239_n690, u1_gt_239_n689, u1_gt_239_n688, u1_gt_239_n687,
         u1_gt_239_n686, u1_gt_239_n685, u1_gt_239_n684, u1_gt_239_n683,
         u1_gt_239_n682, u1_gt_239_n681, u1_gt_239_n680, u1_gt_239_n679,
         u1_gt_239_n678, u1_gt_239_n677, u1_gt_239_n676, u1_gt_239_n675,
         u1_gt_239_n674, u1_gt_239_n673, u1_gt_239_n672, u1_gt_239_n671,
         u1_gt_239_n670, u1_gt_239_n669, u1_gt_239_n668, u1_gt_239_n667,
         u1_gt_239_n666, u1_gt_239_n665, u1_gt_239_n664, u1_gt_239_n663,
         u1_gt_239_n662, u1_gt_239_n661, u1_gt_239_n660, u1_gt_239_n659,
         u1_gt_239_n658, u1_gt_239_n657, u1_gt_239_n656, u1_gt_239_n655,
         u1_gt_239_n654, u1_gt_239_n653, u1_gt_239_n652, u1_gt_239_n651,
         u1_gt_239_n650, u1_gt_239_n649, u1_gt_239_n648, u1_gt_239_n647,
         u1_gt_239_n646, u1_gt_239_n645, u1_gt_239_n644, u1_gt_239_n643,
         u1_gt_239_n642, u1_gt_239_n641, u1_gt_239_n640, u1_gt_239_n639,
         u1_gt_239_n638, u1_gt_239_n637, u1_gt_239_n636, u1_gt_239_n635,
         u1_gt_239_n634, u1_gt_239_n633, u1_gt_239_n632, u1_gt_239_n631,
         u1_gt_239_n630, u1_gt_239_n629, u1_gt_239_n628, u1_gt_239_n627,
         u1_gt_239_n626, u1_gt_239_n625, u1_gt_239_n624, u1_gt_239_n623,
         u1_gt_239_n622, u1_gt_239_n621, u1_gt_239_n620, u1_gt_239_n619,
         u1_gt_239_n618, u1_gt_239_n617, u1_gt_239_n616, u1_gt_239_n615,
         u1_gt_239_n614, u1_gt_239_n613, u1_gt_239_n612, u1_gt_239_n611,
         u1_gt_239_n610, u1_gt_239_n609, u1_gt_239_n608, u1_gt_239_n607,
         u1_gt_239_n606, u1_gt_239_n605, u1_gt_239_n604, u1_gt_239_n603,
         u1_gt_239_n602, u1_gt_239_n601, u1_gt_239_n600, u1_gt_239_n599,
         u1_gt_239_n598, u1_gt_239_n597, u1_gt_239_n596, u1_gt_239_n595,
         u1_gt_239_n594, u1_gt_239_n593, u1_gt_239_n592, u1_gt_239_n591,
         u1_gt_239_n590, u1_gt_239_n589, u1_gt_239_n588, u1_gt_239_n587,
         u1_gt_239_n586, u1_gt_239_n585, u1_gt_239_n584, u1_gt_239_n583,
         u1_gt_239_n582, u1_gt_239_n581, u1_gt_239_n580, u1_gt_239_n579,
         u1_gt_239_n578, u1_gt_239_n577, u1_gt_239_n576, u1_gt_239_n575,
         u1_gt_239_n574, u1_gt_239_n573, u1_gt_239_n572, u1_gt_239_n571,
         u1_gt_239_n570, u1_gt_239_n569, u1_gt_239_n568, u1_gt_239_n567,
         u1_gt_239_n566, u1_gt_239_n565, u1_gt_239_n564, u1_gt_239_n563,
         u1_gt_239_n562, u1_gt_239_n561, u1_gt_239_n560, u1_gt_239_n559,
         u1_gt_239_n558, u1_gt_239_n557, u1_gt_239_n556, u1_gt_239_n555,
         u1_gt_239_n554, u1_gt_239_n553, u1_gt_239_n552, u1_gt_239_n551,
         u1_gt_239_n550, u1_gt_239_n549, u1_gt_239_n548, u1_gt_239_n547,
         u1_gt_239_n546, u1_gt_239_n545, u1_gt_239_n544, u1_gt_239_n543,
         u1_gt_239_n542, u1_gt_239_n541, u1_gt_239_n540, u1_gt_239_n539,
         u1_gt_239_n538, u1_gt_239_n537, u1_gt_239_n536, u1_gt_239_n535,
         u1_gt_239_n534, u1_gt_239_n533, u1_gt_239_n532, u1_gt_239_n531,
         u1_gt_239_n530, u1_gt_239_n529, u1_gt_239_n528, u1_gt_239_n527,
         u1_gt_239_n526, u1_gt_239_n525, u1_gt_239_n524, u1_gt_239_n523,
         u1_gt_239_n522, u1_gt_239_n521, u1_gt_239_n520, u1_gt_239_n519,
         u1_gt_239_n518, u1_gt_239_n517, u1_gt_239_n516, u1_gt_239_n515,
         u1_gt_239_n514, u1_gt_239_n513, u1_gt_239_n512, u1_gt_239_n511,
         u1_gt_239_n510, u1_gt_239_n509, u1_gt_239_n508, u1_gt_239_n507,
         u1_gt_239_n506, u1_gt_239_n505, u1_gt_239_n504, u1_gt_239_n503,
         u1_gt_239_n502, u1_gt_239_n501, u1_gt_239_n500, u1_gt_239_n499,
         u1_gt_239_n498, u1_gt_239_n497, u1_gt_239_n496, u1_gt_239_n495,
         u1_gt_239_n494, u1_gt_239_n493, u1_gt_239_n492, u1_gt_239_n491,
         u1_gt_239_n490, u1_gt_239_n489, u1_gt_239_n488, u1_gt_239_n487,
         u1_gt_239_n486, u1_gt_239_n485, u1_gt_239_n484, u1_gt_239_n483,
         u1_gt_239_n482, u1_gt_239_n481, u1_gt_239_n480, u1_gt_239_n479,
         u1_gt_239_n478, u1_gt_239_n477, u1_gt_239_n476, u1_gt_239_n475,
         u1_gt_239_n474, u1_gt_239_n473, u1_gt_239_n472, u1_gt_239_n471,
         u1_gt_239_n470, u1_gt_239_n469, u1_gt_239_n468, u1_gt_239_n467,
         u1_gt_239_n466, u1_gt_239_n465, u1_gt_239_n464, u1_gt_239_n463,
         u1_gt_239_n462, u1_gt_239_n461, u1_gt_239_n460, u1_gt_239_n459,
         u1_gt_239_n458, u1_gt_239_n457, u1_gt_239_n456, u1_gt_239_n455,
         u1_gt_239_n454, u1_gt_239_n453, u1_gt_239_n452, u1_gt_239_n451,
         u1_gt_239_n450, u1_gt_239_n449, u1_gt_239_n448, u1_gt_239_n447,
         u1_gt_239_n446, u1_gt_239_n445, u1_gt_239_n444, u1_gt_239_n443,
         u1_gt_239_n442, u1_gt_239_n441, u1_gt_239_n440, u1_gt_239_n439,
         u1_gt_239_n438, u1_gt_239_n437, u1_gt_239_n436, u1_gt_239_n435,
         u1_gt_239_n434, u1_gt_239_n433, u1_gt_239_n432, u1_gt_239_n431,
         u1_gt_239_n430, u1_gt_239_n429, u1_gt_239_n428, u1_gt_239_n427,
         u1_gt_239_n426, u1_gt_239_n425, u1_gt_239_n424, u1_gt_239_n423,
         u1_gt_239_n422, u1_gt_239_n421, u1_gt_239_n420, u1_gt_239_n419,
         u1_gt_239_n418, u1_gt_239_n417, u1_gt_239_n416, u1_gt_239_n415,
         u1_gt_239_n414, u1_gt_239_n413, u1_gt_239_n412, u1_gt_239_n411,
         u1_gt_239_n410, u1_gt_239_n409, u1_gt_239_n408, u1_gt_239_n407,
         u1_gt_239_n406, u1_gt_239_n405, u1_gt_239_n404, u1_gt_239_n403,
         u1_gt_239_n402, u1_gt_239_n401, u1_gt_239_n400, u1_gt_239_n399,
         u1_gt_239_n398, u1_gt_239_n397, u1_gt_239_n396, u1_gt_239_n395,
         u1_gt_239_n394, u1_gt_239_n393, u1_gt_239_n392, u1_gt_239_n391,
         u1_gt_239_n390, u1_gt_239_n389, u1_gt_239_n388, u1_gt_239_n387,
         u1_gt_239_n386, u1_gt_239_n385, u1_gt_239_n384, u1_gt_239_n383,
         u1_gt_239_n382, u1_gt_239_n381, u1_gt_239_n380, u1_gt_239_n379,
         u1_gt_239_n378, u1_gt_239_n377, u1_gt_239_n376, u1_gt_239_n375,
         u1_gt_239_n374, u1_gt_239_n373, u1_gt_239_n372, u1_gt_239_n371,
         u1_gt_239_n370, u1_gt_239_n369, u1_gt_239_n368, u1_gt_239_n367,
         u1_gt_239_n366, u1_gt_239_n365, u1_gt_239_n364, u1_gt_239_n363,
         u1_gt_239_n362, u1_gt_239_n361, u1_gt_239_n360, u1_gt_239_n359,
         u1_gt_239_n358, u1_gt_239_n357, u1_gt_239_n356, u1_gt_239_n355,
         u1_gt_239_n354, u1_gt_239_n353, u1_gt_239_n352, u1_gt_239_n351,
         u1_gt_239_n350, u1_gt_239_n349, u1_gt_239_n348, u1_gt_239_n347,
         u1_gt_239_n346, u1_gt_239_n345, u1_gt_239_n344, u1_gt_239_n343,
         u1_gt_239_n342, u1_gt_239_n341, u1_gt_239_n340, u1_gt_239_n339,
         u1_gt_239_n338, u1_gt_239_n337, u1_gt_239_n336, u1_gt_239_n335,
         u1_gt_239_n334, u1_gt_239_n333, u1_gt_239_n332, u1_gt_239_n331,
         u1_gt_239_n330, u1_gt_239_n329, u1_gt_239_n328, u1_gt_239_n327,
         u1_gt_239_n326, u1_gt_239_n325, u1_gt_239_n324, u1_gt_239_n323,
         u1_gt_239_n322, u1_gt_239_n321, u1_gt_239_n320, u1_gt_239_n319,
         u1_gt_239_n318, u1_gt_239_n317, u1_gt_239_n316, u1_gt_239_n315,
         u1_gt_239_n314, u1_gt_239_n313, u1_gt_239_n312, u1_gt_239_n311,
         u1_gt_239_n310, u1_gt_239_n309, u1_gt_239_n308, u1_gt_239_n307,
         u1_gt_239_n306, u1_gt_239_n305, u1_gt_239_n304, u1_gt_239_n303,
         u1_gt_239_n302, u1_gt_239_n301, u1_gt_239_n300, u1_gt_239_n299,
         u1_gt_239_n298, u1_gt_239_n297, u1_gt_239_n296, u1_gt_239_n295,
         u1_gt_239_n294, u1_gt_239_n293, u1_gt_239_n292, u1_gt_239_n291,
         u1_gt_239_n290, u1_gt_239_n289, u1_gt_239_n288, u1_gt_239_n287,
         u1_gt_239_n286, u1_gt_239_n285, u1_gt_239_n284, u1_gt_239_n283,
         u1_gt_239_n282, u1_gt_239_n281, u1_gt_239_n280, u1_gt_239_n279,
         u1_gt_239_n278, u1_gt_239_n277, u1_gt_239_n276, u1_gt_239_n275,
         u1_gt_239_n274, u1_gt_239_n273, u1_gt_239_n272, u1_gt_239_n271,
         u1_gt_239_n270, u1_gt_239_n269, u1_gt_239_n268, u1_gt_239_n267,
         u1_gt_239_n266, u1_gt_239_n265, u1_gt_239_n264, u1_gt_239_n263,
         u1_gt_239_n262, u1_gt_239_n261, u1_gt_239_n260, u1_gt_239_n259,
         u1_gt_239_n258, u1_gt_239_n257, u1_gt_239_n256, u1_gt_239_n255,
         u1_gt_239_n254, u1_gt_239_n253, u1_gt_239_n252, u1_gt_239_n251,
         u1_gt_239_n250, u1_gt_239_n249, u1_gt_239_n248, u1_gt_239_n247,
         u1_gt_239_n246, u1_gt_239_n245, u1_gt_239_n244, u1_gt_239_n243,
         u1_gt_239_n242, u1_gt_239_n241, u1_gt_239_n240, u1_gt_239_n239,
         u1_gt_239_n238, u1_gt_239_n237, u1_gt_239_n236, u1_gt_239_n235,
         u1_gt_239_n234, u1_gt_239_n233, u1_gt_239_n232, u1_gt_239_n231,
         u1_gt_239_n230, u1_gt_239_n229, u1_gt_239_n228, u1_gt_239_n227,
         u1_gt_239_n226, u1_gt_239_n225, u1_gt_239_n224, u1_gt_239_n223,
         u1_gt_239_n222, u1_gt_239_n221, u1_gt_239_n220, u1_gt_239_n219,
         u1_gt_239_n218, u1_gt_239_n217, u1_gt_239_n216, u1_gt_239_n215,
         u1_gt_239_n214, u1_gt_239_n213, u1_gt_239_n212, u1_gt_239_n211,
         u1_gt_239_n210, u1_gt_239_n209, u1_gt_239_n208, u1_gt_239_n207,
         u1_gt_239_n206, u1_gt_239_n205, u1_gt_239_n204, u1_gt_239_n203,
         u1_gt_239_n202, u1_gt_239_n201, u1_gt_239_n200, u1_gt_239_n199,
         u1_gt_239_n198, u1_gt_239_n197, u1_gt_239_n196, u1_gt_239_n195,
         u1_gt_239_n194, u1_gt_239_n193, u1_gt_239_n192, u1_gt_239_n191,
         u1_gt_239_n190, u1_gt_239_n189, u1_gt_239_n188, u1_gt_239_n187,
         u1_gt_239_n186, u1_gt_239_n185, u1_gt_239_n184, u1_gt_239_n183,
         u1_gt_239_n182, u1_gt_239_n181, u1_gt_239_n180, u1_gt_239_n179,
         u1_gt_239_n178, u1_gt_239_n177, u1_gt_239_n176, u1_gt_239_n175,
         u1_gt_239_n174, u1_gt_239_n173, u1_gt_239_n172, u1_gt_239_n171,
         u1_gt_239_n170, u1_gt_239_n169, u1_gt_239_n168, u1_gt_239_n167,
         u1_gt_239_n166, u1_gt_239_n165, u1_gt_239_n164, u1_gt_239_n163,
         u1_gt_239_n162, u1_gt_239_n161, u1_gt_239_n160, u1_gt_239_n159,
         u1_gt_239_n158, u1_gt_239_n157, u1_gt_239_n156, u1_gt_239_n155,
         u1_gt_239_n154, u1_gt_239_n153, u1_gt_239_n152, u1_gt_239_n151,
         u1_gt_239_n150, u1_gt_239_n149, u1_gt_239_n148, u1_gt_239_n147,
         u1_gt_239_n146, u1_gt_239_n145, u1_gt_239_n144, u1_gt_239_n143,
         u1_gt_239_n142, u1_gt_239_n141, u1_gt_239_n140, u1_gt_239_n139,
         u1_gt_239_n138, u1_gt_239_n137, u1_gt_239_n136, u1_gt_239_n135,
         u1_gt_239_n134, u1_gt_239_n133, u1_gt_239_n132, u1_gt_239_n131,
         u1_gt_239_n130, u1_gt_239_n129, u1_gt_239_n128, u1_gt_239_n127,
         u1_gt_239_n126, u1_gt_239_n125, u1_gt_239_n124, u1_gt_239_n123,
         u1_gt_239_n122, u1_gt_239_n121, u1_gt_239_n120, u1_gt_239_n119,
         u1_gt_239_n118, u1_gt_239_n117, u1_gt_239_n116, u1_gt_239_n115,
         u1_gt_239_n114, u1_gt_239_n113, u1_gt_239_n112, u1_gt_239_n111,
         u1_gt_239_n110, u1_gt_239_n109, u1_gt_239_n108, u1_gt_239_n107,
         u1_gt_239_n106, u1_gt_239_n105, u1_gt_239_n104, u1_gt_239_n103,
         u1_gt_239_n102, u1_gt_239_n101, u1_gt_239_n100, u1_gt_239_n99,
         u1_gt_239_n98, u1_gt_239_n97, u1_gt_239_n96, u1_gt_239_n95,
         u1_gt_239_n94, u1_gt_239_n93, u1_gt_239_n92, u1_gt_239_n91,
         u1_gt_239_n90, u1_gt_239_n89, u1_gt_239_n88, u1_gt_239_n87,
         u1_gt_239_n86, u1_gt_239_n85, u1_gt_239_n84, u1_gt_239_n83,
         u1_gt_239_n82, u1_gt_239_n81, u1_gt_239_n80, u1_gt_239_n79,
         u1_gt_239_n78, u1_gt_239_n77, u1_gt_239_n76, u1_gt_239_n75,
         u1_gt_239_n74, u1_gt_239_n73, u1_gt_239_n72, u1_gt_239_n71,
         u1_gt_239_n70, u1_gt_239_n69, u1_gt_239_n68, u1_gt_239_n67,
         u1_gt_239_n66, u1_gt_239_n65, u1_gt_239_n64, u1_gt_239_n63,
         u1_gt_239_n62, u1_gt_239_n61, u1_gt_239_n60, u1_gt_239_n59,
         u1_gt_239_n58, u1_gt_239_n57, u1_gt_239_n56, u1_gt_239_n55,
         u1_gt_239_n54, u1_gt_239_n53, u1_gt_239_n52, u1_gt_239_n51,
         u1_gt_239_n50, u1_gt_239_n49, u1_gt_239_n48, u1_gt_239_n47,
         u1_gt_239_n46, u1_gt_239_n45, u1_gt_239_n44, u1_gt_239_n43,
         u1_gt_239_n42, u1_gt_239_n41, u1_gt_239_n40, u1_gt_239_n39,
         u1_gt_239_n38, u1_gt_239_n37, u1_gt_239_n36, u1_gt_239_n35,
         u1_gt_239_n34, u1_gt_239_n33, u1_gt_239_n32, u1_gt_239_n31,
         u1_gt_239_n30, u1_gt_239_n29, u1_gt_239_n28, u1_gt_239_n27,
         u1_gt_239_n26, u1_gt_239_n25, u1_gt_239_n24, u1_gt_239_n23,
         u1_gt_239_n22, u1_gt_239_n21, u1_gt_239_n20, u1_gt_239_n19,
         u1_gt_239_n18, u1_gt_239_n17, u1_gt_239_n16, u1_gt_239_n15,
         u1_gt_239_n14, u1_gt_239_n13, u1_gt_239_n12, u1_gt_239_n11,
         u1_gt_239_n10, u1_gt_239_n9, u1_gt_239_n8, u1_gt_239_n7, u1_gt_239_n6,
         u1_gt_239_n5, u1_gt_239_n4, u1_gt_239_n3, u1_gt_239_n2, u1_gt_239_n1,
         u4_sub_496_n52, u4_sub_496_n51, u4_sub_496_n50, u4_sub_496_n49,
         u4_sub_496_n48, u4_sub_496_n47, u4_sub_496_n46, u4_sub_496_n45,
         u4_sub_496_n44, u4_sub_496_n43, u4_sub_496_n42, u4_sub_496_n41,
         u4_sub_496_n40, u4_sub_496_n39, u4_sub_496_n38, u4_sub_496_n37,
         u4_sub_496_n36, u4_sub_496_n35, u4_sub_496_n34, u4_sub_496_n33,
         u4_sub_496_n32, u4_sub_496_n31, u4_sub_496_n30, u4_sub_496_n29,
         u4_sub_496_n28, u4_sub_496_n27, u4_sub_496_n26, u4_sub_496_n25,
         u4_sub_496_n24, u4_sub_496_n23, u4_sub_496_n22, u4_sub_496_n21,
         u4_sub_496_n20, u4_sub_496_n19, u4_sub_496_n18, u4_sub_496_n17,
         u4_sub_496_n16, u4_sub_496_n15, u4_sub_496_n14, u4_sub_496_n13,
         u4_sub_496_n12, u4_sub_496_n11, u4_sub_496_n10, u4_sub_496_n9,
         u4_sub_496_n8, u4_sub_496_n7, u4_sub_496_n6, u4_sub_496_n5,
         u4_sub_496_n4, u4_sub_496_n3, u4_sub_496_n2, u4_sub_496_n1,
         u4_sub_496_net61381, u4_sub_496_net61382, u4_sub_496_net61383,
         u4_sub_496_net61374, u4_sub_496_net61376, u4_sub_496_net61379,
         u4_sub_496_net61359, u4_sub_496_net61372, u4_sub_496_net61347,
         u4_sub_496_net61349, u4_sub_496_net61352, u4_sub_496_net61354,
         u4_sub_496_net61355, u4_sub_496_net61358, u4_sub_496_net61360,
         u4_sub_496_net61363, u4_sub_496_net61364, u4_sub_496_net61365,
         u4_sub_496_net61368, u4_sub_496_net61369, u4_sub_496_net61370,
         u4_sub_496_net61385, u4_sub_496_net61386, u4_sub_496_net61387,
         u4_sub_496_net61389, u4_sub_496_net61411, u4_sub_496_net61429,
         u4_sub_496_net61430, u4_sub_496_net61437, u4_sub_496_net61438,
         u4_sll_454_n233, u4_sll_454_n232, u4_sll_454_n231, u4_sll_454_n230,
         u4_sll_454_n229, u4_sll_454_n228, u4_sll_454_n227, u4_sll_454_n226,
         u4_sll_454_n225, u4_sll_454_n224, u4_sll_454_n223, u4_sll_454_n222,
         u4_sll_454_n221, u4_sll_454_n220, u4_sll_454_n219, u4_sll_454_n218,
         u4_sll_454_n217, u4_sll_454_n216, u4_sll_454_n215, u4_sll_454_n214,
         u4_sll_454_n213, u4_sll_454_n212, u4_sll_454_n211, u4_sll_454_n210,
         u4_sll_454_n209, u4_sll_454_n208, u4_sll_454_n207, u4_sll_454_n206,
         u4_sll_454_n205, u4_sll_454_n204, u4_sll_454_n203, u4_sll_454_n202,
         u4_sll_454_n201, u4_sll_454_n200, u4_sll_454_n199, u4_sll_454_n198,
         u4_sll_454_n197, u4_sll_454_n196, u4_sll_454_n195, u4_sll_454_n194,
         u4_sll_454_n193, u4_sll_454_n192, u4_sll_454_n191, u4_sll_454_n190,
         u4_sll_454_n189, u4_sll_454_n188, u4_sll_454_n187, u4_sll_454_n186,
         u4_sll_454_n185, u4_sll_454_n184, u4_sll_454_n183, u4_sll_454_n182,
         u4_sll_454_n181, u4_sll_454_n180, u4_sll_454_n179, u4_sll_454_n178,
         u4_sll_454_n177, u4_sll_454_n176, u4_sll_454_n175, u4_sll_454_n174,
         u4_sll_454_n173, u4_sll_454_n172, u4_sll_454_n171, u4_sll_454_n170,
         u4_sll_454_n169, u4_sll_454_n168, u4_sll_454_n167, u4_sll_454_n166,
         u4_sll_454_n165, u4_sll_454_n164, u4_sll_454_n163, u4_sll_454_n162,
         u4_sll_454_n161, u4_sll_454_n160, u4_sll_454_n159, u4_sll_454_n158,
         u4_sll_454_n157, u4_sll_454_n156, u4_sll_454_n155, u4_sll_454_n154,
         u4_sll_454_n153, u4_sll_454_n152, u4_sll_454_n151, u4_sll_454_n150,
         u4_sll_454_n149, u4_sll_454_n148, u4_sll_454_n147, u4_sll_454_n146,
         u4_sll_454_n145, u4_sll_454_n144, u4_sll_454_n143, u4_sll_454_n142,
         u4_sll_454_n141, u4_sll_454_n140, u4_sll_454_n139, u4_sll_454_n138,
         u4_sll_454_n137, u4_sll_454_n136, u4_sll_454_n135, u4_sll_454_n134,
         u4_sll_454_n133, u4_sll_454_n132, u4_sll_454_n131, u4_sll_454_n130,
         u4_sll_454_n129, u4_sll_454_n128, u4_sll_454_n127, u4_sll_454_n126,
         u4_sll_454_n125, u4_sll_454_n124, u4_sll_454_n123, u4_sll_454_n122,
         u4_sll_454_n121, u4_sll_454_n120, u4_sll_454_n119, u4_sll_454_n118,
         u4_sll_454_n117, u4_sll_454_n116, u4_sll_454_n115, u4_sll_454_n114,
         u4_sll_454_n113, u4_sll_454_n112, u4_sll_454_n111, u4_sll_454_n110,
         u4_sll_454_n109, u4_sll_454_n108, u4_sll_454_n107, u4_sll_454_n106,
         u4_sll_454_n105, u4_sll_454_n104, u4_sll_454_n103, u4_sll_454_n102,
         u4_sll_454_n101, u4_sll_454_n100, u4_sll_454_n99, u4_sll_454_n98,
         u4_sll_454_n97, u4_sll_454_n96, u4_sll_454_n95, u4_sll_454_n94,
         u4_sll_454_n93, u4_sll_454_n92, u4_sll_454_n91, u4_sll_454_n90,
         u4_sll_454_n89, u4_sll_454_n88, u4_sll_454_n87, u4_sll_454_n86,
         u4_sll_454_n85, u4_sll_454_n84, u4_sll_454_n83, u4_sll_454_n82,
         u4_sll_454_n81, u4_sll_454_n80, u4_sll_454_n79, u4_sll_454_n78,
         u4_sll_454_n77, u4_sll_454_n76, u4_sll_454_n75, u4_sll_454_n74,
         u4_sll_454_n73, u4_sll_454_n72, u4_sll_454_n71, u4_sll_454_n70,
         u4_sll_454_n69, u4_sll_454_n68, u4_sll_454_n67, u4_sll_454_n66,
         u4_sll_454_n65, u4_sll_454_n64, u4_sll_454_n63, u4_sll_454_n62,
         u4_sll_454_n61, u4_sll_454_n60, u4_sll_454_n59, u4_sll_454_n58,
         u4_sll_454_n57, u4_sll_454_n56, u4_sll_454_n55, u4_sll_454_n54,
         u4_sll_454_n53, u4_sll_454_n52, u4_sll_454_n51, u4_sll_454_n50,
         u4_sll_454_n49, u4_sll_454_n48, u4_sll_454_n47, u4_sll_454_n46,
         u4_sll_454_n45, u4_sll_454_n44, u4_sll_454_n43, u4_sll_454_n42,
         u4_sll_454_n41, u4_sll_454_n40, u4_sll_454_n39, u4_sll_454_n38,
         u4_sll_454_n37, u4_sll_454_n36, u4_sll_454_n35, u4_sll_454_n34,
         u4_sll_454_n33, u4_sll_454_n32, u4_sll_454_n31, u4_sll_454_n30,
         u4_sll_454_n29, u4_sll_454_n28, u4_sll_454_n27, u4_sll_454_n26,
         u4_sll_454_n25, u4_sll_454_n24, u4_sll_454_n23, u4_sll_454_n22,
         u4_sll_454_n21, u4_sll_454_n20, u4_sll_454_n19, u4_sll_454_n18,
         u4_sll_454_n17, u4_sll_454_n16, u4_sll_454_n15, u4_sll_454_n14,
         u4_sll_454_n13, u4_sll_454_n12, u4_sll_454_n11, u4_sll_454_n10,
         u4_sll_454_n9, u4_sll_454_n8, u4_sll_454_n7, u4_sll_454_n6,
         u4_sll_454_n5, u4_sll_454_n4, u4_sll_454_n3, u4_sll_454_n2,
         u4_sll_454_n1, u4_sll_454__UDW__90155_net73403,
         u4_sll_454_ML_int_6__44_, u4_sll_454_ML_int_7__44_,
         u4_sll_454_SHMAG_5_, u4_sll_454_net61033, u4_sll_454_net66509,
         u4_sll_454_net66537, u4_sll_454__UDW__90347_net74043,
         u4_sll_454_ML_int_5__44_, u4_sll_454_net66565,
         u4_sll_454_ML_int_2__20_, u4_sll_454_ML_int_3__20_,
         u4_sll_454_SHMAG_2_, u4_sll_454_net66697, u4_sll_454_net66701,
         u4_sll_454_net66705, u4_sll_454_net66757, u4_sll_454_ML_int_3__28_,
         u4_sll_454_ML_int_4__28_, u4_sll_454_SHMAG_3_, u4_sll_454_net66621,
         u4_sll_454_net66649, u4_sll_454_net66677, u4_sll_454_ML_int_4__44_,
         u4_sll_454_SHMAG_4_, u4_sll_454_net66585, u4_sll_454_net66589,
         u4_sll_454_net66593, u4_sll_454_ML_int_1__16_,
         u4_sll_454_ML_int_2__16_, u4_sll_454_SHMAG_1_, u4_sll_454_net61034,
         u4_sll_454_net61036, u4_sll_454_net61037, u4_sll_454_net63277,
         u4_sll_454_net66761, u4_sll_454_ML_int_1__14_, u4_sll_454_net61028,
         u4_sll_454_net66379, u4_sll_454_net66383, u4_sll_454_net66387,
         u4_sll_454_temp_int_SH_0_, u4_sll_454__UDW__90011_net72923,
         u4_sll_454__UDW__89963_net72763, u4_sll_454__UDW__89915_net72603,
         u4_sll_454_net66711, u4_sll_454_net66715, u4_sll_454_net66717,
         u4_sll_454_net66719, u4_sll_454_net66721, u4_sll_454_net66723,
         u4_sll_454_net66727, u4_sll_454_net66733, u4_sll_454_net66655,
         u4_sll_454_net66659, u4_sll_454_net66661, u4_sll_454_net66663,
         u4_sll_454_net66667, u4_sll_454_net66673, u4_sll_454_net66675,
         u4_sll_454_net66699, u4_sll_454_net66647, u4_sll_454_net66599,
         u4_sll_454_net66601, u4_sll_454_net66603, u4_sll_454_net66607,
         u4_sll_454_net66609, u4_sll_454_net66611, u4_sll_454_net66613,
         u4_sll_454_net66619, u4_sll_454_net66591, u4_sll_454_net66545,
         u4_sll_454_net66547, u4_sll_454_net66549, u4_sll_454_net66551,
         u4_sll_454_net66555, u4_sll_454_net66557, u4_sll_454_net66563,
         u4_sll_454_net66485, u4_sll_454_net66487, u4_sll_454_net66489,
         u4_sll_454_net66491, u4_sll_454_net66493, u4_sll_454_net66495,
         u4_sll_454_net66497, u4_sll_454_net66499, u4_sll_454_net66501,
         u4_sll_454_net66481, u4_sll_454_net66429, u4_sll_454_net66431,
         u4_sll_454_net66433, u4_sll_454_net66435, u4_sll_454_net66439,
         u4_sll_454_net66441, u4_sll_454_net66443, u4_sll_454_net66445,
         u4_sll_454_net66451, u4_sll_454_net66455, u4_sll_454_net66385,
         u4_sll_454_net66357, u4_sll_454_net66359, u4_sll_454_net66361,
         u4_sll_454_net66363, u4_sll_454_net66365, u4_sll_454_net66367,
         u4_sll_454_net66369, u4_sll_454_net66371, u4_sll_454_net66373,
         u4_sll_454_net66377, u4_sll_454_net63259, u4_sll_454_net63261,
         u4_sll_454_net63265, u4_sll_454_net63267, u4_sll_454_net63269,
         u4_sll_454_net63271, u4_sll_454_net63273, u4_sll_454_net61030,
         u4_sll_454_net61032, u4_sll_454_ML_int_7__0_, u4_sll_454_ML_int_7__1_,
         u4_sll_454_ML_int_7__2_, u4_sll_454_ML_int_7__3_,
         u4_sll_454_ML_int_7__4_, u4_sll_454_ML_int_7__5_,
         u4_sll_454_ML_int_7__6_, u4_sll_454_ML_int_7__7_,
         u4_sll_454_ML_int_7__8_, u4_sll_454_ML_int_7__9_,
         u4_sll_454_ML_int_7__10_, u4_sll_454_ML_int_7__11_,
         u4_sll_454_ML_int_7__12_, u4_sll_454_ML_int_7__13_,
         u4_sll_454_ML_int_7__14_, u4_sll_454_ML_int_7__15_,
         u4_sll_454_ML_int_7__16_, u4_sll_454_ML_int_7__17_,
         u4_sll_454_ML_int_7__18_, u4_sll_454_ML_int_7__19_,
         u4_sll_454_ML_int_7__20_, u4_sll_454_ML_int_7__21_,
         u4_sll_454_ML_int_7__22_, u4_sll_454_ML_int_7__23_,
         u4_sll_454_ML_int_7__24_, u4_sll_454_ML_int_7__25_,
         u4_sll_454_ML_int_7__26_, u4_sll_454_ML_int_7__27_,
         u4_sll_454_ML_int_7__28_, u4_sll_454_ML_int_7__29_,
         u4_sll_454_ML_int_7__30_, u4_sll_454_ML_int_7__31_,
         u4_sll_454_ML_int_7__32_, u4_sll_454_ML_int_7__33_,
         u4_sll_454_ML_int_7__34_, u4_sll_454_ML_int_7__35_,
         u4_sll_454_ML_int_7__36_, u4_sll_454_ML_int_7__37_,
         u4_sll_454_ML_int_7__38_, u4_sll_454_ML_int_7__39_,
         u4_sll_454_ML_int_7__40_, u4_sll_454_ML_int_7__41_,
         u4_sll_454_ML_int_7__42_, u4_sll_454_ML_int_7__43_,
         u4_sll_454_ML_int_7__45_, u4_sll_454_ML_int_7__46_,
         u4_sll_454_ML_int_7__47_, u4_sll_454_ML_int_7__48_,
         u4_sll_454_ML_int_7__49_, u4_sll_454_ML_int_7__50_,
         u4_sll_454_ML_int_7__51_, u4_sll_454_ML_int_7__52_,
         u4_sll_454_ML_int_7__53_, u4_sll_454_ML_int_7__54_,
         u4_sll_454_ML_int_7__55_, u4_sll_454_ML_int_7__56_,
         u4_sll_454_ML_int_7__57_, u4_sll_454_ML_int_7__58_,
         u4_sll_454_ML_int_7__59_, u4_sll_454_ML_int_7__60_,
         u4_sll_454_ML_int_7__61_, u4_sll_454_ML_int_7__62_,
         u4_sll_454_ML_int_7__63_, u4_sll_454_ML_int_7__64_,
         u4_sll_454_ML_int_7__65_, u4_sll_454_ML_int_7__66_,
         u4_sll_454_ML_int_7__67_, u4_sll_454_ML_int_7__68_,
         u4_sll_454_ML_int_7__69_, u4_sll_454_ML_int_7__70_,
         u4_sll_454_ML_int_7__71_, u4_sll_454_ML_int_7__72_,
         u4_sll_454_ML_int_7__73_, u4_sll_454_ML_int_7__74_,
         u4_sll_454_ML_int_7__75_, u4_sll_454_ML_int_7__76_,
         u4_sll_454_ML_int_7__77_, u4_sll_454_ML_int_7__78_,
         u4_sll_454_ML_int_7__79_, u4_sll_454_ML_int_7__80_,
         u4_sll_454_ML_int_7__81_, u4_sll_454_ML_int_7__82_,
         u4_sll_454_ML_int_7__83_, u4_sll_454_ML_int_7__84_,
         u4_sll_454_ML_int_7__85_, u4_sll_454_ML_int_7__86_,
         u4_sll_454_ML_int_7__87_, u4_sll_454_ML_int_7__88_,
         u4_sll_454_ML_int_7__89_, u4_sll_454_ML_int_7__90_,
         u4_sll_454_ML_int_7__91_, u4_sll_454_ML_int_7__92_,
         u4_sll_454_ML_int_7__93_, u4_sll_454_ML_int_7__94_,
         u4_sll_454_ML_int_7__95_, u4_sll_454_ML_int_7__96_,
         u4_sll_454_ML_int_7__97_, u4_sll_454_ML_int_7__98_,
         u4_sll_454_ML_int_7__99_, u4_sll_454_ML_int_7__100_,
         u4_sll_454_ML_int_7__101_, u4_sll_454_ML_int_7__102_,
         u4_sll_454_ML_int_7__103_, u4_sll_454_ML_int_7__104_,
         u4_sll_454_ML_int_7__105_, u4_sll_454_ML_int_6__0_,
         u4_sll_454_ML_int_6__1_, u4_sll_454_ML_int_6__2_,
         u4_sll_454_ML_int_6__3_, u4_sll_454_ML_int_6__4_,
         u4_sll_454_ML_int_6__5_, u4_sll_454_ML_int_6__6_,
         u4_sll_454_ML_int_6__7_, u4_sll_454_ML_int_6__8_,
         u4_sll_454_ML_int_6__9_, u4_sll_454_ML_int_6__10_,
         u4_sll_454_ML_int_6__11_, u4_sll_454_ML_int_6__12_,
         u4_sll_454_ML_int_6__13_, u4_sll_454_ML_int_6__14_,
         u4_sll_454_ML_int_6__15_, u4_sll_454_ML_int_6__16_,
         u4_sll_454_ML_int_6__17_, u4_sll_454_ML_int_6__18_,
         u4_sll_454_ML_int_6__19_, u4_sll_454_ML_int_6__20_,
         u4_sll_454_ML_int_6__21_, u4_sll_454_ML_int_6__22_,
         u4_sll_454_ML_int_6__23_, u4_sll_454_ML_int_6__24_,
         u4_sll_454_ML_int_6__25_, u4_sll_454_ML_int_6__26_,
         u4_sll_454_ML_int_6__27_, u4_sll_454_ML_int_6__28_,
         u4_sll_454_ML_int_6__29_, u4_sll_454_ML_int_6__30_,
         u4_sll_454_ML_int_6__31_, u4_sll_454_ML_int_6__32_,
         u4_sll_454_ML_int_6__33_, u4_sll_454_ML_int_6__34_,
         u4_sll_454_ML_int_6__35_, u4_sll_454_ML_int_6__36_,
         u4_sll_454_ML_int_6__37_, u4_sll_454_ML_int_6__38_,
         u4_sll_454_ML_int_6__39_, u4_sll_454_ML_int_6__40_,
         u4_sll_454_ML_int_6__41_, u4_sll_454_ML_int_6__42_,
         u4_sll_454_ML_int_6__43_, u4_sll_454_ML_int_6__45_,
         u4_sll_454_ML_int_6__46_, u4_sll_454_ML_int_6__47_,
         u4_sll_454_ML_int_6__48_, u4_sll_454_ML_int_6__49_,
         u4_sll_454_ML_int_6__50_, u4_sll_454_ML_int_6__51_,
         u4_sll_454_ML_int_6__52_, u4_sll_454_ML_int_6__53_,
         u4_sll_454_ML_int_6__54_, u4_sll_454_ML_int_6__55_,
         u4_sll_454_ML_int_6__56_, u4_sll_454_ML_int_6__57_,
         u4_sll_454_ML_int_6__58_, u4_sll_454_ML_int_6__59_,
         u4_sll_454_ML_int_6__60_, u4_sll_454_ML_int_6__61_,
         u4_sll_454_ML_int_6__62_, u4_sll_454_ML_int_6__63_,
         u4_sll_454_ML_int_6__64_, u4_sll_454_ML_int_6__65_,
         u4_sll_454_ML_int_6__66_, u4_sll_454_ML_int_6__67_,
         u4_sll_454_ML_int_6__68_, u4_sll_454_ML_int_6__69_,
         u4_sll_454_ML_int_6__70_, u4_sll_454_ML_int_6__71_,
         u4_sll_454_ML_int_6__72_, u4_sll_454_ML_int_6__73_,
         u4_sll_454_ML_int_6__74_, u4_sll_454_ML_int_6__75_,
         u4_sll_454_ML_int_6__76_, u4_sll_454_ML_int_6__77_,
         u4_sll_454_ML_int_6__78_, u4_sll_454_ML_int_6__79_,
         u4_sll_454_ML_int_6__80_, u4_sll_454_ML_int_6__81_,
         u4_sll_454_ML_int_6__82_, u4_sll_454_ML_int_6__83_,
         u4_sll_454_ML_int_6__84_, u4_sll_454_ML_int_6__85_,
         u4_sll_454_ML_int_6__86_, u4_sll_454_ML_int_6__87_,
         u4_sll_454_ML_int_6__88_, u4_sll_454_ML_int_6__89_,
         u4_sll_454_ML_int_6__90_, u4_sll_454_ML_int_6__91_,
         u4_sll_454_ML_int_6__92_, u4_sll_454_ML_int_6__93_,
         u4_sll_454_ML_int_6__94_, u4_sll_454_ML_int_6__95_,
         u4_sll_454_ML_int_6__96_, u4_sll_454_ML_int_6__97_,
         u4_sll_454_ML_int_6__98_, u4_sll_454_ML_int_6__99_,
         u4_sll_454_ML_int_6__100_, u4_sll_454_ML_int_6__101_,
         u4_sll_454_ML_int_6__102_, u4_sll_454_ML_int_6__103_,
         u4_sll_454_ML_int_6__104_, u4_sll_454_ML_int_6__105_,
         u4_sll_454_ML_int_5__0_, u4_sll_454_ML_int_5__1_,
         u4_sll_454_ML_int_5__2_, u4_sll_454_ML_int_5__3_,
         u4_sll_454_ML_int_5__4_, u4_sll_454_ML_int_5__5_,
         u4_sll_454_ML_int_5__6_, u4_sll_454_ML_int_5__7_,
         u4_sll_454_ML_int_5__8_, u4_sll_454_ML_int_5__9_,
         u4_sll_454_ML_int_5__10_, u4_sll_454_ML_int_5__11_,
         u4_sll_454_ML_int_5__12_, u4_sll_454_ML_int_5__13_,
         u4_sll_454_ML_int_5__14_, u4_sll_454_ML_int_5__15_,
         u4_sll_454_ML_int_5__16_, u4_sll_454_ML_int_5__17_,
         u4_sll_454_ML_int_5__18_, u4_sll_454_ML_int_5__19_,
         u4_sll_454_ML_int_5__20_, u4_sll_454_ML_int_5__21_,
         u4_sll_454_ML_int_5__22_, u4_sll_454_ML_int_5__23_,
         u4_sll_454_ML_int_5__24_, u4_sll_454_ML_int_5__25_,
         u4_sll_454_ML_int_5__26_, u4_sll_454_ML_int_5__27_,
         u4_sll_454_ML_int_5__28_, u4_sll_454_ML_int_5__29_,
         u4_sll_454_ML_int_5__30_, u4_sll_454_ML_int_5__31_,
         u4_sll_454_ML_int_5__32_, u4_sll_454_ML_int_5__33_,
         u4_sll_454_ML_int_5__34_, u4_sll_454_ML_int_5__35_,
         u4_sll_454_ML_int_5__36_, u4_sll_454_ML_int_5__37_,
         u4_sll_454_ML_int_5__38_, u4_sll_454_ML_int_5__39_,
         u4_sll_454_ML_int_5__40_, u4_sll_454_ML_int_5__41_,
         u4_sll_454_ML_int_5__42_, u4_sll_454_ML_int_5__43_,
         u4_sll_454_ML_int_5__45_, u4_sll_454_ML_int_5__46_,
         u4_sll_454_ML_int_5__47_, u4_sll_454_ML_int_5__48_,
         u4_sll_454_ML_int_5__49_, u4_sll_454_ML_int_5__50_,
         u4_sll_454_ML_int_5__51_, u4_sll_454_ML_int_5__52_,
         u4_sll_454_ML_int_5__53_, u4_sll_454_ML_int_5__54_,
         u4_sll_454_ML_int_5__55_, u4_sll_454_ML_int_5__56_,
         u4_sll_454_ML_int_5__57_, u4_sll_454_ML_int_5__58_,
         u4_sll_454_ML_int_5__59_, u4_sll_454_ML_int_5__60_,
         u4_sll_454_ML_int_5__61_, u4_sll_454_ML_int_5__62_,
         u4_sll_454_ML_int_5__63_, u4_sll_454_ML_int_5__64_,
         u4_sll_454_ML_int_5__65_, u4_sll_454_ML_int_5__66_,
         u4_sll_454_ML_int_5__67_, u4_sll_454_ML_int_5__68_,
         u4_sll_454_ML_int_5__69_, u4_sll_454_ML_int_5__70_,
         u4_sll_454_ML_int_5__71_, u4_sll_454_ML_int_5__72_,
         u4_sll_454_ML_int_5__73_, u4_sll_454_ML_int_5__74_,
         u4_sll_454_ML_int_5__75_, u4_sll_454_ML_int_5__76_,
         u4_sll_454_ML_int_5__77_, u4_sll_454_ML_int_5__78_,
         u4_sll_454_ML_int_5__79_, u4_sll_454_ML_int_5__80_,
         u4_sll_454_ML_int_5__81_, u4_sll_454_ML_int_5__82_,
         u4_sll_454_ML_int_5__83_, u4_sll_454_ML_int_5__84_,
         u4_sll_454_ML_int_5__85_, u4_sll_454_ML_int_5__86_,
         u4_sll_454_ML_int_5__87_, u4_sll_454_ML_int_5__88_,
         u4_sll_454_ML_int_5__89_, u4_sll_454_ML_int_5__90_,
         u4_sll_454_ML_int_5__91_, u4_sll_454_ML_int_5__92_,
         u4_sll_454_ML_int_5__93_, u4_sll_454_ML_int_5__94_,
         u4_sll_454_ML_int_5__95_, u4_sll_454_ML_int_5__96_,
         u4_sll_454_ML_int_5__97_, u4_sll_454_ML_int_5__98_,
         u4_sll_454_ML_int_5__99_, u4_sll_454_ML_int_5__100_,
         u4_sll_454_ML_int_5__101_, u4_sll_454_ML_int_5__102_,
         u4_sll_454_ML_int_5__103_, u4_sll_454_ML_int_5__104_,
         u4_sll_454_ML_int_5__105_, u4_sll_454_ML_int_4__0_,
         u4_sll_454_ML_int_4__1_, u4_sll_454_ML_int_4__2_,
         u4_sll_454_ML_int_4__3_, u4_sll_454_ML_int_4__4_,
         u4_sll_454_ML_int_4__5_, u4_sll_454_ML_int_4__6_,
         u4_sll_454_ML_int_4__7_, u4_sll_454_ML_int_4__8_,
         u4_sll_454_ML_int_4__9_, u4_sll_454_ML_int_4__10_,
         u4_sll_454_ML_int_4__11_, u4_sll_454_ML_int_4__12_,
         u4_sll_454_ML_int_4__13_, u4_sll_454_ML_int_4__14_,
         u4_sll_454_ML_int_4__15_, u4_sll_454_ML_int_4__16_,
         u4_sll_454_ML_int_4__17_, u4_sll_454_ML_int_4__18_,
         u4_sll_454_ML_int_4__19_, u4_sll_454_ML_int_4__20_,
         u4_sll_454_ML_int_4__21_, u4_sll_454_ML_int_4__22_,
         u4_sll_454_ML_int_4__23_, u4_sll_454_ML_int_4__24_,
         u4_sll_454_ML_int_4__25_, u4_sll_454_ML_int_4__26_,
         u4_sll_454_ML_int_4__27_, u4_sll_454_ML_int_4__29_,
         u4_sll_454_ML_int_4__30_, u4_sll_454_ML_int_4__31_,
         u4_sll_454_ML_int_4__32_, u4_sll_454_ML_int_4__33_,
         u4_sll_454_ML_int_4__34_, u4_sll_454_ML_int_4__35_,
         u4_sll_454_ML_int_4__36_, u4_sll_454_ML_int_4__37_,
         u4_sll_454_ML_int_4__38_, u4_sll_454_ML_int_4__39_,
         u4_sll_454_ML_int_4__40_, u4_sll_454_ML_int_4__41_,
         u4_sll_454_ML_int_4__42_, u4_sll_454_ML_int_4__43_,
         u4_sll_454_ML_int_4__45_, u4_sll_454_ML_int_4__46_,
         u4_sll_454_ML_int_4__47_, u4_sll_454_ML_int_4__48_,
         u4_sll_454_ML_int_4__49_, u4_sll_454_ML_int_4__50_,
         u4_sll_454_ML_int_4__51_, u4_sll_454_ML_int_4__52_,
         u4_sll_454_ML_int_4__53_, u4_sll_454_ML_int_4__54_,
         u4_sll_454_ML_int_4__55_, u4_sll_454_ML_int_4__56_,
         u4_sll_454_ML_int_4__57_, u4_sll_454_ML_int_4__58_,
         u4_sll_454_ML_int_4__59_, u4_sll_454_ML_int_4__60_,
         u4_sll_454_ML_int_4__61_, u4_sll_454_ML_int_4__62_,
         u4_sll_454_ML_int_4__63_, u4_sll_454_ML_int_4__64_,
         u4_sll_454_ML_int_4__65_, u4_sll_454_ML_int_4__66_,
         u4_sll_454_ML_int_4__67_, u4_sll_454_ML_int_4__68_,
         u4_sll_454_ML_int_4__69_, u4_sll_454_ML_int_4__70_,
         u4_sll_454_ML_int_4__71_, u4_sll_454_ML_int_4__72_,
         u4_sll_454_ML_int_4__73_, u4_sll_454_ML_int_4__74_,
         u4_sll_454_ML_int_4__75_, u4_sll_454_ML_int_4__76_,
         u4_sll_454_ML_int_4__77_, u4_sll_454_ML_int_4__78_,
         u4_sll_454_ML_int_4__79_, u4_sll_454_ML_int_4__80_,
         u4_sll_454_ML_int_4__81_, u4_sll_454_ML_int_4__82_,
         u4_sll_454_ML_int_4__83_, u4_sll_454_ML_int_4__84_,
         u4_sll_454_ML_int_4__85_, u4_sll_454_ML_int_4__86_,
         u4_sll_454_ML_int_4__87_, u4_sll_454_ML_int_4__88_,
         u4_sll_454_ML_int_4__89_, u4_sll_454_ML_int_4__90_,
         u4_sll_454_ML_int_4__91_, u4_sll_454_ML_int_4__92_,
         u4_sll_454_ML_int_4__93_, u4_sll_454_ML_int_4__94_,
         u4_sll_454_ML_int_4__95_, u4_sll_454_ML_int_4__96_,
         u4_sll_454_ML_int_4__97_, u4_sll_454_ML_int_4__98_,
         u4_sll_454_ML_int_4__99_, u4_sll_454_ML_int_4__100_,
         u4_sll_454_ML_int_4__101_, u4_sll_454_ML_int_4__102_,
         u4_sll_454_ML_int_4__103_, u4_sll_454_ML_int_4__104_,
         u4_sll_454_ML_int_4__105_, u4_sll_454_ML_int_3__0_,
         u4_sll_454_ML_int_3__1_, u4_sll_454_ML_int_3__2_,
         u4_sll_454_ML_int_3__3_, u4_sll_454_ML_int_3__4_,
         u4_sll_454_ML_int_3__5_, u4_sll_454_ML_int_3__6_,
         u4_sll_454_ML_int_3__7_, u4_sll_454_ML_int_3__8_,
         u4_sll_454_ML_int_3__9_, u4_sll_454_ML_int_3__10_,
         u4_sll_454_ML_int_3__11_, u4_sll_454_ML_int_3__12_,
         u4_sll_454_ML_int_3__13_, u4_sll_454_ML_int_3__14_,
         u4_sll_454_ML_int_3__15_, u4_sll_454_ML_int_3__16_,
         u4_sll_454_ML_int_3__17_, u4_sll_454_ML_int_3__18_,
         u4_sll_454_ML_int_3__19_, u4_sll_454_ML_int_3__21_,
         u4_sll_454_ML_int_3__22_, u4_sll_454_ML_int_3__23_,
         u4_sll_454_ML_int_3__24_, u4_sll_454_ML_int_3__25_,
         u4_sll_454_ML_int_3__26_, u4_sll_454_ML_int_3__27_,
         u4_sll_454_ML_int_3__29_, u4_sll_454_ML_int_3__30_,
         u4_sll_454_ML_int_3__31_, u4_sll_454_ML_int_3__32_,
         u4_sll_454_ML_int_3__33_, u4_sll_454_ML_int_3__34_,
         u4_sll_454_ML_int_3__35_, u4_sll_454_ML_int_3__36_,
         u4_sll_454_ML_int_3__37_, u4_sll_454_ML_int_3__38_,
         u4_sll_454_ML_int_3__39_, u4_sll_454_ML_int_3__40_,
         u4_sll_454_ML_int_3__41_, u4_sll_454_ML_int_3__42_,
         u4_sll_454_ML_int_3__43_, u4_sll_454_ML_int_3__44_,
         u4_sll_454_ML_int_3__45_, u4_sll_454_ML_int_3__46_,
         u4_sll_454_ML_int_3__47_, u4_sll_454_ML_int_3__48_,
         u4_sll_454_ML_int_3__49_, u4_sll_454_ML_int_3__50_,
         u4_sll_454_ML_int_3__51_, u4_sll_454_ML_int_3__52_,
         u4_sll_454_ML_int_3__53_, u4_sll_454_ML_int_3__54_,
         u4_sll_454_ML_int_3__55_, u4_sll_454_ML_int_3__56_,
         u4_sll_454_ML_int_3__57_, u4_sll_454_ML_int_3__58_,
         u4_sll_454_ML_int_3__59_, u4_sll_454_ML_int_3__60_,
         u4_sll_454_ML_int_3__61_, u4_sll_454_ML_int_3__62_,
         u4_sll_454_ML_int_3__63_, u4_sll_454_ML_int_3__64_,
         u4_sll_454_ML_int_3__65_, u4_sll_454_ML_int_3__66_,
         u4_sll_454_ML_int_3__67_, u4_sll_454_ML_int_3__68_,
         u4_sll_454_ML_int_3__69_, u4_sll_454_ML_int_3__70_,
         u4_sll_454_ML_int_3__71_, u4_sll_454_ML_int_3__72_,
         u4_sll_454_ML_int_3__73_, u4_sll_454_ML_int_3__74_,
         u4_sll_454_ML_int_3__75_, u4_sll_454_ML_int_3__76_,
         u4_sll_454_ML_int_3__77_, u4_sll_454_ML_int_3__78_,
         u4_sll_454_ML_int_3__79_, u4_sll_454_ML_int_3__80_,
         u4_sll_454_ML_int_3__81_, u4_sll_454_ML_int_3__82_,
         u4_sll_454_ML_int_3__83_, u4_sll_454_ML_int_3__84_,
         u4_sll_454_ML_int_3__85_, u4_sll_454_ML_int_3__86_,
         u4_sll_454_ML_int_3__87_, u4_sll_454_ML_int_3__88_,
         u4_sll_454_ML_int_3__89_, u4_sll_454_ML_int_3__90_,
         u4_sll_454_ML_int_3__91_, u4_sll_454_ML_int_3__92_,
         u4_sll_454_ML_int_3__93_, u4_sll_454_ML_int_3__94_,
         u4_sll_454_ML_int_3__95_, u4_sll_454_ML_int_3__96_,
         u4_sll_454_ML_int_3__97_, u4_sll_454_ML_int_3__98_,
         u4_sll_454_ML_int_3__99_, u4_sll_454_ML_int_3__100_,
         u4_sll_454_ML_int_3__101_, u4_sll_454_ML_int_3__102_,
         u4_sll_454_ML_int_3__103_, u4_sll_454_ML_int_3__104_,
         u4_sll_454_ML_int_3__105_, u4_sll_454_ML_int_2__0_,
         u4_sll_454_ML_int_2__1_, u4_sll_454_ML_int_2__2_,
         u4_sll_454_ML_int_2__3_, u4_sll_454_ML_int_2__4_,
         u4_sll_454_ML_int_2__5_, u4_sll_454_ML_int_2__6_,
         u4_sll_454_ML_int_2__7_, u4_sll_454_ML_int_2__8_,
         u4_sll_454_ML_int_2__9_, u4_sll_454_ML_int_2__10_,
         u4_sll_454_ML_int_2__11_, u4_sll_454_ML_int_2__12_,
         u4_sll_454_ML_int_2__13_, u4_sll_454_ML_int_2__14_,
         u4_sll_454_ML_int_2__15_, u4_sll_454_ML_int_2__17_,
         u4_sll_454_ML_int_2__18_, u4_sll_454_ML_int_2__19_,
         u4_sll_454_ML_int_2__21_, u4_sll_454_ML_int_2__22_,
         u4_sll_454_ML_int_2__23_, u4_sll_454_ML_int_2__24_,
         u4_sll_454_ML_int_2__25_, u4_sll_454_ML_int_2__26_,
         u4_sll_454_ML_int_2__27_, u4_sll_454_ML_int_2__28_,
         u4_sll_454_ML_int_2__29_, u4_sll_454_ML_int_2__30_,
         u4_sll_454_ML_int_2__31_, u4_sll_454_ML_int_2__32_,
         u4_sll_454_ML_int_2__33_, u4_sll_454_ML_int_2__34_,
         u4_sll_454_ML_int_2__35_, u4_sll_454_ML_int_2__36_,
         u4_sll_454_ML_int_2__37_, u4_sll_454_ML_int_2__38_,
         u4_sll_454_ML_int_2__39_, u4_sll_454_ML_int_2__40_,
         u4_sll_454_ML_int_2__41_, u4_sll_454_ML_int_2__42_,
         u4_sll_454_ML_int_2__43_, u4_sll_454_ML_int_2__44_,
         u4_sll_454_ML_int_2__45_, u4_sll_454_ML_int_2__46_,
         u4_sll_454_ML_int_2__47_, u4_sll_454_ML_int_2__48_,
         u4_sll_454_ML_int_2__49_, u4_sll_454_ML_int_2__50_,
         u4_sll_454_ML_int_2__51_, u4_sll_454_ML_int_2__52_,
         u4_sll_454_ML_int_2__53_, u4_sll_454_ML_int_2__54_,
         u4_sll_454_ML_int_2__55_, u4_sll_454_ML_int_2__56_,
         u4_sll_454_ML_int_2__57_, u4_sll_454_ML_int_2__58_,
         u4_sll_454_ML_int_2__59_, u4_sll_454_ML_int_2__60_,
         u4_sll_454_ML_int_2__61_, u4_sll_454_ML_int_2__62_,
         u4_sll_454_ML_int_2__63_, u4_sll_454_ML_int_2__64_,
         u4_sll_454_ML_int_2__65_, u4_sll_454_ML_int_2__66_,
         u4_sll_454_ML_int_2__67_, u4_sll_454_ML_int_2__68_,
         u4_sll_454_ML_int_2__69_, u4_sll_454_ML_int_2__70_,
         u4_sll_454_ML_int_2__71_, u4_sll_454_ML_int_2__72_,
         u4_sll_454_ML_int_2__73_, u4_sll_454_ML_int_2__74_,
         u4_sll_454_ML_int_2__75_, u4_sll_454_ML_int_2__76_,
         u4_sll_454_ML_int_2__77_, u4_sll_454_ML_int_2__78_,
         u4_sll_454_ML_int_2__79_, u4_sll_454_ML_int_2__80_,
         u4_sll_454_ML_int_2__81_, u4_sll_454_ML_int_2__82_,
         u4_sll_454_ML_int_2__83_, u4_sll_454_ML_int_2__84_,
         u4_sll_454_ML_int_2__85_, u4_sll_454_ML_int_2__86_,
         u4_sll_454_ML_int_2__87_, u4_sll_454_ML_int_2__88_,
         u4_sll_454_ML_int_2__89_, u4_sll_454_ML_int_2__90_,
         u4_sll_454_ML_int_2__91_, u4_sll_454_ML_int_2__92_,
         u4_sll_454_ML_int_2__93_, u4_sll_454_ML_int_2__94_,
         u4_sll_454_ML_int_2__95_, u4_sll_454_ML_int_2__96_,
         u4_sll_454_ML_int_2__97_, u4_sll_454_ML_int_2__98_,
         u4_sll_454_ML_int_2__99_, u4_sll_454_ML_int_2__100_,
         u4_sll_454_ML_int_2__101_, u4_sll_454_ML_int_2__102_,
         u4_sll_454_ML_int_2__103_, u4_sll_454_ML_int_2__104_,
         u4_sll_454_ML_int_2__105_, u4_sll_454_ML_int_1__0_,
         u4_sll_454_ML_int_1__1_, u4_sll_454_ML_int_1__2_,
         u4_sll_454_ML_int_1__3_, u4_sll_454_ML_int_1__4_,
         u4_sll_454_ML_int_1__5_, u4_sll_454_ML_int_1__6_,
         u4_sll_454_ML_int_1__7_, u4_sll_454_ML_int_1__8_,
         u4_sll_454_ML_int_1__9_, u4_sll_454_ML_int_1__10_,
         u4_sll_454_ML_int_1__11_, u4_sll_454_ML_int_1__12_,
         u4_sll_454_ML_int_1__13_, u4_sll_454_ML_int_1__15_,
         u4_sll_454_ML_int_1__17_, u4_sll_454_ML_int_1__18_,
         u4_sll_454_ML_int_1__19_, u4_sll_454_ML_int_1__20_,
         u4_sll_454_ML_int_1__21_, u4_sll_454_ML_int_1__22_,
         u4_sll_454_ML_int_1__23_, u4_sll_454_ML_int_1__24_,
         u4_sll_454_ML_int_1__25_, u4_sll_454_ML_int_1__26_,
         u4_sll_454_ML_int_1__27_, u4_sll_454_ML_int_1__28_,
         u4_sll_454_ML_int_1__29_, u4_sll_454_ML_int_1__30_,
         u4_sll_454_ML_int_1__31_, u4_sll_454_ML_int_1__32_,
         u4_sll_454_ML_int_1__33_, u4_sll_454_ML_int_1__34_,
         u4_sll_454_ML_int_1__35_, u4_sll_454_ML_int_1__36_,
         u4_sll_454_ML_int_1__37_, u4_sll_454_ML_int_1__38_,
         u4_sll_454_ML_int_1__39_, u4_sll_454_ML_int_1__40_,
         u4_sll_454_ML_int_1__41_, u4_sll_454_ML_int_1__42_,
         u4_sll_454_ML_int_1__43_, u4_sll_454_ML_int_1__44_,
         u4_sll_454_ML_int_1__45_, u4_sll_454_ML_int_1__46_,
         u4_sll_454_ML_int_1__47_, u4_sll_454_ML_int_1__48_,
         u4_sll_454_ML_int_1__49_, u4_sll_454_ML_int_1__50_,
         u4_sll_454_ML_int_1__51_, u4_sll_454_ML_int_1__52_,
         u4_sll_454_ML_int_1__53_, u4_sll_454_ML_int_1__54_,
         u4_sll_454_ML_int_1__55_, u4_sll_454_ML_int_1__56_,
         u4_sll_454_ML_int_1__57_, u4_sll_454_ML_int_1__58_,
         u4_sll_454_ML_int_1__59_, u4_sll_454_ML_int_1__60_,
         u4_sll_454_ML_int_1__61_, u4_sll_454_ML_int_1__62_,
         u4_sll_454_ML_int_1__63_, u4_sll_454_ML_int_1__64_,
         u4_sll_454_ML_int_1__65_, u4_sll_454_ML_int_1__66_,
         u4_sll_454_ML_int_1__67_, u4_sll_454_ML_int_1__68_,
         u4_sll_454_ML_int_1__69_, u4_sll_454_ML_int_1__70_,
         u4_sll_454_ML_int_1__71_, u4_sll_454_ML_int_1__72_,
         u4_sll_454_ML_int_1__73_, u4_sll_454_ML_int_1__74_,
         u4_sll_454_ML_int_1__75_, u4_sll_454_ML_int_1__76_,
         u4_sll_454_ML_int_1__77_, u4_sll_454_ML_int_1__78_,
         u4_sll_454_ML_int_1__79_, u4_sll_454_ML_int_1__80_,
         u4_sll_454_ML_int_1__81_, u4_sll_454_ML_int_1__82_,
         u4_sll_454_ML_int_1__83_, u4_sll_454_ML_int_1__84_,
         u4_sll_454_ML_int_1__85_, u4_sll_454_ML_int_1__86_,
         u4_sll_454_ML_int_1__87_, u4_sll_454_ML_int_1__88_,
         u4_sll_454_ML_int_1__89_, u4_sll_454_ML_int_1__90_,
         u4_sll_454_ML_int_1__91_, u4_sll_454_ML_int_1__92_,
         u4_sll_454_ML_int_1__93_, u4_sll_454_ML_int_1__94_,
         u4_sll_454_ML_int_1__95_, u4_sll_454_ML_int_1__96_,
         u4_sll_454_ML_int_1__97_, u4_sll_454_ML_int_1__98_,
         u4_sll_454_ML_int_1__99_, u4_sll_454_ML_int_1__100_,
         u4_sll_454_ML_int_1__101_, u4_sll_454_ML_int_1__102_,
         u4_sll_454_ML_int_1__103_, u4_sll_454_ML_int_1__104_,
         u4_sll_454_ML_int_1__105_, u4_sll_454_SHMAG_6_;
  wire   [63:52] opa_r;
  wire   [63:52] opb_r;
  wire   [1:0] rmode_r1;
  wire   [1:0] rmode_r2;
  wire   [1:0] rmode_r3;
  wire   [2:0] fpu_op_r1;
  wire   [2:0] fpu_op_r2;
  wire   [1:0] fpu_op_r3;
  wire   [55:0] fracta;
  wire   [55:0] fractb;
  wire   [10:0] exp_fasu;
  wire   [51:0] fracta_mul;
  wire   [7:2] exp_mul;
  wire   [1:0] exp_ovf;
  wire   [2:0] underflow_fmul_d;
  wire   [56:0] fract_out_q;
  wire   [105:0] prod;
  wire   [4:0] div_opa_ldz_d;
  wire   [107:0] quo;
  wire   [107:0] remainder;
  wire   [4:0] div_opa_ldz_r1;
  wire   [4:0] div_opa_ldz_r2;
  wire   [9:3] exp_r;
  wire   [59:1] opa_r1;
  wire   [104:0] fract_i2f;
  wire   [104:50] fract_denorm;
  wire   [2:0] underflow_fmul_r;
  wire   [55:0] u1_fractb_s;
  wire   [55:0] u1_fracta_s;
  wire   [10:0] u1_exp_diff2;
  wire   [10:0] u1_exp_small;
  wire   [2:1] u2_underflow_d;
  wire   [105:0] u5_prod1;
  wire   [107:0] u6_remainder;
  wire   [107:0] u6_quo1;
  wire   [10:0] u4_div_exp3;
  wire   [10:0] u4_exp_fix_divb;
  wire   [10:0] u4_exp_fix_diva;
  wire   [6:2] u4_fi_ldz_mi22;
  wire   [8:0] u4_shift_left;
  wire   [10:0] u4_shift_right;
  wire   [6:5] u4_sll_482_SHMAG;
  wire   [10:2] u4_add_466_carry;
  wire   [56:1] u3_sub_63_carry;
  wire   [55:1] u3_add_63_carry;
  wire   [10:2] u2_add_120_carry;
  wire   [10:2] u2_add_118_carry;
  wire   [10:1] u2_add_115_carry;
  wire   [11:1] u2_sub_115_carry;
  wire   [10:1] sub_1_root_u1_sub_133_aco_carry;
  wire   [102:54] u5_mult_82_CLA_SUM;
  wire   [103:53] u5_mult_82_CLA_CARRY;

  OR2_X2 u4_C19042 ( .A1(u4_N6462), .A2(u4_exp_out_0_), .ZN(u4_N6463) );
  OR2_X2 u4_C19043 ( .A1(u4_N6461), .A2(u4_exp_out_1_), .ZN(u4_N6462) );
  OR2_X2 u4_C19044 ( .A1(u4_N6460), .A2(u4_exp_out_2_), .ZN(u4_N6461) );
  OR2_X2 u4_C19045 ( .A1(u4_N6459), .A2(u4_exp_out_3_), .ZN(u4_N6460) );
  OR2_X2 u4_C19048 ( .A1(u4_N6456), .A2(u4_exp_out_6_), .ZN(u4_N6457) );
  OR2_X2 u4_C19049 ( .A1(u4_N6455), .A2(u4_exp_out_7_), .ZN(u4_N6456) );
  OR2_X2 u4_C19050 ( .A1(u4_N6454), .A2(u4_exp_out_8_), .ZN(u4_N6455) );
  OR2_X2 u4_C19051 ( .A1(u4_exp_out_10_), .A2(u4_exp_out_9_), .ZN(u4_N6454) );
  OR2_X2 u4_C19471 ( .A1(u4_shift_right[10]), .A2(u4_shift_right[9]), .ZN(
        u4_N5904) );
  OR2_X2 u4_C19733 ( .A1(net45067), .A2(u4_N6916), .ZN(u4_N6917) );
  AND2_X2 u4_C19735 ( .A1(u4_exp_out_10_), .A2(1'b1), .ZN(u4_N6916) );
  NOR2_X4 U17 ( .A1(net63221), .A2(n2399), .ZN(n2404) );
  AOI22_X2 U18 ( .A1(u4_exp_f2i_1_108_), .A2(1'b0), .B1(net45055), .B2(
        u4_exp_out1_1_), .ZN(n2402) );
  OAI221_X2 U19 ( .B1(n7206), .B2(n2408), .C1(n8244), .C2(net63287), .A(n2409), 
        .ZN(u4_exp_out_2_) );
  OAI221_X2 U21 ( .B1(n7205), .B2(n2408), .C1(net34242), .C2(net63289), .A(
        n2412), .ZN(u4_exp_out_3_) );
  OAI221_X2 U23 ( .B1(n7204), .B2(n2408), .C1(net34243), .C2(net63287), .A(
        n2415), .ZN(u4_exp_out_4_) );
  OAI221_X2 U25 ( .B1(net44770), .B2(n2408), .C1(net34244), .C2(net63287), .A(
        n2417), .ZN(u4_exp_out_5_) );
  OAI221_X2 U27 ( .B1(n7203), .B2(n2408), .C1(n8243), .C2(net63287), .A(n2419), 
        .ZN(u4_exp_out_6_) );
  OAI221_X2 U29 ( .B1(n7202), .B2(n2408), .C1(n8242), .C2(net63287), .A(n2421), 
        .ZN(u4_exp_out_7_) );
  OAI221_X2 U32 ( .B1(n7201), .B2(n2408), .C1(n7199), .C2(net63287), .A(1'b1), 
        .ZN(u4_exp_out_8_) );
  OAI211_X2 U131 ( .C1(net45071), .C2(n2442), .A(n2476), .B(n2477), .ZN(
        u4_shift_right[0]) );
  AND2_X2 U448 ( .A1(opb_r[63]), .A2(opa_r[63]), .ZN(u2_N121) );
  AOI221_X2 U856 ( .B1(opb_nan), .B2(n3063), .C1(n3064), .C2(
        u1_fracta_lt_fractb), .A(u1_signa_r), .ZN(n3060) );
  NAND2_X2 U858 ( .A1(opa_nan), .A2(opb_nan), .ZN(n3063) );
  OAI22_X2 U859 ( .A1(n4493), .A2(n3065), .B1(n3066), .B2(n3067), .ZN(u1_N218)
         );
  XOR2_X2 U860 ( .A(u1_signb_r), .B(u1_add_r), .Z(n3067) );
  AND2_X2 U861 ( .A1(n3065), .A2(n4493), .ZN(n3066) );
  AOI22_X2 U862 ( .A1(u0_snan_r_a), .A2(u0_expa_ff), .B1(u0_snan_r_b), .B2(
        u0_expb_ff), .ZN(n3068) );
  AOI22_X2 U863 ( .A1(u0_qnan_r_a), .A2(u0_expa_ff), .B1(u0_qnan_r_b), .B2(
        u0_expb_ff), .ZN(n3069) );
  NAND2_X2 U864 ( .A1(n3070), .A2(n3071), .ZN(u0_N7) );
  AND2_X2 U868 ( .A1(u0_fractb_00), .A2(u0_expb_00), .ZN(u0_N17) );
  AND2_X2 U869 ( .A1(u0_fracta_00), .A2(u0_expa_00), .ZN(u0_N16) );
  NAND2_X2 U870 ( .A1(u0_infb_f_r), .A2(u0_expb_ff), .ZN(n3070) );
  NAND2_X2 U871 ( .A1(u0_infa_f_r), .A2(u0_expa_ff), .ZN(n3071) );
  OR3_X2 U909 ( .A1(u6_N50), .A2(u6_N5), .A3(u6_N4), .ZN(n3110) );
  OR4_X2 U910 ( .A1(u6_N6), .A2(u6_N7), .A3(u6_N8), .A4(u6_N9), .ZN(n3109) );
  NOR4_X2 U1131 ( .A1(n3293), .A2(n3294), .A3(n4492), .A4(n4359), .ZN(N923) );
  NAND4_X2 U1133 ( .A1(exp_mul[3]), .A2(exp_mul[2]), .A3(exp_mul[4]), .A4(
        n3295), .ZN(n3293) );
  NOR4_X2 U1160 ( .A1(n3358), .A2(prod[21]), .A3(prod[23]), .A4(prod[22]), 
        .ZN(n3357) );
  OR4_X2 U1161 ( .A1(prod[24]), .A2(prod[25]), .A3(prod[26]), .A4(prod[27]), 
        .ZN(n3358) );
  NOR4_X2 U1162 ( .A1(n3359), .A2(prod[16]), .A3(prod[18]), .A4(prod[17]), 
        .ZN(n3356) );
  OR3_X2 U1163 ( .A1(prod[1]), .A2(prod[20]), .A3(prod[19]), .ZN(n3359) );
  NOR4_X2 U1164 ( .A1(n3360), .A2(prod[105]), .A3(prod[11]), .A4(prod[10]), 
        .ZN(n3355) );
  OR4_X2 U1165 ( .A1(prod[12]), .A2(prod[13]), .A3(prod[14]), .A4(prod[15]), 
        .ZN(n3360) );
  NOR4_X2 U1169 ( .A1(n3366), .A2(prod[46]), .A3(prod[48]), .A4(prod[47]), 
        .ZN(n3365) );
  OR4_X2 U1170 ( .A1(prod[49]), .A2(prod[4]), .A3(prod[50]), .A4(prod[51]), 
        .ZN(n3366) );
  NOR4_X2 U1171 ( .A1(n3367), .A2(prod[3]), .A3(prod[41]), .A4(prod[40]), .ZN(
        n3364) );
  OR4_X2 U1172 ( .A1(prod[42]), .A2(prod[43]), .A3(prod[44]), .A4(prod[45]), 
        .ZN(n3367) );
  NOR4_X2 U1173 ( .A1(n3368), .A2(prod[33]), .A3(prod[35]), .A4(prod[34]), 
        .ZN(n3363) );
  OR4_X2 U1174 ( .A1(prod[36]), .A2(prod[37]), .A3(prod[38]), .A4(prod[39]), 
        .ZN(n3368) );
  NOR4_X2 U1175 ( .A1(n3369), .A2(prod[28]), .A3(prod[2]), .A4(prod[29]), .ZN(
        n3362) );
  OR3_X2 U1176 ( .A1(prod[31]), .A2(prod[32]), .A3(prod[30]), .ZN(n3369) );
  NOR4_X2 U1187 ( .A1(n3382), .A2(prod[94]), .A3(prod[96]), .A4(prod[95]), 
        .ZN(n3381) );
  OR4_X2 U1188 ( .A1(prod[97]), .A2(prod[98]), .A3(prod[99]), .A4(prod[9]), 
        .ZN(n3382) );
  NOR4_X2 U1193 ( .A1(n3385), .A2(prod[76]), .A3(prod[78]), .A4(prod[77]), 
        .ZN(n3378) );
  OR3_X2 U1194 ( .A1(prod[7]), .A2(prod[80]), .A3(prod[79]), .ZN(n3385) );
  AOI22_X2 U1762 ( .A1(u4_N5998), .A2(net63325), .B1(u4_N6106), .B2(net63343), 
        .ZN(n3650) );
  AOI22_X2 U1764 ( .A1(u4_N5996), .A2(net63325), .B1(u4_N6104), .B2(net63343), 
        .ZN(n3654) );
  AOI22_X2 U1766 ( .A1(u4_N5995), .A2(net63325), .B1(u4_N6103), .B2(net63343), 
        .ZN(n2528) );
  AOI22_X2 U1767 ( .A1(u4_N5994), .A2(net63325), .B1(u4_N6102), .B2(net63343), 
        .ZN(n2529) );
  AOI22_X2 U1771 ( .A1(u4_N6001), .A2(net63325), .B1(u4_N6109), .B2(net63343), 
        .ZN(n3644) );
  AOI22_X2 U1773 ( .A1(u4_N6002), .A2(net63325), .B1(u4_N6110), .B2(net63343), 
        .ZN(n3641) );
  AOI22_X2 U1775 ( .A1(u4_N6003), .A2(net63323), .B1(u4_N6111), .B2(net63341), 
        .ZN(n3638) );
  AOI22_X2 U1777 ( .A1(u4_N6004), .A2(net63323), .B1(u4_N6112), .B2(net63341), 
        .ZN(n3636) );
  AOI22_X2 U1778 ( .A1(u4_N5999), .A2(net63323), .B1(u4_N6107), .B2(net63341), 
        .ZN(n2527) );
  AOI22_X2 U1779 ( .A1(u4_N6000), .A2(net63323), .B1(u4_N6108), .B2(net63341), 
        .ZN(n2525) );
  AOI22_X2 U1780 ( .A1(u4_N5963), .A2(net63323), .B1(u4_N6071), .B2(net63341), 
        .ZN(n2526) );
  AOI22_X2 U1784 ( .A1(u4_N6009), .A2(net63323), .B1(u4_N6117), .B2(net63341), 
        .ZN(n3626) );
  AOI22_X2 U1786 ( .A1(u4_N5964), .A2(net63323), .B1(u4_N6072), .B2(net63341), 
        .ZN(n3720) );
  AOI22_X2 U1788 ( .A1(u4_N6008), .A2(net63323), .B1(u4_N6116), .B2(net63341), 
        .ZN(n3629) );
  AOI22_X2 U1789 ( .A1(u4_N6005), .A2(net63323), .B1(u4_N6113), .B2(net63341), 
        .ZN(n2524) );
  AOI22_X2 U1790 ( .A1(u4_N6007), .A2(net63323), .B1(u4_N6115), .B2(net63341), 
        .ZN(n2522) );
  AOI22_X2 U1791 ( .A1(u4_N6006), .A2(net63323), .B1(u4_N6114), .B2(net63341), 
        .ZN(n2523) );
  NAND4_X2 U1792 ( .A1(n2520), .A2(n2519), .A3(n2521), .A4(n3897), .ZN(n3888)
         );
  AOI22_X2 U1795 ( .A1(u4_N5966), .A2(net63321), .B1(u4_N6074), .B2(net63339), 
        .ZN(n3717) );
  AOI22_X2 U1797 ( .A1(u4_N5967), .A2(net63321), .B1(u4_N6075), .B2(net63339), 
        .ZN(n3715) );
  AOI22_X2 U1799 ( .A1(u4_N5968), .A2(net63321), .B1(u4_N6076), .B2(net63339), 
        .ZN(n3712) );
  AOI22_X2 U1801 ( .A1(u4_N5969), .A2(net63321), .B1(u4_N6077), .B2(net63339), 
        .ZN(n3709) );
  AOI22_X2 U1802 ( .A1(u4_N6010), .A2(net63321), .B1(u4_N6118), .B2(net63339), 
        .ZN(n2521) );
  AOI22_X2 U1803 ( .A1(u4_N5965), .A2(net63321), .B1(u4_N6073), .B2(net63339), 
        .ZN(n2519) );
  AOI22_X2 U1809 ( .A1(u4_N5973), .A2(net63321), .B1(u4_N6081), .B2(net63339), 
        .ZN(n3702) );
  AOI22_X2 U1811 ( .A1(u4_N5974), .A2(net63321), .B1(u4_N6082), .B2(net63339), 
        .ZN(n3699) );
  AOI22_X2 U1814 ( .A1(u4_N5960), .A2(net63321), .B1(u4_N6068), .B2(net63339), 
        .ZN(n3731) );
  AOI22_X2 U1815 ( .A1(u4_N5971), .A2(net63321), .B1(u4_N6079), .B2(net63339), 
        .ZN(n2540) );
  AOI22_X2 U1820 ( .A1(u4_N5978), .A2(net63319), .B1(u4_N6086), .B2(net63335), 
        .ZN(n3691) );
  AOI22_X2 U1822 ( .A1(u4_N5979), .A2(net63319), .B1(u4_N6087), .B2(net63335), 
        .ZN(n3689) );
  AOI22_X2 U1824 ( .A1(u4_N5961), .A2(net63319), .B1(u4_N6069), .B2(net63335), 
        .ZN(n3727) );
  AOI22_X2 U1826 ( .A1(u4_N5980), .A2(net63319), .B1(u4_N6088), .B2(net63335), 
        .ZN(n3687) );
  AOI22_X2 U1827 ( .A1(u4_N5975), .A2(net63319), .B1(u4_N6083), .B2(net63335), 
        .ZN(n2539) );
  AOI22_X2 U1828 ( .A1(u4_N5977), .A2(net63319), .B1(u4_N6085), .B2(net63335), 
        .ZN(n2537) );
  AOI22_X2 U1829 ( .A1(u4_N5976), .A2(net63319), .B1(u4_N6084), .B2(net63335), 
        .ZN(n2538) );
  AOI22_X2 U1833 ( .A1(u4_N5985), .A2(net63319), .B1(u4_N6093), .B2(net63335), 
        .ZN(n3677) );
  AOI22_X2 U1835 ( .A1(u4_N5986), .A2(net63319), .B1(u4_N6094), .B2(net63335), 
        .ZN(n3675) );
  AOI22_X2 U1837 ( .A1(u4_N5984), .A2(net63319), .B1(u4_N6092), .B2(net63335), 
        .ZN(n3679) );
  AOI22_X2 U1838 ( .A1(u4_N5981), .A2(net63317), .B1(u4_N6089), .B2(net63335), 
        .ZN(n2536) );
  AOI22_X2 U1839 ( .A1(u4_N5983), .A2(net63317), .B1(u4_N6091), .B2(net63335), 
        .ZN(n2534) );
  AOI22_X2 U1840 ( .A1(u4_N5982), .A2(net63317), .B1(u4_N6090), .B2(net63335), 
        .ZN(n2535) );
  AOI22_X2 U1844 ( .A1(u4_N5962), .A2(net63317), .B1(u4_N6070), .B2(net63335), 
        .ZN(n3724) );
  AOI22_X2 U1846 ( .A1(u4_N5990), .A2(net63317), .B1(u4_N6098), .B2(net63335), 
        .ZN(n3666) );
  AOI22_X2 U1848 ( .A1(u4_N5991), .A2(net63317), .B1(u4_N6099), .B2(net63335), 
        .ZN(n3664) );
  AOI22_X2 U1850 ( .A1(u4_N5992), .A2(net63317), .B1(u4_N6100), .B2(net63335), 
        .ZN(n3662) );
  AOI22_X2 U1852 ( .A1(u4_N5989), .A2(net63317), .B1(u4_N6097), .B2(net63335), 
        .ZN(n2531) );
  AOI22_X2 U1853 ( .A1(u4_N5988), .A2(net63317), .B1(u4_N6096), .B2(net63335), 
        .ZN(n2532) );
  AOI22_X2 U1911 ( .A1(u4_N5959), .A2(net63317), .B1(u4_N6067), .B2(net63335), 
        .ZN(n3865) );
  XOR2_X2 U2330 ( .A(n3065), .B(n7196), .Z(N789) );
  NAND2_X2 U2331 ( .A1(rmode_r2[1]), .A2(rmode_r2[0]), .ZN(n3065) );
  OAI221_X2 U2455 ( .B1(n8510), .B2(n4349), .C1(n4490), .C2(n3296), .A(n4253), 
        .ZN(N337) );
  NAND2_X2 U2456 ( .A1(exp_fasu[10]), .A2(n4254), .ZN(n4253) );
  OAI221_X2 U2457 ( .B1(n8510), .B2(n4444), .C1(n4359), .C2(n3296), .A(n4255), 
        .ZN(N336) );
  NAND2_X2 U2458 ( .A1(exp_fasu[9]), .A2(n4254), .ZN(n4255) );
  OAI221_X2 U2459 ( .B1(n8510), .B2(n4317), .C1(n4492), .C2(n3296), .A(n4256), 
        .ZN(N335) );
  NAND2_X2 U2460 ( .A1(exp_fasu[8]), .A2(n4254), .ZN(n4256) );
  OAI221_X2 U2461 ( .B1(n8510), .B2(n4364), .C1(n4499), .C2(n3296), .A(n4257), 
        .ZN(N334) );
  NAND2_X2 U2462 ( .A1(exp_fasu[7]), .A2(n4254), .ZN(n4257) );
  OAI221_X2 U2463 ( .B1(n8510), .B2(n4365), .C1(n4501), .C2(n3296), .A(n4258), 
        .ZN(N333) );
  NAND2_X2 U2464 ( .A1(exp_fasu[6]), .A2(n4254), .ZN(n4258) );
  OAI221_X2 U2465 ( .B1(n8510), .B2(n4363), .C1(n4500), .C2(n3296), .A(n4259), 
        .ZN(N332) );
  NAND2_X2 U2466 ( .A1(exp_fasu[5]), .A2(n4254), .ZN(n4259) );
  OAI221_X2 U2467 ( .B1(n8510), .B2(n4360), .C1(n4502), .C2(n3296), .A(n4260), 
        .ZN(N331) );
  NAND2_X2 U2468 ( .A1(exp_fasu[4]), .A2(n4254), .ZN(n4260) );
  OAI221_X2 U2469 ( .B1(n8510), .B2(n4361), .C1(n4503), .C2(n3296), .A(n4261), 
        .ZN(N330) );
  NAND2_X2 U2470 ( .A1(exp_fasu[3]), .A2(n4254), .ZN(n4261) );
  OAI221_X2 U2473 ( .B1(n4262), .B2(n4362), .C1(n4504), .C2(n4298), .A(n4263), 
        .ZN(N329) );
  NAND2_X2 U2474 ( .A1(exp_fasu[2]), .A2(n4254), .ZN(n4263) );
  OAI221_X2 U2475 ( .B1(n4262), .B2(n4497), .C1(n4358), .C2(n4298), .A(n4264), 
        .ZN(N328) );
  NAND2_X2 U2476 ( .A1(exp_fasu[1]), .A2(n4254), .ZN(n4264) );
  OAI221_X2 U2477 ( .B1(n4262), .B2(n4496), .C1(n4319), .C2(n4298), .A(n4265), 
        .ZN(N327) );
  NAND2_X2 U2478 ( .A1(exp_fasu[0]), .A2(n4254), .ZN(n4265) );
  DFF_X2 opa_r_reg_63_ ( .D(opa[63]), .CK(clk), .Q(opa_r[63]) );
  DFF_X2 opa_r_reg_62_ ( .D(opa[62]), .CK(clk), .QN(n4399) );
  DFF_X2 opa_r_reg_61_ ( .D(opa[61]), .CK(clk), .Q(opa_r[61]), .QN(n4391) );
  DFF_X2 opa_r_reg_60_ ( .D(opa[60]), .CK(clk), .Q(opa_r[60]), .QN(n4394) );
  DFF_X2 opa_r_reg_59_ ( .D(opa[59]), .CK(clk), .Q(opa_r[59]), .QN(n4396) );
  DFF_X2 opa_r_reg_58_ ( .D(opa[58]), .CK(clk), .Q(opa_r[58]), .QN(n4395) );
  DFF_X2 opa_r_reg_57_ ( .D(opa[57]), .CK(clk), .Q(opa_r[57]), .QN(n4393) );
  DFF_X2 opa_r_reg_56_ ( .D(opa[56]), .CK(clk), .Q(opa_r[56]), .QN(n4332) );
  DFF_X2 opa_r_reg_55_ ( .D(opa[55]), .CK(clk), .Q(opa_r[55]), .QN(n4390) );
  DFF_X2 opa_r_reg_54_ ( .D(opa[54]), .CK(clk), .Q(opa_r[54]), .QN(n4331) );
  DFF_X2 opa_r_reg_53_ ( .D(opa[53]), .CK(clk), .Q(opa_r[53]), .QN(n4392) );
  DFF_X2 opa_r_reg_52_ ( .D(opa[52]), .CK(clk), .Q(opa_r[52]), .QN(n4330) );
  DFF_X2 opa_r_reg_51_ ( .D(opa[51]), .CK(clk), .Q(fracta_mul[51]), .QN(n4297)
         );
  DFF_X2 opa_r_reg_50_ ( .D(opa[50]), .CK(clk), .Q(fracta_mul[50]), .QN(n4291)
         );
  DFF_X2 opa_r_reg_49_ ( .D(opa[49]), .CK(clk), .Q(fracta_mul[49]), .QN(n4301)
         );
  DFF_X2 opa_r_reg_48_ ( .D(opa[48]), .CK(clk), .Q(fracta_mul[48]), .QN(n4303)
         );
  DFF_X2 opa_r_reg_47_ ( .D(opa[47]), .CK(clk), .Q(fracta_mul[47]), .QN(n4302)
         );
  DFF_X2 opa_r_reg_46_ ( .D(opa[46]), .CK(clk), .Q(fracta_mul[46]), .QN(n4300)
         );
  DFF_X2 opa_r_reg_45_ ( .D(opa[45]), .CK(clk), .Q(fracta_mul[45]), .QN(n4290)
         );
  DFF_X2 opa_r_reg_44_ ( .D(opa[44]), .CK(clk), .Q(fracta_mul[44]), .QN(n4420)
         );
  DFF_X2 opa_r_reg_43_ ( .D(opa[43]), .CK(clk), .Q(fracta_mul[43]), .QN(n4296)
         );
  DFF_X2 opa_r_reg_42_ ( .D(opa[42]), .CK(clk), .Q(fracta_mul[42]), .QN(n4436)
         );
  DFF_X2 opa_r_reg_41_ ( .D(opa[41]), .CK(clk), .Q(fracta_mul[41]), .QN(n4313)
         );
  DFF_X2 opa_r_reg_40_ ( .D(opa[40]), .CK(clk), .Q(fracta_mul[40]), .QN(n4344)
         );
  DFF_X2 opa_r_reg_39_ ( .D(opa[39]), .CK(clk), .Q(fracta_mul[39]), .QN(n4439)
         );
  DFF_X2 opa_r_reg_38_ ( .D(opa[38]), .CK(clk), .Q(fracta_mul[38]), .QN(n4335)
         );
  DFF_X2 opa_r_reg_37_ ( .D(opa[37]), .CK(clk), .Q(fracta_mul[37]), .QN(n4310)
         );
  DFF_X2 opa_r_reg_36_ ( .D(opa[36]), .CK(clk), .Q(fracta_mul[36]), .QN(n4340)
         );
  DFF_X2 opa_r_reg_35_ ( .D(opa[35]), .CK(clk), .Q(fracta_mul[35]), .QN(n4311)
         );
  DFF_X2 opa_r_reg_34_ ( .D(opa[34]), .CK(clk), .Q(fracta_mul[34]), .QN(n4314)
         );
  DFF_X2 opa_r_reg_33_ ( .D(opa[33]), .CK(clk), .Q(fracta_mul[33]), .QN(n4338)
         );
  DFF_X2 opa_r_reg_32_ ( .D(opa[32]), .CK(clk), .Q(fracta_mul[32]), .QN(n4342)
         );
  DFF_X2 opa_r_reg_31_ ( .D(opa[31]), .CK(clk), .Q(fracta_mul[31]), .QN(n4423)
         );
  DFF_X2 opa_r_reg_30_ ( .D(opa[30]), .CK(clk), .Q(fracta_mul[30]), .QN(n4419)
         );
  DFF_X2 opa_r_reg_29_ ( .D(opa[29]), .CK(clk), .Q(fracta_mul[29]), .QN(n4431)
         );
  DFF_X2 opa_r_reg_28_ ( .D(opa[28]), .CK(clk), .Q(fracta_mul[28]), .QN(n4418)
         );
  DFF_X2 opa_r_reg_27_ ( .D(opa[27]), .CK(clk), .Q(fracta_mul[27]), .QN(n4426)
         );
  DFF_X2 opa_r_reg_26_ ( .D(opa[26]), .CK(clk), .Q(fracta_mul[26]), .QN(n4422)
         );
  DFF_X2 opa_r_reg_25_ ( .D(opa[25]), .CK(clk), .Q(fracta_mul[25]), .QN(n4421)
         );
  DFF_X2 opa_r_reg_24_ ( .D(opa[24]), .CK(clk), .Q(fracta_mul[24]), .QN(n4435)
         );
  DFF_X2 opa_r_reg_23_ ( .D(opa[23]), .CK(clk), .Q(fracta_mul[23]), .QN(n4417)
         );
  DFF_X2 opa_r_reg_22_ ( .D(opa[22]), .CK(clk), .Q(fracta_mul[22]), .QN(n4289)
         );
  DFF_X2 opa_r_reg_21_ ( .D(opa[21]), .CK(clk), .Q(fracta_mul[21]), .QN(n4437)
         );
  DFF_X2 opa_r_reg_20_ ( .D(opa[20]), .CK(clk), .Q(fracta_mul[20]), .QN(n4299)
         );
  DFF_X2 opa_r_reg_19_ ( .D(opa[19]), .CK(clk), .Q(fracta_mul[19]), .QN(n4438)
         );
  DFF_X2 opa_r_reg_18_ ( .D(opa[18]), .CK(clk), .Q(fracta_mul[18]), .QN(n4427)
         );
  DFF_X2 opa_r_reg_17_ ( .D(opa[17]), .CK(clk), .Q(fracta_mul[17]), .QN(n4341)
         );
  DFF_X2 opa_r_reg_16_ ( .D(opa[16]), .CK(clk), .Q(fracta_mul[16]), .QN(n4347)
         );
  DFF_X2 opa_r_reg_15_ ( .D(opa[15]), .CK(clk), .Q(fracta_mul[15]), .QN(n4339)
         );
  DFF_X2 opa_r_reg_14_ ( .D(opa[14]), .CK(clk), .Q(fracta_mul[14]), .QN(n4434)
         );
  DFF_X2 opa_r_reg_13_ ( .D(opa[13]), .CK(clk), .Q(fracta_mul[13]), .QN(n4336)
         );
  DFF_X2 opa_r_reg_12_ ( .D(opa[12]), .CK(clk), .Q(fracta_mul[12]), .QN(n4315)
         );
  DFF_X2 opa_r_reg_11_ ( .D(opa[11]), .CK(clk), .Q(fracta_mul[11]), .QN(n4312)
         );
  DFF_X2 opa_r_reg_10_ ( .D(opa[10]), .CK(clk), .Q(fracta_mul[10]), .QN(n4337)
         );
  DFF_X2 opa_r_reg_9_ ( .D(opa[9]), .CK(clk), .Q(fracta_mul[9]), .QN(n4433) );
  DFF_X2 opa_r_reg_8_ ( .D(opa[8]), .CK(clk), .Q(fracta_mul[8]), .QN(n4430) );
  DFF_X2 opa_r_reg_7_ ( .D(opa[7]), .CK(clk), .Q(fracta_mul[7]), .QN(n4428) );
  DFF_X2 opa_r_reg_6_ ( .D(opa[6]), .CK(clk), .Q(fracta_mul[6]), .QN(n4432) );
  DFF_X2 opa_r_reg_5_ ( .D(opa[5]), .CK(clk), .Q(fracta_mul[5]), .QN(n4343) );
  DFF_X2 opa_r_reg_4_ ( .D(opa[4]), .CK(clk), .Q(fracta_mul[4]), .QN(n4348) );
  DFF_X2 opa_r_reg_3_ ( .D(opa[3]), .CK(clk), .Q(fracta_mul[3]), .QN(n4726) );
  DFF_X2 opa_r_reg_2_ ( .D(opa[2]), .CK(clk), .Q(fracta_mul[2]), .QN(n4801) );
  DFF_X2 opa_r_reg_0_ ( .D(opa[0]), .CK(clk), .Q(fracta_mul[0]), .QN(n4814) );
  DFF_X2 opb_r_reg_63_ ( .D(opb[63]), .CK(clk), .Q(opb_r[63]) );
  DFF_X2 opb_r_reg_62_ ( .D(opb[62]), .CK(clk), .Q(opb_r[62]), .QN(n4828) );
  DFF_X2 opb_r_reg_61_ ( .D(opb[61]), .CK(clk), .Q(opb_r[61]), .QN(n4829) );
  DFF_X2 opb_r_reg_60_ ( .D(opb[60]), .CK(clk), .Q(opb_r[60]), .QN(n4824) );
  DFF_X2 opb_r_reg_57_ ( .D(opb[57]), .CK(clk), .Q(opb_r[57]), .QN(n4827) );
  DFF_X2 opb_r_reg_56_ ( .D(opb[56]), .CK(clk), .Q(opb_r[56]), .QN(n4821) );
  DFF_X2 opb_r_reg_55_ ( .D(opb[55]), .CK(clk), .Q(opb_r[55]), .QN(n4826) );
  DFF_X2 opb_r_reg_54_ ( .D(opb[54]), .CK(clk), .Q(opb_r[54]), .QN(n4832) );
  DFF_X2 opb_r_reg_53_ ( .D(opb[53]), .CK(clk), .Q(opb_r[53]), .QN(n4831) );
  DFF_X2 opb_r_reg_52_ ( .D(opb[52]), .CK(clk), .Q(opb_r[52]), .QN(n4830) );
  DFF_X2 opb_r_reg_51_ ( .D(opb[51]), .CK(clk), .Q(u6_N51), .QN(n4812) );
  DFF_X2 opb_r_reg_50_ ( .D(opb[50]), .CK(clk), .Q(u6_N50), .QN(n4817) );
  DFF_X2 opb_r_reg_49_ ( .D(opb[49]), .CK(clk), .Q(u6_N49), .QN(n4810) );
  DFF_X2 opb_r_reg_48_ ( .D(opb[48]), .CK(clk), .Q(u6_N48), .QN(n4792) );
  DFF_X2 opb_r_reg_46_ ( .D(opb[46]), .CK(clk), .Q(u6_N46), .QN(n4767) );
  DFF_X2 opb_r_reg_45_ ( .D(opb[45]), .CK(clk), .Q(u6_N45), .QN(n4784) );
  DFF_X2 opb_r_reg_43_ ( .D(opb[43]), .CK(clk), .Q(u6_N43), .QN(n4774) );
  DFF_X2 opb_r_reg_40_ ( .D(opb[40]), .CK(clk), .Q(u6_N40), .QN(n4776) );
  DFF_X2 opb_r_reg_39_ ( .D(opb[39]), .CK(clk), .Q(u6_N39), .QN(n4761) );
  DFF_X2 opb_r_reg_37_ ( .D(opb[37]), .CK(clk), .Q(u6_N37), .QN(n4782) );
  DFF_X2 opb_r_reg_36_ ( .D(opb[36]), .CK(clk), .Q(u6_N36), .QN(n4732) );
  DFF_X2 opb_r_reg_35_ ( .D(opb[35]), .CK(clk), .Q(u6_N35), .QN(n4416) );
  DFF_X2 opb_r_reg_33_ ( .D(opb[33]), .CK(clk), .Q(u6_N33), .QN(n4741) );
  DFF_X2 opb_r_reg_32_ ( .D(opb[32]), .CK(clk), .Q(u6_N32), .QN(n4743) );
  DFF_X2 opb_r_reg_31_ ( .D(opb[31]), .CK(clk), .Q(u6_N31), .QN(n4745) );
  DFF_X2 opb_r_reg_30_ ( .D(opb[30]), .CK(clk), .Q(u6_N30), .QN(n4779) );
  DFF_X2 opb_r_reg_29_ ( .D(opb[29]), .CK(clk), .Q(u6_N29), .QN(n4737) );
  DFF_X2 opb_r_reg_27_ ( .D(opb[27]), .CK(clk), .Q(u6_N27), .QN(n4757) );
  DFF_X2 opb_r_reg_26_ ( .D(opb[26]), .CK(clk), .Q(u6_N26), .QN(n4755) );
  DFF_X2 opb_r_reg_25_ ( .D(opb[25]), .CK(clk), .Q(u6_N25), .QN(n4751) );
  DFF_X2 opb_r_reg_24_ ( .D(opb[24]), .CK(clk), .Q(u6_N24), .QN(n4759) );
  DFF_X2 opb_r_reg_23_ ( .D(opb[23]), .CK(clk), .Q(u6_N23), .QN(n4753) );
  DFF_X2 opb_r_reg_22_ ( .D(opb[22]), .CK(clk), .Q(u6_N22), .QN(n4749) );
  DFF_X2 opb_r_reg_21_ ( .D(opb[21]), .CK(clk), .Q(u6_N21), .QN(n4747) );
  DFF_X2 opb_r_reg_20_ ( .D(opb[20]), .CK(clk), .Q(u6_N20), .QN(n4739) );
  DFF_X2 opb_r_reg_19_ ( .D(opb[19]), .CK(clk), .Q(u6_N19), .QN(n4728) );
  DFF_X2 opb_r_reg_18_ ( .D(opb[18]), .CK(clk), .Q(u6_N18), .QN(n4724) );
  DFF_X2 opb_r_reg_17_ ( .D(opb[17]), .CK(clk), .Q(u6_N17), .QN(n4454) );
  DFF_X2 opb_r_reg_16_ ( .D(opb[16]), .CK(clk), .Q(u6_N16), .QN(n4455) );
  DFF_X2 opb_r_reg_15_ ( .D(opb[15]), .CK(clk), .Q(u6_N15), .QN(n4453) );
  DFF_X2 opb_r_reg_14_ ( .D(opb[14]), .CK(clk), .Q(u6_N14), .QN(n4441) );
  DFF_X2 opb_r_reg_13_ ( .D(opb[13]), .CK(clk), .Q(u6_N13), .QN(n4440) );
  DFF_X2 opb_r_reg_12_ ( .D(opb[12]), .CK(clk), .Q(u6_N12), .QN(n4442) );
  DFF_X2 opb_r_reg_11_ ( .D(opb[11]), .CK(clk), .Q(u6_N11), .QN(n4452) );
  DFF_X2 opb_r_reg_10_ ( .D(opb[10]), .CK(clk), .Q(u6_N10), .QN(n4451) );
  DFF_X2 opb_r_reg_9_ ( .D(opb[9]), .CK(clk), .Q(u6_N9), .QN(n4449) );
  DFF_X2 opb_r_reg_8_ ( .D(opb[8]), .CK(clk), .Q(u6_N8), .QN(n4450) );
  DFF_X2 opb_r_reg_7_ ( .D(opb[7]), .CK(clk), .Q(u6_N7), .QN(n4448) );
  DFF_X2 opb_r_reg_6_ ( .D(opb[6]), .CK(clk), .Q(u6_N6), .QN(n4447) );
  DFF_X2 opb_r_reg_5_ ( .D(opb[5]), .CK(clk), .Q(u6_N5), .QN(n4460) );
  DFF_X2 opb_r_reg_4_ ( .D(opb[4]), .CK(clk), .Q(u6_N4), .QN(n4459) );
  DFF_X2 opb_r_reg_3_ ( .D(opb[3]), .CK(clk), .Q(u6_N3), .QN(n4458) );
  DFF_X2 opb_r_reg_2_ ( .D(opb[2]), .CK(clk), .Q(u6_N2), .QN(n4456) );
  DFF_X2 opb_r_reg_1_ ( .D(opb[1]), .CK(clk), .Q(u6_N1), .QN(n4457) );
  DFF_X2 opb_r_reg_0_ ( .D(opb[0]), .CK(clk), .Q(u6_N0), .QN(n4351) );
  DFF_X2 rmode_r1_reg_1_ ( .D(rmode[1]), .CK(clk), .Q(rmode_r1[1]) );
  DFF_X2 rmode_r1_reg_0_ ( .D(rmode[0]), .CK(clk), .Q(rmode_r1[0]) );
  DFF_X2 rmode_r2_reg_1_ ( .D(rmode_r1[1]), .CK(clk), .Q(rmode_r2[1]) );
  DFF_X2 rmode_r2_reg_0_ ( .D(rmode_r1[0]), .CK(clk), .Q(rmode_r2[0]) );
  DFF_X2 rmode_r3_reg_1_ ( .D(rmode_r2[1]), .CK(clk), .Q(rmode_r3[1]), .QN(
        n4334) );
  DFF_X2 rmode_r3_reg_0_ ( .D(rmode_r2[0]), .CK(clk), .Q(rmode_r3[0]), .QN(
        n4401) );
  DFF_X2 fpu_op_r1_reg_2_ ( .D(fpu_op[2]), .CK(clk), .Q(fpu_op_r1[2]), .QN(
        n4352) );
  DFF_X2 fpu_op_r1_reg_1_ ( .D(fpu_op[1]), .CK(clk), .Q(fpu_op_r1[1]) );
  DFF_X2 fpu_op_r1_reg_0_ ( .D(fpu_op[0]), .CK(clk), .Q(fpu_op_r1[0]), .QN(
        n4445) );
  DFF_X2 fpu_op_r2_reg_2_ ( .D(fpu_op_r1[2]), .CK(clk), .Q(fpu_op_r2[2]) );
  DFF_X2 fpu_op_r2_reg_1_ ( .D(fpu_op_r1[1]), .CK(clk), .Q(fpu_op_r2[1]), .QN(
        n4298) );
  DFF_X2 fpu_op_r2_reg_0_ ( .D(fpu_op_r1[0]), .CK(clk), .Q(fpu_op_r2[0]), .QN(
        n4495) );
  DFF_X2 fpu_op_r3_reg_2_ ( .D(fpu_op_r2[2]), .CK(clk), .Q(n4294), .QN(n4376)
         );
  DFF_X2 fpu_op_r3_reg_1_ ( .D(fpu_op_r2[1]), .CK(clk), .Q(fpu_op_r3[1]), .QN(
        n4288) );
  DFF_X2 fpu_op_r3_reg_0_ ( .D(fpu_op_r2[0]), .CK(clk), .Q(fpu_op_r3[0]), .QN(
        n4366) );
  DFF_X2 div_opa_ldz_r1_reg_4_ ( .D(div_opa_ldz_d[4]), .CK(clk), .Q(
        div_opa_ldz_r1[4]) );
  DFF_X2 div_opa_ldz_r1_reg_3_ ( .D(div_opa_ldz_d[3]), .CK(clk), .Q(
        div_opa_ldz_r1[3]) );
  DFF_X2 div_opa_ldz_r1_reg_2_ ( .D(div_opa_ldz_d[2]), .CK(clk), .Q(
        div_opa_ldz_r1[2]) );
  DFF_X2 div_opa_ldz_r1_reg_1_ ( .D(div_opa_ldz_d[1]), .CK(clk), .Q(
        div_opa_ldz_r1[1]) );
  DFF_X2 div_opa_ldz_r1_reg_0_ ( .D(div_opa_ldz_d[0]), .CK(clk), .Q(
        div_opa_ldz_r1[0]) );
  DFF_X2 div_opa_ldz_r2_reg_4_ ( .D(div_opa_ldz_r1[4]), .CK(clk), .Q(
        div_opa_ldz_r2[4]), .QN(n4387) );
  DFF_X2 div_opa_ldz_r2_reg_3_ ( .D(div_opa_ldz_r1[3]), .CK(clk), .Q(
        div_opa_ldz_r2[3]), .QN(n4386) );
  DFF_X2 div_opa_ldz_r2_reg_2_ ( .D(div_opa_ldz_r1[2]), .CK(clk), .Q(
        div_opa_ldz_r2[2]), .QN(n4324) );
  DFF_X2 div_opa_ldz_r2_reg_1_ ( .D(div_opa_ldz_r1[1]), .CK(clk), .Q(
        div_opa_ldz_r2[1]), .QN(n4377) );
  DFF_X2 div_opa_ldz_r2_reg_0_ ( .D(div_opa_ldz_r1[0]), .CK(clk), .Q(
        div_opa_ldz_r2[0]), .QN(n4381) );
  DFF_X2 opa_r1_reg_62_ ( .D(n4853), .CK(clk), .QN(n4349) );
  DFF_X2 opa_r1_reg_61_ ( .D(opa_r[61]), .CK(clk), .QN(n4444) );
  DFF_X2 opa_r1_reg_60_ ( .D(opa_r[60]), .CK(clk), .QN(n4317) );
  DFF_X2 opa_r1_reg_59_ ( .D(opa_r[59]), .CK(clk), .Q(opa_r1[59]), .QN(n4364)
         );
  DFF_X2 opa_r1_reg_58_ ( .D(opa_r[58]), .CK(clk), .Q(opa_r1[58]), .QN(n4365)
         );
  DFF_X2 opa_r1_reg_57_ ( .D(opa_r[57]), .CK(clk), .Q(opa_r1[57]), .QN(n4363)
         );
  DFF_X2 opa_r1_reg_56_ ( .D(opa_r[56]), .CK(clk), .Q(opa_r1[56]), .QN(n4360)
         );
  DFF_X2 opa_r1_reg_55_ ( .D(opa_r[55]), .CK(clk), .Q(opa_r1[55]), .QN(n4361)
         );
  DFF_X2 opa_r1_reg_54_ ( .D(opa_r[54]), .CK(clk), .Q(opa_r1[54]), .QN(n4362)
         );
  DFF_X2 opa_r1_reg_53_ ( .D(opa_r[53]), .CK(clk), .Q(opa_r1[53]), .QN(n4497)
         );
  DFF_X2 opa_r1_reg_52_ ( .D(opa_r[52]), .CK(clk), .Q(opa_r1[52]), .QN(n4496)
         );
  DFF_X2 opa_r1_reg_51_ ( .D(fracta_mul[51]), .CK(clk), .Q(opa_r1[51]) );
  DFF_X2 opa_r1_reg_50_ ( .D(fracta_mul[50]), .CK(clk), .Q(opa_r1[50]) );
  DFF_X2 opa_r1_reg_49_ ( .D(fracta_mul[49]), .CK(clk), .Q(opa_r1[49]) );
  DFF_X2 opa_r1_reg_48_ ( .D(fracta_mul[48]), .CK(clk), .Q(opa_r1[48]) );
  DFF_X2 opa_r1_reg_47_ ( .D(fracta_mul[47]), .CK(clk), .Q(opa_r1[47]) );
  DFF_X2 opa_r1_reg_46_ ( .D(fracta_mul[46]), .CK(clk), .Q(opa_r1[46]) );
  DFF_X2 opa_r1_reg_45_ ( .D(fracta_mul[45]), .CK(clk), .Q(opa_r1[45]) );
  DFF_X2 opa_r1_reg_44_ ( .D(fracta_mul[44]), .CK(clk), .Q(opa_r1[44]) );
  DFF_X2 opa_r1_reg_43_ ( .D(fracta_mul[43]), .CK(clk), .Q(opa_r1[43]) );
  DFF_X2 opa_r1_reg_42_ ( .D(fracta_mul[42]), .CK(clk), .Q(opa_r1[42]) );
  DFF_X2 opa_r1_reg_41_ ( .D(fracta_mul[41]), .CK(clk), .Q(opa_r1[41]) );
  DFF_X2 opa_r1_reg_40_ ( .D(fracta_mul[40]), .CK(clk), .Q(opa_r1[40]) );
  DFF_X2 opa_r1_reg_39_ ( .D(fracta_mul[39]), .CK(clk), .Q(opa_r1[39]) );
  DFF_X2 opa_r1_reg_38_ ( .D(fracta_mul[38]), .CK(clk), .Q(opa_r1[38]) );
  DFF_X2 opa_r1_reg_37_ ( .D(fracta_mul[37]), .CK(clk), .Q(opa_r1[37]) );
  DFF_X2 opa_r1_reg_36_ ( .D(fracta_mul[36]), .CK(clk), .Q(opa_r1[36]) );
  DFF_X2 opa_r1_reg_35_ ( .D(fracta_mul[35]), .CK(clk), .Q(opa_r1[35]) );
  DFF_X2 opa_r1_reg_34_ ( .D(fracta_mul[34]), .CK(clk), .Q(opa_r1[34]) );
  DFF_X2 opa_r1_reg_33_ ( .D(fracta_mul[33]), .CK(clk), .Q(opa_r1[33]) );
  DFF_X2 opa_r1_reg_32_ ( .D(fracta_mul[32]), .CK(clk), .Q(opa_r1[32]) );
  DFF_X2 opa_r1_reg_31_ ( .D(fracta_mul[31]), .CK(clk), .Q(opa_r1[31]) );
  DFF_X2 opa_r1_reg_30_ ( .D(fracta_mul[30]), .CK(clk), .Q(opa_r1[30]) );
  DFF_X2 opa_r1_reg_29_ ( .D(fracta_mul[29]), .CK(clk), .Q(opa_r1[29]) );
  DFF_X2 opa_r1_reg_28_ ( .D(fracta_mul[28]), .CK(clk), .Q(opa_r1[28]) );
  DFF_X2 opa_r1_reg_27_ ( .D(fracta_mul[27]), .CK(clk), .Q(opa_r1[27]) );
  DFF_X2 opa_r1_reg_26_ ( .D(fracta_mul[26]), .CK(clk), .Q(opa_r1[26]) );
  DFF_X2 opa_r1_reg_25_ ( .D(fracta_mul[25]), .CK(clk), .Q(opa_r1[25]) );
  DFF_X2 opa_r1_reg_24_ ( .D(fracta_mul[24]), .CK(clk), .Q(opa_r1[24]) );
  DFF_X2 opa_r1_reg_23_ ( .D(fracta_mul[23]), .CK(clk), .Q(opa_r1[23]) );
  DFF_X2 opa_r1_reg_22_ ( .D(fracta_mul[22]), .CK(clk), .Q(opa_r1[22]) );
  DFF_X2 opa_r1_reg_21_ ( .D(fracta_mul[21]), .CK(clk), .Q(opa_r1[21]) );
  DFF_X2 opa_r1_reg_20_ ( .D(fracta_mul[20]), .CK(clk), .Q(opa_r1[20]) );
  DFF_X2 opa_r1_reg_19_ ( .D(fracta_mul[19]), .CK(clk), .Q(opa_r1[19]) );
  DFF_X2 opa_r1_reg_18_ ( .D(fracta_mul[18]), .CK(clk), .Q(opa_r1[18]) );
  DFF_X2 opa_r1_reg_17_ ( .D(fracta_mul[17]), .CK(clk), .Q(opa_r1[17]) );
  DFF_X2 opa_r1_reg_16_ ( .D(fracta_mul[16]), .CK(clk), .Q(opa_r1[16]) );
  DFF_X2 opa_r1_reg_15_ ( .D(fracta_mul[15]), .CK(clk), .Q(opa_r1[15]) );
  DFF_X2 opa_r1_reg_14_ ( .D(fracta_mul[14]), .CK(clk), .Q(opa_r1[14]) );
  DFF_X2 opa_r1_reg_13_ ( .D(fracta_mul[13]), .CK(clk), .Q(opa_r1[13]) );
  DFF_X2 opa_r1_reg_12_ ( .D(fracta_mul[12]), .CK(clk), .Q(opa_r1[12]) );
  DFF_X2 opa_r1_reg_11_ ( .D(fracta_mul[11]), .CK(clk), .Q(opa_r1[11]) );
  DFF_X2 opa_r1_reg_10_ ( .D(fracta_mul[10]), .CK(clk), .Q(opa_r1[10]) );
  DFF_X2 opa_r1_reg_9_ ( .D(fracta_mul[9]), .CK(clk), .Q(opa_r1[9]) );
  DFF_X2 opa_r1_reg_8_ ( .D(fracta_mul[8]), .CK(clk), .Q(opa_r1[8]) );
  DFF_X2 opa_r1_reg_7_ ( .D(fracta_mul[7]), .CK(clk), .Q(opa_r1[7]) );
  DFF_X2 opa_r1_reg_6_ ( .D(fracta_mul[6]), .CK(clk), .Q(opa_r1[6]) );
  DFF_X2 opa_r1_reg_5_ ( .D(fracta_mul[5]), .CK(clk), .Q(opa_r1[5]) );
  DFF_X2 opa_r1_reg_4_ ( .D(fracta_mul[4]), .CK(clk), .Q(opa_r1[4]) );
  DFF_X2 opa_r1_reg_3_ ( .D(n4727), .CK(clk), .Q(opa_r1[3]) );
  DFF_X2 opa_r1_reg_2_ ( .D(fracta_mul[2]), .CK(clk), .Q(opa_r1[2]) );
  DFF_X2 opa_r1_reg_1_ ( .D(n4799), .CK(clk), .Q(opa_r1[1]) );
  DFF_X2 opa_r1_reg_0_ ( .D(fracta_mul[0]), .CK(clk), .Q(N343), .QN(n4491) );
  DFF_X2 opas_r1_reg ( .D(opa_r[63]), .CK(clk), .Q(opas_r1) );
  DFF_X2 opas_r2_reg ( .D(opas_r1), .CK(clk), .Q(opas_r2) );
  DFF_X2 u0_fractb_00_reg ( .D(n4346), .CK(clk), .Q(u0_fractb_00) );
  DFF_X2 u0_fracta_00_reg ( .D(n7197), .CK(clk), .Q(u0_fracta_00) );
  DFF_X2 u0_expb_00_reg ( .D(n7209), .CK(clk), .Q(u0_expb_00) );
  DFF_X2 u0_opb_dn_reg ( .D(u0_expb_00), .CK(clk), .Q(opb_dn), .QN(n4519) );
  DFF_X2 u0_opb_00_reg ( .D(u0_N17), .CK(clk), .Q(opb_00), .QN(n4461) );
  DFF_X2 u0_expa_00_reg ( .D(n4902), .CK(clk), .Q(u0_expa_00) );
  DFF_X2 u0_opa_dn_reg ( .D(u0_expa_00), .CK(clk), .Q(opa_dn), .QN(n4389) );
  DFF_X2 u0_opa_00_reg ( .D(u0_N16), .CK(clk), .Q(opa_00), .QN(n4446) );
  DFF_X2 u0_opb_nan_reg ( .D(u0_N11), .CK(clk), .Q(opb_nan), .QN(n4494) );
  DFF_X2 u0_opa_nan_reg ( .D(u0_N10), .CK(clk), .Q(opa_nan) );
  DFF_X2 opa_nan_r_reg ( .D(N912), .CK(clk), .Q(opa_nan_r) );
  DFF_X2 u0_snan_r_b_reg ( .D(u0_N5), .CK(clk), .Q(u0_snan_r_b) );
  DFF_X2 u0_qnan_r_b_reg ( .D(u6_N51), .CK(clk), .Q(u0_qnan_r_b) );
  DFF_X2 u0_snan_r_a_reg ( .D(u0_N4), .CK(clk), .Q(u0_snan_r_a) );
  DFF_X2 u0_qnan_r_a_reg ( .D(fracta_mul[51]), .CK(clk), .Q(u0_qnan_r_a) );
  DFF_X2 u0_infb_f_r_reg ( .D(n4346), .CK(clk), .Q(u0_infb_f_r) );
  DFF_X2 u0_infa_f_r_reg ( .D(n7197), .CK(clk), .Q(u0_infa_f_r) );
  DFF_X2 u0_expb_ff_reg ( .D(n8508), .CK(clk), .Q(u0_expb_ff) );
  DFF_X2 u0_opb_inf_reg ( .D(n8528), .CK(clk), .Q(opb_inf), .QN(n4429) );
  DFF_X2 u0_expa_ff_reg ( .D(n7195), .CK(clk), .Q(u0_expa_ff) );
  DFF_X2 u0_snan_reg ( .D(n8526), .CK(clk), .Q(snan_d), .QN(n4355) );
  DFF_X2 snan_reg ( .D(snan_d), .CK(clk), .Q(snan) );
  DFF_X2 u0_qnan_reg ( .D(n8527), .CK(clk), .QN(n4482) );
  DFF_X2 u0_opa_inf_reg ( .D(n8529), .CK(clk), .Q(opa_inf), .QN(n4345) );
  DFF_X2 div_by_zero_reg ( .D(N913), .CK(clk), .Q(div_by_zero) );
  DFF_X2 u0_inf_reg ( .D(u0_N7), .CK(clk), .Q(inf_d), .QN(n4478) );
  DFF_X2 u0_ind_reg ( .D(u0_N6), .CK(clk), .Q(ind_d) );
  DFF_X2 u1_fasu_op_reg ( .D(u1_N232), .CK(clk), .Q(n4287), .QN(n4304) );
  DFF_X2 fasu_op_r1_reg ( .D(n4916), .CK(clk), .Q(fasu_op_r1) );
  DFF_X2 fasu_op_r2_reg ( .D(fasu_op_r1), .CK(clk), .QN(n4484) );
  DFF_X2 qnan_reg ( .D(N904), .CK(clk), .Q(qnan) );
  DFF_X2 u1_fracta_eq_fractb_reg ( .D(u1_N220), .CK(clk), .Q(
        u1_fracta_eq_fractb) );
  DFF_X2 u1_fracta_lt_fractb_reg ( .D(u1_N219), .CK(clk), .Q(
        u1_fracta_lt_fractb) );
  DFF_X2 u1_add_r_reg ( .D(n4445), .CK(clk), .Q(u1_add_r) );
  DFF_X2 u1_signb_r_reg ( .D(opb_r[63]), .CK(clk), .Q(u1_signb_r), .QN(n4498)
         );
  DFF_X2 u1_signa_r_reg ( .D(opa_r[63]), .CK(clk), .Q(u1_signa_r), .QN(n4493)
         );
  DFF_X2 u1_result_zero_sign_reg ( .D(u1_N218), .CK(clk), .Q(
        result_zero_sign_d) );
  DFF_X2 u1_nan_sign_reg ( .D(u1_N229), .CK(clk), .Q(nan_sign_d) );
  DFF_X2 sign_fasu_r_reg ( .D(sign_fasu), .CK(clk), .Q(sign_fasu_r) );
  DFF_X2 u1_fractb_out_reg_0_ ( .D(u1_fractb_s[0]), .CK(clk), .Q(fractb[0]) );
  DFF_X2 u1_fractb_out_reg_1_ ( .D(u1_fractb_s[1]), .CK(clk), .Q(fractb[1]) );
  DFF_X2 u1_fractb_out_reg_2_ ( .D(u1_fractb_s[2]), .CK(clk), .Q(fractb[2]) );
  DFF_X2 u1_fractb_out_reg_3_ ( .D(u1_fractb_s[3]), .CK(clk), .Q(fractb[3]) );
  DFF_X2 u1_fractb_out_reg_4_ ( .D(u1_fractb_s[4]), .CK(clk), .Q(fractb[4]) );
  DFF_X2 u1_fractb_out_reg_5_ ( .D(u1_fractb_s[5]), .CK(clk), .Q(fractb[5]) );
  DFF_X2 u1_fractb_out_reg_6_ ( .D(u1_fractb_s[6]), .CK(clk), .Q(fractb[6]) );
  DFF_X2 u1_fractb_out_reg_7_ ( .D(u1_fractb_s[7]), .CK(clk), .Q(fractb[7]) );
  DFF_X2 u1_fractb_out_reg_8_ ( .D(u1_fractb_s[8]), .CK(clk), .Q(fractb[8]) );
  DFF_X2 u1_fractb_out_reg_9_ ( .D(u1_fractb_s[9]), .CK(clk), .Q(fractb[9]) );
  DFF_X2 u1_fractb_out_reg_10_ ( .D(u1_fractb_s[10]), .CK(clk), .Q(fractb[10])
         );
  DFF_X2 u1_fractb_out_reg_11_ ( .D(u1_fractb_s[11]), .CK(clk), .Q(fractb[11])
         );
  DFF_X2 u1_fractb_out_reg_12_ ( .D(u1_fractb_s[12]), .CK(clk), .Q(fractb[12])
         );
  DFF_X2 u1_fractb_out_reg_13_ ( .D(u1_fractb_s[13]), .CK(clk), .Q(fractb[13])
         );
  DFF_X2 u1_fractb_out_reg_14_ ( .D(u1_fractb_s[14]), .CK(clk), .Q(fractb[14])
         );
  DFF_X2 u1_fractb_out_reg_15_ ( .D(u1_fractb_s[15]), .CK(clk), .Q(fractb[15])
         );
  DFF_X2 u1_fractb_out_reg_16_ ( .D(u1_fractb_s[16]), .CK(clk), .Q(fractb[16])
         );
  DFF_X2 u1_fractb_out_reg_17_ ( .D(u1_fractb_s[17]), .CK(clk), .Q(fractb[17])
         );
  DFF_X2 u1_fractb_out_reg_18_ ( .D(u1_fractb_s[18]), .CK(clk), .Q(fractb[18])
         );
  DFF_X2 u1_fractb_out_reg_19_ ( .D(u1_fractb_s[19]), .CK(clk), .Q(fractb[19])
         );
  DFF_X2 u1_fractb_out_reg_20_ ( .D(u1_fractb_s[20]), .CK(clk), .Q(fractb[20])
         );
  DFF_X2 u1_fractb_out_reg_21_ ( .D(u1_fractb_s[21]), .CK(clk), .Q(fractb[21])
         );
  DFF_X2 u1_fractb_out_reg_22_ ( .D(u1_fractb_s[22]), .CK(clk), .Q(fractb[22])
         );
  DFF_X2 u1_fractb_out_reg_23_ ( .D(u1_fractb_s[23]), .CK(clk), .Q(fractb[23])
         );
  DFF_X2 u1_fractb_out_reg_24_ ( .D(u1_fractb_s[24]), .CK(clk), .Q(fractb[24])
         );
  DFF_X2 u1_fractb_out_reg_25_ ( .D(u1_fractb_s[25]), .CK(clk), .Q(fractb[25])
         );
  DFF_X2 u1_fractb_out_reg_26_ ( .D(u1_fractb_s[26]), .CK(clk), .Q(fractb[26])
         );
  DFF_X2 u1_fractb_out_reg_27_ ( .D(u1_fractb_s[27]), .CK(clk), .Q(fractb[27])
         );
  DFF_X2 u1_fractb_out_reg_28_ ( .D(u1_fractb_s[28]), .CK(clk), .Q(fractb[28])
         );
  DFF_X2 u1_fractb_out_reg_29_ ( .D(u1_fractb_s[29]), .CK(clk), .Q(fractb[29])
         );
  DFF_X2 u1_fractb_out_reg_30_ ( .D(u1_fractb_s[30]), .CK(clk), .Q(fractb[30])
         );
  DFF_X2 u1_fractb_out_reg_31_ ( .D(u1_fractb_s[31]), .CK(clk), .Q(fractb[31])
         );
  DFF_X2 u1_fractb_out_reg_32_ ( .D(u1_fractb_s[32]), .CK(clk), .Q(fractb[32])
         );
  DFF_X2 u1_fractb_out_reg_33_ ( .D(u1_fractb_s[33]), .CK(clk), .Q(fractb[33])
         );
  DFF_X2 u1_fractb_out_reg_34_ ( .D(u1_fractb_s[34]), .CK(clk), .Q(fractb[34])
         );
  DFF_X2 u1_fractb_out_reg_35_ ( .D(u1_fractb_s[35]), .CK(clk), .Q(fractb[35])
         );
  DFF_X2 u1_fractb_out_reg_36_ ( .D(u1_fractb_s[36]), .CK(clk), .Q(fractb[36])
         );
  DFF_X2 u1_fractb_out_reg_37_ ( .D(u1_fractb_s[37]), .CK(clk), .Q(fractb[37])
         );
  DFF_X2 u1_fractb_out_reg_38_ ( .D(u1_fractb_s[38]), .CK(clk), .Q(fractb[38])
         );
  DFF_X2 u1_fractb_out_reg_39_ ( .D(u1_fractb_s[39]), .CK(clk), .Q(fractb[39])
         );
  DFF_X2 u1_fractb_out_reg_40_ ( .D(u1_fractb_s[40]), .CK(clk), .Q(fractb[40])
         );
  DFF_X2 u1_fractb_out_reg_41_ ( .D(u1_fractb_s[41]), .CK(clk), .Q(fractb[41])
         );
  DFF_X2 u1_fractb_out_reg_42_ ( .D(u1_fractb_s[42]), .CK(clk), .Q(fractb[42])
         );
  DFF_X2 u1_fractb_out_reg_43_ ( .D(u1_fractb_s[43]), .CK(clk), .Q(fractb[43])
         );
  DFF_X2 u1_fractb_out_reg_44_ ( .D(u1_fractb_s[44]), .CK(clk), .Q(fractb[44])
         );
  DFF_X2 u1_fractb_out_reg_45_ ( .D(u1_fractb_s[45]), .CK(clk), .Q(fractb[45])
         );
  DFF_X2 u1_fractb_out_reg_46_ ( .D(u1_fractb_s[46]), .CK(clk), .Q(fractb[46])
         );
  DFF_X2 u1_fractb_out_reg_47_ ( .D(u1_fractb_s[47]), .CK(clk), .Q(fractb[47])
         );
  DFF_X2 u1_fractb_out_reg_48_ ( .D(u1_fractb_s[48]), .CK(clk), .Q(fractb[48])
         );
  DFF_X2 u1_fractb_out_reg_49_ ( .D(u1_fractb_s[49]), .CK(clk), .Q(fractb[49])
         );
  DFF_X2 u1_fractb_out_reg_50_ ( .D(u1_fractb_s[50]), .CK(clk), .Q(fractb[50])
         );
  DFF_X2 u1_fractb_out_reg_51_ ( .D(u1_fractb_s[51]), .CK(clk), .Q(fractb[51])
         );
  DFF_X2 u1_fractb_out_reg_52_ ( .D(u1_fractb_s[52]), .CK(clk), .Q(fractb[52])
         );
  DFF_X2 u1_fractb_out_reg_53_ ( .D(u1_fractb_s[53]), .CK(clk), .Q(fractb[53])
         );
  DFF_X2 u1_fractb_out_reg_54_ ( .D(u1_fractb_s[54]), .CK(clk), .Q(fractb[54])
         );
  DFF_X2 u1_fractb_out_reg_55_ ( .D(u1_fractb_s[55]), .CK(clk), .Q(fractb[55])
         );
  DFF_X2 u1_fracta_out_reg_0_ ( .D(u1_fracta_s[0]), .CK(clk), .Q(fracta[0]) );
  DFF_X2 u1_fracta_out_reg_1_ ( .D(u1_fracta_s[1]), .CK(clk), .Q(fracta[1]) );
  DFF_X2 u1_fracta_out_reg_2_ ( .D(u1_fracta_s[2]), .CK(clk), .Q(fracta[2]) );
  DFF_X2 u1_fracta_out_reg_3_ ( .D(u1_fracta_s[3]), .CK(clk), .Q(fracta[3]) );
  DFF_X2 u1_fracta_out_reg_4_ ( .D(u1_fracta_s[4]), .CK(clk), .Q(fracta[4]) );
  DFF_X2 u1_fracta_out_reg_5_ ( .D(u1_fracta_s[5]), .CK(clk), .Q(fracta[5]) );
  DFF_X2 u1_fracta_out_reg_6_ ( .D(u1_fracta_s[6]), .CK(clk), .Q(fracta[6]) );
  DFF_X2 u1_fracta_out_reg_7_ ( .D(u1_fracta_s[7]), .CK(clk), .Q(fracta[7]) );
  DFF_X2 u1_fracta_out_reg_8_ ( .D(u1_fracta_s[8]), .CK(clk), .Q(fracta[8]) );
  DFF_X2 u1_fracta_out_reg_9_ ( .D(u1_fracta_s[9]), .CK(clk), .Q(fracta[9]) );
  DFF_X2 u1_fracta_out_reg_10_ ( .D(u1_fracta_s[10]), .CK(clk), .Q(fracta[10])
         );
  DFF_X2 u1_fracta_out_reg_11_ ( .D(u1_fracta_s[11]), .CK(clk), .Q(fracta[11])
         );
  DFF_X2 u1_fracta_out_reg_12_ ( .D(u1_fracta_s[12]), .CK(clk), .Q(fracta[12])
         );
  DFF_X2 u1_fracta_out_reg_13_ ( .D(u1_fracta_s[13]), .CK(clk), .Q(fracta[13])
         );
  DFF_X2 u1_fracta_out_reg_14_ ( .D(u1_fracta_s[14]), .CK(clk), .Q(fracta[14])
         );
  DFF_X2 u1_fracta_out_reg_15_ ( .D(u1_fracta_s[15]), .CK(clk), .Q(fracta[15])
         );
  DFF_X2 u1_fracta_out_reg_16_ ( .D(u1_fracta_s[16]), .CK(clk), .Q(fracta[16])
         );
  DFF_X2 u1_fracta_out_reg_17_ ( .D(u1_fracta_s[17]), .CK(clk), .Q(fracta[17])
         );
  DFF_X2 u1_fracta_out_reg_18_ ( .D(u1_fracta_s[18]), .CK(clk), .Q(fracta[18])
         );
  DFF_X2 u1_fracta_out_reg_19_ ( .D(u1_fracta_s[19]), .CK(clk), .Q(fracta[19])
         );
  DFF_X2 u1_fracta_out_reg_20_ ( .D(u1_fracta_s[20]), .CK(clk), .Q(fracta[20])
         );
  DFF_X2 u1_fracta_out_reg_21_ ( .D(u1_fracta_s[21]), .CK(clk), .Q(fracta[21])
         );
  DFF_X2 u1_fracta_out_reg_22_ ( .D(u1_fracta_s[22]), .CK(clk), .Q(fracta[22])
         );
  DFF_X2 u1_fracta_out_reg_23_ ( .D(u1_fracta_s[23]), .CK(clk), .Q(fracta[23])
         );
  DFF_X2 u1_fracta_out_reg_24_ ( .D(u1_fracta_s[24]), .CK(clk), .Q(fracta[24])
         );
  DFF_X2 u1_fracta_out_reg_25_ ( .D(u1_fracta_s[25]), .CK(clk), .Q(fracta[25])
         );
  DFF_X2 u1_fracta_out_reg_26_ ( .D(u1_fracta_s[26]), .CK(clk), .Q(fracta[26])
         );
  DFF_X2 u1_fracta_out_reg_27_ ( .D(u1_fracta_s[27]), .CK(clk), .Q(fracta[27])
         );
  DFF_X2 u1_fracta_out_reg_28_ ( .D(u1_fracta_s[28]), .CK(clk), .Q(fracta[28])
         );
  DFF_X2 u1_fracta_out_reg_29_ ( .D(u1_fracta_s[29]), .CK(clk), .Q(fracta[29])
         );
  DFF_X2 u1_fracta_out_reg_30_ ( .D(u1_fracta_s[30]), .CK(clk), .Q(fracta[30])
         );
  DFF_X2 u1_fracta_out_reg_31_ ( .D(u1_fracta_s[31]), .CK(clk), .Q(fracta[31])
         );
  DFF_X2 u1_fracta_out_reg_32_ ( .D(u1_fracta_s[32]), .CK(clk), .Q(fracta[32])
         );
  DFF_X2 u1_fracta_out_reg_33_ ( .D(u1_fracta_s[33]), .CK(clk), .Q(fracta[33])
         );
  DFF_X2 u1_fracta_out_reg_34_ ( .D(u1_fracta_s[34]), .CK(clk), .Q(fracta[34])
         );
  DFF_X2 u1_fracta_out_reg_35_ ( .D(u1_fracta_s[35]), .CK(clk), .Q(fracta[35])
         );
  DFF_X2 u1_fracta_out_reg_36_ ( .D(u1_fracta_s[36]), .CK(clk), .Q(fracta[36])
         );
  DFF_X2 u1_fracta_out_reg_37_ ( .D(u1_fracta_s[37]), .CK(clk), .Q(fracta[37])
         );
  DFF_X2 u1_fracta_out_reg_38_ ( .D(u1_fracta_s[38]), .CK(clk), .Q(fracta[38])
         );
  DFF_X2 u1_fracta_out_reg_39_ ( .D(u1_fracta_s[39]), .CK(clk), .Q(fracta[39])
         );
  DFF_X2 u1_fracta_out_reg_40_ ( .D(u1_fracta_s[40]), .CK(clk), .Q(fracta[40])
         );
  DFF_X2 u1_fracta_out_reg_41_ ( .D(u1_fracta_s[41]), .CK(clk), .Q(fracta[41])
         );
  DFF_X2 u1_fracta_out_reg_42_ ( .D(u1_fracta_s[42]), .CK(clk), .Q(fracta[42])
         );
  DFF_X2 u1_fracta_out_reg_43_ ( .D(u1_fracta_s[43]), .CK(clk), .Q(fracta[43])
         );
  DFF_X2 u1_fracta_out_reg_44_ ( .D(u1_fracta_s[44]), .CK(clk), .Q(fracta[44])
         );
  DFF_X2 u1_fracta_out_reg_45_ ( .D(u1_fracta_s[45]), .CK(clk), .Q(fracta[45])
         );
  DFF_X2 u1_fracta_out_reg_46_ ( .D(u1_fracta_s[46]), .CK(clk), .Q(fracta[46])
         );
  DFF_X2 u1_fracta_out_reg_47_ ( .D(u1_fracta_s[47]), .CK(clk), .Q(fracta[47])
         );
  DFF_X2 u1_fracta_out_reg_48_ ( .D(u1_fracta_s[48]), .CK(clk), .Q(fracta[48])
         );
  DFF_X2 u1_fracta_out_reg_49_ ( .D(u1_fracta_s[49]), .CK(clk), .Q(fracta[49])
         );
  DFF_X2 u1_fracta_out_reg_50_ ( .D(u1_fracta_s[50]), .CK(clk), .Q(fracta[50])
         );
  DFF_X2 u1_fracta_out_reg_51_ ( .D(u1_fracta_s[51]), .CK(clk), .Q(fracta[51])
         );
  DFF_X2 u1_fracta_out_reg_52_ ( .D(u1_fracta_s[52]), .CK(clk), .Q(fracta[52])
         );
  DFF_X2 u1_fracta_out_reg_53_ ( .D(u1_fracta_s[53]), .CK(clk), .Q(fracta[53])
         );
  DFF_X2 u1_fracta_out_reg_54_ ( .D(u1_fracta_s[54]), .CK(clk), .Q(fracta[54])
         );
  DFF_X2 u1_fracta_out_reg_55_ ( .D(u1_fracta_s[55]), .CK(clk), .Q(fracta[55])
         );
  DFF_X2 fract_out_q_reg_0_ ( .D(n8355), .CK(clk), .Q(fract_out_q[0]) );
  DFF_X2 fract_out_q_reg_1_ ( .D(n8354), .CK(clk), .Q(fract_out_q[1]) );
  DFF_X2 fract_out_q_reg_2_ ( .D(n8353), .CK(clk), .Q(fract_out_q[2]) );
  DFF_X2 fract_out_q_reg_3_ ( .D(n8352), .CK(clk), .Q(fract_out_q[3]) );
  DFF_X2 fract_out_q_reg_4_ ( .D(n8351), .CK(clk), .Q(fract_out_q[4]) );
  DFF_X2 fract_out_q_reg_5_ ( .D(n8350), .CK(clk), .Q(fract_out_q[5]) );
  DFF_X2 fract_out_q_reg_6_ ( .D(n8349), .CK(clk), .Q(fract_out_q[6]) );
  DFF_X2 fract_out_q_reg_7_ ( .D(n8348), .CK(clk), .Q(fract_out_q[7]) );
  DFF_X2 fract_out_q_reg_8_ ( .D(n8347), .CK(clk), .Q(fract_out_q[8]) );
  DFF_X2 fract_out_q_reg_9_ ( .D(n8346), .CK(clk), .Q(fract_out_q[9]) );
  DFF_X2 fract_out_q_reg_10_ ( .D(n8345), .CK(clk), .Q(fract_out_q[10]) );
  DFF_X2 fract_out_q_reg_11_ ( .D(n8344), .CK(clk), .Q(fract_out_q[11]) );
  DFF_X2 fract_out_q_reg_12_ ( .D(n8343), .CK(clk), .Q(fract_out_q[12]) );
  DFF_X2 fract_out_q_reg_13_ ( .D(n8342), .CK(clk), .Q(fract_out_q[13]) );
  DFF_X2 fract_out_q_reg_14_ ( .D(n8341), .CK(clk), .Q(fract_out_q[14]) );
  DFF_X2 fract_out_q_reg_15_ ( .D(n8340), .CK(clk), .Q(fract_out_q[15]) );
  DFF_X2 fract_out_q_reg_16_ ( .D(n8339), .CK(clk), .Q(fract_out_q[16]) );
  DFF_X2 fract_out_q_reg_17_ ( .D(n8338), .CK(clk), .Q(fract_out_q[17]) );
  DFF_X2 fract_out_q_reg_18_ ( .D(n8337), .CK(clk), .Q(fract_out_q[18]) );
  DFF_X2 fract_out_q_reg_19_ ( .D(n8336), .CK(clk), .Q(fract_out_q[19]) );
  DFF_X2 fract_out_q_reg_20_ ( .D(n8335), .CK(clk), .Q(fract_out_q[20]) );
  DFF_X2 fract_out_q_reg_21_ ( .D(n8334), .CK(clk), .Q(fract_out_q[21]) );
  DFF_X2 fract_out_q_reg_22_ ( .D(n8333), .CK(clk), .Q(fract_out_q[22]) );
  DFF_X2 fract_out_q_reg_23_ ( .D(n8332), .CK(clk), .Q(fract_out_q[23]) );
  DFF_X2 fract_out_q_reg_24_ ( .D(n8331), .CK(clk), .Q(fract_out_q[24]) );
  DFF_X2 fract_out_q_reg_25_ ( .D(n8330), .CK(clk), .Q(fract_out_q[25]) );
  DFF_X2 fract_out_q_reg_26_ ( .D(n8329), .CK(clk), .Q(fract_out_q[26]) );
  DFF_X2 fract_out_q_reg_27_ ( .D(n8328), .CK(clk), .Q(fract_out_q[27]) );
  DFF_X2 fract_out_q_reg_28_ ( .D(n8327), .CK(clk), .Q(fract_out_q[28]) );
  DFF_X2 fract_out_q_reg_29_ ( .D(n8326), .CK(clk), .Q(fract_out_q[29]) );
  DFF_X2 fract_out_q_reg_30_ ( .D(n8325), .CK(clk), .Q(fract_out_q[30]) );
  DFF_X2 fract_out_q_reg_31_ ( .D(n8324), .CK(clk), .Q(fract_out_q[31]) );
  DFF_X2 fract_out_q_reg_32_ ( .D(n8323), .CK(clk), .Q(fract_out_q[32]) );
  DFF_X2 fract_out_q_reg_33_ ( .D(n8322), .CK(clk), .Q(fract_out_q[33]) );
  DFF_X2 fract_out_q_reg_34_ ( .D(n8321), .CK(clk), .Q(fract_out_q[34]) );
  DFF_X2 fract_out_q_reg_35_ ( .D(n8320), .CK(clk), .Q(fract_out_q[35]) );
  DFF_X2 fract_out_q_reg_36_ ( .D(n8319), .CK(clk), .Q(fract_out_q[36]) );
  DFF_X2 fract_out_q_reg_37_ ( .D(n8318), .CK(clk), .Q(fract_out_q[37]) );
  DFF_X2 fract_out_q_reg_38_ ( .D(n8317), .CK(clk), .Q(fract_out_q[38]) );
  DFF_X2 fract_out_q_reg_39_ ( .D(n8316), .CK(clk), .Q(fract_out_q[39]) );
  DFF_X2 fract_out_q_reg_40_ ( .D(n8315), .CK(clk), .Q(fract_out_q[40]) );
  DFF_X2 fract_out_q_reg_41_ ( .D(n8314), .CK(clk), .Q(fract_out_q[41]) );
  DFF_X2 fract_out_q_reg_42_ ( .D(n8313), .CK(clk), .Q(fract_out_q[42]) );
  DFF_X2 fract_out_q_reg_43_ ( .D(n8312), .CK(clk), .Q(fract_out_q[43]) );
  DFF_X2 fract_out_q_reg_44_ ( .D(n8311), .CK(clk), .Q(fract_out_q[44]) );
  DFF_X2 fract_out_q_reg_45_ ( .D(n8310), .CK(clk), .Q(fract_out_q[45]) );
  DFF_X2 fract_out_q_reg_46_ ( .D(n8309), .CK(clk), .Q(fract_out_q[46]) );
  DFF_X2 fract_out_q_reg_47_ ( .D(n8308), .CK(clk), .Q(fract_out_q[47]) );
  DFF_X2 fract_out_q_reg_48_ ( .D(n8307), .CK(clk), .Q(fract_out_q[48]) );
  DFF_X2 fract_out_q_reg_49_ ( .D(n8306), .CK(clk), .Q(fract_out_q[49]) );
  DFF_X2 fract_out_q_reg_50_ ( .D(n8305), .CK(clk), .Q(fract_out_q[50]) );
  DFF_X2 fract_out_q_reg_51_ ( .D(n8304), .CK(clk), .Q(fract_out_q[51]) );
  DFF_X2 fract_out_q_reg_52_ ( .D(n8303), .CK(clk), .Q(fract_out_q[52]) );
  DFF_X2 fract_out_q_reg_53_ ( .D(n8302), .CK(clk), .Q(fract_out_q[53]) );
  DFF_X2 fract_out_q_reg_54_ ( .D(n8301), .CK(clk), .Q(fract_out_q[54]) );
  DFF_X2 fract_out_q_reg_55_ ( .D(n8300), .CK(clk), .Q(fract_out_q[55]) );
  DFF_X2 fract_out_q_reg_56_ ( .D(n8299), .CK(clk), .Q(fract_out_q[56]) );
  DFF_X2 u1_exp_dn_out_reg_0_ ( .D(u1_N52), .CK(clk), .Q(exp_fasu[0]) );
  DFF_X2 u1_exp_dn_out_reg_1_ ( .D(u1_N53), .CK(clk), .Q(exp_fasu[1]) );
  DFF_X2 u1_exp_dn_out_reg_2_ ( .D(u1_N54), .CK(clk), .Q(exp_fasu[2]) );
  DFF_X2 u1_exp_dn_out_reg_3_ ( .D(u1_N55), .CK(clk), .Q(exp_fasu[3]) );
  DFF_X2 u1_exp_dn_out_reg_4_ ( .D(u1_N56), .CK(clk), .Q(exp_fasu[4]) );
  DFF_X2 u1_exp_dn_out_reg_5_ ( .D(u1_N57), .CK(clk), .Q(exp_fasu[5]) );
  DFF_X2 u1_exp_dn_out_reg_6_ ( .D(u1_N58), .CK(clk), .Q(exp_fasu[6]) );
  DFF_X2 u1_exp_dn_out_reg_7_ ( .D(u1_N59), .CK(clk), .Q(exp_fasu[7]) );
  DFF_X2 u1_exp_dn_out_reg_8_ ( .D(u1_N60), .CK(clk), .Q(exp_fasu[8]) );
  DFF_X2 u1_exp_dn_out_reg_9_ ( .D(u1_N61), .CK(clk), .Q(exp_fasu[9]) );
  DFF_X2 u1_exp_dn_out_reg_10_ ( .D(u1_N62), .CK(clk), .Q(exp_fasu[10]) );
  DFF_X2 u2_sign_exe_reg ( .D(u2_N121), .CK(clk), .Q(sign_exe) );
  DFF_X2 sign_exe_r_reg ( .D(sign_exe), .CK(clk), .Q(sign_exe_r) );
  DFF_X2 u2_sign_reg ( .D(u2_sign_d), .CK(clk), .Q(sign_mul), .QN(n4481) );
  DFF_X2 sign_mul_r_reg ( .D(sign_mul), .CK(clk), .Q(sign_mul_r) );
  DFF_X2 sign_reg ( .D(N789), .CK(clk), .Q(sign), .QN(n4462) );
  DFF_X2 fract_i2f_reg_105_ ( .D(N769), .CK(clk), .QN(n4375) );
  DFF_X2 fract_i2f_reg_104_ ( .D(N768), .CK(clk), .Q(fract_i2f[104]) );
  DFF_X2 fract_i2f_reg_103_ ( .D(N767), .CK(clk), .Q(fract_i2f[103]) );
  DFF_X2 fract_i2f_reg_102_ ( .D(N766), .CK(clk), .Q(fract_i2f[102]) );
  DFF_X2 fract_i2f_reg_101_ ( .D(N765), .CK(clk), .Q(fract_i2f[101]) );
  DFF_X2 fract_i2f_reg_100_ ( .D(N764), .CK(clk), .Q(fract_i2f[100]) );
  DFF_X2 fract_i2f_reg_99_ ( .D(N763), .CK(clk), .Q(fract_i2f[99]) );
  DFF_X2 fract_i2f_reg_98_ ( .D(N762), .CK(clk), .Q(fract_i2f[98]) );
  DFF_X2 fract_i2f_reg_97_ ( .D(N761), .CK(clk), .Q(fract_i2f[97]) );
  DFF_X2 fract_i2f_reg_96_ ( .D(N760), .CK(clk), .Q(fract_i2f[96]) );
  DFF_X2 fract_i2f_reg_95_ ( .D(N759), .CK(clk), .Q(fract_i2f[95]) );
  DFF_X2 fract_i2f_reg_94_ ( .D(N758), .CK(clk), .Q(fract_i2f[94]) );
  DFF_X2 fract_i2f_reg_93_ ( .D(N757), .CK(clk), .Q(fract_i2f[93]) );
  DFF_X2 fract_i2f_reg_92_ ( .D(N756), .CK(clk), .Q(fract_i2f[92]) );
  DFF_X2 fract_i2f_reg_91_ ( .D(N755), .CK(clk), .Q(fract_i2f[91]) );
  DFF_X2 fract_i2f_reg_90_ ( .D(N754), .CK(clk), .Q(fract_i2f[90]) );
  DFF_X2 fract_i2f_reg_89_ ( .D(N753), .CK(clk), .Q(fract_i2f[89]) );
  DFF_X2 fract_i2f_reg_88_ ( .D(N752), .CK(clk), .Q(fract_i2f[88]) );
  DFF_X2 fract_i2f_reg_87_ ( .D(N751), .CK(clk), .Q(fract_i2f[87]) );
  DFF_X2 fract_i2f_reg_86_ ( .D(N750), .CK(clk), .Q(fract_i2f[86]) );
  DFF_X2 fract_i2f_reg_85_ ( .D(N749), .CK(clk), .Q(fract_i2f[85]) );
  DFF_X2 fract_i2f_reg_84_ ( .D(N748), .CK(clk), .Q(fract_i2f[84]) );
  DFF_X2 fract_i2f_reg_83_ ( .D(N747), .CK(clk), .Q(fract_i2f[83]) );
  DFF_X2 fract_i2f_reg_82_ ( .D(N746), .CK(clk), .Q(fract_i2f[82]) );
  DFF_X2 fract_i2f_reg_81_ ( .D(N745), .CK(clk), .Q(fract_i2f[81]) );
  DFF_X2 fract_i2f_reg_80_ ( .D(N744), .CK(clk), .Q(fract_i2f[80]) );
  DFF_X2 fract_i2f_reg_79_ ( .D(N743), .CK(clk), .Q(fract_i2f[79]) );
  DFF_X2 fract_i2f_reg_78_ ( .D(N742), .CK(clk), .Q(fract_i2f[78]) );
  DFF_X2 fract_i2f_reg_77_ ( .D(N741), .CK(clk), .Q(fract_i2f[77]) );
  DFF_X2 fract_i2f_reg_76_ ( .D(N740), .CK(clk), .Q(fract_i2f[76]) );
  DFF_X2 fract_i2f_reg_75_ ( .D(N739), .CK(clk), .Q(fract_i2f[75]) );
  DFF_X2 fract_i2f_reg_74_ ( .D(N738), .CK(clk), .Q(fract_i2f[74]) );
  DFF_X2 fract_i2f_reg_73_ ( .D(N737), .CK(clk), .Q(fract_i2f[73]) );
  DFF_X2 fract_i2f_reg_72_ ( .D(N736), .CK(clk), .Q(fract_i2f[72]) );
  DFF_X2 fract_i2f_reg_71_ ( .D(N735), .CK(clk), .Q(fract_i2f[71]) );
  DFF_X2 fract_i2f_reg_70_ ( .D(N734), .CK(clk), .Q(fract_i2f[70]) );
  DFF_X2 fract_i2f_reg_69_ ( .D(N733), .CK(clk), .Q(fract_i2f[69]) );
  DFF_X2 fract_i2f_reg_68_ ( .D(N732), .CK(clk), .Q(fract_i2f[68]) );
  DFF_X2 fract_i2f_reg_67_ ( .D(N731), .CK(clk), .Q(fract_i2f[67]) );
  DFF_X2 fract_i2f_reg_66_ ( .D(N730), .CK(clk), .Q(fract_i2f[66]) );
  DFF_X2 fract_i2f_reg_65_ ( .D(N729), .CK(clk), .Q(fract_i2f[65]) );
  DFF_X2 fract_i2f_reg_64_ ( .D(N728), .CK(clk), .Q(fract_i2f[64]) );
  DFF_X2 fract_i2f_reg_63_ ( .D(N727), .CK(clk), .Q(fract_i2f[63]) );
  DFF_X2 fract_i2f_reg_62_ ( .D(N726), .CK(clk), .Q(fract_i2f[62]) );
  DFF_X2 fract_i2f_reg_61_ ( .D(N725), .CK(clk), .Q(fract_i2f[61]) );
  DFF_X2 fract_i2f_reg_60_ ( .D(N724), .CK(clk), .Q(fract_i2f[60]) );
  DFF_X2 fract_i2f_reg_59_ ( .D(N723), .CK(clk), .Q(fract_i2f[59]) );
  DFF_X2 fract_i2f_reg_58_ ( .D(N722), .CK(clk), .Q(fract_i2f[58]) );
  DFF_X2 fract_i2f_reg_57_ ( .D(N721), .CK(clk), .Q(fract_i2f[57]) );
  DFF_X2 fract_i2f_reg_56_ ( .D(N720), .CK(clk), .Q(fract_i2f[56]) );
  DFF_X2 fract_i2f_reg_55_ ( .D(N719), .CK(clk), .Q(fract_i2f[55]) );
  DFF_X2 fract_i2f_reg_54_ ( .D(N718), .CK(clk), .Q(fract_i2f[54]) );
  DFF_X2 fract_i2f_reg_53_ ( .D(N717), .CK(clk), .Q(fract_i2f[53]) );
  DFF_X2 fract_i2f_reg_52_ ( .D(N716), .CK(clk), .Q(fract_i2f[52]) );
  DFF_X2 fract_i2f_reg_51_ ( .D(N715), .CK(clk), .Q(fract_i2f[51]) );
  DFF_X2 fract_i2f_reg_50_ ( .D(N714), .CK(clk), .Q(fract_i2f[50]) );
  DFF_X2 fract_i2f_reg_49_ ( .D(N713), .CK(clk), .Q(fract_i2f[49]) );
  DFF_X2 fract_i2f_reg_48_ ( .D(N712), .CK(clk), .Q(fract_i2f[48]) );
  DFF_X2 fract_i2f_reg_47_ ( .D(N711), .CK(clk), .Q(fract_i2f[47]) );
  DFF_X2 fract_i2f_reg_46_ ( .D(N710), .CK(clk), .Q(fract_i2f[46]) );
  DFF_X2 fract_i2f_reg_45_ ( .D(n8245), .CK(clk), .Q(fract_i2f[45]) );
  DFF_X2 fract_i2f_reg_44_ ( .D(n8246), .CK(clk), .Q(fract_i2f[44]) );
  DFF_X2 fract_i2f_reg_43_ ( .D(n8247), .CK(clk), .Q(fract_i2f[43]) );
  DFF_X2 fract_i2f_reg_42_ ( .D(n8248), .CK(clk), .Q(fract_i2f[42]) );
  DFF_X2 fract_i2f_reg_41_ ( .D(n8249), .CK(clk), .Q(fract_i2f[41]) );
  DFF_X2 fract_i2f_reg_40_ ( .D(n8250), .CK(clk), .Q(fract_i2f[40]) );
  DFF_X2 fract_i2f_reg_39_ ( .D(n8251), .CK(clk), .Q(fract_i2f[39]) );
  DFF_X2 fract_i2f_reg_38_ ( .D(n8252), .CK(clk), .Q(fract_i2f[38]) );
  DFF_X2 fract_i2f_reg_37_ ( .D(n8253), .CK(clk), .Q(fract_i2f[37]) );
  DFF_X2 fract_i2f_reg_36_ ( .D(n8254), .CK(clk), .Q(fract_i2f[36]) );
  DFF_X2 fract_i2f_reg_35_ ( .D(n8255), .CK(clk), .Q(fract_i2f[35]) );
  DFF_X2 fract_i2f_reg_34_ ( .D(n8256), .CK(clk), .Q(fract_i2f[34]) );
  DFF_X2 fract_i2f_reg_33_ ( .D(n8257), .CK(clk), .Q(fract_i2f[33]) );
  DFF_X2 fract_i2f_reg_32_ ( .D(n8258), .CK(clk), .Q(fract_i2f[32]) );
  DFF_X2 fract_i2f_reg_31_ ( .D(n8259), .CK(clk), .Q(fract_i2f[31]) );
  DFF_X2 fract_i2f_reg_30_ ( .D(n8260), .CK(clk), .Q(fract_i2f[30]) );
  DFF_X2 fract_i2f_reg_29_ ( .D(n8261), .CK(clk), .Q(fract_i2f[29]) );
  DFF_X2 fract_i2f_reg_28_ ( .D(n8262), .CK(clk), .Q(fract_i2f[28]) );
  DFF_X2 fract_i2f_reg_27_ ( .D(n8263), .CK(clk), .Q(fract_i2f[27]) );
  DFF_X2 fract_i2f_reg_26_ ( .D(n8264), .CK(clk), .Q(fract_i2f[26]) );
  DFF_X2 fract_i2f_reg_25_ ( .D(n8265), .CK(clk), .Q(fract_i2f[25]) );
  DFF_X2 fract_i2f_reg_24_ ( .D(n8266), .CK(clk), .Q(fract_i2f[24]) );
  DFF_X2 fract_i2f_reg_23_ ( .D(n8267), .CK(clk), .Q(fract_i2f[23]) );
  DFF_X2 fract_i2f_reg_22_ ( .D(n8268), .CK(clk), .Q(fract_i2f[22]) );
  DFF_X2 fract_i2f_reg_21_ ( .D(n8269), .CK(clk), .Q(fract_i2f[21]) );
  DFF_X2 fract_i2f_reg_20_ ( .D(n8270), .CK(clk), .Q(fract_i2f[20]) );
  DFF_X2 fract_i2f_reg_19_ ( .D(n8271), .CK(clk), .Q(fract_i2f[19]) );
  DFF_X2 fract_i2f_reg_18_ ( .D(n8272), .CK(clk), .Q(fract_i2f[18]) );
  DFF_X2 fract_i2f_reg_17_ ( .D(n8273), .CK(clk), .Q(fract_i2f[17]) );
  DFF_X2 fract_i2f_reg_16_ ( .D(n8274), .CK(clk), .Q(fract_i2f[16]) );
  DFF_X2 fract_i2f_reg_15_ ( .D(n8275), .CK(clk), .Q(fract_i2f[15]) );
  DFF_X2 fract_i2f_reg_14_ ( .D(n8276), .CK(clk), .Q(fract_i2f[14]) );
  DFF_X2 fract_i2f_reg_13_ ( .D(n8277), .CK(clk), .Q(fract_i2f[13]) );
  DFF_X2 fract_i2f_reg_12_ ( .D(n8278), .CK(clk), .Q(fract_i2f[12]) );
  DFF_X2 fract_i2f_reg_11_ ( .D(n8279), .CK(clk), .Q(fract_i2f[11]) );
  DFF_X2 fract_i2f_reg_10_ ( .D(n8280), .CK(clk), .Q(fract_i2f[10]) );
  DFF_X2 fract_i2f_reg_9_ ( .D(n8281), .CK(clk), .Q(fract_i2f[9]) );
  DFF_X2 fract_i2f_reg_8_ ( .D(n8282), .CK(clk), .Q(fract_i2f[8]) );
  DFF_X2 fract_i2f_reg_7_ ( .D(n8283), .CK(clk), .Q(fract_i2f[7]) );
  DFF_X2 fract_i2f_reg_6_ ( .D(n8284), .CK(clk), .Q(fract_i2f[6]) );
  DFF_X2 fract_i2f_reg_5_ ( .D(n8285), .CK(clk), .Q(fract_i2f[5]) );
  DFF_X2 fract_i2f_reg_4_ ( .D(n8286), .CK(clk), .Q(fract_i2f[4]) );
  DFF_X2 fract_i2f_reg_3_ ( .D(n8287), .CK(clk), .Q(fract_i2f[3]) );
  DFF_X2 fract_i2f_reg_2_ ( .D(n8288), .CK(clk), .Q(fract_i2f[2]) );
  DFF_X2 fract_i2f_reg_1_ ( .D(n8289), .CK(clk), .Q(fract_i2f[1]) );
  DFF_X2 fract_i2f_reg_0_ ( .D(n8509), .CK(clk), .Q(fract_i2f[0]) );
  DFF_X2 u2_inf_reg ( .D(u2_N114), .CK(clk), .Q(inf_mul) );
  DFF_X2 inf_mul_r_reg ( .D(inf_mul), .CK(clk), .QN(n4353) );
  DFF_X2 u2_underflow_reg_0_ ( .D(n4487), .CK(clk), .Q(underflow_fmul_d[0]) );
  DFF_X2 underflow_fmul_r_reg_0_ ( .D(underflow_fmul_d[0]), .CK(clk), .Q(
        underflow_fmul_r[0]) );
  DFF_X2 u2_underflow_reg_1_ ( .D(u2_underflow_d[1]), .CK(clk), .Q(
        underflow_fmul_d[1]) );
  DFF_X2 underflow_fmul_r_reg_1_ ( .D(underflow_fmul_d[1]), .CK(clk), .Q(
        underflow_fmul_r[1]) );
  DFF_X2 u2_underflow_reg_2_ ( .D(u2_underflow_d[2]), .CK(clk), .Q(
        underflow_fmul_d[2]) );
  DFF_X2 underflow_fmul_r_reg_2_ ( .D(underflow_fmul_d[2]), .CK(clk), .Q(
        underflow_fmul_r[2]) );
  DFF_X2 u2_exp_ovf_reg_0_ ( .D(u2_exp_ovf_d_0_), .CK(clk), .Q(exp_ovf[0]) );
  DFF_X2 exp_ovf_r_reg_0_ ( .D(exp_ovf[0]), .CK(clk), .Q(exp_ovf_r_0_), .QN(
        n4404) );
  DFF_X2 u2_exp_ovf_reg_1_ ( .D(u2_exp_ovf_d_1_), .CK(clk), .Q(exp_ovf[1]) );
  DFF_X2 exp_ovf_r_reg_1_ ( .D(exp_ovf[1]), .CK(clk), .QN(n4388) );
  DFF_X2 exp_r_reg_0_ ( .D(N327), .CK(clk), .QN(n4326) );
  DFF_X2 exp_r_reg_1_ ( .D(N328), .CK(clk), .QN(n4379) );
  DFF_X2 exp_r_reg_2_ ( .D(N329), .CK(clk), .QN(n4378) );
  DFF_X2 exp_r_reg_3_ ( .D(N330), .CK(clk), .Q(exp_r[3]), .QN(n4308) );
  DFF_X2 exp_r_reg_4_ ( .D(N331), .CK(clk), .Q(exp_r[4]), .QN(n4328) );
  DFF_X2 exp_r_reg_5_ ( .D(N332), .CK(clk), .Q(exp_r[5]), .QN(n4327) );
  DFF_X2 exp_r_reg_6_ ( .D(N333), .CK(clk), .Q(exp_r[6]), .QN(n4384) );
  DFF_X2 exp_r_reg_7_ ( .D(N334), .CK(clk), .QN(n4307) );
  DFF_X2 exp_r_reg_8_ ( .D(N335), .CK(clk), .QN(n4383) );
  DFF_X2 exp_r_reg_9_ ( .D(N336), .CK(clk), .Q(exp_r[9]), .QN(n4505) );
  DFF_X2 inf_mul2_reg ( .D(N923), .CK(clk), .QN(n4483) );
  DFF_X2 exp_r_reg_10_ ( .D(N337), .CK(clk), .QN(n4306) );
  DFF_X2 u5_prod1_reg_0_ ( .D(u5_N0), .CK(clk), .Q(u5_prod1[0]) );
  DFF_X2 u5_prod_reg_0_ ( .D(u5_prod1[0]), .CK(clk), .Q(prod[0]) );
  DFF_X2 u5_prod1_reg_1_ ( .D(u5_N1), .CK(clk), .Q(u5_prod1[1]) );
  DFF_X2 u5_prod_reg_1_ ( .D(u5_prod1[1]), .CK(clk), .Q(prod[1]) );
  DFF_X2 u5_prod1_reg_2_ ( .D(u5_N2), .CK(clk), .Q(u5_prod1[2]) );
  DFF_X2 u5_prod_reg_2_ ( .D(u5_prod1[2]), .CK(clk), .Q(prod[2]) );
  DFF_X2 u5_prod1_reg_3_ ( .D(u5_N3), .CK(clk), .Q(u5_prod1[3]) );
  DFF_X2 u5_prod_reg_3_ ( .D(u5_prod1[3]), .CK(clk), .Q(prod[3]) );
  DFF_X2 u5_prod1_reg_4_ ( .D(u5_N4), .CK(clk), .Q(u5_prod1[4]) );
  DFF_X2 u5_prod_reg_4_ ( .D(u5_prod1[4]), .CK(clk), .Q(prod[4]) );
  DFF_X2 u5_prod1_reg_5_ ( .D(u5_N5), .CK(clk), .Q(u5_prod1[5]) );
  DFF_X2 u5_prod_reg_5_ ( .D(u5_prod1[5]), .CK(clk), .Q(prod[5]) );
  DFF_X2 u5_prod1_reg_6_ ( .D(u5_N6), .CK(clk), .Q(u5_prod1[6]) );
  DFF_X2 u5_prod_reg_6_ ( .D(u5_prod1[6]), .CK(clk), .Q(prod[6]) );
  DFF_X2 u5_prod1_reg_7_ ( .D(u5_N7), .CK(clk), .Q(u5_prod1[7]) );
  DFF_X2 u5_prod_reg_7_ ( .D(u5_prod1[7]), .CK(clk), .Q(prod[7]) );
  DFF_X2 u5_prod1_reg_8_ ( .D(u5_N8), .CK(clk), .Q(u5_prod1[8]) );
  DFF_X2 u5_prod_reg_8_ ( .D(u5_prod1[8]), .CK(clk), .Q(prod[8]) );
  DFF_X2 u5_prod1_reg_9_ ( .D(u5_N9), .CK(clk), .Q(u5_prod1[9]) );
  DFF_X2 u5_prod_reg_9_ ( .D(u5_prod1[9]), .CK(clk), .Q(prod[9]) );
  DFF_X2 u5_prod1_reg_10_ ( .D(u5_N10), .CK(clk), .Q(u5_prod1[10]) );
  DFF_X2 u5_prod_reg_10_ ( .D(u5_prod1[10]), .CK(clk), .Q(prod[10]) );
  DFF_X2 u5_prod1_reg_11_ ( .D(u5_N11), .CK(clk), .Q(u5_prod1[11]) );
  DFF_X2 u5_prod_reg_11_ ( .D(u5_prod1[11]), .CK(clk), .Q(prod[11]) );
  DFF_X2 u5_prod1_reg_12_ ( .D(u5_N12), .CK(clk), .Q(u5_prod1[12]) );
  DFF_X2 u5_prod_reg_12_ ( .D(u5_prod1[12]), .CK(clk), .Q(prod[12]) );
  DFF_X2 u5_prod1_reg_13_ ( .D(u5_N13), .CK(clk), .Q(u5_prod1[13]) );
  DFF_X2 u5_prod_reg_13_ ( .D(u5_prod1[13]), .CK(clk), .Q(prod[13]) );
  DFF_X2 u5_prod1_reg_14_ ( .D(u5_N14), .CK(clk), .Q(u5_prod1[14]) );
  DFF_X2 u5_prod_reg_14_ ( .D(u5_prod1[14]), .CK(clk), .Q(prod[14]) );
  DFF_X2 u5_prod1_reg_15_ ( .D(u5_N15), .CK(clk), .Q(u5_prod1[15]) );
  DFF_X2 u5_prod_reg_15_ ( .D(u5_prod1[15]), .CK(clk), .Q(prod[15]) );
  DFF_X2 u5_prod1_reg_16_ ( .D(u5_N16), .CK(clk), .Q(u5_prod1[16]) );
  DFF_X2 u5_prod_reg_16_ ( .D(u5_prod1[16]), .CK(clk), .Q(prod[16]) );
  DFF_X2 u5_prod1_reg_17_ ( .D(u5_N17), .CK(clk), .Q(u5_prod1[17]) );
  DFF_X2 u5_prod_reg_17_ ( .D(u5_prod1[17]), .CK(clk), .Q(prod[17]) );
  DFF_X2 u5_prod1_reg_18_ ( .D(u5_N18), .CK(clk), .Q(u5_prod1[18]) );
  DFF_X2 u5_prod_reg_18_ ( .D(u5_prod1[18]), .CK(clk), .Q(prod[18]) );
  DFF_X2 u5_prod1_reg_19_ ( .D(u5_N19), .CK(clk), .Q(u5_prod1[19]) );
  DFF_X2 u5_prod_reg_19_ ( .D(u5_prod1[19]), .CK(clk), .Q(prod[19]) );
  DFF_X2 u5_prod1_reg_20_ ( .D(u5_N20), .CK(clk), .Q(u5_prod1[20]) );
  DFF_X2 u5_prod_reg_20_ ( .D(u5_prod1[20]), .CK(clk), .Q(prod[20]) );
  DFF_X2 u5_prod1_reg_21_ ( .D(u5_N21), .CK(clk), .Q(u5_prod1[21]) );
  DFF_X2 u5_prod_reg_21_ ( .D(u5_prod1[21]), .CK(clk), .Q(prod[21]) );
  DFF_X2 u5_prod1_reg_22_ ( .D(u5_N22), .CK(clk), .Q(u5_prod1[22]) );
  DFF_X2 u5_prod_reg_22_ ( .D(u5_prod1[22]), .CK(clk), .Q(prod[22]) );
  DFF_X2 u5_prod1_reg_23_ ( .D(u5_N23), .CK(clk), .Q(u5_prod1[23]) );
  DFF_X2 u5_prod_reg_23_ ( .D(u5_prod1[23]), .CK(clk), .Q(prod[23]) );
  DFF_X2 u5_prod1_reg_24_ ( .D(u5_N24), .CK(clk), .Q(u5_prod1[24]) );
  DFF_X2 u5_prod_reg_24_ ( .D(u5_prod1[24]), .CK(clk), .Q(prod[24]) );
  DFF_X2 u5_prod1_reg_25_ ( .D(u5_N25), .CK(clk), .Q(u5_prod1[25]) );
  DFF_X2 u5_prod_reg_25_ ( .D(u5_prod1[25]), .CK(clk), .Q(prod[25]) );
  DFF_X2 u5_prod1_reg_26_ ( .D(u5_N26), .CK(clk), .Q(u5_prod1[26]) );
  DFF_X2 u5_prod_reg_26_ ( .D(u5_prod1[26]), .CK(clk), .Q(prod[26]) );
  DFF_X2 u5_prod1_reg_27_ ( .D(u5_N27), .CK(clk), .Q(u5_prod1[27]) );
  DFF_X2 u5_prod_reg_27_ ( .D(u5_prod1[27]), .CK(clk), .Q(prod[27]) );
  DFF_X2 u5_prod1_reg_28_ ( .D(u5_N28), .CK(clk), .Q(u5_prod1[28]) );
  DFF_X2 u5_prod_reg_28_ ( .D(u5_prod1[28]), .CK(clk), .Q(prod[28]) );
  DFF_X2 u5_prod1_reg_29_ ( .D(u5_N29), .CK(clk), .Q(u5_prod1[29]) );
  DFF_X2 u5_prod_reg_29_ ( .D(u5_prod1[29]), .CK(clk), .Q(prod[29]) );
  DFF_X2 u5_prod1_reg_30_ ( .D(u5_N30), .CK(clk), .Q(u5_prod1[30]) );
  DFF_X2 u5_prod_reg_30_ ( .D(u5_prod1[30]), .CK(clk), .Q(prod[30]) );
  DFF_X2 u5_prod1_reg_31_ ( .D(u5_N31), .CK(clk), .Q(u5_prod1[31]) );
  DFF_X2 u5_prod_reg_31_ ( .D(u5_prod1[31]), .CK(clk), .Q(prod[31]) );
  DFF_X2 u5_prod1_reg_32_ ( .D(u5_N32), .CK(clk), .Q(u5_prod1[32]) );
  DFF_X2 u5_prod_reg_32_ ( .D(u5_prod1[32]), .CK(clk), .Q(prod[32]) );
  DFF_X2 u5_prod1_reg_33_ ( .D(u5_N33), .CK(clk), .Q(u5_prod1[33]) );
  DFF_X2 u5_prod_reg_33_ ( .D(u5_prod1[33]), .CK(clk), .Q(prod[33]) );
  DFF_X2 u5_prod1_reg_34_ ( .D(u5_N34), .CK(clk), .Q(u5_prod1[34]) );
  DFF_X2 u5_prod_reg_34_ ( .D(u5_prod1[34]), .CK(clk), .Q(prod[34]) );
  DFF_X2 u5_prod1_reg_35_ ( .D(u5_N35), .CK(clk), .Q(u5_prod1[35]) );
  DFF_X2 u5_prod_reg_35_ ( .D(u5_prod1[35]), .CK(clk), .Q(prod[35]) );
  DFF_X2 u5_prod1_reg_36_ ( .D(u5_N36), .CK(clk), .Q(u5_prod1[36]) );
  DFF_X2 u5_prod_reg_36_ ( .D(u5_prod1[36]), .CK(clk), .Q(prod[36]) );
  DFF_X2 u5_prod1_reg_37_ ( .D(u5_N37), .CK(clk), .Q(u5_prod1[37]) );
  DFF_X2 u5_prod_reg_37_ ( .D(u5_prod1[37]), .CK(clk), .Q(prod[37]) );
  DFF_X2 u5_prod1_reg_38_ ( .D(u5_N38), .CK(clk), .Q(u5_prod1[38]) );
  DFF_X2 u5_prod_reg_38_ ( .D(u5_prod1[38]), .CK(clk), .Q(prod[38]) );
  DFF_X2 u5_prod1_reg_39_ ( .D(u5_N39), .CK(clk), .Q(u5_prod1[39]) );
  DFF_X2 u5_prod_reg_39_ ( .D(u5_prod1[39]), .CK(clk), .Q(prod[39]) );
  DFF_X2 u5_prod1_reg_40_ ( .D(u5_N40), .CK(clk), .Q(u5_prod1[40]) );
  DFF_X2 u5_prod_reg_40_ ( .D(u5_prod1[40]), .CK(clk), .Q(prod[40]) );
  DFF_X2 u5_prod1_reg_41_ ( .D(u5_N41), .CK(clk), .Q(u5_prod1[41]) );
  DFF_X2 u5_prod_reg_41_ ( .D(u5_prod1[41]), .CK(clk), .Q(prod[41]) );
  DFF_X2 u5_prod1_reg_42_ ( .D(u5_N42), .CK(clk), .Q(u5_prod1[42]) );
  DFF_X2 u5_prod_reg_42_ ( .D(u5_prod1[42]), .CK(clk), .Q(prod[42]) );
  DFF_X2 u5_prod1_reg_43_ ( .D(u5_N43), .CK(clk), .Q(u5_prod1[43]) );
  DFF_X2 u5_prod_reg_43_ ( .D(u5_prod1[43]), .CK(clk), .Q(prod[43]) );
  DFF_X2 u5_prod1_reg_44_ ( .D(u5_N44), .CK(clk), .Q(u5_prod1[44]) );
  DFF_X2 u5_prod_reg_44_ ( .D(u5_prod1[44]), .CK(clk), .Q(prod[44]) );
  DFF_X2 u5_prod1_reg_45_ ( .D(u5_N45), .CK(clk), .Q(u5_prod1[45]) );
  DFF_X2 u5_prod_reg_45_ ( .D(u5_prod1[45]), .CK(clk), .Q(prod[45]) );
  DFF_X2 u5_prod_reg_46_ ( .D(u5_prod1[46]), .CK(clk), .Q(prod[46]) );
  DFF_X2 u5_prod_reg_47_ ( .D(u5_prod1[47]), .CK(clk), .Q(prod[47]) );
  DFF_X2 u5_prod1_reg_48_ ( .D(u5_N48), .CK(clk), .Q(u5_prod1[48]) );
  DFF_X2 u5_prod_reg_48_ ( .D(u5_prod1[48]), .CK(clk), .Q(prod[48]) );
  DFF_X2 u5_prod1_reg_49_ ( .D(u5_N49), .CK(clk), .Q(u5_prod1[49]) );
  DFF_X2 u5_prod_reg_49_ ( .D(u5_prod1[49]), .CK(clk), .Q(prod[49]) );
  DFF_X2 u5_prod1_reg_50_ ( .D(u5_N50), .CK(clk), .Q(u5_prod1[50]) );
  DFF_X2 u5_prod_reg_50_ ( .D(u5_prod1[50]), .CK(clk), .Q(prod[50]) );
  DFF_X2 u5_prod1_reg_51_ ( .D(u5_N51), .CK(clk), .Q(u5_prod1[51]) );
  DFF_X2 u5_prod_reg_51_ ( .D(u5_prod1[51]), .CK(clk), .Q(prod[51]) );
  DFF_X2 u5_prod_reg_52_ ( .D(u5_prod1[52]), .CK(clk), .Q(prod[52]) );
  DFF_X2 u5_prod1_reg_53_ ( .D(u5_N53), .CK(clk), .Q(u5_prod1[53]) );
  DFF_X2 u5_prod_reg_53_ ( .D(u5_prod1[53]), .CK(clk), .Q(prod[53]) );
  DFF_X2 u5_prod1_reg_54_ ( .D(u5_N54), .CK(clk), .Q(u5_prod1[54]) );
  DFF_X2 u5_prod_reg_54_ ( .D(u5_prod1[54]), .CK(clk), .Q(prod[54]) );
  DFF_X2 u5_prod1_reg_55_ ( .D(u5_N55), .CK(clk), .Q(u5_prod1[55]) );
  DFF_X2 u5_prod_reg_55_ ( .D(u5_prod1[55]), .CK(clk), .Q(prod[55]) );
  DFF_X2 u5_prod1_reg_56_ ( .D(u5_N56), .CK(clk), .Q(u5_prod1[56]) );
  DFF_X2 u5_prod_reg_56_ ( .D(u5_prod1[56]), .CK(clk), .Q(prod[56]) );
  DFF_X2 u5_prod1_reg_57_ ( .D(u5_N57), .CK(clk), .Q(u5_prod1[57]) );
  DFF_X2 u5_prod_reg_57_ ( .D(u5_prod1[57]), .CK(clk), .Q(prod[57]) );
  DFF_X2 u5_prod1_reg_58_ ( .D(u5_N58), .CK(clk), .Q(u5_prod1[58]) );
  DFF_X2 u5_prod_reg_58_ ( .D(u5_prod1[58]), .CK(clk), .Q(prod[58]) );
  DFF_X2 u5_prod1_reg_59_ ( .D(u5_N59), .CK(clk), .Q(u5_prod1[59]) );
  DFF_X2 u5_prod_reg_59_ ( .D(u5_prod1[59]), .CK(clk), .Q(prod[59]) );
  DFF_X2 u5_prod1_reg_60_ ( .D(u5_N60), .CK(clk), .Q(u5_prod1[60]) );
  DFF_X2 u5_prod_reg_60_ ( .D(u5_prod1[60]), .CK(clk), .Q(prod[60]) );
  DFF_X2 u5_prod1_reg_61_ ( .D(u5_N61), .CK(clk), .Q(u5_prod1[61]) );
  DFF_X2 u5_prod1_reg_62_ ( .D(u5_N62), .CK(clk), .Q(u5_prod1[62]) );
  DFF_X2 u5_prod_reg_62_ ( .D(u5_prod1[62]), .CK(clk), .Q(prod[62]) );
  DFF_X2 u5_prod1_reg_63_ ( .D(u5_N63), .CK(clk), .Q(u5_prod1[63]) );
  DFF_X2 u5_prod_reg_63_ ( .D(u5_prod1[63]), .CK(clk), .Q(prod[63]) );
  DFF_X2 u5_prod1_reg_64_ ( .D(u5_N64), .CK(clk), .Q(u5_prod1[64]) );
  DFF_X2 u5_prod_reg_64_ ( .D(u5_prod1[64]), .CK(clk), .Q(prod[64]) );
  DFF_X2 u5_prod1_reg_65_ ( .D(u5_N65), .CK(clk), .Q(u5_prod1[65]) );
  DFF_X2 u5_prod_reg_65_ ( .D(u5_prod1[65]), .CK(clk), .Q(prod[65]) );
  DFF_X2 u5_prod1_reg_66_ ( .D(u5_N66), .CK(clk), .Q(u5_prod1[66]) );
  DFF_X2 u5_prod_reg_66_ ( .D(u5_prod1[66]), .CK(clk), .Q(prod[66]) );
  DFF_X2 u5_prod1_reg_67_ ( .D(u5_N67), .CK(clk), .Q(u5_prod1[67]) );
  DFF_X2 u5_prod_reg_67_ ( .D(u5_prod1[67]), .CK(clk), .Q(prod[67]) );
  DFF_X2 u5_prod1_reg_68_ ( .D(u5_N68), .CK(clk), .Q(u5_prod1[68]) );
  DFF_X2 u5_prod1_reg_69_ ( .D(u5_N69), .CK(clk), .Q(u5_prod1[69]) );
  DFF_X2 u5_prod_reg_69_ ( .D(u5_prod1[69]), .CK(clk), .Q(prod[69]) );
  DFF_X2 u5_prod1_reg_70_ ( .D(u5_N70), .CK(clk), .Q(u5_prod1[70]) );
  DFF_X2 u5_prod_reg_70_ ( .D(u5_prod1[70]), .CK(clk), .Q(prod[70]) );
  DFF_X2 u5_prod1_reg_71_ ( .D(u5_N71), .CK(clk), .Q(u5_prod1[71]) );
  DFF_X2 u5_prod_reg_71_ ( .D(u5_prod1[71]), .CK(clk), .Q(prod[71]) );
  DFF_X2 u5_prod1_reg_72_ ( .D(u5_N72), .CK(clk), .Q(u5_prod1[72]) );
  DFF_X2 u5_prod_reg_72_ ( .D(u5_prod1[72]), .CK(clk), .Q(prod[72]) );
  DFF_X2 u5_prod1_reg_73_ ( .D(u5_N73), .CK(clk), .Q(u5_prod1[73]) );
  DFF_X2 u5_prod_reg_73_ ( .D(u5_prod1[73]), .CK(clk), .Q(prod[73]) );
  DFF_X2 u5_prod1_reg_74_ ( .D(u5_N74), .CK(clk), .Q(u5_prod1[74]) );
  DFF_X2 u5_prod_reg_74_ ( .D(u5_prod1[74]), .CK(clk), .Q(prod[74]) );
  DFF_X2 u5_prod1_reg_75_ ( .D(u5_N75), .CK(clk), .Q(u5_prod1[75]) );
  DFF_X2 u5_prod_reg_75_ ( .D(u5_prod1[75]), .CK(clk), .Q(prod[75]) );
  DFF_X2 u5_prod1_reg_76_ ( .D(u5_N76), .CK(clk), .Q(u5_prod1[76]) );
  DFF_X2 u5_prod_reg_76_ ( .D(u5_prod1[76]), .CK(clk), .Q(prod[76]) );
  DFF_X2 u5_prod_reg_77_ ( .D(u5_prod1[77]), .CK(clk), .Q(prod[77]) );
  DFF_X2 u5_prod1_reg_78_ ( .D(u5_N78), .CK(clk), .Q(u5_prod1[78]) );
  DFF_X2 u5_prod_reg_78_ ( .D(u5_prod1[78]), .CK(clk), .Q(prod[78]) );
  DFF_X2 u5_prod1_reg_79_ ( .D(u5_N79), .CK(clk), .Q(u5_prod1[79]) );
  DFF_X2 u5_prod_reg_79_ ( .D(u5_prod1[79]), .CK(clk), .Q(prod[79]) );
  DFF_X2 u5_prod1_reg_80_ ( .D(u5_N80), .CK(clk), .Q(u5_prod1[80]) );
  DFF_X2 u5_prod_reg_80_ ( .D(u5_prod1[80]), .CK(clk), .Q(prod[80]) );
  DFF_X2 u5_prod1_reg_81_ ( .D(u5_N81), .CK(clk), .Q(u5_prod1[81]) );
  DFF_X2 u5_prod_reg_81_ ( .D(u5_prod1[81]), .CK(clk), .Q(prod[81]) );
  DFF_X2 u5_prod1_reg_82_ ( .D(u5_N82), .CK(clk), .Q(u5_prod1[82]) );
  DFF_X2 u5_prod_reg_82_ ( .D(u5_prod1[82]), .CK(clk), .Q(prod[82]) );
  DFF_X2 u5_prod_reg_83_ ( .D(u5_prod1[83]), .CK(clk), .Q(prod[83]) );
  DFF_X2 u5_prod1_reg_84_ ( .D(u5_N84), .CK(clk), .Q(u5_prod1[84]) );
  DFF_X2 u5_prod_reg_84_ ( .D(u5_prod1[84]), .CK(clk), .Q(prod[84]) );
  DFF_X2 u5_prod1_reg_85_ ( .D(u5_N85), .CK(clk), .Q(u5_prod1[85]) );
  DFF_X2 u5_prod_reg_85_ ( .D(u5_prod1[85]), .CK(clk), .Q(prod[85]) );
  DFF_X2 u5_prod_reg_86_ ( .D(u5_prod1[86]), .CK(clk), .Q(prod[86]) );
  DFF_X2 u5_prod_reg_87_ ( .D(u5_prod1[87]), .CK(clk), .Q(prod[87]) );
  DFF_X2 u5_prod1_reg_88_ ( .D(u5_N88), .CK(clk), .Q(u5_prod1[88]) );
  DFF_X2 u5_prod_reg_88_ ( .D(u5_prod1[88]), .CK(clk), .Q(prod[88]) );
  DFF_X2 u5_prod_reg_89_ ( .D(u5_prod1[89]), .CK(clk), .Q(prod[89]) );
  DFF_X2 u5_prod_reg_90_ ( .D(u5_prod1[90]), .CK(clk), .Q(prod[90]) );
  DFF_X2 u5_prod1_reg_91_ ( .D(u5_N91), .CK(clk), .Q(u5_prod1[91]) );
  DFF_X2 u5_prod_reg_91_ ( .D(u5_prod1[91]), .CK(clk), .Q(prod[91]) );
  DFF_X2 u5_prod_reg_92_ ( .D(u5_prod1[92]), .CK(clk), .Q(prod[92]) );
  DFF_X2 u5_prod_reg_93_ ( .D(u5_prod1[93]), .CK(clk), .Q(prod[93]) );
  DFF_X2 u5_prod_reg_94_ ( .D(u5_prod1[94]), .CK(clk), .Q(prod[94]) );
  DFF_X2 u5_prod_reg_95_ ( .D(u5_prod1[95]), .CK(clk), .Q(prod[95]) );
  DFF_X2 u5_prod_reg_96_ ( .D(u5_prod1[96]), .CK(clk), .Q(prod[96]) );
  DFF_X2 u5_prod_reg_97_ ( .D(u5_prod1[97]), .CK(clk), .Q(prod[97]) );
  DFF_X2 u5_prod1_reg_98_ ( .D(u5_N98), .CK(clk), .Q(u5_prod1[98]) );
  DFF_X2 u5_prod_reg_98_ ( .D(u5_prod1[98]), .CK(clk), .Q(prod[98]) );
  DFF_X2 u5_prod_reg_99_ ( .D(u5_prod1[99]), .CK(clk), .Q(prod[99]) );
  DFF_X2 u5_prod_reg_100_ ( .D(u5_prod1[100]), .CK(clk), .Q(prod[100]) );
  DFF_X2 u5_prod_reg_101_ ( .D(u5_prod1[101]), .CK(clk), .Q(prod[101]) );
  DFF_X2 u5_prod1_reg_102_ ( .D(u5_N102), .CK(clk), .Q(u5_prod1[102]) );
  DFF_X2 u5_prod_reg_102_ ( .D(u5_prod1[102]), .CK(clk), .Q(prod[102]) );
  DFF_X2 u5_prod_reg_103_ ( .D(u5_prod1[103]), .CK(clk), .Q(prod[103]) );
  DFF_X2 u5_prod_reg_104_ ( .D(u5_prod1[104]), .CK(clk), .Q(prod[104]) );
  DFF_X2 u5_prod1_reg_105_ ( .D(u5_N105), .CK(clk), .Q(u5_prod1[105]) );
  DFF_X2 u5_prod_reg_105_ ( .D(u5_prod1[105]), .CK(clk), .Q(prod[105]) );
  DFF_X2 u6_remainder_reg_0_ ( .D(u6_N0), .CK(clk), .Q(u6_remainder[0]) );
  DFF_X2 u6_rem_reg_0_ ( .D(u6_remainder[0]), .CK(clk), .Q(remainder[0]) );
  DFF_X2 u6_remainder_reg_1_ ( .D(u6_N1), .CK(clk), .Q(u6_remainder[1]) );
  DFF_X2 u6_rem_reg_1_ ( .D(u6_remainder[1]), .CK(clk), .Q(remainder[1]) );
  DFF_X2 u6_remainder_reg_2_ ( .D(u6_N2), .CK(clk), .Q(u6_remainder[2]) );
  DFF_X2 u6_rem_reg_2_ ( .D(u6_remainder[2]), .CK(clk), .Q(remainder[2]) );
  DFF_X2 u6_remainder_reg_3_ ( .D(u6_N3), .CK(clk), .Q(u6_remainder[3]) );
  DFF_X2 u6_rem_reg_3_ ( .D(u6_remainder[3]), .CK(clk), .Q(remainder[3]) );
  DFF_X2 u6_remainder_reg_4_ ( .D(u6_N4), .CK(clk), .Q(u6_remainder[4]) );
  DFF_X2 u6_rem_reg_4_ ( .D(u6_remainder[4]), .CK(clk), .Q(remainder[4]) );
  DFF_X2 u6_remainder_reg_5_ ( .D(u6_N5), .CK(clk), .Q(u6_remainder[5]) );
  DFF_X2 u6_rem_reg_5_ ( .D(u6_remainder[5]), .CK(clk), .Q(remainder[5]) );
  DFF_X2 u6_remainder_reg_6_ ( .D(u6_N6), .CK(clk), .Q(u6_remainder[6]) );
  DFF_X2 u6_rem_reg_6_ ( .D(u6_remainder[6]), .CK(clk), .QN(n4409) );
  DFF_X2 u6_remainder_reg_7_ ( .D(u6_N7), .CK(clk), .Q(u6_remainder[7]) );
  DFF_X2 u6_rem_reg_7_ ( .D(u6_remainder[7]), .CK(clk), .Q(remainder[7]) );
  DFF_X2 u6_remainder_reg_8_ ( .D(u6_N8), .CK(clk), .Q(u6_remainder[8]) );
  DFF_X2 u6_rem_reg_8_ ( .D(u6_remainder[8]), .CK(clk), .Q(remainder[8]) );
  DFF_X2 u6_remainder_reg_9_ ( .D(u6_N9), .CK(clk), .Q(u6_remainder[9]) );
  DFF_X2 u6_rem_reg_9_ ( .D(u6_remainder[9]), .CK(clk), .Q(remainder[9]) );
  DFF_X2 u6_remainder_reg_10_ ( .D(u6_N10), .CK(clk), .Q(u6_remainder[10]) );
  DFF_X2 u6_rem_reg_10_ ( .D(u6_remainder[10]), .CK(clk), .Q(remainder[10]) );
  DFF_X2 u6_remainder_reg_11_ ( .D(u6_N11), .CK(clk), .Q(u6_remainder[11]) );
  DFF_X2 u6_rem_reg_11_ ( .D(u6_remainder[11]), .CK(clk), .Q(remainder[11]) );
  DFF_X2 u6_remainder_reg_12_ ( .D(u6_N12), .CK(clk), .Q(u6_remainder[12]) );
  DFF_X2 u6_rem_reg_12_ ( .D(u6_remainder[12]), .CK(clk), .Q(remainder[12]) );
  DFF_X2 u6_remainder_reg_13_ ( .D(u6_N13), .CK(clk), .Q(u6_remainder[13]) );
  DFF_X2 u6_rem_reg_13_ ( .D(u6_remainder[13]), .CK(clk), .QN(n4408) );
  DFF_X2 u6_remainder_reg_14_ ( .D(u6_N14), .CK(clk), .Q(u6_remainder[14]) );
  DFF_X2 u6_rem_reg_14_ ( .D(u6_remainder[14]), .CK(clk), .Q(remainder[14]) );
  DFF_X2 u6_remainder_reg_15_ ( .D(u6_N15), .CK(clk), .Q(u6_remainder[15]) );
  DFF_X2 u6_rem_reg_15_ ( .D(u6_remainder[15]), .CK(clk), .Q(remainder[15]) );
  DFF_X2 u6_remainder_reg_16_ ( .D(u6_N16), .CK(clk), .Q(u6_remainder[16]) );
  DFF_X2 u6_rem_reg_16_ ( .D(u6_remainder[16]), .CK(clk), .Q(remainder[16]) );
  DFF_X2 u6_remainder_reg_17_ ( .D(u6_N17), .CK(clk), .Q(u6_remainder[17]) );
  DFF_X2 u6_rem_reg_17_ ( .D(u6_remainder[17]), .CK(clk), .Q(remainder[17]) );
  DFF_X2 u6_remainder_reg_18_ ( .D(u6_N18), .CK(clk), .Q(u6_remainder[18]) );
  DFF_X2 u6_rem_reg_18_ ( .D(u6_remainder[18]), .CK(clk), .Q(remainder[18]) );
  DFF_X2 u6_remainder_reg_19_ ( .D(u6_N19), .CK(clk), .Q(u6_remainder[19]) );
  DFF_X2 u6_rem_reg_19_ ( .D(u6_remainder[19]), .CK(clk), .Q(remainder[19]) );
  DFF_X2 u6_remainder_reg_20_ ( .D(u6_N20), .CK(clk), .Q(u6_remainder[20]) );
  DFF_X2 u6_rem_reg_20_ ( .D(u6_remainder[20]), .CK(clk), .Q(remainder[20]) );
  DFF_X2 u6_remainder_reg_21_ ( .D(u6_N21), .CK(clk), .Q(u6_remainder[21]) );
  DFF_X2 u6_rem_reg_21_ ( .D(u6_remainder[21]), .CK(clk), .Q(remainder[21]) );
  DFF_X2 u6_remainder_reg_22_ ( .D(u6_N22), .CK(clk), .Q(u6_remainder[22]) );
  DFF_X2 u6_rem_reg_22_ ( .D(u6_remainder[22]), .CK(clk), .Q(remainder[22]) );
  DFF_X2 u6_remainder_reg_23_ ( .D(u6_N23), .CK(clk), .Q(u6_remainder[23]) );
  DFF_X2 u6_rem_reg_23_ ( .D(u6_remainder[23]), .CK(clk), .Q(remainder[23]) );
  DFF_X2 u6_remainder_reg_24_ ( .D(u6_N24), .CK(clk), .Q(u6_remainder[24]) );
  DFF_X2 u6_rem_reg_24_ ( .D(u6_remainder[24]), .CK(clk), .Q(remainder[24]) );
  DFF_X2 u6_remainder_reg_25_ ( .D(u6_N25), .CK(clk), .Q(u6_remainder[25]) );
  DFF_X2 u6_rem_reg_25_ ( .D(u6_remainder[25]), .CK(clk), .Q(remainder[25]) );
  DFF_X2 u6_remainder_reg_26_ ( .D(u6_N26), .CK(clk), .Q(u6_remainder[26]) );
  DFF_X2 u6_rem_reg_26_ ( .D(u6_remainder[26]), .CK(clk), .Q(remainder[26]) );
  DFF_X2 u6_remainder_reg_27_ ( .D(u6_N27), .CK(clk), .Q(u6_remainder[27]) );
  DFF_X2 u6_rem_reg_27_ ( .D(u6_remainder[27]), .CK(clk), .Q(remainder[27]) );
  DFF_X2 u6_remainder_reg_28_ ( .D(n4764), .CK(clk), .Q(u6_remainder[28]) );
  DFF_X2 u6_rem_reg_28_ ( .D(u6_remainder[28]), .CK(clk), .Q(remainder[28]) );
  DFF_X2 u6_remainder_reg_29_ ( .D(u6_N29), .CK(clk), .Q(u6_remainder[29]) );
  DFF_X2 u6_rem_reg_29_ ( .D(u6_remainder[29]), .CK(clk), .Q(remainder[29]) );
  DFF_X2 u6_remainder_reg_30_ ( .D(u6_N30), .CK(clk), .Q(u6_remainder[30]) );
  DFF_X2 u6_rem_reg_30_ ( .D(u6_remainder[30]), .CK(clk), .Q(remainder[30]) );
  DFF_X2 u6_remainder_reg_31_ ( .D(u6_N31), .CK(clk), .Q(u6_remainder[31]) );
  DFF_X2 u6_rem_reg_31_ ( .D(u6_remainder[31]), .CK(clk), .Q(remainder[31]) );
  DFF_X2 u6_remainder_reg_32_ ( .D(u6_N32), .CK(clk), .Q(u6_remainder[32]) );
  DFF_X2 u6_rem_reg_32_ ( .D(u6_remainder[32]), .CK(clk), .Q(remainder[32]) );
  DFF_X2 u6_remainder_reg_33_ ( .D(u6_N33), .CK(clk), .Q(u6_remainder[33]) );
  DFF_X2 u6_rem_reg_33_ ( .D(u6_remainder[33]), .CK(clk), .QN(n4411) );
  DFF_X2 u6_remainder_reg_34_ ( .D(n4786), .CK(clk), .Q(u6_remainder[34]) );
  DFF_X2 u6_rem_reg_34_ ( .D(u6_remainder[34]), .CK(clk), .Q(remainder[34]) );
  DFF_X2 u6_remainder_reg_35_ ( .D(u6_N35), .CK(clk), .Q(u6_remainder[35]) );
  DFF_X2 u6_rem_reg_35_ ( .D(u6_remainder[35]), .CK(clk), .Q(remainder[35]) );
  DFF_X2 u6_remainder_reg_36_ ( .D(u6_N36), .CK(clk), .Q(u6_remainder[36]) );
  DFF_X2 u6_rem_reg_36_ ( .D(u6_remainder[36]), .CK(clk), .Q(remainder[36]) );
  DFF_X2 u6_remainder_reg_37_ ( .D(u6_N37), .CK(clk), .Q(u6_remainder[37]) );
  DFF_X2 u6_rem_reg_37_ ( .D(u6_remainder[37]), .CK(clk), .Q(remainder[37]) );
  DFF_X2 u6_remainder_reg_38_ ( .D(n4791), .CK(clk), .Q(u6_remainder[38]) );
  DFF_X2 u6_rem_reg_38_ ( .D(u6_remainder[38]), .CK(clk), .Q(remainder[38]) );
  DFF_X2 u6_remainder_reg_39_ ( .D(u6_N39), .CK(clk), .Q(u6_remainder[39]) );
  DFF_X2 u6_rem_reg_39_ ( .D(u6_remainder[39]), .CK(clk), .Q(remainder[39]) );
  DFF_X2 u6_remainder_reg_40_ ( .D(u6_N40), .CK(clk), .Q(u6_remainder[40]) );
  DFF_X2 u6_rem_reg_40_ ( .D(u6_remainder[40]), .CK(clk), .QN(n4410) );
  DFF_X2 u6_remainder_reg_41_ ( .D(n4772), .CK(clk), .Q(u6_remainder[41]) );
  DFF_X2 u6_rem_reg_41_ ( .D(u6_remainder[41]), .CK(clk), .Q(remainder[41]) );
  DFF_X2 u6_remainder_reg_42_ ( .D(n4787), .CK(clk), .Q(u6_remainder[42]) );
  DFF_X2 u6_rem_reg_42_ ( .D(u6_remainder[42]), .CK(clk), .Q(remainder[42]) );
  DFF_X2 u6_remainder_reg_43_ ( .D(u6_N43), .CK(clk), .Q(u6_remainder[43]) );
  DFF_X2 u6_rem_reg_43_ ( .D(u6_remainder[43]), .CK(clk), .Q(remainder[43]) );
  DFF_X2 u6_remainder_reg_44_ ( .D(n4765), .CK(clk), .Q(u6_remainder[44]) );
  DFF_X2 u6_rem_reg_44_ ( .D(u6_remainder[44]), .CK(clk), .Q(remainder[44]) );
  DFF_X2 u6_remainder_reg_45_ ( .D(u6_N45), .CK(clk), .Q(u6_remainder[45]) );
  DFF_X2 u6_rem_reg_45_ ( .D(u6_remainder[45]), .CK(clk), .Q(remainder[45]) );
  DFF_X2 u6_remainder_reg_46_ ( .D(u6_N46), .CK(clk), .Q(u6_remainder[46]) );
  DFF_X2 u6_rem_reg_46_ ( .D(u6_remainder[46]), .CK(clk), .Q(remainder[46]) );
  DFF_X2 u6_remainder_reg_47_ ( .D(n4424), .CK(clk), .Q(u6_remainder[47]) );
  DFF_X2 u6_rem_reg_47_ ( .D(u6_remainder[47]), .CK(clk), .Q(remainder[47]) );
  DFF_X2 u6_remainder_reg_48_ ( .D(u6_N48), .CK(clk), .Q(u6_remainder[48]) );
  DFF_X2 u6_rem_reg_48_ ( .D(u6_remainder[48]), .CK(clk), .Q(remainder[48]) );
  DFF_X2 u6_remainder_reg_49_ ( .D(u6_N49), .CK(clk), .Q(u6_remainder[49]) );
  DFF_X2 u6_rem_reg_49_ ( .D(u6_remainder[49]), .CK(clk), .Q(remainder[49]) );
  DFF_X2 u6_remainder_reg_50_ ( .D(u6_N50), .CK(clk), .Q(u6_remainder[50]) );
  DFF_X2 u6_rem_reg_50_ ( .D(u6_remainder[50]), .CK(clk), .Q(remainder[50]) );
  DFF_X2 u6_remainder_reg_51_ ( .D(u6_N51), .CK(clk), .Q(u6_remainder[51]) );
  DFF_X2 u6_rem_reg_51_ ( .D(u6_remainder[51]), .CK(clk), .Q(remainder[51]) );
  DFF_X2 u6_remainder_reg_52_ ( .D(n4309), .CK(clk), .Q(u6_remainder[52]) );
  DFF_X2 u6_rem_reg_52_ ( .D(u6_remainder[52]), .CK(clk), .Q(remainder[52]) );
  DFF_X2 u6_remainder_reg_55_ ( .D(u6_N55), .CK(clk), .Q(u6_remainder[55]) );
  DFF_X2 u6_rem_reg_55_ ( .D(u6_remainder[55]), .CK(clk), .Q(remainder[55]) );
  DFF_X2 u6_remainder_reg_56_ ( .D(u6_N56), .CK(clk), .Q(u6_remainder[56]) );
  DFF_X2 u6_rem_reg_56_ ( .D(u6_remainder[56]), .CK(clk), .Q(remainder[56]) );
  DFF_X2 u6_remainder_reg_57_ ( .D(u6_N57), .CK(clk), .Q(u6_remainder[57]) );
  DFF_X2 u6_rem_reg_57_ ( .D(u6_remainder[57]), .CK(clk), .Q(remainder[57]) );
  DFF_X2 u6_remainder_reg_58_ ( .D(u6_N58), .CK(clk), .Q(u6_remainder[58]) );
  DFF_X2 u6_rem_reg_58_ ( .D(u6_remainder[58]), .CK(clk), .Q(remainder[58]) );
  DFF_X2 u6_remainder_reg_59_ ( .D(u6_N59), .CK(clk), .Q(u6_remainder[59]) );
  DFF_X2 u6_rem_reg_59_ ( .D(u6_remainder[59]), .CK(clk), .Q(remainder[59]) );
  DFF_X2 u6_remainder_reg_60_ ( .D(u6_N60), .CK(clk), .Q(u6_remainder[60]) );
  DFF_X2 u6_rem_reg_60_ ( .D(u6_remainder[60]), .CK(clk), .QN(n4413) );
  DFF_X2 u6_remainder_reg_61_ ( .D(u6_N61), .CK(clk), .Q(u6_remainder[61]) );
  DFF_X2 u6_rem_reg_61_ ( .D(u6_remainder[61]), .CK(clk), .Q(remainder[61]) );
  DFF_X2 u6_remainder_reg_62_ ( .D(u6_N62), .CK(clk), .Q(u6_remainder[62]) );
  DFF_X2 u6_rem_reg_62_ ( .D(u6_remainder[62]), .CK(clk), .Q(remainder[62]) );
  DFF_X2 u6_remainder_reg_63_ ( .D(u6_N63), .CK(clk), .Q(u6_remainder[63]) );
  DFF_X2 u6_rem_reg_63_ ( .D(u6_remainder[63]), .CK(clk), .Q(remainder[63]) );
  DFF_X2 u6_remainder_reg_64_ ( .D(u6_N64), .CK(clk), .Q(u6_remainder[64]) );
  DFF_X2 u6_rem_reg_64_ ( .D(u6_remainder[64]), .CK(clk), .Q(remainder[64]) );
  DFF_X2 u6_remainder_reg_65_ ( .D(u6_N65), .CK(clk), .Q(u6_remainder[65]) );
  DFF_X2 u6_rem_reg_65_ ( .D(u6_remainder[65]), .CK(clk), .Q(remainder[65]) );
  DFF_X2 u6_remainder_reg_66_ ( .D(u6_N66), .CK(clk), .Q(u6_remainder[66]) );
  DFF_X2 u6_rem_reg_66_ ( .D(u6_remainder[66]), .CK(clk), .Q(remainder[66]) );
  DFF_X2 u6_remainder_reg_67_ ( .D(u6_N67), .CK(clk), .Q(u6_remainder[67]) );
  DFF_X2 u6_rem_reg_67_ ( .D(u6_remainder[67]), .CK(clk), .QN(n4412) );
  DFF_X2 u6_remainder_reg_68_ ( .D(u6_N68), .CK(clk), .Q(u6_remainder[68]) );
  DFF_X2 u6_rem_reg_68_ ( .D(u6_remainder[68]), .CK(clk), .Q(remainder[68]) );
  DFF_X2 u6_remainder_reg_69_ ( .D(u6_N69), .CK(clk), .Q(u6_remainder[69]) );
  DFF_X2 u6_rem_reg_69_ ( .D(u6_remainder[69]), .CK(clk), .Q(remainder[69]) );
  DFF_X2 u6_remainder_reg_70_ ( .D(u6_N70), .CK(clk), .Q(u6_remainder[70]) );
  DFF_X2 u6_rem_reg_70_ ( .D(u6_remainder[70]), .CK(clk), .Q(remainder[70]) );
  DFF_X2 u6_remainder_reg_71_ ( .D(u6_N71), .CK(clk), .Q(u6_remainder[71]) );
  DFF_X2 u6_rem_reg_71_ ( .D(u6_remainder[71]), .CK(clk), .Q(remainder[71]) );
  DFF_X2 u6_remainder_reg_72_ ( .D(u6_N72), .CK(clk), .Q(u6_remainder[72]) );
  DFF_X2 u6_rem_reg_72_ ( .D(u6_remainder[72]), .CK(clk), .Q(remainder[72]) );
  DFF_X2 u6_remainder_reg_73_ ( .D(u6_N73), .CK(clk), .Q(u6_remainder[73]) );
  DFF_X2 u6_rem_reg_73_ ( .D(u6_remainder[73]), .CK(clk), .Q(remainder[73]) );
  DFF_X2 u6_remainder_reg_74_ ( .D(u6_N74), .CK(clk), .Q(u6_remainder[74]) );
  DFF_X2 u6_rem_reg_74_ ( .D(u6_remainder[74]), .CK(clk), .Q(remainder[74]) );
  DFF_X2 u6_remainder_reg_75_ ( .D(u6_N75), .CK(clk), .Q(u6_remainder[75]) );
  DFF_X2 u6_rem_reg_75_ ( .D(u6_remainder[75]), .CK(clk), .Q(remainder[75]) );
  DFF_X2 u6_remainder_reg_76_ ( .D(u6_N76), .CK(clk), .Q(u6_remainder[76]) );
  DFF_X2 u6_rem_reg_76_ ( .D(u6_remainder[76]), .CK(clk), .Q(remainder[76]) );
  DFF_X2 u6_remainder_reg_77_ ( .D(u6_N77), .CK(clk), .Q(u6_remainder[77]) );
  DFF_X2 u6_rem_reg_77_ ( .D(u6_remainder[77]), .CK(clk), .Q(remainder[77]) );
  DFF_X2 u6_remainder_reg_78_ ( .D(u6_N78), .CK(clk), .Q(u6_remainder[78]) );
  DFF_X2 u6_rem_reg_78_ ( .D(u6_remainder[78]), .CK(clk), .Q(remainder[78]) );
  DFF_X2 u6_remainder_reg_79_ ( .D(u6_N79), .CK(clk), .Q(u6_remainder[79]) );
  DFF_X2 u6_rem_reg_79_ ( .D(u6_remainder[79]), .CK(clk), .Q(remainder[79]) );
  DFF_X2 u6_remainder_reg_80_ ( .D(u6_N80), .CK(clk), .Q(u6_remainder[80]) );
  DFF_X2 u6_rem_reg_80_ ( .D(u6_remainder[80]), .CK(clk), .Q(remainder[80]) );
  DFF_X2 u6_remainder_reg_81_ ( .D(u6_N81), .CK(clk), .Q(u6_remainder[81]) );
  DFF_X2 u6_rem_reg_81_ ( .D(u6_remainder[81]), .CK(clk), .Q(remainder[81]) );
  DFF_X2 u6_remainder_reg_82_ ( .D(u6_N82), .CK(clk), .Q(u6_remainder[82]) );
  DFF_X2 u6_rem_reg_82_ ( .D(u6_remainder[82]), .CK(clk), .Q(remainder[82]) );
  DFF_X2 u6_remainder_reg_83_ ( .D(u6_N83), .CK(clk), .Q(u6_remainder[83]) );
  DFF_X2 u6_rem_reg_83_ ( .D(u6_remainder[83]), .CK(clk), .Q(remainder[83]) );
  DFF_X2 u6_remainder_reg_84_ ( .D(u6_N84), .CK(clk), .Q(u6_remainder[84]) );
  DFF_X2 u6_rem_reg_84_ ( .D(u6_remainder[84]), .CK(clk), .Q(remainder[84]) );
  DFF_X2 u6_remainder_reg_85_ ( .D(u6_N85), .CK(clk), .Q(u6_remainder[85]) );
  DFF_X2 u6_rem_reg_85_ ( .D(u6_remainder[85]), .CK(clk), .Q(remainder[85]) );
  DFF_X2 u6_remainder_reg_86_ ( .D(u6_N86), .CK(clk), .Q(u6_remainder[86]) );
  DFF_X2 u6_rem_reg_86_ ( .D(u6_remainder[86]), .CK(clk), .Q(remainder[86]) );
  DFF_X2 u6_remainder_reg_87_ ( .D(u6_N87), .CK(clk), .Q(u6_remainder[87]) );
  DFF_X2 u6_rem_reg_87_ ( .D(u6_remainder[87]), .CK(clk), .QN(n4415) );
  DFF_X2 u6_remainder_reg_88_ ( .D(u6_N88), .CK(clk), .Q(u6_remainder[88]) );
  DFF_X2 u6_rem_reg_88_ ( .D(u6_remainder[88]), .CK(clk), .Q(remainder[88]) );
  DFF_X2 u6_remainder_reg_89_ ( .D(u6_N89), .CK(clk), .Q(u6_remainder[89]) );
  DFF_X2 u6_rem_reg_89_ ( .D(u6_remainder[89]), .CK(clk), .Q(remainder[89]) );
  DFF_X2 u6_remainder_reg_90_ ( .D(u6_N90), .CK(clk), .Q(u6_remainder[90]) );
  DFF_X2 u6_rem_reg_90_ ( .D(u6_remainder[90]), .CK(clk), .Q(remainder[90]) );
  DFF_X2 u6_remainder_reg_91_ ( .D(u6_N91), .CK(clk), .Q(u6_remainder[91]) );
  DFF_X2 u6_rem_reg_91_ ( .D(u6_remainder[91]), .CK(clk), .Q(remainder[91]) );
  DFF_X2 u6_remainder_reg_92_ ( .D(u6_N92), .CK(clk), .Q(u6_remainder[92]) );
  DFF_X2 u6_rem_reg_92_ ( .D(u6_remainder[92]), .CK(clk), .Q(remainder[92]) );
  DFF_X2 u6_remainder_reg_93_ ( .D(u6_N93), .CK(clk), .Q(u6_remainder[93]) );
  DFF_X2 u6_rem_reg_93_ ( .D(u6_remainder[93]), .CK(clk), .Q(remainder[93]) );
  DFF_X2 u6_remainder_reg_94_ ( .D(u6_N94), .CK(clk), .Q(u6_remainder[94]) );
  DFF_X2 u6_rem_reg_94_ ( .D(u6_remainder[94]), .CK(clk), .QN(n4414) );
  DFF_X2 u6_remainder_reg_95_ ( .D(u6_N95), .CK(clk), .Q(u6_remainder[95]) );
  DFF_X2 u6_rem_reg_95_ ( .D(u6_remainder[95]), .CK(clk), .Q(remainder[95]) );
  DFF_X2 u6_remainder_reg_96_ ( .D(u6_N96), .CK(clk), .Q(u6_remainder[96]) );
  DFF_X2 u6_rem_reg_96_ ( .D(u6_remainder[96]), .CK(clk), .Q(remainder[96]) );
  DFF_X2 u6_remainder_reg_97_ ( .D(u6_N97), .CK(clk), .Q(u6_remainder[97]) );
  DFF_X2 u6_rem_reg_97_ ( .D(u6_remainder[97]), .CK(clk), .Q(remainder[97]) );
  DFF_X2 u6_remainder_reg_98_ ( .D(u6_N98), .CK(clk), .Q(u6_remainder[98]) );
  DFF_X2 u6_rem_reg_98_ ( .D(u6_remainder[98]), .CK(clk), .Q(remainder[98]) );
  DFF_X2 u6_remainder_reg_99_ ( .D(u6_N99), .CK(clk), .Q(u6_remainder[99]) );
  DFF_X2 u6_rem_reg_99_ ( .D(u6_remainder[99]), .CK(clk), .Q(remainder[99]) );
  DFF_X2 u6_remainder_reg_100_ ( .D(u6_N100), .CK(clk), .Q(u6_remainder[100])
         );
  DFF_X2 u6_rem_reg_100_ ( .D(u6_remainder[100]), .CK(clk), .Q(remainder[100])
         );
  DFF_X2 u6_remainder_reg_101_ ( .D(u6_N101), .CK(clk), .Q(u6_remainder[101])
         );
  DFF_X2 u6_rem_reg_101_ ( .D(u6_remainder[101]), .CK(clk), .Q(remainder[101])
         );
  DFF_X2 u6_remainder_reg_102_ ( .D(u6_N102), .CK(clk), .Q(u6_remainder[102])
         );
  DFF_X2 u6_rem_reg_102_ ( .D(u6_remainder[102]), .CK(clk), .Q(remainder[102])
         );
  DFF_X2 u6_remainder_reg_103_ ( .D(u6_N103), .CK(clk), .Q(u6_remainder[103])
         );
  DFF_X2 u6_rem_reg_103_ ( .D(u6_remainder[103]), .CK(clk), .Q(remainder[103])
         );
  DFF_X2 u6_remainder_reg_104_ ( .D(u6_N104), .CK(clk), .Q(u6_remainder[104])
         );
  DFF_X2 u6_rem_reg_104_ ( .D(u6_remainder[104]), .CK(clk), .Q(remainder[104])
         );
  DFF_X2 u6_remainder_reg_105_ ( .D(u6_N105), .CK(clk), .Q(u6_remainder[105])
         );
  DFF_X2 u6_rem_reg_105_ ( .D(u6_remainder[105]), .CK(clk), .Q(remainder[105])
         );
  DFF_X2 u6_remainder_reg_106_ ( .D(u6_N106), .CK(clk), .Q(u6_remainder[106])
         );
  DFF_X2 u6_rem_reg_106_ ( .D(u6_remainder[106]), .CK(clk), .Q(remainder[106])
         );
  DFF_X2 u6_remainder_reg_107_ ( .D(u6_N107), .CK(clk), .Q(u6_remainder[107])
         );
  DFF_X2 u6_rem_reg_107_ ( .D(u6_remainder[107]), .CK(clk), .Q(remainder[107])
         );
  DFF_X2 u6_quo1_reg_0_ ( .D(u6_N0), .CK(clk), .Q(u6_quo1[0]) );
  DFF_X2 u6_quo_reg_0_ ( .D(u6_quo1[0]), .CK(clk), .Q(quo[0]) );
  DFF_X2 u6_quo1_reg_1_ ( .D(u6_N1), .CK(clk), .Q(u6_quo1[1]) );
  DFF_X2 u6_quo_reg_1_ ( .D(u6_quo1[1]), .CK(clk), .Q(quo[1]) );
  DFF_X2 u6_quo1_reg_2_ ( .D(u6_N2), .CK(clk), .Q(u6_quo1[2]) );
  DFF_X2 u6_quo_reg_2_ ( .D(u6_quo1[2]), .CK(clk), .Q(quo[2]) );
  DFF_X2 u6_quo1_reg_3_ ( .D(u6_N3), .CK(clk), .Q(u6_quo1[3]) );
  DFF_X2 u6_quo_reg_3_ ( .D(u6_quo1[3]), .CK(clk), .Q(quo[3]) );
  DFF_X2 u6_quo1_reg_4_ ( .D(u6_N4), .CK(clk), .Q(u6_quo1[4]) );
  DFF_X2 u6_quo_reg_4_ ( .D(u6_quo1[4]), .CK(clk), .Q(quo[4]) );
  DFF_X2 u6_quo1_reg_5_ ( .D(u6_N5), .CK(clk), .Q(u6_quo1[5]) );
  DFF_X2 u6_quo_reg_5_ ( .D(u6_quo1[5]), .CK(clk), .Q(quo[5]) );
  DFF_X2 u6_quo1_reg_6_ ( .D(u6_N6), .CK(clk), .Q(u6_quo1[6]) );
  DFF_X2 u6_quo_reg_6_ ( .D(u6_quo1[6]), .CK(clk), .Q(quo[6]) );
  DFF_X2 u6_quo1_reg_7_ ( .D(u6_N7), .CK(clk), .Q(u6_quo1[7]) );
  DFF_X2 u6_quo_reg_7_ ( .D(u6_quo1[7]), .CK(clk), .Q(quo[7]) );
  DFF_X2 u6_quo1_reg_8_ ( .D(u6_N8), .CK(clk), .Q(u6_quo1[8]) );
  DFF_X2 u6_quo_reg_8_ ( .D(u6_quo1[8]), .CK(clk), .Q(quo[8]) );
  DFF_X2 u6_quo1_reg_9_ ( .D(u6_N9), .CK(clk), .Q(u6_quo1[9]) );
  DFF_X2 u6_quo_reg_9_ ( .D(u6_quo1[9]), .CK(clk), .Q(quo[9]) );
  DFF_X2 u6_quo1_reg_10_ ( .D(u6_N10), .CK(clk), .Q(u6_quo1[10]) );
  DFF_X2 u6_quo_reg_10_ ( .D(u6_quo1[10]), .CK(clk), .Q(quo[10]) );
  DFF_X2 u6_quo1_reg_11_ ( .D(u6_N11), .CK(clk), .Q(u6_quo1[11]) );
  DFF_X2 u6_quo_reg_11_ ( .D(u6_quo1[11]), .CK(clk), .Q(quo[11]) );
  DFF_X2 u6_quo1_reg_12_ ( .D(u6_N12), .CK(clk), .Q(u6_quo1[12]) );
  DFF_X2 u6_quo_reg_12_ ( .D(u6_quo1[12]), .CK(clk), .Q(quo[12]) );
  DFF_X2 u6_quo1_reg_13_ ( .D(u6_N13), .CK(clk), .Q(u6_quo1[13]) );
  DFF_X2 u6_quo_reg_13_ ( .D(u6_quo1[13]), .CK(clk), .Q(quo[13]) );
  DFF_X2 u6_quo1_reg_14_ ( .D(u6_N14), .CK(clk), .Q(u6_quo1[14]) );
  DFF_X2 u6_quo_reg_14_ ( .D(u6_quo1[14]), .CK(clk), .Q(quo[14]) );
  DFF_X2 u6_quo1_reg_15_ ( .D(u6_N15), .CK(clk), .Q(u6_quo1[15]) );
  DFF_X2 u6_quo_reg_15_ ( .D(u6_quo1[15]), .CK(clk), .Q(quo[15]) );
  DFF_X2 u6_quo1_reg_16_ ( .D(u6_N16), .CK(clk), .Q(u6_quo1[16]) );
  DFF_X2 u6_quo_reg_16_ ( .D(u6_quo1[16]), .CK(clk), .Q(quo[16]) );
  DFF_X2 u6_quo1_reg_17_ ( .D(u6_N17), .CK(clk), .Q(u6_quo1[17]) );
  DFF_X2 u6_quo_reg_17_ ( .D(u6_quo1[17]), .CK(clk), .Q(quo[17]) );
  DFF_X2 u6_quo1_reg_18_ ( .D(u6_N18), .CK(clk), .Q(u6_quo1[18]) );
  DFF_X2 u6_quo_reg_18_ ( .D(u6_quo1[18]), .CK(clk), .Q(quo[18]) );
  DFF_X2 u6_quo1_reg_19_ ( .D(u6_N19), .CK(clk), .Q(u6_quo1[19]) );
  DFF_X2 u6_quo_reg_19_ ( .D(u6_quo1[19]), .CK(clk), .Q(quo[19]) );
  DFF_X2 u6_quo1_reg_20_ ( .D(u6_N20), .CK(clk), .Q(u6_quo1[20]) );
  DFF_X2 u6_quo_reg_20_ ( .D(u6_quo1[20]), .CK(clk), .Q(quo[20]) );
  DFF_X2 u6_quo1_reg_21_ ( .D(u6_N21), .CK(clk), .Q(u6_quo1[21]) );
  DFF_X2 u6_quo_reg_21_ ( .D(u6_quo1[21]), .CK(clk), .Q(quo[21]) );
  DFF_X2 u6_quo1_reg_22_ ( .D(u6_N22), .CK(clk), .Q(u6_quo1[22]) );
  DFF_X2 u6_quo_reg_22_ ( .D(u6_quo1[22]), .CK(clk), .Q(quo[22]) );
  DFF_X2 u6_quo1_reg_23_ ( .D(u6_N23), .CK(clk), .Q(u6_quo1[23]) );
  DFF_X2 u6_quo_reg_23_ ( .D(u6_quo1[23]), .CK(clk), .Q(quo[23]) );
  DFF_X2 u6_quo1_reg_24_ ( .D(u6_N24), .CK(clk), .Q(u6_quo1[24]) );
  DFF_X2 u6_quo_reg_24_ ( .D(u6_quo1[24]), .CK(clk), .Q(quo[24]) );
  DFF_X2 u6_quo1_reg_25_ ( .D(u6_N25), .CK(clk), .Q(u6_quo1[25]) );
  DFF_X2 u6_quo_reg_25_ ( .D(u6_quo1[25]), .CK(clk), .Q(quo[25]) );
  DFF_X2 u6_quo1_reg_26_ ( .D(u6_N26), .CK(clk), .Q(u6_quo1[26]) );
  DFF_X2 u6_quo_reg_26_ ( .D(u6_quo1[26]), .CK(clk), .Q(quo[26]) );
  DFF_X2 u6_quo1_reg_27_ ( .D(u6_N27), .CK(clk), .Q(u6_quo1[27]) );
  DFF_X2 u6_quo_reg_27_ ( .D(u6_quo1[27]), .CK(clk), .Q(quo[27]) );
  DFF_X2 u6_quo1_reg_28_ ( .D(n4764), .CK(clk), .Q(u6_quo1[28]) );
  DFF_X2 u6_quo_reg_28_ ( .D(u6_quo1[28]), .CK(clk), .Q(quo[28]) );
  DFF_X2 u6_quo1_reg_29_ ( .D(u6_N29), .CK(clk), .Q(u6_quo1[29]) );
  DFF_X2 u6_quo_reg_29_ ( .D(u6_quo1[29]), .CK(clk), .Q(quo[29]) );
  DFF_X2 u6_quo1_reg_30_ ( .D(u6_N30), .CK(clk), .Q(u6_quo1[30]) );
  DFF_X2 u6_quo_reg_30_ ( .D(u6_quo1[30]), .CK(clk), .Q(quo[30]) );
  DFF_X2 u6_quo1_reg_31_ ( .D(u6_N31), .CK(clk), .Q(u6_quo1[31]) );
  DFF_X2 u6_quo_reg_31_ ( .D(u6_quo1[31]), .CK(clk), .Q(quo[31]) );
  DFF_X2 u6_quo1_reg_32_ ( .D(u6_N32), .CK(clk), .Q(u6_quo1[32]) );
  DFF_X2 u6_quo_reg_32_ ( .D(u6_quo1[32]), .CK(clk), .Q(quo[32]) );
  DFF_X2 u6_quo1_reg_33_ ( .D(u6_N33), .CK(clk), .Q(u6_quo1[33]) );
  DFF_X2 u6_quo_reg_33_ ( .D(u6_quo1[33]), .CK(clk), .Q(quo[33]) );
  DFF_X2 u6_quo1_reg_34_ ( .D(n4786), .CK(clk), .Q(u6_quo1[34]) );
  DFF_X2 u6_quo_reg_34_ ( .D(u6_quo1[34]), .CK(clk), .Q(quo[34]) );
  DFF_X2 u6_quo1_reg_35_ ( .D(u6_N35), .CK(clk), .Q(u6_quo1[35]) );
  DFF_X2 u6_quo_reg_35_ ( .D(u6_quo1[35]), .CK(clk), .Q(quo[35]) );
  DFF_X2 u6_quo1_reg_36_ ( .D(u6_N36), .CK(clk), .Q(u6_quo1[36]) );
  DFF_X2 u6_quo_reg_36_ ( .D(u6_quo1[36]), .CK(clk), .Q(quo[36]) );
  DFF_X2 u6_quo1_reg_37_ ( .D(u6_N37), .CK(clk), .Q(u6_quo1[37]) );
  DFF_X2 u6_quo_reg_37_ ( .D(u6_quo1[37]), .CK(clk), .Q(quo[37]) );
  DFF_X2 u6_quo1_reg_38_ ( .D(n4791), .CK(clk), .Q(u6_quo1[38]) );
  DFF_X2 u6_quo_reg_38_ ( .D(u6_quo1[38]), .CK(clk), .Q(quo[38]) );
  DFF_X2 u6_quo1_reg_39_ ( .D(u6_N39), .CK(clk), .Q(u6_quo1[39]) );
  DFF_X2 u6_quo_reg_39_ ( .D(u6_quo1[39]), .CK(clk), .Q(quo[39]) );
  DFF_X2 u6_quo1_reg_40_ ( .D(u6_N40), .CK(clk), .Q(u6_quo1[40]) );
  DFF_X2 u6_quo_reg_40_ ( .D(u6_quo1[40]), .CK(clk), .Q(quo[40]) );
  DFF_X2 u6_quo1_reg_41_ ( .D(n4772), .CK(clk), .Q(u6_quo1[41]) );
  DFF_X2 u6_quo_reg_41_ ( .D(u6_quo1[41]), .CK(clk), .Q(quo[41]) );
  DFF_X2 u6_quo1_reg_42_ ( .D(n4787), .CK(clk), .Q(u6_quo1[42]) );
  DFF_X2 u6_quo_reg_42_ ( .D(u6_quo1[42]), .CK(clk), .Q(quo[42]) );
  DFF_X2 u6_quo1_reg_43_ ( .D(u6_N43), .CK(clk), .Q(u6_quo1[43]) );
  DFF_X2 u6_quo_reg_43_ ( .D(u6_quo1[43]), .CK(clk), .Q(quo[43]) );
  DFF_X2 u6_quo1_reg_44_ ( .D(n4765), .CK(clk), .Q(u6_quo1[44]) );
  DFF_X2 u6_quo_reg_44_ ( .D(u6_quo1[44]), .CK(clk), .Q(quo[44]) );
  DFF_X2 u6_quo1_reg_45_ ( .D(u6_N45), .CK(clk), .Q(u6_quo1[45]) );
  DFF_X2 u6_quo_reg_45_ ( .D(u6_quo1[45]), .CK(clk), .Q(quo[45]) );
  DFF_X2 u6_quo1_reg_46_ ( .D(u6_N46), .CK(clk), .Q(u6_quo1[46]) );
  DFF_X2 u6_quo_reg_46_ ( .D(u6_quo1[46]), .CK(clk), .Q(quo[46]) );
  DFF_X2 u6_quo1_reg_47_ ( .D(n4424), .CK(clk), .Q(u6_quo1[47]) );
  DFF_X2 u6_quo_reg_47_ ( .D(u6_quo1[47]), .CK(clk), .Q(quo[47]) );
  DFF_X2 u6_quo1_reg_48_ ( .D(u6_N48), .CK(clk), .Q(u6_quo1[48]) );
  DFF_X2 u6_quo_reg_48_ ( .D(u6_quo1[48]), .CK(clk), .Q(quo[48]) );
  DFF_X2 u6_quo1_reg_49_ ( .D(u6_N49), .CK(clk), .Q(u6_quo1[49]) );
  DFF_X2 u6_quo_reg_49_ ( .D(u6_quo1[49]), .CK(clk), .Q(quo[49]) );
  DFF_X2 u6_quo1_reg_50_ ( .D(u6_N50), .CK(clk), .Q(u6_quo1[50]) );
  DFF_X2 u6_quo_reg_50_ ( .D(u6_quo1[50]), .CK(clk), .Q(quo[50]) );
  DFF_X2 u6_quo1_reg_51_ ( .D(u6_N51), .CK(clk), .Q(u6_quo1[51]) );
  DFF_X2 u6_quo_reg_51_ ( .D(u6_quo1[51]), .CK(clk), .Q(quo[51]) );
  DFF_X2 u6_quo1_reg_52_ ( .D(n4309), .CK(clk), .Q(u6_quo1[52]) );
  DFF_X2 u6_quo_reg_52_ ( .D(u6_quo1[52]), .CK(clk), .Q(quo[52]) );
  DFF_X2 u6_quo1_reg_55_ ( .D(u6_N55), .CK(clk), .Q(u6_quo1[55]) );
  DFF_X2 u6_quo_reg_55_ ( .D(u6_quo1[55]), .CK(clk), .Q(quo[55]) );
  DFF_X2 u6_quo1_reg_56_ ( .D(u6_N56), .CK(clk), .Q(u6_quo1[56]) );
  DFF_X2 u6_quo_reg_56_ ( .D(u6_quo1[56]), .CK(clk), .Q(quo[56]) );
  DFF_X2 u6_quo1_reg_57_ ( .D(u6_N57), .CK(clk), .Q(u6_quo1[57]) );
  DFF_X2 u6_quo_reg_57_ ( .D(u6_quo1[57]), .CK(clk), .Q(quo[57]) );
  DFF_X2 u6_quo1_reg_58_ ( .D(u6_N58), .CK(clk), .Q(u6_quo1[58]) );
  DFF_X2 u6_quo_reg_58_ ( .D(u6_quo1[58]), .CK(clk), .Q(quo[58]) );
  DFF_X2 u6_quo1_reg_59_ ( .D(u6_N59), .CK(clk), .Q(u6_quo1[59]) );
  DFF_X2 u6_quo_reg_59_ ( .D(u6_quo1[59]), .CK(clk), .Q(quo[59]) );
  DFF_X2 u6_quo1_reg_60_ ( .D(u6_N60), .CK(clk), .Q(u6_quo1[60]) );
  DFF_X2 u6_quo_reg_60_ ( .D(u6_quo1[60]), .CK(clk), .Q(quo[60]) );
  DFF_X2 u6_quo1_reg_61_ ( .D(u6_N61), .CK(clk), .Q(u6_quo1[61]) );
  DFF_X2 u6_quo_reg_61_ ( .D(u6_quo1[61]), .CK(clk), .Q(quo[61]) );
  DFF_X2 u6_quo1_reg_62_ ( .D(u6_N62), .CK(clk), .Q(u6_quo1[62]) );
  DFF_X2 u6_quo_reg_62_ ( .D(u6_quo1[62]), .CK(clk), .Q(quo[62]) );
  DFF_X2 u6_quo1_reg_63_ ( .D(u6_N63), .CK(clk), .Q(u6_quo1[63]) );
  DFF_X2 u6_quo_reg_63_ ( .D(u6_quo1[63]), .CK(clk), .Q(quo[63]) );
  DFF_X2 u6_quo1_reg_64_ ( .D(u6_N64), .CK(clk), .Q(u6_quo1[64]) );
  DFF_X2 u6_quo_reg_64_ ( .D(u6_quo1[64]), .CK(clk), .Q(quo[64]) );
  DFF_X2 u6_quo1_reg_65_ ( .D(u6_N65), .CK(clk), .Q(u6_quo1[65]) );
  DFF_X2 u6_quo_reg_65_ ( .D(u6_quo1[65]), .CK(clk), .Q(quo[65]) );
  DFF_X2 u6_quo1_reg_66_ ( .D(u6_N66), .CK(clk), .Q(u6_quo1[66]) );
  DFF_X2 u6_quo_reg_66_ ( .D(u6_quo1[66]), .CK(clk), .Q(quo[66]) );
  DFF_X2 u6_quo1_reg_67_ ( .D(u6_N67), .CK(clk), .Q(u6_quo1[67]) );
  DFF_X2 u6_quo_reg_67_ ( .D(u6_quo1[67]), .CK(clk), .Q(quo[67]) );
  DFF_X2 u6_quo1_reg_68_ ( .D(u6_N68), .CK(clk), .Q(u6_quo1[68]) );
  DFF_X2 u6_quo_reg_68_ ( .D(u6_quo1[68]), .CK(clk), .Q(quo[68]) );
  DFF_X2 u6_quo1_reg_69_ ( .D(u6_N69), .CK(clk), .Q(u6_quo1[69]) );
  DFF_X2 u6_quo_reg_69_ ( .D(u6_quo1[69]), .CK(clk), .Q(quo[69]) );
  DFF_X2 u6_quo1_reg_70_ ( .D(u6_N70), .CK(clk), .Q(u6_quo1[70]) );
  DFF_X2 u6_quo_reg_70_ ( .D(u6_quo1[70]), .CK(clk), .Q(quo[70]) );
  DFF_X2 u6_quo1_reg_71_ ( .D(u6_N71), .CK(clk), .Q(u6_quo1[71]) );
  DFF_X2 u6_quo_reg_71_ ( .D(u6_quo1[71]), .CK(clk), .Q(quo[71]) );
  DFF_X2 u6_quo1_reg_72_ ( .D(u6_N72), .CK(clk), .Q(u6_quo1[72]) );
  DFF_X2 u6_quo_reg_72_ ( .D(u6_quo1[72]), .CK(clk), .Q(quo[72]) );
  DFF_X2 u6_quo1_reg_73_ ( .D(u6_N73), .CK(clk), .Q(u6_quo1[73]) );
  DFF_X2 u6_quo_reg_73_ ( .D(u6_quo1[73]), .CK(clk), .Q(quo[73]) );
  DFF_X2 u6_quo1_reg_74_ ( .D(u6_N74), .CK(clk), .Q(u6_quo1[74]) );
  DFF_X2 u6_quo_reg_74_ ( .D(u6_quo1[74]), .CK(clk), .Q(quo[74]) );
  DFF_X2 u6_quo1_reg_75_ ( .D(u6_N75), .CK(clk), .Q(u6_quo1[75]) );
  DFF_X2 u6_quo_reg_75_ ( .D(u6_quo1[75]), .CK(clk), .Q(quo[75]) );
  DFF_X2 u6_quo1_reg_76_ ( .D(u6_N76), .CK(clk), .Q(u6_quo1[76]) );
  DFF_X2 u6_quo_reg_76_ ( .D(u6_quo1[76]), .CK(clk), .Q(quo[76]) );
  DFF_X2 u6_quo1_reg_77_ ( .D(u6_N77), .CK(clk), .Q(u6_quo1[77]) );
  DFF_X2 u6_quo_reg_77_ ( .D(u6_quo1[77]), .CK(clk), .Q(quo[77]) );
  DFF_X2 u6_quo1_reg_78_ ( .D(u6_N78), .CK(clk), .Q(u6_quo1[78]) );
  DFF_X2 u6_quo_reg_78_ ( .D(u6_quo1[78]), .CK(clk), .Q(quo[78]) );
  DFF_X2 u6_quo1_reg_79_ ( .D(u6_N79), .CK(clk), .Q(u6_quo1[79]) );
  DFF_X2 u6_quo_reg_79_ ( .D(u6_quo1[79]), .CK(clk), .Q(quo[79]) );
  DFF_X2 u6_quo1_reg_80_ ( .D(u6_N80), .CK(clk), .Q(u6_quo1[80]) );
  DFF_X2 u6_quo_reg_80_ ( .D(u6_quo1[80]), .CK(clk), .Q(quo[80]) );
  DFF_X2 u6_quo1_reg_81_ ( .D(u6_N81), .CK(clk), .Q(u6_quo1[81]) );
  DFF_X2 u6_quo_reg_81_ ( .D(u6_quo1[81]), .CK(clk), .Q(quo[81]) );
  DFF_X2 u6_quo1_reg_82_ ( .D(u6_N82), .CK(clk), .Q(u6_quo1[82]) );
  DFF_X2 u6_quo_reg_82_ ( .D(u6_quo1[82]), .CK(clk), .Q(quo[82]) );
  DFF_X2 u6_quo1_reg_83_ ( .D(u6_N83), .CK(clk), .Q(u6_quo1[83]) );
  DFF_X2 u6_quo_reg_83_ ( .D(u6_quo1[83]), .CK(clk), .Q(quo[83]) );
  DFF_X2 u6_quo1_reg_84_ ( .D(u6_N84), .CK(clk), .Q(u6_quo1[84]) );
  DFF_X2 u6_quo_reg_84_ ( .D(u6_quo1[84]), .CK(clk), .Q(quo[84]) );
  DFF_X2 u6_quo1_reg_85_ ( .D(u6_N85), .CK(clk), .Q(u6_quo1[85]) );
  DFF_X2 u6_quo_reg_85_ ( .D(u6_quo1[85]), .CK(clk), .Q(quo[85]) );
  DFF_X2 u6_quo1_reg_86_ ( .D(u6_N86), .CK(clk), .Q(u6_quo1[86]) );
  DFF_X2 u6_quo_reg_86_ ( .D(u6_quo1[86]), .CK(clk), .Q(quo[86]) );
  DFF_X2 u6_quo1_reg_87_ ( .D(u6_N87), .CK(clk), .Q(u6_quo1[87]) );
  DFF_X2 u6_quo_reg_87_ ( .D(u6_quo1[87]), .CK(clk), .Q(quo[87]) );
  DFF_X2 u6_quo1_reg_88_ ( .D(u6_N88), .CK(clk), .Q(u6_quo1[88]) );
  DFF_X2 u6_quo_reg_88_ ( .D(u6_quo1[88]), .CK(clk), .Q(quo[88]) );
  DFF_X2 u6_quo1_reg_89_ ( .D(u6_N89), .CK(clk), .Q(u6_quo1[89]) );
  DFF_X2 u6_quo_reg_89_ ( .D(u6_quo1[89]), .CK(clk), .Q(quo[89]) );
  DFF_X2 u6_quo1_reg_90_ ( .D(u6_N90), .CK(clk), .Q(u6_quo1[90]) );
  DFF_X2 u6_quo_reg_90_ ( .D(u6_quo1[90]), .CK(clk), .Q(quo[90]) );
  DFF_X2 u6_quo1_reg_91_ ( .D(u6_N91), .CK(clk), .Q(u6_quo1[91]) );
  DFF_X2 u6_quo_reg_91_ ( .D(u6_quo1[91]), .CK(clk), .Q(quo[91]) );
  DFF_X2 u6_quo1_reg_92_ ( .D(u6_N92), .CK(clk), .Q(u6_quo1[92]) );
  DFF_X2 u6_quo_reg_92_ ( .D(u6_quo1[92]), .CK(clk), .Q(quo[92]) );
  DFF_X2 u6_quo1_reg_93_ ( .D(u6_N93), .CK(clk), .Q(u6_quo1[93]) );
  DFF_X2 u6_quo_reg_93_ ( .D(u6_quo1[93]), .CK(clk), .Q(quo[93]) );
  DFF_X2 u6_quo1_reg_94_ ( .D(u6_N94), .CK(clk), .Q(u6_quo1[94]) );
  DFF_X2 u6_quo_reg_94_ ( .D(u6_quo1[94]), .CK(clk), .Q(quo[94]) );
  DFF_X2 u6_quo1_reg_95_ ( .D(u6_N95), .CK(clk), .Q(u6_quo1[95]) );
  DFF_X2 u6_quo_reg_95_ ( .D(u6_quo1[95]), .CK(clk), .Q(quo[95]) );
  DFF_X2 u6_quo1_reg_96_ ( .D(u6_N96), .CK(clk), .Q(u6_quo1[96]) );
  DFF_X2 u6_quo_reg_96_ ( .D(u6_quo1[96]), .CK(clk), .Q(quo[96]) );
  DFF_X2 u6_quo1_reg_97_ ( .D(u6_N97), .CK(clk), .Q(u6_quo1[97]) );
  DFF_X2 u6_quo_reg_97_ ( .D(u6_quo1[97]), .CK(clk), .Q(quo[97]) );
  DFF_X2 u6_quo1_reg_98_ ( .D(u6_N98), .CK(clk), .Q(u6_quo1[98]) );
  DFF_X2 u6_quo_reg_98_ ( .D(u6_quo1[98]), .CK(clk), .Q(quo[98]) );
  DFF_X2 u6_quo1_reg_99_ ( .D(u6_N99), .CK(clk), .Q(u6_quo1[99]) );
  DFF_X2 u6_quo_reg_99_ ( .D(u6_quo1[99]), .CK(clk), .Q(quo[99]) );
  DFF_X2 u6_quo1_reg_100_ ( .D(u6_N100), .CK(clk), .Q(u6_quo1[100]) );
  DFF_X2 u6_quo_reg_100_ ( .D(u6_quo1[100]), .CK(clk), .Q(quo[100]) );
  DFF_X2 u6_quo1_reg_101_ ( .D(u6_N101), .CK(clk), .Q(u6_quo1[101]) );
  DFF_X2 u6_quo_reg_101_ ( .D(u6_quo1[101]), .CK(clk), .Q(quo[101]) );
  DFF_X2 u6_quo1_reg_102_ ( .D(u6_N102), .CK(clk), .Q(u6_quo1[102]) );
  DFF_X2 u6_quo_reg_102_ ( .D(u6_quo1[102]), .CK(clk), .Q(quo[102]) );
  DFF_X2 u6_quo1_reg_103_ ( .D(u6_N103), .CK(clk), .Q(u6_quo1[103]) );
  DFF_X2 u6_quo_reg_103_ ( .D(u6_quo1[103]), .CK(clk), .Q(quo[103]) );
  DFF_X2 u6_quo1_reg_104_ ( .D(u6_N104), .CK(clk), .Q(u6_quo1[104]) );
  DFF_X2 u6_quo_reg_104_ ( .D(u6_quo1[104]), .CK(clk), .Q(quo[104]) );
  DFF_X2 u6_quo1_reg_105_ ( .D(u6_N105), .CK(clk), .Q(u6_quo1[105]) );
  DFF_X2 u6_quo_reg_105_ ( .D(u6_quo1[105]), .CK(clk), .Q(quo[105]) );
  DFF_X2 u6_quo1_reg_106_ ( .D(u6_N106), .CK(clk), .Q(u6_quo1[106]) );
  DFF_X2 u6_quo_reg_106_ ( .D(u6_quo1[106]), .CK(clk), .Q(quo[106]) );
  DFF_X2 out_reg_55_ ( .D(N848), .CK(clk), .Q(out[55]) );
  DFF_X2 out_reg_56_ ( .D(N849), .CK(clk), .Q(out[56]) );
  DFF_X2 out_reg_54_ ( .D(N847), .CK(clk), .Q(out[54]) );
  DFF_X2 out_reg_57_ ( .D(N850), .CK(clk), .Q(out[57]) );
  DFF_X2 out_reg_59_ ( .D(N852), .CK(clk), .Q(out[59]) );
  DFF_X2 out_reg_58_ ( .D(N851), .CK(clk), .Q(out[58]) );
  DFF_X2 out_reg_53_ ( .D(N846), .CK(clk), .Q(out[53]) );
  DFF_X2 out_reg_52_ ( .D(N845), .CK(clk), .Q(out[52]) );
  DFF_X2 out_reg_62_ ( .D(N855), .CK(clk), .Q(out[62]) );
  DFF_X2 out_reg_61_ ( .D(N854), .CK(clk), .Q(out[61]) );
  DFF_X2 out_reg_60_ ( .D(N853), .CK(clk), .Q(out[60]) );
  DFF_X2 overflow_reg ( .D(N899), .CK(clk), .Q(overflow) );
  DFF_X2 out_reg_51_ ( .D(N844), .CK(clk), .Q(out[51]) );
  DFF_X2 out_reg_50_ ( .D(N843), .CK(clk), .Q(out[50]) );
  DFF_X2 out_reg_49_ ( .D(N842), .CK(clk), .Q(out[49]) );
  DFF_X2 out_reg_48_ ( .D(N841), .CK(clk), .Q(out[48]) );
  DFF_X2 out_reg_47_ ( .D(N840), .CK(clk), .Q(out[47]) );
  DFF_X2 out_reg_46_ ( .D(N839), .CK(clk), .Q(out[46]) );
  DFF_X2 out_reg_45_ ( .D(N838), .CK(clk), .Q(out[45]) );
  DFF_X2 out_reg_44_ ( .D(N837), .CK(clk), .Q(out[44]) );
  DFF_X2 out_reg_43_ ( .D(N836), .CK(clk), .Q(out[43]) );
  DFF_X2 out_reg_42_ ( .D(N835), .CK(clk), .Q(out[42]) );
  DFF_X2 out_reg_41_ ( .D(N834), .CK(clk), .Q(out[41]) );
  DFF_X2 out_reg_40_ ( .D(N833), .CK(clk), .Q(out[40]) );
  DFF_X2 out_reg_39_ ( .D(N832), .CK(clk), .Q(out[39]) );
  DFF_X2 out_reg_38_ ( .D(N831), .CK(clk), .Q(out[38]) );
  DFF_X2 out_reg_37_ ( .D(N830), .CK(clk), .Q(out[37]) );
  DFF_X2 out_reg_36_ ( .D(N829), .CK(clk), .Q(out[36]) );
  DFF_X2 out_reg_35_ ( .D(N828), .CK(clk), .Q(out[35]) );
  DFF_X2 out_reg_34_ ( .D(N827), .CK(clk), .Q(out[34]) );
  DFF_X2 out_reg_33_ ( .D(N826), .CK(clk), .Q(out[33]) );
  DFF_X2 out_reg_32_ ( .D(N825), .CK(clk), .Q(out[32]) );
  DFF_X2 out_reg_31_ ( .D(N824), .CK(clk), .Q(out[31]) );
  DFF_X2 out_reg_30_ ( .D(N823), .CK(clk), .Q(out[30]) );
  DFF_X2 out_reg_29_ ( .D(N822), .CK(clk), .Q(out[29]) );
  DFF_X2 out_reg_28_ ( .D(N821), .CK(clk), .Q(out[28]) );
  DFF_X2 out_reg_27_ ( .D(N820), .CK(clk), .Q(out[27]) );
  DFF_X2 out_reg_26_ ( .D(N819), .CK(clk), .Q(out[26]) );
  DFF_X2 out_reg_25_ ( .D(N818), .CK(clk), .Q(out[25]) );
  DFF_X2 out_reg_24_ ( .D(N817), .CK(clk), .Q(out[24]) );
  DFF_X2 out_reg_23_ ( .D(N816), .CK(clk), .Q(out[23]) );
  DFF_X2 out_reg_22_ ( .D(N815), .CK(clk), .Q(out[22]) );
  DFF_X2 out_reg_21_ ( .D(N814), .CK(clk), .Q(out[21]) );
  DFF_X2 out_reg_20_ ( .D(N813), .CK(clk), .Q(out[20]) );
  DFF_X2 out_reg_19_ ( .D(N812), .CK(clk), .Q(out[19]) );
  DFF_X2 out_reg_18_ ( .D(N811), .CK(clk), .Q(out[18]) );
  DFF_X2 out_reg_17_ ( .D(N810), .CK(clk), .Q(out[17]) );
  DFF_X2 out_reg_16_ ( .D(N809), .CK(clk), .Q(out[16]) );
  DFF_X2 out_reg_15_ ( .D(N808), .CK(clk), .Q(out[15]) );
  DFF_X2 out_reg_14_ ( .D(N807), .CK(clk), .Q(out[14]) );
  DFF_X2 out_reg_13_ ( .D(N806), .CK(clk), .Q(out[13]) );
  DFF_X2 out_reg_12_ ( .D(N805), .CK(clk), .Q(out[12]) );
  DFF_X2 out_reg_11_ ( .D(N804), .CK(clk), .Q(out[11]) );
  DFF_X2 out_reg_10_ ( .D(N803), .CK(clk), .Q(out[10]) );
  DFF_X2 out_reg_9_ ( .D(N802), .CK(clk), .Q(out[9]) );
  DFF_X2 out_reg_8_ ( .D(N801), .CK(clk), .Q(out[8]) );
  DFF_X2 out_reg_7_ ( .D(N800), .CK(clk), .Q(out[7]) );
  DFF_X2 out_reg_6_ ( .D(N799), .CK(clk), .Q(out[6]) );
  DFF_X2 out_reg_5_ ( .D(N798), .CK(clk), .Q(out[5]) );
  DFF_X2 out_reg_4_ ( .D(N797), .CK(clk), .Q(out[4]) );
  DFF_X2 out_reg_3_ ( .D(N796), .CK(clk), .Q(out[3]) );
  DFF_X2 out_reg_2_ ( .D(N795), .CK(clk), .Q(out[2]) );
  DFF_X2 out_reg_1_ ( .D(N794), .CK(clk), .Q(out[1]) );
  DFF_X2 inf_reg ( .D(N906), .CK(clk), .Q(inf) );
  DFF_X2 underflow_reg ( .D(N902), .CK(clk), .Q(underflow) );
  DFF_X2 ine_reg ( .D(N889), .CK(clk), .Q(ine) );
  DFF_X2 zero_reg ( .D(N911), .CK(clk), .Q(zero) );
  DFF_X2 out_reg_63_ ( .D(N875), .CK(clk), .Q(out[63]) );
  DFF_X2 out_reg_0_ ( .D(N793), .CK(clk), .Q(out[0]) );
  DFF_X2 u6_quo1_reg_107_ ( .D(u6_N107), .CK(clk), .Q(u6_quo1[107]) );
  DFF_X2 u6_quo_reg_107_ ( .D(u6_quo1[107]), .CK(clk), .Q(quo[107]) );
  DFF_X1 u5_prod1_reg_103_ ( .D(u5_N103), .CK(clk), .Q(u5_prod1[103]) );
  DFF_X1 u5_prod1_reg_89_ ( .D(u5_N89), .CK(clk), .Q(u5_prod1[89]) );
  DFF_X2 opb_r_reg_58_ ( .D(opb[58]), .CK(clk), .Q(n4425), .QN(n4833) );
  DFF_X2 opb_r_reg_59_ ( .D(opb[59]), .CK(clk), .Q(n4819), .QN(n4825) );
  DFF_X2 opa_r_reg_1_ ( .D(opa[1]), .CK(clk), .Q(n4781), .QN(n4816) );
  DFF_X2 opb_r_reg_47_ ( .D(opb[47]), .CK(clk), .Q(n4424), .QN(n4800) );
  DFF_X1 u5_prod1_reg_97_ ( .D(u5_N97), .CK(clk), .Q(u5_prod1[97]) );
  DFF_X1 u5_prod1_reg_104_ ( .D(u5_N104), .CK(clk), .Q(u5_prod1[104]) );
  DFF_X1 u5_prod1_reg_95_ ( .D(u5_N95), .CK(clk), .Q(u5_prod1[95]) );
  DFF_X1 u5_prod1_reg_100_ ( .D(u5_N100), .CK(clk), .Q(u5_prod1[100]) );
  DFF_X1 u5_prod1_reg_90_ ( .D(u5_N90), .CK(clk), .Q(u5_prod1[90]) );
  DFF_X1 u5_prod1_reg_93_ ( .D(u5_N93), .CK(clk), .Q(u5_prod1[93]) );
  DFF_X2 opb_r_reg_38_ ( .D(opb[38]), .CK(clk), .QN(n4788) );
  DFF_X2 opb_r_reg_44_ ( .D(opb[44]), .CK(clk), .Q(n4731), .QN(n4778) );
  DFF_X2 opb_r_reg_34_ ( .D(opb[34]), .CK(clk), .QN(n4771) );
  DFF_X2 opb_r_reg_41_ ( .D(opb[41]), .CK(clk), .QN(n4769) );
  DFF_X1 u5_prod1_reg_96_ ( .D(u5_N96), .CK(clk), .Q(u5_prod1[96]) );
  DFF_X1 opb_r_reg_28_ ( .D(opb[28]), .CK(clk), .QN(n4541) );
  DFF_X2 opb_r_reg_42_ ( .D(opb[42]), .CK(clk), .QN(n4773) );
  DFF_X1 u5_prod1_reg_77_ ( .D(u5_N77), .CK(clk), .Q(u5_prod1[77]) );
  AND4_X2 U1135 ( .A1(opb_00), .A2(opa_nan_r), .A3(n4446), .A4(n4345), .ZN(
        N913) );
  NOR4_X2 U1876 ( .A1(u4_N5931), .A2(u4_N5930), .A3(u4_N5929), .A4(u4_N5928), 
        .ZN(n3927) );
  NOR4_X2 U1871 ( .A1(u4_N5918), .A2(u4_N5917), .A3(u4_N5916), .A4(u4_N5915), 
        .ZN(n3923) );
  NOR4_X2 U1886 ( .A1(u4_N5958), .A2(u4_N5957), .A3(u4_N5956), .A4(u4_N5955), 
        .ZN(n3935) );
  NOR4_X2 U1888 ( .A1(u4_N5951), .A2(u4_N5950), .A3(u4_N5949), .A4(u4_N5948), 
        .ZN(n3933) );
  NOR4_X2 U1881 ( .A1(u4_N5944), .A2(u4_N5943), .A3(u4_N5942), .A4(u4_N5941), 
        .ZN(n3931) );
  AOI22_X2 U1813 ( .A1(u4_N5972), .A2(net63321), .B1(u4_N6080), .B2(net63339), 
        .ZN(n3704) );
  OR2_X2 u4_C19047 ( .A1(u4_exp_out_5_), .A2(u4_N6457), .ZN(u4_N6458) );
  OR2_X2 u4_C19046 ( .A1(u4_N6458), .A2(u4_exp_out_4_), .ZN(u4_N6459) );
  DFF_X1 u5_prod1_reg_83_ ( .D(u5_N83), .CK(clk), .Q(u5_prod1[83]) );
  DFF_X1 u5_prod1_reg_87_ ( .D(u5_N87), .CK(clk), .Q(u5_prod1[87]) );
  DFF_X1 u5_prod1_reg_99_ ( .D(u5_N99), .CK(clk), .Q(u5_prod1[99]) );
  DFF_X1 u5_prod1_reg_92_ ( .D(u5_N92), .CK(clk), .Q(u5_prod1[92]) );
  DFF_X1 u5_prod1_reg_86_ ( .D(u5_N86), .CK(clk), .Q(u5_prod1[86]) );
  DFF_X1 u5_prod1_reg_94_ ( .D(u5_N94), .CK(clk), .Q(u5_prod1[94]) );
  DFF_X1 u5_prod1_reg_47_ ( .D(u5_N47), .CK(clk), .Q(u5_prod1[47]) );
  DFF_X1 u5_prod1_reg_46_ ( .D(u5_N46), .CK(clk), .Q(u5_prod1[46]) );
  DFF_X1 u2_exp_out_reg_2_ ( .D(u2_N78), .CK(clk), .Q(exp_mul[2]), .QN(n4504)
         );
  DFF_X1 u2_exp_out_reg_3_ ( .D(u2_N79), .CK(clk), .Q(exp_mul[3]), .QN(n4503)
         );
  DFF_X1 u2_exp_out_reg_4_ ( .D(u2_N80), .CK(clk), .Q(exp_mul[4]), .QN(n4502)
         );
  DFF_X1 u2_exp_out_reg_6_ ( .D(u2_N82), .CK(clk), .Q(exp_mul[6]), .QN(n4501)
         );
  DFF_X1 u2_exp_out_reg_5_ ( .D(u2_N81), .CK(clk), .Q(exp_mul[5]), .QN(n4500)
         );
  DFF_X1 u2_exp_out_reg_7_ ( .D(u2_N83), .CK(clk), .Q(exp_mul[7]), .QN(n4499)
         );
  DFF_X1 u2_exp_out_reg_8_ ( .D(u2_N84), .CK(clk), .QN(n4492) );
  DFF_X1 u2_exp_out_reg_10_ ( .D(u2_N86), .CK(clk), .QN(n4490) );
  DFF_X1 u5_prod_reg_68_ ( .D(u5_prod1[68]), .CK(clk), .Q(prod[68]), .QN(n4480) );
  DFF_X1 u5_prod_reg_61_ ( .D(u5_prod1[61]), .CK(clk), .Q(prod[61]), .QN(n4479) );
  DFF_X1 u2_exp_out_reg_9_ ( .D(u2_N85), .CK(clk), .QN(n4359) );
  DFF_X1 u2_exp_out_reg_1_ ( .D(u2_N77), .CK(clk), .QN(n4358) );
  DFF_X1 u1_sign_reg ( .D(u1_sign_d), .CK(clk), .Q(sign_fasu), .QN(n4356) );
  DFF_X1 u2_exp_out_reg_0_ ( .D(u2_N76), .CK(clk), .QN(n4319) );
  DFF_X1 u5_prod1_reg_52_ ( .D(u5_N52), .CK(clk), .Q(u5_prod1[52]) );
  DFF_X1 u5_prod1_reg_101_ ( .D(u5_N101), .CK(clk), .Q(u5_prod1[101]) );
  NAND2_X2 U3379 ( .A1(n5232), .A2(n5231), .ZN(fract_denorm[52]) );
  NAND2_X2 U3380 ( .A1(n5230), .A2(n5229), .ZN(fract_denorm[51]) );
  NAND2_X2 U3381 ( .A1(fract_out_q[55]), .A2(net63509), .ZN(n5109) );
  NAND2_X2 U3382 ( .A1(fract_out_q[54]), .A2(net63509), .ZN(n5112) );
  INV_X4 U3383 ( .A(remainder[55]), .ZN(n5757) );
  NOR2_X4 U3384 ( .A1(remainder[52]), .A2(remainder[51]), .ZN(n5735) );
  INV_X8 U3385 ( .A(n6837), .ZN(n4770) );
  BUF_X32 U3386 ( .A(n4805), .Z(n4270) );
  INV_X1 U3387 ( .A(n4820), .ZN(n4271) );
  INV_X4 U3388 ( .A(n4825), .ZN(n4837) );
  INV_X8 U3389 ( .A(n4812), .ZN(n4813) );
  NAND2_X1 U3390 ( .A1(u4_div_exp1_6_), .A2(u4_div_exp1_5_), .ZN(net59064) );
  NAND3_X1 U3391 ( .A1(net58642), .A2(net58643), .A3(net58644), .ZN(net58641)
         );
  NOR3_X2 U3392 ( .A1(net59352), .A2(net58642), .A3(net59356), .ZN(net59348)
         );
  INV_X4 U3393 ( .A(net59503), .ZN(net58642) );
  INV_X4 U3394 ( .A(net60051), .ZN(n4510) );
  NAND2_X1 U3395 ( .A1(n5647), .A2(n5646), .ZN(net59579) );
  NOR2_X1 U3396 ( .A1(net63287), .A2(n5646), .ZN(n5636) );
  INV_X2 U3397 ( .A(u4_div_exp2_5_), .ZN(net58729) );
  INV_X1 U3398 ( .A(net58700), .ZN(net59644) );
  NOR2_X1 U3399 ( .A1(n6010), .A2(net59541), .ZN(n5670) );
  NOR2_X1 U3400 ( .A1(n4308), .A2(net59541), .ZN(n5656) );
  OAI21_X2 U3401 ( .B1(n5622), .B2(net59543), .A(net59541), .ZN(n5629) );
  AOI22_X1 U3402 ( .A1(net59600), .A2(div_opa_ldz_r2[2]), .B1(net59578), .B2(
        u4_fi_ldz_2_), .ZN(n5665) );
  AOI22_X1 U3403 ( .A1(net59600), .A2(div_opa_ldz_r2[4]), .B1(net59578), .B2(
        u4_fi_ldz_4_), .ZN(n5648) );
  OAI221_X4 U3404 ( .B1(net59347), .B2(net59641), .C1(net58440), .C2(net59590), 
        .A(net59642), .ZN(net59578) );
  NAND4_X1 U3405 ( .A1(net58700), .A2(net58701), .A3(n6010), .A4(n6009), .ZN(
        n6017) );
  INV_X4 U3406 ( .A(net59592), .ZN(net59641) );
  INV_X16 U3407 ( .A(net63555), .ZN(net63553) );
  NAND2_X2 U3408 ( .A1(n4273), .A2(n4274), .ZN(n4272) );
  AND3_X4 U3409 ( .A1(n2528), .A2(n2530), .A3(n2529), .ZN(n4273) );
  AND3_X4 U3410 ( .A1(n3650), .A2(n3652), .A3(n3654), .ZN(n4274) );
  NAND3_X4 U3411 ( .A1(n5153), .A2(n5152), .A3(n5151), .ZN(fract_denorm[85])
         );
  NAND3_X2 U3412 ( .A1(n4520), .A2(net60192), .A3(net60196), .ZN(n4533) );
  BUF_X4 U3413 ( .A(net60093), .Z(n4520) );
  OR2_X2 U3414 ( .A1(net33547), .A2(net59322), .ZN(n4275) );
  NOR2_X4 U3415 ( .A1(net60159), .A2(n4277), .ZN(n4276) );
  INV_X32 U3416 ( .A(net60344), .ZN(n4277) );
  INV_X8 U3417 ( .A(net60159), .ZN(net60085) );
  AOI21_X1 U3418 ( .B1(net59589), .B2(net59590), .A(net59591), .ZN(net59582)
         );
  INV_X32 U3419 ( .A(net66894), .ZN(net66897) );
  AOI22_X2 U3420 ( .A1(fract_out_q[53]), .A2(net63507), .B1(quo[52]), .B2(
        net66895), .ZN(n5121) );
  AOI22_X2 U3421 ( .A1(fract_out_q[47]), .A2(net63507), .B1(quo[46]), .B2(
        net66895), .ZN(n4680) );
  NAND2_X4 U3422 ( .A1(net59192), .A2(net59193), .ZN(net59169) );
  OAI21_X2 U3423 ( .B1(net58988), .B2(net58970), .A(net58971), .ZN(net58771)
         );
  INV_X4 U3424 ( .A(net60354), .ZN(net59429) );
  NAND2_X2 U3425 ( .A1(fpu_op_r3[1]), .A2(n4366), .ZN(net60697) );
  NAND4_X2 U3426 ( .A1(n4607), .A2(net58981), .A3(net58983), .A4(net58985), 
        .ZN(net59068) );
  AOI21_X4 U3427 ( .B1(net59342), .B2(net59008), .A(net59343), .ZN(net59311)
         );
  NOR3_X1 U3428 ( .A1(net58987), .A2(net59072), .A3(net58972), .ZN(net59071)
         );
  NAND3_X4 U3429 ( .A1(net58637), .A2(n4279), .A3(n4280), .ZN(n4278) );
  INV_X8 U3430 ( .A(n4278), .ZN(net58950) );
  INV_X32 U3431 ( .A(net58966), .ZN(n4279) );
  INV_X32 U3432 ( .A(n4532), .ZN(n4280) );
  NAND2_X4 U3433 ( .A1(net58991), .A2(net58633), .ZN(n4281) );
  NAND2_X4 U3434 ( .A1(net58991), .A2(net58633), .ZN(n4282) );
  NOR3_X2 U3435 ( .A1(net59981), .A2(net59912), .A3(net59975), .ZN(net60101)
         );
  NAND4_X4 U3436 ( .A1(n4609), .A2(net60119), .A3(net60120), .A4(net60121), 
        .ZN(net59981) );
  NAND2_X2 U3437 ( .A1(net58950), .A2(net58953), .ZN(net58952) );
  NAND2_X1 U3438 ( .A1(u4_exp_in_pl1_8_), .A2(net59568), .ZN(n5625) );
  INV_X1 U3439 ( .A(net59568), .ZN(net59651) );
  INV_X4 U3440 ( .A(net59590), .ZN(net59662) );
  NAND4_X2 U3441 ( .A1(net59641), .A2(net59026), .A3(net58926), .A4(net59664), 
        .ZN(n4552) );
  INV_X32 U3442 ( .A(net66894), .ZN(net66895) );
  INV_X32 U3443 ( .A(net60468), .ZN(net66894) );
  INV_X4 U3444 ( .A(n4749), .ZN(n4750) );
  INV_X2 U3445 ( .A(n4416), .ZN(n4284) );
  AND2_X2 U3446 ( .A1(u1_adj_op_out_sft_1_), .A2(n7138), .ZN(n4285) );
  AND2_X2 U3447 ( .A1(n4406), .A2(n6915), .ZN(n4286) );
  NOR2_X1 U3448 ( .A1(n3731), .A2(net59222), .ZN(net59221) );
  NOR2_X2 U3449 ( .A1(net59208), .A2(net58997), .ZN(n5818) );
  NOR2_X1 U3450 ( .A1(u4_fi_ldz_2_), .A2(u4_fi_ldz_3_), .ZN(net59209) );
  AOI21_X2 U3451 ( .B1(n4645), .B2(net59423), .A(n3865), .ZN(net59243) );
  AOI21_X2 U3452 ( .B1(net59424), .B2(n4646), .A(net59426), .ZN(n4645) );
  AOI211_X2 U3453 ( .C1(net59012), .C2(net59013), .A(net59014), .B(n4704), 
        .ZN(n4703) );
  NOR2_X2 U3454 ( .A1(n4705), .A2(net59017), .ZN(n4704) );
  AOI211_X1 U3455 ( .C1(n4700), .C2(n4701), .A(n4702), .B(n4468), .ZN(n4699)
         );
  NOR2_X1 U3456 ( .A1(u4_exp_out_8_), .A2(net59010), .ZN(n4701) );
  NOR2_X1 U3457 ( .A1(rmode_r3[0]), .A2(net58935), .ZN(n4557) );
  OAI21_X2 U3458 ( .B1(n5524), .B2(n5613), .A(n5523), .ZN(n5525) );
  NOR2_X1 U3459 ( .A1(div_opa_ldz_r2[1]), .A2(n4852), .ZN(n5524) );
  NOR4_X2 U3460 ( .A1(net60305), .A2(fract_denorm[91]), .A3(fract_denorm[90]), 
        .A4(fract_denorm[92]), .ZN(net59428) );
  NAND3_X2 U3461 ( .A1(n5410), .A2(n5412), .A3(n5318), .ZN(net60289) );
  INV_X8 U3462 ( .A(net60006), .ZN(net60022) );
  AOI21_X1 U3463 ( .B1(net58994), .B2(net58995), .A(net58996), .ZN(net58993)
         );
  AOI211_X2 U3464 ( .C1(net58998), .C2(n4697), .A(n4698), .B(n4699), .ZN(n4696) );
  AOI21_X2 U3465 ( .B1(net59093), .B2(net66871), .A(n5860), .ZN(n5861) );
  OAI21_X1 U3466 ( .B1(u4_fi_ldz_3_), .B2(n5496), .A(u4_fi_ldz_4_), .ZN(
        net59901) );
  INV_X4 U3467 ( .A(n4388), .ZN(net66835) );
  NAND3_X2 U3468 ( .A1(n5555), .A2(n5554), .A3(n5553), .ZN(u4_shift_right[6])
         );
  NAND3_X2 U3469 ( .A1(net59020), .A2(net59021), .A3(n4601), .ZN(net59019) );
  NOR2_X1 U3470 ( .A1(n4602), .A2(u4_fi_ldz_2a_5_), .ZN(n4601) );
  NOR2_X2 U3471 ( .A1(div_opa_ldz_r2[3]), .A2(net66851), .ZN(n5530) );
  NOR2_X1 U3472 ( .A1(exp_ovf_r_0_), .A2(net58550), .ZN(n5620) );
  NOR2_X1 U3473 ( .A1(fract_denorm[86]), .A2(n5412), .ZN(n5413) );
  NOR2_X1 U3474 ( .A1(fract_denorm[54]), .A2(n4688), .ZN(net60058) );
  NOR3_X1 U3475 ( .A1(net59923), .A2(fract_denorm[70]), .A3(n4662), .ZN(
        net60060) );
  NOR3_X2 U3476 ( .A1(n5414), .A2(n8514), .A3(net59927), .ZN(n5415) );
  NOR3_X1 U3477 ( .A1(n4843), .A2(n5547), .A3(n4384), .ZN(n5541) );
  AOI21_X1 U3478 ( .B1(n5548), .B2(n4848), .A(n4843), .ZN(n5540) );
  NAND3_X2 U3479 ( .A1(net60236), .A2(net59945), .A3(net60167), .ZN(net60235)
         );
  NOR2_X2 U3480 ( .A1(net59988), .A2(n5435), .ZN(n5440) );
  NAND3_X2 U3481 ( .A1(n5138), .A2(n5137), .A3(n5136), .ZN(fract_denorm[90])
         );
  NAND3_X2 U3482 ( .A1(n5108), .A2(n5107), .A3(n5106), .ZN(fract_denorm[79])
         );
  NOR3_X2 U3483 ( .A1(net58585), .A2(net58586), .A3(net58587), .ZN(n6064) );
  NAND3_X2 U3484 ( .A1(n5010), .A2(n4344), .A3(n4313), .ZN(n6441) );
  NAND3_X2 U3485 ( .A1(n5692), .A2(n5691), .A3(n5778), .ZN(n5693) );
  NOR2_X2 U3486 ( .A1(net66851), .A2(n5493), .ZN(n5491) );
  NAND3_X1 U3487 ( .A1(n8523), .A2(n5461), .A3(n5460), .ZN(n5462) );
  NAND3_X1 U3488 ( .A1(n8519), .A2(n5459), .A3(n4320), .ZN(n5463) );
  NAND3_X1 U3489 ( .A1(net59326), .A2(net60220), .A3(net33552), .ZN(net60215)
         );
  AOI21_X1 U3490 ( .B1(net60173), .B2(net60174), .A(net59697), .ZN(n5391) );
  NOR2_X1 U3491 ( .A1(fract_denorm[99]), .A2(n4597), .ZN(net60173) );
  NAND3_X2 U3492 ( .A1(n5340), .A2(n5339), .A3(net60279), .ZN(n5381) );
  INV_X8 U3493 ( .A(n4379), .ZN(n4852) );
  NAND3_X2 U3494 ( .A1(net58783), .A2(n5966), .A3(n5965), .ZN(n5967) );
  NAND3_X1 U3495 ( .A1(net58787), .A2(net58636), .A3(n4405), .ZN(n5966) );
  NAND3_X1 U3496 ( .A1(n5964), .A2(net58644), .A3(net58636), .ZN(n5965) );
  NOR2_X1 U3497 ( .A1(net58530), .A2(net58475), .ZN(net58529) );
  NAND3_X1 U3498 ( .A1(n6116), .A2(n6115), .A3(n6114), .ZN(n6098) );
  NAND3_X1 U3499 ( .A1(n4854), .A2(u2_exp_tmp4_10_), .A3(n6273), .ZN(n6281) );
  NAND3_X2 U3500 ( .A1(n4927), .A2(n4316), .A3(n4420), .ZN(n4999) );
  INV_X8 U3501 ( .A(n4383), .ZN(n4846) );
  INV_X8 U3502 ( .A(n4307), .ZN(net66863) );
  INV_X16 U3503 ( .A(n4322), .ZN(net63295) );
  NOR2_X2 U3504 ( .A1(exp_ovf_r_0_), .A2(net66835), .ZN(net59054) );
  INV_X4 U3505 ( .A(n4876), .ZN(n4894) );
  NAND3_X2 U3506 ( .A1(n4596), .A2(n4597), .A3(n4595), .ZN(net60354) );
  AOI211_X2 U3507 ( .C1(n5721), .C2(n5720), .A(n5719), .B(n5718), .ZN(net59424) );
  AOI21_X1 U3508 ( .B1(n5716), .B2(n5715), .A(n5714), .ZN(n5721) );
  NOR3_X2 U3509 ( .A1(n5656), .A2(n5655), .A3(n5654), .ZN(n5659) );
  NOR2_X1 U3510 ( .A1(net58935), .A2(n5779), .ZN(n5655) );
  NOR2_X2 U3511 ( .A1(net59982), .A2(net59981), .ZN(net59980) );
  NAND3_X2 U3512 ( .A1(opas_r2), .A2(net58644), .A3(n4405), .ZN(n5872) );
  OAI21_X2 U3513 ( .B1(n5687), .B2(net59551), .A(n5686), .ZN(n5871) );
  NOR2_X2 U3514 ( .A1(n4846), .A2(net59553), .ZN(n5686) );
  NOR2_X2 U3515 ( .A1(n5685), .A2(net59555), .ZN(n5687) );
  NOR2_X1 U3516 ( .A1(n4850), .A2(n4851), .ZN(n6009) );
  NOR2_X2 U3517 ( .A1(n7213), .A2(n7212), .ZN(n6018) );
  NOR2_X1 U3518 ( .A1(n4848), .A2(net58688), .ZN(n6020) );
  NOR3_X2 U3519 ( .A1(net58711), .A2(n8243), .A3(n8242), .ZN(n6005) );
  INV_X16 U3520 ( .A(n4878), .ZN(n4876) );
  INV_X16 U3521 ( .A(net63521), .ZN(net63517) );
  NOR3_X2 U3522 ( .A1(net60151), .A2(net60152), .A3(net60153), .ZN(net60136)
         );
  NAND4_X2 U3523 ( .A1(net60054), .A2(net60055), .A3(net60056), .A4(net60057), 
        .ZN(net59913) );
  NAND3_X1 U3524 ( .A1(n5460), .A2(n8522), .A3(n5408), .ZN(net60054) );
  NOR2_X2 U3525 ( .A1(n4591), .A2(net33647), .ZN(n4592) );
  INV_X8 U3526 ( .A(net59973), .ZN(net60072) );
  NOR2_X1 U3527 ( .A1(n5547), .A2(n4843), .ZN(n5550) );
  NOR2_X1 U3528 ( .A1(n5548), .A2(n4843), .ZN(n5549) );
  INV_X4 U3529 ( .A(net58952), .ZN(net63555) );
  AOI21_X1 U3530 ( .B1(net58932), .B2(net58957), .A(net58624), .ZN(net58956)
         );
  NOR2_X2 U3531 ( .A1(net59171), .A2(n5814), .ZN(n5815) );
  NOR2_X1 U3532 ( .A1(net59112), .A2(net59195), .ZN(net59228) );
  AOI21_X1 U3533 ( .B1(u4_exp_out_8_), .B2(net59084), .A(net59212), .ZN(
        net59201) );
  NOR2_X1 U3534 ( .A1(u4_exp_out_0_), .A2(net59083), .ZN(net59111) );
  NOR2_X2 U3535 ( .A1(net59142), .A2(net59143), .ZN(n5849) );
  NOR2_X2 U3536 ( .A1(net59144), .A2(net59145), .ZN(net59143) );
  AOI21_X1 U3537 ( .B1(u4_exp_out_3_), .B2(net59118), .A(n4369), .ZN(n4615) );
  NAND3_X2 U3538 ( .A1(n4990), .A2(n6833), .A3(n4943), .ZN(n5040) );
  NOR2_X1 U3539 ( .A1(fracta_mul[5]), .A2(fracta_mul[4]), .ZN(n4943) );
  NOR2_X1 U3540 ( .A1(fracta_mul[25]), .A2(fracta_mul[26]), .ZN(n4938) );
  NOR2_X1 U3541 ( .A1(fracta_mul[27]), .A2(fracta_mul[24]), .ZN(n4939) );
  NAND3_X2 U3542 ( .A1(n5639), .A2(n5638), .A3(n5637), .ZN(u4_shift_left[6])
         );
  NOR2_X1 U3543 ( .A1(net59918), .A2(net59919), .ZN(net59917) );
  NOR2_X2 U3544 ( .A1(n5465), .A2(net59927), .ZN(n5466) );
  NOR3_X2 U3545 ( .A1(net59911), .A2(net59912), .A3(net59913), .ZN(net59910)
         );
  NAND3_X2 U3546 ( .A1(net60078), .A2(n5405), .A3(n5404), .ZN(net59974) );
  AOI21_X2 U3547 ( .B1(net60231), .B2(net60106), .A(net60232), .ZN(net60223)
         );
  NAND3_X1 U3548 ( .A1(net60085), .A2(net60230), .A3(net33584), .ZN(n5380) );
  INV_X4 U3549 ( .A(net60696), .ZN(net60695) );
  NOR2_X1 U3550 ( .A1(n5520), .A2(n4843), .ZN(n5522) );
  NOR2_X1 U3551 ( .A1(n5681), .A2(n4843), .ZN(n5521) );
  NOR2_X2 U3552 ( .A1(net58609), .A2(n6095), .ZN(n6041) );
  NOR3_X1 U3553 ( .A1(n4466), .A2(n6442), .A3(n6441), .ZN(n6443) );
  NAND3_X2 U3554 ( .A1(n4996), .A2(n4929), .A3(n4439), .ZN(n4982) );
  NAND3_X1 U3555 ( .A1(fracta_mul[21]), .A2(n4951), .A3(n4289), .ZN(n4992) );
  AOI21_X2 U3556 ( .B1(n5567), .B2(n5566), .A(n5565), .ZN(n5576) );
  INV_X8 U3557 ( .A(net44903), .ZN(net63333) );
  AOI21_X1 U3558 ( .B1(n4657), .B2(net59717), .A(net59863), .ZN(net59715) );
  NOR3_X2 U3559 ( .A1(n4659), .A2(net59555), .A3(net58688), .ZN(net59707) );
  NAND3_X2 U3560 ( .A1(net60311), .A2(net60312), .A3(n5332), .ZN(n5342) );
  AOI21_X2 U3561 ( .B1(n4321), .B2(net60318), .A(n4370), .ZN(net60311) );
  NAND3_X2 U3562 ( .A1(net59826), .A2(n5489), .A3(n5488), .ZN(u4_exp_in_mi1_6_) );
  INV_X4 U3563 ( .A(exp_r[9]), .ZN(net66870) );
  INV_X4 U3564 ( .A(net66875), .ZN(net58636) );
  NOR3_X2 U3565 ( .A1(n6098), .A2(net58533), .A3(n6097), .ZN(n6102) );
  NOR3_X2 U3566 ( .A1(net58523), .A2(net58524), .A3(net58525), .ZN(n6100) );
  OAI21_X2 U3567 ( .B1(n6272), .B2(n6467), .A(n6281), .ZN(n6278) );
  INV_X8 U3568 ( .A(n4326), .ZN(net66839) );
  INV_X4 U3569 ( .A(net59703), .ZN(net58719) );
  OAI21_X2 U3570 ( .B1(n4692), .B2(n4505), .A(net59888), .ZN(u4_exp_in_mi1_9_)
         );
  INV_X8 U3571 ( .A(n4306), .ZN(net66875) );
  INV_X8 U3572 ( .A(u4_exp_out_0_), .ZN(net45071) );
  NOR2_X1 U3573 ( .A1(net63287), .A2(net58506), .ZN(net58818) );
  NOR2_X1 U3574 ( .A1(opb_r[55]), .A2(n4390), .ZN(n6712) );
  NOR2_X1 U3575 ( .A1(u4_exp_in_pl1_1_), .A2(u4_exp_in_mi1_11_), .ZN(net59593)
         );
  NOR3_X1 U3576 ( .A1(net60128), .A2(fract_denorm[92]), .A3(net60094), .ZN(
        n4683) );
  NOR2_X2 U3577 ( .A1(net33565), .A2(net60130), .ZN(n4681) );
  AOI211_X1 U3578 ( .C1(net58651), .C2(n4404), .A(net59354), .B(net59054), 
        .ZN(net59353) );
  OAI21_X1 U3579 ( .B1(net66835), .B2(net59032), .A(net63287), .ZN(net59354)
         );
  NOR2_X1 U3580 ( .A1(net33546), .A2(net59324), .ZN(n4561) );
  NOR2_X1 U3581 ( .A1(net59322), .A2(net59323), .ZN(net59321) );
  NAND3_X2 U3582 ( .A1(net60186), .A2(net59423), .A3(net60187), .ZN(net60182)
         );
  NAND3_X2 U3583 ( .A1(n5418), .A2(n5417), .A3(n8511), .ZN(n5419) );
  NOR2_X2 U3584 ( .A1(fract_denorm[52]), .A2(n4524), .ZN(n5421) );
  NOR2_X1 U3585 ( .A1(n4595), .A2(net60038), .ZN(net60032) );
  NOR2_X1 U3586 ( .A1(net60048), .A2(net59991), .ZN(net60047) );
  NAND3_X2 U3587 ( .A1(net60049), .A2(net60050), .A3(net33573), .ZN(n5424) );
  INV_X16 U3588 ( .A(n7134), .ZN(n4878) );
  NOR2_X1 U3589 ( .A1(div_opa_ldz_r2[2]), .A2(n4851), .ZN(n5527) );
  AOI21_X1 U3590 ( .B1(n4558), .B2(n4559), .A(opas_r2), .ZN(n4556) );
  NOR3_X1 U3591 ( .A1(net59332), .A2(net59333), .A3(net59334), .ZN(n4558) );
  NOR2_X2 U3592 ( .A1(net59318), .A2(n4560), .ZN(n4559) );
  NAND3_X1 U3593 ( .A1(net59335), .A2(net59336), .A3(net59337), .ZN(net59334)
         );
  NOR3_X1 U3594 ( .A1(n5451), .A2(fract_denorm[72]), .A3(n5427), .ZN(n5428) );
  NOR3_X1 U3595 ( .A1(net59952), .A2(fract_denorm[88]), .A3(n5426), .ZN(n5429)
         );
  NOR2_X1 U3596 ( .A1(fract_denorm[56]), .A2(n5425), .ZN(n5430) );
  OAI21_X2 U3597 ( .B1(n5399), .B2(n5398), .A(net60110), .ZN(net60107) );
  NOR2_X1 U3598 ( .A1(fract_denorm[97]), .A2(net60114), .ZN(net60113) );
  NOR2_X1 U3599 ( .A1(net59233), .A2(net59029), .ZN(net59230) );
  NOR3_X1 U3600 ( .A1(n6919), .A2(n6918), .A3(n6928), .ZN(n6924) );
  NOR2_X2 U3601 ( .A1(n6953), .A2(n6979), .ZN(n6958) );
  NOR2_X2 U3602 ( .A1(n6930), .A2(n6985), .ZN(n6937) );
  NOR2_X2 U3603 ( .A1(n6934), .A2(n6983), .ZN(n6935) );
  NOR2_X1 U3604 ( .A1(n6933), .A2(n6941), .ZN(n6936) );
  NOR2_X1 U3605 ( .A1(net59337), .A2(net59328), .ZN(n4562) );
  NOR3_X2 U3606 ( .A1(net59998), .A2(net59999), .A3(n4717), .ZN(net59997) );
  NAND3_X2 U3607 ( .A1(n6332), .A2(n6336), .A3(n6401), .ZN(n6329) );
  NOR2_X1 U3608 ( .A1(prod[63]), .A2(prod[62]), .ZN(n6082) );
  NOR2_X1 U3609 ( .A1(prod[65]), .A2(prod[64]), .ZN(n6083) );
  NOR2_X1 U3610 ( .A1(prod[66]), .A2(prod[67]), .ZN(n6084) );
  NOR2_X1 U3611 ( .A1(prod[103]), .A2(prod[104]), .ZN(n6073) );
  NOR3_X1 U3612 ( .A1(prod[100]), .A2(prod[102]), .A3(prod[101]), .ZN(n6072)
         );
  NOR3_X1 U3613 ( .A1(prod[87]), .A2(prod[88]), .A3(prod[89]), .ZN(n6070) );
  NOR3_X1 U3614 ( .A1(prod[75]), .A2(prod[82]), .A3(prod[81]), .ZN(n6068) );
  NOR3_X1 U3615 ( .A1(prod[54]), .A2(prod[56]), .A3(prod[55]), .ZN(n6080) );
  NOR3_X1 U3616 ( .A1(prod[8]), .A2(prod[52]), .A3(prod[53]), .ZN(n6079) );
  NOR3_X1 U3617 ( .A1(prod[0]), .A2(prod[6]), .A3(prod[5]), .ZN(n6078) );
  NOR2_X1 U3618 ( .A1(prod[74]), .A2(prod[73]), .ZN(n6087) );
  NOR2_X1 U3619 ( .A1(prod[72]), .A2(prod[71]), .ZN(n6086) );
  NOR2_X1 U3620 ( .A1(prod[70]), .A2(prod[69]), .ZN(n6085) );
  AOI21_X2 U3621 ( .B1(n6006), .B2(n6005), .A(n6004), .ZN(n6007) );
  NOR2_X1 U3622 ( .A1(net66835), .A2(net58664), .ZN(n6033) );
  NOR2_X1 U3623 ( .A1(net58550), .A2(n4404), .ZN(net58664) );
  NAND3_X2 U3624 ( .A1(n2534), .A2(n2536), .A3(n2535), .ZN(n5705) );
  NAND3_X2 U3625 ( .A1(n3666), .A2(n3724), .A3(n3664), .ZN(n5706) );
  NAND3_X2 U3626 ( .A1(n3675), .A2(n3677), .A3(n3679), .ZN(n5711) );
  NAND3_X2 U3627 ( .A1(n2537), .A2(n2539), .A3(n2538), .ZN(n5710) );
  NOR2_X1 U3628 ( .A1(net58636), .A2(net59088), .ZN(net59123) );
  NAND3_X2 U3629 ( .A1(net59034), .A2(net63291), .A3(net58932), .ZN(net59033)
         );
  INV_X4 U3630 ( .A(n6708), .ZN(n4868) );
  INV_X16 U3631 ( .A(n4906), .ZN(n4904) );
  NOR2_X1 U3632 ( .A1(fracta_mul[17]), .A2(fracta_mul[16]), .ZN(n4932) );
  NOR2_X1 U3633 ( .A1(fracta_mul[19]), .A2(fracta_mul[18]), .ZN(n4933) );
  NAND3_X2 U3634 ( .A1(n4940), .A2(n6444), .A3(n4417), .ZN(n4941) );
  NAND3_X2 U3635 ( .A1(n5102), .A2(n5101), .A3(n5100), .ZN(fract_denorm[77])
         );
  NOR2_X2 U3636 ( .A1(n5619), .A2(n5618), .ZN(net59679) );
  NOR2_X1 U3637 ( .A1(n4852), .A2(n4843), .ZN(n5618) );
  NOR2_X1 U3638 ( .A1(n5557), .A2(net57241), .ZN(n5558) );
  NOR2_X1 U3639 ( .A1(n6336), .A2(n6409), .ZN(n6331) );
  AOI21_X2 U3640 ( .B1(net58648), .B2(net58649), .A(net58650), .ZN(n6037) );
  NOR2_X1 U3641 ( .A1(net66835), .A2(net58651), .ZN(net58649) );
  NAND3_X2 U3642 ( .A1(net63579), .A2(n5956), .A3(n5955), .ZN(n6058) );
  NOR2_X2 U3643 ( .A1(net59107), .A2(n5853), .ZN(n5856) );
  AOI21_X1 U3644 ( .B1(net59093), .B2(n4851), .A(n5847), .ZN(n5848) );
  NAND3_X2 U3645 ( .A1(n4444), .A2(n4349), .A3(n4317), .ZN(n4252) );
  NOR3_X2 U3646 ( .A1(opa_r1[59]), .A2(opa_r1[55]), .A3(opa_r1[56]), .ZN(n6476) );
  NOR2_X1 U3647 ( .A1(u1_N232), .A2(n6736), .ZN(n6749) );
  NOR2_X1 U3648 ( .A1(fracta_mul[23]), .A2(n6440), .ZN(n6445) );
  NOR3_X1 U3649 ( .A1(fracta_mul[29]), .A2(fracta_mul[28]), .A3(fracta_mul[31]), .ZN(n6447) );
  NOR3_X1 U3650 ( .A1(fracta_mul[37]), .A2(fracta_mul[36]), .A3(fracta_mul[38]), .ZN(n6446) );
  NOR2_X1 U3651 ( .A1(fracta_mul[20]), .A2(fracta_mul[30]), .ZN(n6448) );
  NOR2_X1 U3652 ( .A1(fracta_mul[45]), .A2(n6450), .ZN(n6452) );
  NAND3_X1 U3653 ( .A1(opa_r[61]), .A2(n4853), .A3(opa_r[60]), .ZN(n3081) );
  NAND3_X1 U3654 ( .A1(opa_r[58]), .A2(opa_r[57]), .A3(opa_r[59]), .ZN(n7141)
         );
  NOR2_X2 U3655 ( .A1(n4465), .A2(n4350), .ZN(n6456) );
  NOR3_X2 U3656 ( .A1(n3108), .A2(n3109), .A3(n3110), .ZN(n3098) );
  NOR2_X1 U3657 ( .A1(n5020), .A2(n5068), .ZN(n5021) );
  NOR2_X1 U3658 ( .A1(fracta_mul[14]), .A2(n4336), .ZN(n5022) );
  OAI21_X1 U3659 ( .B1(fracta_mul[46]), .B2(n4290), .A(n4302), .ZN(n5018) );
  NAND3_X2 U3660 ( .A1(n4980), .A2(n5038), .A3(n4998), .ZN(n5035) );
  NOR2_X1 U3661 ( .A1(n4997), .A2(n4433), .ZN(n4998) );
  NAND3_X1 U3662 ( .A1(fracta_mul[41]), .A2(n4996), .A3(n5010), .ZN(n5034) );
  NAND3_X1 U3663 ( .A1(n4924), .A2(n4342), .A3(n4311), .ZN(n6442) );
  NAND3_X1 U3664 ( .A1(fracta_mul[29]), .A2(n4961), .A3(n4419), .ZN(n5033) );
  NOR3_X2 U3665 ( .A1(n4954), .A2(n4953), .A3(n4417), .ZN(n5017) );
  NAND3_X1 U3666 ( .A1(fracta_mul[24]), .A2(n4955), .A3(n4421), .ZN(n5012) );
  NOR2_X2 U3667 ( .A1(n5696), .A2(n5695), .ZN(n5697) );
  OAI21_X2 U3668 ( .B1(n5487), .B2(net59551), .A(n5486), .ZN(u4_exp_in_mi1_7_)
         );
  INV_X4 U3669 ( .A(exp_r[6]), .ZN(n4847) );
  NAND3_X2 U3670 ( .A1(n5345), .A2(n5344), .A3(n5343), .ZN(u4_fi_ldz_4_) );
  AOI211_X1 U3671 ( .C1(n5335), .C2(net60092), .A(net60300), .B(net60301), 
        .ZN(n5345) );
  NOR3_X2 U3672 ( .A1(net60283), .A2(net60284), .A3(net60285), .ZN(n5344) );
  INV_X4 U3673 ( .A(exp_r[4]), .ZN(n4849) );
  AOI211_X2 U3674 ( .C1(net59914), .C2(n5469), .A(n5468), .B(net59917), .ZN(
        n5470) );
  NOR3_X1 U3675 ( .A1(net60221), .A2(n5381), .A3(n5468), .ZN(n5407) );
  INV_X4 U3676 ( .A(exp_r[3]), .ZN(net66850) );
  NOR2_X1 U3677 ( .A1(n4505), .A2(net59433), .ZN(n5717) );
  NAND3_X2 U3678 ( .A1(net59695), .A2(opas_r2), .A3(net58780), .ZN(n7162) );
  NOR2_X2 U3679 ( .A1(net63287), .A2(n6051), .ZN(n6047) );
  INV_X4 U3680 ( .A(n4734), .ZN(n6120) );
  INV_X4 U3681 ( .A(u4_fract_out_pl1_27_), .ZN(n4735) );
  NAND3_X2 U3682 ( .A1(net63577), .A2(n5888), .A3(n5887), .ZN(n5889) );
  NAND3_X2 U3683 ( .A1(net63577), .A2(n5885), .A3(n5884), .ZN(n5886) );
  INV_X4 U3684 ( .A(n4727), .ZN(n6833) );
  NOR2_X1 U3685 ( .A1(u2_N16), .A2(n6427), .ZN(n6435) );
  NOR3_X2 U3686 ( .A1(n6426), .A2(n6425), .A3(n6424), .ZN(n6436) );
  NOR2_X2 U3687 ( .A1(n6433), .A2(n6432), .ZN(n6434) );
  NOR2_X1 U3688 ( .A1(n6430), .A2(n6429), .ZN(n6431) );
  NOR2_X1 U3689 ( .A1(u2_N28), .A2(n6414), .ZN(n6422) );
  NOR3_X2 U3690 ( .A1(n6413), .A2(n6412), .A3(n6411), .ZN(n6423) );
  NOR2_X2 U3691 ( .A1(n6420), .A2(n6419), .ZN(n6421) );
  NOR2_X1 U3692 ( .A1(n6417), .A2(n6416), .ZN(n6418) );
  OAI21_X1 U3693 ( .B1(u2_N157), .B2(n7153), .A(n6462), .ZN(n6465) );
  NOR2_X2 U3694 ( .A1(u1_fracta_eq_fractb), .A2(n3063), .ZN(n3064) );
  NAND3_X2 U3695 ( .A1(net58812), .A2(net58936), .A3(net58937), .ZN(net57282)
         );
  OAI21_X2 U3696 ( .B1(n5877), .B2(n5880), .A(opa_00), .ZN(net58936) );
  AOI21_X2 U3697 ( .B1(net58938), .B2(opa_inf), .A(net58939), .ZN(net58937) );
  AOI21_X1 U3698 ( .B1(n4987), .B2(n4986), .A(n4985), .ZN(n4995) );
  NOR2_X2 U3699 ( .A1(n4999), .A2(n4475), .ZN(n4985) );
  NAND3_X1 U3700 ( .A1(fracta_mul[6]), .A2(n4980), .A3(n4937), .ZN(n4981) );
  NAND3_X1 U3701 ( .A1(n4927), .A2(n4316), .A3(fracta_mul[44]), .ZN(n4973) );
  NAND3_X1 U3702 ( .A1(fracta_mul[28]), .A2(n4972), .A3(n4971), .ZN(n4974) );
  OAI21_X1 U3703 ( .B1(n4969), .B2(n5067), .A(n4968), .ZN(n4978) );
  AOI21_X1 U3704 ( .B1(fracta_mul[8]), .B2(n4433), .A(n4997), .ZN(n4969) );
  NAND3_X1 U3705 ( .A1(n5039), .A2(n4967), .A3(fracta_mul[12]), .ZN(n4968) );
  NOR2_X1 U3706 ( .A1(net58728), .A2(n7203), .ZN(n5994) );
  AOI21_X2 U3707 ( .B1(net59275), .B2(n5799), .A(n5798), .ZN(n5801) );
  NOR2_X2 U3708 ( .A1(net44696), .A2(net57276), .ZN(n4667) );
  NOR2_X1 U3709 ( .A1(n6343), .A2(n6342), .ZN(n6346) );
  AOI21_X1 U3710 ( .B1(n6361), .B2(n6360), .A(n6359), .ZN(n6362) );
  AOI222_X1 U3711 ( .A1(u2_exp_tmp3_7_), .A2(n6399), .B1(n4845), .B2(n8293), 
        .C1(u2_N61), .C2(n4844), .ZN(n6363) );
  OAI21_X1 U3712 ( .B1(n6357), .B2(n6358), .A(n6356), .ZN(n6360) );
  AOI21_X1 U3713 ( .B1(n6361), .B2(n6372), .A(n6371), .ZN(n6373) );
  AOI222_X1 U3714 ( .A1(u2_exp_tmp3_5_), .A2(n6399), .B1(n4845), .B2(n8295), 
        .C1(u2_N59), .C2(n4844), .ZN(n6374) );
  OAI21_X1 U3715 ( .B1(n6369), .B2(n6370), .A(n6368), .ZN(n6372) );
  NOR2_X2 U3716 ( .A1(net58506), .A2(n4548), .ZN(net58805) );
  NOR2_X1 U3717 ( .A1(net63529), .A2(n6114), .ZN(N797) );
  NOR2_X1 U3718 ( .A1(net63529), .A2(n6115), .ZN(N798) );
  NOR2_X1 U3719 ( .A1(net63529), .A2(net58495), .ZN(N802) );
  NOR2_X1 U3720 ( .A1(net63529), .A2(net58493), .ZN(N804) );
  NOR2_X1 U3721 ( .A1(net63527), .A2(net58477), .ZN(N813) );
  NOR2_X1 U3722 ( .A1(net63527), .A2(net58472), .ZN(N817) );
  NOR2_X2 U3723 ( .A1(net63523), .A2(n6124), .ZN(N824) );
  NOR2_X2 U3724 ( .A1(net63523), .A2(n6125), .ZN(N825) );
  NOR2_X2 U3725 ( .A1(net63523), .A2(n6127), .ZN(N827) );
  NOR2_X2 U3726 ( .A1(net63523), .A2(n6132), .ZN(N832) );
  NOR2_X2 U3727 ( .A1(net63523), .A2(n6134), .ZN(N834) );
  NOR2_X2 U3728 ( .A1(net63523), .A2(n6135), .ZN(N835) );
  NOR2_X2 U3729 ( .A1(net63523), .A2(n6137), .ZN(N837) );
  NOR2_X2 U3730 ( .A1(net63523), .A2(n6138), .ZN(N838) );
  NOR2_X2 U3731 ( .A1(net63523), .A2(n6140), .ZN(N840) );
  OAI21_X2 U3732 ( .B1(net58431), .B2(net58432), .A(net58433), .ZN(N899) );
  NAND3_X1 U3733 ( .A1(net58434), .A2(net63089), .A3(n6148), .ZN(net58433) );
  AOI21_X2 U3734 ( .B1(n6148), .B2(net58438), .A(n6147), .ZN(net58431) );
  NOR3_X1 U3735 ( .A1(net58780), .A2(net63293), .A3(net58781), .ZN(n4693) );
  NOR2_X2 U3736 ( .A1(net60202), .A2(n4663), .ZN(net60197) );
  NOR3_X2 U3737 ( .A1(fract_denorm[74]), .A2(fract_denorm[76]), .A3(
        fract_denorm[75]), .ZN(n5387) );
  NOR3_X1 U3738 ( .A1(n5672), .A2(n5671), .A3(n5670), .ZN(n5673) );
  NOR2_X1 U3739 ( .A1(net59588), .A2(net58935), .ZN(n5672) );
  NOR2_X1 U3740 ( .A1(net63287), .A2(net59026), .ZN(n5647) );
  NOR2_X1 U3741 ( .A1(net63293), .A2(net59070), .ZN(net59356) );
  NAND3_X1 U3742 ( .A1(net59325), .A2(net59326), .A3(net59327), .ZN(net59318)
         );
  NOR2_X1 U3743 ( .A1(net59330), .A2(net59331), .ZN(net59325) );
  NOR2_X1 U3744 ( .A1(net59328), .A2(net59329), .ZN(net59327) );
  NAND3_X1 U3745 ( .A1(net59338), .A2(net59339), .A3(net59340), .ZN(net59332)
         );
  NAND3_X2 U3746 ( .A1(n4617), .A2(n4618), .A3(n4619), .ZN(net59480) );
  NAND3_X2 U3747 ( .A1(n4620), .A2(n4621), .A3(n4622), .ZN(net59479) );
  NAND3_X2 U3748 ( .A1(n4632), .A2(n4633), .A3(n4634), .ZN(n4631) );
  NAND3_X2 U3749 ( .A1(n4635), .A2(n4636), .A3(n4637), .ZN(n4630) );
  NAND3_X2 U3750 ( .A1(n4604), .A2(net59021), .A3(net58650), .ZN(net59009) );
  NAND3_X1 U3751 ( .A1(u4_fi_ldz_2a_5_), .A2(u4_fi_ldz_2a_4_), .A3(n4605), 
        .ZN(n4604) );
  NOR2_X1 U3752 ( .A1(net63217), .A2(u4_exp_in_mi1_11_), .ZN(n4705) );
  NAND3_X2 U3753 ( .A1(n5870), .A2(n5797), .A3(net59057), .ZN(net59017) );
  NAND2_X2 U3754 ( .A1(net59101), .A2(net57231), .ZN(n4553) );
  NAND3_X2 U3755 ( .A1(n6899), .A2(n6898), .A3(n6897), .ZN(n6972) );
  NOR2_X2 U3756 ( .A1(n6713), .A2(n6712), .ZN(n6717) );
  OAI21_X1 U3757 ( .B1(n5615), .B2(n5569), .A(n5568), .ZN(n5570) );
  NOR2_X1 U3758 ( .A1(div_opa_ldz_r2[1]), .A2(n6010), .ZN(n5569) );
  NOR2_X1 U3759 ( .A1(n5664), .A2(n5663), .ZN(n5668) );
  NOR2_X1 U3760 ( .A1(net58935), .A2(n5661), .ZN(n5664) );
  INV_X4 U3761 ( .A(net59651), .ZN(n4529) );
  INV_X1 U3762 ( .A(n5791), .ZN(n4530) );
  NOR3_X1 U3763 ( .A1(n5398), .A2(n5395), .A3(fract_denorm[78]), .ZN(net60152)
         );
  NOR3_X2 U3764 ( .A1(net60154), .A2(net59919), .A3(fract_denorm[94]), .ZN(
        net60153) );
  NOR2_X1 U3765 ( .A1(n8519), .A2(n8520), .ZN(n5409) );
  NOR2_X2 U3766 ( .A1(n8525), .A2(n8523), .ZN(n5408) );
  AOI211_X2 U3767 ( .C1(n4681), .C2(n4682), .A(n4683), .B(n4684), .ZN(net60121) );
  NOR2_X2 U3768 ( .A1(net59344), .A2(net59345), .ZN(net59343) );
  NOR2_X2 U3769 ( .A1(div_opa_ldz_r2[4]), .A2(n4850), .ZN(n5532) );
  AOI21_X2 U3770 ( .B1(net60040), .B2(fract_denorm[67]), .A(n4372), .ZN(n5423)
         );
  AOI211_X2 U3771 ( .C1(n5421), .C2(fract_denorm[51]), .A(net60032), .B(n5420), 
        .ZN(n5422) );
  AOI21_X1 U3772 ( .B1(n6023), .B2(n4467), .A(net58681), .ZN(n6024) );
  NOR2_X1 U3773 ( .A1(net66875), .A2(net58673), .ZN(n6004) );
  NOR2_X2 U3774 ( .A1(u4_N6015), .A2(u4_N6014), .ZN(n4668) );
  AOI21_X2 U3775 ( .B1(net59046), .B2(net59047), .A(net58792), .ZN(net59045)
         );
  OAI21_X1 U3776 ( .B1(net66875), .B2(u4_exp_in_mi1_11_), .A(net59034), .ZN(
        net59047) );
  NOR2_X1 U3777 ( .A1(net63287), .A2(net59042), .ZN(net59041) );
  NOR3_X1 U3778 ( .A1(net58932), .A2(net58792), .A3(net58631), .ZN(net58996)
         );
  NOR2_X2 U3779 ( .A1(net59079), .A2(n5817), .ZN(net59212) );
  NOR2_X2 U3780 ( .A1(net59079), .A2(n5857), .ZN(net59097) );
  NAND3_X2 U3781 ( .A1(n6905), .A2(n6981), .A3(n6904), .ZN(n6963) );
  OAI21_X1 U3782 ( .B1(n7191), .B2(n5612), .A(n5611), .ZN(n5617) );
  NOR2_X1 U3783 ( .A1(net57241), .A2(n5715), .ZN(n5599) );
  NOR2_X1 U3784 ( .A1(net60086), .A2(net60159), .ZN(net60163) );
  NOR3_X2 U3785 ( .A1(n5377), .A2(fract_denorm[79]), .A3(n5398), .ZN(net60232)
         );
  NOR2_X1 U3786 ( .A1(fract_denorm[63]), .A2(net60237), .ZN(net60231) );
  NAND3_X2 U3787 ( .A1(n5433), .A2(n5432), .A3(n5431), .ZN(net59976) );
  AOI211_X2 U3788 ( .C1(n5441), .C2(n5430), .A(n5429), .B(n5428), .ZN(n5431)
         );
  AOI21_X1 U3789 ( .B1(net60106), .B2(fract_denorm[63]), .A(net60107), .ZN(
        net60105) );
  NOR2_X1 U3790 ( .A1(n5452), .A2(n5451), .ZN(n5453) );
  OAI21_X2 U3791 ( .B1(net59953), .B2(net59954), .A(net59955), .ZN(net59939)
         );
  NAND3_X1 U3792 ( .A1(n4515), .A2(net59950), .A3(fract_denorm[80]), .ZN(n5449) );
  NAND3_X2 U3793 ( .A1(n5222), .A2(n5221), .A3(n5220), .ZN(fract_denorm[53])
         );
  NOR3_X2 U3794 ( .A1(net58526), .A2(net58592), .A3(net58475), .ZN(net58591)
         );
  NOR3_X2 U3795 ( .A1(n6059), .A2(n6058), .A3(n6097), .ZN(n6062) );
  OAI21_X2 U3796 ( .B1(n6022), .B2(n6021), .A(net58687), .ZN(n6030) );
  AOI211_X2 U3797 ( .C1(n6020), .C2(n6019), .A(n6031), .B(n6018), .ZN(n6021)
         );
  NOR2_X2 U3798 ( .A1(n6028), .A2(n6027), .ZN(n6029) );
  NOR2_X1 U3799 ( .A1(net58673), .A2(net58674), .ZN(n6027) );
  NOR2_X1 U3800 ( .A1(n6026), .A2(net58676), .ZN(n6028) );
  NOR2_X1 U3801 ( .A1(n6025), .A2(n6024), .ZN(n6026) );
  INV_X16 U3802 ( .A(net63573), .ZN(net63571) );
  NAND3_X1 U3803 ( .A1(net58932), .A2(u4_fract_out_pl1_52_), .A3(net58951), 
        .ZN(n4644) );
  NOR2_X1 U3804 ( .A1(n4406), .A2(n6982), .ZN(n6988) );
  NOR2_X2 U3805 ( .A1(n6924), .A2(n6952), .ZN(n6940) );
  NOR2_X2 U3806 ( .A1(fracta_mul[9]), .A2(fracta_mul[8]), .ZN(n6862) );
  NOR2_X1 U3807 ( .A1(net57241), .A2(n5716), .ZN(n5584) );
  NAND3_X2 U3808 ( .A1(n5126), .A2(n5125), .A3(n5124), .ZN(fract_denorm[98])
         );
  NAND3_X2 U3809 ( .A1(n5546), .A2(net59799), .A3(n5545), .ZN(
        u4_shift_right[7]) );
  OAI21_X1 U3810 ( .B1(div_opa_ldz_r2[1]), .B2(n5497), .A(n5508), .ZN(net59721) );
  NOR2_X1 U3811 ( .A1(n4852), .A2(n5512), .ZN(n5497) );
  NAND3_X1 U3812 ( .A1(n4515), .A2(net60276), .A3(fract_denorm[76]), .ZN(
        net60275) );
  OAI21_X2 U3813 ( .B1(net60050), .B2(net60273), .A(n5341), .ZN(n5437) );
  NOR3_X1 U3814 ( .A1(n5337), .A2(fract_denorm[75]), .A3(fract_denorm[81]), 
        .ZN(net60291) );
  NOR3_X1 U3815 ( .A1(fract_denorm[91]), .A2(fract_denorm[92]), .A3(net60306), 
        .ZN(n5335) );
  NAND3_X2 U3816 ( .A1(n5375), .A2(n5374), .A3(n5373), .ZN(net33648) );
  NAND3_X2 U3817 ( .A1(n5515), .A2(n5514), .A3(n5513), .ZN(net33546) );
  NOR2_X1 U3818 ( .A1(net57241), .A2(net59435), .ZN(n5535) );
  NAND3_X1 U3819 ( .A1(opb_inf), .A2(opa_inf), .A3(sign_exe_r), .ZN(net58820)
         );
  NOR3_X2 U3820 ( .A1(n6090), .A2(n6089), .A3(n6088), .ZN(n6091) );
  INV_X16 U3821 ( .A(net63569), .ZN(net63565) );
  NOR2_X1 U3822 ( .A1(net58550), .A2(net58636), .ZN(net58634) );
  INV_X4 U3823 ( .A(net58657), .ZN(net58632) );
  NOR2_X1 U3824 ( .A1(exp_ovf_r_0_), .A2(net63287), .ZN(net59198) );
  INV_X4 U3825 ( .A(n4764), .ZN(n7067) );
  INV_X4 U3826 ( .A(u1_fractb_lt_fracta), .ZN(n4906) );
  NOR2_X2 U3827 ( .A1(opb_r[61]), .A2(n4391), .ZN(n6730) );
  NAND3_X1 U3828 ( .A1(fracta_mul[25]), .A2(n4955), .A3(n4422), .ZN(n5069) );
  NOR3_X1 U3829 ( .A1(fracta_mul[9]), .A2(fracta_mul[8]), .A3(n5068), .ZN(
        n4986) );
  NOR2_X1 U3830 ( .A1(n5068), .A2(n6837), .ZN(n4945) );
  NOR2_X2 U3831 ( .A1(n4946), .A2(n5048), .ZN(n4947) );
  AOI21_X1 U3832 ( .B1(fracta_mul[33]), .B2(n4314), .A(fracta_mul[35]), .ZN(
        n4946) );
  NOR2_X2 U3833 ( .A1(n5989), .A2(n7205), .ZN(n5990) );
  NOR2_X2 U3834 ( .A1(net66871), .A2(n5676), .ZN(n5678) );
  OAI21_X1 U3835 ( .B1(net66871), .B2(n5501), .A(net66875), .ZN(n5499) );
  OAI21_X1 U3836 ( .B1(u2_exp_tmp4_9_), .B2(n6290), .A(n6289), .ZN(n6291) );
  NOR2_X1 U3837 ( .A1(n6341), .A2(n6393), .ZN(n6342) );
  NOR2_X2 U3838 ( .A1(n6340), .A2(n6402), .ZN(n6343) );
  NOR2_X1 U3839 ( .A1(n6358), .A2(n6393), .ZN(n6359) );
  NOR2_X1 U3840 ( .A1(n6370), .A2(n6393), .ZN(n6371) );
  INV_X8 U3841 ( .A(n4354), .ZN(n4845) );
  NOR2_X1 U3842 ( .A1(n6332), .A2(n6409), .ZN(n6333) );
  INV_X8 U3843 ( .A(n4474), .ZN(n4844) );
  NOR2_X2 U3844 ( .A1(net66839), .A2(net58932), .ZN(n5683) );
  INV_X4 U3845 ( .A(net58772), .ZN(net58428) );
  NOR2_X2 U3846 ( .A1(n5880), .A2(net58506), .ZN(n5881) );
  INV_X16 U3847 ( .A(n4903), .ZN(n4901) );
  NAND2_X2 U3848 ( .A1(n6477), .A2(n4298), .ZN(n8510) );
  NOR2_X2 U3849 ( .A1(fpu_op_r2[1]), .A2(fpu_op_r2[2]), .ZN(n4254) );
  NOR2_X2 U3850 ( .A1(opa_r1[57]), .A2(opa_r1[58]), .ZN(n6475) );
  NOR2_X2 U3851 ( .A1(n4252), .A2(opa_r1[52]), .ZN(n6474) );
  NOR2_X2 U3852 ( .A1(opa_r1[53]), .A2(opa_r1[54]), .ZN(n6473) );
  NOR3_X1 U3853 ( .A1(n4398), .A2(n6738), .A3(n6737), .ZN(n6748) );
  NOR2_X2 U3854 ( .A1(n6746), .A2(n6745), .ZN(n6747) );
  NOR3_X2 U3855 ( .A1(n6455), .A2(n6454), .A3(n6453), .ZN(n7198) );
  NAND3_X1 U3856 ( .A1(n4439), .A2(n6452), .A3(n6451), .ZN(n6453) );
  NAND3_X1 U3857 ( .A1(n6445), .A2(n6444), .A3(n6443), .ZN(n6455) );
  NOR2_X1 U3858 ( .A1(n4392), .A2(n4331), .ZN(n7142) );
  NOR2_X1 U3859 ( .A1(n7141), .A2(n4390), .ZN(n7144) );
  NOR2_X1 U3860 ( .A1(n3081), .A2(n4330), .ZN(n7143) );
  NOR2_X1 U3861 ( .A1(n7146), .A2(n7145), .ZN(n7152) );
  NOR2_X1 U3862 ( .A1(n7149), .A2(n7148), .ZN(n7150) );
  NOR2_X1 U3863 ( .A1(n3078), .A2(n7147), .ZN(n7151) );
  NOR3_X2 U3864 ( .A1(n6458), .A2(n4472), .A3(n6457), .ZN(n6459) );
  NOR2_X1 U3865 ( .A1(fracta_mul[50]), .A2(n4301), .ZN(n5071) );
  AOI21_X2 U3866 ( .B1(n4991), .B2(n4990), .A(n4989), .ZN(n4993) );
  NOR2_X1 U3867 ( .A1(n4988), .A2(n4310), .ZN(n4989) );
  NOR2_X1 U3868 ( .A1(n5068), .A2(n4343), .ZN(n4991) );
  NAND3_X1 U3869 ( .A1(n5050), .A2(n5049), .A3(n4311), .ZN(n5051) );
  OAI21_X1 U3870 ( .B1(fracta_mul[17]), .B2(fracta_mul[18]), .A(n4438), .ZN(
        n5044) );
  NAND3_X1 U3871 ( .A1(fracta_mul[10]), .A2(n5038), .A3(n4312), .ZN(n5045) );
  AOI21_X1 U3872 ( .B1(n5019), .B2(n5018), .A(n5017), .ZN(n5028) );
  OAI21_X1 U3873 ( .B1(n5022), .B2(fracta_mul[15]), .A(n5021), .ZN(n5027) );
  NAND3_X2 U3874 ( .A1(n5009), .A2(n5008), .A3(n5007), .ZN(n5015) );
  NAND3_X1 U3875 ( .A1(fracta_mul[16]), .A2(n4341), .A3(n4464), .ZN(n5009) );
  AOI21_X1 U3876 ( .B1(fracta_mul[14]), .B2(n4934), .A(n6439), .ZN(n5007) );
  NOR3_X1 U3877 ( .A1(n5048), .A2(fracta_mul[35]), .A3(n5049), .ZN(n5005) );
  NOR3_X2 U3878 ( .A1(fracta_mul[5]), .A2(n4942), .A3(n5068), .ZN(n4962) );
  OAI21_X1 U3879 ( .B1(n3203), .B2(n5048), .A(n4960), .ZN(n4963) );
  NOR3_X1 U3880 ( .A1(fracta_mul[32]), .A2(fracta_mul[34]), .A3(fracta_mul[28]), .ZN(n3203) );
  NAND3_X1 U3881 ( .A1(fracta_mul[36]), .A2(n4959), .A3(n4310), .ZN(n4960) );
  NOR2_X2 U3882 ( .A1(n5998), .A2(n7202), .ZN(n5999) );
  AOI21_X1 U3883 ( .B1(n4723), .B2(net58733), .A(net58728), .ZN(n4721) );
  NOR2_X2 U3884 ( .A1(net58743), .A2(n5986), .ZN(n5988) );
  NOR2_X1 U3885 ( .A1(n5989), .A2(n5970), .ZN(n5972) );
  NOR2_X1 U3886 ( .A1(n4505), .A2(n7191), .ZN(n7192) );
  NOR2_X1 U3887 ( .A1(net57240), .A2(net57241), .ZN(n7194) );
  NOR2_X1 U3888 ( .A1(n7180), .A2(n4843), .ZN(n7181) );
  NOR2_X1 U3889 ( .A1(net57241), .A2(n7183), .ZN(n7184) );
  AOI21_X1 U3890 ( .B1(u4_exp_out1_1_), .B2(net59258), .A(net59296), .ZN(
        net59701) );
  OAI21_X2 U3891 ( .B1(net58789), .B2(net58506), .A(net58790), .ZN(N911) );
  AOI21_X2 U3892 ( .B1(n6048), .B2(net58613), .A(n6047), .ZN(n6050) );
  OAI21_X2 U3893 ( .B1(opa_00), .B2(n6106), .A(n6105), .ZN(n6107) );
  NOR2_X2 U3894 ( .A1(net63529), .A2(n6116), .ZN(N799) );
  NOR2_X2 U3895 ( .A1(net63529), .A2(n6117), .ZN(N800) );
  NOR2_X1 U3896 ( .A1(net63529), .A2(net58494), .ZN(N803) );
  NAND3_X2 U3897 ( .A1(exp_mul[6]), .A2(exp_mul[5]), .A3(exp_mul[7]), .ZN(
        n3294) );
  NOR3_X2 U3898 ( .A1(n4358), .A2(n4319), .A3(n4490), .ZN(n3295) );
  NOR2_X2 U3899 ( .A1(n6410), .A2(n6711), .ZN(u2_exp_ovf_d_0_) );
  NOR2_X2 U3900 ( .A1(n6463), .A2(n6465), .ZN(u2_underflow_d[2]) );
  NOR2_X1 U3901 ( .A1(n6765), .A2(n6763), .ZN(u1_N54) );
  NOR2_X1 U3902 ( .A1(n6765), .A2(n6764), .ZN(u1_N53) );
  NOR2_X1 U3903 ( .A1(n6766), .A2(n6765), .ZN(u1_N52) );
  OAI21_X2 U3904 ( .B1(n3060), .B2(n4498), .A(n3061), .ZN(u1_N229) );
  OAI21_X2 U3905 ( .B1(n3062), .B2(n4494), .A(u1_signa_r), .ZN(n3061) );
  NOR3_X2 U3906 ( .A1(n3063), .A2(u1_fracta_lt_fractb), .A3(
        u1_fracta_eq_fractb), .ZN(n3062) );
  NOR2_X1 U3907 ( .A1(net63083), .A2(n3341), .ZN(N904) );
  NOR2_X2 U3908 ( .A1(n3071), .A2(n3070), .ZN(u0_N6) );
  NOR2_X1 U3909 ( .A1(fracta_mul[51]), .A2(n7198), .ZN(u0_N4) );
  NOR3_X2 U3910 ( .A1(n4495), .A2(opa_nan), .A3(n3296), .ZN(N912) );
  NOR2_X2 U3911 ( .A1(n7197), .A2(n7154), .ZN(u0_N10) );
  NOR2_X2 U3912 ( .A1(n4346), .A2(n3074), .ZN(u0_N11) );
  INV_X4 U3913 ( .A(n4399), .ZN(n4853) );
  NAND3_X2 U3914 ( .A1(n5032), .A2(n5031), .A3(n5030), .ZN(div_opa_ldz_d[2])
         );
  AOI21_X1 U3915 ( .B1(n5005), .B2(fracta_mul[32]), .A(n5004), .ZN(n5032) );
  AOI211_X1 U3916 ( .C1(n5016), .C2(n5015), .A(n5014), .B(n4463), .ZN(n5031)
         );
  NOR3_X1 U3917 ( .A1(n5060), .A2(n5029), .A3(n5073), .ZN(n5030) );
  AOI211_X1 U3918 ( .C1(n4978), .C2(n4977), .A(n4976), .B(n4975), .ZN(n5002)
         );
  NOR3_X1 U3919 ( .A1(n4983), .A2(n4443), .A3(n5060), .ZN(n5001) );
  NOR2_X1 U3920 ( .A1(n5024), .A2(n5065), .ZN(n5000) );
  INV_X16 U3921 ( .A(net63351), .ZN(net63339) );
  INV_X16 U3922 ( .A(net63351), .ZN(net63343) );
  NOR2_X2 U3923 ( .A1(n7158), .A2(n7157), .ZN(n2476) );
  NOR2_X1 U3924 ( .A1(net57281), .A2(net57241), .ZN(n7157) );
  NOR2_X2 U3925 ( .A1(net57281), .A2(n7191), .ZN(n7158) );
  AOI21_X2 U3926 ( .B1(n5976), .B2(n5975), .A(n5974), .ZN(n5978) );
  AOI21_X1 U3927 ( .B1(n7163), .B2(n7169), .A(n7178), .ZN(n2421) );
  NOR2_X1 U3928 ( .A1(net57276), .A2(n7159), .ZN(n7163) );
  NOR2_X1 U3929 ( .A1(u4_fi_ldz_5_), .A2(n7166), .ZN(n7164) );
  NOR2_X1 U3930 ( .A1(n5998), .A2(n5994), .ZN(n5996) );
  AOI21_X1 U3931 ( .B1(net57252), .B2(n7176), .A(n7178), .ZN(n2412) );
  AOI21_X1 U3932 ( .B1(net57252), .B2(u4_fi_ldz_mi22[2]), .A(n7178), .ZN(n2409) );
  NOR3_X2 U3933 ( .A1(n7194), .A2(n7193), .A3(n7192), .ZN(net57232) );
  NOR2_X1 U3934 ( .A1(n7190), .A2(n4843), .ZN(n7193) );
  NOR2_X2 U3935 ( .A1(n7185), .A2(n7184), .ZN(n7186) );
  NAND3_X1 U3936 ( .A1(net59260), .A2(net59261), .A3(fract_denorm[104]), .ZN(
        n4564) );
  NOR3_X2 U3937 ( .A1(u4_N5938), .A2(u4_N5940), .A3(u4_N5939), .ZN(n3930) );
  NOR3_X2 U3938 ( .A1(u4_N5935), .A2(u4_N5937), .A3(u4_N5936), .ZN(n3929) );
  NOR3_X2 U3939 ( .A1(u4_N5932), .A2(u4_N5934), .A3(u4_N5933), .ZN(n3928) );
  NOR3_X2 U3940 ( .A1(u4_N5945), .A2(u4_N5947), .A3(u4_N5946), .ZN(n3932) );
  NOR3_X2 U3941 ( .A1(u4_N5952), .A2(u4_N5954), .A3(u4_N5953), .ZN(n3934) );
  NOR3_X2 U3942 ( .A1(u4_N5912), .A2(u4_N5914), .A3(u4_N5913), .ZN(n3922) );
  NOR3_X2 U3943 ( .A1(u4_N5909), .A2(u4_N5911), .A3(u4_N5910), .ZN(n3921) );
  NOR3_X2 U3944 ( .A1(u4_N5906), .A2(u4_N5908), .A3(u4_N5907), .ZN(n3920) );
  NOR3_X2 U3945 ( .A1(u4_N5922), .A2(u4_N5924), .A3(u4_N5923), .ZN(n3925) );
  NOR3_X2 U3946 ( .A1(u4_N5919), .A2(u4_N5921), .A3(u4_N5920), .ZN(n3924) );
  NOR3_X2 U3947 ( .A1(u4_N5925), .A2(u4_N5927), .A3(u4_N5926), .ZN(n3926) );
  INV_X4 U3948 ( .A(n6597), .ZN(n4862) );
  AND2_X4 U3949 ( .A1(n8510), .A2(n6578), .ZN(n4292) );
  INV_X1 U3950 ( .A(n7208), .ZN(n4898) );
  INV_X2 U3951 ( .A(u2_N157), .ZN(n7208) );
  OR2_X4 U3952 ( .A1(net60696), .A2(n4519), .ZN(n4293) );
  INV_X4 U3953 ( .A(net59081), .ZN(net59154) );
  XOR2_X2 U3954 ( .A(n5645), .B(n4328), .Z(n4295) );
  INV_X4 U3955 ( .A(n7208), .ZN(n4903) );
  OR2_X4 U3956 ( .A1(net60696), .A2(n4519), .ZN(n4305) );
  NAND2_X2 U3957 ( .A1(n4804), .A2(n4736), .ZN(n4309) );
  INV_X8 U3958 ( .A(n4893), .ZN(n4892) );
  INV_X16 U3959 ( .A(n4897), .ZN(n4879) );
  INV_X16 U3960 ( .A(n4897), .ZN(n4880) );
  AND2_X4 U3961 ( .A1(n4300), .A2(n4290), .ZN(n4316) );
  XOR2_X2 U3962 ( .A(n4854), .B(n6337), .Z(n4318) );
  INV_X4 U3963 ( .A(n6480), .ZN(n4859) );
  INV_X4 U3964 ( .A(n4898), .ZN(n4900) );
  INV_X4 U3965 ( .A(n4903), .ZN(n4899) );
  INV_X1 U3966 ( .A(n4903), .ZN(n4902) );
  NAND2_X1 U3967 ( .A1(net58925), .A2(net58926), .ZN(net58420) );
  AND3_X4 U3968 ( .A1(net60072), .A2(net60073), .A3(net60008), .ZN(n4320) );
  INV_X4 U3969 ( .A(n4305), .ZN(net66912) );
  INV_X4 U3970 ( .A(n4305), .ZN(net66914) );
  INV_X4 U3971 ( .A(n4305), .ZN(net66910) );
  AND2_X4 U3972 ( .A1(net60085), .A2(net60317), .ZN(n4321) );
  AND2_X4 U3973 ( .A1(net60695), .A2(n4376), .ZN(n4322) );
  AND4_X2 U3974 ( .A1(fract_denorm[61]), .A2(net60142), .A3(net60237), .A4(
        net60106), .ZN(n4323) );
  INV_X4 U3975 ( .A(net63515), .ZN(net63513) );
  XOR2_X1 U3976 ( .A(div_opa_ldz_r2[1]), .B(n4852), .Z(n4325) );
  INV_X16 U3977 ( .A(net63351), .ZN(net63349) );
  INV_X16 U3978 ( .A(net44995), .ZN(net63351) );
  XOR2_X2 U3979 ( .A(n5640), .B(n4327), .Z(n4329) );
  AND2_X4 U3980 ( .A1(n7139), .A2(n7138), .ZN(n4333) );
  AND2_X2 U3981 ( .A1(n4473), .A2(n6999), .ZN(n4346) );
  OR3_X1 U3982 ( .A1(u6_N18), .A2(u6_N1), .A3(u6_N19), .ZN(n4350) );
  INV_X4 U3983 ( .A(net58420), .ZN(net63523) );
  OR2_X4 U3984 ( .A1(u2_exp_ovf_d_1_), .A2(u1_N46), .ZN(n4354) );
  INV_X8 U3985 ( .A(n4895), .ZN(n4886) );
  OR2_X4 U3986 ( .A1(net63515), .A2(net58432), .ZN(n4357) );
  INV_X4 U3987 ( .A(n4292), .ZN(n4866) );
  INV_X4 U3988 ( .A(n4304), .ZN(n4917) );
  INV_X4 U3989 ( .A(n4304), .ZN(n4916) );
  AND2_X2 U3990 ( .A1(net58546), .A2(net58781), .ZN(n4367) );
  AND3_X4 U3991 ( .A1(n4624), .A2(n4625), .A3(n4626), .ZN(n4368) );
  AND2_X2 U3992 ( .A1(net59099), .A2(net59161), .ZN(n4369) );
  AND3_X2 U3993 ( .A1(n4520), .A2(net60196), .A3(fract_denorm[58]), .ZN(n4370)
         );
  OR2_X4 U3994 ( .A1(u4_fi_ldz_3_), .A2(u4_fi_ldz_4_), .ZN(n4371) );
  AND3_X4 U3995 ( .A1(n5416), .A2(net60044), .A3(fract_denorm[83]), .ZN(n4372)
         );
  AND3_X4 U3996 ( .A1(net60026), .A2(net59953), .A3(net33642), .ZN(n4373) );
  OR2_X1 U3997 ( .A1(net60011), .A2(n4521), .ZN(n4374) );
  INV_X16 U3998 ( .A(net63573), .ZN(net63569) );
  INV_X16 U3999 ( .A(net63575), .ZN(net63573) );
  INV_X8 U4000 ( .A(net63569), .ZN(net63567) );
  INV_X16 U4001 ( .A(net63571), .ZN(net63559) );
  NAND3_X2 U4002 ( .A1(n4689), .A2(n4688), .A3(n4690), .ZN(net60201) );
  INV_X2 U4003 ( .A(net60201), .ZN(net60316) );
  INV_X1 U4004 ( .A(n4663), .ZN(n4664) );
  NAND3_X2 U4005 ( .A1(net60062), .A2(n4662), .A3(n4665), .ZN(n4663) );
  INV_X8 U4006 ( .A(n4376), .ZN(net63093) );
  INV_X16 U4007 ( .A(fract_denorm_105_), .ZN(net63221) );
  NAND2_X2 U4008 ( .A1(net60219), .A2(net60304), .ZN(net60094) );
  INV_X2 U4009 ( .A(net60094), .ZN(net60092) );
  INV_X8 U4010 ( .A(n4378), .ZN(n4851) );
  AND2_X4 U4011 ( .A1(net59551), .A2(n5534), .ZN(n4380) );
  INV_X2 U4012 ( .A(net59087), .ZN(net59122) );
  AND3_X4 U4013 ( .A1(net60329), .A2(net60167), .A3(net60196), .ZN(n4382) );
  XOR2_X2 U4014 ( .A(n5490), .B(n4327), .Z(n4385) );
  AND2_X4 U4015 ( .A1(u1_adj_op_out_sft_2_), .A2(n7138), .ZN(n4397) );
  AND2_X2 U4016 ( .A1(opb_r[55]), .A2(n4390), .ZN(n4398) );
  OR2_X2 U4017 ( .A1(u4_exp_in_pl1_10_), .A2(u4_exp_in_pl1_9_), .ZN(n4400) );
  AND2_X2 U4018 ( .A1(net59717), .A2(n5577), .ZN(n4402) );
  OR2_X2 U4019 ( .A1(u1_exp_diff2[7]), .A2(u1_exp_diff2[6]), .ZN(n4403) );
  AND2_X4 U4020 ( .A1(rmode_r3[0]), .A2(rmode_r3[1]), .ZN(n4405) );
  AND3_X2 U4021 ( .A1(n6922), .A2(n6914), .A3(n6955), .ZN(n4406) );
  AND3_X2 U4022 ( .A1(n6923), .A2(n6909), .A3(n6953), .ZN(n4407) );
  INV_X4 U4023 ( .A(opb_r[56]), .ZN(n4835) );
  AND3_X4 U4024 ( .A1(fracta_mul[40]), .A2(n4996), .A3(n4313), .ZN(n4443) );
  INV_X4 U4025 ( .A(n4731), .ZN(n7020) );
  NAND3_X2 U4026 ( .A1(u1_N46), .A2(n6409), .A3(u2_exp_ovf_d_1_), .ZN(n6402)
         );
  AND2_X2 U4027 ( .A1(fracta_mul[46]), .A2(n5019), .ZN(n4463) );
  NAND3_X1 U4028 ( .A1(n4936), .A2(n4428), .A3(n6862), .ZN(n4979) );
  NOR2_X1 U4029 ( .A1(fracta_mul[18]), .A2(fracta_mul[19]), .ZN(n4464) );
  INV_X1 U4030 ( .A(n5067), .ZN(n5038) );
  OR3_X1 U4031 ( .A1(u6_N12), .A2(u6_N14), .A3(u6_N13), .ZN(n4465) );
  OR3_X1 U4032 ( .A1(fracta_mul[46]), .A2(fracta_mul[48]), .A3(fracta_mul[47]), 
        .ZN(n4466) );
  AND3_X4 U4033 ( .A1(n7220), .A2(n7219), .A3(n7218), .ZN(n4467) );
  OR2_X4 U4034 ( .A1(exp_ovf_r_0_), .A2(net58932), .ZN(n4468) );
  OR2_X4 U4035 ( .A1(fracta_mul[6]), .A2(fracta_mul[7]), .ZN(n4469) );
  AND2_X2 U4036 ( .A1(net58812), .A2(net58645), .ZN(n4470) );
  AND3_X4 U4037 ( .A1(net63293), .A2(opa_inf), .A3(n4429), .ZN(n4471) );
  OR2_X4 U4038 ( .A1(u6_N10), .A2(u6_N0), .ZN(n4472) );
  AND3_X4 U4039 ( .A1(n6461), .A2(n6460), .A3(n6459), .ZN(n4473) );
  OR3_X4 U4040 ( .A1(n6468), .A2(n6406), .A3(n6409), .ZN(n4474) );
  OR2_X4 U4041 ( .A1(n6441), .A2(n4439), .ZN(n4475) );
  OR2_X1 U4042 ( .A1(n6442), .A2(n4423), .ZN(n4476) );
  AND2_X2 U4043 ( .A1(n6385), .A2(n6409), .ZN(n4477) );
  INV_X1 U4044 ( .A(n6409), .ZN(n6272) );
  OR2_X4 U4045 ( .A1(opb_00), .A2(opb_inf), .ZN(n4485) );
  OR2_X4 U4046 ( .A1(net58650), .A2(net59053), .ZN(n4486) );
  AND3_X4 U4047 ( .A1(n6470), .A2(n6468), .A3(n6469), .ZN(n4487) );
  INV_X4 U4048 ( .A(n6480), .ZN(n4861) );
  INV_X4 U4049 ( .A(n6480), .ZN(n4860) );
  INV_X4 U4050 ( .A(n6480), .ZN(n4858) );
  OR2_X1 U4051 ( .A1(net66835), .A2(net58550), .ZN(n4488) );
  INV_X4 U4052 ( .A(n4866), .ZN(n4864) );
  INV_X4 U4053 ( .A(n4866), .ZN(n4863) );
  INV_X4 U4054 ( .A(n4866), .ZN(n4865) );
  OR2_X4 U4055 ( .A1(n5048), .A2(n4476), .ZN(n4489) );
  INV_X4 U4056 ( .A(n6481), .ZN(n4856) );
  INV_X4 U4057 ( .A(n6481), .ZN(n4857) );
  INV_X4 U4058 ( .A(n6481), .ZN(n4855) );
  INV_X4 U4059 ( .A(net58420), .ZN(net63537) );
  INV_X4 U4060 ( .A(net58420), .ZN(net63529) );
  INV_X4 U4061 ( .A(net58420), .ZN(net63527) );
  INV_X16 U4062 ( .A(net58443), .ZN(net63521) );
  INV_X16 U4063 ( .A(net63521), .ZN(net63515) );
  INV_X4 U4064 ( .A(n4304), .ZN(n4918) );
  INV_X2 U4065 ( .A(net60289), .ZN(net60295) );
  AOI21_X2 U4066 ( .B1(net59958), .B2(net59959), .A(net63217), .ZN(net59957)
         );
  NOR2_X1 U4067 ( .A1(n4366), .A2(net58437), .ZN(net58537) );
  NAND3_X1 U4068 ( .A1(net63083), .A2(n4288), .A3(n4366), .ZN(net58926) );
  NAND3_X1 U4069 ( .A1(n4534), .A2(net58662), .A3(n6033), .ZN(n6034) );
  NOR2_X1 U4070 ( .A1(n4534), .A2(n4488), .ZN(n6025) );
  NAND4_X2 U4071 ( .A1(net33564), .A2(n4694), .A3(n4695), .A4(n4509), .ZN(
        net60137) );
  INV_X4 U4072 ( .A(n4508), .ZN(n4509) );
  OAI21_X2 U4073 ( .B1(net58973), .B2(net58970), .A(net58971), .ZN(net58772)
         );
  INV_X4 U4074 ( .A(net58974), .ZN(net58990) );
  NAND2_X1 U4075 ( .A1(net60022), .A2(net60289), .ZN(net60288) );
  NAND2_X1 U4076 ( .A1(n5410), .A2(net60022), .ZN(n5411) );
  NAND2_X1 U4077 ( .A1(net60022), .A2(net60005), .ZN(net59952) );
  AND2_X2 U4078 ( .A1(net60022), .A2(net60191), .ZN(n4515) );
  NAND2_X1 U4079 ( .A1(net60295), .A2(net60022), .ZN(n5338) );
  NAND3_X1 U4080 ( .A1(net58768), .A2(net58769), .A3(n4709), .ZN(net58653) );
  NAND3_X2 U4081 ( .A1(net59191), .A2(net59234), .A3(net59235), .ZN(net59194)
         );
  OAI21_X1 U4082 ( .B1(net59191), .B2(net59083), .A(net59146), .ZN(net59184)
         );
  OAI21_X1 U4083 ( .B1(net59230), .B2(net59101), .A(net59099), .ZN(net59200)
         );
  AOI22_X2 U4084 ( .A1(net59670), .A2(n5623), .B1(n4846), .B2(n5629), .ZN(
        n5626) );
  INV_X1 U4085 ( .A(net60097), .ZN(n4508) );
  INV_X4 U4086 ( .A(n4510), .ZN(n4511) );
  INV_X8 U4087 ( .A(net59966), .ZN(net60097) );
  INV_X8 U4088 ( .A(net60287), .ZN(net60051) );
  NAND2_X1 U4089 ( .A1(n4509), .A2(net33562), .ZN(n5382) );
  NAND3_X1 U4090 ( .A1(net60187), .A2(net33550), .A3(net60072), .ZN(net60279)
         );
  NAND2_X1 U4091 ( .A1(net60072), .A2(net60290), .ZN(net60273) );
  AOI21_X1 U4092 ( .B1(n4511), .B2(net60186), .A(n5330), .ZN(n5334) );
  NAND3_X1 U4093 ( .A1(n4511), .A2(net59336), .A3(n4562), .ZN(net59995) );
  NAND3_X1 U4094 ( .A1(net33577), .A2(net60145), .A3(n4511), .ZN(n5379) );
  AOI22_X1 U4095 ( .A1(n4592), .A2(net59697), .B1(n4511), .B2(net33575), .ZN(
        net60100) );
  NAND3_X1 U4096 ( .A1(n4511), .A2(net60084), .A3(n8516), .ZN(n5405) );
  NAND3_X1 U4097 ( .A1(net60051), .A2(n8517), .A3(n5396), .ZN(n5401) );
  NAND2_X1 U4098 ( .A1(net60316), .A2(n4522), .ZN(n4524) );
  AOI21_X1 U4099 ( .B1(net60085), .B2(net60314), .A(n5331), .ZN(n5332) );
  NAND3_X1 U4100 ( .A1(net60085), .A2(net60086), .A3(net33583), .ZN(net60078)
         );
  NAND3_X1 U4101 ( .A1(net60085), .A2(n8515), .A3(n5397), .ZN(n5400) );
  NOR3_X2 U4102 ( .A1(net59519), .A2(u4_fract_out_0_), .A3(u4_fract_out_12_), 
        .ZN(n4577) );
  NAND3_X1 U4103 ( .A1(n2523), .A2(n3702), .A3(n3699), .ZN(net59519) );
  NOR2_X2 U4104 ( .A1(n5713), .A2(n5712), .ZN(net59517) );
  NAND3_X1 U4105 ( .A1(n3626), .A2(n2526), .A3(n3720), .ZN(n5712) );
  NAND3_X1 U4106 ( .A1(n3629), .A2(n2524), .A3(n2522), .ZN(n5713) );
  NOR4_X1 U4107 ( .A1(net59592), .A2(net59593), .A3(net58780), .A4(net59347), 
        .ZN(net59591) );
  NOR2_X1 U4108 ( .A1(u4_exp_in_mi1_11_), .A2(net58652), .ZN(net58648) );
  NOR2_X2 U4109 ( .A1(net59260), .A2(net58652), .ZN(net59592) );
  INV_X8 U4110 ( .A(net63589), .ZN(net63583) );
  INV_X16 U4111 ( .A(net63589), .ZN(net63585) );
  NOR2_X2 U4112 ( .A1(n4575), .A2(n4576), .ZN(n4574) );
  NAND3_X1 U4113 ( .A1(n3636), .A2(n2527), .A3(n2525), .ZN(n4575) );
  NAND3_X1 U4114 ( .A1(n4512), .A2(net60193), .A3(fract_denorm[66]), .ZN(
        net60322) );
  NAND3_X2 U4115 ( .A1(n4512), .A2(net60194), .A3(net60193), .ZN(net59946) );
  NOR2_X4 U4116 ( .A1(net60352), .A2(n4663), .ZN(n4512) );
  MUX2_X2 U4117 ( .A(net58821), .B(nan_sign_d), .S(n4513), .Z(net58816) );
  OR2_X4 U4118 ( .A1(ind_d), .A2(net58506), .ZN(n4513) );
  INV_X4 U4119 ( .A(net60352), .ZN(net60004) );
  NAND2_X1 U4120 ( .A1(net60004), .A2(n4664), .ZN(n4517) );
  NAND3_X1 U4121 ( .A1(n4514), .A2(net59990), .A3(net60047), .ZN(net60028) );
  NOR3_X2 U4122 ( .A1(n4521), .A2(net33554), .A3(n8524), .ZN(n5460) );
  NAND2_X4 U4123 ( .A1(n4276), .A2(net59339), .ZN(n4521) );
  NAND3_X2 U4124 ( .A1(n4320), .A2(n8518), .A3(n5409), .ZN(net60055) );
  AOI211_X2 U4125 ( .C1(net59922), .C2(net60058), .A(n5415), .B(net60060), 
        .ZN(net60057) );
  NOR2_X4 U4126 ( .A1(n4275), .A2(net60159), .ZN(n4514) );
  INV_X2 U4127 ( .A(net33547), .ZN(net59339) );
  NOR4_X1 U4128 ( .A1(n6017), .A2(n6016), .A3(u4_ldz_all_6_), .A4(n6015), .ZN(
        n6022) );
  OAI21_X1 U4129 ( .B1(net58634), .B2(exp_ovf_r_0_), .A(net58635), .ZN(
        net58630) );
  NAND4_X2 U4130 ( .A1(net58950), .A2(net58635), .A3(net63289), .A4(net58960), 
        .ZN(net58959) );
  AOI22_X4 U4131 ( .A1(u4_N5970), .A2(net63319), .B1(u4_N6078), .B2(net63335), 
        .ZN(n2541) );
  NAND3_X2 U4132 ( .A1(n2540), .A2(n2541), .A3(n3691), .ZN(n5708) );
  NAND3_X2 U4133 ( .A1(n3689), .A2(n3727), .A3(n3687), .ZN(n5709) );
  NAND3_X2 U4134 ( .A1(n5626), .A2(n5625), .A3(n5624), .ZN(u4_shift_left[8])
         );
  INV_X1 U4135 ( .A(net59946), .ZN(net60236) );
  OAI21_X2 U4136 ( .B1(net60286), .B2(n4510), .A(net60288), .ZN(net60285) );
  AOI21_X1 U4137 ( .B1(net58776), .B2(net58777), .A(net58778), .ZN(net58775)
         );
  NAND2_X1 U4138 ( .A1(net59351), .A2(net59352), .ZN(net59350) );
  INV_X8 U4139 ( .A(n2530), .ZN(u4_fract_out_33_) );
  AOI22_X4 U4140 ( .A1(u4_N5993), .A2(net63325), .B1(u4_N6101), .B2(net63343), 
        .ZN(n2530) );
  NAND3_X2 U4141 ( .A1(n3641), .A2(n3644), .A3(n3638), .ZN(n4576) );
  INV_X8 U4142 ( .A(net59241), .ZN(net59231) );
  OAI21_X1 U4143 ( .B1(net58643), .B2(net59241), .A(n4644), .ZN(net59078) );
  NAND2_X1 U4144 ( .A1(net60085), .A2(net60344), .ZN(n4516) );
  INV_X1 U4145 ( .A(net59543), .ZN(net59670) );
  AOI222_X2 U4146 ( .A1(net59576), .A2(u4_ldz_dif_0_), .B1(net59600), .B2(
        div_opa_ldz_r2[0]), .C1(net59578), .C2(n4526), .ZN(net59573) );
  INV_X8 U4147 ( .A(n4528), .ZN(u4_shift_left[7]) );
  AOI211_X2 U4148 ( .C1(n4529), .C2(n4530), .A(n4531), .B(n5631), .ZN(n4528)
         );
  NAND3_X2 U4149 ( .A1(net59226), .A2(u4_exp_out_0_), .A3(net59225), .ZN(
        net58638) );
  NAND2_X1 U4150 ( .A1(net59578), .A2(u4_fi_ldz_5_), .ZN(n5642) );
  NOR2_X1 U4151 ( .A1(net60303), .A2(net60135), .ZN(net60300) );
  NOR2_X1 U4152 ( .A1(net59026), .A2(net58638), .ZN(net59020) );
  INV_X8 U4153 ( .A(n4554), .ZN(net59101) );
  INV_X8 U4154 ( .A(net58835), .ZN(net63575) );
  NOR3_X4 U4155 ( .A1(n5915), .A2(n5914), .A3(n5913), .ZN(n5919) );
  INV_X8 U4156 ( .A(net63589), .ZN(net63587) );
  OAI211_X1 U4157 ( .C1(net60291), .C2(net60282), .A(net60292), .B(net60293), 
        .ZN(net60283) );
  NOR2_X1 U4158 ( .A1(fract_denorm[103]), .A2(net59920), .ZN(net59914) );
  NOR4_X1 U4159 ( .A1(n5381), .A2(n5342), .A3(net60095), .A4(n5437), .ZN(n5343) );
  INV_X1 U4160 ( .A(net59961), .ZN(net60219) );
  NOR2_X1 U4161 ( .A1(net59961), .A2(net60168), .ZN(net60162) );
  INV_X2 U4162 ( .A(net59269), .ZN(n4518) );
  OAI221_X1 U4163 ( .B1(n5988), .B2(net58714), .C1(net58741), .C2(net58716), 
        .A(n5987), .ZN(net57265) );
  NAND2_X4 U4164 ( .A1(net59239), .A2(n4545), .ZN(n4544) );
  INV_X8 U4165 ( .A(net58638), .ZN(net58635) );
  NOR2_X2 U4166 ( .A1(net58997), .A2(net58638), .ZN(n4698) );
  NOR2_X2 U4167 ( .A1(net58638), .A2(n4462), .ZN(net59215) );
  INV_X8 U4168 ( .A(net59216), .ZN(net59192) );
  OAI21_X4 U4169 ( .B1(net58635), .B2(net59217), .A(net59218), .ZN(net59216)
         );
  OAI21_X2 U4170 ( .B1(net58969), .B2(net58970), .A(net58971), .ZN(net58968)
         );
  NAND2_X4 U4171 ( .A1(net58976), .A2(net58990), .ZN(net58970) );
  INV_X8 U4172 ( .A(net59447), .ZN(net59315) );
  OAI21_X4 U4173 ( .B1(net59448), .B2(net57285), .A(net59449), .ZN(net59447)
         );
  NOR3_X4 U4174 ( .A1(net58422), .A2(net58419), .A3(net58421), .ZN(n4712) );
  OAI221_X1 U4175 ( .B1(n6002), .B2(net58714), .C1(n4656), .C2(net58716), .A(
        n6001), .ZN(n6003) );
  OAI221_X1 U4176 ( .B1(n5972), .B2(net58714), .C1(net58762), .C2(net58716), 
        .A(n5971), .ZN(n7177) );
  AOI21_X1 U4177 ( .B1(fract_denorm[101]), .B2(n5434), .A(fract_denorm[103]), 
        .ZN(net60007) );
  INV_X8 U4178 ( .A(net60694), .ZN(net60468) );
  NAND2_X1 U4179 ( .A1(net60191), .A2(net60192), .ZN(net60190) );
  NOR4_X4 U4180 ( .A1(fract_denorm[84]), .A2(fract_denorm[83]), .A3(
        fract_denorm[82]), .A4(net60289), .ZN(net60191) );
  INV_X16 U4181 ( .A(net60697), .ZN(net59840) );
  NAND4_X4 U4182 ( .A1(net59994), .A2(net59995), .A3(net59996), .A4(net59997), 
        .ZN(net87917) );
  NOR2_X2 U4183 ( .A1(fract_denorm[104]), .A2(net63217), .ZN(n5469) );
  NAND4_X2 U4184 ( .A1(net60101), .A2(net60099), .A3(net60100), .A4(net60098), 
        .ZN(net60053) );
  NAND3_X1 U4185 ( .A1(net58646), .A2(n4519), .A3(n6034), .ZN(n6035) );
  NOR2_X1 U4186 ( .A1(opa_dn), .A2(n4519), .ZN(net59057) );
  NAND2_X1 U4187 ( .A1(opb_dn), .A2(net59703), .ZN(net58752) );
  NAND2_X1 U4188 ( .A1(n4519), .A2(n4389), .ZN(net59070) );
  NAND2_X1 U4189 ( .A1(opa_dn), .A2(opb_dn), .ZN(net59703) );
  NAND2_X4 U4190 ( .A1(net60695), .A2(n4519), .ZN(net60694) );
  INV_X1 U4191 ( .A(net60305), .ZN(net60304) );
  NAND2_X1 U4192 ( .A1(n5448), .A2(fract_denorm[100]), .ZN(net59959) );
  NOR3_X1 U4193 ( .A1(net59966), .A2(net33561), .A3(net59965), .ZN(n5446) );
  NOR2_X1 U4194 ( .A1(n4594), .A2(net59966), .ZN(n4593) );
  NOR2_X1 U4195 ( .A1(net60129), .A2(net59966), .ZN(n4682) );
  AOI22_X4 U4196 ( .A1(fract_out_q[46]), .A2(net63507), .B1(quo[45]), .B2(
        net66895), .ZN(n5130) );
  INV_X16 U4197 ( .A(net66894), .ZN(net66896) );
  INV_X8 U4198 ( .A(net59961), .ZN(net60111) );
  NOR2_X1 U4199 ( .A1(fract_denorm[97]), .A2(net59961), .ZN(net59956) );
  AND2_X2 U4200 ( .A1(net60316), .A2(net60348), .ZN(n4523) );
  INV_X4 U4201 ( .A(net60002), .ZN(n4522) );
  INV_X4 U4202 ( .A(n4524), .ZN(net59986) );
  INV_X1 U4203 ( .A(n4521), .ZN(net60220) );
  NAND4_X1 U4204 ( .A1(net60098), .A2(net60099), .A3(net60100), .A4(net60101), 
        .ZN(n4525) );
  NAND2_X4 U4205 ( .A1(net59344), .A2(net58779), .ZN(net59352) );
  NAND4_X1 U4206 ( .A1(net59994), .A2(net59995), .A3(net59996), .A4(net59997), 
        .ZN(n4526) );
  NAND4_X1 U4207 ( .A1(net59994), .A2(net59995), .A3(net59996), .A4(net59997), 
        .ZN(n4527) );
  NOR3_X1 U4208 ( .A1(n4525), .A2(net59984), .A3(net59974), .ZN(net60077) );
  NOR2_X4 U4209 ( .A1(n5437), .A2(net59984), .ZN(n5438) );
  NOR3_X4 U4210 ( .A1(net59478), .A2(net59479), .A3(net59480), .ZN(net59477)
         );
  NOR2_X2 U4211 ( .A1(net59540), .A2(net59541), .ZN(n5695) );
  AND2_X2 U4212 ( .A1(net58781), .A2(u4_f2i_shft_7_), .ZN(n4531) );
  NAND2_X4 U4213 ( .A1(net59310), .A2(u4_fract_out_pl1_52_), .ZN(net59241) );
  NAND3_X2 U4214 ( .A1(n5843), .A2(n5842), .A3(n5841), .ZN(net58983) );
  INV_X8 U4215 ( .A(net58776), .ZN(net59344) );
  NAND2_X4 U4216 ( .A1(net59421), .A2(net59222), .ZN(net58776) );
  INV_X1 U4217 ( .A(net58955), .ZN(net59224) );
  OAI21_X1 U4218 ( .B1(n4334), .B2(net58955), .A(net58956), .ZN(net58953) );
  AOI21_X1 U4219 ( .B1(n5694), .B2(net58636), .A(net59543), .ZN(n5696) );
  INV_X1 U4220 ( .A(net59543), .ZN(net59645) );
  NOR2_X1 U4221 ( .A1(net59543), .A2(n5653), .ZN(n5654) );
  NOR2_X1 U4222 ( .A1(net59543), .A2(n5662), .ZN(n5663) );
  INV_X1 U4223 ( .A(net59543), .ZN(net59576) );
  NOR2_X1 U4224 ( .A1(n5669), .A2(net59543), .ZN(n5671) );
  INV_X1 U4225 ( .A(net59543), .ZN(net59626) );
  INV_X1 U4226 ( .A(net59543), .ZN(net59632) );
  NOR2_X2 U4227 ( .A1(fract_denorm[102]), .A2(fract_denorm[101]), .ZN(n5448)
         );
  NAND4_X4 U4228 ( .A1(net59124), .A2(net59125), .A3(net59126), .A4(net59127), 
        .ZN(net59031) );
  NAND2_X4 U4229 ( .A1(net59132), .A2(net59099), .ZN(net59125) );
  NOR3_X4 U4230 ( .A1(net58829), .A2(net58830), .A3(net58831), .ZN(net58828)
         );
  NOR2_X1 U4231 ( .A1(net33554), .A2(n4521), .ZN(n5444) );
  NAND2_X1 U4232 ( .A1(net59578), .A2(u4_fi_ldz_1_), .ZN(n5675) );
  NAND2_X4 U4233 ( .A1(net58440), .A2(net63289), .ZN(net59008) );
  NOR2_X2 U4234 ( .A1(net58440), .A2(net59594), .ZN(net59589) );
  NOR2_X1 U4235 ( .A1(net58440), .A2(n4429), .ZN(n5877) );
  NOR2_X1 U4236 ( .A1(net58440), .A2(n6145), .ZN(net58800) );
  NOR2_X1 U4237 ( .A1(opa_00), .A2(net58440), .ZN(n6048) );
  NOR2_X1 U4238 ( .A1(net58440), .A2(net58623), .ZN(n6044) );
  NOR2_X1 U4239 ( .A1(net58440), .A2(n6146), .ZN(n6147) );
  INV_X8 U4240 ( .A(net58440), .ZN(net58645) );
  NAND2_X1 U4241 ( .A1(net60131), .A2(fract_denorm[75]), .ZN(net60120) );
  NAND3_X1 U4242 ( .A1(net60131), .A2(net60325), .A3(fract_denorm[74]), .ZN(
        net60324) );
  NAND4_X1 U4243 ( .A1(fract_denorm[50]), .A2(net60349), .A3(n5384), .A4(
        net59986), .ZN(n5385) );
  NAND2_X1 U4244 ( .A1(net59986), .A2(net59331), .ZN(net60312) );
  AOI22_X1 U4245 ( .A1(n5418), .A2(n8512), .B1(net59986), .B2(fract_denorm[52]), .ZN(n5439) );
  NAND4_X4 U4246 ( .A1(net60088), .A2(n5403), .A3(net60089), .A4(net60090), 
        .ZN(net59984) );
  NAND4_X4 U4247 ( .A1(n5440), .A2(n5439), .A3(n5438), .A4(net59980), .ZN(
        net59911) );
  NOR3_X2 U4248 ( .A1(fpu_op_r3[1]), .A2(net63089), .A3(n4375), .ZN(net60650)
         );
  INV_X16 U4249 ( .A(net58836), .ZN(net63589) );
  INV_X8 U4250 ( .A(n3652), .ZN(u4_fract_out_37_) );
  AOI22_X4 U4251 ( .A1(u4_N5997), .A2(net63325), .B1(u4_N6105), .B2(net63343), 
        .ZN(n3652) );
  AOI21_X1 U4252 ( .B1(net59084), .B2(u4_exp_out_9_), .A(net59097), .ZN(
        net59091) );
  INV_X8 U4253 ( .A(u4_exp_out_9_), .ZN(net57231) );
  NOR3_X2 U4254 ( .A1(net59030), .A2(net58636), .A3(net59031), .ZN(net59012)
         );
  INV_X1 U4255 ( .A(net58632), .ZN(n4532) );
  NAND3_X1 U4256 ( .A1(net58615), .A2(net58617), .A3(net58616), .ZN(net58613)
         );
  NAND2_X4 U4257 ( .A1(net60051), .A2(net60286), .ZN(net60135) );
  OAI21_X1 U4258 ( .B1(net59209), .B2(net59210), .A(n4516), .ZN(net58676) );
  OAI21_X1 U4259 ( .B1(net57268), .B2(net59901), .A(n4516), .ZN(
        u4_fi_ldz_2a_6_) );
  INV_X32 U4260 ( .A(net63517), .ZN(net63507) );
  NAND2_X4 U4261 ( .A1(n4288), .A2(net63089), .ZN(net58443) );
  AOI22_X4 U4262 ( .A1(fract_out_q[51]), .A2(net63507), .B1(quo[50]), .B2(
        net66895), .ZN(n5115) );
  AOI22_X4 U4263 ( .A1(fract_out_q[52]), .A2(net63507), .B1(quo[51]), .B2(
        net66896), .ZN(n5118) );
  NAND3_X1 U4264 ( .A1(u4_ldz_all_5_), .A2(n6013), .A3(u4_ldz_all_4_), .ZN(
        n6014) );
  NAND2_X4 U4265 ( .A1(net59666), .A2(net59026), .ZN(net59590) );
  NAND2_X1 U4266 ( .A1(n4400), .A2(net59568), .ZN(n5699) );
  NOR2_X2 U4267 ( .A1(n5628), .A2(net59543), .ZN(n5630) );
  AOI211_X4 U4268 ( .C1(net59707), .C2(net59708), .A(net59709), .B(n4652), 
        .ZN(net59704) );
  OAI21_X2 U4269 ( .B1(n4282), .B2(net58980), .A(net58976), .ZN(net58424) );
  OAI21_X2 U4270 ( .B1(n4281), .B2(net58975), .A(net58976), .ZN(net58426) );
  OAI21_X2 U4271 ( .B1(n4281), .B2(net58984), .A(net58976), .ZN(net58419) );
  NOR4_X4 U4272 ( .A1(n4656), .A2(n4654), .A3(n4655), .A4(n4653), .ZN(n4652)
         );
  INV_X8 U4273 ( .A(net58989), .ZN(net58991) );
  NAND3_X1 U4274 ( .A1(net58430), .A2(net58419), .A3(net58421), .ZN(net58579)
         );
  NOR4_X4 U4275 ( .A1(n4710), .A2(net58426), .A3(net58428), .A4(net58427), 
        .ZN(net58528) );
  NAND3_X1 U4276 ( .A1(net57265), .A2(net57260), .A3(n4720), .ZN(net58711) );
  INV_X8 U4277 ( .A(n4720), .ZN(net34244) );
  INV_X8 U4278 ( .A(net58652), .ZN(n4534) );
  INV_X8 U4279 ( .A(u4_N6463), .ZN(net58652) );
  NOR2_X2 U4280 ( .A1(n6126), .A2(net63523), .ZN(N826) );
  NAND4_X4 U4281 ( .A1(net58825), .A2(net58826), .A3(net58827), .A4(net58828), 
        .ZN(net58616) );
  NOR2_X1 U4282 ( .A1(net63527), .A2(n6120), .ZN(N820) );
  NAND4_X1 U4283 ( .A1(net58630), .A2(net58631), .A3(net58632), .A4(net58633), 
        .ZN(net58629) );
  INV_X1 U4284 ( .A(net58716), .ZN(net59269) );
  INV_X8 U4285 ( .A(net59220), .ZN(net59421) );
  OAI221_X1 U4286 ( .B1(n5993), .B2(net58714), .C1(net58735), .C2(net58716), 
        .A(n5992), .ZN(net57260) );
  OAI21_X1 U4287 ( .B1(net60193), .B2(n4517), .A(net60324), .ZN(net60310) );
  NOR2_X1 U4288 ( .A1(n4382), .A2(net59946), .ZN(n5330) );
  OAI21_X1 U4289 ( .B1(net59945), .B2(net59946), .A(net60322), .ZN(net60221)
         );
  OAI21_X1 U4290 ( .B1(fract_denorm[94]), .B2(fract_denorm[96]), .A(net60219), 
        .ZN(n5383) );
  NOR3_X1 U4291 ( .A1(net59945), .A2(fract_denorm[65]), .A3(net59946), .ZN(
        net59941) );
  NOR2_X1 U4292 ( .A1(n4517), .A2(net59993), .ZN(net59988) );
  AOI21_X1 U4293 ( .B1(net59956), .B2(fract_denorm[96]), .A(net59957), .ZN(
        net59955) );
  NOR2_X1 U4294 ( .A1(net60167), .A2(net59946), .ZN(net60164) );
  NOR2_X1 U4295 ( .A1(fract_denorm[68]), .A2(n4517), .ZN(net60040) );
  INV_X2 U4296 ( .A(fract_denorm[96]), .ZN(net60112) );
  NAND3_X2 U4297 ( .A1(net60155), .A2(net60154), .A3(net59918), .ZN(net60305)
         );
  OAI221_X4 U4298 ( .B1(net58716), .B2(net58729), .C1(n4721), .C2(net58714), 
        .A(n4722), .ZN(n4720) );
  AOI221_X4 U4299 ( .B1(net63545), .B2(u4_fract_out_32_), .C1(
        u4_fract_out_pl1_32_), .C2(net63559), .A(net63585), .ZN(n6125) );
  NAND4_X1 U4300 ( .A1(net58471), .A2(n4368), .A3(net58472), .A4(net58591), 
        .ZN(net58590) );
  NOR2_X2 U4301 ( .A1(net63527), .A2(net58471), .ZN(N818) );
  AOI221_X4 U4302 ( .B1(net63541), .B2(u4_fract_out_25_), .C1(
        u4_fract_out_pl1_25_), .C2(net63559), .A(net63587), .ZN(net58471) );
  BUF_X32 U4303 ( .A(u4_exp_out_4_), .Z(net96080) );
  BUF_X32 U4304 ( .A(u4_exp_out_5_), .Z(net87237) );
  NAND2_X4 U4305 ( .A1(net58546), .A2(net58610), .ZN(net58823) );
  INV_X4 U4306 ( .A(net58823), .ZN(net58791) );
  INV_X4 U4307 ( .A(net58432), .ZN(net58610) );
  NAND2_X2 U4308 ( .A1(net58610), .A2(n4461), .ZN(net58437) );
  INV_X8 U4309 ( .A(net58616), .ZN(net58546) );
  NAND3_X1 U4310 ( .A1(net58546), .A2(sign), .A3(net58547), .ZN(net58544) );
  NAND3_X1 U4311 ( .A1(net58546), .A2(n4429), .A3(net58800), .ZN(net58799) );
  NAND2_X2 U4312 ( .A1(net58812), .A2(n4478), .ZN(net58432) );
  INV_X4 U4313 ( .A(net58506), .ZN(net58812) );
  NOR3_X1 U4314 ( .A1(n4485), .A2(net63287), .A3(net58616), .ZN(net58795) );
  NAND2_X2 U4315 ( .A1(net58832), .A2(net58593), .ZN(net58831) );
  INV_X4 U4316 ( .A(net58833), .ZN(net58593) );
  NAND4_X2 U4317 ( .A1(net58593), .A2(net58493), .A3(net58495), .A4(net58494), 
        .ZN(net58589) );
  NAND2_X2 U4318 ( .A1(net58492), .A2(net58477), .ZN(net58833) );
  NOR2_X4 U4319 ( .A1(net58475), .A2(net58526), .ZN(net58832) );
  NAND2_X2 U4320 ( .A1(n4542), .A2(n4543), .ZN(net58830) );
  INV_X4 U4321 ( .A(net58524), .ZN(n4543) );
  INV_X4 U4322 ( .A(net58533), .ZN(n4542) );
  NAND4_X2 U4323 ( .A1(n4368), .A2(net58427), .A3(net58846), .A4(net58847), 
        .ZN(net58829) );
  NOR2_X4 U4324 ( .A1(net58530), .A2(net58848), .ZN(net58847) );
  NAND2_X2 U4325 ( .A1(net58471), .A2(net58430), .ZN(net58848) );
  NAND3_X4 U4326 ( .A1(net58632), .A2(net58964), .A3(net59033), .ZN(net58989)
         );
  NAND2_X1 U4327 ( .A1(net58976), .A2(net58989), .ZN(net58971) );
  INV_X8 U4328 ( .A(net59042), .ZN(net58932) );
  INV_X32 U4329 ( .A(net63295), .ZN(net63291) );
  INV_X32 U4330 ( .A(net63295), .ZN(net63293) );
  INV_X32 U4331 ( .A(net63093), .ZN(net63089) );
  INV_X4 U4332 ( .A(net58631), .ZN(net59034) );
  NAND2_X2 U4333 ( .A1(net58781), .A2(net58787), .ZN(net58964) );
  NAND2_X2 U4334 ( .A1(net58633), .A2(net58964), .ZN(net58963) );
  INV_X4 U4335 ( .A(net58935), .ZN(net58781) );
  NAND2_X2 U4336 ( .A1(n4334), .A2(n4401), .ZN(net59042) );
  NAND2_X2 U4337 ( .A1(rmode_r3[0]), .A2(n4334), .ZN(net58962) );
  NAND2_X2 U4338 ( .A1(net59194), .A2(net59195), .ZN(net59189) );
  INV_X4 U4339 ( .A(net59194), .ZN(net59233) );
  INV_X4 U4340 ( .A(u4_exp_out_6_), .ZN(net59235) );
  INV_X4 U4341 ( .A(u4_exp_out_7_), .ZN(net59234) );
  INV_X8 U4342 ( .A(net59170), .ZN(net59191) );
  NAND3_X4 U4343 ( .A1(net59161), .A2(net59236), .A3(net59237), .ZN(net59170)
         );
  NAND2_X1 U4344 ( .A1(net59170), .A2(net59171), .ZN(net59166) );
  NOR2_X1 U4345 ( .A1(net59170), .A2(net59083), .ZN(net59183) );
  INV_X4 U4346 ( .A(net96080), .ZN(net59237) );
  INV_X4 U4347 ( .A(net87237), .ZN(net59236) );
  INV_X8 U4348 ( .A(n4544), .ZN(net59161) );
  INV_X4 U4349 ( .A(u4_exp_out_3_), .ZN(n4545) );
  INV_X4 U4350 ( .A(net59149), .ZN(net59239) );
  AOI21_X1 U4351 ( .B1(net59099), .B2(net59149), .A(net59169), .ZN(net59120)
         );
  AOI21_X1 U4352 ( .B1(net59148), .B2(net59149), .A(net59083), .ZN(net59142)
         );
  NAND3_X2 U4353 ( .A1(net59112), .A2(net45071), .A3(net59145), .ZN(net59149)
         );
  INV_X2 U4354 ( .A(u4_exp_out_2_), .ZN(net59145) );
  MUX2_X2 U4355 ( .A(net59082), .B(net59083), .S(net45071), .Z(net59074) );
  INV_X4 U4356 ( .A(u4_exp_out_1_), .ZN(net59112) );
  OAI221_X2 U4357 ( .B1(net59588), .B2(net57230), .C1(n2442), .C2(net59112), 
        .A(net59679), .ZN(u4_shift_right[1]) );
  MUX2_X2 U4358 ( .A(net59110), .B(net59111), .S(net59112), .Z(net59107) );
  NAND2_X2 U4359 ( .A1(u4_exp_out_2_), .A2(u4_exp_out_1_), .ZN(net59148) );
  INV_X4 U4360 ( .A(fract_denorm[94]), .ZN(net59918) );
  INV_X4 U4361 ( .A(fract_denorm[93]), .ZN(net60154) );
  NOR3_X4 U4362 ( .A1(fract_denorm[97]), .A2(fract_denorm[96]), .A3(
        fract_denorm[95]), .ZN(net60155) );
  NAND2_X1 U4363 ( .A1(net60219), .A2(net60155), .ZN(net59919) );
  NAND3_X4 U4364 ( .A1(net60599), .A2(net60600), .A3(n4546), .ZN(
        fract_denorm[94]) );
  AOI22_X2 U4365 ( .A1(fract_out_q[45]), .A2(net63511), .B1(net66896), .B2(
        quo[44]), .ZN(n4546) );
  INV_X32 U4366 ( .A(net63515), .ZN(net63511) );
  INV_X32 U4367 ( .A(net63515), .ZN(net63509) );
  MUX2_X2 U4368 ( .A(sign_fasu_r), .B(result_zero_sign_d), .S(net58791), .Z(
        net58821) );
  NAND2_X2 U4369 ( .A1(net58791), .A2(net58792), .ZN(net58790) );
  INV_X4 U4370 ( .A(net58771), .ZN(net58430) );
  NAND2_X2 U4371 ( .A1(net58420), .A2(net58430), .ZN(N853) );
  NAND2_X2 U4372 ( .A1(net58472), .A2(n4547), .ZN(net58530) );
  INV_X4 U4373 ( .A(net58592), .ZN(n4547) );
  NOR2_X4 U4374 ( .A1(net63527), .A2(n4547), .ZN(N816) );
  NAND4_X1 U4375 ( .A1(n4368), .A2(net58528), .A3(net58471), .A4(net58529), 
        .ZN(net58523) );
  NAND2_X4 U4376 ( .A1(net58958), .A2(net58959), .ZN(net58836) );
  NAND2_X2 U4377 ( .A1(net58961), .A2(net58962), .ZN(net58960) );
  INV_X32 U4378 ( .A(net63291), .ZN(net63289) );
  MUX2_X2 U4379 ( .A(net58804), .B(net58805), .S(n4367), .Z(N875) );
  AOI211_X4 U4380 ( .C1(net58793), .C2(n4345), .A(n4367), .B(net58795), .ZN(
        net58789) );
  INV_X4 U4381 ( .A(net58808), .ZN(n4548) );
  MUX2_X2 U4382 ( .A(net58809), .B(net58810), .S(n4470), .Z(net58804) );
  NAND3_X2 U4383 ( .A1(net58540), .A2(n4353), .A3(n4470), .ZN(net58535) );
  XNOR2_X2 U4384 ( .A(sign_mul_r), .B(n4549), .ZN(net58810) );
  NAND2_X2 U4385 ( .A1(net58623), .A2(sign_exe_r), .ZN(n4549) );
  MUX2_X2 U4386 ( .A(net58816), .B(net58817), .S(net58818), .Z(net58809) );
  INV_X32 U4387 ( .A(net63291), .ZN(net63287) );
  NAND2_X2 U4388 ( .A1(ind_d), .A2(n4484), .ZN(net58517) );
  NAND2_X2 U4389 ( .A1(n4482), .A2(n4355), .ZN(net58506) );
  MUX2_X2 U4390 ( .A(n4550), .B(net58820), .S(sign_mul_r), .Z(net58817) );
  NAND2_X2 U4391 ( .A1(net58820), .A2(net58802), .ZN(n4550) );
  MUX2_X2 U4392 ( .A(n4551), .B(net59541), .S(net66839), .Z(net59574) );
  NAND2_X2 U4393 ( .A1(net59574), .A2(net59573), .ZN(u4_shift_left[0]) );
  NOR2_X1 U4394 ( .A1(net58781), .A2(net59568), .ZN(n4551) );
  NAND2_X4 U4395 ( .A1(net58700), .A2(net63293), .ZN(net59541) );
  OAI21_X4 U4396 ( .B1(net59662), .B2(net58440), .A(n4552), .ZN(net59568) );
  INV_X4 U4397 ( .A(net59347), .ZN(net59664) );
  NAND3_X1 U4398 ( .A1(net63083), .A2(fpu_op_r3[0]), .A3(n4288), .ZN(net58935)
         );
  XNOR2_X2 U4399 ( .A(n4553), .B(u4_exp_out_10_), .ZN(net59132) );
  NOR2_X4 U4400 ( .A1(net57231), .A2(net45067), .ZN(net59226) );
  XNOR2_X2 U4401 ( .A(net57231), .B(net59101), .ZN(net59100) );
  OAI221_X2 U4402 ( .B1(net57229), .B2(net57230), .C1(n2442), .C2(net57231), 
        .A(net57232), .ZN(u4_shift_right[9]) );
  NAND2_X2 U4403 ( .A1(net59233), .A2(net59029), .ZN(n4554) );
  INV_X4 U4404 ( .A(u4_exp_out_8_), .ZN(net59029) );
  NOR2_X1 U4405 ( .A1(u4_exp_out_10_), .A2(net59029), .ZN(net59027) );
  NOR2_X4 U4406 ( .A1(net59010), .A2(net59029), .ZN(net59225) );
  INV_X4 U4407 ( .A(net59083), .ZN(net59099) );
  OAI21_X4 U4408 ( .B1(n2408), .B2(net59278), .A(n4555), .ZN(u4_exp_out_10_)
         );
  NAND2_X2 U4409 ( .A1(net58707), .A2(net63293), .ZN(n4555) );
  NAND2_X4 U4410 ( .A1(net58955), .A2(rmode_r3[1]), .ZN(net58948) );
  INV_X4 U4411 ( .A(net58948), .ZN(net59310) );
  AOI21_X2 U4412 ( .B1(net58947), .B2(net58948), .A(n4278), .ZN(net58835) );
  OAI21_X4 U4413 ( .B1(net59311), .B2(sign), .A(net59312), .ZN(net58955) );
  OAI21_X4 U4414 ( .B1(n4556), .B2(net58646), .A(n4557), .ZN(net59312) );
  NAND2_X2 U4415 ( .A1(n4561), .A2(net59321), .ZN(n4560) );
  INV_X4 U4416 ( .A(net33548), .ZN(net59337) );
  NAND2_X2 U4417 ( .A1(net59336), .A2(net59337), .ZN(net60204) );
  INV_X4 U4418 ( .A(net33549), .ZN(net59336) );
  INV_X4 U4419 ( .A(net33550), .ZN(net59335) );
  NAND3_X4 U4420 ( .A1(net60072), .A2(net59335), .A3(net60187), .ZN(net60287)
         );
  INV_X4 U4421 ( .A(net60207), .ZN(net59340) );
  NAND2_X2 U4422 ( .A1(net59340), .A2(net60026), .ZN(net59927) );
  NAND2_X2 U4423 ( .A1(net60208), .A2(net59953), .ZN(net60207) );
  INV_X4 U4424 ( .A(net33641), .ZN(net59953) );
  OAI21_X4 U4425 ( .B1(n2408), .B2(net59270), .A(n4563), .ZN(u4_exp_out_9_) );
  NAND2_X2 U4426 ( .A1(net58759), .A2(net63293), .ZN(n4563) );
  MUX2_X2 U4427 ( .A(quo[55]), .B(quo[107]), .S(opb_dn), .Z(net60649) );
  NAND2_X4 U4428 ( .A1(fpu_op_r3[1]), .A2(fpu_op_r3[0]), .ZN(net60696) );
  OAI21_X1 U4429 ( .B1(net63085), .B2(fpu_op_r3[0]), .A(net63515), .ZN(
        net58438) );
  NAND2_X4 U4430 ( .A1(net59258), .A2(net59259), .ZN(n4565) );
  NAND3_X4 U4431 ( .A1(n4565), .A2(n4564), .A3(net59255), .ZN(u4_exp_out_0_)
         );
  INV_X4 U4432 ( .A(n2408), .ZN(net59259) );
  MUX2_X2 U4433 ( .A(net43686), .B(u4_exp_next_mi_0_), .S(net63221), .Z(
        net59258) );
  INV_X4 U4434 ( .A(net59258), .ZN(net59268) );
  NOR2_X4 U4435 ( .A1(u4_exp_out1_1_), .A2(net59258), .ZN(net59296) );
  INV_X4 U4436 ( .A(net66839), .ZN(net43686) );
  NAND2_X4 U4437 ( .A1(net58777), .A2(net59305), .ZN(n2408) );
  INV_X4 U4438 ( .A(n2399), .ZN(net59305) );
  INV_X4 U4439 ( .A(net59260), .ZN(net58777) );
  AOI22_X2 U4440 ( .A1(u4_exp_next_mi_0_), .A2(net59153), .B1(
        u4_exp_out_pl1_0_), .B2(net59078), .ZN(net59076) );
  INV_X2 U4441 ( .A(n2399), .ZN(net59261) );
  AOI21_X4 U4442 ( .B1(n2404), .B2(net59260), .A(net59694), .ZN(net59693) );
  NOR3_X4 U4443 ( .A1(u4_N6060), .A2(u4_N6059), .A3(u4_N6058), .ZN(n4566) );
  NAND3_X2 U4444 ( .A1(net59487), .A2(net59488), .A3(n4566), .ZN(net59478) );
  INV_X4 U4445 ( .A(net59329), .ZN(net60187) );
  NAND2_X2 U4446 ( .A1(n4567), .A2(net60290), .ZN(net59329) );
  NOR2_X4 U4447 ( .A1(net33572), .A2(net33573), .ZN(n4567) );
  NAND3_X4 U4448 ( .A1(n4568), .A2(n4569), .A3(n4570), .ZN(net33550) );
  NAND2_X2 U4449 ( .A1(quo[20]), .A2(net66910), .ZN(n4570) );
  NAND2_X2 U4450 ( .A1(fract_i2f[18]), .A2(net63083), .ZN(n4569) );
  INV_X32 U4451 ( .A(net63089), .ZN(net63083) );
  INV_X32 U4452 ( .A(net63089), .ZN(net63085) );
  NAND2_X2 U4453 ( .A1(prod[18]), .A2(net66928), .ZN(n4568) );
  OAI21_X2 U4454 ( .B1(net59348), .B2(net59349), .A(net59350), .ZN(net59342)
         );
  NAND4_X2 U4455 ( .A1(net59504), .A2(net59505), .A3(net59506), .A4(n4571), 
        .ZN(net59503) );
  NOR3_X4 U4456 ( .A1(n4572), .A2(n4573), .A3(n4272), .ZN(n4571) );
  INV_X4 U4457 ( .A(n4574), .ZN(n4573) );
  NAND2_X2 U4458 ( .A1(net59517), .A2(n4577), .ZN(n4572) );
  INV_X4 U4459 ( .A(n3704), .ZN(u4_fract_out_12_) );
  AOI221_X2 U4460 ( .B1(net63541), .B2(u4_fract_out_12_), .C1(
        u4_fract_out_pl1_12_), .C2(net63559), .A(net63587), .ZN(net58492) );
  INV_X32 U4461 ( .A(net63347), .ZN(net63341) );
  INV_X32 U4462 ( .A(net63349), .ZN(net63347) );
  INV_X4 U4463 ( .A(net57285), .ZN(net44995) );
  INV_X32 U4464 ( .A(net63327), .ZN(net63321) );
  INV_X32 U4465 ( .A(net63331), .ZN(net63327) );
  INV_X32 U4466 ( .A(net63327), .ZN(net63325) );
  NAND3_X4 U4467 ( .A1(net60097), .A2(net60205), .A3(net60184), .ZN(net59973)
         );
  OAI221_X1 U4468 ( .B1(fract_denorm[104]), .B2(net60007), .C1(net60008), .C2(
        net59973), .A(n4374), .ZN(net59998) );
  NOR2_X1 U4469 ( .A1(net33568), .A2(net59973), .ZN(net59962) );
  NOR2_X1 U4470 ( .A1(net60290), .A2(net59973), .ZN(net60284) );
  INV_X4 U4471 ( .A(net59330), .ZN(net60184) );
  NAND3_X1 U4472 ( .A1(net60184), .A2(net33551), .A3(n4509), .ZN(net60302) );
  NAND3_X4 U4473 ( .A1(net60184), .A2(net59326), .A3(net60185), .ZN(net60183)
         );
  INV_X4 U4474 ( .A(net33551), .ZN(net60205) );
  NAND2_X2 U4475 ( .A1(net60205), .A2(net60206), .ZN(net59341) );
  NAND2_X2 U4476 ( .A1(n4578), .A2(net60096), .ZN(net59330) );
  NOR2_X4 U4477 ( .A1(net33565), .A2(net33566), .ZN(n4578) );
  NAND3_X4 U4478 ( .A1(n4579), .A2(n4580), .A3(n4581), .ZN(net33551) );
  NAND2_X2 U4479 ( .A1(quo[28]), .A2(net66912), .ZN(n4581) );
  NAND2_X2 U4480 ( .A1(fract_i2f[26]), .A2(net63083), .ZN(n4580) );
  NAND2_X2 U4481 ( .A1(prod[26]), .A2(net66929), .ZN(n4579) );
  NAND2_X2 U4482 ( .A1(net63325), .A2(n4582), .ZN(net59449) );
  NAND2_X2 U4483 ( .A1(n4583), .A2(n4584), .ZN(n4582) );
  NOR3_X4 U4484 ( .A1(n4585), .A2(n4586), .A3(n4587), .ZN(n4584) );
  NAND2_X2 U4485 ( .A1(n3930), .A2(n3931), .ZN(n4587) );
  NAND2_X2 U4486 ( .A1(n3928), .A2(n3929), .ZN(n4586) );
  NAND4_X2 U4487 ( .A1(n3934), .A2(n3935), .A3(n3932), .A4(n3933), .ZN(n4585)
         );
  NOR3_X4 U4488 ( .A1(n4588), .A2(n4589), .A3(n4590), .ZN(n4583) );
  NAND2_X2 U4489 ( .A1(n3922), .A2(n3923), .ZN(n4590) );
  NAND2_X2 U4490 ( .A1(n3920), .A2(n3921), .ZN(n4589) );
  NAND4_X2 U4491 ( .A1(n3926), .A2(n3927), .A3(n3924), .A4(n3925), .ZN(n4588)
         );
  NOR2_X4 U4492 ( .A1(net60053), .A2(net59913), .ZN(net59994) );
  INV_X4 U4493 ( .A(net33648), .ZN(n4591) );
  NAND2_X2 U4494 ( .A1(net60082), .A2(n4591), .ZN(net59323) );
  NAND2_X2 U4495 ( .A1(n4515), .A2(fract_denorm[81]), .ZN(net60099) );
  NOR4_X2 U4496 ( .A1(net60162), .A2(net60163), .A3(net60164), .A4(n4593), 
        .ZN(net60098) );
  INV_X4 U4497 ( .A(net33561), .ZN(n4594) );
  NAND2_X2 U4498 ( .A1(net59965), .A2(n4594), .ZN(net60340) );
  INV_X4 U4499 ( .A(fract_denorm[65]), .ZN(net60167) );
  INV_X4 U4500 ( .A(net33625), .ZN(net60086) );
  INV_X4 U4501 ( .A(fract_denorm[97]), .ZN(net60168) );
  NAND2_X4 U4502 ( .A1(net60111), .A2(net59428), .ZN(net60006) );
  NOR2_X1 U4503 ( .A1(net60005), .A2(net60006), .ZN(net59999) );
  NOR3_X1 U4504 ( .A1(net60204), .A2(net59322), .A3(net60006), .ZN(net60180)
         );
  NAND3_X1 U4505 ( .A1(net60219), .A2(net60112), .A3(net60113), .ZN(net60110)
         );
  NAND3_X1 U4506 ( .A1(net59428), .A2(net59427), .A3(net59429), .ZN(net59426)
         );
  NAND2_X4 U4507 ( .A1(net59429), .A2(net63221), .ZN(net59961) );
  NAND2_X2 U4508 ( .A1(u4_exp_next_mi_11_), .A2(net63221), .ZN(net59696) );
  MUX2_X2 U4509 ( .A(net59594), .B(net59892), .S(net63221), .Z(net59891) );
  NAND2_X2 U4510 ( .A1(n4596), .A2(net63221), .ZN(net60038) );
  INV_X4 U4511 ( .A(fract_denorm[99]), .ZN(n4595) );
  INV_X4 U4512 ( .A(fract_denorm[98]), .ZN(n4597) );
  INV_X4 U4513 ( .A(n4598), .ZN(n4596) );
  NAND2_X2 U4514 ( .A1(net59920), .A2(net59958), .ZN(n4598) );
  NOR2_X4 U4515 ( .A1(net59123), .A2(net59031), .ZN(net58973) );
  NAND4_X2 U4516 ( .A1(net58973), .A2(net58984), .A3(net58975), .A4(net59071), 
        .ZN(net59069) );
  AOI211_X1 U4517 ( .C1(net59084), .C2(u4_exp_out_10_), .A(net59128), .B(
        net59129), .ZN(net59127) );
  NOR2_X4 U4518 ( .A1(net59081), .A2(n4599), .ZN(net59129) );
  INV_X4 U4519 ( .A(u4_exp_fix_diva[10]), .ZN(n4599) );
  NOR2_X4 U4520 ( .A1(net59087), .A2(n4600), .ZN(net59128) );
  INV_X4 U4521 ( .A(u4_exp_fix_divb[10]), .ZN(n4600) );
  NAND2_X2 U4522 ( .A1(u4_exp_next_mi_10_), .A2(net59117), .ZN(net59126) );
  INV_X4 U4523 ( .A(net59079), .ZN(net59117) );
  OAI21_X4 U4524 ( .B1(net59048), .B2(net59009), .A(net59049), .ZN(net59044)
         );
  AOI21_X4 U4525 ( .B1(net59044), .B2(net63293), .A(net59045), .ZN(net59038)
         );
  NAND2_X2 U4526 ( .A1(net58994), .A2(net59050), .ZN(net59049) );
  NAND2_X2 U4527 ( .A1(n4486), .A2(net58674), .ZN(net59050) );
  INV_X4 U4528 ( .A(net59054), .ZN(net59053) );
  INV_X4 U4529 ( .A(net59017), .ZN(net58994) );
  NAND2_X2 U4530 ( .A1(net59041), .A2(net58994), .ZN(net59040) );
  OAI21_X4 U4531 ( .B1(net59068), .B2(net59069), .A(net59070), .ZN(net59048)
         );
  AND2_X2 U4532 ( .A1(net58980), .A2(net58982), .ZN(n4607) );
  INV_X4 U4533 ( .A(net59009), .ZN(net59007) );
  INV_X4 U4534 ( .A(u4_fi_ldz_2a_6_), .ZN(net59021) );
  NAND2_X2 U4535 ( .A1(n4603), .A2(n4606), .ZN(n4605) );
  INV_X4 U4536 ( .A(u4_fi_ldz_2a_2_), .ZN(n4606) );
  INV_X4 U4537 ( .A(net44706), .ZN(n4603) );
  NOR2_X4 U4538 ( .A1(net59024), .A2(n4603), .ZN(n4602) );
  INV_X4 U4539 ( .A(n4608), .ZN(u4_fi_ldz_2a_5_) );
  XNOR2_X2 U4540 ( .A(net59901), .B(u4_fi_ldz_5_), .ZN(n4608) );
  NAND2_X2 U4541 ( .A1(u4_exp_in_mi1_11_), .A2(net59566), .ZN(net58674) );
  INV_X4 U4542 ( .A(net66835), .ZN(net59566) );
  NOR2_X4 U4543 ( .A1(net58550), .A2(net59566), .ZN(net59674) );
  NOR2_X4 U4544 ( .A1(u4_N6057), .A2(u4_N6056), .ZN(net59488) );
  NOR2_X4 U4545 ( .A1(u4_N6055), .A2(u4_N6054), .ZN(net59487) );
  NAND3_X2 U4546 ( .A1(net60133), .A2(net60134), .A3(net33581), .ZN(n4609) );
  INV_X4 U4547 ( .A(net33579), .ZN(net60134) );
  OAI21_X4 U4548 ( .B1(net60134), .B2(net60135), .A(net60275), .ZN(net60095)
         );
  INV_X4 U4549 ( .A(net60135), .ZN(net60133) );
  NAND3_X4 U4550 ( .A1(n4610), .A2(n4611), .A3(n4612), .ZN(net33581) );
  NAND2_X2 U4551 ( .A1(quo[13]), .A2(net66912), .ZN(n4612) );
  NAND2_X2 U4552 ( .A1(fract_i2f[11]), .A2(net63085), .ZN(n4611) );
  NAND2_X2 U4553 ( .A1(prod[11]), .A2(net66930), .ZN(n4610) );
  INV_X32 U4554 ( .A(net66927), .ZN(net66930) );
  INV_X32 U4555 ( .A(net59840), .ZN(net66927) );
  INV_X32 U4556 ( .A(net66927), .ZN(net66929) );
  INV_X32 U4557 ( .A(net66927), .ZN(net66928) );
  NAND2_X4 U4558 ( .A1(net60191), .A2(net60022), .ZN(net60282) );
  NOR3_X4 U4559 ( .A1(net60282), .A2(fract_denorm[76]), .A3(net60202), .ZN(
        net60131) );
  INV_X4 U4560 ( .A(net59283), .ZN(net59278) );
  OAI21_X2 U4561 ( .B1(net58651), .B2(net58652), .A(net59566), .ZN(net59666)
         );
  OAI21_X4 U4562 ( .B1(exp_ovf_r_0_), .B2(net58662), .A(net59566), .ZN(
        net59563) );
  INV_X4 U4563 ( .A(net59667), .ZN(net58651) );
  NAND2_X2 U4564 ( .A1(net58645), .A2(net58651), .ZN(net59307) );
  MUX2_X2 U4565 ( .A(net59668), .B(net59669), .S(net63221), .Z(net59667) );
  INV_X4 U4566 ( .A(u4_exp_next_mi_11_), .ZN(net59669) );
  INV_X4 U4567 ( .A(u4_exp_in_pl1_11_), .ZN(net59668) );
  NAND3_X4 U4568 ( .A1(net60646), .A2(net60647), .A3(n4613), .ZN(
        fract_denorm_105_) );
  AOI21_X4 U4569 ( .B1(net60649), .B2(net63293), .A(net60650), .ZN(n4613) );
  NOR2_X4 U4570 ( .A1(net59946), .A2(net60200), .ZN(net60093) );
  NAND3_X2 U4571 ( .A1(net60093), .A2(net60192), .A3(net60196), .ZN(net60002)
         );
  AOI22_X1 U4572 ( .A1(fract_denorm[92]), .A2(net60092), .B1(n4520), .B2(
        fract_denorm[60]), .ZN(net60089) );
  NAND3_X1 U4573 ( .A1(n4520), .A2(net60132), .A3(fract_denorm[59]), .ZN(
        net60119) );
  NAND2_X2 U4574 ( .A1(n4614), .A2(net60329), .ZN(net60200) );
  NOR2_X4 U4575 ( .A1(net60200), .A2(net60201), .ZN(net60199) );
  NOR2_X4 U4576 ( .A1(fract_denorm[65]), .A2(fract_denorm[64]), .ZN(n4614) );
  INV_X4 U4577 ( .A(fract_denorm[66]), .ZN(net60194) );
  NAND4_X2 U4578 ( .A1(net60193), .A2(net60194), .A3(net60349), .A4(net60196), 
        .ZN(net60189) );
  NAND4_X2 U4579 ( .A1(net59113), .A2(net59114), .A3(n4615), .A4(n4616), .ZN(
        net58984) );
  AOI22_X2 U4580 ( .A1(u4_exp_next_mi_3_), .A2(net59117), .B1(
        u4_exp_out_pl1_3_), .B2(net59078), .ZN(n4616) );
  MUX2_X2 U4581 ( .A(n4369), .B(net59159), .S(net96080), .Z(net59155) );
  INV_X2 U4582 ( .A(net59120), .ZN(net59118) );
  INV_X4 U4583 ( .A(net59353), .ZN(net59351) );
  NAND2_X2 U4584 ( .A1(net58643), .A2(n4404), .ZN(net59306) );
  NAND2_X2 U4585 ( .A1(net58666), .A2(n4404), .ZN(net58658) );
  OAI21_X4 U4586 ( .B1(net59038), .B2(net59039), .A(net59040), .ZN(net58657)
         );
  INV_X4 U4587 ( .A(net59008), .ZN(net58792) );
  INV_X4 U4588 ( .A(net59026), .ZN(u4_exp_in_mi1_11_) );
  NAND2_X2 U4589 ( .A1(net58650), .A2(net63289), .ZN(net59046) );
  NAND3_X2 U4590 ( .A1(net59477), .A2(net59476), .A3(net59475), .ZN(net59459)
         );
  INV_X4 U4591 ( .A(u4_N6063), .ZN(n4619) );
  INV_X4 U4592 ( .A(u4_N6062), .ZN(n4618) );
  INV_X4 U4593 ( .A(u4_N6061), .ZN(n4617) );
  INV_X4 U4594 ( .A(u4_N6066), .ZN(n4622) );
  INV_X4 U4595 ( .A(u4_N6065), .ZN(n4621) );
  INV_X4 U4596 ( .A(u4_N6064), .ZN(n4620) );
  INV_X4 U4597 ( .A(net58968), .ZN(net58427) );
  INV_X4 U4598 ( .A(net58972), .ZN(net58969) );
  OAI21_X4 U4599 ( .B1(net58986), .B2(net58970), .A(net58971), .ZN(net58581)
         );
  NAND4_X2 U4600 ( .A1(net59073), .A2(net59074), .A3(n4623), .A4(net59076), 
        .ZN(net58972) );
  NAND2_X2 U4601 ( .A1(u4_exp_fix_diva[0]), .A2(net59121), .ZN(n4623) );
  INV_X4 U4602 ( .A(net59084), .ZN(net59082) );
  AOI22_X2 U4603 ( .A1(net59085), .A2(net66839), .B1(u4_exp_fix_divb[0]), .B2(
        net59122), .ZN(net59073) );
  INV_X4 U4604 ( .A(net59088), .ZN(net59085) );
  NOR2_X1 U4605 ( .A1(net58772), .A2(net58581), .ZN(net58846) );
  NOR3_X4 U4606 ( .A1(net58491), .A2(net58489), .A3(net58487), .ZN(n4626) );
  NOR2_X4 U4607 ( .A1(net58485), .A2(net58483), .ZN(n4625) );
  NOR2_X4 U4608 ( .A1(net58481), .A2(net58479), .ZN(n4624) );
  NAND3_X2 U4609 ( .A1(net58476), .A2(net58477), .A3(net58492), .ZN(net58525)
         );
  NOR2_X2 U4610 ( .A1(net63529), .A2(net58492), .ZN(N805) );
  NAND3_X4 U4611 ( .A1(n4514), .A2(net60206), .A3(net59326), .ZN(net59966) );
  INV_X4 U4612 ( .A(net33552), .ZN(net60206) );
  NOR3_X4 U4613 ( .A1(net59991), .A2(net33558), .A3(net33559), .ZN(net59326)
         );
  NAND3_X4 U4614 ( .A1(n4627), .A2(n4628), .A3(n4629), .ZN(net33552) );
  NAND2_X2 U4615 ( .A1(quo[36]), .A2(net66910), .ZN(n4629) );
  NAND2_X2 U4616 ( .A1(fract_i2f[34]), .A2(net63083), .ZN(n4628) );
  NAND2_X2 U4617 ( .A1(prod[34]), .A2(net66930), .ZN(n4627) );
  OAI21_X4 U4618 ( .B1(n3865), .B2(net63287), .A(net59315), .ZN(net59220) );
  OAI21_X1 U4619 ( .B1(u4_fract_out_0_), .B2(net59220), .A(net59243), .ZN(
        net58957) );
  NAND3_X1 U4620 ( .A1(net58650), .A2(net59220), .A3(net59221), .ZN(net59208)
         );
  NAND2_X2 U4621 ( .A1(n3865), .A2(net59315), .ZN(net58646) );
  NAND2_X2 U4622 ( .A1(net58682), .A2(net63293), .ZN(net58779) );
  INV_X4 U4623 ( .A(net58779), .ZN(net58778) );
  INV_X4 U4624 ( .A(net59243), .ZN(net59222) );
  NOR4_X4 U4625 ( .A1(net59459), .A2(net59460), .A3(net59461), .A4(net59462), 
        .ZN(net59448) );
  NOR2_X4 U4626 ( .A1(n4630), .A2(n4631), .ZN(net59476) );
  INV_X4 U4627 ( .A(u4_N6050), .ZN(n4634) );
  INV_X4 U4628 ( .A(u4_N6049), .ZN(n4633) );
  INV_X4 U4629 ( .A(u4_N6048), .ZN(n4632) );
  INV_X4 U4630 ( .A(u4_N6053), .ZN(n4637) );
  INV_X4 U4631 ( .A(u4_N6052), .ZN(n4636) );
  INV_X4 U4632 ( .A(u4_N6051), .ZN(n4635) );
  NOR3_X4 U4633 ( .A1(n4638), .A2(u4_N6047), .A3(n4639), .ZN(net59475) );
  INV_X4 U4634 ( .A(n4640), .ZN(n4639) );
  NOR2_X4 U4635 ( .A1(u4_N6046), .A2(u4_N6045), .ZN(n4640) );
  NAND2_X2 U4636 ( .A1(n4641), .A2(n4642), .ZN(n4638) );
  NOR2_X4 U4637 ( .A1(u4_N6044), .A2(u4_N6043), .ZN(n4642) );
  NOR2_X4 U4638 ( .A1(u4_N6042), .A2(u4_N6041), .ZN(n4641) );
  NAND3_X4 U4639 ( .A1(net58635), .A2(net58624), .A3(net59208), .ZN(net59088)
         );
  NAND2_X2 U4640 ( .A1(net58950), .A2(net58963), .ZN(net58958) );
  NAND2_X2 U4641 ( .A1(sign), .A2(rmode_r3[1]), .ZN(net58961) );
  INV_X4 U4642 ( .A(net58961), .ZN(net58998) );
  INV_X4 U4643 ( .A(net58962), .ZN(net58624) );
  NAND3_X2 U4644 ( .A1(net58528), .A2(net58935), .A3(net58962), .ZN(net58637)
         );
  NOR2_X4 U4645 ( .A1(fract_denorm[68]), .A2(fract_denorm[67]), .ZN(net60193)
         );
  NAND3_X4 U4646 ( .A1(net60536), .A2(net60537), .A3(n4643), .ZN(
        fract_denorm[66]) );
  AOI22_X2 U4647 ( .A1(fract_out_q[17]), .A2(net63503), .B1(quo[16]), .B2(
        net66895), .ZN(n4643) );
  INV_X32 U4648 ( .A(net63517), .ZN(net63503) );
  INV_X4 U4649 ( .A(u4_fract_out_pl1_52_), .ZN(net59219) );
  INV_X4 U4650 ( .A(net57241), .ZN(net59427) );
  NOR3_X4 U4651 ( .A1(net59430), .A2(n4647), .A3(n4648), .ZN(n4646) );
  INV_X4 U4652 ( .A(net57240), .ZN(n4648) );
  INV_X4 U4653 ( .A(n4650), .ZN(n4647) );
  NAND2_X2 U4654 ( .A1(n4647), .A2(net59427), .ZN(net59799) );
  XNOR2_X2 U4655 ( .A(net66863), .B(n4649), .ZN(n4650) );
  INV_X4 U4656 ( .A(n4651), .ZN(n4649) );
  NAND2_X2 U4657 ( .A1(n4649), .A2(net66863), .ZN(net59812) );
  NAND2_X2 U4658 ( .A1(n4649), .A2(net59442), .ZN(net59433) );
  NAND2_X2 U4659 ( .A1(net59678), .A2(net59792), .ZN(n4651) );
  NAND3_X4 U4660 ( .A1(net59704), .A2(net59705), .A3(net59706), .ZN(net58716)
         );
  NOR2_X4 U4661 ( .A1(u4_div_exp2_10_), .A2(u4_div_exp2_9_), .ZN(net59706) );
  INV_X4 U4662 ( .A(u4_div_exp2_8_), .ZN(net59705) );
  INV_X4 U4663 ( .A(u4_div_exp2_7_), .ZN(n4656) );
  INV_X4 U4664 ( .A(u4_div_exp2_6_), .ZN(n4655) );
  NAND2_X2 U4665 ( .A1(u4_div_exp2_5_), .A2(u4_div_exp2_4_), .ZN(n4654) );
  NAND4_X2 U4666 ( .A1(u4_div_exp2_1_), .A2(u4_div_exp2_0_), .A3(
        u4_div_exp2_3_), .A4(u4_div_exp2_2_), .ZN(n4653) );
  NAND2_X2 U4667 ( .A1(opa_dn), .A2(net59703), .ZN(net59709) );
  INV_X4 U4668 ( .A(net59715), .ZN(net59708) );
  OAI211_X2 U4669 ( .C1(n4658), .C2(net59721), .A(net59722), .B(net59723), 
        .ZN(n4657) );
  INV_X4 U4670 ( .A(net59724), .ZN(n4658) );
  INV_X4 U4671 ( .A(net59726), .ZN(n4659) );
  INV_X4 U4672 ( .A(u4_div_exp2_4_), .ZN(net58741) );
  INV_X4 U4673 ( .A(u4_div_exp2_1_), .ZN(net59700) );
  AOI22_X2 U4674 ( .A1(u4_div_exp1_0_), .A2(net58718), .B1(net59269), .B2(
        u4_div_exp2_0_), .ZN(net59265) );
  INV_X4 U4675 ( .A(u4_div_exp2_3_), .ZN(net58735) );
  INV_X4 U4676 ( .A(u4_div_exp2_2_), .ZN(net58762) );
  NAND3_X4 U4677 ( .A1(n4660), .A2(net60607), .A3(net60606), .ZN(
        fract_denorm[97]) );
  AOI22_X2 U4678 ( .A1(fract_out_q[48]), .A2(net63507), .B1(quo[47]), .B2(
        net66896), .ZN(n4660) );
  NAND3_X2 U4679 ( .A1(net60131), .A2(net60353), .A3(net60325), .ZN(net60352)
         );
  INV_X4 U4680 ( .A(fract_denorm[75]), .ZN(net60325) );
  INV_X4 U4681 ( .A(fract_denorm[74]), .ZN(net60353) );
  NAND3_X4 U4682 ( .A1(net60548), .A2(net60549), .A3(n4661), .ZN(
        fract_denorm[75]) );
  AOI22_X2 U4683 ( .A1(fract_out_q[26]), .A2(net63513), .B1(quo[25]), .B2(
        net66895), .ZN(n4661) );
  NAND2_X2 U4684 ( .A1(net60004), .A2(n4663), .ZN(net60308) );
  INV_X4 U4685 ( .A(fract_denorm[70]), .ZN(n4665) );
  INV_X4 U4686 ( .A(fract_denorm[69]), .ZN(n4662) );
  NAND3_X4 U4687 ( .A1(net60136), .A2(net60137), .A3(n4666), .ZN(net59912) );
  NOR2_X4 U4688 ( .A1(net60139), .A2(n4323), .ZN(n4666) );
  AOI21_X4 U4689 ( .B1(net59262), .B2(net63293), .A(n4667), .ZN(net59255) );
  INV_X4 U4690 ( .A(n4527), .ZN(net44696) );
  NAND4_X2 U4691 ( .A1(n4668), .A2(n4669), .A3(n4670), .A4(n4671), .ZN(
        net59462) );
  INV_X4 U4692 ( .A(u4_N6020), .ZN(n4671) );
  NOR2_X4 U4693 ( .A1(u4_N6019), .A2(u4_N6018), .ZN(n4670) );
  NOR2_X4 U4694 ( .A1(u4_N6017), .A2(u4_N6016), .ZN(n4669) );
  NAND4_X2 U4695 ( .A1(n4672), .A2(n4673), .A3(n4674), .A4(n4675), .ZN(
        net59461) );
  INV_X4 U4696 ( .A(u4_N6027), .ZN(n4675) );
  NOR2_X4 U4697 ( .A1(u4_N6026), .A2(u4_N6025), .ZN(n4674) );
  NOR2_X4 U4698 ( .A1(u4_N6024), .A2(u4_N6023), .ZN(n4673) );
  NOR2_X4 U4699 ( .A1(u4_N6022), .A2(u4_N6021), .ZN(n4672) );
  NAND4_X2 U4700 ( .A1(n4676), .A2(n4677), .A3(n4678), .A4(n4679), .ZN(
        net59460) );
  NOR3_X4 U4701 ( .A1(u4_N6040), .A2(u4_N6039), .A3(u4_N6038), .ZN(n4679) );
  NOR3_X4 U4702 ( .A1(u4_N6037), .A2(u4_N6036), .A3(u4_N6035), .ZN(n4678) );
  NOR3_X4 U4703 ( .A1(u4_N6034), .A2(u4_N6033), .A3(u4_N6032), .ZN(n4677) );
  NOR4_X2 U4704 ( .A1(u4_N6031), .A2(u4_N6030), .A3(u4_N6029), .A4(u4_N6028), 
        .ZN(n4676) );
  NAND3_X4 U4705 ( .A1(net60610), .A2(net60611), .A3(n4680), .ZN(
        fract_denorm[96]) );
  NAND2_X2 U4706 ( .A1(quo[98]), .A2(net66907), .ZN(net60611) );
  AOI22_X2 U4707 ( .A1(u4_exp_fix_diva[3]), .A2(net59121), .B1(
        u4_exp_fix_divb[3]), .B2(net59122), .ZN(net59114) );
  INV_X4 U4708 ( .A(net59081), .ZN(net59121) );
  NAND2_X2 U4709 ( .A1(net59093), .A2(net66851), .ZN(net59113) );
  INV_X32 U4710 ( .A(net66850), .ZN(net66851) );
  INV_X4 U4711 ( .A(n4685), .ZN(n4684) );
  NAND3_X4 U4712 ( .A1(n4321), .A2(n4686), .A3(net33587), .ZN(n4685) );
  INV_X4 U4713 ( .A(net33586), .ZN(n4686) );
  NAND2_X2 U4714 ( .A1(net60346), .A2(n4686), .ZN(net60318) );
  NAND2_X2 U4715 ( .A1(n4321), .A2(net33586), .ZN(net60090) );
  INV_X4 U4716 ( .A(fract_denorm[91]), .ZN(net60128) );
  INV_X4 U4717 ( .A(net33566), .ZN(net60129) );
  INV_X4 U4718 ( .A(net60096), .ZN(net60130) );
  INV_X4 U4719 ( .A(fract_denorm[60]), .ZN(net60132) );
  NAND3_X4 U4720 ( .A1(net60461), .A2(net60462), .A3(n4687), .ZN(net33587) );
  NAND2_X2 U4721 ( .A1(quo[45]), .A2(net66910), .ZN(n4687) );
  INV_X4 U4722 ( .A(net58656), .ZN(net58633) );
  NAND2_X4 U4723 ( .A1(net58991), .A2(net58633), .ZN(net58974) );
  NAND4_X2 U4724 ( .A1(net58633), .A2(net58773), .A3(net58774), .A4(net58775), 
        .ZN(net58609) );
  NAND2_X2 U4725 ( .A1(u4_N6917), .A2(net59664), .ZN(net59345) );
  INV_X4 U4726 ( .A(net58926), .ZN(net58780) );
  NAND2_X4 U4727 ( .A1(n4523), .A2(n4522), .ZN(net60159) );
  NOR4_X1 U4728 ( .A1(net60157), .A2(net60158), .A3(net33584), .A4(net60159), 
        .ZN(net60151) );
  INV_X4 U4729 ( .A(net59331), .ZN(net60348) );
  NAND2_X2 U4730 ( .A1(net60185), .A2(net60349), .ZN(net59331) );
  INV_X4 U4731 ( .A(fract_denorm[52]), .ZN(net60349) );
  NOR3_X1 U4732 ( .A1(net58656), .A2(net63287), .A3(net58657), .ZN(net58655)
         );
  NAND2_X2 U4733 ( .A1(rmode_r3[1]), .A2(n4462), .ZN(net59039) );
  INV_X4 U4734 ( .A(fract_denorm[54]), .ZN(n4690) );
  INV_X4 U4735 ( .A(fract_denorm[53]), .ZN(n4688) );
  INV_X4 U4736 ( .A(net60065), .ZN(n4689) );
  INV_X4 U4737 ( .A(fract_denorm[58]), .ZN(net60192) );
  NOR2_X1 U4738 ( .A1(net60065), .A2(n4533), .ZN(net59922) );
  NAND3_X4 U4739 ( .A1(net60652), .A2(net60653), .A3(n4691), .ZN(
        fract_denorm[76]) );
  AOI22_X2 U4740 ( .A1(fract_out_q[27]), .A2(net63509), .B1(quo[26]), .B2(
        net66895), .ZN(n4691) );
  NAND2_X4 U4741 ( .A1(n4692), .A2(net59540), .ZN(net59026) );
  INV_X4 U4742 ( .A(net59553), .ZN(net59540) );
  INV_X4 U4743 ( .A(net59886), .ZN(n4692) );
  NAND2_X2 U4744 ( .A1(n4692), .A2(n4505), .ZN(net59888) );
  OAI211_X4 U4745 ( .C1(net59231), .C2(net59306), .A(net59307), .B(n4693), 
        .ZN(n2399) );
  INV_X4 U4746 ( .A(net60235), .ZN(net60106) );
  INV_X4 U4747 ( .A(fract_denorm[64]), .ZN(net59945) );
  INV_X4 U4748 ( .A(fract_denorm[63]), .ZN(net60142) );
  INV_X4 U4749 ( .A(net60144), .ZN(net60139) );
  NAND4_X2 U4750 ( .A1(net33578), .A2(net60051), .A3(net60146), .A4(net60145), 
        .ZN(net60144) );
  INV_X4 U4751 ( .A(net33577), .ZN(net60146) );
  INV_X4 U4752 ( .A(net60147), .ZN(net60145) );
  INV_X4 U4753 ( .A(net33563), .ZN(n4695) );
  INV_X4 U4754 ( .A(net60150), .ZN(n4694) );
  OAI211_X2 U4755 ( .C1(n4446), .C2(net58792), .A(net58941), .B(net58803), 
        .ZN(net58966) );
  AOI21_X4 U4756 ( .B1(net59198), .B2(net66835), .A(net58966), .ZN(net58976)
         );
  NOR3_X4 U4757 ( .A1(net60147), .A2(net33577), .A3(net33578), .ZN(net60286)
         );
  NAND2_X2 U4758 ( .A1(net60330), .A2(net60286), .ZN(net59328) );
  OAI21_X4 U4759 ( .B1(net66835), .B2(n4696), .A(net58993), .ZN(net58656) );
  INV_X4 U4760 ( .A(net58997), .ZN(net58995) );
  NAND2_X2 U4761 ( .A1(net59007), .A2(net59008), .ZN(n4702) );
  NOR3_X1 U4762 ( .A1(u4_exp_out_10_), .A2(u4_exp_out_0_), .A3(u4_exp_out_9_), 
        .ZN(n4700) );
  NOR2_X4 U4763 ( .A1(net63287), .A2(n4703), .ZN(n4697) );
  NAND3_X4 U4764 ( .A1(n4706), .A2(n4707), .A3(n4708), .ZN(net33547) );
  NAND2_X2 U4765 ( .A1(quo[44]), .A2(net66911), .ZN(n4708) );
  INV_X8 U4766 ( .A(n4305), .ZN(net66911) );
  NAND2_X2 U4767 ( .A1(fract_i2f[42]), .A2(net63083), .ZN(n4707) );
  NAND2_X2 U4768 ( .A1(prod[42]), .A2(net66928), .ZN(n4706) );
  INV_X4 U4769 ( .A(net59322), .ZN(net60344) );
  NAND2_X2 U4770 ( .A1(net60317), .A2(net60345), .ZN(net59322) );
  INV_X4 U4771 ( .A(net60318), .ZN(net60345) );
  INV_X4 U4772 ( .A(net60317), .ZN(net60314) );
  NAND2_X1 U4773 ( .A1(net58638), .A2(net58637), .ZN(net58628) );
  NAND3_X1 U4774 ( .A1(net58428), .A2(net58427), .A3(net58429), .ZN(net58580)
         );
  NAND2_X2 U4775 ( .A1(net58420), .A2(net58428), .ZN(N855) );
  NAND3_X2 U4776 ( .A1(n4709), .A2(net58581), .A3(net58771), .ZN(n4710) );
  INV_X4 U4777 ( .A(n4711), .ZN(n4709) );
  NAND2_X2 U4778 ( .A1(n4712), .A2(n4713), .ZN(n4711) );
  NOR3_X4 U4779 ( .A1(net58425), .A2(net58423), .A3(net58424), .ZN(n4713) );
  NOR3_X1 U4780 ( .A1(net58581), .A2(net58426), .A3(net58772), .ZN(net58768)
         );
  NAND2_X2 U4781 ( .A1(net58426), .A2(net58425), .ZN(net58584) );
  NAND2_X2 U4782 ( .A1(net58420), .A2(net58426), .ZN(N846) );
  NOR2_X4 U4783 ( .A1(fract_denorm[60]), .A2(fract_denorm[59]), .ZN(net60196)
         );
  NAND3_X4 U4784 ( .A1(net60509), .A2(net60510), .A3(n4714), .ZN(
        fract_denorm[58]) );
  AOI22_X2 U4785 ( .A1(fract_out_q[9]), .A2(net63511), .B1(net66896), .B2(
        quo[8]), .ZN(n4714) );
  NAND2_X2 U4786 ( .A1(quo[46]), .A2(net66911), .ZN(net60460) );
  NAND2_X2 U4787 ( .A1(u4_exp_out_pl1_10_), .A2(net59078), .ZN(net59124) );
  OAI21_X4 U4788 ( .B1(net59215), .B2(net59193), .A(net59192), .ZN(net59084)
         );
  NAND2_X4 U4789 ( .A1(net66928), .A2(net63089), .ZN(net58440) );
  NAND3_X4 U4790 ( .A1(net60587), .A2(net60588), .A3(n4715), .ZN(
        fract_denorm[92]) );
  AOI22_X2 U4791 ( .A1(fract_out_q[43]), .A2(net63513), .B1(quo[42]), .B2(
        net66896), .ZN(n4715) );
  NAND2_X2 U4792 ( .A1(net66851), .A2(n4386), .ZN(net59717) );
  OAI21_X4 U4793 ( .B1(net59850), .B2(net59765), .A(net59717), .ZN(net59865)
         );
  NAND2_X2 U4794 ( .A1(net59265), .A2(n4716), .ZN(net59262) );
  AOI22_X2 U4795 ( .A1(net59267), .A2(net59268), .B1(u4_div_exp3[0]), .B2(
        net58719), .ZN(n4716) );
  INV_X4 U4796 ( .A(net58714), .ZN(net59267) );
  INV_X4 U4797 ( .A(net58752), .ZN(net58718) );
  NOR3_X4 U4798 ( .A1(net59982), .A2(net63217), .A3(net59976), .ZN(net59996)
         );
  INV_X32 U4799 ( .A(net63221), .ZN(net63217) );
  OAI21_X1 U4800 ( .B1(n4718), .B2(n4533), .A(n4719), .ZN(n4717) );
  NAND2_X2 U4801 ( .A1(net60004), .A2(fract_denorm[73]), .ZN(n4719) );
  INV_X4 U4802 ( .A(fract_denorm[57]), .ZN(n4718) );
  INV_X4 U4803 ( .A(fract_denorm[89]), .ZN(net60005) );
  AOI22_X2 U4804 ( .A1(u4_div_exp3[5]), .A2(net58719), .B1(u4_div_exp1_5_), 
        .B2(net58718), .ZN(n4722) );
  INV_X4 U4805 ( .A(net44770), .ZN(n4723) );
  NOR2_X4 U4806 ( .A1(n4723), .A2(net58733), .ZN(net58728) );
  NAND2_X4 U4807 ( .A1(net58550), .A2(net58674), .ZN(net58714) );
  INV_X4 U4808 ( .A(net59070), .ZN(net58550) );
  NAND3_X2 U4809 ( .A1(n6121), .A2(n6120), .A3(n6119), .ZN(n5917) );
  NOR2_X2 U4810 ( .A1(net63523), .A2(n6123), .ZN(N823) );
  INV_X2 U4811 ( .A(n4724), .ZN(n4725) );
  INV_X4 U4812 ( .A(n4726), .ZN(n4727) );
  INV_X4 U4813 ( .A(n4728), .ZN(n4729) );
  INV_X8 U4814 ( .A(n4773), .ZN(n4787) );
  NAND3_X1 U4815 ( .A1(n4727), .A2(n4962), .A3(n4348), .ZN(n4950) );
  NAND2_X1 U4816 ( .A1(net58420), .A2(net58427), .ZN(N845) );
  NOR2_X1 U4817 ( .A1(net58427), .A2(net58771), .ZN(net58769) );
  OAI21_X1 U4818 ( .B1(n4276), .B2(n5807), .A(n7159), .ZN(u4_fi_ldz_mi22[6])
         );
  XNOR2_X1 U4819 ( .A(n4276), .B(n7164), .ZN(n7165) );
  OAI221_X1 U4820 ( .B1(n5996), .B2(net58714), .C1(n4655), .C2(n4518), .A(
        n5995), .ZN(n5997) );
  OAI221_X1 U4821 ( .B1(net58716), .B2(net59700), .C1(net59701), .C2(net58714), 
        .A(n5607), .ZN(n5973) );
  NOR2_X1 U4822 ( .A1(u4_fi_ldz_5_), .A2(n4276), .ZN(n5806) );
  OAI21_X1 U4823 ( .B1(u4_fi_ldz_5_), .B2(n5479), .A(n4276), .ZN(n5477) );
  INV_X4 U4824 ( .A(n4817), .ZN(n4818) );
  NOR2_X1 U4825 ( .A1(net63523), .A2(n6133), .ZN(N833) );
  NAND3_X2 U4826 ( .A1(n6134), .A2(n6133), .A3(n6132), .ZN(n5900) );
  INV_X4 U4827 ( .A(n4732), .ZN(n4733) );
  INV_X8 U4828 ( .A(n4541), .ZN(n4764) );
  NAND2_X1 U4829 ( .A1(n4837), .A2(n4396), .ZN(n6742) );
  NOR2_X1 U4830 ( .A1(net63523), .A2(n6121), .ZN(N821) );
  NOR2_X2 U4831 ( .A1(net63527), .A2(n6119), .ZN(N819) );
  OAI221_X2 U4832 ( .B1(net63551), .B2(n2533), .C1(n4735), .C2(net63575), .A(
        net63579), .ZN(n4734) );
  INV_X2 U4833 ( .A(n2533), .ZN(u4_fract_out_27_) );
  AOI22_X4 U4834 ( .A1(u4_N5987), .A2(net63317), .B1(u4_N6095), .B2(net63335), 
        .ZN(n2533) );
  NOR3_X1 U4835 ( .A1(n4823), .A2(n4837), .A3(n4840), .ZN(n4736) );
  INV_X4 U4836 ( .A(n4737), .ZN(n4738) );
  NOR2_X2 U4837 ( .A1(remainder[35]), .A2(remainder[34]), .ZN(n5741) );
  NAND3_X2 U4838 ( .A1(n6945), .A2(n6892), .A3(n6891), .ZN(n6967) );
  INV_X2 U4839 ( .A(n4739), .ZN(n4740) );
  INV_X4 U4840 ( .A(n4741), .ZN(n4742) );
  NOR3_X1 U4841 ( .A1(u6_N19), .A2(u6_N1), .A3(u6_N18), .ZN(n6852) );
  INV_X1 U4842 ( .A(u6_N19), .ZN(n7094) );
  INV_X4 U4843 ( .A(n4743), .ZN(n4744) );
  INV_X4 U4844 ( .A(n4745), .ZN(n4746) );
  INV_X2 U4845 ( .A(n4747), .ZN(n4748) );
  INV_X4 U4846 ( .A(n4751), .ZN(n4752) );
  INV_X4 U4847 ( .A(n4753), .ZN(n4754) );
  INV_X4 U4848 ( .A(n4755), .ZN(n4756) );
  INV_X4 U4849 ( .A(n4757), .ZN(n4758) );
  INV_X4 U4850 ( .A(n4759), .ZN(n4760) );
  INV_X4 U4851 ( .A(n4761), .ZN(n4762) );
  INV_X4 U4852 ( .A(n4800), .ZN(n4809) );
  NOR2_X2 U4853 ( .A1(remainder[32]), .A2(remainder[31]), .ZN(n5742) );
  NOR4_X1 U4854 ( .A1(n3100), .A2(u6_N22), .A3(u6_N21), .A4(u6_N20), .ZN(n6460) );
  NAND3_X2 U4855 ( .A1(n6946), .A2(n6986), .A3(n6885), .ZN(n6886) );
  INV_X4 U4856 ( .A(n7020), .ZN(n4765) );
  INV_X4 U4857 ( .A(n4778), .ZN(n4790) );
  INV_X1 U4858 ( .A(u6_N31), .ZN(n7058) );
  INV_X4 U4859 ( .A(n4767), .ZN(n4768) );
  OR4_X4 U4860 ( .A1(u6_N31), .A2(u6_N30), .A3(u6_N2), .A4(u6_N29), .ZN(n3107)
         );
  INV_X2 U4861 ( .A(u6_N46), .ZN(n7014) );
  INV_X8 U4862 ( .A(n4781), .ZN(n6837) );
  INV_X8 U4863 ( .A(n4769), .ZN(n4772) );
  INV_X1 U4864 ( .A(u6_N27), .ZN(n7070) );
  INV_X1 U4865 ( .A(n4772), .ZN(n7029) );
  INV_X8 U4866 ( .A(n4816), .ZN(n4822) );
  INV_X4 U4867 ( .A(n4787), .ZN(n7026) );
  INV_X2 U4868 ( .A(u6_N24), .ZN(n7079) );
  NOR2_X2 U4869 ( .A1(remainder[37]), .A2(remainder[36]), .ZN(n5740) );
  OR4_X1 U4870 ( .A1(u6_N45), .A2(u6_N46), .A3(n4765), .A4(n3111), .ZN(n3108)
         );
  OR4_X1 U4871 ( .A1(u6_N40), .A2(n4772), .A3(n4787), .A4(u6_N43), .ZN(n3112)
         );
  INV_X8 U4872 ( .A(n4771), .ZN(n4786) );
  INV_X1 U4873 ( .A(u6_N36), .ZN(n7044) );
  INV_X4 U4874 ( .A(n4774), .ZN(n4775) );
  INV_X1 U4875 ( .A(u6_N43), .ZN(n7023) );
  NOR2_X1 U4876 ( .A1(net63523), .A2(n6136), .ZN(N836) );
  INV_X2 U4877 ( .A(n6053), .ZN(n6056) );
  NOR3_X4 U4878 ( .A1(n5922), .A2(net58886), .A3(n6053), .ZN(net58825) );
  NAND3_X2 U4879 ( .A1(n6137), .A2(n6136), .A3(n6135), .ZN(n5899) );
  OAI21_X2 U4880 ( .B1(n4282), .B2(net58982), .A(net58976), .ZN(net58425) );
  OAI21_X2 U4881 ( .B1(n4281), .B2(net58985), .A(net58976), .ZN(net58422) );
  OAI21_X2 U4882 ( .B1(n4282), .B2(net58981), .A(net58976), .ZN(net58423) );
  OAI21_X2 U4883 ( .B1(net58974), .B2(net58983), .A(net58976), .ZN(net58421)
         );
  AOI22_X1 U4884 ( .A1(net59166), .A2(net59099), .B1(net87237), .B2(net59159), 
        .ZN(n5836) );
  INV_X8 U4885 ( .A(u4_exp_out_10_), .ZN(net45067) );
  AOI22_X1 U4886 ( .A1(u4_exp_in_pl1_6_), .A2(net59568), .B1(n4276), .B2(
        net59578), .ZN(n5637) );
  NAND2_X1 U4887 ( .A1(u4_exp_in_pl1_5_), .A2(net59568), .ZN(n5643) );
  NAND2_X1 U4888 ( .A1(u4_exp_in_pl1_4_), .A2(net59568), .ZN(n5649) );
  NAND2_X1 U4889 ( .A1(u4_exp_in_pl1_3_), .A2(net59568), .ZN(n5658) );
  NAND2_X1 U4890 ( .A1(u4_exp_in_pl1_2_), .A2(net59568), .ZN(n5666) );
  NOR2_X1 U4891 ( .A1(net60316), .A2(n4533), .ZN(n5331) );
  NAND3_X1 U4892 ( .A1(net33563), .A2(n4694), .A3(n4509), .ZN(n5378) );
  NAND3_X1 U4893 ( .A1(net60096), .A2(net33565), .A3(n4509), .ZN(n5403) );
  NOR2_X1 U4894 ( .A1(fract_denorm[57]), .A2(n4533), .ZN(n5441) );
  NAND3_X1 U4895 ( .A1(n4509), .A2(n8521), .A3(net60117), .ZN(n5402) );
  INV_X4 U4896 ( .A(n4776), .ZN(n4777) );
  INV_X1 U4897 ( .A(u6_N39), .ZN(n7035) );
  INV_X4 U4898 ( .A(n4779), .ZN(n4780) );
  INV_X1 U4899 ( .A(u6_N30), .ZN(n7061) );
  NOR3_X1 U4900 ( .A1(u6_N23), .A2(u6_N25), .A3(u6_N24), .ZN(n3106) );
  NOR3_X1 U4901 ( .A1(u6_N24), .A2(u6_N2), .A3(u6_N23), .ZN(n6850) );
  INV_X1 U4902 ( .A(u6_N40), .ZN(n7032) );
  OR4_X1 U4903 ( .A1(u6_N27), .A2(n4764), .A3(u6_N26), .A4(n3107), .ZN(n3100)
         );
  NOR2_X1 U4904 ( .A1(net63523), .A2(n6139), .ZN(N839) );
  NOR3_X4 U4905 ( .A1(n5898), .A2(n5897), .A3(n5896), .ZN(n5921) );
  NAND3_X2 U4906 ( .A1(n6140), .A2(n6139), .A3(n6138), .ZN(n5898) );
  NOR2_X1 U4907 ( .A1(u4_fi_ldz_1_), .A2(net87917), .ZN(n5475) );
  NOR3_X1 U4908 ( .A1(net59990), .A2(net59991), .A3(n4521), .ZN(n5435) );
  NAND3_X2 U4909 ( .A1(n6124), .A2(n6123), .A3(n6122), .ZN(n5916) );
  NOR2_X2 U4910 ( .A1(net63523), .A2(n6122), .ZN(N822) );
  INV_X1 U4911 ( .A(u6_N29), .ZN(n7064) );
  INV_X4 U4912 ( .A(n4782), .ZN(n4783) );
  INV_X1 U4913 ( .A(u6_N37), .ZN(n7041) );
  INV_X4 U4914 ( .A(n4784), .ZN(n4785) );
  NAND3_X2 U4915 ( .A1(n6127), .A2(n6126), .A3(n6125), .ZN(n5915) );
  INV_X1 U4916 ( .A(n4786), .ZN(n7049) );
  INV_X2 U4917 ( .A(u6_N33), .ZN(n7052) );
  OR3_X1 U4918 ( .A1(u6_N36), .A2(u6_N37), .A3(u6_N35), .ZN(n3113) );
  NOR4_X1 U4919 ( .A1(n3113), .A2(u6_N32), .A3(n4786), .A4(u6_N33), .ZN(n3096)
         );
  INV_X1 U4920 ( .A(u6_N45), .ZN(n7017) );
  INV_X1 U4921 ( .A(n4791), .ZN(n7038) );
  INV_X8 U4922 ( .A(n4788), .ZN(n4791) );
  INV_X4 U4923 ( .A(n4792), .ZN(n4793) );
  NOR4_X1 U4924 ( .A1(n3112), .A2(n4791), .A3(u6_N3), .A4(u6_N39), .ZN(n3097)
         );
  INV_X4 U4925 ( .A(n6837), .ZN(n4799) );
  NAND2_X4 U4926 ( .A1(n4805), .A2(n4919), .ZN(u6_N52) );
  INV_X4 U4927 ( .A(n4801), .ZN(n4802) );
  INV_X1 U4928 ( .A(n4270), .ZN(n4803) );
  INV_X2 U4929 ( .A(n4803), .ZN(n4804) );
  INV_X4 U4930 ( .A(n4833), .ZN(n4840) );
  NOR3_X4 U4931 ( .A1(n4806), .A2(n4808), .A3(n4807), .ZN(n4805) );
  NAND3_X2 U4932 ( .A1(n4826), .A2(n4821), .A3(n4827), .ZN(n4806) );
  NAND2_X2 U4933 ( .A1(n4828), .A2(n4829), .ZN(n4807) );
  NAND3_X2 U4934 ( .A1(n4830), .A2(n4831), .A3(n4832), .ZN(n4808) );
  INV_X1 U4935 ( .A(n4809), .ZN(n7011) );
  NOR2_X1 U4936 ( .A1(fracta_mul[2]), .A2(n5040), .ZN(n4944) );
  INV_X2 U4937 ( .A(fracta_mul[2]), .ZN(n6835) );
  NOR3_X1 U4938 ( .A1(fracta_mul[24]), .A2(fracta_mul[2]), .A3(fracta_mul[23]), 
        .ZN(n6849) );
  NAND2_X1 U4939 ( .A1(n4395), .A2(n4840), .ZN(n6720) );
  NOR2_X1 U4940 ( .A1(n4840), .A2(n4395), .ZN(n6724) );
  OR3_X1 U4941 ( .A1(n4424), .A2(u6_N49), .A3(u6_N48), .ZN(n3111) );
  INV_X1 U4942 ( .A(u6_N48), .ZN(n7008) );
  INV_X4 U4943 ( .A(n4810), .ZN(n4811) );
  INV_X4 U4944 ( .A(n4814), .ZN(n4815) );
  INV_X1 U4945 ( .A(fracta_mul[0]), .ZN(n6839) );
  NOR3_X1 U4946 ( .A1(fracta_mul[22]), .A2(fracta_mul[0]), .A3(fracta_mul[21]), 
        .ZN(n6449) );
  INV_X1 U4947 ( .A(u6_N51), .ZN(n6999) );
  NOR2_X1 U4948 ( .A1(u6_N51), .A2(n4473), .ZN(u0_N5) );
  INV_X4 U4949 ( .A(n4819), .ZN(n4820) );
  INV_X16 U4950 ( .A(net63553), .ZN(net63543) );
  INV_X16 U4951 ( .A(net63571), .ZN(net63561) );
  INV_X4 U4952 ( .A(n4824), .ZN(n4823) );
  NOR3_X1 U4953 ( .A1(fracta_mul[2]), .A2(n4799), .A3(n5040), .ZN(n6439) );
  OAI21_X1 U4954 ( .B1(fracta_mul[2]), .B2(n4799), .A(n5041), .ZN(n5042) );
  NOR3_X1 U4955 ( .A1(fracta_mul[19]), .A2(fracta_mul[18]), .A3(n4770), .ZN(
        n6851) );
  INV_X4 U4956 ( .A(n4835), .ZN(n4836) );
  INV_X1 U4957 ( .A(n4840), .ZN(n6757) );
  INV_X2 U4958 ( .A(opb_r[53]), .ZN(n7148) );
  NAND2_X1 U4959 ( .A1(opb_r[53]), .A2(n4392), .ZN(n6739) );
  OAI22_X1 U4960 ( .A1(opb_r[52]), .A2(n4330), .B1(opb_r[53]), .B2(n4392), 
        .ZN(n6714) );
  NOR2_X1 U4961 ( .A1(opb_r[60]), .A2(n4394), .ZN(n6729) );
  NAND2_X1 U4962 ( .A1(opb_r[60]), .A2(n4394), .ZN(n6726) );
  INV_X2 U4963 ( .A(opb_r[54]), .ZN(n7149) );
  NOR2_X1 U4964 ( .A1(opb_r[54]), .A2(n4331), .ZN(n6713) );
  NAND2_X1 U4965 ( .A1(opb_r[54]), .A2(n4331), .ZN(n6740) );
  INV_X4 U4966 ( .A(opb_r[57]), .ZN(n4838) );
  INV_X8 U4967 ( .A(n4838), .ZN(n4839) );
  NOR3_X4 U4968 ( .A1(n4823), .A2(n4837), .A3(n4840), .ZN(n4919) );
  OAI221_X1 U4969 ( .B1(n4309), .B2(n4346), .C1(n6466), .C2(n6465), .A(n6464), 
        .ZN(u2_underflow_d[1]) );
  NAND4_X1 U4970 ( .A1(n7152), .A2(n4836), .A3(n7151), .A4(n7150), .ZN(n3074)
         );
  NOR2_X1 U4971 ( .A1(n4836), .A2(n4332), .ZN(n6718) );
  NAND2_X1 U4972 ( .A1(n4836), .A2(n4332), .ZN(n6743) );
  NOR2_X1 U4973 ( .A1(n4853), .A2(opb_r[62]), .ZN(n6466) );
  NAND3_X1 U4974 ( .A1(opb_r[61]), .A2(opb_r[62]), .A3(opb_r[60]), .ZN(n3078)
         );
  NOR2_X1 U4975 ( .A1(opb_r[62]), .A2(n4854), .ZN(n6284) );
  NAND3_X1 U4976 ( .A1(n4425), .A2(n4839), .A3(n4271), .ZN(n7146) );
  NOR2_X1 U4977 ( .A1(n4853), .A2(n4309), .ZN(n6471) );
  NAND2_X1 U4978 ( .A1(u2_N157), .A2(n4309), .ZN(n6916) );
  INV_X8 U4979 ( .A(n4293), .ZN(net66904) );
  INV_X8 U4980 ( .A(n4293), .ZN(net66905) );
  INV_X8 U4981 ( .A(n4293), .ZN(net66906) );
  INV_X8 U4982 ( .A(n4293), .ZN(net66907) );
  INV_X32 U4983 ( .A(n7189), .ZN(n4842) );
  INV_X32 U4984 ( .A(n4842), .ZN(n4843) );
  NAND2_X4 U4985 ( .A1(net59674), .A2(net63293), .ZN(net57241) );
  NAND2_X4 U4986 ( .A1(net59207), .A2(n5818), .ZN(net59087) );
  NAND2_X4 U4987 ( .A1(n5818), .A2(net58676), .ZN(net59081) );
  INV_X8 U4988 ( .A(n6751), .ZN(n6765) );
  INV_X32 U4989 ( .A(net66870), .ZN(net66871) );
  INV_X32 U4990 ( .A(n4847), .ZN(n4848) );
  INV_X32 U4991 ( .A(n4849), .ZN(n4850) );
  OR2_X4 U4992 ( .A1(n4298), .A2(fpu_op_r2[2]), .ZN(n3296) );
  INV_X32 U4993 ( .A(net63583), .ZN(net63577) );
  INV_X32 U4994 ( .A(net63583), .ZN(net63579) );
  INV_X32 U4995 ( .A(net63553), .ZN(net63541) );
  INV_X32 U4996 ( .A(net63551), .ZN(net63545) );
  INV_X32 U4997 ( .A(net63551), .ZN(net63547) );
  INV_X32 U4998 ( .A(net63555), .ZN(net63551) );
  INV_X32 U4999 ( .A(n6409), .ZN(n4854) );
  INV_X32 U5000 ( .A(n4868), .ZN(n4867) );
  INV_X32 U5001 ( .A(n4875), .ZN(n4869) );
  INV_X32 U5002 ( .A(n4875), .ZN(n4870) );
  INV_X32 U5003 ( .A(n4874), .ZN(n4871) );
  INV_X32 U5004 ( .A(n4874), .ZN(n4872) );
  INV_X32 U5005 ( .A(n4874), .ZN(n4873) );
  INV_X32 U5006 ( .A(n4867), .ZN(n4874) );
  INV_X32 U5007 ( .A(n4867), .ZN(n4875) );
  INV_X32 U5008 ( .A(n4878), .ZN(n4877) );
  INV_X32 U5009 ( .A(n4896), .ZN(n4881) );
  INV_X32 U5010 ( .A(n4896), .ZN(n4882) );
  INV_X32 U5011 ( .A(n4896), .ZN(n4883) );
  INV_X32 U5012 ( .A(n4895), .ZN(n4884) );
  INV_X32 U5013 ( .A(n4895), .ZN(n4885) );
  INV_X32 U5014 ( .A(n4894), .ZN(n4887) );
  INV_X32 U5015 ( .A(n4894), .ZN(n4888) );
  INV_X32 U5016 ( .A(n4894), .ZN(n4889) );
  INV_X32 U5017 ( .A(n4893), .ZN(n4890) );
  INV_X32 U5018 ( .A(n4893), .ZN(n4891) );
  INV_X32 U5019 ( .A(n4876), .ZN(n4893) );
  INV_X32 U5020 ( .A(n4877), .ZN(n4895) );
  INV_X32 U5021 ( .A(n4877), .ZN(n4896) );
  INV_X32 U5022 ( .A(n4877), .ZN(n4897) );
  INV_X32 U5023 ( .A(net63347), .ZN(net63335) );
  INV_X32 U5024 ( .A(net63329), .ZN(net63317) );
  INV_X32 U5025 ( .A(net63329), .ZN(net63319) );
  INV_X32 U5026 ( .A(net63327), .ZN(net63323) );
  INV_X32 U5027 ( .A(net63331), .ZN(net63329) );
  INV_X32 U5028 ( .A(net63333), .ZN(net63331) );
  INV_X32 U5029 ( .A(n4906), .ZN(n4905) );
  INV_X32 U5030 ( .A(n4915), .ZN(n4907) );
  INV_X32 U5031 ( .A(n4915), .ZN(n4908) );
  INV_X32 U5032 ( .A(n4915), .ZN(n4909) );
  INV_X32 U5033 ( .A(n4915), .ZN(n4910) );
  INV_X32 U5034 ( .A(n4915), .ZN(n4911) );
  INV_X32 U5035 ( .A(n4915), .ZN(n4912) );
  INV_X32 U5036 ( .A(n4915), .ZN(n4913) );
  INV_X32 U5037 ( .A(n4915), .ZN(n4914) );
  INV_X32 U5038 ( .A(n4904), .ZN(n4915) );
  INV_X32 U5039 ( .A(net63089), .ZN(net63079) );
  NOR3_X4 U5040 ( .A1(opa_r[55]), .A2(opa_r[58]), .A3(opa_r[60]), .ZN(n4923)
         );
  NOR3_X4 U5041 ( .A1(opa_r[56]), .A2(opa_r[54]), .A3(opa_r[53]), .ZN(n4922)
         );
  NOR3_X4 U5042 ( .A1(opa_r[61]), .A2(opa_r[59]), .A3(opa_r[57]), .ZN(n4921)
         );
  NOR2_X4 U5043 ( .A1(opa_r[52]), .A2(n4853), .ZN(n4920) );
  NAND4_X2 U5044 ( .A1(n4923), .A2(n4922), .A3(n4921), .A4(n4920), .ZN(u2_N157) );
  NAND2_X2 U5045 ( .A1(n4314), .A2(n4338), .ZN(n5049) );
  INV_X4 U5046 ( .A(n5049), .ZN(n4924) );
  NAND2_X2 U5047 ( .A1(n4301), .A2(n4291), .ZN(n6450) );
  INV_X4 U5048 ( .A(n6450), .ZN(n5054) );
  NAND2_X2 U5049 ( .A1(n5054), .A2(n4297), .ZN(n5013) );
  INV_X4 U5050 ( .A(n5013), .ZN(n4925) );
  NAND2_X2 U5051 ( .A1(n4925), .A2(n4303), .ZN(n4926) );
  INV_X4 U5052 ( .A(n4926), .ZN(n5019) );
  NAND2_X2 U5053 ( .A1(n5019), .A2(n4302), .ZN(n5055) );
  INV_X4 U5054 ( .A(n5055), .ZN(n4927) );
  INV_X4 U5055 ( .A(n4999), .ZN(n4996) );
  NAND2_X2 U5056 ( .A1(n4436), .A2(n4296), .ZN(n4928) );
  INV_X4 U5057 ( .A(n4928), .ZN(n5010) );
  INV_X4 U5058 ( .A(n6441), .ZN(n4929) );
  INV_X4 U5059 ( .A(n4982), .ZN(n4930) );
  NAND2_X2 U5060 ( .A1(n4930), .A2(n4335), .ZN(n4988) );
  INV_X4 U5061 ( .A(n4988), .ZN(n4959) );
  NAND3_X4 U5062 ( .A1(n4959), .A2(n4340), .A3(n4310), .ZN(n5048) );
  NOR2_X4 U5063 ( .A1(n6442), .A2(n5048), .ZN(n4931) );
  NAND2_X2 U5064 ( .A1(n4931), .A2(n4423), .ZN(n4970) );
  INV_X4 U5065 ( .A(n4970), .ZN(n4961) );
  NAND2_X2 U5066 ( .A1(n5033), .A2(n4489), .ZN(n5023) );
  NAND2_X2 U5067 ( .A1(n4933), .A2(n4932), .ZN(n5020) );
  INV_X4 U5068 ( .A(n5020), .ZN(n4934) );
  NAND2_X2 U5069 ( .A1(n4934), .A2(n4339), .ZN(n4935) );
  INV_X4 U5070 ( .A(n4935), .ZN(n5039) );
  NAND2_X2 U5071 ( .A1(n4434), .A2(n4336), .ZN(n6859) );
  INV_X4 U5072 ( .A(n6859), .ZN(n4967) );
  NAND3_X4 U5073 ( .A1(n5039), .A2(n4967), .A3(n4315), .ZN(n5067) );
  NAND2_X2 U5074 ( .A1(n4337), .A2(n4312), .ZN(n4997) );
  NOR2_X4 U5075 ( .A1(n5067), .A2(n4997), .ZN(n4936) );
  INV_X4 U5076 ( .A(n4979), .ZN(n4937) );
  NAND2_X2 U5077 ( .A1(n4937), .A2(n4432), .ZN(n4942) );
  NOR2_X4 U5078 ( .A1(fracta_mul[30]), .A2(fracta_mul[29]), .ZN(n4971) );
  NAND3_X4 U5079 ( .A1(n4961), .A2(n4418), .A3(n4971), .ZN(n4954) );
  INV_X4 U5080 ( .A(n4954), .ZN(n4940) );
  NAND2_X2 U5081 ( .A1(n4939), .A2(n4938), .ZN(n4953) );
  INV_X4 U5082 ( .A(n4953), .ZN(n6444) );
  INV_X4 U5083 ( .A(n4941), .ZN(n4951) );
  NAND3_X4 U5084 ( .A1(n4951), .A2(n4299), .A3(n4289), .ZN(n5068) );
  INV_X4 U5085 ( .A(n4942), .ZN(n4990) );
  NAND2_X2 U5086 ( .A1(n4945), .A2(n4944), .ZN(n4949) );
  NOR2_X4 U5087 ( .A1(n4954), .A2(n4426), .ZN(n4976) );
  NOR2_X4 U5088 ( .A1(n4947), .A2(n4976), .ZN(n4948) );
  NAND3_X4 U5089 ( .A1(n4950), .A2(n4949), .A3(n4948), .ZN(n5074) );
  NOR2_X4 U5090 ( .A1(n5023), .A2(n5074), .ZN(n4966) );
  INV_X4 U5091 ( .A(n4992), .ZN(n4958) );
  NOR2_X4 U5092 ( .A1(fracta_mul[27]), .A2(n4954), .ZN(n4955) );
  NAND2_X2 U5093 ( .A1(fracta_mul[26]), .A2(n4955), .ZN(n4952) );
  NAND2_X2 U5094 ( .A1(fracta_mul[22]), .A2(n4951), .ZN(n5003) );
  NAND3_X4 U5095 ( .A1(n4952), .A2(n5069), .A3(n5003), .ZN(n5061) );
  INV_X4 U5096 ( .A(n5061), .ZN(n4957) );
  INV_X4 U5097 ( .A(n5017), .ZN(n4956) );
  NAND3_X4 U5098 ( .A1(n4957), .A2(n4956), .A3(n5012), .ZN(n4983) );
  NOR2_X4 U5099 ( .A1(n4958), .A2(n4983), .ZN(n4965) );
  NAND2_X2 U5100 ( .A1(fracta_mul[30]), .A2(n4961), .ZN(n5053) );
  INV_X4 U5101 ( .A(n5053), .ZN(n5029) );
  NOR3_X4 U5102 ( .A1(n4963), .A2(n4962), .A3(n5029), .ZN(n4964) );
  NAND3_X4 U5103 ( .A1(n4966), .A2(n4965), .A3(n4964), .ZN(div_opa_ldz_d[4])
         );
  INV_X4 U5104 ( .A(n5068), .ZN(n4977) );
  INV_X4 U5105 ( .A(n4970), .ZN(n4972) );
  NAND2_X2 U5106 ( .A1(n4974), .A2(n4973), .ZN(n4975) );
  NAND2_X2 U5107 ( .A1(fracta_mul[42]), .A2(n4996), .ZN(n5046) );
  INV_X4 U5108 ( .A(n5068), .ZN(n4980) );
  OAI21_X4 U5109 ( .B1(n4982), .B2(n4335), .A(n4981), .ZN(n5060) );
  INV_X4 U5110 ( .A(n4997), .ZN(n5006) );
  NAND2_X2 U5111 ( .A1(fracta_mul[7]), .A2(n5006), .ZN(n4984) );
  NOR2_X4 U5112 ( .A1(n5067), .A2(n4984), .ZN(n4987) );
  NAND2_X2 U5113 ( .A1(n4993), .A2(n4992), .ZN(n5059) );
  INV_X4 U5114 ( .A(n5059), .ZN(n4994) );
  NAND2_X2 U5115 ( .A1(n4995), .A2(n4994), .ZN(n5024) );
  OAI211_X2 U5116 ( .C1(n4999), .C2(n4296), .A(n5034), .B(n5035), .ZN(n5065)
         );
  NAND4_X2 U5117 ( .A1(n5002), .A2(n5046), .A3(n5001), .A4(n5000), .ZN(
        div_opa_ldz_d[3]) );
  INV_X4 U5118 ( .A(n5003), .ZN(n5004) );
  INV_X4 U5119 ( .A(n5068), .ZN(n5016) );
  NAND4_X2 U5120 ( .A1(fracta_mul[8]), .A2(n5006), .A3(n4433), .A4(n5038), 
        .ZN(n5008) );
  NAND2_X2 U5121 ( .A1(n4443), .A2(n5010), .ZN(n5011) );
  OAI221_X2 U5122 ( .B1(n5013), .B2(n4303), .C1(fracta_mul[26]), .C2(n5012), 
        .A(n5011), .ZN(n5014) );
  INV_X4 U5123 ( .A(n5023), .ZN(n5026) );
  INV_X4 U5124 ( .A(n5024), .ZN(n5025) );
  NAND4_X2 U5125 ( .A1(n5028), .A2(n5027), .A3(n5026), .A4(n5025), .ZN(n5073)
         );
  NAND2_X2 U5126 ( .A1(n5034), .A2(n5033), .ZN(n5037) );
  INV_X4 U5127 ( .A(n5035), .ZN(n5036) );
  NOR2_X4 U5128 ( .A1(n5037), .A2(n5036), .ZN(n5064) );
  NAND2_X2 U5129 ( .A1(n5039), .A2(n6859), .ZN(n5043) );
  INV_X4 U5130 ( .A(n5040), .ZN(n5041) );
  NAND4_X2 U5131 ( .A1(n5045), .A2(n5044), .A3(n5043), .A4(n5042), .ZN(n5058)
         );
  INV_X4 U5132 ( .A(n5046), .ZN(n5047) );
  NAND2_X2 U5133 ( .A1(n5047), .A2(n4296), .ZN(n5052) );
  INV_X4 U5134 ( .A(n5048), .ZN(n5050) );
  NAND3_X4 U5135 ( .A1(n5053), .A2(n5052), .A3(n5051), .ZN(n5057) );
  OAI22_X2 U5136 ( .A1(n4316), .A2(n5055), .B1(fracta_mul[51]), .B2(n5054), 
        .ZN(n5056) );
  AOI211_X4 U5137 ( .C1(n5016), .C2(n5058), .A(n5057), .B(n5056), .ZN(n5063)
         );
  NOR3_X4 U5138 ( .A1(n5061), .A2(n5060), .A3(n5059), .ZN(n5062) );
  NAND3_X4 U5139 ( .A1(n5064), .A2(n5063), .A3(n5062), .ZN(div_opa_ldz_d[1])
         );
  NOR2_X4 U5140 ( .A1(fracta_mul[51]), .A2(n5065), .ZN(n5077) );
  NAND2_X2 U5141 ( .A1(fracta_mul[17]), .A2(n4427), .ZN(n5066) );
  OAI211_X2 U5142 ( .C1(n5067), .C2(n4312), .A(n5066), .B(n4438), .ZN(n5072)
         );
  INV_X4 U5143 ( .A(n5069), .ZN(n5070) );
  AOI211_X4 U5144 ( .C1(n5072), .C2(n4977), .A(n5071), .B(n5070), .ZN(n5076)
         );
  NOR2_X4 U5145 ( .A1(n5074), .A2(n5073), .ZN(n5075) );
  NAND3_X4 U5146 ( .A1(n5077), .A2(n5076), .A3(n5075), .ZN(div_opa_ldz_d[0])
         );
  INV_X4 U5147 ( .A(N308), .ZN(n5078) );
  NAND2_X2 U5148 ( .A1(n5078), .A2(n4900), .ZN(u6_N107) );
  AOI22_X2 U5149 ( .A1(fract_i2f[73]), .A2(net63079), .B1(prod[73]), .B2(
        net66929), .ZN(n5081) );
  NAND2_X2 U5150 ( .A1(quo[75]), .A2(net66905), .ZN(n5080) );
  AOI22_X2 U5151 ( .A1(fract_out_q[24]), .A2(net63503), .B1(quo[23]), .B2(
        net66896), .ZN(n5079) );
  NAND3_X4 U5152 ( .A1(n5081), .A2(n5080), .A3(n5079), .ZN(fract_denorm[73])
         );
  AOI22_X2 U5153 ( .A1(fract_i2f[71]), .A2(n4294), .B1(prod[71]), .B2(net66930), .ZN(n5084) );
  NAND2_X2 U5154 ( .A1(quo[73]), .A2(net66906), .ZN(n5083) );
  AOI22_X2 U5155 ( .A1(fract_out_q[22]), .A2(net63511), .B1(quo[21]), .B2(
        net66895), .ZN(n5082) );
  NAND3_X4 U5156 ( .A1(n5084), .A2(n5083), .A3(n5082), .ZN(fract_denorm[71])
         );
  AOI22_X2 U5157 ( .A1(fract_i2f[72]), .A2(net63083), .B1(prod[72]), .B2(
        net66929), .ZN(n5087) );
  NAND2_X2 U5158 ( .A1(quo[74]), .A2(net66907), .ZN(n5086) );
  AOI22_X2 U5159 ( .A1(fract_out_q[23]), .A2(net63513), .B1(quo[22]), .B2(
        net66897), .ZN(n5085) );
  NAND3_X4 U5160 ( .A1(n5087), .A2(n5086), .A3(n5085), .ZN(fract_denorm[72])
         );
  AOI22_X2 U5161 ( .A1(fract_i2f[69]), .A2(net63083), .B1(prod[69]), .B2(
        net66930), .ZN(n5090) );
  NAND2_X2 U5162 ( .A1(quo[71]), .A2(net66910), .ZN(n5089) );
  AOI22_X2 U5163 ( .A1(fract_out_q[20]), .A2(net63511), .B1(quo[19]), .B2(
        net66897), .ZN(n5088) );
  NAND3_X4 U5164 ( .A1(n5090), .A2(n5089), .A3(n5088), .ZN(fract_denorm[69])
         );
  AOI22_X2 U5165 ( .A1(fract_i2f[70]), .A2(net63083), .B1(prod[70]), .B2(
        net66928), .ZN(n5093) );
  NAND2_X2 U5166 ( .A1(quo[72]), .A2(net66904), .ZN(n5092) );
  AOI22_X2 U5167 ( .A1(fract_out_q[21]), .A2(net63511), .B1(net66896), .B2(
        quo[20]), .ZN(n5091) );
  NAND3_X4 U5168 ( .A1(n5093), .A2(n5092), .A3(n5091), .ZN(fract_denorm[70])
         );
  AOI22_X2 U5169 ( .A1(fract_i2f[80]), .A2(net63083), .B1(prod[80]), .B2(
        net66929), .ZN(n5096) );
  NAND2_X2 U5170 ( .A1(quo[82]), .A2(net66910), .ZN(n5095) );
  AOI22_X2 U5171 ( .A1(fract_out_q[31]), .A2(net63509), .B1(quo[30]), .B2(
        net66895), .ZN(n5094) );
  NAND3_X4 U5172 ( .A1(n5096), .A2(n5095), .A3(n5094), .ZN(fract_denorm[80])
         );
  AOI22_X2 U5173 ( .A1(fract_i2f[81]), .A2(net63083), .B1(prod[81]), .B2(
        net66930), .ZN(n5099) );
  NAND2_X2 U5174 ( .A1(quo[83]), .A2(net66911), .ZN(n5098) );
  AOI22_X2 U5175 ( .A1(fract_out_q[32]), .A2(net63509), .B1(quo[31]), .B2(
        net66897), .ZN(n5097) );
  NAND3_X4 U5176 ( .A1(n5099), .A2(n5098), .A3(n5097), .ZN(fract_denorm[81])
         );
  AOI22_X2 U5177 ( .A1(fract_i2f[77]), .A2(net63083), .B1(prod[77]), .B2(
        net66928), .ZN(n5102) );
  NAND2_X2 U5178 ( .A1(quo[79]), .A2(net66912), .ZN(n5101) );
  AOI22_X2 U5179 ( .A1(fract_out_q[28]), .A2(net63509), .B1(quo[27]), .B2(
        net66896), .ZN(n5100) );
  AOI22_X2 U5180 ( .A1(fract_i2f[78]), .A2(net63083), .B1(prod[78]), .B2(
        net66929), .ZN(n5105) );
  NAND2_X2 U5181 ( .A1(quo[80]), .A2(net66906), .ZN(n5104) );
  AOI22_X2 U5182 ( .A1(fract_out_q[29]), .A2(net63511), .B1(net66896), .B2(
        quo[28]), .ZN(n5103) );
  NAND3_X4 U5183 ( .A1(n5105), .A2(n5104), .A3(n5103), .ZN(fract_denorm[78])
         );
  AOI22_X2 U5184 ( .A1(fract_i2f[79]), .A2(net63083), .B1(prod[79]), .B2(
        net66930), .ZN(n5108) );
  NAND2_X2 U5185 ( .A1(quo[81]), .A2(net66914), .ZN(n5107) );
  AOI22_X2 U5186 ( .A1(fract_out_q[30]), .A2(net63509), .B1(quo[29]), .B2(
        net66895), .ZN(n5106) );
  AOI22_X2 U5187 ( .A1(fract_i2f[76]), .A2(net63083), .B1(prod[76]), .B2(
        net66928), .ZN(net60652) );
  NAND2_X2 U5188 ( .A1(quo[78]), .A2(net66910), .ZN(net60653) );
  NAND2_X2 U5189 ( .A1(prod[105]), .A2(net58645), .ZN(net60646) );
  NAND2_X2 U5190 ( .A1(fract_out_q[56]), .A2(net63513), .ZN(net60647) );
  AOI22_X2 U5191 ( .A1(fract_i2f[104]), .A2(n4294), .B1(prod[104]), .B2(
        net66929), .ZN(n5111) );
  NAND2_X2 U5192 ( .A1(quo[106]), .A2(net66911), .ZN(n5110) );
  NAND3_X4 U5193 ( .A1(n5111), .A2(n5110), .A3(n5109), .ZN(fract_denorm[104])
         );
  AOI22_X2 U5194 ( .A1(fract_i2f[103]), .A2(net63085), .B1(prod[103]), .B2(
        net66930), .ZN(n5114) );
  NAND2_X2 U5195 ( .A1(quo[105]), .A2(net66912), .ZN(n5113) );
  NAND3_X4 U5196 ( .A1(n5114), .A2(n5113), .A3(n5112), .ZN(fract_denorm[103])
         );
  AOI22_X2 U5197 ( .A1(fract_i2f[100]), .A2(n4294), .B1(prod[100]), .B2(
        net66928), .ZN(n5117) );
  NAND2_X2 U5198 ( .A1(quo[102]), .A2(net66912), .ZN(n5116) );
  NAND3_X4 U5199 ( .A1(n5117), .A2(n5116), .A3(n5115), .ZN(fract_denorm[100])
         );
  AOI22_X2 U5200 ( .A1(fract_i2f[101]), .A2(n4294), .B1(prod[101]), .B2(
        net66929), .ZN(n5120) );
  NAND2_X2 U5201 ( .A1(quo[103]), .A2(net66905), .ZN(n5119) );
  NAND3_X4 U5202 ( .A1(n5120), .A2(n5119), .A3(n5118), .ZN(fract_denorm[101])
         );
  AOI22_X2 U5203 ( .A1(fract_i2f[102]), .A2(net63079), .B1(prod[102]), .B2(
        net66930), .ZN(n5123) );
  NAND2_X2 U5204 ( .A1(quo[104]), .A2(net66904), .ZN(n5122) );
  NAND3_X4 U5205 ( .A1(n5123), .A2(n5122), .A3(n5121), .ZN(fract_denorm[102])
         );
  AOI22_X2 U5206 ( .A1(fract_i2f[98]), .A2(net63083), .B1(prod[98]), .B2(
        net66928), .ZN(n5126) );
  NAND2_X2 U5207 ( .A1(quo[100]), .A2(net66905), .ZN(n5125) );
  AOI22_X2 U5208 ( .A1(fract_out_q[49]), .A2(net63507), .B1(quo[48]), .B2(
        net66897), .ZN(n5124) );
  AOI22_X2 U5209 ( .A1(fract_i2f[99]), .A2(net63083), .B1(prod[99]), .B2(
        net66929), .ZN(n5129) );
  NAND2_X2 U5210 ( .A1(quo[101]), .A2(net66906), .ZN(n5128) );
  AOI22_X2 U5211 ( .A1(fract_out_q[50]), .A2(net63507), .B1(quo[49]), .B2(
        net66897), .ZN(n5127) );
  NAND3_X4 U5212 ( .A1(n5129), .A2(n5128), .A3(n5127), .ZN(fract_denorm[99])
         );
  AOI22_X2 U5213 ( .A1(fract_i2f[95]), .A2(net63083), .B1(prod[95]), .B2(
        net66930), .ZN(n5132) );
  NAND2_X2 U5214 ( .A1(quo[97]), .A2(net66907), .ZN(n5131) );
  NAND3_X4 U5215 ( .A1(n5132), .A2(n5131), .A3(n5130), .ZN(fract_denorm[95])
         );
  AOI22_X2 U5216 ( .A1(fract_i2f[96]), .A2(net63083), .B1(prod[96]), .B2(
        net66928), .ZN(net60610) );
  AOI22_X2 U5217 ( .A1(fract_i2f[97]), .A2(net63083), .B1(prod[97]), .B2(
        net66929), .ZN(net60606) );
  NAND2_X2 U5218 ( .A1(quo[99]), .A2(net66914), .ZN(net60607) );
  AOI22_X2 U5219 ( .A1(fract_i2f[93]), .A2(net63079), .B1(prod[93]), .B2(
        net66930), .ZN(n5135) );
  NAND2_X2 U5220 ( .A1(quo[95]), .A2(net66904), .ZN(n5134) );
  AOI22_X2 U5221 ( .A1(fract_out_q[44]), .A2(net63507), .B1(quo[43]), .B2(
        net66897), .ZN(n5133) );
  NAND3_X4 U5222 ( .A1(n5135), .A2(n5134), .A3(n5133), .ZN(fract_denorm[93])
         );
  AOI22_X2 U5223 ( .A1(fract_i2f[94]), .A2(net63079), .B1(prod[94]), .B2(
        net66928), .ZN(net60599) );
  NAND2_X2 U5224 ( .A1(quo[96]), .A2(net66905), .ZN(net60600) );
  AOI22_X2 U5225 ( .A1(fract_i2f[90]), .A2(net63079), .B1(prod[90]), .B2(
        net66929), .ZN(n5138) );
  NAND2_X2 U5226 ( .A1(quo[92]), .A2(net66906), .ZN(n5137) );
  AOI22_X2 U5227 ( .A1(fract_out_q[41]), .A2(net63507), .B1(quo[40]), .B2(
        net66897), .ZN(n5136) );
  AOI22_X2 U5228 ( .A1(fract_i2f[91]), .A2(net63079), .B1(prod[91]), .B2(
        net66930), .ZN(n5141) );
  NAND2_X2 U5229 ( .A1(quo[93]), .A2(net66906), .ZN(n5140) );
  AOI22_X2 U5230 ( .A1(fract_out_q[42]), .A2(net63513), .B1(quo[41]), .B2(
        net66897), .ZN(n5139) );
  NAND3_X4 U5231 ( .A1(n5141), .A2(n5140), .A3(n5139), .ZN(fract_denorm[91])
         );
  AOI22_X2 U5232 ( .A1(fract_i2f[92]), .A2(net63079), .B1(prod[92]), .B2(
        net66928), .ZN(net60587) );
  NAND2_X2 U5233 ( .A1(quo[94]), .A2(net66910), .ZN(net60588) );
  AOI22_X2 U5234 ( .A1(fract_i2f[89]), .A2(net63079), .B1(prod[89]), .B2(
        net66929), .ZN(n5144) );
  NAND2_X2 U5235 ( .A1(quo[91]), .A2(net66911), .ZN(n5143) );
  AOI22_X2 U5236 ( .A1(fract_out_q[40]), .A2(net63503), .B1(quo[39]), .B2(
        net66897), .ZN(n5142) );
  NAND3_X4 U5237 ( .A1(n5144), .A2(n5143), .A3(n5142), .ZN(fract_denorm[89])
         );
  AOI22_X2 U5238 ( .A1(fract_i2f[87]), .A2(net63079), .B1(prod[87]), .B2(
        net66930), .ZN(n5147) );
  NAND2_X2 U5239 ( .A1(quo[89]), .A2(net66912), .ZN(n5146) );
  AOI22_X2 U5240 ( .A1(fract_out_q[38]), .A2(net63503), .B1(quo[37]), .B2(
        net66895), .ZN(n5145) );
  NAND3_X4 U5241 ( .A1(n5147), .A2(n5146), .A3(n5145), .ZN(fract_denorm[87])
         );
  AOI22_X2 U5242 ( .A1(fract_i2f[88]), .A2(net63079), .B1(prod[88]), .B2(
        net66928), .ZN(n5150) );
  NAND2_X2 U5243 ( .A1(quo[90]), .A2(net66914), .ZN(n5149) );
  AOI22_X2 U5244 ( .A1(fract_out_q[39]), .A2(net63513), .B1(quo[38]), .B2(
        net66897), .ZN(n5148) );
  NAND3_X4 U5245 ( .A1(n5150), .A2(n5149), .A3(n5148), .ZN(fract_denorm[88])
         );
  AOI22_X2 U5246 ( .A1(fract_i2f[85]), .A2(net63079), .B1(prod[85]), .B2(
        net66929), .ZN(n5153) );
  NAND2_X2 U5247 ( .A1(quo[87]), .A2(net66914), .ZN(n5152) );
  AOI22_X2 U5248 ( .A1(fract_out_q[36]), .A2(net63513), .B1(quo[35]), .B2(
        net66896), .ZN(n5151) );
  AOI22_X2 U5249 ( .A1(fract_i2f[86]), .A2(net63079), .B1(prod[86]), .B2(
        net66930), .ZN(n5156) );
  NAND2_X2 U5250 ( .A1(quo[88]), .A2(net66907), .ZN(n5155) );
  AOI22_X2 U5251 ( .A1(fract_out_q[37]), .A2(net63511), .B1(net66895), .B2(
        quo[36]), .ZN(n5154) );
  NAND3_X4 U5252 ( .A1(n5156), .A2(n5155), .A3(n5154), .ZN(fract_denorm[86])
         );
  AOI22_X2 U5253 ( .A1(fract_i2f[82]), .A2(net63079), .B1(prod[82]), .B2(
        net66928), .ZN(n5159) );
  NAND2_X2 U5254 ( .A1(quo[84]), .A2(net66910), .ZN(n5158) );
  AOI22_X2 U5255 ( .A1(fract_out_q[33]), .A2(net63513), .B1(quo[32]), .B2(
        net66896), .ZN(n5157) );
  NAND3_X4 U5256 ( .A1(n5159), .A2(n5158), .A3(n5157), .ZN(fract_denorm[82])
         );
  AOI22_X2 U5257 ( .A1(fract_i2f[83]), .A2(net63079), .B1(prod[83]), .B2(
        net66929), .ZN(n5162) );
  NAND2_X2 U5258 ( .A1(quo[85]), .A2(net66910), .ZN(n5161) );
  AOI22_X2 U5259 ( .A1(fract_out_q[34]), .A2(net63513), .B1(quo[33]), .B2(
        net66895), .ZN(n5160) );
  NAND3_X4 U5260 ( .A1(n5162), .A2(n5161), .A3(n5160), .ZN(fract_denorm[83])
         );
  AOI22_X2 U5261 ( .A1(fract_i2f[84]), .A2(net63079), .B1(prod[84]), .B2(
        net66930), .ZN(n5165) );
  NAND2_X2 U5262 ( .A1(quo[86]), .A2(net66911), .ZN(n5164) );
  AOI22_X2 U5263 ( .A1(fract_out_q[35]), .A2(net63503), .B1(quo[34]), .B2(
        net66897), .ZN(n5163) );
  NAND3_X4 U5264 ( .A1(n5165), .A2(n5164), .A3(n5163), .ZN(fract_denorm[84])
         );
  AOI22_X2 U5265 ( .A1(fract_i2f[74]), .A2(net63079), .B1(prod[74]), .B2(
        net66928), .ZN(n5168) );
  NAND2_X2 U5266 ( .A1(quo[76]), .A2(net66907), .ZN(n5167) );
  AOI22_X2 U5267 ( .A1(fract_out_q[25]), .A2(net63503), .B1(quo[24]), .B2(
        net66897), .ZN(n5166) );
  NAND3_X4 U5268 ( .A1(n5168), .A2(n5167), .A3(n5166), .ZN(fract_denorm[74])
         );
  AOI22_X2 U5269 ( .A1(fract_i2f[75]), .A2(net63079), .B1(prod[75]), .B2(
        net66929), .ZN(net60548) );
  NAND2_X2 U5270 ( .A1(quo[77]), .A2(net66904), .ZN(net60549) );
  AOI22_X2 U5271 ( .A1(fract_i2f[67]), .A2(net63079), .B1(prod[67]), .B2(
        net66930), .ZN(n5171) );
  NAND2_X2 U5272 ( .A1(quo[69]), .A2(net66905), .ZN(n5170) );
  AOI22_X2 U5273 ( .A1(fract_out_q[18]), .A2(net63503), .B1(quo[17]), .B2(
        net66895), .ZN(n5169) );
  NAND3_X4 U5274 ( .A1(n5171), .A2(n5170), .A3(n5169), .ZN(fract_denorm[67])
         );
  AOI22_X2 U5275 ( .A1(fract_i2f[68]), .A2(net63079), .B1(prod[68]), .B2(
        net66928), .ZN(n5174) );
  NAND2_X2 U5276 ( .A1(quo[70]), .A2(net66906), .ZN(n5173) );
  AOI22_X2 U5277 ( .A1(fract_out_q[19]), .A2(net63503), .B1(quo[18]), .B2(
        net66895), .ZN(n5172) );
  NAND3_X4 U5278 ( .A1(n5174), .A2(n5173), .A3(n5172), .ZN(fract_denorm[68])
         );
  AOI22_X2 U5279 ( .A1(fract_i2f[66]), .A2(net63079), .B1(prod[66]), .B2(
        net66929), .ZN(net60536) );
  NAND2_X2 U5280 ( .A1(quo[68]), .A2(net66907), .ZN(net60537) );
  AOI22_X2 U5281 ( .A1(fract_i2f[64]), .A2(net63079), .B1(prod[64]), .B2(
        net66930), .ZN(n5177) );
  NAND2_X2 U5282 ( .A1(quo[66]), .A2(net66910), .ZN(n5176) );
  AOI22_X2 U5283 ( .A1(fract_out_q[15]), .A2(net63503), .B1(quo[14]), .B2(
        net66896), .ZN(n5175) );
  NAND3_X4 U5284 ( .A1(n5177), .A2(n5176), .A3(n5175), .ZN(fract_denorm[64])
         );
  AOI22_X2 U5285 ( .A1(fract_i2f[65]), .A2(net63079), .B1(prod[65]), .B2(
        net66928), .ZN(n5180) );
  NAND2_X2 U5286 ( .A1(quo[67]), .A2(net66912), .ZN(n5179) );
  AOI22_X2 U5287 ( .A1(fract_out_q[16]), .A2(net63503), .B1(quo[15]), .B2(
        net66897), .ZN(n5178) );
  NAND3_X4 U5288 ( .A1(n5180), .A2(n5179), .A3(n5178), .ZN(fract_denorm[65])
         );
  AOI22_X2 U5289 ( .A1(fract_i2f[61]), .A2(net63079), .B1(prod[61]), .B2(
        net66929), .ZN(n5183) );
  NAND2_X2 U5290 ( .A1(quo[63]), .A2(net66906), .ZN(n5182) );
  AOI22_X2 U5291 ( .A1(fract_out_q[12]), .A2(net63511), .B1(net66895), .B2(
        quo[11]), .ZN(n5181) );
  NAND3_X4 U5292 ( .A1(n5183), .A2(n5182), .A3(n5181), .ZN(fract_denorm[61])
         );
  AOI22_X2 U5293 ( .A1(fract_i2f[62]), .A2(net63083), .B1(prod[62]), .B2(
        net66930), .ZN(n5186) );
  NAND2_X2 U5294 ( .A1(quo[64]), .A2(net66914), .ZN(n5185) );
  AOI22_X2 U5295 ( .A1(fract_out_q[13]), .A2(net63511), .B1(net66896), .B2(
        quo[12]), .ZN(n5184) );
  NAND3_X4 U5296 ( .A1(n5186), .A2(n5185), .A3(n5184), .ZN(fract_denorm[62])
         );
  AOI22_X2 U5297 ( .A1(fract_i2f[63]), .A2(net63083), .B1(prod[63]), .B2(
        net66928), .ZN(n5189) );
  NAND2_X2 U5298 ( .A1(quo[65]), .A2(net66904), .ZN(n5188) );
  AOI22_X2 U5299 ( .A1(fract_out_q[14]), .A2(net63503), .B1(quo[13]), .B2(
        net66897), .ZN(n5187) );
  NAND3_X4 U5300 ( .A1(n5189), .A2(n5188), .A3(n5187), .ZN(fract_denorm[63])
         );
  AOI22_X2 U5301 ( .A1(fract_i2f[59]), .A2(net63085), .B1(prod[59]), .B2(
        net66929), .ZN(n5192) );
  NAND2_X2 U5302 ( .A1(quo[61]), .A2(net66910), .ZN(n5191) );
  AOI22_X2 U5303 ( .A1(fract_out_q[10]), .A2(net63511), .B1(net66896), .B2(
        quo[9]), .ZN(n5190) );
  NAND3_X4 U5304 ( .A1(n5192), .A2(n5191), .A3(n5190), .ZN(fract_denorm[59])
         );
  AOI22_X2 U5305 ( .A1(fract_i2f[60]), .A2(net63083), .B1(prod[60]), .B2(
        net66930), .ZN(n5195) );
  NAND2_X2 U5306 ( .A1(quo[62]), .A2(net66910), .ZN(n5194) );
  AOI22_X2 U5307 ( .A1(fract_out_q[11]), .A2(net63511), .B1(net66897), .B2(
        quo[10]), .ZN(n5193) );
  NAND3_X4 U5308 ( .A1(n5195), .A2(n5194), .A3(n5193), .ZN(fract_denorm[60])
         );
  AOI22_X2 U5309 ( .A1(fract_i2f[58]), .A2(net63085), .B1(prod[58]), .B2(
        net66928), .ZN(net60509) );
  NAND2_X2 U5310 ( .A1(quo[60]), .A2(net66911), .ZN(net60510) );
  NAND2_X2 U5311 ( .A1(prod[45]), .A2(net66928), .ZN(n5198) );
  NAND2_X2 U5312 ( .A1(fract_i2f[45]), .A2(net63083), .ZN(n5197) );
  NAND2_X2 U5313 ( .A1(quo[47]), .A2(net66912), .ZN(n5196) );
  NAND3_X4 U5314 ( .A1(n5198), .A2(n5197), .A3(n5196), .ZN(net33585) );
  NAND2_X2 U5315 ( .A1(prod[46]), .A2(net66929), .ZN(n5201) );
  NAND2_X2 U5316 ( .A1(fract_i2f[46]), .A2(net63083), .ZN(n5200) );
  NAND2_X2 U5317 ( .A1(quo[48]), .A2(net66910), .ZN(n5199) );
  NAND3_X4 U5318 ( .A1(n5201), .A2(n5200), .A3(n5199), .ZN(net33584) );
  NAND2_X2 U5319 ( .A1(prod[48]), .A2(net66930), .ZN(n5204) );
  NAND2_X2 U5320 ( .A1(fract_i2f[48]), .A2(net63083), .ZN(n5203) );
  NAND2_X2 U5321 ( .A1(quo[50]), .A2(net66914), .ZN(n5202) );
  NAND3_X4 U5322 ( .A1(n5204), .A2(n5203), .A3(n5202), .ZN(net33583) );
  NAND2_X2 U5323 ( .A1(quo[51]), .A2(net66905), .ZN(n5207) );
  NAND2_X2 U5324 ( .A1(prod[49]), .A2(net66928), .ZN(n5206) );
  AOI22_X2 U5325 ( .A1(fract_out_q[0]), .A2(net63509), .B1(fract_i2f[49]), 
        .B2(net63085), .ZN(n5205) );
  NAND3_X4 U5326 ( .A1(n5207), .A2(n5206), .A3(n5205), .ZN(net33625) );
  NAND2_X2 U5327 ( .A1(prod[47]), .A2(net66929), .ZN(n5210) );
  NAND2_X2 U5328 ( .A1(fract_i2f[47]), .A2(net63083), .ZN(n5209) );
  NAND2_X2 U5329 ( .A1(quo[49]), .A2(net66906), .ZN(n5208) );
  NAND3_X4 U5330 ( .A1(n5210), .A2(n5209), .A3(n5208), .ZN(n8515) );
  AOI22_X2 U5331 ( .A1(fract_i2f[57]), .A2(net63083), .B1(prod[57]), .B2(
        net66929), .ZN(n5213) );
  NAND2_X2 U5332 ( .A1(quo[59]), .A2(net66907), .ZN(n5212) );
  AOI22_X2 U5333 ( .A1(fract_out_q[8]), .A2(net63509), .B1(net66896), .B2(
        quo[7]), .ZN(n5211) );
  NAND3_X4 U5334 ( .A1(n5213), .A2(n5212), .A3(n5211), .ZN(fract_denorm[57])
         );
  AOI22_X2 U5335 ( .A1(fract_i2f[55]), .A2(net63083), .B1(prod[55]), .B2(
        net66930), .ZN(n5216) );
  NAND2_X2 U5336 ( .A1(quo[57]), .A2(net66910), .ZN(n5215) );
  AOI22_X2 U5337 ( .A1(fract_out_q[6]), .A2(net63509), .B1(net66897), .B2(
        quo[5]), .ZN(n5214) );
  NAND3_X4 U5338 ( .A1(n5216), .A2(n5215), .A3(n5214), .ZN(fract_denorm[55])
         );
  AOI22_X2 U5339 ( .A1(fract_i2f[56]), .A2(net63083), .B1(prod[56]), .B2(
        net66928), .ZN(n5219) );
  NAND2_X2 U5340 ( .A1(quo[58]), .A2(net66910), .ZN(n5218) );
  AOI22_X2 U5341 ( .A1(fract_out_q[7]), .A2(net63509), .B1(net66895), .B2(
        quo[6]), .ZN(n5217) );
  NAND3_X4 U5342 ( .A1(n5219), .A2(n5218), .A3(n5217), .ZN(fract_denorm[56])
         );
  AOI22_X2 U5343 ( .A1(fract_i2f[53]), .A2(net63083), .B1(prod[53]), .B2(
        net66929), .ZN(n5222) );
  NAND2_X2 U5344 ( .A1(quo[55]), .A2(net66904), .ZN(n5221) );
  AOI22_X2 U5345 ( .A1(fract_out_q[4]), .A2(net63503), .B1(quo[3]), .B2(
        net66896), .ZN(n5220) );
  AOI22_X2 U5346 ( .A1(fract_i2f[54]), .A2(net63085), .B1(prod[54]), .B2(
        net66930), .ZN(n5225) );
  NAND2_X2 U5347 ( .A1(quo[56]), .A2(net66905), .ZN(n5224) );
  AOI22_X2 U5348 ( .A1(fract_out_q[5]), .A2(net63503), .B1(quo[4]), .B2(
        net66896), .ZN(n5223) );
  NAND3_X4 U5349 ( .A1(n5225), .A2(n5224), .A3(n5223), .ZN(fract_denorm[54])
         );
  AOI22_X2 U5350 ( .A1(fract_i2f[50]), .A2(net63085), .B1(prod[50]), .B2(
        net66928), .ZN(n5228) );
  NAND2_X2 U5351 ( .A1(quo[52]), .A2(net66906), .ZN(n5227) );
  AOI22_X2 U5352 ( .A1(fract_out_q[1]), .A2(net63503), .B1(quo[0]), .B2(
        net66895), .ZN(n5226) );
  NAND3_X4 U5353 ( .A1(n5228), .A2(n5227), .A3(n5226), .ZN(fract_denorm[50])
         );
  AOI22_X2 U5354 ( .A1(fract_i2f[51]), .A2(net63083), .B1(prod[51]), .B2(
        net66929), .ZN(n5230) );
  AOI22_X2 U5355 ( .A1(fract_out_q[2]), .A2(net63503), .B1(quo[1]), .B2(
        net66897), .ZN(n5229) );
  AOI22_X2 U5356 ( .A1(fract_i2f[52]), .A2(net63083), .B1(prod[52]), .B2(
        net66930), .ZN(n5232) );
  AOI22_X2 U5357 ( .A1(fract_out_q[3]), .A2(net63507), .B1(quo[2]), .B2(
        net66897), .ZN(n5231) );
  NAND2_X2 U5358 ( .A1(prod[43]), .A2(net66930), .ZN(net60461) );
  NAND2_X2 U5359 ( .A1(fract_i2f[43]), .A2(net63083), .ZN(net60462) );
  NAND2_X2 U5360 ( .A1(prod[44]), .A2(net66928), .ZN(n5234) );
  NAND2_X2 U5361 ( .A1(fract_i2f[44]), .A2(net63083), .ZN(n5233) );
  NAND3_X4 U5362 ( .A1(n5234), .A2(n5233), .A3(net60460), .ZN(net33586) );
  NAND2_X2 U5363 ( .A1(prod[35]), .A2(net66929), .ZN(n5237) );
  NAND2_X2 U5364 ( .A1(fract_i2f[35]), .A2(net63083), .ZN(n5236) );
  NAND2_X2 U5365 ( .A1(quo[37]), .A2(net66910), .ZN(n5235) );
  NAND3_X4 U5366 ( .A1(n5237), .A2(n5236), .A3(n5235), .ZN(net33559) );
  NAND2_X2 U5367 ( .A1(prod[36]), .A2(net66930), .ZN(n5240) );
  NAND2_X2 U5368 ( .A1(fract_i2f[36]), .A2(net63083), .ZN(n5239) );
  NAND2_X2 U5369 ( .A1(quo[38]), .A2(net66911), .ZN(n5238) );
  NAND3_X4 U5370 ( .A1(n5240), .A2(n5239), .A3(n5238), .ZN(net33558) );
  NAND2_X2 U5371 ( .A1(prod[37]), .A2(net66928), .ZN(n5243) );
  NAND2_X2 U5372 ( .A1(fract_i2f[37]), .A2(net63083), .ZN(n5242) );
  NAND2_X2 U5373 ( .A1(quo[39]), .A2(net66912), .ZN(n5241) );
  NAND3_X4 U5374 ( .A1(n5243), .A2(n5242), .A3(n5241), .ZN(n8522) );
  NAND2_X2 U5375 ( .A1(prod[38]), .A2(net66929), .ZN(n5246) );
  NAND2_X2 U5376 ( .A1(fract_i2f[38]), .A2(net63083), .ZN(n5245) );
  NAND2_X2 U5377 ( .A1(quo[40]), .A2(net66906), .ZN(n5244) );
  NAND3_X4 U5378 ( .A1(n5246), .A2(n5245), .A3(n5244), .ZN(n8523) );
  NAND2_X2 U5379 ( .A1(prod[40]), .A2(net66930), .ZN(n5249) );
  NAND2_X2 U5380 ( .A1(fract_i2f[40]), .A2(net63083), .ZN(n5248) );
  NAND2_X2 U5381 ( .A1(quo[42]), .A2(net66914), .ZN(n5247) );
  NAND3_X4 U5382 ( .A1(n5249), .A2(n5248), .A3(n5247), .ZN(n8524) );
  NAND2_X2 U5383 ( .A1(prod[41]), .A2(net66928), .ZN(n5252) );
  NAND2_X2 U5384 ( .A1(fract_i2f[41]), .A2(net63083), .ZN(n5251) );
  NAND2_X2 U5385 ( .A1(quo[43]), .A2(net66914), .ZN(n5250) );
  NAND3_X4 U5386 ( .A1(n5252), .A2(n5251), .A3(n5250), .ZN(net33554) );
  NAND2_X2 U5387 ( .A1(prod[39]), .A2(net66929), .ZN(n5255) );
  NAND2_X2 U5388 ( .A1(fract_i2f[39]), .A2(net63083), .ZN(n5254) );
  NAND2_X2 U5389 ( .A1(quo[41]), .A2(net66904), .ZN(n5253) );
  NAND3_X4 U5390 ( .A1(n5255), .A2(n5254), .A3(n5253), .ZN(n8525) );
  NAND2_X2 U5391 ( .A1(prod[27]), .A2(net66930), .ZN(n5258) );
  NAND2_X2 U5392 ( .A1(fract_i2f[27]), .A2(net63083), .ZN(n5257) );
  NAND2_X2 U5393 ( .A1(quo[29]), .A2(net66905), .ZN(n5256) );
  NAND3_X4 U5394 ( .A1(n5258), .A2(n5257), .A3(n5256), .ZN(net33566) );
  NAND2_X2 U5395 ( .A1(prod[28]), .A2(net66928), .ZN(n5261) );
  NAND2_X2 U5396 ( .A1(fract_i2f[28]), .A2(net63083), .ZN(n5260) );
  NAND2_X2 U5397 ( .A1(quo[30]), .A2(net66906), .ZN(n5259) );
  NAND3_X4 U5398 ( .A1(n5261), .A2(n5260), .A3(n5259), .ZN(net33565) );
  NAND2_X2 U5399 ( .A1(prod[29]), .A2(net66929), .ZN(n5264) );
  NAND2_X2 U5400 ( .A1(fract_i2f[29]), .A2(net63085), .ZN(n5263) );
  NAND2_X2 U5401 ( .A1(quo[31]), .A2(net66912), .ZN(n5262) );
  NAND3_X4 U5402 ( .A1(n5264), .A2(n5263), .A3(n5262), .ZN(net33564) );
  NAND2_X2 U5403 ( .A1(prod[30]), .A2(net66930), .ZN(n5267) );
  NAND2_X2 U5404 ( .A1(fract_i2f[30]), .A2(net63083), .ZN(n5266) );
  NAND2_X2 U5405 ( .A1(quo[32]), .A2(net66904), .ZN(n5265) );
  NAND3_X4 U5406 ( .A1(n5267), .A2(n5266), .A3(n5265), .ZN(net33563) );
  NAND2_X2 U5407 ( .A1(prod[32]), .A2(net66928), .ZN(n5270) );
  NAND2_X2 U5408 ( .A1(fract_i2f[32]), .A2(net63083), .ZN(n5269) );
  NAND2_X2 U5409 ( .A1(quo[34]), .A2(net66905), .ZN(n5268) );
  NAND3_X4 U5410 ( .A1(n5270), .A2(n5269), .A3(n5268), .ZN(net33562) );
  NAND2_X2 U5411 ( .A1(prod[33]), .A2(net66929), .ZN(n5273) );
  NAND2_X2 U5412 ( .A1(fract_i2f[33]), .A2(net63083), .ZN(n5272) );
  NAND2_X2 U5413 ( .A1(quo[35]), .A2(net66906), .ZN(n5271) );
  NAND3_X4 U5414 ( .A1(n5273), .A2(n5272), .A3(n5271), .ZN(net33561) );
  NAND2_X2 U5415 ( .A1(prod[31]), .A2(net66930), .ZN(n5276) );
  NAND2_X2 U5416 ( .A1(fract_i2f[31]), .A2(net63083), .ZN(n5275) );
  NAND2_X2 U5417 ( .A1(quo[33]), .A2(net66907), .ZN(n5274) );
  NAND3_X4 U5418 ( .A1(n5276), .A2(n5275), .A3(n5274), .ZN(n8521) );
  NAND2_X2 U5419 ( .A1(prod[19]), .A2(net66929), .ZN(n5279) );
  NAND2_X2 U5420 ( .A1(fract_i2f[19]), .A2(net63083), .ZN(n5278) );
  NAND2_X2 U5421 ( .A1(quo[21]), .A2(net66907), .ZN(n5277) );
  NAND3_X4 U5422 ( .A1(n5279), .A2(n5278), .A3(n5277), .ZN(net33573) );
  NAND2_X2 U5423 ( .A1(prod[20]), .A2(net66930), .ZN(n5282) );
  NAND2_X2 U5424 ( .A1(fract_i2f[20]), .A2(net63085), .ZN(n5281) );
  NAND2_X2 U5425 ( .A1(quo[22]), .A2(net66910), .ZN(n5280) );
  NAND3_X4 U5426 ( .A1(n5282), .A2(n5281), .A3(n5280), .ZN(net33572) );
  NAND2_X2 U5427 ( .A1(prod[23]), .A2(net66928), .ZN(n5285) );
  NAND2_X2 U5428 ( .A1(fract_i2f[23]), .A2(net63083), .ZN(n5284) );
  NAND2_X2 U5429 ( .A1(quo[25]), .A2(net66910), .ZN(n5283) );
  NAND3_X4 U5430 ( .A1(n5285), .A2(n5284), .A3(n5283), .ZN(n8520) );
  NAND2_X2 U5431 ( .A1(prod[24]), .A2(net66929), .ZN(n5288) );
  NAND2_X2 U5432 ( .A1(fract_i2f[24]), .A2(net63085), .ZN(n5287) );
  NAND2_X2 U5433 ( .A1(quo[26]), .A2(net66911), .ZN(n5286) );
  NAND3_X4 U5434 ( .A1(n5288), .A2(n5287), .A3(n5286), .ZN(net33569) );
  NAND2_X2 U5435 ( .A1(prod[25]), .A2(net66930), .ZN(n5291) );
  NAND2_X2 U5436 ( .A1(fract_i2f[25]), .A2(net63083), .ZN(n5290) );
  NAND2_X2 U5437 ( .A1(quo[27]), .A2(net66906), .ZN(n5289) );
  NAND3_X4 U5438 ( .A1(n5291), .A2(n5290), .A3(n5289), .ZN(net33568) );
  NAND2_X2 U5439 ( .A1(prod[21]), .A2(net66928), .ZN(n5294) );
  NAND2_X2 U5440 ( .A1(fract_i2f[21]), .A2(net63085), .ZN(n5293) );
  NAND2_X2 U5441 ( .A1(quo[23]), .A2(net66910), .ZN(n5292) );
  NAND3_X4 U5442 ( .A1(n5294), .A2(n5293), .A3(n5292), .ZN(n8518) );
  NAND2_X2 U5443 ( .A1(prod[22]), .A2(net66929), .ZN(n5297) );
  NAND2_X2 U5444 ( .A1(fract_i2f[22]), .A2(net63085), .ZN(n5296) );
  NAND2_X2 U5445 ( .A1(quo[24]), .A2(net66911), .ZN(n5295) );
  NAND3_X4 U5446 ( .A1(n5297), .A2(n5296), .A3(n5295), .ZN(n8519) );
  NAND2_X2 U5447 ( .A1(prod[12]), .A2(net66928), .ZN(n5300) );
  NAND2_X2 U5448 ( .A1(fract_i2f[12]), .A2(net63085), .ZN(n5299) );
  NAND2_X2 U5449 ( .A1(quo[14]), .A2(net66906), .ZN(n5298) );
  NAND3_X4 U5450 ( .A1(n5300), .A2(n5299), .A3(n5298), .ZN(net33579) );
  NAND2_X2 U5451 ( .A1(prod[13]), .A2(net66929), .ZN(n5303) );
  NAND2_X2 U5452 ( .A1(fract_i2f[13]), .A2(net63085), .ZN(n5302) );
  NAND2_X2 U5453 ( .A1(quo[15]), .A2(net66914), .ZN(n5301) );
  NAND3_X4 U5454 ( .A1(n5303), .A2(n5302), .A3(n5301), .ZN(net33578) );
  NAND2_X2 U5455 ( .A1(prod[14]), .A2(net66930), .ZN(n5306) );
  NAND2_X2 U5456 ( .A1(fract_i2f[14]), .A2(net63085), .ZN(n5305) );
  NAND2_X2 U5457 ( .A1(quo[16]), .A2(net66912), .ZN(n5304) );
  NAND3_X4 U5458 ( .A1(n5306), .A2(n5305), .A3(n5304), .ZN(net33577) );
  NAND2_X2 U5459 ( .A1(prod[16]), .A2(net66928), .ZN(n5309) );
  NAND2_X2 U5460 ( .A1(fract_i2f[16]), .A2(net63085), .ZN(n5308) );
  NAND2_X2 U5461 ( .A1(quo[18]), .A2(net66906), .ZN(n5307) );
  NAND3_X4 U5462 ( .A1(n5309), .A2(n5308), .A3(n5307), .ZN(n8516) );
  NAND2_X2 U5463 ( .A1(prod[17]), .A2(net66929), .ZN(n5312) );
  NAND2_X2 U5464 ( .A1(fract_i2f[17]), .A2(net63085), .ZN(n5311) );
  NAND2_X2 U5465 ( .A1(quo[19]), .A2(net66914), .ZN(n5310) );
  NAND3_X4 U5466 ( .A1(n5312), .A2(n5311), .A3(n5310), .ZN(net33575) );
  NAND2_X2 U5467 ( .A1(prod[15]), .A2(net66930), .ZN(n5315) );
  NAND2_X2 U5468 ( .A1(fract_i2f[15]), .A2(net63085), .ZN(n5314) );
  NAND2_X2 U5469 ( .A1(quo[17]), .A2(net66904), .ZN(n5313) );
  NAND3_X4 U5470 ( .A1(n5315), .A2(n5314), .A3(n5313), .ZN(n8517) );
  NOR2_X4 U5471 ( .A1(fract_denorm[55]), .A2(fract_denorm[57]), .ZN(n5317) );
  INV_X4 U5472 ( .A(fract_denorm[56]), .ZN(n5316) );
  NAND2_X2 U5473 ( .A1(n5317), .A2(n5316), .ZN(net60065) );
  NOR3_X4 U5474 ( .A1(fract_denorm[63]), .A2(fract_denorm[62]), .A3(
        fract_denorm[61]), .ZN(net60329) );
  NOR3_X4 U5475 ( .A1(fract_denorm[88]), .A2(fract_denorm[87]), .A3(
        fract_denorm[89]), .ZN(n5410) );
  INV_X4 U5476 ( .A(fract_denorm[85]), .ZN(n5412) );
  INV_X4 U5477 ( .A(fract_denorm[86]), .ZN(n5318) );
  NOR2_X4 U5478 ( .A1(fract_denorm[103]), .A2(fract_denorm[104]), .ZN(net59958) );
  NOR3_X4 U5479 ( .A1(fract_denorm[102]), .A2(fract_denorm[101]), .A3(
        fract_denorm[100]), .ZN(net59920) );
  NOR2_X4 U5480 ( .A1(fract_denorm[81]), .A2(fract_denorm[80]), .ZN(n5376) );
  NOR3_X4 U5481 ( .A1(fract_denorm[79]), .A2(fract_denorm[78]), .A3(
        fract_denorm[77]), .ZN(n5336) );
  NAND2_X2 U5482 ( .A1(n5376), .A2(n5336), .ZN(net60202) );
  NOR3_X4 U5483 ( .A1(fract_denorm[72]), .A2(fract_denorm[71]), .A3(
        fract_denorm[73]), .ZN(net60062) );
  NOR2_X4 U5484 ( .A1(fract_denorm[51]), .A2(fract_denorm[50]), .ZN(net60185)
         );
  NOR2_X4 U5485 ( .A1(net33625), .A2(net33583), .ZN(n5397) );
  INV_X4 U5486 ( .A(n8515), .ZN(n5319) );
  NAND2_X2 U5487 ( .A1(n5397), .A2(n5319), .ZN(net60157) );
  NOR3_X4 U5488 ( .A1(net60157), .A2(net33584), .A3(net33585), .ZN(net60317)
         );
  INV_X4 U5489 ( .A(net33587), .ZN(net60346) );
  NOR2_X4 U5490 ( .A1(n8523), .A2(n8522), .ZN(n5322) );
  INV_X4 U5491 ( .A(n8524), .ZN(n5321) );
  NOR2_X4 U5492 ( .A1(n8525), .A2(net33554), .ZN(n5320) );
  NAND3_X4 U5493 ( .A1(n5322), .A2(n5321), .A3(n5320), .ZN(net59991) );
  INV_X4 U5494 ( .A(net33562), .ZN(net59965) );
  INV_X4 U5495 ( .A(net60340), .ZN(net60117) );
  INV_X4 U5496 ( .A(n8521), .ZN(n5323) );
  NAND2_X2 U5497 ( .A1(net60117), .A2(n5323), .ZN(net60150) );
  NOR3_X4 U5498 ( .A1(net60150), .A2(net33563), .A3(net33564), .ZN(net60096)
         );
  INV_X4 U5499 ( .A(n8518), .ZN(n5325) );
  INV_X4 U5500 ( .A(n8519), .ZN(n5324) );
  INV_X4 U5501 ( .A(net33568), .ZN(net60008) );
  NAND3_X4 U5502 ( .A1(n5325), .A2(n5324), .A3(net60008), .ZN(n5326) );
  NOR3_X4 U5503 ( .A1(n5326), .A2(net33569), .A3(n8520), .ZN(net60290) );
  NOR2_X4 U5504 ( .A1(net33579), .A2(net33581), .ZN(net60330) );
  INV_X4 U5505 ( .A(n8516), .ZN(n5327) );
  INV_X4 U5506 ( .A(net33575), .ZN(net60084) );
  NAND2_X2 U5507 ( .A1(n5327), .A2(net60084), .ZN(n5328) );
  INV_X4 U5508 ( .A(n5328), .ZN(n5396) );
  INV_X4 U5509 ( .A(n8517), .ZN(n5329) );
  NAND2_X2 U5510 ( .A1(n5396), .A2(n5329), .ZN(net60147) );
  INV_X4 U5511 ( .A(net59328), .ZN(net60186) );
  NOR3_X4 U5512 ( .A1(net60310), .A2(net60221), .A3(n5342), .ZN(n5333) );
  NAND3_X4 U5513 ( .A1(n5334), .A2(net60308), .A3(n5333), .ZN(u4_fi_ldz_5_) );
  INV_X4 U5514 ( .A(fract_denorm[90]), .ZN(net60306) );
  INV_X4 U5515 ( .A(net33581), .ZN(net60303) );
  INV_X4 U5516 ( .A(net60302), .ZN(net60301) );
  INV_X4 U5517 ( .A(n5336), .ZN(n5337) );
  INV_X4 U5518 ( .A(n5338), .ZN(n5416) );
  NAND2_X2 U5519 ( .A1(n5416), .A2(fract_denorm[83]), .ZN(net60292) );
  INV_X4 U5520 ( .A(net60273), .ZN(net60049) );
  NAND2_X2 U5521 ( .A1(net60049), .A2(net33573), .ZN(net60293) );
  NAND2_X2 U5522 ( .A1(n4515), .A2(fract_denorm[80]), .ZN(n5340) );
  INV_X4 U5523 ( .A(fract_denorm[83]), .ZN(net60281) );
  NAND4_X2 U5524 ( .A1(fract_denorm[82]), .A2(net60044), .A3(net60281), .A4(
        n5416), .ZN(n5339) );
  INV_X4 U5525 ( .A(net60202), .ZN(net60276) );
  NAND2_X2 U5526 ( .A1(n5416), .A2(fract_denorm[84]), .ZN(n5341) );
  NAND2_X2 U5527 ( .A1(prod[2]), .A2(net66928), .ZN(n5348) );
  NAND2_X2 U5528 ( .A1(fract_i2f[2]), .A2(net63085), .ZN(n5347) );
  NAND2_X2 U5529 ( .A1(quo[4]), .A2(net66914), .ZN(n5346) );
  NAND3_X4 U5530 ( .A1(n5348), .A2(n5347), .A3(n5346), .ZN(net33647) );
  NAND2_X2 U5531 ( .A1(prod[3]), .A2(net66929), .ZN(n5351) );
  NAND2_X2 U5532 ( .A1(fract_i2f[3]), .A2(net63085), .ZN(n5350) );
  NAND2_X2 U5533 ( .A1(quo[5]), .A2(net66904), .ZN(n5349) );
  NAND3_X4 U5534 ( .A1(n5351), .A2(n5350), .A3(n5349), .ZN(n8511) );
  NAND2_X2 U5535 ( .A1(prod[4]), .A2(net66930), .ZN(n5354) );
  NAND2_X2 U5536 ( .A1(fract_i2f[4]), .A2(net63085), .ZN(n5353) );
  NAND2_X2 U5537 ( .A1(quo[6]), .A2(net66905), .ZN(n5352) );
  NAND3_X4 U5538 ( .A1(n5354), .A2(n5353), .A3(n5352), .ZN(n8512) );
  NAND2_X2 U5539 ( .A1(prod[5]), .A2(net66928), .ZN(n5357) );
  NAND2_X2 U5540 ( .A1(fract_i2f[5]), .A2(net63085), .ZN(n5356) );
  NAND2_X2 U5541 ( .A1(quo[7]), .A2(net66906), .ZN(n5355) );
  NAND3_X4 U5542 ( .A1(n5357), .A2(n5356), .A3(n5355), .ZN(n8513) );
  NAND2_X2 U5543 ( .A1(prod[6]), .A2(net66929), .ZN(n5360) );
  NAND2_X2 U5544 ( .A1(fract_i2f[6]), .A2(net63085), .ZN(n5359) );
  NAND2_X2 U5545 ( .A1(quo[8]), .A2(net66907), .ZN(n5358) );
  NAND3_X4 U5546 ( .A1(n5360), .A2(n5359), .A3(n5358), .ZN(n8514) );
  NAND2_X2 U5547 ( .A1(prod[7]), .A2(net66930), .ZN(n5363) );
  NAND2_X2 U5548 ( .A1(fract_i2f[7]), .A2(net63085), .ZN(n5362) );
  NAND2_X2 U5549 ( .A1(quo[9]), .A2(net66910), .ZN(n5361) );
  NAND3_X4 U5550 ( .A1(n5363), .A2(n5362), .A3(n5361), .ZN(net33642) );
  NAND2_X2 U5551 ( .A1(prod[8]), .A2(net66928), .ZN(n5366) );
  NAND2_X2 U5552 ( .A1(fract_i2f[8]), .A2(net63085), .ZN(n5365) );
  NAND2_X2 U5553 ( .A1(quo[10]), .A2(net66905), .ZN(n5364) );
  NAND3_X4 U5554 ( .A1(n5366), .A2(n5365), .A3(n5364), .ZN(net33641) );
  NAND2_X2 U5555 ( .A1(prod[10]), .A2(net66929), .ZN(n5369) );
  NAND2_X2 U5556 ( .A1(fract_i2f[10]), .A2(net63085), .ZN(n5368) );
  NAND2_X2 U5557 ( .A1(quo[12]), .A2(net66906), .ZN(n5367) );
  NAND3_X4 U5558 ( .A1(n5369), .A2(n5368), .A3(n5367), .ZN(net33549) );
  NAND2_X2 U5559 ( .A1(prod[9]), .A2(net66930), .ZN(n5372) );
  NAND2_X2 U5560 ( .A1(fract_i2f[9]), .A2(net63085), .ZN(n5371) );
  NAND2_X2 U5561 ( .A1(quo[11]), .A2(net66907), .ZN(n5370) );
  NAND3_X4 U5562 ( .A1(n5372), .A2(n5371), .A3(n5370), .ZN(net33548) );
  NAND2_X2 U5563 ( .A1(prod[1]), .A2(net66928), .ZN(n5375) );
  NAND2_X2 U5564 ( .A1(fract_i2f[1]), .A2(net63085), .ZN(n5374) );
  NAND2_X2 U5565 ( .A1(net66904), .A2(quo[3]), .ZN(n5373) );
  INV_X4 U5566 ( .A(fract_denorm[62]), .ZN(net60237) );
  INV_X4 U5567 ( .A(fract_denorm[78]), .ZN(n5377) );
  NAND2_X2 U5568 ( .A1(n4515), .A2(n5376), .ZN(n5398) );
  INV_X4 U5569 ( .A(net60157), .ZN(net60230) );
  NAND4_X2 U5570 ( .A1(net60223), .A2(n5380), .A3(n5379), .A4(n5378), .ZN(
        n5468) );
  NAND3_X4 U5571 ( .A1(net60215), .A2(n5383), .A3(n5382), .ZN(n5394) );
  INV_X4 U5572 ( .A(fract_denorm[51]), .ZN(n5384) );
  INV_X4 U5573 ( .A(n5385), .ZN(n5393) );
  INV_X4 U5574 ( .A(net60038), .ZN(net60174) );
  INV_X4 U5575 ( .A(n8511), .ZN(n5386) );
  INV_X4 U5576 ( .A(n8512), .ZN(n5417) );
  NAND2_X2 U5577 ( .A1(n5386), .A2(n5417), .ZN(net59333) );
  INV_X4 U5578 ( .A(net59333), .ZN(net60176) );
  INV_X4 U5579 ( .A(n8513), .ZN(n5414) );
  INV_X4 U5580 ( .A(n8514), .ZN(n5465) );
  NAND2_X2 U5581 ( .A1(n5414), .A2(n5465), .ZN(net59324) );
  INV_X4 U5582 ( .A(net59324), .ZN(net60177) );
  INV_X4 U5583 ( .A(net33642), .ZN(net60208) );
  NOR3_X4 U5584 ( .A1(net59341), .A2(net33550), .A3(net33547), .ZN(n5390) );
  NAND3_X4 U5585 ( .A1(net60197), .A2(n5387), .A3(net60199), .ZN(n5388) );
  NOR3_X4 U5586 ( .A1(n5388), .A2(net60189), .A3(net60190), .ZN(net59423) );
  NOR2_X4 U5587 ( .A1(net60182), .A2(net60183), .ZN(n5389) );
  NAND3_X4 U5588 ( .A1(n5390), .A2(net60180), .A3(n5389), .ZN(net59954) );
  INV_X4 U5589 ( .A(net59954), .ZN(net60026) );
  INV_X4 U5590 ( .A(net59927), .ZN(net60178) );
  NAND2_X2 U5591 ( .A1(net60177), .A2(net60178), .ZN(n5436) );
  INV_X4 U5592 ( .A(n5436), .ZN(n5418) );
  NAND2_X2 U5593 ( .A1(net60176), .A2(n5418), .ZN(net60081) );
  INV_X4 U5594 ( .A(n5391), .ZN(n5392) );
  NOR3_X4 U5595 ( .A1(n5394), .A2(n5393), .A3(n5392), .ZN(n5406) );
  INV_X4 U5596 ( .A(net33585), .ZN(net60158) );
  INV_X4 U5597 ( .A(fract_denorm[79]), .ZN(n5399) );
  NAND2_X2 U5598 ( .A1(fract_denorm[77]), .A2(n5399), .ZN(n5395) );
  INV_X4 U5599 ( .A(fract_denorm[95]), .ZN(net60114) );
  NAND4_X2 U5600 ( .A1(n5402), .A2(n5401), .A3(n5400), .A4(net60105), .ZN(
        net59975) );
  INV_X4 U5601 ( .A(net60095), .ZN(net60088) );
  INV_X4 U5602 ( .A(net33647), .ZN(net60082) );
  INV_X4 U5603 ( .A(net59323), .ZN(net59699) );
  INV_X4 U5604 ( .A(net60081), .ZN(net59697) );
  NAND2_X2 U5605 ( .A1(net59699), .A2(net59697), .ZN(n5404) );
  NAND3_X4 U5606 ( .A1(n5407), .A2(n5406), .A3(net60077), .ZN(u4_fi_ldz_3_) );
  INV_X4 U5607 ( .A(net33569), .ZN(net60073) );
  INV_X4 U5608 ( .A(n5411), .ZN(n5458) );
  NAND2_X2 U5609 ( .A1(n5458), .A2(n5413), .ZN(net60056) );
  NAND2_X2 U5610 ( .A1(net60004), .A2(net60062), .ZN(net59923) );
  INV_X4 U5611 ( .A(net33572), .ZN(net60050) );
  INV_X4 U5612 ( .A(net33559), .ZN(net60048) );
  INV_X4 U5613 ( .A(fract_denorm[84]), .ZN(net60044) );
  INV_X4 U5614 ( .A(n5419), .ZN(n5420) );
  NAND4_X2 U5615 ( .A1(n5424), .A2(net60028), .A3(n5423), .A4(n5422), .ZN(
        net59982) );
  AOI21_X4 U5616 ( .B1(n4320), .B2(n8520), .A(n4373), .ZN(n5433) );
  NAND2_X2 U5617 ( .A1(n5460), .A2(n8525), .ZN(n5432) );
  INV_X4 U5618 ( .A(fract_denorm[55]), .ZN(n5425) );
  INV_X4 U5619 ( .A(fract_denorm[87]), .ZN(n5426) );
  INV_X4 U5620 ( .A(fract_denorm[73]), .ZN(net60020) );
  NAND2_X2 U5621 ( .A1(net60004), .A2(net60020), .ZN(n5451) );
  INV_X4 U5622 ( .A(fract_denorm[71]), .ZN(n5427) );
  INV_X4 U5623 ( .A(fract_denorm[102]), .ZN(n5434) );
  INV_X4 U5624 ( .A(net33554), .ZN(net60011) );
  INV_X4 U5625 ( .A(fract_denorm[68]), .ZN(net59993) );
  INV_X4 U5626 ( .A(net33558), .ZN(net59990) );
  NOR4_X2 U5627 ( .A1(net59911), .A2(net59974), .A3(net59975), .A4(net59976), 
        .ZN(n5457) );
  NAND2_X2 U5628 ( .A1(n5441), .A2(fract_denorm[56]), .ZN(n5442) );
  INV_X4 U5629 ( .A(n5442), .ZN(n5443) );
  AOI21_X4 U5630 ( .B1(n5444), .B2(n8524), .A(n5443), .ZN(n5445) );
  INV_X4 U5631 ( .A(n5445), .ZN(n5447) );
  AOI211_X4 U5632 ( .C1(net59962), .C2(net33569), .A(n5447), .B(n5446), .ZN(
        n5456) );
  INV_X4 U5633 ( .A(net59952), .ZN(net59951) );
  NAND2_X2 U5634 ( .A1(net59951), .A2(fract_denorm[88]), .ZN(n5450) );
  INV_X4 U5635 ( .A(fract_denorm[81]), .ZN(net59950) );
  NAND2_X2 U5636 ( .A1(n5450), .A2(n5449), .ZN(n5454) );
  INV_X4 U5637 ( .A(fract_denorm[72]), .ZN(n5452) );
  NOR4_X2 U5638 ( .A1(net59939), .A2(n5454), .A3(net59941), .A4(n5453), .ZN(
        n5455) );
  NAND3_X4 U5639 ( .A1(n5457), .A2(n5456), .A3(n5455), .ZN(u4_fi_ldz_1_) );
  NAND2_X2 U5640 ( .A1(n5458), .A2(fract_denorm[86]), .ZN(n5464) );
  INV_X4 U5641 ( .A(n8520), .ZN(n5459) );
  INV_X4 U5642 ( .A(n8525), .ZN(n5461) );
  NAND3_X4 U5643 ( .A1(n5464), .A2(n5463), .A3(n5462), .ZN(n5467) );
  NOR2_X4 U5644 ( .A1(n5467), .A2(n5466), .ZN(n5472) );
  INV_X4 U5645 ( .A(net59923), .ZN(net59921) );
  AOI22_X2 U5646 ( .A1(net59921), .A2(fract_denorm[70]), .B1(net59922), .B2(
        fract_denorm[54]), .ZN(n5471) );
  NAND4_X2 U5647 ( .A1(n5472), .A2(n5471), .A3(n5470), .A4(net59910), .ZN(
        u4_fi_ldz_2_) );
  INV_X4 U5648 ( .A(n5475), .ZN(n5474) );
  NAND2_X2 U5649 ( .A1(n5474), .A2(u4_fi_ldz_2_), .ZN(n5473) );
  INV_X4 U5650 ( .A(n5473), .ZN(n5496) );
  OAI21_X4 U5651 ( .B1(n5496), .B2(n4371), .A(net59901), .ZN(u4_fi_ldz_2a_4_)
         );
  INV_X4 U5652 ( .A(u4_fi_ldz_2_), .ZN(n5803) );
  NAND2_X2 U5653 ( .A1(n5475), .A2(n5803), .ZN(n5480) );
  NAND2_X2 U5654 ( .A1(n5480), .A2(n5473), .ZN(u4_fi_ldz_2a_2_) );
  NAND2_X2 U5655 ( .A1(n4527), .A2(u4_fi_ldz_1_), .ZN(n5811) );
  NAND2_X2 U5656 ( .A1(n5474), .A2(n5811), .ZN(u4_fi_ldz_mi1_1_) );
  INV_X4 U5657 ( .A(u4_fi_ldz_5_), .ZN(net57268) );
  NAND2_X2 U5658 ( .A1(net59209), .A2(n5475), .ZN(n5482) );
  INV_X4 U5659 ( .A(n5482), .ZN(n5476) );
  INV_X4 U5660 ( .A(u4_fi_ldz_4_), .ZN(n7168) );
  NAND2_X2 U5661 ( .A1(n5476), .A2(n7168), .ZN(n5479) );
  INV_X4 U5662 ( .A(n5477), .ZN(u4_fi_ldz_mi1_6_) );
  XNOR2_X2 U5663 ( .A(n5479), .B(u4_fi_ldz_5_), .ZN(u4_fi_ldz_mi1_5_) );
  NAND2_X2 U5664 ( .A1(n5482), .A2(u4_fi_ldz_4_), .ZN(n5478) );
  NAND2_X2 U5665 ( .A1(n5479), .A2(n5478), .ZN(u4_fi_ldz_mi1_4_) );
  NAND2_X2 U5666 ( .A1(n5480), .A2(u4_fi_ldz_3_), .ZN(n5481) );
  NAND2_X2 U5667 ( .A1(n5482), .A2(n5481), .ZN(u4_fi_ldz_mi1_3_) );
  INV_X4 U5668 ( .A(u4_exp_in_pl1_1_), .ZN(net59594) );
  INV_X4 U5669 ( .A(u4_exp_next_mi_1_), .ZN(net59892) );
  INV_X4 U5670 ( .A(net59891), .ZN(u4_exp_out1_1_) );
  NOR2_X4 U5671 ( .A1(n4852), .A2(net66839), .ZN(n5660) );
  NAND2_X2 U5672 ( .A1(n5660), .A2(n4378), .ZN(n5493) );
  INV_X4 U5673 ( .A(n5493), .ZN(n5483) );
  NAND3_X4 U5674 ( .A1(n5483), .A2(n4328), .A3(n4308), .ZN(n5490) );
  INV_X4 U5675 ( .A(n5490), .ZN(n5484) );
  NAND2_X2 U5676 ( .A1(n4384), .A2(n4327), .ZN(net59555) );
  INV_X4 U5677 ( .A(net59555), .ZN(net58701) );
  NAND2_X2 U5678 ( .A1(n5484), .A2(net58701), .ZN(n5489) );
  INV_X4 U5679 ( .A(n5489), .ZN(n5487) );
  INV_X4 U5680 ( .A(net66863), .ZN(net59551) );
  NAND2_X2 U5681 ( .A1(n5487), .A2(net59551), .ZN(n5486) );
  INV_X4 U5682 ( .A(n5486), .ZN(n5485) );
  INV_X4 U5683 ( .A(n4846), .ZN(n5534) );
  NAND2_X2 U5684 ( .A1(n5485), .A2(n5534), .ZN(net59886) );
  NAND2_X2 U5685 ( .A1(net58636), .A2(n4505), .ZN(net59553) );
  INV_X4 U5686 ( .A(net59888), .ZN(net59355) );
  OAI21_X4 U5687 ( .B1(net59355), .B2(net58636), .A(net59026), .ZN(
        u4_exp_in_mi1_10_) );
  OAI21_X4 U5688 ( .B1(n5485), .B2(n5534), .A(net59886), .ZN(u4_exp_in_mi1_8_)
         );
  NAND2_X2 U5689 ( .A1(exp_r[5]), .A2(n4848), .ZN(net59826) );
  NAND2_X2 U5690 ( .A1(n4848), .A2(n5490), .ZN(n5488) );
  OAI21_X4 U5691 ( .B1(n5491), .B2(n4328), .A(n5490), .ZN(u4_exp_in_mi1_4_) );
  XNOR2_X2 U5692 ( .A(n5493), .B(n4308), .ZN(n5492) );
  INV_X4 U5693 ( .A(n5492), .ZN(u4_exp_in_mi1_3_) );
  NOR2_X4 U5694 ( .A1(n5660), .A2(n4378), .ZN(n5652) );
  INV_X4 U5695 ( .A(n5652), .ZN(n5494) );
  NAND2_X2 U5696 ( .A1(n5494), .A2(n5493), .ZN(u4_exp_in_mi1_2_) );
  INV_X4 U5697 ( .A(n4852), .ZN(n6010) );
  INV_X4 U5698 ( .A(n5660), .ZN(n5495) );
  OAI21_X4 U5699 ( .B1(net43686), .B2(n6010), .A(n5495), .ZN(u4_exp_in_mi1_1_)
         );
  INV_X4 U5700 ( .A(u4_fi_ldz_3_), .ZN(n7172) );
  XNOR2_X2 U5701 ( .A(n7172), .B(n5496), .ZN(net44706) );
  INV_X4 U5702 ( .A(u4_fi_ldz_mi1_1_), .ZN(n7207) );
  NAND2_X2 U5703 ( .A1(div_opa_ldz_r2[0]), .A2(net43686), .ZN(n5512) );
  NAND2_X2 U5704 ( .A1(n4852), .A2(n5512), .ZN(n5508) );
  INV_X4 U5705 ( .A(net59721), .ZN(net59849) );
  NAND2_X2 U5706 ( .A1(div_opa_ldz_r2[2]), .A2(n4378), .ZN(net59723) );
  INV_X4 U5707 ( .A(net59723), .ZN(net59869) );
  NAND2_X2 U5708 ( .A1(n4851), .A2(n4324), .ZN(net59724) );
  OAI21_X4 U5709 ( .B1(net59849), .B2(net59869), .A(net59724), .ZN(net59868)
         );
  INV_X4 U5710 ( .A(net59868), .ZN(net59850) );
  NAND2_X2 U5711 ( .A1(div_opa_ldz_r2[3]), .A2(n4308), .ZN(net59722) );
  INV_X4 U5712 ( .A(net59865), .ZN(net59851) );
  NAND2_X2 U5713 ( .A1(div_opa_ldz_r2[4]), .A2(n4328), .ZN(net59719) );
  INV_X4 U5714 ( .A(net59719), .ZN(net59863) );
  NAND2_X2 U5715 ( .A1(n4850), .A2(n4387), .ZN(net59726) );
  OAI21_X4 U5716 ( .B1(net59851), .B2(net59863), .A(net59726), .ZN(n5498) );
  INV_X4 U5717 ( .A(n5498), .ZN(n5506) );
  NAND2_X2 U5718 ( .A1(n5506), .A2(n4327), .ZN(n5505) );
  INV_X4 U5719 ( .A(n5505), .ZN(n5504) );
  NAND2_X2 U5720 ( .A1(n5504), .A2(n4384), .ZN(n5628) );
  INV_X4 U5721 ( .A(n5628), .ZN(n5622) );
  NAND2_X2 U5722 ( .A1(n5622), .A2(n4380), .ZN(n5501) );
  INV_X4 U5723 ( .A(n5501), .ZN(n5500) );
  NAND2_X2 U5724 ( .A1(net59540), .A2(n5500), .ZN(n5518) );
  NAND2_X2 U5725 ( .A1(n5518), .A2(n5499), .ZN(u4_ldz_dif_10_) );
  XNOR2_X2 U5726 ( .A(net66871), .B(n5500), .ZN(n5694) );
  INV_X4 U5727 ( .A(n5694), .ZN(u4_ldz_dif_9_) );
  NAND2_X2 U5728 ( .A1(n4846), .A2(net66863), .ZN(net59443) );
  NAND2_X2 U5729 ( .A1(net59443), .A2(n5501), .ZN(n5623) );
  INV_X4 U5730 ( .A(n5623), .ZN(n5503) );
  NAND2_X2 U5731 ( .A1(n4846), .A2(n5628), .ZN(n5502) );
  NAND2_X2 U5732 ( .A1(n5503), .A2(n5502), .ZN(u4_ldz_dif_8_) );
  XNOR2_X2 U5733 ( .A(net66863), .B(n5628), .ZN(u4_ldz_dif_7_) );
  OAI21_X4 U5734 ( .B1(n5504), .B2(n4384), .A(n5628), .ZN(u4_ldz_dif_6_) );
  OAI21_X4 U5735 ( .B1(n5506), .B2(n4327), .A(n5505), .ZN(u4_ldz_dif_5_) );
  NAND2_X2 U5736 ( .A1(net59726), .A2(net59719), .ZN(n5572) );
  INV_X4 U5737 ( .A(n5572), .ZN(n5507) );
  XNOR2_X2 U5738 ( .A(net59851), .B(n5507), .ZN(u4_ldz_dif_4_) );
  NAND2_X2 U5739 ( .A1(net59717), .A2(net59722), .ZN(n5580) );
  INV_X4 U5740 ( .A(n5580), .ZN(n5582) );
  XNOR2_X2 U5741 ( .A(div_opa_ldz_r2[3]), .B(net66851), .ZN(n5579) );
  INV_X4 U5742 ( .A(n5579), .ZN(n5583) );
  MUX2_X2 U5743 ( .A(n5582), .B(n5583), .S(net59850), .Z(n5653) );
  INV_X4 U5744 ( .A(n5653), .ZN(u4_ldz_dif_3_) );
  NAND2_X2 U5745 ( .A1(net59724), .A2(net59723), .ZN(n5595) );
  INV_X4 U5746 ( .A(n5595), .ZN(n5597) );
  XNOR2_X2 U5747 ( .A(div_opa_ldz_r2[2]), .B(n4851), .ZN(n5594) );
  INV_X4 U5748 ( .A(n5594), .ZN(n5598) );
  MUX2_X2 U5749 ( .A(n5597), .B(n5598), .S(net59849), .Z(n5662) );
  INV_X4 U5750 ( .A(n5662), .ZN(u4_ldz_dif_2_) );
  NAND2_X2 U5751 ( .A1(div_opa_ldz_r2[1]), .A2(n6010), .ZN(n5568) );
  MUX2_X2 U5752 ( .A(n4325), .B(n5568), .S(n5512), .Z(n5511) );
  INV_X4 U5753 ( .A(n5508), .ZN(n5509) );
  NAND2_X2 U5754 ( .A1(n5509), .A2(n4377), .ZN(n5510) );
  NAND2_X2 U5755 ( .A1(n5511), .A2(n5510), .ZN(u4_ldz_dif_1_) );
  NAND2_X2 U5756 ( .A1(net66839), .A2(n4381), .ZN(n5612) );
  NAND2_X2 U5757 ( .A1(n5612), .A2(n5512), .ZN(u4_ldz_dif_0_) );
  NAND2_X2 U5758 ( .A1(prod[0]), .A2(net66929), .ZN(n5515) );
  NAND2_X2 U5759 ( .A1(fract_i2f[0]), .A2(net63085), .ZN(n5514) );
  NAND2_X2 U5760 ( .A1(quo[2]), .A2(net66910), .ZN(n5513) );
  INV_X4 U5761 ( .A(net58674), .ZN(net59835) );
  NAND2_X2 U5762 ( .A1(net59835), .A2(net63289), .ZN(n2442) );
  INV_X4 U5763 ( .A(n2442), .ZN(net59731) );
  NAND2_X2 U5764 ( .A1(u4_exp_out_8_), .A2(net59731), .ZN(n5539) );
  NAND2_X2 U5765 ( .A1(net58674), .A2(net63289), .ZN(net57230) );
  INV_X4 U5766 ( .A(net57230), .ZN(net59565) );
  NAND2_X2 U5767 ( .A1(net59565), .A2(u4_exp_in_mi1_8_), .ZN(n5538) );
  NAND2_X2 U5768 ( .A1(n4851), .A2(n4852), .ZN(n5587) );
  INV_X4 U5769 ( .A(n5587), .ZN(n5516) );
  NAND2_X2 U5770 ( .A1(n5516), .A2(net66851), .ZN(n5563) );
  INV_X4 U5771 ( .A(n5563), .ZN(n5517) );
  NAND2_X2 U5772 ( .A1(n5517), .A2(n4850), .ZN(n5684) );
  NOR2_X4 U5773 ( .A1(n5684), .A2(n4327), .ZN(n5548) );
  NAND3_X4 U5774 ( .A1(net66863), .A2(n4848), .A3(n5548), .ZN(n5520) );
  INV_X4 U5775 ( .A(n5518), .ZN(n5519) );
  NAND3_X4 U5776 ( .A1(net59026), .A2(net59070), .A3(n5519), .ZN(net58662) );
  INV_X4 U5777 ( .A(net59674), .ZN(net58681) );
  NAND3_X4 U5778 ( .A1(net58662), .A2(net63291), .A3(net58681), .ZN(n7189) );
  INV_X4 U5779 ( .A(n5520), .ZN(n5681) );
  MUX2_X2 U5780 ( .A(n5522), .B(n5521), .S(n4846), .Z(n5536) );
  INV_X4 U5781 ( .A(net59826), .ZN(net59678) );
  NAND2_X2 U5782 ( .A1(div_opa_ldz_r2[0]), .A2(net66839), .ZN(n5613) );
  NAND2_X2 U5783 ( .A1(div_opa_ldz_r2[1]), .A2(n4852), .ZN(n5523) );
  INV_X4 U5784 ( .A(n5525), .ZN(n5596) );
  NAND2_X2 U5785 ( .A1(n4851), .A2(div_opa_ldz_r2[2]), .ZN(n5526) );
  OAI21_X4 U5786 ( .B1(n5596), .B2(n5527), .A(n5526), .ZN(n5528) );
  INV_X4 U5787 ( .A(n5528), .ZN(n5581) );
  NAND2_X2 U5788 ( .A1(net66851), .A2(div_opa_ldz_r2[3]), .ZN(n5529) );
  OAI21_X4 U5789 ( .B1(n5581), .B2(n5530), .A(n5529), .ZN(n5564) );
  INV_X4 U5790 ( .A(n5564), .ZN(n5533) );
  NAND2_X2 U5791 ( .A1(n4850), .A2(div_opa_ldz_r2[4]), .ZN(n5531) );
  OAI21_X4 U5792 ( .B1(n5533), .B2(n5532), .A(n5531), .ZN(net59792) );
  XNOR2_X2 U5793 ( .A(net59812), .B(n5534), .ZN(net59435) );
  NOR2_X4 U5794 ( .A1(n5536), .A2(n5535), .ZN(n5537) );
  NAND3_X4 U5795 ( .A1(n5539), .A2(n5538), .A3(n5537), .ZN(u4_shift_right[8])
         );
  INV_X4 U5796 ( .A(n5548), .ZN(n5547) );
  MUX2_X2 U5797 ( .A(n5541), .B(n5540), .S(net66863), .Z(n5544) );
  INV_X4 U5798 ( .A(u4_exp_in_mi1_7_), .ZN(n5542) );
  NOR2_X4 U5799 ( .A1(net57230), .A2(n5542), .ZN(n5543) );
  NOR2_X4 U5800 ( .A1(n5544), .A2(n5543), .ZN(n5546) );
  NAND2_X2 U5801 ( .A1(u4_exp_out_7_), .A2(net59731), .ZN(n5545) );
  MUX2_X2 U5802 ( .A(n5550), .B(n5549), .S(n4848), .Z(n5551) );
  INV_X4 U5803 ( .A(n5551), .ZN(n5555) );
  NAND2_X2 U5804 ( .A1(exp_r[5]), .A2(n4384), .ZN(n5633) );
  INV_X4 U5805 ( .A(net59792), .ZN(net59785) );
  MUX2_X2 U5806 ( .A(n5633), .B(n4384), .S(net59785), .Z(n5552) );
  NAND2_X2 U5807 ( .A1(n4848), .A2(n4327), .ZN(n5634) );
  NAND2_X2 U5808 ( .A1(n5552), .A2(n5634), .ZN(n5718) );
  AOI22_X2 U5809 ( .A1(u4_exp_in_mi1_6_), .A2(net59565), .B1(net59427), .B2(
        n5718), .ZN(n5554) );
  NAND2_X2 U5810 ( .A1(u4_exp_out_6_), .A2(net59731), .ZN(n5553) );
  NAND2_X2 U5811 ( .A1(net87237), .A2(net59731), .ZN(n5562) );
  NAND2_X2 U5812 ( .A1(n4385), .A2(net59565), .ZN(n5561) );
  XNOR2_X2 U5813 ( .A(n5684), .B(n4327), .ZN(n5556) );
  NOR2_X4 U5814 ( .A1(n4843), .A2(n5556), .ZN(n5559) );
  XNOR2_X2 U5815 ( .A(exp_r[5]), .B(net59785), .ZN(n5720) );
  INV_X4 U5816 ( .A(n5720), .ZN(n5557) );
  NOR2_X4 U5817 ( .A1(n5559), .A2(n5558), .ZN(n5560) );
  NAND3_X2 U5818 ( .A1(n5562), .A2(n5561), .A3(n5560), .ZN(u4_shift_right[5])
         );
  XNOR2_X2 U5819 ( .A(n4850), .B(n5563), .ZN(n5567) );
  INV_X4 U5820 ( .A(n4843), .ZN(n5566) );
  XNOR2_X2 U5821 ( .A(n5572), .B(n5564), .ZN(n5714) );
  NOR2_X4 U5822 ( .A1(n5714), .A2(net57241), .ZN(n5565) );
  INV_X4 U5823 ( .A(n5612), .ZN(n5615) );
  INV_X4 U5824 ( .A(n5570), .ZN(n5593) );
  OAI21_X4 U5825 ( .B1(n4658), .B2(n5593), .A(net59723), .ZN(n5577) );
  INV_X4 U5826 ( .A(net59722), .ZN(net59765) );
  INV_X4 U5827 ( .A(net58662), .ZN(net59768) );
  NAND3_X4 U5828 ( .A1(net59768), .A2(net63291), .A3(net58681), .ZN(n7191) );
  INV_X4 U5829 ( .A(n7191), .ZN(n5571) );
  OAI211_X2 U5830 ( .C1(n4402), .C2(net59765), .A(n5572), .B(n5571), .ZN(n5575) );
  NAND2_X2 U5831 ( .A1(net59565), .A2(u4_exp_in_mi1_4_), .ZN(n5574) );
  NAND2_X2 U5832 ( .A1(net96080), .A2(net59731), .ZN(n5573) );
  NAND4_X2 U5833 ( .A1(n5576), .A2(n5575), .A3(n5574), .A4(n5573), .ZN(
        u4_shift_right[4]) );
  INV_X4 U5834 ( .A(n7191), .ZN(n5586) );
  INV_X4 U5835 ( .A(n5577), .ZN(n5578) );
  MUX2_X2 U5836 ( .A(n5580), .B(n5579), .S(n5578), .Z(n5585) );
  MUX2_X2 U5837 ( .A(n5583), .B(n5582), .S(n5581), .Z(n5716) );
  AOI21_X4 U5838 ( .B1(n5586), .B2(n5585), .A(n5584), .ZN(n5592) );
  XNOR2_X2 U5839 ( .A(n5587), .B(net66851), .ZN(n5588) );
  NAND2_X2 U5840 ( .A1(n5588), .A2(n5602), .ZN(n5591) );
  NAND2_X2 U5841 ( .A1(u4_exp_in_mi1_3_), .A2(net59565), .ZN(n5590) );
  NAND2_X2 U5842 ( .A1(u4_exp_out_3_), .A2(net59731), .ZN(n5589) );
  NAND4_X2 U5843 ( .A1(n5592), .A2(n5591), .A3(n5590), .A4(n5589), .ZN(
        u4_shift_right[3]) );
  MUX2_X2 U5844 ( .A(n5595), .B(n5594), .S(n5593), .Z(n5600) );
  MUX2_X2 U5845 ( .A(n5598), .B(n5597), .S(n5596), .Z(n5715) );
  AOI21_X4 U5846 ( .B1(n5571), .B2(n5600), .A(n5599), .ZN(n5606) );
  INV_X4 U5847 ( .A(n4843), .ZN(n5602) );
  XOR2_X2 U5848 ( .A(n4851), .B(n4852), .Z(n5601) );
  NAND2_X2 U5849 ( .A1(n5602), .A2(n5601), .ZN(n5605) );
  NAND2_X2 U5850 ( .A1(net59565), .A2(u4_exp_in_mi1_2_), .ZN(n5604) );
  NAND2_X2 U5851 ( .A1(u4_exp_out_2_), .A2(net59731), .ZN(n5603) );
  NAND4_X2 U5852 ( .A1(n5606), .A2(n5605), .A3(n5604), .A4(n5603), .ZN(
        u4_shift_right[2]) );
  NAND2_X2 U5853 ( .A1(net59540), .A2(n4380), .ZN(net58688) );
  AOI22_X2 U5854 ( .A1(u4_div_exp3[1]), .A2(net58719), .B1(u4_div_exp1_1_), 
        .B2(net58718), .ZN(n5607) );
  NAND2_X2 U5855 ( .A1(n5973), .A2(net63293), .ZN(n5609) );
  INV_X4 U5856 ( .A(net33546), .ZN(net59698) );
  NAND3_X4 U5857 ( .A1(net59697), .A2(net59698), .A3(net59699), .ZN(net58644)
         );
  NAND2_X2 U5858 ( .A1(net58780), .A2(net58644), .ZN(net57276) );
  INV_X4 U5859 ( .A(net57276), .ZN(net57252) );
  NAND2_X2 U5860 ( .A1(net57252), .A2(u4_fi_ldz_mi1_1_), .ZN(n5608) );
  AOI21_X4 U5861 ( .B1(net59696), .B2(net59026), .A(net59008), .ZN(net59260)
         );
  INV_X4 U5862 ( .A(net58644), .ZN(net59695) );
  NAND2_X2 U5863 ( .A1(n2402), .A2(n7162), .ZN(net59694) );
  NAND3_X4 U5864 ( .A1(n5609), .A2(n5608), .A3(net59693), .ZN(u4_exp_out_1_)
         );
  INV_X4 U5865 ( .A(u4_exp_in_mi1_1_), .ZN(net59588) );
  INV_X4 U5866 ( .A(n5613), .ZN(n5610) );
  NAND2_X2 U5867 ( .A1(net59427), .A2(n5610), .ZN(n5611) );
  NAND2_X2 U5868 ( .A1(net59427), .A2(n5613), .ZN(n5614) );
  OAI21_X4 U5869 ( .B1(n5615), .B2(n7191), .A(n5614), .ZN(n5616) );
  MUX2_X2 U5870 ( .A(n5617), .B(n5616), .S(n4325), .Z(n5619) );
  NAND3_X4 U5871 ( .A1(n4850), .A2(net66851), .A3(n5652), .ZN(n5640) );
  INV_X4 U5872 ( .A(n5640), .ZN(n5632) );
  NAND2_X2 U5873 ( .A1(n5632), .A2(net59678), .ZN(n5627) );
  NAND2_X2 U5874 ( .A1(n4380), .A2(n5627), .ZN(n5676) );
  OAI211_X2 U5875 ( .C1(n4383), .C2(n5627), .A(net59443), .B(n5676), .ZN(
        u4_f2i_shft_8_) );
  NOR2_X4 U5876 ( .A1(net59674), .A2(n5620), .ZN(n5621) );
  NOR2_X4 U5877 ( .A1(n4534), .A2(n5621), .ZN(n5646) );
  NAND3_X4 U5878 ( .A1(n5646), .A2(net63291), .A3(net59026), .ZN(net59543) );
  NOR3_X4 U5879 ( .A1(n4534), .A2(net66835), .A3(net59070), .ZN(net58700) );
  NAND2_X2 U5880 ( .A1(net58792), .A2(net58935), .ZN(net59347) );
  NAND2_X2 U5881 ( .A1(net58781), .A2(u4_f2i_shft_8_), .ZN(n5624) );
  XNOR2_X2 U5882 ( .A(n5627), .B(net59551), .ZN(u4_f2i_shft_7_) );
  INV_X4 U5883 ( .A(u4_exp_in_pl1_7_), .ZN(n5791) );
  MUX2_X2 U5884 ( .A(n5630), .B(n5629), .S(net66863), .Z(n5631) );
  MUX2_X2 U5885 ( .A(n4384), .B(n5633), .S(n5632), .Z(n5635) );
  NAND2_X2 U5886 ( .A1(n5635), .A2(n5634), .ZN(u4_f2i_shft_6_) );
  INV_X4 U5887 ( .A(net59541), .ZN(net59635) );
  AOI22_X2 U5888 ( .A1(u4_f2i_shft_6_), .A2(net58781), .B1(net59635), .B2(
        n4848), .ZN(n5639) );
  NAND2_X2 U5889 ( .A1(u4_ldz_dif_6_), .A2(net59645), .ZN(n5638) );
  AOI21_X4 U5890 ( .B1(n5636), .B2(net59644), .A(net58780), .ZN(net59642) );
  AOI22_X2 U5891 ( .A1(n4329), .A2(net58781), .B1(net59635), .B2(exp_r[5]), 
        .ZN(n5644) );
  NAND2_X2 U5892 ( .A1(u4_ldz_dif_5_), .A2(net59632), .ZN(n5641) );
  NAND4_X2 U5893 ( .A1(n5644), .A2(n5643), .A3(n5642), .A4(n5641), .ZN(
        u4_shift_left[5]) );
  NAND2_X2 U5894 ( .A1(n5652), .A2(net66851), .ZN(n5645) );
  AOI22_X2 U5895 ( .A1(n4295), .A2(net58781), .B1(u4_ldz_dif_4_), .B2(net59626), .ZN(n5651) );
  NAND2_X2 U5896 ( .A1(net59635), .A2(n4850), .ZN(n5650) );
  NAND4_X2 U5897 ( .A1(n5651), .A2(n5650), .A3(n5649), .A4(n5648), .ZN(
        u4_shift_left[4]) );
  XNOR2_X2 U5898 ( .A(net66851), .B(n5652), .ZN(n5779) );
  AOI22_X2 U5899 ( .A1(net59600), .A2(div_opa_ldz_r2[3]), .B1(net59578), .B2(
        u4_fi_ldz_3_), .ZN(n5657) );
  NAND3_X4 U5900 ( .A1(n5659), .A2(n5658), .A3(n5657), .ZN(u4_shift_left[3])
         );
  XNOR2_X2 U5901 ( .A(n4851), .B(n5660), .ZN(u4_f2i_shft_2_) );
  INV_X4 U5902 ( .A(u4_f2i_shft_2_), .ZN(n5661) );
  NAND2_X2 U5903 ( .A1(net59635), .A2(n4851), .ZN(n5667) );
  INV_X4 U5904 ( .A(net59579), .ZN(net59600) );
  NAND4_X2 U5905 ( .A1(n5668), .A2(n5667), .A3(n5666), .A4(n5665), .ZN(
        u4_shift_left[2]) );
  NAND2_X2 U5906 ( .A1(net59600), .A2(div_opa_ldz_r2[1]), .ZN(n5674) );
  INV_X4 U5907 ( .A(u4_ldz_dif_1_), .ZN(n5669) );
  NAND4_X2 U5908 ( .A1(n5675), .A2(n5674), .A3(net59582), .A4(n5673), .ZN(
        u4_shift_left[1]) );
  INV_X4 U5909 ( .A(n5676), .ZN(n5690) );
  NAND2_X2 U5910 ( .A1(n5690), .A2(net59540), .ZN(n5677) );
  OAI21_X4 U5911 ( .B1(n5678), .B2(net58636), .A(n5677), .ZN(u4_f2i_shft_10_)
         );
  NAND2_X2 U5912 ( .A1(net58645), .A2(net66835), .ZN(net59309) );
  NAND2_X2 U5913 ( .A1(net59309), .A2(net63289), .ZN(n5680) );
  NAND2_X2 U5914 ( .A1(net59565), .A2(u4_exp_in_mi1_11_), .ZN(n5679) );
  NAND3_X4 U5915 ( .A1(n5680), .A2(net59563), .A3(n5679), .ZN(n5700) );
  INV_X4 U5916 ( .A(n5872), .ZN(n5689) );
  NAND2_X2 U5917 ( .A1(n4846), .A2(n5681), .ZN(n5682) );
  INV_X4 U5918 ( .A(n5682), .ZN(n7188) );
  NAND2_X2 U5919 ( .A1(n7188), .A2(net66871), .ZN(n7179) );
  OAI21_X4 U5920 ( .B1(n5683), .B2(n7179), .A(net58636), .ZN(net58808) );
  INV_X4 U5921 ( .A(n5684), .ZN(n5685) );
  NAND2_X2 U5922 ( .A1(opas_r2), .A2(n5871), .ZN(n5688) );
  OAI21_X4 U5923 ( .B1(n5689), .B2(net58808), .A(n5688), .ZN(n5964) );
  INV_X4 U5924 ( .A(n5964), .ZN(n5692) );
  INV_X4 U5925 ( .A(u4_f2i_shft_10_), .ZN(n5691) );
  XNOR2_X2 U5926 ( .A(net66871), .B(n5690), .ZN(n5778) );
  NAND2_X2 U5927 ( .A1(net58781), .A2(n5693), .ZN(n5698) );
  NAND4_X2 U5928 ( .A1(n5699), .A2(n5700), .A3(n5698), .A4(n5697), .ZN(
        net57285) );
  INV_X4 U5929 ( .A(u4_N6119), .ZN(n5704) );
  INV_X4 U5930 ( .A(n5700), .ZN(n5702) );
  INV_X4 U5931 ( .A(u4_N5904), .ZN(n5701) );
  NAND2_X2 U5932 ( .A1(n5702), .A2(n5701), .ZN(net59531) );
  INV_X4 U5933 ( .A(net59531), .ZN(net44903) );
  NAND2_X2 U5934 ( .A1(u4_N6011), .A2(net63325), .ZN(n5703) );
  OAI21_X4 U5935 ( .B1(net57285), .B2(n5704), .A(n5703), .ZN(u4_fract_out_51_)
         );
  INV_X4 U5936 ( .A(n2521), .ZN(u4_fract_out_50_) );
  INV_X4 U5937 ( .A(n3626), .ZN(u4_fract_out_49_) );
  INV_X4 U5938 ( .A(n3629), .ZN(u4_fract_out_48_) );
  INV_X4 U5939 ( .A(n2522), .ZN(u4_fract_out_47_) );
  INV_X4 U5940 ( .A(n2523), .ZN(u4_fract_out_46_) );
  INV_X4 U5941 ( .A(n2524), .ZN(u4_fract_out_45_) );
  INV_X4 U5942 ( .A(n3636), .ZN(u4_fract_out_44_) );
  INV_X4 U5943 ( .A(n3638), .ZN(u4_fract_out_43_) );
  INV_X4 U5944 ( .A(n3641), .ZN(u4_fract_out_42_) );
  INV_X4 U5945 ( .A(n3644), .ZN(u4_fract_out_41_) );
  INV_X4 U5946 ( .A(n2525), .ZN(u4_fract_out_40_) );
  INV_X4 U5947 ( .A(n2527), .ZN(u4_fract_out_39_) );
  INV_X4 U5948 ( .A(n3650), .ZN(u4_fract_out_38_) );
  INV_X4 U5949 ( .A(n3654), .ZN(u4_fract_out_36_) );
  INV_X4 U5950 ( .A(n2528), .ZN(u4_fract_out_35_) );
  INV_X4 U5951 ( .A(n2529), .ZN(u4_fract_out_34_) );
  INV_X4 U5952 ( .A(n3662), .ZN(u4_fract_out_32_) );
  INV_X4 U5953 ( .A(n3664), .ZN(u4_fract_out_31_) );
  INV_X4 U5954 ( .A(n3666), .ZN(u4_fract_out_30_) );
  INV_X4 U5955 ( .A(n2531), .ZN(u4_fract_out_29_) );
  INV_X4 U5956 ( .A(n2532), .ZN(u4_fract_out_28_) );
  INV_X4 U5957 ( .A(n3675), .ZN(u4_fract_out_26_) );
  INV_X4 U5958 ( .A(n3677), .ZN(u4_fract_out_25_) );
  INV_X4 U5959 ( .A(n3679), .ZN(u4_fract_out_24_) );
  INV_X4 U5960 ( .A(n2534), .ZN(u4_fract_out_23_) );
  INV_X4 U5961 ( .A(n2535), .ZN(u4_fract_out_22_) );
  INV_X4 U5962 ( .A(n2536), .ZN(u4_fract_out_21_) );
  INV_X4 U5963 ( .A(n3687), .ZN(u4_fract_out_20_) );
  INV_X4 U5964 ( .A(n3689), .ZN(u4_fract_out_19_) );
  INV_X4 U5965 ( .A(n3691), .ZN(u4_fract_out_18_) );
  INV_X4 U5966 ( .A(n2537), .ZN(u4_fract_out_17_) );
  INV_X4 U5967 ( .A(n2538), .ZN(u4_fract_out_16_) );
  INV_X4 U5968 ( .A(n2539), .ZN(u4_fract_out_15_) );
  INV_X4 U5969 ( .A(n3699), .ZN(u4_fract_out_14_) );
  INV_X4 U5970 ( .A(n3702), .ZN(u4_fract_out_13_) );
  INV_X4 U5971 ( .A(n2540), .ZN(u4_fract_out_11_) );
  INV_X4 U5972 ( .A(n2541), .ZN(u4_fract_out_10_) );
  INV_X4 U5973 ( .A(n3709), .ZN(u4_fract_out_9_) );
  INV_X4 U5974 ( .A(n3712), .ZN(u4_fract_out_8_) );
  INV_X4 U5975 ( .A(n3715), .ZN(u4_fract_out_7_) );
  INV_X4 U5976 ( .A(n3717), .ZN(u4_fract_out_6_) );
  INV_X4 U5977 ( .A(n2519), .ZN(u4_fract_out_5_) );
  INV_X4 U5978 ( .A(n3720), .ZN(u4_fract_out_4_) );
  INV_X4 U5979 ( .A(n2526), .ZN(u4_fract_out_3_) );
  INV_X4 U5980 ( .A(n3724), .ZN(u4_fract_out_2_) );
  INV_X4 U5981 ( .A(n3727), .ZN(u4_fract_out_1_) );
  INV_X4 U5982 ( .A(n3731), .ZN(u4_fract_out_0_) );
  NOR2_X4 U5983 ( .A1(n5706), .A2(n5705), .ZN(net59504) );
  NAND2_X2 U5984 ( .A1(n3662), .A2(n2533), .ZN(n5707) );
  NOR4_X2 U5985 ( .A1(n3888), .A2(u4_fract_out_28_), .A3(u4_fract_out_29_), 
        .A4(n5707), .ZN(net59505) );
  NOR4_X2 U5986 ( .A1(n5711), .A2(n5710), .A3(n5709), .A4(n5708), .ZN(net59506) );
  INV_X4 U5987 ( .A(net59443), .ZN(net59442) );
  XNOR2_X2 U5988 ( .A(net66875), .B(n5717), .ZN(n7183) );
  INV_X4 U5989 ( .A(n7183), .ZN(n5719) );
  INV_X4 U5990 ( .A(net59435), .ZN(net59430) );
  XNOR2_X2 U5991 ( .A(net59433), .B(n4505), .ZN(net57240) );
  NOR4_X2 U5992 ( .A1(remainder[17]), .A2(remainder[16]), .A3(remainder[15]), 
        .A4(remainder[14]), .ZN(n5725) );
  NOR3_X4 U5993 ( .A1(remainder[20]), .A2(remainder[19]), .A3(remainder[18]), 
        .ZN(n5724) );
  NOR3_X4 U5994 ( .A1(remainder[23]), .A2(remainder[22]), .A3(remainder[21]), 
        .ZN(n5723) );
  NOR3_X4 U5995 ( .A1(remainder[26]), .A2(remainder[25]), .A3(remainder[24]), 
        .ZN(n5722) );
  NAND4_X2 U5996 ( .A1(n5725), .A2(n5724), .A3(n5723), .A4(n5722), .ZN(n5734)
         );
  NOR2_X4 U5997 ( .A1(remainder[8]), .A2(remainder[7]), .ZN(n5728) );
  NOR2_X4 U5998 ( .A1(remainder[10]), .A2(remainder[9]), .ZN(n5727) );
  NOR2_X4 U5999 ( .A1(remainder[12]), .A2(remainder[11]), .ZN(n5726) );
  NAND4_X2 U6000 ( .A1(n5728), .A2(n5727), .A3(n5726), .A4(n4408), .ZN(n5733)
         );
  NOR2_X4 U6001 ( .A1(remainder[1]), .A2(remainder[0]), .ZN(n5731) );
  NOR2_X4 U6002 ( .A1(remainder[3]), .A2(remainder[2]), .ZN(n5730) );
  NOR2_X4 U6003 ( .A1(remainder[5]), .A2(remainder[4]), .ZN(n5729) );
  NAND4_X2 U6004 ( .A1(n5731), .A2(n5730), .A3(n5729), .A4(n4409), .ZN(n5732)
         );
  NOR3_X4 U6005 ( .A1(n5734), .A2(n5733), .A3(n5732), .ZN(n5777) );
  NOR4_X2 U6006 ( .A1(remainder[44]), .A2(remainder[43]), .A3(remainder[42]), 
        .A4(remainder[41]), .ZN(n5738) );
  NOR3_X4 U6007 ( .A1(remainder[47]), .A2(remainder[46]), .A3(remainder[45]), 
        .ZN(n5737) );
  NOR3_X4 U6008 ( .A1(remainder[50]), .A2(remainder[49]), .A3(remainder[48]), 
        .ZN(n5736) );
  NAND4_X2 U6009 ( .A1(n5738), .A2(n5737), .A3(n5736), .A4(n5735), .ZN(n5747)
         );
  NOR2_X4 U6010 ( .A1(remainder[39]), .A2(remainder[38]), .ZN(n5739) );
  NAND4_X2 U6011 ( .A1(n5741), .A2(n5740), .A3(n5739), .A4(n4410), .ZN(n5746)
         );
  NOR2_X4 U6012 ( .A1(remainder[28]), .A2(remainder[27]), .ZN(n5744) );
  NOR2_X4 U6013 ( .A1(remainder[30]), .A2(remainder[29]), .ZN(n5743) );
  NAND4_X2 U6014 ( .A1(n5744), .A2(n5743), .A3(n5742), .A4(n4411), .ZN(n5745)
         );
  NOR3_X4 U6015 ( .A1(n5747), .A2(n5746), .A3(n5745), .ZN(n5776) );
  NOR4_X2 U6016 ( .A1(remainder[71]), .A2(remainder[70]), .A3(remainder[69]), 
        .A4(remainder[68]), .ZN(n5751) );
  NOR3_X4 U6017 ( .A1(remainder[74]), .A2(remainder[73]), .A3(remainder[72]), 
        .ZN(n5750) );
  NOR3_X4 U6018 ( .A1(remainder[77]), .A2(remainder[76]), .A3(remainder[75]), 
        .ZN(n5749) );
  NOR3_X4 U6019 ( .A1(remainder[80]), .A2(remainder[79]), .A3(remainder[78]), 
        .ZN(n5748) );
  NAND4_X2 U6020 ( .A1(n5751), .A2(n5750), .A3(n5749), .A4(n5748), .ZN(n5760)
         );
  NOR2_X4 U6021 ( .A1(remainder[62]), .A2(remainder[61]), .ZN(n5754) );
  NOR2_X4 U6022 ( .A1(remainder[64]), .A2(remainder[63]), .ZN(n5753) );
  NOR2_X4 U6023 ( .A1(remainder[66]), .A2(remainder[65]), .ZN(n5752) );
  NAND4_X2 U6024 ( .A1(n5754), .A2(n5753), .A3(n5752), .A4(n4412), .ZN(n5759)
         );
  NOR2_X4 U6025 ( .A1(remainder[57]), .A2(remainder[56]), .ZN(n5756) );
  NOR2_X4 U6026 ( .A1(remainder[59]), .A2(remainder[58]), .ZN(n5755) );
  NAND4_X2 U6027 ( .A1(n5757), .A2(n5756), .A3(n5755), .A4(n4413), .ZN(n5758)
         );
  NOR3_X4 U6028 ( .A1(n5760), .A2(n5759), .A3(n5758), .ZN(n5775) );
  NOR4_X2 U6029 ( .A1(remainder[98]), .A2(remainder[97]), .A3(remainder[96]), 
        .A4(remainder[95]), .ZN(n5764) );
  NOR3_X4 U6030 ( .A1(remainder[101]), .A2(remainder[100]), .A3(remainder[99]), 
        .ZN(n5763) );
  NOR3_X4 U6031 ( .A1(remainder[104]), .A2(remainder[103]), .A3(remainder[102]), .ZN(n5762) );
  NOR3_X4 U6032 ( .A1(remainder[107]), .A2(remainder[106]), .A3(remainder[105]), .ZN(n5761) );
  NAND4_X2 U6033 ( .A1(n5764), .A2(n5763), .A3(n5762), .A4(n5761), .ZN(n5773)
         );
  NOR2_X4 U6034 ( .A1(remainder[89]), .A2(remainder[88]), .ZN(n5767) );
  NOR2_X4 U6035 ( .A1(remainder[91]), .A2(remainder[90]), .ZN(n5766) );
  NOR2_X4 U6036 ( .A1(remainder[93]), .A2(remainder[92]), .ZN(n5765) );
  NAND4_X2 U6037 ( .A1(n5767), .A2(n5766), .A3(n5765), .A4(n4414), .ZN(n5772)
         );
  NOR2_X4 U6038 ( .A1(remainder[82]), .A2(remainder[81]), .ZN(n5770) );
  NOR2_X4 U6039 ( .A1(remainder[84]), .A2(remainder[83]), .ZN(n5769) );
  NOR2_X4 U6040 ( .A1(remainder[86]), .A2(remainder[85]), .ZN(n5768) );
  NAND4_X2 U6041 ( .A1(n5770), .A2(n5769), .A3(n5768), .A4(n4415), .ZN(n5771)
         );
  NOR3_X4 U6042 ( .A1(n5773), .A2(n5772), .A3(n5771), .ZN(n5774) );
  NAND4_X2 U6043 ( .A1(n5777), .A2(n5776), .A3(n5775), .A4(n5774), .ZN(
        net58682) );
  NAND2_X2 U6044 ( .A1(net66835), .A2(net58644), .ZN(net59349) );
  NAND2_X2 U6045 ( .A1(net59355), .A2(net66875), .ZN(net59032) );
  INV_X4 U6046 ( .A(net59341), .ZN(net59338) );
  INV_X4 U6047 ( .A(net59309), .ZN(net58643) );
  INV_X4 U6048 ( .A(n5778), .ZN(u4_f2i_shft_9_) );
  INV_X4 U6049 ( .A(n5779), .ZN(u4_f2i_shft_3_) );
  MUX2_X2 U6050 ( .A(u4_exp_in_pl1_10_), .B(u4_exp_next_mi_10_), .S(net63221), 
        .Z(net59283) );
  INV_X4 U6051 ( .A(u4_div_exp1_10_), .ZN(n5797) );
  INV_X4 U6052 ( .A(u4_exp_in_pl1_5_), .ZN(n5781) );
  INV_X4 U6053 ( .A(u4_exp_next_mi_5_), .ZN(n5780) );
  MUX2_X2 U6054 ( .A(n5781), .B(n5780), .S(net63221), .Z(net44770) );
  INV_X4 U6055 ( .A(u4_exp_in_pl1_2_), .ZN(n5783) );
  INV_X4 U6056 ( .A(u4_exp_next_mi_2_), .ZN(n5782) );
  MUX2_X2 U6057 ( .A(n5783), .B(n5782), .S(net63221), .Z(n7206) );
  INV_X4 U6058 ( .A(n7206), .ZN(n5968) );
  INV_X4 U6059 ( .A(net59296), .ZN(net58767) );
  NOR2_X4 U6060 ( .A1(n5968), .A2(net58767), .ZN(n5989) );
  INV_X4 U6061 ( .A(u4_exp_in_pl1_3_), .ZN(n5784) );
  INV_X4 U6062 ( .A(u4_exp_next_mi_3_), .ZN(net59295) );
  MUX2_X2 U6063 ( .A(n5784), .B(net59295), .S(net63221), .Z(n7205) );
  NAND2_X2 U6064 ( .A1(n5989), .A2(n7205), .ZN(n5983) );
  INV_X4 U6065 ( .A(n5983), .ZN(n5991) );
  INV_X4 U6066 ( .A(u4_exp_in_pl1_4_), .ZN(n5786) );
  INV_X4 U6067 ( .A(u4_exp_next_mi_4_), .ZN(n5785) );
  MUX2_X2 U6068 ( .A(n5786), .B(n5785), .S(net63221), .Z(n7204) );
  NAND2_X2 U6069 ( .A1(n5991), .A2(n7204), .ZN(net58733) );
  INV_X4 U6070 ( .A(u4_exp_in_pl1_6_), .ZN(n5788) );
  INV_X4 U6071 ( .A(u4_exp_next_mi_6_), .ZN(n5787) );
  MUX2_X2 U6072 ( .A(n5788), .B(n5787), .S(net63221), .Z(n7203) );
  NAND2_X2 U6073 ( .A1(net58728), .A2(n7203), .ZN(n5789) );
  INV_X4 U6074 ( .A(n5789), .ZN(n5998) );
  INV_X4 U6075 ( .A(u4_exp_next_mi_7_), .ZN(n5790) );
  MUX2_X2 U6076 ( .A(n5791), .B(n5790), .S(net63221), .Z(n7202) );
  NAND2_X2 U6077 ( .A1(n5998), .A2(n7202), .ZN(n5975) );
  INV_X4 U6078 ( .A(n5975), .ZN(n6000) );
  INV_X4 U6079 ( .A(u4_exp_in_pl1_8_), .ZN(n5792) );
  INV_X4 U6080 ( .A(u4_exp_next_mi_8_), .ZN(n5817) );
  MUX2_X2 U6081 ( .A(n5792), .B(n5817), .S(net63221), .Z(n7201) );
  NAND2_X2 U6082 ( .A1(n6000), .A2(n7201), .ZN(n5799) );
  INV_X4 U6083 ( .A(n5799), .ZN(n5974) );
  INV_X4 U6084 ( .A(u4_exp_in_pl1_9_), .ZN(n5793) );
  INV_X4 U6085 ( .A(u4_exp_next_mi_9_), .ZN(n5857) );
  MUX2_X2 U6086 ( .A(n5793), .B(n5857), .S(net63221), .Z(net59270) );
  NAND2_X2 U6087 ( .A1(n5974), .A2(net59270), .ZN(n5794) );
  INV_X4 U6088 ( .A(n5794), .ZN(n5798) );
  XNOR2_X2 U6089 ( .A(n5798), .B(net59283), .ZN(n5796) );
  NAND2_X2 U6090 ( .A1(u4_div_exp3[10]), .A2(net58719), .ZN(n5795) );
  OAI221_X2 U6091 ( .B1(net58752), .B2(n5797), .C1(n5796), .C2(net58714), .A(
        n5795), .ZN(net58707) );
  INV_X4 U6092 ( .A(u4_div_exp1_9_), .ZN(n5802) );
  INV_X4 U6093 ( .A(net59270), .ZN(net59275) );
  NAND2_X2 U6094 ( .A1(u4_div_exp3[9]), .A2(net58719), .ZN(n5800) );
  OAI221_X2 U6095 ( .B1(net58752), .B2(n5802), .C1(n5801), .C2(net58714), .A(
        n5800), .ZN(net58759) );
  NAND2_X2 U6096 ( .A1(n5811), .A2(n5803), .ZN(n5813) );
  INV_X4 U6097 ( .A(n5813), .ZN(n5804) );
  NAND2_X2 U6098 ( .A1(n5804), .A2(n7172), .ZN(n5810) );
  NAND2_X2 U6099 ( .A1(n5810), .A2(u4_fi_ldz_4_), .ZN(n5805) );
  INV_X4 U6100 ( .A(n5805), .ZN(n5807) );
  INV_X4 U6101 ( .A(n5806), .ZN(n7159) );
  XNOR2_X2 U6102 ( .A(net57268), .B(n5807), .ZN(u4_fi_ldz_mi22[5]) );
  INV_X4 U6103 ( .A(n5810), .ZN(n5808) );
  XNOR2_X2 U6104 ( .A(n5808), .B(u4_fi_ldz_4_), .ZN(u4_fi_ldz_mi22[4]) );
  NAND2_X2 U6105 ( .A1(u4_fi_ldz_3_), .A2(n5813), .ZN(n5809) );
  NAND2_X2 U6106 ( .A1(n5810), .A2(n5809), .ZN(u4_fi_ldz_mi22[3]) );
  INV_X4 U6107 ( .A(n5811), .ZN(n5812) );
  NAND2_X2 U6108 ( .A1(n5812), .A2(u4_fi_ldz_2_), .ZN(n7173) );
  NAND2_X2 U6109 ( .A1(n7173), .A2(n5813), .ZN(u4_fi_ldz_mi22[2]) );
  INV_X4 U6110 ( .A(net58957), .ZN(net58951) );
  NAND2_X2 U6111 ( .A1(u4_exp_out_pl1_8_), .A2(net59078), .ZN(n5823) );
  NAND2_X2 U6112 ( .A1(net59231), .A2(net58643), .ZN(net59083) );
  NAND2_X2 U6113 ( .A1(net96080), .A2(net87237), .ZN(net59171) );
  NAND2_X2 U6114 ( .A1(u4_exp_out_2_), .A2(u4_exp_out_3_), .ZN(n5814) );
  NAND2_X2 U6115 ( .A1(u4_exp_out_6_), .A2(u4_exp_out_7_), .ZN(net59195) );
  NAND2_X2 U6116 ( .A1(n5815), .A2(net59228), .ZN(net59010) );
  OAI21_X4 U6117 ( .B1(net59224), .B2(net59219), .A(rmode_r3[1]), .ZN(net59193) );
  NAND2_X2 U6118 ( .A1(net66875), .A2(net66839), .ZN(n5816) );
  NOR2_X4 U6119 ( .A1(n7179), .A2(n5816), .ZN(net58650) );
  NAND2_X2 U6120 ( .A1(net58624), .A2(net59208), .ZN(net59217) );
  OAI21_X4 U6121 ( .B1(net59219), .B2(net58957), .A(net58932), .ZN(net59218)
         );
  INV_X4 U6122 ( .A(net59208), .ZN(net59214) );
  NAND3_X4 U6123 ( .A1(net59214), .A2(net58624), .A3(net63287), .ZN(net59079)
         );
  INV_X4 U6124 ( .A(net59088), .ZN(net59093) );
  NAND2_X2 U6125 ( .A1(u4_fi_ldz_5_), .A2(u4_fi_ldz_4_), .ZN(net59210) );
  INV_X4 U6126 ( .A(net58676), .ZN(net59207) );
  NAND2_X2 U6127 ( .A1(net58624), .A2(net63293), .ZN(net58997) );
  INV_X4 U6128 ( .A(u4_exp_fix_divb[8]), .ZN(n5820) );
  INV_X4 U6129 ( .A(u4_exp_fix_diva[8]), .ZN(n5819) );
  OAI22_X2 U6130 ( .A1(net59087), .A2(n5820), .B1(net59081), .B2(n5819), .ZN(
        n5821) );
  AOI21_X4 U6131 ( .B1(net59093), .B2(n4846), .A(n5821), .ZN(n5822) );
  NAND4_X2 U6132 ( .A1(n5823), .A2(net59200), .A3(net59201), .A4(n5822), .ZN(
        net59072) );
  INV_X4 U6133 ( .A(net59072), .ZN(net58988) );
  NAND2_X2 U6134 ( .A1(opb_00), .A2(net58645), .ZN(net58941) );
  NAND2_X2 U6135 ( .A1(opb_inf), .A2(net63293), .ZN(net58803) );
  NAND2_X2 U6136 ( .A1(net59093), .A2(net66863), .ZN(n5827) );
  AOI22_X2 U6137 ( .A1(u4_exp_fix_diva[7]), .A2(net59154), .B1(
        u4_exp_fix_divb[7]), .B2(net59122), .ZN(n5826) );
  INV_X4 U6138 ( .A(net59169), .ZN(net59146) );
  AOI22_X2 U6139 ( .A1(net59189), .A2(net59099), .B1(net59184), .B2(
        u4_exp_out_7_), .ZN(n5825) );
  AOI22_X2 U6140 ( .A1(u4_exp_next_mi_7_), .A2(net59117), .B1(
        u4_exp_out_pl1_7_), .B2(net59078), .ZN(n5824) );
  NAND4_X2 U6141 ( .A1(n5827), .A2(n5826), .A3(n5825), .A4(n5824), .ZN(
        net58980) );
  MUX2_X2 U6142 ( .A(net59183), .B(net59184), .S(u4_exp_out_6_), .Z(n5830) );
  INV_X4 U6143 ( .A(u4_exp_fix_divb[6]), .ZN(n5828) );
  OAI22_X2 U6144 ( .A1(net59087), .A2(n5828), .B1(n4384), .B2(net59088), .ZN(
        n5829) );
  NOR2_X4 U6145 ( .A1(n5830), .A2(n5829), .ZN(n5833) );
  NAND2_X2 U6146 ( .A1(u4_exp_fix_diva[6]), .A2(net59121), .ZN(n5832) );
  AOI22_X2 U6147 ( .A1(u4_exp_next_mi_6_), .A2(net59153), .B1(
        u4_exp_out_pl1_6_), .B2(net59078), .ZN(n5831) );
  NAND3_X4 U6148 ( .A1(n5833), .A2(n5832), .A3(n5831), .ZN(net58982) );
  NAND2_X2 U6149 ( .A1(net59093), .A2(exp_r[5]), .ZN(n5838) );
  AOI22_X2 U6150 ( .A1(u4_exp_fix_diva[5]), .A2(net59154), .B1(
        u4_exp_fix_divb[5]), .B2(net59122), .ZN(n5837) );
  NAND2_X2 U6151 ( .A1(u4_exp_out_3_), .A2(net59099), .ZN(n5834) );
  NAND2_X2 U6152 ( .A1(net59120), .A2(n5834), .ZN(net59159) );
  AOI22_X2 U6153 ( .A1(u4_exp_next_mi_5_), .A2(net59117), .B1(
        u4_exp_out_pl1_5_), .B2(net59078), .ZN(n5835) );
  NAND4_X2 U6154 ( .A1(n5838), .A2(n5837), .A3(n5836), .A4(n5835), .ZN(
        net58981) );
  INV_X4 U6155 ( .A(u4_exp_fix_divb[4]), .ZN(n5839) );
  OAI22_X2 U6156 ( .A1(net59087), .A2(n5839), .B1(n4328), .B2(net59088), .ZN(
        n5840) );
  NOR2_X4 U6157 ( .A1(net59155), .A2(n5840), .ZN(n5843) );
  NAND2_X2 U6158 ( .A1(u4_exp_fix_diva[4]), .A2(net59154), .ZN(n5842) );
  INV_X4 U6159 ( .A(net59079), .ZN(net59153) );
  AOI22_X2 U6160 ( .A1(u4_exp_next_mi_4_), .A2(net59153), .B1(
        u4_exp_out_pl1_4_), .B2(net59078), .ZN(n5841) );
  NAND2_X2 U6161 ( .A1(u4_exp_next_mi_2_), .A2(net59117), .ZN(n5851) );
  NAND2_X2 U6162 ( .A1(u4_exp_out_pl1_2_), .A2(net59078), .ZN(n5850) );
  NAND2_X2 U6163 ( .A1(net59099), .A2(u4_exp_out_0_), .ZN(n5844) );
  NAND2_X2 U6164 ( .A1(net59146), .A2(n5844), .ZN(net59110) );
  INV_X4 U6165 ( .A(net59110), .ZN(net59144) );
  INV_X4 U6166 ( .A(u4_exp_fix_divb[2]), .ZN(n5846) );
  INV_X4 U6167 ( .A(u4_exp_fix_diva[2]), .ZN(n5845) );
  OAI22_X2 U6168 ( .A1(net59087), .A2(n5846), .B1(net59081), .B2(n5845), .ZN(
        n5847) );
  NAND4_X2 U6169 ( .A1(n5851), .A2(n5850), .A3(n5849), .A4(n5848), .ZN(
        net58985) );
  INV_X4 U6170 ( .A(u4_exp_fix_divb[1]), .ZN(n5852) );
  OAI22_X2 U6171 ( .A1(net59087), .A2(n5852), .B1(n6010), .B2(net59088), .ZN(
        n5853) );
  NAND2_X2 U6172 ( .A1(u4_exp_fix_diva[1]), .A2(net59154), .ZN(n5855) );
  AOI22_X2 U6173 ( .A1(u4_exp_next_mi_1_), .A2(net59153), .B1(
        u4_exp_out_pl1_1_), .B2(net59078), .ZN(n5854) );
  NAND3_X4 U6174 ( .A1(n5856), .A2(n5855), .A3(n5854), .ZN(net58975) );
  NAND2_X2 U6175 ( .A1(u4_exp_out_pl1_9_), .A2(net59078), .ZN(n5863) );
  NAND2_X2 U6176 ( .A1(net59099), .A2(net59100), .ZN(n5862) );
  INV_X4 U6177 ( .A(u4_exp_fix_divb[9]), .ZN(n5859) );
  INV_X4 U6178 ( .A(u4_exp_fix_diva[9]), .ZN(n5858) );
  OAI22_X2 U6179 ( .A1(net59087), .A2(n5859), .B1(net59081), .B2(n5858), .ZN(
        n5860) );
  NAND4_X2 U6180 ( .A1(n5863), .A2(n5862), .A3(net59091), .A4(n5861), .ZN(
        net58987) );
  INV_X4 U6181 ( .A(u4_div_exp1_7_), .ZN(n5864) );
  NOR2_X4 U6182 ( .A1(n5864), .A2(net59064), .ZN(n5869) );
  NAND2_X2 U6183 ( .A1(u4_div_exp1_4_), .A2(u4_div_exp1_3_), .ZN(n5867) );
  AND2_X2 U6184 ( .A1(u4_div_exp1_1_), .A2(u4_div_exp1_0_), .ZN(n5865) );
  NAND2_X2 U6185 ( .A1(n5865), .A2(u4_div_exp1_2_), .ZN(n5866) );
  NOR2_X4 U6186 ( .A1(n5867), .A2(n5866), .ZN(n5868) );
  NAND4_X2 U6187 ( .A1(u4_div_exp1_8_), .A2(u4_div_exp1_9_), .A3(n5869), .A4(
        n5868), .ZN(n5870) );
  NAND2_X2 U6188 ( .A1(exp_ovf_r_0_), .A2(net66835), .ZN(net58631) );
  INV_X4 U6189 ( .A(n5871), .ZN(n5873) );
  OAI22_X2 U6190 ( .A1(opas_r2), .A2(n5873), .B1(net58808), .B2(n5872), .ZN(
        net58787) );
  INV_X4 U6191 ( .A(net59032), .ZN(net59030) );
  INV_X4 U6192 ( .A(net59010), .ZN(net59028) );
  NAND4_X2 U6193 ( .A1(net59027), .A2(net59028), .A3(u4_exp_out_0_), .A4(
        u4_exp_out_9_), .ZN(net59013) );
  NAND2_X2 U6194 ( .A1(net58650), .A2(net63217), .ZN(n5874) );
  INV_X4 U6195 ( .A(u4_fi_ldz_2a_4_), .ZN(net59024) );
  NAND2_X2 U6196 ( .A1(n5874), .A2(net59019), .ZN(net59014) );
  INV_X4 U6197 ( .A(net58987), .ZN(net58986) );
  NAND2_X2 U6198 ( .A1(net63545), .A2(u4_fract_out_0_), .ZN(n5876) );
  NAND2_X2 U6199 ( .A1(net58932), .A2(net58951), .ZN(net58947) );
  NAND2_X2 U6200 ( .A1(u4_fract_out_pl1_0_), .A2(net63559), .ZN(n5875) );
  NAND3_X4 U6201 ( .A1(net63577), .A2(n5876), .A3(n5875), .ZN(n6052) );
  NAND2_X2 U6202 ( .A1(opb_00), .A2(net63293), .ZN(n6106) );
  INV_X4 U6203 ( .A(n6106), .ZN(n5880) );
  INV_X4 U6204 ( .A(net58941), .ZN(net58938) );
  INV_X4 U6205 ( .A(net58517), .ZN(net58939) );
  NAND2_X2 U6206 ( .A1(inf_d), .A2(net58935), .ZN(n5878) );
  MUX2_X2 U6207 ( .A(n5878), .B(n4345), .S(net63293), .Z(n5883) );
  NAND2_X2 U6208 ( .A1(n4483), .A2(n4353), .ZN(n6145) );
  NAND2_X2 U6209 ( .A1(net58932), .A2(n6145), .ZN(n6042) );
  INV_X4 U6210 ( .A(n6042), .ZN(n5879) );
  NAND2_X2 U6211 ( .A1(n5879), .A2(net58645), .ZN(n5882) );
  NAND3_X2 U6212 ( .A1(n5883), .A2(n5882), .A3(n5881), .ZN(net58925) );
  MUX2_X2 U6213 ( .A(n6052), .B(net57282), .S(net63537), .Z(N793) );
  NAND2_X2 U6214 ( .A1(net58422), .A2(net58421), .ZN(n5922) );
  INV_X4 U6215 ( .A(net58419), .ZN(net58886) );
  AOI221_X2 U6216 ( .B1(net63541), .B2(u4_fract_out_47_), .C1(
        u4_fract_out_pl1_47_), .C2(net63559), .A(net63585), .ZN(n6140) );
  AOI221_X2 U6217 ( .B1(net63541), .B2(u4_fract_out_46_), .C1(
        u4_fract_out_pl1_46_), .C2(net63559), .A(net63585), .ZN(n6139) );
  AOI221_X2 U6218 ( .B1(net63541), .B2(u4_fract_out_45_), .C1(
        u4_fract_out_pl1_45_), .C2(net63559), .A(net63585), .ZN(n6138) );
  NAND2_X2 U6219 ( .A1(net63541), .A2(u4_fract_out_49_), .ZN(n5885) );
  NAND2_X2 U6220 ( .A1(u4_fract_out_pl1_49_), .A2(net63559), .ZN(n5884) );
  INV_X4 U6221 ( .A(n5886), .ZN(n6142) );
  NAND2_X2 U6222 ( .A1(net63545), .A2(u4_fract_out_48_), .ZN(n5888) );
  NAND2_X2 U6223 ( .A1(u4_fract_out_pl1_48_), .A2(net63559), .ZN(n5887) );
  INV_X4 U6224 ( .A(n5889), .ZN(n6141) );
  NAND2_X2 U6225 ( .A1(n6142), .A2(n6141), .ZN(n5897) );
  NAND2_X2 U6226 ( .A1(net63543), .A2(u4_fract_out_51_), .ZN(n5891) );
  NAND2_X2 U6227 ( .A1(u4_fract_out_pl1_51_), .A2(net63561), .ZN(n5890) );
  NAND3_X4 U6228 ( .A1(net63577), .A2(n5891), .A3(n5890), .ZN(n5892) );
  INV_X4 U6229 ( .A(n5892), .ZN(n6144) );
  NAND2_X2 U6230 ( .A1(net63545), .A2(u4_fract_out_50_), .ZN(n5894) );
  NAND2_X2 U6231 ( .A1(u4_fract_out_pl1_50_), .A2(net63567), .ZN(n5893) );
  NAND3_X4 U6232 ( .A1(net63577), .A2(n5894), .A3(n5893), .ZN(n5895) );
  INV_X4 U6233 ( .A(n5895), .ZN(n6143) );
  NAND2_X2 U6234 ( .A1(n6144), .A2(n6143), .ZN(n5896) );
  AOI221_X2 U6235 ( .B1(net63543), .B2(u4_fract_out_41_), .C1(
        u4_fract_out_pl1_41_), .C2(net63561), .A(net63585), .ZN(n6134) );
  AOI221_X2 U6236 ( .B1(net63543), .B2(u4_fract_out_40_), .C1(
        u4_fract_out_pl1_40_), .C2(net63561), .A(net63585), .ZN(n6133) );
  AOI221_X2 U6237 ( .B1(net63543), .B2(u4_fract_out_39_), .C1(
        u4_fract_out_pl1_39_), .C2(net63561), .A(net63585), .ZN(n6132) );
  AOI221_X2 U6238 ( .B1(net63543), .B2(u4_fract_out_44_), .C1(
        u4_fract_out_pl1_44_), .C2(net63561), .A(net63585), .ZN(n6137) );
  AOI221_X2 U6239 ( .B1(net63543), .B2(u4_fract_out_43_), .C1(
        u4_fract_out_pl1_43_), .C2(net63561), .A(net63585), .ZN(n6136) );
  AOI221_X2 U6240 ( .B1(net63543), .B2(u4_fract_out_42_), .C1(
        u4_fract_out_pl1_42_), .C2(net63561), .A(net63585), .ZN(n6135) );
  NOR2_X4 U6241 ( .A1(n5900), .A2(n5899), .ZN(n5920) );
  AOI221_X2 U6242 ( .B1(net63543), .B2(u4_fract_out_34_), .C1(
        u4_fract_out_pl1_34_), .C2(net63561), .A(net63585), .ZN(n6127) );
  AOI221_X2 U6243 ( .B1(net63543), .B2(u4_fract_out_33_), .C1(
        u4_fract_out_pl1_33_), .C2(net63561), .A(net63585), .ZN(n6126) );
  NAND2_X2 U6244 ( .A1(net63545), .A2(u4_fract_out_36_), .ZN(n5902) );
  NAND2_X2 U6245 ( .A1(u4_fract_out_pl1_36_), .A2(net63567), .ZN(n5901) );
  NAND3_X4 U6246 ( .A1(net63577), .A2(n5902), .A3(n5901), .ZN(n5903) );
  INV_X4 U6247 ( .A(n5903), .ZN(n6129) );
  NAND2_X2 U6248 ( .A1(net63545), .A2(u4_fract_out_35_), .ZN(n5905) );
  NAND2_X2 U6249 ( .A1(u4_fract_out_pl1_35_), .A2(net63567), .ZN(n5904) );
  NAND3_X4 U6250 ( .A1(net63577), .A2(n5905), .A3(n5904), .ZN(n5906) );
  INV_X4 U6251 ( .A(n5906), .ZN(n6128) );
  NAND2_X2 U6252 ( .A1(n6129), .A2(n6128), .ZN(n5914) );
  NAND2_X2 U6253 ( .A1(net63545), .A2(u4_fract_out_38_), .ZN(n5908) );
  NAND2_X2 U6254 ( .A1(u4_fract_out_pl1_38_), .A2(net63573), .ZN(n5907) );
  NAND3_X4 U6255 ( .A1(net63577), .A2(n5908), .A3(n5907), .ZN(n5909) );
  INV_X4 U6256 ( .A(n5909), .ZN(n6131) );
  NAND2_X2 U6257 ( .A1(net63547), .A2(u4_fract_out_37_), .ZN(n5911) );
  NAND2_X2 U6258 ( .A1(u4_fract_out_pl1_37_), .A2(net63573), .ZN(n5910) );
  NAND3_X4 U6259 ( .A1(net63577), .A2(n5911), .A3(n5910), .ZN(n5912) );
  INV_X4 U6260 ( .A(n5912), .ZN(n6130) );
  NAND2_X2 U6261 ( .A1(n6131), .A2(n6130), .ZN(n5913) );
  AOI221_X2 U6262 ( .B1(net63545), .B2(u4_fract_out_28_), .C1(
        u4_fract_out_pl1_28_), .C2(net63567), .A(net63585), .ZN(n6121) );
  AOI221_X2 U6263 ( .B1(net63543), .B2(u4_fract_out_26_), .C1(
        u4_fract_out_pl1_26_), .C2(net63561), .A(net63585), .ZN(n6119) );
  AOI221_X2 U6264 ( .B1(net63545), .B2(u4_fract_out_31_), .C1(
        u4_fract_out_pl1_31_), .C2(net63559), .A(net63585), .ZN(n6124) );
  AOI221_X2 U6265 ( .B1(net63543), .B2(u4_fract_out_30_), .C1(
        u4_fract_out_pl1_30_), .C2(net63561), .A(net63585), .ZN(n6123) );
  AOI221_X2 U6266 ( .B1(net63545), .B2(u4_fract_out_29_), .C1(
        u4_fract_out_pl1_29_), .C2(net63559), .A(net63585), .ZN(n6122) );
  NOR2_X4 U6267 ( .A1(n5916), .A2(n5917), .ZN(n5918) );
  NAND4_X2 U6268 ( .A1(n5921), .A2(n5920), .A3(n5919), .A4(n5918), .ZN(n6053)
         );
  INV_X4 U6269 ( .A(net58423), .ZN(net58587) );
  INV_X4 U6270 ( .A(net58424), .ZN(net58585) );
  NOR3_X4 U6271 ( .A1(net58584), .A2(net58587), .A3(net58585), .ZN(net58826)
         );
  NAND2_X2 U6272 ( .A1(net63547), .A2(u4_fract_out_1_), .ZN(n5924) );
  NAND2_X2 U6273 ( .A1(u4_fract_out_pl1_1_), .A2(net63565), .ZN(n5923) );
  NAND3_X4 U6274 ( .A1(net63577), .A2(n5924), .A3(n5923), .ZN(n6110) );
  NOR2_X4 U6275 ( .A1(n6110), .A2(n6052), .ZN(n5932) );
  NAND2_X2 U6276 ( .A1(net63547), .A2(u4_fract_out_3_), .ZN(n5926) );
  NAND2_X2 U6277 ( .A1(u4_fract_out_pl1_3_), .A2(net63565), .ZN(n5925) );
  NAND3_X4 U6278 ( .A1(net63577), .A2(n5926), .A3(n5925), .ZN(n5927) );
  INV_X4 U6279 ( .A(n5927), .ZN(n6113) );
  NAND2_X2 U6280 ( .A1(net63547), .A2(u4_fract_out_2_), .ZN(n5929) );
  NAND2_X2 U6281 ( .A1(u4_fract_out_pl1_2_), .A2(net63565), .ZN(n5928) );
  NAND3_X4 U6282 ( .A1(net63577), .A2(n5929), .A3(n5928), .ZN(n5930) );
  INV_X4 U6283 ( .A(n5930), .ZN(n6112) );
  NAND2_X2 U6284 ( .A1(n6113), .A2(n6112), .ZN(n6054) );
  INV_X4 U6285 ( .A(n6054), .ZN(n5931) );
  NAND2_X2 U6286 ( .A1(n5932), .A2(n5931), .ZN(n5938) );
  AOI221_X2 U6287 ( .B1(net63543), .B2(u4_fract_out_4_), .C1(
        u4_fract_out_pl1_4_), .C2(net63561), .A(net63585), .ZN(n6114) );
  AOI221_X2 U6288 ( .B1(net63541), .B2(u4_fract_out_5_), .C1(
        u4_fract_out_pl1_5_), .C2(net63559), .A(net63587), .ZN(n6115) );
  NAND2_X2 U6289 ( .A1(n6114), .A2(n6115), .ZN(n6060) );
  NAND2_X2 U6290 ( .A1(net63547), .A2(u4_fract_out_6_), .ZN(n5934) );
  NAND2_X2 U6291 ( .A1(u4_fract_out_pl1_6_), .A2(net63565), .ZN(n5933) );
  NAND3_X4 U6292 ( .A1(net63579), .A2(n5934), .A3(n5933), .ZN(n6059) );
  INV_X4 U6293 ( .A(n6059), .ZN(n6116) );
  NAND2_X2 U6294 ( .A1(net63547), .A2(u4_fract_out_7_), .ZN(n5936) );
  NAND2_X2 U6295 ( .A1(u4_fract_out_pl1_7_), .A2(net63565), .ZN(n5935) );
  NAND3_X4 U6296 ( .A1(net63579), .A2(n5936), .A3(n5935), .ZN(n6097) );
  INV_X4 U6297 ( .A(n6097), .ZN(n6117) );
  NAND2_X2 U6298 ( .A1(n6116), .A2(n6117), .ZN(n5937) );
  NOR3_X4 U6299 ( .A1(n5938), .A2(n6060), .A3(n5937), .ZN(net58827) );
  NAND2_X2 U6300 ( .A1(net63547), .A2(u4_fract_out_18_), .ZN(n5940) );
  NAND2_X2 U6301 ( .A1(u4_fract_out_pl1_18_), .A2(net63565), .ZN(n5939) );
  NAND3_X4 U6302 ( .A1(net63579), .A2(n5940), .A3(n5939), .ZN(net58481) );
  NAND2_X2 U6303 ( .A1(net63547), .A2(u4_fract_out_19_), .ZN(n5942) );
  NAND2_X2 U6304 ( .A1(u4_fract_out_pl1_19_), .A2(net63565), .ZN(n5941) );
  NAND3_X4 U6305 ( .A1(net63579), .A2(n5942), .A3(n5941), .ZN(net58479) );
  NAND2_X2 U6306 ( .A1(net63547), .A2(u4_fract_out_16_), .ZN(n5944) );
  NAND2_X2 U6307 ( .A1(u4_fract_out_pl1_16_), .A2(net63565), .ZN(n5943) );
  NAND3_X4 U6308 ( .A1(net63579), .A2(n5944), .A3(n5943), .ZN(net58485) );
  NAND2_X2 U6309 ( .A1(net63547), .A2(u4_fract_out_17_), .ZN(n5946) );
  NAND2_X2 U6310 ( .A1(u4_fract_out_pl1_17_), .A2(net63565), .ZN(n5945) );
  NAND3_X4 U6311 ( .A1(net63579), .A2(n5946), .A3(n5945), .ZN(net58483) );
  NAND2_X2 U6312 ( .A1(net63547), .A2(u4_fract_out_13_), .ZN(n5948) );
  NAND2_X2 U6313 ( .A1(u4_fract_out_pl1_13_), .A2(net63565), .ZN(n5947) );
  NAND3_X4 U6314 ( .A1(net63579), .A2(n5948), .A3(n5947), .ZN(net58491) );
  NAND2_X2 U6315 ( .A1(net63547), .A2(u4_fract_out_14_), .ZN(n5950) );
  NAND2_X2 U6316 ( .A1(u4_fract_out_pl1_14_), .A2(net63565), .ZN(n5949) );
  NAND3_X4 U6317 ( .A1(net63579), .A2(n5950), .A3(n5949), .ZN(net58489) );
  NAND2_X2 U6318 ( .A1(net63547), .A2(u4_fract_out_15_), .ZN(n5952) );
  NAND2_X2 U6319 ( .A1(u4_fract_out_pl1_15_), .A2(net63565), .ZN(n5951) );
  NAND3_X4 U6320 ( .A1(net63579), .A2(n5952), .A3(n5951), .ZN(net58487) );
  AOI221_X2 U6321 ( .B1(net63541), .B2(u4_fract_out_24_), .C1(
        u4_fract_out_pl1_24_), .C2(net63559), .A(net63587), .ZN(net58472) );
  NAND2_X2 U6322 ( .A1(net63547), .A2(u4_fract_out_23_), .ZN(n5954) );
  NAND2_X2 U6323 ( .A1(u4_fract_out_pl1_23_), .A2(net63565), .ZN(n5953) );
  NAND3_X4 U6324 ( .A1(net63579), .A2(n5954), .A3(n5953), .ZN(net58592) );
  AOI221_X2 U6325 ( .B1(net63541), .B2(u4_fract_out_9_), .C1(
        u4_fract_out_pl1_9_), .C2(net63559), .A(net63587), .ZN(net58495) );
  NAND2_X2 U6326 ( .A1(net63547), .A2(u4_fract_out_8_), .ZN(n5956) );
  NAND2_X2 U6327 ( .A1(u4_fract_out_pl1_8_), .A2(net63565), .ZN(n5955) );
  INV_X4 U6328 ( .A(n6058), .ZN(n6118) );
  NAND2_X2 U6329 ( .A1(net58495), .A2(n6118), .ZN(net58533) );
  AOI221_X2 U6330 ( .B1(net63541), .B2(u4_fract_out_11_), .C1(
        u4_fract_out_pl1_11_), .C2(net63559), .A(net63587), .ZN(net58493) );
  AOI221_X2 U6331 ( .B1(net63541), .B2(u4_fract_out_10_), .C1(
        u4_fract_out_pl1_10_), .C2(net63559), .A(net63587), .ZN(net58494) );
  NAND2_X2 U6332 ( .A1(net58493), .A2(net58494), .ZN(net58524) );
  NAND2_X2 U6333 ( .A1(net63547), .A2(u4_fract_out_22_), .ZN(n5958) );
  NAND2_X2 U6334 ( .A1(u4_fract_out_pl1_22_), .A2(net63567), .ZN(n5957) );
  NAND3_X4 U6335 ( .A1(net63579), .A2(n5958), .A3(n5957), .ZN(net58475) );
  NAND2_X2 U6336 ( .A1(net63545), .A2(u4_fract_out_21_), .ZN(n5960) );
  NAND2_X2 U6337 ( .A1(u4_fract_out_pl1_21_), .A2(net63559), .ZN(n5959) );
  NAND3_X4 U6338 ( .A1(net63577), .A2(n5960), .A3(n5959), .ZN(net58526) );
  AOI221_X2 U6339 ( .B1(net63541), .B2(u4_fract_out_20_), .C1(
        u4_fract_out_pl1_20_), .C2(net63559), .A(net63587), .ZN(net58477) );
  NAND2_X2 U6340 ( .A1(opb_00), .A2(opa_00), .ZN(net58802) );
  NAND2_X2 U6341 ( .A1(opb_inf), .A2(opa_00), .ZN(n5962) );
  NAND2_X2 U6342 ( .A1(opb_00), .A2(opa_inf), .ZN(n5961) );
  NAND2_X2 U6343 ( .A1(n5962), .A2(n5961), .ZN(net58623) );
  INV_X4 U6344 ( .A(net58803), .ZN(net58801) );
  NAND2_X2 U6345 ( .A1(net58801), .A2(net58802), .ZN(n5963) );
  NAND2_X2 U6346 ( .A1(n5963), .A2(net58799), .ZN(net58793) );
  INV_X4 U6347 ( .A(net58646), .ZN(net58783) );
  NAND2_X2 U6348 ( .A1(net58781), .A2(n5967), .ZN(net58773) );
  NAND2_X2 U6349 ( .A1(net58780), .A2(net58646), .ZN(net58774) );
  NAND2_X2 U6350 ( .A1(net66875), .A2(net58682), .ZN(n6008) );
  NAND2_X2 U6351 ( .A1(n5968), .A2(net58767), .ZN(n5969) );
  INV_X4 U6352 ( .A(n5969), .ZN(n5970) );
  AOI22_X2 U6353 ( .A1(u4_div_exp1_2_), .A2(net58718), .B1(u4_div_exp3[2]), 
        .B2(net58719), .ZN(n5971) );
  NAND2_X2 U6354 ( .A1(n5973), .A2(n7177), .ZN(n5982) );
  INV_X4 U6355 ( .A(net58759), .ZN(net58750) );
  INV_X4 U6356 ( .A(u4_div_exp1_8_), .ZN(n5979) );
  INV_X4 U6357 ( .A(n7201), .ZN(n5976) );
  NAND2_X2 U6358 ( .A1(u4_div_exp3[8]), .A2(net58719), .ZN(n5977) );
  OAI221_X2 U6359 ( .B1(net58752), .B2(n5979), .C1(n5978), .C2(net58714), .A(
        n5977), .ZN(n5980) );
  INV_X4 U6360 ( .A(n5980), .ZN(n7199) );
  NAND3_X2 U6361 ( .A1(net58750), .A2(u4_exp_in_mi1_11_), .A3(n7199), .ZN(
        n5981) );
  NOR2_X4 U6362 ( .A1(n5982), .A2(n5981), .ZN(n6006) );
  INV_X4 U6363 ( .A(net58733), .ZN(net58743) );
  INV_X4 U6364 ( .A(n7204), .ZN(n5984) );
  NAND2_X2 U6365 ( .A1(n5984), .A2(n5983), .ZN(n5985) );
  INV_X4 U6366 ( .A(n5985), .ZN(n5986) );
  AOI22_X2 U6367 ( .A1(u4_div_exp1_4_), .A2(net58718), .B1(u4_div_exp3[4]), 
        .B2(net58719), .ZN(n5987) );
  NOR2_X4 U6368 ( .A1(n5991), .A2(n5990), .ZN(n5993) );
  AOI22_X2 U6369 ( .A1(u4_div_exp1_3_), .A2(net58718), .B1(u4_div_exp3[3]), 
        .B2(net58719), .ZN(n5992) );
  AOI22_X2 U6370 ( .A1(u4_div_exp1_6_), .A2(net58718), .B1(u4_div_exp3[6]), 
        .B2(net58719), .ZN(n5995) );
  INV_X4 U6371 ( .A(n5997), .ZN(n8243) );
  NOR2_X4 U6372 ( .A1(n6000), .A2(n5999), .ZN(n6002) );
  AOI22_X2 U6373 ( .A1(u4_div_exp1_7_), .A2(net58718), .B1(u4_div_exp3[7]), 
        .B2(net58719), .ZN(n6001) );
  INV_X4 U6374 ( .A(n6003), .ZN(n8242) );
  INV_X4 U6375 ( .A(net58682), .ZN(net58673) );
  INV_X4 U6376 ( .A(net58707), .ZN(net58706) );
  MUX2_X2 U6377 ( .A(n6008), .B(n6007), .S(net58706), .Z(n6032) );
  NAND2_X2 U6378 ( .A1(net58550), .A2(net66835), .ZN(n6031) );
  NAND2_X2 U6379 ( .A1(net58682), .A2(n4308), .ZN(n6016) );
  INV_X4 U6380 ( .A(u4_ldz_all_3_), .ZN(n6012) );
  INV_X4 U6381 ( .A(u4_ldz_all_2_), .ZN(n6011) );
  NAND2_X2 U6382 ( .A1(n6012), .A2(n6011), .ZN(n6013) );
  INV_X4 U6383 ( .A(n6014), .ZN(n6015) );
  NAND2_X2 U6384 ( .A1(n7211), .A2(exp_r[5]), .ZN(n6019) );
  INV_X4 U6385 ( .A(net58688), .ZN(net58687) );
  NAND2_X2 U6386 ( .A1(u4_N6280), .A2(net58682), .ZN(n6023) );
  OAI211_X2 U6387 ( .C1(n6032), .C2(n6031), .A(n6030), .B(n6029), .ZN(net58666) );
  NAND2_X2 U6388 ( .A1(net58658), .A2(n6035), .ZN(n6036) );
  NAND4_X2 U6389 ( .A1(net58653), .A2(n6036), .A3(net58631), .A4(net58655), 
        .ZN(n6039) );
  NAND3_X2 U6390 ( .A1(net58645), .A2(net58646), .A3(n6037), .ZN(n6038) );
  NAND3_X2 U6391 ( .A1(n6039), .A2(n6038), .A3(net58641), .ZN(n6095) );
  MUX2_X2 U6392 ( .A(net58628), .B(net58629), .S(net63293), .Z(n6148) );
  INV_X4 U6393 ( .A(n6148), .ZN(n6040) );
  NAND2_X2 U6394 ( .A1(n6041), .A2(n6040), .ZN(n6045) );
  INV_X4 U6395 ( .A(n6045), .ZN(n6051) );
  NAND2_X2 U6396 ( .A1(net58624), .A2(n6145), .ZN(net58615) );
  NAND3_X2 U6397 ( .A1(n6042), .A2(n4345), .A3(n4429), .ZN(n6043) );
  NAND2_X2 U6398 ( .A1(n6044), .A2(n6043), .ZN(n6103) );
  INV_X4 U6399 ( .A(n6103), .ZN(n6046) );
  NOR2_X4 U6400 ( .A1(n6046), .A2(n6045), .ZN(net58617) );
  NAND2_X2 U6401 ( .A1(net63083), .A2(net58609), .ZN(n6049) );
  OAI221_X2 U6402 ( .B1(n6051), .B2(n4357), .C1(n6050), .C2(net58437), .A(
        n6049), .ZN(N889) );
  INV_X4 U6403 ( .A(n6052), .ZN(n6057) );
  NOR2_X4 U6404 ( .A1(n6054), .A2(n6110), .ZN(n6055) );
  NAND3_X4 U6405 ( .A1(n6057), .A2(n6056), .A3(n6055), .ZN(n6099) );
  INV_X4 U6406 ( .A(n6060), .ZN(n6061) );
  NAND2_X2 U6407 ( .A1(n6062), .A2(n6061), .ZN(n6063) );
  NOR4_X2 U6408 ( .A1(n6099), .A2(n6063), .A3(net58589), .A4(net58590), .ZN(
        n6067) );
  INV_X4 U6409 ( .A(net58422), .ZN(net58586) );
  INV_X4 U6410 ( .A(net58584), .ZN(net58583) );
  NAND2_X2 U6411 ( .A1(n6064), .A2(net58583), .ZN(n6065) );
  INV_X4 U6412 ( .A(net58581), .ZN(net58429) );
  NOR3_X4 U6413 ( .A1(n6065), .A2(net58579), .A3(net58580), .ZN(n6066) );
  OAI21_X4 U6414 ( .B1(n6067), .B2(n6066), .A(underflow_fmul_r[2]), .ZN(n6094)
         );
  NOR4_X2 U6415 ( .A1(prod[91]), .A2(prod[90]), .A3(prod[92]), .A4(prod[93]), 
        .ZN(n6071) );
  NOR4_X2 U6416 ( .A1(prod[84]), .A2(prod[83]), .A3(prod[86]), .A4(prod[85]), 
        .ZN(n6069) );
  NAND4_X2 U6417 ( .A1(n6071), .A2(n6070), .A3(n6069), .A4(n6068), .ZN(n6077)
         );
  NAND4_X2 U6418 ( .A1(n3378), .A2(n3381), .A3(n6073), .A4(n6072), .ZN(n6076)
         );
  NAND3_X2 U6419 ( .A1(n3363), .A2(n3364), .A3(n3362), .ZN(n6075) );
  NAND4_X2 U6420 ( .A1(n3356), .A2(n3357), .A3(n3365), .A4(n3355), .ZN(n6074)
         );
  NOR4_X2 U6421 ( .A1(n6077), .A2(n6076), .A3(n6075), .A4(n6074), .ZN(n6092)
         );
  NOR4_X2 U6422 ( .A1(prod[57]), .A2(prod[58]), .A3(prod[60]), .A4(prod[59]), 
        .ZN(n6081) );
  NAND4_X2 U6423 ( .A1(n6081), .A2(n6080), .A3(n6079), .A4(n6078), .ZN(n6090)
         );
  NAND4_X2 U6424 ( .A1(n6084), .A2(n6083), .A3(n6082), .A4(n4479), .ZN(n6089)
         );
  NAND4_X2 U6425 ( .A1(n6087), .A2(n6086), .A3(n6085), .A4(n4480), .ZN(n6088)
         );
  AOI21_X2 U6426 ( .B1(n6092), .B2(n6091), .A(net58550), .ZN(net58547) );
  AOI21_X2 U6427 ( .B1(underflow_fmul_r[1]), .B2(n6095), .A(
        underflow_fmul_r[0]), .ZN(n6093) );
  NAND3_X2 U6428 ( .A1(n6094), .A2(net58544), .A3(n6093), .ZN(net58540) );
  NAND2_X2 U6429 ( .A1(net58537), .A2(n6095), .ZN(n6096) );
  NAND2_X2 U6430 ( .A1(net58535), .A2(n6096), .ZN(N902) );
  INV_X4 U6431 ( .A(n6099), .ZN(n6101) );
  INV_X4 U6432 ( .A(net58526), .ZN(net58476) );
  NAND3_X4 U6433 ( .A1(n6102), .A2(n6101), .A3(n6100), .ZN(n6104) );
  NAND2_X2 U6434 ( .A1(n6104), .A2(n6103), .ZN(n6108) );
  NAND3_X2 U6435 ( .A1(inf_d), .A2(net63513), .A3(net58517), .ZN(n6105) );
  AOI211_X4 U6436 ( .C1(n6108), .C2(net63089), .A(n6107), .B(n4471), .ZN(n6109) );
  NOR2_X4 U6437 ( .A1(n6109), .A2(net58506), .ZN(N906) );
  INV_X4 U6438 ( .A(n6110), .ZN(n6111) );
  NOR2_X4 U6439 ( .A1(net63529), .A2(n6111), .ZN(N794) );
  NOR2_X4 U6440 ( .A1(net63527), .A2(n6112), .ZN(N795) );
  NOR2_X4 U6441 ( .A1(net63529), .A2(n6113), .ZN(N796) );
  NOR2_X4 U6442 ( .A1(net63529), .A2(n6118), .ZN(N801) );
  INV_X4 U6443 ( .A(net58491), .ZN(net58490) );
  NOR2_X4 U6444 ( .A1(net63529), .A2(net58490), .ZN(N806) );
  INV_X4 U6445 ( .A(net58489), .ZN(net58488) );
  NOR2_X4 U6446 ( .A1(net63529), .A2(net58488), .ZN(N807) );
  INV_X4 U6447 ( .A(net58487), .ZN(net58486) );
  NOR2_X4 U6448 ( .A1(net63529), .A2(net58486), .ZN(N808) );
  INV_X4 U6449 ( .A(net58485), .ZN(net58484) );
  NOR2_X4 U6450 ( .A1(net63527), .A2(net58484), .ZN(N809) );
  INV_X4 U6451 ( .A(net58483), .ZN(net58482) );
  NOR2_X4 U6452 ( .A1(net63527), .A2(net58482), .ZN(N810) );
  INV_X4 U6453 ( .A(net58481), .ZN(net58480) );
  NOR2_X4 U6454 ( .A1(net63527), .A2(net58480), .ZN(N811) );
  INV_X4 U6455 ( .A(net58479), .ZN(net58478) );
  NOR2_X4 U6456 ( .A1(net63527), .A2(net58478), .ZN(N812) );
  NOR2_X4 U6457 ( .A1(net63527), .A2(net58476), .ZN(N814) );
  INV_X4 U6458 ( .A(net58475), .ZN(net58474) );
  NOR2_X4 U6459 ( .A1(net63527), .A2(net58474), .ZN(N815) );
  NOR2_X4 U6460 ( .A1(net63523), .A2(n6128), .ZN(N828) );
  NOR2_X4 U6461 ( .A1(net63523), .A2(n6129), .ZN(N829) );
  NOR2_X4 U6462 ( .A1(net63523), .A2(n6130), .ZN(N830) );
  NOR2_X4 U6463 ( .A1(net63523), .A2(n6131), .ZN(N831) );
  NOR2_X4 U6464 ( .A1(net63523), .A2(n6141), .ZN(N841) );
  NOR2_X4 U6465 ( .A1(net63523), .A2(n6142), .ZN(N842) );
  NOR2_X4 U6466 ( .A1(net63523), .A2(n6143), .ZN(N843) );
  NOR2_X4 U6467 ( .A1(net63523), .A2(n6144), .ZN(N844) );
  INV_X4 U6468 ( .A(n6145), .ZN(n6146) );
  INV_X4 U6469 ( .A(net58437), .ZN(net58434) );
  NAND2_X2 U6470 ( .A1(net58420), .A2(net58429), .ZN(N854) );
  NAND2_X2 U6471 ( .A1(net58420), .A2(net58425), .ZN(N851) );
  NAND2_X2 U6472 ( .A1(net58420), .A2(net58424), .ZN(N852) );
  NAND2_X2 U6473 ( .A1(net58420), .A2(net58423), .ZN(N850) );
  NAND2_X2 U6474 ( .A1(net58420), .A2(net58422), .ZN(N847) );
  NAND2_X2 U6475 ( .A1(net58420), .A2(net58421), .ZN(N849) );
  NAND2_X2 U6476 ( .A1(net58419), .A2(net58420), .ZN(N848) );
  INV_X4 U6477 ( .A(N307), .ZN(n6149) );
  MUX2_X2 U6478 ( .A(n4297), .B(n6149), .S(n4900), .Z(n6150) );
  INV_X4 U6479 ( .A(n6150), .ZN(u6_N106) );
  INV_X4 U6480 ( .A(N306), .ZN(n6151) );
  MUX2_X2 U6481 ( .A(n4291), .B(n6151), .S(n4902), .Z(n6152) );
  INV_X4 U6482 ( .A(n6152), .ZN(u6_N105) );
  INV_X4 U6483 ( .A(N305), .ZN(n6153) );
  MUX2_X2 U6484 ( .A(n4301), .B(n6153), .S(n4899), .Z(n6154) );
  INV_X4 U6485 ( .A(n6154), .ZN(u6_N104) );
  INV_X4 U6486 ( .A(N304), .ZN(n6155) );
  MUX2_X2 U6487 ( .A(n4303), .B(n6155), .S(n4899), .Z(n6156) );
  INV_X4 U6488 ( .A(n6156), .ZN(u6_N103) );
  INV_X4 U6489 ( .A(N303), .ZN(n6157) );
  MUX2_X2 U6490 ( .A(n4302), .B(n6157), .S(n4900), .Z(n6158) );
  INV_X4 U6491 ( .A(n6158), .ZN(u6_N102) );
  INV_X4 U6492 ( .A(N302), .ZN(n6159) );
  MUX2_X2 U6493 ( .A(n4300), .B(n6159), .S(n4900), .Z(n6160) );
  INV_X4 U6494 ( .A(n6160), .ZN(u6_N101) );
  INV_X4 U6495 ( .A(N301), .ZN(n6161) );
  MUX2_X2 U6496 ( .A(n4290), .B(n6161), .S(n4902), .Z(n6162) );
  INV_X4 U6497 ( .A(n6162), .ZN(u6_N100) );
  INV_X4 U6498 ( .A(N300), .ZN(n6163) );
  MUX2_X2 U6499 ( .A(n6451), .B(n6163), .S(n4902), .Z(n6164) );
  INV_X4 U6500 ( .A(n6164), .ZN(u6_N99) );
  INV_X4 U6501 ( .A(N299), .ZN(n6165) );
  MUX2_X2 U6502 ( .A(n4296), .B(n6165), .S(n4899), .Z(n6166) );
  INV_X4 U6503 ( .A(n6166), .ZN(u6_N98) );
  INV_X4 U6504 ( .A(N298), .ZN(n6167) );
  MUX2_X2 U6505 ( .A(n4436), .B(n6167), .S(n4902), .Z(n6168) );
  INV_X4 U6506 ( .A(n6168), .ZN(u6_N97) );
  INV_X4 U6507 ( .A(N297), .ZN(n6169) );
  MUX2_X2 U6508 ( .A(n4313), .B(n6169), .S(n4902), .Z(n6170) );
  INV_X4 U6509 ( .A(n6170), .ZN(u6_N96) );
  INV_X4 U6510 ( .A(N296), .ZN(n6171) );
  MUX2_X2 U6511 ( .A(n4344), .B(n6171), .S(n4902), .Z(n6172) );
  INV_X4 U6512 ( .A(n6172), .ZN(u6_N95) );
  INV_X4 U6513 ( .A(N295), .ZN(n6173) );
  MUX2_X2 U6514 ( .A(n4439), .B(n6173), .S(n4902), .Z(n6174) );
  INV_X4 U6515 ( .A(n6174), .ZN(u6_N94) );
  INV_X4 U6516 ( .A(N294), .ZN(n6175) );
  MUX2_X2 U6517 ( .A(n4335), .B(n6175), .S(n4902), .Z(n6176) );
  INV_X4 U6518 ( .A(n6176), .ZN(u6_N93) );
  INV_X4 U6519 ( .A(N293), .ZN(n6177) );
  MUX2_X2 U6520 ( .A(n4310), .B(n6177), .S(n4902), .Z(n6178) );
  INV_X4 U6521 ( .A(n6178), .ZN(u6_N92) );
  INV_X4 U6522 ( .A(N292), .ZN(n6179) );
  MUX2_X2 U6523 ( .A(n4340), .B(n6179), .S(n4902), .Z(n6180) );
  INV_X4 U6524 ( .A(n6180), .ZN(u6_N91) );
  INV_X4 U6525 ( .A(N291), .ZN(n6181) );
  MUX2_X2 U6526 ( .A(n4311), .B(n6181), .S(n4902), .Z(n6182) );
  INV_X4 U6527 ( .A(n6182), .ZN(u6_N90) );
  INV_X4 U6528 ( .A(N290), .ZN(n6183) );
  MUX2_X2 U6529 ( .A(n4314), .B(n6183), .S(n4902), .Z(n6184) );
  INV_X4 U6530 ( .A(n6184), .ZN(u6_N89) );
  INV_X4 U6531 ( .A(N289), .ZN(n6185) );
  MUX2_X2 U6532 ( .A(n4338), .B(n6185), .S(n4902), .Z(n6186) );
  INV_X4 U6533 ( .A(n6186), .ZN(u6_N88) );
  INV_X4 U6534 ( .A(N288), .ZN(n6187) );
  MUX2_X2 U6535 ( .A(n4342), .B(n6187), .S(n4901), .Z(n6188) );
  INV_X4 U6536 ( .A(n6188), .ZN(u6_N87) );
  INV_X4 U6537 ( .A(N287), .ZN(n6189) );
  MUX2_X2 U6538 ( .A(n4423), .B(n6189), .S(n4901), .Z(n6190) );
  INV_X4 U6539 ( .A(n6190), .ZN(u6_N86) );
  INV_X4 U6540 ( .A(N286), .ZN(n6191) );
  MUX2_X2 U6541 ( .A(n4419), .B(n6191), .S(n4901), .Z(n6192) );
  INV_X4 U6542 ( .A(n6192), .ZN(u6_N85) );
  INV_X4 U6543 ( .A(N285), .ZN(n6193) );
  MUX2_X2 U6544 ( .A(n4431), .B(n6193), .S(n4901), .Z(n6194) );
  INV_X4 U6545 ( .A(n6194), .ZN(u6_N84) );
  INV_X4 U6546 ( .A(N284), .ZN(n6195) );
  MUX2_X2 U6547 ( .A(n4418), .B(n6195), .S(n4901), .Z(n6196) );
  INV_X4 U6548 ( .A(n6196), .ZN(u6_N83) );
  INV_X4 U6549 ( .A(N283), .ZN(n6197) );
  MUX2_X2 U6550 ( .A(n4426), .B(n6197), .S(n4901), .Z(n6198) );
  INV_X4 U6551 ( .A(n6198), .ZN(u6_N82) );
  INV_X4 U6552 ( .A(N282), .ZN(n6199) );
  MUX2_X2 U6553 ( .A(n4422), .B(n6199), .S(n4901), .Z(n6200) );
  INV_X4 U6554 ( .A(n6200), .ZN(u6_N81) );
  INV_X4 U6555 ( .A(N281), .ZN(n6201) );
  MUX2_X2 U6556 ( .A(n4421), .B(n6201), .S(n4901), .Z(n6202) );
  INV_X4 U6557 ( .A(n6202), .ZN(u6_N80) );
  INV_X4 U6558 ( .A(N280), .ZN(n6203) );
  MUX2_X2 U6559 ( .A(n4435), .B(n6203), .S(n4901), .Z(n6204) );
  INV_X4 U6560 ( .A(n6204), .ZN(u6_N79) );
  INV_X4 U6561 ( .A(N279), .ZN(n6205) );
  MUX2_X2 U6562 ( .A(n4417), .B(n6205), .S(n4901), .Z(n6206) );
  INV_X4 U6563 ( .A(n6206), .ZN(u6_N78) );
  INV_X4 U6564 ( .A(N278), .ZN(n6207) );
  MUX2_X2 U6565 ( .A(n4289), .B(n6207), .S(n4900), .Z(n6208) );
  INV_X4 U6566 ( .A(n6208), .ZN(u6_N77) );
  INV_X4 U6567 ( .A(N277), .ZN(n6209) );
  MUX2_X2 U6568 ( .A(n4437), .B(n6209), .S(n4900), .Z(n6210) );
  INV_X4 U6569 ( .A(n6210), .ZN(u6_N76) );
  INV_X4 U6570 ( .A(N276), .ZN(n6211) );
  MUX2_X2 U6571 ( .A(n4299), .B(n6211), .S(n4900), .Z(n6212) );
  INV_X4 U6572 ( .A(n6212), .ZN(u6_N75) );
  INV_X4 U6573 ( .A(N275), .ZN(n6213) );
  MUX2_X2 U6574 ( .A(n4438), .B(n6213), .S(n4900), .Z(n6214) );
  INV_X4 U6575 ( .A(n6214), .ZN(u6_N74) );
  INV_X4 U6576 ( .A(N274), .ZN(n6215) );
  MUX2_X2 U6577 ( .A(n4427), .B(n6215), .S(n4900), .Z(n6216) );
  INV_X4 U6578 ( .A(n6216), .ZN(u6_N73) );
  INV_X4 U6579 ( .A(N273), .ZN(n6217) );
  MUX2_X2 U6580 ( .A(n4341), .B(n6217), .S(n4900), .Z(n6218) );
  INV_X4 U6581 ( .A(n6218), .ZN(u6_N72) );
  INV_X4 U6582 ( .A(N272), .ZN(n6219) );
  MUX2_X2 U6583 ( .A(n4347), .B(n6219), .S(n4900), .Z(n6220) );
  INV_X4 U6584 ( .A(n6220), .ZN(u6_N71) );
  INV_X4 U6585 ( .A(N271), .ZN(n6221) );
  MUX2_X2 U6586 ( .A(n4339), .B(n6221), .S(n4900), .Z(n6222) );
  INV_X4 U6587 ( .A(n6222), .ZN(u6_N70) );
  INV_X4 U6588 ( .A(N270), .ZN(n6223) );
  MUX2_X2 U6589 ( .A(n4434), .B(n6223), .S(n4900), .Z(n6224) );
  INV_X4 U6590 ( .A(n6224), .ZN(u6_N69) );
  INV_X4 U6591 ( .A(N269), .ZN(n6225) );
  MUX2_X2 U6592 ( .A(n4336), .B(n6225), .S(n4900), .Z(n6226) );
  INV_X4 U6593 ( .A(n6226), .ZN(u6_N68) );
  INV_X4 U6594 ( .A(N268), .ZN(n6227) );
  MUX2_X2 U6595 ( .A(n4315), .B(n6227), .S(n4900), .Z(n6228) );
  INV_X4 U6596 ( .A(n6228), .ZN(u6_N67) );
  INV_X4 U6597 ( .A(N267), .ZN(n6229) );
  MUX2_X2 U6598 ( .A(n4312), .B(n6229), .S(n4901), .Z(n6230) );
  INV_X4 U6599 ( .A(n6230), .ZN(u6_N66) );
  INV_X4 U6600 ( .A(N266), .ZN(n6231) );
  MUX2_X2 U6601 ( .A(n4337), .B(n6231), .S(n4899), .Z(n6232) );
  INV_X4 U6602 ( .A(n6232), .ZN(u6_N65) );
  INV_X4 U6603 ( .A(N265), .ZN(n6233) );
  MUX2_X2 U6604 ( .A(n4433), .B(n6233), .S(n4899), .Z(n6234) );
  INV_X4 U6605 ( .A(n6234), .ZN(u6_N64) );
  INV_X4 U6606 ( .A(N264), .ZN(n6235) );
  MUX2_X2 U6607 ( .A(n4430), .B(n6235), .S(n4899), .Z(n6236) );
  INV_X4 U6608 ( .A(n6236), .ZN(u6_N63) );
  INV_X4 U6609 ( .A(N263), .ZN(n6237) );
  MUX2_X2 U6610 ( .A(n4428), .B(n6237), .S(n4899), .Z(n6238) );
  INV_X4 U6611 ( .A(n6238), .ZN(u6_N62) );
  INV_X4 U6612 ( .A(N262), .ZN(n6239) );
  MUX2_X2 U6613 ( .A(n4432), .B(n6239), .S(n4899), .Z(n6240) );
  INV_X4 U6614 ( .A(n6240), .ZN(u6_N61) );
  INV_X4 U6615 ( .A(N261), .ZN(n6241) );
  MUX2_X2 U6616 ( .A(n4343), .B(n6241), .S(n4899), .Z(n6242) );
  INV_X4 U6617 ( .A(n6242), .ZN(u6_N60) );
  INV_X4 U6618 ( .A(N260), .ZN(n6243) );
  MUX2_X2 U6619 ( .A(n4348), .B(n6243), .S(n4899), .Z(n6244) );
  INV_X4 U6620 ( .A(n6244), .ZN(u6_N59) );
  INV_X4 U6621 ( .A(N259), .ZN(n6245) );
  MUX2_X2 U6622 ( .A(n6833), .B(n6245), .S(n4899), .Z(n6246) );
  INV_X4 U6623 ( .A(n6246), .ZN(u6_N58) );
  INV_X4 U6624 ( .A(N258), .ZN(n6247) );
  MUX2_X2 U6625 ( .A(n6835), .B(n6247), .S(n4899), .Z(n6248) );
  INV_X4 U6626 ( .A(n6248), .ZN(u6_N57) );
  INV_X4 U6627 ( .A(N257), .ZN(n6249) );
  MUX2_X2 U6628 ( .A(n6837), .B(n6249), .S(n4899), .Z(n6250) );
  INV_X4 U6629 ( .A(n6250), .ZN(u6_N56) );
  INV_X4 U6630 ( .A(N256), .ZN(n6251) );
  MUX2_X2 U6631 ( .A(n6839), .B(n6251), .S(n4899), .Z(n6252) );
  INV_X4 U6632 ( .A(n6252), .ZN(u6_N55) );
  NAND2_X2 U6633 ( .A1(u2_N157), .A2(n4309), .ZN(u1_N46) );
  INV_X4 U6634 ( .A(u2_N28), .ZN(n6254) );
  INV_X4 U6635 ( .A(u2_N16), .ZN(n6253) );
  NAND3_X4 U6636 ( .A1(fpu_op_r1[1]), .A2(fpu_op_r1[0]), .A3(n4352), .ZN(n6409) );
  MUX2_X2 U6637 ( .A(n6254), .B(n6253), .S(n4854), .Z(n6341) );
  INV_X4 U6638 ( .A(n6341), .ZN(u2_exp_tmp4_10_) );
  INV_X4 U6639 ( .A(u2_N20), .ZN(n6256) );
  INV_X4 U6640 ( .A(u2_N8), .ZN(n6255) );
  MUX2_X2 U6641 ( .A(n6256), .B(n6255), .S(n4854), .Z(u2_exp_tmp4_2_) );
  INV_X4 U6642 ( .A(u2_exp_tmp4_2_), .ZN(n6332) );
  INV_X4 U6643 ( .A(u2_N19), .ZN(n6417) );
  INV_X4 U6644 ( .A(u2_N7), .ZN(n6430) );
  MUX2_X2 U6645 ( .A(n6417), .B(n6430), .S(n4854), .Z(u2_exp_tmp4_1_) );
  INV_X4 U6646 ( .A(u2_exp_tmp4_1_), .ZN(n6336) );
  INV_X4 U6647 ( .A(u2_N18), .ZN(n6416) );
  INV_X4 U6648 ( .A(u2_N6), .ZN(n6429) );
  MUX2_X2 U6649 ( .A(n6416), .B(n6429), .S(n4854), .Z(u2_exp_tmp4_0_) );
  INV_X4 U6650 ( .A(u2_exp_tmp4_0_), .ZN(n6401) );
  INV_X4 U6651 ( .A(n6329), .ZN(n6322) );
  INV_X4 U6652 ( .A(u2_N21), .ZN(n6258) );
  INV_X4 U6653 ( .A(u2_N9), .ZN(n6257) );
  MUX2_X2 U6654 ( .A(n6258), .B(n6257), .S(n4854), .Z(u2_exp_tmp4_3_) );
  INV_X4 U6655 ( .A(u2_exp_tmp4_3_), .ZN(n6323) );
  NAND2_X2 U6656 ( .A1(n6322), .A2(n6323), .ZN(n6315) );
  INV_X4 U6657 ( .A(n6315), .ZN(n6261) );
  INV_X4 U6658 ( .A(u2_N22), .ZN(n6260) );
  INV_X4 U6659 ( .A(u2_N10), .ZN(n6259) );
  MUX2_X2 U6660 ( .A(n6260), .B(n6259), .S(n4854), .Z(u2_exp_tmp4_4_) );
  INV_X4 U6661 ( .A(u2_exp_tmp4_4_), .ZN(n6319) );
  NAND2_X2 U6662 ( .A1(n6261), .A2(n6319), .ZN(n6316) );
  INV_X4 U6663 ( .A(n6316), .ZN(n6369) );
  INV_X4 U6664 ( .A(u2_N23), .ZN(n6263) );
  INV_X4 U6665 ( .A(u2_N11), .ZN(n6262) );
  MUX2_X2 U6666 ( .A(n6263), .B(n6262), .S(n4854), .Z(u2_exp_tmp4_5_) );
  INV_X4 U6667 ( .A(u2_exp_tmp4_5_), .ZN(n6370) );
  NAND2_X2 U6668 ( .A1(n6369), .A2(n6370), .ZN(n6368) );
  INV_X4 U6669 ( .A(n6368), .ZN(n6264) );
  INV_X4 U6670 ( .A(u2_N24), .ZN(n6412) );
  INV_X4 U6671 ( .A(u2_N12), .ZN(n6425) );
  MUX2_X2 U6672 ( .A(n6412), .B(n6425), .S(n4854), .Z(u2_exp_tmp4_6_) );
  INV_X4 U6673 ( .A(u2_exp_tmp4_6_), .ZN(n6306) );
  NAND2_X2 U6674 ( .A1(n6264), .A2(n6306), .ZN(n6304) );
  INV_X4 U6675 ( .A(n6304), .ZN(n6357) );
  INV_X4 U6676 ( .A(u2_N25), .ZN(n6411) );
  INV_X4 U6677 ( .A(u2_N13), .ZN(n6424) );
  MUX2_X2 U6678 ( .A(n6411), .B(n6424), .S(n4854), .Z(u2_exp_tmp4_7_) );
  INV_X4 U6679 ( .A(u2_exp_tmp4_7_), .ZN(n6358) );
  NAND2_X2 U6680 ( .A1(n6357), .A2(n6358), .ZN(n6356) );
  INV_X4 U6681 ( .A(n6356), .ZN(n6265) );
  INV_X4 U6682 ( .A(u2_N26), .ZN(n6413) );
  INV_X4 U6683 ( .A(u2_N14), .ZN(n6426) );
  MUX2_X2 U6684 ( .A(n6413), .B(n6426), .S(n4854), .Z(u2_exp_tmp4_8_) );
  INV_X4 U6685 ( .A(u2_exp_tmp4_8_), .ZN(n6295) );
  NAND2_X2 U6686 ( .A1(n6265), .A2(n6295), .ZN(n6293) );
  INV_X4 U6687 ( .A(n6293), .ZN(n6286) );
  INV_X4 U6688 ( .A(u2_N27), .ZN(n6414) );
  INV_X4 U6689 ( .A(u2_N15), .ZN(n6427) );
  MUX2_X2 U6690 ( .A(n6414), .B(n6427), .S(n4854), .Z(u2_exp_tmp4_9_) );
  INV_X4 U6691 ( .A(u2_exp_tmp4_9_), .ZN(n6287) );
  NAND2_X2 U6692 ( .A1(n6286), .A2(n6287), .ZN(n6338) );
  NAND2_X2 U6693 ( .A1(n6341), .A2(n6338), .ZN(n6467) );
  NAND2_X2 U6694 ( .A1(u2_exp_tmp4_2_), .A2(u2_exp_tmp4_1_), .ZN(n6330) );
  INV_X4 U6695 ( .A(n6330), .ZN(n6266) );
  NAND2_X2 U6696 ( .A1(n6266), .A2(u2_exp_tmp4_0_), .ZN(n6324) );
  NOR2_X4 U6697 ( .A1(n6323), .A2(n6324), .ZN(n6318) );
  INV_X4 U6698 ( .A(n6318), .ZN(n6325) );
  NOR2_X4 U6699 ( .A1(n6319), .A2(n6325), .ZN(n6309) );
  INV_X4 U6700 ( .A(n6309), .ZN(n6267) );
  NOR2_X4 U6701 ( .A1(n6370), .A2(n6267), .ZN(n6312) );
  INV_X4 U6702 ( .A(n6312), .ZN(n6268) );
  NOR2_X4 U6703 ( .A1(n6306), .A2(n6268), .ZN(n6298) );
  INV_X4 U6704 ( .A(n6298), .ZN(n6269) );
  NOR2_X4 U6705 ( .A1(n6358), .A2(n6269), .ZN(n6301) );
  INV_X4 U6706 ( .A(n6301), .ZN(n6270) );
  NOR2_X4 U6707 ( .A1(n6295), .A2(n6270), .ZN(n6290) );
  INV_X4 U6708 ( .A(n6290), .ZN(n6271) );
  NOR2_X4 U6709 ( .A1(n6287), .A2(n6271), .ZN(n6288) );
  INV_X4 U6710 ( .A(n6288), .ZN(n6273) );
  XNOR2_X2 U6711 ( .A(n4854), .B(u2_exp_tmp4_10_), .ZN(n6274) );
  MUX2_X2 U6712 ( .A(n6338), .B(n6273), .S(n4854), .Z(n6280) );
  NAND2_X2 U6713 ( .A1(n6274), .A2(n6280), .ZN(n6277) );
  INV_X4 U6714 ( .A(u2_N29), .ZN(n6276) );
  INV_X4 U6715 ( .A(u2_N17), .ZN(n6275) );
  MUX2_X2 U6716 ( .A(n6276), .B(n6275), .S(n4854), .Z(n6469) );
  MUX2_X2 U6717 ( .A(n6278), .B(n6277), .S(n6469), .Z(n6406) );
  NAND2_X2 U6718 ( .A1(n6338), .A2(n6409), .ZN(n6279) );
  MUX2_X2 U6719 ( .A(n6280), .B(n6279), .S(u2_exp_tmp4_10_), .Z(n6282) );
  NAND2_X2 U6720 ( .A1(n6282), .A2(n6281), .ZN(n6283) );
  INV_X4 U6721 ( .A(n6283), .ZN(n8290) );
  INV_X4 U6722 ( .A(n4853), .ZN(n6711) );
  NAND3_X2 U6723 ( .A1(n8290), .A2(n6711), .A3(n6284), .ZN(n6285) );
  NAND2_X2 U6724 ( .A1(n6406), .A2(n6285), .ZN(u2_exp_ovf_d_1_) );
  XNOR2_X2 U6725 ( .A(n6287), .B(n6286), .ZN(n6347) );
  INV_X4 U6726 ( .A(n6347), .ZN(n6292) );
  INV_X4 U6727 ( .A(n6288), .ZN(n6289) );
  MUX2_X2 U6728 ( .A(n6292), .B(n6291), .S(n6272), .Z(n8291) );
  NAND2_X2 U6729 ( .A1(u2_exp_tmp4_8_), .A2(n6356), .ZN(n6294) );
  NAND2_X2 U6730 ( .A1(n6294), .A2(n6293), .ZN(n6352) );
  XNOR2_X2 U6731 ( .A(n6295), .B(n6301), .ZN(n6296) );
  MUX2_X2 U6732 ( .A(n6352), .B(n6296), .S(n6272), .Z(n6297) );
  INV_X4 U6733 ( .A(n6297), .ZN(n8292) );
  NAND2_X2 U6734 ( .A1(n6357), .A2(n6409), .ZN(n6300) );
  MUX2_X2 U6735 ( .A(n6357), .B(n6298), .S(n6272), .Z(n6299) );
  MUX2_X2 U6736 ( .A(n6300), .B(n6299), .S(n6358), .Z(n6303) );
  NAND2_X2 U6737 ( .A1(n6272), .A2(n6301), .ZN(n6302) );
  NAND2_X2 U6738 ( .A1(n6303), .A2(n6302), .ZN(n8293) );
  NAND2_X2 U6739 ( .A1(u2_exp_tmp4_6_), .A2(n6368), .ZN(n6305) );
  NAND2_X2 U6740 ( .A1(n6305), .A2(n6304), .ZN(n6364) );
  XNOR2_X2 U6741 ( .A(n6306), .B(n6312), .ZN(n6307) );
  MUX2_X2 U6742 ( .A(n6364), .B(n6307), .S(n6272), .Z(n6308) );
  INV_X4 U6743 ( .A(n6308), .ZN(n8294) );
  NAND2_X2 U6744 ( .A1(n6369), .A2(n6409), .ZN(n6311) );
  MUX2_X2 U6745 ( .A(n6369), .B(n6309), .S(n6272), .Z(n6310) );
  MUX2_X2 U6746 ( .A(n6311), .B(n6310), .S(n6370), .Z(n6314) );
  NAND2_X2 U6747 ( .A1(n6272), .A2(n6312), .ZN(n6313) );
  NAND2_X2 U6748 ( .A1(n6314), .A2(n6313), .ZN(n8295) );
  NAND2_X2 U6749 ( .A1(u2_exp_tmp4_4_), .A2(n6315), .ZN(n6317) );
  NAND2_X2 U6750 ( .A1(n6317), .A2(n6316), .ZN(n6375) );
  XNOR2_X2 U6751 ( .A(n6319), .B(n6318), .ZN(n6320) );
  MUX2_X2 U6752 ( .A(n6375), .B(n6320), .S(n6272), .Z(n6321) );
  INV_X4 U6753 ( .A(n6321), .ZN(n8296) );
  XNOR2_X2 U6754 ( .A(n6323), .B(n6322), .ZN(n6380) );
  INV_X4 U6755 ( .A(n6380), .ZN(n6328) );
  NAND2_X2 U6756 ( .A1(n6324), .A2(n6323), .ZN(n6326) );
  NAND2_X2 U6757 ( .A1(n6326), .A2(n6325), .ZN(n6327) );
  MUX2_X2 U6758 ( .A(n6328), .B(n6327), .S(n6272), .Z(n8297) );
  NAND2_X2 U6759 ( .A1(n6330), .A2(n6329), .ZN(n6385) );
  MUX2_X2 U6760 ( .A(n6336), .B(n6331), .S(n6332), .Z(n6334) );
  MUX2_X2 U6761 ( .A(n6334), .B(n6333), .S(n6401), .Z(n6335) );
  NOR2_X4 U6762 ( .A1(n4477), .A2(n6335), .ZN(n8298) );
  XNOR2_X2 U6763 ( .A(n6401), .B(n6336), .ZN(n6394) );
  INV_X4 U6764 ( .A(n6394), .ZN(n6337) );
  INV_X4 U6765 ( .A(n6338), .ZN(n6339) );
  XNOR2_X2 U6766 ( .A(n6339), .B(u2_exp_tmp4_10_), .ZN(n6340) );
  INV_X4 U6767 ( .A(u1_N46), .ZN(n6468) );
  NAND2_X2 U6768 ( .A1(u2_exp_ovf_d_1_), .A2(n6468), .ZN(n6393) );
  NOR2_X4 U6769 ( .A1(u2_exp_ovf_d_1_), .A2(n6468), .ZN(n6399) );
  NAND2_X2 U6770 ( .A1(u2_exp_tmp3_10_), .A2(n6399), .ZN(n6345) );
  AOI22_X2 U6771 ( .A1(u2_N64), .A2(n4844), .B1(n4845), .B2(n8290), .ZN(n6344)
         );
  NAND3_X2 U6772 ( .A1(n6346), .A2(n6345), .A3(n6344), .ZN(u2_N86) );
  AOI22_X2 U6773 ( .A1(n6347), .A2(n6361), .B1(n6379), .B2(u2_exp_tmp4_9_), 
        .ZN(n6351) );
  NAND2_X2 U6774 ( .A1(u2_exp_tmp3_9_), .A2(n6399), .ZN(n6350) );
  NAND2_X2 U6775 ( .A1(u2_N63), .A2(n4844), .ZN(n6349) );
  NAND2_X2 U6776 ( .A1(n8291), .A2(n4845), .ZN(n6348) );
  NAND4_X2 U6777 ( .A1(n6351), .A2(n6350), .A3(n6349), .A4(n6348), .ZN(u2_N85)
         );
  INV_X4 U6778 ( .A(n6402), .ZN(n6389) );
  AOI22_X2 U6779 ( .A1(n6389), .A2(n6352), .B1(n8292), .B2(n4845), .ZN(n6355)
         );
  INV_X4 U6780 ( .A(n6393), .ZN(n6400) );
  NAND2_X2 U6781 ( .A1(n6400), .A2(u2_exp_tmp4_8_), .ZN(n6354) );
  AOI22_X2 U6782 ( .A1(u2_exp_tmp3_8_), .A2(n6399), .B1(u2_N62), .B2(n4844), 
        .ZN(n6353) );
  NAND3_X2 U6783 ( .A1(n6355), .A2(n6354), .A3(n6353), .ZN(u2_N84) );
  INV_X4 U6784 ( .A(n6402), .ZN(n6361) );
  NAND2_X2 U6785 ( .A1(n6363), .A2(n6362), .ZN(u2_N83) );
  AOI22_X2 U6786 ( .A1(n6389), .A2(n6364), .B1(n8294), .B2(n4845), .ZN(n6367)
         );
  NAND2_X2 U6787 ( .A1(n6400), .A2(u2_exp_tmp4_6_), .ZN(n6366) );
  AOI22_X2 U6788 ( .A1(u2_exp_tmp3_6_), .A2(n6399), .B1(u2_N60), .B2(n4844), 
        .ZN(n6365) );
  NAND3_X2 U6789 ( .A1(n6367), .A2(n6366), .A3(n6365), .ZN(u2_N82) );
  NAND2_X2 U6790 ( .A1(n6374), .A2(n6373), .ZN(u2_N81) );
  AOI22_X2 U6791 ( .A1(n6389), .A2(n6375), .B1(n4845), .B2(n8296), .ZN(n6378)
         );
  NAND2_X2 U6792 ( .A1(n6400), .A2(u2_exp_tmp4_4_), .ZN(n6377) );
  AOI22_X2 U6793 ( .A1(u2_exp_tmp3_4_), .A2(n6399), .B1(u2_N58), .B2(n4844), 
        .ZN(n6376) );
  NAND3_X2 U6794 ( .A1(n6378), .A2(n6377), .A3(n6376), .ZN(u2_N80) );
  AOI22_X2 U6795 ( .A1(n4845), .A2(n8297), .B1(u2_N57), .B2(n4844), .ZN(n6384)
         );
  NAND2_X2 U6796 ( .A1(u2_exp_tmp3_3_), .A2(n6399), .ZN(n6383) );
  INV_X4 U6797 ( .A(n6393), .ZN(n6379) );
  NAND2_X2 U6798 ( .A1(n6379), .A2(u2_exp_tmp4_3_), .ZN(n6382) );
  NAND2_X2 U6799 ( .A1(n6361), .A2(n6380), .ZN(n6381) );
  NAND4_X2 U6800 ( .A1(n6384), .A2(n6383), .A3(n6382), .A4(n6381), .ZN(u2_N79)
         );
  INV_X4 U6801 ( .A(n6385), .ZN(n6387) );
  NAND2_X2 U6802 ( .A1(u2_exp_tmp4_2_), .A2(u2_exp_tmp4_0_), .ZN(n6386) );
  NAND2_X2 U6803 ( .A1(n6387), .A2(n6386), .ZN(n6388) );
  AOI22_X2 U6804 ( .A1(n6389), .A2(n6388), .B1(n8298), .B2(n4845), .ZN(n6392)
         );
  NAND2_X2 U6805 ( .A1(n6400), .A2(u2_exp_tmp4_2_), .ZN(n6391) );
  AOI22_X2 U6806 ( .A1(u2_exp_tmp3_2_), .A2(n6399), .B1(u2_N56), .B2(n4844), 
        .ZN(n6390) );
  NAND3_X2 U6807 ( .A1(n6392), .A2(n6391), .A3(n6390), .ZN(u2_N78) );
  AOI22_X2 U6808 ( .A1(n4845), .A2(n4318), .B1(u2_N55), .B2(n4844), .ZN(n6398)
         );
  NAND2_X2 U6809 ( .A1(u2_exp_tmp3_1_), .A2(n6399), .ZN(n6397) );
  NAND2_X2 U6810 ( .A1(n6379), .A2(u2_exp_tmp4_1_), .ZN(n6396) );
  NAND2_X2 U6811 ( .A1(n6389), .A2(n6394), .ZN(n6395) );
  NAND4_X2 U6812 ( .A1(n6398), .A2(n6397), .A3(n6396), .A4(n6395), .ZN(u2_N77)
         );
  AOI22_X2 U6813 ( .A1(u2_exp_tmp3_0_), .A2(n6399), .B1(u2_N54), .B2(n4844), 
        .ZN(n6405) );
  NOR2_X4 U6814 ( .A1(n6400), .A2(n4845), .ZN(n6403) );
  MUX2_X2 U6815 ( .A(n6403), .B(n6402), .S(n6401), .Z(n6404) );
  NAND2_X2 U6816 ( .A1(n6405), .A2(n6404), .ZN(u2_N76) );
  INV_X4 U6817 ( .A(n6406), .ZN(n6407) );
  NAND2_X2 U6818 ( .A1(n6407), .A2(n6409), .ZN(n6408) );
  MUX2_X2 U6819 ( .A(n6409), .B(n6408), .S(opb_r[62]), .Z(n6410) );
  AND2_X2 U6820 ( .A1(u2_N22), .A2(u2_N21), .ZN(n6415) );
  NAND2_X2 U6821 ( .A1(u2_N23), .A2(n6415), .ZN(n6420) );
  NAND2_X2 U6822 ( .A1(u2_N20), .A2(n6418), .ZN(n6419) );
  NAND3_X2 U6823 ( .A1(n6423), .A2(n6422), .A3(n6421), .ZN(n6438) );
  AND2_X2 U6824 ( .A1(u2_N10), .A2(u2_N9), .ZN(n6428) );
  NAND2_X2 U6825 ( .A1(u2_N11), .A2(n6428), .ZN(n6433) );
  NAND2_X2 U6826 ( .A1(u2_N8), .A2(n6431), .ZN(n6432) );
  NAND3_X2 U6827 ( .A1(n6436), .A2(n6435), .A3(n6434), .ZN(n6437) );
  MUX2_X2 U6828 ( .A(n6438), .B(n6437), .S(n6272), .Z(n6463) );
  INV_X4 U6829 ( .A(n6439), .ZN(n6440) );
  NAND4_X2 U6830 ( .A1(n6449), .A2(n6448), .A3(n6447), .A4(n6446), .ZN(n6454)
         );
  INV_X4 U6831 ( .A(fracta_mul[44]), .ZN(n6451) );
  NAND2_X2 U6832 ( .A1(n7198), .A2(n4297), .ZN(n7153) );
  NOR4_X2 U6833 ( .A1(u6_N17), .A2(u6_N16), .A3(u6_N15), .A4(u6_N11), .ZN(
        n6461) );
  NAND3_X2 U6834 ( .A1(n3098), .A2(n3106), .A3(n6456), .ZN(n6458) );
  NAND2_X2 U6835 ( .A1(n3096), .A2(n3097), .ZN(n6457) );
  INV_X4 U6836 ( .A(n4309), .ZN(n7209) );
  NAND2_X2 U6837 ( .A1(n4346), .A2(n7209), .ZN(n6462) );
  NAND2_X2 U6838 ( .A1(n7153), .A2(n4899), .ZN(n6464) );
  INV_X4 U6839 ( .A(n6467), .ZN(n6470) );
  NOR2_X4 U6840 ( .A1(n6470), .A2(n6469), .ZN(n6472) );
  MUX2_X2 U6841 ( .A(n6472), .B(n6471), .S(n4854), .Z(u2_N114) );
  NAND4_X2 U6842 ( .A1(n6476), .A2(n6475), .A3(n6474), .A4(n6473), .ZN(N340)
         );
  NAND2_X2 U6843 ( .A1(fpu_op_r2[0]), .A2(fpu_op_r2[2]), .ZN(n4262) );
  INV_X4 U6844 ( .A(n4262), .ZN(n6477) );
  MUX2_X2 U6845 ( .A(n4356), .B(n4481), .S(fpu_op_r2[1]), .Z(n7196) );
  INV_X4 U6846 ( .A(n7196), .ZN(n6578) );
  INV_X4 U6847 ( .A(n8510), .ZN(n6478) );
  NAND2_X2 U6848 ( .A1(n6578), .A2(n6478), .ZN(n6480) );
  INV_X4 U6849 ( .A(N343), .ZN(n6479) );
  NAND2_X2 U6850 ( .A1(n7196), .A2(n6478), .ZN(n6481) );
  OAI22_X2 U6851 ( .A1(n6480), .A2(n6479), .B1(n6481), .B2(n4491), .ZN(n8509)
         );
  NAND2_X2 U6852 ( .A1(N344), .A2(n4860), .ZN(n6483) );
  INV_X4 U6853 ( .A(n6481), .ZN(n6599) );
  NAND2_X2 U6854 ( .A1(opa_r1[1]), .A2(n4857), .ZN(n6482) );
  NAND2_X2 U6855 ( .A1(n6483), .A2(n6482), .ZN(n8289) );
  NAND2_X2 U6856 ( .A1(N345), .A2(n4860), .ZN(n6485) );
  NAND2_X2 U6857 ( .A1(opa_r1[2]), .A2(n4856), .ZN(n6484) );
  NAND2_X2 U6858 ( .A1(n6485), .A2(n6484), .ZN(n8288) );
  NAND2_X2 U6859 ( .A1(N346), .A2(n4860), .ZN(n6487) );
  NAND2_X2 U6860 ( .A1(opa_r1[3]), .A2(n4855), .ZN(n6486) );
  NAND2_X2 U6861 ( .A1(n6487), .A2(n6486), .ZN(n8287) );
  NAND2_X2 U6862 ( .A1(N347), .A2(n4860), .ZN(n6489) );
  NAND2_X2 U6863 ( .A1(opa_r1[4]), .A2(n4856), .ZN(n6488) );
  NAND2_X2 U6864 ( .A1(n6489), .A2(n6488), .ZN(n8286) );
  NAND2_X2 U6865 ( .A1(N348), .A2(n4860), .ZN(n6491) );
  NAND2_X2 U6866 ( .A1(opa_r1[5]), .A2(n4857), .ZN(n6490) );
  NAND2_X2 U6867 ( .A1(n6491), .A2(n6490), .ZN(n8285) );
  NAND2_X2 U6868 ( .A1(N349), .A2(n4860), .ZN(n6493) );
  NAND2_X2 U6869 ( .A1(n4855), .A2(opa_r1[6]), .ZN(n6492) );
  NAND2_X2 U6870 ( .A1(n6493), .A2(n6492), .ZN(n8284) );
  NAND2_X2 U6871 ( .A1(N350), .A2(n4860), .ZN(n6495) );
  NAND2_X2 U6872 ( .A1(n4856), .A2(opa_r1[7]), .ZN(n6494) );
  NAND2_X2 U6873 ( .A1(n6495), .A2(n6494), .ZN(n8283) );
  NAND2_X2 U6874 ( .A1(N351), .A2(n4860), .ZN(n6497) );
  NAND2_X2 U6875 ( .A1(n4857), .A2(opa_r1[8]), .ZN(n6496) );
  NAND2_X2 U6876 ( .A1(n6497), .A2(n6496), .ZN(n8282) );
  NAND2_X2 U6877 ( .A1(N352), .A2(n4860), .ZN(n6499) );
  NAND2_X2 U6878 ( .A1(n4857), .A2(opa_r1[9]), .ZN(n6498) );
  NAND2_X2 U6879 ( .A1(n6499), .A2(n6498), .ZN(n8281) );
  NAND2_X2 U6880 ( .A1(N353), .A2(n4859), .ZN(n6501) );
  NAND2_X2 U6881 ( .A1(n4857), .A2(opa_r1[10]), .ZN(n6500) );
  NAND2_X2 U6882 ( .A1(n6501), .A2(n6500), .ZN(n8280) );
  NAND2_X2 U6883 ( .A1(N354), .A2(n4859), .ZN(n6503) );
  NAND2_X2 U6884 ( .A1(n4857), .A2(opa_r1[11]), .ZN(n6502) );
  NAND2_X2 U6885 ( .A1(n6503), .A2(n6502), .ZN(n8279) );
  NAND2_X2 U6886 ( .A1(N355), .A2(n4859), .ZN(n6505) );
  NAND2_X2 U6887 ( .A1(n4857), .A2(opa_r1[12]), .ZN(n6504) );
  NAND2_X2 U6888 ( .A1(n6505), .A2(n6504), .ZN(n8278) );
  NAND2_X2 U6889 ( .A1(N356), .A2(n4859), .ZN(n6507) );
  NAND2_X2 U6890 ( .A1(n4857), .A2(opa_r1[13]), .ZN(n6506) );
  NAND2_X2 U6891 ( .A1(n6507), .A2(n6506), .ZN(n8277) );
  NAND2_X2 U6892 ( .A1(N357), .A2(n4859), .ZN(n6509) );
  NAND2_X2 U6893 ( .A1(n4857), .A2(opa_r1[14]), .ZN(n6508) );
  NAND2_X2 U6894 ( .A1(n6509), .A2(n6508), .ZN(n8276) );
  NAND2_X2 U6895 ( .A1(N358), .A2(n4859), .ZN(n6511) );
  NAND2_X2 U6896 ( .A1(n4857), .A2(opa_r1[15]), .ZN(n6510) );
  NAND2_X2 U6897 ( .A1(n6511), .A2(n6510), .ZN(n8275) );
  NAND2_X2 U6898 ( .A1(N359), .A2(n4859), .ZN(n6513) );
  NAND2_X2 U6899 ( .A1(n4857), .A2(opa_r1[16]), .ZN(n6512) );
  NAND2_X2 U6900 ( .A1(n6513), .A2(n6512), .ZN(n8274) );
  NAND2_X2 U6901 ( .A1(N360), .A2(n4859), .ZN(n6515) );
  NAND2_X2 U6902 ( .A1(n4857), .A2(opa_r1[17]), .ZN(n6514) );
  NAND2_X2 U6903 ( .A1(n6515), .A2(n6514), .ZN(n8273) );
  NAND2_X2 U6904 ( .A1(N361), .A2(n4859), .ZN(n6517) );
  NAND2_X2 U6905 ( .A1(n4857), .A2(opa_r1[18]), .ZN(n6516) );
  NAND2_X2 U6906 ( .A1(n6517), .A2(n6516), .ZN(n8272) );
  NAND2_X2 U6907 ( .A1(N362), .A2(n4859), .ZN(n6519) );
  NAND2_X2 U6908 ( .A1(n4857), .A2(opa_r1[19]), .ZN(n6518) );
  NAND2_X2 U6909 ( .A1(n6519), .A2(n6518), .ZN(n8271) );
  NAND2_X2 U6910 ( .A1(N363), .A2(n4859), .ZN(n6521) );
  NAND2_X2 U6911 ( .A1(n4856), .A2(opa_r1[20]), .ZN(n6520) );
  NAND2_X2 U6912 ( .A1(n6521), .A2(n6520), .ZN(n8270) );
  NAND2_X2 U6913 ( .A1(N364), .A2(n4859), .ZN(n6523) );
  NAND2_X2 U6914 ( .A1(n4856), .A2(opa_r1[21]), .ZN(n6522) );
  NAND2_X2 U6915 ( .A1(n6523), .A2(n6522), .ZN(n8269) );
  NAND2_X2 U6916 ( .A1(N365), .A2(n4859), .ZN(n6525) );
  NAND2_X2 U6917 ( .A1(n4856), .A2(opa_r1[22]), .ZN(n6524) );
  NAND2_X2 U6918 ( .A1(n6525), .A2(n6524), .ZN(n8268) );
  NAND2_X2 U6919 ( .A1(N366), .A2(n4859), .ZN(n6527) );
  NAND2_X2 U6920 ( .A1(n4856), .A2(opa_r1[23]), .ZN(n6526) );
  NAND2_X2 U6921 ( .A1(n6527), .A2(n6526), .ZN(n8267) );
  NAND2_X2 U6922 ( .A1(N367), .A2(n4859), .ZN(n6529) );
  NAND2_X2 U6923 ( .A1(n4856), .A2(opa_r1[24]), .ZN(n6528) );
  NAND2_X2 U6924 ( .A1(n6529), .A2(n6528), .ZN(n8266) );
  NAND2_X2 U6925 ( .A1(N368), .A2(n4859), .ZN(n6531) );
  NAND2_X2 U6926 ( .A1(n4856), .A2(opa_r1[25]), .ZN(n6530) );
  NAND2_X2 U6927 ( .A1(n6531), .A2(n6530), .ZN(n8265) );
  NAND2_X2 U6928 ( .A1(N369), .A2(n4859), .ZN(n6533) );
  NAND2_X2 U6929 ( .A1(n4856), .A2(opa_r1[26]), .ZN(n6532) );
  NAND2_X2 U6930 ( .A1(n6533), .A2(n6532), .ZN(n8264) );
  NAND2_X2 U6931 ( .A1(N370), .A2(n4859), .ZN(n6535) );
  NAND2_X2 U6932 ( .A1(n4856), .A2(opa_r1[27]), .ZN(n6534) );
  NAND2_X2 U6933 ( .A1(n6535), .A2(n6534), .ZN(n8263) );
  NAND2_X2 U6934 ( .A1(N371), .A2(n4859), .ZN(n6537) );
  NAND2_X2 U6935 ( .A1(n4856), .A2(opa_r1[28]), .ZN(n6536) );
  NAND2_X2 U6936 ( .A1(n6537), .A2(n6536), .ZN(n8262) );
  NAND2_X2 U6937 ( .A1(N372), .A2(n4859), .ZN(n6539) );
  NAND2_X2 U6938 ( .A1(n4856), .A2(opa_r1[29]), .ZN(n6538) );
  NAND2_X2 U6939 ( .A1(n6539), .A2(n6538), .ZN(n8261) );
  NAND2_X2 U6940 ( .A1(N373), .A2(n4859), .ZN(n6541) );
  NAND2_X2 U6941 ( .A1(n4856), .A2(opa_r1[30]), .ZN(n6540) );
  NAND2_X2 U6942 ( .A1(n6541), .A2(n6540), .ZN(n8260) );
  NAND2_X2 U6943 ( .A1(N374), .A2(n4859), .ZN(n6543) );
  NAND2_X2 U6944 ( .A1(n4855), .A2(opa_r1[31]), .ZN(n6542) );
  NAND2_X2 U6945 ( .A1(n6543), .A2(n6542), .ZN(n8259) );
  NAND2_X2 U6946 ( .A1(N375), .A2(n4858), .ZN(n6545) );
  NAND2_X2 U6947 ( .A1(n4855), .A2(opa_r1[32]), .ZN(n6544) );
  NAND2_X2 U6948 ( .A1(n6545), .A2(n6544), .ZN(n8258) );
  NAND2_X2 U6949 ( .A1(N376), .A2(n4858), .ZN(n6547) );
  NAND2_X2 U6950 ( .A1(n4855), .A2(opa_r1[33]), .ZN(n6546) );
  NAND2_X2 U6951 ( .A1(n6547), .A2(n6546), .ZN(n8257) );
  NAND2_X2 U6952 ( .A1(N377), .A2(n4858), .ZN(n6549) );
  NAND2_X2 U6953 ( .A1(n4855), .A2(opa_r1[34]), .ZN(n6548) );
  NAND2_X2 U6954 ( .A1(n6549), .A2(n6548), .ZN(n8256) );
  NAND2_X2 U6955 ( .A1(N378), .A2(n4858), .ZN(n6551) );
  NAND2_X2 U6956 ( .A1(n4855), .A2(opa_r1[35]), .ZN(n6550) );
  NAND2_X2 U6957 ( .A1(n6551), .A2(n6550), .ZN(n8255) );
  NAND2_X2 U6958 ( .A1(N379), .A2(n4858), .ZN(n6553) );
  NAND2_X2 U6959 ( .A1(n4855), .A2(opa_r1[36]), .ZN(n6552) );
  NAND2_X2 U6960 ( .A1(n6553), .A2(n6552), .ZN(n8254) );
  NAND2_X2 U6961 ( .A1(N380), .A2(n4858), .ZN(n6555) );
  NAND2_X2 U6962 ( .A1(n4855), .A2(opa_r1[37]), .ZN(n6554) );
  NAND2_X2 U6963 ( .A1(n6555), .A2(n6554), .ZN(n8253) );
  NAND2_X2 U6964 ( .A1(N381), .A2(n4858), .ZN(n6557) );
  NAND2_X2 U6965 ( .A1(n4855), .A2(opa_r1[38]), .ZN(n6556) );
  NAND2_X2 U6966 ( .A1(n6557), .A2(n6556), .ZN(n8252) );
  NAND2_X2 U6967 ( .A1(N382), .A2(n4858), .ZN(n6559) );
  NAND2_X2 U6968 ( .A1(n4855), .A2(opa_r1[39]), .ZN(n6558) );
  NAND2_X2 U6969 ( .A1(n6559), .A2(n6558), .ZN(n8251) );
  NAND2_X2 U6970 ( .A1(N383), .A2(n4858), .ZN(n6561) );
  NAND2_X2 U6971 ( .A1(n4855), .A2(opa_r1[40]), .ZN(n6560) );
  NAND2_X2 U6972 ( .A1(n6561), .A2(n6560), .ZN(n8250) );
  NAND2_X2 U6973 ( .A1(N384), .A2(n4858), .ZN(n6563) );
  NAND2_X2 U6974 ( .A1(n4855), .A2(opa_r1[41]), .ZN(n6562) );
  NAND2_X2 U6975 ( .A1(n6563), .A2(n6562), .ZN(n8249) );
  NAND2_X2 U6976 ( .A1(N385), .A2(n4858), .ZN(n6565) );
  NAND2_X2 U6977 ( .A1(n6599), .A2(opa_r1[42]), .ZN(n6564) );
  NAND2_X2 U6978 ( .A1(n6565), .A2(n6564), .ZN(n8248) );
  NAND2_X2 U6979 ( .A1(N386), .A2(n4859), .ZN(n6567) );
  NAND2_X2 U6980 ( .A1(n6599), .A2(opa_r1[43]), .ZN(n6566) );
  NAND2_X2 U6981 ( .A1(n6567), .A2(n6566), .ZN(n8247) );
  NAND2_X2 U6982 ( .A1(N387), .A2(n4859), .ZN(n6569) );
  NAND2_X2 U6983 ( .A1(n6599), .A2(opa_r1[44]), .ZN(n6568) );
  NAND2_X2 U6984 ( .A1(n6569), .A2(n6568), .ZN(n8246) );
  NAND2_X2 U6985 ( .A1(N388), .A2(n4859), .ZN(n6571) );
  NAND2_X2 U6986 ( .A1(n6599), .A2(opa_r1[45]), .ZN(n6570) );
  NAND2_X2 U6987 ( .A1(n6571), .A2(n6570), .ZN(n8245) );
  NAND2_X2 U6988 ( .A1(N389), .A2(n4859), .ZN(n6574) );
  NAND2_X2 U6989 ( .A1(n7196), .A2(n8510), .ZN(n6597) );
  NAND2_X2 U6990 ( .A1(N343), .A2(n4862), .ZN(n6573) );
  NAND2_X2 U6991 ( .A1(n6599), .A2(opa_r1[46]), .ZN(n6572) );
  NAND3_X2 U6992 ( .A1(n6574), .A2(n6573), .A3(n6572), .ZN(N710) );
  NAND2_X2 U6993 ( .A1(N390), .A2(n4859), .ZN(n6577) );
  NAND2_X2 U6994 ( .A1(opa_r1[1]), .A2(n6587), .ZN(n6576) );
  NAND2_X2 U6995 ( .A1(n6599), .A2(opa_r1[47]), .ZN(n6575) );
  NAND3_X2 U6996 ( .A1(n6577), .A2(n6576), .A3(n6575), .ZN(N711) );
  NAND2_X2 U6997 ( .A1(n6599), .A2(opa_r1[48]), .ZN(n6581) );
  NAND2_X2 U6998 ( .A1(N391), .A2(n4860), .ZN(n6580) );
  AOI22_X2 U6999 ( .A1(N343), .A2(n4864), .B1(opa_r1[2]), .B2(n6587), .ZN(
        n6579) );
  NAND3_X2 U7000 ( .A1(n6581), .A2(n6580), .A3(n6579), .ZN(N712) );
  NAND2_X2 U7001 ( .A1(N501), .A2(n4864), .ZN(n6586) );
  INV_X4 U7002 ( .A(n6597), .ZN(n6582) );
  NAND2_X2 U7003 ( .A1(opa_r1[3]), .A2(n6582), .ZN(n6585) );
  NAND2_X2 U7004 ( .A1(N392), .A2(n4858), .ZN(n6584) );
  NAND2_X2 U7005 ( .A1(n4855), .A2(opa_r1[49]), .ZN(n6583) );
  NAND4_X2 U7006 ( .A1(n6586), .A2(n6585), .A3(n6584), .A4(n6583), .ZN(N713)
         );
  NAND2_X2 U7007 ( .A1(N502), .A2(n4292), .ZN(n6591) );
  INV_X4 U7008 ( .A(n6597), .ZN(n6587) );
  NAND2_X2 U7009 ( .A1(opa_r1[4]), .A2(n6587), .ZN(n6590) );
  NAND2_X2 U7010 ( .A1(N393), .A2(n4858), .ZN(n6589) );
  NAND2_X2 U7011 ( .A1(n4855), .A2(opa_r1[50]), .ZN(n6588) );
  NAND4_X2 U7012 ( .A1(n6591), .A2(n6590), .A3(n6589), .A4(n6588), .ZN(N714)
         );
  NAND2_X2 U7013 ( .A1(N503), .A2(n4865), .ZN(n6596) );
  INV_X4 U7014 ( .A(n6597), .ZN(n6592) );
  NAND2_X2 U7015 ( .A1(opa_r1[5]), .A2(n6592), .ZN(n6595) );
  NAND2_X2 U7016 ( .A1(N394), .A2(n4858), .ZN(n6594) );
  NAND2_X2 U7017 ( .A1(n6599), .A2(opa_r1[51]), .ZN(n6593) );
  NAND4_X2 U7018 ( .A1(n6596), .A2(n6595), .A3(n6594), .A4(n6593), .ZN(N715)
         );
  NAND2_X2 U7019 ( .A1(N504), .A2(n4865), .ZN(n6603) );
  INV_X4 U7020 ( .A(n6597), .ZN(n6598) );
  NAND2_X2 U7021 ( .A1(opa_r1[6]), .A2(n6598), .ZN(n6602) );
  NAND2_X2 U7022 ( .A1(N395), .A2(n4858), .ZN(n6601) );
  NAND2_X2 U7023 ( .A1(n4855), .A2(N340), .ZN(n6600) );
  NAND4_X2 U7024 ( .A1(n6603), .A2(n6602), .A3(n6601), .A4(n6600), .ZN(N716)
         );
  NAND2_X2 U7025 ( .A1(N505), .A2(n4292), .ZN(n6605) );
  NAND2_X2 U7026 ( .A1(N396), .A2(n4861), .ZN(n6708) );
  NAND2_X2 U7027 ( .A1(opa_r1[7]), .A2(n6587), .ZN(n6604) );
  NAND3_X2 U7028 ( .A1(n6605), .A2(n4873), .A3(n6604), .ZN(N717) );
  NAND2_X2 U7029 ( .A1(N506), .A2(n4292), .ZN(n6607) );
  NAND2_X2 U7030 ( .A1(opa_r1[8]), .A2(n6592), .ZN(n6606) );
  NAND3_X2 U7031 ( .A1(n6607), .A2(n4873), .A3(n6606), .ZN(N718) );
  NAND2_X2 U7032 ( .A1(N507), .A2(n4292), .ZN(n6609) );
  NAND2_X2 U7033 ( .A1(opa_r1[9]), .A2(n6598), .ZN(n6608) );
  NAND3_X2 U7034 ( .A1(n6609), .A2(n4873), .A3(n6608), .ZN(N719) );
  NAND2_X2 U7035 ( .A1(N508), .A2(n4292), .ZN(n6611) );
  NAND2_X2 U7036 ( .A1(opa_r1[10]), .A2(n6592), .ZN(n6610) );
  NAND3_X2 U7037 ( .A1(n6611), .A2(n4873), .A3(n6610), .ZN(N720) );
  NAND2_X2 U7038 ( .A1(N509), .A2(n4292), .ZN(n6613) );
  NAND2_X2 U7039 ( .A1(opa_r1[11]), .A2(n6598), .ZN(n6612) );
  NAND3_X2 U7040 ( .A1(n6613), .A2(n4873), .A3(n6612), .ZN(N721) );
  NAND2_X2 U7041 ( .A1(N510), .A2(n4292), .ZN(n6615) );
  NAND2_X2 U7042 ( .A1(opa_r1[12]), .A2(n6592), .ZN(n6614) );
  NAND3_X2 U7043 ( .A1(n6615), .A2(n4873), .A3(n6614), .ZN(N722) );
  NAND2_X2 U7044 ( .A1(N511), .A2(n4292), .ZN(n6617) );
  NAND2_X2 U7045 ( .A1(opa_r1[13]), .A2(n6598), .ZN(n6616) );
  NAND3_X2 U7046 ( .A1(n6617), .A2(n4873), .A3(n6616), .ZN(N723) );
  NAND2_X2 U7047 ( .A1(N512), .A2(n4863), .ZN(n6619) );
  NAND2_X2 U7048 ( .A1(opa_r1[14]), .A2(n6592), .ZN(n6618) );
  NAND3_X2 U7049 ( .A1(n6619), .A2(n4873), .A3(n6618), .ZN(N724) );
  NAND2_X2 U7050 ( .A1(N513), .A2(n4863), .ZN(n6621) );
  NAND2_X2 U7051 ( .A1(opa_r1[15]), .A2(n6598), .ZN(n6620) );
  NAND3_X2 U7052 ( .A1(n6621), .A2(n4873), .A3(n6620), .ZN(N725) );
  NAND2_X2 U7053 ( .A1(N514), .A2(n4863), .ZN(n6623) );
  NAND2_X2 U7054 ( .A1(opa_r1[16]), .A2(n6592), .ZN(n6622) );
  NAND3_X2 U7055 ( .A1(n6623), .A2(n4872), .A3(n6622), .ZN(N726) );
  NAND2_X2 U7056 ( .A1(N515), .A2(n4863), .ZN(n6625) );
  NAND2_X2 U7057 ( .A1(opa_r1[17]), .A2(n6598), .ZN(n6624) );
  NAND3_X2 U7058 ( .A1(n6625), .A2(n4872), .A3(n6624), .ZN(N727) );
  NAND2_X2 U7059 ( .A1(N516), .A2(n4863), .ZN(n6627) );
  NAND2_X2 U7060 ( .A1(opa_r1[18]), .A2(n6592), .ZN(n6626) );
  NAND3_X2 U7061 ( .A1(n6627), .A2(n4872), .A3(n6626), .ZN(N728) );
  NAND2_X2 U7062 ( .A1(N517), .A2(n4863), .ZN(n6629) );
  NAND2_X2 U7063 ( .A1(opa_r1[19]), .A2(n6598), .ZN(n6628) );
  NAND3_X2 U7064 ( .A1(n6629), .A2(n4872), .A3(n6628), .ZN(N729) );
  NAND2_X2 U7065 ( .A1(N518), .A2(n4863), .ZN(n6631) );
  NAND2_X2 U7066 ( .A1(opa_r1[20]), .A2(n4862), .ZN(n6630) );
  NAND3_X2 U7067 ( .A1(n6631), .A2(n4872), .A3(n6630), .ZN(N730) );
  NAND2_X2 U7068 ( .A1(N519), .A2(n4863), .ZN(n6633) );
  NAND2_X2 U7069 ( .A1(opa_r1[21]), .A2(n4862), .ZN(n6632) );
  NAND3_X2 U7070 ( .A1(n6633), .A2(n4872), .A3(n6632), .ZN(N731) );
  NAND2_X2 U7071 ( .A1(N520), .A2(n4863), .ZN(n6635) );
  NAND2_X2 U7072 ( .A1(opa_r1[22]), .A2(n4862), .ZN(n6634) );
  NAND3_X2 U7073 ( .A1(n6635), .A2(n4872), .A3(n6634), .ZN(N732) );
  NAND2_X2 U7074 ( .A1(N521), .A2(n4863), .ZN(n6637) );
  NAND2_X2 U7075 ( .A1(opa_r1[23]), .A2(n4862), .ZN(n6636) );
  NAND3_X2 U7076 ( .A1(n6637), .A2(n4872), .A3(n6636), .ZN(N733) );
  NAND2_X2 U7077 ( .A1(N522), .A2(n4863), .ZN(n6639) );
  NAND2_X2 U7078 ( .A1(opa_r1[24]), .A2(n4862), .ZN(n6638) );
  NAND3_X2 U7079 ( .A1(n6639), .A2(n4872), .A3(n6638), .ZN(N734) );
  NAND2_X2 U7080 ( .A1(N523), .A2(n4863), .ZN(n6641) );
  NAND2_X2 U7081 ( .A1(opa_r1[25]), .A2(n4862), .ZN(n6640) );
  NAND3_X2 U7082 ( .A1(n6641), .A2(n4872), .A3(n6640), .ZN(N735) );
  NAND2_X2 U7083 ( .A1(N524), .A2(n4864), .ZN(n6643) );
  NAND2_X2 U7084 ( .A1(opa_r1[26]), .A2(n4862), .ZN(n6642) );
  NAND3_X2 U7085 ( .A1(n6643), .A2(n4872), .A3(n6642), .ZN(N736) );
  NAND2_X2 U7086 ( .A1(N525), .A2(n4864), .ZN(n6645) );
  NAND2_X2 U7087 ( .A1(opa_r1[27]), .A2(n4862), .ZN(n6644) );
  NAND3_X2 U7088 ( .A1(n6645), .A2(n4871), .A3(n6644), .ZN(N737) );
  NAND2_X2 U7089 ( .A1(N526), .A2(n4864), .ZN(n6647) );
  NAND2_X2 U7090 ( .A1(opa_r1[28]), .A2(n4862), .ZN(n6646) );
  NAND3_X2 U7091 ( .A1(n6647), .A2(n4871), .A3(n6646), .ZN(N738) );
  NAND2_X2 U7092 ( .A1(N527), .A2(n4864), .ZN(n6649) );
  NAND2_X2 U7093 ( .A1(opa_r1[29]), .A2(n4862), .ZN(n6648) );
  NAND3_X2 U7094 ( .A1(n6649), .A2(n4871), .A3(n6648), .ZN(N739) );
  NAND2_X2 U7095 ( .A1(N528), .A2(n4864), .ZN(n6651) );
  NAND2_X2 U7096 ( .A1(opa_r1[30]), .A2(n4862), .ZN(n6650) );
  NAND3_X2 U7097 ( .A1(n6651), .A2(n4871), .A3(n6650), .ZN(N740) );
  NAND2_X2 U7098 ( .A1(N529), .A2(n4864), .ZN(n6653) );
  NAND2_X2 U7099 ( .A1(opa_r1[31]), .A2(n6582), .ZN(n6652) );
  NAND3_X2 U7100 ( .A1(n6653), .A2(n4871), .A3(n6652), .ZN(N741) );
  NAND2_X2 U7101 ( .A1(N530), .A2(n4864), .ZN(n6655) );
  NAND2_X2 U7102 ( .A1(opa_r1[32]), .A2(n4862), .ZN(n6654) );
  NAND3_X2 U7103 ( .A1(n6655), .A2(n4871), .A3(n6654), .ZN(N742) );
  NAND2_X2 U7104 ( .A1(N531), .A2(n4864), .ZN(n6657) );
  NAND2_X2 U7105 ( .A1(opa_r1[33]), .A2(n4862), .ZN(n6656) );
  NAND3_X2 U7106 ( .A1(n6657), .A2(n4871), .A3(n6656), .ZN(N743) );
  NAND2_X2 U7107 ( .A1(N532), .A2(n4864), .ZN(n6659) );
  NAND2_X2 U7108 ( .A1(opa_r1[34]), .A2(n4862), .ZN(n6658) );
  NAND3_X2 U7109 ( .A1(n6659), .A2(n4871), .A3(n6658), .ZN(N744) );
  NAND2_X2 U7110 ( .A1(N533), .A2(n4864), .ZN(n6661) );
  NAND2_X2 U7111 ( .A1(opa_r1[35]), .A2(n4862), .ZN(n6660) );
  NAND3_X2 U7112 ( .A1(n6661), .A2(n4871), .A3(n6660), .ZN(N745) );
  NAND2_X2 U7113 ( .A1(N534), .A2(n4864), .ZN(n6663) );
  NAND2_X2 U7114 ( .A1(opa_r1[36]), .A2(n6598), .ZN(n6662) );
  NAND3_X2 U7115 ( .A1(n6663), .A2(n4871), .A3(n6662), .ZN(N746) );
  NAND2_X2 U7116 ( .A1(N535), .A2(n4864), .ZN(n6665) );
  NAND2_X2 U7117 ( .A1(opa_r1[37]), .A2(n6592), .ZN(n6664) );
  NAND3_X2 U7118 ( .A1(n6665), .A2(n4871), .A3(n6664), .ZN(N747) );
  NAND2_X2 U7119 ( .A1(N536), .A2(n4865), .ZN(n6667) );
  NAND2_X2 U7120 ( .A1(opa_r1[38]), .A2(n4862), .ZN(n6666) );
  NAND3_X2 U7121 ( .A1(n6667), .A2(n4870), .A3(n6666), .ZN(N748) );
  NAND2_X2 U7122 ( .A1(N537), .A2(n4865), .ZN(n6669) );
  NAND2_X2 U7123 ( .A1(opa_r1[39]), .A2(n6587), .ZN(n6668) );
  NAND3_X2 U7124 ( .A1(n6669), .A2(n4870), .A3(n6668), .ZN(N749) );
  NAND2_X2 U7125 ( .A1(N538), .A2(n4865), .ZN(n6671) );
  NAND2_X2 U7126 ( .A1(opa_r1[40]), .A2(n6598), .ZN(n6670) );
  NAND3_X2 U7127 ( .A1(n6671), .A2(n4870), .A3(n6670), .ZN(N750) );
  NAND2_X2 U7128 ( .A1(N539), .A2(n4865), .ZN(n6673) );
  NAND2_X2 U7129 ( .A1(opa_r1[41]), .A2(n6592), .ZN(n6672) );
  NAND3_X2 U7130 ( .A1(n6673), .A2(n4870), .A3(n6672), .ZN(N751) );
  NAND2_X2 U7131 ( .A1(N540), .A2(n4865), .ZN(n6675) );
  NAND2_X2 U7132 ( .A1(opa_r1[42]), .A2(n6592), .ZN(n6674) );
  NAND3_X2 U7133 ( .A1(n6675), .A2(n4870), .A3(n6674), .ZN(N752) );
  NAND2_X2 U7134 ( .A1(N541), .A2(n4865), .ZN(n6677) );
  NAND2_X2 U7135 ( .A1(opa_r1[43]), .A2(n6592), .ZN(n6676) );
  NAND3_X2 U7136 ( .A1(n6677), .A2(n4870), .A3(n6676), .ZN(N753) );
  NAND2_X2 U7137 ( .A1(N542), .A2(n4865), .ZN(n6679) );
  NAND2_X2 U7138 ( .A1(opa_r1[44]), .A2(n6587), .ZN(n6678) );
  NAND3_X2 U7139 ( .A1(n6679), .A2(n4870), .A3(n6678), .ZN(N754) );
  NAND2_X2 U7140 ( .A1(N543), .A2(n4865), .ZN(n6681) );
  NAND2_X2 U7141 ( .A1(opa_r1[45]), .A2(n6582), .ZN(n6680) );
  NAND3_X2 U7142 ( .A1(n6681), .A2(n4870), .A3(n6680), .ZN(N755) );
  NAND2_X2 U7143 ( .A1(N544), .A2(n4865), .ZN(n6683) );
  NAND2_X2 U7144 ( .A1(opa_r1[46]), .A2(n6598), .ZN(n6682) );
  NAND3_X2 U7145 ( .A1(n6683), .A2(n4870), .A3(n6682), .ZN(N756) );
  NAND2_X2 U7146 ( .A1(N545), .A2(n4865), .ZN(n6685) );
  NAND2_X2 U7147 ( .A1(opa_r1[47]), .A2(n6592), .ZN(n6684) );
  NAND3_X2 U7148 ( .A1(n6685), .A2(n4870), .A3(n6684), .ZN(N757) );
  NAND2_X2 U7149 ( .A1(N546), .A2(n4865), .ZN(n6687) );
  NAND2_X2 U7150 ( .A1(opa_r1[48]), .A2(n6587), .ZN(n6686) );
  NAND3_X2 U7151 ( .A1(n6687), .A2(n4870), .A3(n6686), .ZN(N758) );
  NAND2_X2 U7152 ( .A1(N547), .A2(n4865), .ZN(n6689) );
  NAND2_X2 U7153 ( .A1(opa_r1[49]), .A2(n6582), .ZN(n6688) );
  NAND3_X2 U7154 ( .A1(n6689), .A2(n4869), .A3(n6688), .ZN(N759) );
  NAND2_X2 U7155 ( .A1(N548), .A2(n4863), .ZN(n6691) );
  NAND2_X2 U7156 ( .A1(opa_r1[50]), .A2(n6598), .ZN(n6690) );
  NAND3_X2 U7157 ( .A1(n6691), .A2(n4869), .A3(n6690), .ZN(N760) );
  NAND2_X2 U7158 ( .A1(N549), .A2(n4865), .ZN(n6693) );
  NAND2_X2 U7159 ( .A1(opa_r1[51]), .A2(n6587), .ZN(n6692) );
  NAND3_X2 U7160 ( .A1(n6693), .A2(n4869), .A3(n6692), .ZN(N761) );
  NAND2_X2 U7161 ( .A1(N550), .A2(n4863), .ZN(n6695) );
  NAND2_X2 U7162 ( .A1(n6598), .A2(opa_r1[52]), .ZN(n6694) );
  NAND3_X2 U7163 ( .A1(n6695), .A2(n4869), .A3(n6694), .ZN(N762) );
  NAND2_X2 U7164 ( .A1(N551), .A2(n4865), .ZN(n6697) );
  NAND2_X2 U7165 ( .A1(n6598), .A2(opa_r1[53]), .ZN(n6696) );
  NAND3_X2 U7166 ( .A1(n6697), .A2(n4869), .A3(n6696), .ZN(N763) );
  NAND2_X2 U7167 ( .A1(N552), .A2(n4863), .ZN(n6699) );
  NAND2_X2 U7168 ( .A1(n6592), .A2(opa_r1[54]), .ZN(n6698) );
  NAND3_X2 U7169 ( .A1(n6699), .A2(n4869), .A3(n6698), .ZN(N764) );
  NAND2_X2 U7170 ( .A1(N553), .A2(n4865), .ZN(n6701) );
  NAND2_X2 U7171 ( .A1(n6587), .A2(opa_r1[55]), .ZN(n6700) );
  NAND3_X2 U7172 ( .A1(n6701), .A2(n4869), .A3(n6700), .ZN(N765) );
  NAND2_X2 U7173 ( .A1(N554), .A2(n4863), .ZN(n6703) );
  NAND2_X2 U7174 ( .A1(n6587), .A2(opa_r1[56]), .ZN(n6702) );
  NAND3_X2 U7175 ( .A1(n6703), .A2(n4869), .A3(n6702), .ZN(N766) );
  NAND2_X2 U7176 ( .A1(N555), .A2(n4865), .ZN(n6705) );
  NAND2_X2 U7177 ( .A1(n6592), .A2(opa_r1[57]), .ZN(n6704) );
  NAND3_X2 U7178 ( .A1(n6705), .A2(n4869), .A3(n6704), .ZN(N767) );
  NAND2_X2 U7179 ( .A1(N556), .A2(n4863), .ZN(n6707) );
  NAND2_X2 U7180 ( .A1(n6587), .A2(opa_r1[58]), .ZN(n6706) );
  NAND3_X2 U7181 ( .A1(n6707), .A2(n4869), .A3(n6706), .ZN(N768) );
  NAND2_X2 U7182 ( .A1(n6598), .A2(opa_r1[59]), .ZN(n6710) );
  NAND2_X2 U7183 ( .A1(N557), .A2(n4864), .ZN(n6709) );
  NAND3_X2 U7184 ( .A1(n6710), .A2(n6709), .A3(n4869), .ZN(N769) );
  XNOR2_X2 U7185 ( .A(opb_r[63]), .B(opa_r[63]), .ZN(n6735) );
  INV_X4 U7186 ( .A(n6735), .ZN(u2_sign_d) );
  INV_X4 U7187 ( .A(opb_r[62]), .ZN(n6732) );
  NAND2_X2 U7188 ( .A1(n6732), .A2(n6711), .ZN(u1_exp_large_10_) );
  NAND3_X2 U7189 ( .A1(n6739), .A2(n6714), .A3(n6740), .ZN(n6716) );
  INV_X4 U7190 ( .A(n6743), .ZN(n6715) );
  AOI211_X4 U7191 ( .C1(n6717), .C2(n6716), .A(n6715), .B(n4398), .ZN(n6719)
         );
  NOR2_X4 U7192 ( .A1(n6719), .A2(n6718), .ZN(n6723) );
  INV_X4 U7193 ( .A(n4839), .ZN(n6759) );
  NAND2_X2 U7194 ( .A1(opa_r[57]), .A2(n6759), .ZN(n6722) );
  NAND2_X2 U7195 ( .A1(n4839), .A2(n4393), .ZN(n6744) );
  INV_X4 U7196 ( .A(n6744), .ZN(n6721) );
  INV_X4 U7197 ( .A(n6720), .ZN(n6737) );
  AOI211_X4 U7198 ( .C1(n6723), .C2(n6722), .A(n6721), .B(n6737), .ZN(n6725)
         );
  NOR2_X4 U7199 ( .A1(n6725), .A2(n6724), .ZN(n6728) );
  NAND2_X2 U7200 ( .A1(opa_r[59]), .A2(n4820), .ZN(n6727) );
  INV_X4 U7201 ( .A(n6726), .ZN(n6738) );
  AOI21_X4 U7202 ( .B1(n6728), .B2(n6727), .A(n6738), .ZN(n6731) );
  AOI211_X4 U7203 ( .C1(n6731), .C2(n6742), .A(n6730), .B(n6729), .ZN(n6734)
         );
  INV_X4 U7204 ( .A(opb_r[61]), .ZN(n6753) );
  OAI22_X2 U7205 ( .A1(n4853), .A2(n6732), .B1(opa_r[61]), .B2(n6753), .ZN(
        n6736) );
  NAND2_X2 U7206 ( .A1(n4853), .A2(n6732), .ZN(n6733) );
  OAI21_X4 U7207 ( .B1(n6734), .B2(n6736), .A(n6733), .ZN(n7138) );
  INV_X4 U7208 ( .A(n7138), .ZN(n7134) );
  AND2_X2 U7209 ( .A1(u1_N220), .A2(n4882), .ZN(n6750) );
  XNOR2_X2 U7210 ( .A(n6735), .B(n4445), .ZN(u1_N232) );
  NAND2_X2 U7211 ( .A1(opb_r[52]), .A2(n4330), .ZN(n6741) );
  NAND3_X2 U7212 ( .A1(n6741), .A2(n6740), .A3(n6739), .ZN(n6746) );
  NAND3_X2 U7213 ( .A1(n6744), .A2(n6743), .A3(n6742), .ZN(n6745) );
  NAND4_X2 U7214 ( .A1(n6750), .A2(n6749), .A3(n6748), .A4(n6747), .ZN(n6751)
         );
  INV_X4 U7215 ( .A(u1_exp_large_10_), .ZN(n6752) );
  NOR2_X4 U7216 ( .A1(n6765), .A2(n6752), .ZN(u1_N62) );
  MUX2_X2 U7217 ( .A(n4391), .B(n6753), .S(n4892), .Z(n6754) );
  INV_X4 U7218 ( .A(n6754), .ZN(n8506) );
  NOR2_X4 U7219 ( .A1(n6765), .A2(n6754), .ZN(u1_N61) );
  MUX2_X2 U7220 ( .A(n4394), .B(n4824), .S(n4892), .Z(n6755) );
  INV_X4 U7221 ( .A(n6755), .ZN(n8507) );
  NOR2_X4 U7222 ( .A1(n6765), .A2(n6755), .ZN(u1_N60) );
  MUX2_X2 U7223 ( .A(n4396), .B(n4820), .S(n4892), .Z(n6756) );
  INV_X4 U7224 ( .A(n6756), .ZN(u1_exp_large_7_) );
  NOR2_X4 U7225 ( .A1(n6765), .A2(n6756), .ZN(u1_N59) );
  MUX2_X2 U7226 ( .A(n4395), .B(n6757), .S(n4892), .Z(n6758) );
  INV_X4 U7227 ( .A(n6758), .ZN(u1_exp_large_6_) );
  NOR2_X4 U7228 ( .A1(n6765), .A2(n6758), .ZN(u1_N58) );
  MUX2_X2 U7229 ( .A(n4393), .B(n6759), .S(n4892), .Z(n6760) );
  INV_X4 U7230 ( .A(n6760), .ZN(u1_exp_large_5_) );
  NOR2_X4 U7231 ( .A1(n6765), .A2(n6760), .ZN(u1_N57) );
  MUX2_X2 U7232 ( .A(n4332), .B(n4835), .S(n4892), .Z(n6761) );
  INV_X4 U7233 ( .A(n6761), .ZN(u1_exp_large_4_) );
  NOR2_X4 U7234 ( .A1(n6765), .A2(n6761), .ZN(u1_N56) );
  INV_X4 U7235 ( .A(opb_r[55]), .ZN(n7145) );
  MUX2_X2 U7236 ( .A(n4390), .B(n7145), .S(n4891), .Z(n6762) );
  INV_X4 U7237 ( .A(n6762), .ZN(u1_exp_large_3_) );
  NOR2_X4 U7238 ( .A1(n6765), .A2(n6762), .ZN(u1_N55) );
  MUX2_X2 U7239 ( .A(n4331), .B(n7149), .S(n4891), .Z(n6763) );
  INV_X4 U7240 ( .A(n6763), .ZN(u1_exp_large_2_) );
  MUX2_X2 U7241 ( .A(n4392), .B(n7148), .S(n4891), .Z(n6764) );
  INV_X4 U7242 ( .A(n6764), .ZN(u1_exp_large_1_) );
  INV_X4 U7243 ( .A(opb_r[52]), .ZN(n7147) );
  MUX2_X2 U7244 ( .A(n4330), .B(n7147), .S(n4891), .Z(n6766) );
  INV_X4 U7245 ( .A(n6766), .ZN(u1_exp_large_0_) );
  MUX2_X2 U7246 ( .A(u3_N116), .B(u3_N59), .S(n4916), .Z(n8299) );
  MUX2_X2 U7247 ( .A(u3_N115), .B(u3_N58), .S(n4916), .Z(n8300) );
  MUX2_X2 U7248 ( .A(u3_N114), .B(u3_N57), .S(n4916), .Z(n8301) );
  MUX2_X2 U7249 ( .A(u3_N113), .B(u3_N56), .S(n4916), .Z(n8302) );
  MUX2_X2 U7250 ( .A(u3_N112), .B(u3_N55), .S(n4916), .Z(n8303) );
  MUX2_X2 U7251 ( .A(u3_N111), .B(u3_N54), .S(n4916), .Z(n8304) );
  MUX2_X2 U7252 ( .A(u3_N110), .B(u3_N53), .S(n4916), .Z(n8305) );
  MUX2_X2 U7253 ( .A(u3_N109), .B(u3_N52), .S(n4916), .Z(n8306) );
  MUX2_X2 U7254 ( .A(u3_N108), .B(u3_N51), .S(n4916), .Z(n8307) );
  MUX2_X2 U7255 ( .A(u3_N107), .B(u3_N50), .S(n4916), .Z(n8308) );
  MUX2_X2 U7256 ( .A(u3_N106), .B(u3_N49), .S(n4916), .Z(n8309) );
  MUX2_X2 U7257 ( .A(u3_N105), .B(u3_N48), .S(n4917), .Z(n8310) );
  MUX2_X2 U7258 ( .A(u3_N104), .B(u3_N47), .S(n4917), .Z(n8311) );
  MUX2_X2 U7259 ( .A(u3_N103), .B(u3_N46), .S(n4917), .Z(n8312) );
  MUX2_X2 U7260 ( .A(u3_N102), .B(u3_N45), .S(n4917), .Z(n8313) );
  MUX2_X2 U7261 ( .A(u3_N101), .B(u3_N44), .S(n4917), .Z(n8314) );
  MUX2_X2 U7262 ( .A(u3_N100), .B(u3_N43), .S(n4917), .Z(n8315) );
  MUX2_X2 U7263 ( .A(u3_N99), .B(u3_N42), .S(n4917), .Z(n8316) );
  MUX2_X2 U7264 ( .A(u3_N98), .B(u3_N41), .S(n4917), .Z(n8317) );
  MUX2_X2 U7265 ( .A(u3_N97), .B(u3_N40), .S(n4917), .Z(n8318) );
  MUX2_X2 U7266 ( .A(u3_N96), .B(u3_N39), .S(n4917), .Z(n8319) );
  MUX2_X2 U7267 ( .A(u3_N95), .B(u3_N38), .S(n4917), .Z(n8320) );
  MUX2_X2 U7268 ( .A(u3_N94), .B(u3_N37), .S(n4917), .Z(n8321) );
  MUX2_X2 U7269 ( .A(u3_N93), .B(u3_N36), .S(n4916), .Z(n8322) );
  MUX2_X2 U7270 ( .A(u3_N92), .B(u3_N35), .S(n4917), .Z(n8323) );
  MUX2_X2 U7271 ( .A(u3_N91), .B(u3_N34), .S(n4916), .Z(n8324) );
  MUX2_X2 U7272 ( .A(u3_N90), .B(u3_N33), .S(n4917), .Z(n8325) );
  MUX2_X2 U7273 ( .A(u3_N89), .B(u3_N32), .S(n4916), .Z(n8326) );
  MUX2_X2 U7274 ( .A(u3_N88), .B(u3_N31), .S(n4917), .Z(n8327) );
  MUX2_X2 U7275 ( .A(u3_N87), .B(u3_N30), .S(n4916), .Z(n8328) );
  MUX2_X2 U7276 ( .A(u3_N86), .B(u3_N29), .S(n4917), .Z(n8329) );
  MUX2_X2 U7277 ( .A(u3_N85), .B(u3_N28), .S(n4916), .Z(n8330) );
  MUX2_X2 U7278 ( .A(u3_N84), .B(u3_N27), .S(n4917), .Z(n8331) );
  MUX2_X2 U7279 ( .A(u3_N83), .B(u3_N26), .S(n4918), .Z(n8332) );
  MUX2_X2 U7280 ( .A(u3_N82), .B(u3_N25), .S(n4918), .Z(n8333) );
  MUX2_X2 U7281 ( .A(u3_N81), .B(u3_N24), .S(n4918), .Z(n8334) );
  MUX2_X2 U7282 ( .A(u3_N80), .B(u3_N23), .S(n4918), .Z(n8335) );
  MUX2_X2 U7283 ( .A(u3_N79), .B(u3_N22), .S(n4918), .Z(n8336) );
  MUX2_X2 U7284 ( .A(u3_N78), .B(u3_N21), .S(n4918), .Z(n8337) );
  MUX2_X2 U7285 ( .A(u3_N77), .B(u3_N20), .S(n4918), .Z(n8338) );
  MUX2_X2 U7286 ( .A(u3_N76), .B(u3_N19), .S(n4918), .Z(n8339) );
  MUX2_X2 U7287 ( .A(u3_N75), .B(u3_N18), .S(n4918), .Z(n8340) );
  MUX2_X2 U7288 ( .A(u3_N74), .B(u3_N17), .S(n4918), .Z(n8341) );
  MUX2_X2 U7289 ( .A(u3_N73), .B(u3_N16), .S(n4918), .Z(n8342) );
  MUX2_X2 U7290 ( .A(u3_N72), .B(u3_N15), .S(n4918), .Z(n8343) );
  MUX2_X2 U7291 ( .A(u3_N71), .B(u3_N14), .S(n4918), .Z(n8344) );
  MUX2_X2 U7292 ( .A(u3_N70), .B(u3_N13), .S(n4287), .Z(n8345) );
  MUX2_X2 U7293 ( .A(u3_N69), .B(u3_N12), .S(n4287), .Z(n8346) );
  MUX2_X2 U7294 ( .A(u3_N68), .B(u3_N11), .S(n4287), .Z(n8347) );
  MUX2_X2 U7295 ( .A(u3_N67), .B(u3_N10), .S(n4287), .Z(n8348) );
  MUX2_X2 U7296 ( .A(u3_N66), .B(u3_N9), .S(n4287), .Z(n8349) );
  MUX2_X2 U7297 ( .A(u3_N65), .B(u3_N8), .S(n4287), .Z(n8350) );
  MUX2_X2 U7298 ( .A(u3_N64), .B(u3_N7), .S(n4287), .Z(n8351) );
  MUX2_X2 U7299 ( .A(u3_N63), .B(u3_N6), .S(n4287), .Z(n8352) );
  MUX2_X2 U7300 ( .A(u3_N62), .B(u3_N5), .S(n4287), .Z(n8353) );
  MUX2_X2 U7301 ( .A(u3_N61), .B(u3_N4), .S(n4287), .Z(n8354) );
  MUX2_X2 U7302 ( .A(u3_N60), .B(u3_N3), .S(n4918), .Z(n8355) );
  MUX2_X2 U7303 ( .A(n6999), .B(n4297), .S(n4891), .Z(n6915) );
  INV_X4 U7304 ( .A(n6915), .ZN(u1_adj_op_51_) );
  INV_X4 U7305 ( .A(u6_N50), .ZN(n7002) );
  MUX2_X2 U7306 ( .A(n7002), .B(n4291), .S(n4891), .Z(n6914) );
  INV_X4 U7307 ( .A(n6914), .ZN(n8478) );
  INV_X4 U7308 ( .A(u6_N49), .ZN(n7005) );
  MUX2_X2 U7309 ( .A(n7005), .B(n4301), .S(n4891), .Z(n6955) );
  INV_X4 U7310 ( .A(n6955), .ZN(n8480) );
  MUX2_X2 U7311 ( .A(n7008), .B(n4303), .S(n4891), .Z(n6911) );
  INV_X4 U7312 ( .A(n6911), .ZN(n8481) );
  MUX2_X2 U7313 ( .A(n7011), .B(n4302), .S(n4891), .Z(n6910) );
  INV_X4 U7314 ( .A(n6910), .ZN(n8482) );
  MUX2_X2 U7315 ( .A(n7014), .B(n4300), .S(n4891), .Z(n6909) );
  INV_X4 U7316 ( .A(n6909), .ZN(n8483) );
  MUX2_X2 U7317 ( .A(n7017), .B(n4290), .S(n4891), .Z(n6953) );
  INV_X4 U7318 ( .A(n6953), .ZN(n8484) );
  MUX2_X2 U7319 ( .A(n7020), .B(n6451), .S(n4890), .Z(n6906) );
  INV_X4 U7320 ( .A(n6906), .ZN(u1_adj_op_44_) );
  MUX2_X2 U7321 ( .A(n7023), .B(n4296), .S(n4887), .Z(n6904) );
  INV_X4 U7322 ( .A(n6904), .ZN(n8485) );
  MUX2_X2 U7323 ( .A(n7026), .B(n4436), .S(n4890), .Z(n6981) );
  INV_X4 U7324 ( .A(n6981), .ZN(u1_adj_op_42_) );
  MUX2_X2 U7325 ( .A(n7029), .B(n4313), .S(n4890), .Z(n6902) );
  INV_X4 U7326 ( .A(n6902), .ZN(n8486) );
  MUX2_X2 U7327 ( .A(n7032), .B(n4344), .S(n4890), .Z(n6900) );
  INV_X4 U7328 ( .A(n6900), .ZN(n8487) );
  MUX2_X2 U7329 ( .A(n7035), .B(n4439), .S(n4890), .Z(n6897) );
  INV_X4 U7330 ( .A(n6897), .ZN(n8488) );
  MUX2_X2 U7331 ( .A(n7038), .B(n4335), .S(n4890), .Z(n6898) );
  INV_X4 U7332 ( .A(n6898), .ZN(u1_adj_op_38_) );
  MUX2_X2 U7333 ( .A(n7041), .B(n4310), .S(n4890), .Z(n6896) );
  INV_X4 U7334 ( .A(n6896), .ZN(u1_adj_op_37_) );
  MUX2_X2 U7335 ( .A(n7044), .B(n4340), .S(n4890), .Z(n6893) );
  INV_X4 U7336 ( .A(n6893), .ZN(u1_adj_op_36_) );
  MUX2_X2 U7337 ( .A(n4416), .B(n4311), .S(n4890), .Z(n6891) );
  INV_X4 U7338 ( .A(n6891), .ZN(n8489) );
  MUX2_X2 U7339 ( .A(n7049), .B(n4314), .S(n4890), .Z(n6892) );
  INV_X4 U7340 ( .A(n6892), .ZN(n8490) );
  MUX2_X2 U7341 ( .A(n7052), .B(n4338), .S(n4890), .Z(n6888) );
  INV_X4 U7342 ( .A(n6888), .ZN(n8491) );
  INV_X4 U7343 ( .A(u6_N32), .ZN(n7055) );
  MUX2_X2 U7344 ( .A(n7055), .B(n4342), .S(n4889), .Z(n6887) );
  INV_X4 U7345 ( .A(n6887), .ZN(u1_adj_op_32_) );
  MUX2_X2 U7346 ( .A(n7058), .B(n4423), .S(n4889), .Z(n6885) );
  INV_X4 U7347 ( .A(n6885), .ZN(n8492) );
  MUX2_X2 U7348 ( .A(n7061), .B(n4419), .S(n4889), .Z(n6986) );
  INV_X4 U7349 ( .A(n6986), .ZN(n8493) );
  MUX2_X2 U7350 ( .A(n7064), .B(n4431), .S(n4889), .Z(n6883) );
  INV_X4 U7351 ( .A(n6883), .ZN(n8495) );
  MUX2_X2 U7352 ( .A(n7067), .B(n4418), .S(n4889), .Z(n6880) );
  INV_X4 U7353 ( .A(n6880), .ZN(u1_adj_op_28_) );
  MUX2_X2 U7354 ( .A(n7070), .B(n4426), .S(n4889), .Z(n6879) );
  INV_X4 U7355 ( .A(n6879), .ZN(u1_adj_op_27_) );
  INV_X4 U7356 ( .A(u6_N26), .ZN(n7073) );
  MUX2_X2 U7357 ( .A(n7073), .B(n4422), .S(n4889), .Z(n6877) );
  INV_X4 U7358 ( .A(n6877), .ZN(n8496) );
  INV_X4 U7359 ( .A(u6_N25), .ZN(n7076) );
  MUX2_X2 U7360 ( .A(n7076), .B(n4421), .S(n4889), .Z(n6875) );
  INV_X4 U7361 ( .A(n6875), .ZN(n8497) );
  MUX2_X2 U7362 ( .A(u6_N24), .B(fracta_mul[24]), .S(n4880), .Z(n8498) );
  MUX2_X2 U7363 ( .A(u6_N23), .B(fracta_mul[23]), .S(n4889), .Z(n8499) );
  INV_X4 U7364 ( .A(u6_N22), .ZN(n7085) );
  MUX2_X2 U7365 ( .A(n7085), .B(n4289), .S(n4889), .Z(n6857) );
  INV_X4 U7366 ( .A(n6857), .ZN(u1_adj_op_22_) );
  INV_X4 U7367 ( .A(u6_N21), .ZN(n7088) );
  MUX2_X2 U7368 ( .A(n7088), .B(n4437), .S(n4889), .Z(n6858) );
  INV_X4 U7369 ( .A(n6858), .ZN(u1_adj_op_21_) );
  INV_X4 U7370 ( .A(u6_N20), .ZN(n7091) );
  MUX2_X2 U7371 ( .A(n7091), .B(n4299), .S(n4888), .Z(n6767) );
  INV_X4 U7372 ( .A(n6767), .ZN(u1_adj_op_20_) );
  MUX2_X2 U7373 ( .A(u6_N19), .B(fracta_mul[19]), .S(n4888), .Z(n8501) );
  MUX2_X2 U7374 ( .A(u6_N18), .B(fracta_mul[18]), .S(n4888), .Z(n8502) );
  MUX2_X2 U7375 ( .A(n4454), .B(n4341), .S(n4888), .Z(n6768) );
  INV_X4 U7376 ( .A(n6768), .ZN(u1_adj_op_17_) );
  MUX2_X2 U7377 ( .A(n4455), .B(n4347), .S(n4888), .Z(n6843) );
  INV_X4 U7378 ( .A(n6843), .ZN(u1_adj_op_16_) );
  MUX2_X2 U7379 ( .A(n4453), .B(n4339), .S(n4888), .Z(n6844) );
  INV_X4 U7380 ( .A(n6844), .ZN(u1_adj_op_15_) );
  MUX2_X2 U7381 ( .A(u6_N14), .B(fracta_mul[14]), .S(n4888), .Z(n8503) );
  MUX2_X2 U7382 ( .A(u6_N13), .B(fracta_mul[13]), .S(n4888), .Z(n8504) );
  MUX2_X2 U7383 ( .A(u6_N12), .B(fracta_mul[12]), .S(n4888), .Z(n8505) );
  MUX2_X2 U7384 ( .A(n4452), .B(n4312), .S(n4888), .Z(n6769) );
  INV_X4 U7385 ( .A(n6769), .ZN(u1_adj_op_11_) );
  MUX2_X2 U7386 ( .A(n4451), .B(n4337), .S(n4888), .Z(n6770) );
  INV_X4 U7387 ( .A(n6770), .ZN(u1_adj_op_10_) );
  MUX2_X2 U7388 ( .A(u6_N9), .B(fracta_mul[9]), .S(n4887), .Z(n8473) );
  MUX2_X2 U7389 ( .A(u6_N8), .B(fracta_mul[8]), .S(n4887), .Z(n8474) );
  MUX2_X2 U7390 ( .A(u6_N7), .B(fracta_mul[7]), .S(n4887), .Z(n8475) );
  MUX2_X2 U7391 ( .A(u6_N6), .B(fracta_mul[6]), .S(n4887), .Z(n8476) );
  MUX2_X2 U7392 ( .A(n4460), .B(n4343), .S(n4887), .Z(n6855) );
  INV_X4 U7393 ( .A(n6855), .ZN(n8477) );
  MUX2_X2 U7394 ( .A(n4459), .B(n4348), .S(n4887), .Z(n6856) );
  INV_X4 U7395 ( .A(n6856), .ZN(n8479) );
  MUX2_X2 U7396 ( .A(n4458), .B(n6833), .S(n4887), .Z(n6846) );
  INV_X4 U7397 ( .A(n6846), .ZN(u1_adj_op_3_) );
  MUX2_X2 U7398 ( .A(u6_N2), .B(fracta_mul[2]), .S(n4887), .Z(n8494) );
  MUX2_X2 U7399 ( .A(u6_N1), .B(n4799), .S(n4887), .Z(n8500) );
  MUX2_X2 U7400 ( .A(n4351), .B(n6839), .S(n4887), .Z(n6847) );
  INV_X4 U7401 ( .A(n6847), .ZN(u1_adj_op_0_) );
  MUX2_X2 U7402 ( .A(opb_r[62]), .B(n4853), .S(n4882), .Z(u1_exp_small[10]) );
  MUX2_X2 U7403 ( .A(opb_r[61]), .B(opa_r[61]), .S(n4883), .Z(n8471) );
  MUX2_X2 U7404 ( .A(n4823), .B(opa_r[60]), .S(n4884), .Z(n8472) );
  MUX2_X2 U7405 ( .A(n4837), .B(opa_r[59]), .S(n4890), .Z(u1_exp_small[7]) );
  MUX2_X2 U7406 ( .A(n4425), .B(opa_r[58]), .S(n4888), .Z(u1_exp_small[6]) );
  MUX2_X2 U7407 ( .A(n4839), .B(opa_r[57]), .S(n4887), .Z(u1_exp_small[5]) );
  MUX2_X2 U7408 ( .A(n4836), .B(opa_r[56]), .S(n4889), .Z(u1_exp_small[4]) );
  MUX2_X2 U7409 ( .A(opb_r[55]), .B(opa_r[55]), .S(n4880), .Z(u1_exp_small[3])
         );
  MUX2_X2 U7410 ( .A(opb_r[54]), .B(opa_r[54]), .S(n4879), .Z(u1_exp_small[2])
         );
  MUX2_X2 U7411 ( .A(opb_r[53]), .B(opa_r[53]), .S(n4892), .Z(u1_exp_small[1])
         );
  MUX2_X2 U7412 ( .A(opb_r[52]), .B(opa_r[52]), .S(n4877), .Z(u1_exp_small[0])
         );
  NAND2_X2 U7413 ( .A1(n7209), .A2(n4901), .ZN(n6779) );
  INV_X4 U7414 ( .A(n6779), .ZN(n6777) );
  INV_X4 U7415 ( .A(u1_exp_diff2[5]), .ZN(n6775) );
  NOR4_X2 U7416 ( .A1(u1_exp_diff2[10]), .A2(u1_exp_diff2[9]), .A3(
        u1_exp_diff2[8]), .A4(n4403), .ZN(n6773) );
  NAND2_X2 U7417 ( .A1(u1_exp_diff2[3]), .A2(n6779), .ZN(n6778) );
  INV_X4 U7418 ( .A(n6778), .ZN(n6771) );
  NAND3_X2 U7419 ( .A1(u1_exp_diff2[5]), .A2(u1_exp_diff2[4]), .A3(n6771), 
        .ZN(n6772) );
  OAI21_X4 U7420 ( .B1(n6777), .B2(n6773), .A(n6772), .ZN(n6774) );
  INV_X4 U7421 ( .A(n6774), .ZN(n6780) );
  OAI21_X4 U7422 ( .B1(n6777), .B2(n6775), .A(n6780), .ZN(n8470) );
  INV_X4 U7423 ( .A(u1_exp_diff2[4]), .ZN(n6776) );
  OAI21_X4 U7424 ( .B1(n6777), .B2(n6776), .A(n6780), .ZN(n8469) );
  NAND2_X2 U7425 ( .A1(n6780), .A2(n6778), .ZN(n8468) );
  NAND2_X2 U7426 ( .A1(n6780), .A2(n6779), .ZN(n6781) );
  INV_X4 U7427 ( .A(n6781), .ZN(n6783) );
  NAND2_X2 U7428 ( .A1(u1_exp_diff2[2]), .A2(n6783), .ZN(n6931) );
  INV_X4 U7429 ( .A(n6931), .ZN(n8465) );
  NAND2_X2 U7430 ( .A1(u1_exp_diff2[1]), .A2(n6783), .ZN(n6782) );
  INV_X4 U7431 ( .A(n6782), .ZN(n8466) );
  NAND2_X2 U7432 ( .A1(u1_exp_diff2[0]), .A2(n6783), .ZN(n6784) );
  INV_X4 U7433 ( .A(n6784), .ZN(n8467) );
  INV_X4 U7434 ( .A(u1_adj_op_out_sft_55_), .ZN(n6997) );
  NAND2_X2 U7435 ( .A1(n6997), .A2(n4880), .ZN(n8414) );
  INV_X4 U7436 ( .A(u1_adj_op_out_sft_54_), .ZN(n7000) );
  MUX2_X2 U7437 ( .A(n4297), .B(n7000), .S(n4885), .Z(n6785) );
  INV_X4 U7438 ( .A(n6785), .ZN(n8415) );
  INV_X4 U7439 ( .A(u1_adj_op_out_sft_53_), .ZN(n7003) );
  MUX2_X2 U7440 ( .A(n4291), .B(n7003), .S(n4885), .Z(n6786) );
  INV_X4 U7441 ( .A(n6786), .ZN(n8416) );
  INV_X4 U7442 ( .A(u1_adj_op_out_sft_52_), .ZN(n7006) );
  MUX2_X2 U7443 ( .A(n4301), .B(n7006), .S(n4885), .Z(n6787) );
  INV_X4 U7444 ( .A(n6787), .ZN(n8417) );
  INV_X4 U7445 ( .A(u1_adj_op_out_sft_51_), .ZN(n7009) );
  MUX2_X2 U7446 ( .A(n4303), .B(n7009), .S(n4885), .Z(n6788) );
  INV_X4 U7447 ( .A(n6788), .ZN(n8418) );
  INV_X4 U7448 ( .A(u1_adj_op_out_sft_50_), .ZN(n7012) );
  MUX2_X2 U7449 ( .A(n4302), .B(n7012), .S(n4885), .Z(n6789) );
  INV_X4 U7450 ( .A(n6789), .ZN(n8419) );
  INV_X4 U7451 ( .A(u1_adj_op_out_sft_49_), .ZN(n7015) );
  MUX2_X2 U7452 ( .A(n4300), .B(n7015), .S(n4885), .Z(n6790) );
  INV_X4 U7453 ( .A(n6790), .ZN(n8421) );
  INV_X4 U7454 ( .A(u1_adj_op_out_sft_48_), .ZN(n7018) );
  MUX2_X2 U7455 ( .A(n4290), .B(n7018), .S(n4885), .Z(n6791) );
  INV_X4 U7456 ( .A(n6791), .ZN(n8422) );
  INV_X4 U7457 ( .A(u1_adj_op_out_sft_47_), .ZN(n7021) );
  MUX2_X2 U7458 ( .A(n6451), .B(n7021), .S(n4886), .Z(n6792) );
  INV_X4 U7459 ( .A(n6792), .ZN(n8423) );
  INV_X4 U7460 ( .A(u1_adj_op_out_sft_46_), .ZN(n7024) );
  MUX2_X2 U7461 ( .A(n4296), .B(n7024), .S(n4885), .Z(n6793) );
  INV_X4 U7462 ( .A(n6793), .ZN(n8424) );
  INV_X4 U7463 ( .A(u1_adj_op_out_sft_45_), .ZN(n7027) );
  MUX2_X2 U7464 ( .A(n4436), .B(n7027), .S(n4885), .Z(n6794) );
  INV_X4 U7465 ( .A(n6794), .ZN(n8425) );
  INV_X4 U7466 ( .A(u1_adj_op_out_sft_44_), .ZN(n7030) );
  MUX2_X2 U7467 ( .A(n4313), .B(n7030), .S(n4886), .Z(n6795) );
  INV_X4 U7468 ( .A(n6795), .ZN(n8426) );
  INV_X4 U7469 ( .A(u1_adj_op_out_sft_43_), .ZN(n7033) );
  MUX2_X2 U7470 ( .A(n4344), .B(n7033), .S(n4885), .Z(n6796) );
  INV_X4 U7471 ( .A(n6796), .ZN(n8427) );
  INV_X4 U7472 ( .A(u1_adj_op_out_sft_42_), .ZN(n7036) );
  MUX2_X2 U7473 ( .A(n4439), .B(n7036), .S(n4885), .Z(n6797) );
  INV_X4 U7474 ( .A(n6797), .ZN(n8428) );
  INV_X4 U7475 ( .A(u1_adj_op_out_sft_41_), .ZN(n7039) );
  MUX2_X2 U7476 ( .A(n4335), .B(n7039), .S(n4885), .Z(n6798) );
  INV_X4 U7477 ( .A(n6798), .ZN(n8429) );
  INV_X4 U7478 ( .A(u1_adj_op_out_sft_40_), .ZN(n7042) );
  MUX2_X2 U7479 ( .A(n4310), .B(n7042), .S(n4885), .Z(n6799) );
  INV_X4 U7480 ( .A(n6799), .ZN(n8430) );
  INV_X4 U7481 ( .A(u1_adj_op_out_sft_39_), .ZN(n7045) );
  MUX2_X2 U7482 ( .A(n4340), .B(n7045), .S(n4885), .Z(n6800) );
  INV_X4 U7483 ( .A(n6800), .ZN(n8432) );
  INV_X4 U7484 ( .A(u1_adj_op_out_sft_38_), .ZN(n7047) );
  MUX2_X2 U7485 ( .A(n4311), .B(n7047), .S(n4885), .Z(n6801) );
  INV_X4 U7486 ( .A(n6801), .ZN(n8433) );
  INV_X4 U7487 ( .A(u1_adj_op_out_sft_37_), .ZN(n7050) );
  MUX2_X2 U7488 ( .A(n4314), .B(n7050), .S(n4885), .Z(n6802) );
  INV_X4 U7489 ( .A(n6802), .ZN(n8434) );
  INV_X4 U7490 ( .A(u1_adj_op_out_sft_36_), .ZN(n7053) );
  MUX2_X2 U7491 ( .A(n4338), .B(n7053), .S(n4885), .Z(n6803) );
  INV_X4 U7492 ( .A(n6803), .ZN(n8435) );
  INV_X4 U7493 ( .A(u1_adj_op_out_sft_35_), .ZN(n7056) );
  MUX2_X2 U7494 ( .A(n4342), .B(n7056), .S(n4885), .Z(n6804) );
  INV_X4 U7495 ( .A(n6804), .ZN(n8436) );
  INV_X4 U7496 ( .A(u1_adj_op_out_sft_34_), .ZN(n7059) );
  MUX2_X2 U7497 ( .A(n4423), .B(n7059), .S(n4886), .Z(n6805) );
  INV_X4 U7498 ( .A(n6805), .ZN(n8437) );
  INV_X4 U7499 ( .A(u1_adj_op_out_sft_33_), .ZN(n7062) );
  MUX2_X2 U7500 ( .A(n4419), .B(n7062), .S(n4886), .Z(n6806) );
  INV_X4 U7501 ( .A(n6806), .ZN(n8438) );
  INV_X4 U7502 ( .A(u1_adj_op_out_sft_32_), .ZN(n7065) );
  MUX2_X2 U7503 ( .A(n4431), .B(n7065), .S(n4886), .Z(n6807) );
  INV_X4 U7504 ( .A(n6807), .ZN(n8439) );
  INV_X4 U7505 ( .A(u1_adj_op_out_sft_31_), .ZN(n7068) );
  MUX2_X2 U7506 ( .A(n4418), .B(n7068), .S(n4886), .Z(n6808) );
  INV_X4 U7507 ( .A(n6808), .ZN(n8440) );
  INV_X4 U7508 ( .A(u1_adj_op_out_sft_30_), .ZN(n7071) );
  MUX2_X2 U7509 ( .A(n4426), .B(n7071), .S(n4886), .Z(n6809) );
  INV_X4 U7510 ( .A(n6809), .ZN(n8441) );
  INV_X4 U7511 ( .A(u1_adj_op_out_sft_29_), .ZN(n7074) );
  MUX2_X2 U7512 ( .A(n4422), .B(n7074), .S(n4886), .Z(n6810) );
  INV_X4 U7513 ( .A(n6810), .ZN(n8443) );
  INV_X4 U7514 ( .A(u1_adj_op_out_sft_28_), .ZN(n7077) );
  MUX2_X2 U7515 ( .A(n4421), .B(n7077), .S(n4886), .Z(n6811) );
  INV_X4 U7516 ( .A(n6811), .ZN(n8444) );
  INV_X4 U7517 ( .A(u1_adj_op_out_sft_27_), .ZN(n7080) );
  MUX2_X2 U7518 ( .A(n4435), .B(n7080), .S(n4886), .Z(n6812) );
  INV_X4 U7519 ( .A(n6812), .ZN(n8445) );
  INV_X4 U7520 ( .A(u1_adj_op_out_sft_26_), .ZN(n7083) );
  MUX2_X2 U7521 ( .A(n4417), .B(n7083), .S(n4886), .Z(n6813) );
  INV_X4 U7522 ( .A(n6813), .ZN(n8446) );
  INV_X4 U7523 ( .A(u1_adj_op_out_sft_25_), .ZN(n7086) );
  MUX2_X2 U7524 ( .A(n4289), .B(n7086), .S(n4886), .Z(n6814) );
  INV_X4 U7525 ( .A(n6814), .ZN(n8447) );
  INV_X4 U7526 ( .A(u1_adj_op_out_sft_24_), .ZN(n7089) );
  MUX2_X2 U7527 ( .A(n4437), .B(n7089), .S(n4886), .Z(n6815) );
  INV_X4 U7528 ( .A(n6815), .ZN(n8448) );
  INV_X4 U7529 ( .A(u1_adj_op_out_sft_23_), .ZN(n7092) );
  MUX2_X2 U7530 ( .A(n4299), .B(n7092), .S(n4885), .Z(n6816) );
  INV_X4 U7531 ( .A(n6816), .ZN(n8449) );
  INV_X4 U7532 ( .A(u1_adj_op_out_sft_22_), .ZN(n7095) );
  MUX2_X2 U7533 ( .A(n4438), .B(n7095), .S(n4885), .Z(n6817) );
  INV_X4 U7534 ( .A(n6817), .ZN(n8450) );
  INV_X4 U7535 ( .A(u1_adj_op_out_sft_21_), .ZN(n7098) );
  MUX2_X2 U7536 ( .A(n4427), .B(n7098), .S(n4885), .Z(n6818) );
  INV_X4 U7537 ( .A(n6818), .ZN(n8451) );
  INV_X4 U7538 ( .A(u1_adj_op_out_sft_20_), .ZN(n7100) );
  MUX2_X2 U7539 ( .A(n4341), .B(n7100), .S(n4885), .Z(n6819) );
  INV_X4 U7540 ( .A(n6819), .ZN(n8452) );
  INV_X4 U7541 ( .A(u1_adj_op_out_sft_19_), .ZN(n7102) );
  MUX2_X2 U7542 ( .A(n4347), .B(n7102), .S(n4885), .Z(n6820) );
  INV_X4 U7543 ( .A(n6820), .ZN(n8454) );
  INV_X4 U7544 ( .A(u1_adj_op_out_sft_18_), .ZN(n7104) );
  MUX2_X2 U7545 ( .A(n4339), .B(n7104), .S(n4885), .Z(n6821) );
  INV_X4 U7546 ( .A(n6821), .ZN(n8455) );
  INV_X4 U7547 ( .A(u1_adj_op_out_sft_17_), .ZN(n7106) );
  MUX2_X2 U7548 ( .A(n4434), .B(n7106), .S(n4885), .Z(n6822) );
  INV_X4 U7549 ( .A(n6822), .ZN(n8456) );
  INV_X4 U7550 ( .A(u1_adj_op_out_sft_16_), .ZN(n7108) );
  MUX2_X2 U7551 ( .A(n4336), .B(n7108), .S(n4885), .Z(n6823) );
  INV_X4 U7552 ( .A(n6823), .ZN(n8457) );
  INV_X4 U7553 ( .A(u1_adj_op_out_sft_15_), .ZN(n7110) );
  MUX2_X2 U7554 ( .A(n4315), .B(n7110), .S(n4885), .Z(n6824) );
  INV_X4 U7555 ( .A(n6824), .ZN(n8458) );
  INV_X4 U7556 ( .A(u1_adj_op_out_sft_14_), .ZN(n7112) );
  MUX2_X2 U7557 ( .A(n4312), .B(n7112), .S(n4885), .Z(n6825) );
  INV_X4 U7558 ( .A(n6825), .ZN(n8459) );
  INV_X4 U7559 ( .A(u1_adj_op_out_sft_13_), .ZN(n7114) );
  MUX2_X2 U7560 ( .A(n4337), .B(n7114), .S(n4885), .Z(n6826) );
  INV_X4 U7561 ( .A(n6826), .ZN(n8460) );
  INV_X4 U7562 ( .A(u1_adj_op_out_sft_12_), .ZN(n7116) );
  MUX2_X2 U7563 ( .A(n4433), .B(n7116), .S(n4884), .Z(n6827) );
  INV_X4 U7564 ( .A(n6827), .ZN(n8461) );
  INV_X4 U7565 ( .A(u1_adj_op_out_sft_11_), .ZN(n7118) );
  MUX2_X2 U7566 ( .A(n4430), .B(n7118), .S(n4884), .Z(n6828) );
  INV_X4 U7567 ( .A(n6828), .ZN(n8462) );
  INV_X4 U7568 ( .A(u1_adj_op_out_sft_10_), .ZN(n7120) );
  MUX2_X2 U7569 ( .A(n4428), .B(n7120), .S(n4884), .Z(n6829) );
  INV_X4 U7570 ( .A(n6829), .ZN(n8463) );
  INV_X4 U7571 ( .A(u1_adj_op_out_sft_9_), .ZN(n7122) );
  MUX2_X2 U7572 ( .A(n4432), .B(n7122), .S(n4884), .Z(n6830) );
  INV_X4 U7573 ( .A(n6830), .ZN(n8409) );
  INV_X4 U7574 ( .A(u1_adj_op_out_sft_8_), .ZN(n7124) );
  MUX2_X2 U7575 ( .A(n4343), .B(n7124), .S(n4884), .Z(n6831) );
  INV_X4 U7576 ( .A(n6831), .ZN(n8410) );
  INV_X4 U7577 ( .A(u1_adj_op_out_sft_7_), .ZN(n7126) );
  MUX2_X2 U7578 ( .A(n4348), .B(n7126), .S(n4884), .Z(n6832) );
  INV_X4 U7579 ( .A(n6832), .ZN(n8411) );
  INV_X4 U7580 ( .A(u1_adj_op_out_sft_6_), .ZN(n7128) );
  MUX2_X2 U7581 ( .A(n6833), .B(n7128), .S(n4884), .Z(n6834) );
  INV_X4 U7582 ( .A(n6834), .ZN(n8412) );
  INV_X4 U7583 ( .A(u1_adj_op_out_sft_5_), .ZN(n7130) );
  MUX2_X2 U7584 ( .A(n6835), .B(n7130), .S(n4884), .Z(n6836) );
  INV_X4 U7585 ( .A(n6836), .ZN(n8413) );
  INV_X4 U7586 ( .A(u1_adj_op_out_sft_4_), .ZN(n7132) );
  MUX2_X2 U7587 ( .A(n6837), .B(n7132), .S(n4884), .Z(n6838) );
  INV_X4 U7588 ( .A(n6838), .ZN(n8420) );
  INV_X4 U7589 ( .A(u1_adj_op_out_sft_3_), .ZN(n7135) );
  MUX2_X2 U7590 ( .A(n6839), .B(n7135), .S(n4884), .Z(n6840) );
  INV_X4 U7591 ( .A(n6840), .ZN(n8431) );
  NAND2_X2 U7592 ( .A1(u1_adj_op_out_sft_2_), .A2(n4879), .ZN(n6841) );
  INV_X4 U7593 ( .A(n6841), .ZN(n8442) );
  NAND2_X2 U7594 ( .A1(u1_adj_op_out_sft_1_), .A2(n4881), .ZN(n6842) );
  INV_X4 U7595 ( .A(n6842), .ZN(n8453) );
  NAND2_X2 U7596 ( .A1(n6844), .A2(n6843), .ZN(n6845) );
  NOR3_X4 U7597 ( .A1(n6845), .A2(u1_adj_op_20_), .A3(u1_adj_op_17_), .ZN(
        n6873) );
  NAND2_X2 U7598 ( .A1(n6847), .A2(n6846), .ZN(n6848) );
  NOR3_X4 U7599 ( .A1(n6848), .A2(u1_adj_op_11_), .A3(u1_adj_op_10_), .ZN(
        n6872) );
  MUX2_X2 U7600 ( .A(n6850), .B(n6849), .S(n4884), .Z(n6854) );
  MUX2_X2 U7601 ( .A(n6852), .B(n6851), .S(n4883), .Z(n6853) );
  NAND4_X2 U7602 ( .A1(n6856), .A2(n6855), .A3(n6854), .A4(n6853), .ZN(n6870)
         );
  NAND2_X2 U7603 ( .A1(n6858), .A2(n6857), .ZN(n6869) );
  NOR3_X4 U7604 ( .A1(u6_N14), .A2(u6_N12), .A3(u6_N13), .ZN(n6861) );
  NOR2_X4 U7605 ( .A1(fracta_mul[12]), .A2(n6859), .ZN(n6860) );
  MUX2_X2 U7606 ( .A(n6861), .B(n6860), .S(n4883), .Z(n6867) );
  NOR4_X2 U7607 ( .A1(u6_N8), .A2(u6_N9), .A3(u6_N6), .A4(u6_N7), .ZN(n6865)
         );
  INV_X4 U7608 ( .A(n6862), .ZN(n6863) );
  NOR2_X4 U7609 ( .A1(n6863), .A2(n4469), .ZN(n6864) );
  MUX2_X2 U7610 ( .A(n6865), .B(n6864), .S(n4883), .Z(n6866) );
  NAND2_X2 U7611 ( .A1(n6867), .A2(n6866), .ZN(n6868) );
  NOR3_X4 U7612 ( .A1(n6870), .A2(n6869), .A3(n6868), .ZN(n6871) );
  NAND3_X4 U7613 ( .A1(n6873), .A2(n6872), .A3(n6871), .ZN(n6874) );
  INV_X4 U7614 ( .A(n6874), .ZN(n6934) );
  NAND2_X2 U7615 ( .A1(n6934), .A2(n6875), .ZN(n6876) );
  INV_X4 U7616 ( .A(n6876), .ZN(n6954) );
  NAND2_X2 U7617 ( .A1(n6954), .A2(n6877), .ZN(n6878) );
  INV_X4 U7618 ( .A(n6878), .ZN(n6984) );
  NAND2_X2 U7619 ( .A1(n6984), .A2(n6879), .ZN(n6970) );
  INV_X4 U7620 ( .A(n6970), .ZN(n6881) );
  NAND2_X2 U7621 ( .A1(n6881), .A2(n6880), .ZN(n6882) );
  INV_X4 U7622 ( .A(n6882), .ZN(n6930) );
  NAND2_X2 U7623 ( .A1(n6930), .A2(n6883), .ZN(n6884) );
  INV_X4 U7624 ( .A(n6884), .ZN(n6946) );
  INV_X4 U7625 ( .A(n6886), .ZN(n6966) );
  NAND2_X2 U7626 ( .A1(n6966), .A2(n6887), .ZN(n6926) );
  INV_X4 U7627 ( .A(n6926), .ZN(n6889) );
  NAND2_X2 U7628 ( .A1(n6889), .A2(n6888), .ZN(n6890) );
  INV_X4 U7629 ( .A(n6890), .ZN(n6945) );
  INV_X4 U7630 ( .A(n6967), .ZN(n6894) );
  NAND2_X2 U7631 ( .A1(n6894), .A2(n6893), .ZN(n6895) );
  INV_X4 U7632 ( .A(n6895), .ZN(n6933) );
  NAND2_X2 U7633 ( .A1(n6933), .A2(n6896), .ZN(n6943) );
  INV_X4 U7634 ( .A(n6943), .ZN(n6899) );
  INV_X4 U7635 ( .A(n6972), .ZN(n6901) );
  NAND2_X2 U7636 ( .A1(n6901), .A2(n6900), .ZN(n6927) );
  INV_X4 U7637 ( .A(n6927), .ZN(n6903) );
  NAND2_X2 U7638 ( .A1(n6903), .A2(n6902), .ZN(n6942) );
  INV_X4 U7639 ( .A(n6942), .ZN(n6905) );
  INV_X4 U7640 ( .A(n6963), .ZN(n6907) );
  NAND2_X2 U7641 ( .A1(n6907), .A2(n6906), .ZN(n6908) );
  INV_X4 U7642 ( .A(n6908), .ZN(n6923) );
  NAND2_X2 U7643 ( .A1(n4407), .A2(n6910), .ZN(n6968) );
  INV_X4 U7644 ( .A(n6968), .ZN(n6912) );
  NAND2_X2 U7645 ( .A1(n6912), .A2(n6911), .ZN(n6913) );
  INV_X4 U7646 ( .A(n6913), .ZN(n6922) );
  NAND2_X2 U7647 ( .A1(n4286), .A2(n6916), .ZN(n6917) );
  NAND2_X2 U7648 ( .A1(n6917), .A2(n8468), .ZN(n6919) );
  INV_X4 U7649 ( .A(n8470), .ZN(n6918) );
  INV_X4 U7650 ( .A(n8469), .ZN(n6928) );
  INV_X4 U7651 ( .A(n8468), .ZN(n6920) );
  NAND2_X2 U7652 ( .A1(n8470), .A2(n6920), .ZN(n6921) );
  INV_X4 U7653 ( .A(n6921), .ZN(n6929) );
  NAND3_X4 U7654 ( .A1(n6929), .A2(n8469), .A3(n6931), .ZN(n6979) );
  NAND3_X4 U7655 ( .A1(n8465), .A2(n6929), .A3(n8469), .ZN(n6982) );
  OAI22_X2 U7656 ( .A1(n6923), .A2(n6979), .B1(n6922), .B2(n6982), .ZN(n6952)
         );
  NAND3_X2 U7657 ( .A1(n8470), .A2(n6928), .A3(n8468), .ZN(n6925) );
  INV_X4 U7658 ( .A(n6925), .ZN(n6932) );
  NAND2_X2 U7659 ( .A1(n6932), .A2(n8465), .ZN(n6980) );
  INV_X4 U7660 ( .A(n6980), .ZN(n6964) );
  NAND3_X4 U7661 ( .A1(n8465), .A2(n6928), .A3(n6929), .ZN(n6944) );
  INV_X4 U7662 ( .A(n6944), .ZN(n6978) );
  AOI22_X2 U7663 ( .A1(n6964), .A2(n6927), .B1(n6978), .B2(n6926), .ZN(n6939)
         );
  NAND3_X4 U7664 ( .A1(n6929), .A2(n6928), .A3(n6931), .ZN(n6985) );
  NAND2_X2 U7665 ( .A1(n6932), .A2(n6931), .ZN(n6941) );
  NAND3_X4 U7666 ( .A1(n8469), .A2(n8468), .A3(n8465), .ZN(n6983) );
  NOR3_X4 U7667 ( .A1(n6937), .A2(n6936), .A3(n6935), .ZN(n6938) );
  NAND3_X2 U7668 ( .A1(n6940), .A2(n6939), .A3(n6938), .ZN(n6962) );
  INV_X4 U7669 ( .A(n6941), .ZN(n6977) );
  AOI22_X2 U7670 ( .A1(n6977), .A2(n6943), .B1(n6964), .B2(n6942), .ZN(n6950)
         );
  NOR2_X4 U7671 ( .A1(n6945), .A2(n6944), .ZN(n6948) );
  NOR2_X4 U7672 ( .A1(n6946), .A2(n6985), .ZN(n6947) );
  NOR2_X4 U7673 ( .A1(n6948), .A2(n6947), .ZN(n6949) );
  NAND2_X2 U7674 ( .A1(n6950), .A2(n6949), .ZN(n6951) );
  INV_X4 U7675 ( .A(n6951), .ZN(n6993) );
  INV_X4 U7676 ( .A(n6952), .ZN(n6960) );
  NOR2_X4 U7677 ( .A1(n6954), .A2(n6983), .ZN(n6957) );
  NOR2_X4 U7678 ( .A1(n6955), .A2(n6982), .ZN(n6956) );
  NOR3_X4 U7679 ( .A1(n6958), .A2(n6957), .A3(n6956), .ZN(n6959) );
  NAND3_X2 U7680 ( .A1(n6993), .A2(n6960), .A3(n6959), .ZN(n6961) );
  MUX2_X2 U7681 ( .A(n6962), .B(n6961), .S(n8467), .Z(n6995) );
  NAND2_X2 U7682 ( .A1(n6964), .A2(n6963), .ZN(n6965) );
  OAI221_X2 U7683 ( .B1(n6966), .B2(n6985), .C1(n4286), .C2(n6982), .A(n6965), 
        .ZN(n6976) );
  INV_X4 U7684 ( .A(n6979), .ZN(n6969) );
  AOI22_X2 U7685 ( .A1(n6969), .A2(n6968), .B1(n6978), .B2(n6967), .ZN(n6974)
         );
  INV_X4 U7686 ( .A(n6983), .ZN(n6971) );
  AOI22_X2 U7687 ( .A1(n6977), .A2(n6972), .B1(n6971), .B2(n6970), .ZN(n6973)
         );
  NAND2_X2 U7688 ( .A1(n6974), .A2(n6973), .ZN(n6975) );
  OAI21_X2 U7689 ( .B1(n6976), .B2(n6975), .A(n8467), .ZN(n6992) );
  AOI22_X2 U7690 ( .A1(n6978), .A2(n8490), .B1(n6977), .B2(u1_adj_op_38_), 
        .ZN(n6991) );
  OAI22_X2 U7691 ( .A1(n6981), .A2(n6980), .B1(n4407), .B2(n6979), .ZN(n6989)
         );
  OAI22_X2 U7692 ( .A1(n6986), .A2(n6985), .B1(n6984), .B2(n6983), .ZN(n6987)
         );
  NOR3_X2 U7693 ( .A1(n6989), .A2(n6988), .A3(n6987), .ZN(n6990) );
  NAND4_X2 U7694 ( .A1(n6993), .A2(n6992), .A3(n6991), .A4(n6990), .ZN(n6994)
         );
  MUX2_X2 U7695 ( .A(n6995), .B(n6994), .S(n8466), .Z(n6996) );
  NOR2_X4 U7696 ( .A1(u1_adj_op_out_sft_0_), .A2(n6996), .ZN(n7137) );
  NOR2_X4 U7697 ( .A1(n7137), .A2(n7138), .ZN(n8464) );
  MUX2_X2 U7698 ( .A(n6997), .B(n7209), .S(n4883), .Z(n6998) );
  INV_X4 U7699 ( .A(n6998), .ZN(n8361) );
  MUX2_X2 U7700 ( .A(n7000), .B(n6999), .S(n4883), .Z(n7001) );
  INV_X4 U7701 ( .A(n7001), .ZN(n8362) );
  MUX2_X2 U7702 ( .A(n7003), .B(n7002), .S(n4883), .Z(n7004) );
  INV_X4 U7703 ( .A(n7004), .ZN(n8363) );
  MUX2_X2 U7704 ( .A(n7006), .B(n7005), .S(n4883), .Z(n7007) );
  INV_X4 U7705 ( .A(n7007), .ZN(n8364) );
  MUX2_X2 U7706 ( .A(n7009), .B(n7008), .S(n4883), .Z(n7010) );
  INV_X4 U7707 ( .A(n7010), .ZN(n8365) );
  MUX2_X2 U7708 ( .A(n7012), .B(n7011), .S(n4883), .Z(n7013) );
  INV_X4 U7709 ( .A(n7013), .ZN(n8366) );
  MUX2_X2 U7710 ( .A(n7015), .B(n7014), .S(n4883), .Z(n7016) );
  INV_X4 U7711 ( .A(n7016), .ZN(n8368) );
  MUX2_X2 U7712 ( .A(n7018), .B(n7017), .S(n4883), .Z(n7019) );
  INV_X4 U7713 ( .A(n7019), .ZN(n8369) );
  MUX2_X2 U7714 ( .A(n7021), .B(n7020), .S(n4882), .Z(n7022) );
  INV_X4 U7715 ( .A(n7022), .ZN(n8370) );
  MUX2_X2 U7716 ( .A(n7024), .B(n7023), .S(n4882), .Z(n7025) );
  INV_X4 U7717 ( .A(n7025), .ZN(n8371) );
  MUX2_X2 U7718 ( .A(n7027), .B(n7026), .S(n4882), .Z(n7028) );
  INV_X4 U7719 ( .A(n7028), .ZN(n8372) );
  MUX2_X2 U7720 ( .A(n7030), .B(n7029), .S(n4882), .Z(n7031) );
  INV_X4 U7721 ( .A(n7031), .ZN(n8373) );
  MUX2_X2 U7722 ( .A(n7033), .B(n7032), .S(n4882), .Z(n7034) );
  INV_X4 U7723 ( .A(n7034), .ZN(n8374) );
  MUX2_X2 U7724 ( .A(n7036), .B(n7035), .S(n4882), .Z(n7037) );
  INV_X4 U7725 ( .A(n7037), .ZN(n8375) );
  MUX2_X2 U7726 ( .A(n7039), .B(n7038), .S(n4882), .Z(n7040) );
  INV_X4 U7727 ( .A(n7040), .ZN(n8376) );
  MUX2_X2 U7728 ( .A(n7042), .B(n7041), .S(n4882), .Z(n7043) );
  INV_X4 U7729 ( .A(n7043), .ZN(n8377) );
  MUX2_X2 U7730 ( .A(n7045), .B(n7044), .S(n4882), .Z(n7046) );
  INV_X4 U7731 ( .A(n7046), .ZN(n8379) );
  MUX2_X2 U7732 ( .A(n7047), .B(n4416), .S(n4882), .Z(n7048) );
  INV_X4 U7733 ( .A(n7048), .ZN(n8380) );
  MUX2_X2 U7734 ( .A(n7050), .B(n7049), .S(n4882), .Z(n7051) );
  INV_X4 U7735 ( .A(n7051), .ZN(n8381) );
  MUX2_X2 U7736 ( .A(n7053), .B(n7052), .S(n4881), .Z(n7054) );
  INV_X4 U7737 ( .A(n7054), .ZN(n8382) );
  MUX2_X2 U7738 ( .A(n7056), .B(n7055), .S(n4881), .Z(n7057) );
  INV_X4 U7739 ( .A(n7057), .ZN(n8383) );
  MUX2_X2 U7740 ( .A(n7059), .B(n7058), .S(n4881), .Z(n7060) );
  INV_X4 U7741 ( .A(n7060), .ZN(n8384) );
  MUX2_X2 U7742 ( .A(n7062), .B(n7061), .S(n4881), .Z(n7063) );
  INV_X4 U7743 ( .A(n7063), .ZN(n8385) );
  MUX2_X2 U7744 ( .A(n7065), .B(n7064), .S(n4881), .Z(n7066) );
  INV_X4 U7745 ( .A(n7066), .ZN(n8386) );
  MUX2_X2 U7746 ( .A(n7068), .B(n7067), .S(n4881), .Z(n7069) );
  INV_X4 U7747 ( .A(n7069), .ZN(n8387) );
  MUX2_X2 U7748 ( .A(n7071), .B(n7070), .S(n4881), .Z(n7072) );
  INV_X4 U7749 ( .A(n7072), .ZN(n8388) );
  MUX2_X2 U7750 ( .A(n7074), .B(n7073), .S(n4881), .Z(n7075) );
  INV_X4 U7751 ( .A(n7075), .ZN(n8389) );
  MUX2_X2 U7752 ( .A(n7077), .B(n7076), .S(n4881), .Z(n7078) );
  INV_X4 U7753 ( .A(n7078), .ZN(n8390) );
  MUX2_X2 U7754 ( .A(n7080), .B(n7079), .S(n4881), .Z(n7081) );
  INV_X4 U7755 ( .A(n7081), .ZN(n8391) );
  INV_X4 U7756 ( .A(u6_N23), .ZN(n7082) );
  MUX2_X2 U7757 ( .A(n7083), .B(n7082), .S(n4881), .Z(n7084) );
  INV_X4 U7758 ( .A(n7084), .ZN(n8392) );
  MUX2_X2 U7759 ( .A(n7086), .B(n7085), .S(n4880), .Z(n7087) );
  INV_X4 U7760 ( .A(n7087), .ZN(n8393) );
  MUX2_X2 U7761 ( .A(n7089), .B(n7088), .S(n4880), .Z(n7090) );
  INV_X4 U7762 ( .A(n7090), .ZN(n8394) );
  MUX2_X2 U7763 ( .A(n7092), .B(n7091), .S(n4880), .Z(n7093) );
  INV_X4 U7764 ( .A(n7093), .ZN(n8395) );
  MUX2_X2 U7765 ( .A(n7095), .B(n7094), .S(n4880), .Z(n7096) );
  INV_X4 U7766 ( .A(n7096), .ZN(n8396) );
  INV_X4 U7767 ( .A(u6_N18), .ZN(n7097) );
  MUX2_X2 U7768 ( .A(n7098), .B(n7097), .S(n4880), .Z(n7099) );
  INV_X4 U7769 ( .A(n7099), .ZN(n8397) );
  MUX2_X2 U7770 ( .A(n7100), .B(n4454), .S(n4880), .Z(n7101) );
  INV_X4 U7771 ( .A(n7101), .ZN(n8398) );
  MUX2_X2 U7772 ( .A(n7102), .B(n4455), .S(n4880), .Z(n7103) );
  INV_X4 U7773 ( .A(n7103), .ZN(n8399) );
  MUX2_X2 U7774 ( .A(n7104), .B(n4453), .S(n4880), .Z(n7105) );
  INV_X4 U7775 ( .A(n7105), .ZN(n8400) );
  MUX2_X2 U7776 ( .A(n7106), .B(n4441), .S(n4880), .Z(n7107) );
  INV_X4 U7777 ( .A(n7107), .ZN(n8401) );
  MUX2_X2 U7778 ( .A(n7108), .B(n4440), .S(n4880), .Z(n7109) );
  INV_X4 U7779 ( .A(n7109), .ZN(n8402) );
  MUX2_X2 U7780 ( .A(n7110), .B(n4442), .S(n4880), .Z(n7111) );
  INV_X4 U7781 ( .A(n7111), .ZN(n8403) );
  MUX2_X2 U7782 ( .A(n7112), .B(n4452), .S(n4879), .Z(n7113) );
  INV_X4 U7783 ( .A(n7113), .ZN(n8404) );
  MUX2_X2 U7784 ( .A(n7114), .B(n4451), .S(n4879), .Z(n7115) );
  INV_X4 U7785 ( .A(n7115), .ZN(n8405) );
  MUX2_X2 U7786 ( .A(n7116), .B(n4449), .S(n4879), .Z(n7117) );
  INV_X4 U7787 ( .A(n7117), .ZN(n8406) );
  MUX2_X2 U7788 ( .A(n7118), .B(n4450), .S(n4879), .Z(n7119) );
  INV_X4 U7789 ( .A(n7119), .ZN(n8407) );
  MUX2_X2 U7790 ( .A(n7120), .B(n4448), .S(n4879), .Z(n7121) );
  INV_X4 U7791 ( .A(n7121), .ZN(n8408) );
  MUX2_X2 U7792 ( .A(n7122), .B(n4447), .S(n4879), .Z(n7123) );
  INV_X4 U7793 ( .A(n7123), .ZN(n8356) );
  MUX2_X2 U7794 ( .A(n7124), .B(n4460), .S(n4879), .Z(n7125) );
  INV_X4 U7795 ( .A(n7125), .ZN(n8357) );
  MUX2_X2 U7796 ( .A(n7126), .B(n4459), .S(n4879), .Z(n7127) );
  INV_X4 U7797 ( .A(n7127), .ZN(n8358) );
  MUX2_X2 U7798 ( .A(n7128), .B(n4458), .S(n4879), .Z(n7129) );
  INV_X4 U7799 ( .A(n7129), .ZN(n8359) );
  MUX2_X2 U7800 ( .A(n7130), .B(n4456), .S(n4879), .Z(n7131) );
  INV_X4 U7801 ( .A(n7131), .ZN(n8360) );
  MUX2_X2 U7802 ( .A(n7132), .B(n4457), .S(n4879), .Z(n7133) );
  INV_X4 U7803 ( .A(n7133), .ZN(n8367) );
  MUX2_X2 U7804 ( .A(n7135), .B(n4351), .S(n4885), .Z(n7136) );
  INV_X4 U7805 ( .A(n7136), .ZN(n8378) );
  INV_X4 U7806 ( .A(n7137), .ZN(n7139) );
  MUX2_X2 U7807 ( .A(n8414), .B(n8361), .S(n4905), .Z(u1_fracta_s[55]) );
  MUX2_X2 U7808 ( .A(n8415), .B(n8362), .S(n4905), .Z(u1_fracta_s[54]) );
  MUX2_X2 U7809 ( .A(n8416), .B(n8363), .S(n4905), .Z(u1_fracta_s[53]) );
  MUX2_X2 U7810 ( .A(n8417), .B(n8364), .S(n4905), .Z(u1_fracta_s[52]) );
  MUX2_X2 U7811 ( .A(n8418), .B(n8365), .S(n4905), .Z(u1_fracta_s[51]) );
  MUX2_X2 U7812 ( .A(n8419), .B(n8366), .S(n4905), .Z(u1_fracta_s[50]) );
  MUX2_X2 U7813 ( .A(n8421), .B(n8368), .S(n4905), .Z(u1_fracta_s[49]) );
  MUX2_X2 U7814 ( .A(n8422), .B(n8369), .S(n4905), .Z(u1_fracta_s[48]) );
  MUX2_X2 U7815 ( .A(n8423), .B(n8370), .S(n4905), .Z(u1_fracta_s[47]) );
  MUX2_X2 U7816 ( .A(n8424), .B(n8371), .S(n4905), .Z(u1_fracta_s[46]) );
  MUX2_X2 U7817 ( .A(n8425), .B(n8372), .S(n4905), .Z(u1_fracta_s[45]) );
  MUX2_X2 U7818 ( .A(n8426), .B(n8373), .S(n4905), .Z(u1_fracta_s[44]) );
  MUX2_X2 U7819 ( .A(n8427), .B(n8374), .S(n4905), .Z(u1_fracta_s[43]) );
  MUX2_X2 U7820 ( .A(n8428), .B(n8375), .S(n4905), .Z(u1_fracta_s[42]) );
  MUX2_X2 U7821 ( .A(n8429), .B(n8376), .S(n4905), .Z(u1_fracta_s[41]) );
  MUX2_X2 U7822 ( .A(n8430), .B(n8377), .S(n4905), .Z(u1_fracta_s[40]) );
  MUX2_X2 U7823 ( .A(n8432), .B(n8379), .S(n4905), .Z(u1_fracta_s[39]) );
  MUX2_X2 U7824 ( .A(n8433), .B(n8380), .S(n4905), .Z(u1_fracta_s[38]) );
  MUX2_X2 U7825 ( .A(n8434), .B(n8381), .S(n4905), .Z(u1_fracta_s[37]) );
  MUX2_X2 U7826 ( .A(n8435), .B(n8382), .S(n4905), .Z(u1_fracta_s[36]) );
  MUX2_X2 U7827 ( .A(n8436), .B(n8383), .S(n4905), .Z(u1_fracta_s[35]) );
  MUX2_X2 U7828 ( .A(n8437), .B(n8384), .S(n4905), .Z(u1_fracta_s[34]) );
  MUX2_X2 U7829 ( .A(n8438), .B(n8385), .S(n4907), .Z(u1_fracta_s[33]) );
  MUX2_X2 U7830 ( .A(n8439), .B(n8386), .S(n4907), .Z(u1_fracta_s[32]) );
  MUX2_X2 U7831 ( .A(n8440), .B(n8387), .S(n4907), .Z(u1_fracta_s[31]) );
  MUX2_X2 U7832 ( .A(n8441), .B(n8388), .S(n4907), .Z(u1_fracta_s[30]) );
  MUX2_X2 U7833 ( .A(n8443), .B(n8389), .S(n4907), .Z(u1_fracta_s[29]) );
  MUX2_X2 U7834 ( .A(n8444), .B(n8390), .S(n4907), .Z(u1_fracta_s[28]) );
  MUX2_X2 U7835 ( .A(n8445), .B(n8391), .S(n4907), .Z(u1_fracta_s[27]) );
  MUX2_X2 U7836 ( .A(n8446), .B(n8392), .S(n4907), .Z(u1_fracta_s[26]) );
  MUX2_X2 U7837 ( .A(n8447), .B(n8393), .S(n4907), .Z(u1_fracta_s[25]) );
  MUX2_X2 U7838 ( .A(n8448), .B(n8394), .S(n4907), .Z(u1_fracta_s[24]) );
  MUX2_X2 U7839 ( .A(n8449), .B(n8395), .S(n4907), .Z(u1_fracta_s[23]) );
  MUX2_X2 U7840 ( .A(n8450), .B(n8396), .S(n4908), .Z(u1_fracta_s[22]) );
  MUX2_X2 U7841 ( .A(n8451), .B(n8397), .S(n4908), .Z(u1_fracta_s[21]) );
  MUX2_X2 U7842 ( .A(n8452), .B(n8398), .S(n4908), .Z(u1_fracta_s[20]) );
  MUX2_X2 U7843 ( .A(n8454), .B(n8399), .S(n4908), .Z(u1_fracta_s[19]) );
  MUX2_X2 U7844 ( .A(n8455), .B(n8400), .S(n4908), .Z(u1_fracta_s[18]) );
  MUX2_X2 U7845 ( .A(n8456), .B(n8401), .S(n4908), .Z(u1_fracta_s[17]) );
  MUX2_X2 U7846 ( .A(n8457), .B(n8402), .S(n4908), .Z(u1_fracta_s[16]) );
  MUX2_X2 U7847 ( .A(n8458), .B(n8403), .S(n4908), .Z(u1_fracta_s[15]) );
  MUX2_X2 U7848 ( .A(n8459), .B(n8404), .S(n4908), .Z(u1_fracta_s[14]) );
  MUX2_X2 U7849 ( .A(n8460), .B(n8405), .S(n4908), .Z(u1_fracta_s[13]) );
  MUX2_X2 U7850 ( .A(n8461), .B(n8406), .S(n4908), .Z(u1_fracta_s[12]) );
  MUX2_X2 U7851 ( .A(n8462), .B(n8407), .S(n4909), .Z(u1_fracta_s[11]) );
  MUX2_X2 U7852 ( .A(n8463), .B(n8408), .S(n4909), .Z(u1_fracta_s[10]) );
  MUX2_X2 U7853 ( .A(n8409), .B(n8356), .S(n4909), .Z(u1_fracta_s[9]) );
  MUX2_X2 U7854 ( .A(n8410), .B(n8357), .S(n4909), .Z(u1_fracta_s[8]) );
  MUX2_X2 U7855 ( .A(n8411), .B(n8358), .S(n4909), .Z(u1_fracta_s[7]) );
  MUX2_X2 U7856 ( .A(n8412), .B(n8359), .S(n4909), .Z(u1_fracta_s[6]) );
  MUX2_X2 U7857 ( .A(n8413), .B(n8360), .S(n4909), .Z(u1_fracta_s[5]) );
  MUX2_X2 U7858 ( .A(n8420), .B(n8367), .S(n4909), .Z(u1_fracta_s[4]) );
  MUX2_X2 U7859 ( .A(n8431), .B(n8378), .S(n4909), .Z(u1_fracta_s[3]) );
  MUX2_X2 U7860 ( .A(n8442), .B(n4397), .S(n4909), .Z(u1_fracta_s[2]) );
  MUX2_X2 U7861 ( .A(n8453), .B(n4285), .S(n4909), .Z(u1_fracta_s[1]) );
  MUX2_X2 U7862 ( .A(n8464), .B(n4333), .S(n4910), .Z(u1_fracta_s[0]) );
  MUX2_X2 U7863 ( .A(n8361), .B(n8414), .S(n4910), .Z(u1_fractb_s[55]) );
  MUX2_X2 U7864 ( .A(n8362), .B(n8415), .S(n4910), .Z(u1_fractb_s[54]) );
  MUX2_X2 U7865 ( .A(n8363), .B(n8416), .S(n4910), .Z(u1_fractb_s[53]) );
  MUX2_X2 U7866 ( .A(n8364), .B(n8417), .S(n4910), .Z(u1_fractb_s[52]) );
  MUX2_X2 U7867 ( .A(n8365), .B(n8418), .S(n4910), .Z(u1_fractb_s[51]) );
  MUX2_X2 U7868 ( .A(n8366), .B(n8419), .S(n4910), .Z(u1_fractb_s[50]) );
  MUX2_X2 U7869 ( .A(n8368), .B(n8421), .S(n4910), .Z(u1_fractb_s[49]) );
  MUX2_X2 U7870 ( .A(n8369), .B(n8422), .S(n4910), .Z(u1_fractb_s[48]) );
  MUX2_X2 U7871 ( .A(n8370), .B(n8423), .S(n4910), .Z(u1_fractb_s[47]) );
  MUX2_X2 U7872 ( .A(n8371), .B(n8424), .S(n4910), .Z(u1_fractb_s[46]) );
  MUX2_X2 U7873 ( .A(n8372), .B(n8425), .S(n4911), .Z(u1_fractb_s[45]) );
  MUX2_X2 U7874 ( .A(n8373), .B(n8426), .S(n4911), .Z(u1_fractb_s[44]) );
  MUX2_X2 U7875 ( .A(n8374), .B(n8427), .S(n4911), .Z(u1_fractb_s[43]) );
  MUX2_X2 U7876 ( .A(n8375), .B(n8428), .S(n4911), .Z(u1_fractb_s[42]) );
  MUX2_X2 U7877 ( .A(n8376), .B(n8429), .S(n4911), .Z(u1_fractb_s[41]) );
  MUX2_X2 U7878 ( .A(n8377), .B(n8430), .S(n4911), .Z(u1_fractb_s[40]) );
  MUX2_X2 U7879 ( .A(n8379), .B(n8432), .S(n4911), .Z(u1_fractb_s[39]) );
  MUX2_X2 U7880 ( .A(n8380), .B(n8433), .S(n4911), .Z(u1_fractb_s[38]) );
  MUX2_X2 U7881 ( .A(n8381), .B(n8434), .S(n4911), .Z(u1_fractb_s[37]) );
  MUX2_X2 U7882 ( .A(n8382), .B(n8435), .S(n4911), .Z(u1_fractb_s[36]) );
  MUX2_X2 U7883 ( .A(n8383), .B(n8436), .S(n4911), .Z(u1_fractb_s[35]) );
  MUX2_X2 U7884 ( .A(n8384), .B(n8437), .S(n4912), .Z(u1_fractb_s[34]) );
  MUX2_X2 U7885 ( .A(n8385), .B(n8438), .S(n4912), .Z(u1_fractb_s[33]) );
  MUX2_X2 U7886 ( .A(n8386), .B(n8439), .S(n4912), .Z(u1_fractb_s[32]) );
  MUX2_X2 U7887 ( .A(n8387), .B(n8440), .S(n4912), .Z(u1_fractb_s[31]) );
  MUX2_X2 U7888 ( .A(n8388), .B(n8441), .S(n4912), .Z(u1_fractb_s[30]) );
  MUX2_X2 U7889 ( .A(n8389), .B(n8443), .S(n4912), .Z(u1_fractb_s[29]) );
  MUX2_X2 U7890 ( .A(n8390), .B(n8444), .S(n4912), .Z(u1_fractb_s[28]) );
  MUX2_X2 U7891 ( .A(n8391), .B(n8445), .S(n4912), .Z(u1_fractb_s[27]) );
  MUX2_X2 U7892 ( .A(n8392), .B(n8446), .S(n4912), .Z(u1_fractb_s[26]) );
  MUX2_X2 U7893 ( .A(n8393), .B(n8447), .S(n4912), .Z(u1_fractb_s[25]) );
  MUX2_X2 U7894 ( .A(n8394), .B(n8448), .S(n4912), .Z(u1_fractb_s[24]) );
  MUX2_X2 U7895 ( .A(n8395), .B(n8449), .S(n4913), .Z(u1_fractb_s[23]) );
  MUX2_X2 U7896 ( .A(n8396), .B(n8450), .S(n4913), .Z(u1_fractb_s[22]) );
  MUX2_X2 U7897 ( .A(n8397), .B(n8451), .S(n4913), .Z(u1_fractb_s[21]) );
  MUX2_X2 U7898 ( .A(n8398), .B(n8452), .S(n4913), .Z(u1_fractb_s[20]) );
  MUX2_X2 U7899 ( .A(n8399), .B(n8454), .S(n4913), .Z(u1_fractb_s[19]) );
  MUX2_X2 U7900 ( .A(n8400), .B(n8455), .S(n4913), .Z(u1_fractb_s[18]) );
  MUX2_X2 U7901 ( .A(n8401), .B(n8456), .S(n4913), .Z(u1_fractb_s[17]) );
  MUX2_X2 U7902 ( .A(n8402), .B(n8457), .S(n4913), .Z(u1_fractb_s[16]) );
  MUX2_X2 U7903 ( .A(n8403), .B(n8458), .S(n4913), .Z(u1_fractb_s[15]) );
  MUX2_X2 U7904 ( .A(n8404), .B(n8459), .S(n4913), .Z(u1_fractb_s[14]) );
  MUX2_X2 U7905 ( .A(n8405), .B(n8460), .S(n4913), .Z(u1_fractb_s[13]) );
  MUX2_X2 U7906 ( .A(n8406), .B(n8461), .S(n4914), .Z(u1_fractb_s[12]) );
  MUX2_X2 U7907 ( .A(n8407), .B(n8462), .S(n4914), .Z(u1_fractb_s[11]) );
  MUX2_X2 U7908 ( .A(n8408), .B(n8463), .S(n4914), .Z(u1_fractb_s[10]) );
  MUX2_X2 U7909 ( .A(n8356), .B(n8409), .S(n4914), .Z(u1_fractb_s[9]) );
  MUX2_X2 U7910 ( .A(n8357), .B(n8410), .S(n4905), .Z(u1_fractb_s[8]) );
  MUX2_X2 U7911 ( .A(n8358), .B(n8411), .S(n4914), .Z(u1_fractb_s[7]) );
  MUX2_X2 U7912 ( .A(n8359), .B(n8412), .S(n4914), .Z(u1_fractb_s[6]) );
  MUX2_X2 U7913 ( .A(n8360), .B(n8413), .S(n4913), .Z(u1_fractb_s[5]) );
  MUX2_X2 U7914 ( .A(n8367), .B(n8420), .S(n4914), .Z(u1_fractb_s[4]) );
  MUX2_X2 U7915 ( .A(n8378), .B(n8431), .S(n4914), .Z(u1_fractb_s[3]) );
  MUX2_X2 U7916 ( .A(n4397), .B(n8442), .S(n4914), .Z(u1_fractb_s[2]) );
  MUX2_X2 U7917 ( .A(n4285), .B(n8453), .S(n4914), .Z(u1_fractb_s[1]) );
  MUX2_X2 U7918 ( .A(n4333), .B(n8464), .S(n4914), .Z(u1_fractb_s[0]) );
  XOR2_X2 U7919 ( .A(opb_r[63]), .B(fpu_op_r1[0]), .Z(n7140) );
  MUX2_X2 U7920 ( .A(opa_r[63]), .B(n7140), .S(n4914), .Z(u1_sign_d) );
  NAND4_X2 U7921 ( .A1(n7144), .A2(opa_r[56]), .A3(n7143), .A4(n7142), .ZN(
        n7154) );
  INV_X4 U7922 ( .A(n7154), .ZN(n7195) );
  INV_X4 U7923 ( .A(n3074), .ZN(n8508) );
  INV_X4 U7924 ( .A(n7153), .ZN(n7197) );
  INV_X4 U7925 ( .A(u4_fract_out_51_), .ZN(n2520) );
  NAND2_X2 U7926 ( .A1(n3709), .A2(n3712), .ZN(n7156) );
  NAND2_X2 U7927 ( .A1(n3715), .A2(n3717), .ZN(n7155) );
  NOR2_X2 U7928 ( .A1(n7156), .A2(n7155), .ZN(n3897) );
  INV_X4 U7929 ( .A(net57282), .ZN(n3341) );
  INV_X4 U7930 ( .A(u4_ldz_dif_0_), .ZN(net57281) );
  MUX2_X2 U7931 ( .A(net57230), .B(n4843), .S(net66839), .Z(n2477) );
  INV_X4 U7933 ( .A(n7173), .ZN(n7160) );
  NAND2_X2 U7934 ( .A1(n7160), .A2(u4_fi_ldz_3_), .ZN(n7174) );
  INV_X4 U7935 ( .A(n7174), .ZN(n7161) );
  NAND2_X2 U7936 ( .A1(n7161), .A2(u4_fi_ldz_4_), .ZN(n7169) );
  INV_X4 U7937 ( .A(n7162), .ZN(n7178) );
  INV_X4 U7938 ( .A(n7169), .ZN(n7166) );
  NAND2_X2 U7939 ( .A1(net57252), .A2(n7165), .ZN(n2419) );
  XNOR2_X2 U7940 ( .A(n7166), .B(net57268), .ZN(n7167) );
  NAND2_X2 U7941 ( .A1(net57252), .A2(n7167), .ZN(n2417) );
  INV_X4 U7942 ( .A(net57265), .ZN(net34243) );
  NAND2_X2 U7943 ( .A1(n7174), .A2(n7168), .ZN(n7170) );
  NAND2_X2 U7944 ( .A1(n7170), .A2(n7169), .ZN(n7171) );
  AOI21_X4 U7945 ( .B1(net57252), .B2(n7171), .A(n7178), .ZN(n2415) );
  INV_X4 U7946 ( .A(net57260), .ZN(net34242) );
  NAND2_X2 U7947 ( .A1(n7173), .A2(n7172), .ZN(n7175) );
  NAND2_X2 U7948 ( .A1(n7175), .A2(n7174), .ZN(n7176) );
  INV_X4 U7949 ( .A(n7177), .ZN(n8244) );
  INV_X4 U7951 ( .A(n2408), .ZN(net45055) );
  INV_X4 U7952 ( .A(u4_exp_in_mi1_10_), .ZN(n7187) );
  OAI22_X2 U7953 ( .A1(n4843), .A2(n7179), .B1(n4505), .B2(n7191), .ZN(n7182)
         );
  INV_X4 U7954 ( .A(n7179), .ZN(n7180) );
  MUX2_X2 U7955 ( .A(n7182), .B(n7181), .S(net66875), .Z(n7185) );
  OAI221_X2 U7956 ( .B1(n7187), .B2(net57230), .C1(n2442), .C2(net45067), .A(
        n7186), .ZN(u4_shift_right[10]) );
  INV_X4 U7957 ( .A(u4_exp_in_mi1_9_), .ZN(net57229) );
  XNOR2_X2 U7958 ( .A(net66871), .B(n7188), .ZN(n7190) );
  OR3_X1 U7959 ( .A1(n4850), .A2(net66851), .A3(n4851), .ZN(n7210) );
  OR3_X1 U7960 ( .A1(n4852), .A2(net66839), .A3(n7210), .ZN(n7211) );
  NAND4_X1 U7961 ( .A1(net66851), .A2(n4851), .A3(n4852), .A4(net66839), .ZN(
        n7213) );
  NAND3_X1 U7962 ( .A1(exp_r[5]), .A2(n4850), .A3(n4848), .ZN(n7212) );
  NOR2_X1 U7963 ( .A1(n4848), .A2(net66875), .ZN(n7215) );
  OAI211_X1 U7964 ( .C1(net66851), .C2(n4851), .A(n4850), .B(exp_r[5]), .ZN(
        n7214) );
  NAND2_X1 U7965 ( .A1(n7215), .A2(n7214), .ZN(n7216) );
  NOR4_X1 U7966 ( .A1(n7216), .A2(net66863), .A3(net66871), .A4(n4846), .ZN(
        u4_N6280) );
  NOR2_X1 U7967 ( .A1(exp_r[5]), .A2(net66875), .ZN(n7220) );
  AND3_X1 U7968 ( .A1(n4852), .A2(net66839), .A3(n4851), .ZN(n7217) );
  OAI21_X1 U7969 ( .B1(n7217), .B2(net66851), .A(n4850), .ZN(n7219) );
  NOR4_X1 U7970 ( .A1(net66871), .A2(n4846), .A3(net66863), .A4(n4848), .ZN(
        n7218) );
  INV_X4 U7971 ( .A(n3068), .ZN(n8526) );
  INV_X4 U7972 ( .A(n3069), .ZN(n8527) );
  INV_X4 U7973 ( .A(n3070), .ZN(n8528) );
  INV_X4 U7974 ( .A(n3071), .ZN(n8529) );
  INV_X4 u4_sub_473_U23 ( .A(u4_fi_ldz_mi1_1_), .ZN(u4_sub_473_n13) );
  INV_X4 u4_sub_473_U22 ( .A(u4_fi_ldz_mi1_6_), .ZN(u4_sub_473_n12) );
  INV_X4 u4_sub_473_U21 ( .A(u4_fi_ldz_mi1_5_), .ZN(u4_sub_473_n11) );
  INV_X4 u4_sub_473_U20 ( .A(u4_fi_ldz_mi1_4_), .ZN(u4_sub_473_n10) );
  INV_X4 u4_sub_473_U19 ( .A(u4_fi_ldz_mi1_3_), .ZN(u4_sub_473_n9) );
  INV_X4 u4_sub_473_U18 ( .A(u4_fi_ldz_2a_2_), .ZN(u4_sub_473_n8) );
  INV_X4 u4_sub_473_U17 ( .A(net66839), .ZN(u4_sub_473_n7) );
  XNOR2_X2 u4_sub_473_U16 ( .A(u4_sub_473_n14), .B(net66839), .ZN(
        u4_exp_fix_divb[0]) );
  NAND2_X2 u4_sub_473_U15 ( .A1(net44696), .A2(u4_sub_473_n7), .ZN(
        u4_sub_473_carry_1_) );
  INV_X4 u4_sub_473_U14 ( .A(u4_sub_473_carry_9_), .ZN(u4_sub_473_n6) );
  INV_X4 u4_sub_473_U13 ( .A(net66871), .ZN(u4_sub_473_n5) );
  XNOR2_X2 u4_sub_473_U12 ( .A(net66871), .B(u4_sub_473_carry_9_), .ZN(
        u4_exp_fix_divb[9]) );
  NAND2_X2 u4_sub_473_U11 ( .A1(u4_sub_473_n5), .A2(u4_sub_473_n6), .ZN(
        u4_sub_473_carry_10_) );
  INV_X4 u4_sub_473_U10 ( .A(u4_sub_473_carry_8_), .ZN(u4_sub_473_n4) );
  INV_X4 u4_sub_473_U9 ( .A(n4846), .ZN(u4_sub_473_n3) );
  XNOR2_X2 u4_sub_473_U8 ( .A(n4846), .B(u4_sub_473_carry_8_), .ZN(
        u4_exp_fix_divb[8]) );
  NAND2_X2 u4_sub_473_U7 ( .A1(u4_sub_473_n3), .A2(u4_sub_473_n4), .ZN(
        u4_sub_473_carry_9_) );
  INV_X4 u4_sub_473_U6 ( .A(u4_sub_473_carry_7_), .ZN(u4_sub_473_n2) );
  INV_X4 u4_sub_473_U5 ( .A(net66863), .ZN(u4_sub_473_n1) );
  XNOR2_X2 u4_sub_473_U4 ( .A(net66863), .B(u4_sub_473_carry_7_), .ZN(
        u4_exp_fix_divb[7]) );
  NAND2_X2 u4_sub_473_U3 ( .A1(u4_sub_473_n1), .A2(u4_sub_473_n2), .ZN(
        u4_sub_473_carry_8_) );
  XNOR2_X2 u4_sub_473_U2 ( .A(net66875), .B(u4_sub_473_carry_10_), .ZN(
        u4_exp_fix_divb[10]) );
  INV_X2 u4_sub_473_U1 ( .A(net44696), .ZN(u4_sub_473_n14) );
  FA_X1 u4_sub_473_U2_1 ( .A(n4852), .B(u4_sub_473_n13), .CI(
        u4_sub_473_carry_1_), .CO(u4_sub_473_carry_2_), .S(u4_exp_fix_divb[1])
         );
  FA_X1 u4_sub_473_U2_2 ( .A(n4851), .B(u4_sub_473_n8), .CI(
        u4_sub_473_carry_2_), .CO(u4_sub_473_carry_3_), .S(u4_exp_fix_divb[2])
         );
  FA_X1 u4_sub_473_U2_3 ( .A(net66851), .B(u4_sub_473_n9), .CI(
        u4_sub_473_carry_3_), .CO(u4_sub_473_carry_4_), .S(u4_exp_fix_divb[3])
         );
  FA_X1 u4_sub_473_U2_4 ( .A(n4850), .B(u4_sub_473_n10), .CI(
        u4_sub_473_carry_4_), .CO(u4_sub_473_carry_5_), .S(u4_exp_fix_divb[4])
         );
  FA_X1 u4_sub_473_U2_5 ( .A(exp_r[5]), .B(u4_sub_473_n11), .CI(
        u4_sub_473_carry_5_), .CO(u4_sub_473_carry_6_), .S(u4_exp_fix_divb[5])
         );
  FA_X1 u4_sub_473_U2_6 ( .A(n4848), .B(u4_sub_473_n12), .CI(
        u4_sub_473_carry_6_), .CO(u4_sub_473_carry_7_), .S(u4_exp_fix_divb[6])
         );
  INV_X4 u4_sub_472_U23 ( .A(n7207), .ZN(u4_sub_472_n13) );
  INV_X4 u4_sub_472_U22 ( .A(u4_fi_ldz_mi22[2]), .ZN(u4_sub_472_n12) );
  INV_X4 u4_sub_472_U21 ( .A(u4_fi_ldz_mi22[3]), .ZN(u4_sub_472_n11) );
  INV_X4 u4_sub_472_U20 ( .A(u4_fi_ldz_mi22[4]), .ZN(u4_sub_472_n10) );
  INV_X4 u4_sub_472_U19 ( .A(u4_fi_ldz_mi22[5]), .ZN(u4_sub_472_n9) );
  INV_X4 u4_sub_472_U18 ( .A(u4_fi_ldz_mi22[6]), .ZN(u4_sub_472_n8) );
  INV_X4 u4_sub_472_U17 ( .A(net66839), .ZN(u4_sub_472_n7) );
  XNOR2_X2 u4_sub_472_U16 ( .A(u4_sub_472_n14), .B(net66839), .ZN(
        u4_exp_fix_diva[0]) );
  NAND2_X2 u4_sub_472_U15 ( .A1(net44696), .A2(u4_sub_472_n7), .ZN(
        u4_sub_472_carry_1_) );
  INV_X4 u4_sub_472_U14 ( .A(u4_sub_472_carry_9_), .ZN(u4_sub_472_n6) );
  INV_X4 u4_sub_472_U13 ( .A(net66871), .ZN(u4_sub_472_n5) );
  XNOR2_X2 u4_sub_472_U12 ( .A(net66871), .B(u4_sub_472_carry_9_), .ZN(
        u4_exp_fix_diva[9]) );
  NAND2_X2 u4_sub_472_U11 ( .A1(u4_sub_472_n5), .A2(u4_sub_472_n6), .ZN(
        u4_sub_472_carry_10_) );
  INV_X4 u4_sub_472_U10 ( .A(u4_sub_472_carry_8_), .ZN(u4_sub_472_n4) );
  INV_X4 u4_sub_472_U9 ( .A(n4846), .ZN(u4_sub_472_n3) );
  XNOR2_X2 u4_sub_472_U8 ( .A(n4846), .B(u4_sub_472_carry_8_), .ZN(
        u4_exp_fix_diva[8]) );
  NAND2_X2 u4_sub_472_U7 ( .A1(u4_sub_472_n3), .A2(u4_sub_472_n4), .ZN(
        u4_sub_472_carry_9_) );
  INV_X4 u4_sub_472_U6 ( .A(u4_sub_472_carry_7_), .ZN(u4_sub_472_n2) );
  INV_X4 u4_sub_472_U5 ( .A(net66863), .ZN(u4_sub_472_n1) );
  XNOR2_X2 u4_sub_472_U4 ( .A(net66863), .B(u4_sub_472_carry_7_), .ZN(
        u4_exp_fix_diva[7]) );
  NAND2_X2 u4_sub_472_U3 ( .A1(u4_sub_472_n1), .A2(u4_sub_472_n2), .ZN(
        u4_sub_472_carry_8_) );
  XNOR2_X2 u4_sub_472_U2 ( .A(net66875), .B(u4_sub_472_carry_10_), .ZN(
        u4_exp_fix_diva[10]) );
  INV_X2 u4_sub_472_U1 ( .A(net44696), .ZN(u4_sub_472_n14) );
  FA_X1 u4_sub_472_U2_1 ( .A(n4852), .B(u4_sub_472_n13), .CI(
        u4_sub_472_carry_1_), .CO(u4_sub_472_carry_2_), .S(u4_exp_fix_diva[1])
         );
  FA_X1 u4_sub_472_U2_2 ( .A(n4851), .B(u4_sub_472_n12), .CI(
        u4_sub_472_carry_2_), .CO(u4_sub_472_carry_3_), .S(u4_exp_fix_diva[2])
         );
  FA_X1 u4_sub_472_U2_3 ( .A(net66851), .B(u4_sub_472_n11), .CI(
        u4_sub_472_carry_3_), .CO(u4_sub_472_carry_4_), .S(u4_exp_fix_diva[3])
         );
  FA_X1 u4_sub_472_U2_4 ( .A(n4850), .B(u4_sub_472_n10), .CI(
        u4_sub_472_carry_4_), .CO(u4_sub_472_carry_5_), .S(u4_exp_fix_diva[4])
         );
  FA_X1 u4_sub_472_U2_5 ( .A(exp_r[5]), .B(u4_sub_472_n9), .CI(
        u4_sub_472_carry_5_), .CO(u4_sub_472_carry_6_), .S(u4_exp_fix_diva[5])
         );
  FA_X1 u4_sub_472_U2_6 ( .A(n4848), .B(u4_sub_472_n8), .CI(
        u4_sub_472_carry_6_), .CO(u4_sub_472_carry_7_), .S(u4_exp_fix_diva[6])
         );
  NOR2_X1 u4_srl_453_U1019 ( .A1(u4_shift_right[1]), .A2(u4_shift_right[7]), 
        .ZN(u4_srl_453_n910) );
  NAND2_X1 u4_srl_453_U1018 ( .A1(u4_srl_453_n910), .A2(u4_shift_right[0]), 
        .ZN(u4_srl_453_n426) );
  INV_X1 u4_srl_453_U1017 ( .A(u4_shift_right[0]), .ZN(u4_srl_453_n911) );
  NOR2_X1 u4_srl_453_U1016 ( .A1(u4_srl_453_n911), .A2(u4_srl_453_n910), .ZN(
        u4_srl_453_n428) );
  AOI22_X1 u4_srl_453_U1015 ( .A1(fract_denorm[71]), .A2(u4_srl_453_n69), .B1(
        fract_denorm[70]), .B2(u4_srl_453_n78), .ZN(u4_srl_453_n909) );
  OAI221_X1 u4_srl_453_U1014 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n142), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n141), .A(u4_srl_453_n909), .ZN(
        u4_srl_453_n536) );
  INV_X1 u4_srl_453_U1013 ( .A(u4_srl_453_n536), .ZN(u4_srl_453_n631) );
  NOR2_X1 u4_srl_453_U1012 ( .A1(u4_shift_right[3]), .A2(u4_shift_right[7]), 
        .ZN(u4_srl_453_n865) );
  INV_X1 u4_srl_453_U1011 ( .A(u4_srl_453_n865), .ZN(u4_srl_453_n760) );
  INV_X1 u4_srl_453_U1010 ( .A(u4_shift_right[2]), .ZN(u4_srl_453_n866) );
  AOI22_X1 u4_srl_453_U1009 ( .A1(fract_denorm[67]), .A2(u4_srl_453_n71), .B1(
        fract_denorm[66]), .B2(u4_srl_453_n85), .ZN(u4_srl_453_n908) );
  OAI221_X1 u4_srl_453_U1008 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n138), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n137), .A(u4_srl_453_n908), .ZN(
        u4_srl_453_n537) );
  INV_X1 u4_srl_453_U1007 ( .A(u4_srl_453_n537), .ZN(u4_srl_453_n778) );
  NOR2_X1 u4_srl_453_U1006 ( .A1(u4_srl_453_n866), .A2(u4_srl_453_n865), .ZN(
        u4_srl_453_n425) );
  AOI22_X1 u4_srl_453_U1005 ( .A1(fract_denorm[79]), .A2(u4_srl_453_n75), .B1(
        fract_denorm[78]), .B2(u4_srl_453_n85), .ZN(u4_srl_453_n907) );
  OAI221_X1 u4_srl_453_U1004 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n128), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n127), .A(u4_srl_453_n907), .ZN(
        u4_srl_453_n633) );
  AOI22_X1 u4_srl_453_U1003 ( .A1(fract_denorm[75]), .A2(u4_srl_453_n75), .B1(
        fract_denorm[74]), .B2(u4_srl_453_n84), .ZN(u4_srl_453_n906) );
  OAI221_X1 u4_srl_453_U1002 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n145), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n144), .A(u4_srl_453_n906), .ZN(
        u4_srl_453_n634) );
  AOI22_X1 u4_srl_453_U1001 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n633), .B1(
        u4_srl_453_n41), .B2(u4_srl_453_n634), .ZN(u4_srl_453_n905) );
  OAI221_X1 u4_srl_453_U1000 ( .B1(u4_srl_453_n631), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n778), .C2(u4_srl_453_n89), .A(u4_srl_453_n905), .ZN(
        u4_srl_453_n455) );
  NOR2_X1 u4_srl_453_U999 ( .A1(u4_shift_right[5]), .A2(u4_shift_right[7]), 
        .ZN(u4_srl_453_n299) );
  INV_X1 u4_srl_453_U998 ( .A(u4_srl_453_n271), .ZN(u4_srl_453_n432) );
  AOI22_X1 u4_srl_453_U997 ( .A1(fract_denorm[103]), .A2(u4_srl_453_n75), .B1(
        fract_denorm[102]), .B2(u4_srl_453_n84), .ZN(u4_srl_453_n904) );
  OAI221_X1 u4_srl_453_U996 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n109), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n111), .A(u4_srl_453_n904), .ZN(
        u4_srl_453_n531) );
  INV_X1 u4_srl_453_U995 ( .A(u4_srl_453_n277), .ZN(u4_srl_453_n412) );
  AOI22_X1 u4_srl_453_U994 ( .A1(fract_denorm[99]), .A2(u4_srl_453_n75), .B1(
        fract_denorm[98]), .B2(u4_srl_453_n84), .ZN(u4_srl_453_n903) );
  OAI221_X1 u4_srl_453_U993 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n105), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n104), .A(u4_srl_453_n903), .ZN(
        u4_srl_453_n532) );
  AOI222_X1 u4_srl_453_U992 ( .A1(u4_srl_453_n531), .A2(u4_srl_453_n25), .B1(
        u4_srl_453_n412), .B2(u4_srl_453_n40), .C1(u4_srl_453_n532), .C2(
        u4_srl_453_n87), .ZN(u4_srl_453_n217) );
  INV_X1 u4_srl_453_U991 ( .A(u4_srl_453_n217), .ZN(u4_srl_453_n378) );
  NOR2_X1 u4_srl_453_U990 ( .A1(u4_shift_right[4]), .A2(u4_srl_453_n299), .ZN(
        u4_srl_453_n368) );
  AOI22_X1 u4_srl_453_U989 ( .A1(fract_denorm[87]), .A2(u4_srl_453_n75), .B1(
        fract_denorm[86]), .B2(u4_srl_453_n84), .ZN(u4_srl_453_n902) );
  OAI221_X1 u4_srl_453_U988 ( .B1(u4_srl_453_n52), .B2(u4_srl_453_n121), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n120), .A(u4_srl_453_n902), .ZN(
        u4_srl_453_n526) );
  INV_X1 u4_srl_453_U987 ( .A(u4_srl_453_n526), .ZN(u4_srl_453_n635) );
  AOI22_X1 u4_srl_453_U986 ( .A1(fract_denorm[83]), .A2(u4_srl_453_n75), .B1(
        fract_denorm[82]), .B2(u4_srl_453_n84), .ZN(u4_srl_453_n901) );
  OAI221_X1 u4_srl_453_U985 ( .B1(u4_srl_453_n52), .B2(u4_srl_453_n131), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n130), .A(u4_srl_453_n901), .ZN(
        u4_srl_453_n527) );
  INV_X1 u4_srl_453_U984 ( .A(u4_srl_453_n527), .ZN(u4_srl_453_n780) );
  AOI22_X1 u4_srl_453_U983 ( .A1(fract_denorm[95]), .A2(u4_srl_453_n75), .B1(
        fract_denorm[94]), .B2(u4_srl_453_n84), .ZN(u4_srl_453_n900) );
  OAI221_X1 u4_srl_453_U982 ( .B1(u4_srl_453_n52), .B2(u4_srl_453_n102), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n101), .A(u4_srl_453_n900), .ZN(
        u4_srl_453_n637) );
  AOI22_X1 u4_srl_453_U981 ( .A1(fract_denorm[91]), .A2(u4_srl_453_n75), .B1(
        fract_denorm[90]), .B2(u4_srl_453_n84), .ZN(u4_srl_453_n899) );
  OAI221_X1 u4_srl_453_U980 ( .B1(u4_srl_453_n52), .B2(u4_srl_453_n124), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n123), .A(u4_srl_453_n899), .ZN(
        u4_srl_453_n638) );
  AOI22_X1 u4_srl_453_U979 ( .A1(u4_srl_453_n36), .A2(u4_srl_453_n637), .B1(
        u4_srl_453_n45), .B2(u4_srl_453_n638), .ZN(u4_srl_453_n898) );
  OAI221_X1 u4_srl_453_U978 ( .B1(u4_srl_453_n635), .B2(u4_srl_453_n30), .C1(
        u4_srl_453_n780), .C2(u4_srl_453_n89), .A(u4_srl_453_n898), .ZN(
        u4_srl_453_n379) );
  INV_X1 u4_srl_453_U977 ( .A(u4_srl_453_n275), .ZN(u4_srl_453_n433) );
  AOI222_X1 u4_srl_453_U976 ( .A1(u4_srl_453_n455), .A2(u4_srl_453_n432), .B1(
        u4_srl_453_n378), .B2(u4_srl_453_n368), .C1(u4_srl_453_n379), .C2(
        u4_srl_453_n433), .ZN(u4_srl_453_n305) );
  NOR2_X1 u4_srl_453_U975 ( .A1(u4_shift_right[6]), .A2(u4_shift_right[7]), 
        .ZN(u4_srl_453_n891) );
  NOR2_X1 u4_srl_453_U974 ( .A1(u4_srl_453_n891), .A2(u4_shift_right[8]), .ZN(
        u4_srl_453_n408) );
  AOI22_X1 u4_srl_453_U973 ( .A1(fract_denorm[55]), .A2(u4_srl_453_n75), .B1(
        fract_denorm[54]), .B2(u4_srl_453_n84), .ZN(u4_srl_453_n897) );
  OAI221_X1 u4_srl_453_U972 ( .B1(u4_srl_453_n52), .B2(u4_srl_453_n114), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n147), .A(u4_srl_453_n897), .ZN(
        u4_srl_453_n549) );
  AOI22_X1 u4_srl_453_U971 ( .A1(fract_denorm[51]), .A2(u4_srl_453_n75), .B1(
        fract_denorm[50]), .B2(u4_srl_453_n84), .ZN(u4_srl_453_n896) );
  OAI221_X1 u4_srl_453_U970 ( .B1(u4_srl_453_n52), .B2(u4_srl_453_n113), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n158), .A(u4_srl_453_n896), .ZN(
        u4_srl_453_n550) );
  AOI22_X1 u4_srl_453_U969 ( .A1(fract_denorm[63]), .A2(u4_srl_453_n75), .B1(
        fract_denorm[62]), .B2(u4_srl_453_n84), .ZN(u4_srl_453_n895) );
  OAI221_X1 u4_srl_453_U968 ( .B1(u4_srl_453_n52), .B2(u4_srl_453_n135), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n134), .A(u4_srl_453_n895), .ZN(
        u4_srl_453_n641) );
  AOI22_X1 u4_srl_453_U967 ( .A1(fract_denorm[59]), .A2(u4_srl_453_n75), .B1(
        fract_denorm[58]), .B2(u4_srl_453_n84), .ZN(u4_srl_453_n894) );
  OAI221_X1 u4_srl_453_U966 ( .B1(u4_srl_453_n52), .B2(u4_srl_453_n117), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n116), .A(u4_srl_453_n894), .ZN(
        u4_srl_453_n538) );
  AOI22_X1 u4_srl_453_U965 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n641), .B1(
        u4_srl_453_n45), .B2(u4_srl_453_n538), .ZN(u4_srl_453_n893) );
  INV_X1 u4_srl_453_U964 ( .A(u4_srl_453_n893), .ZN(u4_srl_453_n892) );
  AOI221_X1 u4_srl_453_U963 ( .B1(u4_srl_453_n549), .B2(u4_srl_453_n26), .C1(
        u4_srl_453_n550), .C2(u4_srl_453_n88), .A(u4_srl_453_n892), .ZN(
        u4_srl_453_n376) );
  NOR2_X1 u4_srl_453_U962 ( .A1(u4_srl_453_n207), .A2(u4_srl_453_n299), .ZN(
        u4_srl_453_n833) );
  INV_X1 u4_srl_453_U961 ( .A(u4_shift_right[8]), .ZN(u4_srl_453_n890) );
  NAND2_X1 u4_srl_453_U960 ( .A1(u4_srl_453_n833), .A2(u4_srl_453_n890), .ZN(
        u4_srl_453_n332) );
  AOI22_X1 u4_srl_453_U959 ( .A1(n8525), .A2(u4_srl_453_n74), .B1(n8523), .B2(
        u4_srl_453_n84), .ZN(u4_srl_453_n889) );
  OAI221_X1 u4_srl_453_U958 ( .B1(u4_srl_453_n52), .B2(u4_srl_453_n182), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n181), .A(u4_srl_453_n889), .ZN(
        u4_srl_453_n542) );
  AOI22_X1 u4_srl_453_U957 ( .A1(net33559), .A2(u4_srl_453_n74), .B1(net33552), 
        .B2(u4_srl_453_n83), .ZN(u4_srl_453_n888) );
  OAI221_X1 u4_srl_453_U956 ( .B1(u4_srl_453_n52), .B2(u4_srl_453_n178), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n177), .A(u4_srl_453_n888), .ZN(
        u4_srl_453_n543) );
  AOI22_X1 u4_srl_453_U955 ( .A1(n8515), .A2(u4_srl_453_n74), .B1(net33584), 
        .B2(u4_srl_453_n83), .ZN(u4_srl_453_n887) );
  OAI221_X1 u4_srl_453_U954 ( .B1(u4_srl_453_n52), .B2(u4_srl_453_n156), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n155), .A(u4_srl_453_n887), .ZN(
        u4_srl_453_n545) );
  AOI22_X1 u4_srl_453_U953 ( .A1(net33587), .A2(u4_srl_453_n74), .B1(net33547), 
        .B2(u4_srl_453_n83), .ZN(u4_srl_453_n886) );
  OAI221_X1 u4_srl_453_U952 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n185), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n184), .A(u4_srl_453_n886), .ZN(
        u4_srl_453_n546) );
  AOI22_X1 u4_srl_453_U951 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n545), .B1(
        u4_srl_453_n45), .B2(u4_srl_453_n546), .ZN(u4_srl_453_n885) );
  INV_X1 u4_srl_453_U950 ( .A(u4_srl_453_n885), .ZN(u4_srl_453_n884) );
  AOI221_X1 u4_srl_453_U949 ( .B1(u4_srl_453_n542), .B2(u4_srl_453_n28), .C1(
        u4_srl_453_n543), .C2(u4_srl_453_n91), .A(u4_srl_453_n884), .ZN(
        u4_srl_453_n453) );
  INV_X1 u4_srl_453_U948 ( .A(u4_srl_453_n453), .ZN(u4_srl_453_n869) );
  NAND2_X1 u4_srl_453_U947 ( .A1(u4_srl_453_n243), .A2(u4_srl_453_n299), .ZN(
        u4_srl_453_n237) );
  INV_X1 u4_srl_453_U946 ( .A(u4_srl_453_n237), .ZN(u4_srl_453_n418) );
  OAI22_X1 u4_srl_453_U945 ( .A1(u4_srl_453_n86), .A2(u4_srl_453_n93), .B1(
        u4_srl_453_n76), .B2(u4_srl_453_n94), .ZN(u4_srl_453_n883) );
  AOI221_X1 u4_srl_453_U944 ( .B1(net33648), .B2(u4_srl_453_n54), .C1(net33546), .C2(u4_srl_453_n67), .A(u4_srl_453_n883), .ZN(u4_srl_453_n871) );
  NAND2_X1 u4_srl_453_U943 ( .A1(u4_srl_453_n91), .A2(u4_srl_453_n424), .ZN(
        u4_srl_453_n298) );
  OAI22_X1 u4_srl_453_U942 ( .A1(u4_srl_453_n172), .A2(u4_srl_453_n76), .B1(
        u4_srl_453_n169), .B2(u4_srl_453_n86), .ZN(u4_srl_453_n882) );
  AOI221_X1 u4_srl_453_U941 ( .B1(u4_srl_453_n54), .B2(n8518), .C1(
        u4_srl_453_n67), .C2(net33572), .A(u4_srl_453_n882), .ZN(
        u4_srl_453_n230) );
  AOI22_X1 u4_srl_453_U940 ( .A1(net33573), .A2(u4_srl_453_n74), .B1(net33550), 
        .B2(u4_srl_453_n83), .ZN(u4_srl_453_n881) );
  OAI221_X1 u4_srl_453_U939 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n165), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n164), .A(u4_srl_453_n881), .ZN(
        u4_srl_453_n359) );
  INV_X1 u4_srl_453_U938 ( .A(u4_srl_453_n359), .ZN(u4_srl_453_n229) );
  AOI22_X1 u4_srl_453_U937 ( .A1(n8521), .A2(u4_srl_453_n74), .B1(net33563), 
        .B2(u4_srl_453_n83), .ZN(u4_srl_453_n880) );
  OAI221_X1 u4_srl_453_U936 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n175), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n174), .A(u4_srl_453_n880), .ZN(
        u4_srl_453_n544) );
  AOI22_X1 u4_srl_453_U935 ( .A1(net33566), .A2(u4_srl_453_n74), .B1(net33551), 
        .B2(u4_srl_453_n83), .ZN(u4_srl_453_n879) );
  OAI221_X1 u4_srl_453_U934 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n171), .C1(
        u4_srl_453_n170), .C2(u4_srl_453_n59), .A(u4_srl_453_n879), .ZN(
        u4_srl_453_n773) );
  AOI22_X1 u4_srl_453_U933 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n544), .B1(
        u4_srl_453_n45), .B2(u4_srl_453_n773), .ZN(u4_srl_453_n878) );
  OAI221_X1 u4_srl_453_U932 ( .B1(u4_srl_453_n230), .B2(u4_srl_453_n30), .C1(
        u4_srl_453_n229), .C2(u4_srl_453_n89), .A(u4_srl_453_n878), .ZN(
        u4_srl_453_n877) );
  INV_X1 u4_srl_453_U931 ( .A(u4_srl_453_n877), .ZN(u4_srl_453_n705) );
  AOI22_X1 u4_srl_453_U930 ( .A1(net33642), .A2(u4_srl_453_n74), .B1(n8514), 
        .B2(u4_srl_453_n83), .ZN(u4_srl_453_n876) );
  OAI221_X1 u4_srl_453_U929 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n96), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n95), .A(u4_srl_453_n876), .ZN(
        u4_srl_453_n362) );
  AOI22_X1 u4_srl_453_U928 ( .A1(n8517), .A2(u4_srl_453_n74), .B1(net33577), 
        .B2(u4_srl_453_n83), .ZN(u4_srl_453_n875) );
  OAI221_X1 u4_srl_453_U927 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n162), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n161), .A(u4_srl_453_n875), .ZN(
        u4_srl_453_n226) );
  AOI22_X1 u4_srl_453_U926 ( .A1(net33581), .A2(u4_srl_453_n74), .B1(net33549), 
        .B2(u4_srl_453_n83), .ZN(u4_srl_453_n874) );
  OAI221_X1 u4_srl_453_U925 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n191), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n99), .A(u4_srl_453_n874), .ZN(
        u4_srl_453_n227) );
  AOI222_X1 u4_srl_453_U924 ( .A1(u4_srl_453_n25), .A2(u4_srl_453_n362), .B1(
        u4_srl_453_n35), .B2(u4_srl_453_n226), .C1(u4_srl_453_n40), .C2(
        u4_srl_453_n227), .ZN(u4_srl_453_n873) );
  MUX2_X1 u4_srl_453_U923 ( .A(u4_srl_453_n705), .B(u4_srl_453_n873), .S(
        u4_srl_453_n424), .Z(u4_srl_453_n872) );
  OAI21_X1 u4_srl_453_U922 ( .B1(u4_srl_453_n871), .B2(u4_srl_453_n298), .A(
        u4_srl_453_n872), .ZN(u4_srl_453_n870) );
  AOI22_X1 u4_srl_453_U921 ( .A1(u4_srl_453_n23), .A2(u4_srl_453_n869), .B1(
        u4_srl_453_n418), .B2(u4_srl_453_n870), .ZN(u4_srl_453_n868) );
  OAI221_X1 u4_srl_453_U920 ( .B1(u4_srl_453_n305), .B2(u4_srl_453_n415), .C1(
        u4_srl_453_n376), .C2(u4_srl_453_n2), .A(u4_srl_453_n868), .ZN(
        u4_N5906) );
  AOI22_X1 u4_srl_453_U919 ( .A1(u4_srl_453_n531), .A2(u4_srl_453_n91), .B1(
        u4_srl_453_n412), .B2(u4_srl_453_n28), .ZN(u4_srl_453_n366) );
  NOR2_X1 u4_srl_453_U918 ( .A1(u4_srl_453_n366), .A2(u4_srl_453_n11), .ZN(
        u4_N6006) );
  NAND2_X1 u4_srl_453_U917 ( .A1(net63217), .A2(u4_srl_453_n67), .ZN(
        u4_srl_453_n273) );
  INV_X1 u4_srl_453_U916 ( .A(u4_srl_453_n273), .ZN(u4_srl_453_n697) );
  AOI22_X1 u4_srl_453_U915 ( .A1(fract_denorm[104]), .A2(u4_srl_453_n74), .B1(
        fract_denorm[103]), .B2(u4_srl_453_n83), .ZN(u4_srl_453_n867) );
  OAI221_X1 u4_srl_453_U914 ( .B1(u4_srl_453_n57), .B2(u4_srl_453_n110), .C1(
        u4_srl_453_n60), .C2(u4_srl_453_n109), .A(u4_srl_453_n867), .ZN(
        u4_srl_453_n501) );
  MUX2_X1 u4_srl_453_U913 ( .A(u4_srl_453_n697), .B(u4_srl_453_n501), .S(
        u4_srl_453_n866), .Z(u4_srl_453_n761) );
  NAND2_X1 u4_srl_453_U912 ( .A1(u4_srl_453_n865), .A2(u4_srl_453_n761), .ZN(
        u4_srl_453_n325) );
  NOR2_X1 u4_srl_453_U911 ( .A1(u4_srl_453_n11), .A2(u4_srl_453_n325), .ZN(
        u4_N6007) );
  AOI22_X1 u4_srl_453_U910 ( .A1(net63217), .A2(u4_srl_453_n74), .B1(
        fract_denorm[104]), .B2(u4_srl_453_n83), .ZN(u4_srl_453_n864) );
  INV_X1 u4_srl_453_U909 ( .A(u4_srl_453_n864), .ZN(u4_srl_453_n863) );
  AOI221_X1 u4_srl_453_U908 ( .B1(u4_srl_453_n58), .B2(fract_denorm[103]), 
        .C1(u4_srl_453_n67), .C2(fract_denorm[102]), .A(u4_srl_453_n863), .ZN(
        u4_srl_453_n296) );
  OR2_X1 u4_srl_453_U907 ( .A1(u4_srl_453_n11), .A2(u4_srl_453_n90), .ZN(
        u4_srl_453_n862) );
  NOR2_X1 u4_srl_453_U906 ( .A1(u4_srl_453_n296), .A2(u4_srl_453_n862), .ZN(
        u4_N6008) );
  AOI222_X1 u4_srl_453_U905 ( .A1(u4_srl_453_n58), .A2(fract_denorm[104]), 
        .B1(u4_srl_453_n78), .B2(net63217), .C1(u4_srl_453_n67), .C2(
        fract_denorm[103]), .ZN(u4_srl_453_n280) );
  NOR2_X1 u4_srl_453_U904 ( .A1(u4_srl_453_n280), .A2(u4_srl_453_n862), .ZN(
        u4_N6009) );
  NOR2_X1 u4_srl_453_U903 ( .A1(u4_srl_453_n277), .A2(u4_srl_453_n862), .ZN(
        u4_N6010) );
  NOR3_X1 u4_srl_453_U902 ( .A1(u4_srl_453_n89), .A2(u4_srl_453_n271), .A3(
        u4_srl_453_n273), .ZN(u4_srl_453_n407) );
  AND2_X1 u4_srl_453_U901 ( .A1(u4_srl_453_n243), .A2(u4_srl_453_n407), .ZN(
        u4_N6011) );
  AOI22_X1 u4_srl_453_U900 ( .A1(net33561), .A2(u4_srl_453_n73), .B1(net33562), 
        .B2(u4_srl_453_n83), .ZN(u4_srl_453_n861) );
  OAI221_X1 u4_srl_453_U899 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n179), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n176), .A(u4_srl_453_n861), .ZN(
        u4_srl_453_n606) );
  AOI22_X1 u4_srl_453_U898 ( .A1(net33564), .A2(u4_srl_453_n73), .B1(net33565), 
        .B2(u4_srl_453_n82), .ZN(u4_srl_453_n860) );
  OAI221_X1 u4_srl_453_U897 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n173), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n188), .A(u4_srl_453_n860), .ZN(
        u4_srl_453_n687) );
  AOI22_X1 u4_srl_453_U896 ( .A1(net33554), .A2(u4_srl_453_n73), .B1(n8524), 
        .B2(u4_srl_453_n82), .ZN(u4_srl_453_n859) );
  OAI221_X1 u4_srl_453_U895 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n186), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n183), .A(u4_srl_453_n859), .ZN(
        u4_srl_453_n608) );
  AOI22_X1 u4_srl_453_U894 ( .A1(n8522), .A2(u4_srl_453_n73), .B1(net33558), 
        .B2(u4_srl_453_n82), .ZN(u4_srl_453_n858) );
  OAI221_X1 u4_srl_453_U893 ( .B1(u4_srl_453_n51), .B2(u4_srl_453_n180), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n187), .A(u4_srl_453_n858), .ZN(
        u4_srl_453_n605) );
  AOI22_X1 u4_srl_453_U892 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n608), .B1(
        u4_srl_453_n45), .B2(u4_srl_453_n605), .ZN(u4_srl_453_n857) );
  INV_X1 u4_srl_453_U891 ( .A(u4_srl_453_n857), .ZN(u4_srl_453_n856) );
  AOI221_X1 u4_srl_453_U890 ( .B1(u4_srl_453_n606), .B2(u4_srl_453_n28), .C1(
        u4_srl_453_n687), .C2(u4_srl_453_n91), .A(u4_srl_453_n856), .ZN(
        u4_srl_453_n484) );
  INV_X1 u4_srl_453_U889 ( .A(u4_srl_453_n484), .ZN(u4_srl_453_n831) );
  AOI22_X1 u4_srl_453_U888 ( .A1(fract_denorm[97]), .A2(u4_srl_453_n73), .B1(
        fract_denorm[96]), .B2(u4_srl_453_n82), .ZN(u4_srl_453_n855) );
  OAI221_X1 u4_srl_453_U887 ( .B1(u4_srl_453_n51), .B2(u4_srl_453_n106), .C1(
        u4_srl_453_n64), .C2(u4_srl_453_n103), .A(u4_srl_453_n855), .ZN(
        u4_srl_453_n595) );
  AOI22_X1 u4_srl_453_U886 ( .A1(fract_denorm[93]), .A2(u4_srl_453_n73), .B1(
        fract_denorm[92]), .B2(u4_srl_453_n82), .ZN(u4_srl_453_n854) );
  OAI221_X1 u4_srl_453_U885 ( .B1(u4_srl_453_n51), .B2(u4_srl_453_n100), .C1(
        u4_srl_453_n64), .C2(u4_srl_453_n107), .A(u4_srl_453_n854), .ZN(
        u4_srl_453_n590) );
  INV_X1 u4_srl_453_U884 ( .A(u4_srl_453_n296), .ZN(u4_srl_453_n438) );
  OAI221_X1 u4_srl_453_U883 ( .B1(u4_srl_453_n51), .B2(u4_srl_453_n108), .C1(
        u4_srl_453_n64), .C2(u4_srl_453_n112), .A(u4_srl_453_n853), .ZN(
        u4_srl_453_n594) );
  AOI22_X1 u4_srl_453_U882 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n438), .B1(
        u4_srl_453_n45), .B2(u4_srl_453_n594), .ZN(u4_srl_453_n852) );
  INV_X1 u4_srl_453_U881 ( .A(u4_srl_453_n852), .ZN(u4_srl_453_n851) );
  AOI221_X1 u4_srl_453_U880 ( .B1(u4_srl_453_n595), .B2(u4_srl_453_n28), .C1(
        u4_srl_453_n590), .C2(u4_srl_453_n91), .A(u4_srl_453_n851), .ZN(
        u4_srl_453_n223) );
  AOI22_X1 u4_srl_453_U879 ( .A1(fract_denorm[81]), .A2(u4_srl_453_n73), .B1(
        fract_denorm[80]), .B2(u4_srl_453_n82), .ZN(u4_srl_453_n850) );
  OAI221_X1 u4_srl_453_U878 ( .B1(u4_srl_453_n51), .B2(u4_srl_453_n132), .C1(
        u4_srl_453_n64), .C2(u4_srl_453_n129), .A(u4_srl_453_n850), .ZN(
        u4_srl_453_n589) );
  INV_X1 u4_srl_453_U877 ( .A(u4_srl_453_n589), .ZN(u4_srl_453_n730) );
  AOI22_X1 u4_srl_453_U876 ( .A1(fract_denorm[77]), .A2(u4_srl_453_n73), .B1(
        fract_denorm[76]), .B2(u4_srl_453_n82), .ZN(u4_srl_453_n849) );
  OAI221_X1 u4_srl_453_U875 ( .B1(u4_srl_453_n51), .B2(u4_srl_453_n126), .C1(
        u4_srl_453_n64), .C2(u4_srl_453_n151), .A(u4_srl_453_n849), .ZN(
        u4_srl_453_n677) );
  INV_X1 u4_srl_453_U874 ( .A(u4_srl_453_n677), .ZN(u4_srl_453_n585) );
  AOI22_X1 u4_srl_453_U873 ( .A1(fract_denorm[89]), .A2(u4_srl_453_n73), .B1(
        fract_denorm[88]), .B2(u4_srl_453_n82), .ZN(u4_srl_453_n848) );
  OAI221_X1 u4_srl_453_U872 ( .B1(u4_srl_453_n51), .B2(u4_srl_453_n125), .C1(
        u4_srl_453_n64), .C2(u4_srl_453_n122), .A(u4_srl_453_n848), .ZN(
        u4_srl_453_n591) );
  AOI22_X1 u4_srl_453_U871 ( .A1(fract_denorm[85]), .A2(u4_srl_453_n73), .B1(
        fract_denorm[84]), .B2(u4_srl_453_n82), .ZN(u4_srl_453_n847) );
  OAI221_X1 u4_srl_453_U870 ( .B1(u4_srl_453_n51), .B2(u4_srl_453_n119), .C1(
        u4_srl_453_n64), .C2(u4_srl_453_n150), .A(u4_srl_453_n847), .ZN(
        u4_srl_453_n588) );
  AOI22_X1 u4_srl_453_U869 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n591), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n588), .ZN(u4_srl_453_n846) );
  OAI221_X1 u4_srl_453_U868 ( .B1(u4_srl_453_n730), .B2(u4_srl_453_n30), .C1(
        u4_srl_453_n585), .C2(u4_srl_453_n89), .A(u4_srl_453_n846), .ZN(
        u4_srl_453_n403) );
  INV_X1 u4_srl_453_U867 ( .A(u4_srl_453_n403), .ZN(u4_srl_453_n330) );
  OAI22_X1 u4_srl_453_U866 ( .A1(u4_srl_453_n223), .A2(u4_srl_453_n275), .B1(
        u4_srl_453_n330), .B2(u4_srl_453_n271), .ZN(u4_srl_453_n269) );
  AOI22_X1 u4_srl_453_U865 ( .A1(fract_denorm[65]), .A2(u4_srl_453_n73), .B1(
        fract_denorm[64]), .B2(u4_srl_453_n82), .ZN(u4_srl_453_n845) );
  OAI221_X1 u4_srl_453_U864 ( .B1(u4_srl_453_n51), .B2(u4_srl_453_n139), .C1(
        u4_srl_453_n64), .C2(u4_srl_453_n136), .A(u4_srl_453_n845), .ZN(
        u4_srl_453_n601) );
  AOI22_X1 u4_srl_453_U863 ( .A1(fract_denorm[61]), .A2(u4_srl_453_n72), .B1(
        fract_denorm[60]), .B2(u4_srl_453_n82), .ZN(u4_srl_453_n844) );
  OAI221_X1 u4_srl_453_U862 ( .B1(u4_srl_453_n51), .B2(u4_srl_453_n133), .C1(
        u4_srl_453_n64), .C2(u4_srl_453_n148), .A(u4_srl_453_n844), .ZN(
        u4_srl_453_n596) );
  AOI22_X1 u4_srl_453_U861 ( .A1(fract_denorm[73]), .A2(u4_srl_453_n72), .B1(
        fract_denorm[72]), .B2(u4_srl_453_n81), .ZN(u4_srl_453_n843) );
  OAI221_X1 u4_srl_453_U860 ( .B1(u4_srl_453_n51), .B2(u4_srl_453_n146), .C1(
        u4_srl_453_n64), .C2(u4_srl_453_n143), .A(u4_srl_453_n843), .ZN(
        u4_srl_453_n678) );
  AOI22_X1 u4_srl_453_U859 ( .A1(fract_denorm[69]), .A2(u4_srl_453_n72), .B1(
        fract_denorm[68]), .B2(u4_srl_453_n81), .ZN(u4_srl_453_n842) );
  OAI221_X1 u4_srl_453_U858 ( .B1(u4_srl_453_n50), .B2(u4_srl_453_n140), .C1(
        u4_srl_453_n64), .C2(u4_srl_453_n149), .A(u4_srl_453_n842), .ZN(
        u4_srl_453_n600) );
  AOI22_X1 u4_srl_453_U857 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n678), .B1(
        u4_srl_453_n45), .B2(u4_srl_453_n600), .ZN(u4_srl_453_n841) );
  INV_X1 u4_srl_453_U856 ( .A(u4_srl_453_n841), .ZN(u4_srl_453_n840) );
  AOI221_X1 u4_srl_453_U855 ( .B1(u4_srl_453_n601), .B2(u4_srl_453_n28), .C1(
        u4_srl_453_n596), .C2(u4_srl_453_n91), .A(u4_srl_453_n840), .ZN(
        u4_srl_453_n331) );
  AOI22_X1 u4_srl_453_U854 ( .A1(net33625), .A2(u4_srl_453_n72), .B1(net33583), 
        .B2(u4_srl_453_n81), .ZN(u4_srl_453_n839) );
  OAI221_X1 u4_srl_453_U853 ( .B1(u4_srl_453_n50), .B2(u4_srl_453_n159), .C1(
        u4_srl_453_n63), .C2(u4_srl_453_n157), .A(u4_srl_453_n839), .ZN(
        u4_srl_453_n612) );
  AOI22_X1 u4_srl_453_U852 ( .A1(net33585), .A2(u4_srl_453_n72), .B1(net33586), 
        .B2(u4_srl_453_n81), .ZN(u4_srl_453_n838) );
  OAI221_X1 u4_srl_453_U851 ( .B1(u4_srl_453_n50), .B2(u4_srl_453_n154), .C1(
        u4_srl_453_n63), .C2(u4_srl_453_n192), .A(u4_srl_453_n838), .ZN(
        u4_srl_453_n607) );
  AOI22_X1 u4_srl_453_U850 ( .A1(fract_denorm[57]), .A2(u4_srl_453_n72), .B1(
        fract_denorm[56]), .B2(u4_srl_453_n81), .ZN(u4_srl_453_n837) );
  OAI221_X1 u4_srl_453_U849 ( .B1(u4_srl_453_n50), .B2(u4_srl_453_n118), .C1(
        u4_srl_453_n63), .C2(u4_srl_453_n115), .A(u4_srl_453_n837), .ZN(
        u4_srl_453_n597) );
  AOI22_X1 u4_srl_453_U848 ( .A1(fract_denorm[53]), .A2(u4_srl_453_n72), .B1(
        fract_denorm[52]), .B2(u4_srl_453_n81), .ZN(u4_srl_453_n836) );
  OAI221_X1 u4_srl_453_U847 ( .B1(u4_srl_453_n50), .B2(u4_srl_453_n152), .C1(
        u4_srl_453_n63), .C2(u4_srl_453_n153), .A(u4_srl_453_n836), .ZN(
        u4_srl_453_n611) );
  AOI22_X1 u4_srl_453_U846 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n597), .B1(
        u4_srl_453_n45), .B2(u4_srl_453_n611), .ZN(u4_srl_453_n835) );
  INV_X1 u4_srl_453_U845 ( .A(u4_srl_453_n835), .ZN(u4_srl_453_n834) );
  AOI221_X1 u4_srl_453_U844 ( .B1(u4_srl_453_n612), .B2(u4_srl_453_n28), .C1(
        u4_srl_453_n607), .C2(u4_srl_453_n91), .A(u4_srl_453_n834), .ZN(
        u4_srl_453_n405) );
  OAI22_X1 u4_srl_453_U843 ( .A1(u4_srl_453_n331), .A2(u4_srl_453_n210), .B1(
        u4_srl_453_n405), .B2(u4_srl_453_n212), .ZN(u4_srl_453_n832) );
  AOI221_X1 u4_srl_453_U842 ( .B1(u4_srl_453_n204), .B2(u4_srl_453_n831), .C1(
        u4_srl_453_n269), .C2(u4_srl_453_n207), .A(u4_srl_453_n832), .ZN(
        u4_srl_453_n823) );
  NOR2_X1 u4_srl_453_U841 ( .A1(u4_srl_453_n271), .A2(u4_srl_453_n207), .ZN(
        u4_srl_453_n826) );
  AOI22_X1 u4_srl_453_U840 ( .A1(net33575), .A2(u4_srl_453_n72), .B1(n8516), 
        .B2(u4_srl_453_n81), .ZN(u4_srl_453_n830) );
  OAI221_X1 u4_srl_453_U839 ( .B1(u4_srl_453_n50), .B2(u4_srl_453_n166), .C1(
        u4_srl_453_n63), .C2(u4_srl_453_n163), .A(u4_srl_453_n830), .ZN(
        u4_srl_453_n286) );
  AOI22_X1 u4_srl_453_U838 ( .A1(net33578), .A2(u4_srl_453_n72), .B1(net33579), 
        .B2(u4_srl_453_n81), .ZN(u4_srl_453_n829) );
  OAI221_X1 u4_srl_453_U837 ( .B1(u4_srl_453_n50), .B2(u4_srl_453_n160), .C1(
        u4_srl_453_n63), .C2(u4_srl_453_n190), .A(u4_srl_453_n829), .ZN(
        u4_srl_453_n290) );
  AOI22_X1 u4_srl_453_U836 ( .A1(n8518), .A2(u4_srl_453_n72), .B1(net33572), 
        .B2(u4_srl_453_n81), .ZN(u4_srl_453_n828) );
  OAI221_X1 u4_srl_453_U835 ( .B1(u4_srl_453_n50), .B2(u4_srl_453_n167), .C1(
        u4_srl_453_n63), .C2(u4_srl_453_n189), .A(u4_srl_453_n828), .ZN(
        u4_srl_453_n285) );
  INV_X1 u4_srl_453_U834 ( .A(u4_srl_453_n285), .ZN(u4_srl_453_n685) );
  OAI22_X1 u4_srl_453_U833 ( .A1(u4_srl_453_n171), .A2(u4_srl_453_n76), .B1(
        u4_srl_453_n86), .B2(u4_srl_453_n170), .ZN(u4_srl_453_n827) );
  AOI221_X1 u4_srl_453_U832 ( .B1(n8520), .B2(u4_srl_453_n54), .C1(n8519), 
        .C2(u4_srl_453_n67), .A(u4_srl_453_n827), .ZN(u4_srl_453_n603) );
  OAI22_X1 u4_srl_453_U831 ( .A1(u4_srl_453_n685), .A2(u4_srl_453_n201), .B1(
        u4_srl_453_n603), .B2(u4_srl_453_n203), .ZN(u4_srl_453_n825) );
  AOI221_X1 u4_srl_453_U830 ( .B1(u4_srl_453_n195), .B2(u4_srl_453_n286), .C1(
        u4_srl_453_n197), .C2(u4_srl_453_n290), .A(u4_srl_453_n825), .ZN(
        u4_srl_453_n824) );
  AOI21_X1 u4_srl_453_U829 ( .B1(u4_srl_453_n823), .B2(u4_srl_453_n824), .A(
        u4_shift_right[8]), .ZN(u4_N5916) );
  AOI22_X1 u4_srl_453_U828 ( .A1(net33552), .A2(u4_srl_453_n72), .B1(net33561), 
        .B2(u4_srl_453_n81), .ZN(u4_srl_453_n822) );
  OAI221_X1 u4_srl_453_U827 ( .B1(u4_srl_453_n50), .B2(u4_srl_453_n177), .C1(
        u4_srl_453_n63), .C2(u4_srl_453_n179), .A(u4_srl_453_n822), .ZN(
        u4_srl_453_n575) );
  AOI22_X1 u4_srl_453_U826 ( .A1(net33563), .A2(u4_srl_453_n71), .B1(net33564), 
        .B2(u4_srl_453_n81), .ZN(u4_srl_453_n821) );
  OAI221_X1 u4_srl_453_U825 ( .B1(u4_srl_453_n50), .B2(u4_srl_453_n174), .C1(
        u4_srl_453_n63), .C2(u4_srl_453_n173), .A(u4_srl_453_n821), .ZN(
        u4_srl_453_n670) );
  AOI22_X1 u4_srl_453_U824 ( .A1(net33547), .A2(u4_srl_453_n71), .B1(net33554), 
        .B2(u4_srl_453_n80), .ZN(u4_srl_453_n820) );
  OAI221_X1 u4_srl_453_U823 ( .B1(u4_srl_453_n49), .B2(u4_srl_453_n184), .C1(
        u4_srl_453_n63), .C2(u4_srl_453_n186), .A(u4_srl_453_n820), .ZN(
        u4_srl_453_n577) );
  AOI22_X1 u4_srl_453_U822 ( .A1(n8523), .A2(u4_srl_453_n71), .B1(n8522), .B2(
        u4_srl_453_n80), .ZN(u4_srl_453_n819) );
  OAI221_X1 u4_srl_453_U821 ( .B1(u4_srl_453_n49), .B2(u4_srl_453_n181), .C1(
        u4_srl_453_n62), .C2(u4_srl_453_n180), .A(u4_srl_453_n819), .ZN(
        u4_srl_453_n574) );
  AOI22_X1 u4_srl_453_U820 ( .A1(u4_srl_453_n36), .A2(u4_srl_453_n577), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n574), .ZN(u4_srl_453_n818) );
  INV_X1 u4_srl_453_U819 ( .A(u4_srl_453_n818), .ZN(u4_srl_453_n817) );
  AOI221_X1 u4_srl_453_U818 ( .B1(u4_srl_453_n575), .B2(u4_srl_453_n28), .C1(
        u4_srl_453_n670), .C2(u4_srl_453_n91), .A(u4_srl_453_n817), .ZN(
        u4_srl_453_n481) );
  INV_X1 u4_srl_453_U817 ( .A(u4_srl_453_n481), .ZN(u4_srl_453_n793) );
  AOI22_X1 u4_srl_453_U816 ( .A1(fract_denorm[98]), .A2(u4_srl_453_n72), .B1(
        fract_denorm[97]), .B2(u4_srl_453_n80), .ZN(u4_srl_453_n816) );
  OAI221_X1 u4_srl_453_U815 ( .B1(u4_srl_453_n49), .B2(u4_srl_453_n104), .C1(
        u4_srl_453_n62), .C2(u4_srl_453_n106), .A(u4_srl_453_n816), .ZN(
        u4_srl_453_n564) );
  AOI22_X1 u4_srl_453_U814 ( .A1(fract_denorm[94]), .A2(u4_srl_453_n71), .B1(
        fract_denorm[93]), .B2(u4_srl_453_n80), .ZN(u4_srl_453_n815) );
  OAI221_X1 u4_srl_453_U813 ( .B1(u4_srl_453_n49), .B2(u4_srl_453_n101), .C1(
        u4_srl_453_n62), .C2(u4_srl_453_n100), .A(u4_srl_453_n815), .ZN(
        u4_srl_453_n559) );
  INV_X1 u4_srl_453_U812 ( .A(u4_srl_453_n280), .ZN(u4_srl_453_n435) );
  OAI221_X1 u4_srl_453_U811 ( .B1(u4_srl_453_n49), .B2(u4_srl_453_n111), .C1(
        u4_srl_453_n62), .C2(u4_srl_453_n108), .A(u4_srl_453_n814), .ZN(
        u4_srl_453_n563) );
  AOI22_X1 u4_srl_453_U810 ( .A1(u4_srl_453_n36), .A2(u4_srl_453_n435), .B1(
        u4_srl_453_n45), .B2(u4_srl_453_n563), .ZN(u4_srl_453_n813) );
  INV_X1 u4_srl_453_U809 ( .A(u4_srl_453_n813), .ZN(u4_srl_453_n812) );
  AOI221_X1 u4_srl_453_U808 ( .B1(u4_srl_453_n564), .B2(u4_srl_453_n28), .C1(
        u4_srl_453_n559), .C2(u4_srl_453_n88), .A(u4_srl_453_n812), .ZN(
        u4_srl_453_n222) );
  AOI22_X1 u4_srl_453_U807 ( .A1(fract_denorm[82]), .A2(u4_srl_453_n71), .B1(
        fract_denorm[81]), .B2(u4_srl_453_n80), .ZN(u4_srl_453_n811) );
  OAI221_X1 u4_srl_453_U806 ( .B1(u4_srl_453_n49), .B2(u4_srl_453_n130), .C1(
        u4_srl_453_n62), .C2(u4_srl_453_n132), .A(u4_srl_453_n811), .ZN(
        u4_srl_453_n558) );
  INV_X1 u4_srl_453_U805 ( .A(u4_srl_453_n558), .ZN(u4_srl_453_n717) );
  AOI22_X1 u4_srl_453_U804 ( .A1(fract_denorm[78]), .A2(u4_srl_453_n71), .B1(
        fract_denorm[77]), .B2(u4_srl_453_n80), .ZN(u4_srl_453_n810) );
  OAI221_X1 u4_srl_453_U803 ( .B1(u4_srl_453_n49), .B2(u4_srl_453_n127), .C1(
        u4_srl_453_n62), .C2(u4_srl_453_n126), .A(u4_srl_453_n810), .ZN(
        u4_srl_453_n660) );
  INV_X1 u4_srl_453_U802 ( .A(u4_srl_453_n660), .ZN(u4_srl_453_n554) );
  AOI22_X1 u4_srl_453_U801 ( .A1(fract_denorm[90]), .A2(u4_srl_453_n71), .B1(
        fract_denorm[89]), .B2(u4_srl_453_n80), .ZN(u4_srl_453_n809) );
  OAI221_X1 u4_srl_453_U800 ( .B1(u4_srl_453_n49), .B2(u4_srl_453_n123), .C1(
        u4_srl_453_n62), .C2(u4_srl_453_n125), .A(u4_srl_453_n809), .ZN(
        u4_srl_453_n560) );
  AOI22_X1 u4_srl_453_U799 ( .A1(fract_denorm[86]), .A2(u4_srl_453_n71), .B1(
        fract_denorm[85]), .B2(u4_srl_453_n80), .ZN(u4_srl_453_n808) );
  OAI221_X1 u4_srl_453_U798 ( .B1(u4_srl_453_n49), .B2(u4_srl_453_n120), .C1(
        u4_srl_453_n62), .C2(u4_srl_453_n119), .A(u4_srl_453_n808), .ZN(
        u4_srl_453_n557) );
  AOI22_X1 u4_srl_453_U797 ( .A1(u4_srl_453_n36), .A2(u4_srl_453_n560), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n557), .ZN(u4_srl_453_n807) );
  OAI221_X1 u4_srl_453_U796 ( .B1(u4_srl_453_n717), .B2(u4_srl_453_n30), .C1(
        u4_srl_453_n554), .C2(u4_srl_453_n89), .A(u4_srl_453_n807), .ZN(
        u4_srl_453_n398) );
  INV_X1 u4_srl_453_U795 ( .A(u4_srl_453_n398), .ZN(u4_srl_453_n328) );
  OAI22_X1 u4_srl_453_U794 ( .A1(u4_srl_453_n222), .A2(u4_srl_453_n275), .B1(
        u4_srl_453_n328), .B2(u4_srl_453_n271), .ZN(u4_srl_453_n268) );
  AOI22_X1 u4_srl_453_U793 ( .A1(fract_denorm[66]), .A2(u4_srl_453_n71), .B1(
        fract_denorm[65]), .B2(u4_srl_453_n80), .ZN(u4_srl_453_n806) );
  OAI221_X1 u4_srl_453_U792 ( .B1(u4_srl_453_n49), .B2(u4_srl_453_n137), .C1(
        u4_srl_453_n62), .C2(u4_srl_453_n139), .A(u4_srl_453_n806), .ZN(
        u4_srl_453_n570) );
  AOI22_X1 u4_srl_453_U791 ( .A1(fract_denorm[62]), .A2(u4_srl_453_n71), .B1(
        fract_denorm[61]), .B2(u4_srl_453_n80), .ZN(u4_srl_453_n805) );
  OAI221_X1 u4_srl_453_U790 ( .B1(u4_srl_453_n49), .B2(u4_srl_453_n134), .C1(
        u4_srl_453_n62), .C2(u4_srl_453_n133), .A(u4_srl_453_n805), .ZN(
        u4_srl_453_n565) );
  AOI22_X1 u4_srl_453_U789 ( .A1(fract_denorm[74]), .A2(u4_srl_453_n71), .B1(
        fract_denorm[73]), .B2(u4_srl_453_n80), .ZN(u4_srl_453_n804) );
  OAI221_X1 u4_srl_453_U788 ( .B1(u4_srl_453_n48), .B2(u4_srl_453_n144), .C1(
        u4_srl_453_n62), .C2(u4_srl_453_n146), .A(u4_srl_453_n804), .ZN(
        u4_srl_453_n661) );
  AOI22_X1 u4_srl_453_U787 ( .A1(fract_denorm[70]), .A2(u4_srl_453_n71), .B1(
        fract_denorm[69]), .B2(u4_srl_453_n85), .ZN(u4_srl_453_n803) );
  OAI221_X1 u4_srl_453_U786 ( .B1(u4_srl_453_n48), .B2(u4_srl_453_n141), .C1(
        u4_srl_453_n61), .C2(u4_srl_453_n140), .A(u4_srl_453_n803), .ZN(
        u4_srl_453_n569) );
  AOI22_X1 u4_srl_453_U785 ( .A1(u4_srl_453_n36), .A2(u4_srl_453_n661), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n569), .ZN(u4_srl_453_n802) );
  INV_X1 u4_srl_453_U784 ( .A(u4_srl_453_n802), .ZN(u4_srl_453_n801) );
  AOI221_X1 u4_srl_453_U783 ( .B1(u4_srl_453_n570), .B2(u4_srl_453_n28), .C1(
        u4_srl_453_n565), .C2(u4_srl_453_n91), .A(u4_srl_453_n801), .ZN(
        u4_srl_453_n329) );
  AOI22_X1 u4_srl_453_U782 ( .A1(fract_denorm[50]), .A2(u4_srl_453_n71), .B1(
        net33625), .B2(u4_srl_453_n85), .ZN(u4_srl_453_n800) );
  OAI221_X1 u4_srl_453_U781 ( .B1(u4_srl_453_n48), .B2(u4_srl_453_n158), .C1(
        u4_srl_453_n61), .C2(u4_srl_453_n159), .A(u4_srl_453_n800), .ZN(
        u4_srl_453_n581) );
  AOI22_X1 u4_srl_453_U780 ( .A1(net33584), .A2(u4_srl_453_n71), .B1(net33585), 
        .B2(u4_srl_453_n85), .ZN(u4_srl_453_n799) );
  OAI221_X1 u4_srl_453_U779 ( .B1(u4_srl_453_n48), .B2(u4_srl_453_n155), .C1(
        u4_srl_453_n61), .C2(u4_srl_453_n154), .A(u4_srl_453_n799), .ZN(
        u4_srl_453_n576) );
  AOI22_X1 u4_srl_453_U778 ( .A1(fract_denorm[58]), .A2(u4_srl_453_n71), .B1(
        fract_denorm[57]), .B2(u4_srl_453_n85), .ZN(u4_srl_453_n798) );
  OAI221_X1 u4_srl_453_U777 ( .B1(u4_srl_453_n48), .B2(u4_srl_453_n116), .C1(
        u4_srl_453_n61), .C2(u4_srl_453_n118), .A(u4_srl_453_n798), .ZN(
        u4_srl_453_n566) );
  AOI22_X1 u4_srl_453_U776 ( .A1(fract_denorm[54]), .A2(u4_srl_453_n71), .B1(
        fract_denorm[53]), .B2(u4_srl_453_n85), .ZN(u4_srl_453_n797) );
  OAI221_X1 u4_srl_453_U775 ( .B1(u4_srl_453_n48), .B2(u4_srl_453_n147), .C1(
        u4_srl_453_n61), .C2(u4_srl_453_n152), .A(u4_srl_453_n797), .ZN(
        u4_srl_453_n580) );
  AOI22_X1 u4_srl_453_U774 ( .A1(u4_srl_453_n36), .A2(u4_srl_453_n566), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n580), .ZN(u4_srl_453_n796) );
  INV_X1 u4_srl_453_U773 ( .A(u4_srl_453_n796), .ZN(u4_srl_453_n795) );
  AOI221_X1 u4_srl_453_U772 ( .B1(u4_srl_453_n581), .B2(u4_srl_453_n28), .C1(
        u4_srl_453_n576), .C2(u4_srl_453_n91), .A(u4_srl_453_n795), .ZN(
        u4_srl_453_n400) );
  OAI22_X1 u4_srl_453_U771 ( .A1(u4_srl_453_n329), .A2(u4_srl_453_n210), .B1(
        u4_srl_453_n400), .B2(u4_srl_453_n212), .ZN(u4_srl_453_n794) );
  AOI221_X1 u4_srl_453_U770 ( .B1(u4_srl_453_n204), .B2(u4_srl_453_n793), .C1(
        u4_srl_453_n268), .C2(u4_srl_453_n207), .A(u4_srl_453_n794), .ZN(
        u4_srl_453_n786) );
  AOI22_X1 u4_srl_453_U769 ( .A1(net33550), .A2(u4_srl_453_n71), .B1(net33575), 
        .B2(u4_srl_453_n85), .ZN(u4_srl_453_n792) );
  OAI221_X1 u4_srl_453_U768 ( .B1(u4_srl_453_n48), .B2(u4_srl_453_n164), .C1(
        u4_srl_453_n61), .C2(u4_srl_453_n166), .A(u4_srl_453_n792), .ZN(
        u4_srl_453_n254) );
  AOI22_X1 u4_srl_453_U767 ( .A1(net33577), .A2(u4_srl_453_n71), .B1(net33578), 
        .B2(u4_srl_453_n85), .ZN(u4_srl_453_n791) );
  OAI221_X1 u4_srl_453_U766 ( .B1(u4_srl_453_n48), .B2(u4_srl_453_n161), .C1(
        u4_srl_453_n61), .C2(u4_srl_453_n160), .A(u4_srl_453_n791), .ZN(
        u4_srl_453_n258) );
  OAI22_X1 u4_srl_453_U765 ( .A1(u4_srl_453_n169), .A2(u4_srl_453_n76), .B1(
        u4_srl_453_n168), .B2(u4_srl_453_n86), .ZN(u4_srl_453_n790) );
  AOI221_X1 u4_srl_453_U764 ( .B1(u4_srl_453_n54), .B2(net33572), .C1(
        u4_srl_453_n67), .C2(net33573), .A(u4_srl_453_n790), .ZN(
        u4_srl_453_n668) );
  OAI22_X1 u4_srl_453_U763 ( .A1(u4_srl_453_n188), .A2(u4_srl_453_n76), .B1(
        u4_srl_453_n171), .B2(u4_srl_453_n86), .ZN(u4_srl_453_n789) );
  AOI221_X1 u4_srl_453_U762 ( .B1(net33569), .B2(u4_srl_453_n54), .C1(n8520), 
        .C2(u4_srl_453_n67), .A(u4_srl_453_n789), .ZN(u4_srl_453_n572) );
  OAI22_X1 u4_srl_453_U761 ( .A1(u4_srl_453_n668), .A2(u4_srl_453_n201), .B1(
        u4_srl_453_n572), .B2(u4_srl_453_n203), .ZN(u4_srl_453_n788) );
  AOI221_X1 u4_srl_453_U760 ( .B1(u4_srl_453_n195), .B2(u4_srl_453_n254), .C1(
        u4_srl_453_n197), .C2(u4_srl_453_n258), .A(u4_srl_453_n788), .ZN(
        u4_srl_453_n787) );
  AOI21_X1 u4_srl_453_U759 ( .B1(u4_srl_453_n786), .B2(u4_srl_453_n787), .A(
        u4_shift_right[8]), .ZN(u4_N5917) );
  AOI22_X1 u4_srl_453_U758 ( .A1(u4_srl_453_n36), .A2(u4_srl_453_n546), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n542), .ZN(u4_srl_453_n785) );
  INV_X1 u4_srl_453_U757 ( .A(u4_srl_453_n785), .ZN(u4_srl_453_n784) );
  AOI221_X1 u4_srl_453_U756 ( .B1(u4_srl_453_n543), .B2(u4_srl_453_n28), .C1(
        u4_srl_453_n544), .C2(u4_srl_453_n91), .A(u4_srl_453_n784), .ZN(
        u4_srl_453_n478) );
  INV_X1 u4_srl_453_U755 ( .A(u4_srl_453_n478), .ZN(u4_srl_453_n774) );
  INV_X1 u4_srl_453_U754 ( .A(u4_srl_453_n532), .ZN(u4_srl_453_n782) );
  INV_X1 u4_srl_453_U753 ( .A(u4_srl_453_n637), .ZN(u4_srl_453_n528) );
  AOI22_X1 u4_srl_453_U752 ( .A1(u4_srl_453_n36), .A2(u4_srl_453_n412), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n531), .ZN(u4_srl_453_n783) );
  OAI221_X1 u4_srl_453_U751 ( .B1(u4_srl_453_n782), .B2(u4_srl_453_n30), .C1(
        u4_srl_453_n528), .C2(u4_srl_453_n89), .A(u4_srl_453_n783), .ZN(
        u4_srl_453_n392) );
  INV_X1 u4_srl_453_U750 ( .A(u4_srl_453_n392), .ZN(u4_srl_453_n221) );
  INV_X1 u4_srl_453_U749 ( .A(u4_srl_453_n633), .ZN(u4_srl_453_n523) );
  AOI22_X1 u4_srl_453_U748 ( .A1(u4_srl_453_n36), .A2(u4_srl_453_n638), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n526), .ZN(u4_srl_453_n781) );
  OAI221_X1 u4_srl_453_U747 ( .B1(u4_srl_453_n780), .B2(u4_srl_453_n30), .C1(
        u4_srl_453_n523), .C2(u4_srl_453_n89), .A(u4_srl_453_n781), .ZN(
        u4_srl_453_n393) );
  INV_X1 u4_srl_453_U746 ( .A(u4_srl_453_n393), .ZN(u4_srl_453_n312) );
  OAI22_X1 u4_srl_453_U745 ( .A1(u4_srl_453_n221), .A2(u4_srl_453_n275), .B1(
        u4_srl_453_n312), .B2(u4_srl_453_n271), .ZN(u4_srl_453_n267) );
  INV_X1 u4_srl_453_U744 ( .A(u4_srl_453_n641), .ZN(u4_srl_453_n533) );
  AOI22_X1 u4_srl_453_U743 ( .A1(u4_srl_453_n36), .A2(u4_srl_453_n634), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n536), .ZN(u4_srl_453_n779) );
  OAI221_X1 u4_srl_453_U742 ( .B1(u4_srl_453_n778), .B2(u4_srl_453_n30), .C1(
        u4_srl_453_n533), .C2(u4_srl_453_n89), .A(u4_srl_453_n779), .ZN(
        u4_srl_453_n480) );
  INV_X1 u4_srl_453_U741 ( .A(u4_srl_453_n480), .ZN(u4_srl_453_n313) );
  AOI22_X1 u4_srl_453_U740 ( .A1(u4_srl_453_n36), .A2(u4_srl_453_n538), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n549), .ZN(u4_srl_453_n777) );
  INV_X1 u4_srl_453_U739 ( .A(u4_srl_453_n777), .ZN(u4_srl_453_n776) );
  AOI221_X1 u4_srl_453_U738 ( .B1(u4_srl_453_n550), .B2(u4_srl_453_n28), .C1(
        u4_srl_453_n545), .C2(u4_srl_453_n91), .A(u4_srl_453_n776), .ZN(
        u4_srl_453_n395) );
  OAI22_X1 u4_srl_453_U737 ( .A1(u4_srl_453_n313), .A2(u4_srl_453_n210), .B1(
        u4_srl_453_n395), .B2(u4_srl_453_n212), .ZN(u4_srl_453_n775) );
  AOI221_X1 u4_srl_453_U736 ( .B1(u4_srl_453_n204), .B2(u4_srl_453_n774), .C1(
        u4_srl_453_n267), .C2(u4_srl_453_n207), .A(u4_srl_453_n775), .ZN(
        u4_srl_453_n770) );
  INV_X1 u4_srl_453_U735 ( .A(u4_srl_453_n773), .ZN(u4_srl_453_n540) );
  OAI22_X1 u4_srl_453_U734 ( .A1(u4_srl_453_n230), .A2(u4_srl_453_n201), .B1(
        u4_srl_453_n540), .B2(u4_srl_453_n203), .ZN(u4_srl_453_n772) );
  AOI221_X1 u4_srl_453_U733 ( .B1(u4_srl_453_n195), .B2(u4_srl_453_n359), .C1(
        u4_srl_453_n197), .C2(u4_srl_453_n226), .A(u4_srl_453_n772), .ZN(
        u4_srl_453_n771) );
  AOI21_X1 u4_srl_453_U732 ( .B1(u4_srl_453_n770), .B2(u4_srl_453_n771), .A(
        u4_shift_right[8]), .ZN(u4_N5918) );
  AOI22_X1 u4_srl_453_U731 ( .A1(net33558), .A2(u4_srl_453_n71), .B1(net33559), 
        .B2(u4_srl_453_n85), .ZN(u4_srl_453_n769) );
  OAI221_X1 u4_srl_453_U730 ( .B1(u4_srl_453_n48), .B2(u4_srl_453_n187), .C1(
        u4_srl_453_n61), .C2(u4_srl_453_n178), .A(u4_srl_453_n769), .ZN(
        u4_srl_453_n513) );
  AOI22_X1 u4_srl_453_U729 ( .A1(net33562), .A2(u4_srl_453_n71), .B1(n8521), 
        .B2(u4_srl_453_n85), .ZN(u4_srl_453_n768) );
  OAI221_X1 u4_srl_453_U728 ( .B1(u4_srl_453_n48), .B2(u4_srl_453_n176), .C1(
        u4_srl_453_n61), .C2(u4_srl_453_n175), .A(u4_srl_453_n768), .ZN(
        u4_srl_453_n514) );
  AOI22_X1 u4_srl_453_U727 ( .A1(net33586), .A2(u4_srl_453_n71), .B1(net33587), 
        .B2(u4_srl_453_n85), .ZN(u4_srl_453_n767) );
  OAI221_X1 u4_srl_453_U726 ( .B1(u4_srl_453_n48), .B2(u4_srl_453_n192), .C1(
        u4_srl_453_n61), .C2(u4_srl_453_n185), .A(u4_srl_453_n767), .ZN(
        u4_srl_453_n516) );
  AOI22_X1 u4_srl_453_U725 ( .A1(n8524), .A2(u4_srl_453_n71), .B1(n8525), .B2(
        u4_srl_453_n85), .ZN(u4_srl_453_n766) );
  OAI221_X1 u4_srl_453_U724 ( .B1(u4_srl_453_n48), .B2(u4_srl_453_n183), .C1(
        u4_srl_453_n61), .C2(u4_srl_453_n182), .A(u4_srl_453_n766), .ZN(
        u4_srl_453_n512) );
  AOI22_X1 u4_srl_453_U723 ( .A1(u4_srl_453_n36), .A2(u4_srl_453_n516), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n512), .ZN(u4_srl_453_n765) );
  INV_X1 u4_srl_453_U722 ( .A(u4_srl_453_n765), .ZN(u4_srl_453_n764) );
  AOI221_X1 u4_srl_453_U721 ( .B1(u4_srl_453_n513), .B2(u4_srl_453_n27), .C1(
        u4_srl_453_n514), .C2(u4_srl_453_n91), .A(u4_srl_453_n764), .ZN(
        u4_srl_453_n475) );
  INV_X1 u4_srl_453_U720 ( .A(u4_srl_453_n475), .ZN(u4_srl_453_n741) );
  AOI22_X1 u4_srl_453_U719 ( .A1(fract_denorm[96]), .A2(u4_srl_453_n70), .B1(
        fract_denorm[95]), .B2(u4_srl_453_n79), .ZN(u4_srl_453_n763) );
  OAI221_X1 u4_srl_453_U718 ( .B1(u4_srl_453_n57), .B2(u4_srl_453_n103), .C1(
        u4_srl_453_n60), .C2(u4_srl_453_n102), .A(u4_srl_453_n763), .ZN(
        u4_srl_453_n497) );
  AOI22_X1 u4_srl_453_U717 ( .A1(fract_denorm[100]), .A2(u4_srl_453_n70), .B1(
        fract_denorm[99]), .B2(u4_srl_453_n79), .ZN(u4_srl_453_n762) );
  OAI221_X1 u4_srl_453_U716 ( .B1(u4_srl_453_n57), .B2(u4_srl_453_n112), .C1(
        u4_srl_453_n60), .C2(u4_srl_453_n105), .A(u4_srl_453_n762), .ZN(
        u4_srl_453_n502) );
  AOI222_X1 u4_srl_453_U715 ( .A1(u4_srl_453_n497), .A2(u4_srl_453_n88), .B1(
        u4_srl_453_n502), .B2(u4_srl_453_n28), .C1(u4_srl_453_n760), .C2(
        u4_srl_453_n761), .ZN(u4_srl_453_n220) );
  AOI22_X1 u4_srl_453_U714 ( .A1(fract_denorm[84]), .A2(u4_srl_453_n70), .B1(
        fract_denorm[83]), .B2(u4_srl_453_n79), .ZN(u4_srl_453_n759) );
  OAI221_X1 u4_srl_453_U713 ( .B1(u4_srl_453_n48), .B2(u4_srl_453_n150), .C1(
        u4_srl_453_n60), .C2(u4_srl_453_n131), .A(u4_srl_453_n759), .ZN(
        u4_srl_453_n495) );
  INV_X1 u4_srl_453_U712 ( .A(u4_srl_453_n495), .ZN(u4_srl_453_n695) );
  AOI22_X1 u4_srl_453_U711 ( .A1(fract_denorm[80]), .A2(u4_srl_453_n70), .B1(
        fract_denorm[79]), .B2(u4_srl_453_n79), .ZN(u4_srl_453_n758) );
  OAI221_X1 u4_srl_453_U710 ( .B1(u4_srl_453_n48), .B2(u4_srl_453_n129), .C1(
        u4_srl_453_n60), .C2(u4_srl_453_n128), .A(u4_srl_453_n758), .ZN(
        u4_srl_453_n619) );
  INV_X1 u4_srl_453_U709 ( .A(u4_srl_453_n619), .ZN(u4_srl_453_n491) );
  AOI22_X1 u4_srl_453_U708 ( .A1(fract_denorm[92]), .A2(u4_srl_453_n70), .B1(
        fract_denorm[91]), .B2(u4_srl_453_n79), .ZN(u4_srl_453_n757) );
  OAI221_X1 u4_srl_453_U707 ( .B1(u4_srl_453_n48), .B2(u4_srl_453_n107), .C1(
        u4_srl_453_n60), .C2(u4_srl_453_n124), .A(u4_srl_453_n757), .ZN(
        u4_srl_453_n498) );
  AOI22_X1 u4_srl_453_U706 ( .A1(fract_denorm[88]), .A2(u4_srl_453_n70), .B1(
        fract_denorm[87]), .B2(u4_srl_453_n79), .ZN(u4_srl_453_n756) );
  OAI221_X1 u4_srl_453_U705 ( .B1(u4_srl_453_n48), .B2(u4_srl_453_n122), .C1(
        u4_srl_453_n60), .C2(u4_srl_453_n121), .A(u4_srl_453_n756), .ZN(
        u4_srl_453_n494) );
  AOI22_X1 u4_srl_453_U704 ( .A1(u4_srl_453_n36), .A2(u4_srl_453_n498), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n494), .ZN(u4_srl_453_n755) );
  OAI221_X1 u4_srl_453_U703 ( .B1(u4_srl_453_n695), .B2(u4_srl_453_n30), .C1(
        u4_srl_453_n491), .C2(u4_srl_453_n89), .A(u4_srl_453_n755), .ZN(
        u4_srl_453_n388) );
  INV_X1 u4_srl_453_U702 ( .A(u4_srl_453_n388), .ZN(u4_srl_453_n310) );
  OAI22_X1 u4_srl_453_U701 ( .A1(u4_srl_453_n220), .A2(u4_srl_453_n275), .B1(
        u4_srl_453_n310), .B2(u4_srl_453_n271), .ZN(u4_srl_453_n266) );
  AOI22_X1 u4_srl_453_U700 ( .A1(fract_denorm[68]), .A2(u4_srl_453_n70), .B1(
        fract_denorm[67]), .B2(u4_srl_453_n79), .ZN(u4_srl_453_n754) );
  OAI221_X1 u4_srl_453_U699 ( .B1(u4_srl_453_n57), .B2(u4_srl_453_n149), .C1(
        u4_srl_453_n60), .C2(u4_srl_453_n138), .A(u4_srl_453_n754), .ZN(
        u4_srl_453_n508) );
  AOI22_X1 u4_srl_453_U698 ( .A1(fract_denorm[64]), .A2(u4_srl_453_n70), .B1(
        fract_denorm[63]), .B2(u4_srl_453_n79), .ZN(u4_srl_453_n753) );
  OAI221_X1 u4_srl_453_U697 ( .B1(u4_srl_453_n48), .B2(u4_srl_453_n136), .C1(
        u4_srl_453_n60), .C2(u4_srl_453_n135), .A(u4_srl_453_n753), .ZN(
        u4_srl_453_n503) );
  AOI22_X1 u4_srl_453_U696 ( .A1(fract_denorm[76]), .A2(u4_srl_453_n70), .B1(
        fract_denorm[75]), .B2(u4_srl_453_n79), .ZN(u4_srl_453_n752) );
  OAI221_X1 u4_srl_453_U695 ( .B1(u4_srl_453_n48), .B2(u4_srl_453_n151), .C1(
        u4_srl_453_n60), .C2(u4_srl_453_n145), .A(u4_srl_453_n752), .ZN(
        u4_srl_453_n620) );
  AOI22_X1 u4_srl_453_U694 ( .A1(fract_denorm[72]), .A2(u4_srl_453_n70), .B1(
        fract_denorm[71]), .B2(u4_srl_453_n79), .ZN(u4_srl_453_n751) );
  OAI221_X1 u4_srl_453_U693 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n143), .C1(
        u4_srl_453_n60), .C2(u4_srl_453_n142), .A(u4_srl_453_n751), .ZN(
        u4_srl_453_n507) );
  AOI22_X1 u4_srl_453_U692 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n620), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n507), .ZN(u4_srl_453_n750) );
  INV_X1 u4_srl_453_U691 ( .A(u4_srl_453_n750), .ZN(u4_srl_453_n749) );
  AOI221_X1 u4_srl_453_U690 ( .B1(u4_srl_453_n508), .B2(u4_srl_453_n27), .C1(
        u4_srl_453_n503), .C2(u4_srl_453_n91), .A(u4_srl_453_n749), .ZN(
        u4_srl_453_n311) );
  AOI22_X1 u4_srl_453_U689 ( .A1(fract_denorm[52]), .A2(u4_srl_453_n70), .B1(
        fract_denorm[51]), .B2(u4_srl_453_n79), .ZN(u4_srl_453_n748) );
  OAI221_X1 u4_srl_453_U688 ( .B1(u4_srl_453_n52), .B2(u4_srl_453_n153), .C1(
        u4_srl_453_n60), .C2(u4_srl_453_n113), .A(u4_srl_453_n748), .ZN(
        u4_srl_453_n520) );
  AOI22_X1 u4_srl_453_U687 ( .A1(net33583), .A2(u4_srl_453_n70), .B1(n8515), 
        .B2(u4_srl_453_n79), .ZN(u4_srl_453_n747) );
  OAI221_X1 u4_srl_453_U686 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n157), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n156), .A(u4_srl_453_n747), .ZN(
        u4_srl_453_n515) );
  AOI22_X1 u4_srl_453_U685 ( .A1(fract_denorm[60]), .A2(u4_srl_453_n69), .B1(
        fract_denorm[59]), .B2(u4_srl_453_n79), .ZN(u4_srl_453_n746) );
  OAI221_X1 u4_srl_453_U684 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n148), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n117), .A(u4_srl_453_n746), .ZN(
        u4_srl_453_n504) );
  AOI22_X1 u4_srl_453_U683 ( .A1(fract_denorm[56]), .A2(u4_srl_453_n69), .B1(
        fract_denorm[55]), .B2(u4_srl_453_n78), .ZN(u4_srl_453_n745) );
  OAI221_X1 u4_srl_453_U682 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n115), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n114), .A(u4_srl_453_n745), .ZN(
        u4_srl_453_n519) );
  AOI22_X1 u4_srl_453_U681 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n504), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n519), .ZN(u4_srl_453_n744) );
  INV_X1 u4_srl_453_U680 ( .A(u4_srl_453_n744), .ZN(u4_srl_453_n743) );
  AOI221_X1 u4_srl_453_U679 ( .B1(u4_srl_453_n520), .B2(u4_srl_453_n28), .C1(
        u4_srl_453_n515), .C2(u4_srl_453_n91), .A(u4_srl_453_n743), .ZN(
        u4_srl_453_n390) );
  OAI22_X1 u4_srl_453_U678 ( .A1(u4_srl_453_n311), .A2(u4_srl_453_n210), .B1(
        u4_srl_453_n390), .B2(u4_srl_453_n212), .ZN(u4_srl_453_n742) );
  AOI221_X1 u4_srl_453_U677 ( .B1(u4_srl_453_n204), .B2(u4_srl_453_n741), .C1(
        u4_srl_453_n266), .C2(u4_srl_453_n207), .A(u4_srl_453_n742), .ZN(
        u4_srl_453_n734) );
  AOI22_X1 u4_srl_453_U676 ( .A1(net33572), .A2(u4_srl_453_n69), .B1(net33573), 
        .B2(u4_srl_453_n78), .ZN(u4_srl_453_n740) );
  OAI221_X1 u4_srl_453_U675 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n189), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n165), .A(u4_srl_453_n740), .ZN(
        u4_srl_453_n316) );
  AOI22_X1 u4_srl_453_U674 ( .A1(n8516), .A2(u4_srl_453_n69), .B1(n8517), .B2(
        u4_srl_453_n78), .ZN(u4_srl_453_n739) );
  OAI221_X1 u4_srl_453_U673 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n163), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n162), .A(u4_srl_453_n739), .ZN(
        u4_srl_453_n196) );
  OAI22_X1 u4_srl_453_U672 ( .A1(u4_srl_453_n170), .A2(u4_srl_453_n76), .B1(
        u4_srl_453_n172), .B2(u4_srl_453_n86), .ZN(u4_srl_453_n738) );
  AOI221_X1 u4_srl_453_U671 ( .B1(u4_srl_453_n54), .B2(n8519), .C1(
        u4_srl_453_n67), .C2(n8518), .A(u4_srl_453_n738), .ZN(u4_srl_453_n202)
         );
  AOI22_X1 u4_srl_453_U670 ( .A1(net33565), .A2(u4_srl_453_n69), .B1(net33566), 
        .B2(u4_srl_453_n78), .ZN(u4_srl_453_n737) );
  OAI221_X1 u4_srl_453_U669 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n188), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n171), .A(u4_srl_453_n737), .ZN(
        u4_srl_453_n702) );
  INV_X1 u4_srl_453_U668 ( .A(u4_srl_453_n702), .ZN(u4_srl_453_n510) );
  OAI22_X1 u4_srl_453_U667 ( .A1(u4_srl_453_n202), .A2(u4_srl_453_n201), .B1(
        u4_srl_453_n510), .B2(u4_srl_453_n203), .ZN(u4_srl_453_n736) );
  AOI221_X1 u4_srl_453_U666 ( .B1(u4_srl_453_n195), .B2(u4_srl_453_n316), .C1(
        u4_srl_453_n197), .C2(u4_srl_453_n196), .A(u4_srl_453_n736), .ZN(
        u4_srl_453_n735) );
  AOI21_X1 u4_srl_453_U665 ( .B1(u4_srl_453_n734), .B2(u4_srl_453_n735), .A(
        u4_shift_right[8]), .ZN(u4_N5919) );
  AOI22_X1 u4_srl_453_U664 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n607), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n608), .ZN(u4_srl_453_n733) );
  INV_X1 u4_srl_453_U663 ( .A(u4_srl_453_n733), .ZN(u4_srl_453_n732) );
  AOI221_X1 u4_srl_453_U662 ( .B1(u4_srl_453_n605), .B2(u4_srl_453_n27), .C1(
        u4_srl_453_n606), .C2(u4_srl_453_n88), .A(u4_srl_453_n732), .ZN(
        u4_srl_453_n461) );
  INV_X1 u4_srl_453_U661 ( .A(u4_srl_453_n461), .ZN(u4_srl_453_n724) );
  AOI222_X1 u4_srl_453_U660 ( .A1(u4_srl_453_n594), .A2(u4_srl_453_n25), .B1(
        u4_srl_453_n438), .B2(u4_srl_453_n40), .C1(u4_srl_453_n595), .C2(
        u4_srl_453_n441), .ZN(u4_srl_453_n219) );
  INV_X1 u4_srl_453_U659 ( .A(u4_srl_453_n588), .ZN(u4_srl_453_n680) );
  AOI22_X1 u4_srl_453_U658 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n590), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n591), .ZN(u4_srl_453_n731) );
  OAI221_X1 u4_srl_453_U657 ( .B1(u4_srl_453_n680), .B2(u4_srl_453_n30), .C1(
        u4_srl_453_n730), .C2(u4_srl_453_n89), .A(u4_srl_453_n731), .ZN(
        u4_srl_453_n464) );
  INV_X1 u4_srl_453_U656 ( .A(u4_srl_453_n464), .ZN(u4_srl_453_n308) );
  OAI22_X1 u4_srl_453_U655 ( .A1(u4_srl_453_n219), .A2(u4_srl_453_n275), .B1(
        u4_srl_453_n308), .B2(u4_srl_453_n271), .ZN(u4_srl_453_n265) );
  AOI22_X1 u4_srl_453_U654 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n677), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n678), .ZN(u4_srl_453_n729) );
  INV_X1 u4_srl_453_U653 ( .A(u4_srl_453_n729), .ZN(u4_srl_453_n728) );
  AOI221_X1 u4_srl_453_U652 ( .B1(u4_srl_453_n600), .B2(u4_srl_453_n28), .C1(
        u4_srl_453_n601), .C2(u4_srl_453_n88), .A(u4_srl_453_n728), .ZN(
        u4_srl_453_n309) );
  AOI22_X1 u4_srl_453_U651 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n596), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n597), .ZN(u4_srl_453_n727) );
  INV_X1 u4_srl_453_U650 ( .A(u4_srl_453_n727), .ZN(u4_srl_453_n726) );
  AOI221_X1 u4_srl_453_U649 ( .B1(u4_srl_453_n611), .B2(u4_srl_453_n27), .C1(
        u4_srl_453_n612), .C2(u4_srl_453_n88), .A(u4_srl_453_n726), .ZN(
        u4_srl_453_n385) );
  OAI22_X1 u4_srl_453_U648 ( .A1(u4_srl_453_n309), .A2(u4_srl_453_n210), .B1(
        u4_srl_453_n385), .B2(u4_srl_453_n212), .ZN(u4_srl_453_n725) );
  AOI221_X1 u4_srl_453_U647 ( .B1(u4_srl_453_n204), .B2(u4_srl_453_n724), .C1(
        u4_srl_453_n265), .C2(u4_srl_453_n207), .A(u4_srl_453_n725), .ZN(
        u4_srl_453_n721) );
  INV_X1 u4_srl_453_U646 ( .A(u4_srl_453_n687), .ZN(u4_srl_453_n602) );
  OAI22_X1 u4_srl_453_U645 ( .A1(u4_srl_453_n603), .A2(u4_srl_453_n201), .B1(
        u4_srl_453_n602), .B2(u4_srl_453_n203), .ZN(u4_srl_453_n723) );
  AOI221_X1 u4_srl_453_U644 ( .B1(u4_srl_453_n195), .B2(u4_srl_453_n285), .C1(
        u4_srl_453_n197), .C2(u4_srl_453_n286), .A(u4_srl_453_n723), .ZN(
        u4_srl_453_n722) );
  AOI21_X1 u4_srl_453_U643 ( .B1(u4_srl_453_n721), .B2(u4_srl_453_n722), .A(
        u4_shift_right[8]), .ZN(u4_N5920) );
  AOI22_X1 u4_srl_453_U642 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n576), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n577), .ZN(u4_srl_453_n720) );
  INV_X1 u4_srl_453_U641 ( .A(u4_srl_453_n720), .ZN(u4_srl_453_n719) );
  AOI221_X1 u4_srl_453_U640 ( .B1(u4_srl_453_n574), .B2(u4_srl_453_n27), .C1(
        u4_srl_453_n575), .C2(u4_srl_453_n88), .A(u4_srl_453_n719), .ZN(
        u4_srl_453_n456) );
  INV_X1 u4_srl_453_U639 ( .A(u4_srl_453_n456), .ZN(u4_srl_453_n711) );
  AOI222_X1 u4_srl_453_U638 ( .A1(u4_srl_453_n563), .A2(u4_srl_453_n25), .B1(
        u4_srl_453_n435), .B2(u4_srl_453_n40), .C1(u4_srl_453_n564), .C2(
        u4_srl_453_n91), .ZN(u4_srl_453_n218) );
  INV_X1 u4_srl_453_U637 ( .A(u4_srl_453_n557), .ZN(u4_srl_453_n663) );
  AOI22_X1 u4_srl_453_U636 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n559), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n560), .ZN(u4_srl_453_n718) );
  OAI221_X1 u4_srl_453_U635 ( .B1(u4_srl_453_n663), .B2(u4_srl_453_n30), .C1(
        u4_srl_453_n717), .C2(u4_srl_453_n89), .A(u4_srl_453_n718), .ZN(
        u4_srl_453_n459) );
  INV_X1 u4_srl_453_U634 ( .A(u4_srl_453_n459), .ZN(u4_srl_453_n306) );
  OAI22_X1 u4_srl_453_U633 ( .A1(u4_srl_453_n218), .A2(u4_srl_453_n275), .B1(
        u4_srl_453_n306), .B2(u4_srl_453_n271), .ZN(u4_srl_453_n264) );
  INV_X1 u4_srl_453_U632 ( .A(u4_srl_453_n569), .ZN(u4_srl_453_n658) );
  INV_X1 u4_srl_453_U631 ( .A(u4_srl_453_n570), .ZN(u4_srl_453_n715) );
  AOI22_X1 u4_srl_453_U630 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n660), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n661), .ZN(u4_srl_453_n716) );
  OAI221_X1 u4_srl_453_U629 ( .B1(u4_srl_453_n658), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n715), .C2(u4_srl_453_n89), .A(u4_srl_453_n716), .ZN(
        u4_srl_453_n458) );
  INV_X1 u4_srl_453_U628 ( .A(u4_srl_453_n458), .ZN(u4_srl_453_n307) );
  AOI22_X1 u4_srl_453_U627 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n565), .B1(
        u4_srl_453_n44), .B2(u4_srl_453_n566), .ZN(u4_srl_453_n714) );
  INV_X1 u4_srl_453_U626 ( .A(u4_srl_453_n714), .ZN(u4_srl_453_n713) );
  AOI221_X1 u4_srl_453_U625 ( .B1(u4_srl_453_n580), .B2(u4_srl_453_n27), .C1(
        u4_srl_453_n581), .C2(u4_srl_453_n88), .A(u4_srl_453_n713), .ZN(
        u4_srl_453_n382) );
  OAI22_X1 u4_srl_453_U624 ( .A1(u4_srl_453_n307), .A2(u4_srl_453_n210), .B1(
        u4_srl_453_n382), .B2(u4_srl_453_n212), .ZN(u4_srl_453_n712) );
  AOI221_X1 u4_srl_453_U623 ( .B1(u4_srl_453_n204), .B2(u4_srl_453_n711), .C1(
        u4_srl_453_n264), .C2(u4_srl_453_n207), .A(u4_srl_453_n712), .ZN(
        u4_srl_453_n708) );
  INV_X1 u4_srl_453_U622 ( .A(u4_srl_453_n668), .ZN(u4_srl_453_n252) );
  INV_X1 u4_srl_453_U621 ( .A(u4_srl_453_n670), .ZN(u4_srl_453_n571) );
  OAI22_X1 u4_srl_453_U620 ( .A1(u4_srl_453_n572), .A2(u4_srl_453_n201), .B1(
        u4_srl_453_n571), .B2(u4_srl_453_n203), .ZN(u4_srl_453_n710) );
  AOI221_X1 u4_srl_453_U619 ( .B1(u4_srl_453_n195), .B2(u4_srl_453_n252), .C1(
        u4_srl_453_n197), .C2(u4_srl_453_n254), .A(u4_srl_453_n710), .ZN(
        u4_srl_453_n709) );
  AOI21_X1 u4_srl_453_U618 ( .B1(u4_srl_453_n708), .B2(u4_srl_453_n709), .A(
        u4_shift_right[8]), .ZN(u4_N5921) );
  AOI22_X1 u4_srl_453_U617 ( .A1(u4_srl_453_n378), .A2(u4_srl_453_n433), .B1(
        u4_srl_453_n379), .B2(u4_srl_453_n432), .ZN(u4_srl_453_n248) );
  INV_X1 u4_srl_453_U616 ( .A(u4_srl_453_n455), .ZN(u4_srl_453_n375) );
  OAI222_X1 u4_srl_453_U615 ( .A1(u4_srl_453_n4), .A2(u4_srl_453_n376), .B1(
        u4_srl_453_n415), .B2(u4_srl_453_n248), .C1(u4_srl_453_n2), .C2(
        u4_srl_453_n375), .ZN(u4_srl_453_n707) );
  INV_X1 u4_srl_453_U614 ( .A(u4_srl_453_n707), .ZN(u4_srl_453_n706) );
  OAI221_X1 u4_srl_453_U613 ( .B1(u4_srl_453_n453), .B2(u4_srl_453_n15), .C1(
        u4_srl_453_n705), .C2(u4_srl_453_n10), .A(u4_srl_453_n706), .ZN(
        u4_N5922) );
  AOI22_X1 u4_srl_453_U612 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n515), .B1(
        u4_srl_453_n44), .B2(u4_srl_453_n516), .ZN(u4_srl_453_n704) );
  INV_X1 u4_srl_453_U611 ( .A(u4_srl_453_n704), .ZN(u4_srl_453_n703) );
  AOI221_X1 u4_srl_453_U610 ( .B1(u4_srl_453_n512), .B2(u4_srl_453_n27), .C1(
        u4_srl_453_n513), .C2(u4_srl_453_n88), .A(u4_srl_453_n703), .ZN(
        u4_srl_453_n450) );
  INV_X1 u4_srl_453_U609 ( .A(u4_srl_453_n316), .ZN(u4_srl_453_n200) );
  AOI22_X1 u4_srl_453_U608 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n514), .B1(
        u4_srl_453_n44), .B2(u4_srl_453_n702), .ZN(u4_srl_453_n701) );
  OAI221_X1 u4_srl_453_U607 ( .B1(u4_srl_453_n202), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n200), .C2(u4_srl_453_n89), .A(u4_srl_453_n701), .ZN(
        u4_srl_453_n700) );
  INV_X1 u4_srl_453_U606 ( .A(u4_srl_453_n700), .ZN(u4_srl_453_n650) );
  AOI22_X1 u4_srl_453_U605 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n503), .B1(
        u4_srl_453_n44), .B2(u4_srl_453_n504), .ZN(u4_srl_453_n699) );
  INV_X1 u4_srl_453_U604 ( .A(u4_srl_453_n699), .ZN(u4_srl_453_n698) );
  AOI221_X1 u4_srl_453_U603 ( .B1(u4_srl_453_n519), .B2(u4_srl_453_n27), .C1(
        u4_srl_453_n520), .C2(u4_srl_453_n88), .A(u4_srl_453_n698), .ZN(
        u4_srl_453_n371) );
  AOI222_X1 u4_srl_453_U602 ( .A1(u4_srl_453_n501), .A2(u4_srl_453_n25), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n697), .C1(u4_srl_453_n502), .C2(
        u4_srl_453_n91), .ZN(u4_srl_453_n216) );
  INV_X1 u4_srl_453_U601 ( .A(u4_srl_453_n216), .ZN(u4_srl_453_n373) );
  INV_X1 u4_srl_453_U600 ( .A(u4_srl_453_n494), .ZN(u4_srl_453_n694) );
  AOI22_X1 u4_srl_453_U599 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n497), .B1(
        u4_srl_453_n44), .B2(u4_srl_453_n498), .ZN(u4_srl_453_n696) );
  OAI221_X1 u4_srl_453_U598 ( .B1(u4_srl_453_n694), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n695), .C2(u4_srl_453_n89), .A(u4_srl_453_n696), .ZN(
        u4_srl_453_n374) );
  AOI22_X1 u4_srl_453_U597 ( .A1(u4_srl_453_n373), .A2(u4_srl_453_n433), .B1(
        u4_srl_453_n374), .B2(u4_srl_453_n432), .ZN(u4_srl_453_n247) );
  AOI22_X1 u4_srl_453_U596 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n619), .B1(
        u4_srl_453_n44), .B2(u4_srl_453_n620), .ZN(u4_srl_453_n693) );
  INV_X1 u4_srl_453_U595 ( .A(u4_srl_453_n693), .ZN(u4_srl_453_n692) );
  AOI221_X1 u4_srl_453_U594 ( .B1(u4_srl_453_n507), .B2(u4_srl_453_n27), .C1(
        u4_srl_453_n508), .C2(u4_srl_453_n88), .A(u4_srl_453_n692), .ZN(
        u4_srl_453_n370) );
  OAI222_X1 u4_srl_453_U593 ( .A1(u4_srl_453_n4), .A2(u4_srl_453_n371), .B1(
        u4_srl_453_n415), .B2(u4_srl_453_n247), .C1(u4_srl_453_n2), .C2(
        u4_srl_453_n370), .ZN(u4_srl_453_n691) );
  INV_X1 u4_srl_453_U592 ( .A(u4_srl_453_n691), .ZN(u4_srl_453_n690) );
  OAI221_X1 u4_srl_453_U591 ( .B1(u4_srl_453_n450), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n650), .C2(u4_srl_453_n10), .A(u4_srl_453_n690), .ZN(
        u4_N5923) );
  AOI22_X1 u4_srl_453_U590 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n612), .B1(
        u4_srl_453_n44), .B2(u4_srl_453_n607), .ZN(u4_srl_453_n689) );
  INV_X1 u4_srl_453_U589 ( .A(u4_srl_453_n689), .ZN(u4_srl_453_n688) );
  AOI221_X1 u4_srl_453_U588 ( .B1(u4_srl_453_n608), .B2(u4_srl_453_n27), .C1(
        u4_srl_453_n605), .C2(u4_srl_453_n88), .A(u4_srl_453_n688), .ZN(
        u4_srl_453_n447) );
  AOI22_X1 u4_srl_453_U587 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n606), .B1(
        u4_srl_453_n44), .B2(u4_srl_453_n687), .ZN(u4_srl_453_n686) );
  OAI221_X1 u4_srl_453_U586 ( .B1(u4_srl_453_n603), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n685), .C2(u4_srl_453_n89), .A(u4_srl_453_n686), .ZN(
        u4_srl_453_n684) );
  INV_X1 u4_srl_453_U585 ( .A(u4_srl_453_n684), .ZN(u4_srl_453_n471) );
  AOI22_X1 u4_srl_453_U584 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n601), .B1(
        u4_srl_453_n44), .B2(u4_srl_453_n596), .ZN(u4_srl_453_n683) );
  INV_X1 u4_srl_453_U583 ( .A(u4_srl_453_n683), .ZN(u4_srl_453_n682) );
  AOI221_X1 u4_srl_453_U582 ( .B1(u4_srl_453_n597), .B2(u4_srl_453_n27), .C1(
        u4_srl_453_n611), .C2(u4_srl_453_n87), .A(u4_srl_453_n682), .ZN(
        u4_srl_453_n353) );
  AOI22_X1 u4_srl_453_U581 ( .A1(u4_srl_453_n594), .A2(u4_srl_453_n91), .B1(
        u4_srl_453_n438), .B2(u4_srl_453_n28), .ZN(u4_srl_453_n215) );
  INV_X1 u4_srl_453_U580 ( .A(u4_srl_453_n215), .ZN(u4_srl_453_n355) );
  INV_X1 u4_srl_453_U579 ( .A(u4_srl_453_n591), .ZN(u4_srl_453_n679) );
  AOI22_X1 u4_srl_453_U578 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n595), .B1(
        u4_srl_453_n44), .B2(u4_srl_453_n590), .ZN(u4_srl_453_n681) );
  OAI221_X1 u4_srl_453_U577 ( .B1(u4_srl_453_n679), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n680), .C2(u4_srl_453_n89), .A(u4_srl_453_n681), .ZN(
        u4_srl_453_n356) );
  AOI22_X1 u4_srl_453_U576 ( .A1(u4_srl_453_n355), .A2(u4_srl_453_n433), .B1(
        u4_srl_453_n356), .B2(u4_srl_453_n432), .ZN(u4_srl_453_n246) );
  INV_X1 u4_srl_453_U575 ( .A(u4_srl_453_n678), .ZN(u4_srl_453_n586) );
  INV_X1 u4_srl_453_U574 ( .A(u4_srl_453_n600), .ZN(u4_srl_453_n675) );
  AOI22_X1 u4_srl_453_U573 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n589), .B1(
        u4_srl_453_n43), .B2(u4_srl_453_n677), .ZN(u4_srl_453_n676) );
  OAI221_X1 u4_srl_453_U572 ( .B1(u4_srl_453_n586), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n675), .C2(u4_srl_453_n89), .A(u4_srl_453_n676), .ZN(
        u4_srl_453_n449) );
  INV_X1 u4_srl_453_U571 ( .A(u4_srl_453_n449), .ZN(u4_srl_453_n352) );
  OAI222_X1 u4_srl_453_U570 ( .A1(u4_srl_453_n4), .A2(u4_srl_453_n353), .B1(
        u4_srl_453_n415), .B2(u4_srl_453_n246), .C1(u4_srl_453_n2), .C2(
        u4_srl_453_n352), .ZN(u4_srl_453_n674) );
  INV_X1 u4_srl_453_U569 ( .A(u4_srl_453_n674), .ZN(u4_srl_453_n673) );
  OAI221_X1 u4_srl_453_U568 ( .B1(u4_srl_453_n447), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n471), .C2(u4_srl_453_n10), .A(u4_srl_453_n673), .ZN(
        u4_N5924) );
  AOI22_X1 u4_srl_453_U567 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n581), .B1(
        u4_srl_453_n43), .B2(u4_srl_453_n576), .ZN(u4_srl_453_n672) );
  INV_X1 u4_srl_453_U566 ( .A(u4_srl_453_n672), .ZN(u4_srl_453_n671) );
  AOI221_X1 u4_srl_453_U565 ( .B1(u4_srl_453_n577), .B2(u4_srl_453_n27), .C1(
        u4_srl_453_n574), .C2(u4_srl_453_n87), .A(u4_srl_453_n671), .ZN(
        u4_srl_453_n430) );
  AOI22_X1 u4_srl_453_U564 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n575), .B1(
        u4_srl_453_n43), .B2(u4_srl_453_n670), .ZN(u4_srl_453_n669) );
  OAI221_X1 u4_srl_453_U563 ( .B1(u4_srl_453_n572), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n668), .C2(u4_srl_453_n89), .A(u4_srl_453_n669), .ZN(
        u4_srl_453_n667) );
  INV_X1 u4_srl_453_U562 ( .A(u4_srl_453_n667), .ZN(u4_srl_453_n422) );
  AOI22_X1 u4_srl_453_U561 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n570), .B1(
        u4_srl_453_n43), .B2(u4_srl_453_n565), .ZN(u4_srl_453_n666) );
  INV_X1 u4_srl_453_U560 ( .A(u4_srl_453_n666), .ZN(u4_srl_453_n665) );
  AOI221_X1 u4_srl_453_U559 ( .B1(u4_srl_453_n566), .B2(u4_srl_453_n26), .C1(
        u4_srl_453_n580), .C2(u4_srl_453_n88), .A(u4_srl_453_n665), .ZN(
        u4_srl_453_n348) );
  AOI22_X1 u4_srl_453_U558 ( .A1(u4_srl_453_n563), .A2(u4_srl_453_n91), .B1(
        u4_srl_453_n435), .B2(u4_srl_453_n28), .ZN(u4_srl_453_n213) );
  INV_X1 u4_srl_453_U557 ( .A(u4_srl_453_n213), .ZN(u4_srl_453_n350) );
  INV_X1 u4_srl_453_U556 ( .A(u4_srl_453_n560), .ZN(u4_srl_453_n662) );
  AOI22_X1 u4_srl_453_U555 ( .A1(u4_srl_453_n34), .A2(u4_srl_453_n564), .B1(
        u4_srl_453_n43), .B2(u4_srl_453_n559), .ZN(u4_srl_453_n664) );
  OAI221_X1 u4_srl_453_U554 ( .B1(u4_srl_453_n662), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n663), .C2(u4_srl_453_n89), .A(u4_srl_453_n664), .ZN(
        u4_srl_453_n351) );
  AOI22_X1 u4_srl_453_U553 ( .A1(u4_srl_453_n350), .A2(u4_srl_453_n433), .B1(
        u4_srl_453_n351), .B2(u4_srl_453_n432), .ZN(u4_srl_453_n244) );
  INV_X1 u4_srl_453_U552 ( .A(u4_srl_453_n661), .ZN(u4_srl_453_n555) );
  AOI22_X1 u4_srl_453_U551 ( .A1(u4_srl_453_n34), .A2(u4_srl_453_n558), .B1(
        u4_srl_453_n43), .B2(u4_srl_453_n660), .ZN(u4_srl_453_n659) );
  OAI221_X1 u4_srl_453_U550 ( .B1(u4_srl_453_n555), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n658), .C2(u4_srl_453_n89), .A(u4_srl_453_n659), .ZN(
        u4_srl_453_n431) );
  INV_X1 u4_srl_453_U549 ( .A(u4_srl_453_n431), .ZN(u4_srl_453_n347) );
  OAI222_X1 u4_srl_453_U548 ( .A1(u4_srl_453_n4), .A2(u4_srl_453_n348), .B1(
        u4_srl_453_n415), .B2(u4_srl_453_n244), .C1(u4_srl_453_n2), .C2(
        u4_srl_453_n347), .ZN(u4_srl_453_n657) );
  INV_X1 u4_srl_453_U547 ( .A(u4_srl_453_n657), .ZN(u4_srl_453_n656) );
  OAI221_X1 u4_srl_453_U546 ( .B1(u4_srl_453_n430), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n422), .C2(u4_srl_453_n9), .A(u4_srl_453_n656), .ZN(
        u4_N5925) );
  INV_X1 u4_srl_453_U545 ( .A(u4_srl_453_n370), .ZN(u4_srl_453_n452) );
  AOI222_X1 u4_srl_453_U544 ( .A1(u4_srl_453_n452), .A2(u4_srl_453_n432), .B1(
        u4_srl_453_n373), .B2(u4_srl_453_n368), .C1(u4_srl_453_n374), .C2(
        u4_srl_453_n433), .ZN(u4_srl_453_n304) );
  INV_X1 u4_srl_453_U543 ( .A(u4_srl_453_n450), .ZN(u4_srl_453_n646) );
  AOI22_X1 u4_srl_453_U542 ( .A1(u4_srl_453_n67), .A2(net33648), .B1(
        u4_srl_453_n54), .B2(net33647), .ZN(u4_srl_453_n655) );
  INV_X1 u4_srl_453_U541 ( .A(u4_srl_453_n655), .ZN(u4_srl_453_n654) );
  AOI221_X1 u4_srl_453_U540 ( .B1(n8512), .B2(u4_srl_453_n69), .C1(n8511), 
        .C2(u4_srl_453_n78), .A(u4_srl_453_n654), .ZN(u4_srl_453_n648) );
  AOI22_X1 u4_srl_453_U539 ( .A1(net33641), .A2(u4_srl_453_n69), .B1(net33642), 
        .B2(u4_srl_453_n78), .ZN(u4_srl_453_n653) );
  OAI221_X1 u4_srl_453_U538 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n97), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n96), .A(u4_srl_453_n653), .ZN(
        u4_srl_453_n319) );
  AOI22_X1 u4_srl_453_U537 ( .A1(net33579), .A2(u4_srl_453_n69), .B1(net33581), 
        .B2(u4_srl_453_n78), .ZN(u4_srl_453_n652) );
  OAI221_X1 u4_srl_453_U536 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n190), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n191), .A(u4_srl_453_n652), .ZN(
        u4_srl_453_n198) );
  AOI222_X1 u4_srl_453_U535 ( .A1(u4_srl_453_n25), .A2(u4_srl_453_n319), .B1(
        u4_srl_453_n35), .B2(u4_srl_453_n196), .C1(u4_srl_453_n40), .C2(
        u4_srl_453_n198), .ZN(u4_srl_453_n651) );
  MUX2_X1 u4_srl_453_U534 ( .A(u4_srl_453_n650), .B(u4_srl_453_n651), .S(
        u4_srl_453_n424), .Z(u4_srl_453_n649) );
  OAI21_X1 u4_srl_453_U533 ( .B1(u4_srl_453_n648), .B2(u4_srl_453_n298), .A(
        u4_srl_453_n649), .ZN(u4_srl_453_n647) );
  AOI22_X1 u4_srl_453_U532 ( .A1(u4_srl_453_n23), .A2(u4_srl_453_n646), .B1(
        u4_srl_453_n418), .B2(u4_srl_453_n647), .ZN(u4_srl_453_n645) );
  OAI221_X1 u4_srl_453_U531 ( .B1(u4_srl_453_n304), .B2(u4_srl_453_n415), .C1(
        u4_srl_453_n371), .C2(u4_srl_453_n2), .A(u4_srl_453_n645), .ZN(
        u4_N5907) );
  AOI22_X1 u4_srl_453_U530 ( .A1(u4_srl_453_n34), .A2(u4_srl_453_n550), .B1(
        u4_srl_453_n43), .B2(u4_srl_453_n545), .ZN(u4_srl_453_n644) );
  INV_X1 u4_srl_453_U529 ( .A(u4_srl_453_n644), .ZN(u4_srl_453_n643) );
  AOI221_X1 u4_srl_453_U528 ( .B1(u4_srl_453_n546), .B2(u4_srl_453_n26), .C1(
        u4_srl_453_n542), .C2(u4_srl_453_n87), .A(u4_srl_453_n643), .ZN(
        u4_srl_453_n365) );
  AOI22_X1 u4_srl_453_U527 ( .A1(u4_srl_453_n34), .A2(u4_srl_453_n543), .B1(
        u4_srl_453_n43), .B2(u4_srl_453_n544), .ZN(u4_srl_453_n642) );
  OAI221_X1 u4_srl_453_U526 ( .B1(u4_srl_453_n540), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n230), .C2(u4_srl_453_n89), .A(u4_srl_453_n642), .ZN(
        u4_srl_453_n363) );
  INV_X1 u4_srl_453_U525 ( .A(u4_srl_453_n363), .ZN(u4_srl_453_n628) );
  AOI22_X1 u4_srl_453_U524 ( .A1(u4_srl_453_n34), .A2(u4_srl_453_n537), .B1(
        u4_srl_453_n43), .B2(u4_srl_453_n641), .ZN(u4_srl_453_n640) );
  INV_X1 u4_srl_453_U523 ( .A(u4_srl_453_n640), .ZN(u4_srl_453_n639) );
  AOI221_X1 u4_srl_453_U522 ( .B1(u4_srl_453_n538), .B2(u4_srl_453_n27), .C1(
        u4_srl_453_n549), .C2(u4_srl_453_n87), .A(u4_srl_453_n639), .ZN(
        u4_srl_453_n343) );
  INV_X1 u4_srl_453_U521 ( .A(u4_srl_453_n343), .ZN(u4_srl_453_n630) );
  INV_X1 u4_srl_453_U520 ( .A(u4_srl_453_n638), .ZN(u4_srl_453_n529) );
  AOI22_X1 u4_srl_453_U519 ( .A1(u4_srl_453_n34), .A2(u4_srl_453_n532), .B1(
        u4_srl_453_n42), .B2(u4_srl_453_n637), .ZN(u4_srl_453_n636) );
  OAI221_X1 u4_srl_453_U518 ( .B1(u4_srl_453_n529), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n635), .C2(u4_srl_453_n89), .A(u4_srl_453_n636), .ZN(
        u4_srl_453_n346) );
  INV_X1 u4_srl_453_U517 ( .A(u4_srl_453_n346), .ZN(u4_srl_453_n367) );
  OAI22_X1 u4_srl_453_U516 ( .A1(u4_srl_453_n366), .A2(u4_srl_453_n275), .B1(
        u4_srl_453_n367), .B2(u4_srl_453_n271), .ZN(u4_srl_453_n242) );
  INV_X1 u4_srl_453_U515 ( .A(u4_srl_453_n634), .ZN(u4_srl_453_n524) );
  AOI22_X1 u4_srl_453_U514 ( .A1(u4_srl_453_n34), .A2(u4_srl_453_n527), .B1(
        u4_srl_453_n42), .B2(u4_srl_453_n633), .ZN(u4_srl_453_n632) );
  OAI221_X1 u4_srl_453_U513 ( .B1(u4_srl_453_n524), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n631), .C2(u4_srl_453_n89), .A(u4_srl_453_n632), .ZN(
        u4_srl_453_n369) );
  AOI222_X1 u4_srl_453_U512 ( .A1(u4_srl_453_n24), .A2(u4_srl_453_n630), .B1(
        u4_srl_453_n408), .B2(u4_srl_453_n242), .C1(u4_srl_453_n22), .C2(
        u4_srl_453_n369), .ZN(u4_srl_453_n629) );
  OAI221_X1 u4_srl_453_U511 ( .B1(u4_srl_453_n365), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n628), .C2(u4_srl_453_n10), .A(u4_srl_453_n629), .ZN(
        u4_N5926) );
  AOI22_X1 u4_srl_453_U510 ( .A1(u4_srl_453_n34), .A2(u4_srl_453_n520), .B1(
        u4_srl_453_n42), .B2(u4_srl_453_n515), .ZN(u4_srl_453_n627) );
  INV_X1 u4_srl_453_U509 ( .A(u4_srl_453_n627), .ZN(u4_srl_453_n626) );
  AOI221_X1 u4_srl_453_U508 ( .B1(u4_srl_453_n516), .B2(u4_srl_453_n26), .C1(
        u4_srl_453_n512), .C2(u4_srl_453_n87), .A(u4_srl_453_n626), .ZN(
        u4_srl_453_n323) );
  AOI22_X1 u4_srl_453_U507 ( .A1(u4_srl_453_n34), .A2(u4_srl_453_n513), .B1(
        u4_srl_453_n42), .B2(u4_srl_453_n514), .ZN(u4_srl_453_n625) );
  OAI221_X1 u4_srl_453_U506 ( .B1(u4_srl_453_n510), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n202), .C2(u4_srl_453_n89), .A(u4_srl_453_n625), .ZN(
        u4_srl_453_n320) );
  INV_X1 u4_srl_453_U505 ( .A(u4_srl_453_n320), .ZN(u4_srl_453_n613) );
  AOI22_X1 u4_srl_453_U504 ( .A1(u4_srl_453_n34), .A2(u4_srl_453_n508), .B1(
        u4_srl_453_n42), .B2(u4_srl_453_n503), .ZN(u4_srl_453_n624) );
  INV_X1 u4_srl_453_U503 ( .A(u4_srl_453_n624), .ZN(u4_srl_453_n623) );
  AOI221_X1 u4_srl_453_U502 ( .B1(u4_srl_453_n504), .B2(u4_srl_453_n27), .C1(
        u4_srl_453_n519), .C2(u4_srl_453_n87), .A(u4_srl_453_n623), .ZN(
        u4_srl_453_n322) );
  INV_X1 u4_srl_453_U501 ( .A(u4_srl_453_n322), .ZN(u4_srl_453_n615) );
  AND2_X1 u4_srl_453_U500 ( .A1(u4_srl_453_n408), .A2(u4_srl_453_n299), .ZN(
        u4_srl_453_n490) );
  AOI22_X1 u4_srl_453_U499 ( .A1(u4_srl_453_n34), .A2(u4_srl_453_n502), .B1(
        u4_srl_453_n42), .B2(u4_srl_453_n497), .ZN(u4_srl_453_n622) );
  INV_X1 u4_srl_453_U498 ( .A(u4_srl_453_n622), .ZN(u4_srl_453_n621) );
  AOI221_X1 u4_srl_453_U497 ( .B1(u4_srl_453_n498), .B2(u4_srl_453_n27), .C1(
        u4_srl_453_n494), .C2(u4_srl_453_n88), .A(u4_srl_453_n621), .ZN(
        u4_srl_453_n327) );
  MUX2_X1 u4_srl_453_U496 ( .A(u4_srl_453_n325), .B(u4_srl_453_n327), .S(
        u4_srl_453_n424), .Z(u4_srl_453_n241) );
  INV_X1 u4_srl_453_U495 ( .A(u4_srl_453_n241), .ZN(u4_srl_453_n616) );
  INV_X1 u4_srl_453_U494 ( .A(u4_srl_453_n620), .ZN(u4_srl_453_n492) );
  INV_X1 u4_srl_453_U493 ( .A(u4_srl_453_n507), .ZN(u4_srl_453_n617) );
  AOI22_X1 u4_srl_453_U492 ( .A1(u4_srl_453_n34), .A2(u4_srl_453_n495), .B1(
        u4_srl_453_n43), .B2(u4_srl_453_n619), .ZN(u4_srl_453_n618) );
  OAI221_X1 u4_srl_453_U491 ( .B1(u4_srl_453_n492), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n617), .C2(u4_srl_453_n89), .A(u4_srl_453_n618), .ZN(
        u4_srl_453_n341) );
  AOI222_X1 u4_srl_453_U490 ( .A1(u4_srl_453_n24), .A2(u4_srl_453_n615), .B1(
        u4_srl_453_n490), .B2(u4_srl_453_n616), .C1(u4_srl_453_n22), .C2(
        u4_srl_453_n341), .ZN(u4_srl_453_n614) );
  OAI221_X1 u4_srl_453_U489 ( .B1(u4_srl_453_n323), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n613), .C2(u4_srl_453_n10), .A(u4_srl_453_n614), .ZN(
        u4_N5927) );
  AOI22_X1 u4_srl_453_U488 ( .A1(u4_srl_453_n33), .A2(u4_srl_453_n611), .B1(
        u4_srl_453_n42), .B2(u4_srl_453_n612), .ZN(u4_srl_453_n610) );
  INV_X1 u4_srl_453_U487 ( .A(u4_srl_453_n610), .ZN(u4_srl_453_n609) );
  AOI221_X1 u4_srl_453_U486 ( .B1(u4_srl_453_n607), .B2(u4_srl_453_n26), .C1(
        u4_srl_453_n608), .C2(u4_srl_453_n87), .A(u4_srl_453_n609), .ZN(
        u4_srl_453_n294) );
  AOI22_X1 u4_srl_453_U485 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n605), .B1(
        u4_srl_453_n44), .B2(u4_srl_453_n606), .ZN(u4_srl_453_n604) );
  OAI221_X1 u4_srl_453_U484 ( .B1(u4_srl_453_n602), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n603), .C2(u4_srl_453_n89), .A(u4_srl_453_n604), .ZN(
        u4_srl_453_n291) );
  INV_X1 u4_srl_453_U483 ( .A(u4_srl_453_n291), .ZN(u4_srl_453_n582) );
  AOI22_X1 u4_srl_453_U482 ( .A1(u4_srl_453_n33), .A2(u4_srl_453_n600), .B1(
        u4_srl_453_n42), .B2(u4_srl_453_n601), .ZN(u4_srl_453_n599) );
  INV_X1 u4_srl_453_U481 ( .A(u4_srl_453_n599), .ZN(u4_srl_453_n598) );
  AOI221_X1 u4_srl_453_U480 ( .B1(u4_srl_453_n596), .B2(u4_srl_453_n26), .C1(
        u4_srl_453_n597), .C2(u4_srl_453_n87), .A(u4_srl_453_n598), .ZN(
        u4_srl_453_n293) );
  INV_X1 u4_srl_453_U479 ( .A(u4_srl_453_n293), .ZN(u4_srl_453_n584) );
  AOI22_X1 u4_srl_453_U478 ( .A1(u4_srl_453_n33), .A2(u4_srl_453_n594), .B1(
        u4_srl_453_n43), .B2(u4_srl_453_n595), .ZN(u4_srl_453_n593) );
  INV_X1 u4_srl_453_U477 ( .A(u4_srl_453_n593), .ZN(u4_srl_453_n592) );
  AOI221_X1 u4_srl_453_U476 ( .B1(u4_srl_453_n590), .B2(u4_srl_453_n26), .C1(
        u4_srl_453_n591), .C2(u4_srl_453_n87), .A(u4_srl_453_n592), .ZN(
        u4_srl_453_n297) );
  NAND2_X1 u4_srl_453_U475 ( .A1(u4_srl_453_n91), .A2(u4_shift_right[4]), .ZN(
        u4_srl_453_n496) );
  OAI22_X1 u4_srl_453_U474 ( .A1(u4_shift_right[4]), .A2(u4_srl_453_n297), 
        .B1(u4_srl_453_n296), .B2(u4_srl_453_n496), .ZN(u4_srl_453_n339) );
  AOI22_X1 u4_srl_453_U473 ( .A1(u4_srl_453_n33), .A2(u4_srl_453_n588), .B1(
        u4_srl_453_n41), .B2(u4_srl_453_n589), .ZN(u4_srl_453_n587) );
  OAI221_X1 u4_srl_453_U472 ( .B1(u4_srl_453_n585), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n586), .C2(u4_srl_453_n89), .A(u4_srl_453_n587), .ZN(
        u4_srl_453_n340) );
  AOI222_X1 u4_srl_453_U471 ( .A1(u4_srl_453_n24), .A2(u4_srl_453_n584), .B1(
        u4_srl_453_n490), .B2(u4_srl_453_n339), .C1(u4_srl_453_n22), .C2(
        u4_srl_453_n340), .ZN(u4_srl_453_n583) );
  OAI221_X1 u4_srl_453_U470 ( .B1(u4_srl_453_n294), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n582), .C2(u4_srl_453_n10), .A(u4_srl_453_n583), .ZN(
        u4_N5928) );
  AOI22_X1 u4_srl_453_U469 ( .A1(u4_srl_453_n33), .A2(u4_srl_453_n580), .B1(
        u4_srl_453_n41), .B2(u4_srl_453_n581), .ZN(u4_srl_453_n579) );
  INV_X1 u4_srl_453_U468 ( .A(u4_srl_453_n579), .ZN(u4_srl_453_n578) );
  AOI221_X1 u4_srl_453_U467 ( .B1(u4_srl_453_n576), .B2(u4_srl_453_n26), .C1(
        u4_srl_453_n577), .C2(u4_srl_453_n87), .A(u4_srl_453_n578), .ZN(
        u4_srl_453_n263) );
  AOI22_X1 u4_srl_453_U466 ( .A1(u4_srl_453_n33), .A2(u4_srl_453_n574), .B1(
        u4_srl_453_n41), .B2(u4_srl_453_n575), .ZN(u4_srl_453_n573) );
  OAI221_X1 u4_srl_453_U465 ( .B1(u4_srl_453_n571), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n572), .C2(u4_srl_453_n90), .A(u4_srl_453_n573), .ZN(
        u4_srl_453_n259) );
  INV_X1 u4_srl_453_U464 ( .A(u4_srl_453_n259), .ZN(u4_srl_453_n551) );
  AOI22_X1 u4_srl_453_U463 ( .A1(u4_srl_453_n33), .A2(u4_srl_453_n569), .B1(
        u4_srl_453_n42), .B2(u4_srl_453_n570), .ZN(u4_srl_453_n568) );
  INV_X1 u4_srl_453_U462 ( .A(u4_srl_453_n568), .ZN(u4_srl_453_n567) );
  AOI221_X1 u4_srl_453_U461 ( .B1(u4_srl_453_n565), .B2(u4_srl_453_n26), .C1(
        u4_srl_453_n566), .C2(u4_srl_453_n88), .A(u4_srl_453_n567), .ZN(
        u4_srl_453_n262) );
  INV_X1 u4_srl_453_U460 ( .A(u4_srl_453_n262), .ZN(u4_srl_453_n553) );
  AOI22_X1 u4_srl_453_U459 ( .A1(u4_srl_453_n33), .A2(u4_srl_453_n563), .B1(
        u4_srl_453_n41), .B2(u4_srl_453_n564), .ZN(u4_srl_453_n562) );
  INV_X1 u4_srl_453_U458 ( .A(u4_srl_453_n562), .ZN(u4_srl_453_n561) );
  AOI221_X1 u4_srl_453_U457 ( .B1(u4_srl_453_n559), .B2(u4_srl_453_n25), .C1(
        u4_srl_453_n560), .C2(u4_srl_453_n87), .A(u4_srl_453_n561), .ZN(
        u4_srl_453_n281) );
  OAI22_X1 u4_srl_453_U456 ( .A1(u4_shift_right[4]), .A2(u4_srl_453_n281), 
        .B1(u4_srl_453_n280), .B2(u4_srl_453_n496), .ZN(u4_srl_453_n337) );
  AOI22_X1 u4_srl_453_U455 ( .A1(u4_srl_453_n33), .A2(u4_srl_453_n557), .B1(
        u4_srl_453_n41), .B2(u4_srl_453_n558), .ZN(u4_srl_453_n556) );
  OAI221_X1 u4_srl_453_U454 ( .B1(u4_srl_453_n554), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n555), .C2(u4_srl_453_n89), .A(u4_srl_453_n556), .ZN(
        u4_srl_453_n338) );
  AOI222_X1 u4_srl_453_U453 ( .A1(u4_srl_453_n24), .A2(u4_srl_453_n553), .B1(
        u4_srl_453_n490), .B2(u4_srl_453_n337), .C1(u4_srl_453_n22), .C2(
        u4_srl_453_n338), .ZN(u4_srl_453_n552) );
  OAI221_X1 u4_srl_453_U452 ( .B1(u4_srl_453_n263), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n551), .C2(u4_srl_453_n10), .A(u4_srl_453_n552), .ZN(
        u4_N5929) );
  AOI22_X1 u4_srl_453_U451 ( .A1(u4_srl_453_n33), .A2(u4_srl_453_n549), .B1(
        u4_srl_453_n41), .B2(u4_srl_453_n550), .ZN(u4_srl_453_n548) );
  INV_X1 u4_srl_453_U450 ( .A(u4_srl_453_n548), .ZN(u4_srl_453_n547) );
  AOI221_X1 u4_srl_453_U449 ( .B1(u4_srl_453_n545), .B2(u4_srl_453_n26), .C1(
        u4_srl_453_n546), .C2(u4_srl_453_n88), .A(u4_srl_453_n547), .ZN(
        u4_srl_453_n235) );
  INV_X1 u4_srl_453_U448 ( .A(u4_srl_453_n544), .ZN(u4_srl_453_n539) );
  AOI22_X1 u4_srl_453_U447 ( .A1(u4_srl_453_n33), .A2(u4_srl_453_n542), .B1(
        u4_srl_453_n42), .B2(u4_srl_453_n543), .ZN(u4_srl_453_n541) );
  OAI221_X1 u4_srl_453_U446 ( .B1(u4_srl_453_n539), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n540), .C2(u4_srl_453_n89), .A(u4_srl_453_n541), .ZN(
        u4_srl_453_n231) );
  INV_X1 u4_srl_453_U445 ( .A(u4_srl_453_n231), .ZN(u4_srl_453_n521) );
  INV_X1 u4_srl_453_U444 ( .A(u4_srl_453_n538), .ZN(u4_srl_453_n534) );
  AOI22_X1 u4_srl_453_U443 ( .A1(u4_srl_453_n33), .A2(u4_srl_453_n536), .B1(
        u4_srl_453_n41), .B2(u4_srl_453_n537), .ZN(u4_srl_453_n535) );
  OAI221_X1 u4_srl_453_U442 ( .B1(u4_srl_453_n533), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n534), .C2(u4_srl_453_n89), .A(u4_srl_453_n535), .ZN(
        u4_srl_453_n414) );
  AOI22_X1 u4_srl_453_U441 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n531), .B1(
        u4_srl_453_n41), .B2(u4_srl_453_n532), .ZN(u4_srl_453_n530) );
  OAI221_X1 u4_srl_453_U440 ( .B1(u4_srl_453_n528), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n529), .C2(u4_srl_453_n89), .A(u4_srl_453_n530), .ZN(
        u4_srl_453_n413) );
  INV_X1 u4_srl_453_U439 ( .A(u4_srl_453_n413), .ZN(u4_srl_453_n278) );
  OAI22_X1 u4_srl_453_U438 ( .A1(u4_shift_right[4]), .A2(u4_srl_453_n278), 
        .B1(u4_srl_453_n277), .B2(u4_srl_453_n496), .ZN(u4_srl_453_n335) );
  AOI22_X1 u4_srl_453_U437 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n526), .B1(
        u4_srl_453_n41), .B2(u4_srl_453_n527), .ZN(u4_srl_453_n525) );
  OAI221_X1 u4_srl_453_U436 ( .B1(u4_srl_453_n523), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n524), .C2(u4_srl_453_n89), .A(u4_srl_453_n525), .ZN(
        u4_srl_453_n336) );
  AOI222_X1 u4_srl_453_U435 ( .A1(u4_srl_453_n24), .A2(u4_srl_453_n414), .B1(
        u4_srl_453_n490), .B2(u4_srl_453_n335), .C1(u4_srl_453_n22), .C2(
        u4_srl_453_n336), .ZN(u4_srl_453_n522) );
  OAI221_X1 u4_srl_453_U434 ( .B1(u4_srl_453_n235), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n521), .C2(u4_srl_453_n10), .A(u4_srl_453_n522), .ZN(
        u4_N5930) );
  AOI22_X1 u4_srl_453_U433 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n519), .B1(
        u4_srl_453_n42), .B2(u4_srl_453_n520), .ZN(u4_srl_453_n518) );
  INV_X1 u4_srl_453_U432 ( .A(u4_srl_453_n518), .ZN(u4_srl_453_n517) );
  AOI221_X1 u4_srl_453_U431 ( .B1(u4_srl_453_n515), .B2(u4_srl_453_n25), .C1(
        u4_srl_453_n516), .C2(u4_srl_453_n88), .A(u4_srl_453_n517), .ZN(
        u4_srl_453_n211) );
  INV_X1 u4_srl_453_U430 ( .A(u4_srl_453_n514), .ZN(u4_srl_453_n509) );
  AOI22_X1 u4_srl_453_U429 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n512), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n513), .ZN(u4_srl_453_n511) );
  OAI221_X1 u4_srl_453_U428 ( .B1(u4_srl_453_n509), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n510), .C2(u4_srl_453_n89), .A(u4_srl_453_n511), .ZN(
        u4_srl_453_n205) );
  INV_X1 u4_srl_453_U427 ( .A(u4_srl_453_n205), .ZN(u4_srl_453_n487) );
  AOI22_X1 u4_srl_453_U426 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n507), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n508), .ZN(u4_srl_453_n506) );
  INV_X1 u4_srl_453_U425 ( .A(u4_srl_453_n506), .ZN(u4_srl_453_n505) );
  AOI221_X1 u4_srl_453_U424 ( .B1(u4_srl_453_n503), .B2(u4_srl_453_n26), .C1(
        u4_srl_453_n504), .C2(u4_srl_453_n88), .A(u4_srl_453_n505), .ZN(
        u4_srl_453_n209) );
  INV_X1 u4_srl_453_U423 ( .A(u4_srl_453_n209), .ZN(u4_srl_453_n489) );
  AOI22_X1 u4_srl_453_U422 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n501), .B1(
        u4_srl_453_n41), .B2(u4_srl_453_n502), .ZN(u4_srl_453_n500) );
  INV_X1 u4_srl_453_U421 ( .A(u4_srl_453_n500), .ZN(u4_srl_453_n499) );
  AOI221_X1 u4_srl_453_U420 ( .B1(u4_srl_453_n497), .B2(u4_srl_453_n25), .C1(
        u4_srl_453_n498), .C2(u4_srl_453_n88), .A(u4_srl_453_n499), .ZN(
        u4_srl_453_n274) );
  OAI22_X1 u4_srl_453_U419 ( .A1(u4_srl_453_n274), .A2(u4_shift_right[4]), 
        .B1(u4_srl_453_n273), .B2(u4_srl_453_n496), .ZN(u4_srl_453_n333) );
  AOI22_X1 u4_srl_453_U418 ( .A1(u4_srl_453_n35), .A2(u4_srl_453_n494), .B1(
        u4_srl_453_n40), .B2(u4_srl_453_n495), .ZN(u4_srl_453_n493) );
  OAI221_X1 u4_srl_453_U417 ( .B1(u4_srl_453_n491), .B2(u4_srl_453_n31), .C1(
        u4_srl_453_n492), .C2(u4_srl_453_n89), .A(u4_srl_453_n493), .ZN(
        u4_srl_453_n334) );
  AOI222_X1 u4_srl_453_U416 ( .A1(u4_srl_453_n24), .A2(u4_srl_453_n489), .B1(
        u4_srl_453_n490), .B2(u4_srl_453_n333), .C1(u4_srl_453_n22), .C2(
        u4_srl_453_n334), .ZN(u4_srl_453_n488) );
  OAI221_X1 u4_srl_453_U415 ( .B1(u4_srl_453_n211), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n487), .C2(u4_srl_453_n10), .A(u4_srl_453_n488), .ZN(
        u4_N5931) );
  INV_X1 u4_srl_453_U414 ( .A(u4_srl_453_n331), .ZN(u4_srl_453_n486) );
  INV_X1 u4_srl_453_U413 ( .A(u4_srl_453_n223), .ZN(u4_srl_453_n402) );
  AOI222_X1 u4_srl_453_U412 ( .A1(u4_srl_453_n24), .A2(u4_srl_453_n486), .B1(
        u4_srl_453_n22), .B2(u4_srl_453_n403), .C1(u4_srl_453_n440), .C2(
        u4_srl_453_n402), .ZN(u4_srl_453_n485) );
  OAI221_X1 u4_srl_453_U411 ( .B1(u4_srl_453_n405), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n484), .C2(u4_srl_453_n9), .A(u4_srl_453_n485), .ZN(
        u4_N5932) );
  INV_X1 u4_srl_453_U410 ( .A(u4_srl_453_n329), .ZN(u4_srl_453_n483) );
  INV_X1 u4_srl_453_U409 ( .A(u4_srl_453_n222), .ZN(u4_srl_453_n397) );
  AOI222_X1 u4_srl_453_U408 ( .A1(u4_srl_453_n24), .A2(u4_srl_453_n483), .B1(
        u4_srl_453_n22), .B2(u4_srl_453_n398), .C1(u4_srl_453_n440), .C2(
        u4_srl_453_n397), .ZN(u4_srl_453_n482) );
  OAI221_X1 u4_srl_453_U407 ( .B1(u4_srl_453_n400), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n481), .C2(u4_srl_453_n9), .A(u4_srl_453_n482), .ZN(
        u4_N5933) );
  AOI222_X1 u4_srl_453_U406 ( .A1(u4_srl_453_n24), .A2(u4_srl_453_n480), .B1(
        u4_srl_453_n22), .B2(u4_srl_453_n393), .C1(u4_srl_453_n440), .C2(
        u4_srl_453_n392), .ZN(u4_srl_453_n479) );
  OAI221_X1 u4_srl_453_U405 ( .B1(u4_srl_453_n395), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n478), .C2(u4_srl_453_n9), .A(u4_srl_453_n479), .ZN(
        u4_N5934) );
  INV_X1 u4_srl_453_U404 ( .A(u4_srl_453_n311), .ZN(u4_srl_453_n477) );
  INV_X1 u4_srl_453_U403 ( .A(u4_srl_453_n220), .ZN(u4_srl_453_n387) );
  AOI222_X1 u4_srl_453_U402 ( .A1(u4_srl_453_n24), .A2(u4_srl_453_n477), .B1(
        u4_srl_453_n22), .B2(u4_srl_453_n388), .C1(u4_srl_453_n440), .C2(
        u4_srl_453_n387), .ZN(u4_srl_453_n476) );
  OAI221_X1 u4_srl_453_U401 ( .B1(u4_srl_453_n390), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n475), .C2(u4_srl_453_n9), .A(u4_srl_453_n476), .ZN(
        u4_N5935) );
  AOI222_X1 u4_srl_453_U400 ( .A1(u4_srl_453_n449), .A2(u4_srl_453_n432), .B1(
        u4_srl_453_n355), .B2(u4_srl_453_n368), .C1(u4_srl_453_n356), .C2(
        u4_srl_453_n433), .ZN(u4_srl_453_n303) );
  INV_X1 u4_srl_453_U399 ( .A(u4_srl_453_n447), .ZN(u4_srl_453_n467) );
  OAI22_X1 u4_srl_453_U398 ( .A1(u4_srl_453_n59), .A2(u4_srl_453_n93), .B1(
        u4_srl_453_n53), .B2(u4_srl_453_n94), .ZN(u4_srl_453_n474) );
  AOI221_X1 u4_srl_453_U397 ( .B1(n8513), .B2(u4_srl_453_n69), .C1(n8512), 
        .C2(u4_srl_453_n78), .A(u4_srl_453_n474), .ZN(u4_srl_453_n469) );
  AOI22_X1 u4_srl_453_U396 ( .A1(net33548), .A2(u4_srl_453_n69), .B1(net33641), 
        .B2(u4_srl_453_n78), .ZN(u4_srl_453_n473) );
  OAI221_X1 u4_srl_453_U395 ( .B1(u4_srl_453_n53), .B2(u4_srl_453_n98), .C1(
        u4_srl_453_n59), .C2(u4_srl_453_n97), .A(u4_srl_453_n473), .ZN(
        u4_srl_453_n289) );
  AOI222_X1 u4_srl_453_U394 ( .A1(u4_srl_453_n25), .A2(u4_srl_453_n289), .B1(
        u4_srl_453_n35), .B2(u4_srl_453_n286), .C1(u4_srl_453_n40), .C2(
        u4_srl_453_n290), .ZN(u4_srl_453_n472) );
  MUX2_X1 u4_srl_453_U393 ( .A(u4_srl_453_n471), .B(u4_srl_453_n472), .S(
        u4_srl_453_n424), .Z(u4_srl_453_n470) );
  OAI21_X1 u4_srl_453_U392 ( .B1(u4_srl_453_n469), .B2(u4_srl_453_n298), .A(
        u4_srl_453_n470), .ZN(u4_srl_453_n468) );
  AOI22_X1 u4_srl_453_U391 ( .A1(u4_srl_453_n23), .A2(u4_srl_453_n467), .B1(
        u4_srl_453_n418), .B2(u4_srl_453_n468), .ZN(u4_srl_453_n466) );
  OAI221_X1 u4_srl_453_U390 ( .B1(u4_srl_453_n303), .B2(u4_srl_453_n415), .C1(
        u4_srl_453_n353), .C2(u4_srl_453_n2), .A(u4_srl_453_n466), .ZN(
        u4_N5908) );
  INV_X1 u4_srl_453_U389 ( .A(u4_srl_453_n309), .ZN(u4_srl_453_n463) );
  INV_X1 u4_srl_453_U388 ( .A(u4_srl_453_n219), .ZN(u4_srl_453_n465) );
  AOI222_X1 u4_srl_453_U387 ( .A1(u4_srl_453_n24), .A2(u4_srl_453_n463), .B1(
        u4_srl_453_n22), .B2(u4_srl_453_n464), .C1(u4_srl_453_n440), .C2(
        u4_srl_453_n465), .ZN(u4_srl_453_n462) );
  OAI221_X1 u4_srl_453_U386 ( .B1(u4_srl_453_n385), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n461), .C2(u4_srl_453_n9), .A(u4_srl_453_n462), .ZN(
        u4_N5936) );
  INV_X1 u4_srl_453_U385 ( .A(u4_srl_453_n218), .ZN(u4_srl_453_n460) );
  AOI222_X1 u4_srl_453_U384 ( .A1(u4_srl_453_n24), .A2(u4_srl_453_n458), .B1(
        u4_srl_453_n22), .B2(u4_srl_453_n459), .C1(u4_srl_453_n440), .C2(
        u4_srl_453_n460), .ZN(u4_srl_453_n457) );
  OAI221_X1 u4_srl_453_U383 ( .B1(u4_srl_453_n382), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n456), .C2(u4_srl_453_n9), .A(u4_srl_453_n457), .ZN(
        u4_N5937) );
  AOI222_X1 u4_srl_453_U382 ( .A1(u4_srl_453_n24), .A2(u4_srl_453_n455), .B1(
        u4_srl_453_n22), .B2(u4_srl_453_n379), .C1(u4_srl_453_n440), .C2(
        u4_srl_453_n378), .ZN(u4_srl_453_n454) );
  OAI221_X1 u4_srl_453_U381 ( .B1(u4_srl_453_n376), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n453), .C2(u4_srl_453_n9), .A(u4_srl_453_n454), .ZN(
        u4_N5938) );
  AOI222_X1 u4_srl_453_U380 ( .A1(u4_srl_453_n24), .A2(u4_srl_453_n452), .B1(
        u4_srl_453_n22), .B2(u4_srl_453_n374), .C1(u4_srl_453_n440), .C2(
        u4_srl_453_n373), .ZN(u4_srl_453_n451) );
  OAI221_X1 u4_srl_453_U379 ( .B1(u4_srl_453_n371), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n450), .C2(u4_srl_453_n9), .A(u4_srl_453_n451), .ZN(
        u4_N5939) );
  AOI222_X1 u4_srl_453_U378 ( .A1(u4_srl_453_n24), .A2(u4_srl_453_n449), .B1(
        u4_srl_453_n22), .B2(u4_srl_453_n356), .C1(u4_srl_453_n440), .C2(
        u4_srl_453_n355), .ZN(u4_srl_453_n448) );
  OAI221_X1 u4_srl_453_U377 ( .B1(u4_srl_453_n353), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n447), .C2(u4_srl_453_n9), .A(u4_srl_453_n448), .ZN(
        u4_N5940) );
  AOI222_X1 u4_srl_453_U376 ( .A1(u4_srl_453_n24), .A2(u4_srl_453_n431), .B1(
        u4_srl_453_n22), .B2(u4_srl_453_n351), .C1(u4_srl_453_n440), .C2(
        u4_srl_453_n350), .ZN(u4_srl_453_n446) );
  OAI221_X1 u4_srl_453_U375 ( .B1(u4_srl_453_n348), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n430), .C2(u4_srl_453_n9), .A(u4_srl_453_n446), .ZN(
        u4_N5941) );
  INV_X1 u4_srl_453_U374 ( .A(u4_srl_453_n366), .ZN(u4_srl_453_n345) );
  AOI222_X1 u4_srl_453_U373 ( .A1(u4_srl_453_n24), .A2(u4_srl_453_n369), .B1(
        u4_srl_453_n22), .B2(u4_srl_453_n346), .C1(u4_srl_453_n440), .C2(
        u4_srl_453_n345), .ZN(u4_srl_453_n445) );
  OAI221_X1 u4_srl_453_U372 ( .B1(u4_srl_453_n343), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n365), .C2(u4_srl_453_n8), .A(u4_srl_453_n445), .ZN(
        u4_N5942) );
  INV_X1 u4_srl_453_U371 ( .A(u4_srl_453_n325), .ZN(u4_srl_453_n443) );
  INV_X1 u4_srl_453_U370 ( .A(u4_srl_453_n327), .ZN(u4_srl_453_n444) );
  AOI222_X1 u4_srl_453_U369 ( .A1(u4_srl_453_n24), .A2(u4_srl_453_n341), .B1(
        u4_srl_453_n440), .B2(u4_srl_453_n443), .C1(u4_srl_453_n22), .C2(
        u4_srl_453_n444), .ZN(u4_srl_453_n442) );
  OAI221_X1 u4_srl_453_U368 ( .B1(u4_srl_453_n322), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n323), .C2(u4_srl_453_n8), .A(u4_srl_453_n442), .ZN(
        u4_N5943) );
  AND2_X1 u4_srl_453_U367 ( .A1(u4_srl_453_n440), .A2(u4_srl_453_n91), .ZN(
        u4_srl_453_n411) );
  INV_X1 u4_srl_453_U366 ( .A(u4_srl_453_n297), .ZN(u4_srl_453_n439) );
  AOI222_X1 u4_srl_453_U365 ( .A1(u4_srl_453_n24), .A2(u4_srl_453_n340), .B1(
        u4_srl_453_n411), .B2(u4_srl_453_n438), .C1(u4_srl_453_n22), .C2(
        u4_srl_453_n439), .ZN(u4_srl_453_n437) );
  OAI221_X1 u4_srl_453_U364 ( .B1(u4_srl_453_n293), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n294), .C2(u4_srl_453_n8), .A(u4_srl_453_n437), .ZN(
        u4_N5944) );
  INV_X1 u4_srl_453_U363 ( .A(u4_srl_453_n281), .ZN(u4_srl_453_n436) );
  AOI222_X1 u4_srl_453_U362 ( .A1(u4_srl_453_n24), .A2(u4_srl_453_n338), .B1(
        u4_srl_453_n411), .B2(u4_srl_453_n435), .C1(u4_srl_453_n22), .C2(
        u4_srl_453_n436), .ZN(u4_srl_453_n434) );
  OAI221_X1 u4_srl_453_U361 ( .B1(u4_srl_453_n262), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n263), .C2(u4_srl_453_n8), .A(u4_srl_453_n434), .ZN(
        u4_N5945) );
  AOI222_X1 u4_srl_453_U360 ( .A1(u4_srl_453_n431), .A2(u4_srl_453_n432), .B1(
        u4_srl_453_n350), .B2(u4_srl_453_n368), .C1(u4_srl_453_n351), .C2(
        u4_srl_453_n433), .ZN(u4_srl_453_n302) );
  INV_X1 u4_srl_453_U359 ( .A(u4_srl_453_n430), .ZN(u4_srl_453_n417) );
  OAI22_X1 u4_srl_453_U358 ( .A1(u4_srl_453_n59), .A2(u4_srl_453_n94), .B1(
        u4_srl_453_n53), .B2(u4_srl_453_n95), .ZN(u4_srl_453_n429) );
  AOI221_X1 u4_srl_453_U357 ( .B1(n8514), .B2(u4_srl_453_n69), .C1(n8513), 
        .C2(u4_srl_453_n78), .A(u4_srl_453_n429), .ZN(u4_srl_453_n420) );
  AOI22_X1 u4_srl_453_U356 ( .A1(net33549), .A2(u4_srl_453_n72), .B1(net33548), 
        .B2(u4_srl_453_n81), .ZN(u4_srl_453_n427) );
  OAI221_X1 u4_srl_453_U355 ( .B1(u4_srl_453_n50), .B2(u4_srl_453_n99), .C1(
        u4_srl_453_n63), .C2(u4_srl_453_n98), .A(u4_srl_453_n427), .ZN(
        u4_srl_453_n257) );
  AOI222_X1 u4_srl_453_U354 ( .A1(u4_srl_453_n25), .A2(u4_srl_453_n257), .B1(
        u4_srl_453_n35), .B2(u4_srl_453_n254), .C1(u4_srl_453_n40), .C2(
        u4_srl_453_n258), .ZN(u4_srl_453_n423) );
  MUX2_X1 u4_srl_453_U353 ( .A(u4_srl_453_n422), .B(u4_srl_453_n423), .S(
        u4_srl_453_n424), .Z(u4_srl_453_n421) );
  OAI21_X1 u4_srl_453_U352 ( .B1(u4_srl_453_n420), .B2(u4_srl_453_n298), .A(
        u4_srl_453_n421), .ZN(u4_srl_453_n419) );
  AOI22_X1 u4_srl_453_U351 ( .A1(u4_srl_453_n23), .A2(u4_srl_453_n417), .B1(
        u4_srl_453_n418), .B2(u4_srl_453_n419), .ZN(u4_srl_453_n416) );
  OAI221_X1 u4_srl_453_U350 ( .B1(u4_srl_453_n302), .B2(u4_srl_453_n415), .C1(
        u4_srl_453_n348), .C2(u4_srl_453_n2), .A(u4_srl_453_n416), .ZN(
        u4_N5909) );
  INV_X1 u4_srl_453_U349 ( .A(u4_srl_453_n414), .ZN(u4_srl_453_n234) );
  AOI222_X1 u4_srl_453_U348 ( .A1(u4_srl_453_n24), .A2(u4_srl_453_n336), .B1(
        u4_srl_453_n411), .B2(u4_srl_453_n412), .C1(u4_srl_453_n22), .C2(
        u4_srl_453_n413), .ZN(u4_srl_453_n410) );
  OAI221_X1 u4_srl_453_U347 ( .B1(u4_srl_453_n234), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n235), .C2(u4_srl_453_n8), .A(u4_srl_453_n410), .ZN(
        u4_N5946) );
  INV_X1 u4_srl_453_U346 ( .A(u4_srl_453_n274), .ZN(u4_srl_453_n409) );
  AOI222_X1 u4_srl_453_U345 ( .A1(u4_srl_453_n24), .A2(u4_srl_453_n334), .B1(
        u4_srl_453_n407), .B2(u4_srl_453_n408), .C1(u4_srl_453_n22), .C2(
        u4_srl_453_n409), .ZN(u4_srl_453_n406) );
  OAI221_X1 u4_srl_453_U344 ( .B1(u4_srl_453_n209), .B2(u4_srl_453_n15), .C1(
        u4_srl_453_n211), .C2(u4_srl_453_n8), .A(u4_srl_453_n406), .ZN(
        u4_N5947) );
  OAI22_X1 u4_srl_453_U343 ( .A1(u4_srl_453_n18), .A2(u4_srl_453_n331), .B1(
        u4_srl_453_n214), .B2(u4_srl_453_n405), .ZN(u4_srl_453_n404) );
  AOI221_X1 u4_srl_453_U342 ( .B1(u4_srl_453_n402), .B2(u4_srl_453_n22), .C1(
        u4_srl_453_n403), .C2(u4_srl_453_n23), .A(u4_srl_453_n404), .ZN(
        u4_srl_453_n401) );
  INV_X1 u4_srl_453_U341 ( .A(u4_srl_453_n401), .ZN(u4_N5948) );
  OAI22_X1 u4_srl_453_U340 ( .A1(u4_srl_453_n19), .A2(u4_srl_453_n329), .B1(
        u4_srl_453_n214), .B2(u4_srl_453_n400), .ZN(u4_srl_453_n399) );
  AOI221_X1 u4_srl_453_U339 ( .B1(u4_srl_453_n397), .B2(u4_srl_453_n22), .C1(
        u4_srl_453_n398), .C2(u4_srl_453_n23), .A(u4_srl_453_n399), .ZN(
        u4_srl_453_n396) );
  INV_X1 u4_srl_453_U338 ( .A(u4_srl_453_n396), .ZN(u4_N5949) );
  OAI22_X1 u4_srl_453_U337 ( .A1(u4_srl_453_n18), .A2(u4_srl_453_n313), .B1(
        u4_srl_453_n11), .B2(u4_srl_453_n395), .ZN(u4_srl_453_n394) );
  AOI221_X1 u4_srl_453_U336 ( .B1(u4_srl_453_n392), .B2(u4_srl_453_n22), .C1(
        u4_srl_453_n393), .C2(u4_srl_453_n23), .A(u4_srl_453_n394), .ZN(
        u4_srl_453_n391) );
  INV_X1 u4_srl_453_U335 ( .A(u4_srl_453_n391), .ZN(u4_N5950) );
  OAI22_X1 u4_srl_453_U334 ( .A1(u4_srl_453_n19), .A2(u4_srl_453_n311), .B1(
        u4_srl_453_n10), .B2(u4_srl_453_n390), .ZN(u4_srl_453_n389) );
  AOI221_X1 u4_srl_453_U333 ( .B1(u4_srl_453_n387), .B2(u4_srl_453_n22), .C1(
        u4_srl_453_n388), .C2(u4_srl_453_n23), .A(u4_srl_453_n389), .ZN(
        u4_srl_453_n386) );
  INV_X1 u4_srl_453_U332 ( .A(u4_srl_453_n386), .ZN(u4_N5951) );
  OAI22_X1 u4_srl_453_U331 ( .A1(u4_srl_453_n19), .A2(u4_srl_453_n309), .B1(
        u4_srl_453_n9), .B2(u4_srl_453_n385), .ZN(u4_srl_453_n384) );
  INV_X1 u4_srl_453_U330 ( .A(u4_srl_453_n384), .ZN(u4_srl_453_n383) );
  OAI221_X1 u4_srl_453_U329 ( .B1(u4_srl_453_n219), .B2(u4_srl_453_n2), .C1(
        u4_srl_453_n308), .C2(u4_srl_453_n4), .A(u4_srl_453_n383), .ZN(
        u4_N5952) );
  OAI22_X1 u4_srl_453_U328 ( .A1(u4_srl_453_n19), .A2(u4_srl_453_n307), .B1(
        u4_srl_453_n8), .B2(u4_srl_453_n382), .ZN(u4_srl_453_n381) );
  INV_X1 u4_srl_453_U327 ( .A(u4_srl_453_n381), .ZN(u4_srl_453_n380) );
  OAI221_X1 u4_srl_453_U326 ( .B1(u4_srl_453_n218), .B2(u4_srl_453_n2), .C1(
        u4_srl_453_n306), .C2(u4_srl_453_n4), .A(u4_srl_453_n380), .ZN(
        u4_N5953) );
  AOI22_X1 u4_srl_453_U325 ( .A1(u4_srl_453_n22), .A2(u4_srl_453_n378), .B1(
        u4_srl_453_n23), .B2(u4_srl_453_n379), .ZN(u4_srl_453_n377) );
  OAI221_X1 u4_srl_453_U324 ( .B1(u4_srl_453_n375), .B2(u4_srl_453_n15), .C1(
        u4_srl_453_n376), .C2(u4_srl_453_n8), .A(u4_srl_453_n377), .ZN(
        u4_N5954) );
  AOI22_X1 u4_srl_453_U323 ( .A1(u4_srl_453_n22), .A2(u4_srl_453_n373), .B1(
        u4_srl_453_n23), .B2(u4_srl_453_n374), .ZN(u4_srl_453_n372) );
  OAI221_X1 u4_srl_453_U322 ( .B1(u4_srl_453_n370), .B2(u4_srl_453_n15), .C1(
        u4_srl_453_n371), .C2(u4_srl_453_n8), .A(u4_srl_453_n372), .ZN(
        u4_N5955) );
  INV_X1 u4_srl_453_U321 ( .A(u4_srl_453_n369), .ZN(u4_srl_453_n342) );
  INV_X1 u4_srl_453_U320 ( .A(u4_srl_453_n368), .ZN(u4_srl_453_n326) );
  OAI222_X1 u4_srl_453_U319 ( .A1(u4_srl_453_n342), .A2(u4_srl_453_n271), .B1(
        u4_srl_453_n366), .B2(u4_srl_453_n326), .C1(u4_srl_453_n367), .C2(
        u4_srl_453_n275), .ZN(u4_srl_453_n301) );
  OAI22_X1 u4_srl_453_U318 ( .A1(u4_srl_453_n343), .A2(u4_srl_453_n210), .B1(
        u4_srl_453_n365), .B2(u4_srl_453_n212), .ZN(u4_srl_453_n364) );
  AOI221_X1 u4_srl_453_U317 ( .B1(u4_srl_453_n204), .B2(u4_srl_453_n363), .C1(
        u4_srl_453_n301), .C2(u4_srl_453_n207), .A(u4_srl_453_n364), .ZN(
        u4_srl_453_n357) );
  INV_X1 u4_srl_453_U316 ( .A(u4_srl_453_n203), .ZN(u4_srl_453_n251) );
  INV_X1 u4_srl_453_U315 ( .A(u4_srl_453_n201), .ZN(u4_srl_453_n253) );
  AOI22_X1 u4_srl_453_U314 ( .A1(u4_srl_453_n362), .A2(u4_srl_453_n197), .B1(
        u4_srl_453_n227), .B2(u4_srl_453_n195), .ZN(u4_srl_453_n361) );
  INV_X1 u4_srl_453_U313 ( .A(u4_srl_453_n361), .ZN(u4_srl_453_n360) );
  AOI221_X1 u4_srl_453_U312 ( .B1(u4_srl_453_n251), .B2(u4_srl_453_n359), .C1(
        u4_srl_453_n253), .C2(u4_srl_453_n226), .A(u4_srl_453_n360), .ZN(
        u4_srl_453_n358) );
  AOI21_X1 u4_srl_453_U311 ( .B1(u4_srl_453_n357), .B2(u4_srl_453_n358), .A(
        u4_shift_right[8]), .ZN(u4_N5910) );
  AOI22_X1 u4_srl_453_U310 ( .A1(u4_srl_453_n22), .A2(u4_srl_453_n355), .B1(
        u4_srl_453_n23), .B2(u4_srl_453_n356), .ZN(u4_srl_453_n354) );
  OAI221_X1 u4_srl_453_U309 ( .B1(u4_srl_453_n352), .B2(u4_srl_453_n15), .C1(
        u4_srl_453_n353), .C2(u4_srl_453_n8), .A(u4_srl_453_n354), .ZN(
        u4_N5956) );
  AOI22_X1 u4_srl_453_U308 ( .A1(u4_srl_453_n22), .A2(u4_srl_453_n350), .B1(
        u4_srl_453_n23), .B2(u4_srl_453_n351), .ZN(u4_srl_453_n349) );
  OAI221_X1 u4_srl_453_U307 ( .B1(u4_srl_453_n347), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n348), .C2(u4_srl_453_n8), .A(u4_srl_453_n349), .ZN(
        u4_N5957) );
  AOI22_X1 u4_srl_453_U306 ( .A1(u4_srl_453_n22), .A2(u4_srl_453_n345), .B1(
        u4_srl_453_n23), .B2(u4_srl_453_n346), .ZN(u4_srl_453_n344) );
  OAI221_X1 u4_srl_453_U305 ( .B1(u4_srl_453_n342), .B2(u4_srl_453_n15), .C1(
        u4_srl_453_n343), .C2(u4_srl_453_n8), .A(u4_srl_453_n344), .ZN(
        u4_N5958) );
  INV_X1 u4_srl_453_U304 ( .A(u4_srl_453_n341), .ZN(u4_srl_453_n324) );
  OAI222_X1 u4_srl_453_U303 ( .A1(u4_srl_453_n322), .A2(u4_srl_453_n11), .B1(
        u4_srl_453_n324), .B2(u4_srl_453_n15), .C1(u4_srl_453_n241), .C2(
        u4_srl_453_n332), .ZN(u4_N5959) );
  INV_X1 u4_srl_453_U302 ( .A(u4_srl_453_n340), .ZN(u4_srl_453_n295) );
  INV_X1 u4_srl_453_U301 ( .A(u4_srl_453_n339), .ZN(u4_srl_453_n240) );
  OAI222_X1 u4_srl_453_U300 ( .A1(u4_srl_453_n293), .A2(u4_srl_453_n11), .B1(
        u4_srl_453_n295), .B2(u4_srl_453_n15), .C1(u4_srl_453_n240), .C2(
        u4_srl_453_n332), .ZN(u4_N5960) );
  INV_X1 u4_srl_453_U299 ( .A(u4_srl_453_n338), .ZN(u4_srl_453_n279) );
  INV_X1 u4_srl_453_U298 ( .A(u4_srl_453_n337), .ZN(u4_srl_453_n239) );
  OAI222_X1 u4_srl_453_U297 ( .A1(u4_srl_453_n262), .A2(u4_srl_453_n11), .B1(
        u4_srl_453_n279), .B2(u4_srl_453_n15), .C1(u4_srl_453_n239), .C2(
        u4_srl_453_n332), .ZN(u4_N5961) );
  INV_X1 u4_srl_453_U296 ( .A(u4_srl_453_n336), .ZN(u4_srl_453_n276) );
  INV_X1 u4_srl_453_U295 ( .A(u4_srl_453_n335), .ZN(u4_srl_453_n238) );
  OAI222_X1 u4_srl_453_U294 ( .A1(u4_srl_453_n234), .A2(u4_srl_453_n11), .B1(
        u4_srl_453_n276), .B2(u4_srl_453_n15), .C1(u4_srl_453_n238), .C2(
        u4_srl_453_n332), .ZN(u4_N5962) );
  INV_X1 u4_srl_453_U293 ( .A(u4_srl_453_n334), .ZN(u4_srl_453_n270) );
  INV_X1 u4_srl_453_U292 ( .A(u4_srl_453_n333), .ZN(u4_srl_453_n236) );
  OAI222_X1 u4_srl_453_U291 ( .A1(u4_srl_453_n209), .A2(u4_srl_453_n11), .B1(
        u4_srl_453_n270), .B2(u4_srl_453_n15), .C1(u4_srl_453_n236), .C2(
        u4_srl_453_n332), .ZN(u4_N5963) );
  OAI222_X1 u4_srl_453_U290 ( .A1(u4_srl_453_n330), .A2(u4_srl_453_n18), .B1(
        u4_srl_453_n223), .B2(u4_srl_453_n4), .C1(u4_srl_453_n331), .C2(
        u4_srl_453_n10), .ZN(u4_N5964) );
  OAI222_X1 u4_srl_453_U289 ( .A1(u4_srl_453_n328), .A2(u4_srl_453_n18), .B1(
        u4_srl_453_n222), .B2(u4_srl_453_n4), .C1(u4_srl_453_n329), .C2(
        u4_srl_453_n11), .ZN(u4_N5965) );
  OAI222_X1 u4_srl_453_U288 ( .A1(u4_srl_453_n324), .A2(u4_srl_453_n271), .B1(
        u4_srl_453_n325), .B2(u4_srl_453_n326), .C1(u4_srl_453_n327), .C2(
        u4_srl_453_n275), .ZN(u4_srl_453_n300) );
  OAI22_X1 u4_srl_453_U287 ( .A1(u4_srl_453_n322), .A2(u4_srl_453_n210), .B1(
        u4_srl_453_n323), .B2(u4_srl_453_n212), .ZN(u4_srl_453_n321) );
  AOI221_X1 u4_srl_453_U286 ( .B1(u4_srl_453_n204), .B2(u4_srl_453_n320), .C1(
        u4_srl_453_n300), .C2(u4_srl_453_n207), .A(u4_srl_453_n321), .ZN(
        u4_srl_453_n314) );
  AOI22_X1 u4_srl_453_U285 ( .A1(u4_srl_453_n319), .A2(u4_srl_453_n197), .B1(
        u4_srl_453_n198), .B2(u4_srl_453_n195), .ZN(u4_srl_453_n318) );
  INV_X1 u4_srl_453_U284 ( .A(u4_srl_453_n318), .ZN(u4_srl_453_n317) );
  AOI221_X1 u4_srl_453_U283 ( .B1(u4_srl_453_n251), .B2(u4_srl_453_n316), .C1(
        u4_srl_453_n253), .C2(u4_srl_453_n196), .A(u4_srl_453_n317), .ZN(
        u4_srl_453_n315) );
  AOI21_X1 u4_srl_453_U282 ( .B1(u4_srl_453_n314), .B2(u4_srl_453_n315), .A(
        u4_shift_right[8]), .ZN(u4_N5911) );
  OAI222_X1 u4_srl_453_U281 ( .A1(u4_srl_453_n312), .A2(u4_srl_453_n18), .B1(
        u4_srl_453_n221), .B2(u4_srl_453_n4), .C1(u4_srl_453_n313), .C2(
        u4_srl_453_n11), .ZN(u4_N5966) );
  OAI222_X1 u4_srl_453_U280 ( .A1(u4_srl_453_n310), .A2(u4_srl_453_n18), .B1(
        u4_srl_453_n220), .B2(u4_srl_453_n4), .C1(u4_srl_453_n311), .C2(
        u4_srl_453_n10), .ZN(u4_N5967) );
  OAI222_X1 u4_srl_453_U279 ( .A1(u4_srl_453_n308), .A2(u4_srl_453_n18), .B1(
        u4_srl_453_n219), .B2(u4_srl_453_n4), .C1(u4_srl_453_n309), .C2(
        u4_srl_453_n11), .ZN(u4_N5968) );
  OAI222_X1 u4_srl_453_U278 ( .A1(u4_srl_453_n306), .A2(u4_srl_453_n18), .B1(
        u4_srl_453_n218), .B2(u4_srl_453_n4), .C1(u4_srl_453_n307), .C2(
        u4_srl_453_n11), .ZN(u4_N5969) );
  INV_X1 u4_srl_453_U277 ( .A(u4_srl_453_n243), .ZN(u4_srl_453_n245) );
  NOR2_X1 u4_srl_453_U276 ( .A1(u4_srl_453_n305), .A2(u4_srl_453_n245), .ZN(
        u4_N5970) );
  NOR2_X1 u4_srl_453_U275 ( .A1(u4_srl_453_n304), .A2(u4_srl_453_n245), .ZN(
        u4_N5971) );
  NOR2_X1 u4_srl_453_U274 ( .A1(u4_srl_453_n303), .A2(u4_srl_453_n245), .ZN(
        u4_N5972) );
  NOR2_X1 u4_srl_453_U273 ( .A1(u4_srl_453_n302), .A2(u4_srl_453_n245), .ZN(
        u4_N5973) );
  AND2_X1 u4_srl_453_U272 ( .A1(u4_srl_453_n301), .A2(u4_srl_453_n243), .ZN(
        u4_N5974) );
  AND2_X1 u4_srl_453_U271 ( .A1(u4_srl_453_n300), .A2(u4_srl_453_n243), .ZN(
        u4_N5975) );
  OR2_X1 u4_srl_453_U270 ( .A1(u4_srl_453_n298), .A2(u4_srl_453_n299), .ZN(
        u4_srl_453_n272) );
  OAI222_X1 u4_srl_453_U269 ( .A1(u4_srl_453_n295), .A2(u4_srl_453_n271), .B1(
        u4_srl_453_n296), .B2(u4_srl_453_n272), .C1(u4_srl_453_n297), .C2(
        u4_srl_453_n275), .ZN(u4_srl_453_n282) );
  OAI22_X1 u4_srl_453_U268 ( .A1(u4_srl_453_n293), .A2(u4_srl_453_n210), .B1(
        u4_srl_453_n294), .B2(u4_srl_453_n212), .ZN(u4_srl_453_n292) );
  AOI221_X1 u4_srl_453_U267 ( .B1(u4_srl_453_n204), .B2(u4_srl_453_n291), .C1(
        u4_srl_453_n282), .C2(u4_srl_453_n207), .A(u4_srl_453_n292), .ZN(
        u4_srl_453_n283) );
  AOI22_X1 u4_srl_453_U266 ( .A1(u4_srl_453_n289), .A2(u4_srl_453_n197), .B1(
        u4_srl_453_n290), .B2(u4_srl_453_n195), .ZN(u4_srl_453_n288) );
  INV_X1 u4_srl_453_U265 ( .A(u4_srl_453_n288), .ZN(u4_srl_453_n287) );
  AOI221_X1 u4_srl_453_U264 ( .B1(u4_srl_453_n251), .B2(u4_srl_453_n285), .C1(
        u4_srl_453_n253), .C2(u4_srl_453_n286), .A(u4_srl_453_n287), .ZN(
        u4_srl_453_n284) );
  AOI21_X1 u4_srl_453_U263 ( .B1(u4_srl_453_n283), .B2(u4_srl_453_n284), .A(
        u4_shift_right[8]), .ZN(u4_N5912) );
  AND2_X1 u4_srl_453_U262 ( .A1(u4_srl_453_n282), .A2(u4_srl_453_n243), .ZN(
        u4_N5976) );
  OAI222_X1 u4_srl_453_U261 ( .A1(u4_srl_453_n279), .A2(u4_srl_453_n271), .B1(
        u4_srl_453_n280), .B2(u4_srl_453_n272), .C1(u4_srl_453_n281), .C2(
        u4_srl_453_n275), .ZN(u4_srl_453_n260) );
  AND2_X1 u4_srl_453_U260 ( .A1(u4_srl_453_n260), .A2(u4_srl_453_n243), .ZN(
        u4_N5977) );
  OAI222_X1 u4_srl_453_U259 ( .A1(u4_srl_453_n276), .A2(u4_srl_453_n271), .B1(
        u4_srl_453_n277), .B2(u4_srl_453_n272), .C1(u4_srl_453_n278), .C2(
        u4_srl_453_n275), .ZN(u4_srl_453_n232) );
  AND2_X1 u4_srl_453_U258 ( .A1(u4_srl_453_n232), .A2(u4_srl_453_n243), .ZN(
        u4_N5978) );
  OAI222_X1 u4_srl_453_U257 ( .A1(u4_srl_453_n270), .A2(u4_srl_453_n271), .B1(
        u4_srl_453_n272), .B2(u4_srl_453_n273), .C1(u4_srl_453_n274), .C2(
        u4_srl_453_n275), .ZN(u4_srl_453_n206) );
  AND2_X1 u4_srl_453_U256 ( .A1(u4_srl_453_n206), .A2(u4_srl_453_n243), .ZN(
        u4_N5979) );
  AND2_X1 u4_srl_453_U255 ( .A1(u4_srl_453_n269), .A2(u4_srl_453_n243), .ZN(
        u4_N5980) );
  AND2_X1 u4_srl_453_U254 ( .A1(u4_srl_453_n268), .A2(u4_srl_453_n243), .ZN(
        u4_N5981) );
  AND2_X1 u4_srl_453_U253 ( .A1(u4_srl_453_n267), .A2(u4_srl_453_n243), .ZN(
        u4_N5982) );
  AND2_X1 u4_srl_453_U252 ( .A1(u4_srl_453_n266), .A2(u4_srl_453_n243), .ZN(
        u4_N5983) );
  AND2_X1 u4_srl_453_U251 ( .A1(u4_srl_453_n265), .A2(u4_srl_453_n243), .ZN(
        u4_N5984) );
  AND2_X1 u4_srl_453_U250 ( .A1(u4_srl_453_n264), .A2(u4_srl_453_n243), .ZN(
        u4_N5985) );
  OAI22_X1 u4_srl_453_U249 ( .A1(u4_srl_453_n262), .A2(u4_srl_453_n210), .B1(
        u4_srl_453_n263), .B2(u4_srl_453_n212), .ZN(u4_srl_453_n261) );
  AOI221_X1 u4_srl_453_U248 ( .B1(u4_srl_453_n204), .B2(u4_srl_453_n259), .C1(
        u4_srl_453_n260), .C2(u4_srl_453_n207), .A(u4_srl_453_n261), .ZN(
        u4_srl_453_n249) );
  AOI22_X1 u4_srl_453_U247 ( .A1(u4_srl_453_n257), .A2(u4_srl_453_n197), .B1(
        u4_srl_453_n258), .B2(u4_srl_453_n195), .ZN(u4_srl_453_n256) );
  INV_X1 u4_srl_453_U246 ( .A(u4_srl_453_n256), .ZN(u4_srl_453_n255) );
  AOI221_X1 u4_srl_453_U245 ( .B1(u4_srl_453_n251), .B2(u4_srl_453_n252), .C1(
        u4_srl_453_n253), .C2(u4_srl_453_n254), .A(u4_srl_453_n255), .ZN(
        u4_srl_453_n250) );
  AOI21_X1 u4_srl_453_U244 ( .B1(u4_srl_453_n249), .B2(u4_srl_453_n250), .A(
        u4_shift_right[8]), .ZN(u4_N5913) );
  NOR2_X1 u4_srl_453_U243 ( .A1(u4_srl_453_n248), .A2(u4_srl_453_n245), .ZN(
        u4_N5986) );
  NOR2_X1 u4_srl_453_U242 ( .A1(u4_srl_453_n247), .A2(u4_srl_453_n245), .ZN(
        u4_N5987) );
  NOR2_X1 u4_srl_453_U241 ( .A1(u4_srl_453_n246), .A2(u4_srl_453_n245), .ZN(
        u4_N5988) );
  NOR2_X1 u4_srl_453_U240 ( .A1(u4_srl_453_n244), .A2(u4_srl_453_n245), .ZN(
        u4_N5989) );
  AND2_X1 u4_srl_453_U239 ( .A1(u4_srl_453_n242), .A2(u4_srl_453_n243), .ZN(
        u4_N5990) );
  NOR2_X1 u4_srl_453_U238 ( .A1(u4_srl_453_n241), .A2(u4_srl_453_n237), .ZN(
        u4_N5991) );
  NOR2_X1 u4_srl_453_U237 ( .A1(u4_srl_453_n240), .A2(u4_srl_453_n237), .ZN(
        u4_N5992) );
  NOR2_X1 u4_srl_453_U236 ( .A1(u4_srl_453_n239), .A2(u4_srl_453_n237), .ZN(
        u4_N5993) );
  NOR2_X1 u4_srl_453_U235 ( .A1(u4_srl_453_n238), .A2(u4_srl_453_n237), .ZN(
        u4_N5994) );
  NOR2_X1 u4_srl_453_U234 ( .A1(u4_srl_453_n236), .A2(u4_srl_453_n237), .ZN(
        u4_N5995) );
  OAI22_X1 u4_srl_453_U233 ( .A1(u4_srl_453_n234), .A2(u4_srl_453_n210), .B1(
        u4_srl_453_n235), .B2(u4_srl_453_n212), .ZN(u4_srl_453_n233) );
  AOI221_X1 u4_srl_453_U232 ( .B1(u4_srl_453_n204), .B2(u4_srl_453_n231), .C1(
        u4_srl_453_n232), .C2(u4_srl_453_n207), .A(u4_srl_453_n233), .ZN(
        u4_srl_453_n224) );
  OAI22_X1 u4_srl_453_U231 ( .A1(u4_srl_453_n229), .A2(u4_srl_453_n201), .B1(
        u4_srl_453_n230), .B2(u4_srl_453_n203), .ZN(u4_srl_453_n228) );
  AOI221_X1 u4_srl_453_U230 ( .B1(u4_srl_453_n195), .B2(u4_srl_453_n226), .C1(
        u4_srl_453_n197), .C2(u4_srl_453_n227), .A(u4_srl_453_n228), .ZN(
        u4_srl_453_n225) );
  AOI21_X1 u4_srl_453_U229 ( .B1(u4_srl_453_n224), .B2(u4_srl_453_n225), .A(
        u4_shift_right[8]), .ZN(u4_N5914) );
  NOR2_X1 u4_srl_453_U228 ( .A1(u4_srl_453_n223), .A2(u4_srl_453_n9), .ZN(
        u4_N5996) );
  NOR2_X1 u4_srl_453_U227 ( .A1(u4_srl_453_n222), .A2(u4_srl_453_n9), .ZN(
        u4_N5997) );
  NOR2_X1 u4_srl_453_U226 ( .A1(u4_srl_453_n221), .A2(u4_srl_453_n9), .ZN(
        u4_N5998) );
  NOR2_X1 u4_srl_453_U225 ( .A1(u4_srl_453_n220), .A2(u4_srl_453_n9), .ZN(
        u4_N5999) );
  NOR2_X1 u4_srl_453_U224 ( .A1(u4_srl_453_n219), .A2(u4_srl_453_n9), .ZN(
        u4_N6000) );
  NOR2_X1 u4_srl_453_U223 ( .A1(u4_srl_453_n218), .A2(u4_srl_453_n11), .ZN(
        u4_N6001) );
  NOR2_X1 u4_srl_453_U222 ( .A1(u4_srl_453_n217), .A2(u4_srl_453_n11), .ZN(
        u4_N6002) );
  NOR2_X1 u4_srl_453_U221 ( .A1(u4_srl_453_n216), .A2(u4_srl_453_n11), .ZN(
        u4_N6003) );
  NOR2_X1 u4_srl_453_U220 ( .A1(u4_srl_453_n215), .A2(u4_srl_453_n11), .ZN(
        u4_N6004) );
  NOR2_X1 u4_srl_453_U219 ( .A1(u4_srl_453_n213), .A2(u4_srl_453_n9), .ZN(
        u4_N6005) );
  OAI22_X1 u4_srl_453_U218 ( .A1(u4_srl_453_n209), .A2(u4_srl_453_n210), .B1(
        u4_srl_453_n211), .B2(u4_srl_453_n212), .ZN(u4_srl_453_n208) );
  AOI221_X1 u4_srl_453_U217 ( .B1(u4_srl_453_n204), .B2(u4_srl_453_n205), .C1(
        u4_srl_453_n206), .C2(u4_srl_453_n207), .A(u4_srl_453_n208), .ZN(
        u4_srl_453_n193) );
  OAI22_X1 u4_srl_453_U216 ( .A1(u4_srl_453_n200), .A2(u4_srl_453_n201), .B1(
        u4_srl_453_n202), .B2(u4_srl_453_n203), .ZN(u4_srl_453_n199) );
  AOI221_X1 u4_srl_453_U215 ( .B1(u4_srl_453_n195), .B2(u4_srl_453_n196), .C1(
        u4_srl_453_n197), .C2(u4_srl_453_n198), .A(u4_srl_453_n199), .ZN(
        u4_srl_453_n194) );
  AOI21_X1 u4_srl_453_U214 ( .B1(u4_srl_453_n193), .B2(u4_srl_453_n194), .A(
        u4_shift_right[8]), .ZN(u4_N5915) );
  INV_X4 u4_srl_453_U213 ( .A(net33547), .ZN(u4_srl_453_n192) );
  INV_X4 u4_srl_453_U212 ( .A(net33548), .ZN(u4_srl_453_n191) );
  INV_X4 u4_srl_453_U211 ( .A(net33549), .ZN(u4_srl_453_n190) );
  INV_X4 u4_srl_453_U210 ( .A(net33550), .ZN(u4_srl_453_n189) );
  INV_X4 u4_srl_453_U209 ( .A(net33551), .ZN(u4_srl_453_n188) );
  INV_X4 u4_srl_453_U208 ( .A(net33552), .ZN(u4_srl_453_n187) );
  INV_X4 u4_srl_453_U207 ( .A(n8525), .ZN(u4_srl_453_n186) );
  INV_X4 u4_srl_453_U206 ( .A(net33554), .ZN(u4_srl_453_n185) );
  INV_X4 u4_srl_453_U205 ( .A(n8524), .ZN(u4_srl_453_n184) );
  INV_X4 u4_srl_453_U204 ( .A(n8523), .ZN(u4_srl_453_n183) );
  INV_X4 u4_srl_453_U203 ( .A(n8522), .ZN(u4_srl_453_n182) );
  INV_X4 u4_srl_453_U202 ( .A(net33558), .ZN(u4_srl_453_n181) );
  INV_X4 u4_srl_453_U201 ( .A(net33559), .ZN(u4_srl_453_n180) );
  INV_X4 u4_srl_453_U200 ( .A(n8521), .ZN(u4_srl_453_n179) );
  INV_X4 u4_srl_453_U199 ( .A(net33561), .ZN(u4_srl_453_n178) );
  INV_X4 u4_srl_453_U198 ( .A(net33562), .ZN(u4_srl_453_n177) );
  INV_X4 u4_srl_453_U197 ( .A(net33563), .ZN(u4_srl_453_n176) );
  INV_X4 u4_srl_453_U196 ( .A(net33564), .ZN(u4_srl_453_n175) );
  INV_X4 u4_srl_453_U195 ( .A(net33565), .ZN(u4_srl_453_n174) );
  INV_X4 u4_srl_453_U194 ( .A(net33566), .ZN(u4_srl_453_n173) );
  INV_X4 u4_srl_453_U193 ( .A(n8520), .ZN(u4_srl_453_n172) );
  INV_X4 u4_srl_453_U192 ( .A(net33568), .ZN(u4_srl_453_n171) );
  INV_X4 u4_srl_453_U191 ( .A(net33569), .ZN(u4_srl_453_n170) );
  INV_X4 u4_srl_453_U190 ( .A(n8519), .ZN(u4_srl_453_n169) );
  INV_X4 u4_srl_453_U189 ( .A(n8518), .ZN(u4_srl_453_n168) );
  INV_X4 u4_srl_453_U188 ( .A(net33573), .ZN(u4_srl_453_n167) );
  INV_X4 u4_srl_453_U187 ( .A(n8517), .ZN(u4_srl_453_n166) );
  INV_X4 u4_srl_453_U186 ( .A(net33575), .ZN(u4_srl_453_n165) );
  INV_X4 u4_srl_453_U185 ( .A(n8516), .ZN(u4_srl_453_n164) );
  INV_X4 u4_srl_453_U184 ( .A(net33577), .ZN(u4_srl_453_n163) );
  INV_X4 u4_srl_453_U183 ( .A(net33578), .ZN(u4_srl_453_n162) );
  INV_X4 u4_srl_453_U182 ( .A(net33579), .ZN(u4_srl_453_n161) );
  INV_X4 u4_srl_453_U181 ( .A(net33581), .ZN(u4_srl_453_n160) );
  INV_X4 u4_srl_453_U180 ( .A(n8515), .ZN(u4_srl_453_n159) );
  INV_X4 u4_srl_453_U179 ( .A(net33583), .ZN(u4_srl_453_n158) );
  INV_X4 u4_srl_453_U178 ( .A(net33584), .ZN(u4_srl_453_n157) );
  INV_X4 u4_srl_453_U177 ( .A(net33585), .ZN(u4_srl_453_n156) );
  INV_X4 u4_srl_453_U176 ( .A(net33586), .ZN(u4_srl_453_n155) );
  INV_X4 u4_srl_453_U175 ( .A(net33587), .ZN(u4_srl_453_n154) );
  INV_X4 u4_srl_453_U174 ( .A(fract_denorm[50]), .ZN(u4_srl_453_n153) );
  INV_X4 u4_srl_453_U173 ( .A(fract_denorm[51]), .ZN(u4_srl_453_n152) );
  INV_X4 u4_srl_453_U172 ( .A(fract_denorm[74]), .ZN(u4_srl_453_n151) );
  INV_X4 u4_srl_453_U171 ( .A(fract_denorm[82]), .ZN(u4_srl_453_n150) );
  INV_X4 u4_srl_453_U170 ( .A(fract_denorm[66]), .ZN(u4_srl_453_n149) );
  INV_X4 u4_srl_453_U169 ( .A(fract_denorm[58]), .ZN(u4_srl_453_n148) );
  INV_X4 u4_srl_453_U168 ( .A(fract_denorm[52]), .ZN(u4_srl_453_n147) );
  INV_X4 u4_srl_453_U167 ( .A(fract_denorm[71]), .ZN(u4_srl_453_n146) );
  INV_X4 u4_srl_453_U166 ( .A(fract_denorm[73]), .ZN(u4_srl_453_n145) );
  INV_X4 u4_srl_453_U165 ( .A(fract_denorm[72]), .ZN(u4_srl_453_n144) );
  INV_X4 u4_srl_453_U164 ( .A(fract_denorm[70]), .ZN(u4_srl_453_n143) );
  INV_X4 u4_srl_453_U163 ( .A(fract_denorm[69]), .ZN(u4_srl_453_n142) );
  INV_X4 u4_srl_453_U162 ( .A(fract_denorm[68]), .ZN(u4_srl_453_n141) );
  INV_X4 u4_srl_453_U161 ( .A(fract_denorm[67]), .ZN(u4_srl_453_n140) );
  INV_X4 u4_srl_453_U160 ( .A(fract_denorm[63]), .ZN(u4_srl_453_n139) );
  INV_X4 u4_srl_453_U159 ( .A(fract_denorm[65]), .ZN(u4_srl_453_n138) );
  INV_X4 u4_srl_453_U158 ( .A(fract_denorm[64]), .ZN(u4_srl_453_n137) );
  INV_X4 u4_srl_453_U157 ( .A(fract_denorm[62]), .ZN(u4_srl_453_n136) );
  INV_X4 u4_srl_453_U156 ( .A(fract_denorm[61]), .ZN(u4_srl_453_n135) );
  INV_X4 u4_srl_453_U155 ( .A(fract_denorm[60]), .ZN(u4_srl_453_n134) );
  INV_X4 u4_srl_453_U154 ( .A(fract_denorm[59]), .ZN(u4_srl_453_n133) );
  INV_X4 u4_srl_453_U153 ( .A(fract_denorm[79]), .ZN(u4_srl_453_n132) );
  INV_X4 u4_srl_453_U152 ( .A(fract_denorm[81]), .ZN(u4_srl_453_n131) );
  INV_X4 u4_srl_453_U151 ( .A(fract_denorm[80]), .ZN(u4_srl_453_n130) );
  INV_X4 u4_srl_453_U150 ( .A(fract_denorm[78]), .ZN(u4_srl_453_n129) );
  INV_X4 u4_srl_453_U149 ( .A(fract_denorm[77]), .ZN(u4_srl_453_n128) );
  INV_X4 u4_srl_453_U148 ( .A(fract_denorm[76]), .ZN(u4_srl_453_n127) );
  INV_X4 u4_srl_453_U147 ( .A(fract_denorm[75]), .ZN(u4_srl_453_n126) );
  INV_X4 u4_srl_453_U146 ( .A(fract_denorm[87]), .ZN(u4_srl_453_n125) );
  INV_X4 u4_srl_453_U145 ( .A(fract_denorm[89]), .ZN(u4_srl_453_n124) );
  INV_X4 u4_srl_453_U144 ( .A(fract_denorm[88]), .ZN(u4_srl_453_n123) );
  INV_X4 u4_srl_453_U143 ( .A(fract_denorm[86]), .ZN(u4_srl_453_n122) );
  INV_X4 u4_srl_453_U142 ( .A(fract_denorm[85]), .ZN(u4_srl_453_n121) );
  INV_X4 u4_srl_453_U141 ( .A(fract_denorm[84]), .ZN(u4_srl_453_n120) );
  INV_X4 u4_srl_453_U140 ( .A(fract_denorm[83]), .ZN(u4_srl_453_n119) );
  INV_X4 u4_srl_453_U139 ( .A(fract_denorm[55]), .ZN(u4_srl_453_n118) );
  INV_X4 u4_srl_453_U138 ( .A(fract_denorm[57]), .ZN(u4_srl_453_n117) );
  INV_X4 u4_srl_453_U137 ( .A(fract_denorm[56]), .ZN(u4_srl_453_n116) );
  INV_X4 u4_srl_453_U136 ( .A(fract_denorm[54]), .ZN(u4_srl_453_n115) );
  INV_X4 u4_srl_453_U135 ( .A(fract_denorm[53]), .ZN(u4_srl_453_n114) );
  INV_X4 u4_srl_453_U134 ( .A(net33625), .ZN(u4_srl_453_n113) );
  INV_X4 u4_srl_453_U133 ( .A(fract_denorm[98]), .ZN(u4_srl_453_n112) );
  INV_X4 u4_srl_453_U132 ( .A(fract_denorm[102]), .ZN(u4_srl_453_n110) );
  INV_X4 u4_srl_453_U131 ( .A(fract_denorm[99]), .ZN(u4_srl_453_n108) );
  INV_X4 u4_srl_453_U130 ( .A(fract_denorm[90]), .ZN(u4_srl_453_n107) );
  INV_X4 u4_srl_453_U129 ( .A(fract_denorm[95]), .ZN(u4_srl_453_n106) );
  INV_X4 u4_srl_453_U128 ( .A(fract_denorm[97]), .ZN(u4_srl_453_n105) );
  INV_X4 u4_srl_453_U127 ( .A(fract_denorm[94]), .ZN(u4_srl_453_n103) );
  INV_X4 u4_srl_453_U126 ( .A(fract_denorm[93]), .ZN(u4_srl_453_n102) );
  INV_X4 u4_srl_453_U125 ( .A(fract_denorm[92]), .ZN(u4_srl_453_n101) );
  INV_X4 u4_srl_453_U124 ( .A(fract_denorm[91]), .ZN(u4_srl_453_n100) );
  INV_X4 u4_srl_453_U123 ( .A(net33641), .ZN(u4_srl_453_n99) );
  INV_X4 u4_srl_453_U122 ( .A(net33642), .ZN(u4_srl_453_n98) );
  INV_X4 u4_srl_453_U121 ( .A(n8514), .ZN(u4_srl_453_n97) );
  INV_X4 u4_srl_453_U120 ( .A(n8513), .ZN(u4_srl_453_n96) );
  INV_X4 u4_srl_453_U119 ( .A(n8512), .ZN(u4_srl_453_n95) );
  INV_X4 u4_srl_453_U118 ( .A(n8511), .ZN(u4_srl_453_n94) );
  INV_X4 u4_srl_453_U117 ( .A(net33647), .ZN(u4_srl_453_n93) );
  INV_X32 u4_srl_453_U116 ( .A(u4_srl_453_n83), .ZN(u4_srl_453_n86) );
  INV_X32 u4_srl_453_U115 ( .A(u4_srl_453_n86), .ZN(u4_srl_453_n84) );
  INV_X32 u4_srl_453_U114 ( .A(u4_srl_453_n86), .ZN(u4_srl_453_n82) );
  INV_X32 u4_srl_453_U113 ( .A(u4_srl_453_n86), .ZN(u4_srl_453_n81) );
  INV_X32 u4_srl_453_U112 ( .A(u4_srl_453_n86), .ZN(u4_srl_453_n80) );
  INV_X32 u4_srl_453_U111 ( .A(u4_srl_453_n86), .ZN(u4_srl_453_n79) );
  INV_X32 u4_srl_453_U110 ( .A(u4_srl_453_n86), .ZN(u4_srl_453_n78) );
  INV_X32 u4_srl_453_U109 ( .A(u4_srl_453_n76), .ZN(u4_srl_453_n73) );
  INV_X32 u4_srl_453_U108 ( .A(u4_srl_453_n76), .ZN(u4_srl_453_n71) );
  INV_X32 u4_srl_453_U107 ( .A(u4_srl_453_n68), .ZN(u4_srl_453_n67) );
  INV_X32 u4_srl_453_U106 ( .A(u4_srl_453_n68), .ZN(u4_srl_453_n65) );
  INV_X32 u4_srl_453_U105 ( .A(u4_srl_453_n65), .ZN(u4_srl_453_n64) );
  INV_X32 u4_srl_453_U104 ( .A(u4_srl_453_n65), .ZN(u4_srl_453_n63) );
  INV_X32 u4_srl_453_U103 ( .A(u4_srl_453_n65), .ZN(u4_srl_453_n62) );
  INV_X32 u4_srl_453_U102 ( .A(u4_srl_453_n66), .ZN(u4_srl_453_n59) );
  INV_X32 u4_srl_453_U101 ( .A(u4_srl_453_n54), .ZN(u4_srl_453_n53) );
  INV_X32 u4_srl_453_U100 ( .A(u4_srl_453_n5), .ZN(u4_srl_453_n40) );
  INV_X32 u4_srl_453_U99 ( .A(u4_srl_453_n32), .ZN(u4_srl_453_n31) );
  INV_X32 u4_srl_453_U98 ( .A(u4_srl_453_n32), .ZN(u4_srl_453_n30) );
  INV_X32 u4_srl_453_U97 ( .A(u4_srl_453_n32), .ZN(u4_srl_453_n29) );
  INV_X32 u4_srl_453_U96 ( .A(u4_srl_453_n30), .ZN(u4_srl_453_n26) );
  INV_X32 u4_srl_453_U95 ( .A(u4_srl_453_n14), .ZN(u4_srl_453_n21) );
  INV_X32 u4_srl_453_U94 ( .A(u4_srl_453_n14), .ZN(u4_srl_453_n20) );
  INV_X32 u4_srl_453_U93 ( .A(u4_srl_453_n20), .ZN(u4_srl_453_n18) );
  INV_X32 u4_srl_453_U92 ( .A(u4_srl_453_n20), .ZN(u4_srl_453_n17) );
  INV_X32 u4_srl_453_U91 ( .A(u4_srl_453_n21), .ZN(u4_srl_453_n16) );
  INV_X32 u4_srl_453_U90 ( .A(u4_srl_453_n21), .ZN(u4_srl_453_n15) );
  INV_X32 u4_srl_453_U89 ( .A(u4_srl_453_n13), .ZN(u4_srl_453_n9) );
  INV_X32 u4_srl_453_U88 ( .A(u4_srl_453_n13), .ZN(u4_srl_453_n8) );
  INV_X8 u4_srl_453_U87 ( .A(u4_shift_right[4]), .ZN(u4_srl_453_n424) );
  NAND2_X4 u4_srl_453_U86 ( .A1(u4_srl_453_n299), .A2(u4_srl_453_n424), .ZN(
        u4_srl_453_n271) );
  NAND2_X4 u4_srl_453_U85 ( .A1(u4_srl_453_n299), .A2(u4_shift_right[4]), .ZN(
        u4_srl_453_n275) );
  INV_X4 u4_srl_453_U84 ( .A(u4_srl_453_n408), .ZN(u4_srl_453_n415) );
  INV_X4 u4_srl_453_U83 ( .A(u4_srl_453_n891), .ZN(u4_srl_453_n207) );
  NOR2_X4 u4_srl_453_U82 ( .A1(u4_srl_453_n207), .A2(u4_shift_right[8]), .ZN(
        u4_srl_453_n243) );
  NOR2_X4 u4_srl_453_U81 ( .A1(u4_srl_453_n275), .A2(u4_srl_453_n207), .ZN(
        u4_srl_453_n204) );
  NAND2_X4 u4_srl_453_U80 ( .A1(u4_srl_453_n833), .A2(u4_shift_right[4]), .ZN(
        u4_srl_453_n210) );
  NAND2_X4 u4_srl_453_U79 ( .A1(u4_srl_453_n833), .A2(u4_srl_453_n424), .ZN(
        u4_srl_453_n212) );
  AND2_X4 u4_srl_453_U78 ( .A1(u4_srl_453_n28), .A2(u4_srl_453_n826), .ZN(
        u4_srl_453_n195) );
  AND2_X4 u4_srl_453_U77 ( .A1(u4_srl_453_n91), .A2(u4_srl_453_n826), .ZN(
        u4_srl_453_n197) );
  NAND2_X4 u4_srl_453_U76 ( .A1(u4_srl_453_n45), .A2(u4_srl_453_n826), .ZN(
        u4_srl_453_n201) );
  NAND2_X4 u4_srl_453_U75 ( .A1(u4_srl_453_n826), .A2(u4_srl_453_n35), .ZN(
        u4_srl_453_n203) );
  NOR2_X4 u4_srl_453_U74 ( .A1(u4_srl_453_n415), .A2(u4_srl_453_n271), .ZN(
        u4_srl_453_n440) );
  INV_X2 u4_srl_453_U73 ( .A(fract_denorm[96]), .ZN(u4_srl_453_n104) );
  AOI22_X1 u4_srl_453_U72 ( .A1(fract_denorm[101]), .A2(u4_srl_453_n73), .B1(
        fract_denorm[100]), .B2(u4_srl_453_n82), .ZN(u4_srl_453_n853) );
  INV_X2 u4_srl_453_U71 ( .A(fract_denorm[100]), .ZN(u4_srl_453_n111) );
  AOI22_X2 u4_srl_453_U70 ( .A1(u4_srl_453_n67), .A2(fract_denorm[104]), .B1(
        u4_srl_453_n54), .B2(net63217), .ZN(u4_srl_453_n277) );
  AOI22_X1 u4_srl_453_U69 ( .A1(fract_denorm[102]), .A2(u4_srl_453_n69), .B1(
        fract_denorm[101]), .B2(u4_srl_453_n80), .ZN(u4_srl_453_n814) );
  INV_X1 u4_srl_453_U68 ( .A(fract_denorm[101]), .ZN(u4_srl_453_n109) );
  INV_X8 u4_srl_453_U67 ( .A(u4_srl_453_n46), .ZN(u4_srl_453_n45) );
  INV_X16 u4_srl_453_U66 ( .A(u4_srl_453_n29), .ZN(u4_srl_453_n27) );
  INV_X16 u4_srl_453_U65 ( .A(u4_srl_453_n29), .ZN(u4_srl_453_n28) );
  AND2_X4 u4_srl_453_U64 ( .A1(u4_srl_453_n418), .A2(u4_shift_right[4]), .ZN(
        u4_srl_453_n7) );
  INV_X8 u4_srl_453_U63 ( .A(u4_srl_453_n37), .ZN(u4_srl_453_n36) );
  INV_X8 u4_srl_453_U62 ( .A(u4_srl_453_n90), .ZN(u4_srl_453_n88) );
  INV_X8 u4_srl_453_U61 ( .A(u4_srl_453_n4), .ZN(u4_srl_453_n23) );
  OR2_X4 u4_srl_453_U60 ( .A1(u4_srl_453_n760), .A2(u4_srl_453_n866), .ZN(
        u4_srl_453_n6) );
  INV_X16 u4_srl_453_U59 ( .A(u4_srl_453_n13), .ZN(u4_srl_453_n10) );
  INV_X16 u4_srl_453_U58 ( .A(u4_srl_453_n54), .ZN(u4_srl_453_n52) );
  INV_X16 u4_srl_453_U57 ( .A(u4_srl_453_n76), .ZN(u4_srl_453_n69) );
  INV_X16 u4_srl_453_U56 ( .A(u4_srl_453_n76), .ZN(u4_srl_453_n72) );
  INV_X16 u4_srl_453_U55 ( .A(u4_srl_453_n86), .ZN(u4_srl_453_n85) );
  INV_X8 u4_srl_453_U54 ( .A(u4_srl_453_n4), .ZN(u4_srl_453_n24) );
  INV_X4 u4_srl_453_U53 ( .A(u4_srl_453_n87), .ZN(u4_srl_453_n90) );
  NAND2_X2 u4_srl_453_U52 ( .A1(u4_srl_453_n418), .A2(u4_srl_453_n424), .ZN(
        u4_srl_453_n214) );
  INV_X4 u4_srl_453_U51 ( .A(u4_srl_453_n425), .ZN(u4_srl_453_n39) );
  INV_X4 u4_srl_453_U50 ( .A(u4_srl_453_n39), .ZN(u4_srl_453_n38) );
  INV_X4 u4_srl_453_U49 ( .A(u4_srl_453_n57), .ZN(u4_srl_453_n54) );
  INV_X4 u4_srl_453_U48 ( .A(u4_srl_453_n426), .ZN(u4_srl_453_n58) );
  INV_X4 u4_srl_453_U47 ( .A(u4_srl_453_n58), .ZN(u4_srl_453_n56) );
  INV_X4 u4_srl_453_U46 ( .A(u4_srl_453_n66), .ZN(u4_srl_453_n61) );
  INV_X4 u4_srl_453_U45 ( .A(u4_srl_453_n66), .ZN(u4_srl_453_n60) );
  INV_X16 u4_srl_453_U44 ( .A(u4_srl_453_n92), .ZN(u4_srl_453_n91) );
  INV_X16 u4_srl_453_U43 ( .A(u4_srl_453_n47), .ZN(u4_srl_453_n46) );
  INV_X4 u4_srl_453_U42 ( .A(u4_srl_453_n5), .ZN(u4_srl_453_n47) );
  INV_X8 u4_srl_453_U41 ( .A(u4_srl_453_n39), .ZN(u4_srl_453_n35) );
  INV_X4 u4_srl_453_U40 ( .A(u4_srl_453_n38), .ZN(u4_srl_453_n37) );
  INV_X4 u4_srl_453_U39 ( .A(u4_srl_453_n55), .ZN(u4_srl_453_n48) );
  INV_X4 u4_srl_453_U38 ( .A(u4_srl_453_n58), .ZN(u4_srl_453_n57) );
  INV_X4 u4_srl_453_U37 ( .A(u4_srl_453_n441), .ZN(u4_srl_453_n89) );
  INV_X4 u4_srl_453_U36 ( .A(u4_srl_453_n441), .ZN(u4_srl_453_n92) );
  OR2_X4 u4_srl_453_U35 ( .A1(u4_shift_right[2]), .A2(u4_srl_453_n865), .ZN(
        u4_srl_453_n5) );
  OR2_X4 u4_srl_453_U34 ( .A1(u4_srl_453_n332), .A2(u4_shift_right[4]), .ZN(
        u4_srl_453_n4) );
  INV_X8 u4_srl_453_U33 ( .A(u4_srl_453_n56), .ZN(u4_srl_453_n55) );
  INV_X16 u4_srl_453_U32 ( .A(u4_srl_453_n74), .ZN(u4_srl_453_n76) );
  INV_X4 u4_srl_453_U31 ( .A(u4_srl_453_n428), .ZN(u4_srl_453_n77) );
  INV_X4 u4_srl_453_U30 ( .A(u4_srl_453_n1), .ZN(u4_srl_453_n83) );
  AND2_X4 u4_srl_453_U29 ( .A1(u4_srl_453_n910), .A2(u4_srl_453_n911), .ZN(
        u4_srl_453_n3) );
  INV_X4 u4_srl_453_U28 ( .A(u4_srl_453_n92), .ZN(u4_srl_453_n87) );
  NOR2_X2 u4_srl_453_U27 ( .A1(u4_srl_453_n760), .A2(u4_shift_right[2]), .ZN(
        u4_srl_453_n441) );
  OR2_X4 u4_srl_453_U26 ( .A1(u4_srl_453_n332), .A2(u4_srl_453_n424), .ZN(
        u4_srl_453_n2) );
  OR2_X4 u4_srl_453_U25 ( .A1(u4_shift_right[0]), .A2(u4_srl_453_n910), .ZN(
        u4_srl_453_n1) );
  INV_X4 u4_srl_453_U24 ( .A(u4_srl_453_n77), .ZN(u4_srl_453_n74) );
  INV_X4 u4_srl_453_U23 ( .A(u4_srl_453_n214), .ZN(u4_srl_453_n12) );
  INV_X16 u4_srl_453_U22 ( .A(u4_srl_453_n12), .ZN(u4_srl_453_n11) );
  INV_X16 u4_srl_453_U21 ( .A(u4_srl_453_n2), .ZN(u4_srl_453_n22) );
  INV_X16 u4_srl_453_U20 ( .A(u4_srl_453_n20), .ZN(u4_srl_453_n19) );
  INV_X4 u4_srl_453_U19 ( .A(u4_srl_453_n214), .ZN(u4_srl_453_n13) );
  INV_X16 u4_srl_453_U18 ( .A(u4_srl_453_n30), .ZN(u4_srl_453_n25) );
  INV_X4 u4_srl_453_U17 ( .A(u4_srl_453_n37), .ZN(u4_srl_453_n33) );
  INV_X16 u4_srl_453_U16 ( .A(u4_srl_453_n46), .ZN(u4_srl_453_n42) );
  INV_X4 u4_srl_453_U15 ( .A(u4_srl_453_n37), .ZN(u4_srl_453_n34) );
  INV_X16 u4_srl_453_U14 ( .A(u4_srl_453_n46), .ZN(u4_srl_453_n43) );
  INV_X16 u4_srl_453_U13 ( .A(u4_srl_453_n46), .ZN(u4_srl_453_n41) );
  INV_X16 u4_srl_453_U12 ( .A(u4_srl_453_n46), .ZN(u4_srl_453_n44) );
  INV_X16 u4_srl_453_U11 ( .A(u4_srl_453_n55), .ZN(u4_srl_453_n50) );
  INV_X16 u4_srl_453_U10 ( .A(u4_srl_453_n55), .ZN(u4_srl_453_n51) );
  INV_X16 u4_srl_453_U9 ( .A(u4_srl_453_n55), .ZN(u4_srl_453_n49) );
  INV_X16 u4_srl_453_U8 ( .A(u4_srl_453_n76), .ZN(u4_srl_453_n75) );
  INV_X16 u4_srl_453_U7 ( .A(u4_srl_453_n76), .ZN(u4_srl_453_n70) );
  INV_X8 u4_srl_453_U6 ( .A(u4_srl_453_n6), .ZN(u4_srl_453_n32) );
  INV_X16 u4_srl_453_U5 ( .A(u4_srl_453_n3), .ZN(u4_srl_453_n68) );
  INV_X16 u4_srl_453_U4 ( .A(u4_srl_453_n68), .ZN(u4_srl_453_n66) );
  INV_X16 u4_srl_453_U3 ( .A(u4_srl_453_n7), .ZN(u4_srl_453_n14) );
  OR3_X1 u4_sll_482_U69 ( .A1(u4_f2i_shft_8_), .A2(u4_f2i_shft_9_), .A3(
        u4_f2i_shft_7_), .ZN(u4_sll_482_n59) );
  NAND2_X1 u4_sll_482_U68 ( .A1(u4_sll_482_n59), .A2(u4_sll_482_n50), .ZN(
        u4_sll_482_n52) );
  NAND3_X1 u4_sll_482_U67 ( .A1(u4_f2i_shft_8_), .A2(u4_f2i_shft_7_), .A3(
        u4_f2i_shft_9_), .ZN(u4_sll_482_n58) );
  NAND2_X1 u4_sll_482_U66 ( .A1(u4_f2i_shft_10_), .A2(u4_sll_482_n58), .ZN(
        u4_sll_482_n51) );
  NAND2_X1 u4_sll_482_U65 ( .A1(net43686), .A2(u4_sll_482_n51), .ZN(
        u4_sll_482_n57) );
  NAND2_X1 u4_sll_482_U64 ( .A1(u4_sll_482_n52), .A2(u4_sll_482_n57), .ZN(
        u4_sll_482_temp_int_SH_0_) );
  AND2_X1 u4_sll_482_U63 ( .A1(net33546), .A2(u4_sll_482_n9), .ZN(
        u4_sll_482_ML_int_1__0_) );
  NAND2_X1 u4_sll_482_U62 ( .A1(u4_exp_in_mi1_1_), .A2(u4_sll_482_n51), .ZN(
        u4_sll_482_n56) );
  NAND2_X1 u4_sll_482_U61 ( .A1(u4_f2i_shft_2_), .A2(u4_sll_482_n51), .ZN(
        u4_sll_482_n55) );
  NAND2_X1 u4_sll_482_U60 ( .A1(u4_sll_482_n52), .A2(u4_sll_482_n55), .ZN(
        u4_sll_482_temp_int_SH_2_) );
  NAND2_X1 u4_sll_482_U59 ( .A1(u4_f2i_shft_3_), .A2(u4_sll_482_n51), .ZN(
        u4_sll_482_n54) );
  NAND2_X1 u4_sll_482_U58 ( .A1(u4_sll_482_n52), .A2(u4_sll_482_n54), .ZN(
        u4_sll_482_temp_int_SH_3_) );
  NAND2_X1 u4_sll_482_U57 ( .A1(n4295), .A2(u4_sll_482_n51), .ZN(
        u4_sll_482_n53) );
  AND2_X1 u4_sll_482_U56 ( .A1(u4_sll_482_ML_int_4__12_), .A2(u4_sll_482_n46), 
        .ZN(u4_sll_482_ML_int_5__12_) );
  AND2_X1 u4_sll_482_U55 ( .A1(u4_sll_482_ML_int_7__108_), .A2(u4_sll_482_n50), 
        .ZN(u4_exp_f2i_1_108_) );
  OAI21_X1 u4_sll_482_U54 ( .B1(n4329), .B2(u4_sll_482_n49), .A(u4_sll_482_n51), .ZN(u4_sll_482_SHMAG[5]) );
  OAI21_X1 u4_sll_482_U53 ( .B1(u4_f2i_shft_6_), .B2(u4_sll_482_n49), .A(
        u4_sll_482_n51), .ZN(u4_sll_482_SHMAG[6]) );
  INV_X4 u4_sll_482_U52 ( .A(u4_sll_482_n52), .ZN(u4_sll_482_n49) );
  INV_X4 u4_sll_482_U51 ( .A(u4_sll_482_SHMAG[6]), .ZN(u4_sll_482_n48) );
  INV_X32 u4_sll_482_U50 ( .A(u4_sll_482_n26), .ZN(u4_sll_482_n25) );
  INV_X32 u4_sll_482_U49 ( .A(u4_sll_482_n18), .ZN(u4_sll_482_n15) );
  INV_X16 u4_sll_482_U48 ( .A(u4_sll_482_n15), .ZN(u4_sll_482_n14) );
  INV_X16 u4_sll_482_U47 ( .A(u4_sll_482_n15), .ZN(u4_sll_482_n13) );
  INV_X16 u4_sll_482_U46 ( .A(u4_sll_482_n16), .ZN(u4_sll_482_n12) );
  INV_X16 u4_sll_482_U45 ( .A(u4_sll_482_n16), .ZN(u4_sll_482_n11) );
  INV_X16 u4_sll_482_U44 ( .A(u4_sll_482_n16), .ZN(u4_sll_482_n10) );
  INV_X32 u4_sll_482_U43 ( .A(u4_sll_482_n11), .ZN(u4_sll_482_n7) );
  INV_X32 u4_sll_482_U42 ( .A(u4_sll_482_n12), .ZN(u4_sll_482_n6) );
  INV_X32 u4_sll_482_U41 ( .A(u4_sll_482_n13), .ZN(u4_sll_482_n5) );
  INV_X32 u4_sll_482_U40 ( .A(u4_sll_482_n14), .ZN(u4_sll_482_n4) );
  INV_X4 u4_sll_482_U39 ( .A(u4_sll_482_n2), .ZN(u4_sll_482_n45) );
  INV_X1 u4_sll_482_U38 ( .A(u4_sll_482_n45), .ZN(u4_sll_482_n46) );
  INV_X4 u4_sll_482_U37 ( .A(u4_sll_482_n18), .ZN(u4_sll_482_n17) );
  INV_X2 u4_sll_482_U36 ( .A(u4_sll_482_n17), .ZN(u4_sll_482_n9) );
  INV_X8 u4_sll_482_U35 ( .A(u4_sll_482_n42), .ZN(u4_sll_482_n41) );
  INV_X16 u4_sll_482_U34 ( .A(u4_sll_482_n40), .ZN(u4_sll_482_n39) );
  INV_X2 u4_sll_482_U33 ( .A(u4_sll_482_SHMAG[5]), .ZN(u4_sll_482_n47) );
  AND2_X2 u4_sll_482_U32 ( .A1(u4_sll_482_ML_int_1__0_), .A2(u4_sll_482_n28), 
        .ZN(u4_sll_482_n3) );
  INV_X8 u4_sll_482_U31 ( .A(u4_sll_482_n34), .ZN(u4_sll_482_n30) );
  INV_X4 u4_sll_482_U30 ( .A(u4_sll_482_n38), .ZN(u4_sll_482_n37) );
  INV_X4 u4_sll_482_U29 ( .A(u4_sll_482_n29), .ZN(u4_sll_482_n28) );
  INV_X4 u4_sll_482_U28 ( .A(u4_sll_482_n38), .ZN(u4_sll_482_n35) );
  INV_X4 u4_sll_482_U27 ( .A(u4_sll_482_n27), .ZN(u4_sll_482_n19) );
  INV_X4 u4_sll_482_U26 ( .A(u4_sll_482_n1), .ZN(u4_sll_482_n22) );
  INV_X4 u4_sll_482_U25 ( .A(u4_sll_482_n1), .ZN(u4_sll_482_n29) );
  AND2_X2 u4_sll_482_U24 ( .A1(u4_sll_482_n52), .A2(u4_sll_482_n53), .ZN(
        u4_sll_482_n2) );
  INV_X16 u4_sll_482_U23 ( .A(u4_sll_482_n40), .ZN(u4_sll_482_n38) );
  INV_X4 u4_sll_482_U22 ( .A(u4_sll_482_n38), .ZN(u4_sll_482_n36) );
  INV_X8 u4_sll_482_U21 ( .A(u4_sll_482_n43), .ZN(u4_sll_482_n42) );
  AND2_X2 u4_sll_482_U20 ( .A1(u4_sll_482_n52), .A2(u4_sll_482_n56), .ZN(
        u4_sll_482_n1) );
  INV_X2 u4_sll_482_U19 ( .A(u4_sll_482_temp_int_SH_3_), .ZN(u4_sll_482_n44)
         );
  INV_X4 u4_sll_482_U18 ( .A(u4_sll_482_n44), .ZN(u4_sll_482_n43) );
  INV_X4 u4_sll_482_U17 ( .A(u4_sll_482_n39), .ZN(u4_sll_482_n34) );
  INV_X8 u4_sll_482_U16 ( .A(u4_sll_482_n29), .ZN(u4_sll_482_n27) );
  INV_X4 u4_sll_482_U15 ( .A(u4_f2i_shft_10_), .ZN(u4_sll_482_n50) );
  INV_X4 u4_sll_482_U14 ( .A(u4_sll_482_n35), .ZN(u4_sll_482_n31) );
  INV_X8 u4_sll_482_U13 ( .A(u4_sll_482_n22), .ZN(u4_sll_482_n26) );
  INV_X4 u4_sll_482_U12 ( .A(u4_sll_482_n37), .ZN(u4_sll_482_n33) );
  INV_X4 u4_sll_482_U11 ( .A(u4_sll_482_n28), .ZN(u4_sll_482_n24) );
  INV_X4 u4_sll_482_U10 ( .A(u4_sll_482_n36), .ZN(u4_sll_482_n32) );
  INV_X8 u4_sll_482_U9 ( .A(u4_sll_482_n27), .ZN(u4_sll_482_n21) );
  INV_X4 u4_sll_482_U8 ( .A(u4_sll_482_n27), .ZN(u4_sll_482_n23) );
  INV_X16 u4_sll_482_U7 ( .A(u4_sll_482_n10), .ZN(u4_sll_482_n8) );
  INV_X4 u4_sll_482_U6 ( .A(u4_sll_482_temp_int_SH_2_), .ZN(u4_sll_482_n40) );
  INV_X4 u4_sll_482_U5 ( .A(u4_sll_482_n27), .ZN(u4_sll_482_n20) );
  INV_X4 u4_sll_482_U4 ( .A(u4_sll_482_temp_int_SH_0_), .ZN(u4_sll_482_n18) );
  INV_X16 u4_sll_482_U3 ( .A(u4_sll_482_n18), .ZN(u4_sll_482_n16) );
  MUX2_X2 u4_sll_482_M1_0_2 ( .A(net33647), .B(net33648), .S(u4_sll_482_n17), 
        .Z(u4_sll_482_ML_int_1__2_) );
  MUX2_X2 u4_sll_482_M1_0_4 ( .A(n8512), .B(n8511), .S(u4_sll_482_n8), .Z(
        u4_sll_482_ML_int_1__4_) );
  MUX2_X2 u4_sll_482_M1_0_6 ( .A(n8514), .B(n8513), .S(u4_sll_482_n8), .Z(
        u4_sll_482_ML_int_1__6_) );
  MUX2_X2 u4_sll_482_M1_0_8 ( .A(net33641), .B(net33642), .S(u4_sll_482_n8), 
        .Z(u4_sll_482_ML_int_1__8_) );
  MUX2_X2 u4_sll_482_M1_0_10 ( .A(net33549), .B(net33548), .S(u4_sll_482_n8), 
        .Z(u4_sll_482_ML_int_1__10_) );
  MUX2_X2 u4_sll_482_M1_0_12 ( .A(net33579), .B(net33581), .S(u4_sll_482_n8), 
        .Z(u4_sll_482_ML_int_1__12_) );
  MUX2_X2 u4_sll_482_M1_0_14 ( .A(net33577), .B(net33578), .S(u4_sll_482_n8), 
        .Z(u4_sll_482_ML_int_1__14_) );
  MUX2_X2 u4_sll_482_M1_0_16 ( .A(n8516), .B(n8517), .S(u4_sll_482_n15), .Z(
        u4_sll_482_ML_int_1__16_) );
  MUX2_X2 u4_sll_482_M1_0_18 ( .A(net33550), .B(net33575), .S(u4_sll_482_n15), 
        .Z(u4_sll_482_ML_int_1__18_) );
  MUX2_X2 u4_sll_482_M1_0_20 ( .A(net33572), .B(net33573), .S(u4_sll_482_n4), 
        .Z(u4_sll_482_ML_int_1__20_) );
  MUX2_X2 u4_sll_482_M1_0_22 ( .A(n8519), .B(n8518), .S(u4_sll_482_n5), .Z(
        u4_sll_482_ML_int_1__22_) );
  MUX2_X2 u4_sll_482_M1_0_24 ( .A(net33569), .B(n8520), .S(u4_sll_482_n17), 
        .Z(u4_sll_482_ML_int_1__24_) );
  MUX2_X2 u4_sll_482_M1_0_26 ( .A(net33551), .B(net33568), .S(u4_sll_482_n7), 
        .Z(u4_sll_482_ML_int_1__26_) );
  MUX2_X2 u4_sll_482_M1_0_28 ( .A(net33565), .B(net33566), .S(u4_sll_482_n7), 
        .Z(u4_sll_482_ML_int_1__28_) );
  MUX2_X2 u4_sll_482_M1_0_30 ( .A(net33563), .B(net33564), .S(u4_sll_482_n7), 
        .Z(u4_sll_482_ML_int_1__30_) );
  MUX2_X2 u4_sll_482_M1_0_32 ( .A(net33562), .B(n8521), .S(u4_sll_482_n7), .Z(
        u4_sll_482_ML_int_1__32_) );
  MUX2_X2 u4_sll_482_M1_0_34 ( .A(net33552), .B(net33561), .S(u4_sll_482_n7), 
        .Z(u4_sll_482_ML_int_1__34_) );
  MUX2_X2 u4_sll_482_M1_0_36 ( .A(net33558), .B(net33559), .S(u4_sll_482_n7), 
        .Z(u4_sll_482_ML_int_1__36_) );
  MUX2_X2 u4_sll_482_M1_0_38 ( .A(n8523), .B(n8522), .S(u4_sll_482_n4), .Z(
        u4_sll_482_ML_int_1__38_) );
  MUX2_X2 u4_sll_482_M1_0_40 ( .A(n8524), .B(n8525), .S(u4_sll_482_n4), .Z(
        u4_sll_482_ML_int_1__40_) );
  MUX2_X2 u4_sll_482_M1_0_42 ( .A(net33547), .B(net33554), .S(u4_sll_482_n4), 
        .Z(u4_sll_482_ML_int_1__42_) );
  MUX2_X2 u4_sll_482_M1_0_44 ( .A(net33586), .B(net33587), .S(u4_sll_482_n4), 
        .Z(u4_sll_482_ML_int_1__44_) );
  MUX2_X2 u4_sll_482_M1_0_46 ( .A(net33584), .B(net33585), .S(u4_sll_482_n15), 
        .Z(u4_sll_482_ML_int_1__46_) );
  MUX2_X2 u4_sll_482_M1_0_48 ( .A(net33583), .B(n8515), .S(u4_sll_482_n6), .Z(
        u4_sll_482_ML_int_1__48_) );
  MUX2_X2 u4_sll_482_M1_0_50 ( .A(fract_denorm[50]), .B(net33625), .S(
        u4_sll_482_n6), .Z(u4_sll_482_ML_int_1__50_) );
  MUX2_X2 u4_sll_482_M1_0_52 ( .A(fract_denorm[52]), .B(fract_denorm[51]), .S(
        u4_sll_482_n6), .Z(u4_sll_482_ML_int_1__52_) );
  MUX2_X2 u4_sll_482_M1_0_54 ( .A(fract_denorm[54]), .B(fract_denorm[53]), .S(
        u4_sll_482_n6), .Z(u4_sll_482_ML_int_1__54_) );
  MUX2_X2 u4_sll_482_M1_0_56 ( .A(fract_denorm[56]), .B(fract_denorm[55]), .S(
        u4_sll_482_n6), .Z(u4_sll_482_ML_int_1__56_) );
  MUX2_X2 u4_sll_482_M1_0_58 ( .A(fract_denorm[58]), .B(fract_denorm[57]), .S(
        u4_sll_482_n6), .Z(u4_sll_482_ML_int_1__58_) );
  MUX2_X2 u4_sll_482_M1_0_60 ( .A(fract_denorm[60]), .B(fract_denorm[59]), .S(
        u4_sll_482_n4), .Z(u4_sll_482_ML_int_1__60_) );
  MUX2_X2 u4_sll_482_M1_0_62 ( .A(fract_denorm[62]), .B(fract_denorm[61]), .S(
        u4_sll_482_n5), .Z(u4_sll_482_ML_int_1__62_) );
  MUX2_X2 u4_sll_482_M1_0_64 ( .A(fract_denorm[64]), .B(fract_denorm[63]), .S(
        u4_sll_482_n4), .Z(u4_sll_482_ML_int_1__64_) );
  MUX2_X2 u4_sll_482_M1_0_66 ( .A(fract_denorm[66]), .B(fract_denorm[65]), .S(
        u4_sll_482_n4), .Z(u4_sll_482_ML_int_1__66_) );
  MUX2_X2 u4_sll_482_M1_0_68 ( .A(fract_denorm[68]), .B(fract_denorm[67]), .S(
        u4_sll_482_n4), .Z(u4_sll_482_ML_int_1__68_) );
  MUX2_X2 u4_sll_482_M1_0_70 ( .A(fract_denorm[70]), .B(fract_denorm[69]), .S(
        u4_sll_482_n5), .Z(u4_sll_482_ML_int_1__70_) );
  MUX2_X2 u4_sll_482_M1_0_72 ( .A(fract_denorm[72]), .B(fract_denorm[71]), .S(
        u4_sll_482_n5), .Z(u4_sll_482_ML_int_1__72_) );
  MUX2_X2 u4_sll_482_M1_0_74 ( .A(fract_denorm[74]), .B(fract_denorm[73]), .S(
        u4_sll_482_n5), .Z(u4_sll_482_ML_int_1__74_) );
  MUX2_X2 u4_sll_482_M1_0_76 ( .A(fract_denorm[76]), .B(fract_denorm[75]), .S(
        u4_sll_482_n5), .Z(u4_sll_482_ML_int_1__76_) );
  MUX2_X2 u4_sll_482_M1_0_78 ( .A(fract_denorm[78]), .B(fract_denorm[77]), .S(
        u4_sll_482_n5), .Z(u4_sll_482_ML_int_1__78_) );
  MUX2_X2 u4_sll_482_M1_0_80 ( .A(fract_denorm[80]), .B(fract_denorm[79]), .S(
        u4_sll_482_n5), .Z(u4_sll_482_ML_int_1__80_) );
  MUX2_X2 u4_sll_482_M1_0_82 ( .A(fract_denorm[82]), .B(fract_denorm[81]), .S(
        u4_sll_482_n17), .Z(u4_sll_482_ML_int_1__82_) );
  MUX2_X2 u4_sll_482_M1_0_84 ( .A(fract_denorm[84]), .B(fract_denorm[83]), .S(
        u4_sll_482_n4), .Z(u4_sll_482_ML_int_1__84_) );
  MUX2_X2 u4_sll_482_M1_0_86 ( .A(fract_denorm[86]), .B(fract_denorm[85]), .S(
        u4_sll_482_n4), .Z(u4_sll_482_ML_int_1__86_) );
  MUX2_X2 u4_sll_482_M1_0_88 ( .A(fract_denorm[88]), .B(fract_denorm[87]), .S(
        u4_sll_482_n4), .Z(u4_sll_482_ML_int_1__88_) );
  MUX2_X2 u4_sll_482_M1_0_90 ( .A(fract_denorm[90]), .B(fract_denorm[89]), .S(
        u4_sll_482_n4), .Z(u4_sll_482_ML_int_1__90_) );
  MUX2_X2 u4_sll_482_M1_0_92 ( .A(fract_denorm[92]), .B(fract_denorm[91]), .S(
        u4_sll_482_n4), .Z(u4_sll_482_ML_int_1__92_) );
  MUX2_X2 u4_sll_482_M1_0_94 ( .A(fract_denorm[94]), .B(fract_denorm[93]), .S(
        u4_sll_482_n4), .Z(u4_sll_482_ML_int_1__94_) );
  MUX2_X2 u4_sll_482_M1_0_96 ( .A(fract_denorm[96]), .B(fract_denorm[95]), .S(
        u4_sll_482_n4), .Z(u4_sll_482_ML_int_1__96_) );
  MUX2_X2 u4_sll_482_M1_0_98 ( .A(fract_denorm[98]), .B(fract_denorm[97]), .S(
        u4_sll_482_n4), .Z(u4_sll_482_ML_int_1__98_) );
  MUX2_X2 u4_sll_482_M1_0_100 ( .A(fract_denorm[100]), .B(fract_denorm[99]), 
        .S(u4_sll_482_n4), .Z(u4_sll_482_ML_int_1__100_) );
  MUX2_X2 u4_sll_482_M1_0_102 ( .A(fract_denorm[102]), .B(fract_denorm[101]), 
        .S(u4_sll_482_n4), .Z(u4_sll_482_ML_int_1__102_) );
  MUX2_X2 u4_sll_482_M1_0_104 ( .A(fract_denorm[104]), .B(fract_denorm[103]), 
        .S(u4_sll_482_n17), .Z(u4_sll_482_ML_int_1__104_) );
  MUX2_X2 u4_sll_482_M1_0_106 ( .A(net63217), .B(net63217), .S(u4_sll_482_n17), 
        .Z(u4_sll_482_ML_int_1__106_) );
  MUX2_X2 u4_sll_482_M1_0_108 ( .A(net63217), .B(net63217), .S(u4_sll_482_n17), 
        .Z(u4_sll_482_ML_int_1__108_) );
  MUX2_X2 u4_sll_482_M1_1_4 ( .A(u4_sll_482_ML_int_1__4_), .B(
        u4_sll_482_ML_int_1__2_), .S(u4_sll_482_n25), .Z(
        u4_sll_482_ML_int_2__4_) );
  MUX2_X2 u4_sll_482_M1_1_8 ( .A(u4_sll_482_ML_int_1__8_), .B(
        u4_sll_482_ML_int_1__6_), .S(u4_sll_482_n25), .Z(
        u4_sll_482_ML_int_2__8_) );
  MUX2_X2 u4_sll_482_M1_1_12 ( .A(u4_sll_482_ML_int_1__12_), .B(
        u4_sll_482_ML_int_1__10_), .S(u4_sll_482_n25), .Z(
        u4_sll_482_ML_int_2__12_) );
  MUX2_X2 u4_sll_482_M1_1_16 ( .A(u4_sll_482_ML_int_1__16_), .B(
        u4_sll_482_ML_int_1__14_), .S(u4_sll_482_n29), .Z(
        u4_sll_482_ML_int_2__16_) );
  MUX2_X2 u4_sll_482_M1_1_20 ( .A(u4_sll_482_ML_int_1__20_), .B(
        u4_sll_482_ML_int_1__18_), .S(u4_sll_482_n19), .Z(
        u4_sll_482_ML_int_2__20_) );
  MUX2_X2 u4_sll_482_M1_1_24 ( .A(u4_sll_482_ML_int_1__24_), .B(
        u4_sll_482_ML_int_1__22_), .S(u4_sll_482_n19), .Z(
        u4_sll_482_ML_int_2__24_) );
  MUX2_X2 u4_sll_482_M1_1_28 ( .A(u4_sll_482_ML_int_1__28_), .B(
        u4_sll_482_ML_int_1__26_), .S(u4_sll_482_n19), .Z(
        u4_sll_482_ML_int_2__28_) );
  MUX2_X2 u4_sll_482_M1_1_32 ( .A(u4_sll_482_ML_int_1__32_), .B(
        u4_sll_482_ML_int_1__30_), .S(u4_sll_482_n19), .Z(
        u4_sll_482_ML_int_2__32_) );
  MUX2_X2 u4_sll_482_M1_1_36 ( .A(u4_sll_482_ML_int_1__36_), .B(
        u4_sll_482_ML_int_1__34_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__36_) );
  MUX2_X2 u4_sll_482_M1_1_40 ( .A(u4_sll_482_ML_int_1__40_), .B(
        u4_sll_482_ML_int_1__38_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__40_) );
  MUX2_X2 u4_sll_482_M1_1_44 ( .A(u4_sll_482_ML_int_1__44_), .B(
        u4_sll_482_ML_int_1__42_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__44_) );
  MUX2_X2 u4_sll_482_M1_1_48 ( .A(u4_sll_482_ML_int_1__48_), .B(
        u4_sll_482_ML_int_1__46_), .S(u4_sll_482_n21), .Z(
        u4_sll_482_ML_int_2__48_) );
  MUX2_X2 u4_sll_482_M1_1_52 ( .A(u4_sll_482_ML_int_1__52_), .B(
        u4_sll_482_ML_int_1__50_), .S(u4_sll_482_n21), .Z(
        u4_sll_482_ML_int_2__52_) );
  MUX2_X2 u4_sll_482_M1_1_56 ( .A(u4_sll_482_ML_int_1__56_), .B(
        u4_sll_482_ML_int_1__54_), .S(u4_sll_482_n21), .Z(
        u4_sll_482_ML_int_2__56_) );
  MUX2_X2 u4_sll_482_M1_1_60 ( .A(u4_sll_482_ML_int_1__60_), .B(
        u4_sll_482_ML_int_1__58_), .S(u4_sll_482_n22), .Z(
        u4_sll_482_ML_int_2__60_) );
  MUX2_X2 u4_sll_482_M1_1_64 ( .A(u4_sll_482_ML_int_1__64_), .B(
        u4_sll_482_ML_int_1__62_), .S(u4_sll_482_n22), .Z(
        u4_sll_482_ML_int_2__64_) );
  MUX2_X2 u4_sll_482_M1_1_68 ( .A(u4_sll_482_ML_int_1__68_), .B(
        u4_sll_482_ML_int_1__66_), .S(u4_sll_482_n23), .Z(
        u4_sll_482_ML_int_2__68_) );
  MUX2_X2 u4_sll_482_M1_1_72 ( .A(u4_sll_482_ML_int_1__72_), .B(
        u4_sll_482_ML_int_1__70_), .S(u4_sll_482_n23), .Z(
        u4_sll_482_ML_int_2__72_) );
  MUX2_X2 u4_sll_482_M1_1_76 ( .A(u4_sll_482_ML_int_1__76_), .B(
        u4_sll_482_ML_int_1__74_), .S(u4_sll_482_n23), .Z(
        u4_sll_482_ML_int_2__76_) );
  MUX2_X2 u4_sll_482_M1_1_80 ( .A(u4_sll_482_ML_int_1__80_), .B(
        u4_sll_482_ML_int_1__78_), .S(u4_sll_482_n24), .Z(
        u4_sll_482_ML_int_2__80_) );
  MUX2_X2 u4_sll_482_M1_1_84 ( .A(u4_sll_482_ML_int_1__84_), .B(
        u4_sll_482_ML_int_1__82_), .S(u4_sll_482_n24), .Z(
        u4_sll_482_ML_int_2__84_) );
  MUX2_X2 u4_sll_482_M1_1_88 ( .A(u4_sll_482_ML_int_1__88_), .B(
        u4_sll_482_ML_int_1__86_), .S(u4_sll_482_n24), .Z(
        u4_sll_482_ML_int_2__88_) );
  MUX2_X2 u4_sll_482_M1_1_92 ( .A(u4_sll_482_ML_int_1__92_), .B(
        u4_sll_482_ML_int_1__90_), .S(u4_sll_482_n25), .Z(
        u4_sll_482_ML_int_2__92_) );
  MUX2_X2 u4_sll_482_M1_1_96 ( .A(u4_sll_482_ML_int_1__96_), .B(
        u4_sll_482_ML_int_1__94_), .S(u4_sll_482_n25), .Z(
        u4_sll_482_ML_int_2__96_) );
  MUX2_X2 u4_sll_482_M1_1_100 ( .A(u4_sll_482_ML_int_1__100_), .B(
        u4_sll_482_ML_int_1__98_), .S(u4_sll_482_n25), .Z(
        u4_sll_482_ML_int_2__100_) );
  MUX2_X2 u4_sll_482_M1_1_104 ( .A(u4_sll_482_ML_int_1__104_), .B(
        u4_sll_482_ML_int_1__102_), .S(u4_sll_482_n25), .Z(
        u4_sll_482_ML_int_2__104_) );
  MUX2_X2 u4_sll_482_M1_1_108 ( .A(u4_sll_482_ML_int_1__108_), .B(
        u4_sll_482_ML_int_1__106_), .S(u4_sll_482_n25), .Z(
        u4_sll_482_ML_int_2__108_) );
  MUX2_X2 u4_sll_482_M1_2_4 ( .A(u4_sll_482_ML_int_2__4_), .B(u4_sll_482_n3), 
        .S(u4_sll_482_n30), .Z(u4_sll_482_ML_int_3__4_) );
  MUX2_X2 u4_sll_482_M1_2_12 ( .A(u4_sll_482_ML_int_2__12_), .B(
        u4_sll_482_ML_int_2__8_), .S(u4_sll_482_n30), .Z(
        u4_sll_482_ML_int_3__12_) );
  MUX2_X2 u4_sll_482_M1_2_20 ( .A(u4_sll_482_ML_int_2__20_), .B(
        u4_sll_482_ML_int_2__16_), .S(u4_sll_482_n39), .Z(
        u4_sll_482_ML_int_3__20_) );
  MUX2_X2 u4_sll_482_M1_2_28 ( .A(u4_sll_482_ML_int_2__28_), .B(
        u4_sll_482_ML_int_2__24_), .S(u4_sll_482_n39), .Z(
        u4_sll_482_ML_int_3__28_) );
  MUX2_X2 u4_sll_482_M1_2_36 ( .A(u4_sll_482_ML_int_2__36_), .B(
        u4_sll_482_ML_int_2__32_), .S(u4_sll_482_n39), .Z(
        u4_sll_482_ML_int_3__36_) );
  MUX2_X2 u4_sll_482_M1_2_44 ( .A(u4_sll_482_ML_int_2__44_), .B(
        u4_sll_482_ML_int_2__40_), .S(u4_sll_482_n31), .Z(
        u4_sll_482_ML_int_3__44_) );
  MUX2_X2 u4_sll_482_M1_2_52 ( .A(u4_sll_482_ML_int_2__52_), .B(
        u4_sll_482_ML_int_2__48_), .S(u4_sll_482_n39), .Z(
        u4_sll_482_ML_int_3__52_) );
  MUX2_X2 u4_sll_482_M1_2_60 ( .A(u4_sll_482_ML_int_2__60_), .B(
        u4_sll_482_ML_int_2__56_), .S(u4_sll_482_n38), .Z(
        u4_sll_482_ML_int_3__60_) );
  MUX2_X2 u4_sll_482_M1_2_68 ( .A(u4_sll_482_ML_int_2__68_), .B(
        u4_sll_482_ML_int_2__64_), .S(u4_sll_482_n38), .Z(
        u4_sll_482_ML_int_3__68_) );
  MUX2_X2 u4_sll_482_M1_2_76 ( .A(u4_sll_482_ML_int_2__76_), .B(
        u4_sll_482_ML_int_2__72_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_3__76_) );
  MUX2_X2 u4_sll_482_M1_2_84 ( .A(u4_sll_482_ML_int_2__84_), .B(
        u4_sll_482_ML_int_2__80_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_3__84_) );
  MUX2_X2 u4_sll_482_M1_2_92 ( .A(u4_sll_482_ML_int_2__92_), .B(
        u4_sll_482_ML_int_2__88_), .S(u4_sll_482_n33), .Z(
        u4_sll_482_ML_int_3__92_) );
  MUX2_X2 u4_sll_482_M1_2_100 ( .A(u4_sll_482_ML_int_2__100_), .B(
        u4_sll_482_ML_int_2__96_), .S(u4_sll_482_n33), .Z(
        u4_sll_482_ML_int_3__100_) );
  MUX2_X2 u4_sll_482_M1_2_108 ( .A(u4_sll_482_ML_int_2__108_), .B(
        u4_sll_482_ML_int_2__104_), .S(u4_sll_482_n30), .Z(
        u4_sll_482_ML_int_3__108_) );
  MUX2_X2 u4_sll_482_M1_3_12 ( .A(u4_sll_482_ML_int_3__12_), .B(
        u4_sll_482_ML_int_3__4_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_4__12_) );
  MUX2_X2 u4_sll_482_M1_3_28 ( .A(u4_sll_482_ML_int_3__28_), .B(
        u4_sll_482_ML_int_3__20_), .S(u4_sll_482_n43), .Z(
        u4_sll_482_ML_int_4__28_) );
  MUX2_X2 u4_sll_482_M1_3_44 ( .A(u4_sll_482_ML_int_3__44_), .B(
        u4_sll_482_ML_int_3__36_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_4__44_) );
  MUX2_X2 u4_sll_482_M1_3_60 ( .A(u4_sll_482_ML_int_3__60_), .B(
        u4_sll_482_ML_int_3__52_), .S(u4_sll_482_n43), .Z(
        u4_sll_482_ML_int_4__60_) );
  MUX2_X2 u4_sll_482_M1_3_76 ( .A(u4_sll_482_ML_int_3__76_), .B(
        u4_sll_482_ML_int_3__68_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_4__76_) );
  MUX2_X2 u4_sll_482_M1_3_92 ( .A(u4_sll_482_ML_int_3__92_), .B(
        u4_sll_482_ML_int_3__84_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_4__92_) );
  MUX2_X2 u4_sll_482_M1_3_108 ( .A(u4_sll_482_ML_int_3__108_), .B(
        u4_sll_482_ML_int_3__100_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_4__108_) );
  MUX2_X2 u4_sll_482_M1_4_44 ( .A(u4_sll_482_ML_int_4__44_), .B(
        u4_sll_482_ML_int_4__28_), .S(u4_sll_482_n45), .Z(
        u4_sll_482_ML_int_5__44_) );
  MUX2_X2 u4_sll_482_M1_4_76 ( .A(u4_sll_482_ML_int_4__76_), .B(
        u4_sll_482_ML_int_4__60_), .S(u4_sll_482_n45), .Z(
        u4_sll_482_ML_int_5__76_) );
  MUX2_X2 u4_sll_482_M1_4_108 ( .A(u4_sll_482_ML_int_4__108_), .B(
        u4_sll_482_ML_int_4__92_), .S(u4_sll_482_n45), .Z(
        u4_sll_482_ML_int_5__108_) );
  MUX2_X2 u4_sll_482_M1_5_44 ( .A(u4_sll_482_ML_int_5__44_), .B(
        u4_sll_482_ML_int_5__12_), .S(u4_sll_482_n47), .Z(
        u4_sll_482_ML_int_6__44_) );
  MUX2_X2 u4_sll_482_M1_5_108 ( .A(u4_sll_482_ML_int_5__108_), .B(
        u4_sll_482_ML_int_5__76_), .S(u4_sll_482_n47), .Z(
        u4_sll_482_ML_int_6__108_) );
  MUX2_X2 u4_sll_482_M1_6_108 ( .A(u4_sll_482_ML_int_6__108_), .B(
        u4_sll_482_ML_int_6__44_), .S(u4_sll_482_n48), .Z(
        u4_sll_482_ML_int_7__108_) );
  INV_X4 u4_add_489_U8 ( .A(u4_add_489__UDW__88319_net67884), .ZN(
        u4_ldz_all_0_) );
  NAND2_X2 u4_add_489_U7 ( .A1(u4_fi_ldz_5_), .A2(u4_add_489_carry_5_), .ZN(
        u4_add_489__UDW__88324_net67896) );
  INV_X4 u4_add_489_U6 ( .A(u4_add_489__UDW__88324_net67898), .ZN(
        u4_ldz_all_5_) );
  XNOR2_X2 u4_add_489_U5 ( .A(u4_fi_ldz_5_), .B(u4_add_489_carry_5_), .ZN(
        u4_add_489__UDW__88324_net67898) );
  XNOR2_X1 u4_add_489_U4 ( .A(net87917), .B(div_opa_ldz_r2[0]), .ZN(
        u4_add_489__UDW__88319_net67884) );
  INV_X4 u4_add_489_U3 ( .A(u4_add_489_n2), .ZN(u4_add_489_carry_1_) );
  NAND2_X4 u4_add_489_U2 ( .A1(net87917), .A2(div_opa_ldz_r2[0]), .ZN(
        u4_add_489_n2) );
  XNOR2_X2 u4_add_489_U1 ( .A(n4276), .B(u4_add_489__UDW__88324_net67896), 
        .ZN(u4_ldz_all_6_) );
  FA_X1 u4_add_489_U1_4 ( .A(div_opa_ldz_r2[4]), .B(u4_fi_ldz_4_), .CI(
        u4_add_489_carry_4_), .CO(u4_add_489_carry_5_), .S(u4_ldz_all_4_) );
  FA_X1 u4_add_489_U1_3 ( .A(div_opa_ldz_r2[3]), .B(u4_fi_ldz_3_), .CI(
        u4_add_489_carry_3_), .CO(u4_add_489_carry_4_), .S(u4_ldz_all_3_) );
  FA_X1 u4_add_489_U1_2 ( .A(div_opa_ldz_r2[2]), .B(u4_fi_ldz_2_), .CI(
        u4_add_489_carry_2_), .CO(u4_add_489_carry_3_), .S(u4_ldz_all_2_) );
  FA_X1 u4_add_489_U1_1 ( .A(div_opa_ldz_r2[1]), .B(u4_fi_ldz_1_), .CI(
        u4_add_489_carry_1_), .CO(u4_add_489_carry_2_), .S(u4_ldz_all_1_) );
  INV_X4 u4_add_466_U1 ( .A(net66839), .ZN(u4_exp_in_pl1_0_) );
  HA_X1 u4_add_466_U1_1_1 ( .A(n4852), .B(net66839), .CO(u4_add_466_carry[2]), 
        .S(u4_exp_in_pl1_1_) );
  HA_X1 u4_add_466_U1_1_2 ( .A(n4851), .B(u4_add_466_carry[2]), .CO(
        u4_add_466_carry[3]), .S(u4_exp_in_pl1_2_) );
  HA_X1 u4_add_466_U1_1_3 ( .A(net66851), .B(u4_add_466_carry[3]), .CO(
        u4_add_466_carry[4]), .S(u4_exp_in_pl1_3_) );
  HA_X1 u4_add_466_U1_1_4 ( .A(n4850), .B(u4_add_466_carry[4]), .CO(
        u4_add_466_carry[5]), .S(u4_exp_in_pl1_4_) );
  HA_X1 u4_add_466_U1_1_5 ( .A(exp_r[5]), .B(u4_add_466_carry[5]), .CO(
        u4_add_466_carry[6]), .S(u4_exp_in_pl1_5_) );
  HA_X1 u4_add_466_U1_1_6 ( .A(n4848), .B(u4_add_466_carry[6]), .CO(
        u4_add_466_carry[7]), .S(u4_exp_in_pl1_6_) );
  HA_X1 u4_add_466_U1_1_7 ( .A(net66863), .B(u4_add_466_carry[7]), .CO(
        u4_add_466_carry[8]), .S(u4_exp_in_pl1_7_) );
  HA_X1 u4_add_466_U1_1_8 ( .A(n4846), .B(u4_add_466_carry[8]), .CO(
        u4_add_466_carry[9]), .S(u4_exp_in_pl1_8_) );
  HA_X1 u4_add_466_U1_1_9 ( .A(net66871), .B(u4_add_466_carry[9]), .CO(
        u4_add_466_carry[10]), .S(u4_exp_in_pl1_9_) );
  HA_X1 u4_add_466_U1_1_10 ( .A(net66875), .B(u4_add_466_carry[10]), .CO(
        u4_exp_in_pl1_11_), .S(u4_exp_in_pl1_10_) );
  INV_X4 u4_add_494_U9 ( .A(u4_add_494_n7), .ZN(u4_add_494_carry_9_) );
  NAND2_X2 u4_add_494_U8 ( .A1(u4_exp_in_mi1_8_), .A2(u4_add_494_carry_8_), 
        .ZN(u4_add_494_n7) );
  INV_X4 u4_add_494_U7 ( .A(u4_add_494_n6), .ZN(u4_add_494_carry_10_) );
  NAND2_X2 u4_add_494_U6 ( .A1(u4_exp_in_mi1_9_), .A2(u4_add_494_carry_9_), 
        .ZN(u4_add_494_n6) );
  XOR2_X1 u4_add_494_U5 ( .A(n4526), .B(net43686), .Z(u4_div_exp1_0_) );
  XOR2_X2 u4_add_494_U4 ( .A(u4_exp_in_mi1_9_), .B(u4_add_494_carry_9_), .Z(
        u4_div_exp1_9_) );
  AND2_X2 u4_add_494_U3 ( .A1(n4526), .A2(net43686), .ZN(u4_add_494_n3) );
  XOR2_X2 u4_add_494_U2 ( .A(u4_exp_in_mi1_10_), .B(u4_add_494_carry_10_), .Z(
        u4_div_exp1_10_) );
  XOR2_X2 u4_add_494_U1 ( .A(u4_exp_in_mi1_8_), .B(u4_add_494_carry_8_), .Z(
        u4_div_exp1_8_) );
  FA_X1 u4_add_494_U1_1 ( .A(u4_exp_in_mi1_1_), .B(n7207), .CI(u4_add_494_n3), 
        .CO(u4_add_494_carry_2_), .S(u4_div_exp1_1_) );
  FA_X1 u4_add_494_U1_2 ( .A(u4_exp_in_mi1_2_), .B(u4_fi_ldz_2a_2_), .CI(
        u4_add_494_carry_2_), .CO(u4_add_494_carry_3_), .S(u4_div_exp1_2_) );
  FA_X1 u4_add_494_U1_3 ( .A(u4_exp_in_mi1_3_), .B(net44706), .CI(
        u4_add_494_carry_3_), .CO(u4_add_494_carry_4_), .S(u4_div_exp1_3_) );
  FA_X1 u4_add_494_U1_4 ( .A(u4_exp_in_mi1_4_), .B(u4_fi_ldz_2a_4_), .CI(
        u4_add_494_carry_4_), .CO(u4_add_494_carry_5_), .S(u4_div_exp1_4_) );
  FA_X1 u4_add_494_U1_5 ( .A(n4385), .B(u4_fi_ldz_2a_5_), .CI(
        u4_add_494_carry_5_), .CO(u4_add_494_carry_6_), .S(u4_div_exp1_5_) );
  FA_X1 u4_add_494_U1_6 ( .A(u4_exp_in_mi1_6_), .B(u4_fi_ldz_2a_6_), .CI(
        u4_add_494_carry_6_), .CO(u4_add_494_carry_7_), .S(u4_div_exp1_6_) );
  FA_X1 u4_add_494_U1_7 ( .A(u4_exp_in_mi1_7_), .B(u4_fi_ldz_2a_6_), .CI(
        u4_add_494_carry_7_), .CO(u4_add_494_carry_8_), .S(u4_div_exp1_7_) );
  INV_X4 u3_sub_63_U61 ( .A(fractb[55]), .ZN(u3_sub_63_n59) );
  INV_X4 u3_sub_63_U60 ( .A(fractb[54]), .ZN(u3_sub_63_n58) );
  INV_X4 u3_sub_63_U59 ( .A(fractb[53]), .ZN(u3_sub_63_n57) );
  INV_X4 u3_sub_63_U58 ( .A(fractb[52]), .ZN(u3_sub_63_n56) );
  INV_X4 u3_sub_63_U57 ( .A(fractb[51]), .ZN(u3_sub_63_n55) );
  INV_X4 u3_sub_63_U56 ( .A(fractb[50]), .ZN(u3_sub_63_n54) );
  INV_X4 u3_sub_63_U55 ( .A(fractb[49]), .ZN(u3_sub_63_n53) );
  INV_X4 u3_sub_63_U54 ( .A(fractb[48]), .ZN(u3_sub_63_n52) );
  INV_X4 u3_sub_63_U53 ( .A(fractb[47]), .ZN(u3_sub_63_n51) );
  INV_X4 u3_sub_63_U52 ( .A(fractb[46]), .ZN(u3_sub_63_n50) );
  INV_X4 u3_sub_63_U51 ( .A(fractb[45]), .ZN(u3_sub_63_n49) );
  INV_X4 u3_sub_63_U50 ( .A(fractb[44]), .ZN(u3_sub_63_n48) );
  INV_X4 u3_sub_63_U49 ( .A(fractb[43]), .ZN(u3_sub_63_n47) );
  INV_X4 u3_sub_63_U48 ( .A(fractb[42]), .ZN(u3_sub_63_n46) );
  INV_X4 u3_sub_63_U47 ( .A(fractb[41]), .ZN(u3_sub_63_n45) );
  INV_X4 u3_sub_63_U46 ( .A(fractb[40]), .ZN(u3_sub_63_n44) );
  INV_X4 u3_sub_63_U45 ( .A(fractb[39]), .ZN(u3_sub_63_n43) );
  INV_X4 u3_sub_63_U44 ( .A(fractb[38]), .ZN(u3_sub_63_n42) );
  INV_X4 u3_sub_63_U43 ( .A(fractb[37]), .ZN(u3_sub_63_n41) );
  INV_X4 u3_sub_63_U42 ( .A(fractb[36]), .ZN(u3_sub_63_n40) );
  INV_X4 u3_sub_63_U41 ( .A(fractb[35]), .ZN(u3_sub_63_n39) );
  INV_X4 u3_sub_63_U40 ( .A(fractb[34]), .ZN(u3_sub_63_n38) );
  INV_X4 u3_sub_63_U39 ( .A(fractb[33]), .ZN(u3_sub_63_n37) );
  INV_X4 u3_sub_63_U38 ( .A(fractb[32]), .ZN(u3_sub_63_n36) );
  INV_X4 u3_sub_63_U37 ( .A(fractb[31]), .ZN(u3_sub_63_n35) );
  INV_X4 u3_sub_63_U36 ( .A(fractb[30]), .ZN(u3_sub_63_n34) );
  INV_X4 u3_sub_63_U35 ( .A(fractb[29]), .ZN(u3_sub_63_n33) );
  INV_X4 u3_sub_63_U34 ( .A(fractb[28]), .ZN(u3_sub_63_n32) );
  INV_X4 u3_sub_63_U33 ( .A(fractb[27]), .ZN(u3_sub_63_n31) );
  INV_X4 u3_sub_63_U32 ( .A(fractb[26]), .ZN(u3_sub_63_n30) );
  INV_X4 u3_sub_63_U31 ( .A(fractb[25]), .ZN(u3_sub_63_n29) );
  INV_X4 u3_sub_63_U30 ( .A(fractb[24]), .ZN(u3_sub_63_n28) );
  INV_X4 u3_sub_63_U29 ( .A(fractb[23]), .ZN(u3_sub_63_n27) );
  INV_X4 u3_sub_63_U28 ( .A(fractb[22]), .ZN(u3_sub_63_n26) );
  INV_X4 u3_sub_63_U27 ( .A(fractb[21]), .ZN(u3_sub_63_n25) );
  INV_X4 u3_sub_63_U26 ( .A(fractb[20]), .ZN(u3_sub_63_n24) );
  INV_X4 u3_sub_63_U25 ( .A(fractb[19]), .ZN(u3_sub_63_n23) );
  INV_X4 u3_sub_63_U24 ( .A(fractb[18]), .ZN(u3_sub_63_n22) );
  INV_X4 u3_sub_63_U23 ( .A(fractb[17]), .ZN(u3_sub_63_n21) );
  INV_X4 u3_sub_63_U22 ( .A(fractb[16]), .ZN(u3_sub_63_n20) );
  INV_X4 u3_sub_63_U21 ( .A(fractb[15]), .ZN(u3_sub_63_n19) );
  INV_X4 u3_sub_63_U20 ( .A(fractb[14]), .ZN(u3_sub_63_n18) );
  INV_X4 u3_sub_63_U19 ( .A(fractb[13]), .ZN(u3_sub_63_n17) );
  INV_X4 u3_sub_63_U18 ( .A(fractb[12]), .ZN(u3_sub_63_n16) );
  INV_X4 u3_sub_63_U17 ( .A(fractb[11]), .ZN(u3_sub_63_n15) );
  INV_X4 u3_sub_63_U16 ( .A(fractb[10]), .ZN(u3_sub_63_n14) );
  INV_X4 u3_sub_63_U15 ( .A(fractb[9]), .ZN(u3_sub_63_n13) );
  INV_X4 u3_sub_63_U14 ( .A(fractb[8]), .ZN(u3_sub_63_n12) );
  INV_X4 u3_sub_63_U13 ( .A(fractb[7]), .ZN(u3_sub_63_n11) );
  INV_X4 u3_sub_63_U12 ( .A(fractb[6]), .ZN(u3_sub_63_n10) );
  INV_X4 u3_sub_63_U11 ( .A(fractb[5]), .ZN(u3_sub_63_n9) );
  INV_X4 u3_sub_63_U10 ( .A(fractb[4]), .ZN(u3_sub_63_n8) );
  INV_X4 u3_sub_63_U9 ( .A(fractb[3]), .ZN(u3_sub_63_n7) );
  INV_X4 u3_sub_63_U8 ( .A(fractb[2]), .ZN(u3_sub_63_n6) );
  INV_X4 u3_sub_63_U7 ( .A(fractb[1]), .ZN(u3_sub_63_n5) );
  INV_X4 u3_sub_63_U6 ( .A(fractb[0]), .ZN(u3_sub_63_n4) );
  INV_X4 u3_sub_63_U5 ( .A(u3_sub_63_carry[56]), .ZN(u3_N116) );
  INV_X4 u3_sub_63_U4 ( .A(fracta[0]), .ZN(u3_sub_63_n2) );
  INV_X4 u3_sub_63_U3 ( .A(u3_sub_63_n4), .ZN(u3_sub_63_n1) );
  XNOR2_X2 u3_sub_63_U2 ( .A(u3_sub_63_n4), .B(fracta[0]), .ZN(u3_N60) );
  NAND2_X2 u3_sub_63_U1 ( .A1(u3_sub_63_n1), .A2(u3_sub_63_n2), .ZN(
        u3_sub_63_carry[1]) );
  FA_X1 u3_sub_63_U2_1 ( .A(fracta[1]), .B(u3_sub_63_n5), .CI(
        u3_sub_63_carry[1]), .CO(u3_sub_63_carry[2]), .S(u3_N61) );
  FA_X1 u3_sub_63_U2_2 ( .A(fracta[2]), .B(u3_sub_63_n6), .CI(
        u3_sub_63_carry[2]), .CO(u3_sub_63_carry[3]), .S(u3_N62) );
  FA_X1 u3_sub_63_U2_3 ( .A(fracta[3]), .B(u3_sub_63_n7), .CI(
        u3_sub_63_carry[3]), .CO(u3_sub_63_carry[4]), .S(u3_N63) );
  FA_X1 u3_sub_63_U2_4 ( .A(fracta[4]), .B(u3_sub_63_n8), .CI(
        u3_sub_63_carry[4]), .CO(u3_sub_63_carry[5]), .S(u3_N64) );
  FA_X1 u3_sub_63_U2_5 ( .A(fracta[5]), .B(u3_sub_63_n9), .CI(
        u3_sub_63_carry[5]), .CO(u3_sub_63_carry[6]), .S(u3_N65) );
  FA_X1 u3_sub_63_U2_6 ( .A(fracta[6]), .B(u3_sub_63_n10), .CI(
        u3_sub_63_carry[6]), .CO(u3_sub_63_carry[7]), .S(u3_N66) );
  FA_X1 u3_sub_63_U2_7 ( .A(fracta[7]), .B(u3_sub_63_n11), .CI(
        u3_sub_63_carry[7]), .CO(u3_sub_63_carry[8]), .S(u3_N67) );
  FA_X1 u3_sub_63_U2_8 ( .A(fracta[8]), .B(u3_sub_63_n12), .CI(
        u3_sub_63_carry[8]), .CO(u3_sub_63_carry[9]), .S(u3_N68) );
  FA_X1 u3_sub_63_U2_9 ( .A(fracta[9]), .B(u3_sub_63_n13), .CI(
        u3_sub_63_carry[9]), .CO(u3_sub_63_carry[10]), .S(u3_N69) );
  FA_X1 u3_sub_63_U2_10 ( .A(fracta[10]), .B(u3_sub_63_n14), .CI(
        u3_sub_63_carry[10]), .CO(u3_sub_63_carry[11]), .S(u3_N70) );
  FA_X1 u3_sub_63_U2_11 ( .A(fracta[11]), .B(u3_sub_63_n15), .CI(
        u3_sub_63_carry[11]), .CO(u3_sub_63_carry[12]), .S(u3_N71) );
  FA_X1 u3_sub_63_U2_12 ( .A(fracta[12]), .B(u3_sub_63_n16), .CI(
        u3_sub_63_carry[12]), .CO(u3_sub_63_carry[13]), .S(u3_N72) );
  FA_X1 u3_sub_63_U2_13 ( .A(fracta[13]), .B(u3_sub_63_n17), .CI(
        u3_sub_63_carry[13]), .CO(u3_sub_63_carry[14]), .S(u3_N73) );
  FA_X1 u3_sub_63_U2_14 ( .A(fracta[14]), .B(u3_sub_63_n18), .CI(
        u3_sub_63_carry[14]), .CO(u3_sub_63_carry[15]), .S(u3_N74) );
  FA_X1 u3_sub_63_U2_15 ( .A(fracta[15]), .B(u3_sub_63_n19), .CI(
        u3_sub_63_carry[15]), .CO(u3_sub_63_carry[16]), .S(u3_N75) );
  FA_X1 u3_sub_63_U2_16 ( .A(fracta[16]), .B(u3_sub_63_n20), .CI(
        u3_sub_63_carry[16]), .CO(u3_sub_63_carry[17]), .S(u3_N76) );
  FA_X1 u3_sub_63_U2_17 ( .A(fracta[17]), .B(u3_sub_63_n21), .CI(
        u3_sub_63_carry[17]), .CO(u3_sub_63_carry[18]), .S(u3_N77) );
  FA_X1 u3_sub_63_U2_18 ( .A(fracta[18]), .B(u3_sub_63_n22), .CI(
        u3_sub_63_carry[18]), .CO(u3_sub_63_carry[19]), .S(u3_N78) );
  FA_X1 u3_sub_63_U2_19 ( .A(fracta[19]), .B(u3_sub_63_n23), .CI(
        u3_sub_63_carry[19]), .CO(u3_sub_63_carry[20]), .S(u3_N79) );
  FA_X1 u3_sub_63_U2_20 ( .A(fracta[20]), .B(u3_sub_63_n24), .CI(
        u3_sub_63_carry[20]), .CO(u3_sub_63_carry[21]), .S(u3_N80) );
  FA_X1 u3_sub_63_U2_21 ( .A(fracta[21]), .B(u3_sub_63_n25), .CI(
        u3_sub_63_carry[21]), .CO(u3_sub_63_carry[22]), .S(u3_N81) );
  FA_X1 u3_sub_63_U2_22 ( .A(fracta[22]), .B(u3_sub_63_n26), .CI(
        u3_sub_63_carry[22]), .CO(u3_sub_63_carry[23]), .S(u3_N82) );
  FA_X1 u3_sub_63_U2_23 ( .A(fracta[23]), .B(u3_sub_63_n27), .CI(
        u3_sub_63_carry[23]), .CO(u3_sub_63_carry[24]), .S(u3_N83) );
  FA_X1 u3_sub_63_U2_24 ( .A(fracta[24]), .B(u3_sub_63_n28), .CI(
        u3_sub_63_carry[24]), .CO(u3_sub_63_carry[25]), .S(u3_N84) );
  FA_X1 u3_sub_63_U2_25 ( .A(fracta[25]), .B(u3_sub_63_n29), .CI(
        u3_sub_63_carry[25]), .CO(u3_sub_63_carry[26]), .S(u3_N85) );
  FA_X1 u3_sub_63_U2_26 ( .A(fracta[26]), .B(u3_sub_63_n30), .CI(
        u3_sub_63_carry[26]), .CO(u3_sub_63_carry[27]), .S(u3_N86) );
  FA_X1 u3_sub_63_U2_27 ( .A(fracta[27]), .B(u3_sub_63_n31), .CI(
        u3_sub_63_carry[27]), .CO(u3_sub_63_carry[28]), .S(u3_N87) );
  FA_X1 u3_sub_63_U2_28 ( .A(fracta[28]), .B(u3_sub_63_n32), .CI(
        u3_sub_63_carry[28]), .CO(u3_sub_63_carry[29]), .S(u3_N88) );
  FA_X1 u3_sub_63_U2_29 ( .A(fracta[29]), .B(u3_sub_63_n33), .CI(
        u3_sub_63_carry[29]), .CO(u3_sub_63_carry[30]), .S(u3_N89) );
  FA_X1 u3_sub_63_U2_30 ( .A(fracta[30]), .B(u3_sub_63_n34), .CI(
        u3_sub_63_carry[30]), .CO(u3_sub_63_carry[31]), .S(u3_N90) );
  FA_X1 u3_sub_63_U2_31 ( .A(fracta[31]), .B(u3_sub_63_n35), .CI(
        u3_sub_63_carry[31]), .CO(u3_sub_63_carry[32]), .S(u3_N91) );
  FA_X1 u3_sub_63_U2_32 ( .A(fracta[32]), .B(u3_sub_63_n36), .CI(
        u3_sub_63_carry[32]), .CO(u3_sub_63_carry[33]), .S(u3_N92) );
  FA_X1 u3_sub_63_U2_33 ( .A(fracta[33]), .B(u3_sub_63_n37), .CI(
        u3_sub_63_carry[33]), .CO(u3_sub_63_carry[34]), .S(u3_N93) );
  FA_X1 u3_sub_63_U2_34 ( .A(fracta[34]), .B(u3_sub_63_n38), .CI(
        u3_sub_63_carry[34]), .CO(u3_sub_63_carry[35]), .S(u3_N94) );
  FA_X1 u3_sub_63_U2_35 ( .A(fracta[35]), .B(u3_sub_63_n39), .CI(
        u3_sub_63_carry[35]), .CO(u3_sub_63_carry[36]), .S(u3_N95) );
  FA_X1 u3_sub_63_U2_36 ( .A(fracta[36]), .B(u3_sub_63_n40), .CI(
        u3_sub_63_carry[36]), .CO(u3_sub_63_carry[37]), .S(u3_N96) );
  FA_X1 u3_sub_63_U2_37 ( .A(fracta[37]), .B(u3_sub_63_n41), .CI(
        u3_sub_63_carry[37]), .CO(u3_sub_63_carry[38]), .S(u3_N97) );
  FA_X1 u3_sub_63_U2_38 ( .A(fracta[38]), .B(u3_sub_63_n42), .CI(
        u3_sub_63_carry[38]), .CO(u3_sub_63_carry[39]), .S(u3_N98) );
  FA_X1 u3_sub_63_U2_39 ( .A(fracta[39]), .B(u3_sub_63_n43), .CI(
        u3_sub_63_carry[39]), .CO(u3_sub_63_carry[40]), .S(u3_N99) );
  FA_X1 u3_sub_63_U2_40 ( .A(fracta[40]), .B(u3_sub_63_n44), .CI(
        u3_sub_63_carry[40]), .CO(u3_sub_63_carry[41]), .S(u3_N100) );
  FA_X1 u3_sub_63_U2_41 ( .A(fracta[41]), .B(u3_sub_63_n45), .CI(
        u3_sub_63_carry[41]), .CO(u3_sub_63_carry[42]), .S(u3_N101) );
  FA_X1 u3_sub_63_U2_42 ( .A(fracta[42]), .B(u3_sub_63_n46), .CI(
        u3_sub_63_carry[42]), .CO(u3_sub_63_carry[43]), .S(u3_N102) );
  FA_X1 u3_sub_63_U2_43 ( .A(fracta[43]), .B(u3_sub_63_n47), .CI(
        u3_sub_63_carry[43]), .CO(u3_sub_63_carry[44]), .S(u3_N103) );
  FA_X1 u3_sub_63_U2_44 ( .A(fracta[44]), .B(u3_sub_63_n48), .CI(
        u3_sub_63_carry[44]), .CO(u3_sub_63_carry[45]), .S(u3_N104) );
  FA_X1 u3_sub_63_U2_45 ( .A(fracta[45]), .B(u3_sub_63_n49), .CI(
        u3_sub_63_carry[45]), .CO(u3_sub_63_carry[46]), .S(u3_N105) );
  FA_X1 u3_sub_63_U2_46 ( .A(fracta[46]), .B(u3_sub_63_n50), .CI(
        u3_sub_63_carry[46]), .CO(u3_sub_63_carry[47]), .S(u3_N106) );
  FA_X1 u3_sub_63_U2_47 ( .A(fracta[47]), .B(u3_sub_63_n51), .CI(
        u3_sub_63_carry[47]), .CO(u3_sub_63_carry[48]), .S(u3_N107) );
  FA_X1 u3_sub_63_U2_48 ( .A(fracta[48]), .B(u3_sub_63_n52), .CI(
        u3_sub_63_carry[48]), .CO(u3_sub_63_carry[49]), .S(u3_N108) );
  FA_X1 u3_sub_63_U2_49 ( .A(fracta[49]), .B(u3_sub_63_n53), .CI(
        u3_sub_63_carry[49]), .CO(u3_sub_63_carry[50]), .S(u3_N109) );
  FA_X1 u3_sub_63_U2_50 ( .A(fracta[50]), .B(u3_sub_63_n54), .CI(
        u3_sub_63_carry[50]), .CO(u3_sub_63_carry[51]), .S(u3_N110) );
  FA_X1 u3_sub_63_U2_51 ( .A(fracta[51]), .B(u3_sub_63_n55), .CI(
        u3_sub_63_carry[51]), .CO(u3_sub_63_carry[52]), .S(u3_N111) );
  FA_X1 u3_sub_63_U2_52 ( .A(fracta[52]), .B(u3_sub_63_n56), .CI(
        u3_sub_63_carry[52]), .CO(u3_sub_63_carry[53]), .S(u3_N112) );
  FA_X1 u3_sub_63_U2_53 ( .A(fracta[53]), .B(u3_sub_63_n57), .CI(
        u3_sub_63_carry[53]), .CO(u3_sub_63_carry[54]), .S(u3_N113) );
  FA_X1 u3_sub_63_U2_54 ( .A(fracta[54]), .B(u3_sub_63_n58), .CI(
        u3_sub_63_carry[54]), .CO(u3_sub_63_carry[55]), .S(u3_N114) );
  FA_X1 u3_sub_63_U2_55 ( .A(fracta[55]), .B(u3_sub_63_n59), .CI(
        u3_sub_63_carry[55]), .CO(u3_sub_63_carry[56]), .S(u3_N115) );
  INV_X4 u3_add_63_U3 ( .A(u3_add_63_n2), .ZN(u3_add_63_carry[1]) );
  NAND2_X2 u3_add_63_U2 ( .A1(fractb[0]), .A2(fracta[0]), .ZN(u3_add_63_n2) );
  XOR2_X1 u3_add_63_U1 ( .A(fractb[0]), .B(fracta[0]), .Z(u3_N3) );
  FA_X1 u3_add_63_U1_1 ( .A(fracta[1]), .B(fractb[1]), .CI(u3_add_63_carry[1]), 
        .CO(u3_add_63_carry[2]), .S(u3_N4) );
  FA_X1 u3_add_63_U1_2 ( .A(fracta[2]), .B(fractb[2]), .CI(u3_add_63_carry[2]), 
        .CO(u3_add_63_carry[3]), .S(u3_N5) );
  FA_X1 u3_add_63_U1_3 ( .A(fracta[3]), .B(fractb[3]), .CI(u3_add_63_carry[3]), 
        .CO(u3_add_63_carry[4]), .S(u3_N6) );
  FA_X1 u3_add_63_U1_4 ( .A(fracta[4]), .B(fractb[4]), .CI(u3_add_63_carry[4]), 
        .CO(u3_add_63_carry[5]), .S(u3_N7) );
  FA_X1 u3_add_63_U1_5 ( .A(fracta[5]), .B(fractb[5]), .CI(u3_add_63_carry[5]), 
        .CO(u3_add_63_carry[6]), .S(u3_N8) );
  FA_X1 u3_add_63_U1_6 ( .A(fracta[6]), .B(fractb[6]), .CI(u3_add_63_carry[6]), 
        .CO(u3_add_63_carry[7]), .S(u3_N9) );
  FA_X1 u3_add_63_U1_7 ( .A(fracta[7]), .B(fractb[7]), .CI(u3_add_63_carry[7]), 
        .CO(u3_add_63_carry[8]), .S(u3_N10) );
  FA_X1 u3_add_63_U1_8 ( .A(fracta[8]), .B(fractb[8]), .CI(u3_add_63_carry[8]), 
        .CO(u3_add_63_carry[9]), .S(u3_N11) );
  FA_X1 u3_add_63_U1_9 ( .A(fracta[9]), .B(fractb[9]), .CI(u3_add_63_carry[9]), 
        .CO(u3_add_63_carry[10]), .S(u3_N12) );
  FA_X1 u3_add_63_U1_10 ( .A(fracta[10]), .B(fractb[10]), .CI(
        u3_add_63_carry[10]), .CO(u3_add_63_carry[11]), .S(u3_N13) );
  FA_X1 u3_add_63_U1_11 ( .A(fracta[11]), .B(fractb[11]), .CI(
        u3_add_63_carry[11]), .CO(u3_add_63_carry[12]), .S(u3_N14) );
  FA_X1 u3_add_63_U1_12 ( .A(fracta[12]), .B(fractb[12]), .CI(
        u3_add_63_carry[12]), .CO(u3_add_63_carry[13]), .S(u3_N15) );
  FA_X1 u3_add_63_U1_13 ( .A(fracta[13]), .B(fractb[13]), .CI(
        u3_add_63_carry[13]), .CO(u3_add_63_carry[14]), .S(u3_N16) );
  FA_X1 u3_add_63_U1_14 ( .A(fracta[14]), .B(fractb[14]), .CI(
        u3_add_63_carry[14]), .CO(u3_add_63_carry[15]), .S(u3_N17) );
  FA_X1 u3_add_63_U1_15 ( .A(fracta[15]), .B(fractb[15]), .CI(
        u3_add_63_carry[15]), .CO(u3_add_63_carry[16]), .S(u3_N18) );
  FA_X1 u3_add_63_U1_16 ( .A(fracta[16]), .B(fractb[16]), .CI(
        u3_add_63_carry[16]), .CO(u3_add_63_carry[17]), .S(u3_N19) );
  FA_X1 u3_add_63_U1_17 ( .A(fracta[17]), .B(fractb[17]), .CI(
        u3_add_63_carry[17]), .CO(u3_add_63_carry[18]), .S(u3_N20) );
  FA_X1 u3_add_63_U1_18 ( .A(fracta[18]), .B(fractb[18]), .CI(
        u3_add_63_carry[18]), .CO(u3_add_63_carry[19]), .S(u3_N21) );
  FA_X1 u3_add_63_U1_19 ( .A(fracta[19]), .B(fractb[19]), .CI(
        u3_add_63_carry[19]), .CO(u3_add_63_carry[20]), .S(u3_N22) );
  FA_X1 u3_add_63_U1_20 ( .A(fracta[20]), .B(fractb[20]), .CI(
        u3_add_63_carry[20]), .CO(u3_add_63_carry[21]), .S(u3_N23) );
  FA_X1 u3_add_63_U1_21 ( .A(fracta[21]), .B(fractb[21]), .CI(
        u3_add_63_carry[21]), .CO(u3_add_63_carry[22]), .S(u3_N24) );
  FA_X1 u3_add_63_U1_22 ( .A(fracta[22]), .B(fractb[22]), .CI(
        u3_add_63_carry[22]), .CO(u3_add_63_carry[23]), .S(u3_N25) );
  FA_X1 u3_add_63_U1_23 ( .A(fracta[23]), .B(fractb[23]), .CI(
        u3_add_63_carry[23]), .CO(u3_add_63_carry[24]), .S(u3_N26) );
  FA_X1 u3_add_63_U1_24 ( .A(fracta[24]), .B(fractb[24]), .CI(
        u3_add_63_carry[24]), .CO(u3_add_63_carry[25]), .S(u3_N27) );
  FA_X1 u3_add_63_U1_25 ( .A(fracta[25]), .B(fractb[25]), .CI(
        u3_add_63_carry[25]), .CO(u3_add_63_carry[26]), .S(u3_N28) );
  FA_X1 u3_add_63_U1_26 ( .A(fracta[26]), .B(fractb[26]), .CI(
        u3_add_63_carry[26]), .CO(u3_add_63_carry[27]), .S(u3_N29) );
  FA_X1 u3_add_63_U1_27 ( .A(fracta[27]), .B(fractb[27]), .CI(
        u3_add_63_carry[27]), .CO(u3_add_63_carry[28]), .S(u3_N30) );
  FA_X1 u3_add_63_U1_28 ( .A(fracta[28]), .B(fractb[28]), .CI(
        u3_add_63_carry[28]), .CO(u3_add_63_carry[29]), .S(u3_N31) );
  FA_X1 u3_add_63_U1_29 ( .A(fracta[29]), .B(fractb[29]), .CI(
        u3_add_63_carry[29]), .CO(u3_add_63_carry[30]), .S(u3_N32) );
  FA_X1 u3_add_63_U1_30 ( .A(fracta[30]), .B(fractb[30]), .CI(
        u3_add_63_carry[30]), .CO(u3_add_63_carry[31]), .S(u3_N33) );
  FA_X1 u3_add_63_U1_31 ( .A(fracta[31]), .B(fractb[31]), .CI(
        u3_add_63_carry[31]), .CO(u3_add_63_carry[32]), .S(u3_N34) );
  FA_X1 u3_add_63_U1_32 ( .A(fracta[32]), .B(fractb[32]), .CI(
        u3_add_63_carry[32]), .CO(u3_add_63_carry[33]), .S(u3_N35) );
  FA_X1 u3_add_63_U1_33 ( .A(fracta[33]), .B(fractb[33]), .CI(
        u3_add_63_carry[33]), .CO(u3_add_63_carry[34]), .S(u3_N36) );
  FA_X1 u3_add_63_U1_34 ( .A(fracta[34]), .B(fractb[34]), .CI(
        u3_add_63_carry[34]), .CO(u3_add_63_carry[35]), .S(u3_N37) );
  FA_X1 u3_add_63_U1_35 ( .A(fracta[35]), .B(fractb[35]), .CI(
        u3_add_63_carry[35]), .CO(u3_add_63_carry[36]), .S(u3_N38) );
  FA_X1 u3_add_63_U1_36 ( .A(fracta[36]), .B(fractb[36]), .CI(
        u3_add_63_carry[36]), .CO(u3_add_63_carry[37]), .S(u3_N39) );
  FA_X1 u3_add_63_U1_37 ( .A(fracta[37]), .B(fractb[37]), .CI(
        u3_add_63_carry[37]), .CO(u3_add_63_carry[38]), .S(u3_N40) );
  FA_X1 u3_add_63_U1_38 ( .A(fracta[38]), .B(fractb[38]), .CI(
        u3_add_63_carry[38]), .CO(u3_add_63_carry[39]), .S(u3_N41) );
  FA_X1 u3_add_63_U1_39 ( .A(fracta[39]), .B(fractb[39]), .CI(
        u3_add_63_carry[39]), .CO(u3_add_63_carry[40]), .S(u3_N42) );
  FA_X1 u3_add_63_U1_40 ( .A(fracta[40]), .B(fractb[40]), .CI(
        u3_add_63_carry[40]), .CO(u3_add_63_carry[41]), .S(u3_N43) );
  FA_X1 u3_add_63_U1_41 ( .A(fracta[41]), .B(fractb[41]), .CI(
        u3_add_63_carry[41]), .CO(u3_add_63_carry[42]), .S(u3_N44) );
  FA_X1 u3_add_63_U1_42 ( .A(fracta[42]), .B(fractb[42]), .CI(
        u3_add_63_carry[42]), .CO(u3_add_63_carry[43]), .S(u3_N45) );
  FA_X1 u3_add_63_U1_43 ( .A(fracta[43]), .B(fractb[43]), .CI(
        u3_add_63_carry[43]), .CO(u3_add_63_carry[44]), .S(u3_N46) );
  FA_X1 u3_add_63_U1_44 ( .A(fracta[44]), .B(fractb[44]), .CI(
        u3_add_63_carry[44]), .CO(u3_add_63_carry[45]), .S(u3_N47) );
  FA_X1 u3_add_63_U1_45 ( .A(fracta[45]), .B(fractb[45]), .CI(
        u3_add_63_carry[45]), .CO(u3_add_63_carry[46]), .S(u3_N48) );
  FA_X1 u3_add_63_U1_46 ( .A(fracta[46]), .B(fractb[46]), .CI(
        u3_add_63_carry[46]), .CO(u3_add_63_carry[47]), .S(u3_N49) );
  FA_X1 u3_add_63_U1_47 ( .A(fracta[47]), .B(fractb[47]), .CI(
        u3_add_63_carry[47]), .CO(u3_add_63_carry[48]), .S(u3_N50) );
  FA_X1 u3_add_63_U1_48 ( .A(fracta[48]), .B(fractb[48]), .CI(
        u3_add_63_carry[48]), .CO(u3_add_63_carry[49]), .S(u3_N51) );
  FA_X1 u3_add_63_U1_49 ( .A(fracta[49]), .B(fractb[49]), .CI(
        u3_add_63_carry[49]), .CO(u3_add_63_carry[50]), .S(u3_N52) );
  FA_X1 u3_add_63_U1_50 ( .A(fracta[50]), .B(fractb[50]), .CI(
        u3_add_63_carry[50]), .CO(u3_add_63_carry[51]), .S(u3_N53) );
  FA_X1 u3_add_63_U1_51 ( .A(fracta[51]), .B(fractb[51]), .CI(
        u3_add_63_carry[51]), .CO(u3_add_63_carry[52]), .S(u3_N54) );
  FA_X1 u3_add_63_U1_52 ( .A(fracta[52]), .B(fractb[52]), .CI(
        u3_add_63_carry[52]), .CO(u3_add_63_carry[53]), .S(u3_N55) );
  FA_X1 u3_add_63_U1_53 ( .A(fracta[53]), .B(fractb[53]), .CI(
        u3_add_63_carry[53]), .CO(u3_add_63_carry[54]), .S(u3_N56) );
  FA_X1 u3_add_63_U1_54 ( .A(fracta[54]), .B(fractb[54]), .CI(
        u3_add_63_carry[54]), .CO(u3_add_63_carry[55]), .S(u3_N57) );
  FA_X1 u3_add_63_U1_55 ( .A(fracta[55]), .B(fractb[55]), .CI(
        u3_add_63_carry[55]), .CO(u3_N59), .S(u3_N58) );
  XOR2_X1 u2_add_120_U2 ( .A(u2_add_120_carry[10]), .B(u2_exp_tmp4_10_), .Z(
        u2_N64) );
  INV_X4 u2_add_120_U1 ( .A(u2_exp_tmp4_0_), .ZN(u2_N54) );
  HA_X1 u2_add_120_U1_1_1 ( .A(u2_exp_tmp4_1_), .B(u2_exp_tmp4_0_), .CO(
        u2_add_120_carry[2]), .S(u2_N55) );
  HA_X1 u2_add_120_U1_1_2 ( .A(u2_exp_tmp4_2_), .B(u2_add_120_carry[2]), .CO(
        u2_add_120_carry[3]), .S(u2_N56) );
  HA_X1 u2_add_120_U1_1_3 ( .A(u2_exp_tmp4_3_), .B(u2_add_120_carry[3]), .CO(
        u2_add_120_carry[4]), .S(u2_N57) );
  HA_X1 u2_add_120_U1_1_4 ( .A(u2_exp_tmp4_4_), .B(u2_add_120_carry[4]), .CO(
        u2_add_120_carry[5]), .S(u2_N58) );
  HA_X1 u2_add_120_U1_1_5 ( .A(u2_exp_tmp4_5_), .B(u2_add_120_carry[5]), .CO(
        u2_add_120_carry[6]), .S(u2_N59) );
  HA_X1 u2_add_120_U1_1_6 ( .A(u2_exp_tmp4_6_), .B(u2_add_120_carry[6]), .CO(
        u2_add_120_carry[7]), .S(u2_N60) );
  HA_X1 u2_add_120_U1_1_7 ( .A(u2_exp_tmp4_7_), .B(u2_add_120_carry[7]), .CO(
        u2_add_120_carry[8]), .S(u2_N61) );
  HA_X1 u2_add_120_U1_1_8 ( .A(u2_exp_tmp4_8_), .B(u2_add_120_carry[8]), .CO(
        u2_add_120_carry[9]), .S(u2_N62) );
  HA_X1 u2_add_120_U1_1_9 ( .A(u2_exp_tmp4_9_), .B(u2_add_120_carry[9]), .CO(
        u2_add_120_carry[10]), .S(u2_N63) );
  XOR2_X1 u2_add_118_U2 ( .A(u2_add_118_carry[10]), .B(n8290), .Z(
        u2_exp_tmp3_10_) );
  INV_X4 u2_add_118_U1 ( .A(u2_exp_tmp4_0_), .ZN(u2_exp_tmp3_0_) );
  HA_X1 u2_add_118_U1_1_1 ( .A(n4318), .B(u2_exp_tmp4_0_), .CO(
        u2_add_118_carry[2]), .S(u2_exp_tmp3_1_) );
  HA_X1 u2_add_118_U1_1_2 ( .A(n8298), .B(u2_add_118_carry[2]), .CO(
        u2_add_118_carry[3]), .S(u2_exp_tmp3_2_) );
  HA_X1 u2_add_118_U1_1_3 ( .A(n8297), .B(u2_add_118_carry[3]), .CO(
        u2_add_118_carry[4]), .S(u2_exp_tmp3_3_) );
  HA_X1 u2_add_118_U1_1_4 ( .A(n8296), .B(u2_add_118_carry[4]), .CO(
        u2_add_118_carry[5]), .S(u2_exp_tmp3_4_) );
  HA_X1 u2_add_118_U1_1_5 ( .A(n8295), .B(u2_add_118_carry[5]), .CO(
        u2_add_118_carry[6]), .S(u2_exp_tmp3_5_) );
  HA_X1 u2_add_118_U1_1_6 ( .A(n8294), .B(u2_add_118_carry[6]), .CO(
        u2_add_118_carry[7]), .S(u2_exp_tmp3_6_) );
  HA_X1 u2_add_118_U1_1_7 ( .A(n8293), .B(u2_add_118_carry[7]), .CO(
        u2_add_118_carry[8]), .S(u2_exp_tmp3_7_) );
  HA_X1 u2_add_118_U1_1_8 ( .A(n8292), .B(u2_add_118_carry[8]), .CO(
        u2_add_118_carry[9]), .S(u2_exp_tmp3_8_) );
  HA_X1 u2_add_118_U1_1_9 ( .A(n8291), .B(u2_add_118_carry[9]), .CO(
        u2_add_118_carry[10]), .S(u2_exp_tmp3_9_) );
  INV_X4 u2_add_115_U3 ( .A(u2_add_115_n2), .ZN(u2_add_115_carry[1]) );
  NAND2_X2 u2_add_115_U2 ( .A1(opb_r[52]), .A2(opa_r[52]), .ZN(u2_add_115_n2)
         );
  XOR2_X1 u2_add_115_U1 ( .A(opb_r[52]), .B(opa_r[52]), .Z(u2_N18) );
  FA_X1 u2_add_115_U1_1 ( .A(opa_r[53]), .B(opb_r[53]), .CI(
        u2_add_115_carry[1]), .CO(u2_add_115_carry[2]), .S(u2_N19) );
  FA_X1 u2_add_115_U1_2 ( .A(opa_r[54]), .B(opb_r[54]), .CI(
        u2_add_115_carry[2]), .CO(u2_add_115_carry[3]), .S(u2_N20) );
  FA_X1 u2_add_115_U1_3 ( .A(opa_r[55]), .B(opb_r[55]), .CI(
        u2_add_115_carry[3]), .CO(u2_add_115_carry[4]), .S(u2_N21) );
  FA_X1 u2_add_115_U1_4 ( .A(opa_r[56]), .B(n4836), .CI(u2_add_115_carry[4]), 
        .CO(u2_add_115_carry[5]), .S(u2_N22) );
  FA_X1 u2_add_115_U1_5 ( .A(opa_r[57]), .B(n4839), .CI(u2_add_115_carry[5]), 
        .CO(u2_add_115_carry[6]), .S(u2_N23) );
  FA_X1 u2_add_115_U1_6 ( .A(opa_r[58]), .B(n4425), .CI(u2_add_115_carry[6]), 
        .CO(u2_add_115_carry[7]), .S(u2_N24) );
  FA_X1 u2_add_115_U1_7 ( .A(opa_r[59]), .B(n4271), .CI(u2_add_115_carry[7]), 
        .CO(u2_add_115_carry[8]), .S(u2_N25) );
  FA_X1 u2_add_115_U1_8 ( .A(opa_r[60]), .B(n4823), .CI(u2_add_115_carry[8]), 
        .CO(u2_add_115_carry[9]), .S(u2_N26) );
  FA_X1 u2_add_115_U1_9 ( .A(opa_r[61]), .B(opb_r[61]), .CI(
        u2_add_115_carry[9]), .CO(u2_add_115_carry[10]), .S(u2_N27) );
  FA_X1 u2_add_115_U1_10 ( .A(n4853), .B(opb_r[62]), .CI(u2_add_115_carry[10]), 
        .CO(u2_N29), .S(u2_N28) );
  INV_X4 u2_sub_115_U16 ( .A(opb_r[52]), .ZN(u2_sub_115_n14) );
  INV_X4 u2_sub_115_U15 ( .A(opb_r[55]), .ZN(u2_sub_115_n11) );
  INV_X4 u2_sub_115_U14 ( .A(n4839), .ZN(u2_sub_115_n9) );
  INV_X4 u2_sub_115_U13 ( .A(opb_r[61]), .ZN(u2_sub_115_n5) );
  INV_X4 u2_sub_115_U12 ( .A(u2_sub_115_carry[11]), .ZN(u2_N17) );
  INV_X2 u2_sub_115_U11 ( .A(opb_r[62]), .ZN(u2_sub_115_n4) );
  INV_X2 u2_sub_115_U10 ( .A(n4836), .ZN(u2_sub_115_n10) );
  INV_X2 u2_sub_115_U9 ( .A(opb_r[54]), .ZN(u2_sub_115_n12) );
  INV_X2 u2_sub_115_U8 ( .A(n4823), .ZN(u2_sub_115_n6) );
  INV_X2 u2_sub_115_U7 ( .A(opb_r[53]), .ZN(u2_sub_115_n13) );
  INV_X1 u2_sub_115_U6 ( .A(n4425), .ZN(u2_sub_115_n8) );
  INV_X4 u2_sub_115_U5 ( .A(opa_r[52]), .ZN(u2_sub_115_n2) );
  INV_X4 u2_sub_115_U4 ( .A(u2_sub_115_n14), .ZN(u2_sub_115_n1) );
  XNOR2_X2 u2_sub_115_U3 ( .A(u2_sub_115_n14), .B(opa_r[52]), .ZN(u2_N6) );
  NAND2_X2 u2_sub_115_U2 ( .A1(u2_sub_115_n1), .A2(u2_sub_115_n2), .ZN(
        u2_sub_115_carry[1]) );
  INV_X1 u2_sub_115_U1 ( .A(n4837), .ZN(u2_sub_115_n7) );
  FA_X1 u2_sub_115_U2_1 ( .A(opa_r[53]), .B(u2_sub_115_n13), .CI(
        u2_sub_115_carry[1]), .CO(u2_sub_115_carry[2]), .S(u2_N7) );
  FA_X1 u2_sub_115_U2_2 ( .A(opa_r[54]), .B(u2_sub_115_n12), .CI(
        u2_sub_115_carry[2]), .CO(u2_sub_115_carry[3]), .S(u2_N8) );
  FA_X1 u2_sub_115_U2_3 ( .A(opa_r[55]), .B(u2_sub_115_n11), .CI(
        u2_sub_115_carry[3]), .CO(u2_sub_115_carry[4]), .S(u2_N9) );
  FA_X1 u2_sub_115_U2_4 ( .A(opa_r[56]), .B(u2_sub_115_n10), .CI(
        u2_sub_115_carry[4]), .CO(u2_sub_115_carry[5]), .S(u2_N10) );
  FA_X1 u2_sub_115_U2_5 ( .A(opa_r[57]), .B(u2_sub_115_n9), .CI(
        u2_sub_115_carry[5]), .CO(u2_sub_115_carry[6]), .S(u2_N11) );
  FA_X1 u2_sub_115_U2_6 ( .A(opa_r[58]), .B(u2_sub_115_n8), .CI(
        u2_sub_115_carry[6]), .CO(u2_sub_115_carry[7]), .S(u2_N12) );
  FA_X1 u2_sub_115_U2_7 ( .A(opa_r[59]), .B(u2_sub_115_n7), .CI(
        u2_sub_115_carry[7]), .CO(u2_sub_115_carry[8]), .S(u2_N13) );
  FA_X1 u2_sub_115_U2_8 ( .A(opa_r[60]), .B(u2_sub_115_n6), .CI(
        u2_sub_115_carry[8]), .CO(u2_sub_115_carry[9]), .S(u2_N14) );
  FA_X1 u2_sub_115_U2_9 ( .A(opa_r[61]), .B(u2_sub_115_n5), .CI(
        u2_sub_115_carry[9]), .CO(u2_sub_115_carry[10]), .S(u2_N15) );
  FA_X1 u2_sub_115_U2_10 ( .A(n4853), .B(u2_sub_115_n4), .CI(
        u2_sub_115_carry[10]), .CO(u2_sub_115_carry[11]), .S(u2_N16) );
  NOR2_X1 u1_srl_151_U433 ( .A1(u1_srl_151_n111), .A2(n8470), .ZN(
        u1_srl_151_n177) );
  NAND2_X1 u1_srl_151_U432 ( .A1(n8466), .A2(u1_srl_151_n107), .ZN(
        u1_srl_151_n211) );
  AOI22_X1 u1_srl_151_U431 ( .A1(u1_adj_op_28_), .A2(u1_srl_151_n17), .B1(
        n8497), .B2(u1_srl_151_n27), .ZN(u1_srl_151_n375) );
  OAI221_X1 u1_srl_151_U430 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n132), .C1(
        u1_srl_151_n14), .C2(u1_srl_151_n131), .A(u1_srl_151_n375), .ZN(
        u1_srl_151_n257) );
  AOI22_X1 u1_srl_151_U429 ( .A1(n8498), .A2(u1_srl_151_n21), .B1(
        u1_srl_151_n27), .B2(u1_adj_op_21_), .ZN(u1_srl_151_n374) );
  OAI221_X1 u1_srl_151_U428 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n136), .C1(
        u1_srl_151_n14), .C2(u1_srl_151_n135), .A(u1_srl_151_n374), .ZN(
        u1_srl_151_n258) );
  AOI22_X1 u1_srl_151_U427 ( .A1(u1_srl_151_n17), .A2(u1_adj_op_20_), .B1(
        u1_adj_op_17_), .B2(u1_srl_151_n27), .ZN(u1_srl_151_n373) );
  OAI221_X1 u1_srl_151_U426 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n141), .C1(
        u1_srl_151_n140), .C2(u1_srl_151_n14), .A(u1_srl_151_n373), .ZN(
        u1_srl_151_n167) );
  AOI22_X1 u1_srl_151_U425 ( .A1(u1_adj_op_16_), .A2(u1_srl_151_n21), .B1(
        n8504), .B2(u1_srl_151_n27), .ZN(u1_srl_151_n372) );
  OAI221_X1 u1_srl_151_U424 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n145), .C1(
        u1_srl_151_n14), .C2(u1_srl_151_n144), .A(u1_srl_151_n372), .ZN(
        u1_srl_151_n168) );
  AOI22_X1 u1_srl_151_U423 ( .A1(u1_srl_151_n13), .A2(u1_srl_151_n167), .B1(
        u1_srl_151_n31), .B2(u1_srl_151_n168), .ZN(u1_srl_151_n371) );
  AOI221_X1 u1_srl_151_U422 ( .B1(u1_srl_151_n257), .B2(u1_srl_151_n252), .C1(
        u1_srl_151_n258), .C2(u1_srl_151_n5), .A(u1_srl_151_n35), .ZN(
        u1_srl_151_n304) );
  AOI22_X1 u1_srl_151_U421 ( .A1(n8479), .A2(u1_srl_151_n21), .B1(n8500), .B2(
        u1_srl_151_n27), .ZN(u1_srl_151_n370) );
  OAI221_X1 u1_srl_151_U420 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n128), .C1(
        u1_srl_151_n14), .C2(u1_srl_151_n119), .A(u1_srl_151_n370), .ZN(
        u1_srl_151_n198) );
  AOI22_X1 u1_srl_151_U419 ( .A1(u1_adj_op_36_), .A2(u1_srl_151_n21), .B1(
        n8491), .B2(u1_srl_151_n26), .ZN(u1_srl_151_n369) );
  OAI221_X1 u1_srl_151_U418 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n123), .C1(
        u1_srl_151_n14), .C2(u1_srl_151_n122), .A(u1_srl_151_n369), .ZN(
        u1_srl_151_n260) );
  AOI22_X1 u1_srl_151_U417 ( .A1(u1_adj_op_32_), .A2(u1_srl_151_n21), .B1(
        n8495), .B2(u1_srl_151_n26), .ZN(u1_srl_151_n368) );
  OAI221_X1 u1_srl_151_U416 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n127), .C1(
        u1_srl_151_n14), .C2(u1_srl_151_n126), .A(u1_srl_151_n368), .ZN(
        u1_srl_151_n261) );
  AOI22_X1 u1_srl_151_U415 ( .A1(u1_adj_op_44_), .A2(u1_srl_151_n20), .B1(
        n8486), .B2(u1_srl_151_n26), .ZN(u1_srl_151_n367) );
  AOI221_X1 u1_srl_151_U414 ( .B1(u1_srl_151_n6), .B2(u1_adj_op_42_), .C1(
        u1_srl_151_n16), .C2(n8485), .A(u1_srl_151_n75), .ZN(u1_srl_151_n285)
         );
  AOI22_X1 u1_srl_151_U413 ( .A1(n8487), .A2(u1_srl_151_n20), .B1(
        u1_adj_op_37_), .B2(u1_srl_151_n26), .ZN(u1_srl_151_n366) );
  AOI221_X1 u1_srl_151_U412 ( .B1(u1_srl_151_n6), .B2(u1_adj_op_38_), .C1(
        u1_srl_151_n16), .C2(n8488), .A(u1_srl_151_n77), .ZN(u1_srl_151_n327)
         );
  OAI22_X1 u1_srl_151_U411 ( .A1(u1_srl_151_n72), .A2(u1_srl_151_n285), .B1(
        u1_srl_151_n4), .B2(u1_srl_151_n327), .ZN(u1_srl_151_n365) );
  AOI221_X1 u1_srl_151_U410 ( .B1(u1_srl_151_n260), .B2(u1_srl_151_n13), .C1(
        u1_srl_151_n261), .C2(u1_srl_151_n31), .A(u1_srl_151_n365), .ZN(
        u1_srl_151_n230) );
  AOI222_X1 u1_srl_151_U409 ( .A1(u1_srl_151_n177), .A2(u1_srl_151_n34), .B1(
        u1_srl_151_n153), .B2(u1_srl_151_n198), .C1(u1_srl_151_n159), .C2(
        u1_srl_151_n36), .ZN(u1_srl_151_n357) );
  NAND2_X1 u1_srl_151_U408 ( .A1(n8469), .A2(n8470), .ZN(u1_srl_151_n238) );
  AOI22_X1 u1_srl_151_U407 ( .A1(n8481), .A2(u1_srl_151_n20), .B1(n8484), .B2(
        u1_srl_151_n26), .ZN(u1_srl_151_n364) );
  AOI221_X1 u1_srl_151_U406 ( .B1(u1_srl_151_n6), .B2(n8483), .C1(
        u1_srl_151_n16), .C2(n8482), .A(u1_srl_151_n79), .ZN(u1_srl_151_n256)
         );
  AOI22_X1 u1_srl_151_U405 ( .A1(n6468), .A2(u1_srl_151_n20), .B1(n8480), .B2(
        u1_srl_151_n26), .ZN(u1_srl_151_n363) );
  AOI221_X1 u1_srl_151_U404 ( .B1(u1_srl_151_n6), .B2(n8478), .C1(
        u1_srl_151_n16), .C2(u1_adj_op_51_), .A(u1_srl_151_n81), .ZN(
        u1_srl_151_n193) );
  AOI22_X1 u1_srl_151_U403 ( .A1(u1_srl_151_n78), .A2(u1_srl_151_n31), .B1(
        u1_srl_151_n80), .B2(u1_srl_151_n13), .ZN(u1_srl_151_n201) );
  AOI22_X1 u1_srl_151_U402 ( .A1(n8474), .A2(u1_srl_151_n20), .B1(n8477), .B2(
        u1_srl_151_n26), .ZN(u1_srl_151_n362) );
  OAI221_X1 u1_srl_151_U401 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n116), .C1(
        u1_srl_151_n14), .C2(u1_srl_151_n115), .A(u1_srl_151_n362), .ZN(
        u1_srl_151_n169) );
  AOI22_X1 u1_srl_151_U400 ( .A1(n8505), .A2(u1_srl_151_n20), .B1(n8473), .B2(
        u1_srl_151_n26), .ZN(u1_srl_151_n361) );
  OAI221_X1 u1_srl_151_U399 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n149), .C1(
        u1_srl_151_n14), .C2(u1_srl_151_n148), .A(u1_srl_151_n361), .ZN(
        u1_srl_151_n166) );
  AOI22_X1 u1_srl_151_U398 ( .A1(u1_srl_151_n169), .A2(u1_srl_151_n157), .B1(
        u1_srl_151_n166), .B2(u1_srl_151_n155), .ZN(u1_srl_151_n359) );
  NAND3_X1 u1_srl_151_U397 ( .A1(u1_adj_op_0_), .A2(u1_srl_151_n17), .A3(
        u1_srl_151_n160), .ZN(u1_srl_151_n360) );
  OAI211_X1 u1_srl_151_U396 ( .C1(u1_srl_151_n238), .C2(u1_srl_151_n201), .A(
        u1_srl_151_n359), .B(u1_srl_151_n360), .ZN(u1_srl_151_n358) );
  NAND2_X1 u1_srl_151_U395 ( .A1(u1_srl_151_n357), .A2(u1_srl_151_n37), .ZN(
        u1_adj_op_out_sft_0_) );
  AOI22_X1 u1_srl_151_U394 ( .A1(n8493), .A2(u1_srl_151_n20), .B1(
        u1_adj_op_27_), .B2(u1_srl_151_n26), .ZN(u1_srl_151_n356) );
  OAI221_X1 u1_srl_151_U393 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n130), .C1(
        u1_srl_151_n14), .C2(u1_srl_151_n129), .A(u1_srl_151_n356), .ZN(
        u1_srl_151_n274) );
  AOI22_X1 u1_srl_151_U392 ( .A1(n8496), .A2(u1_srl_151_n20), .B1(n8499), .B2(
        u1_srl_151_n26), .ZN(u1_srl_151_n355) );
  OAI221_X1 u1_srl_151_U391 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n134), .C1(
        u1_srl_151_n14), .C2(u1_srl_151_n133), .A(u1_srl_151_n355), .ZN(
        u1_srl_151_n270) );
  AOI22_X1 u1_srl_151_U390 ( .A1(u1_adj_op_38_), .A2(u1_srl_151_n20), .B1(
        n8489), .B2(u1_srl_151_n26), .ZN(u1_srl_151_n354) );
  OAI221_X1 u1_srl_151_U389 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n121), .C1(
        u1_srl_151_n14), .C2(u1_srl_151_n120), .A(u1_srl_151_n354), .ZN(
        u1_srl_151_n275) );
  AOI22_X1 u1_srl_151_U388 ( .A1(n8490), .A2(u1_srl_151_n20), .B1(n8492), .B2(
        u1_srl_151_n26), .ZN(u1_srl_151_n353) );
  OAI221_X1 u1_srl_151_U387 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n125), .C1(
        u1_srl_151_n14), .C2(u1_srl_151_n124), .A(u1_srl_151_n353), .ZN(
        u1_srl_151_n273) );
  AOI22_X1 u1_srl_151_U386 ( .A1(u1_srl_151_n252), .A2(u1_srl_151_n275), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n273), .ZN(u1_srl_151_n352) );
  AOI221_X1 u1_srl_151_U385 ( .B1(u1_srl_151_n274), .B2(u1_srl_151_n13), .C1(
        u1_srl_151_n270), .C2(u1_srl_151_n31), .A(u1_srl_151_n62), .ZN(
        u1_srl_151_n246) );
  AOI22_X1 u1_srl_151_U384 ( .A1(n8483), .A2(u1_srl_151_n20), .B1(n8485), .B2(
        u1_srl_151_n25), .ZN(u1_srl_151_n351) );
  AOI221_X1 u1_srl_151_U383 ( .B1(u1_srl_151_n6), .B2(u1_adj_op_44_), .C1(
        u1_srl_151_n16), .C2(n8484), .A(u1_srl_151_n83), .ZN(u1_srl_151_n278)
         );
  AOI22_X1 u1_srl_151_U382 ( .A1(u1_adj_op_42_), .A2(u1_srl_151_n20), .B1(
        n8488), .B2(u1_srl_151_n25), .ZN(u1_srl_151_n350) );
  AOI221_X1 u1_srl_151_U381 ( .B1(u1_srl_151_n6), .B2(n8487), .C1(
        u1_srl_151_n16), .C2(n8486), .A(u1_srl_151_n85), .ZN(u1_srl_151_n301)
         );
  AOI22_X1 u1_srl_151_U380 ( .A1(u1_srl_151_n27), .A2(u1_adj_op_51_), .B1(
        u1_srl_151_n6), .B2(n6468), .ZN(u1_srl_151_n191) );
  AOI22_X1 u1_srl_151_U379 ( .A1(n8478), .A2(u1_srl_151_n19), .B1(n8482), .B2(
        u1_srl_151_n25), .ZN(u1_srl_151_n349) );
  AOI221_X1 u1_srl_151_U378 ( .B1(u1_srl_151_n6), .B2(n8481), .C1(
        u1_srl_151_n16), .C2(n8480), .A(u1_srl_151_n88), .ZN(u1_srl_151_n277)
         );
  OAI22_X1 u1_srl_151_U377 ( .A1(u1_srl_151_n72), .A2(u1_srl_151_n191), .B1(
        u1_srl_151_n4), .B2(u1_srl_151_n277), .ZN(u1_srl_151_n348) );
  AOI221_X1 u1_srl_151_U376 ( .B1(u1_srl_151_n82), .B2(u1_srl_151_n13), .C1(
        u1_srl_151_n84), .C2(u1_srl_151_n31), .A(u1_srl_151_n348), .ZN(
        u1_srl_151_n205) );
  AOI22_X1 u1_srl_151_U375 ( .A1(u1_adj_op_10_), .A2(u1_srl_151_n19), .B1(
        n8475), .B2(u1_srl_151_n25), .ZN(u1_srl_151_n347) );
  OAI221_X1 u1_srl_151_U374 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n114), .C1(
        u1_srl_151_n14), .C2(u1_srl_151_n113), .A(u1_srl_151_n347), .ZN(
        u1_srl_151_n181) );
  AOI22_X1 u1_srl_151_U373 ( .A1(u1_srl_151_n159), .A2(u1_srl_151_n42), .B1(
        u1_srl_151_n160), .B2(u1_srl_151_n181), .ZN(u1_srl_151_n342) );
  AOI22_X1 u1_srl_151_U372 ( .A1(n8503), .A2(u1_srl_151_n19), .B1(
        u1_adj_op_11_), .B2(u1_srl_151_n25), .ZN(u1_srl_151_n346) );
  OAI221_X1 u1_srl_151_U371 ( .B1(u1_srl_151_n7), .B2(u1_srl_151_n147), .C1(
        u1_srl_151_n14), .C2(u1_srl_151_n146), .A(u1_srl_151_n346), .ZN(
        u1_srl_151_n183) );
  AOI22_X1 u1_srl_151_U370 ( .A1(u1_adj_op_22_), .A2(u1_srl_151_n19), .B1(
        u1_srl_151_n27), .B2(n8501), .ZN(u1_srl_151_n345) );
  OAI221_X1 u1_srl_151_U369 ( .B1(u1_srl_151_n7), .B2(u1_srl_151_n138), .C1(
        u1_srl_151_n15), .C2(u1_srl_151_n137), .A(u1_srl_151_n345), .ZN(
        u1_srl_151_n271) );
  AOI22_X1 u1_srl_151_U368 ( .A1(n8502), .A2(u1_srl_151_n19), .B1(
        u1_adj_op_15_), .B2(u1_srl_151_n25), .ZN(u1_srl_151_n344) );
  OAI221_X1 u1_srl_151_U367 ( .B1(u1_srl_151_n7), .B2(u1_srl_151_n143), .C1(
        u1_srl_151_n15), .C2(u1_srl_151_n142), .A(u1_srl_151_n344), .ZN(
        u1_srl_151_n182) );
  AOI222_X1 u1_srl_151_U366 ( .A1(u1_srl_151_n153), .A2(u1_srl_151_n183), .B1(
        u1_srl_151_n155), .B2(u1_srl_151_n271), .C1(u1_srl_151_n157), .C2(
        u1_srl_151_n182), .ZN(u1_srl_151_n343) );
  OAI211_X1 u1_srl_151_U365 ( .C1(u1_srl_151_n246), .C2(u1_srl_151_n110), .A(
        u1_srl_151_n342), .B(u1_srl_151_n343), .ZN(u1_adj_op_out_sft_10_) );
  AOI22_X1 u1_srl_151_U364 ( .A1(n8492), .A2(u1_srl_151_n19), .B1(
        u1_adj_op_28_), .B2(u1_srl_151_n25), .ZN(u1_srl_151_n341) );
  OAI221_X1 u1_srl_151_U363 ( .B1(u1_srl_151_n7), .B2(u1_srl_151_n129), .C1(
        u1_srl_151_n15), .C2(u1_srl_151_n127), .A(u1_srl_151_n341), .ZN(
        u1_srl_151_n294) );
  AOI22_X1 u1_srl_151_U362 ( .A1(u1_adj_op_27_), .A2(u1_srl_151_n19), .B1(
        n8498), .B2(u1_srl_151_n25), .ZN(u1_srl_151_n340) );
  OAI221_X1 u1_srl_151_U361 ( .B1(u1_srl_151_n7), .B2(u1_srl_151_n133), .C1(
        u1_srl_151_n15), .C2(u1_srl_151_n132), .A(u1_srl_151_n340), .ZN(
        u1_srl_151_n263) );
  AOI22_X1 u1_srl_151_U360 ( .A1(n8488), .A2(u1_srl_151_n19), .B1(
        u1_adj_op_36_), .B2(u1_srl_151_n25), .ZN(u1_srl_151_n339) );
  AOI221_X1 u1_srl_151_U359 ( .B1(u1_srl_151_n6), .B2(u1_adj_op_37_), .C1(
        u1_srl_151_n16), .C2(u1_adj_op_38_), .A(u1_srl_151_n92), .ZN(
        u1_srl_151_n298) );
  AOI22_X1 u1_srl_151_U358 ( .A1(n8489), .A2(u1_srl_151_n19), .B1(
        u1_adj_op_32_), .B2(u1_srl_151_n25), .ZN(u1_srl_151_n338) );
  OAI221_X1 u1_srl_151_U357 ( .B1(u1_srl_151_n7), .B2(u1_srl_151_n124), .C1(
        u1_srl_151_n15), .C2(u1_srl_151_n123), .A(u1_srl_151_n338), .ZN(
        u1_srl_151_n296) );
  OAI22_X1 u1_srl_151_U356 ( .A1(u1_srl_151_n72), .A2(u1_srl_151_n298), .B1(
        u1_srl_151_n4), .B2(u1_srl_151_n93), .ZN(u1_srl_151_n337) );
  AOI221_X1 u1_srl_151_U355 ( .B1(u1_srl_151_n294), .B2(u1_srl_151_n13), .C1(
        u1_srl_151_n263), .C2(u1_srl_151_n31), .A(u1_srl_151_n337), .ZN(
        u1_srl_151_n244) );
  AOI22_X1 u1_srl_151_U354 ( .A1(n8485), .A2(u1_srl_151_n19), .B1(n8487), .B2(
        u1_srl_151_n25), .ZN(u1_srl_151_n336) );
  AOI221_X1 u1_srl_151_U353 ( .B1(u1_srl_151_n6), .B2(n8486), .C1(
        u1_srl_151_n16), .C2(u1_adj_op_42_), .A(u1_srl_151_n95), .ZN(
        u1_srl_151_n269) );
  AOI22_X1 u1_srl_151_U352 ( .A1(n8482), .A2(u1_srl_151_n19), .B1(
        u1_adj_op_44_), .B2(u1_srl_151_n24), .ZN(u1_srl_151_n335) );
  AOI221_X1 u1_srl_151_U351 ( .B1(u1_srl_151_n6), .B2(n8484), .C1(
        u1_srl_151_n16), .C2(n8483), .A(u1_srl_151_n96), .ZN(u1_srl_151_n268)
         );
  NAND2_X1 u1_srl_151_U350 ( .A1(n6468), .A2(u1_srl_151_n27), .ZN(
        u1_srl_151_n190) );
  AOI22_X1 u1_srl_151_U349 ( .A1(u1_adj_op_51_), .A2(u1_srl_151_n18), .B1(
        n8481), .B2(u1_srl_151_n24), .ZN(u1_srl_151_n334) );
  AOI221_X1 u1_srl_151_U348 ( .B1(u1_srl_151_n6), .B2(n8480), .C1(
        u1_srl_151_n16), .C2(n8478), .A(u1_srl_151_n97), .ZN(u1_srl_151_n267)
         );
  MUX2_X1 u1_srl_151_U347 ( .A(u1_srl_151_n190), .B(u1_srl_151_n267), .S(
        u1_srl_151_n73), .Z(u1_srl_151_n295) );
  OAI222_X1 u1_srl_151_U346 ( .A1(u1_srl_151_n269), .A2(u1_srl_151_n32), .B1(
        u1_srl_151_n268), .B2(u1_srl_151_n1), .C1(u1_srl_151_n295), .C2(
        u1_srl_151_n108), .ZN(u1_srl_151_n245) );
  AOI22_X1 u1_srl_151_U345 ( .A1(u1_adj_op_11_), .A2(u1_srl_151_n18), .B1(
        n8474), .B2(u1_srl_151_n24), .ZN(u1_srl_151_n333) );
  OAI221_X1 u1_srl_151_U344 ( .B1(u1_srl_151_n7), .B2(u1_srl_151_n113), .C1(
        u1_srl_151_n15), .C2(u1_srl_151_n149), .A(u1_srl_151_n333), .ZN(
        u1_srl_151_n173) );
  AOI22_X1 u1_srl_151_U343 ( .A1(u1_srl_151_n159), .A2(u1_srl_151_n245), .B1(
        u1_srl_151_n160), .B2(u1_srl_151_n173), .ZN(u1_srl_151_n328) );
  AOI22_X1 u1_srl_151_U342 ( .A1(u1_adj_op_15_), .A2(u1_srl_151_n18), .B1(
        n8505), .B2(u1_srl_151_n24), .ZN(u1_srl_151_n332) );
  OAI221_X1 u1_srl_151_U341 ( .B1(u1_srl_151_n7), .B2(u1_srl_151_n146), .C1(
        u1_srl_151_n15), .C2(u1_srl_151_n145), .A(u1_srl_151_n332), .ZN(
        u1_srl_151_n175) );
  AOI22_X1 u1_srl_151_U340 ( .A1(n8499), .A2(u1_srl_151_n18), .B1(
        u1_srl_151_n27), .B2(u1_adj_op_20_), .ZN(u1_srl_151_n331) );
  OAI221_X1 u1_srl_151_U339 ( .B1(u1_srl_151_n7), .B2(u1_srl_151_n137), .C1(
        u1_srl_151_n15), .C2(u1_srl_151_n136), .A(u1_srl_151_n331), .ZN(
        u1_srl_151_n264) );
  AOI22_X1 u1_srl_151_U338 ( .A1(u1_srl_151_n17), .A2(n8501), .B1(
        u1_adj_op_16_), .B2(u1_srl_151_n24), .ZN(u1_srl_151_n330) );
  OAI221_X1 u1_srl_151_U337 ( .B1(u1_srl_151_n7), .B2(u1_srl_151_n142), .C1(
        u1_srl_151_n15), .C2(u1_srl_151_n141), .A(u1_srl_151_n330), .ZN(
        u1_srl_151_n174) );
  AOI222_X1 u1_srl_151_U336 ( .A1(u1_srl_151_n153), .A2(u1_srl_151_n175), .B1(
        u1_srl_151_n155), .B2(u1_srl_151_n264), .C1(u1_srl_151_n157), .C2(
        u1_srl_151_n174), .ZN(u1_srl_151_n329) );
  OAI211_X1 u1_srl_151_U335 ( .C1(u1_srl_151_n244), .C2(u1_srl_151_n110), .A(
        u1_srl_151_n328), .B(u1_srl_151_n329), .ZN(u1_adj_op_out_sft_11_) );
  AOI22_X1 u1_srl_151_U334 ( .A1(u1_srl_151_n252), .A2(u1_srl_151_n76), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n260), .ZN(u1_srl_151_n326) );
  AOI221_X1 u1_srl_151_U333 ( .B1(u1_srl_151_n261), .B2(u1_srl_151_n13), .C1(
        u1_srl_151_n257), .C2(u1_srl_151_n31), .A(u1_srl_151_n63), .ZN(
        u1_srl_151_n243) );
  AOI222_X1 u1_srl_151_U332 ( .A1(u1_srl_151_n78), .A2(u1_srl_151_n12), .B1(
        u1_srl_151_n80), .B2(u1_srl_151_n5), .C1(u1_srl_151_n74), .C2(
        u1_srl_151_n29), .ZN(u1_srl_151_n204) );
  AOI22_X1 u1_srl_151_U331 ( .A1(u1_srl_151_n159), .A2(u1_srl_151_n43), .B1(
        u1_srl_151_n160), .B2(u1_srl_151_n166), .ZN(u1_srl_151_n324) );
  AOI222_X1 u1_srl_151_U330 ( .A1(u1_srl_151_n153), .A2(u1_srl_151_n168), .B1(
        u1_srl_151_n155), .B2(u1_srl_151_n258), .C1(u1_srl_151_n157), .C2(
        u1_srl_151_n167), .ZN(u1_srl_151_n325) );
  OAI211_X1 u1_srl_151_U329 ( .C1(u1_srl_151_n243), .C2(u1_srl_151_n110), .A(
        u1_srl_151_n324), .B(u1_srl_151_n325), .ZN(u1_adj_op_out_sft_12_) );
  AOI22_X1 u1_srl_151_U328 ( .A1(n8491), .A2(u1_srl_151_n18), .B1(n8493), .B2(
        u1_srl_151_n24), .ZN(u1_srl_151_n323) );
  OAI221_X1 u1_srl_151_U327 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n126), .C1(
        u1_srl_151_n15), .C2(u1_srl_151_n125), .A(u1_srl_151_n323), .ZN(
        u1_srl_151_n254) );
  AOI22_X1 u1_srl_151_U326 ( .A1(n8495), .A2(u1_srl_151_n18), .B1(n8496), .B2(
        u1_srl_151_n24), .ZN(u1_srl_151_n322) );
  OAI221_X1 u1_srl_151_U325 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n131), .C1(
        u1_srl_151_n14), .C2(u1_srl_151_n130), .A(u1_srl_151_n322), .ZN(
        u1_srl_151_n249) );
  AOI22_X1 u1_srl_151_U324 ( .A1(n8486), .A2(u1_srl_151_n18), .B1(
        u1_adj_op_38_), .B2(u1_srl_151_n24), .ZN(u1_srl_151_n321) );
  AOI221_X1 u1_srl_151_U323 ( .B1(u1_srl_151_n6), .B2(n8488), .C1(
        u1_srl_151_n16), .C2(n8487), .A(u1_srl_151_n100), .ZN(u1_srl_151_n282)
         );
  AOI22_X1 u1_srl_151_U322 ( .A1(u1_adj_op_37_), .A2(u1_srl_151_n18), .B1(
        n8490), .B2(u1_srl_151_n24), .ZN(u1_srl_151_n320) );
  OAI221_X1 u1_srl_151_U321 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n122), .C1(
        u1_srl_151_n14), .C2(u1_srl_151_n121), .A(u1_srl_151_n320), .ZN(
        u1_srl_151_n253) );
  OAI22_X1 u1_srl_151_U320 ( .A1(u1_srl_151_n72), .A2(u1_srl_151_n282), .B1(
        u1_srl_151_n4), .B2(u1_srl_151_n101), .ZN(u1_srl_151_n319) );
  AOI221_X1 u1_srl_151_U319 ( .B1(u1_srl_151_n254), .B2(u1_srl_151_n13), .C1(
        u1_srl_151_n249), .C2(u1_srl_151_n31), .A(u1_srl_151_n319), .ZN(
        u1_srl_151_n242) );
  AOI22_X1 u1_srl_151_U318 ( .A1(n8480), .A2(u1_srl_151_n18), .B1(n8483), .B2(
        u1_srl_151_n24), .ZN(u1_srl_151_n318) );
  AOI221_X1 u1_srl_151_U317 ( .B1(u1_srl_151_n6), .B2(n8482), .C1(
        u1_srl_151_n16), .C2(n8481), .A(u1_srl_151_n103), .ZN(u1_srl_151_n248)
         );
  AOI222_X1 u1_srl_151_U316 ( .A1(u1_srl_151_n16), .A2(n6468), .B1(
        u1_srl_151_n6), .B2(u1_adj_op_51_), .C1(u1_srl_151_n27), .C2(n8478), 
        .ZN(u1_srl_151_n192) );
  AOI22_X1 u1_srl_151_U315 ( .A1(n8484), .A2(u1_srl_151_n18), .B1(
        u1_adj_op_42_), .B2(u1_srl_151_n24), .ZN(u1_srl_151_n317) );
  AOI221_X1 u1_srl_151_U314 ( .B1(u1_srl_151_n6), .B2(n8485), .C1(
        u1_srl_151_n16), .C2(u1_adj_op_44_), .A(u1_srl_151_n106), .ZN(
        u1_srl_151_n281) );
  AOI222_X1 u1_srl_151_U313 ( .A1(u1_srl_151_n102), .A2(u1_srl_151_n12), .B1(
        u1_srl_151_n104), .B2(u1_srl_151_n5), .C1(u1_srl_151_n105), .C2(
        u1_srl_151_n29), .ZN(u1_srl_151_n203) );
  AOI22_X1 u1_srl_151_U312 ( .A1(n8504), .A2(u1_srl_151_n18), .B1(
        u1_adj_op_10_), .B2(u1_srl_151_n27), .ZN(u1_srl_151_n316) );
  OAI221_X1 u1_srl_151_U311 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n148), .C1(
        u1_srl_151_n14), .C2(u1_srl_151_n147), .A(u1_srl_151_n316), .ZN(
        u1_srl_151_n154) );
  AOI22_X1 u1_srl_151_U310 ( .A1(u1_srl_151_n159), .A2(u1_srl_151_n44), .B1(
        u1_srl_151_n160), .B2(u1_srl_151_n154), .ZN(u1_srl_151_n311) );
  AOI22_X1 u1_srl_151_U309 ( .A1(u1_adj_op_17_), .A2(u1_srl_151_n18), .B1(
        n8503), .B2(u1_srl_151_n27), .ZN(u1_srl_151_n315) );
  OAI221_X1 u1_srl_151_U308 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n144), .C1(
        u1_srl_151_n14), .C2(u1_srl_151_n143), .A(u1_srl_151_n315), .ZN(
        u1_srl_151_n158) );
  AOI22_X1 u1_srl_151_U307 ( .A1(n8497), .A2(u1_srl_151_n17), .B1(
        u1_adj_op_22_), .B2(u1_srl_151_n27), .ZN(u1_srl_151_n314) );
  OAI221_X1 u1_srl_151_U306 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n135), .C1(
        u1_srl_151_n14), .C2(u1_srl_151_n134), .A(u1_srl_151_n314), .ZN(
        u1_srl_151_n250) );
  AOI22_X1 u1_srl_151_U305 ( .A1(u1_adj_op_21_), .A2(u1_srl_151_n17), .B1(
        n8502), .B2(u1_srl_151_n24), .ZN(u1_srl_151_n313) );
  OAI221_X1 u1_srl_151_U304 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n140), .C1(
        u1_srl_151_n14), .C2(u1_srl_151_n138), .A(u1_srl_151_n313), .ZN(
        u1_srl_151_n156) );
  AOI222_X1 u1_srl_151_U303 ( .A1(u1_srl_151_n153), .A2(u1_srl_151_n158), .B1(
        u1_srl_151_n155), .B2(u1_srl_151_n250), .C1(u1_srl_151_n157), .C2(
        u1_srl_151_n156), .ZN(u1_srl_151_n312) );
  OAI211_X1 u1_srl_151_U302 ( .C1(u1_srl_151_n242), .C2(u1_srl_151_n110), .A(
        u1_srl_151_n311), .B(u1_srl_151_n312), .ZN(u1_adj_op_out_sft_13_) );
  AOI22_X1 u1_srl_151_U301 ( .A1(u1_srl_151_n252), .A2(u1_srl_151_n84), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n275), .ZN(u1_srl_151_n310) );
  AOI221_X1 u1_srl_151_U300 ( .B1(u1_srl_151_n273), .B2(u1_srl_151_n13), .C1(
        u1_srl_151_n274), .C2(u1_srl_151_n30), .A(u1_srl_151_n64), .ZN(
        u1_srl_151_n233) );
  AOI222_X1 u1_srl_151_U299 ( .A1(u1_srl_151_n87), .A2(u1_srl_151_n12), .B1(
        u1_srl_151_n86), .B2(u1_srl_151_n5), .C1(u1_srl_151_n82), .C2(
        u1_srl_151_n29), .ZN(u1_srl_151_n202) );
  AOI22_X1 u1_srl_151_U298 ( .A1(u1_srl_151_n159), .A2(u1_srl_151_n45), .B1(
        u1_srl_151_n160), .B2(u1_srl_151_n183), .ZN(u1_srl_151_n308) );
  AOI222_X1 u1_srl_151_U297 ( .A1(u1_srl_151_n153), .A2(u1_srl_151_n182), .B1(
        u1_srl_151_n155), .B2(u1_srl_151_n270), .C1(u1_srl_151_n157), .C2(
        u1_srl_151_n271), .ZN(u1_srl_151_n309) );
  OAI211_X1 u1_srl_151_U296 ( .C1(u1_srl_151_n233), .C2(u1_srl_151_n110), .A(
        u1_srl_151_n308), .B(u1_srl_151_n309), .ZN(u1_adj_op_out_sft_14_) );
  OAI22_X1 u1_srl_151_U295 ( .A1(u1_srl_151_n72), .A2(u1_srl_151_n269), .B1(
        u1_srl_151_n4), .B2(u1_srl_151_n298), .ZN(u1_srl_151_n307) );
  AOI221_X1 u1_srl_151_U294 ( .B1(u1_srl_151_n296), .B2(u1_srl_151_n13), .C1(
        u1_srl_151_n294), .C2(u1_srl_151_n31), .A(u1_srl_151_n307), .ZN(
        u1_srl_151_n231) );
  OAI222_X1 u1_srl_151_U293 ( .A1(u1_srl_151_n267), .A2(u1_srl_151_n1), .B1(
        u1_srl_151_n4), .B2(u1_srl_151_n190), .C1(u1_srl_151_n268), .C2(
        u1_srl_151_n33), .ZN(u1_srl_151_n232) );
  AOI22_X1 u1_srl_151_U292 ( .A1(u1_srl_151_n159), .A2(u1_srl_151_n232), .B1(
        u1_srl_151_n160), .B2(u1_srl_151_n175), .ZN(u1_srl_151_n305) );
  AOI222_X1 u1_srl_151_U291 ( .A1(u1_srl_151_n153), .A2(u1_srl_151_n174), .B1(
        u1_srl_151_n155), .B2(u1_srl_151_n263), .C1(u1_srl_151_n157), .C2(
        u1_srl_151_n264), .ZN(u1_srl_151_n306) );
  OAI211_X1 u1_srl_151_U290 ( .C1(u1_srl_151_n231), .C2(u1_srl_151_n110), .A(
        u1_srl_151_n305), .B(u1_srl_151_n306), .ZN(u1_adj_op_out_sft_15_) );
  OAI222_X1 u1_srl_151_U289 ( .A1(u1_srl_151_n230), .A2(u1_srl_151_n110), .B1(
        u1_srl_151_n201), .B2(u1_srl_151_n109), .C1(u1_srl_151_n304), .C2(
        u1_srl_151_n11), .ZN(u1_adj_op_out_sft_16_) );
  OAI22_X1 u1_srl_151_U288 ( .A1(u1_srl_151_n72), .A2(u1_srl_151_n281), .B1(
        u1_srl_151_n4), .B2(u1_srl_151_n282), .ZN(u1_srl_151_n303) );
  AOI221_X1 u1_srl_151_U287 ( .B1(u1_srl_151_n253), .B2(u1_srl_151_n13), .C1(
        u1_srl_151_n254), .C2(u1_srl_151_n30), .A(u1_srl_151_n303), .ZN(
        u1_srl_151_n229) );
  AOI22_X1 u1_srl_151_U286 ( .A1(u1_srl_151_n102), .A2(u1_srl_151_n31), .B1(
        u1_srl_151_n104), .B2(u1_srl_151_n13), .ZN(u1_srl_151_n200) );
  AOI22_X1 u1_srl_151_U285 ( .A1(u1_srl_151_n252), .A2(u1_srl_151_n249), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n250), .ZN(u1_srl_151_n302) );
  AOI221_X1 u1_srl_151_U284 ( .B1(u1_srl_151_n156), .B2(u1_srl_151_n13), .C1(
        u1_srl_151_n158), .C2(u1_srl_151_n30), .A(u1_srl_151_n65), .ZN(
        u1_srl_151_n292) );
  OAI222_X1 u1_srl_151_U283 ( .A1(u1_srl_151_n229), .A2(u1_srl_151_n110), .B1(
        u1_srl_151_n200), .B2(u1_srl_151_n109), .C1(u1_srl_151_n292), .C2(
        u1_srl_151_n11), .ZN(u1_adj_op_out_sft_17_) );
  OAI22_X1 u1_srl_151_U282 ( .A1(u1_srl_151_n72), .A2(u1_srl_151_n278), .B1(
        u1_srl_151_n4), .B2(u1_srl_151_n301), .ZN(u1_srl_151_n300) );
  AOI221_X1 u1_srl_151_U281 ( .B1(u1_srl_151_n275), .B2(u1_srl_151_n13), .C1(
        u1_srl_151_n273), .C2(u1_srl_151_n30), .A(u1_srl_151_n300), .ZN(
        u1_srl_151_n228) );
  AOI22_X1 u1_srl_151_U280 ( .A1(u1_srl_151_n87), .A2(u1_srl_151_n31), .B1(
        u1_srl_151_n86), .B2(u1_srl_151_n13), .ZN(u1_srl_151_n195) );
  AOI22_X1 u1_srl_151_U279 ( .A1(u1_srl_151_n252), .A2(u1_srl_151_n274), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n270), .ZN(u1_srl_151_n299) );
  AOI221_X1 u1_srl_151_U278 ( .B1(u1_srl_151_n271), .B2(u1_srl_151_n13), .C1(
        u1_srl_151_n182), .C2(u1_srl_151_n30), .A(u1_srl_151_n66), .ZN(
        u1_srl_151_n241) );
  OAI222_X1 u1_srl_151_U277 ( .A1(u1_srl_151_n228), .A2(u1_srl_151_n110), .B1(
        u1_srl_151_n195), .B2(u1_srl_151_n109), .C1(u1_srl_151_n241), .C2(
        u1_srl_151_n11), .ZN(u1_adj_op_out_sft_18_) );
  OAI22_X1 u1_srl_151_U276 ( .A1(u1_srl_151_n72), .A2(u1_srl_151_n268), .B1(
        u1_srl_151_n4), .B2(u1_srl_151_n269), .ZN(u1_srl_151_n297) );
  AOI221_X1 u1_srl_151_U275 ( .B1(u1_srl_151_n91), .B2(u1_srl_151_n13), .C1(
        u1_srl_151_n296), .C2(u1_srl_151_n30), .A(u1_srl_151_n297), .ZN(
        u1_srl_151_n227) );
  OR2_X1 u1_srl_151_U274 ( .A1(u1_srl_151_n295), .A2(n8468), .ZN(
        u1_srl_151_n194) );
  OAI22_X1 u1_srl_151_U273 ( .A1(u1_srl_151_n72), .A2(u1_srl_151_n89), .B1(
        u1_srl_151_n4), .B2(u1_srl_151_n90), .ZN(u1_srl_151_n293) );
  AOI221_X1 u1_srl_151_U272 ( .B1(u1_srl_151_n264), .B2(u1_srl_151_n13), .C1(
        u1_srl_151_n174), .C2(u1_srl_151_n30), .A(u1_srl_151_n293), .ZN(
        u1_srl_151_n215) );
  OAI222_X1 u1_srl_151_U271 ( .A1(u1_srl_151_n227), .A2(u1_srl_151_n110), .B1(
        u1_srl_151_n109), .B2(u1_srl_151_n194), .C1(u1_srl_151_n215), .C2(
        u1_srl_151_n11), .ZN(u1_adj_op_out_sft_19_) );
  AOI22_X1 u1_srl_151_U270 ( .A1(n8477), .A2(u1_srl_151_n17), .B1(n8494), .B2(
        u1_srl_151_n27), .ZN(u1_srl_151_n291) );
  OAI221_X1 u1_srl_151_U269 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n119), .C1(
        u1_srl_151_n14), .C2(u1_srl_151_n118), .A(u1_srl_151_n291), .ZN(
        u1_srl_151_n188) );
  AOI222_X1 u1_srl_151_U268 ( .A1(u1_srl_151_n177), .A2(u1_srl_151_n47), .B1(
        u1_srl_151_n153), .B2(u1_srl_151_n188), .C1(u1_srl_151_n159), .C2(
        u1_srl_151_n46), .ZN(u1_srl_151_n286) );
  AOI22_X1 u1_srl_151_U267 ( .A1(u1_srl_151_n17), .A2(n8500), .B1(
        u1_srl_151_n16), .B2(u1_adj_op_0_), .ZN(u1_srl_151_n288) );
  AOI22_X1 u1_srl_151_U266 ( .A1(n8473), .A2(u1_srl_151_n17), .B1(n8476), .B2(
        u1_srl_151_n27), .ZN(u1_srl_151_n290) );
  OAI221_X1 u1_srl_151_U265 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n115), .C1(
        u1_srl_151_n14), .C2(u1_srl_151_n114), .A(u1_srl_151_n290), .ZN(
        u1_srl_151_n161) );
  AOI22_X1 u1_srl_151_U264 ( .A1(u1_srl_151_n161), .A2(u1_srl_151_n157), .B1(
        u1_srl_151_n154), .B2(u1_srl_151_n155), .ZN(u1_srl_151_n289) );
  OAI221_X1 u1_srl_151_U263 ( .B1(u1_srl_151_n39), .B2(u1_srl_151_n288), .C1(
        u1_srl_151_n238), .C2(u1_srl_151_n200), .A(u1_srl_151_n289), .ZN(
        u1_srl_151_n287) );
  NAND2_X1 u1_srl_151_U262 ( .A1(u1_srl_151_n286), .A2(u1_srl_151_n38), .ZN(
        u1_adj_op_out_sft_1_) );
  OAI22_X1 u1_srl_151_U261 ( .A1(u1_srl_151_n72), .A2(u1_srl_151_n256), .B1(
        u1_srl_151_n4), .B2(u1_srl_151_n285), .ZN(u1_srl_151_n284) );
  AOI221_X1 u1_srl_151_U260 ( .B1(u1_srl_151_n76), .B2(u1_srl_151_n13), .C1(
        u1_srl_151_n260), .C2(u1_srl_151_n30), .A(u1_srl_151_n284), .ZN(
        u1_srl_151_n225) );
  NAND2_X1 u1_srl_151_U259 ( .A1(u1_srl_151_n159), .A2(u1_srl_151_n30), .ZN(
        u1_srl_151_n262) );
  AOI22_X1 u1_srl_151_U258 ( .A1(u1_srl_151_n252), .A2(u1_srl_151_n261), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n257), .ZN(u1_srl_151_n283) );
  AOI221_X1 u1_srl_151_U257 ( .B1(u1_srl_151_n258), .B2(u1_srl_151_n13), .C1(
        u1_srl_151_n167), .C2(u1_srl_151_n30), .A(u1_srl_151_n67), .ZN(
        u1_srl_151_n199) );
  OAI222_X1 u1_srl_151_U256 ( .A1(u1_srl_151_n225), .A2(u1_srl_151_n110), .B1(
        u1_srl_151_n193), .B2(u1_srl_151_n262), .C1(u1_srl_151_n199), .C2(
        u1_srl_151_n11), .ZN(u1_adj_op_out_sft_20_) );
  OAI22_X1 u1_srl_151_U255 ( .A1(u1_srl_151_n72), .A2(u1_srl_151_n248), .B1(
        u1_srl_151_n4), .B2(u1_srl_151_n281), .ZN(u1_srl_151_n280) );
  AOI221_X1 u1_srl_151_U254 ( .B1(u1_srl_151_n99), .B2(u1_srl_151_n13), .C1(
        u1_srl_151_n253), .C2(u1_srl_151_n30), .A(u1_srl_151_n280), .ZN(
        u1_srl_151_n223) );
  AOI22_X1 u1_srl_151_U253 ( .A1(u1_srl_151_n252), .A2(u1_srl_151_n254), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n249), .ZN(u1_srl_151_n279) );
  AOI221_X1 u1_srl_151_U252 ( .B1(u1_srl_151_n250), .B2(u1_srl_151_n12), .C1(
        u1_srl_151_n156), .C2(u1_srl_151_n29), .A(u1_srl_151_n68), .ZN(
        u1_srl_151_n189) );
  OAI222_X1 u1_srl_151_U251 ( .A1(u1_srl_151_n223), .A2(u1_srl_151_n110), .B1(
        u1_srl_151_n192), .B2(u1_srl_151_n262), .C1(u1_srl_151_n189), .C2(
        u1_srl_151_n11), .ZN(u1_adj_op_out_sft_21_) );
  OAI22_X1 u1_srl_151_U250 ( .A1(u1_srl_151_n72), .A2(u1_srl_151_n277), .B1(
        u1_srl_151_n4), .B2(u1_srl_151_n278), .ZN(u1_srl_151_n276) );
  AOI221_X1 u1_srl_151_U249 ( .B1(u1_srl_151_n84), .B2(u1_srl_151_n13), .C1(
        u1_srl_151_n275), .C2(u1_srl_151_n30), .A(u1_srl_151_n276), .ZN(
        u1_srl_151_n221) );
  AOI22_X1 u1_srl_151_U248 ( .A1(u1_srl_151_n252), .A2(u1_srl_151_n273), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n274), .ZN(u1_srl_151_n272) );
  AOI221_X1 u1_srl_151_U247 ( .B1(u1_srl_151_n270), .B2(u1_srl_151_n12), .C1(
        u1_srl_151_n271), .C2(u1_srl_151_n29), .A(u1_srl_151_n69), .ZN(
        u1_srl_151_n185) );
  OAI222_X1 u1_srl_151_U246 ( .A1(u1_srl_151_n221), .A2(u1_srl_151_n110), .B1(
        u1_srl_151_n191), .B2(u1_srl_151_n262), .C1(u1_srl_151_n185), .C2(
        u1_srl_151_n11), .ZN(u1_adj_op_out_sft_22_) );
  OAI22_X1 u1_srl_151_U245 ( .A1(u1_srl_151_n72), .A2(u1_srl_151_n267), .B1(
        u1_srl_151_n4), .B2(u1_srl_151_n268), .ZN(u1_srl_151_n266) );
  AOI221_X1 u1_srl_151_U244 ( .B1(u1_srl_151_n94), .B2(u1_srl_151_n12), .C1(
        u1_srl_151_n91), .C2(u1_srl_151_n29), .A(u1_srl_151_n266), .ZN(
        u1_srl_151_n218) );
  OAI22_X1 u1_srl_151_U243 ( .A1(u1_srl_151_n72), .A2(u1_srl_151_n93), .B1(
        u1_srl_151_n4), .B2(u1_srl_151_n89), .ZN(u1_srl_151_n265) );
  AOI221_X1 u1_srl_151_U242 ( .B1(u1_srl_151_n263), .B2(u1_srl_151_n12), .C1(
        u1_srl_151_n264), .C2(u1_srl_151_n29), .A(u1_srl_151_n265), .ZN(
        u1_srl_151_n178) );
  OAI222_X1 u1_srl_151_U241 ( .A1(u1_srl_151_n218), .A2(u1_srl_151_n110), .B1(
        u1_srl_151_n190), .B2(u1_srl_151_n262), .C1(u1_srl_151_n178), .C2(
        u1_srl_151_n11), .ZN(u1_adj_op_out_sft_23_) );
  AOI22_X1 u1_srl_151_U240 ( .A1(u1_srl_151_n252), .A2(u1_srl_151_n260), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n261), .ZN(u1_srl_151_n259) );
  AOI221_X1 u1_srl_151_U239 ( .B1(u1_srl_151_n257), .B2(u1_srl_151_n12), .C1(
        u1_srl_151_n258), .C2(u1_srl_151_n29), .A(u1_srl_151_n70), .ZN(
        u1_srl_151_n163) );
  OAI22_X1 u1_srl_151_U238 ( .A1(u1_srl_151_n72), .A2(u1_srl_151_n193), .B1(
        u1_srl_151_n4), .B2(u1_srl_151_n256), .ZN(u1_srl_151_n255) );
  AOI221_X1 u1_srl_151_U237 ( .B1(u1_srl_151_n74), .B2(u1_srl_151_n12), .C1(
        u1_srl_151_n76), .C2(u1_srl_151_n29), .A(u1_srl_151_n255), .ZN(
        u1_srl_151_n170) );
  OAI22_X1 u1_srl_151_U236 ( .A1(u1_srl_151_n163), .A2(u1_srl_151_n10), .B1(
        u1_srl_151_n170), .B2(u1_srl_151_n110), .ZN(u1_adj_op_out_sft_24_) );
  AOI22_X1 u1_srl_151_U235 ( .A1(u1_srl_151_n252), .A2(u1_srl_151_n253), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n254), .ZN(u1_srl_151_n251) );
  AOI221_X1 u1_srl_151_U234 ( .B1(u1_srl_151_n249), .B2(u1_srl_151_n12), .C1(
        u1_srl_151_n250), .C2(u1_srl_151_n29), .A(u1_srl_151_n71), .ZN(
        u1_srl_151_n150) );
  OAI22_X1 u1_srl_151_U233 ( .A1(u1_srl_151_n72), .A2(u1_srl_151_n192), .B1(
        u1_srl_151_n4), .B2(u1_srl_151_n248), .ZN(u1_srl_151_n247) );
  AOI221_X1 u1_srl_151_U232 ( .B1(u1_srl_151_n105), .B2(u1_srl_151_n12), .C1(
        u1_srl_151_n99), .C2(u1_srl_151_n29), .A(u1_srl_151_n247), .ZN(
        u1_srl_151_n162) );
  OAI22_X1 u1_srl_151_U231 ( .A1(u1_srl_151_n150), .A2(u1_srl_151_n10), .B1(
        u1_srl_151_n162), .B2(u1_srl_151_n110), .ZN(u1_adj_op_out_sft_25_) );
  OAI22_X1 u1_srl_151_U230 ( .A1(u1_srl_151_n246), .A2(u1_srl_151_n10), .B1(
        u1_srl_151_n205), .B2(u1_srl_151_n110), .ZN(u1_adj_op_out_sft_26_) );
  OAI22_X1 u1_srl_151_U229 ( .A1(u1_srl_151_n244), .A2(u1_srl_151_n10), .B1(
        u1_srl_151_n40), .B2(u1_srl_151_n110), .ZN(u1_adj_op_out_sft_27_) );
  OAI22_X1 u1_srl_151_U228 ( .A1(u1_srl_151_n243), .A2(u1_srl_151_n10), .B1(
        u1_srl_151_n204), .B2(u1_srl_151_n110), .ZN(u1_adj_op_out_sft_28_) );
  OAI22_X1 u1_srl_151_U227 ( .A1(u1_srl_151_n242), .A2(u1_srl_151_n10), .B1(
        u1_srl_151_n203), .B2(u1_srl_151_n110), .ZN(u1_adj_op_out_sft_29_) );
  AOI22_X1 u1_srl_151_U226 ( .A1(n8476), .A2(u1_srl_151_n17), .B1(u1_adj_op_3_), .B2(u1_srl_151_n27), .ZN(u1_srl_151_n240) );
  OAI221_X1 u1_srl_151_U225 ( .B1(u1_srl_151_n8), .B2(u1_srl_151_n118), .C1(
        u1_srl_151_n14), .C2(u1_srl_151_n117), .A(u1_srl_151_n240), .ZN(
        u1_srl_151_n184) );
  AOI222_X1 u1_srl_151_U224 ( .A1(u1_srl_151_n177), .A2(u1_srl_151_n49), .B1(
        u1_srl_151_n153), .B2(u1_srl_151_n184), .C1(u1_srl_151_n159), .C2(
        u1_srl_151_n48), .ZN(u1_srl_151_n234) );
  AOI222_X1 u1_srl_151_U223 ( .A1(n8494), .A2(u1_srl_151_n17), .B1(
        u1_adj_op_0_), .B2(u1_srl_151_n6), .C1(n8500), .C2(u1_srl_151_n16), 
        .ZN(u1_srl_151_n237) );
  OAI22_X1 u1_srl_151_U222 ( .A1(u1_srl_151_n237), .A2(u1_srl_151_n39), .B1(
        u1_srl_151_n195), .B2(u1_srl_151_n238), .ZN(u1_srl_151_n236) );
  AOI221_X1 u1_srl_151_U221 ( .B1(u1_srl_151_n155), .B2(u1_srl_151_n183), .C1(
        u1_srl_151_n157), .C2(u1_srl_151_n181), .A(u1_srl_151_n236), .ZN(
        u1_srl_151_n235) );
  NAND2_X1 u1_srl_151_U220 ( .A1(u1_srl_151_n234), .A2(u1_srl_151_n235), .ZN(
        u1_adj_op_out_sft_2_) );
  OAI22_X1 u1_srl_151_U219 ( .A1(u1_srl_151_n233), .A2(u1_srl_151_n10), .B1(
        u1_srl_151_n202), .B2(u1_srl_151_n110), .ZN(u1_adj_op_out_sft_30_) );
  OAI22_X1 u1_srl_151_U218 ( .A1(u1_srl_151_n231), .A2(u1_srl_151_n11), .B1(
        u1_srl_151_n41), .B2(u1_srl_151_n110), .ZN(u1_adj_op_out_sft_31_) );
  OAI22_X1 u1_srl_151_U217 ( .A1(u1_srl_151_n230), .A2(u1_srl_151_n10), .B1(
        u1_srl_151_n201), .B2(u1_srl_151_n110), .ZN(u1_adj_op_out_sft_32_) );
  OAI22_X1 u1_srl_151_U216 ( .A1(u1_srl_151_n229), .A2(u1_srl_151_n11), .B1(
        u1_srl_151_n200), .B2(u1_srl_151_n110), .ZN(u1_adj_op_out_sft_33_) );
  OAI22_X1 u1_srl_151_U215 ( .A1(u1_srl_151_n228), .A2(u1_srl_151_n11), .B1(
        u1_srl_151_n195), .B2(u1_srl_151_n110), .ZN(u1_adj_op_out_sft_34_) );
  MUX2_X1 u1_srl_151_U214 ( .A(u1_srl_151_n194), .B(u1_srl_151_n227), .S(
        u1_srl_151_n111), .Z(u1_srl_151_n216) );
  NOR2_X1 u1_srl_151_U213 ( .A1(n8470), .A2(u1_srl_151_n216), .ZN(
        u1_adj_op_out_sft_35_) );
  NAND2_X1 u1_srl_151_U212 ( .A1(n8469), .A2(u1_srl_151_n31), .ZN(
        u1_srl_151_n219) );
  OAI22_X1 u1_srl_151_U211 ( .A1(n8469), .A2(u1_srl_151_n225), .B1(
        u1_srl_151_n193), .B2(u1_srl_151_n219), .ZN(u1_srl_151_n224) );
  NOR2_X1 u1_srl_151_U210 ( .A1(n8470), .A2(u1_srl_151_n52), .ZN(
        u1_adj_op_out_sft_36_) );
  OAI22_X1 u1_srl_151_U209 ( .A1(n8469), .A2(u1_srl_151_n223), .B1(
        u1_srl_151_n192), .B2(u1_srl_151_n219), .ZN(u1_srl_151_n222) );
  NOR2_X1 u1_srl_151_U208 ( .A1(n8470), .A2(u1_srl_151_n54), .ZN(
        u1_adj_op_out_sft_37_) );
  OAI22_X1 u1_srl_151_U207 ( .A1(n8469), .A2(u1_srl_151_n221), .B1(
        u1_srl_151_n191), .B2(u1_srl_151_n219), .ZN(u1_srl_151_n220) );
  NOR2_X1 u1_srl_151_U206 ( .A1(n8470), .A2(u1_srl_151_n56), .ZN(
        u1_adj_op_out_sft_38_) );
  OAI22_X1 u1_srl_151_U205 ( .A1(n8469), .A2(u1_srl_151_n218), .B1(
        u1_srl_151_n219), .B2(u1_srl_151_n190), .ZN(u1_srl_151_n217) );
  NOR2_X1 u1_srl_151_U204 ( .A1(n8470), .A2(u1_srl_151_n58), .ZN(
        u1_adj_op_out_sft_39_) );
  OAI22_X1 u1_srl_151_U203 ( .A1(u1_srl_151_n14), .A2(u1_srl_151_n128), .B1(
        u1_srl_151_n8), .B2(u1_srl_151_n139), .ZN(u1_srl_151_n214) );
  AOI221_X1 u1_srl_151_U202 ( .B1(u1_adj_op_3_), .B2(u1_srl_151_n17), .C1(
        u1_adj_op_0_), .C2(u1_srl_151_n27), .A(u1_srl_151_n214), .ZN(
        u1_srl_151_n208) );
  AOI22_X1 u1_srl_151_U201 ( .A1(n8475), .A2(u1_srl_151_n19), .B1(n8479), .B2(
        u1_srl_151_n25), .ZN(u1_srl_151_n212) );
  OAI221_X1 u1_srl_151_U200 ( .B1(u1_srl_151_n7), .B2(u1_srl_151_n117), .C1(
        u1_srl_151_n15), .C2(u1_srl_151_n116), .A(u1_srl_151_n212), .ZN(
        u1_srl_151_n176) );
  AOI22_X1 u1_srl_151_U199 ( .A1(u1_srl_151_n5), .A2(u1_srl_151_n173), .B1(
        u1_srl_151_n13), .B2(u1_srl_151_n176), .ZN(u1_srl_151_n209) );
  OAI221_X1 u1_srl_151_U198 ( .B1(u1_srl_151_n208), .B2(u1_srl_151_n32), .C1(
        u1_srl_151_n98), .C2(u1_srl_151_n72), .A(u1_srl_151_n209), .ZN(
        u1_srl_151_n207) );
  MUX2_X1 u1_srl_151_U197 ( .A(u1_srl_151_n51), .B(u1_srl_151_n207), .S(
        u1_srl_151_n111), .Z(u1_srl_151_n206) );
  MUX2_X1 u1_srl_151_U196 ( .A(u1_srl_151_n50), .B(u1_srl_151_n206), .S(
        u1_srl_151_n112), .Z(u1_adj_op_out_sft_3_) );
  NOR2_X1 u1_srl_151_U195 ( .A1(u1_srl_151_n170), .A2(u1_srl_151_n11), .ZN(
        u1_adj_op_out_sft_40_) );
  NOR2_X1 u1_srl_151_U194 ( .A1(u1_srl_151_n162), .A2(u1_srl_151_n11), .ZN(
        u1_adj_op_out_sft_41_) );
  NOR2_X1 u1_srl_151_U193 ( .A1(u1_srl_151_n205), .A2(u1_srl_151_n11), .ZN(
        u1_adj_op_out_sft_42_) );
  NOR2_X1 u1_srl_151_U192 ( .A1(u1_srl_151_n40), .A2(u1_srl_151_n11), .ZN(
        u1_adj_op_out_sft_43_) );
  NOR2_X1 u1_srl_151_U191 ( .A1(u1_srl_151_n204), .A2(u1_srl_151_n11), .ZN(
        u1_adj_op_out_sft_44_) );
  NOR2_X1 u1_srl_151_U190 ( .A1(u1_srl_151_n203), .A2(u1_srl_151_n11), .ZN(
        u1_adj_op_out_sft_45_) );
  NOR2_X1 u1_srl_151_U189 ( .A1(u1_srl_151_n202), .A2(u1_srl_151_n11), .ZN(
        u1_adj_op_out_sft_46_) );
  NOR2_X1 u1_srl_151_U188 ( .A1(u1_srl_151_n41), .A2(u1_srl_151_n11), .ZN(
        u1_adj_op_out_sft_47_) );
  NOR2_X1 u1_srl_151_U187 ( .A1(u1_srl_151_n201), .A2(u1_srl_151_n11), .ZN(
        u1_adj_op_out_sft_48_) );
  NOR2_X1 u1_srl_151_U186 ( .A1(u1_srl_151_n200), .A2(u1_srl_151_n11), .ZN(
        u1_adj_op_out_sft_49_) );
  AOI22_X1 u1_srl_151_U185 ( .A1(u1_srl_151_n160), .A2(u1_srl_151_n198), .B1(
        u1_srl_151_n177), .B2(u1_srl_151_n53), .ZN(u1_srl_151_n196) );
  AOI222_X1 u1_srl_151_U184 ( .A1(u1_srl_151_n153), .A2(u1_srl_151_n169), .B1(
        u1_srl_151_n155), .B2(u1_srl_151_n168), .C1(u1_srl_151_n157), .C2(
        u1_srl_151_n166), .ZN(u1_srl_151_n197) );
  OAI211_X1 u1_srl_151_U183 ( .C1(u1_srl_151_n52), .C2(u1_srl_151_n112), .A(
        u1_srl_151_n196), .B(u1_srl_151_n197), .ZN(u1_adj_op_out_sft_4_) );
  NOR2_X1 u1_srl_151_U182 ( .A1(u1_srl_151_n195), .A2(u1_srl_151_n11), .ZN(
        u1_adj_op_out_sft_50_) );
  NOR2_X1 u1_srl_151_U181 ( .A1(u1_srl_151_n10), .A2(u1_srl_151_n194), .ZN(
        u1_adj_op_out_sft_51_) );
  NOR2_X1 u1_srl_151_U180 ( .A1(u1_srl_151_n193), .A2(u1_srl_151_n39), .ZN(
        u1_adj_op_out_sft_52_) );
  NOR2_X1 u1_srl_151_U179 ( .A1(u1_srl_151_n192), .A2(u1_srl_151_n39), .ZN(
        u1_adj_op_out_sft_53_) );
  NOR2_X1 u1_srl_151_U178 ( .A1(u1_srl_151_n191), .A2(u1_srl_151_n39), .ZN(
        u1_adj_op_out_sft_54_) );
  NOR2_X1 u1_srl_151_U177 ( .A1(u1_srl_151_n39), .A2(u1_srl_151_n190), .ZN(
        u1_adj_op_out_sft_55_) );
  AOI22_X1 u1_srl_151_U176 ( .A1(u1_srl_151_n160), .A2(u1_srl_151_n188), .B1(
        u1_srl_151_n177), .B2(u1_srl_151_n55), .ZN(u1_srl_151_n186) );
  AOI222_X1 u1_srl_151_U175 ( .A1(u1_srl_151_n153), .A2(u1_srl_151_n161), .B1(
        u1_srl_151_n155), .B2(u1_srl_151_n158), .C1(u1_srl_151_n157), .C2(
        u1_srl_151_n154), .ZN(u1_srl_151_n187) );
  OAI211_X1 u1_srl_151_U174 ( .C1(u1_srl_151_n54), .C2(u1_srl_151_n112), .A(
        u1_srl_151_n186), .B(u1_srl_151_n187), .ZN(u1_adj_op_out_sft_5_) );
  AOI22_X1 u1_srl_151_U173 ( .A1(u1_srl_151_n160), .A2(u1_srl_151_n184), .B1(
        u1_srl_151_n177), .B2(u1_srl_151_n57), .ZN(u1_srl_151_n179) );
  AOI222_X1 u1_srl_151_U172 ( .A1(u1_srl_151_n153), .A2(u1_srl_151_n181), .B1(
        u1_srl_151_n155), .B2(u1_srl_151_n182), .C1(u1_srl_151_n157), .C2(
        u1_srl_151_n183), .ZN(u1_srl_151_n180) );
  OAI211_X1 u1_srl_151_U171 ( .C1(u1_srl_151_n56), .C2(u1_srl_151_n112), .A(
        u1_srl_151_n179), .B(u1_srl_151_n180), .ZN(u1_adj_op_out_sft_6_) );
  AOI22_X1 u1_srl_151_U170 ( .A1(u1_srl_151_n160), .A2(u1_srl_151_n176), .B1(
        u1_srl_151_n177), .B2(u1_srl_151_n59), .ZN(u1_srl_151_n171) );
  AOI222_X1 u1_srl_151_U169 ( .A1(u1_srl_151_n153), .A2(u1_srl_151_n173), .B1(
        u1_srl_151_n155), .B2(u1_srl_151_n174), .C1(u1_srl_151_n157), .C2(
        u1_srl_151_n175), .ZN(u1_srl_151_n172) );
  OAI211_X1 u1_srl_151_U168 ( .C1(u1_srl_151_n58), .C2(u1_srl_151_n112), .A(
        u1_srl_151_n171), .B(u1_srl_151_n172), .ZN(u1_adj_op_out_sft_7_) );
  AOI22_X1 u1_srl_151_U167 ( .A1(u1_srl_151_n159), .A2(u1_srl_151_n60), .B1(
        u1_srl_151_n160), .B2(u1_srl_151_n169), .ZN(u1_srl_151_n164) );
  AOI222_X1 u1_srl_151_U166 ( .A1(u1_srl_151_n153), .A2(u1_srl_151_n166), .B1(
        u1_srl_151_n155), .B2(u1_srl_151_n167), .C1(u1_srl_151_n157), .C2(
        u1_srl_151_n168), .ZN(u1_srl_151_n165) );
  OAI211_X1 u1_srl_151_U165 ( .C1(u1_srl_151_n163), .C2(u1_srl_151_n110), .A(
        u1_srl_151_n164), .B(u1_srl_151_n165), .ZN(u1_adj_op_out_sft_8_) );
  AOI22_X1 u1_srl_151_U164 ( .A1(u1_srl_151_n159), .A2(u1_srl_151_n61), .B1(
        u1_srl_151_n160), .B2(u1_srl_151_n161), .ZN(u1_srl_151_n151) );
  AOI222_X1 u1_srl_151_U163 ( .A1(u1_srl_151_n153), .A2(u1_srl_151_n154), .B1(
        u1_srl_151_n155), .B2(u1_srl_151_n156), .C1(u1_srl_151_n157), .C2(
        u1_srl_151_n158), .ZN(u1_srl_151_n152) );
  OAI211_X1 u1_srl_151_U162 ( .C1(u1_srl_151_n150), .C2(u1_srl_151_n110), .A(
        u1_srl_151_n151), .B(u1_srl_151_n152), .ZN(u1_adj_op_out_sft_9_) );
  INV_X4 u1_srl_151_U161 ( .A(u1_adj_op_10_), .ZN(u1_srl_151_n149) );
  INV_X4 u1_srl_151_U160 ( .A(u1_adj_op_11_), .ZN(u1_srl_151_n148) );
  INV_X4 u1_srl_151_U159 ( .A(n8505), .ZN(u1_srl_151_n147) );
  INV_X4 u1_srl_151_U158 ( .A(n8504), .ZN(u1_srl_151_n146) );
  INV_X4 u1_srl_151_U157 ( .A(n8503), .ZN(u1_srl_151_n145) );
  INV_X4 u1_srl_151_U156 ( .A(u1_adj_op_15_), .ZN(u1_srl_151_n144) );
  INV_X4 u1_srl_151_U155 ( .A(u1_adj_op_16_), .ZN(u1_srl_151_n143) );
  INV_X4 u1_srl_151_U154 ( .A(u1_adj_op_17_), .ZN(u1_srl_151_n142) );
  INV_X4 u1_srl_151_U153 ( .A(n8502), .ZN(u1_srl_151_n141) );
  INV_X4 u1_srl_151_U152 ( .A(n8501), .ZN(u1_srl_151_n140) );
  INV_X4 u1_srl_151_U151 ( .A(n8500), .ZN(u1_srl_151_n139) );
  INV_X4 u1_srl_151_U150 ( .A(u1_adj_op_20_), .ZN(u1_srl_151_n138) );
  INV_X4 u1_srl_151_U149 ( .A(u1_adj_op_21_), .ZN(u1_srl_151_n137) );
  INV_X4 u1_srl_151_U148 ( .A(u1_adj_op_22_), .ZN(u1_srl_151_n136) );
  INV_X4 u1_srl_151_U147 ( .A(n8499), .ZN(u1_srl_151_n135) );
  INV_X4 u1_srl_151_U146 ( .A(n8498), .ZN(u1_srl_151_n134) );
  INV_X4 u1_srl_151_U145 ( .A(n8497), .ZN(u1_srl_151_n133) );
  INV_X4 u1_srl_151_U144 ( .A(n8496), .ZN(u1_srl_151_n132) );
  INV_X4 u1_srl_151_U143 ( .A(u1_adj_op_27_), .ZN(u1_srl_151_n131) );
  INV_X4 u1_srl_151_U142 ( .A(u1_adj_op_28_), .ZN(u1_srl_151_n130) );
  INV_X4 u1_srl_151_U141 ( .A(n8495), .ZN(u1_srl_151_n129) );
  INV_X4 u1_srl_151_U140 ( .A(n8494), .ZN(u1_srl_151_n128) );
  INV_X4 u1_srl_151_U139 ( .A(n8493), .ZN(u1_srl_151_n127) );
  INV_X4 u1_srl_151_U138 ( .A(n8492), .ZN(u1_srl_151_n126) );
  INV_X4 u1_srl_151_U137 ( .A(u1_adj_op_32_), .ZN(u1_srl_151_n125) );
  INV_X4 u1_srl_151_U136 ( .A(n8491), .ZN(u1_srl_151_n124) );
  INV_X4 u1_srl_151_U135 ( .A(n8490), .ZN(u1_srl_151_n123) );
  INV_X4 u1_srl_151_U134 ( .A(n8489), .ZN(u1_srl_151_n122) );
  INV_X4 u1_srl_151_U133 ( .A(u1_adj_op_36_), .ZN(u1_srl_151_n121) );
  INV_X4 u1_srl_151_U132 ( .A(u1_adj_op_37_), .ZN(u1_srl_151_n120) );
  INV_X4 u1_srl_151_U131 ( .A(u1_adj_op_3_), .ZN(u1_srl_151_n119) );
  INV_X4 u1_srl_151_U130 ( .A(n8479), .ZN(u1_srl_151_n118) );
  INV_X4 u1_srl_151_U129 ( .A(n8477), .ZN(u1_srl_151_n117) );
  INV_X4 u1_srl_151_U128 ( .A(n8476), .ZN(u1_srl_151_n116) );
  INV_X4 u1_srl_151_U127 ( .A(n8475), .ZN(u1_srl_151_n115) );
  INV_X4 u1_srl_151_U126 ( .A(n8474), .ZN(u1_srl_151_n114) );
  INV_X4 u1_srl_151_U125 ( .A(n8473), .ZN(u1_srl_151_n113) );
  INV_X4 u1_srl_151_U124 ( .A(n8470), .ZN(u1_srl_151_n112) );
  INV_X4 u1_srl_151_U123 ( .A(n8469), .ZN(u1_srl_151_n111) );
  INV_X4 u1_srl_151_U122 ( .A(u1_srl_151_n159), .ZN(u1_srl_151_n109) );
  INV_X4 u1_srl_151_U121 ( .A(n8468), .ZN(u1_srl_151_n108) );
  INV_X4 u1_srl_151_U120 ( .A(n8467), .ZN(u1_srl_151_n107) );
  INV_X4 u1_srl_151_U119 ( .A(u1_srl_151_n317), .ZN(u1_srl_151_n106) );
  INV_X4 u1_srl_151_U118 ( .A(u1_srl_151_n281), .ZN(u1_srl_151_n105) );
  INV_X4 u1_srl_151_U117 ( .A(u1_srl_151_n192), .ZN(u1_srl_151_n104) );
  INV_X4 u1_srl_151_U116 ( .A(u1_srl_151_n318), .ZN(u1_srl_151_n103) );
  INV_X4 u1_srl_151_U115 ( .A(u1_srl_151_n248), .ZN(u1_srl_151_n102) );
  INV_X4 u1_srl_151_U114 ( .A(u1_srl_151_n253), .ZN(u1_srl_151_n101) );
  INV_X4 u1_srl_151_U113 ( .A(u1_srl_151_n321), .ZN(u1_srl_151_n100) );
  INV_X4 u1_srl_151_U112 ( .A(u1_srl_151_n282), .ZN(u1_srl_151_n99) );
  INV_X4 u1_srl_151_U111 ( .A(u1_srl_151_n175), .ZN(u1_srl_151_n98) );
  INV_X4 u1_srl_151_U110 ( .A(u1_srl_151_n334), .ZN(u1_srl_151_n97) );
  INV_X4 u1_srl_151_U109 ( .A(u1_srl_151_n335), .ZN(u1_srl_151_n96) );
  INV_X4 u1_srl_151_U108 ( .A(u1_srl_151_n336), .ZN(u1_srl_151_n95) );
  INV_X4 u1_srl_151_U107 ( .A(u1_srl_151_n269), .ZN(u1_srl_151_n94) );
  INV_X4 u1_srl_151_U106 ( .A(u1_srl_151_n296), .ZN(u1_srl_151_n93) );
  INV_X4 u1_srl_151_U105 ( .A(u1_srl_151_n339), .ZN(u1_srl_151_n92) );
  INV_X4 u1_srl_151_U104 ( .A(u1_srl_151_n298), .ZN(u1_srl_151_n91) );
  INV_X4 u1_srl_151_U103 ( .A(u1_srl_151_n263), .ZN(u1_srl_151_n90) );
  INV_X4 u1_srl_151_U102 ( .A(u1_srl_151_n294), .ZN(u1_srl_151_n89) );
  INV_X4 u1_srl_151_U101 ( .A(u1_srl_151_n349), .ZN(u1_srl_151_n88) );
  INV_X4 u1_srl_151_U100 ( .A(u1_srl_151_n277), .ZN(u1_srl_151_n87) );
  INV_X4 u1_srl_151_U99 ( .A(u1_srl_151_n191), .ZN(u1_srl_151_n86) );
  INV_X4 u1_srl_151_U98 ( .A(u1_srl_151_n350), .ZN(u1_srl_151_n85) );
  INV_X4 u1_srl_151_U97 ( .A(u1_srl_151_n301), .ZN(u1_srl_151_n84) );
  INV_X4 u1_srl_151_U96 ( .A(u1_srl_151_n351), .ZN(u1_srl_151_n83) );
  INV_X4 u1_srl_151_U95 ( .A(u1_srl_151_n278), .ZN(u1_srl_151_n82) );
  INV_X4 u1_srl_151_U94 ( .A(u1_srl_151_n363), .ZN(u1_srl_151_n81) );
  INV_X4 u1_srl_151_U93 ( .A(u1_srl_151_n193), .ZN(u1_srl_151_n80) );
  INV_X4 u1_srl_151_U92 ( .A(u1_srl_151_n364), .ZN(u1_srl_151_n79) );
  INV_X4 u1_srl_151_U91 ( .A(u1_srl_151_n256), .ZN(u1_srl_151_n78) );
  INV_X4 u1_srl_151_U90 ( .A(u1_srl_151_n366), .ZN(u1_srl_151_n77) );
  INV_X4 u1_srl_151_U89 ( .A(u1_srl_151_n327), .ZN(u1_srl_151_n76) );
  INV_X4 u1_srl_151_U88 ( .A(u1_srl_151_n367), .ZN(u1_srl_151_n75) );
  INV_X4 u1_srl_151_U87 ( .A(u1_srl_151_n285), .ZN(u1_srl_151_n74) );
  INV_X4 u1_srl_151_U86 ( .A(n8465), .ZN(u1_srl_151_n73) );
  INV_X4 u1_srl_151_U85 ( .A(u1_srl_151_n251), .ZN(u1_srl_151_n71) );
  INV_X4 u1_srl_151_U84 ( .A(u1_srl_151_n259), .ZN(u1_srl_151_n70) );
  INV_X4 u1_srl_151_U83 ( .A(u1_srl_151_n272), .ZN(u1_srl_151_n69) );
  INV_X4 u1_srl_151_U82 ( .A(u1_srl_151_n279), .ZN(u1_srl_151_n68) );
  INV_X4 u1_srl_151_U81 ( .A(u1_srl_151_n283), .ZN(u1_srl_151_n67) );
  INV_X4 u1_srl_151_U80 ( .A(u1_srl_151_n299), .ZN(u1_srl_151_n66) );
  INV_X4 u1_srl_151_U79 ( .A(u1_srl_151_n302), .ZN(u1_srl_151_n65) );
  INV_X4 u1_srl_151_U78 ( .A(u1_srl_151_n310), .ZN(u1_srl_151_n64) );
  INV_X4 u1_srl_151_U77 ( .A(u1_srl_151_n326), .ZN(u1_srl_151_n63) );
  INV_X4 u1_srl_151_U76 ( .A(u1_srl_151_n352), .ZN(u1_srl_151_n62) );
  INV_X4 u1_srl_151_U75 ( .A(u1_srl_151_n162), .ZN(u1_srl_151_n61) );
  INV_X4 u1_srl_151_U74 ( .A(u1_srl_151_n170), .ZN(u1_srl_151_n60) );
  INV_X4 u1_srl_151_U73 ( .A(u1_srl_151_n178), .ZN(u1_srl_151_n59) );
  INV_X4 u1_srl_151_U72 ( .A(u1_srl_151_n217), .ZN(u1_srl_151_n58) );
  INV_X4 u1_srl_151_U71 ( .A(u1_srl_151_n185), .ZN(u1_srl_151_n57) );
  INV_X4 u1_srl_151_U70 ( .A(u1_srl_151_n220), .ZN(u1_srl_151_n56) );
  INV_X4 u1_srl_151_U69 ( .A(u1_srl_151_n189), .ZN(u1_srl_151_n55) );
  INV_X4 u1_srl_151_U68 ( .A(u1_srl_151_n222), .ZN(u1_srl_151_n54) );
  INV_X4 u1_srl_151_U67 ( .A(u1_srl_151_n199), .ZN(u1_srl_151_n53) );
  INV_X4 u1_srl_151_U66 ( .A(u1_srl_151_n224), .ZN(u1_srl_151_n52) );
  INV_X4 u1_srl_151_U65 ( .A(u1_srl_151_n215), .ZN(u1_srl_151_n51) );
  INV_X4 u1_srl_151_U64 ( .A(u1_srl_151_n216), .ZN(u1_srl_151_n50) );
  INV_X4 u1_srl_151_U63 ( .A(u1_srl_151_n241), .ZN(u1_srl_151_n49) );
  INV_X4 u1_srl_151_U62 ( .A(u1_srl_151_n228), .ZN(u1_srl_151_n48) );
  INV_X4 u1_srl_151_U61 ( .A(u1_srl_151_n292), .ZN(u1_srl_151_n47) );
  INV_X4 u1_srl_151_U60 ( .A(u1_srl_151_n229), .ZN(u1_srl_151_n46) );
  INV_X4 u1_srl_151_U59 ( .A(u1_srl_151_n202), .ZN(u1_srl_151_n45) );
  INV_X4 u1_srl_151_U58 ( .A(u1_srl_151_n203), .ZN(u1_srl_151_n44) );
  INV_X4 u1_srl_151_U57 ( .A(u1_srl_151_n204), .ZN(u1_srl_151_n43) );
  INV_X4 u1_srl_151_U56 ( .A(u1_srl_151_n205), .ZN(u1_srl_151_n42) );
  INV_X4 u1_srl_151_U55 ( .A(u1_srl_151_n232), .ZN(u1_srl_151_n41) );
  INV_X4 u1_srl_151_U54 ( .A(u1_srl_151_n245), .ZN(u1_srl_151_n40) );
  INV_X4 u1_srl_151_U53 ( .A(u1_srl_151_n160), .ZN(u1_srl_151_n39) );
  INV_X4 u1_srl_151_U52 ( .A(u1_srl_151_n287), .ZN(u1_srl_151_n38) );
  INV_X4 u1_srl_151_U51 ( .A(u1_srl_151_n358), .ZN(u1_srl_151_n37) );
  INV_X4 u1_srl_151_U50 ( .A(u1_srl_151_n230), .ZN(u1_srl_151_n36) );
  INV_X4 u1_srl_151_U49 ( .A(u1_srl_151_n371), .ZN(u1_srl_151_n35) );
  INV_X4 u1_srl_151_U48 ( .A(u1_srl_151_n304), .ZN(u1_srl_151_n34) );
  INV_X32 u1_srl_151_U47 ( .A(u1_srl_151_n28), .ZN(u1_srl_151_n25) );
  INV_X32 u1_srl_151_U46 ( .A(u1_srl_151_n22), .ZN(u1_srl_151_n20) );
  INV_X32 u1_srl_151_U45 ( .A(u1_srl_151_n22), .ZN(u1_srl_151_n19) );
  INV_X32 u1_srl_151_U44 ( .A(u1_srl_151_n22), .ZN(u1_srl_151_n17) );
  NOR2_X4 u1_srl_151_U43 ( .A1(u1_srl_151_n107), .A2(n8466), .ZN(
        u1_srl_151_n239) );
  NOR2_X4 u1_srl_151_U42 ( .A1(u1_srl_151_n108), .A2(u1_srl_151_n73), .ZN(
        u1_srl_151_n252) );
  NOR2_X4 u1_srl_151_U41 ( .A1(u1_srl_151_n108), .A2(n8465), .ZN(
        u1_srl_151_n210) );
  NOR2_X4 u1_srl_151_U40 ( .A1(u1_srl_151_n1), .A2(u1_srl_151_n11), .ZN(
        u1_srl_151_n153) );
  NOR2_X4 u1_srl_151_U39 ( .A1(u1_srl_151_n112), .A2(n8469), .ZN(
        u1_srl_151_n159) );
  NOR2_X4 u1_srl_151_U38 ( .A1(u1_srl_151_n4), .A2(u1_srl_151_n9), .ZN(
        u1_srl_151_n157) );
  NOR2_X4 u1_srl_151_U37 ( .A1(u1_srl_151_n10), .A2(u1_srl_151_n72), .ZN(
        u1_srl_151_n155) );
  NOR2_X4 u1_srl_151_U36 ( .A1(u1_srl_151_n32), .A2(u1_srl_151_n10), .ZN(
        u1_srl_151_n160) );
  INV_X8 u1_srl_151_U35 ( .A(u1_srl_151_n177), .ZN(u1_srl_151_n110) );
  INV_X16 u1_srl_151_U34 ( .A(u1_srl_151_n252), .ZN(u1_srl_151_n72) );
  INV_X16 u1_srl_151_U33 ( .A(u1_srl_151_n213), .ZN(u1_srl_151_n22) );
  INV_X8 u1_srl_151_U32 ( .A(u1_srl_151_n23), .ZN(u1_srl_151_n28) );
  INV_X4 u1_srl_151_U31 ( .A(u1_srl_151_n3), .ZN(u1_srl_151_n23) );
  INV_X8 u1_srl_151_U30 ( .A(u1_srl_151_n210), .ZN(u1_srl_151_n4) );
  INV_X4 u1_srl_151_U29 ( .A(u1_srl_151_n4), .ZN(u1_srl_151_n5) );
  INV_X8 u1_srl_151_U28 ( .A(u1_srl_151_n211), .ZN(u1_srl_151_n16) );
  NOR2_X2 u1_srl_151_U27 ( .A1(n8465), .A2(n8468), .ZN(u1_srl_151_n226) );
  AND2_X2 u1_srl_151_U26 ( .A1(n8466), .A2(n8467), .ZN(u1_srl_151_n213) );
  OR2_X4 u1_srl_151_U25 ( .A1(n8467), .A2(n8466), .ZN(u1_srl_151_n3) );
  INV_X4 u1_srl_151_U24 ( .A(u1_srl_151_n2), .ZN(u1_srl_151_n9) );
  INV_X16 u1_srl_151_U23 ( .A(u1_srl_151_n28), .ZN(u1_srl_151_n27) );
  INV_X4 u1_srl_151_U22 ( .A(u1_srl_151_n226), .ZN(u1_srl_151_n32) );
  INV_X4 u1_srl_151_U21 ( .A(u1_srl_151_n226), .ZN(u1_srl_151_n33) );
  INV_X16 u1_srl_151_U20 ( .A(u1_srl_151_n16), .ZN(u1_srl_151_n14) );
  INV_X16 u1_srl_151_U19 ( .A(u1_srl_151_n8), .ZN(u1_srl_151_n6) );
  AND2_X4 u1_srl_151_U18 ( .A1(u1_srl_151_n111), .A2(u1_srl_151_n112), .ZN(
        u1_srl_151_n2) );
  INV_X8 u1_srl_151_U17 ( .A(u1_srl_151_n239), .ZN(u1_srl_151_n8) );
  OR2_X4 u1_srl_151_U16 ( .A1(u1_srl_151_n73), .A2(n8468), .ZN(u1_srl_151_n1)
         );
  INV_X8 u1_srl_151_U15 ( .A(u1_srl_151_n2), .ZN(u1_srl_151_n11) );
  INV_X4 u1_srl_151_U14 ( .A(u1_srl_151_n2), .ZN(u1_srl_151_n10) );
  INV_X16 u1_srl_151_U13 ( .A(u1_srl_151_n1), .ZN(u1_srl_151_n13) );
  INV_X8 u1_srl_151_U12 ( .A(u1_srl_151_n33), .ZN(u1_srl_151_n31) );
  INV_X16 u1_srl_151_U11 ( .A(u1_srl_151_n6), .ZN(u1_srl_151_n7) );
  INV_X16 u1_srl_151_U10 ( .A(u1_srl_151_n28), .ZN(u1_srl_151_n26) );
  INV_X8 u1_srl_151_U9 ( .A(u1_srl_151_n22), .ZN(u1_srl_151_n21) );
  INV_X16 u1_srl_151_U8 ( .A(u1_srl_151_n22), .ZN(u1_srl_151_n18) );
  INV_X16 u1_srl_151_U7 ( .A(u1_srl_151_n16), .ZN(u1_srl_151_n15) );
  INV_X16 u1_srl_151_U6 ( .A(u1_srl_151_n28), .ZN(u1_srl_151_n24) );
  INV_X8 u1_srl_151_U5 ( .A(u1_srl_151_n1), .ZN(u1_srl_151_n12) );
  INV_X8 u1_srl_151_U4 ( .A(u1_srl_151_n32), .ZN(u1_srl_151_n29) );
  INV_X8 u1_srl_151_U3 ( .A(u1_srl_151_n32), .ZN(u1_srl_151_n30) );
  INV_X4 sub_1_root_u1_sub_133_aco_U12 ( .A(u1_N46), .ZN(
        sub_1_root_u1_sub_133_aco_n12) );
  INV_X4 sub_1_root_u1_sub_133_aco_U11 ( .A(u1_exp_small[0]), .ZN(
        sub_1_root_u1_sub_133_aco_n11) );
  INV_X4 sub_1_root_u1_sub_133_aco_U10 ( .A(u1_exp_small[10]), .ZN(
        sub_1_root_u1_sub_133_aco_n10) );
  INV_X4 sub_1_root_u1_sub_133_aco_U9 ( .A(u1_exp_small[1]), .ZN(
        sub_1_root_u1_sub_133_aco_n9) );
  INV_X4 sub_1_root_u1_sub_133_aco_U8 ( .A(u1_exp_small[2]), .ZN(
        sub_1_root_u1_sub_133_aco_n8) );
  INV_X4 sub_1_root_u1_sub_133_aco_U7 ( .A(u1_exp_small[3]), .ZN(
        sub_1_root_u1_sub_133_aco_n7) );
  INV_X4 sub_1_root_u1_sub_133_aco_U6 ( .A(u1_exp_small[4]), .ZN(
        sub_1_root_u1_sub_133_aco_n6) );
  INV_X4 sub_1_root_u1_sub_133_aco_U5 ( .A(u1_exp_small[5]), .ZN(
        sub_1_root_u1_sub_133_aco_n5) );
  INV_X4 sub_1_root_u1_sub_133_aco_U4 ( .A(u1_exp_small[6]), .ZN(
        sub_1_root_u1_sub_133_aco_n4) );
  INV_X4 sub_1_root_u1_sub_133_aco_U3 ( .A(u1_exp_small[7]), .ZN(
        sub_1_root_u1_sub_133_aco_n3) );
  INV_X4 sub_1_root_u1_sub_133_aco_U2 ( .A(n8472), .ZN(
        sub_1_root_u1_sub_133_aco_n2) );
  INV_X4 sub_1_root_u1_sub_133_aco_U1 ( .A(n8471), .ZN(
        sub_1_root_u1_sub_133_aco_n1) );
  FA_X1 sub_1_root_u1_sub_133_aco_U2_0 ( .A(u1_exp_large_0_), .B(
        sub_1_root_u1_sub_133_aco_n11), .CI(sub_1_root_u1_sub_133_aco_n12), 
        .CO(sub_1_root_u1_sub_133_aco_carry[1]), .S(u1_exp_diff2[0]) );
  FA_X1 sub_1_root_u1_sub_133_aco_U2_1 ( .A(u1_exp_large_1_), .B(
        sub_1_root_u1_sub_133_aco_n9), .CI(sub_1_root_u1_sub_133_aco_carry[1]), 
        .CO(sub_1_root_u1_sub_133_aco_carry[2]), .S(u1_exp_diff2[1]) );
  FA_X1 sub_1_root_u1_sub_133_aco_U2_2 ( .A(u1_exp_large_2_), .B(
        sub_1_root_u1_sub_133_aco_n8), .CI(sub_1_root_u1_sub_133_aco_carry[2]), 
        .CO(sub_1_root_u1_sub_133_aco_carry[3]), .S(u1_exp_diff2[2]) );
  FA_X1 sub_1_root_u1_sub_133_aco_U2_3 ( .A(u1_exp_large_3_), .B(
        sub_1_root_u1_sub_133_aco_n7), .CI(sub_1_root_u1_sub_133_aco_carry[3]), 
        .CO(sub_1_root_u1_sub_133_aco_carry[4]), .S(u1_exp_diff2[3]) );
  FA_X1 sub_1_root_u1_sub_133_aco_U2_4 ( .A(u1_exp_large_4_), .B(
        sub_1_root_u1_sub_133_aco_n6), .CI(sub_1_root_u1_sub_133_aco_carry[4]), 
        .CO(sub_1_root_u1_sub_133_aco_carry[5]), .S(u1_exp_diff2[4]) );
  FA_X1 sub_1_root_u1_sub_133_aco_U2_5 ( .A(u1_exp_large_5_), .B(
        sub_1_root_u1_sub_133_aco_n5), .CI(sub_1_root_u1_sub_133_aco_carry[5]), 
        .CO(sub_1_root_u1_sub_133_aco_carry[6]), .S(u1_exp_diff2[5]) );
  FA_X1 sub_1_root_u1_sub_133_aco_U2_6 ( .A(u1_exp_large_6_), .B(
        sub_1_root_u1_sub_133_aco_n4), .CI(sub_1_root_u1_sub_133_aco_carry[6]), 
        .CO(sub_1_root_u1_sub_133_aco_carry[7]), .S(u1_exp_diff2[6]) );
  FA_X1 sub_1_root_u1_sub_133_aco_U2_7 ( .A(u1_exp_large_7_), .B(
        sub_1_root_u1_sub_133_aco_n3), .CI(sub_1_root_u1_sub_133_aco_carry[7]), 
        .CO(sub_1_root_u1_sub_133_aco_carry[8]), .S(u1_exp_diff2[7]) );
  FA_X1 sub_1_root_u1_sub_133_aco_U2_8 ( .A(n8507), .B(
        sub_1_root_u1_sub_133_aco_n2), .CI(sub_1_root_u1_sub_133_aco_carry[8]), 
        .CO(sub_1_root_u1_sub_133_aco_carry[9]), .S(u1_exp_diff2[8]) );
  FA_X1 sub_1_root_u1_sub_133_aco_U2_9 ( .A(n8506), .B(
        sub_1_root_u1_sub_133_aco_n1), .CI(sub_1_root_u1_sub_133_aco_carry[9]), 
        .CO(sub_1_root_u1_sub_133_aco_carry[10]), .S(u1_exp_diff2[9]) );
  FA_X1 sub_1_root_u1_sub_133_aco_U2_10 ( .A(u1_exp_large_10_), .B(
        sub_1_root_u1_sub_133_aco_n10), .CI(
        sub_1_root_u1_sub_133_aco_carry[10]), .S(u1_exp_diff2[10]) );
  INV_X4 sub_436_3_U259 ( .A(N343), .ZN(sub_436_3_n171) );
  INV_X4 sub_436_3_U258 ( .A(opa_r1[1]), .ZN(sub_436_3_n170) );
  INV_X4 sub_436_3_U257 ( .A(opa_r1[2]), .ZN(sub_436_3_n169) );
  INV_X4 sub_436_3_U256 ( .A(opa_r1[3]), .ZN(sub_436_3_n168) );
  INV_X4 sub_436_3_U255 ( .A(opa_r1[4]), .ZN(sub_436_3_n167) );
  INV_X4 sub_436_3_U254 ( .A(opa_r1[5]), .ZN(sub_436_3_n166) );
  INV_X4 sub_436_3_U253 ( .A(opa_r1[6]), .ZN(sub_436_3_n165) );
  INV_X4 sub_436_3_U252 ( .A(opa_r1[7]), .ZN(sub_436_3_n164) );
  INV_X4 sub_436_3_U251 ( .A(opa_r1[8]), .ZN(sub_436_3_n163) );
  INV_X4 sub_436_3_U250 ( .A(opa_r1[9]), .ZN(sub_436_3_n162) );
  INV_X4 sub_436_3_U249 ( .A(opa_r1[10]), .ZN(sub_436_3_n161) );
  INV_X4 sub_436_3_U248 ( .A(opa_r1[11]), .ZN(sub_436_3_n160) );
  INV_X4 sub_436_3_U247 ( .A(opa_r1[12]), .ZN(sub_436_3_n159) );
  INV_X4 sub_436_3_U246 ( .A(opa_r1[13]), .ZN(sub_436_3_n158) );
  INV_X4 sub_436_3_U245 ( .A(opa_r1[14]), .ZN(sub_436_3_n157) );
  INV_X4 sub_436_3_U244 ( .A(opa_r1[15]), .ZN(sub_436_3_n156) );
  INV_X4 sub_436_3_U243 ( .A(opa_r1[16]), .ZN(sub_436_3_n155) );
  INV_X4 sub_436_3_U242 ( .A(opa_r1[17]), .ZN(sub_436_3_n154) );
  INV_X4 sub_436_3_U241 ( .A(opa_r1[18]), .ZN(sub_436_3_n153) );
  INV_X4 sub_436_3_U240 ( .A(opa_r1[19]), .ZN(sub_436_3_n152) );
  INV_X4 sub_436_3_U239 ( .A(opa_r1[20]), .ZN(sub_436_3_n151) );
  INV_X4 sub_436_3_U238 ( .A(opa_r1[21]), .ZN(sub_436_3_n150) );
  INV_X4 sub_436_3_U237 ( .A(opa_r1[22]), .ZN(sub_436_3_n149) );
  INV_X4 sub_436_3_U236 ( .A(opa_r1[23]), .ZN(sub_436_3_n148) );
  INV_X4 sub_436_3_U235 ( .A(opa_r1[24]), .ZN(sub_436_3_n147) );
  INV_X4 sub_436_3_U234 ( .A(opa_r1[25]), .ZN(sub_436_3_n146) );
  INV_X4 sub_436_3_U233 ( .A(opa_r1[26]), .ZN(sub_436_3_n145) );
  INV_X4 sub_436_3_U232 ( .A(opa_r1[27]), .ZN(sub_436_3_n144) );
  INV_X4 sub_436_3_U231 ( .A(opa_r1[28]), .ZN(sub_436_3_n143) );
  INV_X4 sub_436_3_U230 ( .A(opa_r1[29]), .ZN(sub_436_3_n142) );
  INV_X4 sub_436_3_U229 ( .A(opa_r1[30]), .ZN(sub_436_3_n141) );
  INV_X4 sub_436_3_U228 ( .A(opa_r1[31]), .ZN(sub_436_3_n140) );
  INV_X4 sub_436_3_U227 ( .A(opa_r1[32]), .ZN(sub_436_3_n139) );
  INV_X4 sub_436_3_U226 ( .A(opa_r1[33]), .ZN(sub_436_3_n138) );
  INV_X4 sub_436_3_U225 ( .A(opa_r1[34]), .ZN(sub_436_3_n137) );
  INV_X4 sub_436_3_U224 ( .A(opa_r1[35]), .ZN(sub_436_3_n136) );
  INV_X4 sub_436_3_U223 ( .A(opa_r1[36]), .ZN(sub_436_3_n135) );
  INV_X4 sub_436_3_U222 ( .A(opa_r1[37]), .ZN(sub_436_3_n134) );
  INV_X4 sub_436_3_U221 ( .A(opa_r1[38]), .ZN(sub_436_3_n133) );
  INV_X4 sub_436_3_U220 ( .A(opa_r1[39]), .ZN(sub_436_3_n132) );
  INV_X4 sub_436_3_U219 ( .A(opa_r1[40]), .ZN(sub_436_3_n131) );
  INV_X4 sub_436_3_U218 ( .A(opa_r1[41]), .ZN(sub_436_3_n130) );
  INV_X4 sub_436_3_U217 ( .A(opa_r1[42]), .ZN(sub_436_3_n129) );
  INV_X4 sub_436_3_U216 ( .A(opa_r1[43]), .ZN(sub_436_3_n128) );
  INV_X4 sub_436_3_U215 ( .A(opa_r1[44]), .ZN(sub_436_3_n127) );
  INV_X4 sub_436_3_U214 ( .A(opa_r1[45]), .ZN(sub_436_3_n126) );
  INV_X4 sub_436_3_U213 ( .A(opa_r1[46]), .ZN(sub_436_3_n125) );
  INV_X4 sub_436_3_U212 ( .A(opa_r1[47]), .ZN(sub_436_3_n124) );
  INV_X4 sub_436_3_U211 ( .A(opa_r1[48]), .ZN(sub_436_3_n123) );
  INV_X4 sub_436_3_U210 ( .A(opa_r1[49]), .ZN(sub_436_3_n122) );
  INV_X4 sub_436_3_U209 ( .A(opa_r1[50]), .ZN(sub_436_3_n121) );
  INV_X4 sub_436_3_U208 ( .A(opa_r1[51]), .ZN(sub_436_3_n120) );
  INV_X4 sub_436_3_U207 ( .A(opa_r1[52]), .ZN(sub_436_3_n119) );
  INV_X4 sub_436_3_U206 ( .A(opa_r1[53]), .ZN(sub_436_3_n118) );
  INV_X4 sub_436_3_U205 ( .A(opa_r1[54]), .ZN(sub_436_3_n117) );
  INV_X4 sub_436_3_U204 ( .A(opa_r1[55]), .ZN(sub_436_3_n116) );
  INV_X4 sub_436_3_U203 ( .A(opa_r1[56]), .ZN(sub_436_3_n115) );
  INV_X4 sub_436_3_U202 ( .A(opa_r1[57]), .ZN(sub_436_3_n114) );
  INV_X4 sub_436_3_U201 ( .A(sub_436_3_n113), .ZN(sub_436_3_carry_50_) );
  NAND2_X2 sub_436_3_U200 ( .A1(sub_436_3_n170), .A2(sub_436_3_n171), .ZN(
        sub_436_3_n113) );
  INV_X4 sub_436_3_U199 ( .A(sub_436_3_n112), .ZN(sub_436_3_carry_51_) );
  NAND2_X2 sub_436_3_U198 ( .A1(sub_436_3_n169), .A2(sub_436_3_carry_50_), 
        .ZN(sub_436_3_n112) );
  INV_X4 sub_436_3_U197 ( .A(sub_436_3_n111), .ZN(sub_436_3_carry_52_) );
  NAND2_X2 sub_436_3_U196 ( .A1(sub_436_3_n168), .A2(sub_436_3_carry_51_), 
        .ZN(sub_436_3_n111) );
  INV_X4 sub_436_3_U195 ( .A(sub_436_3_n110), .ZN(sub_436_3_carry_53_) );
  NAND2_X2 sub_436_3_U194 ( .A1(sub_436_3_n167), .A2(sub_436_3_carry_52_), 
        .ZN(sub_436_3_n110) );
  INV_X4 sub_436_3_U193 ( .A(sub_436_3_n109), .ZN(sub_436_3_carry_54_) );
  NAND2_X2 sub_436_3_U192 ( .A1(sub_436_3_n166), .A2(sub_436_3_carry_53_), 
        .ZN(sub_436_3_n109) );
  INV_X4 sub_436_3_U191 ( .A(sub_436_3_n108), .ZN(sub_436_3_carry_55_) );
  NAND2_X2 sub_436_3_U190 ( .A1(sub_436_3_n165), .A2(sub_436_3_carry_54_), 
        .ZN(sub_436_3_n108) );
  INV_X4 sub_436_3_U189 ( .A(sub_436_3_n107), .ZN(sub_436_3_carry_56_) );
  NAND2_X2 sub_436_3_U188 ( .A1(sub_436_3_n164), .A2(sub_436_3_carry_55_), 
        .ZN(sub_436_3_n107) );
  INV_X4 sub_436_3_U187 ( .A(sub_436_3_n106), .ZN(sub_436_3_carry_57_) );
  NAND2_X2 sub_436_3_U186 ( .A1(sub_436_3_n163), .A2(sub_436_3_carry_56_), 
        .ZN(sub_436_3_n106) );
  INV_X4 sub_436_3_U185 ( .A(sub_436_3_n105), .ZN(sub_436_3_carry_58_) );
  NAND2_X2 sub_436_3_U184 ( .A1(sub_436_3_n162), .A2(sub_436_3_carry_57_), 
        .ZN(sub_436_3_n105) );
  INV_X4 sub_436_3_U183 ( .A(sub_436_3_n104), .ZN(sub_436_3_carry_59_) );
  NAND2_X2 sub_436_3_U182 ( .A1(sub_436_3_n161), .A2(sub_436_3_carry_58_), 
        .ZN(sub_436_3_n104) );
  INV_X4 sub_436_3_U181 ( .A(sub_436_3_n103), .ZN(sub_436_3_carry_60_) );
  NAND2_X2 sub_436_3_U180 ( .A1(sub_436_3_n160), .A2(sub_436_3_carry_59_), 
        .ZN(sub_436_3_n103) );
  INV_X4 sub_436_3_U179 ( .A(sub_436_3_n102), .ZN(sub_436_3_carry_61_) );
  NAND2_X2 sub_436_3_U178 ( .A1(sub_436_3_n159), .A2(sub_436_3_carry_60_), 
        .ZN(sub_436_3_n102) );
  INV_X4 sub_436_3_U177 ( .A(sub_436_3_n101), .ZN(sub_436_3_carry_62_) );
  NAND2_X2 sub_436_3_U176 ( .A1(sub_436_3_n158), .A2(sub_436_3_carry_61_), 
        .ZN(sub_436_3_n101) );
  INV_X4 sub_436_3_U175 ( .A(sub_436_3_n100), .ZN(sub_436_3_carry_63_) );
  NAND2_X2 sub_436_3_U174 ( .A1(sub_436_3_n157), .A2(sub_436_3_carry_62_), 
        .ZN(sub_436_3_n100) );
  INV_X4 sub_436_3_U173 ( .A(sub_436_3_n99), .ZN(sub_436_3_carry_64_) );
  NAND2_X2 sub_436_3_U172 ( .A1(sub_436_3_n156), .A2(sub_436_3_carry_63_), 
        .ZN(sub_436_3_n99) );
  INV_X4 sub_436_3_U171 ( .A(sub_436_3_n98), .ZN(sub_436_3_carry_65_) );
  NAND2_X2 sub_436_3_U170 ( .A1(sub_436_3_n155), .A2(sub_436_3_carry_64_), 
        .ZN(sub_436_3_n98) );
  INV_X4 sub_436_3_U169 ( .A(sub_436_3_n97), .ZN(sub_436_3_carry_66_) );
  NAND2_X2 sub_436_3_U168 ( .A1(sub_436_3_n154), .A2(sub_436_3_carry_65_), 
        .ZN(sub_436_3_n97) );
  INV_X4 sub_436_3_U167 ( .A(sub_436_3_n96), .ZN(sub_436_3_carry_67_) );
  NAND2_X2 sub_436_3_U166 ( .A1(sub_436_3_n153), .A2(sub_436_3_carry_66_), 
        .ZN(sub_436_3_n96) );
  INV_X4 sub_436_3_U165 ( .A(sub_436_3_n95), .ZN(sub_436_3_carry_68_) );
  NAND2_X2 sub_436_3_U164 ( .A1(sub_436_3_n152), .A2(sub_436_3_carry_67_), 
        .ZN(sub_436_3_n95) );
  INV_X4 sub_436_3_U163 ( .A(sub_436_3_n94), .ZN(sub_436_3_carry_69_) );
  NAND2_X2 sub_436_3_U162 ( .A1(sub_436_3_n151), .A2(sub_436_3_carry_68_), 
        .ZN(sub_436_3_n94) );
  INV_X4 sub_436_3_U161 ( .A(sub_436_3_n93), .ZN(sub_436_3_carry_70_) );
  NAND2_X2 sub_436_3_U160 ( .A1(sub_436_3_n150), .A2(sub_436_3_carry_69_), 
        .ZN(sub_436_3_n93) );
  INV_X4 sub_436_3_U159 ( .A(sub_436_3_n92), .ZN(sub_436_3_carry_71_) );
  NAND2_X2 sub_436_3_U158 ( .A1(sub_436_3_n149), .A2(sub_436_3_carry_70_), 
        .ZN(sub_436_3_n92) );
  INV_X4 sub_436_3_U157 ( .A(sub_436_3_n91), .ZN(sub_436_3_carry_72_) );
  NAND2_X2 sub_436_3_U156 ( .A1(sub_436_3_n148), .A2(sub_436_3_carry_71_), 
        .ZN(sub_436_3_n91) );
  INV_X4 sub_436_3_U155 ( .A(sub_436_3_n90), .ZN(sub_436_3_carry_73_) );
  NAND2_X2 sub_436_3_U154 ( .A1(sub_436_3_n147), .A2(sub_436_3_carry_72_), 
        .ZN(sub_436_3_n90) );
  INV_X4 sub_436_3_U153 ( .A(sub_436_3_n89), .ZN(N525) );
  XNOR2_X2 sub_436_3_U152 ( .A(sub_436_3_n146), .B(sub_436_3_carry_73_), .ZN(
        sub_436_3_n89) );
  INV_X4 sub_436_3_U151 ( .A(sub_436_3_n88), .ZN(sub_436_3_carry_74_) );
  NAND2_X2 sub_436_3_U150 ( .A1(sub_436_3_n146), .A2(sub_436_3_carry_73_), 
        .ZN(sub_436_3_n88) );
  INV_X4 sub_436_3_U149 ( .A(sub_436_3_n87), .ZN(N526) );
  XNOR2_X2 sub_436_3_U148 ( .A(sub_436_3_n145), .B(sub_436_3_carry_74_), .ZN(
        sub_436_3_n87) );
  INV_X4 sub_436_3_U147 ( .A(sub_436_3_n86), .ZN(sub_436_3_carry_75_) );
  NAND2_X2 sub_436_3_U146 ( .A1(sub_436_3_n145), .A2(sub_436_3_carry_74_), 
        .ZN(sub_436_3_n86) );
  INV_X4 sub_436_3_U145 ( .A(sub_436_3_n85), .ZN(N527) );
  XNOR2_X2 sub_436_3_U144 ( .A(sub_436_3_n144), .B(sub_436_3_carry_75_), .ZN(
        sub_436_3_n85) );
  INV_X4 sub_436_3_U143 ( .A(sub_436_3_n84), .ZN(sub_436_3_carry_76_) );
  NAND2_X2 sub_436_3_U142 ( .A1(sub_436_3_n144), .A2(sub_436_3_carry_75_), 
        .ZN(sub_436_3_n84) );
  INV_X4 sub_436_3_U141 ( .A(sub_436_3_n83), .ZN(N528) );
  XNOR2_X2 sub_436_3_U140 ( .A(sub_436_3_n143), .B(sub_436_3_carry_76_), .ZN(
        sub_436_3_n83) );
  INV_X4 sub_436_3_U139 ( .A(sub_436_3_n82), .ZN(sub_436_3_carry_77_) );
  NAND2_X2 sub_436_3_U138 ( .A1(sub_436_3_n143), .A2(sub_436_3_carry_76_), 
        .ZN(sub_436_3_n82) );
  INV_X4 sub_436_3_U137 ( .A(sub_436_3_n81), .ZN(N529) );
  XNOR2_X2 sub_436_3_U136 ( .A(sub_436_3_n142), .B(sub_436_3_carry_77_), .ZN(
        sub_436_3_n81) );
  INV_X4 sub_436_3_U135 ( .A(sub_436_3_n80), .ZN(sub_436_3_carry_78_) );
  NAND2_X2 sub_436_3_U134 ( .A1(sub_436_3_n142), .A2(sub_436_3_carry_77_), 
        .ZN(sub_436_3_n80) );
  INV_X4 sub_436_3_U133 ( .A(sub_436_3_n79), .ZN(N530) );
  XNOR2_X2 sub_436_3_U132 ( .A(sub_436_3_n141), .B(sub_436_3_carry_78_), .ZN(
        sub_436_3_n79) );
  INV_X4 sub_436_3_U131 ( .A(sub_436_3_n78), .ZN(sub_436_3_carry_79_) );
  NAND2_X2 sub_436_3_U130 ( .A1(sub_436_3_n141), .A2(sub_436_3_carry_78_), 
        .ZN(sub_436_3_n78) );
  INV_X4 sub_436_3_U129 ( .A(sub_436_3_n77), .ZN(N531) );
  XNOR2_X2 sub_436_3_U128 ( .A(sub_436_3_n140), .B(sub_436_3_carry_79_), .ZN(
        sub_436_3_n77) );
  INV_X4 sub_436_3_U127 ( .A(sub_436_3_n76), .ZN(sub_436_3_carry_80_) );
  NAND2_X2 sub_436_3_U126 ( .A1(sub_436_3_n140), .A2(sub_436_3_carry_79_), 
        .ZN(sub_436_3_n76) );
  INV_X4 sub_436_3_U125 ( .A(sub_436_3_n75), .ZN(N532) );
  XNOR2_X2 sub_436_3_U124 ( .A(sub_436_3_n139), .B(sub_436_3_carry_80_), .ZN(
        sub_436_3_n75) );
  INV_X4 sub_436_3_U123 ( .A(sub_436_3_n74), .ZN(sub_436_3_carry_81_) );
  NAND2_X2 sub_436_3_U122 ( .A1(sub_436_3_n139), .A2(sub_436_3_carry_80_), 
        .ZN(sub_436_3_n74) );
  INV_X4 sub_436_3_U121 ( .A(sub_436_3_n73), .ZN(N533) );
  XNOR2_X2 sub_436_3_U120 ( .A(sub_436_3_n138), .B(sub_436_3_carry_81_), .ZN(
        sub_436_3_n73) );
  INV_X4 sub_436_3_U119 ( .A(sub_436_3_n72), .ZN(sub_436_3_carry_82_) );
  NAND2_X2 sub_436_3_U118 ( .A1(sub_436_3_n138), .A2(sub_436_3_carry_81_), 
        .ZN(sub_436_3_n72) );
  INV_X4 sub_436_3_U117 ( .A(sub_436_3_n71), .ZN(N534) );
  XNOR2_X2 sub_436_3_U116 ( .A(sub_436_3_n137), .B(sub_436_3_carry_82_), .ZN(
        sub_436_3_n71) );
  INV_X4 sub_436_3_U115 ( .A(sub_436_3_n70), .ZN(sub_436_3_carry_83_) );
  NAND2_X2 sub_436_3_U114 ( .A1(sub_436_3_n137), .A2(sub_436_3_carry_82_), 
        .ZN(sub_436_3_n70) );
  INV_X4 sub_436_3_U113 ( .A(sub_436_3_n69), .ZN(N535) );
  XNOR2_X2 sub_436_3_U112 ( .A(sub_436_3_n136), .B(sub_436_3_carry_83_), .ZN(
        sub_436_3_n69) );
  INV_X4 sub_436_3_U111 ( .A(sub_436_3_n68), .ZN(sub_436_3_carry_84_) );
  NAND2_X2 sub_436_3_U110 ( .A1(sub_436_3_n136), .A2(sub_436_3_carry_83_), 
        .ZN(sub_436_3_n68) );
  INV_X4 sub_436_3_U109 ( .A(sub_436_3_n67), .ZN(N536) );
  XNOR2_X2 sub_436_3_U108 ( .A(sub_436_3_n135), .B(sub_436_3_carry_84_), .ZN(
        sub_436_3_n67) );
  INV_X4 sub_436_3_U107 ( .A(sub_436_3_n66), .ZN(sub_436_3_carry_85_) );
  NAND2_X2 sub_436_3_U106 ( .A1(sub_436_3_n135), .A2(sub_436_3_carry_84_), 
        .ZN(sub_436_3_n66) );
  INV_X4 sub_436_3_U105 ( .A(sub_436_3_n65), .ZN(N537) );
  XNOR2_X2 sub_436_3_U104 ( .A(sub_436_3_n134), .B(sub_436_3_carry_85_), .ZN(
        sub_436_3_n65) );
  INV_X4 sub_436_3_U103 ( .A(sub_436_3_n64), .ZN(sub_436_3_carry_86_) );
  NAND2_X2 sub_436_3_U102 ( .A1(sub_436_3_n134), .A2(sub_436_3_carry_85_), 
        .ZN(sub_436_3_n64) );
  INV_X4 sub_436_3_U101 ( .A(sub_436_3_n63), .ZN(N538) );
  XNOR2_X2 sub_436_3_U100 ( .A(sub_436_3_n133), .B(sub_436_3_carry_86_), .ZN(
        sub_436_3_n63) );
  INV_X4 sub_436_3_U99 ( .A(sub_436_3_n62), .ZN(sub_436_3_carry_87_) );
  NAND2_X2 sub_436_3_U98 ( .A1(sub_436_3_n133), .A2(sub_436_3_carry_86_), .ZN(
        sub_436_3_n62) );
  INV_X4 sub_436_3_U97 ( .A(sub_436_3_n61), .ZN(N539) );
  XNOR2_X2 sub_436_3_U96 ( .A(sub_436_3_n132), .B(sub_436_3_carry_87_), .ZN(
        sub_436_3_n61) );
  INV_X4 sub_436_3_U95 ( .A(sub_436_3_n60), .ZN(sub_436_3_carry_88_) );
  NAND2_X2 sub_436_3_U94 ( .A1(sub_436_3_n132), .A2(sub_436_3_carry_87_), .ZN(
        sub_436_3_n60) );
  INV_X4 sub_436_3_U93 ( .A(sub_436_3_n59), .ZN(N540) );
  XNOR2_X2 sub_436_3_U92 ( .A(sub_436_3_n131), .B(sub_436_3_carry_88_), .ZN(
        sub_436_3_n59) );
  INV_X4 sub_436_3_U91 ( .A(sub_436_3_n58), .ZN(sub_436_3_carry_89_) );
  NAND2_X2 sub_436_3_U90 ( .A1(sub_436_3_n131), .A2(sub_436_3_carry_88_), .ZN(
        sub_436_3_n58) );
  INV_X4 sub_436_3_U89 ( .A(sub_436_3_n57), .ZN(N541) );
  XNOR2_X2 sub_436_3_U88 ( .A(sub_436_3_n130), .B(sub_436_3_carry_89_), .ZN(
        sub_436_3_n57) );
  INV_X4 sub_436_3_U87 ( .A(sub_436_3_n56), .ZN(sub_436_3_carry_90_) );
  NAND2_X2 sub_436_3_U86 ( .A1(sub_436_3_n130), .A2(sub_436_3_carry_89_), .ZN(
        sub_436_3_n56) );
  INV_X4 sub_436_3_U85 ( .A(sub_436_3_n55), .ZN(N542) );
  XNOR2_X2 sub_436_3_U84 ( .A(sub_436_3_n129), .B(sub_436_3_carry_90_), .ZN(
        sub_436_3_n55) );
  INV_X4 sub_436_3_U83 ( .A(sub_436_3_n54), .ZN(sub_436_3_carry_91_) );
  NAND2_X2 sub_436_3_U82 ( .A1(sub_436_3_n129), .A2(sub_436_3_carry_90_), .ZN(
        sub_436_3_n54) );
  INV_X4 sub_436_3_U81 ( .A(sub_436_3_n53), .ZN(N543) );
  XNOR2_X2 sub_436_3_U80 ( .A(sub_436_3_n128), .B(sub_436_3_carry_91_), .ZN(
        sub_436_3_n53) );
  INV_X4 sub_436_3_U79 ( .A(sub_436_3_n52), .ZN(sub_436_3_carry_92_) );
  NAND2_X2 sub_436_3_U78 ( .A1(sub_436_3_n128), .A2(sub_436_3_carry_91_), .ZN(
        sub_436_3_n52) );
  INV_X4 sub_436_3_U77 ( .A(sub_436_3_n51), .ZN(N544) );
  XNOR2_X2 sub_436_3_U76 ( .A(sub_436_3_n127), .B(sub_436_3_carry_92_), .ZN(
        sub_436_3_n51) );
  INV_X4 sub_436_3_U75 ( .A(sub_436_3_n50), .ZN(sub_436_3_carry_93_) );
  NAND2_X2 sub_436_3_U74 ( .A1(sub_436_3_n127), .A2(sub_436_3_carry_92_), .ZN(
        sub_436_3_n50) );
  INV_X4 sub_436_3_U73 ( .A(sub_436_3_n49), .ZN(N545) );
  XNOR2_X2 sub_436_3_U72 ( .A(sub_436_3_n126), .B(sub_436_3_carry_93_), .ZN(
        sub_436_3_n49) );
  INV_X4 sub_436_3_U71 ( .A(sub_436_3_n48), .ZN(sub_436_3_carry_94_) );
  NAND2_X2 sub_436_3_U70 ( .A1(sub_436_3_n126), .A2(sub_436_3_carry_93_), .ZN(
        sub_436_3_n48) );
  INV_X4 sub_436_3_U69 ( .A(sub_436_3_n47), .ZN(N546) );
  XNOR2_X2 sub_436_3_U68 ( .A(sub_436_3_n125), .B(sub_436_3_carry_94_), .ZN(
        sub_436_3_n47) );
  INV_X4 sub_436_3_U67 ( .A(sub_436_3_n46), .ZN(sub_436_3_carry_95_) );
  NAND2_X2 sub_436_3_U66 ( .A1(sub_436_3_n125), .A2(sub_436_3_carry_94_), .ZN(
        sub_436_3_n46) );
  INV_X4 sub_436_3_U65 ( .A(sub_436_3_n45), .ZN(N547) );
  XNOR2_X2 sub_436_3_U64 ( .A(sub_436_3_n124), .B(sub_436_3_carry_95_), .ZN(
        sub_436_3_n45) );
  INV_X4 sub_436_3_U63 ( .A(sub_436_3_n44), .ZN(sub_436_3_carry_96_) );
  NAND2_X2 sub_436_3_U62 ( .A1(sub_436_3_n124), .A2(sub_436_3_carry_95_), .ZN(
        sub_436_3_n44) );
  INV_X4 sub_436_3_U61 ( .A(sub_436_3_n43), .ZN(N548) );
  XNOR2_X2 sub_436_3_U60 ( .A(sub_436_3_n123), .B(sub_436_3_carry_96_), .ZN(
        sub_436_3_n43) );
  INV_X4 sub_436_3_U59 ( .A(sub_436_3_n42), .ZN(sub_436_3_carry_97_) );
  NAND2_X2 sub_436_3_U58 ( .A1(sub_436_3_n123), .A2(sub_436_3_carry_96_), .ZN(
        sub_436_3_n42) );
  INV_X4 sub_436_3_U57 ( .A(sub_436_3_n41), .ZN(N549) );
  XNOR2_X2 sub_436_3_U56 ( .A(sub_436_3_n122), .B(sub_436_3_carry_97_), .ZN(
        sub_436_3_n41) );
  INV_X4 sub_436_3_U55 ( .A(sub_436_3_n40), .ZN(sub_436_3_carry_98_) );
  NAND2_X2 sub_436_3_U54 ( .A1(sub_436_3_n122), .A2(sub_436_3_carry_97_), .ZN(
        sub_436_3_n40) );
  INV_X4 sub_436_3_U53 ( .A(sub_436_3_n39), .ZN(N550) );
  XNOR2_X2 sub_436_3_U52 ( .A(sub_436_3_n121), .B(sub_436_3_carry_98_), .ZN(
        sub_436_3_n39) );
  INV_X4 sub_436_3_U51 ( .A(sub_436_3_n38), .ZN(sub_436_3_carry_99_) );
  NAND2_X2 sub_436_3_U50 ( .A1(sub_436_3_n121), .A2(sub_436_3_carry_98_), .ZN(
        sub_436_3_n38) );
  INV_X4 sub_436_3_U49 ( .A(sub_436_3_n37), .ZN(N551) );
  XNOR2_X2 sub_436_3_U48 ( .A(sub_436_3_n120), .B(sub_436_3_carry_99_), .ZN(
        sub_436_3_n37) );
  INV_X4 sub_436_3_U47 ( .A(sub_436_3_n36), .ZN(sub_436_3_carry_100_) );
  NAND2_X2 sub_436_3_U46 ( .A1(sub_436_3_n120), .A2(sub_436_3_carry_99_), .ZN(
        sub_436_3_n36) );
  INV_X4 sub_436_3_U45 ( .A(sub_436_3_n35), .ZN(N552) );
  XNOR2_X2 sub_436_3_U44 ( .A(sub_436_3_n119), .B(sub_436_3_carry_100_), .ZN(
        sub_436_3_n35) );
  INV_X4 sub_436_3_U43 ( .A(sub_436_3_n34), .ZN(sub_436_3_carry_101_) );
  NAND2_X2 sub_436_3_U42 ( .A1(sub_436_3_n119), .A2(sub_436_3_carry_100_), 
        .ZN(sub_436_3_n34) );
  INV_X4 sub_436_3_U41 ( .A(sub_436_3_n33), .ZN(N553) );
  XNOR2_X2 sub_436_3_U40 ( .A(sub_436_3_n118), .B(sub_436_3_carry_101_), .ZN(
        sub_436_3_n33) );
  INV_X4 sub_436_3_U39 ( .A(sub_436_3_n32), .ZN(sub_436_3_carry_102_) );
  NAND2_X2 sub_436_3_U38 ( .A1(sub_436_3_n118), .A2(sub_436_3_carry_101_), 
        .ZN(sub_436_3_n32) );
  INV_X4 sub_436_3_U37 ( .A(sub_436_3_n31), .ZN(N554) );
  XNOR2_X2 sub_436_3_U36 ( .A(sub_436_3_n117), .B(sub_436_3_carry_102_), .ZN(
        sub_436_3_n31) );
  INV_X4 sub_436_3_U35 ( .A(sub_436_3_n30), .ZN(sub_436_3_carry_103_) );
  NAND2_X2 sub_436_3_U34 ( .A1(sub_436_3_n117), .A2(sub_436_3_carry_102_), 
        .ZN(sub_436_3_n30) );
  INV_X4 sub_436_3_U33 ( .A(sub_436_3_n29), .ZN(N555) );
  XNOR2_X2 sub_436_3_U32 ( .A(sub_436_3_n116), .B(sub_436_3_carry_103_), .ZN(
        sub_436_3_n29) );
  INV_X4 sub_436_3_U31 ( .A(sub_436_3_n28), .ZN(sub_436_3_carry_104_) );
  NAND2_X2 sub_436_3_U30 ( .A1(sub_436_3_n116), .A2(sub_436_3_carry_103_), 
        .ZN(sub_436_3_n28) );
  INV_X4 sub_436_3_U29 ( .A(sub_436_3_n27), .ZN(N556) );
  XNOR2_X2 sub_436_3_U28 ( .A(sub_436_3_n115), .B(sub_436_3_carry_104_), .ZN(
        sub_436_3_n27) );
  INV_X4 sub_436_3_U27 ( .A(sub_436_3_n26), .ZN(sub_436_3_carry_105_) );
  NAND2_X2 sub_436_3_U26 ( .A1(sub_436_3_n115), .A2(sub_436_3_carry_104_), 
        .ZN(sub_436_3_n26) );
  XOR2_X1 sub_436_3_U25 ( .A(sub_436_3_n147), .B(sub_436_3_carry_72_), .Z(N524) );
  XOR2_X1 sub_436_3_U24 ( .A(sub_436_3_n148), .B(sub_436_3_carry_71_), .Z(N523) );
  XOR2_X1 sub_436_3_U23 ( .A(sub_436_3_n149), .B(sub_436_3_carry_70_), .Z(N522) );
  XOR2_X1 sub_436_3_U22 ( .A(sub_436_3_n150), .B(sub_436_3_carry_69_), .Z(N521) );
  XOR2_X1 sub_436_3_U21 ( .A(sub_436_3_n151), .B(sub_436_3_carry_68_), .Z(N520) );
  XOR2_X1 sub_436_3_U20 ( .A(sub_436_3_n152), .B(sub_436_3_carry_67_), .Z(N519) );
  XOR2_X1 sub_436_3_U19 ( .A(sub_436_3_n153), .B(sub_436_3_carry_66_), .Z(N518) );
  XOR2_X1 sub_436_3_U18 ( .A(sub_436_3_n154), .B(sub_436_3_carry_65_), .Z(N517) );
  XOR2_X1 sub_436_3_U17 ( .A(sub_436_3_n155), .B(sub_436_3_carry_64_), .Z(N516) );
  XOR2_X1 sub_436_3_U16 ( .A(sub_436_3_n156), .B(sub_436_3_carry_63_), .Z(N515) );
  XOR2_X1 sub_436_3_U15 ( .A(sub_436_3_n157), .B(sub_436_3_carry_62_), .Z(N514) );
  XOR2_X1 sub_436_3_U14 ( .A(sub_436_3_n158), .B(sub_436_3_carry_61_), .Z(N513) );
  XOR2_X1 sub_436_3_U13 ( .A(sub_436_3_n159), .B(sub_436_3_carry_60_), .Z(N512) );
  XOR2_X1 sub_436_3_U12 ( .A(sub_436_3_n160), .B(sub_436_3_carry_59_), .Z(N511) );
  XOR2_X1 sub_436_3_U11 ( .A(sub_436_3_n161), .B(sub_436_3_carry_58_), .Z(N510) );
  XOR2_X1 sub_436_3_U10 ( .A(sub_436_3_n162), .B(sub_436_3_carry_57_), .Z(N509) );
  XOR2_X1 sub_436_3_U9 ( .A(sub_436_3_n163), .B(sub_436_3_carry_56_), .Z(N508)
         );
  XOR2_X1 sub_436_3_U8 ( .A(sub_436_3_n164), .B(sub_436_3_carry_55_), .Z(N507)
         );
  XOR2_X1 sub_436_3_U7 ( .A(sub_436_3_n165), .B(sub_436_3_carry_54_), .Z(N506)
         );
  XOR2_X1 sub_436_3_U6 ( .A(sub_436_3_n166), .B(sub_436_3_carry_53_), .Z(N505)
         );
  XOR2_X1 sub_436_3_U5 ( .A(sub_436_3_n167), .B(sub_436_3_carry_52_), .Z(N504)
         );
  XOR2_X1 sub_436_3_U4 ( .A(sub_436_3_n168), .B(sub_436_3_carry_51_), .Z(N503)
         );
  XOR2_X1 sub_436_3_U3 ( .A(sub_436_3_n169), .B(sub_436_3_carry_50_), .Z(N502)
         );
  XOR2_X1 sub_436_3_U2 ( .A(sub_436_3_n170), .B(sub_436_3_n171), .Z(N501) );
  XOR2_X1 sub_436_3_U1 ( .A(sub_436_3_n114), .B(sub_436_3_carry_105_), .Z(N557) );
  INV_X4 sub_436_b0_U231 ( .A(N343), .ZN(sub_436_b0_n157) );
  INV_X4 sub_436_b0_U230 ( .A(opa_r1[1]), .ZN(sub_436_b0_n156) );
  INV_X4 sub_436_b0_U229 ( .A(opa_r1[2]), .ZN(sub_436_b0_n155) );
  INV_X4 sub_436_b0_U228 ( .A(opa_r1[3]), .ZN(sub_436_b0_n154) );
  INV_X4 sub_436_b0_U227 ( .A(opa_r1[4]), .ZN(sub_436_b0_n153) );
  INV_X4 sub_436_b0_U226 ( .A(opa_r1[5]), .ZN(sub_436_b0_n152) );
  INV_X4 sub_436_b0_U225 ( .A(opa_r1[6]), .ZN(sub_436_b0_n151) );
  INV_X4 sub_436_b0_U224 ( .A(opa_r1[7]), .ZN(sub_436_b0_n150) );
  INV_X4 sub_436_b0_U223 ( .A(opa_r1[8]), .ZN(sub_436_b0_n149) );
  INV_X4 sub_436_b0_U222 ( .A(opa_r1[9]), .ZN(sub_436_b0_n148) );
  INV_X4 sub_436_b0_U221 ( .A(opa_r1[10]), .ZN(sub_436_b0_n147) );
  INV_X4 sub_436_b0_U220 ( .A(opa_r1[11]), .ZN(sub_436_b0_n146) );
  INV_X4 sub_436_b0_U219 ( .A(opa_r1[12]), .ZN(sub_436_b0_n145) );
  INV_X4 sub_436_b0_U218 ( .A(opa_r1[13]), .ZN(sub_436_b0_n144) );
  INV_X4 sub_436_b0_U217 ( .A(opa_r1[14]), .ZN(sub_436_b0_n143) );
  INV_X4 sub_436_b0_U216 ( .A(opa_r1[15]), .ZN(sub_436_b0_n142) );
  INV_X4 sub_436_b0_U215 ( .A(opa_r1[16]), .ZN(sub_436_b0_n141) );
  INV_X4 sub_436_b0_U214 ( .A(opa_r1[17]), .ZN(sub_436_b0_n140) );
  INV_X4 sub_436_b0_U213 ( .A(opa_r1[18]), .ZN(sub_436_b0_n139) );
  INV_X4 sub_436_b0_U212 ( .A(opa_r1[19]), .ZN(sub_436_b0_n138) );
  INV_X4 sub_436_b0_U211 ( .A(opa_r1[20]), .ZN(sub_436_b0_n137) );
  INV_X4 sub_436_b0_U210 ( .A(opa_r1[21]), .ZN(sub_436_b0_n136) );
  INV_X4 sub_436_b0_U209 ( .A(opa_r1[22]), .ZN(sub_436_b0_n135) );
  INV_X4 sub_436_b0_U208 ( .A(opa_r1[23]), .ZN(sub_436_b0_n134) );
  INV_X4 sub_436_b0_U207 ( .A(opa_r1[24]), .ZN(sub_436_b0_n133) );
  INV_X4 sub_436_b0_U206 ( .A(opa_r1[25]), .ZN(sub_436_b0_n132) );
  INV_X4 sub_436_b0_U205 ( .A(opa_r1[26]), .ZN(sub_436_b0_n131) );
  INV_X4 sub_436_b0_U204 ( .A(opa_r1[27]), .ZN(sub_436_b0_n130) );
  INV_X4 sub_436_b0_U203 ( .A(opa_r1[28]), .ZN(sub_436_b0_n129) );
  INV_X4 sub_436_b0_U202 ( .A(opa_r1[29]), .ZN(sub_436_b0_n128) );
  INV_X4 sub_436_b0_U201 ( .A(opa_r1[30]), .ZN(sub_436_b0_n127) );
  INV_X4 sub_436_b0_U200 ( .A(opa_r1[31]), .ZN(sub_436_b0_n126) );
  INV_X4 sub_436_b0_U199 ( .A(opa_r1[32]), .ZN(sub_436_b0_n125) );
  INV_X4 sub_436_b0_U198 ( .A(opa_r1[33]), .ZN(sub_436_b0_n124) );
  INV_X4 sub_436_b0_U197 ( .A(opa_r1[34]), .ZN(sub_436_b0_n123) );
  INV_X4 sub_436_b0_U196 ( .A(opa_r1[35]), .ZN(sub_436_b0_n122) );
  INV_X4 sub_436_b0_U195 ( .A(opa_r1[36]), .ZN(sub_436_b0_n121) );
  INV_X4 sub_436_b0_U194 ( .A(opa_r1[37]), .ZN(sub_436_b0_n120) );
  INV_X4 sub_436_b0_U193 ( .A(opa_r1[38]), .ZN(sub_436_b0_n119) );
  INV_X4 sub_436_b0_U192 ( .A(opa_r1[39]), .ZN(sub_436_b0_n118) );
  INV_X4 sub_436_b0_U191 ( .A(opa_r1[40]), .ZN(sub_436_b0_n117) );
  INV_X4 sub_436_b0_U190 ( .A(opa_r1[41]), .ZN(sub_436_b0_n116) );
  INV_X4 sub_436_b0_U189 ( .A(opa_r1[42]), .ZN(sub_436_b0_n115) );
  INV_X4 sub_436_b0_U188 ( .A(opa_r1[43]), .ZN(sub_436_b0_n114) );
  INV_X4 sub_436_b0_U187 ( .A(opa_r1[44]), .ZN(sub_436_b0_n113) );
  INV_X4 sub_436_b0_U186 ( .A(opa_r1[45]), .ZN(sub_436_b0_n112) );
  INV_X4 sub_436_b0_U185 ( .A(opa_r1[46]), .ZN(sub_436_b0_n111) );
  INV_X4 sub_436_b0_U184 ( .A(opa_r1[47]), .ZN(sub_436_b0_n110) );
  INV_X4 sub_436_b0_U183 ( .A(opa_r1[48]), .ZN(sub_436_b0_n109) );
  INV_X4 sub_436_b0_U182 ( .A(opa_r1[49]), .ZN(sub_436_b0_n108) );
  INV_X4 sub_436_b0_U181 ( .A(opa_r1[50]), .ZN(sub_436_b0_n107) );
  INV_X4 sub_436_b0_U180 ( .A(opa_r1[51]), .ZN(sub_436_b0_n106) );
  INV_X4 sub_436_b0_U179 ( .A(N340), .ZN(sub_436_b0_n105) );
  INV_X4 sub_436_b0_U178 ( .A(sub_436_b0_n104), .ZN(sub_436_b0_carry_2_) );
  NAND2_X2 sub_436_b0_U177 ( .A1(sub_436_b0_n156), .A2(sub_436_b0_n157), .ZN(
        sub_436_b0_n104) );
  INV_X4 sub_436_b0_U176 ( .A(sub_436_b0_n103), .ZN(sub_436_b0_carry_3_) );
  NAND2_X2 sub_436_b0_U175 ( .A1(sub_436_b0_n155), .A2(sub_436_b0_carry_2_), 
        .ZN(sub_436_b0_n103) );
  INV_X4 sub_436_b0_U174 ( .A(sub_436_b0_n102), .ZN(sub_436_b0_carry_4_) );
  NAND2_X2 sub_436_b0_U173 ( .A1(sub_436_b0_n154), .A2(sub_436_b0_carry_3_), 
        .ZN(sub_436_b0_n102) );
  INV_X4 sub_436_b0_U172 ( .A(sub_436_b0_n101), .ZN(sub_436_b0_carry_5_) );
  NAND2_X2 sub_436_b0_U171 ( .A1(sub_436_b0_n153), .A2(sub_436_b0_carry_4_), 
        .ZN(sub_436_b0_n101) );
  INV_X4 sub_436_b0_U170 ( .A(sub_436_b0_n100), .ZN(sub_436_b0_carry_6_) );
  NAND2_X2 sub_436_b0_U169 ( .A1(sub_436_b0_n152), .A2(sub_436_b0_carry_5_), 
        .ZN(sub_436_b0_n100) );
  INV_X4 sub_436_b0_U168 ( .A(sub_436_b0_n99), .ZN(sub_436_b0_carry_7_) );
  NAND2_X2 sub_436_b0_U167 ( .A1(sub_436_b0_n151), .A2(sub_436_b0_carry_6_), 
        .ZN(sub_436_b0_n99) );
  INV_X4 sub_436_b0_U166 ( .A(sub_436_b0_n98), .ZN(sub_436_b0_carry_8_) );
  NAND2_X2 sub_436_b0_U165 ( .A1(sub_436_b0_n150), .A2(sub_436_b0_carry_7_), 
        .ZN(sub_436_b0_n98) );
  INV_X4 sub_436_b0_U164 ( .A(sub_436_b0_n97), .ZN(sub_436_b0_carry_9_) );
  NAND2_X2 sub_436_b0_U163 ( .A1(sub_436_b0_n149), .A2(sub_436_b0_carry_8_), 
        .ZN(sub_436_b0_n97) );
  INV_X4 sub_436_b0_U162 ( .A(sub_436_b0_n96), .ZN(sub_436_b0_carry_10_) );
  NAND2_X2 sub_436_b0_U161 ( .A1(sub_436_b0_n148), .A2(sub_436_b0_carry_9_), 
        .ZN(sub_436_b0_n96) );
  INV_X4 sub_436_b0_U160 ( .A(sub_436_b0_n95), .ZN(sub_436_b0_carry_11_) );
  NAND2_X2 sub_436_b0_U159 ( .A1(sub_436_b0_n147), .A2(sub_436_b0_carry_10_), 
        .ZN(sub_436_b0_n95) );
  INV_X4 sub_436_b0_U158 ( .A(sub_436_b0_n94), .ZN(sub_436_b0_carry_12_) );
  NAND2_X2 sub_436_b0_U157 ( .A1(sub_436_b0_n146), .A2(sub_436_b0_carry_11_), 
        .ZN(sub_436_b0_n94) );
  INV_X4 sub_436_b0_U156 ( .A(sub_436_b0_n93), .ZN(sub_436_b0_carry_13_) );
  NAND2_X2 sub_436_b0_U155 ( .A1(sub_436_b0_n145), .A2(sub_436_b0_carry_12_), 
        .ZN(sub_436_b0_n93) );
  INV_X4 sub_436_b0_U154 ( .A(sub_436_b0_n92), .ZN(sub_436_b0_carry_14_) );
  NAND2_X2 sub_436_b0_U153 ( .A1(sub_436_b0_n144), .A2(sub_436_b0_carry_13_), 
        .ZN(sub_436_b0_n92) );
  INV_X4 sub_436_b0_U152 ( .A(sub_436_b0_n91), .ZN(sub_436_b0_carry_15_) );
  NAND2_X2 sub_436_b0_U151 ( .A1(sub_436_b0_n143), .A2(sub_436_b0_carry_14_), 
        .ZN(sub_436_b0_n91) );
  INV_X4 sub_436_b0_U150 ( .A(sub_436_b0_n90), .ZN(sub_436_b0_carry_16_) );
  NAND2_X2 sub_436_b0_U149 ( .A1(sub_436_b0_n142), .A2(sub_436_b0_carry_15_), 
        .ZN(sub_436_b0_n90) );
  INV_X4 sub_436_b0_U148 ( .A(sub_436_b0_n89), .ZN(sub_436_b0_carry_17_) );
  NAND2_X2 sub_436_b0_U147 ( .A1(sub_436_b0_n141), .A2(sub_436_b0_carry_16_), 
        .ZN(sub_436_b0_n89) );
  INV_X4 sub_436_b0_U146 ( .A(sub_436_b0_n88), .ZN(sub_436_b0_carry_18_) );
  NAND2_X2 sub_436_b0_U145 ( .A1(sub_436_b0_n140), .A2(sub_436_b0_carry_17_), 
        .ZN(sub_436_b0_n88) );
  INV_X4 sub_436_b0_U144 ( .A(sub_436_b0_n87), .ZN(sub_436_b0_carry_19_) );
  NAND2_X2 sub_436_b0_U143 ( .A1(sub_436_b0_n139), .A2(sub_436_b0_carry_18_), 
        .ZN(sub_436_b0_n87) );
  INV_X4 sub_436_b0_U142 ( .A(sub_436_b0_n86), .ZN(sub_436_b0_carry_20_) );
  NAND2_X2 sub_436_b0_U141 ( .A1(sub_436_b0_n138), .A2(sub_436_b0_carry_19_), 
        .ZN(sub_436_b0_n86) );
  INV_X4 sub_436_b0_U140 ( .A(sub_436_b0_n85), .ZN(sub_436_b0_carry_21_) );
  NAND2_X2 sub_436_b0_U139 ( .A1(sub_436_b0_n137), .A2(sub_436_b0_carry_20_), 
        .ZN(sub_436_b0_n85) );
  INV_X4 sub_436_b0_U138 ( .A(sub_436_b0_n84), .ZN(sub_436_b0_carry_22_) );
  NAND2_X2 sub_436_b0_U137 ( .A1(sub_436_b0_n136), .A2(sub_436_b0_carry_21_), 
        .ZN(sub_436_b0_n84) );
  INV_X4 sub_436_b0_U136 ( .A(sub_436_b0_n83), .ZN(sub_436_b0_carry_23_) );
  NAND2_X2 sub_436_b0_U135 ( .A1(sub_436_b0_n135), .A2(sub_436_b0_carry_22_), 
        .ZN(sub_436_b0_n83) );
  INV_X4 sub_436_b0_U134 ( .A(sub_436_b0_n82), .ZN(sub_436_b0_carry_24_) );
  NAND2_X2 sub_436_b0_U133 ( .A1(sub_436_b0_n134), .A2(sub_436_b0_carry_23_), 
        .ZN(sub_436_b0_n82) );
  INV_X4 sub_436_b0_U132 ( .A(sub_436_b0_n81), .ZN(sub_436_b0_carry_25_) );
  NAND2_X2 sub_436_b0_U131 ( .A1(sub_436_b0_n133), .A2(sub_436_b0_carry_24_), 
        .ZN(sub_436_b0_n81) );
  INV_X4 sub_436_b0_U130 ( .A(sub_436_b0_n80), .ZN(N368) );
  XNOR2_X2 sub_436_b0_U129 ( .A(sub_436_b0_n132), .B(sub_436_b0_carry_25_), 
        .ZN(sub_436_b0_n80) );
  INV_X4 sub_436_b0_U128 ( .A(sub_436_b0_n79), .ZN(sub_436_b0_carry_26_) );
  NAND2_X2 sub_436_b0_U127 ( .A1(sub_436_b0_n132), .A2(sub_436_b0_carry_25_), 
        .ZN(sub_436_b0_n79) );
  INV_X4 sub_436_b0_U126 ( .A(sub_436_b0_n78), .ZN(N369) );
  XNOR2_X2 sub_436_b0_U125 ( .A(sub_436_b0_n131), .B(sub_436_b0_carry_26_), 
        .ZN(sub_436_b0_n78) );
  INV_X4 sub_436_b0_U124 ( .A(sub_436_b0_n77), .ZN(sub_436_b0_carry_27_) );
  NAND2_X2 sub_436_b0_U123 ( .A1(sub_436_b0_n131), .A2(sub_436_b0_carry_26_), 
        .ZN(sub_436_b0_n77) );
  INV_X4 sub_436_b0_U122 ( .A(sub_436_b0_n76), .ZN(N370) );
  XNOR2_X2 sub_436_b0_U121 ( .A(sub_436_b0_n130), .B(sub_436_b0_carry_27_), 
        .ZN(sub_436_b0_n76) );
  INV_X4 sub_436_b0_U120 ( .A(sub_436_b0_n75), .ZN(sub_436_b0_carry_28_) );
  NAND2_X2 sub_436_b0_U119 ( .A1(sub_436_b0_n130), .A2(sub_436_b0_carry_27_), 
        .ZN(sub_436_b0_n75) );
  INV_X4 sub_436_b0_U118 ( .A(sub_436_b0_n74), .ZN(N371) );
  XNOR2_X2 sub_436_b0_U117 ( .A(sub_436_b0_n129), .B(sub_436_b0_carry_28_), 
        .ZN(sub_436_b0_n74) );
  INV_X4 sub_436_b0_U116 ( .A(sub_436_b0_n73), .ZN(sub_436_b0_carry_29_) );
  NAND2_X2 sub_436_b0_U115 ( .A1(sub_436_b0_n129), .A2(sub_436_b0_carry_28_), 
        .ZN(sub_436_b0_n73) );
  INV_X4 sub_436_b0_U114 ( .A(sub_436_b0_n72), .ZN(N372) );
  XNOR2_X2 sub_436_b0_U113 ( .A(sub_436_b0_n128), .B(sub_436_b0_carry_29_), 
        .ZN(sub_436_b0_n72) );
  INV_X4 sub_436_b0_U112 ( .A(sub_436_b0_n71), .ZN(sub_436_b0_carry_30_) );
  NAND2_X2 sub_436_b0_U111 ( .A1(sub_436_b0_n128), .A2(sub_436_b0_carry_29_), 
        .ZN(sub_436_b0_n71) );
  INV_X4 sub_436_b0_U110 ( .A(sub_436_b0_n70), .ZN(N373) );
  XNOR2_X2 sub_436_b0_U109 ( .A(sub_436_b0_n127), .B(sub_436_b0_carry_30_), 
        .ZN(sub_436_b0_n70) );
  INV_X4 sub_436_b0_U108 ( .A(sub_436_b0_n69), .ZN(sub_436_b0_carry_31_) );
  NAND2_X2 sub_436_b0_U107 ( .A1(sub_436_b0_n127), .A2(sub_436_b0_carry_30_), 
        .ZN(sub_436_b0_n69) );
  INV_X4 sub_436_b0_U106 ( .A(sub_436_b0_n68), .ZN(N374) );
  XNOR2_X2 sub_436_b0_U105 ( .A(sub_436_b0_n126), .B(sub_436_b0_carry_31_), 
        .ZN(sub_436_b0_n68) );
  INV_X4 sub_436_b0_U104 ( .A(sub_436_b0_n67), .ZN(sub_436_b0_carry_32_) );
  NAND2_X2 sub_436_b0_U103 ( .A1(sub_436_b0_n126), .A2(sub_436_b0_carry_31_), 
        .ZN(sub_436_b0_n67) );
  INV_X4 sub_436_b0_U102 ( .A(sub_436_b0_n66), .ZN(N375) );
  XNOR2_X2 sub_436_b0_U101 ( .A(sub_436_b0_n125), .B(sub_436_b0_carry_32_), 
        .ZN(sub_436_b0_n66) );
  INV_X4 sub_436_b0_U100 ( .A(sub_436_b0_n65), .ZN(sub_436_b0_carry_33_) );
  NAND2_X2 sub_436_b0_U99 ( .A1(sub_436_b0_n125), .A2(sub_436_b0_carry_32_), 
        .ZN(sub_436_b0_n65) );
  INV_X4 sub_436_b0_U98 ( .A(sub_436_b0_n64), .ZN(N376) );
  XNOR2_X2 sub_436_b0_U97 ( .A(sub_436_b0_n124), .B(sub_436_b0_carry_33_), 
        .ZN(sub_436_b0_n64) );
  INV_X4 sub_436_b0_U96 ( .A(sub_436_b0_n63), .ZN(sub_436_b0_carry_34_) );
  NAND2_X2 sub_436_b0_U95 ( .A1(sub_436_b0_n124), .A2(sub_436_b0_carry_33_), 
        .ZN(sub_436_b0_n63) );
  INV_X4 sub_436_b0_U94 ( .A(sub_436_b0_n62), .ZN(N377) );
  XNOR2_X2 sub_436_b0_U93 ( .A(sub_436_b0_n123), .B(sub_436_b0_carry_34_), 
        .ZN(sub_436_b0_n62) );
  INV_X4 sub_436_b0_U92 ( .A(sub_436_b0_n61), .ZN(sub_436_b0_carry_35_) );
  NAND2_X2 sub_436_b0_U91 ( .A1(sub_436_b0_n123), .A2(sub_436_b0_carry_34_), 
        .ZN(sub_436_b0_n61) );
  INV_X4 sub_436_b0_U90 ( .A(sub_436_b0_n60), .ZN(N378) );
  XNOR2_X2 sub_436_b0_U89 ( .A(sub_436_b0_n122), .B(sub_436_b0_carry_35_), 
        .ZN(sub_436_b0_n60) );
  INV_X4 sub_436_b0_U88 ( .A(sub_436_b0_n59), .ZN(sub_436_b0_carry_36_) );
  NAND2_X2 sub_436_b0_U87 ( .A1(sub_436_b0_n122), .A2(sub_436_b0_carry_35_), 
        .ZN(sub_436_b0_n59) );
  INV_X4 sub_436_b0_U86 ( .A(sub_436_b0_n58), .ZN(N379) );
  XNOR2_X2 sub_436_b0_U85 ( .A(sub_436_b0_n121), .B(sub_436_b0_carry_36_), 
        .ZN(sub_436_b0_n58) );
  INV_X4 sub_436_b0_U84 ( .A(sub_436_b0_n57), .ZN(sub_436_b0_carry_37_) );
  NAND2_X2 sub_436_b0_U83 ( .A1(sub_436_b0_n121), .A2(sub_436_b0_carry_36_), 
        .ZN(sub_436_b0_n57) );
  INV_X4 sub_436_b0_U82 ( .A(sub_436_b0_n56), .ZN(N380) );
  XNOR2_X2 sub_436_b0_U81 ( .A(sub_436_b0_n120), .B(sub_436_b0_carry_37_), 
        .ZN(sub_436_b0_n56) );
  INV_X4 sub_436_b0_U80 ( .A(sub_436_b0_n55), .ZN(sub_436_b0_carry_38_) );
  NAND2_X2 sub_436_b0_U79 ( .A1(sub_436_b0_n120), .A2(sub_436_b0_carry_37_), 
        .ZN(sub_436_b0_n55) );
  INV_X4 sub_436_b0_U78 ( .A(sub_436_b0_n54), .ZN(N381) );
  XNOR2_X2 sub_436_b0_U77 ( .A(sub_436_b0_n119), .B(sub_436_b0_carry_38_), 
        .ZN(sub_436_b0_n54) );
  INV_X4 sub_436_b0_U76 ( .A(sub_436_b0_n53), .ZN(sub_436_b0_carry_39_) );
  NAND2_X2 sub_436_b0_U75 ( .A1(sub_436_b0_n119), .A2(sub_436_b0_carry_38_), 
        .ZN(sub_436_b0_n53) );
  INV_X4 sub_436_b0_U74 ( .A(sub_436_b0_n52), .ZN(N382) );
  XNOR2_X2 sub_436_b0_U73 ( .A(sub_436_b0_n118), .B(sub_436_b0_carry_39_), 
        .ZN(sub_436_b0_n52) );
  INV_X4 sub_436_b0_U72 ( .A(sub_436_b0_n51), .ZN(sub_436_b0_carry_40_) );
  NAND2_X2 sub_436_b0_U71 ( .A1(sub_436_b0_n118), .A2(sub_436_b0_carry_39_), 
        .ZN(sub_436_b0_n51) );
  INV_X4 sub_436_b0_U70 ( .A(sub_436_b0_n50), .ZN(N383) );
  XNOR2_X2 sub_436_b0_U69 ( .A(sub_436_b0_n117), .B(sub_436_b0_carry_40_), 
        .ZN(sub_436_b0_n50) );
  INV_X4 sub_436_b0_U68 ( .A(sub_436_b0_n49), .ZN(sub_436_b0_carry_41_) );
  NAND2_X2 sub_436_b0_U67 ( .A1(sub_436_b0_n117), .A2(sub_436_b0_carry_40_), 
        .ZN(sub_436_b0_n49) );
  INV_X4 sub_436_b0_U66 ( .A(sub_436_b0_n48), .ZN(N384) );
  XNOR2_X2 sub_436_b0_U65 ( .A(sub_436_b0_n116), .B(sub_436_b0_carry_41_), 
        .ZN(sub_436_b0_n48) );
  INV_X4 sub_436_b0_U64 ( .A(sub_436_b0_n47), .ZN(sub_436_b0_carry_42_) );
  NAND2_X2 sub_436_b0_U63 ( .A1(sub_436_b0_n116), .A2(sub_436_b0_carry_41_), 
        .ZN(sub_436_b0_n47) );
  INV_X4 sub_436_b0_U62 ( .A(sub_436_b0_n46), .ZN(N385) );
  XNOR2_X2 sub_436_b0_U61 ( .A(sub_436_b0_n115), .B(sub_436_b0_carry_42_), 
        .ZN(sub_436_b0_n46) );
  INV_X4 sub_436_b0_U60 ( .A(sub_436_b0_n45), .ZN(sub_436_b0_carry_43_) );
  NAND2_X2 sub_436_b0_U59 ( .A1(sub_436_b0_n115), .A2(sub_436_b0_carry_42_), 
        .ZN(sub_436_b0_n45) );
  INV_X4 sub_436_b0_U58 ( .A(sub_436_b0_n44), .ZN(N386) );
  XNOR2_X2 sub_436_b0_U57 ( .A(sub_436_b0_n114), .B(sub_436_b0_carry_43_), 
        .ZN(sub_436_b0_n44) );
  INV_X4 sub_436_b0_U56 ( .A(sub_436_b0_n43), .ZN(sub_436_b0_carry_44_) );
  NAND2_X2 sub_436_b0_U55 ( .A1(sub_436_b0_n114), .A2(sub_436_b0_carry_43_), 
        .ZN(sub_436_b0_n43) );
  INV_X4 sub_436_b0_U54 ( .A(sub_436_b0_n42), .ZN(N387) );
  XNOR2_X2 sub_436_b0_U53 ( .A(sub_436_b0_n113), .B(sub_436_b0_carry_44_), 
        .ZN(sub_436_b0_n42) );
  INV_X4 sub_436_b0_U52 ( .A(sub_436_b0_n41), .ZN(sub_436_b0_carry_45_) );
  NAND2_X2 sub_436_b0_U51 ( .A1(sub_436_b0_n113), .A2(sub_436_b0_carry_44_), 
        .ZN(sub_436_b0_n41) );
  INV_X4 sub_436_b0_U50 ( .A(sub_436_b0_n40), .ZN(N388) );
  XNOR2_X2 sub_436_b0_U49 ( .A(sub_436_b0_n112), .B(sub_436_b0_carry_45_), 
        .ZN(sub_436_b0_n40) );
  INV_X4 sub_436_b0_U48 ( .A(sub_436_b0_n39), .ZN(sub_436_b0_carry_46_) );
  NAND2_X2 sub_436_b0_U47 ( .A1(sub_436_b0_n112), .A2(sub_436_b0_carry_45_), 
        .ZN(sub_436_b0_n39) );
  INV_X4 sub_436_b0_U46 ( .A(sub_436_b0_n38), .ZN(N389) );
  XNOR2_X2 sub_436_b0_U45 ( .A(sub_436_b0_n111), .B(sub_436_b0_carry_46_), 
        .ZN(sub_436_b0_n38) );
  INV_X4 sub_436_b0_U44 ( .A(sub_436_b0_n37), .ZN(sub_436_b0_carry_47_) );
  NAND2_X2 sub_436_b0_U43 ( .A1(sub_436_b0_n111), .A2(sub_436_b0_carry_46_), 
        .ZN(sub_436_b0_n37) );
  INV_X4 sub_436_b0_U42 ( .A(sub_436_b0_n36), .ZN(N390) );
  XNOR2_X2 sub_436_b0_U41 ( .A(sub_436_b0_n110), .B(sub_436_b0_carry_47_), 
        .ZN(sub_436_b0_n36) );
  INV_X4 sub_436_b0_U40 ( .A(sub_436_b0_n35), .ZN(sub_436_b0_carry_48_) );
  NAND2_X2 sub_436_b0_U39 ( .A1(sub_436_b0_n110), .A2(sub_436_b0_carry_47_), 
        .ZN(sub_436_b0_n35) );
  INV_X4 sub_436_b0_U38 ( .A(sub_436_b0_n34), .ZN(sub_436_b0_carry_49_) );
  NAND2_X2 sub_436_b0_U37 ( .A1(sub_436_b0_n109), .A2(sub_436_b0_carry_48_), 
        .ZN(sub_436_b0_n34) );
  INV_X4 sub_436_b0_U36 ( .A(sub_436_b0_n33), .ZN(sub_436_b0_carry_50_) );
  NAND2_X2 sub_436_b0_U35 ( .A1(sub_436_b0_n108), .A2(sub_436_b0_carry_49_), 
        .ZN(sub_436_b0_n33) );
  INV_X4 sub_436_b0_U34 ( .A(sub_436_b0_n32), .ZN(sub_436_b0_carry_51_) );
  NAND2_X2 sub_436_b0_U33 ( .A1(sub_436_b0_n107), .A2(sub_436_b0_carry_50_), 
        .ZN(sub_436_b0_n32) );
  INV_X4 sub_436_b0_U32 ( .A(sub_436_b0_n31), .ZN(sub_436_b0_carry_52_) );
  NAND2_X2 sub_436_b0_U31 ( .A1(sub_436_b0_n106), .A2(sub_436_b0_carry_51_), 
        .ZN(sub_436_b0_n31) );
  NAND2_X2 sub_436_b0_U30 ( .A1(sub_436_b0_n105), .A2(sub_436_b0_carry_52_), 
        .ZN(N396) );
  XOR2_X1 sub_436_b0_U29 ( .A(sub_436_b0_n156), .B(sub_436_b0_n157), .Z(N344)
         );
  XOR2_X1 sub_436_b0_U28 ( .A(sub_436_b0_n133), .B(sub_436_b0_carry_24_), .Z(
        N367) );
  XOR2_X1 sub_436_b0_U27 ( .A(sub_436_b0_n134), .B(sub_436_b0_carry_23_), .Z(
        N366) );
  XOR2_X1 sub_436_b0_U26 ( .A(sub_436_b0_n135), .B(sub_436_b0_carry_22_), .Z(
        N365) );
  XOR2_X1 sub_436_b0_U25 ( .A(sub_436_b0_n136), .B(sub_436_b0_carry_21_), .Z(
        N364) );
  XOR2_X1 sub_436_b0_U24 ( .A(sub_436_b0_n137), .B(sub_436_b0_carry_20_), .Z(
        N363) );
  XOR2_X1 sub_436_b0_U23 ( .A(sub_436_b0_n138), .B(sub_436_b0_carry_19_), .Z(
        N362) );
  XOR2_X1 sub_436_b0_U22 ( .A(sub_436_b0_n139), .B(sub_436_b0_carry_18_), .Z(
        N361) );
  XOR2_X1 sub_436_b0_U21 ( .A(sub_436_b0_n140), .B(sub_436_b0_carry_17_), .Z(
        N360) );
  XOR2_X1 sub_436_b0_U20 ( .A(sub_436_b0_n141), .B(sub_436_b0_carry_16_), .Z(
        N359) );
  XOR2_X1 sub_436_b0_U19 ( .A(sub_436_b0_n142), .B(sub_436_b0_carry_15_), .Z(
        N358) );
  XOR2_X1 sub_436_b0_U18 ( .A(sub_436_b0_n143), .B(sub_436_b0_carry_14_), .Z(
        N357) );
  XOR2_X1 sub_436_b0_U17 ( .A(sub_436_b0_n144), .B(sub_436_b0_carry_13_), .Z(
        N356) );
  XOR2_X1 sub_436_b0_U16 ( .A(sub_436_b0_n145), .B(sub_436_b0_carry_12_), .Z(
        N355) );
  XOR2_X1 sub_436_b0_U15 ( .A(sub_436_b0_n146), .B(sub_436_b0_carry_11_), .Z(
        N354) );
  XOR2_X1 sub_436_b0_U14 ( .A(sub_436_b0_n147), .B(sub_436_b0_carry_10_), .Z(
        N353) );
  XOR2_X1 sub_436_b0_U13 ( .A(sub_436_b0_n148), .B(sub_436_b0_carry_9_), .Z(
        N352) );
  XOR2_X1 sub_436_b0_U12 ( .A(sub_436_b0_n149), .B(sub_436_b0_carry_8_), .Z(
        N351) );
  XOR2_X1 sub_436_b0_U11 ( .A(sub_436_b0_n150), .B(sub_436_b0_carry_7_), .Z(
        N350) );
  XOR2_X1 sub_436_b0_U10 ( .A(sub_436_b0_n151), .B(sub_436_b0_carry_6_), .Z(
        N349) );
  XOR2_X1 sub_436_b0_U9 ( .A(sub_436_b0_n152), .B(sub_436_b0_carry_5_), .Z(
        N348) );
  XOR2_X1 sub_436_b0_U8 ( .A(sub_436_b0_n153), .B(sub_436_b0_carry_4_), .Z(
        N347) );
  XOR2_X1 sub_436_b0_U7 ( .A(sub_436_b0_n154), .B(sub_436_b0_carry_3_), .Z(
        N346) );
  XOR2_X1 sub_436_b0_U6 ( .A(sub_436_b0_n155), .B(sub_436_b0_carry_2_), .Z(
        N345) );
  XOR2_X1 sub_436_b0_U5 ( .A(sub_436_b0_n105), .B(sub_436_b0_carry_52_), .Z(
        N395) );
  XOR2_X1 sub_436_b0_U4 ( .A(sub_436_b0_n106), .B(sub_436_b0_carry_51_), .Z(
        N394) );
  XOR2_X1 sub_436_b0_U3 ( .A(sub_436_b0_n107), .B(sub_436_b0_carry_50_), .Z(
        N393) );
  XOR2_X1 sub_436_b0_U2 ( .A(sub_436_b0_n108), .B(sub_436_b0_carry_49_), .Z(
        N392) );
  XOR2_X1 sub_436_b0_U1 ( .A(sub_436_b0_n109), .B(sub_436_b0_carry_48_), .Z(
        N391) );
  AND2_X1 sll_386_U66 ( .A1(fracta_mul[0]), .A2(sll_386_n2), .ZN(
        sll_386_ML_int_1__0_) );
  AND2_X1 sll_386_U65 ( .A1(sll_386_ML_int_1__0_), .A2(sll_386_n8), .ZN(
        sll_386_ML_int_2__0_) );
  AND2_X1 sll_386_U64 ( .A1(sll_386_ML_int_1__1_), .A2(sll_386_n8), .ZN(
        sll_386_ML_int_2__1_) );
  AND2_X1 sll_386_U63 ( .A1(sll_386_ML_int_2__0_), .A2(sll_386_n13), .ZN(
        sll_386_ML_int_3__0_) );
  AND2_X1 sll_386_U62 ( .A1(sll_386_ML_int_2__1_), .A2(sll_386_n13), .ZN(
        sll_386_ML_int_3__1_) );
  AND2_X1 sll_386_U61 ( .A1(sll_386_ML_int_2__2_), .A2(sll_386_n13), .ZN(
        sll_386_ML_int_3__2_) );
  AND2_X1 sll_386_U60 ( .A1(sll_386_ML_int_2__3_), .A2(sll_386_n13), .ZN(
        sll_386_ML_int_3__3_) );
  NAND2_X1 sll_386_U59 ( .A1(sll_386_ML_int_3__0_), .A2(sll_386_n21), .ZN(
        sll_386_n41) );
  NAND2_X1 sll_386_U58 ( .A1(sll_386_ML_int_3__1_), .A2(sll_386_n21), .ZN(
        sll_386_n40) );
  NAND2_X1 sll_386_U57 ( .A1(sll_386_ML_int_3__2_), .A2(sll_386_n21), .ZN(
        sll_386_n39) );
  NAND2_X1 sll_386_U56 ( .A1(sll_386_ML_int_3__3_), .A2(sll_386_n21), .ZN(
        sll_386_n38) );
  NAND2_X1 sll_386_U55 ( .A1(sll_386_ML_int_3__4_), .A2(sll_386_n21), .ZN(
        sll_386_n37) );
  NAND2_X1 sll_386_U54 ( .A1(sll_386_ML_int_3__5_), .A2(sll_386_n21), .ZN(
        sll_386_n36) );
  NAND2_X1 sll_386_U53 ( .A1(sll_386_ML_int_3__6_), .A2(sll_386_n21), .ZN(
        sll_386_n35) );
  NAND2_X1 sll_386_U52 ( .A1(sll_386_ML_int_3__7_), .A2(sll_386_n21), .ZN(
        sll_386_n34) );
  NOR2_X1 sll_386_U51 ( .A1(sll_386_n22), .A2(sll_386_n41), .ZN(N256) );
  AND2_X1 sll_386_U50 ( .A1(sll_386_ML_int_4__10_), .A2(sll_386_n25), .ZN(N266) );
  AND2_X1 sll_386_U49 ( .A1(sll_386_ML_int_4__11_), .A2(sll_386_n25), .ZN(N267) );
  AND2_X1 sll_386_U48 ( .A1(sll_386_ML_int_4__12_), .A2(sll_386_n25), .ZN(N268) );
  AND2_X1 sll_386_U47 ( .A1(sll_386_ML_int_4__13_), .A2(sll_386_n25), .ZN(N269) );
  AND2_X1 sll_386_U46 ( .A1(sll_386_ML_int_4__14_), .A2(sll_386_n25), .ZN(N270) );
  AND2_X1 sll_386_U45 ( .A1(sll_386_ML_int_4__15_), .A2(sll_386_n25), .ZN(N271) );
  NOR2_X1 sll_386_U44 ( .A1(sll_386_n23), .A2(sll_386_n40), .ZN(N257) );
  NOR2_X1 sll_386_U43 ( .A1(sll_386_n24), .A2(sll_386_n39), .ZN(N258) );
  NOR2_X1 sll_386_U42 ( .A1(div_opa_ldz_d[4]), .A2(sll_386_n38), .ZN(N259) );
  NOR2_X1 sll_386_U41 ( .A1(div_opa_ldz_d[4]), .A2(sll_386_n37), .ZN(N260) );
  NOR2_X1 sll_386_U40 ( .A1(div_opa_ldz_d[4]), .A2(sll_386_n36), .ZN(N261) );
  NOR2_X1 sll_386_U39 ( .A1(div_opa_ldz_d[4]), .A2(sll_386_n35), .ZN(N262) );
  NOR2_X1 sll_386_U38 ( .A1(div_opa_ldz_d[4]), .A2(sll_386_n34), .ZN(N263) );
  AND2_X1 sll_386_U37 ( .A1(sll_386_ML_int_4__8_), .A2(sll_386_n25), .ZN(N264)
         );
  AND2_X1 sll_386_U36 ( .A1(sll_386_ML_int_4__9_), .A2(sll_386_n25), .ZN(N265)
         );
  INV_X4 sll_386_U35 ( .A(sll_386_n34), .ZN(sll_386_n33) );
  INV_X4 sll_386_U34 ( .A(sll_386_n35), .ZN(sll_386_n32) );
  INV_X4 sll_386_U33 ( .A(sll_386_n36), .ZN(sll_386_n31) );
  INV_X4 sll_386_U32 ( .A(sll_386_n37), .ZN(sll_386_n30) );
  INV_X4 sll_386_U31 ( .A(sll_386_n41), .ZN(sll_386_n29) );
  INV_X4 sll_386_U30 ( .A(sll_386_n40), .ZN(sll_386_n28) );
  INV_X4 sll_386_U29 ( .A(sll_386_n39), .ZN(sll_386_n27) );
  INV_X4 sll_386_U28 ( .A(sll_386_n38), .ZN(sll_386_n26) );
  INV_X32 sll_386_U27 ( .A(sll_386_n14), .ZN(sll_386_n21) );
  INV_X32 sll_386_U26 ( .A(sll_386_n14), .ZN(sll_386_n20) );
  INV_X32 sll_386_U25 ( .A(sll_386_n20), .ZN(sll_386_n19) );
  INV_X32 sll_386_U24 ( .A(sll_386_n20), .ZN(sll_386_n18) );
  INV_X32 sll_386_U23 ( .A(sll_386_n21), .ZN(sll_386_n17) );
  INV_X32 sll_386_U22 ( .A(sll_386_n21), .ZN(sll_386_n16) );
  INV_X32 sll_386_U21 ( .A(sll_386_n15), .ZN(sll_386_n14) );
  INV_X32 sll_386_U20 ( .A(sll_386_n13), .ZN(sll_386_n12) );
  INV_X16 sll_386_U19 ( .A(div_opa_ldz_d[1]), .ZN(sll_386_n8) );
  INV_X32 sll_386_U18 ( .A(sll_386_n8), .ZN(sll_386_n7) );
  INV_X32 sll_386_U17 ( .A(sll_386_n8), .ZN(sll_386_n6) );
  INV_X32 sll_386_U16 ( .A(sll_386_n8), .ZN(sll_386_n5) );
  INV_X32 sll_386_U15 ( .A(sll_386_n2), .ZN(sll_386_n4) );
  INV_X32 sll_386_U14 ( .A(sll_386_n2), .ZN(sll_386_n3) );
  INV_X32 sll_386_U13 ( .A(sll_386_n2), .ZN(sll_386_n1) );
  INV_X16 sll_386_U12 ( .A(div_opa_ldz_d[0]), .ZN(sll_386_n2) );
  INV_X8 sll_386_U11 ( .A(sll_386_n25), .ZN(sll_386_n22) );
  INV_X8 sll_386_U10 ( .A(sll_386_n25), .ZN(sll_386_n23) );
  INV_X4 sll_386_U9 ( .A(div_opa_ldz_d[4]), .ZN(sll_386_n25) );
  INV_X4 sll_386_U8 ( .A(div_opa_ldz_d[2]), .ZN(sll_386_n13) );
  INV_X4 sll_386_U7 ( .A(sll_386_n13), .ZN(sll_386_n9) );
  INV_X4 sll_386_U6 ( .A(sll_386_n13), .ZN(sll_386_n10) );
  INV_X4 sll_386_U5 ( .A(sll_386_n13), .ZN(sll_386_n11) );
  INV_X4 sll_386_U4 ( .A(div_opa_ldz_d[3]), .ZN(sll_386_n15) );
  INV_X4 sll_386_U3 ( .A(sll_386_n25), .ZN(sll_386_n24) );
  MUX2_X2 sll_386_M1_0_1 ( .A(n4799), .B(fracta_mul[0]), .S(sll_386_n1), .Z(
        sll_386_ML_int_1__1_) );
  MUX2_X2 sll_386_M1_0_2 ( .A(fracta_mul[2]), .B(n4799), .S(sll_386_n1), .Z(
        sll_386_ML_int_1__2_) );
  MUX2_X2 sll_386_M1_0_3 ( .A(n4727), .B(fracta_mul[2]), .S(sll_386_n1), .Z(
        sll_386_ML_int_1__3_) );
  MUX2_X2 sll_386_M1_0_4 ( .A(fracta_mul[4]), .B(n4727), .S(sll_386_n1), .Z(
        sll_386_ML_int_1__4_) );
  MUX2_X2 sll_386_M1_0_5 ( .A(fracta_mul[5]), .B(fracta_mul[4]), .S(sll_386_n1), .Z(sll_386_ML_int_1__5_) );
  MUX2_X2 sll_386_M1_0_6 ( .A(fracta_mul[6]), .B(fracta_mul[5]), .S(sll_386_n1), .Z(sll_386_ML_int_1__6_) );
  MUX2_X2 sll_386_M1_0_7 ( .A(fracta_mul[7]), .B(fracta_mul[6]), .S(sll_386_n1), .Z(sll_386_ML_int_1__7_) );
  MUX2_X2 sll_386_M1_0_8 ( .A(fracta_mul[8]), .B(fracta_mul[7]), .S(sll_386_n1), .Z(sll_386_ML_int_1__8_) );
  MUX2_X2 sll_386_M1_0_9 ( .A(fracta_mul[9]), .B(fracta_mul[8]), .S(sll_386_n1), .Z(sll_386_ML_int_1__9_) );
  MUX2_X2 sll_386_M1_0_10 ( .A(fracta_mul[10]), .B(fracta_mul[9]), .S(
        sll_386_n1), .Z(sll_386_ML_int_1__10_) );
  MUX2_X2 sll_386_M1_0_11 ( .A(fracta_mul[11]), .B(fracta_mul[10]), .S(
        sll_386_n1), .Z(sll_386_ML_int_1__11_) );
  MUX2_X2 sll_386_M1_0_12 ( .A(fracta_mul[12]), .B(fracta_mul[11]), .S(
        sll_386_n1), .Z(sll_386_ML_int_1__12_) );
  MUX2_X2 sll_386_M1_0_13 ( .A(fracta_mul[13]), .B(fracta_mul[12]), .S(
        sll_386_n1), .Z(sll_386_ML_int_1__13_) );
  MUX2_X2 sll_386_M1_0_14 ( .A(fracta_mul[14]), .B(fracta_mul[13]), .S(
        sll_386_n1), .Z(sll_386_ML_int_1__14_) );
  MUX2_X2 sll_386_M1_0_15 ( .A(fracta_mul[15]), .B(fracta_mul[14]), .S(
        sll_386_n1), .Z(sll_386_ML_int_1__15_) );
  MUX2_X2 sll_386_M1_0_16 ( .A(fracta_mul[16]), .B(fracta_mul[15]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__16_) );
  MUX2_X2 sll_386_M1_0_17 ( .A(fracta_mul[17]), .B(fracta_mul[16]), .S(
        sll_386_n1), .Z(sll_386_ML_int_1__17_) );
  MUX2_X2 sll_386_M1_0_18 ( .A(fracta_mul[18]), .B(fracta_mul[17]), .S(
        sll_386_n1), .Z(sll_386_ML_int_1__18_) );
  MUX2_X2 sll_386_M1_0_19 ( .A(fracta_mul[19]), .B(fracta_mul[18]), .S(
        sll_386_n1), .Z(sll_386_ML_int_1__19_) );
  MUX2_X2 sll_386_M1_0_20 ( .A(fracta_mul[20]), .B(fracta_mul[19]), .S(
        sll_386_n1), .Z(sll_386_ML_int_1__20_) );
  MUX2_X2 sll_386_M1_0_21 ( .A(fracta_mul[21]), .B(fracta_mul[20]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__21_) );
  MUX2_X2 sll_386_M1_0_22 ( .A(fracta_mul[22]), .B(fracta_mul[21]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__22_) );
  MUX2_X2 sll_386_M1_0_23 ( .A(fracta_mul[23]), .B(fracta_mul[22]), .S(
        sll_386_n4), .Z(sll_386_ML_int_1__23_) );
  MUX2_X2 sll_386_M1_0_24 ( .A(fracta_mul[24]), .B(fracta_mul[23]), .S(
        sll_386_n4), .Z(sll_386_ML_int_1__24_) );
  MUX2_X2 sll_386_M1_0_25 ( .A(fracta_mul[25]), .B(fracta_mul[24]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__25_) );
  MUX2_X2 sll_386_M1_0_26 ( .A(fracta_mul[26]), .B(fracta_mul[25]), .S(
        sll_386_n4), .Z(sll_386_ML_int_1__26_) );
  MUX2_X2 sll_386_M1_0_27 ( .A(fracta_mul[27]), .B(fracta_mul[26]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__27_) );
  MUX2_X2 sll_386_M1_0_28 ( .A(fracta_mul[28]), .B(fracta_mul[27]), .S(
        sll_386_n4), .Z(sll_386_ML_int_1__28_) );
  MUX2_X2 sll_386_M1_0_29 ( .A(fracta_mul[29]), .B(fracta_mul[28]), .S(
        sll_386_n4), .Z(sll_386_ML_int_1__29_) );
  MUX2_X2 sll_386_M1_0_30 ( .A(fracta_mul[30]), .B(fracta_mul[29]), .S(
        sll_386_n4), .Z(sll_386_ML_int_1__30_) );
  MUX2_X2 sll_386_M1_0_31 ( .A(fracta_mul[31]), .B(fracta_mul[30]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__31_) );
  MUX2_X2 sll_386_M1_0_32 ( .A(fracta_mul[32]), .B(fracta_mul[31]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__32_) );
  MUX2_X2 sll_386_M1_0_33 ( .A(fracta_mul[33]), .B(fracta_mul[32]), .S(
        sll_386_n4), .Z(sll_386_ML_int_1__33_) );
  MUX2_X2 sll_386_M1_0_34 ( .A(fracta_mul[34]), .B(fracta_mul[33]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__34_) );
  MUX2_X2 sll_386_M1_0_35 ( .A(fracta_mul[35]), .B(fracta_mul[34]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__35_) );
  MUX2_X2 sll_386_M1_0_36 ( .A(fracta_mul[36]), .B(fracta_mul[35]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__36_) );
  MUX2_X2 sll_386_M1_0_37 ( .A(fracta_mul[37]), .B(fracta_mul[36]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__37_) );
  MUX2_X2 sll_386_M1_0_38 ( .A(fracta_mul[38]), .B(fracta_mul[37]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__38_) );
  MUX2_X2 sll_386_M1_0_39 ( .A(fracta_mul[39]), .B(fracta_mul[38]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__39_) );
  MUX2_X2 sll_386_M1_0_40 ( .A(fracta_mul[40]), .B(fracta_mul[39]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__40_) );
  MUX2_X2 sll_386_M1_0_41 ( .A(fracta_mul[41]), .B(fracta_mul[40]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__41_) );
  MUX2_X2 sll_386_M1_0_42 ( .A(fracta_mul[42]), .B(fracta_mul[41]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__42_) );
  MUX2_X2 sll_386_M1_0_43 ( .A(fracta_mul[43]), .B(fracta_mul[42]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__43_) );
  MUX2_X2 sll_386_M1_0_44 ( .A(fracta_mul[44]), .B(fracta_mul[43]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__44_) );
  MUX2_X2 sll_386_M1_0_45 ( .A(fracta_mul[45]), .B(fracta_mul[44]), .S(
        sll_386_n4), .Z(sll_386_ML_int_1__45_) );
  MUX2_X2 sll_386_M1_0_46 ( .A(fracta_mul[46]), .B(fracta_mul[45]), .S(
        sll_386_n4), .Z(sll_386_ML_int_1__46_) );
  MUX2_X2 sll_386_M1_0_47 ( .A(fracta_mul[47]), .B(fracta_mul[46]), .S(
        sll_386_n4), .Z(sll_386_ML_int_1__47_) );
  MUX2_X2 sll_386_M1_0_48 ( .A(fracta_mul[48]), .B(fracta_mul[47]), .S(
        sll_386_n4), .Z(sll_386_ML_int_1__48_) );
  MUX2_X2 sll_386_M1_0_49 ( .A(fracta_mul[49]), .B(fracta_mul[48]), .S(
        sll_386_n4), .Z(sll_386_ML_int_1__49_) );
  MUX2_X2 sll_386_M1_0_50 ( .A(fracta_mul[50]), .B(fracta_mul[49]), .S(
        sll_386_n4), .Z(sll_386_ML_int_1__50_) );
  MUX2_X2 sll_386_M1_0_51 ( .A(fracta_mul[51]), .B(fracta_mul[50]), .S(
        sll_386_n4), .Z(sll_386_ML_int_1__51_) );
  MUX2_X2 sll_386_M1_0_52 ( .A(u2_N157), .B(fracta_mul[51]), .S(sll_386_n4), 
        .Z(sll_386_ML_int_1__52_) );
  MUX2_X2 sll_386_M1_1_2 ( .A(sll_386_ML_int_1__2_), .B(sll_386_ML_int_1__0_), 
        .S(sll_386_n5), .Z(sll_386_ML_int_2__2_) );
  MUX2_X2 sll_386_M1_1_3 ( .A(sll_386_ML_int_1__3_), .B(sll_386_ML_int_1__1_), 
        .S(sll_386_n5), .Z(sll_386_ML_int_2__3_) );
  MUX2_X2 sll_386_M1_1_4 ( .A(sll_386_ML_int_1__4_), .B(sll_386_ML_int_1__2_), 
        .S(sll_386_n5), .Z(sll_386_ML_int_2__4_) );
  MUX2_X2 sll_386_M1_1_5 ( .A(sll_386_ML_int_1__5_), .B(sll_386_ML_int_1__3_), 
        .S(sll_386_n5), .Z(sll_386_ML_int_2__5_) );
  MUX2_X2 sll_386_M1_1_6 ( .A(sll_386_ML_int_1__6_), .B(sll_386_ML_int_1__4_), 
        .S(sll_386_n5), .Z(sll_386_ML_int_2__6_) );
  MUX2_X2 sll_386_M1_1_7 ( .A(sll_386_ML_int_1__7_), .B(sll_386_ML_int_1__5_), 
        .S(sll_386_n5), .Z(sll_386_ML_int_2__7_) );
  MUX2_X2 sll_386_M1_1_8 ( .A(sll_386_ML_int_1__8_), .B(sll_386_ML_int_1__6_), 
        .S(sll_386_n5), .Z(sll_386_ML_int_2__8_) );
  MUX2_X2 sll_386_M1_1_9 ( .A(sll_386_ML_int_1__9_), .B(sll_386_ML_int_1__7_), 
        .S(sll_386_n5), .Z(sll_386_ML_int_2__9_) );
  MUX2_X2 sll_386_M1_1_10 ( .A(sll_386_ML_int_1__10_), .B(sll_386_ML_int_1__8_), .S(sll_386_n5), .Z(sll_386_ML_int_2__10_) );
  MUX2_X2 sll_386_M1_1_11 ( .A(sll_386_ML_int_1__11_), .B(sll_386_ML_int_1__9_), .S(sll_386_n5), .Z(sll_386_ML_int_2__11_) );
  MUX2_X2 sll_386_M1_1_12 ( .A(sll_386_ML_int_1__12_), .B(
        sll_386_ML_int_1__10_), .S(sll_386_n5), .Z(sll_386_ML_int_2__12_) );
  MUX2_X2 sll_386_M1_1_13 ( .A(sll_386_ML_int_1__13_), .B(
        sll_386_ML_int_1__11_), .S(sll_386_n6), .Z(sll_386_ML_int_2__13_) );
  MUX2_X2 sll_386_M1_1_14 ( .A(sll_386_ML_int_1__14_), .B(
        sll_386_ML_int_1__12_), .S(sll_386_n6), .Z(sll_386_ML_int_2__14_) );
  MUX2_X2 sll_386_M1_1_15 ( .A(sll_386_ML_int_1__15_), .B(
        sll_386_ML_int_1__13_), .S(sll_386_n6), .Z(sll_386_ML_int_2__15_) );
  MUX2_X2 sll_386_M1_1_16 ( .A(sll_386_ML_int_1__16_), .B(
        sll_386_ML_int_1__14_), .S(sll_386_n6), .Z(sll_386_ML_int_2__16_) );
  MUX2_X2 sll_386_M1_1_17 ( .A(sll_386_ML_int_1__17_), .B(
        sll_386_ML_int_1__15_), .S(sll_386_n6), .Z(sll_386_ML_int_2__17_) );
  MUX2_X2 sll_386_M1_1_18 ( .A(sll_386_ML_int_1__18_), .B(
        sll_386_ML_int_1__16_), .S(sll_386_n6), .Z(sll_386_ML_int_2__18_) );
  MUX2_X2 sll_386_M1_1_19 ( .A(sll_386_ML_int_1__19_), .B(
        sll_386_ML_int_1__17_), .S(sll_386_n6), .Z(sll_386_ML_int_2__19_) );
  MUX2_X2 sll_386_M1_1_20 ( .A(sll_386_ML_int_1__20_), .B(
        sll_386_ML_int_1__18_), .S(sll_386_n6), .Z(sll_386_ML_int_2__20_) );
  MUX2_X2 sll_386_M1_1_21 ( .A(sll_386_ML_int_1__21_), .B(
        sll_386_ML_int_1__19_), .S(sll_386_n6), .Z(sll_386_ML_int_2__21_) );
  MUX2_X2 sll_386_M1_1_22 ( .A(sll_386_ML_int_1__22_), .B(
        sll_386_ML_int_1__20_), .S(sll_386_n6), .Z(sll_386_ML_int_2__22_) );
  MUX2_X2 sll_386_M1_1_23 ( .A(sll_386_ML_int_1__23_), .B(
        sll_386_ML_int_1__21_), .S(sll_386_n6), .Z(sll_386_ML_int_2__23_) );
  MUX2_X2 sll_386_M1_1_24 ( .A(sll_386_ML_int_1__24_), .B(
        sll_386_ML_int_1__22_), .S(sll_386_n7), .Z(sll_386_ML_int_2__24_) );
  MUX2_X2 sll_386_M1_1_25 ( .A(sll_386_ML_int_1__25_), .B(
        sll_386_ML_int_1__23_), .S(sll_386_n7), .Z(sll_386_ML_int_2__25_) );
  MUX2_X2 sll_386_M1_1_26 ( .A(sll_386_ML_int_1__26_), .B(
        sll_386_ML_int_1__24_), .S(sll_386_n7), .Z(sll_386_ML_int_2__26_) );
  MUX2_X2 sll_386_M1_1_27 ( .A(sll_386_ML_int_1__27_), .B(
        sll_386_ML_int_1__25_), .S(sll_386_n7), .Z(sll_386_ML_int_2__27_) );
  MUX2_X2 sll_386_M1_1_28 ( .A(sll_386_ML_int_1__28_), .B(
        sll_386_ML_int_1__26_), .S(sll_386_n7), .Z(sll_386_ML_int_2__28_) );
  MUX2_X2 sll_386_M1_1_29 ( .A(sll_386_ML_int_1__29_), .B(
        sll_386_ML_int_1__27_), .S(sll_386_n7), .Z(sll_386_ML_int_2__29_) );
  MUX2_X2 sll_386_M1_1_30 ( .A(sll_386_ML_int_1__30_), .B(
        sll_386_ML_int_1__28_), .S(sll_386_n7), .Z(sll_386_ML_int_2__30_) );
  MUX2_X2 sll_386_M1_1_31 ( .A(sll_386_ML_int_1__31_), .B(
        sll_386_ML_int_1__29_), .S(sll_386_n7), .Z(sll_386_ML_int_2__31_) );
  MUX2_X2 sll_386_M1_1_32 ( .A(sll_386_ML_int_1__32_), .B(
        sll_386_ML_int_1__30_), .S(sll_386_n7), .Z(sll_386_ML_int_2__32_) );
  MUX2_X2 sll_386_M1_1_33 ( .A(sll_386_ML_int_1__33_), .B(
        sll_386_ML_int_1__31_), .S(sll_386_n7), .Z(sll_386_ML_int_2__33_) );
  MUX2_X2 sll_386_M1_1_34 ( .A(sll_386_ML_int_1__34_), .B(
        sll_386_ML_int_1__32_), .S(sll_386_n7), .Z(sll_386_ML_int_2__34_) );
  MUX2_X2 sll_386_M1_1_35 ( .A(sll_386_ML_int_1__35_), .B(
        sll_386_ML_int_1__33_), .S(sll_386_n7), .Z(sll_386_ML_int_2__35_) );
  MUX2_X2 sll_386_M1_1_36 ( .A(sll_386_ML_int_1__36_), .B(
        sll_386_ML_int_1__34_), .S(sll_386_n7), .Z(sll_386_ML_int_2__36_) );
  MUX2_X2 sll_386_M1_1_37 ( .A(sll_386_ML_int_1__37_), .B(
        sll_386_ML_int_1__35_), .S(sll_386_n7), .Z(sll_386_ML_int_2__37_) );
  MUX2_X2 sll_386_M1_1_38 ( .A(sll_386_ML_int_1__38_), .B(
        sll_386_ML_int_1__36_), .S(sll_386_n7), .Z(sll_386_ML_int_2__38_) );
  MUX2_X2 sll_386_M1_1_39 ( .A(sll_386_ML_int_1__39_), .B(
        sll_386_ML_int_1__37_), .S(sll_386_n7), .Z(sll_386_ML_int_2__39_) );
  MUX2_X2 sll_386_M1_1_40 ( .A(sll_386_ML_int_1__40_), .B(
        sll_386_ML_int_1__38_), .S(sll_386_n7), .Z(sll_386_ML_int_2__40_) );
  MUX2_X2 sll_386_M1_1_41 ( .A(sll_386_ML_int_1__41_), .B(
        sll_386_ML_int_1__39_), .S(sll_386_n7), .Z(sll_386_ML_int_2__41_) );
  MUX2_X2 sll_386_M1_1_42 ( .A(sll_386_ML_int_1__42_), .B(
        sll_386_ML_int_1__40_), .S(sll_386_n7), .Z(sll_386_ML_int_2__42_) );
  MUX2_X2 sll_386_M1_1_43 ( .A(sll_386_ML_int_1__43_), .B(
        sll_386_ML_int_1__41_), .S(sll_386_n7), .Z(sll_386_ML_int_2__43_) );
  MUX2_X2 sll_386_M1_1_44 ( .A(sll_386_ML_int_1__44_), .B(
        sll_386_ML_int_1__42_), .S(sll_386_n7), .Z(sll_386_ML_int_2__44_) );
  MUX2_X2 sll_386_M1_1_45 ( .A(sll_386_ML_int_1__45_), .B(
        sll_386_ML_int_1__43_), .S(sll_386_n7), .Z(sll_386_ML_int_2__45_) );
  MUX2_X2 sll_386_M1_1_46 ( .A(sll_386_ML_int_1__46_), .B(
        sll_386_ML_int_1__44_), .S(sll_386_n7), .Z(sll_386_ML_int_2__46_) );
  MUX2_X2 sll_386_M1_1_47 ( .A(sll_386_ML_int_1__47_), .B(
        sll_386_ML_int_1__45_), .S(sll_386_n7), .Z(sll_386_ML_int_2__47_) );
  MUX2_X2 sll_386_M1_1_48 ( .A(sll_386_ML_int_1__48_), .B(
        sll_386_ML_int_1__46_), .S(sll_386_n7), .Z(sll_386_ML_int_2__48_) );
  MUX2_X2 sll_386_M1_1_49 ( .A(sll_386_ML_int_1__49_), .B(
        sll_386_ML_int_1__47_), .S(sll_386_n7), .Z(sll_386_ML_int_2__49_) );
  MUX2_X2 sll_386_M1_1_50 ( .A(sll_386_ML_int_1__50_), .B(
        sll_386_ML_int_1__48_), .S(sll_386_n7), .Z(sll_386_ML_int_2__50_) );
  MUX2_X2 sll_386_M1_1_51 ( .A(sll_386_ML_int_1__51_), .B(
        sll_386_ML_int_1__49_), .S(sll_386_n7), .Z(sll_386_ML_int_2__51_) );
  MUX2_X2 sll_386_M1_1_52 ( .A(sll_386_ML_int_1__52_), .B(
        sll_386_ML_int_1__50_), .S(sll_386_n7), .Z(sll_386_ML_int_2__52_) );
  MUX2_X2 sll_386_M1_2_4 ( .A(sll_386_ML_int_2__4_), .B(sll_386_ML_int_2__0_), 
        .S(sll_386_n9), .Z(sll_386_ML_int_3__4_) );
  MUX2_X2 sll_386_M1_2_5 ( .A(sll_386_ML_int_2__5_), .B(sll_386_ML_int_2__1_), 
        .S(sll_386_n9), .Z(sll_386_ML_int_3__5_) );
  MUX2_X2 sll_386_M1_2_6 ( .A(sll_386_ML_int_2__6_), .B(sll_386_ML_int_2__2_), 
        .S(sll_386_n9), .Z(sll_386_ML_int_3__6_) );
  MUX2_X2 sll_386_M1_2_7 ( .A(sll_386_ML_int_2__7_), .B(sll_386_ML_int_2__3_), 
        .S(sll_386_n9), .Z(sll_386_ML_int_3__7_) );
  MUX2_X2 sll_386_M1_2_8 ( .A(sll_386_ML_int_2__8_), .B(sll_386_ML_int_2__4_), 
        .S(sll_386_n9), .Z(sll_386_ML_int_3__8_) );
  MUX2_X2 sll_386_M1_2_9 ( .A(sll_386_ML_int_2__9_), .B(sll_386_ML_int_2__5_), 
        .S(sll_386_n9), .Z(sll_386_ML_int_3__9_) );
  MUX2_X2 sll_386_M1_2_10 ( .A(sll_386_ML_int_2__10_), .B(sll_386_ML_int_2__6_), .S(sll_386_n9), .Z(sll_386_ML_int_3__10_) );
  MUX2_X2 sll_386_M1_2_11 ( .A(sll_386_ML_int_2__11_), .B(sll_386_ML_int_2__7_), .S(sll_386_n9), .Z(sll_386_ML_int_3__11_) );
  MUX2_X2 sll_386_M1_2_12 ( .A(sll_386_ML_int_2__12_), .B(sll_386_ML_int_2__8_), .S(sll_386_n9), .Z(sll_386_ML_int_3__12_) );
  MUX2_X2 sll_386_M1_2_13 ( .A(sll_386_ML_int_2__13_), .B(sll_386_ML_int_2__9_), .S(sll_386_n9), .Z(sll_386_ML_int_3__13_) );
  MUX2_X2 sll_386_M1_2_14 ( .A(sll_386_ML_int_2__14_), .B(
        sll_386_ML_int_2__10_), .S(sll_386_n9), .Z(sll_386_ML_int_3__14_) );
  MUX2_X2 sll_386_M1_2_15 ( .A(sll_386_ML_int_2__15_), .B(
        sll_386_ML_int_2__11_), .S(sll_386_n10), .Z(sll_386_ML_int_3__15_) );
  MUX2_X2 sll_386_M1_2_16 ( .A(sll_386_ML_int_2__16_), .B(
        sll_386_ML_int_2__12_), .S(sll_386_n10), .Z(sll_386_ML_int_3__16_) );
  MUX2_X2 sll_386_M1_2_17 ( .A(sll_386_ML_int_2__17_), .B(
        sll_386_ML_int_2__13_), .S(sll_386_n10), .Z(sll_386_ML_int_3__17_) );
  MUX2_X2 sll_386_M1_2_18 ( .A(sll_386_ML_int_2__18_), .B(
        sll_386_ML_int_2__14_), .S(sll_386_n10), .Z(sll_386_ML_int_3__18_) );
  MUX2_X2 sll_386_M1_2_19 ( .A(sll_386_ML_int_2__19_), .B(
        sll_386_ML_int_2__15_), .S(sll_386_n10), .Z(sll_386_ML_int_3__19_) );
  MUX2_X2 sll_386_M1_2_20 ( .A(sll_386_ML_int_2__20_), .B(
        sll_386_ML_int_2__16_), .S(sll_386_n10), .Z(sll_386_ML_int_3__20_) );
  MUX2_X2 sll_386_M1_2_21 ( .A(sll_386_ML_int_2__21_), .B(
        sll_386_ML_int_2__17_), .S(sll_386_n10), .Z(sll_386_ML_int_3__21_) );
  MUX2_X2 sll_386_M1_2_22 ( .A(sll_386_ML_int_2__22_), .B(
        sll_386_ML_int_2__18_), .S(sll_386_n10), .Z(sll_386_ML_int_3__22_) );
  MUX2_X2 sll_386_M1_2_23 ( .A(sll_386_ML_int_2__23_), .B(
        sll_386_ML_int_2__19_), .S(sll_386_n10), .Z(sll_386_ML_int_3__23_) );
  MUX2_X2 sll_386_M1_2_24 ( .A(sll_386_ML_int_2__24_), .B(
        sll_386_ML_int_2__20_), .S(sll_386_n10), .Z(sll_386_ML_int_3__24_) );
  MUX2_X2 sll_386_M1_2_25 ( .A(sll_386_ML_int_2__25_), .B(
        sll_386_ML_int_2__21_), .S(sll_386_n10), .Z(sll_386_ML_int_3__25_) );
  MUX2_X2 sll_386_M1_2_26 ( .A(sll_386_ML_int_2__26_), .B(
        sll_386_ML_int_2__22_), .S(sll_386_n11), .Z(sll_386_ML_int_3__26_) );
  MUX2_X2 sll_386_M1_2_27 ( .A(sll_386_ML_int_2__27_), .B(
        sll_386_ML_int_2__23_), .S(sll_386_n11), .Z(sll_386_ML_int_3__27_) );
  MUX2_X2 sll_386_M1_2_28 ( .A(sll_386_ML_int_2__28_), .B(
        sll_386_ML_int_2__24_), .S(sll_386_n11), .Z(sll_386_ML_int_3__28_) );
  MUX2_X2 sll_386_M1_2_29 ( .A(sll_386_ML_int_2__29_), .B(
        sll_386_ML_int_2__25_), .S(sll_386_n11), .Z(sll_386_ML_int_3__29_) );
  MUX2_X2 sll_386_M1_2_30 ( .A(sll_386_ML_int_2__30_), .B(
        sll_386_ML_int_2__26_), .S(sll_386_n11), .Z(sll_386_ML_int_3__30_) );
  MUX2_X2 sll_386_M1_2_31 ( .A(sll_386_ML_int_2__31_), .B(
        sll_386_ML_int_2__27_), .S(sll_386_n11), .Z(sll_386_ML_int_3__31_) );
  MUX2_X2 sll_386_M1_2_32 ( .A(sll_386_ML_int_2__32_), .B(
        sll_386_ML_int_2__28_), .S(sll_386_n11), .Z(sll_386_ML_int_3__32_) );
  MUX2_X2 sll_386_M1_2_33 ( .A(sll_386_ML_int_2__33_), .B(
        sll_386_ML_int_2__29_), .S(sll_386_n11), .Z(sll_386_ML_int_3__33_) );
  MUX2_X2 sll_386_M1_2_34 ( .A(sll_386_ML_int_2__34_), .B(
        sll_386_ML_int_2__30_), .S(sll_386_n11), .Z(sll_386_ML_int_3__34_) );
  MUX2_X2 sll_386_M1_2_35 ( .A(sll_386_ML_int_2__35_), .B(
        sll_386_ML_int_2__31_), .S(sll_386_n11), .Z(sll_386_ML_int_3__35_) );
  MUX2_X2 sll_386_M1_2_36 ( .A(sll_386_ML_int_2__36_), .B(
        sll_386_ML_int_2__32_), .S(sll_386_n11), .Z(sll_386_ML_int_3__36_) );
  MUX2_X2 sll_386_M1_2_37 ( .A(sll_386_ML_int_2__37_), .B(
        sll_386_ML_int_2__33_), .S(sll_386_n12), .Z(sll_386_ML_int_3__37_) );
  MUX2_X2 sll_386_M1_2_38 ( .A(sll_386_ML_int_2__38_), .B(
        sll_386_ML_int_2__34_), .S(sll_386_n12), .Z(sll_386_ML_int_3__38_) );
  MUX2_X2 sll_386_M1_2_39 ( .A(sll_386_ML_int_2__39_), .B(
        sll_386_ML_int_2__35_), .S(sll_386_n12), .Z(sll_386_ML_int_3__39_) );
  MUX2_X2 sll_386_M1_2_40 ( .A(sll_386_ML_int_2__40_), .B(
        sll_386_ML_int_2__36_), .S(sll_386_n12), .Z(sll_386_ML_int_3__40_) );
  MUX2_X2 sll_386_M1_2_41 ( .A(sll_386_ML_int_2__41_), .B(
        sll_386_ML_int_2__37_), .S(sll_386_n12), .Z(sll_386_ML_int_3__41_) );
  MUX2_X2 sll_386_M1_2_42 ( .A(sll_386_ML_int_2__42_), .B(
        sll_386_ML_int_2__38_), .S(sll_386_n12), .Z(sll_386_ML_int_3__42_) );
  MUX2_X2 sll_386_M1_2_43 ( .A(sll_386_ML_int_2__43_), .B(
        sll_386_ML_int_2__39_), .S(sll_386_n12), .Z(sll_386_ML_int_3__43_) );
  MUX2_X2 sll_386_M1_2_44 ( .A(sll_386_ML_int_2__44_), .B(
        sll_386_ML_int_2__40_), .S(sll_386_n12), .Z(sll_386_ML_int_3__44_) );
  MUX2_X2 sll_386_M1_2_45 ( .A(sll_386_ML_int_2__45_), .B(
        sll_386_ML_int_2__41_), .S(sll_386_n12), .Z(sll_386_ML_int_3__45_) );
  MUX2_X2 sll_386_M1_2_46 ( .A(sll_386_ML_int_2__46_), .B(
        sll_386_ML_int_2__42_), .S(sll_386_n12), .Z(sll_386_ML_int_3__46_) );
  MUX2_X2 sll_386_M1_2_47 ( .A(sll_386_ML_int_2__47_), .B(
        sll_386_ML_int_2__43_), .S(sll_386_n12), .Z(sll_386_ML_int_3__47_) );
  MUX2_X2 sll_386_M1_2_48 ( .A(sll_386_ML_int_2__48_), .B(
        sll_386_ML_int_2__44_), .S(sll_386_n12), .Z(sll_386_ML_int_3__48_) );
  MUX2_X2 sll_386_M1_2_49 ( .A(sll_386_ML_int_2__49_), .B(
        sll_386_ML_int_2__45_), .S(sll_386_n12), .Z(sll_386_ML_int_3__49_) );
  MUX2_X2 sll_386_M1_2_50 ( .A(sll_386_ML_int_2__50_), .B(
        sll_386_ML_int_2__46_), .S(sll_386_n12), .Z(sll_386_ML_int_3__50_) );
  MUX2_X2 sll_386_M1_2_51 ( .A(sll_386_ML_int_2__51_), .B(
        sll_386_ML_int_2__47_), .S(sll_386_n12), .Z(sll_386_ML_int_3__51_) );
  MUX2_X2 sll_386_M1_2_52 ( .A(sll_386_ML_int_2__52_), .B(
        sll_386_ML_int_2__48_), .S(sll_386_n12), .Z(sll_386_ML_int_3__52_) );
  MUX2_X2 sll_386_M1_3_8 ( .A(sll_386_ML_int_3__8_), .B(sll_386_ML_int_3__0_), 
        .S(sll_386_n16), .Z(sll_386_ML_int_4__8_) );
  MUX2_X2 sll_386_M1_3_9 ( .A(sll_386_ML_int_3__9_), .B(sll_386_ML_int_3__1_), 
        .S(sll_386_n16), .Z(sll_386_ML_int_4__9_) );
  MUX2_X2 sll_386_M1_3_10 ( .A(sll_386_ML_int_3__10_), .B(sll_386_ML_int_3__2_), .S(sll_386_n16), .Z(sll_386_ML_int_4__10_) );
  MUX2_X2 sll_386_M1_3_11 ( .A(sll_386_ML_int_3__11_), .B(sll_386_ML_int_3__3_), .S(sll_386_n16), .Z(sll_386_ML_int_4__11_) );
  MUX2_X2 sll_386_M1_3_12 ( .A(sll_386_ML_int_3__12_), .B(sll_386_ML_int_3__4_), .S(sll_386_n16), .Z(sll_386_ML_int_4__12_) );
  MUX2_X2 sll_386_M1_3_13 ( .A(sll_386_ML_int_3__13_), .B(sll_386_ML_int_3__5_), .S(sll_386_n16), .Z(sll_386_ML_int_4__13_) );
  MUX2_X2 sll_386_M1_3_14 ( .A(sll_386_ML_int_3__14_), .B(sll_386_ML_int_3__6_), .S(sll_386_n16), .Z(sll_386_ML_int_4__14_) );
  MUX2_X2 sll_386_M1_3_15 ( .A(sll_386_ML_int_3__15_), .B(sll_386_ML_int_3__7_), .S(sll_386_n16), .Z(sll_386_ML_int_4__15_) );
  MUX2_X2 sll_386_M1_3_16 ( .A(sll_386_ML_int_3__16_), .B(sll_386_ML_int_3__8_), .S(sll_386_n16), .Z(sll_386_ML_int_4__16_) );
  MUX2_X2 sll_386_M1_3_17 ( .A(sll_386_ML_int_3__17_), .B(sll_386_ML_int_3__9_), .S(sll_386_n16), .Z(sll_386_ML_int_4__17_) );
  MUX2_X2 sll_386_M1_3_18 ( .A(sll_386_ML_int_3__18_), .B(
        sll_386_ML_int_3__10_), .S(sll_386_n16), .Z(sll_386_ML_int_4__18_) );
  MUX2_X2 sll_386_M1_3_19 ( .A(sll_386_ML_int_3__19_), .B(
        sll_386_ML_int_3__11_), .S(sll_386_n17), .Z(sll_386_ML_int_4__19_) );
  MUX2_X2 sll_386_M1_3_20 ( .A(sll_386_ML_int_3__20_), .B(
        sll_386_ML_int_3__12_), .S(sll_386_n17), .Z(sll_386_ML_int_4__20_) );
  MUX2_X2 sll_386_M1_3_21 ( .A(sll_386_ML_int_3__21_), .B(
        sll_386_ML_int_3__13_), .S(sll_386_n17), .Z(sll_386_ML_int_4__21_) );
  MUX2_X2 sll_386_M1_3_22 ( .A(sll_386_ML_int_3__22_), .B(
        sll_386_ML_int_3__14_), .S(sll_386_n17), .Z(sll_386_ML_int_4__22_) );
  MUX2_X2 sll_386_M1_3_23 ( .A(sll_386_ML_int_3__23_), .B(
        sll_386_ML_int_3__15_), .S(sll_386_n17), .Z(sll_386_ML_int_4__23_) );
  MUX2_X2 sll_386_M1_3_24 ( .A(sll_386_ML_int_3__24_), .B(
        sll_386_ML_int_3__16_), .S(sll_386_n17), .Z(sll_386_ML_int_4__24_) );
  MUX2_X2 sll_386_M1_3_25 ( .A(sll_386_ML_int_3__25_), .B(
        sll_386_ML_int_3__17_), .S(sll_386_n17), .Z(sll_386_ML_int_4__25_) );
  MUX2_X2 sll_386_M1_3_26 ( .A(sll_386_ML_int_3__26_), .B(
        sll_386_ML_int_3__18_), .S(sll_386_n17), .Z(sll_386_ML_int_4__26_) );
  MUX2_X2 sll_386_M1_3_27 ( .A(sll_386_ML_int_3__27_), .B(
        sll_386_ML_int_3__19_), .S(sll_386_n17), .Z(sll_386_ML_int_4__27_) );
  MUX2_X2 sll_386_M1_3_28 ( .A(sll_386_ML_int_3__28_), .B(
        sll_386_ML_int_3__20_), .S(sll_386_n17), .Z(sll_386_ML_int_4__28_) );
  MUX2_X2 sll_386_M1_3_29 ( .A(sll_386_ML_int_3__29_), .B(
        sll_386_ML_int_3__21_), .S(sll_386_n17), .Z(sll_386_ML_int_4__29_) );
  MUX2_X2 sll_386_M1_3_30 ( .A(sll_386_ML_int_3__30_), .B(
        sll_386_ML_int_3__22_), .S(sll_386_n18), .Z(sll_386_ML_int_4__30_) );
  MUX2_X2 sll_386_M1_3_31 ( .A(sll_386_ML_int_3__31_), .B(
        sll_386_ML_int_3__23_), .S(sll_386_n18), .Z(sll_386_ML_int_4__31_) );
  MUX2_X2 sll_386_M1_3_32 ( .A(sll_386_ML_int_3__32_), .B(
        sll_386_ML_int_3__24_), .S(sll_386_n18), .Z(sll_386_ML_int_4__32_) );
  MUX2_X2 sll_386_M1_3_33 ( .A(sll_386_ML_int_3__33_), .B(
        sll_386_ML_int_3__25_), .S(sll_386_n18), .Z(sll_386_ML_int_4__33_) );
  MUX2_X2 sll_386_M1_3_34 ( .A(sll_386_ML_int_3__34_), .B(
        sll_386_ML_int_3__26_), .S(sll_386_n18), .Z(sll_386_ML_int_4__34_) );
  MUX2_X2 sll_386_M1_3_35 ( .A(sll_386_ML_int_3__35_), .B(
        sll_386_ML_int_3__27_), .S(sll_386_n18), .Z(sll_386_ML_int_4__35_) );
  MUX2_X2 sll_386_M1_3_36 ( .A(sll_386_ML_int_3__36_), .B(
        sll_386_ML_int_3__28_), .S(sll_386_n18), .Z(sll_386_ML_int_4__36_) );
  MUX2_X2 sll_386_M1_3_37 ( .A(sll_386_ML_int_3__37_), .B(
        sll_386_ML_int_3__29_), .S(sll_386_n18), .Z(sll_386_ML_int_4__37_) );
  MUX2_X2 sll_386_M1_3_38 ( .A(sll_386_ML_int_3__38_), .B(
        sll_386_ML_int_3__30_), .S(sll_386_n18), .Z(sll_386_ML_int_4__38_) );
  MUX2_X2 sll_386_M1_3_39 ( .A(sll_386_ML_int_3__39_), .B(
        sll_386_ML_int_3__31_), .S(sll_386_n18), .Z(sll_386_ML_int_4__39_) );
  MUX2_X2 sll_386_M1_3_40 ( .A(sll_386_ML_int_3__40_), .B(
        sll_386_ML_int_3__32_), .S(sll_386_n18), .Z(sll_386_ML_int_4__40_) );
  MUX2_X2 sll_386_M1_3_41 ( .A(sll_386_ML_int_3__41_), .B(
        sll_386_ML_int_3__33_), .S(sll_386_n19), .Z(sll_386_ML_int_4__41_) );
  MUX2_X2 sll_386_M1_3_42 ( .A(sll_386_ML_int_3__42_), .B(
        sll_386_ML_int_3__34_), .S(sll_386_n19), .Z(sll_386_ML_int_4__42_) );
  MUX2_X2 sll_386_M1_3_43 ( .A(sll_386_ML_int_3__43_), .B(
        sll_386_ML_int_3__35_), .S(sll_386_n19), .Z(sll_386_ML_int_4__43_) );
  MUX2_X2 sll_386_M1_3_44 ( .A(sll_386_ML_int_3__44_), .B(
        sll_386_ML_int_3__36_), .S(sll_386_n19), .Z(sll_386_ML_int_4__44_) );
  MUX2_X2 sll_386_M1_3_45 ( .A(sll_386_ML_int_3__45_), .B(
        sll_386_ML_int_3__37_), .S(sll_386_n19), .Z(sll_386_ML_int_4__45_) );
  MUX2_X2 sll_386_M1_3_46 ( .A(sll_386_ML_int_3__46_), .B(
        sll_386_ML_int_3__38_), .S(sll_386_n19), .Z(sll_386_ML_int_4__46_) );
  MUX2_X2 sll_386_M1_3_47 ( .A(sll_386_ML_int_3__47_), .B(
        sll_386_ML_int_3__39_), .S(sll_386_n19), .Z(sll_386_ML_int_4__47_) );
  MUX2_X2 sll_386_M1_3_48 ( .A(sll_386_ML_int_3__48_), .B(
        sll_386_ML_int_3__40_), .S(sll_386_n19), .Z(sll_386_ML_int_4__48_) );
  MUX2_X2 sll_386_M1_3_49 ( .A(sll_386_ML_int_3__49_), .B(
        sll_386_ML_int_3__41_), .S(sll_386_n19), .Z(sll_386_ML_int_4__49_) );
  MUX2_X2 sll_386_M1_3_50 ( .A(sll_386_ML_int_3__50_), .B(
        sll_386_ML_int_3__42_), .S(sll_386_n19), .Z(sll_386_ML_int_4__50_) );
  MUX2_X2 sll_386_M1_3_51 ( .A(sll_386_ML_int_3__51_), .B(
        sll_386_ML_int_3__43_), .S(sll_386_n19), .Z(sll_386_ML_int_4__51_) );
  MUX2_X2 sll_386_M1_3_52 ( .A(sll_386_ML_int_3__52_), .B(
        sll_386_ML_int_3__44_), .S(sll_386_n19), .Z(sll_386_ML_int_4__52_) );
  MUX2_X2 sll_386_M1_4_16 ( .A(sll_386_ML_int_4__16_), .B(sll_386_n29), .S(
        sll_386_n24), .Z(N272) );
  MUX2_X2 sll_386_M1_4_17 ( .A(sll_386_ML_int_4__17_), .B(sll_386_n28), .S(
        div_opa_ldz_d[4]), .Z(N273) );
  MUX2_X2 sll_386_M1_4_18 ( .A(sll_386_ML_int_4__18_), .B(sll_386_n27), .S(
        div_opa_ldz_d[4]), .Z(N274) );
  MUX2_X2 sll_386_M1_4_19 ( .A(sll_386_ML_int_4__19_), .B(sll_386_n26), .S(
        div_opa_ldz_d[4]), .Z(N275) );
  MUX2_X2 sll_386_M1_4_20 ( .A(sll_386_ML_int_4__20_), .B(sll_386_n30), .S(
        sll_386_n24), .Z(N276) );
  MUX2_X2 sll_386_M1_4_21 ( .A(sll_386_ML_int_4__21_), .B(sll_386_n31), .S(
        sll_386_n24), .Z(N277) );
  MUX2_X2 sll_386_M1_4_22 ( .A(sll_386_ML_int_4__22_), .B(sll_386_n32), .S(
        sll_386_n24), .Z(N278) );
  MUX2_X2 sll_386_M1_4_23 ( .A(sll_386_ML_int_4__23_), .B(sll_386_n33), .S(
        sll_386_n24), .Z(N279) );
  MUX2_X2 sll_386_M1_4_24 ( .A(sll_386_ML_int_4__24_), .B(sll_386_ML_int_4__8_), .S(sll_386_n24), .Z(N280) );
  MUX2_X2 sll_386_M1_4_25 ( .A(sll_386_ML_int_4__25_), .B(sll_386_ML_int_4__9_), .S(sll_386_n24), .Z(N281) );
  MUX2_X2 sll_386_M1_4_26 ( .A(sll_386_ML_int_4__26_), .B(
        sll_386_ML_int_4__10_), .S(sll_386_n24), .Z(N282) );
  MUX2_X2 sll_386_M1_4_27 ( .A(sll_386_ML_int_4__27_), .B(
        sll_386_ML_int_4__11_), .S(sll_386_n24), .Z(N283) );
  MUX2_X2 sll_386_M1_4_28 ( .A(sll_386_ML_int_4__28_), .B(
        sll_386_ML_int_4__12_), .S(sll_386_n24), .Z(N284) );
  MUX2_X2 sll_386_M1_4_29 ( .A(sll_386_ML_int_4__29_), .B(
        sll_386_ML_int_4__13_), .S(sll_386_n24), .Z(N285) );
  MUX2_X2 sll_386_M1_4_30 ( .A(sll_386_ML_int_4__30_), .B(
        sll_386_ML_int_4__14_), .S(sll_386_n24), .Z(N286) );
  MUX2_X2 sll_386_M1_4_31 ( .A(sll_386_ML_int_4__31_), .B(
        sll_386_ML_int_4__15_), .S(sll_386_n23), .Z(N287) );
  MUX2_X2 sll_386_M1_4_32 ( .A(sll_386_ML_int_4__32_), .B(
        sll_386_ML_int_4__16_), .S(sll_386_n23), .Z(N288) );
  MUX2_X2 sll_386_M1_4_33 ( .A(sll_386_ML_int_4__33_), .B(
        sll_386_ML_int_4__17_), .S(sll_386_n23), .Z(N289) );
  MUX2_X2 sll_386_M1_4_34 ( .A(sll_386_ML_int_4__34_), .B(
        sll_386_ML_int_4__18_), .S(sll_386_n23), .Z(N290) );
  MUX2_X2 sll_386_M1_4_35 ( .A(sll_386_ML_int_4__35_), .B(
        sll_386_ML_int_4__19_), .S(sll_386_n23), .Z(N291) );
  MUX2_X2 sll_386_M1_4_36 ( .A(sll_386_ML_int_4__36_), .B(
        sll_386_ML_int_4__20_), .S(sll_386_n23), .Z(N292) );
  MUX2_X2 sll_386_M1_4_37 ( .A(sll_386_ML_int_4__37_), .B(
        sll_386_ML_int_4__21_), .S(sll_386_n23), .Z(N293) );
  MUX2_X2 sll_386_M1_4_38 ( .A(sll_386_ML_int_4__38_), .B(
        sll_386_ML_int_4__22_), .S(sll_386_n23), .Z(N294) );
  MUX2_X2 sll_386_M1_4_39 ( .A(sll_386_ML_int_4__39_), .B(
        sll_386_ML_int_4__23_), .S(sll_386_n23), .Z(N295) );
  MUX2_X2 sll_386_M1_4_40 ( .A(sll_386_ML_int_4__40_), .B(
        sll_386_ML_int_4__24_), .S(sll_386_n23), .Z(N296) );
  MUX2_X2 sll_386_M1_4_41 ( .A(sll_386_ML_int_4__41_), .B(
        sll_386_ML_int_4__25_), .S(sll_386_n23), .Z(N297) );
  MUX2_X2 sll_386_M1_4_42 ( .A(sll_386_ML_int_4__42_), .B(
        sll_386_ML_int_4__26_), .S(sll_386_n22), .Z(N298) );
  MUX2_X2 sll_386_M1_4_43 ( .A(sll_386_ML_int_4__43_), .B(
        sll_386_ML_int_4__27_), .S(sll_386_n22), .Z(N299) );
  MUX2_X2 sll_386_M1_4_44 ( .A(sll_386_ML_int_4__44_), .B(
        sll_386_ML_int_4__28_), .S(sll_386_n22), .Z(N300) );
  MUX2_X2 sll_386_M1_4_45 ( .A(sll_386_ML_int_4__45_), .B(
        sll_386_ML_int_4__29_), .S(sll_386_n22), .Z(N301) );
  MUX2_X2 sll_386_M1_4_46 ( .A(sll_386_ML_int_4__46_), .B(
        sll_386_ML_int_4__30_), .S(sll_386_n22), .Z(N302) );
  MUX2_X2 sll_386_M1_4_47 ( .A(sll_386_ML_int_4__47_), .B(
        sll_386_ML_int_4__31_), .S(sll_386_n22), .Z(N303) );
  MUX2_X2 sll_386_M1_4_48 ( .A(sll_386_ML_int_4__48_), .B(
        sll_386_ML_int_4__32_), .S(sll_386_n22), .Z(N304) );
  MUX2_X2 sll_386_M1_4_49 ( .A(sll_386_ML_int_4__49_), .B(
        sll_386_ML_int_4__33_), .S(sll_386_n22), .Z(N305) );
  MUX2_X2 sll_386_M1_4_50 ( .A(sll_386_ML_int_4__50_), .B(
        sll_386_ML_int_4__34_), .S(sll_386_n22), .Z(N306) );
  MUX2_X2 sll_386_M1_4_51 ( .A(sll_386_ML_int_4__51_), .B(
        sll_386_ML_int_4__35_), .S(sll_386_n22), .Z(N307) );
  MUX2_X2 sll_386_M1_4_52 ( .A(sll_386_ML_int_4__52_), .B(
        sll_386_ML_int_4__36_), .S(sll_386_n22), .Z(N308) );
  NAND2_X1 r471_U180 ( .A1(fracta_mul[49]), .A2(r471_n7), .ZN(r471_n168) );
  OR2_X1 r471_U179 ( .A1(r471_n1), .A2(u6_N50), .ZN(r471_n167) );
  AND2_X1 r471_U178 ( .A1(fracta_mul[0]), .A2(r471_n56), .ZN(r471_n178) );
  OAI22_X1 r471_U177 ( .A1(n4770), .A2(r471_n178), .B1(r471_n178), .B2(
        r471_n55), .ZN(r471_n177) );
  AND3_X1 r471_U176 ( .A1(r471_n168), .A2(r471_n167), .A3(r471_n177), .ZN(
        r471_n176) );
  NAND2_X1 r471_U175 ( .A1(fracta_mul[48]), .A2(r471_n8), .ZN(r471_n93) );
  NAND2_X1 r471_U174 ( .A1(fracta_mul[46]), .A2(r471_n10), .ZN(r471_n97) );
  NAND2_X1 r471_U173 ( .A1(fracta_mul[47]), .A2(r471_n9), .ZN(r471_n94) );
  AND4_X1 r471_U172 ( .A1(r471_n176), .A2(r471_n93), .A3(r471_n97), .A4(
        r471_n94), .ZN(r471_n169) );
  NAND2_X1 r471_U171 ( .A1(fracta_mul[42]), .A2(r471_n14), .ZN(r471_n105) );
  NAND2_X1 r471_U170 ( .A1(fracta_mul[41]), .A2(r471_n15), .ZN(r471_n106) );
  NAND2_X1 r471_U169 ( .A1(fracta_mul[40]), .A2(r471_n16), .ZN(r471_n109) );
  NAND2_X1 r471_U168 ( .A1(fracta_mul[39]), .A2(r471_n17), .ZN(r471_n110) );
  AND4_X1 r471_U167 ( .A1(r471_n105), .A2(r471_n106), .A3(r471_n109), .A4(
        r471_n110), .ZN(r471_n175) );
  NAND2_X1 r471_U166 ( .A1(fracta_mul[45]), .A2(r471_n11), .ZN(r471_n98) );
  NAND2_X1 r471_U165 ( .A1(fracta_mul[43]), .A2(r471_n13), .ZN(r471_n102) );
  NAND2_X1 r471_U164 ( .A1(fracta_mul[44]), .A2(r471_n12), .ZN(r471_n101) );
  AND4_X1 r471_U163 ( .A1(r471_n175), .A2(r471_n98), .A3(r471_n102), .A4(
        r471_n101), .ZN(r471_n170) );
  NAND2_X1 r471_U162 ( .A1(fracta_mul[34]), .A2(r471_n22), .ZN(r471_n121) );
  NAND2_X1 r471_U161 ( .A1(fracta_mul[33]), .A2(r471_n23), .ZN(r471_n122) );
  NAND2_X1 r471_U160 ( .A1(fracta_mul[35]), .A2(r471_n21), .ZN(r471_n118) );
  AND3_X1 r471_U159 ( .A1(r471_n121), .A2(r471_n122), .A3(r471_n118), .ZN(
        r471_n174) );
  NAND2_X1 r471_U158 ( .A1(fracta_mul[38]), .A2(r471_n18), .ZN(r471_n113) );
  NAND2_X1 r471_U157 ( .A1(fracta_mul[36]), .A2(r471_n20), .ZN(r471_n117) );
  NAND2_X1 r471_U156 ( .A1(fracta_mul[37]), .A2(r471_n19), .ZN(r471_n114) );
  AND4_X1 r471_U155 ( .A1(r471_n174), .A2(r471_n113), .A3(r471_n117), .A4(
        r471_n114), .ZN(r471_n171) );
  NAND2_X1 r471_U154 ( .A1(fracta_mul[29]), .A2(r471_n27), .ZN(r471_n130) );
  NAND2_X1 r471_U153 ( .A1(fracta_mul[28]), .A2(r471_n28), .ZN(r471_n133) );
  NAND2_X1 r471_U152 ( .A1(fracta_mul[27]), .A2(r471_n29), .ZN(r471_n134) );
  NAND2_X1 r471_U151 ( .A1(fracta_mul[26]), .A2(r471_n30), .ZN(r471_n137) );
  AND4_X1 r471_U150 ( .A1(r471_n130), .A2(r471_n133), .A3(r471_n134), .A4(
        r471_n137), .ZN(r471_n173) );
  NAND2_X1 r471_U149 ( .A1(fracta_mul[32]), .A2(r471_n24), .ZN(r471_n125) );
  NAND2_X1 r471_U148 ( .A1(fracta_mul[30]), .A2(r471_n26), .ZN(r471_n129) );
  NAND2_X1 r471_U147 ( .A1(fracta_mul[31]), .A2(r471_n25), .ZN(r471_n126) );
  AND4_X1 r471_U146 ( .A1(r471_n173), .A2(r471_n125), .A3(r471_n129), .A4(
        r471_n126), .ZN(r471_n172) );
  NAND4_X1 r471_U145 ( .A1(r471_n169), .A2(r471_n170), .A3(r471_n171), .A4(
        r471_n172), .ZN(r471_n57) );
  NAND2_X1 r471_U144 ( .A1(fracta_mul[6]), .A2(r471_n50), .ZN(r471_n158) );
  NAND2_X1 r471_U143 ( .A1(fracta_mul[4]), .A2(r471_n52), .ZN(r471_n162) );
  NAND2_X1 r471_U142 ( .A1(fracta_mul[5]), .A2(r471_n51), .ZN(r471_n159) );
  AND3_X1 r471_U141 ( .A1(r471_n158), .A2(r471_n162), .A3(r471_n159), .ZN(
        r471_n76) );
  AND2_X1 r471_U140 ( .A1(fracta_mul[51]), .A2(r471_n6), .ZN(r471_n86) );
  AND2_X1 r471_U139 ( .A1(r471_n167), .A2(r471_n168), .ZN(r471_n90) );
  NAND2_X1 r471_U138 ( .A1(fracta_mul[25]), .A2(r471_n31), .ZN(r471_n63) );
  NAND2_X1 r471_U137 ( .A1(fracta_mul[24]), .A2(r471_n32), .ZN(r471_n61) );
  NAND2_X1 r471_U136 ( .A1(fracta_mul[23]), .A2(r471_n33), .ZN(r471_n62) );
  NAND2_X1 r471_U135 ( .A1(fracta_mul[22]), .A2(r471_n34), .ZN(r471_n65) );
  NAND2_X1 r471_U134 ( .A1(fracta_mul[21]), .A2(r471_n35), .ZN(r471_n67) );
  NAND2_X1 r471_U133 ( .A1(fracta_mul[20]), .A2(r471_n36), .ZN(r471_n66) );
  NAND2_X1 r471_U132 ( .A1(fracta_mul[19]), .A2(r471_n37), .ZN(r471_n70) );
  NAND2_X1 r471_U131 ( .A1(fracta_mul[18]), .A2(r471_n38), .ZN(r471_n68) );
  NAND2_X1 r471_U130 ( .A1(fracta_mul[17]), .A2(r471_n39), .ZN(r471_n69) );
  NAND2_X1 r471_U129 ( .A1(fracta_mul[16]), .A2(r471_n40), .ZN(r471_n75) );
  NAND2_X1 r471_U128 ( .A1(fracta_mul[15]), .A2(r471_n41), .ZN(r471_n74) );
  NAND2_X1 r471_U127 ( .A1(fracta_mul[14]), .A2(r471_n42), .ZN(r471_n73) );
  NAND2_X1 r471_U126 ( .A1(fracta_mul[13]), .A2(r471_n43), .ZN(r471_n72) );
  NAND2_X1 r471_U125 ( .A1(fracta_mul[12]), .A2(r471_n44), .ZN(r471_n80) );
  NAND2_X1 r471_U124 ( .A1(fracta_mul[11]), .A2(r471_n45), .ZN(r471_n82) );
  NAND2_X1 r471_U123 ( .A1(fracta_mul[10]), .A2(r471_n46), .ZN(r471_n81) );
  NAND2_X1 r471_U122 ( .A1(fracta_mul[9]), .A2(r471_n47), .ZN(r471_n85) );
  NAND2_X1 r471_U121 ( .A1(fracta_mul[8]), .A2(r471_n48), .ZN(r471_n83) );
  NAND2_X1 r471_U120 ( .A1(fracta_mul[7]), .A2(r471_n49), .ZN(r471_n84) );
  NAND2_X1 r471_U119 ( .A1(n4727), .A2(r471_n53), .ZN(r471_n87) );
  NOR2_X1 r471_U118 ( .A1(r471_n56), .A2(fracta_mul[0]), .ZN(r471_n165) );
  OAI211_X1 r471_U117 ( .C1(r471_n165), .C2(r471_n4), .A(r471_n166), .B(
        r471_n88), .ZN(r471_n164) );
  NAND3_X1 r471_U116 ( .A1(r471_n162), .A2(r471_n87), .A3(r471_n163), .ZN(
        r471_n161) );
  OAI221_X1 r471_U115 ( .B1(fracta_mul[4]), .B2(r471_n52), .C1(fracta_mul[5]), 
        .C2(r471_n51), .A(r471_n161), .ZN(r471_n160) );
  NAND3_X1 r471_U114 ( .A1(r471_n158), .A2(r471_n159), .A3(r471_n160), .ZN(
        r471_n157) );
  OAI221_X1 r471_U113 ( .B1(fracta_mul[6]), .B2(r471_n50), .C1(fracta_mul[7]), 
        .C2(r471_n49), .A(r471_n157), .ZN(r471_n156) );
  NAND3_X1 r471_U112 ( .A1(r471_n83), .A2(r471_n84), .A3(r471_n156), .ZN(
        r471_n155) );
  OAI221_X1 r471_U111 ( .B1(fracta_mul[8]), .B2(r471_n48), .C1(fracta_mul[9]), 
        .C2(r471_n47), .A(r471_n155), .ZN(r471_n154) );
  NAND3_X1 r471_U110 ( .A1(r471_n81), .A2(r471_n85), .A3(r471_n154), .ZN(
        r471_n153) );
  OAI221_X1 r471_U109 ( .B1(fracta_mul[10]), .B2(r471_n46), .C1(fracta_mul[11]), .C2(r471_n45), .A(r471_n153), .ZN(r471_n152) );
  NAND3_X1 r471_U108 ( .A1(r471_n80), .A2(r471_n82), .A3(r471_n152), .ZN(
        r471_n151) );
  OAI221_X1 r471_U107 ( .B1(fracta_mul[12]), .B2(r471_n44), .C1(fracta_mul[13]), .C2(r471_n43), .A(r471_n151), .ZN(r471_n150) );
  NAND3_X1 r471_U106 ( .A1(r471_n73), .A2(r471_n72), .A3(r471_n150), .ZN(
        r471_n149) );
  OAI221_X1 r471_U105 ( .B1(fracta_mul[14]), .B2(r471_n42), .C1(fracta_mul[15]), .C2(r471_n41), .A(r471_n149), .ZN(r471_n148) );
  NAND3_X1 r471_U104 ( .A1(r471_n75), .A2(r471_n74), .A3(r471_n148), .ZN(
        r471_n147) );
  OAI221_X1 r471_U103 ( .B1(fracta_mul[16]), .B2(r471_n40), .C1(fracta_mul[17]), .C2(r471_n39), .A(r471_n147), .ZN(r471_n146) );
  NAND3_X1 r471_U102 ( .A1(r471_n68), .A2(r471_n69), .A3(r471_n146), .ZN(
        r471_n145) );
  OAI221_X1 r471_U101 ( .B1(fracta_mul[18]), .B2(r471_n38), .C1(fracta_mul[19]), .C2(r471_n37), .A(r471_n145), .ZN(r471_n144) );
  NAND3_X1 r471_U100 ( .A1(r471_n66), .A2(r471_n70), .A3(r471_n144), .ZN(
        r471_n143) );
  OAI221_X1 r471_U99 ( .B1(fracta_mul[20]), .B2(r471_n36), .C1(fracta_mul[21]), 
        .C2(r471_n35), .A(r471_n143), .ZN(r471_n142) );
  NAND3_X1 r471_U98 ( .A1(r471_n65), .A2(r471_n67), .A3(r471_n142), .ZN(
        r471_n141) );
  OAI221_X1 r471_U97 ( .B1(fracta_mul[22]), .B2(r471_n34), .C1(fracta_mul[23]), 
        .C2(r471_n33), .A(r471_n141), .ZN(r471_n140) );
  NAND3_X1 r471_U96 ( .A1(r471_n61), .A2(r471_n62), .A3(r471_n140), .ZN(
        r471_n139) );
  OAI221_X1 r471_U95 ( .B1(fracta_mul[24]), .B2(r471_n32), .C1(fracta_mul[25]), 
        .C2(r471_n31), .A(r471_n139), .ZN(r471_n138) );
  NAND3_X1 r471_U94 ( .A1(r471_n137), .A2(r471_n63), .A3(r471_n138), .ZN(
        r471_n136) );
  OAI221_X1 r471_U93 ( .B1(fracta_mul[26]), .B2(r471_n30), .C1(fracta_mul[27]), 
        .C2(r471_n29), .A(r471_n136), .ZN(r471_n135) );
  NAND3_X1 r471_U92 ( .A1(r471_n133), .A2(r471_n134), .A3(r471_n135), .ZN(
        r471_n132) );
  OAI221_X1 r471_U91 ( .B1(fracta_mul[28]), .B2(r471_n28), .C1(fracta_mul[29]), 
        .C2(r471_n27), .A(r471_n132), .ZN(r471_n131) );
  NAND3_X1 r471_U90 ( .A1(r471_n129), .A2(r471_n130), .A3(r471_n131), .ZN(
        r471_n128) );
  OAI221_X1 r471_U89 ( .B1(fracta_mul[30]), .B2(r471_n26), .C1(fracta_mul[31]), 
        .C2(r471_n25), .A(r471_n128), .ZN(r471_n127) );
  NAND3_X1 r471_U88 ( .A1(r471_n125), .A2(r471_n126), .A3(r471_n127), .ZN(
        r471_n124) );
  OAI221_X1 r471_U87 ( .B1(fracta_mul[32]), .B2(r471_n24), .C1(fracta_mul[33]), 
        .C2(r471_n23), .A(r471_n124), .ZN(r471_n123) );
  NAND3_X1 r471_U86 ( .A1(r471_n121), .A2(r471_n122), .A3(r471_n123), .ZN(
        r471_n120) );
  OAI221_X1 r471_U85 ( .B1(fracta_mul[34]), .B2(r471_n22), .C1(fracta_mul[35]), 
        .C2(r471_n21), .A(r471_n120), .ZN(r471_n119) );
  NAND3_X1 r471_U84 ( .A1(r471_n117), .A2(r471_n118), .A3(r471_n119), .ZN(
        r471_n116) );
  OAI221_X1 r471_U83 ( .B1(fracta_mul[36]), .B2(r471_n20), .C1(fracta_mul[37]), 
        .C2(r471_n19), .A(r471_n116), .ZN(r471_n115) );
  NAND3_X1 r471_U82 ( .A1(r471_n113), .A2(r471_n114), .A3(r471_n115), .ZN(
        r471_n112) );
  OAI221_X1 r471_U81 ( .B1(fracta_mul[38]), .B2(r471_n18), .C1(fracta_mul[39]), 
        .C2(r471_n17), .A(r471_n112), .ZN(r471_n111) );
  NAND3_X1 r471_U80 ( .A1(r471_n109), .A2(r471_n110), .A3(r471_n111), .ZN(
        r471_n108) );
  OAI221_X1 r471_U79 ( .B1(fracta_mul[40]), .B2(r471_n16), .C1(fracta_mul[41]), 
        .C2(r471_n15), .A(r471_n108), .ZN(r471_n107) );
  NAND3_X1 r471_U78 ( .A1(r471_n105), .A2(r471_n106), .A3(r471_n107), .ZN(
        r471_n104) );
  OAI221_X1 r471_U77 ( .B1(fracta_mul[42]), .B2(r471_n14), .C1(fracta_mul[43]), 
        .C2(r471_n13), .A(r471_n104), .ZN(r471_n103) );
  NAND3_X1 r471_U76 ( .A1(r471_n101), .A2(r471_n102), .A3(r471_n103), .ZN(
        r471_n100) );
  OAI221_X1 r471_U75 ( .B1(fracta_mul[44]), .B2(r471_n12), .C1(fracta_mul[45]), 
        .C2(r471_n11), .A(r471_n100), .ZN(r471_n99) );
  NAND3_X1 r471_U74 ( .A1(r471_n97), .A2(r471_n98), .A3(r471_n99), .ZN(
        r471_n96) );
  OAI221_X1 r471_U73 ( .B1(fracta_mul[46]), .B2(r471_n10), .C1(fracta_mul[47]), 
        .C2(r471_n9), .A(r471_n96), .ZN(r471_n95) );
  NAND3_X1 r471_U72 ( .A1(r471_n93), .A2(r471_n94), .A3(r471_n95), .ZN(
        r471_n92) );
  OAI221_X1 r471_U71 ( .B1(fracta_mul[48]), .B2(r471_n8), .C1(fracta_mul[49]), 
        .C2(r471_n7), .A(r471_n92), .ZN(r471_n91) );
  AOI22_X1 r471_U70 ( .A1(u6_N50), .A2(r471_n1), .B1(r471_n90), .B2(r471_n91), 
        .ZN(r471_n89) );
  OAI22_X1 r471_U69 ( .A1(fracta_mul[51]), .A2(r471_n6), .B1(r471_n86), .B2(
        r471_n89), .ZN(u1_N219) );
  NOR4_X1 r471_U68 ( .A1(u1_N219), .A2(r471_n86), .A3(r471_n3), .A4(r471_n2), 
        .ZN(r471_n77) );
  AND3_X1 r471_U67 ( .A1(r471_n83), .A2(r471_n84), .A3(r471_n85), .ZN(r471_n79) );
  AND4_X1 r471_U66 ( .A1(r471_n79), .A2(r471_n80), .A3(r471_n81), .A4(r471_n82), .ZN(r471_n78) );
  NAND3_X1 r471_U65 ( .A1(r471_n76), .A2(r471_n77), .A3(r471_n78), .ZN(
        r471_n58) );
  AND4_X1 r471_U64 ( .A1(r471_n72), .A2(r471_n73), .A3(r471_n74), .A4(r471_n75), .ZN(r471_n71) );
  NAND4_X1 r471_U63 ( .A1(r471_n68), .A2(r471_n69), .A3(r471_n70), .A4(
        r471_n71), .ZN(r471_n59) );
  AND3_X1 r471_U62 ( .A1(r471_n65), .A2(r471_n66), .A3(r471_n67), .ZN(r471_n64) );
  NAND4_X1 r471_U61 ( .A1(r471_n61), .A2(r471_n62), .A3(r471_n63), .A4(
        r471_n64), .ZN(r471_n60) );
  NOR4_X1 r471_U60 ( .A1(r471_n57), .A2(r471_n58), .A3(r471_n59), .A4(r471_n60), .ZN(u1_N220) );
  INV_X4 r471_U59 ( .A(u6_N0), .ZN(r471_n56) );
  INV_X4 r471_U58 ( .A(u6_N1), .ZN(r471_n55) );
  INV_X4 r471_U57 ( .A(u6_N2), .ZN(r471_n54) );
  INV_X4 r471_U56 ( .A(u6_N3), .ZN(r471_n53) );
  INV_X4 r471_U55 ( .A(u6_N4), .ZN(r471_n52) );
  INV_X4 r471_U54 ( .A(u6_N5), .ZN(r471_n51) );
  INV_X4 r471_U53 ( .A(u6_N6), .ZN(r471_n50) );
  INV_X4 r471_U52 ( .A(u6_N7), .ZN(r471_n49) );
  INV_X4 r471_U51 ( .A(u6_N8), .ZN(r471_n48) );
  INV_X4 r471_U50 ( .A(u6_N9), .ZN(r471_n47) );
  INV_X4 r471_U49 ( .A(u6_N10), .ZN(r471_n46) );
  INV_X4 r471_U48 ( .A(u6_N11), .ZN(r471_n45) );
  INV_X4 r471_U47 ( .A(u6_N12), .ZN(r471_n44) );
  INV_X4 r471_U46 ( .A(u6_N13), .ZN(r471_n43) );
  INV_X4 r471_U45 ( .A(u6_N14), .ZN(r471_n42) );
  INV_X4 r471_U44 ( .A(u6_N15), .ZN(r471_n41) );
  INV_X4 r471_U43 ( .A(u6_N16), .ZN(r471_n40) );
  INV_X4 r471_U42 ( .A(u6_N17), .ZN(r471_n39) );
  INV_X4 r471_U41 ( .A(u6_N18), .ZN(r471_n38) );
  INV_X4 r471_U40 ( .A(u6_N20), .ZN(r471_n36) );
  INV_X4 r471_U39 ( .A(u6_N21), .ZN(r471_n35) );
  INV_X4 r471_U38 ( .A(u6_N22), .ZN(r471_n34) );
  INV_X4 r471_U37 ( .A(u6_N23), .ZN(r471_n33) );
  INV_X4 r471_U36 ( .A(u6_N26), .ZN(r471_n30) );
  INV_X4 r471_U35 ( .A(u6_N27), .ZN(r471_n29) );
  INV_X4 r471_U34 ( .A(u6_N49), .ZN(r471_n7) );
  INV_X4 r471_U33 ( .A(r471_n165), .ZN(r471_n5) );
  INV_X4 r471_U32 ( .A(r471_n88), .ZN(r471_n3) );
  INV_X4 r471_U31 ( .A(r471_n87), .ZN(r471_n2) );
  INV_X4 r471_U30 ( .A(fracta_mul[50]), .ZN(r471_n1) );
  INV_X1 r471_U29 ( .A(u6_N51), .ZN(r471_n6) );
  INV_X1 r471_U28 ( .A(n4770), .ZN(r471_n4) );
  OAI21_X1 r471_U27 ( .B1(n4770), .B2(r471_n5), .A(r471_n55), .ZN(r471_n166)
         );
  INV_X1 r471_U26 ( .A(u6_N48), .ZN(r471_n8) );
  NAND2_X2 r471_U25 ( .A1(fracta_mul[2]), .A2(r471_n54), .ZN(r471_n88) );
  INV_X1 r471_U24 ( .A(n4424), .ZN(r471_n9) );
  INV_X1 r471_U23 ( .A(u6_N43), .ZN(r471_n13) );
  INV_X1 r471_U22 ( .A(u6_N46), .ZN(r471_n10) );
  INV_X1 r471_U21 ( .A(u6_N45), .ZN(r471_n11) );
  INV_X1 r471_U20 ( .A(n4765), .ZN(r471_n12) );
  INV_X1 r471_U19 ( .A(n4787), .ZN(r471_n14) );
  INV_X1 r471_U18 ( .A(u6_N37), .ZN(r471_n19) );
  INV_X1 r471_U17 ( .A(u6_N40), .ZN(r471_n16) );
  INV_X1 r471_U16 ( .A(u6_N35), .ZN(r471_n21) );
  INV_X1 r471_U15 ( .A(n4786), .ZN(r471_n22) );
  INV_X2 r471_U14 ( .A(u6_N33), .ZN(r471_n23) );
  INV_X1 r471_U13 ( .A(n4772), .ZN(r471_n15) );
  INV_X1 r471_U12 ( .A(u6_N29), .ZN(r471_n27) );
  INV_X1 r471_U11 ( .A(u6_N30), .ZN(r471_n26) );
  INV_X1 r471_U10 ( .A(u6_N39), .ZN(r471_n17) );
  INV_X1 r471_U9 ( .A(u6_N36), .ZN(r471_n20) );
  INV_X2 r471_U8 ( .A(u6_N24), .ZN(r471_n32) );
  INV_X1 r471_U7 ( .A(u6_N32), .ZN(r471_n24) );
  INV_X2 r471_U6 ( .A(u6_N25), .ZN(r471_n31) );
  INV_X1 r471_U5 ( .A(u6_N31), .ZN(r471_n25) );
  INV_X2 r471_U4 ( .A(u6_N19), .ZN(r471_n37) );
  OAI221_X2 r471_U3 ( .B1(fracta_mul[2]), .B2(r471_n54), .C1(n4727), .C2(
        r471_n53), .A(r471_n164), .ZN(r471_n163) );
  INV_X4 r471_U2 ( .A(n4791), .ZN(r471_n18) );
  INV_X4 r471_U1 ( .A(n4764), .ZN(r471_n28) );
  INV_X4 add_0_root_sub_0_root_u4_add_497_U10 ( .A(
        add_0_root_sub_0_root_u4_add_497_n7), .ZN(u4_div_exp3[0]) );
  INV_X4 add_0_root_sub_0_root_u4_add_497_U9 ( .A(
        add_0_root_sub_0_root_u4_add_497_n6), .ZN(
        add_0_root_sub_0_root_u4_add_497_carry_9_) );
  NAND2_X2 add_0_root_sub_0_root_u4_add_497_U8 ( .A1(u4_ldz_dif_8_), .A2(
        add_0_root_sub_0_root_u4_add_497_carry_8_), .ZN(
        add_0_root_sub_0_root_u4_add_497_n6) );
  INV_X4 add_0_root_sub_0_root_u4_add_497_U7 ( .A(
        add_0_root_sub_0_root_u4_add_497_n5), .ZN(
        add_0_root_sub_0_root_u4_add_497_carry_10_) );
  NAND2_X2 add_0_root_sub_0_root_u4_add_497_U6 ( .A1(u4_ldz_dif_9_), .A2(
        add_0_root_sub_0_root_u4_add_497_carry_9_), .ZN(
        add_0_root_sub_0_root_u4_add_497_n5) );
  XNOR2_X1 add_0_root_sub_0_root_u4_add_497_U5 ( .A(n4526), .B(u4_ldz_dif_0_), 
        .ZN(add_0_root_sub_0_root_u4_add_497_n7) );
  XOR2_X2 add_0_root_sub_0_root_u4_add_497_U4 ( .A(u4_ldz_dif_9_), .B(
        add_0_root_sub_0_root_u4_add_497_carry_9_), .Z(u4_div_exp3[9]) );
  XOR2_X2 add_0_root_sub_0_root_u4_add_497_U3 ( .A(u4_ldz_dif_10_), .B(
        add_0_root_sub_0_root_u4_add_497_carry_10_), .Z(u4_div_exp3[10]) );
  XOR2_X2 add_0_root_sub_0_root_u4_add_497_U2 ( .A(u4_ldz_dif_8_), .B(
        add_0_root_sub_0_root_u4_add_497_carry_8_), .Z(u4_div_exp3[8]) );
  AND2_X2 add_0_root_sub_0_root_u4_add_497_U1 ( .A1(n4526), .A2(u4_ldz_dif_0_), 
        .ZN(add_0_root_sub_0_root_u4_add_497_n1) );
  FA_X1 add_0_root_sub_0_root_u4_add_497_U1_1 ( .A(u4_ldz_dif_1_), .B(n7207), 
        .CI(add_0_root_sub_0_root_u4_add_497_n1), .CO(
        add_0_root_sub_0_root_u4_add_497_carry_2_), .S(u4_div_exp3[1]) );
  FA_X1 add_0_root_sub_0_root_u4_add_497_U1_2 ( .A(u4_ldz_dif_2_), .B(
        u4_fi_ldz_2a_2_), .CI(add_0_root_sub_0_root_u4_add_497_carry_2_), .CO(
        add_0_root_sub_0_root_u4_add_497_carry_3_), .S(u4_div_exp3[2]) );
  FA_X1 add_0_root_sub_0_root_u4_add_497_U1_3 ( .A(u4_ldz_dif_3_), .B(net44706), .CI(add_0_root_sub_0_root_u4_add_497_carry_3_), .CO(
        add_0_root_sub_0_root_u4_add_497_carry_4_), .S(u4_div_exp3[3]) );
  FA_X1 add_0_root_sub_0_root_u4_add_497_U1_4 ( .A(u4_ldz_dif_4_), .B(
        u4_fi_ldz_2a_4_), .CI(add_0_root_sub_0_root_u4_add_497_carry_4_), .CO(
        add_0_root_sub_0_root_u4_add_497_carry_5_), .S(u4_div_exp3[4]) );
  FA_X1 add_0_root_sub_0_root_u4_add_497_U1_5 ( .A(u4_ldz_dif_5_), .B(
        u4_fi_ldz_2a_5_), .CI(add_0_root_sub_0_root_u4_add_497_carry_5_), .CO(
        add_0_root_sub_0_root_u4_add_497_carry_6_), .S(u4_div_exp3[5]) );
  FA_X1 add_0_root_sub_0_root_u4_add_497_U1_6 ( .A(u4_ldz_dif_6_), .B(
        u4_fi_ldz_2a_6_), .CI(add_0_root_sub_0_root_u4_add_497_carry_6_), .CO(
        add_0_root_sub_0_root_u4_add_497_carry_7_), .S(u4_div_exp3[6]) );
  FA_X1 add_0_root_sub_0_root_u4_add_497_U1_7 ( .A(u4_ldz_dif_7_), .B(
        u4_fi_ldz_2a_6_), .CI(add_0_root_sub_0_root_u4_add_497_carry_7_), .CO(
        add_0_root_sub_0_root_u4_add_497_carry_8_), .S(u4_div_exp3[7]) );
  NOR2_X4 u5_mult_82_U12973 ( .A1(u5_mult_82_net64899), .A2(
        u5_mult_82_net65225), .ZN(u5_mult_82_ab_50__35_) );
  NOR2_X4 u5_mult_82_U12972 ( .A1(u5_mult_82_net64379), .A2(u5_mult_82_n6755), 
        .ZN(u5_mult_82_ab_49__6_) );
  NOR2_X4 u5_mult_82_U12971 ( .A1(u5_mult_82_n6940), .A2(u5_mult_82_n6755), 
        .ZN(u5_mult_82_ab_49__7_) );
  NOR2_X4 u5_mult_82_U12970 ( .A1(u5_mult_82_net64455), .A2(u5_mult_82_n6755), 
        .ZN(u5_mult_82_ab_49__10_) );
  NOR2_X4 u5_mult_82_U12969 ( .A1(u5_mult_82_net64469), .A2(u5_mult_82_n6755), 
        .ZN(u5_mult_82_ab_49__11_) );
  NOR2_X4 u5_mult_82_U12968 ( .A1(u5_mult_82_net64505), .A2(u5_mult_82_n6755), 
        .ZN(u5_mult_82_ab_49__13_) );
  NOR2_X4 u5_mult_82_U12967 ( .A1(u5_mult_82_n6933), .A2(u5_mult_82_n6755), 
        .ZN(u5_mult_82_ab_49__15_) );
  NOR2_X4 u5_mult_82_U12966 ( .A1(u5_mult_82_net64559), .A2(u5_mult_82_n6754), 
        .ZN(u5_mult_82_ab_49__16_) );
  NOR2_X4 u5_mult_82_U12965 ( .A1(u5_mult_82_n6919), .A2(u5_mult_82_n6754), 
        .ZN(u5_mult_82_ab_49__18_) );
  NOR2_X4 u5_mult_82_U12964 ( .A1(u5_mult_82_net64665), .A2(u5_mult_82_n6754), 
        .ZN(u5_mult_82_ab_49__22_) );
  NOR2_X4 u5_mult_82_U12963 ( .A1(u5_mult_82_n6891), .A2(u5_mult_82_n6754), 
        .ZN(u5_mult_82_ab_49__24_) );
  NOR2_X4 u5_mult_82_U12962 ( .A1(u5_mult_82_n6884), .A2(u5_mult_82_n6754), 
        .ZN(u5_mult_82_ab_49__25_) );
  NOR2_X4 u5_mult_82_U12961 ( .A1(u5_mult_82_n6849), .A2(u5_mult_82_n6753), 
        .ZN(u5_mult_82_ab_49__31_) );
  NOR2_X4 u5_mult_82_U12960 ( .A1(u5_mult_82_n6837), .A2(u5_mult_82_n6753), 
        .ZN(u5_mult_82_ab_49__33_) );
  NOR2_X4 u5_mult_82_U12959 ( .A1(u5_mult_82_net64935), .A2(u5_mult_82_n6753), 
        .ZN(u5_mult_82_ab_49__37_) );
  NOR2_X4 u5_mult_82_U12958 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6753), 
        .ZN(u5_mult_82_ab_49__38_) );
  INV_X4 u5_mult_82_U12957 ( .A(fracta_mul[49]), .ZN(u5_mult_82_n7005) );
  NOR2_X4 u5_mult_82_U12956 ( .A1(u5_mult_82_n6967), .A2(u5_mult_82_n6749), 
        .ZN(u5_mult_82_ab_48__1_) );
  NOR2_X4 u5_mult_82_U12955 ( .A1(u5_mult_82_n6940), .A2(u5_mult_82_n6748), 
        .ZN(u5_mult_82_ab_48__7_) );
  NOR2_X4 u5_mult_82_U12954 ( .A1(u5_mult_82_net64415), .A2(u5_mult_82_n6748), 
        .ZN(u5_mult_82_ab_48__8_) );
  NOR2_X4 u5_mult_82_U12953 ( .A1(u5_mult_82_net64433), .A2(u5_mult_82_n6748), 
        .ZN(u5_mult_82_ab_48__9_) );
  NOR2_X4 u5_mult_82_U12952 ( .A1(u5_mult_82_net64455), .A2(u5_mult_82_n6748), 
        .ZN(u5_mult_82_ab_48__10_) );
  NOR2_X4 u5_mult_82_U12951 ( .A1(u5_mult_82_net64469), .A2(u5_mult_82_n6748), 
        .ZN(u5_mult_82_ab_48__11_) );
  NOR2_X4 u5_mult_82_U12950 ( .A1(u5_mult_82_net64487), .A2(u5_mult_82_n6748), 
        .ZN(u5_mult_82_ab_48__12_) );
  NOR2_X4 u5_mult_82_U12949 ( .A1(u5_mult_82_net64523), .A2(u5_mult_82_n6748), 
        .ZN(u5_mult_82_ab_48__14_) );
  NOR2_X4 u5_mult_82_U12948 ( .A1(u5_mult_82_n6933), .A2(u5_mult_82_n6748), 
        .ZN(u5_mult_82_ab_48__15_) );
  NOR2_X4 u5_mult_82_U12947 ( .A1(u5_mult_82_n6927), .A2(u5_mult_82_n6749), 
        .ZN(u5_mult_82_ab_48__17_) );
  NOR2_X4 u5_mult_82_U12946 ( .A1(u5_mult_82_n6919), .A2(u5_mult_82_n6749), 
        .ZN(u5_mult_82_ab_48__18_) );
  NOR2_X4 u5_mult_82_U12945 ( .A1(u5_mult_82_n6912), .A2(u5_mult_82_n6749), 
        .ZN(u5_mult_82_ab_48__19_) );
  NOR2_X4 u5_mult_82_U12944 ( .A1(u5_mult_82_n6903), .A2(u5_mult_82_n6749), 
        .ZN(u5_mult_82_ab_48__20_) );
  NOR2_X4 u5_mult_82_U12943 ( .A1(u5_mult_82_net64665), .A2(u5_mult_82_n6749), 
        .ZN(u5_mult_82_ab_48__22_) );
  NOR2_X4 u5_mult_82_U12942 ( .A1(u5_mult_82_n6891), .A2(u5_mult_82_n6749), 
        .ZN(u5_mult_82_ab_48__24_) );
  NOR2_X4 u5_mult_82_U12941 ( .A1(u5_mult_82_n6884), .A2(u5_mult_82_n6749), 
        .ZN(u5_mult_82_ab_48__25_) );
  NOR2_X4 u5_mult_82_U12940 ( .A1(u5_mult_82_n6856), .A2(u5_mult_82_n6747), 
        .ZN(u5_mult_82_ab_48__30_) );
  NOR2_X4 u5_mult_82_U12939 ( .A1(u5_mult_82_n6849), .A2(u5_mult_82_n6747), 
        .ZN(u5_mult_82_ab_48__31_) );
  NOR2_X4 u5_mult_82_U12938 ( .A1(u5_mult_82_n6842), .A2(u5_mult_82_n6747), 
        .ZN(u5_mult_82_ab_48__32_) );
  NOR2_X4 u5_mult_82_U12937 ( .A1(u5_mult_82_n6837), .A2(u5_mult_82_n6747), 
        .ZN(u5_mult_82_ab_48__33_) );
  NOR2_X4 u5_mult_82_U12936 ( .A1(u5_mult_82_net64881), .A2(u5_mult_82_n6747), 
        .ZN(u5_mult_82_ab_48__34_) );
  NOR2_X4 u5_mult_82_U12935 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6747), 
        .ZN(u5_mult_82_ab_48__38_) );
  NOR2_X4 u5_mult_82_U12934 ( .A1(u5_mult_82_n6826), .A2(u5_mult_82_n6746), 
        .ZN(u5_mult_82_ab_48__40_) );
  INV_X4 u5_mult_82_U12933 ( .A(fracta_mul[48]), .ZN(u5_mult_82_n7004) );
  NOR2_X4 u5_mult_82_U12932 ( .A1(u5_mult_82_n6967), .A2(u5_mult_82_net65285), 
        .ZN(u5_mult_82_ab_47__1_) );
  NOR2_X4 u5_mult_82_U12931 ( .A1(u5_mult_82_n6960), .A2(u5_mult_82_net65285), 
        .ZN(u5_mult_82_ab_47__2_) );
  NOR2_X4 u5_mult_82_U12930 ( .A1(u5_mult_82_net64361), .A2(
        u5_mult_82_net65283), .ZN(u5_mult_82_ab_47__5_) );
  NOR2_X4 u5_mult_82_U12929 ( .A1(u5_mult_82_n6940), .A2(u5_mult_82_net65283), 
        .ZN(u5_mult_82_ab_47__7_) );
  NOR2_X4 u5_mult_82_U12928 ( .A1(u5_mult_82_net64433), .A2(
        u5_mult_82_net65283), .ZN(u5_mult_82_ab_47__9_) );
  NOR2_X4 u5_mult_82_U12927 ( .A1(u5_mult_82_net64469), .A2(
        u5_mult_82_net65283), .ZN(u5_mult_82_ab_47__11_) );
  NOR2_X4 u5_mult_82_U12926 ( .A1(u5_mult_82_net64523), .A2(
        u5_mult_82_net65283), .ZN(u5_mult_82_ab_47__14_) );
  NOR2_X4 u5_mult_82_U12925 ( .A1(u5_mult_82_n6933), .A2(u5_mult_82_net65283), 
        .ZN(u5_mult_82_ab_47__15_) );
  NOR2_X4 u5_mult_82_U12924 ( .A1(u5_mult_82_net64559), .A2(
        u5_mult_82_net65285), .ZN(u5_mult_82_ab_47__16_) );
  NOR2_X4 u5_mult_82_U12923 ( .A1(u5_mult_82_n6927), .A2(u5_mult_82_net65285), 
        .ZN(u5_mult_82_ab_47__17_) );
  NOR2_X4 u5_mult_82_U12922 ( .A1(u5_mult_82_n6912), .A2(u5_mult_82_net65285), 
        .ZN(u5_mult_82_ab_47__19_) );
  NOR2_X4 u5_mult_82_U12921 ( .A1(u5_mult_82_n6903), .A2(u5_mult_82_net65285), 
        .ZN(u5_mult_82_ab_47__20_) );
  NOR2_X4 u5_mult_82_U12920 ( .A1(u5_mult_82_n6895), .A2(u5_mult_82_net65285), 
        .ZN(u5_mult_82_ab_47__21_) );
  NOR2_X4 u5_mult_82_U12919 ( .A1(u5_mult_82_n6861), .A2(u5_mult_82_net65279), 
        .ZN(u5_mult_82_ab_47__29_) );
  NOR2_X4 u5_mult_82_U12918 ( .A1(u5_mult_82_n6842), .A2(u5_mult_82_net65279), 
        .ZN(u5_mult_82_ab_47__32_) );
  NOR2_X4 u5_mult_82_U12917 ( .A1(u5_mult_82_net64881), .A2(
        u5_mult_82_net65279), .ZN(u5_mult_82_ab_47__34_) );
  NOR2_X4 u5_mult_82_U12916 ( .A1(u5_mult_82_net64935), .A2(
        u5_mult_82_net65279), .ZN(u5_mult_82_ab_47__37_) );
  INV_X4 u5_mult_82_U12915 ( .A(fracta_mul[47]), .ZN(u5_mult_82_net57182) );
  NOR2_X4 u5_mult_82_U12914 ( .A1(u5_mult_82_n6952), .A2(u5_mult_82_n6743), 
        .ZN(u5_mult_82_ab_46__3_) );
  NOR2_X4 u5_mult_82_U12913 ( .A1(u5_mult_82_n6946), .A2(u5_mult_82_n6742), 
        .ZN(u5_mult_82_ab_46__4_) );
  NOR2_X4 u5_mult_82_U12912 ( .A1(u5_mult_82_net64361), .A2(u5_mult_82_n6742), 
        .ZN(u5_mult_82_ab_46__5_) );
  NOR2_X4 u5_mult_82_U12911 ( .A1(u5_mult_82_net64379), .A2(u5_mult_82_n6742), 
        .ZN(u5_mult_82_ab_46__6_) );
  NOR2_X4 u5_mult_82_U12910 ( .A1(u5_mult_82_n6940), .A2(u5_mult_82_n6742), 
        .ZN(u5_mult_82_ab_46__7_) );
  NOR2_X4 u5_mult_82_U12909 ( .A1(u5_mult_82_net64415), .A2(u5_mult_82_n6742), 
        .ZN(u5_mult_82_ab_46__8_) );
  NOR2_X4 u5_mult_82_U12908 ( .A1(u5_mult_82_net64433), .A2(u5_mult_82_n6742), 
        .ZN(u5_mult_82_ab_46__9_) );
  NOR2_X4 u5_mult_82_U12907 ( .A1(u5_mult_82_net64455), .A2(u5_mult_82_n6742), 
        .ZN(u5_mult_82_ab_46__10_) );
  NOR2_X4 u5_mult_82_U12906 ( .A1(u5_mult_82_net64487), .A2(u5_mult_82_n6742), 
        .ZN(u5_mult_82_ab_46__12_) );
  NOR2_X4 u5_mult_82_U12905 ( .A1(u5_mult_82_net64505), .A2(u5_mult_82_n6742), 
        .ZN(u5_mult_82_ab_46__13_) );
  NOR2_X4 u5_mult_82_U12904 ( .A1(u5_mult_82_n6927), .A2(u5_mult_82_n6741), 
        .ZN(u5_mult_82_ab_46__17_) );
  NOR2_X4 u5_mult_82_U12903 ( .A1(u5_mult_82_n6919), .A2(u5_mult_82_n6741), 
        .ZN(u5_mult_82_ab_46__18_) );
  NOR2_X4 u5_mult_82_U12902 ( .A1(u5_mult_82_n6912), .A2(u5_mult_82_n6741), 
        .ZN(u5_mult_82_ab_46__19_) );
  NOR2_X4 u5_mult_82_U12901 ( .A1(u5_mult_82_net64683), .A2(u5_mult_82_n6741), 
        .ZN(u5_mult_82_ab_46__23_) );
  NOR2_X4 u5_mult_82_U12900 ( .A1(u5_mult_82_n6884), .A2(u5_mult_82_n6741), 
        .ZN(u5_mult_82_ab_46__25_) );
  NOR2_X4 u5_mult_82_U12899 ( .A1(u5_mult_82_n6879), .A2(u5_mult_82_n6741), 
        .ZN(u5_mult_82_ab_46__26_) );
  NOR2_X4 u5_mult_82_U12898 ( .A1(u5_mult_82_n6874), .A2(u5_mult_82_n6741), 
        .ZN(u5_mult_82_ab_46__27_) );
  NOR2_X4 u5_mult_82_U12897 ( .A1(u5_mult_82_n6867), .A2(u5_mult_82_n6742), 
        .ZN(u5_mult_82_ab_46__28_) );
  NOR2_X4 u5_mult_82_U12896 ( .A1(u5_mult_82_n6856), .A2(u5_mult_82_n6741), 
        .ZN(u5_mult_82_ab_46__30_) );
  NOR2_X4 u5_mult_82_U12895 ( .A1(u5_mult_82_n6849), .A2(u5_mult_82_n6741), 
        .ZN(u5_mult_82_ab_46__31_) );
  NOR2_X4 u5_mult_82_U12894 ( .A1(u5_mult_82_n6842), .A2(u5_mult_82_n6742), 
        .ZN(u5_mult_82_ab_46__32_) );
  NOR2_X4 u5_mult_82_U12893 ( .A1(u5_mult_82_n6960), .A2(u5_mult_82_net65321), 
        .ZN(u5_mult_82_ab_45__2_) );
  NOR2_X4 u5_mult_82_U12892 ( .A1(u5_mult_82_n6952), .A2(u5_mult_82_net65321), 
        .ZN(u5_mult_82_ab_45__3_) );
  NOR2_X4 u5_mult_82_U12891 ( .A1(u5_mult_82_net64361), .A2(
        u5_mult_82_net65319), .ZN(u5_mult_82_ab_45__5_) );
  NOR2_X4 u5_mult_82_U12890 ( .A1(u5_mult_82_net64379), .A2(
        u5_mult_82_net65319), .ZN(u5_mult_82_ab_45__6_) );
  NOR2_X4 u5_mult_82_U12889 ( .A1(u5_mult_82_n6940), .A2(u5_mult_82_net65319), 
        .ZN(u5_mult_82_ab_45__7_) );
  NOR2_X4 u5_mult_82_U12888 ( .A1(u5_mult_82_net64455), .A2(
        u5_mult_82_net65319), .ZN(u5_mult_82_ab_45__10_) );
  NOR2_X4 u5_mult_82_U12887 ( .A1(u5_mult_82_net64469), .A2(
        u5_mult_82_net65319), .ZN(u5_mult_82_ab_45__11_) );
  NOR2_X4 u5_mult_82_U12886 ( .A1(u5_mult_82_net64487), .A2(
        u5_mult_82_net65319), .ZN(u5_mult_82_ab_45__12_) );
  NOR2_X4 u5_mult_82_U12885 ( .A1(u5_mult_82_net64505), .A2(
        u5_mult_82_net65319), .ZN(u5_mult_82_ab_45__13_) );
  NOR2_X4 u5_mult_82_U12884 ( .A1(u5_mult_82_net64523), .A2(
        u5_mult_82_net65319), .ZN(u5_mult_82_ab_45__14_) );
  NOR2_X4 u5_mult_82_U12883 ( .A1(u5_mult_82_n6933), .A2(u5_mult_82_net65319), 
        .ZN(u5_mult_82_ab_45__15_) );
  NOR2_X4 u5_mult_82_U12882 ( .A1(u5_mult_82_n6903), .A2(u5_mult_82_net65321), 
        .ZN(u5_mult_82_ab_45__20_) );
  NOR2_X4 u5_mult_82_U12881 ( .A1(u5_mult_82_n6891), .A2(u5_mult_82_net65321), 
        .ZN(u5_mult_82_ab_45__24_) );
  NOR2_X4 u5_mult_82_U12880 ( .A1(u5_mult_82_n6879), .A2(u5_mult_82_net65321), 
        .ZN(u5_mult_82_ab_45__26_) );
  NOR2_X4 u5_mult_82_U12879 ( .A1(u5_mult_82_n6874), .A2(u5_mult_82_net65321), 
        .ZN(u5_mult_82_ab_45__27_) );
  NOR2_X4 u5_mult_82_U12878 ( .A1(u5_mult_82_n6867), .A2(u5_mult_82_net65315), 
        .ZN(u5_mult_82_ab_45__28_) );
  NOR2_X4 u5_mult_82_U12877 ( .A1(u5_mult_82_n6861), .A2(u5_mult_82_net65315), 
        .ZN(u5_mult_82_ab_45__29_) );
  NOR2_X4 u5_mult_82_U12876 ( .A1(u5_mult_82_n6856), .A2(u5_mult_82_net65315), 
        .ZN(u5_mult_82_ab_45__30_) );
  NOR2_X4 u5_mult_82_U12875 ( .A1(u5_mult_82_n6842), .A2(u5_mult_82_net65315), 
        .ZN(u5_mult_82_ab_45__32_) );
  NOR2_X4 u5_mult_82_U12874 ( .A1(u5_mult_82_n6837), .A2(u5_mult_82_net65315), 
        .ZN(u5_mult_82_ab_45__33_) );
  NOR2_X4 u5_mult_82_U12873 ( .A1(u5_mult_82_net64881), .A2(
        u5_mult_82_net65315), .ZN(u5_mult_82_ab_45__34_) );
  NOR2_X4 u5_mult_82_U12872 ( .A1(u5_mult_82_net64913), .A2(
        u5_mult_82_net65315), .ZN(u5_mult_82_ab_45__35_) );
  NOR2_X4 u5_mult_82_U12871 ( .A1(u5_mult_82_n6946), .A2(u5_mult_82_n6736), 
        .ZN(u5_mult_82_ab_44__4_) );
  NOR2_X4 u5_mult_82_U12870 ( .A1(u5_mult_82_net64379), .A2(u5_mult_82_n6736), 
        .ZN(u5_mult_82_ab_44__6_) );
  NOR2_X4 u5_mult_82_U12869 ( .A1(u5_mult_82_net64415), .A2(u5_mult_82_n6736), 
        .ZN(u5_mult_82_ab_44__8_) );
  NOR2_X4 u5_mult_82_U12868 ( .A1(u5_mult_82_net64433), .A2(u5_mult_82_n6736), 
        .ZN(u5_mult_82_ab_44__9_) );
  NOR2_X4 u5_mult_82_U12867 ( .A1(u5_mult_82_net64455), .A2(u5_mult_82_n6736), 
        .ZN(u5_mult_82_ab_44__10_) );
  NOR2_X4 u5_mult_82_U12866 ( .A1(u5_mult_82_net64487), .A2(u5_mult_82_n6736), 
        .ZN(u5_mult_82_ab_44__12_) );
  NOR2_X4 u5_mult_82_U12865 ( .A1(u5_mult_82_net64559), .A2(u5_mult_82_n6735), 
        .ZN(u5_mult_82_ab_44__16_) );
  NOR2_X4 u5_mult_82_U12864 ( .A1(u5_mult_82_n6919), .A2(u5_mult_82_n6735), 
        .ZN(u5_mult_82_ab_44__18_) );
  NOR2_X4 u5_mult_82_U12863 ( .A1(u5_mult_82_n6895), .A2(u5_mult_82_n6735), 
        .ZN(u5_mult_82_ab_44__21_) );
  NOR2_X4 u5_mult_82_U12862 ( .A1(u5_mult_82_n6849), .A2(u5_mult_82_n6734), 
        .ZN(u5_mult_82_ab_44__31_) );
  NOR2_X4 u5_mult_82_U12861 ( .A1(u5_mult_82_n6842), .A2(u5_mult_82_n6734), 
        .ZN(u5_mult_82_ab_44__32_) );
  NOR2_X4 u5_mult_82_U12860 ( .A1(u5_mult_82_n6816), .A2(u5_mult_82_n6736), 
        .ZN(u5_mult_82_ab_44__42_) );
  NOR2_X4 u5_mult_82_U12859 ( .A1(u5_mult_82_n6810), .A2(u5_mult_82_n6735), 
        .ZN(u5_mult_82_ab_44__43_) );
  NOR2_X4 u5_mult_82_U12858 ( .A1(u5_mult_82_n6803), .A2(u5_mult_82_n6736), 
        .ZN(u5_mult_82_ab_44__44_) );
  NOR2_X4 u5_mult_82_U12857 ( .A1(u5_mult_82_net64379), .A2(
        u5_mult_82_net65355), .ZN(u5_mult_82_ab_43__6_) );
  NOR2_X4 u5_mult_82_U12856 ( .A1(u5_mult_82_n6940), .A2(u5_mult_82_net65355), 
        .ZN(u5_mult_82_ab_43__7_) );
  NOR2_X4 u5_mult_82_U12855 ( .A1(u5_mult_82_net64433), .A2(
        u5_mult_82_net65355), .ZN(u5_mult_82_ab_43__9_) );
  NOR2_X4 u5_mult_82_U12854 ( .A1(u5_mult_82_net64487), .A2(
        u5_mult_82_net65355), .ZN(u5_mult_82_ab_43__12_) );
  NOR2_X4 u5_mult_82_U12853 ( .A1(u5_mult_82_net64505), .A2(
        u5_mult_82_net65355), .ZN(u5_mult_82_ab_43__13_) );
  NOR2_X4 u5_mult_82_U12852 ( .A1(u5_mult_82_net64523), .A2(
        u5_mult_82_net65355), .ZN(u5_mult_82_ab_43__14_) );
  NOR2_X4 u5_mult_82_U12851 ( .A1(u5_mult_82_n6919), .A2(u5_mult_82_net65353), 
        .ZN(u5_mult_82_ab_43__18_) );
  NOR2_X4 u5_mult_82_U12850 ( .A1(u5_mult_82_n6912), .A2(u5_mult_82_net65353), 
        .ZN(u5_mult_82_ab_43__19_) );
  NOR2_X4 u5_mult_82_U12849 ( .A1(u5_mult_82_n6903), .A2(u5_mult_82_net65353), 
        .ZN(u5_mult_82_ab_43__20_) );
  NOR2_X4 u5_mult_82_U12848 ( .A1(u5_mult_82_n6895), .A2(u5_mult_82_net65353), 
        .ZN(u5_mult_82_ab_43__21_) );
  NOR2_X4 u5_mult_82_U12847 ( .A1(u5_mult_82_n6837), .A2(u5_mult_82_net65351), 
        .ZN(u5_mult_82_ab_43__33_) );
  NOR2_X4 u5_mult_82_U12846 ( .A1(u5_mult_82_n6826), .A2(u5_mult_82_net65349), 
        .ZN(u5_mult_82_ab_43__40_) );
  NOR2_X4 u5_mult_82_U12845 ( .A1(u5_mult_82_n6810), .A2(u5_mult_82_net65349), 
        .ZN(u5_mult_82_ab_43__43_) );
  NOR2_X4 u5_mult_82_U12844 ( .A1(u5_mult_82_n6803), .A2(u5_mult_82_net65349), 
        .ZN(u5_mult_82_ab_43__44_) );
  NOR2_X4 u5_mult_82_U12843 ( .A1(u5_mult_82_n6967), .A2(u5_mult_82_net65375), 
        .ZN(u5_mult_82_ab_42__1_) );
  NOR2_X4 u5_mult_82_U12842 ( .A1(u5_mult_82_n6946), .A2(u5_mult_82_net65373), 
        .ZN(u5_mult_82_ab_42__4_) );
  NOR2_X4 u5_mult_82_U12841 ( .A1(u5_mult_82_net64379), .A2(
        u5_mult_82_net65373), .ZN(u5_mult_82_ab_42__6_) );
  NOR2_X4 u5_mult_82_U12840 ( .A1(u5_mult_82_n6940), .A2(u5_mult_82_net65373), 
        .ZN(u5_mult_82_ab_42__7_) );
  NOR2_X4 u5_mult_82_U12839 ( .A1(u5_mult_82_net64505), .A2(
        u5_mult_82_net65373), .ZN(u5_mult_82_ab_42__13_) );
  NOR2_X4 u5_mult_82_U12838 ( .A1(u5_mult_82_net64523), .A2(
        u5_mult_82_net65373), .ZN(u5_mult_82_ab_42__14_) );
  NOR2_X4 u5_mult_82_U12837 ( .A1(u5_mult_82_n6933), .A2(u5_mult_82_net65373), 
        .ZN(u5_mult_82_ab_42__15_) );
  NOR2_X4 u5_mult_82_U12836 ( .A1(u5_mult_82_n6927), .A2(u5_mult_82_net65371), 
        .ZN(u5_mult_82_ab_42__17_) );
  NOR2_X4 u5_mult_82_U12835 ( .A1(u5_mult_82_n6912), .A2(u5_mult_82_net65371), 
        .ZN(u5_mult_82_ab_42__19_) );
  NOR2_X4 u5_mult_82_U12834 ( .A1(u5_mult_82_n6895), .A2(u5_mult_82_net65371), 
        .ZN(u5_mult_82_ab_42__21_) );
  NOR2_X4 u5_mult_82_U12833 ( .A1(u5_mult_82_n6891), .A2(u5_mult_82_net65371), 
        .ZN(u5_mult_82_ab_42__24_) );
  NOR2_X4 u5_mult_82_U12832 ( .A1(u5_mult_82_n6879), .A2(u5_mult_82_net65371), 
        .ZN(u5_mult_82_ab_42__26_) );
  NOR2_X4 u5_mult_82_U12831 ( .A1(u5_mult_82_n6874), .A2(u5_mult_82_net65371), 
        .ZN(u5_mult_82_ab_42__27_) );
  NOR2_X4 u5_mult_82_U12830 ( .A1(u5_mult_82_n6861), .A2(u5_mult_82_net65369), 
        .ZN(u5_mult_82_ab_42__29_) );
  NOR2_X4 u5_mult_82_U12829 ( .A1(u5_mult_82_n6849), .A2(u5_mult_82_net65369), 
        .ZN(u5_mult_82_ab_42__31_) );
  NOR2_X4 u5_mult_82_U12828 ( .A1(u5_mult_82_n6837), .A2(u5_mult_82_net65369), 
        .ZN(u5_mult_82_ab_42__33_) );
  NOR2_X4 u5_mult_82_U12827 ( .A1(u5_mult_82_n6784), .A2(u5_mult_82_n1321), 
        .ZN(u5_mult_82_ab_42__47_) );
  NOR2_X4 u5_mult_82_U12826 ( .A1(u5_mult_82_n6960), .A2(u5_mult_82_net65393), 
        .ZN(u5_mult_82_ab_41__2_) );
  NOR2_X4 u5_mult_82_U12825 ( .A1(u5_mult_82_n6946), .A2(u5_mult_82_net65391), 
        .ZN(u5_mult_82_ab_41__4_) );
  NOR2_X4 u5_mult_82_U12824 ( .A1(u5_mult_82_net64361), .A2(
        u5_mult_82_net65391), .ZN(u5_mult_82_ab_41__5_) );
  NOR2_X4 u5_mult_82_U12823 ( .A1(u5_mult_82_n6940), .A2(u5_mult_82_net65391), 
        .ZN(u5_mult_82_ab_41__7_) );
  NOR2_X4 u5_mult_82_U12822 ( .A1(u5_mult_82_net64415), .A2(
        u5_mult_82_net65391), .ZN(u5_mult_82_ab_41__8_) );
  NOR2_X4 u5_mult_82_U12821 ( .A1(u5_mult_82_net64451), .A2(
        u5_mult_82_net65391), .ZN(u5_mult_82_ab_41__10_) );
  NOR2_X4 u5_mult_82_U12820 ( .A1(u5_mult_82_net64523), .A2(
        u5_mult_82_net65391), .ZN(u5_mult_82_ab_41__14_) );
  NOR2_X4 u5_mult_82_U12819 ( .A1(u5_mult_82_n6933), .A2(u5_mult_82_net65391), 
        .ZN(u5_mult_82_ab_41__15_) );
  NOR2_X4 u5_mult_82_U12818 ( .A1(u5_mult_82_n6927), .A2(u5_mult_82_net65389), 
        .ZN(u5_mult_82_ab_41__17_) );
  NOR2_X4 u5_mult_82_U12817 ( .A1(u5_mult_82_n6920), .A2(u5_mult_82_net65389), 
        .ZN(u5_mult_82_ab_41__18_) );
  NOR2_X4 u5_mult_82_U12816 ( .A1(u5_mult_82_n6913), .A2(u5_mult_82_net65389), 
        .ZN(u5_mult_82_ab_41__19_) );
  NOR2_X4 u5_mult_82_U12815 ( .A1(u5_mult_82_net64667), .A2(
        u5_mult_82_net65389), .ZN(u5_mult_82_ab_41__22_) );
  NOR2_X4 u5_mult_82_U12814 ( .A1(u5_mult_82_net64685), .A2(
        u5_mult_82_net65389), .ZN(u5_mult_82_ab_41__23_) );
  NOR2_X4 u5_mult_82_U12813 ( .A1(u5_mult_82_n6885), .A2(u5_mult_82_net65389), 
        .ZN(u5_mult_82_ab_41__25_) );
  NOR2_X4 u5_mult_82_U12812 ( .A1(u5_mult_82_n6880), .A2(u5_mult_82_net65389), 
        .ZN(u5_mult_82_ab_41__26_) );
  NOR2_X4 u5_mult_82_U12811 ( .A1(u5_mult_82_n6875), .A2(u5_mult_82_net65389), 
        .ZN(u5_mult_82_ab_41__27_) );
  NOR2_X4 u5_mult_82_U12810 ( .A1(u5_mult_82_n6868), .A2(u5_mult_82_net65387), 
        .ZN(u5_mult_82_ab_41__28_) );
  NOR2_X4 u5_mult_82_U12809 ( .A1(u5_mult_82_n6857), .A2(u5_mult_82_net65387), 
        .ZN(u5_mult_82_ab_41__30_) );
  NOR2_X4 u5_mult_82_U12808 ( .A1(u5_mult_82_n6843), .A2(u5_mult_82_net65387), 
        .ZN(u5_mult_82_ab_41__32_) );
  NOR2_X4 u5_mult_82_U12807 ( .A1(u5_mult_82_net64883), .A2(
        u5_mult_82_net65387), .ZN(u5_mult_82_ab_41__34_) );
  NOR2_X4 u5_mult_82_U12806 ( .A1(u5_mult_82_net64937), .A2(
        u5_mult_82_net65387), .ZN(u5_mult_82_ab_41__37_) );
  NOR2_X4 u5_mult_82_U12805 ( .A1(u5_mult_82_net64957), .A2(
        u5_mult_82_net65387), .ZN(u5_mult_82_ab_41__38_) );
  NOR2_X4 u5_mult_82_U12804 ( .A1(u5_mult_82_n6968), .A2(u5_mult_82_net65411), 
        .ZN(u5_mult_82_ab_40__1_) );
  NOR2_X4 u5_mult_82_U12803 ( .A1(u5_mult_82_n6954), .A2(u5_mult_82_net65411), 
        .ZN(u5_mult_82_ab_40__3_) );
  NOR2_X4 u5_mult_82_U12802 ( .A1(u5_mult_82_net64435), .A2(
        u5_mult_82_net65409), .ZN(u5_mult_82_ab_40__9_) );
  NOR2_X4 u5_mult_82_U12801 ( .A1(u5_mult_82_net64471), .A2(
        u5_mult_82_net65409), .ZN(u5_mult_82_ab_40__11_) );
  NOR2_X4 u5_mult_82_U12800 ( .A1(u5_mult_82_net64507), .A2(
        u5_mult_82_net65409), .ZN(u5_mult_82_ab_40__13_) );
  NOR2_X4 u5_mult_82_U12799 ( .A1(u5_mult_82_net64525), .A2(
        u5_mult_82_net65409), .ZN(u5_mult_82_ab_40__14_) );
  NOR2_X4 u5_mult_82_U12798 ( .A1(u5_mult_82_n6934), .A2(u5_mult_82_net65409), 
        .ZN(u5_mult_82_ab_40__15_) );
  NOR2_X4 u5_mult_82_U12797 ( .A1(u5_mult_82_net64561), .A2(
        u5_mult_82_net65407), .ZN(u5_mult_82_ab_40__16_) );
  NOR2_X4 u5_mult_82_U12796 ( .A1(u5_mult_82_n6928), .A2(u5_mult_82_net65407), 
        .ZN(u5_mult_82_ab_40__17_) );
  NOR2_X4 u5_mult_82_U12795 ( .A1(u5_mult_82_n6914), .A2(u5_mult_82_net65407), 
        .ZN(u5_mult_82_ab_40__19_) );
  NOR2_X4 u5_mult_82_U12794 ( .A1(u5_mult_82_n6905), .A2(u5_mult_82_net65407), 
        .ZN(u5_mult_82_ab_40__20_) );
  NOR2_X4 u5_mult_82_U12793 ( .A1(u5_mult_82_net64687), .A2(
        u5_mult_82_net65407), .ZN(u5_mult_82_ab_40__23_) );
  NOR2_X4 u5_mult_82_U12792 ( .A1(u5_mult_82_n6892), .A2(u5_mult_82_net65407), 
        .ZN(u5_mult_82_ab_40__24_) );
  NOR2_X4 u5_mult_82_U12791 ( .A1(u5_mult_82_n6886), .A2(u5_mult_82_net65407), 
        .ZN(u5_mult_82_ab_40__25_) );
  NOR2_X4 u5_mult_82_U12790 ( .A1(u5_mult_82_n6876), .A2(u5_mult_82_net65407), 
        .ZN(u5_mult_82_ab_40__27_) );
  NOR2_X4 u5_mult_82_U12789 ( .A1(u5_mult_82_n6858), .A2(u5_mult_82_net65405), 
        .ZN(u5_mult_82_ab_40__30_) );
  NOR2_X4 u5_mult_82_U12788 ( .A1(u5_mult_82_n6844), .A2(u5_mult_82_net65405), 
        .ZN(u5_mult_82_ab_40__32_) );
  NOR2_X4 u5_mult_82_U12787 ( .A1(u5_mult_82_net64885), .A2(
        u5_mult_82_net65405), .ZN(u5_mult_82_ab_40__34_) );
  NOR2_X4 u5_mult_82_U12786 ( .A1(u5_mult_82_n6828), .A2(u5_mult_82_net65403), 
        .ZN(u5_mult_82_ab_40__40_) );
  NOR2_X4 u5_mult_82_U12785 ( .A1(u5_mult_82_n6967), .A2(u5_mult_82_n6730), 
        .ZN(u5_mult_82_ab_39__1_) );
  NOR2_X4 u5_mult_82_U12784 ( .A1(u5_mult_82_net64379), .A2(u5_mult_82_n6729), 
        .ZN(u5_mult_82_ab_39__6_) );
  NOR2_X4 u5_mult_82_U12783 ( .A1(u5_mult_82_n6940), .A2(u5_mult_82_n6729), 
        .ZN(u5_mult_82_ab_39__7_) );
  NOR2_X4 u5_mult_82_U12782 ( .A1(u5_mult_82_net64415), .A2(u5_mult_82_n6729), 
        .ZN(u5_mult_82_ab_39__8_) );
  NOR2_X4 u5_mult_82_U12781 ( .A1(u5_mult_82_net64433), .A2(u5_mult_82_n6729), 
        .ZN(u5_mult_82_ab_39__9_) );
  NOR2_X4 u5_mult_82_U12780 ( .A1(u5_mult_82_net64469), .A2(u5_mult_82_n6729), 
        .ZN(u5_mult_82_ab_39__11_) );
  NOR2_X4 u5_mult_82_U12779 ( .A1(u5_mult_82_net64487), .A2(u5_mult_82_n6729), 
        .ZN(u5_mult_82_ab_39__12_) );
  NOR2_X4 u5_mult_82_U12778 ( .A1(u5_mult_82_net64523), .A2(u5_mult_82_n6729), 
        .ZN(u5_mult_82_ab_39__14_) );
  NOR2_X4 u5_mult_82_U12777 ( .A1(u5_mult_82_n6933), .A2(u5_mult_82_n6729), 
        .ZN(u5_mult_82_ab_39__15_) );
  NOR2_X4 u5_mult_82_U12776 ( .A1(u5_mult_82_net64559), .A2(u5_mult_82_n6728), 
        .ZN(u5_mult_82_ab_39__16_) );
  NOR2_X4 u5_mult_82_U12775 ( .A1(u5_mult_82_n6927), .A2(u5_mult_82_n6728), 
        .ZN(u5_mult_82_ab_39__17_) );
  NOR2_X4 u5_mult_82_U12774 ( .A1(u5_mult_82_n6920), .A2(u5_mult_82_n6728), 
        .ZN(u5_mult_82_ab_39__18_) );
  NOR2_X4 u5_mult_82_U12773 ( .A1(u5_mult_82_n6913), .A2(u5_mult_82_n6728), 
        .ZN(u5_mult_82_ab_39__19_) );
  NOR2_X4 u5_mult_82_U12772 ( .A1(u5_mult_82_n6891), .A2(u5_mult_82_n6728), 
        .ZN(u5_mult_82_ab_39__24_) );
  NOR2_X4 u5_mult_82_U12771 ( .A1(u5_mult_82_n6880), .A2(u5_mult_82_n6728), 
        .ZN(u5_mult_82_ab_39__26_) );
  NOR2_X4 u5_mult_82_U12770 ( .A1(u5_mult_82_n6862), .A2(u5_mult_82_n6727), 
        .ZN(u5_mult_82_ab_39__29_) );
  NOR2_X4 u5_mult_82_U12769 ( .A1(u5_mult_82_n6857), .A2(u5_mult_82_n6727), 
        .ZN(u5_mult_82_ab_39__30_) );
  NOR2_X4 u5_mult_82_U12768 ( .A1(u5_mult_82_n6850), .A2(u5_mult_82_n6727), 
        .ZN(u5_mult_82_ab_39__31_) );
  NOR2_X4 u5_mult_82_U12767 ( .A1(u5_mult_82_n6838), .A2(u5_mult_82_n6727), 
        .ZN(u5_mult_82_ab_39__33_) );
  NOR2_X4 u5_mult_82_U12766 ( .A1(u5_mult_82_net64883), .A2(u5_mult_82_n6727), 
        .ZN(u5_mult_82_ab_39__34_) );
  NOR2_X4 u5_mult_82_U12765 ( .A1(u5_mult_82_net64901), .A2(u5_mult_82_n6727), 
        .ZN(u5_mult_82_ab_39__35_) );
  NOR2_X4 u5_mult_82_U12764 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6727), 
        .ZN(u5_mult_82_ab_39__36_) );
  NOR2_X4 u5_mult_82_U12763 ( .A1(u5_mult_82_n6773), .A2(u5_mult_82_n6727), 
        .ZN(u5_mult_82_ab_39__49_) );
  NOR2_X4 u5_mult_82_U12762 ( .A1(u5_mult_82_n6767), .A2(u5_mult_82_n6726), 
        .ZN(u5_mult_82_ab_39__50_) );
  NOR2_X4 u5_mult_82_U12761 ( .A1(u5_mult_82_n6967), .A2(u5_mult_82_net65447), 
        .ZN(u5_mult_82_ab_38__1_) );
  NOR2_X4 u5_mult_82_U12760 ( .A1(u5_mult_82_n6960), .A2(u5_mult_82_net65447), 
        .ZN(u5_mult_82_ab_38__2_) );
  NOR2_X4 u5_mult_82_U12759 ( .A1(u5_mult_82_n6940), .A2(u5_mult_82_net65445), 
        .ZN(u5_mult_82_ab_38__7_) );
  NOR2_X4 u5_mult_82_U12758 ( .A1(u5_mult_82_net64415), .A2(
        u5_mult_82_net65445), .ZN(u5_mult_82_ab_38__8_) );
  NOR2_X4 u5_mult_82_U12757 ( .A1(u5_mult_82_net64433), .A2(
        u5_mult_82_net65445), .ZN(u5_mult_82_ab_38__9_) );
  NOR2_X4 u5_mult_82_U12756 ( .A1(u5_mult_82_net64451), .A2(
        u5_mult_82_net65445), .ZN(u5_mult_82_ab_38__10_) );
  NOR2_X4 u5_mult_82_U12755 ( .A1(u5_mult_82_net64487), .A2(
        u5_mult_82_net65445), .ZN(u5_mult_82_ab_38__12_) );
  NOR2_X4 u5_mult_82_U12754 ( .A1(u5_mult_82_net64505), .A2(
        u5_mult_82_net65445), .ZN(u5_mult_82_ab_38__13_) );
  NOR2_X4 u5_mult_82_U12753 ( .A1(u5_mult_82_n6933), .A2(u5_mult_82_net65445), 
        .ZN(u5_mult_82_ab_38__15_) );
  NOR2_X4 u5_mult_82_U12752 ( .A1(u5_mult_82_n6927), .A2(u5_mult_82_net65443), 
        .ZN(u5_mult_82_ab_38__17_) );
  NOR2_X4 u5_mult_82_U12751 ( .A1(u5_mult_82_n6920), .A2(u5_mult_82_net65443), 
        .ZN(u5_mult_82_ab_38__18_) );
  NOR2_X4 u5_mult_82_U12750 ( .A1(u5_mult_82_n6904), .A2(u5_mult_82_net65443), 
        .ZN(u5_mult_82_ab_38__20_) );
  NOR2_X4 u5_mult_82_U12749 ( .A1(u5_mult_82_n6868), .A2(u5_mult_82_net65441), 
        .ZN(u5_mult_82_ab_38__28_) );
  NOR2_X4 u5_mult_82_U12748 ( .A1(u5_mult_82_n6857), .A2(u5_mult_82_net65441), 
        .ZN(u5_mult_82_ab_38__30_) );
  NOR2_X4 u5_mult_82_U12747 ( .A1(u5_mult_82_n6850), .A2(u5_mult_82_net65441), 
        .ZN(u5_mult_82_ab_38__31_) );
  NOR2_X4 u5_mult_82_U12746 ( .A1(u5_mult_82_n6843), .A2(u5_mult_82_net65441), 
        .ZN(u5_mult_82_ab_38__32_) );
  NOR2_X4 u5_mult_82_U12745 ( .A1(u5_mult_82_n6838), .A2(u5_mult_82_net65441), 
        .ZN(u5_mult_82_ab_38__33_) );
  NOR2_X4 u5_mult_82_U12744 ( .A1(u5_mult_82_net64901), .A2(
        u5_mult_82_net65441), .ZN(u5_mult_82_ab_38__35_) );
  NOR2_X4 u5_mult_82_U12743 ( .A1(u5_mult_82_net64937), .A2(
        u5_mult_82_net65441), .ZN(u5_mult_82_ab_38__37_) );
  NOR2_X4 u5_mult_82_U12742 ( .A1(u5_mult_82_n6832), .A2(u5_mult_82_net65441), 
        .ZN(u5_mult_82_ab_38__39_) );
  NOR2_X4 u5_mult_82_U12741 ( .A1(u5_mult_82_n6953), .A2(u5_mult_82_n6723), 
        .ZN(u5_mult_82_ab_37__3_) );
  NOR2_X4 u5_mult_82_U12740 ( .A1(u5_mult_82_net64451), .A2(u5_mult_82_n6722), 
        .ZN(u5_mult_82_ab_37__10_) );
  NOR2_X4 u5_mult_82_U12739 ( .A1(u5_mult_82_net64523), .A2(u5_mult_82_n6722), 
        .ZN(u5_mult_82_ab_37__14_) );
  NOR2_X4 u5_mult_82_U12738 ( .A1(u5_mult_82_n6933), .A2(u5_mult_82_n6722), 
        .ZN(u5_mult_82_ab_37__15_) );
  NOR2_X4 u5_mult_82_U12737 ( .A1(u5_mult_82_n6927), .A2(u5_mult_82_n6721), 
        .ZN(u5_mult_82_ab_37__17_) );
  NOR2_X4 u5_mult_82_U12736 ( .A1(u5_mult_82_net64685), .A2(u5_mult_82_n6721), 
        .ZN(u5_mult_82_ab_37__23_) );
  NOR2_X4 u5_mult_82_U12735 ( .A1(u5_mult_82_n6862), .A2(u5_mult_82_n6720), 
        .ZN(u5_mult_82_ab_37__29_) );
  NOR2_X4 u5_mult_82_U12734 ( .A1(u5_mult_82_n6850), .A2(u5_mult_82_n6720), 
        .ZN(u5_mult_82_ab_37__31_) );
  NOR2_X4 u5_mult_82_U12733 ( .A1(u5_mult_82_n6838), .A2(u5_mult_82_n6720), 
        .ZN(u5_mult_82_ab_37__33_) );
  NOR2_X4 u5_mult_82_U12732 ( .A1(u5_mult_82_net64883), .A2(u5_mult_82_n6720), 
        .ZN(u5_mult_82_ab_37__34_) );
  NOR2_X4 u5_mult_82_U12731 ( .A1(u5_mult_82_net64901), .A2(u5_mult_82_n6720), 
        .ZN(u5_mult_82_ab_37__35_) );
  NOR2_X4 u5_mult_82_U12730 ( .A1(u5_mult_82_n6827), .A2(u5_mult_82_n6721), 
        .ZN(u5_mult_82_ab_37__40_) );
  NOR2_X4 u5_mult_82_U12729 ( .A1(u5_mult_82_n6811), .A2(u5_mult_82_n6721), 
        .ZN(u5_mult_82_ab_37__43_) );
  NOR2_X4 u5_mult_82_U12728 ( .A1(u5_mult_82_n6804), .A2(u5_mult_82_n6721), 
        .ZN(u5_mult_82_ab_37__44_) );
  NOR2_X4 u5_mult_82_U12727 ( .A1(u5_mult_82_n6784), .A2(u5_mult_82_n6722), 
        .ZN(u5_mult_82_ab_37__47_) );
  NOR2_X4 u5_mult_82_U12726 ( .A1(u5_mult_82_net64415), .A2(u5_mult_82_n6716), 
        .ZN(u5_mult_82_ab_36__8_) );
  NOR2_X4 u5_mult_82_U12725 ( .A1(u5_mult_82_net64469), .A2(u5_mult_82_n6716), 
        .ZN(u5_mult_82_ab_36__11_) );
  NOR2_X4 u5_mult_82_U12724 ( .A1(u5_mult_82_n6933), .A2(u5_mult_82_n6716), 
        .ZN(u5_mult_82_ab_36__15_) );
  NOR2_X4 u5_mult_82_U12723 ( .A1(u5_mult_82_net64559), .A2(u5_mult_82_n6715), 
        .ZN(u5_mult_82_ab_36__16_) );
  NOR2_X4 u5_mult_82_U12722 ( .A1(u5_mult_82_n6920), .A2(u5_mult_82_n6715), 
        .ZN(u5_mult_82_ab_36__18_) );
  NOR2_X4 u5_mult_82_U12721 ( .A1(u5_mult_82_net64667), .A2(u5_mult_82_n6715), 
        .ZN(u5_mult_82_ab_36__22_) );
  NOR2_X4 u5_mult_82_U12720 ( .A1(u5_mult_82_net64685), .A2(u5_mult_82_n6715), 
        .ZN(u5_mult_82_ab_36__23_) );
  NOR2_X4 u5_mult_82_U12719 ( .A1(u5_mult_82_n6891), .A2(u5_mult_82_n6715), 
        .ZN(u5_mult_82_ab_36__24_) );
  NOR2_X4 u5_mult_82_U12718 ( .A1(u5_mult_82_n6880), .A2(u5_mult_82_n6715), 
        .ZN(u5_mult_82_ab_36__26_) );
  NOR2_X4 u5_mult_82_U12717 ( .A1(u5_mult_82_n6862), .A2(u5_mult_82_n6714), 
        .ZN(u5_mult_82_ab_36__29_) );
  NOR2_X4 u5_mult_82_U12716 ( .A1(u5_mult_82_n6850), .A2(u5_mult_82_n6714), 
        .ZN(u5_mult_82_ab_36__31_) );
  NOR2_X4 u5_mult_82_U12715 ( .A1(u5_mult_82_n6843), .A2(u5_mult_82_n6714), 
        .ZN(u5_mult_82_ab_36__32_) );
  NOR2_X4 u5_mult_82_U12714 ( .A1(u5_mult_82_n6838), .A2(u5_mult_82_n6714), 
        .ZN(u5_mult_82_ab_36__33_) );
  NOR2_X4 u5_mult_82_U12713 ( .A1(u5_mult_82_net64883), .A2(u5_mult_82_n6714), 
        .ZN(u5_mult_82_ab_36__34_) );
  NOR2_X4 u5_mult_82_U12712 ( .A1(u5_mult_82_net64901), .A2(u5_mult_82_n6714), 
        .ZN(u5_mult_82_ab_36__35_) );
  NOR2_X4 u5_mult_82_U12711 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6714), 
        .ZN(u5_mult_82_ab_36__36_) );
  NOR2_X4 u5_mult_82_U12710 ( .A1(u5_mult_82_n6778), .A2(u5_mult_82_n6713), 
        .ZN(u5_mult_82_ab_36__48_) );
  INV_X4 u5_mult_82_U12709 ( .A(fracta_mul[36]), .ZN(u5_mult_82_n7003) );
  NOR2_X4 u5_mult_82_U12708 ( .A1(u5_mult_82_n6946), .A2(u5_mult_82_n6709), 
        .ZN(u5_mult_82_ab_35__4_) );
  NOR2_X4 u5_mult_82_U12707 ( .A1(u5_mult_82_net64433), .A2(u5_mult_82_n6709), 
        .ZN(u5_mult_82_ab_35__9_) );
  NOR2_X4 u5_mult_82_U12706 ( .A1(u5_mult_82_net64505), .A2(u5_mult_82_n6709), 
        .ZN(u5_mult_82_ab_35__13_) );
  NOR2_X4 u5_mult_82_U12705 ( .A1(u5_mult_82_net64523), .A2(u5_mult_82_n6709), 
        .ZN(u5_mult_82_ab_35__14_) );
  NOR2_X4 u5_mult_82_U12704 ( .A1(u5_mult_82_n6913), .A2(u5_mult_82_n6708), 
        .ZN(u5_mult_82_ab_35__19_) );
  NOR2_X4 u5_mult_82_U12703 ( .A1(u5_mult_82_n6904), .A2(u5_mult_82_n6708), 
        .ZN(u5_mult_82_ab_35__20_) );
  NOR2_X4 u5_mult_82_U12702 ( .A1(u5_mult_82_n6896), .A2(u5_mult_82_n6708), 
        .ZN(u5_mult_82_ab_35__21_) );
  NOR2_X4 u5_mult_82_U12701 ( .A1(u5_mult_82_net64685), .A2(u5_mult_82_n6708), 
        .ZN(u5_mult_82_ab_35__23_) );
  NOR2_X4 u5_mult_82_U12700 ( .A1(u5_mult_82_n6885), .A2(u5_mult_82_n6708), 
        .ZN(u5_mult_82_ab_35__25_) );
  NOR2_X4 u5_mult_82_U12699 ( .A1(u5_mult_82_n6875), .A2(u5_mult_82_n6708), 
        .ZN(u5_mult_82_ab_35__27_) );
  NOR2_X4 u5_mult_82_U12698 ( .A1(u5_mult_82_n6868), .A2(u5_mult_82_n6707), 
        .ZN(u5_mult_82_ab_35__28_) );
  NOR2_X4 u5_mult_82_U12697 ( .A1(u5_mult_82_n6857), .A2(u5_mult_82_n6707), 
        .ZN(u5_mult_82_ab_35__30_) );
  NOR2_X4 u5_mult_82_U12696 ( .A1(u5_mult_82_n6850), .A2(u5_mult_82_n6707), 
        .ZN(u5_mult_82_ab_35__31_) );
  NOR2_X4 u5_mult_82_U12695 ( .A1(u5_mult_82_n6843), .A2(u5_mult_82_n6707), 
        .ZN(u5_mult_82_ab_35__32_) );
  NOR2_X4 u5_mult_82_U12694 ( .A1(u5_mult_82_net64883), .A2(u5_mult_82_n6707), 
        .ZN(u5_mult_82_ab_35__34_) );
  NOR2_X4 u5_mult_82_U12693 ( .A1(u5_mult_82_net64901), .A2(u5_mult_82_n6707), 
        .ZN(u5_mult_82_ab_35__35_) );
  NOR2_X4 u5_mult_82_U12692 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6707), 
        .ZN(u5_mult_82_ab_35__36_) );
  NOR2_X4 u5_mult_82_U12691 ( .A1(u5_mult_82_n6821), .A2(u5_mult_82_n6706), 
        .ZN(u5_mult_82_ab_35__41_) );
  NOR2_X4 u5_mult_82_U12690 ( .A1(u5_mult_82_n6816), .A2(u5_mult_82_n6706), 
        .ZN(u5_mult_82_ab_35__42_) );
  NOR2_X4 u5_mult_82_U12689 ( .A1(u5_mult_82_n6811), .A2(u5_mult_82_n6706), 
        .ZN(u5_mult_82_ab_35__43_) );
  INV_X4 u5_mult_82_U12688 ( .A(fracta_mul[35]), .ZN(u5_mult_82_n7002) );
  NOR2_X4 u5_mult_82_U12687 ( .A1(u5_mult_82_n6946), .A2(u5_mult_82_net65517), 
        .ZN(u5_mult_82_ab_34__4_) );
  NOR2_X4 u5_mult_82_U12686 ( .A1(u5_mult_82_net64361), .A2(
        u5_mult_82_net65517), .ZN(u5_mult_82_ab_34__5_) );
  NOR2_X4 u5_mult_82_U12685 ( .A1(u5_mult_82_net64379), .A2(
        u5_mult_82_net65517), .ZN(u5_mult_82_ab_34__6_) );
  NOR2_X4 u5_mult_82_U12684 ( .A1(u5_mult_82_n6940), .A2(u5_mult_82_net65517), 
        .ZN(u5_mult_82_ab_34__7_) );
  NOR2_X4 u5_mult_82_U12683 ( .A1(u5_mult_82_net64415), .A2(
        u5_mult_82_net65517), .ZN(u5_mult_82_ab_34__8_) );
  NOR2_X4 u5_mult_82_U12682 ( .A1(u5_mult_82_net64433), .A2(
        u5_mult_82_net65517), .ZN(u5_mult_82_ab_34__9_) );
  NOR2_X4 u5_mult_82_U12681 ( .A1(u5_mult_82_net64505), .A2(
        u5_mult_82_net65517), .ZN(u5_mult_82_ab_34__13_) );
  NOR2_X4 u5_mult_82_U12680 ( .A1(u5_mult_82_net64523), .A2(
        u5_mult_82_net65517), .ZN(u5_mult_82_ab_34__14_) );
  NOR2_X4 u5_mult_82_U12679 ( .A1(u5_mult_82_n6933), .A2(u5_mult_82_net65517), 
        .ZN(u5_mult_82_ab_34__15_) );
  NOR2_X4 u5_mult_82_U12678 ( .A1(u5_mult_82_n6904), .A2(u5_mult_82_net65515), 
        .ZN(u5_mult_82_ab_34__20_) );
  NOR2_X4 u5_mult_82_U12677 ( .A1(u5_mult_82_n6896), .A2(u5_mult_82_net65515), 
        .ZN(u5_mult_82_ab_34__21_) );
  NOR2_X4 u5_mult_82_U12676 ( .A1(u5_mult_82_net64667), .A2(
        u5_mult_82_net65515), .ZN(u5_mult_82_ab_34__22_) );
  NOR2_X4 u5_mult_82_U12675 ( .A1(u5_mult_82_n6885), .A2(u5_mult_82_net65515), 
        .ZN(u5_mult_82_ab_34__25_) );
  NOR2_X4 u5_mult_82_U12674 ( .A1(u5_mult_82_n6862), .A2(u5_mult_82_net65513), 
        .ZN(u5_mult_82_ab_34__29_) );
  NOR2_X4 u5_mult_82_U12673 ( .A1(u5_mult_82_n6857), .A2(u5_mult_82_net65513), 
        .ZN(u5_mult_82_ab_34__30_) );
  NOR2_X4 u5_mult_82_U12672 ( .A1(u5_mult_82_n6850), .A2(u5_mult_82_net65513), 
        .ZN(u5_mult_82_ab_34__31_) );
  NOR2_X4 u5_mult_82_U12671 ( .A1(u5_mult_82_n6843), .A2(u5_mult_82_net65513), 
        .ZN(u5_mult_82_ab_34__32_) );
  NOR2_X4 u5_mult_82_U12670 ( .A1(u5_mult_82_n6827), .A2(u5_mult_82_net65515), 
        .ZN(u5_mult_82_ab_34__40_) );
  NOR2_X4 u5_mult_82_U12669 ( .A1(u5_mult_82_n6816), .A2(u5_mult_82_net65515), 
        .ZN(u5_mult_82_ab_34__42_) );
  NOR2_X4 u5_mult_82_U12668 ( .A1(u5_mult_82_n6811), .A2(u5_mult_82_net65515), 
        .ZN(u5_mult_82_ab_34__43_) );
  NOR2_X4 u5_mult_82_U12667 ( .A1(u5_mult_82_n6946), .A2(u5_mult_82_n6701), 
        .ZN(u5_mult_82_ab_33__4_) );
  NOR2_X4 u5_mult_82_U12666 ( .A1(u5_mult_82_net64361), .A2(u5_mult_82_n6701), 
        .ZN(u5_mult_82_ab_33__5_) );
  NOR2_X4 u5_mult_82_U12665 ( .A1(u5_mult_82_n6940), .A2(u5_mult_82_n6701), 
        .ZN(u5_mult_82_ab_33__7_) );
  NOR2_X4 u5_mult_82_U12664 ( .A1(u5_mult_82_net64415), .A2(u5_mult_82_n6701), 
        .ZN(u5_mult_82_ab_33__8_) );
  NOR2_X4 u5_mult_82_U12663 ( .A1(u5_mult_82_net64433), .A2(u5_mult_82_n6701), 
        .ZN(u5_mult_82_ab_33__9_) );
  NOR2_X4 u5_mult_82_U12662 ( .A1(u5_mult_82_net64451), .A2(u5_mult_82_n6701), 
        .ZN(u5_mult_82_ab_33__10_) );
  NOR2_X4 u5_mult_82_U12661 ( .A1(u5_mult_82_net64469), .A2(u5_mult_82_n6701), 
        .ZN(u5_mult_82_ab_33__11_) );
  NOR2_X4 u5_mult_82_U12660 ( .A1(u5_mult_82_net64523), .A2(u5_mult_82_n6701), 
        .ZN(u5_mult_82_ab_33__14_) );
  NOR2_X4 u5_mult_82_U12659 ( .A1(u5_mult_82_n6913), .A2(u5_mult_82_n6700), 
        .ZN(u5_mult_82_ab_33__19_) );
  NOR2_X4 u5_mult_82_U12658 ( .A1(u5_mult_82_n6891), .A2(u5_mult_82_n6700), 
        .ZN(u5_mult_82_ab_33__24_) );
  NOR2_X4 u5_mult_82_U12657 ( .A1(u5_mult_82_n6885), .A2(u5_mult_82_n6700), 
        .ZN(u5_mult_82_ab_33__25_) );
  NOR2_X4 u5_mult_82_U12656 ( .A1(u5_mult_82_n6880), .A2(u5_mult_82_n6700), 
        .ZN(u5_mult_82_ab_33__26_) );
  NOR2_X4 u5_mult_82_U12655 ( .A1(u5_mult_82_n6857), .A2(u5_mult_82_n6699), 
        .ZN(u5_mult_82_ab_33__30_) );
  NOR2_X4 u5_mult_82_U12654 ( .A1(u5_mult_82_n6850), .A2(u5_mult_82_n6699), 
        .ZN(u5_mult_82_ab_33__31_) );
  NOR2_X4 u5_mult_82_U12653 ( .A1(u5_mult_82_n6843), .A2(u5_mult_82_n6699), 
        .ZN(u5_mult_82_ab_33__32_) );
  NOR2_X4 u5_mult_82_U12652 ( .A1(u5_mult_82_n6821), .A2(u5_mult_82_n6701), 
        .ZN(u5_mult_82_ab_33__41_) );
  NOR2_X4 u5_mult_82_U12651 ( .A1(u5_mult_82_n6816), .A2(u5_mult_82_n6701), 
        .ZN(u5_mult_82_ab_33__42_) );
  NOR2_X4 u5_mult_82_U12650 ( .A1(u5_mult_82_n6811), .A2(u5_mult_82_n6701), 
        .ZN(u5_mult_82_ab_33__43_) );
  NOR2_X4 u5_mult_82_U12649 ( .A1(u5_mult_82_n6784), .A2(u5_mult_82_n6700), 
        .ZN(u5_mult_82_ab_33__47_) );
  NOR2_X4 u5_mult_82_U12648 ( .A1(u5_mult_82_n6778), .A2(u5_mult_82_n6702), 
        .ZN(u5_mult_82_ab_33__48_) );
  NOR2_X4 u5_mult_82_U12647 ( .A1(u5_mult_82_n6982), .A2(u5_mult_82_n6696), 
        .ZN(u5_mult_82_ab_32__52_) );
  NOR2_X4 u5_mult_82_U12646 ( .A1(u5_mult_82_n6760), .A2(u5_mult_82_n6698), 
        .ZN(u5_mult_82_ab_33__51_) );
  NOR2_X4 u5_mult_82_U12645 ( .A1(u5_mult_82_net64361), .A2(u5_mult_82_n6695), 
        .ZN(u5_mult_82_ab_32__5_) );
  NOR2_X4 u5_mult_82_U12644 ( .A1(u5_mult_82_n6940), .A2(u5_mult_82_n6695), 
        .ZN(u5_mult_82_ab_32__7_) );
  NOR2_X4 u5_mult_82_U12643 ( .A1(u5_mult_82_net64469), .A2(u5_mult_82_n6695), 
        .ZN(u5_mult_82_ab_32__11_) );
  NOR2_X4 u5_mult_82_U12642 ( .A1(u5_mult_82_net64487), .A2(u5_mult_82_n6695), 
        .ZN(u5_mult_82_ab_32__12_) );
  NOR2_X4 u5_mult_82_U12641 ( .A1(u5_mult_82_n6927), .A2(u5_mult_82_n6694), 
        .ZN(u5_mult_82_ab_32__17_) );
  NOR2_X4 u5_mult_82_U12640 ( .A1(u5_mult_82_n6904), .A2(u5_mult_82_n6694), 
        .ZN(u5_mult_82_ab_32__20_) );
  NOR2_X4 u5_mult_82_U12639 ( .A1(u5_mult_82_net64667), .A2(u5_mult_82_n6694), 
        .ZN(u5_mult_82_ab_32__22_) );
  NOR2_X4 u5_mult_82_U12638 ( .A1(u5_mult_82_n6891), .A2(u5_mult_82_n6694), 
        .ZN(u5_mult_82_ab_32__24_) );
  NOR2_X4 u5_mult_82_U12637 ( .A1(u5_mult_82_n6885), .A2(u5_mult_82_n6694), 
        .ZN(u5_mult_82_ab_32__25_) );
  NOR2_X4 u5_mult_82_U12636 ( .A1(u5_mult_82_n6880), .A2(u5_mult_82_n6694), 
        .ZN(u5_mult_82_ab_32__26_) );
  NOR2_X4 u5_mult_82_U12635 ( .A1(u5_mult_82_n6875), .A2(u5_mult_82_n6694), 
        .ZN(u5_mult_82_ab_32__27_) );
  NOR2_X4 u5_mult_82_U12634 ( .A1(u5_mult_82_n6862), .A2(u5_mult_82_n6693), 
        .ZN(u5_mult_82_ab_32__29_) );
  NOR2_X4 u5_mult_82_U12633 ( .A1(u5_mult_82_n6850), .A2(u5_mult_82_n6693), 
        .ZN(u5_mult_82_ab_32__31_) );
  NOR2_X4 u5_mult_82_U12632 ( .A1(u5_mult_82_n6827), .A2(u5_mult_82_n6692), 
        .ZN(u5_mult_82_ab_32__40_) );
  NOR2_X4 u5_mult_82_U12631 ( .A1(u5_mult_82_n6821), .A2(u5_mult_82_n6692), 
        .ZN(u5_mult_82_ab_32__41_) );
  NOR2_X4 u5_mult_82_U12630 ( .A1(u5_mult_82_n6811), .A2(u5_mult_82_n6692), 
        .ZN(u5_mult_82_ab_32__43_) );
  NOR2_X4 u5_mult_82_U12629 ( .A1(u5_mult_82_n6773), .A2(u5_mult_82_n6692), 
        .ZN(u5_mult_82_ab_32__49_) );
  NOR2_X4 u5_mult_82_U12628 ( .A1(u5_mult_82_n6767), .A2(u5_mult_82_n6692), 
        .ZN(u5_mult_82_ab_32__50_) );
  NOR2_X4 u5_mult_82_U12627 ( .A1(u5_mult_82_n6982), .A2(u5_mult_82_n6687), 
        .ZN(u5_mult_82_ab_31__52_) );
  NOR2_X4 u5_mult_82_U12626 ( .A1(u5_mult_82_n6760), .A2(u5_mult_82_n6692), 
        .ZN(u5_mult_82_ab_32__51_) );
  INV_X4 u5_mult_82_U12625 ( .A(fracta_mul[32]), .ZN(u5_mult_82_n7001) );
  NOR2_X4 u5_mult_82_U12624 ( .A1(u5_mult_82_n6946), .A2(u5_mult_82_n6686), 
        .ZN(u5_mult_82_ab_31__4_) );
  NOR2_X4 u5_mult_82_U12623 ( .A1(u5_mult_82_net64415), .A2(u5_mult_82_n6686), 
        .ZN(u5_mult_82_ab_31__8_) );
  NOR2_X4 u5_mult_82_U12622 ( .A1(u5_mult_82_net64451), .A2(u5_mult_82_n6686), 
        .ZN(u5_mult_82_ab_31__10_) );
  NOR2_X4 u5_mult_82_U12621 ( .A1(u5_mult_82_net64487), .A2(u5_mult_82_n6686), 
        .ZN(u5_mult_82_ab_31__12_) );
  NOR2_X4 u5_mult_82_U12620 ( .A1(u5_mult_82_net64505), .A2(u5_mult_82_n6686), 
        .ZN(u5_mult_82_ab_31__13_) );
  NOR2_X4 u5_mult_82_U12619 ( .A1(u5_mult_82_net64523), .A2(u5_mult_82_n6686), 
        .ZN(u5_mult_82_ab_31__14_) );
  NOR2_X4 u5_mult_82_U12618 ( .A1(u5_mult_82_n6927), .A2(u5_mult_82_n6685), 
        .ZN(u5_mult_82_ab_31__17_) );
  NOR2_X4 u5_mult_82_U12617 ( .A1(u5_mult_82_n6920), .A2(u5_mult_82_n6685), 
        .ZN(u5_mult_82_ab_31__18_) );
  NOR2_X4 u5_mult_82_U12616 ( .A1(u5_mult_82_n6913), .A2(u5_mult_82_n6685), 
        .ZN(u5_mult_82_ab_31__19_) );
  NOR2_X4 u5_mult_82_U12615 ( .A1(u5_mult_82_net64667), .A2(u5_mult_82_n6685), 
        .ZN(u5_mult_82_ab_31__22_) );
  NOR2_X4 u5_mult_82_U12614 ( .A1(u5_mult_82_net64685), .A2(u5_mult_82_n6685), 
        .ZN(u5_mult_82_ab_31__23_) );
  NOR2_X4 u5_mult_82_U12613 ( .A1(u5_mult_82_n6885), .A2(u5_mult_82_n6685), 
        .ZN(u5_mult_82_ab_31__25_) );
  NOR2_X4 u5_mult_82_U12612 ( .A1(u5_mult_82_n6868), .A2(u5_mult_82_n6684), 
        .ZN(u5_mult_82_ab_31__28_) );
  NOR2_X4 u5_mult_82_U12611 ( .A1(u5_mult_82_n6857), .A2(u5_mult_82_n6684), 
        .ZN(u5_mult_82_ab_31__30_) );
  NOR2_X4 u5_mult_82_U12610 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6684), 
        .ZN(u5_mult_82_ab_31__36_) );
  NOR2_X4 u5_mult_82_U12609 ( .A1(u5_mult_82_n6791), .A2(u5_mult_82_n6685), 
        .ZN(u5_mult_82_ab_31__46_) );
  NOR2_X4 u5_mult_82_U12608 ( .A1(u5_mult_82_n6784), .A2(u5_mult_82_n6686), 
        .ZN(u5_mult_82_ab_31__47_) );
  NOR2_X4 u5_mult_82_U12607 ( .A1(u5_mult_82_net64379), .A2(u5_mult_82_n6680), 
        .ZN(u5_mult_82_ab_30__6_) );
  NOR2_X4 u5_mult_82_U12606 ( .A1(u5_mult_82_net64415), .A2(u5_mult_82_n6680), 
        .ZN(u5_mult_82_ab_30__8_) );
  NOR2_X4 u5_mult_82_U12605 ( .A1(u5_mult_82_net64469), .A2(u5_mult_82_n6680), 
        .ZN(u5_mult_82_ab_30__11_) );
  NOR2_X4 u5_mult_82_U12604 ( .A1(u5_mult_82_n6933), .A2(u5_mult_82_n6680), 
        .ZN(u5_mult_82_ab_30__15_) );
  NOR2_X4 u5_mult_82_U12603 ( .A1(u5_mult_82_net64559), .A2(u5_mult_82_n6679), 
        .ZN(u5_mult_82_ab_30__16_) );
  NOR2_X4 u5_mult_82_U12602 ( .A1(u5_mult_82_n6927), .A2(u5_mult_82_n6679), 
        .ZN(u5_mult_82_ab_30__17_) );
  NOR2_X4 u5_mult_82_U12601 ( .A1(u5_mult_82_n6920), .A2(u5_mult_82_n6679), 
        .ZN(u5_mult_82_ab_30__18_) );
  NOR2_X4 u5_mult_82_U12600 ( .A1(u5_mult_82_n6913), .A2(u5_mult_82_n6679), 
        .ZN(u5_mult_82_ab_30__19_) );
  NOR2_X4 u5_mult_82_U12599 ( .A1(u5_mult_82_n6904), .A2(u5_mult_82_n6679), 
        .ZN(u5_mult_82_ab_30__20_) );
  NOR2_X4 u5_mult_82_U12598 ( .A1(u5_mult_82_net64667), .A2(u5_mult_82_n6679), 
        .ZN(u5_mult_82_ab_30__22_) );
  NOR2_X4 u5_mult_82_U12597 ( .A1(u5_mult_82_net64685), .A2(u5_mult_82_n6679), 
        .ZN(u5_mult_82_ab_30__23_) );
  NOR2_X4 u5_mult_82_U12596 ( .A1(u5_mult_82_n6891), .A2(u5_mult_82_n6679), 
        .ZN(u5_mult_82_ab_30__24_) );
  NOR2_X4 u5_mult_82_U12595 ( .A1(u5_mult_82_n6880), .A2(u5_mult_82_n6679), 
        .ZN(u5_mult_82_ab_30__26_) );
  NOR2_X4 u5_mult_82_U12594 ( .A1(u5_mult_82_n6875), .A2(u5_mult_82_n6679), 
        .ZN(u5_mult_82_ab_30__27_) );
  NOR2_X4 u5_mult_82_U12593 ( .A1(u5_mult_82_n6862), .A2(u5_mult_82_n6678), 
        .ZN(u5_mult_82_ab_30__29_) );
  NOR2_X4 u5_mult_82_U12592 ( .A1(u5_mult_82_n6857), .A2(u5_mult_82_n6678), 
        .ZN(u5_mult_82_ab_30__30_) );
  NOR2_X4 u5_mult_82_U12591 ( .A1(u5_mult_82_n6843), .A2(u5_mult_82_n6678), 
        .ZN(u5_mult_82_ab_30__32_) );
  NOR2_X4 u5_mult_82_U12590 ( .A1(u5_mult_82_net64901), .A2(u5_mult_82_n6678), 
        .ZN(u5_mult_82_ab_30__35_) );
  NOR2_X4 u5_mult_82_U12589 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6678), 
        .ZN(u5_mult_82_ab_30__36_) );
  NOR2_X4 u5_mult_82_U12588 ( .A1(u5_mult_82_net64937), .A2(u5_mult_82_n6678), 
        .ZN(u5_mult_82_ab_30__37_) );
  NOR2_X4 u5_mult_82_U12587 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6678), 
        .ZN(u5_mult_82_ab_30__38_) );
  NOR2_X4 u5_mult_82_U12586 ( .A1(u5_mult_82_n6791), .A2(u5_mult_82_n6677), 
        .ZN(u5_mult_82_ab_30__46_) );
  NOR2_X4 u5_mult_82_U12585 ( .A1(u5_mult_82_n6784), .A2(u5_mult_82_n6677), 
        .ZN(u5_mult_82_ab_30__47_) );
  INV_X4 u5_mult_82_U12584 ( .A(fracta_mul[30]), .ZN(u5_mult_82_n7000) );
  NOR2_X4 u5_mult_82_U12583 ( .A1(u5_mult_82_net64379), .A2(u5_mult_82_n6673), 
        .ZN(u5_mult_82_ab_29__6_) );
  NOR2_X4 u5_mult_82_U12582 ( .A1(u5_mult_82_net64433), .A2(u5_mult_82_n6673), 
        .ZN(u5_mult_82_ab_29__9_) );
  NOR2_X4 u5_mult_82_U12581 ( .A1(u5_mult_82_net64451), .A2(u5_mult_82_n6673), 
        .ZN(u5_mult_82_ab_29__10_) );
  NOR2_X4 u5_mult_82_U12580 ( .A1(u5_mult_82_net64469), .A2(u5_mult_82_n6673), 
        .ZN(u5_mult_82_ab_29__11_) );
  NOR2_X4 u5_mult_82_U12579 ( .A1(u5_mult_82_net64487), .A2(u5_mult_82_n6673), 
        .ZN(u5_mult_82_ab_29__12_) );
  NOR2_X4 u5_mult_82_U12578 ( .A1(u5_mult_82_net64505), .A2(u5_mult_82_n6673), 
        .ZN(u5_mult_82_ab_29__13_) );
  NOR2_X4 u5_mult_82_U12577 ( .A1(u5_mult_82_n6933), .A2(u5_mult_82_n6673), 
        .ZN(u5_mult_82_ab_29__15_) );
  NOR2_X4 u5_mult_82_U12576 ( .A1(u5_mult_82_n6927), .A2(u5_mult_82_n6672), 
        .ZN(u5_mult_82_ab_29__17_) );
  NOR2_X4 u5_mult_82_U12575 ( .A1(u5_mult_82_n6920), .A2(u5_mult_82_n6672), 
        .ZN(u5_mult_82_ab_29__18_) );
  NOR2_X4 u5_mult_82_U12574 ( .A1(u5_mult_82_n6904), .A2(u5_mult_82_n6672), 
        .ZN(u5_mult_82_ab_29__20_) );
  NOR2_X4 u5_mult_82_U12573 ( .A1(u5_mult_82_net64685), .A2(u5_mult_82_n6672), 
        .ZN(u5_mult_82_ab_29__23_) );
  NOR2_X4 u5_mult_82_U12572 ( .A1(u5_mult_82_n6885), .A2(u5_mult_82_n6672), 
        .ZN(u5_mult_82_ab_29__25_) );
  NOR2_X4 u5_mult_82_U12571 ( .A1(u5_mult_82_n6880), .A2(u5_mult_82_n6672), 
        .ZN(u5_mult_82_ab_29__26_) );
  NOR2_X4 u5_mult_82_U12570 ( .A1(u5_mult_82_n6875), .A2(u5_mult_82_n6672), 
        .ZN(u5_mult_82_ab_29__27_) );
  NOR2_X4 u5_mult_82_U12569 ( .A1(u5_mult_82_n6868), .A2(u5_mult_82_n6671), 
        .ZN(u5_mult_82_ab_29__28_) );
  NOR2_X4 u5_mult_82_U12568 ( .A1(u5_mult_82_n6862), .A2(u5_mult_82_n6671), 
        .ZN(u5_mult_82_ab_29__29_) );
  NOR2_X4 u5_mult_82_U12567 ( .A1(u5_mult_82_n6857), .A2(u5_mult_82_n6671), 
        .ZN(u5_mult_82_ab_29__30_) );
  NOR2_X4 u5_mult_82_U12566 ( .A1(u5_mult_82_n6850), .A2(u5_mult_82_n6671), 
        .ZN(u5_mult_82_ab_29__31_) );
  NOR2_X4 u5_mult_82_U12565 ( .A1(u5_mult_82_n6843), .A2(u5_mult_82_n6671), 
        .ZN(u5_mult_82_ab_29__32_) );
  NOR2_X4 u5_mult_82_U12564 ( .A1(u5_mult_82_n6838), .A2(u5_mult_82_n6671), 
        .ZN(u5_mult_82_ab_29__33_) );
  NOR2_X4 u5_mult_82_U12563 ( .A1(u5_mult_82_net64883), .A2(u5_mult_82_n6671), 
        .ZN(u5_mult_82_ab_29__34_) );
  NOR2_X4 u5_mult_82_U12562 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6671), 
        .ZN(u5_mult_82_ab_29__36_) );
  NOR2_X4 u5_mult_82_U12561 ( .A1(u5_mult_82_net64937), .A2(u5_mult_82_n6671), 
        .ZN(u5_mult_82_ab_29__37_) );
  NOR2_X4 u5_mult_82_U12560 ( .A1(u5_mult_82_n6827), .A2(u5_mult_82_n6670), 
        .ZN(u5_mult_82_ab_29__40_) );
  NOR2_X4 u5_mult_82_U12559 ( .A1(u5_mult_82_n6821), .A2(u5_mult_82_n6670), 
        .ZN(u5_mult_82_ab_29__41_) );
  NOR2_X4 u5_mult_82_U12558 ( .A1(u5_mult_82_n6804), .A2(u5_mult_82_n6670), 
        .ZN(u5_mult_82_ab_29__44_) );
  NOR2_X4 u5_mult_82_U12557 ( .A1(u5_mult_82_n6797), .A2(u5_mult_82_n6670), 
        .ZN(u5_mult_82_ab_29__45_) );
  INV_X4 u5_mult_82_U12556 ( .A(fracta_mul[29]), .ZN(u5_mult_82_n6999) );
  NOR2_X4 u5_mult_82_U12555 ( .A1(u5_mult_82_net64415), .A2(u5_mult_82_n6665), 
        .ZN(u5_mult_82_ab_28__8_) );
  NOR2_X4 u5_mult_82_U12554 ( .A1(u5_mult_82_net64469), .A2(u5_mult_82_n6665), 
        .ZN(u5_mult_82_ab_28__11_) );
  NOR2_X4 u5_mult_82_U12553 ( .A1(u5_mult_82_net64487), .A2(u5_mult_82_n6665), 
        .ZN(u5_mult_82_ab_28__12_) );
  NOR2_X4 u5_mult_82_U12552 ( .A1(u5_mult_82_net64505), .A2(u5_mult_82_n6665), 
        .ZN(u5_mult_82_ab_28__13_) );
  NOR2_X4 u5_mult_82_U12551 ( .A1(u5_mult_82_net64523), .A2(u5_mult_82_n6665), 
        .ZN(u5_mult_82_ab_28__14_) );
  NOR2_X4 u5_mult_82_U12550 ( .A1(u5_mult_82_n6933), .A2(u5_mult_82_n6665), 
        .ZN(u5_mult_82_ab_28__15_) );
  NOR2_X4 u5_mult_82_U12549 ( .A1(u5_mult_82_net64559), .A2(u5_mult_82_n6664), 
        .ZN(u5_mult_82_ab_28__16_) );
  NOR2_X4 u5_mult_82_U12548 ( .A1(u5_mult_82_net64667), .A2(u5_mult_82_n6664), 
        .ZN(u5_mult_82_ab_28__22_) );
  NOR2_X4 u5_mult_82_U12547 ( .A1(u5_mult_82_net64685), .A2(u5_mult_82_n6664), 
        .ZN(u5_mult_82_ab_28__23_) );
  NOR2_X4 u5_mult_82_U12546 ( .A1(u5_mult_82_n6885), .A2(u5_mult_82_n6664), 
        .ZN(u5_mult_82_ab_28__25_) );
  NOR2_X4 u5_mult_82_U12545 ( .A1(u5_mult_82_n6875), .A2(u5_mult_82_n6664), 
        .ZN(u5_mult_82_ab_28__27_) );
  NOR2_X4 u5_mult_82_U12544 ( .A1(u5_mult_82_n6857), .A2(u5_mult_82_n6663), 
        .ZN(u5_mult_82_ab_28__30_) );
  NOR2_X4 u5_mult_82_U12543 ( .A1(u5_mult_82_n6850), .A2(u5_mult_82_n6663), 
        .ZN(u5_mult_82_ab_28__31_) );
  NOR2_X4 u5_mult_82_U12542 ( .A1(u5_mult_82_n6838), .A2(u5_mult_82_n6663), 
        .ZN(u5_mult_82_ab_28__33_) );
  NOR2_X4 u5_mult_82_U12541 ( .A1(u5_mult_82_net64901), .A2(u5_mult_82_n6663), 
        .ZN(u5_mult_82_ab_28__35_) );
  NOR2_X4 u5_mult_82_U12540 ( .A1(u5_mult_82_net64937), .A2(u5_mult_82_n6663), 
        .ZN(u5_mult_82_ab_28__37_) );
  NOR2_X4 u5_mult_82_U12539 ( .A1(u5_mult_82_n6821), .A2(u5_mult_82_n6664), 
        .ZN(u5_mult_82_ab_28__41_) );
  NOR2_X4 u5_mult_82_U12538 ( .A1(u5_mult_82_n6816), .A2(u5_mult_82_n6664), 
        .ZN(u5_mult_82_ab_28__42_) );
  NOR2_X4 u5_mult_82_U12537 ( .A1(u5_mult_82_n6804), .A2(u5_mult_82_n6664), 
        .ZN(u5_mult_82_ab_28__44_) );
  NOR2_X4 u5_mult_82_U12536 ( .A1(u5_mult_82_n6797), .A2(u5_mult_82_n6664), 
        .ZN(u5_mult_82_ab_28__45_) );
  NOR2_X4 u5_mult_82_U12535 ( .A1(u5_mult_82_n6791), .A2(u5_mult_82_n6665), 
        .ZN(u5_mult_82_ab_28__46_) );
  NOR2_X4 u5_mult_82_U12534 ( .A1(u5_mult_82_n6784), .A2(u5_mult_82_n6664), 
        .ZN(u5_mult_82_ab_28__47_) );
  NOR2_X4 u5_mult_82_U12533 ( .A1(u5_mult_82_n6778), .A2(u5_mult_82_n6666), 
        .ZN(u5_mult_82_ab_28__48_) );
  NOR2_X4 u5_mult_82_U12532 ( .A1(u5_mult_82_n6773), .A2(u5_mult_82_n6663), 
        .ZN(u5_mult_82_ab_28__49_) );
  NOR2_X4 u5_mult_82_U12531 ( .A1(u5_mult_82_n6941), .A2(u5_mult_82_n6658), 
        .ZN(u5_mult_82_ab_27__7_) );
  NOR2_X4 u5_mult_82_U12530 ( .A1(u5_mult_82_net64417), .A2(u5_mult_82_n6658), 
        .ZN(u5_mult_82_ab_27__8_) );
  NOR2_X4 u5_mult_82_U12529 ( .A1(u5_mult_82_net64471), .A2(u5_mult_82_n6658), 
        .ZN(u5_mult_82_ab_27__11_) );
  NOR2_X4 u5_mult_82_U12528 ( .A1(u5_mult_82_n6934), .A2(u5_mult_82_n6658), 
        .ZN(u5_mult_82_ab_27__15_) );
  NOR2_X4 u5_mult_82_U12527 ( .A1(u5_mult_82_net64561), .A2(u5_mult_82_n6657), 
        .ZN(u5_mult_82_ab_27__16_) );
  NOR2_X4 u5_mult_82_U12526 ( .A1(u5_mult_82_n6921), .A2(u5_mult_82_n6657), 
        .ZN(u5_mult_82_ab_27__18_) );
  NOR2_X4 u5_mult_82_U12525 ( .A1(u5_mult_82_net64687), .A2(u5_mult_82_n6657), 
        .ZN(u5_mult_82_ab_27__23_) );
  NOR2_X4 u5_mult_82_U12524 ( .A1(u5_mult_82_n6892), .A2(u5_mult_82_n6657), 
        .ZN(u5_mult_82_ab_27__24_) );
  NOR2_X4 u5_mult_82_U12523 ( .A1(u5_mult_82_n6886), .A2(u5_mult_82_n6657), 
        .ZN(u5_mult_82_ab_27__25_) );
  NOR2_X4 u5_mult_82_U12522 ( .A1(u5_mult_82_n6881), .A2(u5_mult_82_n6657), 
        .ZN(u5_mult_82_ab_27__26_) );
  NOR2_X4 u5_mult_82_U12521 ( .A1(u5_mult_82_n6863), .A2(u5_mult_82_n6656), 
        .ZN(u5_mult_82_ab_27__29_) );
  NOR2_X4 u5_mult_82_U12520 ( .A1(u5_mult_82_n6844), .A2(u5_mult_82_n6656), 
        .ZN(u5_mult_82_ab_27__32_) );
  NOR2_X4 u5_mult_82_U12519 ( .A1(u5_mult_82_net64885), .A2(u5_mult_82_n6656), 
        .ZN(u5_mult_82_ab_27__34_) );
  NOR2_X4 u5_mult_82_U12518 ( .A1(u5_mult_82_n6828), .A2(u5_mult_82_n6655), 
        .ZN(u5_mult_82_ab_27__40_) );
  NOR2_X4 u5_mult_82_U12517 ( .A1(u5_mult_82_n6947), .A2(u5_mult_82_n6651), 
        .ZN(u5_mult_82_ab_26__4_) );
  NOR2_X4 u5_mult_82_U12516 ( .A1(u5_mult_82_net64381), .A2(u5_mult_82_n6651), 
        .ZN(u5_mult_82_ab_26__6_) );
  NOR2_X4 u5_mult_82_U12515 ( .A1(u5_mult_82_net64417), .A2(u5_mult_82_n6651), 
        .ZN(u5_mult_82_ab_26__8_) );
  NOR2_X4 u5_mult_82_U12514 ( .A1(u5_mult_82_net64435), .A2(u5_mult_82_n6651), 
        .ZN(u5_mult_82_ab_26__9_) );
  NOR2_X4 u5_mult_82_U12513 ( .A1(u5_mult_82_net64489), .A2(u5_mult_82_n6651), 
        .ZN(u5_mult_82_ab_26__12_) );
  NOR2_X4 u5_mult_82_U12512 ( .A1(u5_mult_82_net64507), .A2(u5_mult_82_n6651), 
        .ZN(u5_mult_82_ab_26__13_) );
  NOR2_X4 u5_mult_82_U12511 ( .A1(u5_mult_82_n6934), .A2(u5_mult_82_n6651), 
        .ZN(u5_mult_82_ab_26__15_) );
  NOR2_X4 u5_mult_82_U12510 ( .A1(u5_mult_82_net64561), .A2(u5_mult_82_n6650), 
        .ZN(u5_mult_82_ab_26__16_) );
  NOR2_X4 u5_mult_82_U12509 ( .A1(u5_mult_82_n6928), .A2(u5_mult_82_n6650), 
        .ZN(u5_mult_82_ab_26__17_) );
  NOR2_X4 u5_mult_82_U12508 ( .A1(u5_mult_82_n6914), .A2(u5_mult_82_n6650), 
        .ZN(u5_mult_82_ab_26__19_) );
  NOR2_X4 u5_mult_82_U12507 ( .A1(u5_mult_82_n6881), .A2(u5_mult_82_n6650), 
        .ZN(u5_mult_82_ab_26__26_) );
  NOR2_X4 u5_mult_82_U12506 ( .A1(u5_mult_82_n6869), .A2(u5_mult_82_n6649), 
        .ZN(u5_mult_82_ab_26__28_) );
  NOR2_X4 u5_mult_82_U12505 ( .A1(u5_mult_82_n6858), .A2(u5_mult_82_n6649), 
        .ZN(u5_mult_82_ab_26__30_) );
  NOR2_X4 u5_mult_82_U12504 ( .A1(u5_mult_82_n6839), .A2(u5_mult_82_n6649), 
        .ZN(u5_mult_82_ab_26__33_) );
  NOR2_X4 u5_mult_82_U12503 ( .A1(u5_mult_82_net64903), .A2(u5_mult_82_n6649), 
        .ZN(u5_mult_82_ab_26__35_) );
  NOR2_X4 u5_mult_82_U12502 ( .A1(u5_mult_82_n6828), .A2(u5_mult_82_n6651), 
        .ZN(u5_mult_82_ab_26__40_) );
  NOR2_X4 u5_mult_82_U12501 ( .A1(u5_mult_82_n6817), .A2(u5_mult_82_n6651), 
        .ZN(u5_mult_82_ab_26__42_) );
  NOR2_X4 u5_mult_82_U12500 ( .A1(u5_mult_82_n6812), .A2(u5_mult_82_n6651), 
        .ZN(u5_mult_82_ab_26__43_) );
  NOR2_X4 u5_mult_82_U12499 ( .A1(u5_mult_82_n6798), .A2(u5_mult_82_n6651), 
        .ZN(u5_mult_82_ab_26__45_) );
  NOR2_X4 u5_mult_82_U12498 ( .A1(u5_mult_82_n6792), .A2(u5_mult_82_n6650), 
        .ZN(u5_mult_82_ab_26__46_) );
  NOR2_X4 u5_mult_82_U12497 ( .A1(u5_mult_82_net64363), .A2(
        u5_mult_82_net65679), .ZN(u5_mult_82_ab_25__5_) );
  NOR2_X4 u5_mult_82_U12496 ( .A1(u5_mult_82_net64381), .A2(
        u5_mult_82_net65679), .ZN(u5_mult_82_ab_25__6_) );
  NOR2_X4 u5_mult_82_U12495 ( .A1(u5_mult_82_n6941), .A2(u5_mult_82_net65679), 
        .ZN(u5_mult_82_ab_25__7_) );
  NOR2_X4 u5_mult_82_U12494 ( .A1(u5_mult_82_net64417), .A2(
        u5_mult_82_net65679), .ZN(u5_mult_82_ab_25__8_) );
  NOR2_X4 u5_mult_82_U12493 ( .A1(u5_mult_82_net64435), .A2(
        u5_mult_82_net65679), .ZN(u5_mult_82_ab_25__9_) );
  NOR2_X4 u5_mult_82_U12492 ( .A1(u5_mult_82_net64471), .A2(
        u5_mult_82_net65679), .ZN(u5_mult_82_ab_25__11_) );
  NOR2_X4 u5_mult_82_U12491 ( .A1(u5_mult_82_net64489), .A2(
        u5_mult_82_net65679), .ZN(u5_mult_82_ab_25__12_) );
  NOR2_X4 u5_mult_82_U12490 ( .A1(u5_mult_82_net64525), .A2(
        u5_mult_82_net65679), .ZN(u5_mult_82_ab_25__14_) );
  NOR2_X4 u5_mult_82_U12489 ( .A1(u5_mult_82_net64561), .A2(
        u5_mult_82_net65677), .ZN(u5_mult_82_ab_25__16_) );
  NOR2_X4 u5_mult_82_U12488 ( .A1(u5_mult_82_n6928), .A2(u5_mult_82_net65677), 
        .ZN(u5_mult_82_ab_25__17_) );
  NOR2_X4 u5_mult_82_U12487 ( .A1(u5_mult_82_n6905), .A2(u5_mult_82_net65677), 
        .ZN(u5_mult_82_ab_25__20_) );
  NOR2_X4 u5_mult_82_U12486 ( .A1(u5_mult_82_n6881), .A2(u5_mult_82_net65677), 
        .ZN(u5_mult_82_ab_25__26_) );
  NOR2_X4 u5_mult_82_U12485 ( .A1(u5_mult_82_n6869), .A2(u5_mult_82_net65675), 
        .ZN(u5_mult_82_ab_25__28_) );
  NOR2_X4 u5_mult_82_U12484 ( .A1(u5_mult_82_n6863), .A2(u5_mult_82_net65675), 
        .ZN(u5_mult_82_ab_25__29_) );
  NOR2_X4 u5_mult_82_U12483 ( .A1(u5_mult_82_n6844), .A2(u5_mult_82_net65675), 
        .ZN(u5_mult_82_ab_25__32_) );
  NOR2_X4 u5_mult_82_U12482 ( .A1(u5_mult_82_n6839), .A2(u5_mult_82_net65675), 
        .ZN(u5_mult_82_ab_25__33_) );
  NOR2_X4 u5_mult_82_U12481 ( .A1(u5_mult_82_net64885), .A2(
        u5_mult_82_net65675), .ZN(u5_mult_82_ab_25__34_) );
  NOR2_X4 u5_mult_82_U12480 ( .A1(u5_mult_82_n6831), .A2(u5_mult_82_net65675), 
        .ZN(u5_mult_82_ab_25__39_) );
  NOR2_X4 u5_mult_82_U12479 ( .A1(u5_mult_82_n6828), .A2(u5_mult_82_net65677), 
        .ZN(u5_mult_82_ab_25__40_) );
  NOR2_X4 u5_mult_82_U12478 ( .A1(u5_mult_82_n6822), .A2(u5_mult_82_net65677), 
        .ZN(u5_mult_82_ab_25__41_) );
  NOR2_X4 u5_mult_82_U12477 ( .A1(u5_mult_82_n6812), .A2(u5_mult_82_net65677), 
        .ZN(u5_mult_82_ab_25__43_) );
  NOR2_X4 u5_mult_82_U12476 ( .A1(u5_mult_82_n6792), .A2(u5_mult_82_net65679), 
        .ZN(u5_mult_82_ab_25__46_) );
  NOR2_X4 u5_mult_82_U12475 ( .A1(u5_mult_82_n6947), .A2(u5_mult_82_n6644), 
        .ZN(u5_mult_82_ab_24__4_) );
  NOR2_X4 u5_mult_82_U12474 ( .A1(u5_mult_82_net64489), .A2(u5_mult_82_n6644), 
        .ZN(u5_mult_82_ab_24__12_) );
  NOR2_X4 u5_mult_82_U12473 ( .A1(u5_mult_82_net64507), .A2(u5_mult_82_n6644), 
        .ZN(u5_mult_82_ab_24__13_) );
  NOR2_X4 u5_mult_82_U12472 ( .A1(u5_mult_82_n6928), .A2(u5_mult_82_n6643), 
        .ZN(u5_mult_82_ab_24__17_) );
  NOR2_X4 u5_mult_82_U12471 ( .A1(u5_mult_82_n6921), .A2(u5_mult_82_n6643), 
        .ZN(u5_mult_82_ab_24__18_) );
  NOR2_X4 u5_mult_82_U12470 ( .A1(u5_mult_82_n6905), .A2(u5_mult_82_n6643), 
        .ZN(u5_mult_82_ab_24__20_) );
  NOR2_X4 u5_mult_82_U12469 ( .A1(u5_mult_82_n6897), .A2(u5_mult_82_n6643), 
        .ZN(u5_mult_82_ab_24__21_) );
  NOR2_X4 u5_mult_82_U12468 ( .A1(u5_mult_82_n6863), .A2(u5_mult_82_n6642), 
        .ZN(u5_mult_82_ab_24__29_) );
  NOR2_X4 u5_mult_82_U12467 ( .A1(u5_mult_82_n6851), .A2(u5_mult_82_n6642), 
        .ZN(u5_mult_82_ab_24__31_) );
  NOR2_X4 u5_mult_82_U12466 ( .A1(u5_mult_82_n6839), .A2(u5_mult_82_n6642), 
        .ZN(u5_mult_82_ab_24__33_) );
  NOR2_X4 u5_mult_82_U12465 ( .A1(u5_mult_82_net64885), .A2(u5_mult_82_n6642), 
        .ZN(u5_mult_82_ab_24__34_) );
  NOR2_X4 u5_mult_82_U12464 ( .A1(u5_mult_82_n6822), .A2(u5_mult_82_n6644), 
        .ZN(u5_mult_82_ab_24__41_) );
  NOR2_X4 u5_mult_82_U12463 ( .A1(u5_mult_82_n6812), .A2(u5_mult_82_n6644), 
        .ZN(u5_mult_82_ab_24__43_) );
  NOR2_X4 u5_mult_82_U12462 ( .A1(u5_mult_82_n6785), .A2(u5_mult_82_n6645), 
        .ZN(u5_mult_82_ab_24__47_) );
  NOR2_X4 u5_mult_82_U12461 ( .A1(u5_mult_82_n6941), .A2(u5_mult_82_net65713), 
        .ZN(u5_mult_82_ab_23__7_) );
  NOR2_X4 u5_mult_82_U12460 ( .A1(u5_mult_82_net64417), .A2(
        u5_mult_82_net65717), .ZN(u5_mult_82_ab_23__8_) );
  NOR2_X4 u5_mult_82_U12459 ( .A1(u5_mult_82_net64471), .A2(
        u5_mult_82_net65717), .ZN(u5_mult_82_ab_23__11_) );
  NOR2_X4 u5_mult_82_U12458 ( .A1(u5_mult_82_n6921), .A2(u5_mult_82_net65713), 
        .ZN(u5_mult_82_ab_23__18_) );
  NOR2_X4 u5_mult_82_U12457 ( .A1(u5_mult_82_n6897), .A2(u5_mult_82_net65713), 
        .ZN(u5_mult_82_ab_23__21_) );
  NOR2_X4 u5_mult_82_U12456 ( .A1(u5_mult_82_n6892), .A2(u5_mult_82_net65713), 
        .ZN(u5_mult_82_ab_23__24_) );
  NOR2_X4 u5_mult_82_U12455 ( .A1(u5_mult_82_n6886), .A2(u5_mult_82_net65713), 
        .ZN(u5_mult_82_ab_23__25_) );
  NOR2_X4 u5_mult_82_U12454 ( .A1(u5_mult_82_n6881), .A2(u5_mult_82_net65713), 
        .ZN(u5_mult_82_ab_23__26_) );
  NOR2_X4 u5_mult_82_U12453 ( .A1(u5_mult_82_n6869), .A2(u5_mult_82_net65711), 
        .ZN(u5_mult_82_ab_23__28_) );
  NOR2_X4 u5_mult_82_U12452 ( .A1(u5_mult_82_n6863), .A2(u5_mult_82_net65711), 
        .ZN(u5_mult_82_ab_23__29_) );
  NOR2_X4 u5_mult_82_U12451 ( .A1(u5_mult_82_n6858), .A2(u5_mult_82_net65711), 
        .ZN(u5_mult_82_ab_23__30_) );
  NOR2_X4 u5_mult_82_U12450 ( .A1(u5_mult_82_n6851), .A2(u5_mult_82_net65711), 
        .ZN(u5_mult_82_ab_23__31_) );
  NOR2_X4 u5_mult_82_U12449 ( .A1(u5_mult_82_n6844), .A2(u5_mult_82_net65711), 
        .ZN(u5_mult_82_ab_23__32_) );
  NOR2_X4 u5_mult_82_U12448 ( .A1(u5_mult_82_net64885), .A2(
        u5_mult_82_net65711), .ZN(u5_mult_82_ab_23__34_) );
  NOR2_X4 u5_mult_82_U12447 ( .A1(u5_mult_82_net64939), .A2(
        u5_mult_82_net65711), .ZN(u5_mult_82_ab_23__37_) );
  NOR2_X4 u5_mult_82_U12446 ( .A1(u5_mult_82_n6831), .A2(u5_mult_82_net65711), 
        .ZN(u5_mult_82_ab_23__39_) );
  NOR2_X4 u5_mult_82_U12445 ( .A1(u5_mult_82_n6812), .A2(u5_mult_82_net65717), 
        .ZN(u5_mult_82_ab_23__43_) );
  NOR2_X4 u5_mult_82_U12444 ( .A1(u5_mult_82_n6779), .A2(u5_mult_82_net65713), 
        .ZN(u5_mult_82_ab_23__48_) );
  NOR2_X4 u5_mult_82_U12443 ( .A1(u5_mult_82_n6761), .A2(u5_mult_82_n1344), 
        .ZN(u5_mult_82_ab_23__51_) );
  NOR2_X4 u5_mult_82_U12442 ( .A1(u5_mult_82_net64417), .A2(u5_mult_82_n6637), 
        .ZN(u5_mult_82_ab_22__8_) );
  NOR2_X4 u5_mult_82_U12441 ( .A1(u5_mult_82_net64453), .A2(u5_mult_82_n6637), 
        .ZN(u5_mult_82_ab_22__10_) );
  NOR2_X4 u5_mult_82_U12440 ( .A1(u5_mult_82_net64489), .A2(u5_mult_82_n6637), 
        .ZN(u5_mult_82_ab_22__12_) );
  NOR2_X4 u5_mult_82_U12439 ( .A1(u5_mult_82_net64507), .A2(u5_mult_82_n6637), 
        .ZN(u5_mult_82_ab_22__13_) );
  NOR2_X4 u5_mult_82_U12438 ( .A1(u5_mult_82_n6921), .A2(u5_mult_82_n6636), 
        .ZN(u5_mult_82_ab_22__18_) );
  NOR2_X4 u5_mult_82_U12437 ( .A1(u5_mult_82_net64669), .A2(u5_mult_82_n6636), 
        .ZN(u5_mult_82_ab_22__22_) );
  NOR2_X4 u5_mult_82_U12436 ( .A1(u5_mult_82_n6886), .A2(u5_mult_82_n6636), 
        .ZN(u5_mult_82_ab_22__25_) );
  NOR2_X4 u5_mult_82_U12435 ( .A1(u5_mult_82_n6881), .A2(u5_mult_82_n6636), 
        .ZN(u5_mult_82_ab_22__26_) );
  NOR2_X4 u5_mult_82_U12434 ( .A1(u5_mult_82_n6876), .A2(u5_mult_82_n6636), 
        .ZN(u5_mult_82_ab_22__27_) );
  NOR2_X4 u5_mult_82_U12433 ( .A1(u5_mult_82_n6863), .A2(u5_mult_82_n6635), 
        .ZN(u5_mult_82_ab_22__29_) );
  NOR2_X4 u5_mult_82_U12432 ( .A1(u5_mult_82_n6858), .A2(u5_mult_82_n6635), 
        .ZN(u5_mult_82_ab_22__30_) );
  NOR2_X4 u5_mult_82_U12431 ( .A1(u5_mult_82_n6851), .A2(u5_mult_82_n6635), 
        .ZN(u5_mult_82_ab_22__31_) );
  NOR2_X4 u5_mult_82_U12430 ( .A1(u5_mult_82_n6844), .A2(u5_mult_82_n6635), 
        .ZN(u5_mult_82_ab_22__32_) );
  NOR2_X4 u5_mult_82_U12429 ( .A1(u5_mult_82_net64885), .A2(u5_mult_82_n6635), 
        .ZN(u5_mult_82_ab_22__34_) );
  NOR2_X4 u5_mult_82_U12428 ( .A1(u5_mult_82_net64903), .A2(u5_mult_82_n6635), 
        .ZN(u5_mult_82_ab_22__35_) );
  NOR2_X4 u5_mult_82_U12427 ( .A1(u5_mult_82_net64939), .A2(u5_mult_82_n6635), 
        .ZN(u5_mult_82_ab_22__37_) );
  NOR2_X4 u5_mult_82_U12426 ( .A1(u5_mult_82_n6828), .A2(u5_mult_82_n6636), 
        .ZN(u5_mult_82_ab_22__40_) );
  NOR2_X4 u5_mult_82_U12425 ( .A1(u5_mult_82_n6805), .A2(u5_mult_82_n6636), 
        .ZN(u5_mult_82_ab_22__44_) );
  NOR2_X4 u5_mult_82_U12424 ( .A1(u5_mult_82_net64471), .A2(u5_mult_82_n6630), 
        .ZN(u5_mult_82_ab_21__11_) );
  NOR2_X4 u5_mult_82_U12423 ( .A1(u5_mult_82_net64507), .A2(u5_mult_82_n6630), 
        .ZN(u5_mult_82_ab_21__13_) );
  NOR2_X4 u5_mult_82_U12422 ( .A1(u5_mult_82_net64525), .A2(u5_mult_82_n6630), 
        .ZN(u5_mult_82_ab_21__14_) );
  NOR2_X4 u5_mult_82_U12421 ( .A1(u5_mult_82_n6934), .A2(u5_mult_82_n6630), 
        .ZN(u5_mult_82_ab_21__15_) );
  NOR2_X4 u5_mult_82_U12420 ( .A1(u5_mult_82_n6921), .A2(u5_mult_82_n6629), 
        .ZN(u5_mult_82_ab_21__18_) );
  NOR2_X4 u5_mult_82_U12419 ( .A1(u5_mult_82_n6914), .A2(u5_mult_82_n6629), 
        .ZN(u5_mult_82_ab_21__19_) );
  NOR2_X4 u5_mult_82_U12418 ( .A1(u5_mult_82_net64669), .A2(u5_mult_82_n6629), 
        .ZN(u5_mult_82_ab_21__22_) );
  NOR2_X4 u5_mult_82_U12417 ( .A1(u5_mult_82_n6886), .A2(u5_mult_82_n6629), 
        .ZN(u5_mult_82_ab_21__25_) );
  NOR2_X4 u5_mult_82_U12416 ( .A1(u5_mult_82_n6881), .A2(u5_mult_82_n6629), 
        .ZN(u5_mult_82_ab_21__26_) );
  NOR2_X4 u5_mult_82_U12415 ( .A1(u5_mult_82_n6876), .A2(u5_mult_82_n6629), 
        .ZN(u5_mult_82_ab_21__27_) );
  NOR2_X4 u5_mult_82_U12414 ( .A1(u5_mult_82_n6869), .A2(u5_mult_82_n6628), 
        .ZN(u5_mult_82_ab_21__28_) );
  NOR2_X4 u5_mult_82_U12413 ( .A1(u5_mult_82_n6858), .A2(u5_mult_82_n6628), 
        .ZN(u5_mult_82_ab_21__30_) );
  NOR2_X4 u5_mult_82_U12412 ( .A1(u5_mult_82_n6839), .A2(u5_mult_82_n6628), 
        .ZN(u5_mult_82_ab_21__33_) );
  NOR2_X4 u5_mult_82_U12411 ( .A1(u5_mult_82_net64903), .A2(u5_mult_82_n6628), 
        .ZN(u5_mult_82_ab_21__35_) );
  NOR2_X4 u5_mult_82_U12410 ( .A1(u5_mult_82_net64939), .A2(u5_mult_82_n6628), 
        .ZN(u5_mult_82_ab_21__37_) );
  NOR2_X4 u5_mult_82_U12409 ( .A1(u5_mult_82_n6832), .A2(u5_mult_82_n6628), 
        .ZN(u5_mult_82_ab_21__39_) );
  NOR2_X4 u5_mult_82_U12408 ( .A1(u5_mult_82_n6828), .A2(u5_mult_82_n6630), 
        .ZN(u5_mult_82_ab_21__40_) );
  NOR2_X4 u5_mult_82_U12407 ( .A1(u5_mult_82_n6817), .A2(u5_mult_82_n6630), 
        .ZN(u5_mult_82_ab_21__42_) );
  NOR2_X4 u5_mult_82_U12406 ( .A1(u5_mult_82_n6779), .A2(u5_mult_82_n6629), 
        .ZN(u5_mult_82_ab_21__48_) );
  NOR2_X4 u5_mult_82_U12405 ( .A1(u5_mult_82_n6954), .A2(u5_mult_82_n6624), 
        .ZN(u5_mult_82_ab_20__3_) );
  NOR2_X4 u5_mult_82_U12404 ( .A1(u5_mult_82_n6947), .A2(u5_mult_82_n6623), 
        .ZN(u5_mult_82_ab_20__4_) );
  NOR2_X4 u5_mult_82_U12403 ( .A1(u5_mult_82_net64561), .A2(u5_mult_82_n6622), 
        .ZN(u5_mult_82_ab_20__16_) );
  NOR2_X4 u5_mult_82_U12402 ( .A1(u5_mult_82_n6914), .A2(u5_mult_82_n6622), 
        .ZN(u5_mult_82_ab_20__19_) );
  NOR2_X4 u5_mult_82_U12401 ( .A1(u5_mult_82_n6905), .A2(u5_mult_82_n6622), 
        .ZN(u5_mult_82_ab_20__20_) );
  NOR2_X4 u5_mult_82_U12400 ( .A1(u5_mult_82_n6897), .A2(u5_mult_82_n6622), 
        .ZN(u5_mult_82_ab_20__21_) );
  NOR2_X4 u5_mult_82_U12399 ( .A1(u5_mult_82_net64669), .A2(u5_mult_82_n6622), 
        .ZN(u5_mult_82_ab_20__22_) );
  NOR2_X4 u5_mult_82_U12398 ( .A1(u5_mult_82_net64687), .A2(u5_mult_82_n6622), 
        .ZN(u5_mult_82_ab_20__23_) );
  NOR2_X4 u5_mult_82_U12397 ( .A1(u5_mult_82_n6892), .A2(u5_mult_82_n6622), 
        .ZN(u5_mult_82_ab_20__24_) );
  NOR2_X4 u5_mult_82_U12396 ( .A1(u5_mult_82_n6881), .A2(u5_mult_82_n6622), 
        .ZN(u5_mult_82_ab_20__26_) );
  NOR2_X4 u5_mult_82_U12395 ( .A1(u5_mult_82_n6876), .A2(u5_mult_82_n6622), 
        .ZN(u5_mult_82_ab_20__27_) );
  NOR2_X4 u5_mult_82_U12394 ( .A1(u5_mult_82_n6863), .A2(u5_mult_82_n6621), 
        .ZN(u5_mult_82_ab_20__29_) );
  NOR2_X4 u5_mult_82_U12393 ( .A1(u5_mult_82_n6851), .A2(u5_mult_82_n6621), 
        .ZN(u5_mult_82_ab_20__31_) );
  NOR2_X4 u5_mult_82_U12392 ( .A1(u5_mult_82_n6844), .A2(u5_mult_82_n6621), 
        .ZN(u5_mult_82_ab_20__32_) );
  NOR2_X4 u5_mult_82_U12391 ( .A1(u5_mult_82_n6839), .A2(u5_mult_82_n6621), 
        .ZN(u5_mult_82_ab_20__33_) );
  NOR2_X4 u5_mult_82_U12390 ( .A1(u5_mult_82_net64885), .A2(u5_mult_82_n6621), 
        .ZN(u5_mult_82_ab_20__34_) );
  NOR2_X4 u5_mult_82_U12389 ( .A1(u5_mult_82_n6828), .A2(u5_mult_82_n6622), 
        .ZN(u5_mult_82_ab_20__40_) );
  NOR2_X4 u5_mult_82_U12388 ( .A1(u5_mult_82_n6822), .A2(u5_mult_82_n6623), 
        .ZN(u5_mult_82_ab_20__41_) );
  NOR2_X4 u5_mult_82_U12387 ( .A1(u5_mult_82_n6817), .A2(u5_mult_82_n6622), 
        .ZN(u5_mult_82_ab_20__42_) );
  NOR2_X4 u5_mult_82_U12386 ( .A1(u5_mult_82_n6812), .A2(u5_mult_82_n6622), 
        .ZN(u5_mult_82_ab_20__43_) );
  NOR2_X4 u5_mult_82_U12385 ( .A1(u5_mult_82_n6779), .A2(u5_mult_82_n6622), 
        .ZN(u5_mult_82_ab_20__48_) );
  NOR2_X4 u5_mult_82_U12384 ( .A1(u5_mult_82_n6774), .A2(u5_mult_82_n6621), 
        .ZN(u5_mult_82_ab_20__49_) );
  NOR2_X4 u5_mult_82_U12383 ( .A1(u5_mult_82_n6947), .A2(u5_mult_82_n6616), 
        .ZN(u5_mult_82_ab_19__4_) );
  NOR2_X4 u5_mult_82_U12382 ( .A1(u5_mult_82_net64363), .A2(u5_mult_82_n6616), 
        .ZN(u5_mult_82_ab_19__5_) );
  NOR2_X4 u5_mult_82_U12381 ( .A1(u5_mult_82_net64381), .A2(u5_mult_82_n6616), 
        .ZN(u5_mult_82_ab_19__6_) );
  NOR2_X4 u5_mult_82_U12380 ( .A1(u5_mult_82_n6905), .A2(u5_mult_82_n6615), 
        .ZN(u5_mult_82_ab_19__20_) );
  NOR2_X4 u5_mult_82_U12379 ( .A1(u5_mult_82_n6897), .A2(u5_mult_82_n6615), 
        .ZN(u5_mult_82_ab_19__21_) );
  NOR2_X4 u5_mult_82_U12378 ( .A1(u5_mult_82_net64669), .A2(u5_mult_82_n6615), 
        .ZN(u5_mult_82_ab_19__22_) );
  NOR2_X4 u5_mult_82_U12377 ( .A1(u5_mult_82_net64687), .A2(u5_mult_82_n6615), 
        .ZN(u5_mult_82_ab_19__23_) );
  NOR2_X4 u5_mult_82_U12376 ( .A1(u5_mult_82_n6886), .A2(u5_mult_82_n6615), 
        .ZN(u5_mult_82_ab_19__25_) );
  NOR2_X4 u5_mult_82_U12375 ( .A1(u5_mult_82_n6876), .A2(u5_mult_82_n6615), 
        .ZN(u5_mult_82_ab_19__27_) );
  NOR2_X4 u5_mult_82_U12374 ( .A1(u5_mult_82_n6869), .A2(u5_mult_82_n6614), 
        .ZN(u5_mult_82_ab_19__28_) );
  NOR2_X4 u5_mult_82_U12373 ( .A1(u5_mult_82_n6863), .A2(u5_mult_82_n6614), 
        .ZN(u5_mult_82_ab_19__29_) );
  NOR2_X4 u5_mult_82_U12372 ( .A1(u5_mult_82_n6839), .A2(u5_mult_82_n6614), 
        .ZN(u5_mult_82_ab_19__33_) );
  NOR2_X4 u5_mult_82_U12371 ( .A1(u5_mult_82_net64903), .A2(u5_mult_82_n6614), 
        .ZN(u5_mult_82_ab_19__35_) );
  NOR2_X4 u5_mult_82_U12370 ( .A1(u5_mult_82_net64939), .A2(u5_mult_82_n6614), 
        .ZN(u5_mult_82_ab_19__37_) );
  NOR2_X4 u5_mult_82_U12369 ( .A1(u5_mult_82_n6812), .A2(u5_mult_82_n6615), 
        .ZN(u5_mult_82_ab_19__43_) );
  NOR2_X4 u5_mult_82_U12368 ( .A1(u5_mult_82_n6774), .A2(u5_mult_82_n6614), 
        .ZN(u5_mult_82_ab_19__49_) );
  NOR2_X4 u5_mult_82_U12367 ( .A1(u5_mult_82_n6941), .A2(u5_mult_82_n6610), 
        .ZN(u5_mult_82_ab_18__7_) );
  NOR2_X4 u5_mult_82_U12366 ( .A1(u5_mult_82_n6934), .A2(u5_mult_82_n6610), 
        .ZN(u5_mult_82_ab_18__15_) );
  NOR2_X4 u5_mult_82_U12365 ( .A1(u5_mult_82_net64561), .A2(u5_mult_82_n6609), 
        .ZN(u5_mult_82_ab_18__16_) );
  NOR2_X4 u5_mult_82_U12364 ( .A1(u5_mult_82_n6928), .A2(u5_mult_82_n6609), 
        .ZN(u5_mult_82_ab_18__17_) );
  NOR2_X4 u5_mult_82_U12363 ( .A1(u5_mult_82_n6921), .A2(u5_mult_82_n6609), 
        .ZN(u5_mult_82_ab_18__18_) );
  NOR2_X4 u5_mult_82_U12362 ( .A1(u5_mult_82_n6905), .A2(u5_mult_82_n6609), 
        .ZN(u5_mult_82_ab_18__20_) );
  NOR2_X4 u5_mult_82_U12361 ( .A1(u5_mult_82_net64687), .A2(u5_mult_82_n6609), 
        .ZN(u5_mult_82_ab_18__23_) );
  NOR2_X4 u5_mult_82_U12360 ( .A1(u5_mult_82_n6886), .A2(u5_mult_82_n6609), 
        .ZN(u5_mult_82_ab_18__25_) );
  NOR2_X4 u5_mult_82_U12359 ( .A1(u5_mult_82_n6876), .A2(u5_mult_82_n6609), 
        .ZN(u5_mult_82_ab_18__27_) );
  NOR2_X4 u5_mult_82_U12358 ( .A1(u5_mult_82_n6869), .A2(u5_mult_82_n6608), 
        .ZN(u5_mult_82_ab_18__28_) );
  NOR2_X4 u5_mult_82_U12357 ( .A1(u5_mult_82_n6863), .A2(u5_mult_82_n6608), 
        .ZN(u5_mult_82_ab_18__29_) );
  NOR2_X4 u5_mult_82_U12356 ( .A1(u5_mult_82_n6858), .A2(u5_mult_82_n6608), 
        .ZN(u5_mult_82_ab_18__30_) );
  NOR2_X4 u5_mult_82_U12355 ( .A1(u5_mult_82_net64903), .A2(u5_mult_82_n6608), 
        .ZN(u5_mult_82_ab_18__35_) );
  NOR2_X4 u5_mult_82_U12354 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6608), 
        .ZN(u5_mult_82_ab_18__36_) );
  NOR2_X4 u5_mult_82_U12353 ( .A1(u5_mult_82_net64939), .A2(u5_mult_82_n6608), 
        .ZN(u5_mult_82_ab_18__37_) );
  NOR2_X4 u5_mult_82_U12352 ( .A1(u5_mult_82_n6832), .A2(u5_mult_82_n6608), 
        .ZN(u5_mult_82_ab_18__39_) );
  NOR2_X4 u5_mult_82_U12351 ( .A1(u5_mult_82_n6812), .A2(u5_mult_82_n6607), 
        .ZN(u5_mult_82_ab_18__43_) );
  NOR2_X4 u5_mult_82_U12350 ( .A1(u5_mult_82_n6792), .A2(u5_mult_82_n6607), 
        .ZN(u5_mult_82_ab_18__46_) );
  NOR2_X4 u5_mult_82_U12349 ( .A1(u5_mult_82_n6785), .A2(u5_mult_82_n6607), 
        .ZN(u5_mult_82_ab_18__47_) );
  INV_X4 u5_mult_82_U12348 ( .A(fracta_mul[18]), .ZN(u5_mult_82_n6998) );
  NOR2_X4 u5_mult_82_U12347 ( .A1(u5_mult_82_net64417), .A2(u5_mult_82_n6603), 
        .ZN(u5_mult_82_ab_17__8_) );
  NOR2_X4 u5_mult_82_U12346 ( .A1(u5_mult_82_net64525), .A2(u5_mult_82_n6603), 
        .ZN(u5_mult_82_ab_17__14_) );
  NOR2_X4 u5_mult_82_U12345 ( .A1(u5_mult_82_n6934), .A2(u5_mult_82_n6603), 
        .ZN(u5_mult_82_ab_17__15_) );
  NOR2_X4 u5_mult_82_U12344 ( .A1(u5_mult_82_n6928), .A2(u5_mult_82_n6602), 
        .ZN(u5_mult_82_ab_17__17_) );
  NOR2_X4 u5_mult_82_U12343 ( .A1(u5_mult_82_n6921), .A2(u5_mult_82_n6602), 
        .ZN(u5_mult_82_ab_17__18_) );
  NOR2_X4 u5_mult_82_U12342 ( .A1(u5_mult_82_n6914), .A2(u5_mult_82_n6602), 
        .ZN(u5_mult_82_ab_17__19_) );
  NOR2_X4 u5_mult_82_U12341 ( .A1(u5_mult_82_n6897), .A2(u5_mult_82_n6602), 
        .ZN(u5_mult_82_ab_17__21_) );
  NOR2_X4 u5_mult_82_U12340 ( .A1(u5_mult_82_n6892), .A2(u5_mult_82_n6602), 
        .ZN(u5_mult_82_ab_17__24_) );
  NOR2_X4 u5_mult_82_U12339 ( .A1(u5_mult_82_n6886), .A2(u5_mult_82_n6602), 
        .ZN(u5_mult_82_ab_17__25_) );
  NOR2_X4 u5_mult_82_U12338 ( .A1(u5_mult_82_n6881), .A2(u5_mult_82_n6602), 
        .ZN(u5_mult_82_ab_17__26_) );
  NOR2_X4 u5_mult_82_U12337 ( .A1(u5_mult_82_n6869), .A2(u5_mult_82_n6601), 
        .ZN(u5_mult_82_ab_17__28_) );
  NOR2_X4 u5_mult_82_U12336 ( .A1(u5_mult_82_n6851), .A2(u5_mult_82_n6601), 
        .ZN(u5_mult_82_ab_17__31_) );
  NOR2_X4 u5_mult_82_U12335 ( .A1(u5_mult_82_n6844), .A2(u5_mult_82_n6601), 
        .ZN(u5_mult_82_ab_17__32_) );
  NOR2_X4 u5_mult_82_U12334 ( .A1(u5_mult_82_net64903), .A2(u5_mult_82_n6601), 
        .ZN(u5_mult_82_ab_17__35_) );
  NOR2_X4 u5_mult_82_U12333 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6601), 
        .ZN(u5_mult_82_ab_17__36_) );
  NOR2_X4 u5_mult_82_U12332 ( .A1(u5_mult_82_net64939), .A2(u5_mult_82_n6601), 
        .ZN(u5_mult_82_ab_17__37_) );
  NOR2_X4 u5_mult_82_U12331 ( .A1(u5_mult_82_n6832), .A2(u5_mult_82_n6601), 
        .ZN(u5_mult_82_ab_17__39_) );
  NOR2_X4 u5_mult_82_U12330 ( .A1(u5_mult_82_n6817), .A2(u5_mult_82_n6600), 
        .ZN(u5_mult_82_ab_17__42_) );
  NOR2_X4 u5_mult_82_U12329 ( .A1(u5_mult_82_n6805), .A2(u5_mult_82_n6600), 
        .ZN(u5_mult_82_ab_17__44_) );
  NOR2_X4 u5_mult_82_U12328 ( .A1(u5_mult_82_n6785), .A2(u5_mult_82_n6600), 
        .ZN(u5_mult_82_ab_17__47_) );
  NOR2_X4 u5_mult_82_U12327 ( .A1(u5_mult_82_n6779), .A2(u5_mult_82_n6600), 
        .ZN(u5_mult_82_ab_17__48_) );
  INV_X4 u5_mult_82_U12326 ( .A(fracta_mul[17]), .ZN(u5_mult_82_n6997) );
  NOR2_X4 u5_mult_82_U12325 ( .A1(u5_mult_82_net64381), .A2(u5_mult_82_n6596), 
        .ZN(u5_mult_82_ab_16__6_) );
  NOR2_X4 u5_mult_82_U12324 ( .A1(u5_mult_82_net64435), .A2(u5_mult_82_n6596), 
        .ZN(u5_mult_82_ab_16__9_) );
  NOR2_X4 u5_mult_82_U12323 ( .A1(u5_mult_82_net64489), .A2(u5_mult_82_n6596), 
        .ZN(u5_mult_82_ab_16__12_) );
  NOR2_X4 u5_mult_82_U12322 ( .A1(u5_mult_82_net64507), .A2(u5_mult_82_n6596), 
        .ZN(u5_mult_82_ab_16__13_) );
  NOR2_X4 u5_mult_82_U12321 ( .A1(u5_mult_82_n6934), .A2(u5_mult_82_n6596), 
        .ZN(u5_mult_82_ab_16__15_) );
  NOR2_X4 u5_mult_82_U12320 ( .A1(u5_mult_82_net64561), .A2(u5_mult_82_n6595), 
        .ZN(u5_mult_82_ab_16__16_) );
  NOR2_X4 u5_mult_82_U12319 ( .A1(u5_mult_82_n6914), .A2(u5_mult_82_n6595), 
        .ZN(u5_mult_82_ab_16__19_) );
  NOR2_X4 u5_mult_82_U12318 ( .A1(u5_mult_82_n6905), .A2(u5_mult_82_n6595), 
        .ZN(u5_mult_82_ab_16__20_) );
  NOR2_X4 u5_mult_82_U12317 ( .A1(u5_mult_82_n6886), .A2(u5_mult_82_n6595), 
        .ZN(u5_mult_82_ab_16__25_) );
  NOR2_X4 u5_mult_82_U12316 ( .A1(u5_mult_82_n6881), .A2(u5_mult_82_n6595), 
        .ZN(u5_mult_82_ab_16__26_) );
  NOR2_X4 u5_mult_82_U12315 ( .A1(u5_mult_82_n6863), .A2(u5_mult_82_n6594), 
        .ZN(u5_mult_82_ab_16__29_) );
  NOR2_X4 u5_mult_82_U12314 ( .A1(u5_mult_82_n6851), .A2(u5_mult_82_n6594), 
        .ZN(u5_mult_82_ab_16__31_) );
  NOR2_X4 u5_mult_82_U12313 ( .A1(u5_mult_82_n6844), .A2(u5_mult_82_n6594), 
        .ZN(u5_mult_82_ab_16__32_) );
  NOR2_X4 u5_mult_82_U12312 ( .A1(u5_mult_82_n6839), .A2(u5_mult_82_n6594), 
        .ZN(u5_mult_82_ab_16__33_) );
  NOR2_X4 u5_mult_82_U12311 ( .A1(u5_mult_82_net64885), .A2(u5_mult_82_n6594), 
        .ZN(u5_mult_82_ab_16__34_) );
  NOR2_X4 u5_mult_82_U12310 ( .A1(u5_mult_82_net64903), .A2(u5_mult_82_n6594), 
        .ZN(u5_mult_82_ab_16__35_) );
  NOR2_X4 u5_mult_82_U12309 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6594), 
        .ZN(u5_mult_82_ab_16__36_) );
  NOR2_X4 u5_mult_82_U12308 ( .A1(u5_mult_82_n6822), .A2(u5_mult_82_n6593), 
        .ZN(u5_mult_82_ab_16__41_) );
  NOR2_X4 u5_mult_82_U12307 ( .A1(u5_mult_82_n6812), .A2(u5_mult_82_n6593), 
        .ZN(u5_mult_82_ab_16__43_) );
  NOR2_X4 u5_mult_82_U12306 ( .A1(u5_mult_82_n6805), .A2(u5_mult_82_n6593), 
        .ZN(u5_mult_82_ab_16__44_) );
  NOR2_X4 u5_mult_82_U12305 ( .A1(u5_mult_82_n6798), .A2(u5_mult_82_n6593), 
        .ZN(u5_mult_82_ab_16__45_) );
  NOR2_X4 u5_mult_82_U12304 ( .A1(u5_mult_82_n6792), .A2(u5_mult_82_n6593), 
        .ZN(u5_mult_82_ab_16__46_) );
  NOR2_X4 u5_mult_82_U12303 ( .A1(u5_mult_82_n6761), .A2(u5_mult_82_n6593), 
        .ZN(u5_mult_82_ab_16__51_) );
  INV_X4 u5_mult_82_U12302 ( .A(fracta_mul[16]), .ZN(u5_mult_82_n6996) );
  NOR2_X4 u5_mult_82_U12301 ( .A1(u5_mult_82_net64455), .A2(u5_mult_82_n6588), 
        .ZN(u5_mult_82_ab_15__10_) );
  NOR2_X4 u5_mult_82_U12300 ( .A1(u5_mult_82_net64509), .A2(u5_mult_82_n6588), 
        .ZN(u5_mult_82_ab_15__13_) );
  NOR2_X4 u5_mult_82_U12299 ( .A1(u5_mult_82_net64527), .A2(u5_mult_82_n6588), 
        .ZN(u5_mult_82_ab_15__14_) );
  NOR2_X4 u5_mult_82_U12298 ( .A1(u5_mult_82_n6893), .A2(u5_mult_82_n6587), 
        .ZN(u5_mult_82_ab_15__24_) );
  NOR2_X4 u5_mult_82_U12297 ( .A1(u5_mult_82_n6887), .A2(u5_mult_82_n6587), 
        .ZN(u5_mult_82_ab_15__25_) );
  NOR2_X4 u5_mult_82_U12296 ( .A1(u5_mult_82_n6859), .A2(u5_mult_82_n6586), 
        .ZN(u5_mult_82_ab_15__30_) );
  NOR2_X4 u5_mult_82_U12295 ( .A1(u5_mult_82_n6840), .A2(u5_mult_82_n6586), 
        .ZN(u5_mult_82_ab_15__33_) );
  NOR2_X4 u5_mult_82_U12294 ( .A1(u5_mult_82_net64905), .A2(u5_mult_82_n6586), 
        .ZN(u5_mult_82_ab_15__35_) );
  NOR2_X4 u5_mult_82_U12293 ( .A1(u5_mult_82_net64923), .A2(u5_mult_82_n6586), 
        .ZN(u5_mult_82_ab_15__36_) );
  NOR2_X4 u5_mult_82_U12292 ( .A1(u5_mult_82_n6833), .A2(u5_mult_82_n6586), 
        .ZN(u5_mult_82_ab_15__39_) );
  NOR2_X4 u5_mult_82_U12291 ( .A1(u5_mult_82_n6829), .A2(u5_mult_82_n6585), 
        .ZN(u5_mult_82_ab_15__40_) );
  NOR2_X4 u5_mult_82_U12290 ( .A1(u5_mult_82_n6818), .A2(u5_mult_82_n6585), 
        .ZN(u5_mult_82_ab_15__42_) );
  NOR2_X4 u5_mult_82_U12289 ( .A1(u5_mult_82_n6799), .A2(u5_mult_82_n6585), 
        .ZN(u5_mult_82_ab_15__45_) );
  NOR2_X4 u5_mult_82_U12288 ( .A1(u5_mult_82_n6793), .A2(u5_mult_82_n6585), 
        .ZN(u5_mult_82_ab_15__46_) );
  NOR2_X4 u5_mult_82_U12287 ( .A1(u5_mult_82_n6786), .A2(u5_mult_82_n6585), 
        .ZN(u5_mult_82_ab_15__47_) );
  NOR2_X4 u5_mult_82_U12286 ( .A1(u5_mult_82_n6780), .A2(u5_mult_82_n6585), 
        .ZN(u5_mult_82_ab_15__48_) );
  NOR2_X4 u5_mult_82_U12285 ( .A1(u5_mult_82_net64383), .A2(u5_mult_82_n6580), 
        .ZN(u5_mult_82_ab_14__6_) );
  NOR2_X4 u5_mult_82_U12284 ( .A1(u5_mult_82_n6942), .A2(u5_mult_82_n6580), 
        .ZN(u5_mult_82_ab_14__7_) );
  NOR2_X4 u5_mult_82_U12283 ( .A1(u5_mult_82_net64491), .A2(u5_mult_82_n6580), 
        .ZN(u5_mult_82_ab_14__12_) );
  NOR2_X4 u5_mult_82_U12282 ( .A1(u5_mult_82_n6935), .A2(u5_mult_82_n6580), 
        .ZN(u5_mult_82_ab_14__15_) );
  NOR2_X4 u5_mult_82_U12281 ( .A1(u5_mult_82_n6929), .A2(u5_mult_82_n6579), 
        .ZN(u5_mult_82_ab_14__17_) );
  NOR2_X4 u5_mult_82_U12280 ( .A1(u5_mult_82_n6922), .A2(u5_mult_82_n6579), 
        .ZN(u5_mult_82_ab_14__18_) );
  NOR2_X4 u5_mult_82_U12279 ( .A1(u5_mult_82_n6906), .A2(u5_mult_82_n6579), 
        .ZN(u5_mult_82_ab_14__20_) );
  NOR2_X4 u5_mult_82_U12278 ( .A1(u5_mult_82_n6833), .A2(u5_mult_82_n6578), 
        .ZN(u5_mult_82_ab_14__39_) );
  NOR2_X4 u5_mult_82_U12277 ( .A1(u5_mult_82_n6823), .A2(u5_mult_82_n6580), 
        .ZN(u5_mult_82_ab_14__41_) );
  NOR2_X4 u5_mult_82_U12276 ( .A1(u5_mult_82_n6806), .A2(u5_mult_82_n6580), 
        .ZN(u5_mult_82_ab_14__44_) );
  NOR2_X4 u5_mult_82_U12275 ( .A1(u5_mult_82_n6775), .A2(u5_mult_82_n6579), 
        .ZN(u5_mult_82_ab_14__49_) );
  NOR2_X4 u5_mult_82_U12274 ( .A1(u5_mult_82_n6762), .A2(u5_mult_82_n6577), 
        .ZN(u5_mult_82_ab_14__51_) );
  NOR2_X4 u5_mult_82_U12273 ( .A1(u5_mult_82_net64383), .A2(u5_mult_82_n6573), 
        .ZN(u5_mult_82_ab_13__6_) );
  NOR2_X4 u5_mult_82_U12272 ( .A1(u5_mult_82_n6942), .A2(u5_mult_82_n6573), 
        .ZN(u5_mult_82_ab_13__7_) );
  NOR2_X4 u5_mult_82_U12271 ( .A1(u5_mult_82_net64419), .A2(u5_mult_82_n6573), 
        .ZN(u5_mult_82_ab_13__8_) );
  NOR2_X4 u5_mult_82_U12270 ( .A1(u5_mult_82_net64437), .A2(u5_mult_82_n6573), 
        .ZN(u5_mult_82_ab_13__9_) );
  NOR2_X4 u5_mult_82_U12269 ( .A1(u5_mult_82_net64509), .A2(u5_mult_82_n6573), 
        .ZN(u5_mult_82_ab_13__13_) );
  NOR2_X4 u5_mult_82_U12268 ( .A1(u5_mult_82_n6935), .A2(u5_mult_82_n6573), 
        .ZN(u5_mult_82_ab_13__15_) );
  NOR2_X4 u5_mult_82_U12267 ( .A1(u5_mult_82_n6922), .A2(u5_mult_82_n6572), 
        .ZN(u5_mult_82_ab_13__18_) );
  NOR2_X4 u5_mult_82_U12266 ( .A1(u5_mult_82_n6906), .A2(u5_mult_82_n6572), 
        .ZN(u5_mult_82_ab_13__20_) );
  NOR2_X4 u5_mult_82_U12265 ( .A1(u5_mult_82_n6898), .A2(u5_mult_82_n6572), 
        .ZN(u5_mult_82_ab_13__21_) );
  NOR2_X4 u5_mult_82_U12264 ( .A1(u5_mult_82_net64671), .A2(u5_mult_82_n6572), 
        .ZN(u5_mult_82_ab_13__22_) );
  NOR2_X4 u5_mult_82_U12263 ( .A1(u5_mult_82_net64689), .A2(u5_mult_82_n6572), 
        .ZN(u5_mult_82_ab_13__23_) );
  NOR2_X4 u5_mult_82_U12262 ( .A1(u5_mult_82_n6893), .A2(u5_mult_82_n6572), 
        .ZN(u5_mult_82_ab_13__24_) );
  NOR2_X4 u5_mult_82_U12261 ( .A1(u5_mult_82_n6887), .A2(u5_mult_82_n6572), 
        .ZN(u5_mult_82_ab_13__25_) );
  NOR2_X4 u5_mult_82_U12260 ( .A1(u5_mult_82_n6845), .A2(u5_mult_82_n6571), 
        .ZN(u5_mult_82_ab_13__32_) );
  NOR2_X4 u5_mult_82_U12259 ( .A1(u5_mult_82_net64887), .A2(u5_mult_82_n6571), 
        .ZN(u5_mult_82_ab_13__34_) );
  NOR2_X4 u5_mult_82_U12258 ( .A1(u5_mult_82_net64941), .A2(u5_mult_82_n6571), 
        .ZN(u5_mult_82_ab_13__37_) );
  NOR2_X4 u5_mult_82_U12257 ( .A1(u5_mult_82_net64959), .A2(u5_mult_82_n6571), 
        .ZN(u5_mult_82_ab_13__38_) );
  NOR2_X4 u5_mult_82_U12256 ( .A1(u5_mult_82_n6818), .A2(u5_mult_82_n6573), 
        .ZN(u5_mult_82_ab_13__42_) );
  NOR2_X4 u5_mult_82_U12255 ( .A1(u5_mult_82_n6813), .A2(u5_mult_82_n6573), 
        .ZN(u5_mult_82_ab_13__43_) );
  NOR2_X4 u5_mult_82_U12254 ( .A1(u5_mult_82_n6806), .A2(u5_mult_82_n6573), 
        .ZN(u5_mult_82_ab_13__44_) );
  NOR2_X4 u5_mult_82_U12253 ( .A1(u5_mult_82_n6799), .A2(u5_mult_82_n6573), 
        .ZN(u5_mult_82_ab_13__45_) );
  NOR2_X4 u5_mult_82_U12252 ( .A1(u5_mult_82_n6780), .A2(u5_mult_82_n6573), 
        .ZN(u5_mult_82_ab_13__48_) );
  NOR2_X4 u5_mult_82_U12251 ( .A1(u5_mult_82_n6762), .A2(u5_mult_82_n6570), 
        .ZN(u5_mult_82_ab_13__51_) );
  NOR2_X4 u5_mult_82_U12250 ( .A1(u5_mult_82_net64419), .A2(u5_mult_82_n6567), 
        .ZN(u5_mult_82_ab_12__8_) );
  NOR2_X4 u5_mult_82_U12249 ( .A1(u5_mult_82_net64437), .A2(u5_mult_82_n6567), 
        .ZN(u5_mult_82_ab_12__9_) );
  NOR2_X4 u5_mult_82_U12248 ( .A1(u5_mult_82_net64491), .A2(u5_mult_82_n6567), 
        .ZN(u5_mult_82_ab_12__12_) );
  NOR2_X4 u5_mult_82_U12247 ( .A1(u5_mult_82_net64509), .A2(u5_mult_82_n6567), 
        .ZN(u5_mult_82_ab_12__13_) );
  NOR2_X4 u5_mult_82_U12246 ( .A1(u5_mult_82_net64527), .A2(u5_mult_82_n6567), 
        .ZN(u5_mult_82_ab_12__14_) );
  NOR2_X4 u5_mult_82_U12245 ( .A1(u5_mult_82_n6922), .A2(u5_mult_82_n6566), 
        .ZN(u5_mult_82_ab_12__18_) );
  NOR2_X4 u5_mult_82_U12244 ( .A1(u5_mult_82_n6915), .A2(u5_mult_82_n6566), 
        .ZN(u5_mult_82_ab_12__19_) );
  NOR2_X4 u5_mult_82_U12243 ( .A1(u5_mult_82_n6898), .A2(u5_mult_82_n6566), 
        .ZN(u5_mult_82_ab_12__21_) );
  NOR2_X4 u5_mult_82_U12242 ( .A1(u5_mult_82_n6887), .A2(u5_mult_82_n6566), 
        .ZN(u5_mult_82_ab_12__25_) );
  NOR2_X4 u5_mult_82_U12241 ( .A1(u5_mult_82_n6882), .A2(u5_mult_82_n6566), 
        .ZN(u5_mult_82_ab_12__26_) );
  NOR2_X4 u5_mult_82_U12240 ( .A1(u5_mult_82_n6864), .A2(u5_mult_82_n6565), 
        .ZN(u5_mult_82_ab_12__29_) );
  NOR2_X4 u5_mult_82_U12239 ( .A1(u5_mult_82_n6859), .A2(u5_mult_82_n6565), 
        .ZN(u5_mult_82_ab_12__30_) );
  NOR2_X4 u5_mult_82_U12238 ( .A1(u5_mult_82_n6845), .A2(u5_mult_82_n6565), 
        .ZN(u5_mult_82_ab_12__32_) );
  NOR2_X4 u5_mult_82_U12237 ( .A1(u5_mult_82_n6840), .A2(u5_mult_82_n6565), 
        .ZN(u5_mult_82_ab_12__33_) );
  NOR2_X4 u5_mult_82_U12236 ( .A1(u5_mult_82_net64905), .A2(u5_mult_82_n6565), 
        .ZN(u5_mult_82_ab_12__35_) );
  NOR2_X4 u5_mult_82_U12235 ( .A1(u5_mult_82_net64941), .A2(u5_mult_82_n6565), 
        .ZN(u5_mult_82_ab_12__37_) );
  NOR2_X4 u5_mult_82_U12234 ( .A1(u5_mult_82_n6833), .A2(u5_mult_82_n6565), 
        .ZN(u5_mult_82_ab_12__39_) );
  NOR2_X4 u5_mult_82_U12233 ( .A1(u5_mult_82_n6829), .A2(u5_mult_82_n6564), 
        .ZN(u5_mult_82_ab_12__40_) );
  NOR2_X4 u5_mult_82_U12232 ( .A1(u5_mult_82_n6823), .A2(u5_mult_82_n6564), 
        .ZN(u5_mult_82_ab_12__41_) );
  NOR2_X4 u5_mult_82_U12231 ( .A1(u5_mult_82_n6818), .A2(u5_mult_82_n6564), 
        .ZN(u5_mult_82_ab_12__42_) );
  NOR2_X4 u5_mult_82_U12230 ( .A1(u5_mult_82_n6806), .A2(u5_mult_82_n6564), 
        .ZN(u5_mult_82_ab_12__44_) );
  NOR2_X4 u5_mult_82_U12229 ( .A1(u5_mult_82_n6799), .A2(u5_mult_82_n6564), 
        .ZN(u5_mult_82_ab_12__45_) );
  NOR2_X4 u5_mult_82_U12228 ( .A1(u5_mult_82_n6786), .A2(u5_mult_82_n6564), 
        .ZN(u5_mult_82_ab_12__47_) );
  NOR2_X4 u5_mult_82_U12227 ( .A1(u5_mult_82_n6769), .A2(u5_mult_82_n6564), 
        .ZN(u5_mult_82_ab_12__50_) );
  NOR2_X4 u5_mult_82_U12226 ( .A1(u5_mult_82_n6762), .A2(u5_mult_82_n6564), 
        .ZN(u5_mult_82_ab_12__51_) );
  INV_X4 u5_mult_82_U12225 ( .A(fracta_mul[12]), .ZN(u5_mult_82_n6995) );
  NOR2_X4 u5_mult_82_U12224 ( .A1(u5_mult_82_net64473), .A2(u5_mult_82_n6559), 
        .ZN(u5_mult_82_ab_11__11_) );
  NOR2_X4 u5_mult_82_U12223 ( .A1(u5_mult_82_n6935), .A2(u5_mult_82_n6559), 
        .ZN(u5_mult_82_ab_11__15_) );
  NOR2_X4 u5_mult_82_U12222 ( .A1(u5_mult_82_net64563), .A2(u5_mult_82_n6558), 
        .ZN(u5_mult_82_ab_11__16_) );
  NOR2_X4 u5_mult_82_U12221 ( .A1(u5_mult_82_n6929), .A2(u5_mult_82_n6558), 
        .ZN(u5_mult_82_ab_11__17_) );
  NOR2_X4 u5_mult_82_U12220 ( .A1(u5_mult_82_n6906), .A2(u5_mult_82_n6558), 
        .ZN(u5_mult_82_ab_11__20_) );
  NOR2_X4 u5_mult_82_U12219 ( .A1(u5_mult_82_net64689), .A2(u5_mult_82_n6558), 
        .ZN(u5_mult_82_ab_11__23_) );
  NOR2_X4 u5_mult_82_U12218 ( .A1(u5_mult_82_n6893), .A2(u5_mult_82_n6558), 
        .ZN(u5_mult_82_ab_11__24_) );
  NOR2_X4 u5_mult_82_U12217 ( .A1(u5_mult_82_n6877), .A2(u5_mult_82_n6558), 
        .ZN(u5_mult_82_ab_11__27_) );
  NOR2_X4 u5_mult_82_U12216 ( .A1(u5_mult_82_n6870), .A2(u5_mult_82_n6557), 
        .ZN(u5_mult_82_ab_11__28_) );
  NOR2_X4 u5_mult_82_U12215 ( .A1(u5_mult_82_n6864), .A2(u5_mult_82_n6557), 
        .ZN(u5_mult_82_ab_11__29_) );
  NOR2_X4 u5_mult_82_U12214 ( .A1(u5_mult_82_n6859), .A2(u5_mult_82_n6557), 
        .ZN(u5_mult_82_ab_11__30_) );
  NOR2_X4 u5_mult_82_U12213 ( .A1(u5_mult_82_n6852), .A2(u5_mult_82_n6557), 
        .ZN(u5_mult_82_ab_11__31_) );
  NOR2_X4 u5_mult_82_U12212 ( .A1(u5_mult_82_net64905), .A2(u5_mult_82_n6557), 
        .ZN(u5_mult_82_ab_11__35_) );
  NOR2_X4 u5_mult_82_U12211 ( .A1(u5_mult_82_net64923), .A2(u5_mult_82_n6557), 
        .ZN(u5_mult_82_ab_11__36_) );
  NOR2_X4 u5_mult_82_U12210 ( .A1(u5_mult_82_n6823), .A2(u5_mult_82_n6559), 
        .ZN(u5_mult_82_ab_11__41_) );
  NOR2_X4 u5_mult_82_U12209 ( .A1(u5_mult_82_n6818), .A2(u5_mult_82_n6559), 
        .ZN(u5_mult_82_ab_11__42_) );
  NOR2_X4 u5_mult_82_U12208 ( .A1(u5_mult_82_n6813), .A2(u5_mult_82_n6559), 
        .ZN(u5_mult_82_ab_11__43_) );
  NOR2_X4 u5_mult_82_U12207 ( .A1(u5_mult_82_n6799), .A2(u5_mult_82_n6559), 
        .ZN(u5_mult_82_ab_11__45_) );
  NOR2_X4 u5_mult_82_U12206 ( .A1(u5_mult_82_n6769), .A2(u5_mult_82_n6557), 
        .ZN(u5_mult_82_ab_11__50_) );
  NOR2_X4 u5_mult_82_U12205 ( .A1(u5_mult_82_n6762), .A2(u5_mult_82_n6556), 
        .ZN(u5_mult_82_ab_11__51_) );
  NOR2_X4 u5_mult_82_U12204 ( .A1(u5_mult_82_net64491), .A2(u5_mult_82_n6552), 
        .ZN(u5_mult_82_ab_10__12_) );
  NOR2_X4 u5_mult_82_U12203 ( .A1(u5_mult_82_n6935), .A2(u5_mult_82_n6552), 
        .ZN(u5_mult_82_ab_10__15_) );
  NOR2_X4 u5_mult_82_U12202 ( .A1(u5_mult_82_n6929), .A2(u5_mult_82_n6551), 
        .ZN(u5_mult_82_ab_10__17_) );
  NOR2_X4 u5_mult_82_U12201 ( .A1(u5_mult_82_n6922), .A2(u5_mult_82_n6551), 
        .ZN(u5_mult_82_ab_10__18_) );
  NOR2_X4 u5_mult_82_U12200 ( .A1(u5_mult_82_n6906), .A2(u5_mult_82_n6551), 
        .ZN(u5_mult_82_ab_10__20_) );
  NOR2_X4 u5_mult_82_U12199 ( .A1(u5_mult_82_n6887), .A2(u5_mult_82_n6551), 
        .ZN(u5_mult_82_ab_10__25_) );
  NOR2_X4 u5_mult_82_U12198 ( .A1(u5_mult_82_n6877), .A2(u5_mult_82_n6551), 
        .ZN(u5_mult_82_ab_10__27_) );
  NOR2_X4 u5_mult_82_U12197 ( .A1(u5_mult_82_n6870), .A2(u5_mult_82_n6550), 
        .ZN(u5_mult_82_ab_10__28_) );
  NOR2_X4 u5_mult_82_U12196 ( .A1(u5_mult_82_n6859), .A2(u5_mult_82_n6550), 
        .ZN(u5_mult_82_ab_10__30_) );
  NOR2_X4 u5_mult_82_U12195 ( .A1(u5_mult_82_n6840), .A2(u5_mult_82_n6550), 
        .ZN(u5_mult_82_ab_10__33_) );
  NOR2_X4 u5_mult_82_U12194 ( .A1(u5_mult_82_net64905), .A2(u5_mult_82_n6550), 
        .ZN(u5_mult_82_ab_10__35_) );
  NOR2_X4 u5_mult_82_U12193 ( .A1(u5_mult_82_net64923), .A2(u5_mult_82_n6550), 
        .ZN(u5_mult_82_ab_10__36_) );
  NOR2_X4 u5_mult_82_U12192 ( .A1(u5_mult_82_net64941), .A2(u5_mult_82_n6550), 
        .ZN(u5_mult_82_ab_10__37_) );
  NOR2_X4 u5_mult_82_U12191 ( .A1(u5_mult_82_n6813), .A2(u5_mult_82_n6552), 
        .ZN(u5_mult_82_ab_10__43_) );
  NOR2_X4 u5_mult_82_U12190 ( .A1(u5_mult_82_n6806), .A2(u5_mult_82_n6552), 
        .ZN(u5_mult_82_ab_10__44_) );
  NOR2_X4 u5_mult_82_U12189 ( .A1(u5_mult_82_n6799), .A2(u5_mult_82_n6552), 
        .ZN(u5_mult_82_ab_10__45_) );
  NOR2_X4 u5_mult_82_U12188 ( .A1(u5_mult_82_n6793), .A2(u5_mult_82_n6552), 
        .ZN(u5_mult_82_ab_10__46_) );
  NOR2_X4 u5_mult_82_U12187 ( .A1(u5_mult_82_n6769), .A2(u5_mult_82_n6553), 
        .ZN(u5_mult_82_ab_10__50_) );
  NOR2_X4 u5_mult_82_U12186 ( .A1(u5_mult_82_n6762), .A2(u5_mult_82_n6549), 
        .ZN(u5_mult_82_ab_10__51_) );
  NOR2_X4 u5_mult_82_U12185 ( .A1(u5_mult_82_net64527), .A2(u5_mult_82_n6546), 
        .ZN(u5_mult_82_ab_9__14_) );
  NOR2_X4 u5_mult_82_U12184 ( .A1(u5_mult_82_net64563), .A2(u5_mult_82_n6545), 
        .ZN(u5_mult_82_ab_9__16_) );
  NOR2_X4 u5_mult_82_U12183 ( .A1(u5_mult_82_n6922), .A2(u5_mult_82_n6545), 
        .ZN(u5_mult_82_ab_9__18_) );
  NOR2_X4 u5_mult_82_U12182 ( .A1(u5_mult_82_n6898), .A2(u5_mult_82_n6545), 
        .ZN(u5_mult_82_ab_9__21_) );
  NOR2_X4 u5_mult_82_U12181 ( .A1(u5_mult_82_n6893), .A2(u5_mult_82_n6545), 
        .ZN(u5_mult_82_ab_9__24_) );
  NOR2_X4 u5_mult_82_U12180 ( .A1(u5_mult_82_n6882), .A2(u5_mult_82_n6545), 
        .ZN(u5_mult_82_ab_9__26_) );
  NOR2_X4 u5_mult_82_U12179 ( .A1(u5_mult_82_n6870), .A2(u5_mult_82_n6544), 
        .ZN(u5_mult_82_ab_9__28_) );
  NOR2_X4 u5_mult_82_U12178 ( .A1(u5_mult_82_n6864), .A2(u5_mult_82_n6544), 
        .ZN(u5_mult_82_ab_9__29_) );
  NOR2_X4 u5_mult_82_U12177 ( .A1(u5_mult_82_n6845), .A2(u5_mult_82_n6544), 
        .ZN(u5_mult_82_ab_9__32_) );
  NOR2_X4 u5_mult_82_U12176 ( .A1(u5_mult_82_n6840), .A2(u5_mult_82_n6544), 
        .ZN(u5_mult_82_ab_9__33_) );
  NOR2_X4 u5_mult_82_U12175 ( .A1(u5_mult_82_net64923), .A2(u5_mult_82_n6544), 
        .ZN(u5_mult_82_ab_9__36_) );
  NOR2_X4 u5_mult_82_U12174 ( .A1(u5_mult_82_n6823), .A2(u5_mult_82_n6543), 
        .ZN(u5_mult_82_ab_9__41_) );
  NOR2_X4 u5_mult_82_U12173 ( .A1(u5_mult_82_n6818), .A2(u5_mult_82_n6543), 
        .ZN(u5_mult_82_ab_9__42_) );
  NOR2_X4 u5_mult_82_U12172 ( .A1(u5_mult_82_n6799), .A2(u5_mult_82_n6543), 
        .ZN(u5_mult_82_ab_9__45_) );
  NOR2_X4 u5_mult_82_U12171 ( .A1(u5_mult_82_n6793), .A2(u5_mult_82_n6543), 
        .ZN(u5_mult_82_ab_9__46_) );
  NOR2_X4 u5_mult_82_U12170 ( .A1(u5_mult_82_n6786), .A2(u5_mult_82_n6543), 
        .ZN(u5_mult_82_ab_9__47_) );
  NOR2_X4 u5_mult_82_U12169 ( .A1(u5_mult_82_n6762), .A2(u5_mult_82_n6543), 
        .ZN(u5_mult_82_ab_9__51_) );
  INV_X4 u5_mult_82_U12168 ( .A(fracta_mul[9]), .ZN(u5_mult_82_n6994) );
  NOR2_X4 u5_mult_82_U12167 ( .A1(u5_mult_82_net64473), .A2(u5_mult_82_n6537), 
        .ZN(u5_mult_82_ab_8__11_) );
  NOR2_X4 u5_mult_82_U12166 ( .A1(u5_mult_82_net64491), .A2(u5_mult_82_n6537), 
        .ZN(u5_mult_82_ab_8__12_) );
  NOR2_X4 u5_mult_82_U12165 ( .A1(u5_mult_82_net64509), .A2(u5_mult_82_n6537), 
        .ZN(u5_mult_82_ab_8__13_) );
  NOR2_X4 u5_mult_82_U12164 ( .A1(u5_mult_82_n6922), .A2(u5_mult_82_n6536), 
        .ZN(u5_mult_82_ab_8__18_) );
  NOR2_X4 u5_mult_82_U12163 ( .A1(u5_mult_82_n6915), .A2(u5_mult_82_n6536), 
        .ZN(u5_mult_82_ab_8__19_) );
  NOR2_X4 u5_mult_82_U12162 ( .A1(u5_mult_82_n6893), .A2(u5_mult_82_n6536), 
        .ZN(u5_mult_82_ab_8__24_) );
  NOR2_X4 u5_mult_82_U12161 ( .A1(u5_mult_82_n6887), .A2(u5_mult_82_n6536), 
        .ZN(u5_mult_82_ab_8__25_) );
  NOR2_X4 u5_mult_82_U12160 ( .A1(u5_mult_82_n6877), .A2(u5_mult_82_n6536), 
        .ZN(u5_mult_82_ab_8__27_) );
  NOR2_X4 u5_mult_82_U12159 ( .A1(u5_mult_82_n6864), .A2(u5_mult_82_n6535), 
        .ZN(u5_mult_82_ab_8__29_) );
  NOR2_X4 u5_mult_82_U12158 ( .A1(u5_mult_82_n6859), .A2(u5_mult_82_n6535), 
        .ZN(u5_mult_82_ab_8__30_) );
  NOR2_X4 u5_mult_82_U12157 ( .A1(u5_mult_82_net64887), .A2(u5_mult_82_n6535), 
        .ZN(u5_mult_82_ab_8__34_) );
  NOR2_X4 u5_mult_82_U12156 ( .A1(u5_mult_82_net64905), .A2(u5_mult_82_n6535), 
        .ZN(u5_mult_82_ab_8__35_) );
  NOR2_X4 u5_mult_82_U12155 ( .A1(u5_mult_82_net64923), .A2(u5_mult_82_n6535), 
        .ZN(u5_mult_82_ab_8__36_) );
  NOR2_X4 u5_mult_82_U12154 ( .A1(u5_mult_82_n6829), .A2(u5_mult_82_n6537), 
        .ZN(u5_mult_82_ab_8__40_) );
  NOR2_X4 u5_mult_82_U12153 ( .A1(u5_mult_82_n6823), .A2(u5_mult_82_n6537), 
        .ZN(u5_mult_82_ab_8__41_) );
  NOR2_X4 u5_mult_82_U12152 ( .A1(u5_mult_82_n6818), .A2(u5_mult_82_n6537), 
        .ZN(u5_mult_82_ab_8__42_) );
  NOR2_X4 u5_mult_82_U12151 ( .A1(u5_mult_82_n6786), .A2(u5_mult_82_n6537), 
        .ZN(u5_mult_82_ab_8__47_) );
  NOR2_X4 u5_mult_82_U12150 ( .A1(u5_mult_82_net64491), .A2(u5_mult_82_n6530), 
        .ZN(u5_mult_82_ab_7__12_) );
  NOR2_X4 u5_mult_82_U12149 ( .A1(u5_mult_82_n6935), .A2(u5_mult_82_n6530), 
        .ZN(u5_mult_82_ab_7__15_) );
  NOR2_X4 u5_mult_82_U12148 ( .A1(u5_mult_82_n6893), .A2(u5_mult_82_n6529), 
        .ZN(u5_mult_82_ab_7__24_) );
  NOR2_X4 u5_mult_82_U12147 ( .A1(u5_mult_82_n6887), .A2(u5_mult_82_n6529), 
        .ZN(u5_mult_82_ab_7__25_) );
  NOR2_X4 u5_mult_82_U12146 ( .A1(u5_mult_82_n6877), .A2(u5_mult_82_n6529), 
        .ZN(u5_mult_82_ab_7__27_) );
  NOR2_X4 u5_mult_82_U12145 ( .A1(u5_mult_82_n6859), .A2(u5_mult_82_n6528), 
        .ZN(u5_mult_82_ab_7__30_) );
  NOR2_X4 u5_mult_82_U12144 ( .A1(u5_mult_82_n6852), .A2(u5_mult_82_n6528), 
        .ZN(u5_mult_82_ab_7__31_) );
  NOR2_X4 u5_mult_82_U12143 ( .A1(u5_mult_82_net64905), .A2(u5_mult_82_n6528), 
        .ZN(u5_mult_82_ab_7__35_) );
  NOR2_X4 u5_mult_82_U12142 ( .A1(u5_mult_82_net64923), .A2(u5_mult_82_n6528), 
        .ZN(u5_mult_82_ab_7__36_) );
  NOR2_X4 u5_mult_82_U12141 ( .A1(u5_mult_82_net64941), .A2(u5_mult_82_n6528), 
        .ZN(u5_mult_82_ab_7__37_) );
  NOR2_X4 u5_mult_82_U12140 ( .A1(u5_mult_82_n6833), .A2(u5_mult_82_n6528), 
        .ZN(u5_mult_82_ab_7__39_) );
  NOR2_X4 u5_mult_82_U12139 ( .A1(u5_mult_82_n6823), .A2(u5_mult_82_n6530), 
        .ZN(u5_mult_82_ab_7__41_) );
  NOR2_X4 u5_mult_82_U12138 ( .A1(u5_mult_82_n6818), .A2(u5_mult_82_n6530), 
        .ZN(u5_mult_82_ab_7__42_) );
  NOR2_X4 u5_mult_82_U12137 ( .A1(u5_mult_82_n6806), .A2(u5_mult_82_n6529), 
        .ZN(u5_mult_82_ab_7__44_) );
  NOR2_X4 u5_mult_82_U12136 ( .A1(u5_mult_82_n6793), .A2(u5_mult_82_n6530), 
        .ZN(u5_mult_82_ab_7__46_) );
  NOR2_X4 u5_mult_82_U12135 ( .A1(u5_mult_82_n6780), .A2(u5_mult_82_n6530), 
        .ZN(u5_mult_82_ab_7__48_) );
  NOR2_X4 u5_mult_82_U12134 ( .A1(u5_mult_82_net64527), .A2(
        u5_mult_82_net66021), .ZN(u5_mult_82_ab_6__14_) );
  NOR2_X4 u5_mult_82_U12133 ( .A1(u5_mult_82_net64563), .A2(
        u5_mult_82_net66019), .ZN(u5_mult_82_ab_6__16_) );
  NOR2_X4 u5_mult_82_U12132 ( .A1(u5_mult_82_n6922), .A2(u5_mult_82_net66019), 
        .ZN(u5_mult_82_ab_6__18_) );
  NOR2_X4 u5_mult_82_U12131 ( .A1(u5_mult_82_n6906), .A2(u5_mult_82_net66019), 
        .ZN(u5_mult_82_ab_6__20_) );
  NOR2_X4 u5_mult_82_U12130 ( .A1(u5_mult_82_n6898), .A2(u5_mult_82_net66019), 
        .ZN(u5_mult_82_ab_6__21_) );
  NOR2_X4 u5_mult_82_U12129 ( .A1(u5_mult_82_n6887), .A2(u5_mult_82_net66019), 
        .ZN(u5_mult_82_ab_6__25_) );
  NOR2_X4 u5_mult_82_U12128 ( .A1(u5_mult_82_n6870), .A2(u5_mult_82_net66017), 
        .ZN(u5_mult_82_ab_6__28_) );
  NOR2_X4 u5_mult_82_U12127 ( .A1(u5_mult_82_n6864), .A2(u5_mult_82_net66017), 
        .ZN(u5_mult_82_ab_6__29_) );
  NOR2_X4 u5_mult_82_U12126 ( .A1(u5_mult_82_n6845), .A2(u5_mult_82_net66017), 
        .ZN(u5_mult_82_ab_6__32_) );
  NOR2_X4 u5_mult_82_U12125 ( .A1(u5_mult_82_net64923), .A2(
        u5_mult_82_net66017), .ZN(u5_mult_82_ab_6__36_) );
  NOR2_X4 u5_mult_82_U12124 ( .A1(u5_mult_82_net64941), .A2(
        u5_mult_82_net66017), .ZN(u5_mult_82_ab_6__37_) );
  NOR2_X4 u5_mult_82_U12123 ( .A1(u5_mult_82_n6833), .A2(u5_mult_82_net66017), 
        .ZN(u5_mult_82_ab_6__39_) );
  NOR2_X4 u5_mult_82_U12122 ( .A1(u5_mult_82_n6813), .A2(u5_mult_82_net66019), 
        .ZN(u5_mult_82_ab_6__43_) );
  NOR2_X4 u5_mult_82_U12121 ( .A1(u5_mult_82_n6806), .A2(u5_mult_82_net66019), 
        .ZN(u5_mult_82_ab_6__44_) );
  NOR2_X4 u5_mult_82_U12120 ( .A1(u5_mult_82_n6799), .A2(u5_mult_82_net66019), 
        .ZN(u5_mult_82_ab_6__45_) );
  NOR2_X4 u5_mult_82_U12119 ( .A1(u5_mult_82_n6786), .A2(u5_mult_82_net66019), 
        .ZN(u5_mult_82_ab_6__47_) );
  NOR2_X4 u5_mult_82_U12118 ( .A1(u5_mult_82_n6780), .A2(u5_mult_82_net66019), 
        .ZN(u5_mult_82_ab_6__48_) );
  NOR2_X4 u5_mult_82_U12117 ( .A1(u5_mult_82_n6915), .A2(u5_mult_82_net66037), 
        .ZN(u5_mult_82_ab_5__19_) );
  NOR2_X4 u5_mult_82_U12116 ( .A1(u5_mult_82_n6898), .A2(u5_mult_82_net66037), 
        .ZN(u5_mult_82_ab_5__21_) );
  NOR2_X4 u5_mult_82_U12115 ( .A1(u5_mult_82_net64671), .A2(
        u5_mult_82_net66037), .ZN(u5_mult_82_ab_5__22_) );
  NOR2_X4 u5_mult_82_U12114 ( .A1(u5_mult_82_net64689), .A2(
        u5_mult_82_net66037), .ZN(u5_mult_82_ab_5__23_) );
  NOR2_X4 u5_mult_82_U12113 ( .A1(u5_mult_82_n6887), .A2(u5_mult_82_net66037), 
        .ZN(u5_mult_82_ab_5__25_) );
  NOR2_X4 u5_mult_82_U12112 ( .A1(u5_mult_82_n6877), .A2(u5_mult_82_net66037), 
        .ZN(u5_mult_82_ab_5__27_) );
  NOR2_X4 u5_mult_82_U12111 ( .A1(u5_mult_82_n6870), .A2(u5_mult_82_net66035), 
        .ZN(u5_mult_82_ab_5__28_) );
  NOR2_X4 u5_mult_82_U12110 ( .A1(u5_mult_82_n6859), .A2(u5_mult_82_net66035), 
        .ZN(u5_mult_82_ab_5__30_) );
  NOR2_X4 u5_mult_82_U12109 ( .A1(u5_mult_82_net64905), .A2(
        u5_mult_82_net66035), .ZN(u5_mult_82_ab_5__35_) );
  NOR2_X4 u5_mult_82_U12108 ( .A1(u5_mult_82_net64923), .A2(
        u5_mult_82_net66035), .ZN(u5_mult_82_ab_5__36_) );
  NOR2_X4 u5_mult_82_U12107 ( .A1(u5_mult_82_net64941), .A2(
        u5_mult_82_net66035), .ZN(u5_mult_82_ab_5__37_) );
  NOR2_X4 u5_mult_82_U12106 ( .A1(u5_mult_82_n6829), .A2(u5_mult_82_net66033), 
        .ZN(u5_mult_82_ab_5__40_) );
  NOR2_X4 u5_mult_82_U12105 ( .A1(u5_mult_82_n6806), .A2(u5_mult_82_net66033), 
        .ZN(u5_mult_82_ab_5__44_) );
  NOR2_X4 u5_mult_82_U12104 ( .A1(u5_mult_82_n6799), .A2(u5_mult_82_net66033), 
        .ZN(u5_mult_82_ab_5__45_) );
  NOR2_X4 u5_mult_82_U12103 ( .A1(u5_mult_82_n6775), .A2(u5_mult_82_net66033), 
        .ZN(u5_mult_82_ab_5__49_) );
  NOR2_X4 u5_mult_82_U12102 ( .A1(u5_mult_82_n6935), .A2(u5_mult_82_n6523), 
        .ZN(u5_mult_82_ab_4__15_) );
  NOR2_X4 u5_mult_82_U12101 ( .A1(u5_mult_82_net64689), .A2(u5_mult_82_n6522), 
        .ZN(u5_mult_82_ab_4__23_) );
  NOR2_X4 u5_mult_82_U12100 ( .A1(u5_mult_82_n6887), .A2(u5_mult_82_n6522), 
        .ZN(u5_mult_82_ab_4__25_) );
  NOR2_X4 u5_mult_82_U12099 ( .A1(u5_mult_82_n6882), .A2(u5_mult_82_n6522), 
        .ZN(u5_mult_82_ab_4__26_) );
  NOR2_X4 u5_mult_82_U12098 ( .A1(u5_mult_82_n6870), .A2(u5_mult_82_n6521), 
        .ZN(u5_mult_82_ab_4__28_) );
  NOR2_X4 u5_mult_82_U12097 ( .A1(u5_mult_82_n6864), .A2(u5_mult_82_n6521), 
        .ZN(u5_mult_82_ab_4__29_) );
  NOR2_X4 u5_mult_82_U12096 ( .A1(u5_mult_82_n6840), .A2(u5_mult_82_n6521), 
        .ZN(u5_mult_82_ab_4__33_) );
  NOR2_X4 u5_mult_82_U12095 ( .A1(u5_mult_82_net64905), .A2(u5_mult_82_n6521), 
        .ZN(u5_mult_82_ab_4__35_) );
  NOR2_X4 u5_mult_82_U12094 ( .A1(u5_mult_82_net64923), .A2(u5_mult_82_n6521), 
        .ZN(u5_mult_82_ab_4__36_) );
  NOR2_X4 u5_mult_82_U12093 ( .A1(u5_mult_82_net64941), .A2(u5_mult_82_n6521), 
        .ZN(u5_mult_82_ab_4__37_) );
  NOR2_X4 u5_mult_82_U12092 ( .A1(u5_mult_82_n6833), .A2(u5_mult_82_n6521), 
        .ZN(u5_mult_82_ab_4__39_) );
  NOR2_X4 u5_mult_82_U12091 ( .A1(u5_mult_82_n6823), .A2(u5_mult_82_n6520), 
        .ZN(u5_mult_82_ab_4__41_) );
  NOR2_X4 u5_mult_82_U12090 ( .A1(u5_mult_82_n6793), .A2(u5_mult_82_n6520), 
        .ZN(u5_mult_82_ab_4__46_) );
  INV_X4 u5_mult_82_U12089 ( .A(fracta_mul[4]), .ZN(u5_mult_82_n6993) );
  NOR2_X4 u5_mult_82_U12088 ( .A1(u5_mult_82_net64509), .A2(u5_mult_82_n6516), 
        .ZN(u5_mult_82_ab_3__13_) );
  NOR2_X4 u5_mult_82_U12087 ( .A1(u5_mult_82_net64527), .A2(u5_mult_82_n6516), 
        .ZN(u5_mult_82_ab_3__14_) );
  NOR2_X4 u5_mult_82_U12086 ( .A1(u5_mult_82_n6935), .A2(u5_mult_82_n6516), 
        .ZN(u5_mult_82_ab_3__15_) );
  NOR2_X4 u5_mult_82_U12085 ( .A1(u5_mult_82_n6929), .A2(u5_mult_82_n6515), 
        .ZN(u5_mult_82_ab_3__17_) );
  NOR2_X4 u5_mult_82_U12084 ( .A1(u5_mult_82_n6887), .A2(u5_mult_82_n6515), 
        .ZN(u5_mult_82_ab_3__25_) );
  NOR2_X4 u5_mult_82_U12083 ( .A1(u5_mult_82_n6882), .A2(u5_mult_82_n6515), 
        .ZN(u5_mult_82_ab_3__26_) );
  NOR2_X4 u5_mult_82_U12082 ( .A1(u5_mult_82_n6870), .A2(u5_mult_82_n6514), 
        .ZN(u5_mult_82_ab_3__28_) );
  NOR2_X4 u5_mult_82_U12081 ( .A1(u5_mult_82_n6864), .A2(u5_mult_82_n6514), 
        .ZN(u5_mult_82_ab_3__29_) );
  NOR2_X4 u5_mult_82_U12080 ( .A1(u5_mult_82_n6852), .A2(u5_mult_82_n6514), 
        .ZN(u5_mult_82_ab_3__31_) );
  NOR2_X4 u5_mult_82_U12079 ( .A1(u5_mult_82_net64887), .A2(u5_mult_82_n6514), 
        .ZN(u5_mult_82_ab_3__34_) );
  NOR2_X4 u5_mult_82_U12078 ( .A1(u5_mult_82_net64905), .A2(u5_mult_82_n6514), 
        .ZN(u5_mult_82_ab_3__35_) );
  NOR2_X4 u5_mult_82_U12077 ( .A1(u5_mult_82_net64923), .A2(u5_mult_82_n6514), 
        .ZN(u5_mult_82_ab_3__36_) );
  NOR2_X4 u5_mult_82_U12076 ( .A1(u5_mult_82_net64959), .A2(u5_mult_82_n6514), 
        .ZN(u5_mult_82_ab_3__38_) );
  NOR2_X4 u5_mult_82_U12075 ( .A1(u5_mult_82_n6833), .A2(u5_mult_82_n6514), 
        .ZN(u5_mult_82_ab_3__39_) );
  NOR2_X4 u5_mult_82_U12074 ( .A1(u5_mult_82_n6829), .A2(u5_mult_82_n6513), 
        .ZN(u5_mult_82_ab_3__40_) );
  NOR2_X4 u5_mult_82_U12073 ( .A1(u5_mult_82_n6823), .A2(u5_mult_82_n6513), 
        .ZN(u5_mult_82_ab_3__41_) );
  NOR2_X4 u5_mult_82_U12072 ( .A1(u5_mult_82_n6793), .A2(u5_mult_82_n6513), 
        .ZN(u5_mult_82_ab_3__46_) );
  NOR2_X4 u5_mult_82_U12071 ( .A1(u5_mult_82_n6786), .A2(u5_mult_82_n6513), 
        .ZN(u5_mult_82_ab_3__47_) );
  NOR2_X4 u5_mult_82_U12070 ( .A1(u5_mult_82_n6769), .A2(u5_mult_82_n6513), 
        .ZN(u5_mult_82_ab_3__50_) );
  NOR2_X4 u5_mult_82_U12069 ( .A1(u5_mult_82_net64489), .A2(
        u5_mult_82_net66093), .ZN(u5_mult_82_ab_2__12_) );
  NOR2_X4 u5_mult_82_U12068 ( .A1(u5_mult_82_net64511), .A2(
        u5_mult_82_net66093), .ZN(u5_mult_82_ab_2__13_) );
  NOR2_X4 u5_mult_82_U12067 ( .A1(u5_mult_82_net64525), .A2(
        u5_mult_82_net66093), .ZN(u5_mult_82_ab_2__14_) );
  NOR2_X4 u5_mult_82_U12066 ( .A1(u5_mult_82_n6936), .A2(u5_mult_82_net66093), 
        .ZN(u5_mult_82_ab_2__15_) );
  NOR2_X4 u5_mult_82_U12065 ( .A1(u5_mult_82_n6914), .A2(u5_mult_82_net66091), 
        .ZN(u5_mult_82_ab_2__19_) );
  NOR2_X4 u5_mult_82_U12064 ( .A1(u5_mult_82_n6899), .A2(u5_mult_82_net66091), 
        .ZN(u5_mult_82_ab_2__21_) );
  NOR2_X4 u5_mult_82_U12063 ( .A1(u5_mult_82_n6882), .A2(u5_mult_82_net66091), 
        .ZN(u5_mult_82_ab_2__26_) );
  NOR2_X4 u5_mult_82_U12062 ( .A1(u5_mult_82_n6876), .A2(u5_mult_82_net66091), 
        .ZN(u5_mult_82_ab_2__27_) );
  NOR2_X4 u5_mult_82_U12061 ( .A1(u5_mult_82_n6870), .A2(u5_mult_82_net66089), 
        .ZN(u5_mult_82_ab_2__28_) );
  NOR2_X4 u5_mult_82_U12060 ( .A1(u5_mult_82_n6864), .A2(u5_mult_82_net66089), 
        .ZN(u5_mult_82_ab_2__29_) );
  NOR2_X4 u5_mult_82_U12059 ( .A1(u5_mult_82_n6859), .A2(u5_mult_82_net66089), 
        .ZN(u5_mult_82_ab_2__30_) );
  NOR2_X4 u5_mult_82_U12058 ( .A1(u5_mult_82_n6846), .A2(u5_mult_82_net66089), 
        .ZN(u5_mult_82_ab_2__32_) );
  NOR2_X4 u5_mult_82_U12057 ( .A1(u5_mult_82_net64943), .A2(
        u5_mult_82_net66089), .ZN(u5_mult_82_ab_2__37_) );
  NOR2_X4 u5_mult_82_U12056 ( .A1(u5_mult_82_n6818), .A2(u5_mult_82_net66087), 
        .ZN(u5_mult_82_ab_2__42_) );
  NOR2_X4 u5_mult_82_U12055 ( .A1(u5_mult_82_n6786), .A2(u5_mult_82_net66087), 
        .ZN(u5_mult_82_ab_2__47_) );
  NOR2_X4 u5_mult_82_U12054 ( .A1(u5_mult_82_n6762), .A2(u5_mult_82_net66087), 
        .ZN(u5_mult_82_ab_2__51_) );
  NOR2_X4 u5_mult_82_U12053 ( .A1(u5_mult_82_n6985), .A2(u5_mult_82_net66111), 
        .ZN(u5_mult_82_ab_1__0_) );
  NOR2_X4 u5_mult_82_U12052 ( .A1(u5_mult_82_n6966), .A2(u5_mult_82_net66111), 
        .ZN(u5_mult_82_ab_1__1_) );
  NOR2_X4 u5_mult_82_U12051 ( .A1(u5_mult_82_n6959), .A2(u5_mult_82_net66111), 
        .ZN(u5_mult_82_ab_1__2_) );
  NOR2_X4 u5_mult_82_U12050 ( .A1(u5_mult_82_n6952), .A2(u5_mult_82_net66111), 
        .ZN(u5_mult_82_ab_1__3_) );
  NOR2_X4 u5_mult_82_U12049 ( .A1(u5_mult_82_n6945), .A2(u5_mult_82_net66111), 
        .ZN(u5_mult_82_ab_1__4_) );
  NOR2_X4 u5_mult_82_U12048 ( .A1(u5_mult_82_net64373), .A2(
        u5_mult_82_net66111), .ZN(u5_mult_82_ab_1__5_) );
  NOR2_X4 u5_mult_82_U12047 ( .A1(u5_mult_82_n1271), .A2(u5_mult_82_net66111), 
        .ZN(u5_mult_82_ab_1__6_) );
  NOR2_X4 u5_mult_82_U12046 ( .A1(u5_mult_82_n6939), .A2(u5_mult_82_net66111), 
        .ZN(u5_mult_82_ab_1__7_) );
  NOR2_X4 u5_mult_82_U12045 ( .A1(u5_mult_82_net64427), .A2(
        u5_mult_82_net66111), .ZN(u5_mult_82_ab_1__8_) );
  NOR2_X4 u5_mult_82_U12044 ( .A1(u5_mult_82_net64223), .A2(u5_mult_82_n1289), 
        .ZN(u5_mult_82_ab_0__9_) );
  NOR2_X4 u5_mult_82_U12043 ( .A1(u5_mult_82_n1289), .A2(u5_mult_82_net66111), 
        .ZN(u5_mult_82_ab_1__9_) );
  NOR2_X4 u5_mult_82_U12042 ( .A1(u5_mult_82_n1373), .A2(u5_mult_82_net66111), 
        .ZN(u5_mult_82_ab_1__10_) );
  NOR2_X4 u5_mult_82_U12041 ( .A1(u5_mult_82_n1319), .A2(u5_mult_82_net66111), 
        .ZN(u5_mult_82_ab_1__11_) );
  NOR2_X4 u5_mult_82_U12040 ( .A1(u5_mult_82_net64223), .A2(
        u5_mult_82_net64499), .ZN(u5_mult_82_ab_0__12_) );
  NOR2_X4 u5_mult_82_U12039 ( .A1(u5_mult_82_net64499), .A2(
        u5_mult_82_net66111), .ZN(u5_mult_82_ab_1__12_) );
  NOR2_X4 u5_mult_82_U12038 ( .A1(u5_mult_82_net64223), .A2(
        u5_mult_82_net64517), .ZN(u5_mult_82_ab_0__13_) );
  NOR2_X4 u5_mult_82_U12037 ( .A1(u5_mult_82_net64517), .A2(
        u5_mult_82_net66111), .ZN(u5_mult_82_ab_1__13_) );
  NOR2_X4 u5_mult_82_U12036 ( .A1(u5_mult_82_net64535), .A2(
        u5_mult_82_net66111), .ZN(u5_mult_82_ab_1__14_) );
  NOR2_X4 u5_mult_82_U12035 ( .A1(u5_mult_82_n6932), .A2(u5_mult_82_net66111), 
        .ZN(u5_mult_82_ab_1__15_) );
  NOR2_X4 u5_mult_82_U12034 ( .A1(u5_mult_82_net64571), .A2(
        u5_mult_82_net66109), .ZN(u5_mult_82_ab_1__16_) );
  NOR2_X4 u5_mult_82_U12033 ( .A1(u5_mult_82_n6926), .A2(u5_mult_82_net66109), 
        .ZN(u5_mult_82_ab_1__17_) );
  NOR2_X4 u5_mult_82_U12032 ( .A1(u5_mult_82_net64219), .A2(u5_mult_82_n6919), 
        .ZN(u5_mult_82_ab_0__18_) );
  NOR2_X4 u5_mult_82_U12031 ( .A1(u5_mult_82_n6919), .A2(u5_mult_82_net66109), 
        .ZN(u5_mult_82_ab_1__18_) );
  INV_X4 u5_mult_82_U12030 ( .A(n4725), .ZN(u5_mult_82_n7021) );
  NOR2_X4 u5_mult_82_U12029 ( .A1(u5_mult_82_net64219), .A2(u5_mult_82_n6912), 
        .ZN(u5_mult_82_ab_0__19_) );
  NOR2_X4 u5_mult_82_U12028 ( .A1(u5_mult_82_n6912), .A2(u5_mult_82_net66109), 
        .ZN(u5_mult_82_ab_1__19_) );
  NOR2_X4 u5_mult_82_U12027 ( .A1(u5_mult_82_net64219), .A2(u5_mult_82_n6903), 
        .ZN(u5_mult_82_ab_0__20_) );
  NOR2_X4 u5_mult_82_U12026 ( .A1(u5_mult_82_n6903), .A2(u5_mult_82_net66109), 
        .ZN(u5_mult_82_ab_1__20_) );
  NOR2_X4 u5_mult_82_U12025 ( .A1(u5_mult_82_net64219), .A2(u5_mult_82_n6895), 
        .ZN(u5_mult_82_ab_0__21_) );
  NOR2_X4 u5_mult_82_U12024 ( .A1(u5_mult_82_n6895), .A2(u5_mult_82_net66109), 
        .ZN(u5_mult_82_ab_1__21_) );
  NOR2_X4 u5_mult_82_U12023 ( .A1(u5_mult_82_net64219), .A2(
        u5_mult_82_net64665), .ZN(u5_mult_82_ab_0__22_) );
  NOR2_X4 u5_mult_82_U12022 ( .A1(u5_mult_82_net64665), .A2(
        u5_mult_82_net66109), .ZN(u5_mult_82_ab_1__22_) );
  NOR2_X4 u5_mult_82_U12021 ( .A1(u5_mult_82_net64219), .A2(
        u5_mult_82_net64683), .ZN(u5_mult_82_ab_0__23_) );
  NOR2_X4 u5_mult_82_U12020 ( .A1(u5_mult_82_net64683), .A2(
        u5_mult_82_net66109), .ZN(u5_mult_82_ab_1__23_) );
  NOR2_X4 u5_mult_82_U12019 ( .A1(u5_mult_82_net64219), .A2(u5_mult_82_n7019), 
        .ZN(u5_mult_82_ab_0__24_) );
  NOR2_X4 u5_mult_82_U12018 ( .A1(u5_mult_82_n7019), .A2(u5_mult_82_net66109), 
        .ZN(u5_mult_82_ab_1__24_) );
  NOR2_X4 u5_mult_82_U12017 ( .A1(u5_mult_82_net64219), .A2(u5_mult_82_n6884), 
        .ZN(u5_mult_82_ab_0__25_) );
  NOR2_X4 u5_mult_82_U12016 ( .A1(u5_mult_82_n6884), .A2(u5_mult_82_net66109), 
        .ZN(u5_mult_82_ab_1__25_) );
  NOR2_X4 u5_mult_82_U12015 ( .A1(u5_mult_82_net64219), .A2(u5_mult_82_n6879), 
        .ZN(u5_mult_82_ab_0__26_) );
  NOR2_X4 u5_mult_82_U12014 ( .A1(u5_mult_82_n6879), .A2(u5_mult_82_net66109), 
        .ZN(u5_mult_82_ab_1__26_) );
  NOR2_X4 u5_mult_82_U12013 ( .A1(u5_mult_82_net64219), .A2(u5_mult_82_n6874), 
        .ZN(u5_mult_82_ab_0__27_) );
  NOR2_X4 u5_mult_82_U12012 ( .A1(u5_mult_82_n6874), .A2(u5_mult_82_net66109), 
        .ZN(u5_mult_82_ab_1__27_) );
  NOR2_X4 u5_mult_82_U12011 ( .A1(u5_mult_82_net64219), .A2(u5_mult_82_n6867), 
        .ZN(u5_mult_82_ab_0__28_) );
  NOR2_X4 u5_mult_82_U12010 ( .A1(u5_mult_82_n6867), .A2(u5_mult_82_n1262), 
        .ZN(u5_mult_82_ab_1__28_) );
  NOR2_X4 u5_mult_82_U12009 ( .A1(u5_mult_82_net64219), .A2(u5_mult_82_n6861), 
        .ZN(u5_mult_82_ab_0__29_) );
  NOR2_X4 u5_mult_82_U12008 ( .A1(u5_mult_82_n6861), .A2(u5_mult_82_n1262), 
        .ZN(u5_mult_82_ab_1__29_) );
  NOR2_X4 u5_mult_82_U12007 ( .A1(u5_mult_82_net64219), .A2(u5_mult_82_n6856), 
        .ZN(u5_mult_82_ab_0__30_) );
  NOR2_X4 u5_mult_82_U12006 ( .A1(u5_mult_82_n6856), .A2(u5_mult_82_n1262), 
        .ZN(u5_mult_82_ab_1__30_) );
  NOR2_X4 u5_mult_82_U12005 ( .A1(u5_mult_82_net64219), .A2(u5_mult_82_n6837), 
        .ZN(u5_mult_82_ab_0__33_) );
  NOR2_X4 u5_mult_82_U12004 ( .A1(u5_mult_82_n6837), .A2(u5_mult_82_n1262), 
        .ZN(u5_mult_82_ab_1__33_) );
  NOR2_X4 u5_mult_82_U12003 ( .A1(u5_mult_82_net64219), .A2(
        u5_mult_82_net64881), .ZN(u5_mult_82_ab_0__34_) );
  NOR2_X4 u5_mult_82_U12002 ( .A1(u5_mult_82_net64881), .A2(u5_mult_82_n1262), 
        .ZN(u5_mult_82_ab_1__34_) );
  NOR2_X4 u5_mult_82_U12001 ( .A1(u5_mult_82_net64219), .A2(
        u5_mult_82_net64913), .ZN(u5_mult_82_ab_0__35_) );
  NOR2_X4 u5_mult_82_U12000 ( .A1(u5_mult_82_net64217), .A2(u5_mult_82_n6826), 
        .ZN(u5_mult_82_ab_0__40_) );
  NOR2_X4 u5_mult_82_U11999 ( .A1(u5_mult_82_net64217), .A2(u5_mult_82_n6810), 
        .ZN(u5_mult_82_ab_0__43_) );
  NOR2_X4 u5_mult_82_U11998 ( .A1(u5_mult_82_net66107), .A2(u5_mult_82_n7008), 
        .ZN(u5_mult_82_ab_1__45_) );
  NOR2_X4 u5_mult_82_U11997 ( .A1(u5_mult_82_net64217), .A2(u5_mult_82_n6777), 
        .ZN(u5_mult_82_ab_0__48_) );
  NOR2_X4 u5_mult_82_U11996 ( .A1(u5_mult_82_net64217), .A2(u5_mult_82_n6766), 
        .ZN(u5_mult_82_ab_0__50_) );
  NOR2_X4 u5_mult_82_U11995 ( .A1(u5_mult_82_n6766), .A2(u5_mult_82_net66107), 
        .ZN(u5_mult_82_ab_1__50_) );
  NOR2_X4 u5_mult_82_U11994 ( .A1(u5_mult_82_net64217), .A2(u5_mult_82_n6759), 
        .ZN(u5_mult_82_ab_0__51_) );
  INV_X32 u5_mult_82_U11993 ( .A(u5_mult_82_net64225), .ZN(u5_mult_82_net64219) );
  INV_X32 u5_mult_82_U11992 ( .A(u5_mult_82_n6990), .ZN(u5_mult_82_n6989) );
  INV_X32 u5_mult_82_U11991 ( .A(u5_mult_82_n6990), .ZN(u5_mult_82_n6988) );
  INV_X32 u5_mult_82_U11990 ( .A(u5_mult_82_n6991), .ZN(u5_mult_82_n6987) );
  INV_X32 u5_mult_82_U11989 ( .A(u5_mult_82_n6991), .ZN(u5_mult_82_n6986) );
  INV_X32 u5_mult_82_U11988 ( .A(u5_mult_82_n6971), .ZN(u5_mult_82_n6969) );
  INV_X32 u5_mult_82_U11987 ( .A(u5_mult_82_n6971), .ZN(u5_mult_82_n6968) );
  INV_X32 u5_mult_82_U11986 ( .A(u5_mult_82_n6972), .ZN(u5_mult_82_n6967) );
  INV_X32 u5_mult_82_U11985 ( .A(u5_mult_82_n6964), .ZN(u5_mult_82_n6962) );
  INV_X32 u5_mult_82_U11984 ( .A(u5_mult_82_n6964), .ZN(u5_mult_82_n6961) );
  INV_X32 u5_mult_82_U11983 ( .A(u5_mult_82_n6951), .ZN(u5_mult_82_n6958) );
  INV_X32 u5_mult_82_U11982 ( .A(u5_mult_82_n6951), .ZN(u5_mult_82_n6957) );
  INV_X32 u5_mult_82_U11981 ( .A(u5_mult_82_n6957), .ZN(u5_mult_82_n6955) );
  INV_X32 u5_mult_82_U11980 ( .A(u5_mult_82_n6957), .ZN(u5_mult_82_n6954) );
  INV_X32 u5_mult_82_U11979 ( .A(u5_mult_82_n6958), .ZN(u5_mult_82_n6953) );
  INV_X32 u5_mult_82_U11978 ( .A(u5_mult_82_n6958), .ZN(u5_mult_82_n6952) );
  INV_X32 u5_mult_82_U11977 ( .A(u6_N3), .ZN(u5_mult_82_n6951) );
  INV_X32 u5_mult_82_U11976 ( .A(u5_mult_82_n6945), .ZN(u5_mult_82_n6949) );
  INV_X32 u5_mult_82_U11975 ( .A(u5_mult_82_n6949), .ZN(u5_mult_82_n6948) );
  INV_X32 u5_mult_82_U11974 ( .A(u5_mult_82_n6949), .ZN(u5_mult_82_n6947) );
  INV_X32 u5_mult_82_U11973 ( .A(u5_mult_82_n6950), .ZN(u5_mult_82_n6946) );
  INV_X32 u5_mult_82_U11972 ( .A(u5_mult_82_net64373), .ZN(u5_mult_82_net64369) );
  INV_X32 u5_mult_82_U11971 ( .A(u5_mult_82_net64369), .ZN(u5_mult_82_net64365) );
  INV_X32 u5_mult_82_U11970 ( .A(u5_mult_82_net64369), .ZN(u5_mult_82_net64363) );
  INV_X32 u5_mult_82_U11969 ( .A(u5_mult_82_net64371), .ZN(u5_mult_82_net64361) );
  INV_X32 u5_mult_82_U11968 ( .A(u5_mult_82_net64387), .ZN(u5_mult_82_net64383) );
  INV_X32 u5_mult_82_U11967 ( .A(u5_mult_82_net64387), .ZN(u5_mult_82_net64381) );
  INV_X32 u5_mult_82_U11966 ( .A(u5_mult_82_n6939), .ZN(u5_mult_82_n6943) );
  INV_X32 u5_mult_82_U11965 ( .A(u5_mult_82_n6943), .ZN(u5_mult_82_n6942) );
  INV_X32 u5_mult_82_U11964 ( .A(u5_mult_82_n6943), .ZN(u5_mult_82_n6941) );
  INV_X32 u5_mult_82_U11963 ( .A(u5_mult_82_n6944), .ZN(u5_mult_82_n6940) );
  INV_X32 u5_mult_82_U11962 ( .A(u5_mult_82_net64423), .ZN(u5_mult_82_net64419) );
  INV_X32 u5_mult_82_U11961 ( .A(u5_mult_82_net64423), .ZN(u5_mult_82_net64417) );
  INV_X32 u5_mult_82_U11960 ( .A(u5_mult_82_net64425), .ZN(u5_mult_82_net64415) );
  INV_X32 u5_mult_82_U11959 ( .A(u5_mult_82_net64441), .ZN(u5_mult_82_net64437) );
  INV_X32 u5_mult_82_U11958 ( .A(u5_mult_82_net64441), .ZN(u5_mult_82_net64435) );
  INV_X32 u5_mult_82_U11957 ( .A(u5_mult_82_net64459), .ZN(u5_mult_82_net64455) );
  INV_X32 u5_mult_82_U11956 ( .A(u5_mult_82_net64477), .ZN(u5_mult_82_net64473) );
  INV_X32 u5_mult_82_U11955 ( .A(u5_mult_82_net64477), .ZN(u5_mult_82_net64471) );
  INV_X32 u5_mult_82_U11954 ( .A(u5_mult_82_net64513), .ZN(u5_mult_82_net64509) );
  INV_X32 u5_mult_82_U11953 ( .A(u5_mult_82_net64513), .ZN(u5_mult_82_net64507) );
  INV_X32 u5_mult_82_U11952 ( .A(u5_mult_82_net64531), .ZN(u5_mult_82_net64527) );
  INV_X32 u5_mult_82_U11951 ( .A(u5_mult_82_net64531), .ZN(u5_mult_82_net64525) );
  INV_X32 u5_mult_82_U11950 ( .A(u5_mult_82_net64533), .ZN(u5_mult_82_net64523) );
  INV_X32 u5_mult_82_U11949 ( .A(u5_mult_82_n6937), .ZN(u5_mult_82_n6934) );
  INV_X32 u5_mult_82_U11948 ( .A(u5_mult_82_n6938), .ZN(u5_mult_82_n6933) );
  INV_X32 u5_mult_82_U11947 ( .A(u5_mult_82_net64567), .ZN(u5_mult_82_net64563) );
  INV_X32 u5_mult_82_U11946 ( .A(u5_mult_82_net64567), .ZN(u5_mult_82_net64561) );
  INV_X32 u5_mult_82_U11945 ( .A(u5_mult_82_n6930), .ZN(u5_mult_82_n6928) );
  INV_X32 u5_mult_82_U11944 ( .A(u5_mult_82_n6931), .ZN(u5_mult_82_n6927) );
  INV_X32 u5_mult_82_U11943 ( .A(u5_mult_82_n6917), .ZN(u5_mult_82_n6925) );
  INV_X32 u5_mult_82_U11942 ( .A(u5_mult_82_n6917), .ZN(u5_mult_82_n6924) );
  INV_X32 u5_mult_82_U11941 ( .A(u5_mult_82_n6924), .ZN(u5_mult_82_n6922) );
  INV_X32 u5_mult_82_U11940 ( .A(u5_mult_82_n6924), .ZN(u5_mult_82_n6921) );
  INV_X32 u5_mult_82_U11939 ( .A(u5_mult_82_n6925), .ZN(u5_mult_82_n6920) );
  INV_X32 u5_mult_82_U11938 ( .A(u5_mult_82_n6925), .ZN(u5_mult_82_n6919) );
  INV_X32 u5_mult_82_U11937 ( .A(u5_mult_82_n6918), .ZN(u5_mult_82_n6917) );
  INV_X32 u5_mult_82_U11936 ( .A(u5_mult_82_n6910), .ZN(u5_mult_82_n6916) );
  INV_X32 u5_mult_82_U11935 ( .A(u5_mult_82_n6916), .ZN(u5_mult_82_n6915) );
  INV_X32 u5_mult_82_U11934 ( .A(u5_mult_82_n6916), .ZN(u5_mult_82_n6914) );
  INV_X32 u5_mult_82_U11933 ( .A(u5_mult_82_n6916), .ZN(u5_mult_82_n6913) );
  INV_X32 u5_mult_82_U11932 ( .A(u5_mult_82_n6911), .ZN(u5_mult_82_n6912) );
  INV_X32 u5_mult_82_U11931 ( .A(u5_mult_82_n6911), .ZN(u5_mult_82_n6910) );
  INV_X32 u5_mult_82_U11930 ( .A(u5_mult_82_n6902), .ZN(u5_mult_82_n6909) );
  INV_X32 u5_mult_82_U11929 ( .A(u5_mult_82_n6902), .ZN(u5_mult_82_n6908) );
  INV_X32 u5_mult_82_U11928 ( .A(u5_mult_82_n6908), .ZN(u5_mult_82_n6906) );
  INV_X32 u5_mult_82_U11927 ( .A(u5_mult_82_n6908), .ZN(u5_mult_82_n6905) );
  INV_X32 u5_mult_82_U11926 ( .A(u5_mult_82_n6909), .ZN(u5_mult_82_n6904) );
  INV_X32 u5_mult_82_U11925 ( .A(u5_mult_82_n6909), .ZN(u5_mult_82_n6903) );
  INV_X32 u5_mult_82_U11924 ( .A(u5_mult_82_n6894), .ZN(u5_mult_82_n6900) );
  INV_X32 u5_mult_82_U11923 ( .A(u5_mult_82_n6900), .ZN(u5_mult_82_n6898) );
  INV_X32 u5_mult_82_U11922 ( .A(u5_mult_82_n6900), .ZN(u5_mult_82_n6897) );
  INV_X32 u5_mult_82_U11921 ( .A(u5_mult_82_n6901), .ZN(u5_mult_82_n6896) );
  INV_X32 u5_mult_82_U11920 ( .A(u5_mult_82_n6901), .ZN(u5_mult_82_n6895) );
  INV_X32 u5_mult_82_U11919 ( .A(u5_mult_82_net64677), .ZN(u5_mult_82_net64667) );
  INV_X32 u5_mult_82_U11918 ( .A(u5_mult_82_net64677), .ZN(u5_mult_82_net64665) );
  INV_X32 u5_mult_82_U11917 ( .A(u5_mult_82_net64695), .ZN(u5_mult_82_net64685) );
  INV_X32 u5_mult_82_U11916 ( .A(u5_mult_82_net64695), .ZN(u5_mult_82_net64683) );
  INV_X32 u5_mult_82_U11915 ( .A(u5_mult_82_n6890), .ZN(u5_mult_82_n6893) );
  INV_X32 u5_mult_82_U11914 ( .A(u5_mult_82_n6890), .ZN(u5_mult_82_n6892) );
  INV_X32 u5_mult_82_U11913 ( .A(u5_mult_82_n6890), .ZN(u5_mult_82_n6891) );
  INV_X32 u5_mult_82_U11912 ( .A(u5_mult_82_n6888), .ZN(u5_mult_82_n6887) );
  INV_X32 u5_mult_82_U11911 ( .A(u5_mult_82_n6888), .ZN(u5_mult_82_n6886) );
  INV_X32 u5_mult_82_U11910 ( .A(u5_mult_82_n6889), .ZN(u5_mult_82_n6885) );
  INV_X32 u5_mult_82_U11909 ( .A(u5_mult_82_n6889), .ZN(u5_mult_82_n6884) );
  INV_X32 u5_mult_82_U11908 ( .A(u5_mult_82_n7017), .ZN(u5_mult_82_n6883) );
  INV_X32 u5_mult_82_U11907 ( .A(u5_mult_82_n6883), .ZN(u5_mult_82_n6882) );
  INV_X32 u5_mult_82_U11906 ( .A(u5_mult_82_n6883), .ZN(u5_mult_82_n6881) );
  INV_X32 u5_mult_82_U11905 ( .A(u5_mult_82_n6883), .ZN(u5_mult_82_n6880) );
  INV_X32 u5_mult_82_U11904 ( .A(u5_mult_82_n6883), .ZN(u5_mult_82_n6879) );
  INV_X32 u5_mult_82_U11903 ( .A(u5_mult_82_n6872), .ZN(u5_mult_82_n6878) );
  INV_X32 u5_mult_82_U11902 ( .A(u5_mult_82_n6878), .ZN(u5_mult_82_n6877) );
  INV_X32 u5_mult_82_U11901 ( .A(u5_mult_82_n6878), .ZN(u5_mult_82_n6876) );
  INV_X32 u5_mult_82_U11900 ( .A(u5_mult_82_n6878), .ZN(u5_mult_82_n6875) );
  INV_X32 u5_mult_82_U11899 ( .A(u5_mult_82_n6873), .ZN(u5_mult_82_n6874) );
  INV_X32 u5_mult_82_U11898 ( .A(u5_mult_82_n7015), .ZN(u5_mult_82_n6871) );
  INV_X32 u5_mult_82_U11897 ( .A(u5_mult_82_n6871), .ZN(u5_mult_82_n6870) );
  INV_X32 u5_mult_82_U11896 ( .A(u5_mult_82_n6871), .ZN(u5_mult_82_n6869) );
  INV_X32 u5_mult_82_U11895 ( .A(u5_mult_82_n6871), .ZN(u5_mult_82_n6868) );
  INV_X32 u5_mult_82_U11894 ( .A(u5_mult_82_n6871), .ZN(u5_mult_82_n6867) );
  INV_X32 u5_mult_82_U11893 ( .A(u5_mult_82_n6865), .ZN(u5_mult_82_n6864) );
  INV_X32 u5_mult_82_U11892 ( .A(u5_mult_82_n6865), .ZN(u5_mult_82_n6863) );
  INV_X32 u5_mult_82_U11891 ( .A(u5_mult_82_n6866), .ZN(u5_mult_82_n6862) );
  INV_X32 u5_mult_82_U11890 ( .A(u5_mult_82_n6866), .ZN(u5_mult_82_n6861) );
  INV_X32 u5_mult_82_U11889 ( .A(u5_mult_82_n7013), .ZN(u5_mult_82_n6860) );
  INV_X32 u5_mult_82_U11888 ( .A(u5_mult_82_n6860), .ZN(u5_mult_82_n6859) );
  INV_X32 u5_mult_82_U11887 ( .A(u5_mult_82_n6860), .ZN(u5_mult_82_n6858) );
  INV_X32 u5_mult_82_U11886 ( .A(u5_mult_82_n6860), .ZN(u5_mult_82_n6857) );
  INV_X32 u5_mult_82_U11885 ( .A(u5_mult_82_n6860), .ZN(u5_mult_82_n6856) );
  INV_X32 u5_mult_82_U11884 ( .A(u5_mult_82_n6855), .ZN(u5_mult_82_n6850) );
  INV_X32 u5_mult_82_U11883 ( .A(u5_mult_82_n6847), .ZN(u5_mult_82_n6845) );
  INV_X32 u5_mult_82_U11882 ( .A(u5_mult_82_n6847), .ZN(u5_mult_82_n6844) );
  INV_X32 u5_mult_82_U11881 ( .A(u5_mult_82_n6848), .ZN(u5_mult_82_n6843) );
  INV_X32 u5_mult_82_U11880 ( .A(u5_mult_82_n6848), .ZN(u5_mult_82_n6842) );
  INV_X32 u5_mult_82_U11879 ( .A(u5_mult_82_n6836), .ZN(u5_mult_82_n6841) );
  INV_X32 u5_mult_82_U11878 ( .A(u5_mult_82_n6841), .ZN(u5_mult_82_n6840) );
  INV_X32 u5_mult_82_U11877 ( .A(u5_mult_82_n6841), .ZN(u5_mult_82_n6839) );
  INV_X32 u5_mult_82_U11876 ( .A(u5_mult_82_n6841), .ZN(u5_mult_82_n6838) );
  INV_X32 u5_mult_82_U11875 ( .A(u5_mult_82_n6841), .ZN(u5_mult_82_n6837) );
  INV_X32 u5_mult_82_U11874 ( .A(u5_mult_82_net64893), .ZN(u5_mult_82_net64883) );
  INV_X32 u5_mult_82_U11873 ( .A(u5_mult_82_net64893), .ZN(u5_mult_82_net64881) );
  INV_X32 u5_mult_82_U11872 ( .A(u5_mult_82_net64911), .ZN(u5_mult_82_net64901) );
  INV_X32 u5_mult_82_U11871 ( .A(u5_mult_82_net64915), .ZN(u5_mult_82_net64913) );
  INV_X32 u5_mult_82_U11870 ( .A(u5_mult_82_net64949), .ZN(u5_mult_82_net64945) );
  INV_X32 u5_mult_82_U11869 ( .A(u5_mult_82_net64945), .ZN(u5_mult_82_net64941) );
  INV_X32 u5_mult_82_U11868 ( .A(u5_mult_82_net64945), .ZN(u5_mult_82_net64939) );
  INV_X32 u5_mult_82_U11867 ( .A(u5_mult_82_net64947), .ZN(u5_mult_82_net64937) );
  INV_X32 u5_mult_82_U11866 ( .A(u5_mult_82_net64947), .ZN(u5_mult_82_net64935) );
  INV_X32 u5_mult_82_U11865 ( .A(u5_mult_82_n6834), .ZN(u5_mult_82_n6833) );
  INV_X32 u5_mult_82_U11864 ( .A(u5_mult_82_n6825), .ZN(u5_mult_82_n6830) );
  INV_X32 u5_mult_82_U11863 ( .A(u5_mult_82_n6830), .ZN(u5_mult_82_n6829) );
  INV_X32 u5_mult_82_U11862 ( .A(u5_mult_82_n6830), .ZN(u5_mult_82_n6828) );
  INV_X32 u5_mult_82_U11861 ( .A(u5_mult_82_n6830), .ZN(u5_mult_82_n6827) );
  INV_X32 u5_mult_82_U11860 ( .A(u5_mult_82_n6830), .ZN(u5_mult_82_n6826) );
  INV_X32 u5_mult_82_U11859 ( .A(u5_mult_82_n2480), .ZN(u5_mult_82_n6823) );
  INV_X32 u5_mult_82_U11858 ( .A(u5_mult_82_n2480), .ZN(u5_mult_82_n6822) );
  INV_X32 u5_mult_82_U11857 ( .A(u5_mult_82_n2480), .ZN(u5_mult_82_n6821) );
  INV_X32 u5_mult_82_U11856 ( .A(u5_mult_82_n6815), .ZN(u5_mult_82_n6819) );
  INV_X32 u5_mult_82_U11855 ( .A(u5_mult_82_n6819), .ZN(u5_mult_82_n6818) );
  INV_X32 u5_mult_82_U11854 ( .A(u5_mult_82_n6819), .ZN(u5_mult_82_n6817) );
  INV_X32 u5_mult_82_U11853 ( .A(u5_mult_82_n6819), .ZN(u5_mult_82_n6816) );
  INV_X32 u5_mult_82_U11852 ( .A(u5_mult_82_n6809), .ZN(u5_mult_82_n6814) );
  INV_X32 u5_mult_82_U11851 ( .A(u5_mult_82_n6814), .ZN(u5_mult_82_n6812) );
  INV_X32 u5_mult_82_U11850 ( .A(u5_mult_82_n6808), .ZN(u5_mult_82_n6803) );
  INV_X32 u5_mult_82_U11849 ( .A(u5_mult_82_n6801), .ZN(u5_mult_82_n6799) );
  INV_X32 u5_mult_82_U11848 ( .A(u5_mult_82_n6801), .ZN(u5_mult_82_n6798) );
  INV_X32 u5_mult_82_U11847 ( .A(u5_mult_82_n6795), .ZN(u5_mult_82_n6793) );
  INV_X32 u5_mult_82_U11846 ( .A(u5_mult_82_n6795), .ZN(u5_mult_82_n6792) );
  INV_X32 u5_mult_82_U11845 ( .A(u5_mult_82_n6796), .ZN(u5_mult_82_n6791) );
  INV_X32 u5_mult_82_U11844 ( .A(u5_mult_82_n6787), .ZN(u5_mult_82_n6786) );
  INV_X32 u5_mult_82_U11843 ( .A(u5_mult_82_n6787), .ZN(u5_mult_82_n6785) );
  INV_X32 u5_mult_82_U11842 ( .A(u5_mult_82_n6788), .ZN(u5_mult_82_n6784) );
  INV_X32 u5_mult_82_U11841 ( .A(u5_mult_82_n7006), .ZN(u5_mult_82_n6782) );
  INV_X32 u5_mult_82_U11840 ( .A(u5_mult_82_n6782), .ZN(u5_mult_82_n6780) );
  INV_X32 u5_mult_82_U11839 ( .A(u5_mult_82_n6782), .ZN(u5_mult_82_n6779) );
  INV_X32 u5_mult_82_U11838 ( .A(u5_mult_82_n6782), .ZN(u5_mult_82_n6778) );
  INV_X32 u5_mult_82_U11837 ( .A(u5_mult_82_n6782), .ZN(u5_mult_82_n6777) );
  INV_X32 u5_mult_82_U11836 ( .A(u5_mult_82_n6771), .ZN(u5_mult_82_n6776) );
  INV_X32 u5_mult_82_U11835 ( .A(u5_mult_82_n6776), .ZN(u5_mult_82_n6775) );
  INV_X32 u5_mult_82_U11834 ( .A(u5_mult_82_n6776), .ZN(u5_mult_82_n6774) );
  INV_X32 u5_mult_82_U11833 ( .A(u5_mult_82_n6776), .ZN(u5_mult_82_n6773) );
  INV_X32 u5_mult_82_U11832 ( .A(u5_mult_82_n6776), .ZN(u5_mult_82_n6772) );
  INV_X32 u5_mult_82_U11831 ( .A(u5_mult_82_n6765), .ZN(u5_mult_82_n6770) );
  INV_X32 u5_mult_82_U11830 ( .A(u5_mult_82_n6770), .ZN(u5_mult_82_n6769) );
  INV_X32 u5_mult_82_U11829 ( .A(u5_mult_82_n6770), .ZN(u5_mult_82_n6768) );
  INV_X32 u5_mult_82_U11828 ( .A(u5_mult_82_n6770), .ZN(u5_mult_82_n6767) );
  INV_X32 u5_mult_82_U11827 ( .A(u5_mult_82_n6770), .ZN(u5_mult_82_n6766) );
  INV_X32 u5_mult_82_U11826 ( .A(u5_mult_82_n6758), .ZN(u5_mult_82_n6764) );
  INV_X32 u5_mult_82_U11825 ( .A(u5_mult_82_n6764), .ZN(u5_mult_82_n6759) );
  INV_X32 u5_mult_82_U11824 ( .A(u5_mult_82_n1272), .ZN(u5_mult_82_net65223)
         );
  INV_X32 u5_mult_82_U11823 ( .A(u5_mult_82_n6750), .ZN(u5_mult_82_n6757) );
  INV_X32 u5_mult_82_U11822 ( .A(u5_mult_82_n6750), .ZN(u5_mult_82_n6756) );
  INV_X32 u5_mult_82_U11821 ( .A(u5_mult_82_n6756), .ZN(u5_mult_82_n6755) );
  INV_X32 u5_mult_82_U11820 ( .A(u5_mult_82_n6756), .ZN(u5_mult_82_n6754) );
  INV_X32 u5_mult_82_U11819 ( .A(u5_mult_82_n6757), .ZN(u5_mult_82_n6753) );
  INV_X32 u5_mult_82_U11818 ( .A(u5_mult_82_n6757), .ZN(u5_mult_82_n6752) );
  INV_X32 u5_mult_82_U11817 ( .A(u5_mult_82_n6751), .ZN(u5_mult_82_n6750) );
  INV_X32 u5_mult_82_U11816 ( .A(u5_mult_82_n6745), .ZN(u5_mult_82_n6749) );
  INV_X32 u5_mult_82_U11815 ( .A(u5_mult_82_n6745), .ZN(u5_mult_82_n6748) );
  INV_X32 u5_mult_82_U11814 ( .A(u5_mult_82_n6745), .ZN(u5_mult_82_n6747) );
  INV_X32 u5_mult_82_U11813 ( .A(u5_mult_82_n6745), .ZN(u5_mult_82_n6746) );
  INV_X32 u5_mult_82_U11812 ( .A(u5_mult_82_net65287), .ZN(u5_mult_82_net65285) );
  INV_X32 u5_mult_82_U11811 ( .A(u5_mult_82_net65287), .ZN(u5_mult_82_net65279) );
  INV_X32 u5_mult_82_U11810 ( .A(u5_mult_82_net65293), .ZN(u5_mult_82_net65277) );
  INV_X32 u5_mult_82_U11809 ( .A(u5_mult_82_n6744), .ZN(u5_mult_82_n6741) );
  INV_X32 u5_mult_82_U11808 ( .A(u5_mult_82_n1290), .ZN(u5_mult_82_net65315)
         );
  INV_X32 u5_mult_82_U11807 ( .A(u5_mult_82_n6738), .ZN(u5_mult_82_n6736) );
  INV_X32 u5_mult_82_U11806 ( .A(u5_mult_82_n6738), .ZN(u5_mult_82_n6735) );
  INV_X32 u5_mult_82_U11805 ( .A(u5_mult_82_n6739), .ZN(u5_mult_82_n6734) );
  INV_X32 u5_mult_82_U11804 ( .A(u5_mult_82_net65361), .ZN(u5_mult_82_net65351) );
  INV_X32 u5_mult_82_U11803 ( .A(u5_mult_82_net65361), .ZN(u5_mult_82_net65349) );
  INV_X32 u5_mult_82_U11802 ( .A(u5_mult_82_net65379), .ZN(u5_mult_82_net65369) );
  INV_X32 u5_mult_82_U11801 ( .A(u5_mult_82_n1326), .ZN(u5_mult_82_net65387)
         );
  INV_X32 u5_mult_82_U11800 ( .A(u5_mult_82_n1328), .ZN(u5_mult_82_net65385)
         );
  INV_X32 u5_mult_82_U11799 ( .A(u5_mult_82_n1278), .ZN(u5_mult_82_net65405)
         );
  INV_X32 u5_mult_82_U11798 ( .A(u5_mult_82_n1280), .ZN(u5_mult_82_net65403)
         );
  INV_X32 u5_mult_82_U11797 ( .A(u5_mult_82_n6731), .ZN(u5_mult_82_n6728) );
  INV_X32 u5_mult_82_U11796 ( .A(u5_mult_82_net65451), .ZN(u5_mult_82_net65441) );
  INV_X32 u5_mult_82_U11795 ( .A(u5_mult_82_n6724), .ZN(u5_mult_82_n6722) );
  INV_X32 u5_mult_82_U11794 ( .A(u5_mult_82_n6724), .ZN(u5_mult_82_n6721) );
  INV_X32 u5_mult_82_U11793 ( .A(u5_mult_82_n6725), .ZN(u5_mult_82_n6720) );
  INV_X32 u5_mult_82_U11792 ( .A(u5_mult_82_n6718), .ZN(u5_mult_82_n6717) );
  INV_X32 u5_mult_82_U11791 ( .A(u5_mult_82_n6718), .ZN(u5_mult_82_n6716) );
  INV_X32 u5_mult_82_U11790 ( .A(u5_mult_82_n6718), .ZN(u5_mult_82_n6715) );
  INV_X32 u5_mult_82_U11789 ( .A(u5_mult_82_n6718), .ZN(u5_mult_82_n6714) );
  INV_X32 u5_mult_82_U11788 ( .A(u5_mult_82_n6712), .ZN(u5_mult_82_n6713) );
  INV_X32 u5_mult_82_U11787 ( .A(u5_mult_82_n6711), .ZN(u5_mult_82_n6710) );
  INV_X32 u5_mult_82_U11786 ( .A(u5_mult_82_n6711), .ZN(u5_mult_82_n6709) );
  INV_X32 u5_mult_82_U11785 ( .A(u5_mult_82_n6711), .ZN(u5_mult_82_n6708) );
  INV_X32 u5_mult_82_U11784 ( .A(u5_mult_82_n6711), .ZN(u5_mult_82_n6707) );
  INV_X32 u5_mult_82_U11783 ( .A(u5_mult_82_n6705), .ZN(u5_mult_82_n6706) );
  INV_X32 u5_mult_82_U11782 ( .A(u5_mult_82_net65523), .ZN(u5_mult_82_net65513) );
  INV_X32 u5_mult_82_U11781 ( .A(u5_mult_82_n6703), .ZN(u5_mult_82_n6700) );
  INV_X32 u5_mult_82_U11780 ( .A(u5_mult_82_n6697), .ZN(u5_mult_82_n6696) );
  INV_X32 u5_mult_82_U11779 ( .A(u5_mult_82_n6697), .ZN(u5_mult_82_n6695) );
  INV_X32 u5_mult_82_U11778 ( .A(u5_mult_82_n6697), .ZN(u5_mult_82_n6694) );
  INV_X32 u5_mult_82_U11777 ( .A(u5_mult_82_n6697), .ZN(u5_mult_82_n6693) );
  INV_X32 u5_mult_82_U11776 ( .A(u5_mult_82_n6691), .ZN(u5_mult_82_n6692) );
  INV_X32 u5_mult_82_U11775 ( .A(u5_mult_82_n6688), .ZN(u5_mult_82_n6686) );
  INV_X32 u5_mult_82_U11774 ( .A(u5_mult_82_n6688), .ZN(u5_mult_82_n6685) );
  INV_X32 u5_mult_82_U11773 ( .A(u5_mult_82_n6689), .ZN(u5_mult_82_n6684) );
  INV_X32 u5_mult_82_U11772 ( .A(u5_mult_82_n6682), .ZN(u5_mult_82_n6681) );
  INV_X32 u5_mult_82_U11771 ( .A(u5_mult_82_n6682), .ZN(u5_mult_82_n6680) );
  INV_X32 u5_mult_82_U11770 ( .A(u5_mult_82_n6682), .ZN(u5_mult_82_n6679) );
  INV_X32 u5_mult_82_U11769 ( .A(u5_mult_82_n6682), .ZN(u5_mult_82_n6678) );
  INV_X32 u5_mult_82_U11768 ( .A(u5_mult_82_n6676), .ZN(u5_mult_82_n6677) );
  INV_X32 u5_mult_82_U11767 ( .A(u5_mult_82_n6675), .ZN(u5_mult_82_n6674) );
  INV_X32 u5_mult_82_U11766 ( .A(u5_mult_82_n6675), .ZN(u5_mult_82_n6673) );
  INV_X32 u5_mult_82_U11765 ( .A(u5_mult_82_n6675), .ZN(u5_mult_82_n6672) );
  INV_X32 u5_mult_82_U11764 ( .A(u5_mult_82_n6675), .ZN(u5_mult_82_n6671) );
  INV_X32 u5_mult_82_U11763 ( .A(u5_mult_82_n6669), .ZN(u5_mult_82_n6670) );
  INV_X32 u5_mult_82_U11762 ( .A(u5_mult_82_n6667), .ZN(u5_mult_82_n6665) );
  INV_X32 u5_mult_82_U11761 ( .A(u5_mult_82_n6667), .ZN(u5_mult_82_n6664) );
  INV_X32 u5_mult_82_U11760 ( .A(u5_mult_82_n6654), .ZN(u5_mult_82_n6661) );
  INV_X32 u5_mult_82_U11759 ( .A(u5_mult_82_n6660), .ZN(u5_mult_82_n6659) );
  INV_X32 u5_mult_82_U11758 ( .A(u5_mult_82_n6660), .ZN(u5_mult_82_n6658) );
  INV_X32 u5_mult_82_U11757 ( .A(u5_mult_82_n6661), .ZN(u5_mult_82_n6656) );
  INV_X32 u5_mult_82_U11756 ( .A(u5_mult_82_n6661), .ZN(u5_mult_82_n6655) );
  INV_X32 u5_mult_82_U11755 ( .A(u5_mult_82_n6653), .ZN(u5_mult_82_n6651) );
  INV_X32 u5_mult_82_U11754 ( .A(u5_mult_82_n6653), .ZN(u5_mult_82_n6650) );
  INV_X32 u5_mult_82_U11753 ( .A(u5_mult_82_n6653), .ZN(u5_mult_82_n6649) );
  INV_X32 u5_mult_82_U11752 ( .A(u5_mult_82_net65685), .ZN(u5_mult_82_net65675) );
  INV_X32 u5_mult_82_U11751 ( .A(u5_mult_82_n6646), .ZN(u5_mult_82_n6645) );
  INV_X32 u5_mult_82_U11750 ( .A(u5_mult_82_n6647), .ZN(u5_mult_82_n6642) );
  INV_X32 u5_mult_82_U11749 ( .A(u5_mult_82_n6639), .ZN(u5_mult_82_n6637) );
  INV_X32 u5_mult_82_U11748 ( .A(u5_mult_82_n6639), .ZN(u5_mult_82_n6636) );
  INV_X32 u5_mult_82_U11747 ( .A(u5_mult_82_n6640), .ZN(u5_mult_82_n6635) );
  INV_X32 u5_mult_82_U11746 ( .A(u5_mult_82_n6632), .ZN(u5_mult_82_n6630) );
  INV_X32 u5_mult_82_U11745 ( .A(u5_mult_82_n6625), .ZN(u5_mult_82_n6623) );
  INV_X32 u5_mult_82_U11744 ( .A(u5_mult_82_n6625), .ZN(u5_mult_82_n6622) );
  INV_X32 u5_mult_82_U11743 ( .A(u5_mult_82_n6618), .ZN(u5_mult_82_n6617) );
  INV_X32 u5_mult_82_U11742 ( .A(u5_mult_82_n6618), .ZN(u5_mult_82_n6615) );
  INV_X32 u5_mult_82_U11741 ( .A(u5_mult_82_n6612), .ZN(u5_mult_82_n6611) );
  INV_X32 u5_mult_82_U11740 ( .A(u5_mult_82_n6612), .ZN(u5_mult_82_n6610) );
  INV_X32 u5_mult_82_U11739 ( .A(u5_mult_82_n6612), .ZN(u5_mult_82_n6609) );
  INV_X32 u5_mult_82_U11738 ( .A(u5_mult_82_n6612), .ZN(u5_mult_82_n6608) );
  INV_X32 u5_mult_82_U11737 ( .A(u5_mult_82_n6606), .ZN(u5_mult_82_n6607) );
  INV_X32 u5_mult_82_U11736 ( .A(u5_mult_82_n6605), .ZN(u5_mult_82_n6603) );
  INV_X32 u5_mult_82_U11735 ( .A(u5_mult_82_n6605), .ZN(u5_mult_82_n6602) );
  INV_X32 u5_mult_82_U11734 ( .A(u5_mult_82_n6605), .ZN(u5_mult_82_n6601) );
  INV_X32 u5_mult_82_U11733 ( .A(u5_mult_82_n6599), .ZN(u5_mult_82_n6600) );
  INV_X32 u5_mult_82_U11732 ( .A(u5_mult_82_n6598), .ZN(u5_mult_82_n6597) );
  INV_X32 u5_mult_82_U11731 ( .A(u5_mult_82_n6598), .ZN(u5_mult_82_n6596) );
  INV_X32 u5_mult_82_U11730 ( .A(u5_mult_82_n6598), .ZN(u5_mult_82_n6595) );
  INV_X32 u5_mult_82_U11729 ( .A(u5_mult_82_n6598), .ZN(u5_mult_82_n6594) );
  INV_X32 u5_mult_82_U11728 ( .A(u5_mult_82_n6592), .ZN(u5_mult_82_n6593) );
  INV_X32 u5_mult_82_U11727 ( .A(u5_mult_82_n6584), .ZN(u5_mult_82_n6590) );
  INV_X32 u5_mult_82_U11726 ( .A(u5_mult_82_n6590), .ZN(u5_mult_82_n6589) );
  INV_X32 u5_mult_82_U11725 ( .A(u5_mult_82_n6590), .ZN(u5_mult_82_n6588) );
  INV_X32 u5_mult_82_U11724 ( .A(u5_mult_82_n6590), .ZN(u5_mult_82_n6587) );
  INV_X32 u5_mult_82_U11723 ( .A(u5_mult_82_n6591), .ZN(u5_mult_82_n6586) );
  INV_X32 u5_mult_82_U11722 ( .A(u5_mult_82_n6591), .ZN(u5_mult_82_n6585) );
  INV_X32 u5_mult_82_U11721 ( .A(u5_mult_82_n6582), .ZN(u5_mult_82_n6581) );
  INV_X32 u5_mult_82_U11720 ( .A(u5_mult_82_n6583), .ZN(u5_mult_82_n6578) );
  INV_X32 u5_mult_82_U11719 ( .A(u5_mult_82_n6575), .ZN(u5_mult_82_n6574) );
  INV_X32 u5_mult_82_U11718 ( .A(u5_mult_82_n6569), .ZN(u5_mult_82_n6567) );
  INV_X32 u5_mult_82_U11717 ( .A(u5_mult_82_n6569), .ZN(u5_mult_82_n6566) );
  INV_X32 u5_mult_82_U11716 ( .A(u5_mult_82_n6569), .ZN(u5_mult_82_n6565) );
  INV_X32 u5_mult_82_U11715 ( .A(u5_mult_82_n6563), .ZN(u5_mult_82_n6564) );
  INV_X32 u5_mult_82_U11714 ( .A(u5_mult_82_n6561), .ZN(u5_mult_82_n6559) );
  INV_X32 u5_mult_82_U11713 ( .A(u5_mult_82_n6554), .ZN(u5_mult_82_n6552) );
  INV_X32 u5_mult_82_U11712 ( .A(u5_mult_82_n6554), .ZN(u5_mult_82_n6551) );
  INV_X32 u5_mult_82_U11711 ( .A(u5_mult_82_n6541), .ZN(u5_mult_82_n6548) );
  INV_X32 u5_mult_82_U11710 ( .A(u5_mult_82_n6548), .ZN(u5_mult_82_n6547) );
  INV_X32 u5_mult_82_U11709 ( .A(u5_mult_82_n6548), .ZN(u5_mult_82_n6546) );
  INV_X32 u5_mult_82_U11708 ( .A(u5_mult_82_n6548), .ZN(u5_mult_82_n6545) );
  INV_X32 u5_mult_82_U11707 ( .A(u5_mult_82_n6548), .ZN(u5_mult_82_n6544) );
  INV_X32 u5_mult_82_U11706 ( .A(u5_mult_82_n6542), .ZN(u5_mult_82_n6543) );
  INV_X32 u5_mult_82_U11705 ( .A(u5_mult_82_n6534), .ZN(u5_mult_82_n6539) );
  INV_X32 u5_mult_82_U11704 ( .A(u5_mult_82_n6539), .ZN(u5_mult_82_n6537) );
  INV_X32 u5_mult_82_U11703 ( .A(u5_mult_82_n6539), .ZN(u5_mult_82_n6536) );
  INV_X32 u5_mult_82_U11702 ( .A(u5_mult_82_n6532), .ZN(u5_mult_82_n6530) );
  INV_X32 u5_mult_82_U11701 ( .A(u5_mult_82_n6532), .ZN(u5_mult_82_n6529) );
  INV_X32 u5_mult_82_U11700 ( .A(u5_mult_82_n6533), .ZN(u5_mult_82_n6528) );
  INV_X32 u5_mult_82_U11699 ( .A(u5_mult_82_net66025), .ZN(u5_mult_82_net66019) );
  INV_X32 u5_mult_82_U11698 ( .A(u5_mult_82_net66043), .ZN(u5_mult_82_net66041) );
  INV_X32 u5_mult_82_U11697 ( .A(u5_mult_82_net66043), .ZN(u5_mult_82_net66039) );
  INV_X32 u5_mult_82_U11696 ( .A(u5_mult_82_net66043), .ZN(u5_mult_82_net66037) );
  INV_X32 u5_mult_82_U11695 ( .A(u5_mult_82_n6518), .ZN(u5_mult_82_n6526) );
  INV_X32 u5_mult_82_U11694 ( .A(u5_mult_82_n6518), .ZN(u5_mult_82_n6525) );
  INV_X32 u5_mult_82_U11693 ( .A(u5_mult_82_n6525), .ZN(u5_mult_82_n6524) );
  INV_X32 u5_mult_82_U11692 ( .A(u5_mult_82_n6525), .ZN(u5_mult_82_n6523) );
  INV_X32 u5_mult_82_U11691 ( .A(u5_mult_82_n6525), .ZN(u5_mult_82_n6522) );
  INV_X32 u5_mult_82_U11690 ( .A(u5_mult_82_n6526), .ZN(u5_mult_82_n6521) );
  INV_X32 u5_mult_82_U11689 ( .A(u5_mult_82_n6526), .ZN(u5_mult_82_n6520) );
  INV_X32 u5_mult_82_U11688 ( .A(u5_mult_82_n6519), .ZN(u5_mult_82_n6518) );
  INV_X32 u5_mult_82_U11687 ( .A(u5_mult_82_n6517), .ZN(u5_mult_82_n6516) );
  INV_X32 u5_mult_82_U11686 ( .A(u5_mult_82_n6517), .ZN(u5_mult_82_n6515) );
  INV_X32 u5_mult_82_U11685 ( .A(u5_mult_82_n6517), .ZN(u5_mult_82_n6514) );
  INV_X32 u5_mult_82_U11684 ( .A(u5_mult_82_n6517), .ZN(u5_mult_82_n6513) );
  INV_X32 u5_mult_82_U11683 ( .A(u5_mult_82_net66097), .ZN(u5_mult_82_net66093) );
  INV_X32 u5_mult_82_U11682 ( .A(u5_mult_82_net66097), .ZN(u5_mult_82_net66091) );
  INV_X32 u5_mult_82_U11681 ( .A(u5_mult_82_net66121), .ZN(u5_mult_82_net66111) );
  INV_X32 u5_mult_82_U11680 ( .A(u5_mult_82_net66121), .ZN(u5_mult_82_net66109) );
  INV_X8 u5_mult_82_U11679 ( .A(u5_mult_82_n6984), .ZN(u5_mult_82_n6982) );
  INV_X8 u5_mult_82_U11678 ( .A(u5_mult_82_n6984), .ZN(u5_mult_82_n6983) );
  INV_X8 u5_mult_82_U11677 ( .A(n4793), .ZN(u5_mult_82_n7006) );
  INV_X4 u5_mult_82_U11676 ( .A(u5_mult_82_n6511), .ZN(u5_mult_82_SUMB_1__50_)
         );
  XNOR2_X2 u5_mult_82_U11675 ( .A(u5_mult_82_ab_1__50_), .B(
        u5_mult_82_ab_0__51_), .ZN(u5_mult_82_n6511) );
  XNOR2_X2 u5_mult_82_U11674 ( .A(u5_mult_82_ab_1__49_), .B(
        u5_mult_82_ab_0__50_), .ZN(u5_mult_82_n6509) );
  INV_X4 u5_mult_82_U11673 ( .A(u5_mult_82_n6508), .ZN(
        u5_mult_82_CARRYB_1__49_) );
  INV_X4 u5_mult_82_U11672 ( .A(u5_mult_82_n6507), .ZN(u5_mult_82_SUMB_1__48_)
         );
  XNOR2_X2 u5_mult_82_U11671 ( .A(u5_mult_82_ab_1__48_), .B(
        u5_mult_82_ab_0__49_), .ZN(u5_mult_82_n6507) );
  INV_X4 u5_mult_82_U11670 ( .A(u5_mult_82_n6506), .ZN(
        u5_mult_82_CARRYB_1__48_) );
  XNOR2_X2 u5_mult_82_U11669 ( .A(u5_mult_82_ab_1__47_), .B(
        u5_mult_82_ab_0__48_), .ZN(u5_mult_82_n6505) );
  INV_X4 u5_mult_82_U11668 ( .A(u5_mult_82_n6501), .ZN(u5_mult_82_SUMB_1__45_)
         );
  XNOR2_X2 u5_mult_82_U11667 ( .A(u5_mult_82_n68), .B(u5_mult_82_n64), .ZN(
        u5_mult_82_n6501) );
  INV_X4 u5_mult_82_U11666 ( .A(u5_mult_82_n6499), .ZN(u5_mult_82_SUMB_1__44_)
         );
  XNOR2_X2 u5_mult_82_U11665 ( .A(u5_mult_82_ab_1__44_), .B(
        u5_mult_82_ab_0__45_), .ZN(u5_mult_82_n6499) );
  INV_X4 u5_mult_82_U11664 ( .A(u5_mult_82_n6498), .ZN(
        u5_mult_82_CARRYB_1__44_) );
  INV_X4 u5_mult_82_U11663 ( .A(u5_mult_82_n6497), .ZN(
        u5_mult_82_CARRYB_1__43_) );
  INV_X4 u5_mult_82_U11662 ( .A(u5_mult_82_n6496), .ZN(u5_mult_82_SUMB_1__42_)
         );
  XNOR2_X2 u5_mult_82_U11661 ( .A(u5_mult_82_ab_1__42_), .B(
        u5_mult_82_ab_0__43_), .ZN(u5_mult_82_n6496) );
  INV_X4 u5_mult_82_U11660 ( .A(u5_mult_82_n6495), .ZN(
        u5_mult_82_CARRYB_1__42_) );
  NAND2_X2 u5_mult_82_U11659 ( .A1(u5_mult_82_ab_0__43_), .A2(
        u5_mult_82_ab_1__42_), .ZN(u5_mult_82_n6495) );
  INV_X4 u5_mult_82_U11658 ( .A(u5_mult_82_n6494), .ZN(
        u5_mult_82_CARRYB_1__41_) );
  INV_X4 u5_mult_82_U11657 ( .A(u5_mult_82_n6493), .ZN(u5_mult_82_SUMB_1__40_)
         );
  XNOR2_X2 u5_mult_82_U11656 ( .A(u5_mult_82_n3280), .B(u5_mult_82_ab_0__41_), 
        .ZN(u5_mult_82_n6493) );
  INV_X4 u5_mult_82_U11655 ( .A(u5_mult_82_n6492), .ZN(u5_mult_82_SUMB_1__38_)
         );
  XNOR2_X2 u5_mult_82_U11654 ( .A(u5_mult_82_ab_1__38_), .B(
        u5_mult_82_ab_0__39_), .ZN(u5_mult_82_n6492) );
  INV_X4 u5_mult_82_U11653 ( .A(u5_mult_82__UDW__88983_net69746), .ZN(
        u5_mult_82_CARRYB_1__37_) );
  INV_X4 u5_mult_82_U11652 ( .A(u5_mult_82_n6491), .ZN(u5_mult_82_SUMB_1__36_)
         );
  INV_X4 u5_mult_82_U11651 ( .A(u5_mult_82_n6490), .ZN(u5_mult_82_SUMB_1__35_)
         );
  XNOR2_X2 u5_mult_82_U11650 ( .A(u5_mult_82_n2748), .B(u5_mult_82_ab_0__36_), 
        .ZN(u5_mult_82_n6490) );
  INV_X4 u5_mult_82_U11649 ( .A(u5_mult_82_n6489), .ZN(
        u5_mult_82_CARRYB_1__34_) );
  INV_X4 u5_mult_82_U11648 ( .A(u5_mult_82_n6488), .ZN(u5_mult_82_SUMB_1__33_)
         );
  XNOR2_X2 u5_mult_82_U11647 ( .A(u5_mult_82_ab_1__33_), .B(
        u5_mult_82_ab_0__34_), .ZN(u5_mult_82_n6488) );
  INV_X4 u5_mult_82_U11646 ( .A(u5_mult_82_n6487), .ZN(
        u5_mult_82_CARRYB_1__32_) );
  NAND2_X2 u5_mult_82_U11645 ( .A1(u5_mult_82_ab_0__33_), .A2(
        u5_mult_82_ab_1__32_), .ZN(u5_mult_82_n6487) );
  INV_X4 u5_mult_82_U11644 ( .A(u5_mult_82_n6486), .ZN(u5_mult_82_SUMB_1__31_)
         );
  XNOR2_X2 u5_mult_82_U11643 ( .A(u5_mult_82_ab_1__31_), .B(
        u5_mult_82_ab_0__32_), .ZN(u5_mult_82_n6486) );
  INV_X4 u5_mult_82_U11642 ( .A(u5_mult_82_n6485), .ZN(u5_mult_82_SUMB_1__30_)
         );
  INV_X4 u5_mult_82_U11641 ( .A(u5_mult_82_n6484), .ZN(
        u5_mult_82_CARRYB_1__30_) );
  INV_X4 u5_mult_82_U11640 ( .A(u5_mult_82_n6483), .ZN(u5_mult_82_SUMB_1__29_)
         );
  XNOR2_X2 u5_mult_82_U11639 ( .A(u5_mult_82_ab_1__29_), .B(
        u5_mult_82_ab_0__30_), .ZN(u5_mult_82_n6483) );
  INV_X4 u5_mult_82_U11638 ( .A(u5_mult_82_n6482), .ZN(
        u5_mult_82_CARRYB_1__29_) );
  INV_X4 u5_mult_82_U11637 ( .A(u5_mult_82_n6481), .ZN(u5_mult_82_SUMB_1__27_)
         );
  XNOR2_X2 u5_mult_82_U11636 ( .A(u5_mult_82_ab_1__27_), .B(
        u5_mult_82_ab_0__28_), .ZN(u5_mult_82_n6481) );
  INV_X4 u5_mult_82_U11635 ( .A(u5_mult_82_n6480), .ZN(
        u5_mult_82_CARRYB_1__27_) );
  INV_X4 u5_mult_82_U11634 ( .A(u5_mult_82_n6479), .ZN(u5_mult_82_SUMB_1__26_)
         );
  XNOR2_X2 u5_mult_82_U11633 ( .A(u5_mult_82_ab_1__26_), .B(
        u5_mult_82_ab_0__27_), .ZN(u5_mult_82_n6479) );
  NAND2_X2 u5_mult_82_U11632 ( .A1(u5_mult_82_ab_0__27_), .A2(
        u5_mult_82_ab_1__26_), .ZN(u5_mult_82_n6478) );
  INV_X4 u5_mult_82_U11631 ( .A(u5_mult_82_n6477), .ZN(u5_mult_82_SUMB_1__25_)
         );
  XNOR2_X2 u5_mult_82_U11630 ( .A(u5_mult_82_ab_1__25_), .B(
        u5_mult_82_ab_0__26_), .ZN(u5_mult_82_n6477) );
  INV_X4 u5_mult_82_U11629 ( .A(u5_mult_82_n6476), .ZN(
        u5_mult_82_CARRYB_1__25_) );
  NAND2_X2 u5_mult_82_U11628 ( .A1(u5_mult_82_ab_0__26_), .A2(
        u5_mult_82_ab_1__25_), .ZN(u5_mult_82_n6476) );
  INV_X4 u5_mult_82_U11627 ( .A(u5_mult_82_n6475), .ZN(u5_mult_82_SUMB_1__24_)
         );
  XNOR2_X2 u5_mult_82_U11626 ( .A(u5_mult_82_ab_1__24_), .B(
        u5_mult_82_ab_0__25_), .ZN(u5_mult_82_n6475) );
  INV_X4 u5_mult_82_U11625 ( .A(u5_mult_82_n6474), .ZN(
        u5_mult_82_CARRYB_1__24_) );
  NAND2_X2 u5_mult_82_U11624 ( .A1(u5_mult_82_ab_0__25_), .A2(
        u5_mult_82_ab_1__24_), .ZN(u5_mult_82_n6474) );
  INV_X4 u5_mult_82_U11623 ( .A(u5_mult_82_n6473), .ZN(u5_mult_82_SUMB_1__23_)
         );
  XNOR2_X2 u5_mult_82_U11622 ( .A(u5_mult_82_ab_1__23_), .B(
        u5_mult_82_ab_0__24_), .ZN(u5_mult_82_n6473) );
  INV_X4 u5_mult_82_U11621 ( .A(u5_mult_82_n6472), .ZN(
        u5_mult_82_CARRYB_1__23_) );
  NAND2_X2 u5_mult_82_U11620 ( .A1(u5_mult_82_ab_0__24_), .A2(
        u5_mult_82_ab_1__23_), .ZN(u5_mult_82_n6472) );
  INV_X4 u5_mult_82_U11619 ( .A(u5_mult_82_n6471), .ZN(u5_mult_82_SUMB_1__22_)
         );
  XNOR2_X2 u5_mult_82_U11618 ( .A(u5_mult_82_ab_1__22_), .B(
        u5_mult_82_ab_0__23_), .ZN(u5_mult_82_n6471) );
  INV_X4 u5_mult_82_U11617 ( .A(u5_mult_82_n6470), .ZN(
        u5_mult_82_CARRYB_1__21_) );
  NAND2_X2 u5_mult_82_U11616 ( .A1(u5_mult_82_ab_0__22_), .A2(
        u5_mult_82_ab_1__21_), .ZN(u5_mult_82_n6470) );
  INV_X4 u5_mult_82_U11615 ( .A(u5_mult_82_n6469), .ZN(u5_mult_82_SUMB_1__20_)
         );
  XNOR2_X2 u5_mult_82_U11614 ( .A(u5_mult_82_ab_1__20_), .B(
        u5_mult_82_ab_0__21_), .ZN(u5_mult_82_n6469) );
  INV_X4 u5_mult_82_U11613 ( .A(u5_mult_82_n6468), .ZN(u5_mult_82_SUMB_1__19_)
         );
  XNOR2_X2 u5_mult_82_U11612 ( .A(u5_mult_82_ab_1__19_), .B(
        u5_mult_82_ab_0__20_), .ZN(u5_mult_82_n6468) );
  INV_X4 u5_mult_82_U11611 ( .A(u5_mult_82_n6467), .ZN(
        u5_mult_82_CARRYB_1__19_) );
  NAND2_X2 u5_mult_82_U11610 ( .A1(u5_mult_82_ab_0__20_), .A2(
        u5_mult_82_ab_1__19_), .ZN(u5_mult_82_n6467) );
  INV_X4 u5_mult_82_U11609 ( .A(u5_mult_82_n6466), .ZN(
        u5_mult_82_CARRYB_1__18_) );
  NAND2_X2 u5_mult_82_U11608 ( .A1(u5_mult_82_ab_0__19_), .A2(
        u5_mult_82_ab_1__18_), .ZN(u5_mult_82_n6466) );
  INV_X4 u5_mult_82_U11607 ( .A(u5_mult_82_n6465), .ZN(u5_mult_82_SUMB_1__17_)
         );
  XNOR2_X2 u5_mult_82_U11606 ( .A(u5_mult_82_ab_1__17_), .B(
        u5_mult_82_ab_0__18_), .ZN(u5_mult_82_n6465) );
  INV_X4 u5_mult_82_U11605 ( .A(u5_mult_82_n6464), .ZN(u5_mult_82_SUMB_1__16_)
         );
  XNOR2_X2 u5_mult_82_U11604 ( .A(u5_mult_82_ab_1__16_), .B(
        u5_mult_82_ab_0__17_), .ZN(u5_mult_82_n6464) );
  INV_X4 u5_mult_82_U11603 ( .A(u5_mult_82_n6463), .ZN(
        u5_mult_82_CARRYB_1__16_) );
  NAND2_X2 u5_mult_82_U11602 ( .A1(u5_mult_82_ab_0__17_), .A2(
        u5_mult_82_ab_1__16_), .ZN(u5_mult_82_n6463) );
  INV_X4 u5_mult_82_U11601 ( .A(u5_mult_82_n6462), .ZN(u5_mult_82_SUMB_1__15_)
         );
  XNOR2_X2 u5_mult_82_U11600 ( .A(u5_mult_82_ab_1__15_), .B(
        u5_mult_82_ab_0__16_), .ZN(u5_mult_82_n6462) );
  INV_X4 u5_mult_82_U11599 ( .A(u5_mult_82_n6461), .ZN(u5_mult_82_SUMB_1__14_)
         );
  XNOR2_X2 u5_mult_82_U11598 ( .A(u5_mult_82_ab_1__14_), .B(
        u5_mult_82_ab_0__15_), .ZN(u5_mult_82_n6461) );
  INV_X4 u5_mult_82_U11597 ( .A(u5_mult_82_n6460), .ZN(
        u5_mult_82_CARRYB_1__14_) );
  NAND2_X2 u5_mult_82_U11596 ( .A1(u5_mult_82_ab_0__15_), .A2(
        u5_mult_82_ab_1__14_), .ZN(u5_mult_82_n6460) );
  INV_X4 u5_mult_82_U11595 ( .A(u5_mult_82_n6459), .ZN(u5_mult_82_SUMB_1__13_)
         );
  XNOR2_X2 u5_mult_82_U11594 ( .A(u5_mult_82_ab_1__13_), .B(
        u5_mult_82_ab_0__14_), .ZN(u5_mult_82_n6459) );
  INV_X4 u5_mult_82_U11593 ( .A(u5_mult_82_n6458), .ZN(
        u5_mult_82_CARRYB_1__13_) );
  NAND2_X2 u5_mult_82_U11592 ( .A1(u5_mult_82_ab_0__14_), .A2(
        u5_mult_82_ab_1__13_), .ZN(u5_mult_82_n6458) );
  INV_X4 u5_mult_82_U11591 ( .A(u5_mult_82_n6457), .ZN(u5_mult_82_SUMB_1__12_)
         );
  XNOR2_X2 u5_mult_82_U11590 ( .A(u5_mult_82_ab_1__12_), .B(
        u5_mult_82_ab_0__13_), .ZN(u5_mult_82_n6457) );
  INV_X4 u5_mult_82_U11589 ( .A(u5_mult_82_n6456), .ZN(
        u5_mult_82_CARRYB_1__12_) );
  NAND2_X2 u5_mult_82_U11588 ( .A1(u5_mult_82_ab_0__13_), .A2(
        u5_mult_82_ab_1__12_), .ZN(u5_mult_82_n6456) );
  INV_X4 u5_mult_82_U11587 ( .A(u5_mult_82_n6455), .ZN(u5_mult_82_SUMB_1__11_)
         );
  XNOR2_X2 u5_mult_82_U11586 ( .A(u5_mult_82_ab_1__11_), .B(
        u5_mult_82_ab_0__12_), .ZN(u5_mult_82_n6455) );
  INV_X4 u5_mult_82_U11585 ( .A(u5_mult_82_n6454), .ZN(
        u5_mult_82_CARRYB_1__11_) );
  NAND2_X2 u5_mult_82_U11584 ( .A1(u5_mult_82_ab_0__12_), .A2(
        u5_mult_82_ab_1__11_), .ZN(u5_mult_82_n6454) );
  INV_X4 u5_mult_82_U11583 ( .A(u5_mult_82_n6453), .ZN(u5_mult_82_SUMB_1__9_)
         );
  XNOR2_X2 u5_mult_82_U11582 ( .A(u5_mult_82_ab_1__9_), .B(
        u5_mult_82_ab_0__10_), .ZN(u5_mult_82_n6453) );
  INV_X4 u5_mult_82_U11581 ( .A(u5_mult_82_n6452), .ZN(u5_mult_82_CARRYB_1__9_) );
  NAND2_X2 u5_mult_82_U11580 ( .A1(u5_mult_82_ab_0__10_), .A2(
        u5_mult_82_ab_1__9_), .ZN(u5_mult_82_n6452) );
  INV_X4 u5_mult_82_U11579 ( .A(u5_mult_82_n6451), .ZN(u5_mult_82_SUMB_1__8_)
         );
  XNOR2_X2 u5_mult_82_U11578 ( .A(u5_mult_82_ab_1__8_), .B(u5_mult_82_ab_0__9_), .ZN(u5_mult_82_n6451) );
  INV_X4 u5_mult_82_U11577 ( .A(u5_mult_82_n6450), .ZN(u5_mult_82_SUMB_1__7_)
         );
  XNOR2_X2 u5_mult_82_U11576 ( .A(u5_mult_82_ab_1__7_), .B(u5_mult_82_ab_0__8_), .ZN(u5_mult_82_n6450) );
  INV_X4 u5_mult_82_U11575 ( .A(u5_mult_82_n6449), .ZN(u5_mult_82_CARRYB_1__7_) );
  NAND2_X2 u5_mult_82_U11574 ( .A1(u5_mult_82_ab_0__8_), .A2(
        u5_mult_82_ab_1__7_), .ZN(u5_mult_82_n6449) );
  INV_X4 u5_mult_82_U11573 ( .A(u5_mult_82_n6448), .ZN(u5_mult_82_SUMB_1__6_)
         );
  XNOR2_X2 u5_mult_82_U11572 ( .A(u5_mult_82_ab_1__6_), .B(u5_mult_82_ab_0__7_), .ZN(u5_mult_82_n6448) );
  INV_X4 u5_mult_82_U11571 ( .A(u5_mult_82_n6447), .ZN(u5_mult_82_CARRYB_1__6_) );
  NAND2_X2 u5_mult_82_U11570 ( .A1(u5_mult_82_ab_0__7_), .A2(
        u5_mult_82_ab_1__6_), .ZN(u5_mult_82_n6447) );
  INV_X4 u5_mult_82_U11569 ( .A(u5_mult_82_n6446), .ZN(u5_mult_82_SUMB_1__5_)
         );
  XNOR2_X2 u5_mult_82_U11568 ( .A(u5_mult_82_ab_1__5_), .B(u5_mult_82_ab_0__6_), .ZN(u5_mult_82_n6446) );
  INV_X4 u5_mult_82_U11567 ( .A(u5_mult_82_n6445), .ZN(u5_mult_82_CARRYB_1__5_) );
  NAND2_X2 u5_mult_82_U11566 ( .A1(u5_mult_82_ab_0__6_), .A2(
        u5_mult_82_ab_1__5_), .ZN(u5_mult_82_n6445) );
  INV_X4 u5_mult_82_U11565 ( .A(u5_mult_82_n6444), .ZN(u5_mult_82_SUMB_1__3_)
         );
  XNOR2_X2 u5_mult_82_U11564 ( .A(u5_mult_82_ab_1__3_), .B(u5_mult_82_ab_0__4_), .ZN(u5_mult_82_n6444) );
  INV_X4 u5_mult_82_U11563 ( .A(u5_mult_82_n6443), .ZN(u5_mult_82_CARRYB_1__3_) );
  NAND2_X2 u5_mult_82_U11562 ( .A1(u5_mult_82_ab_0__4_), .A2(
        u5_mult_82_ab_1__3_), .ZN(u5_mult_82_n6443) );
  INV_X4 u5_mult_82_U11561 ( .A(u5_mult_82_n6442), .ZN(u5_mult_82_SUMB_1__2_)
         );
  XNOR2_X2 u5_mult_82_U11560 ( .A(u5_mult_82_ab_1__2_), .B(u5_mult_82_ab_0__3_), .ZN(u5_mult_82_n6442) );
  INV_X4 u5_mult_82_U11559 ( .A(u5_mult_82_n6441), .ZN(u5_mult_82_CARRYB_1__2_) );
  NAND2_X2 u5_mult_82_U11558 ( .A1(u5_mult_82_ab_0__3_), .A2(
        u5_mult_82_ab_1__2_), .ZN(u5_mult_82_n6441) );
  INV_X4 u5_mult_82_U11557 ( .A(u5_mult_82_n6440), .ZN(u5_mult_82_CARRYB_1__0_) );
  NAND2_X2 u5_mult_82_U11556 ( .A1(u5_mult_82_ab_0__1_), .A2(
        u5_mult_82_ab_1__0_), .ZN(u5_mult_82_n6440) );
  INV_X4 u5_mult_82_U11555 ( .A(u5_mult_82_n6439), .ZN(
        u5_mult_82_CLA_CARRY[103]) );
  NAND2_X2 u5_mult_82_U11554 ( .A1(u5_mult_82_SUMB_52__51_), .A2(
        u5_mult_82_CARRYB_52__50_), .ZN(u5_mult_82_n6439) );
  INV_X4 u5_mult_82_U11553 ( .A(u5_mult_82_n6438), .ZN(u5_mult_82_CLA_SUM[102]) );
  XNOR2_X2 u5_mult_82_U11552 ( .A(u5_mult_82_CARRYB_52__49_), .B(
        u5_mult_82_SUMB_52__50_), .ZN(u5_mult_82_n6438) );
  INV_X4 u5_mult_82_U11551 ( .A(u5_mult_82_n6437), .ZN(
        u5_mult_82_CLA_CARRY[102]) );
  NAND2_X2 u5_mult_82_U11550 ( .A1(u5_mult_82_SUMB_52__50_), .A2(
        u5_mult_82_CARRYB_52__49_), .ZN(u5_mult_82_n6437) );
  INV_X4 u5_mult_82_U11549 ( .A(u5_mult_82_n6436), .ZN(u5_mult_82_CLA_SUM[101]) );
  XNOR2_X2 u5_mult_82_U11548 ( .A(u5_mult_82_CARRYB_52__48_), .B(
        u5_mult_82_SUMB_52__49_), .ZN(u5_mult_82_n6436) );
  INV_X4 u5_mult_82_U11547 ( .A(u5_mult_82_n6435), .ZN(u5_mult_82_CLA_SUM[100]) );
  XNOR2_X2 u5_mult_82_U11546 ( .A(u5_mult_82_CARRYB_52__47_), .B(
        u5_mult_82_SUMB_52__48_), .ZN(u5_mult_82_n6435) );
  INV_X4 u5_mult_82_U11545 ( .A(u5_mult_82_n6434), .ZN(u5_mult_82_CLA_SUM[99])
         );
  XNOR2_X2 u5_mult_82_U11544 ( .A(u5_mult_82_CARRYB_52__46_), .B(
        u5_mult_82_SUMB_52__47_), .ZN(u5_mult_82_n6434) );
  INV_X4 u5_mult_82_U11543 ( .A(u5_mult_82_n6433), .ZN(u5_mult_82_CLA_SUM[98])
         );
  XNOR2_X2 u5_mult_82_U11542 ( .A(u5_mult_82_CARRYB_52__45_), .B(
        u5_mult_82_SUMB_52__46_), .ZN(u5_mult_82_n6433) );
  INV_X4 u5_mult_82_U11541 ( .A(u5_mult_82_n6432), .ZN(u5_mult_82_CLA_SUM[97])
         );
  XNOR2_X2 u5_mult_82_U11540 ( .A(u5_mult_82_CARRYB_52__44_), .B(
        u5_mult_82_SUMB_52__45_), .ZN(u5_mult_82_n6432) );
  INV_X4 u5_mult_82_U11539 ( .A(u5_mult_82_n6431), .ZN(u5_mult_82_CLA_SUM[96])
         );
  XNOR2_X2 u5_mult_82_U11538 ( .A(u5_mult_82_CARRYB_52__43_), .B(
        u5_mult_82_SUMB_52__44_), .ZN(u5_mult_82_n6431) );
  INV_X4 u5_mult_82_U11537 ( .A(u5_mult_82_n6430), .ZN(u5_mult_82_CLA_SUM[95])
         );
  XNOR2_X2 u5_mult_82_U11536 ( .A(u5_mult_82_CARRYB_52__42_), .B(
        u5_mult_82_SUMB_52__43_), .ZN(u5_mult_82_n6430) );
  INV_X4 u5_mult_82_U11535 ( .A(u5_mult_82_n6429), .ZN(u5_mult_82_CLA_SUM[94])
         );
  XNOR2_X2 u5_mult_82_U11534 ( .A(u5_mult_82_CARRYB_52__41_), .B(
        u5_mult_82_SUMB_52__42_), .ZN(u5_mult_82_n6429) );
  INV_X4 u5_mult_82_U11533 ( .A(u5_mult_82_n6428), .ZN(u5_mult_82_CLA_SUM[93])
         );
  XNOR2_X2 u5_mult_82_U11532 ( .A(u5_mult_82_CARRYB_52__40_), .B(
        u5_mult_82_SUMB_52__41_), .ZN(u5_mult_82_n6428) );
  INV_X4 u5_mult_82_U11531 ( .A(u5_mult_82_n6427), .ZN(u5_mult_82_CLA_SUM[92])
         );
  XNOR2_X2 u5_mult_82_U11530 ( .A(u5_mult_82_CARRYB_52__39_), .B(
        u5_mult_82_SUMB_52__40_), .ZN(u5_mult_82_n6427) );
  INV_X4 u5_mult_82_U11529 ( .A(u5_mult_82_n6426), .ZN(u5_mult_82_CLA_SUM[91])
         );
  XNOR2_X2 u5_mult_82_U11528 ( .A(u5_mult_82_CARRYB_52__38_), .B(
        u5_mult_82_SUMB_52__39_), .ZN(u5_mult_82_n6426) );
  INV_X4 u5_mult_82_U11527 ( .A(u5_mult_82_n6425), .ZN(u5_mult_82_CLA_SUM[90])
         );
  XNOR2_X2 u5_mult_82_U11526 ( .A(u5_mult_82_CARRYB_52__37_), .B(
        u5_mult_82_SUMB_52__38_), .ZN(u5_mult_82_n6425) );
  INV_X4 u5_mult_82_U11525 ( .A(u5_mult_82_n6424), .ZN(u5_mult_82_CLA_SUM[89])
         );
  XNOR2_X2 u5_mult_82_U11524 ( .A(u5_mult_82_CARRYB_52__36_), .B(
        u5_mult_82_SUMB_52__37_), .ZN(u5_mult_82_n6424) );
  INV_X4 u5_mult_82_U11523 ( .A(u5_mult_82_n6422), .ZN(u5_mult_82_CLA_SUM[87])
         );
  XNOR2_X2 u5_mult_82_U11522 ( .A(u5_mult_82_CARRYB_52__34_), .B(
        u5_mult_82_SUMB_52__35_), .ZN(u5_mult_82_n6422) );
  INV_X4 u5_mult_82_U11521 ( .A(u5_mult_82_n6421), .ZN(u5_mult_82_CLA_SUM[85])
         );
  XNOR2_X2 u5_mult_82_U11520 ( .A(u5_mult_82_SUMB_52__33_), .B(
        u5_mult_82_CARRYB_52__32_), .ZN(u5_mult_82_n6421) );
  INV_X4 u5_mult_82_U11519 ( .A(u5_mult_82_n6420), .ZN(u5_mult_82_CLA_SUM[84])
         );
  XNOR2_X2 u5_mult_82_U11518 ( .A(u5_mult_82_CARRYB_52__31_), .B(
        u5_mult_82_SUMB_52__32_), .ZN(u5_mult_82_n6420) );
  XNOR2_X2 u5_mult_82_U11517 ( .A(u5_mult_82_CARRYB_52__30_), .B(
        u5_mult_82_SUMB_52__31_), .ZN(u5_mult_82_n6419) );
  XNOR2_X2 u5_mult_82_U11516 ( .A(u5_mult_82_CARRYB_52__29_), .B(
        u5_mult_82_SUMB_52__30_), .ZN(u5_mult_82_n6418) );
  INV_X4 u5_mult_82_U11515 ( .A(u5_mult_82_n6417), .ZN(
        u5_mult_82_CLA_CARRY[82]) );
  NAND2_X2 u5_mult_82_U11514 ( .A1(u5_mult_82_SUMB_52__30_), .A2(
        u5_mult_82_CARRYB_52__29_), .ZN(u5_mult_82_n6417) );
  INV_X4 u5_mult_82_U11513 ( .A(u5_mult_82_n6416), .ZN(u5_mult_82_CLA_SUM[81])
         );
  XNOR2_X2 u5_mult_82_U11512 ( .A(u5_mult_82_CARRYB_52__28_), .B(
        u5_mult_82_SUMB_52__29_), .ZN(u5_mult_82_n6416) );
  NAND2_X2 u5_mult_82_U11511 ( .A1(u5_mult_82_SUMB_52__29_), .A2(
        u5_mult_82_CARRYB_52__28_), .ZN(u5_mult_82_n6415) );
  INV_X4 u5_mult_82_U11510 ( .A(u5_mult_82_n6414), .ZN(u5_mult_82_CLA_SUM[80])
         );
  XNOR2_X2 u5_mult_82_U11509 ( .A(u5_mult_82_CARRYB_52__27_), .B(
        u5_mult_82_SUMB_52__28_), .ZN(u5_mult_82_n6414) );
  XNOR2_X2 u5_mult_82_U11508 ( .A(u5_mult_82_CARRYB_52__26_), .B(
        u5_mult_82_SUMB_52__27_), .ZN(u5_mult_82_n6413) );
  INV_X4 u5_mult_82_U11507 ( .A(u5_mult_82_n6412), .ZN(u5_mult_82_CLA_SUM[78])
         );
  XNOR2_X2 u5_mult_82_U11506 ( .A(u5_mult_82_CARRYB_52__25_), .B(
        u5_mult_82_SUMB_52__26_), .ZN(u5_mult_82_n6412) );
  INV_X4 u5_mult_82_U11505 ( .A(u5_mult_82_n6411), .ZN(u5_mult_82_CLA_SUM[77])
         );
  XNOR2_X2 u5_mult_82_U11504 ( .A(u5_mult_82_CARRYB_52__24_), .B(
        u5_mult_82_SUMB_52__25_), .ZN(u5_mult_82_n6411) );
  XNOR2_X2 u5_mult_82_U11503 ( .A(u5_mult_82_SUMB_52__24_), .B(
        u5_mult_82_CARRYB_52__23_), .ZN(u5_mult_82_n6410) );
  XNOR2_X2 u5_mult_82_U11502 ( .A(u5_mult_82_SUMB_52__23_), .B(
        u5_mult_82_CARRYB_52__22_), .ZN(u5_mult_82_n6409) );
  XNOR2_X2 u5_mult_82_U11501 ( .A(u5_mult_82_CARRYB_52__21_), .B(
        u5_mult_82_SUMB_52__22_), .ZN(u5_mult_82_n6408) );
  XNOR2_X2 u5_mult_82_U11500 ( .A(u5_mult_82_CARRYB_52__20_), .B(
        u5_mult_82_SUMB_52__21_), .ZN(u5_mult_82_n6407) );
  INV_X4 u5_mult_82_U11499 ( .A(u5_mult_82_n6406), .ZN(u5_mult_82_CLA_SUM[72])
         );
  XNOR2_X2 u5_mult_82_U11498 ( .A(u5_mult_82_CARRYB_52__19_), .B(
        u5_mult_82_SUMB_52__20_), .ZN(u5_mult_82_n6406) );
  XNOR2_X2 u5_mult_82_U11497 ( .A(u5_mult_82_CARRYB_52__18_), .B(
        u5_mult_82_SUMB_52__19_), .ZN(u5_mult_82_n6405) );
  INV_X4 u5_mult_82_U11496 ( .A(u5_mult_82_n6404), .ZN(
        u5_mult_82_CLA_CARRY[71]) );
  NAND2_X2 u5_mult_82_U11495 ( .A1(u5_mult_82_SUMB_52__19_), .A2(
        u5_mult_82_CARRYB_52__18_), .ZN(u5_mult_82_n6404) );
  XNOR2_X2 u5_mult_82_U11494 ( .A(u5_mult_82_SUMB_52__18_), .B(
        u5_mult_82_CARRYB_52__17_), .ZN(u5_mult_82_n6403) );
  INV_X4 u5_mult_82_U11493 ( .A(u5_mult_82_n6402), .ZN(u5_mult_82_CLA_SUM[68])
         );
  XNOR2_X2 u5_mult_82_U11492 ( .A(u5_mult_82_SUMB_52__16_), .B(
        u5_mult_82_CARRYB_52__15_), .ZN(u5_mult_82_n6402) );
  INV_X4 u5_mult_82_U11491 ( .A(u5_mult_82_n6401), .ZN(u5_mult_82_CLA_SUM[67])
         );
  XNOR2_X2 u5_mult_82_U11490 ( .A(u5_mult_82_CARRYB_52__14_), .B(
        u5_mult_82_SUMB_52__15_), .ZN(u5_mult_82_n6401) );
  INV_X4 u5_mult_82_U11489 ( .A(u5_mult_82_n6400), .ZN(u5_mult_82_CLA_SUM[66])
         );
  XNOR2_X2 u5_mult_82_U11488 ( .A(u5_mult_82_CARRYB_52__13_), .B(
        u5_mult_82_SUMB_52__14_), .ZN(u5_mult_82_n6400) );
  INV_X4 u5_mult_82_U11487 ( .A(u5_mult_82_n6399), .ZN(
        u5_mult_82_CLA_CARRY[66]) );
  XNOR2_X2 u5_mult_82_U11486 ( .A(u5_mult_82_SUMB_52__12_), .B(
        u5_mult_82_CARRYB_52__11_), .ZN(u5_mult_82_n6398) );
  INV_X4 u5_mult_82_U11485 ( .A(u5_mult_82_n6396), .ZN(u5_mult_82_CLA_SUM[62])
         );
  XNOR2_X2 u5_mult_82_U11484 ( .A(u5_mult_82_SUMB_52__10_), .B(
        u5_mult_82_CARRYB_52__9_), .ZN(u5_mult_82_n6396) );
  XNOR2_X2 u5_mult_82_U11483 ( .A(u5_mult_82_SUMB_52__9_), .B(
        u5_mult_82_CARRYB_52__8_), .ZN(u5_mult_82_n6395) );
  INV_X4 u5_mult_82_U11482 ( .A(u5_mult_82_n6394), .ZN(u5_mult_82_CLA_SUM[60])
         );
  XNOR2_X2 u5_mult_82_U11481 ( .A(u5_mult_82_CARRYB_52__7_), .B(
        u5_mult_82_SUMB_52__8_), .ZN(u5_mult_82_n6394) );
  INV_X4 u5_mult_82_U11480 ( .A(u5_mult_82_n6393), .ZN(u5_mult_82_CLA_SUM[58])
         );
  INV_X4 u5_mult_82_U11479 ( .A(u5_mult_82__UDW__89408_net70938), .ZN(
        u5_mult_82_CLA_SUM[57]) );
  INV_X4 u5_mult_82_U11478 ( .A(u5_mult_82_n6392), .ZN(u5_mult_82_CLA_SUM[56])
         );
  XNOR2_X2 u5_mult_82_U11477 ( .A(u5_mult_82_SUMB_52__4_), .B(
        u5_mult_82_CARRYB_52__3_), .ZN(u5_mult_82_n6392) );
  XNOR2_X2 u5_mult_82_U11476 ( .A(u5_mult_82_SUMB_52__3_), .B(
        u5_mult_82_CARRYB_52__2_), .ZN(u5_mult_82_n6391) );
  NAND2_X2 u5_mult_82_U11475 ( .A1(u5_mult_82_SUMB_52__1_), .A2(
        u5_mult_82_CARRYB_52__0_), .ZN(u5_mult_82_n6389) );
  NOR2_X1 u5_mult_82_U11474 ( .A1(u5_mult_82_n6974), .A2(u5_mult_82_net64361), 
        .ZN(u5_mult_82_ab_52__5_) );
  NOR2_X1 u5_mult_82_U11473 ( .A1(u5_mult_82_n6980), .A2(u5_mult_82_n6524), 
        .ZN(u5_mult_82_ab_4__52_) );
  NAND3_X2 u5_mult_82_U11472 ( .A1(u5_mult_82_net78790), .A2(
        u5_mult_82_net78791), .A3(u5_mult_82_net78792), .ZN(
        u5_mult_82_CARRYB_52__5_) );
  NAND3_X2 u5_mult_82_U11471 ( .A1(u5_mult_82_n6386), .A2(u5_mult_82_n6387), 
        .A3(u5_mult_82_n6388), .ZN(u5_mult_82_CARRYB_5__51_) );
  NAND2_X2 u5_mult_82_U11470 ( .A1(u5_mult_82_ab_5__51_), .A2(
        u5_mult_82_ab_4__52_), .ZN(u5_mult_82_n6388) );
  NAND2_X2 u5_mult_82_U11469 ( .A1(u5_mult_82_ab_5__51_), .A2(
        u5_mult_82_CARRYB_4__51_), .ZN(u5_mult_82_n6387) );
  NAND2_X2 u5_mult_82_U11468 ( .A1(u5_mult_82_ab_4__52_), .A2(
        u5_mult_82_CARRYB_4__51_), .ZN(u5_mult_82_n6386) );
  XOR2_X2 u5_mult_82_U11467 ( .A(u5_mult_82_ab_4__52_), .B(
        u5_mult_82_ab_5__51_), .Z(u5_mult_82_n6385) );
  NAND3_X2 u5_mult_82_U11466 ( .A1(u5_mult_82_n6382), .A2(u5_mult_82_n6383), 
        .A3(u5_mult_82_n6384), .ZN(u5_mult_82_CARRYB_13__44_) );
  NAND2_X1 u5_mult_82_U11465 ( .A1(u5_mult_82_CARRYB_12__44_), .A2(
        u5_mult_82_SUMB_12__45_), .ZN(u5_mult_82_n6384) );
  NAND2_X1 u5_mult_82_U11464 ( .A1(u5_mult_82_ab_13__44_), .A2(
        u5_mult_82_SUMB_12__45_), .ZN(u5_mult_82_n6383) );
  NAND2_X1 u5_mult_82_U11463 ( .A1(u5_mult_82_ab_13__44_), .A2(
        u5_mult_82_CARRYB_12__44_), .ZN(u5_mult_82_n6382) );
  NAND2_X2 u5_mult_82_U11462 ( .A1(u5_mult_82_ab_12__45_), .A2(
        u5_mult_82_n1635), .ZN(u5_mult_82_n6380) );
  NAND2_X1 u5_mult_82_U11461 ( .A1(u5_mult_82_ab_12__45_), .A2(
        u5_mult_82_CARRYB_11__45_), .ZN(u5_mult_82_n6379) );
  XOR2_X2 u5_mult_82_U11460 ( .A(u5_mult_82_n6378), .B(u5_mult_82_n1635), .Z(
        u5_mult_82_SUMB_12__45_) );
  NAND2_X1 u5_mult_82_U11459 ( .A1(u5_mult_82_ab_23__34_), .A2(
        u5_mult_82_n5507), .ZN(u5_mult_82_n6375) );
  NAND2_X2 u5_mult_82_U11458 ( .A1(u5_mult_82_CARRYB_21__35_), .A2(
        u5_mult_82_SUMB_21__36_), .ZN(u5_mult_82_n6374) );
  NAND2_X2 u5_mult_82_U11457 ( .A1(u5_mult_82_ab_22__35_), .A2(
        u5_mult_82_SUMB_21__36_), .ZN(u5_mult_82_n6373) );
  NAND2_X1 u5_mult_82_U11456 ( .A1(u5_mult_82_ab_22__35_), .A2(
        u5_mult_82_CARRYB_21__35_), .ZN(u5_mult_82_n6372) );
  NAND3_X2 u5_mult_82_U11455 ( .A1(u5_mult_82_n6368), .A2(u5_mult_82_n6369), 
        .A3(u5_mult_82_n6370), .ZN(u5_mult_82_CARRYB_33__24_) );
  NAND2_X1 u5_mult_82_U11454 ( .A1(u5_mult_82_CARRYB_32__24_), .A2(
        u5_mult_82_SUMB_32__25_), .ZN(u5_mult_82_n6370) );
  NAND2_X1 u5_mult_82_U11453 ( .A1(u5_mult_82_ab_33__24_), .A2(
        u5_mult_82_SUMB_32__25_), .ZN(u5_mult_82_n6369) );
  NAND2_X1 u5_mult_82_U11452 ( .A1(u5_mult_82_ab_33__24_), .A2(
        u5_mult_82_CARRYB_32__24_), .ZN(u5_mult_82_n6368) );
  NAND2_X2 u5_mult_82_U11451 ( .A1(u5_mult_82_SUMB_31__26_), .A2(
        u5_mult_82_CARRYB_31__25_), .ZN(u5_mult_82_n6367) );
  NAND2_X2 u5_mult_82_U11450 ( .A1(u5_mult_82_ab_32__25_), .A2(
        u5_mult_82_SUMB_31__26_), .ZN(u5_mult_82_n6366) );
  NAND2_X1 u5_mult_82_U11449 ( .A1(u5_mult_82_ab_32__25_), .A2(
        u5_mult_82_CARRYB_31__25_), .ZN(u5_mult_82_n6365) );
  XOR2_X2 u5_mult_82_U11448 ( .A(u5_mult_82_n6364), .B(u5_mult_82_n1564), .Z(
        u5_mult_82_SUMB_32__25_) );
  XOR2_X2 u5_mult_82_U11447 ( .A(u5_mult_82_ab_32__25_), .B(
        u5_mult_82_CARRYB_31__25_), .Z(u5_mult_82_n6364) );
  NAND2_X1 u5_mult_82_U11446 ( .A1(u5_mult_82_ab_43__14_), .A2(
        u5_mult_82_CARRYB_42__14_), .ZN(u5_mult_82_n6361) );
  NAND2_X2 u5_mult_82_U11445 ( .A1(u5_mult_82_CARRYB_41__15_), .A2(
        u5_mult_82_SUMB_41__16_), .ZN(u5_mult_82_n6360) );
  NAND2_X2 u5_mult_82_U11444 ( .A1(u5_mult_82_ab_42__15_), .A2(
        u5_mult_82_SUMB_41__16_), .ZN(u5_mult_82_n6359) );
  NAND3_X2 u5_mult_82_U11443 ( .A1(u5_mult_82_n6357), .A2(u5_mult_82_n6356), 
        .A3(u5_mult_82_n6355), .ZN(u5_mult_82_CARRYB_10__44_) );
  NAND2_X1 u5_mult_82_U11442 ( .A1(u5_mult_82_CARRYB_9__44_), .A2(
        u5_mult_82_SUMB_9__45_), .ZN(u5_mult_82_n6357) );
  NAND2_X1 u5_mult_82_U11441 ( .A1(u5_mult_82_ab_10__44_), .A2(
        u5_mult_82_CARRYB_9__44_), .ZN(u5_mult_82_n6355) );
  NAND3_X2 u5_mult_82_U11440 ( .A1(u5_mult_82_n6352), .A2(u5_mult_82_n6353), 
        .A3(u5_mult_82_n6354), .ZN(u5_mult_82_CARRYB_9__45_) );
  NAND2_X2 u5_mult_82_U11439 ( .A1(u5_mult_82_ab_9__45_), .A2(u5_mult_82_n1853), .ZN(u5_mult_82_n6353) );
  XOR2_X2 u5_mult_82_U11438 ( .A(u5_mult_82_n6351), .B(u5_mult_82_n1853), .Z(
        u5_mult_82_SUMB_9__45_) );
  XOR2_X2 u5_mult_82_U11437 ( .A(u5_mult_82_ab_9__45_), .B(
        u5_mult_82_CARRYB_8__45_), .Z(u5_mult_82_n6351) );
  NAND3_X2 u5_mult_82_U11436 ( .A1(u5_mult_82_n6348), .A2(u5_mult_82_n6349), 
        .A3(u5_mult_82_n6350), .ZN(u5_mult_82_CARRYB_6__48_) );
  NAND2_X1 u5_mult_82_U11435 ( .A1(u5_mult_82_SUMB_5__49_), .A2(
        u5_mult_82_CARRYB_5__48_), .ZN(u5_mult_82_n6350) );
  NAND2_X1 u5_mult_82_U11434 ( .A1(u5_mult_82_ab_6__48_), .A2(
        u5_mult_82_CARRYB_5__48_), .ZN(u5_mult_82_n6348) );
  NAND3_X2 u5_mult_82_U11433 ( .A1(u5_mult_82_n6345), .A2(u5_mult_82_n6346), 
        .A3(u5_mult_82_n6347), .ZN(u5_mult_82_CARRYB_5__49_) );
  NAND2_X1 u5_mult_82_U11432 ( .A1(u5_mult_82_ab_23__31_), .A2(
        u5_mult_82_CARRYB_22__31_), .ZN(u5_mult_82_n6342) );
  NAND2_X2 u5_mult_82_U11431 ( .A1(u5_mult_82_SUMB_21__33_), .A2(
        u5_mult_82_CARRYB_21__32_), .ZN(u5_mult_82_n6341) );
  NAND2_X2 u5_mult_82_U11430 ( .A1(u5_mult_82_ab_22__32_), .A2(
        u5_mult_82_SUMB_21__33_), .ZN(u5_mult_82_n6340) );
  NAND2_X1 u5_mult_82_U11429 ( .A1(u5_mult_82_ab_22__32_), .A2(
        u5_mult_82_CARRYB_21__32_), .ZN(u5_mult_82_n6339) );
  NAND3_X2 u5_mult_82_U11428 ( .A1(u5_mult_82_n6338), .A2(u5_mult_82_n6337), 
        .A3(u5_mult_82_n6336), .ZN(u5_mult_82_CARRYB_35__19_) );
  NAND2_X2 u5_mult_82_U11427 ( .A1(u5_mult_82_CARRYB_33__20_), .A2(
        u5_mult_82_n1399), .ZN(u5_mult_82_n6335) );
  NAND2_X2 u5_mult_82_U11426 ( .A1(u5_mult_82_ab_34__20_), .A2(
        u5_mult_82_n1399), .ZN(u5_mult_82_n6334) );
  XOR2_X2 u5_mult_82_U11425 ( .A(u5_mult_82_n6332), .B(u5_mult_82_SUMB_34__20_), .Z(u5_mult_82_SUMB_35__19_) );
  XOR2_X2 u5_mult_82_U11424 ( .A(u5_mult_82_n6331), .B(u5_mult_82_n1399), .Z(
        u5_mult_82_SUMB_34__20_) );
  XOR2_X2 u5_mult_82_U11423 ( .A(u5_mult_82_ab_34__20_), .B(
        u5_mult_82_CARRYB_33__20_), .Z(u5_mult_82_n6331) );
  NAND3_X2 u5_mult_82_U11422 ( .A1(u5_mult_82_n6329), .A2(u5_mult_82_n6328), 
        .A3(u5_mult_82_n6330), .ZN(u5_mult_82_CARRYB_50__4_) );
  NAND2_X1 u5_mult_82_U11421 ( .A1(u5_mult_82_CARRYB_49__4_), .A2(
        u5_mult_82_SUMB_49__5_), .ZN(u5_mult_82_n6330) );
  NAND2_X1 u5_mult_82_U11420 ( .A1(u5_mult_82_ab_50__4_), .A2(
        u5_mult_82_SUMB_49__5_), .ZN(u5_mult_82_n6329) );
  NAND2_X1 u5_mult_82_U11419 ( .A1(u5_mult_82_ab_50__4_), .A2(
        u5_mult_82_CARRYB_49__4_), .ZN(u5_mult_82_n6328) );
  NAND2_X2 u5_mult_82_U11418 ( .A1(u5_mult_82_CARRYB_48__5_), .A2(
        u5_mult_82_SUMB_48__6_), .ZN(u5_mult_82_n6327) );
  NAND2_X1 u5_mult_82_U11417 ( .A1(u5_mult_82_ab_49__5_), .A2(
        u5_mult_82_CARRYB_48__5_), .ZN(u5_mult_82_n6325) );
  NAND2_X2 u5_mult_82_U11416 ( .A1(u5_mult_82_ab_5__49_), .A2(
        u5_mult_82_CARRYB_4__49_), .ZN(u5_mult_82_n6345) );
  NOR2_X2 u5_mult_82_U11415 ( .A1(u5_mult_82_n6775), .A2(u5_mult_82_n6520), 
        .ZN(u5_mult_82_ab_4__49_) );
  NOR2_X1 u5_mult_82_U11414 ( .A1(u5_mult_82_net64939), .A2(u5_mult_82_n6594), 
        .ZN(u5_mult_82_ab_16__37_) );
  NOR2_X1 u5_mult_82_U11413 ( .A1(u5_mult_82_n6891), .A2(u5_mult_82_n6672), 
        .ZN(u5_mult_82_ab_29__24_) );
  NAND3_X2 u5_mult_82_U11412 ( .A1(u5_mult_82_n6322), .A2(u5_mult_82_n6323), 
        .A3(u5_mult_82_n6324), .ZN(u5_mult_82_CARRYB_7__46_) );
  NAND2_X1 u5_mult_82_U11411 ( .A1(u5_mult_82_CARRYB_6__46_), .A2(
        u5_mult_82_SUMB_6__47_), .ZN(u5_mult_82_n6324) );
  NAND2_X1 u5_mult_82_U11410 ( .A1(u5_mult_82_ab_7__46_), .A2(
        u5_mult_82_SUMB_6__47_), .ZN(u5_mult_82_n6323) );
  NAND2_X2 u5_mult_82_U11409 ( .A1(u5_mult_82_ab_6__47_), .A2(u5_mult_82_n1822), .ZN(u5_mult_82_n6320) );
  NAND3_X2 u5_mult_82_U11408 ( .A1(u5_mult_82_n6316), .A2(u5_mult_82_n6317), 
        .A3(u5_mult_82_n6318), .ZN(u5_mult_82_CARRYB_4__49_) );
  NAND2_X1 u5_mult_82_U11407 ( .A1(u5_mult_82_ab_18__35_), .A2(
        u5_mult_82_CARRYB_17__35_), .ZN(u5_mult_82_n6313) );
  NAND2_X2 u5_mult_82_U11406 ( .A1(u5_mult_82_SUMB_16__37_), .A2(
        u5_mult_82_CARRYB_16__36_), .ZN(u5_mult_82_n6312) );
  NAND2_X2 u5_mult_82_U11405 ( .A1(u5_mult_82_ab_17__36_), .A2(
        u5_mult_82_SUMB_16__37_), .ZN(u5_mult_82_n6311) );
  XOR2_X2 u5_mult_82_U11404 ( .A(u5_mult_82_n6309), .B(u5_mult_82_SUMB_17__36_), .Z(u5_mult_82_SUMB_18__35_) );
  NAND3_X2 u5_mult_82_U11403 ( .A1(u5_mult_82_n6305), .A2(u5_mult_82_n6306), 
        .A3(u5_mult_82_n6307), .ZN(u5_mult_82_CARRYB_16__37_) );
  NAND2_X1 u5_mult_82_U11402 ( .A1(u5_mult_82_ab_31__22_), .A2(
        u5_mult_82_CARRYB_30__22_), .ZN(u5_mult_82_n6302) );
  NAND2_X2 u5_mult_82_U11401 ( .A1(u5_mult_82_CARRYB_29__23_), .A2(
        u5_mult_82_SUMB_29__24_), .ZN(u5_mult_82_n6301) );
  NAND2_X2 u5_mult_82_U11400 ( .A1(u5_mult_82_ab_30__23_), .A2(
        u5_mult_82_SUMB_29__24_), .ZN(u5_mult_82_n6300) );
  NAND2_X1 u5_mult_82_U11399 ( .A1(u5_mult_82_ab_30__23_), .A2(
        u5_mult_82_CARRYB_29__23_), .ZN(u5_mult_82_n6299) );
  NAND3_X2 u5_mult_82_U11398 ( .A1(u5_mult_82_n6295), .A2(u5_mult_82_n6296), 
        .A3(u5_mult_82_n6297), .ZN(u5_mult_82_CARRYB_29__24_) );
  NAND2_X1 u5_mult_82_U11397 ( .A1(u5_mult_82_ab_29__24_), .A2(
        u5_mult_82_CARRYB_28__24_), .ZN(u5_mult_82_n6297) );
  XOR2_X2 u5_mult_82_U11396 ( .A(u5_mult_82_SUMB_28__25_), .B(u5_mult_82_n6294), .Z(u5_mult_82_SUMB_29__24_) );
  XOR2_X2 u5_mult_82_U11395 ( .A(u5_mult_82_CARRYB_28__24_), .B(
        u5_mult_82_ab_29__24_), .Z(u5_mult_82_n6294) );
  NAND3_X2 u5_mult_82_U11394 ( .A1(u5_mult_82_net78850), .A2(
        u5_mult_82_net78851), .A3(u5_mult_82_net78852), .ZN(
        u5_mult_82_CARRYB_42__11_) );
  NOR2_X2 u5_mult_82_U11393 ( .A1(u5_mult_82_n6769), .A2(u5_mult_82_net66033), 
        .ZN(u5_mult_82_ab_5__50_) );
  NOR2_X1 u5_mult_82_U11392 ( .A1(u5_mult_82_n6769), .A2(u5_mult_82_n1359), 
        .ZN(u5_mult_82_ab_6__50_) );
  NOR2_X1 u5_mult_82_U11391 ( .A1(u5_mult_82_n6828), .A2(u5_mult_82_n6593), 
        .ZN(u5_mult_82_ab_16__40_) );
  NOR2_X1 u5_mult_82_U11390 ( .A1(u5_mult_82_n6904), .A2(u5_mult_82_n6715), 
        .ZN(u5_mult_82_ab_36__20_) );
  NAND2_X1 u5_mult_82_U11389 ( .A1(u5_mult_82_CARRYB_4__50_), .A2(
        u5_mult_82_SUMB_4__51_), .ZN(u5_mult_82_n6291) );
  NAND3_X2 u5_mult_82_U11388 ( .A1(u5_mult_82_n6288), .A2(u5_mult_82_n6289), 
        .A3(u5_mult_82_n6290), .ZN(u5_mult_82_CARRYB_6__50_) );
  NAND2_X2 u5_mult_82_U11387 ( .A1(u5_mult_82_ab_6__50_), .A2(
        u5_mult_82_SUMB_5__51_), .ZN(u5_mult_82_n6290) );
  NAND2_X2 u5_mult_82_U11386 ( .A1(u5_mult_82_ab_6__50_), .A2(
        u5_mult_82_CARRYB_5__50_), .ZN(u5_mult_82_n6289) );
  NAND3_X2 u5_mult_82_U11385 ( .A1(u5_mult_82_n6285), .A2(u5_mult_82_n6286), 
        .A3(u5_mult_82_n6287), .ZN(u5_mult_82_CARRYB_16__40_) );
  NAND2_X2 u5_mult_82_U11384 ( .A1(u5_mult_82_ab_16__40_), .A2(
        u5_mult_82_SUMB_15__41_), .ZN(u5_mult_82_n6286) );
  NAND2_X1 u5_mult_82_U11383 ( .A1(u5_mult_82_CARRYB_15__40_), .A2(
        u5_mult_82_SUMB_15__41_), .ZN(u5_mult_82_n6285) );
  NAND3_X2 u5_mult_82_U11382 ( .A1(u5_mult_82_n6279), .A2(u5_mult_82_n6280), 
        .A3(u5_mult_82_n6281), .ZN(u5_mult_82_CARRYB_26__30_) );
  NAND2_X2 u5_mult_82_U11381 ( .A1(u5_mult_82_ab_26__30_), .A2(
        u5_mult_82_SUMB_25__31_), .ZN(u5_mult_82_n6280) );
  NAND2_X1 u5_mult_82_U11380 ( .A1(u5_mult_82_ab_26__30_), .A2(
        u5_mult_82_CARRYB_25__30_), .ZN(u5_mult_82_n6279) );
  XOR2_X2 u5_mult_82_U11379 ( .A(u5_mult_82_n6278), .B(u5_mult_82_SUMB_25__31_), .Z(u5_mult_82_SUMB_26__30_) );
  NAND3_X2 u5_mult_82_U11378 ( .A1(u5_mult_82_n6275), .A2(u5_mult_82_n6276), 
        .A3(u5_mult_82_n6277), .ZN(u5_mult_82_CARRYB_36__20_) );
  NAND2_X2 u5_mult_82_U11377 ( .A1(u5_mult_82_ab_36__20_), .A2(
        u5_mult_82_SUMB_35__21_), .ZN(u5_mult_82_n6276) );
  NAND2_X1 u5_mult_82_U11376 ( .A1(u5_mult_82_CARRYB_35__20_), .A2(
        u5_mult_82_SUMB_35__21_), .ZN(u5_mult_82_n6275) );
  XOR2_X2 u5_mult_82_U11375 ( .A(u5_mult_82_SUMB_35__21_), .B(u5_mult_82_n6274), .Z(u5_mult_82_SUMB_36__20_) );
  XOR2_X2 u5_mult_82_U11374 ( .A(u5_mult_82_CARRYB_35__20_), .B(
        u5_mult_82_ab_36__20_), .Z(u5_mult_82_n6274) );
  NAND3_X2 u5_mult_82_U11373 ( .A1(u5_mult_82_n6270), .A2(u5_mult_82_n6269), 
        .A3(u5_mult_82_n6268), .ZN(u5_mult_82_CARRYB_29__27_) );
  NAND2_X2 u5_mult_82_U11372 ( .A1(u5_mult_82_n20), .A2(u5_mult_82_ab_29__27_), 
        .ZN(u5_mult_82_n6269) );
  NAND2_X1 u5_mult_82_U11371 ( .A1(u5_mult_82_ab_29__27_), .A2(
        u5_mult_82_CARRYB_28__27_), .ZN(u5_mult_82_n6268) );
  NAND3_X2 u5_mult_82_U11370 ( .A1(u5_mult_82_n6265), .A2(u5_mult_82_n6266), 
        .A3(u5_mult_82_n6267), .ZN(u5_mult_82_CARRYB_47__9_) );
  NAND2_X1 u5_mult_82_U11369 ( .A1(u5_mult_82_CARRYB_46__9_), .A2(
        u5_mult_82_SUMB_46__10_), .ZN(u5_mult_82_n6267) );
  NAND2_X1 u5_mult_82_U11368 ( .A1(u5_mult_82_ab_47__9_), .A2(
        u5_mult_82_SUMB_46__10_), .ZN(u5_mult_82_n6266) );
  NAND2_X1 u5_mult_82_U11367 ( .A1(u5_mult_82_ab_47__9_), .A2(
        u5_mult_82_CARRYB_46__9_), .ZN(u5_mult_82_n6265) );
  NAND3_X2 u5_mult_82_U11366 ( .A1(u5_mult_82_n534), .A2(u5_mult_82_n6259), 
        .A3(u5_mult_82_n6260), .ZN(u5_mult_82_CARRYB_43__13_) );
  NAND2_X1 u5_mult_82_U11365 ( .A1(u5_mult_82_CARRYB_42__13_), .A2(
        u5_mult_82_SUMB_42__14_), .ZN(u5_mult_82_n6260) );
  NAND2_X1 u5_mult_82_U11364 ( .A1(u5_mult_82_ab_43__13_), .A2(
        u5_mult_82_SUMB_42__14_), .ZN(u5_mult_82_n6259) );
  NAND3_X4 u5_mult_82_U11363 ( .A1(u5_mult_82_n6256), .A2(u5_mult_82_n6257), 
        .A3(u5_mult_82_n6258), .ZN(u5_mult_82_CARRYB_42__14_) );
  NAND2_X2 u5_mult_82_U11362 ( .A1(u5_mult_82_CARRYB_41__14_), .A2(
        u5_mult_82_SUMB_41__15_), .ZN(u5_mult_82_n6258) );
  NAND2_X2 u5_mult_82_U11361 ( .A1(u5_mult_82_ab_42__14_), .A2(
        u5_mult_82_SUMB_41__15_), .ZN(u5_mult_82_n6257) );
  NAND2_X1 u5_mult_82_U11360 ( .A1(u5_mult_82_ab_42__14_), .A2(
        u5_mult_82_CARRYB_41__14_), .ZN(u5_mult_82_n6256) );
  NAND3_X2 u5_mult_82_U11359 ( .A1(u5_mult_82_n6253), .A2(u5_mult_82_n6254), 
        .A3(u5_mult_82_n6255), .ZN(u5_mult_82_CARRYB_29__26_) );
  NAND2_X1 u5_mult_82_U11358 ( .A1(u5_mult_82_SUMB_28__27_), .A2(
        u5_mult_82_n1515), .ZN(u5_mult_82_n6255) );
  NAND2_X1 u5_mult_82_U11357 ( .A1(u5_mult_82_ab_29__26_), .A2(
        u5_mult_82_SUMB_28__27_), .ZN(u5_mult_82_n6254) );
  NAND2_X1 u5_mult_82_U11356 ( .A1(u5_mult_82_ab_29__26_), .A2(
        u5_mult_82_n1515), .ZN(u5_mult_82_n6253) );
  NAND2_X2 u5_mult_82_U11355 ( .A1(u5_mult_82_n1715), .A2(
        u5_mult_82_SUMB_27__28_), .ZN(u5_mult_82_n6252) );
  NAND2_X2 u5_mult_82_U11354 ( .A1(u5_mult_82_ab_28__27_), .A2(
        u5_mult_82_SUMB_27__28_), .ZN(u5_mult_82_n6251) );
  NAND2_X1 u5_mult_82_U11353 ( .A1(u5_mult_82_ab_28__27_), .A2(
        u5_mult_82_CARRYB_27__27_), .ZN(u5_mult_82_n6250) );
  XOR2_X2 u5_mult_82_U11352 ( .A(u5_mult_82_n6249), .B(u5_mult_82_SUMB_28__27_), .Z(u5_mult_82_SUMB_29__26_) );
  XOR2_X2 u5_mult_82_U11351 ( .A(u5_mult_82_n6248), .B(u5_mult_82_SUMB_27__28_), .Z(u5_mult_82_SUMB_28__27_) );
  XOR2_X2 u5_mult_82_U11350 ( .A(u5_mult_82_ab_28__27_), .B(
        u5_mult_82_CARRYB_27__27_), .Z(u5_mult_82_n6248) );
  NAND2_X1 u5_mult_82_U11349 ( .A1(u5_mult_82_ab_48__7_), .A2(
        u5_mult_82_CARRYB_47__7_), .ZN(u5_mult_82_net78954) );
  XNOR2_X2 u5_mult_82_U11348 ( .A(u5_mult_82_CARRYB_52__5_), .B(
        u5_mult_82_SUMB_52__6_), .ZN(u5_mult_82_n6393) );
  XNOR2_X2 u5_mult_82_U11347 ( .A(u5_mult_82_CARRYB_49__4_), .B(
        u5_mult_82_ab_50__4_), .ZN(u5_mult_82_n6247) );
  XNOR2_X2 u5_mult_82_U11346 ( .A(u5_mult_82_n6247), .B(u5_mult_82_SUMB_49__5_), .ZN(u5_mult_82_SUMB_50__4_) );
  NOR2_X2 u5_mult_82_U11345 ( .A1(u5_mult_82_net64487), .A2(
        u5_mult_82_net65283), .ZN(u5_mult_82_ab_47__12_) );
  NAND2_X1 u5_mult_82_U11344 ( .A1(u5_mult_82_ab_15__40_), .A2(
        u5_mult_82_CARRYB_14__40_), .ZN(u5_mult_82_n6244) );
  NAND3_X2 u5_mult_82_U11343 ( .A1(u5_mult_82_n6243), .A2(u5_mult_82_n6242), 
        .A3(u5_mult_82_n6241), .ZN(u5_mult_82_CARRYB_14__41_) );
  NAND2_X2 u5_mult_82_U11342 ( .A1(u5_mult_82_CARRYB_13__41_), .A2(
        u5_mult_82_SUMB_13__42_), .ZN(u5_mult_82_n6243) );
  NAND2_X2 u5_mult_82_U11341 ( .A1(u5_mult_82_ab_14__41_), .A2(
        u5_mult_82_SUMB_13__42_), .ZN(u5_mult_82_n6242) );
  NAND2_X1 u5_mult_82_U11340 ( .A1(u5_mult_82_ab_14__41_), .A2(
        u5_mult_82_CARRYB_13__41_), .ZN(u5_mult_82_n6241) );
  XOR2_X2 u5_mult_82_U11339 ( .A(u5_mult_82_n6240), .B(u5_mult_82_n745), .Z(
        u5_mult_82_SUMB_14__41_) );
  XOR2_X2 u5_mult_82_U11338 ( .A(u5_mult_82_ab_14__41_), .B(
        u5_mult_82_CARRYB_13__41_), .Z(u5_mult_82_n6240) );
  NAND3_X2 u5_mult_82_U11337 ( .A1(u5_mult_82_n6237), .A2(u5_mult_82_n6238), 
        .A3(u5_mult_82_n6239), .ZN(u5_mult_82_CARRYB_49__10_) );
  NAND2_X1 u5_mult_82_U11336 ( .A1(u5_mult_82_ab_49__10_), .A2(
        u5_mult_82_SUMB_48__11_), .ZN(u5_mult_82_n6238) );
  NAND2_X1 u5_mult_82_U11335 ( .A1(u5_mult_82_ab_49__10_), .A2(
        u5_mult_82_CARRYB_48__10_), .ZN(u5_mult_82_n6237) );
  NAND2_X2 u5_mult_82_U11334 ( .A1(u5_mult_82_CARRYB_47__11_), .A2(
        u5_mult_82_SUMB_47__12_), .ZN(u5_mult_82_n6236) );
  NAND2_X2 u5_mult_82_U11333 ( .A1(u5_mult_82_ab_48__11_), .A2(
        u5_mult_82_CARRYB_47__11_), .ZN(u5_mult_82_n6234) );
  NAND2_X1 u5_mult_82_U11332 ( .A1(u5_mult_82_n369), .A2(
        u5_mult_82_SUMB_46__13_), .ZN(u5_mult_82_n6231) );
  XOR2_X2 u5_mult_82_U11331 ( .A(u5_mult_82_SUMB_46__13_), .B(u5_mult_82_n6230), .Z(u5_mult_82_SUMB_47__12_) );
  NOR2_X1 u5_mult_82_U11330 ( .A1(u5_mult_82_n6817), .A2(u5_mult_82_n6593), 
        .ZN(u5_mult_82_ab_16__42_) );
  NAND2_X2 u5_mult_82_U11329 ( .A1(u5_mult_82_ab_24__34_), .A2(
        u5_mult_82_CARRYB_23__34_), .ZN(u5_mult_82_n6224) );
  NAND3_X2 u5_mult_82_U11328 ( .A1(u5_mult_82_n6220), .A2(u5_mult_82_n6221), 
        .A3(u5_mult_82_n6222), .ZN(u5_mult_82_CARRYB_16__42_) );
  NAND2_X2 u5_mult_82_U11327 ( .A1(u5_mult_82_ab_16__42_), .A2(
        u5_mult_82_SUMB_15__43_), .ZN(u5_mult_82_n6221) );
  NAND2_X1 u5_mult_82_U11326 ( .A1(u5_mult_82_CARRYB_15__42_), .A2(
        u5_mult_82_SUMB_15__43_), .ZN(u5_mult_82_n6220) );
  XOR2_X2 u5_mult_82_U11325 ( .A(u5_mult_82_SUMB_15__43_), .B(u5_mult_82_n6219), .Z(u5_mult_82_SUMB_16__42_) );
  NAND3_X2 u5_mult_82_U11324 ( .A1(u5_mult_82_n6216), .A2(u5_mult_82_n6217), 
        .A3(u5_mult_82_n6218), .ZN(u5_mult_82_CARRYB_36__22_) );
  NAND3_X2 u5_mult_82_U11323 ( .A1(u5_mult_82_n6215), .A2(u5_mult_82_n6214), 
        .A3(u5_mult_82_n6213), .ZN(u5_mult_82_CARRYB_35__23_) );
  NAND2_X1 u5_mult_82_U11322 ( .A1(u5_mult_82_ab_35__23_), .A2(
        u5_mult_82_CARRYB_34__23_), .ZN(u5_mult_82_n6213) );
  XOR2_X2 u5_mult_82_U11321 ( .A(u5_mult_82_n6212), .B(u5_mult_82_n82), .Z(
        u5_mult_82_SUMB_35__23_) );
  NAND3_X2 u5_mult_82_U11320 ( .A1(u5_mult_82_n6209), .A2(u5_mult_82_n6210), 
        .A3(u5_mult_82_n6211), .ZN(u5_mult_82_CARRYB_48__10_) );
  NAND2_X1 u5_mult_82_U11319 ( .A1(u5_mult_82_ab_48__10_), .A2(
        u5_mult_82_SUMB_47__11_), .ZN(u5_mult_82_n6210) );
  NAND2_X1 u5_mult_82_U11318 ( .A1(u5_mult_82_ab_47__11_), .A2(
        u5_mult_82_CARRYB_46__11_), .ZN(u5_mult_82_n6206) );
  NAND3_X2 u5_mult_82_U11317 ( .A1(u5_mult_82_n6202), .A2(u5_mult_82_n6203), 
        .A3(u5_mult_82_n6204), .ZN(u5_mult_82_CARRYB_51__7_) );
  NAND2_X1 u5_mult_82_U11316 ( .A1(u5_mult_82_CARRYB_50__7_), .A2(
        u5_mult_82_SUMB_50__8_), .ZN(u5_mult_82_n6204) );
  NAND2_X1 u5_mult_82_U11315 ( .A1(u5_mult_82_ab_51__7_), .A2(
        u5_mult_82_SUMB_50__8_), .ZN(u5_mult_82_n6203) );
  NAND2_X2 u5_mult_82_U11314 ( .A1(u5_mult_82_CARRYB_49__8_), .A2(
        u5_mult_82_SUMB_49__9_), .ZN(u5_mult_82_n6201) );
  NAND2_X1 u5_mult_82_U11313 ( .A1(u5_mult_82_ab_50__8_), .A2(
        u5_mult_82_CARRYB_49__8_), .ZN(u5_mult_82_n6199) );
  NAND2_X2 u5_mult_82_U11312 ( .A1(u5_mult_82_ab_7__46_), .A2(
        u5_mult_82_CARRYB_6__46_), .ZN(u5_mult_82_n6322) );
  NOR2_X2 u5_mult_82_U11311 ( .A1(u5_mult_82_n6793), .A2(u5_mult_82_net66021), 
        .ZN(u5_mult_82_ab_6__46_) );
  NAND2_X2 u5_mult_82_U11310 ( .A1(u5_mult_82_ab_6__47_), .A2(
        u5_mult_82_CARRYB_5__47_), .ZN(u5_mult_82_n6319) );
  NOR2_X2 u5_mult_82_U11309 ( .A1(u5_mult_82_n6786), .A2(u5_mult_82_net66033), 
        .ZN(u5_mult_82_ab_5__47_) );
  NOR2_X2 u5_mult_82_U11308 ( .A1(u5_mult_82_net64455), .A2(
        u5_mult_82_net65373), .ZN(u5_mult_82_ab_42__10_) );
  NAND3_X4 u5_mult_82_U11307 ( .A1(u5_mult_82_n6196), .A2(u5_mult_82_n6197), 
        .A3(u5_mult_82_n6198), .ZN(u5_mult_82_CARRYB_6__46_) );
  NAND2_X2 u5_mult_82_U11306 ( .A1(u5_mult_82_ab_6__46_), .A2(
        u5_mult_82_CARRYB_5__46_), .ZN(u5_mult_82_n6198) );
  NAND2_X2 u5_mult_82_U11305 ( .A1(u5_mult_82_ab_6__46_), .A2(
        u5_mult_82_SUMB_5__47_), .ZN(u5_mult_82_n6197) );
  NAND2_X2 u5_mult_82_U11304 ( .A1(u5_mult_82_n736), .A2(
        u5_mult_82_SUMB_5__47_), .ZN(u5_mult_82_n6196) );
  NAND3_X2 u5_mult_82_U11303 ( .A1(u5_mult_82_n6193), .A2(u5_mult_82_n6194), 
        .A3(u5_mult_82_n6195), .ZN(u5_mult_82_CARRYB_5__47_) );
  NAND2_X1 u5_mult_82_U11302 ( .A1(u5_mult_82_CARRYB_4__47_), .A2(
        u5_mult_82_SUMB_4__48_), .ZN(u5_mult_82_n6193) );
  NAND3_X2 u5_mult_82_U11301 ( .A1(u5_mult_82_n6190), .A2(u5_mult_82_n6191), 
        .A3(u5_mult_82_n6192), .ZN(u5_mult_82_CARRYB_17__35_) );
  NAND2_X1 u5_mult_82_U11300 ( .A1(u5_mult_82_ab_17__35_), .A2(
        u5_mult_82_SUMB_16__36_), .ZN(u5_mult_82_n6191) );
  NAND2_X1 u5_mult_82_U11299 ( .A1(u5_mult_82_ab_17__35_), .A2(
        u5_mult_82_CARRYB_16__35_), .ZN(u5_mult_82_n6190) );
  NAND3_X2 u5_mult_82_U11298 ( .A1(u5_mult_82_n6180), .A2(u5_mult_82_n6181), 
        .A3(u5_mult_82_n6182), .ZN(u5_mult_82_CARRYB_26__26_) );
  NAND2_X2 u5_mult_82_U11297 ( .A1(u5_mult_82_CARRYB_25__26_), .A2(
        u5_mult_82_SUMB_25__27_), .ZN(u5_mult_82_n6182) );
  NAND2_X2 u5_mult_82_U11296 ( .A1(u5_mult_82_ab_26__26_), .A2(
        u5_mult_82_SUMB_25__27_), .ZN(u5_mult_82_n6181) );
  NAND2_X1 u5_mult_82_U11295 ( .A1(u5_mult_82_ab_26__26_), .A2(
        u5_mult_82_CARRYB_25__26_), .ZN(u5_mult_82_n6180) );
  XOR2_X2 u5_mult_82_U11294 ( .A(u5_mult_82_n6179), .B(u5_mult_82_n60), .Z(
        u5_mult_82_SUMB_26__26_) );
  XOR2_X2 u5_mult_82_U11293 ( .A(u5_mult_82_ab_26__26_), .B(
        u5_mult_82_CARRYB_25__26_), .Z(u5_mult_82_n6179) );
  NAND2_X1 u5_mult_82_U11292 ( .A1(u5_mult_82_ab_36__16_), .A2(
        u5_mult_82_CARRYB_35__16_), .ZN(u5_mult_82_n6173) );
  XOR2_X2 u5_mult_82_U11291 ( .A(u5_mult_82_n6172), .B(u5_mult_82_SUMB_35__17_), .Z(u5_mult_82_SUMB_36__16_) );
  XOR2_X2 u5_mult_82_U11290 ( .A(u5_mult_82_ab_36__16_), .B(
        u5_mult_82_CARRYB_35__16_), .Z(u5_mult_82_n6172) );
  NAND2_X1 u5_mult_82_U11289 ( .A1(u5_mult_82_ab_47__5_), .A2(
        u5_mult_82_CARRYB_46__5_), .ZN(u5_mult_82_n6169) );
  NAND2_X1 u5_mult_82_U11288 ( .A1(u5_mult_82_ab_46__6_), .A2(
        u5_mult_82_CARRYB_45__6_), .ZN(u5_mult_82_n6166) );
  XOR2_X2 u5_mult_82_U11287 ( .A(u5_mult_82_n6165), .B(u5_mult_82_SUMB_45__7_), 
        .Z(u5_mult_82_SUMB_46__6_) );
  NOR2_X1 u5_mult_82_U11286 ( .A1(u5_mult_82_n6946), .A2(u5_mult_82_net65283), 
        .ZN(u5_mult_82_ab_47__4_) );
  NAND3_X2 u5_mult_82_U11285 ( .A1(u5_mult_82_n6159), .A2(u5_mult_82_n6160), 
        .A3(u5_mult_82_n6161), .ZN(u5_mult_82_CARRYB_13__38_) );
  NAND2_X1 u5_mult_82_U11284 ( .A1(u5_mult_82_ab_13__38_), .A2(
        u5_mult_82_CARRYB_12__38_), .ZN(u5_mult_82_n6159) );
  NAND3_X2 u5_mult_82_U11283 ( .A1(u5_mult_82_n6156), .A2(u5_mult_82_n6157), 
        .A3(u5_mult_82_n6158), .ZN(u5_mult_82_CARRYB_12__39_) );
  NAND2_X2 u5_mult_82_U11282 ( .A1(u5_mult_82_ab_12__39_), .A2(
        u5_mult_82_SUMB_11__40_), .ZN(u5_mult_82_n6157) );
  NAND2_X1 u5_mult_82_U11281 ( .A1(u5_mult_82_ab_12__39_), .A2(
        u5_mult_82_CARRYB_11__39_), .ZN(u5_mult_82_n6156) );
  XOR2_X2 u5_mult_82_U11280 ( .A(u5_mult_82_n6155), .B(u5_mult_82_SUMB_12__39_), .Z(u5_mult_82_SUMB_13__38_) );
  NAND3_X2 u5_mult_82_U11279 ( .A1(u5_mult_82_n6152), .A2(u5_mult_82_n6153), 
        .A3(u5_mult_82_n6154), .ZN(u5_mult_82_CARRYB_7__44_) );
  NAND2_X1 u5_mult_82_U11278 ( .A1(u5_mult_82_CARRYB_6__44_), .A2(
        u5_mult_82_SUMB_6__45_), .ZN(u5_mult_82_n6154) );
  NAND2_X1 u5_mult_82_U11277 ( .A1(u5_mult_82_ab_7__44_), .A2(
        u5_mult_82_SUMB_6__45_), .ZN(u5_mult_82_n6153) );
  NAND3_X2 u5_mult_82_U11276 ( .A1(u5_mult_82_n6151), .A2(u5_mult_82_n6150), 
        .A3(u5_mult_82_n6149), .ZN(u5_mult_82_CARRYB_6__45_) );
  NAND2_X2 u5_mult_82_U11275 ( .A1(u5_mult_82_SUMB_5__46_), .A2(
        u5_mult_82_ab_6__45_), .ZN(u5_mult_82_n6150) );
  NAND2_X1 u5_mult_82_U11274 ( .A1(u5_mult_82_ab_6__45_), .A2(
        u5_mult_82_CARRYB_5__45_), .ZN(u5_mult_82_n6149) );
  XOR2_X2 u5_mult_82_U11273 ( .A(u5_mult_82_n6148), .B(u5_mult_82_SUMB_6__45_), 
        .Z(u5_mult_82_SUMB_7__44_) );
  XOR2_X2 u5_mult_82_U11272 ( .A(u5_mult_82_n6147), .B(u5_mult_82_SUMB_5__46_), 
        .Z(u5_mult_82_SUMB_6__45_) );
  XOR2_X2 u5_mult_82_U11271 ( .A(u5_mult_82_ab_6__45_), .B(
        u5_mult_82_CARRYB_5__45_), .Z(u5_mult_82_n6147) );
  NAND2_X1 u5_mult_82_U11270 ( .A1(u5_mult_82_ab_25__26_), .A2(
        u5_mult_82_CARRYB_24__26_), .ZN(u5_mult_82_n6144) );
  NAND3_X2 u5_mult_82_U11269 ( .A1(u5_mult_82_n6143), .A2(u5_mult_82_n6142), 
        .A3(u5_mult_82_n6141), .ZN(u5_mult_82_CARRYB_24__27_) );
  XOR2_X2 u5_mult_82_U11268 ( .A(u5_mult_82_n6140), .B(u5_mult_82_SUMB_24__27_), .Z(u5_mult_82_SUMB_25__26_) );
  XOR2_X2 u5_mult_82_U11267 ( .A(u5_mult_82_ab_25__26_), .B(
        u5_mult_82_CARRYB_24__26_), .Z(u5_mult_82_n6140) );
  XOR2_X2 u5_mult_82_U11266 ( .A(u5_mult_82_n6139), .B(u5_mult_82_n1538), .Z(
        u5_mult_82_SUMB_24__27_) );
  NAND3_X2 u5_mult_82_U11265 ( .A1(u5_mult_82_n6135), .A2(u5_mult_82_n6136), 
        .A3(u5_mult_82_n6137), .ZN(u5_mult_82_CARRYB_47__4_) );
  NAND2_X1 u5_mult_82_U11264 ( .A1(u5_mult_82_ab_47__4_), .A2(
        u5_mult_82_CARRYB_46__4_), .ZN(u5_mult_82_n6137) );
  NAND2_X1 u5_mult_82_U11263 ( .A1(u5_mult_82_CARRYB_46__4_), .A2(
        u5_mult_82_SUMB_46__5_), .ZN(u5_mult_82_n6135) );
  XOR2_X2 u5_mult_82_U11262 ( .A(u5_mult_82_SUMB_46__5_), .B(u5_mult_82_n6134), 
        .Z(u5_mult_82_SUMB_47__4_) );
  NAND2_X2 u5_mult_82_U11261 ( .A1(u5_mult_82_ab_42__9_), .A2(
        u5_mult_82_SUMB_41__10_), .ZN(u5_mult_82_n6132) );
  NOR2_X1 u5_mult_82_U11260 ( .A1(u5_mult_82_n6843), .A2(u5_mult_82_n6663), 
        .ZN(u5_mult_82_ab_28__32_) );
  NAND3_X2 u5_mult_82_U11259 ( .A1(u5_mult_82_n6128), .A2(u5_mult_82_n6129), 
        .A3(u5_mult_82_n6130), .ZN(u5_mult_82_CARRYB_16__44_) );
  NAND2_X1 u5_mult_82_U11258 ( .A1(u5_mult_82_ab_16__44_), .A2(
        u5_mult_82_SUMB_15__45_), .ZN(u5_mult_82_n6129) );
  NAND2_X1 u5_mult_82_U11257 ( .A1(u5_mult_82_ab_16__44_), .A2(
        u5_mult_82_n5552), .ZN(u5_mult_82_n6128) );
  NAND3_X2 u5_mult_82_U11256 ( .A1(u5_mult_82_n6125), .A2(u5_mult_82_n6126), 
        .A3(u5_mult_82_n6127), .ZN(u5_mult_82_CARRYB_15__45_) );
  NAND2_X2 u5_mult_82_U11255 ( .A1(u5_mult_82_ab_15__45_), .A2(
        u5_mult_82_n1639), .ZN(u5_mult_82_n6126) );
  XOR2_X2 u5_mult_82_U11254 ( .A(u5_mult_82_n6124), .B(u5_mult_82_n1639), .Z(
        u5_mult_82_SUMB_15__45_) );
  XOR2_X2 u5_mult_82_U11253 ( .A(u5_mult_82_ab_15__45_), .B(
        u5_mult_82_CARRYB_14__45_), .Z(u5_mult_82_n6124) );
  NAND3_X2 u5_mult_82_U11252 ( .A1(u5_mult_82_n6121), .A2(u5_mult_82_n6122), 
        .A3(u5_mult_82_n6123), .ZN(u5_mult_82_CARRYB_30__30_) );
  NAND2_X1 u5_mult_82_U11251 ( .A1(u5_mult_82_CARRYB_29__30_), .A2(
        u5_mult_82_SUMB_29__31_), .ZN(u5_mult_82_n6123) );
  NAND2_X1 u5_mult_82_U11250 ( .A1(u5_mult_82_ab_30__30_), .A2(
        u5_mult_82_SUMB_29__31_), .ZN(u5_mult_82_n6122) );
  NAND3_X2 u5_mult_82_U11249 ( .A1(u5_mult_82_n6118), .A2(u5_mult_82_n6119), 
        .A3(u5_mult_82_n6120), .ZN(u5_mult_82_CARRYB_29__31_) );
  NAND2_X1 u5_mult_82_U11248 ( .A1(u5_mult_82_ab_29__31_), .A2(u5_mult_82_n349), .ZN(u5_mult_82_n6118) );
  XOR2_X2 u5_mult_82_U11247 ( .A(u5_mult_82_n6117), .B(u5_mult_82_SUMB_28__32_), .Z(u5_mult_82_SUMB_29__31_) );
  NAND3_X2 u5_mult_82_U11246 ( .A1(u5_mult_82_n6114), .A2(u5_mult_82_n6115), 
        .A3(u5_mult_82_n6116), .ZN(u5_mult_82_CARRYB_28__32_) );
  NAND2_X1 u5_mult_82_U11245 ( .A1(u5_mult_82_ab_28__32_), .A2(
        u5_mult_82_CARRYB_27__32_), .ZN(u5_mult_82_n6116) );
  NAND2_X2 u5_mult_82_U11244 ( .A1(u5_mult_82_ab_28__32_), .A2(
        u5_mult_82_n1415), .ZN(u5_mult_82_n6115) );
  NAND3_X4 u5_mult_82_U11243 ( .A1(u5_mult_82_n6111), .A2(u5_mult_82_n6112), 
        .A3(u5_mult_82_n6113), .ZN(u5_mult_82_CARRYB_49__11_) );
  NAND2_X2 u5_mult_82_U11242 ( .A1(u5_mult_82_CARRYB_48__11_), .A2(
        u5_mult_82_SUMB_48__12_), .ZN(u5_mult_82_n6113) );
  NAND2_X2 u5_mult_82_U11241 ( .A1(u5_mult_82_ab_49__11_), .A2(
        u5_mult_82_SUMB_48__12_), .ZN(u5_mult_82_n6112) );
  NAND2_X1 u5_mult_82_U11240 ( .A1(u5_mult_82_ab_48__12_), .A2(
        u5_mult_82_CARRYB_47__12_), .ZN(u5_mult_82_n6108) );
  XOR2_X2 u5_mult_82_U11239 ( .A(u5_mult_82_n6107), .B(u5_mult_82_SUMB_48__12_), .Z(u5_mult_82_SUMB_49__11_) );
  NOR2_X2 u5_mult_82_U11238 ( .A1(u5_mult_82_n6781), .A2(u5_mult_82_net66087), 
        .ZN(u5_mult_82_ab_2__48_) );
  XNOR2_X2 u5_mult_82_U11237 ( .A(u5_mult_82_CARRYB_41__10_), .B(
        u5_mult_82_ab_42__10_), .ZN(u5_mult_82_n6106) );
  XNOR2_X2 u5_mult_82_U11236 ( .A(u5_mult_82_n6106), .B(
        u5_mult_82_SUMB_41__11_), .ZN(u5_mult_82_SUMB_42__10_) );
  NOR2_X1 u5_mult_82_U11235 ( .A1(u5_mult_82_n6813), .A2(u5_mult_82_n6527), 
        .ZN(u5_mult_82_ab_7__43_) );
  NOR2_X2 u5_mult_82_U11234 ( .A1(u5_mult_82_net64433), .A2(
        u5_mult_82_net65391), .ZN(u5_mult_82_ab_41__9_) );
  NAND3_X2 u5_mult_82_U11233 ( .A1(u5_mult_82_n6103), .A2(u5_mult_82_n6104), 
        .A3(u5_mult_82_n6105), .ZN(u5_mult_82_CARRYB_9__41_) );
  NAND2_X1 u5_mult_82_U11232 ( .A1(u5_mult_82_ab_9__41_), .A2(
        u5_mult_82_CARRYB_8__41_), .ZN(u5_mult_82_n6103) );
  NAND2_X2 u5_mult_82_U11231 ( .A1(u5_mult_82_CARRYB_7__42_), .A2(
        u5_mult_82_SUMB_7__43_), .ZN(u5_mult_82_n6102) );
  NAND2_X2 u5_mult_82_U11230 ( .A1(u5_mult_82_ab_8__42_), .A2(
        u5_mult_82_SUMB_7__43_), .ZN(u5_mult_82_n6101) );
  NAND2_X1 u5_mult_82_U11229 ( .A1(u5_mult_82_ab_8__42_), .A2(
        u5_mult_82_CARRYB_7__42_), .ZN(u5_mult_82_n6100) );
  XOR2_X2 u5_mult_82_U11228 ( .A(u5_mult_82_n6099), .B(u5_mult_82_SUMB_8__42_), 
        .Z(u5_mult_82_SUMB_9__41_) );
  XOR2_X2 u5_mult_82_U11227 ( .A(u5_mult_82_ab_9__41_), .B(
        u5_mult_82_CARRYB_8__41_), .Z(u5_mult_82_n6099) );
  NAND2_X1 u5_mult_82_U11226 ( .A1(u5_mult_82_ab_7__43_), .A2(
        u5_mult_82_CARRYB_6__43_), .ZN(u5_mult_82_n6098) );
  NAND2_X2 u5_mult_82_U11225 ( .A1(u5_mult_82_ab_7__43_), .A2(
        u5_mult_82_SUMB_6__44_), .ZN(u5_mult_82_n6097) );
  NAND2_X1 u5_mult_82_U11224 ( .A1(u5_mult_82_CARRYB_6__43_), .A2(
        u5_mult_82_SUMB_6__44_), .ZN(u5_mult_82_n6096) );
  XOR2_X2 u5_mult_82_U11223 ( .A(u5_mult_82_SUMB_6__44_), .B(u5_mult_82_n6095), 
        .Z(u5_mult_82_SUMB_7__43_) );
  NAND3_X2 u5_mult_82_U11222 ( .A1(u5_mult_82_n6092), .A2(u5_mult_82_n6093), 
        .A3(u5_mult_82_n6094), .ZN(u5_mult_82_CARRYB_13__37_) );
  NAND2_X1 u5_mult_82_U11221 ( .A1(u5_mult_82_ab_13__37_), .A2(
        u5_mult_82_CARRYB_12__37_), .ZN(u5_mult_82_n6092) );
  NAND2_X1 u5_mult_82_U11220 ( .A1(u5_mult_82_ab_12__38_), .A2(
        u5_mult_82_CARRYB_11__38_), .ZN(u5_mult_82_n6089) );
  NAND3_X2 u5_mult_82_U11219 ( .A1(u5_mult_82_n2756), .A2(u5_mult_82_n6087), 
        .A3(u5_mult_82_n6088), .ZN(u5_mult_82_CARRYB_31__19_) );
  NAND2_X1 u5_mult_82_U11218 ( .A1(u5_mult_82_CARRYB_30__19_), .A2(
        u5_mult_82_SUMB_30__20_), .ZN(u5_mult_82_n6088) );
  NAND2_X1 u5_mult_82_U11217 ( .A1(u5_mult_82_ab_31__19_), .A2(
        u5_mult_82_SUMB_30__20_), .ZN(u5_mult_82_n6087) );
  NAND3_X2 u5_mult_82_U11216 ( .A1(u5_mult_82_n6084), .A2(u5_mult_82_n6085), 
        .A3(u5_mult_82_n6086), .ZN(u5_mult_82_CARRYB_30__20_) );
  NAND2_X2 u5_mult_82_U11215 ( .A1(u5_mult_82_CARRYB_29__20_), .A2(
        u5_mult_82_SUMB_29__21_), .ZN(u5_mult_82_n6086) );
  NAND2_X2 u5_mult_82_U11214 ( .A1(u5_mult_82_ab_30__20_), .A2(
        u5_mult_82_SUMB_29__21_), .ZN(u5_mult_82_n6085) );
  NAND2_X1 u5_mult_82_U11213 ( .A1(u5_mult_82_ab_30__20_), .A2(
        u5_mult_82_CARRYB_29__20_), .ZN(u5_mult_82_n6084) );
  XOR2_X2 u5_mult_82_U11212 ( .A(u5_mult_82_n6083), .B(u5_mult_82_SUMB_29__21_), .Z(u5_mult_82_SUMB_30__20_) );
  XOR2_X2 u5_mult_82_U11211 ( .A(u5_mult_82_ab_30__20_), .B(
        u5_mult_82_CARRYB_29__20_), .Z(u5_mult_82_n6083) );
  NAND3_X2 u5_mult_82_U11210 ( .A1(u5_mult_82_n6080), .A2(u5_mult_82_n6081), 
        .A3(u5_mult_82_n6082), .ZN(u5_mult_82_CARRYB_28__22_) );
  NAND2_X1 u5_mult_82_U11209 ( .A1(u5_mult_82_CARRYB_27__22_), .A2(
        u5_mult_82_SUMB_27__23_), .ZN(u5_mult_82_n6082) );
  NAND2_X1 u5_mult_82_U11208 ( .A1(u5_mult_82_ab_28__22_), .A2(
        u5_mult_82_SUMB_27__23_), .ZN(u5_mult_82_n6081) );
  NAND2_X1 u5_mult_82_U11207 ( .A1(u5_mult_82_CARRYB_27__22_), .A2(
        u5_mult_82_ab_28__22_), .ZN(u5_mult_82_n6080) );
  NAND2_X2 u5_mult_82_U11206 ( .A1(u5_mult_82_CARRYB_26__23_), .A2(
        u5_mult_82_SUMB_26__24_), .ZN(u5_mult_82_n6079) );
  NAND2_X2 u5_mult_82_U11205 ( .A1(u5_mult_82_ab_27__23_), .A2(
        u5_mult_82_SUMB_26__24_), .ZN(u5_mult_82_n6078) );
  NAND2_X1 u5_mult_82_U11204 ( .A1(u5_mult_82_ab_27__23_), .A2(
        u5_mult_82_CARRYB_26__23_), .ZN(u5_mult_82_n6077) );
  NAND3_X2 u5_mult_82_U11203 ( .A1(u5_mult_82_n6074), .A2(u5_mult_82_n6075), 
        .A3(u5_mult_82_n6076), .ZN(u5_mult_82_CARRYB_44__6_) );
  NAND2_X1 u5_mult_82_U11202 ( .A1(u5_mult_82_CARRYB_43__6_), .A2(
        u5_mult_82_SUMB_43__7_), .ZN(u5_mult_82_n6076) );
  NAND2_X1 u5_mult_82_U11201 ( .A1(u5_mult_82_ab_44__6_), .A2(
        u5_mult_82_SUMB_43__7_), .ZN(u5_mult_82_n6075) );
  NAND2_X1 u5_mult_82_U11200 ( .A1(u5_mult_82_ab_44__6_), .A2(
        u5_mult_82_CARRYB_43__6_), .ZN(u5_mult_82_n6074) );
  NAND2_X2 u5_mult_82_U11199 ( .A1(u5_mult_82_ab_43__7_), .A2(
        u5_mult_82_SUMB_42__8_), .ZN(u5_mult_82_n6072) );
  XOR2_X2 u5_mult_82_U11198 ( .A(u5_mult_82_n6070), .B(u5_mult_82_SUMB_42__8_), 
        .Z(u5_mult_82_SUMB_43__7_) );
  XOR2_X2 u5_mult_82_U11197 ( .A(u5_mult_82_ab_43__7_), .B(
        u5_mult_82_CARRYB_42__7_), .Z(u5_mult_82_n6070) );
  NAND2_X1 u5_mult_82_U11196 ( .A1(u5_mult_82_ab_41__9_), .A2(
        u5_mult_82_CARRYB_40__9_), .ZN(u5_mult_82_n6069) );
  NOR2_X1 u5_mult_82_U11195 ( .A1(u5_mult_82_n6952), .A2(u5_mult_82_net65285), 
        .ZN(u5_mult_82_ab_47__3_) );
  NOR2_X1 u5_mult_82_U11194 ( .A1(u5_mult_82_net64361), .A2(u5_mult_82_n6736), 
        .ZN(u5_mult_82_ab_44__5_) );
  NAND3_X2 u5_mult_82_U11193 ( .A1(u5_mult_82_n6064), .A2(u5_mult_82_n6065), 
        .A3(u5_mult_82_n6066), .ZN(u5_mult_82_CARRYB_47__3_) );
  NAND2_X1 u5_mult_82_U11192 ( .A1(u5_mult_82_ab_47__3_), .A2(
        u5_mult_82_CARRYB_46__3_), .ZN(u5_mult_82_n6066) );
  NAND2_X2 u5_mult_82_U11191 ( .A1(u5_mult_82_ab_47__3_), .A2(
        u5_mult_82_SUMB_46__4_), .ZN(u5_mult_82_n6065) );
  NAND2_X1 u5_mult_82_U11190 ( .A1(u5_mult_82_CARRYB_46__3_), .A2(
        u5_mult_82_SUMB_46__4_), .ZN(u5_mult_82_n6064) );
  NAND3_X2 u5_mult_82_U11189 ( .A1(u5_mult_82_n6061), .A2(u5_mult_82_n6062), 
        .A3(u5_mult_82_n6063), .ZN(u5_mult_82_CARRYB_6__43_) );
  NAND2_X1 u5_mult_82_U11188 ( .A1(u5_mult_82_ab_6__43_), .A2(
        u5_mult_82_SUMB_5__44_), .ZN(u5_mult_82_n6062) );
  NAND3_X2 u5_mult_82_U11187 ( .A1(u5_mult_82_n6058), .A2(u5_mult_82_n6059), 
        .A3(u5_mult_82_n6060), .ZN(u5_mult_82_CARRYB_5__44_) );
  NAND2_X1 u5_mult_82_U11186 ( .A1(u5_mult_82_CARRYB_4__44_), .A2(
        u5_mult_82_SUMB_4__45_), .ZN(u5_mult_82_n6060) );
  NAND2_X1 u5_mult_82_U11185 ( .A1(u5_mult_82_ab_5__44_), .A2(
        u5_mult_82_SUMB_4__45_), .ZN(u5_mult_82_n6059) );
  NAND2_X1 u5_mult_82_U11184 ( .A1(u5_mult_82_ab_5__44_), .A2(
        u5_mult_82_CARRYB_4__44_), .ZN(u5_mult_82_n6058) );
  NAND3_X2 u5_mult_82_U11183 ( .A1(u5_mult_82_n6055), .A2(u5_mult_82_n6056), 
        .A3(u5_mult_82_n6057), .ZN(u5_mult_82_CARRYB_25__24_) );
  NAND2_X1 u5_mult_82_U11182 ( .A1(u5_mult_82_CARRYB_24__24_), .A2(
        u5_mult_82_SUMB_24__25_), .ZN(u5_mult_82_n6057) );
  NAND2_X1 u5_mult_82_U11181 ( .A1(u5_mult_82_ab_25__24_), .A2(
        u5_mult_82_SUMB_24__25_), .ZN(u5_mult_82_n6056) );
  NAND2_X2 u5_mult_82_U11180 ( .A1(u5_mult_82_n70), .A2(
        u5_mult_82_CARRYB_23__25_), .ZN(u5_mult_82_n6054) );
  NAND2_X2 u5_mult_82_U11179 ( .A1(u5_mult_82_ab_24__25_), .A2(
        u5_mult_82_SUMB_23__26_), .ZN(u5_mult_82_n6053) );
  NAND2_X1 u5_mult_82_U11178 ( .A1(u5_mult_82_ab_24__25_), .A2(
        u5_mult_82_CARRYB_23__25_), .ZN(u5_mult_82_n6052) );
  XOR2_X2 u5_mult_82_U11177 ( .A(u5_mult_82_n6051), .B(u5_mult_82_SUMB_24__25_), .Z(u5_mult_82_SUMB_25__24_) );
  NAND3_X2 u5_mult_82_U11176 ( .A1(u5_mult_82_n6048), .A2(u5_mult_82_n6049), 
        .A3(u5_mult_82_n6050), .ZN(u5_mult_82_CARRYB_17__32_) );
  NAND2_X1 u5_mult_82_U11175 ( .A1(u5_mult_82_CARRYB_16__32_), .A2(
        u5_mult_82_SUMB_16__33_), .ZN(u5_mult_82_n6050) );
  NAND2_X1 u5_mult_82_U11174 ( .A1(u5_mult_82_ab_17__32_), .A2(
        u5_mult_82_SUMB_16__33_), .ZN(u5_mult_82_n6049) );
  NAND2_X1 u5_mult_82_U11173 ( .A1(u5_mult_82_ab_17__32_), .A2(
        u5_mult_82_CARRYB_16__32_), .ZN(u5_mult_82_n6048) );
  NAND2_X1 u5_mult_82_U11172 ( .A1(u5_mult_82_ab_16__33_), .A2(
        u5_mult_82_CARRYB_15__33_), .ZN(u5_mult_82_n6045) );
  XOR2_X2 u5_mult_82_U11171 ( .A(u5_mult_82_n6044), .B(u5_mult_82_SUMB_16__33_), .Z(u5_mult_82_SUMB_17__32_) );
  XOR2_X2 u5_mult_82_U11170 ( .A(u5_mult_82_n6043), .B(u5_mult_82_SUMB_15__34_), .Z(u5_mult_82_SUMB_16__33_) );
  XOR2_X2 u5_mult_82_U11169 ( .A(u5_mult_82_ab_16__33_), .B(
        u5_mult_82_CARRYB_15__33_), .Z(u5_mult_82_n6043) );
  NAND3_X2 u5_mult_82_U11168 ( .A1(u5_mult_82_n6040), .A2(u5_mult_82_n6041), 
        .A3(u5_mult_82_n6042), .ZN(u5_mult_82_CARRYB_35__14_) );
  NAND2_X1 u5_mult_82_U11167 ( .A1(u5_mult_82_SUMB_34__15_), .A2(
        u5_mult_82_CARRYB_34__14_), .ZN(u5_mult_82_n6042) );
  NAND2_X1 u5_mult_82_U11166 ( .A1(u5_mult_82_ab_35__14_), .A2(
        u5_mult_82_SUMB_34__15_), .ZN(u5_mult_82_n6041) );
  NAND2_X1 u5_mult_82_U11165 ( .A1(u5_mult_82_ab_35__14_), .A2(
        u5_mult_82_CARRYB_34__14_), .ZN(u5_mult_82_n6040) );
  NAND3_X2 u5_mult_82_U11164 ( .A1(u5_mult_82_n6037), .A2(u5_mult_82_n6038), 
        .A3(u5_mult_82_n6039), .ZN(u5_mult_82_CARRYB_34__15_) );
  NAND2_X2 u5_mult_82_U11163 ( .A1(u5_mult_82_ab_34__15_), .A2(
        u5_mult_82_SUMB_33__16_), .ZN(u5_mult_82_n6038) );
  NAND2_X2 u5_mult_82_U11162 ( .A1(u5_mult_82_ab_29__20_), .A2(
        u5_mult_82_SUMB_28__21_), .ZN(u5_mult_82_n6036) );
  NAND2_X2 u5_mult_82_U11161 ( .A1(u5_mult_82_ab_44__5_), .A2(
        u5_mult_82_SUMB_43__6_), .ZN(u5_mult_82_n6034) );
  NAND2_X1 u5_mult_82_U11160 ( .A1(u5_mult_82_ab_43__6_), .A2(
        u5_mult_82_CARRYB_42__6_), .ZN(u5_mult_82_n6030) );
  NAND2_X2 u5_mult_82_U11159 ( .A1(u5_mult_82_CARRYB_41__7_), .A2(
        u5_mult_82_SUMB_41__8_), .ZN(u5_mult_82_n6029) );
  NAND2_X2 u5_mult_82_U11158 ( .A1(u5_mult_82_ab_42__7_), .A2(
        u5_mult_82_SUMB_41__8_), .ZN(u5_mult_82_n6028) );
  INV_X8 u5_mult_82_U11157 ( .A(n4768), .ZN(u5_mult_82_n7007) );
  NOR2_X1 u5_mult_82_U11156 ( .A1(u5_mult_82_n6946), .A2(u5_mult_82_net65319), 
        .ZN(u5_mult_82_ab_45__4_) );
  NAND3_X2 u5_mult_82_U11155 ( .A1(u5_mult_82_n6025), .A2(u5_mult_82_n6024), 
        .A3(u5_mult_82_n6026), .ZN(u5_mult_82_CARRYB_45__4_) );
  NAND2_X2 u5_mult_82_U11154 ( .A1(u5_mult_82_ab_45__4_), .A2(
        u5_mult_82_SUMB_44__5_), .ZN(u5_mult_82_n6025) );
  NAND3_X2 u5_mult_82_U11153 ( .A1(u5_mult_82_n6021), .A2(u5_mult_82_n6022), 
        .A3(u5_mult_82_n6023), .ZN(u5_mult_82_CARRYB_8__40_) );
  NAND2_X1 u5_mult_82_U11152 ( .A1(u5_mult_82_ab_8__40_), .A2(
        u5_mult_82_SUMB_7__41_), .ZN(u5_mult_82_n6022) );
  NAND3_X2 u5_mult_82_U11151 ( .A1(u5_mult_82_n6015), .A2(u5_mult_82_n6016), 
        .A3(u5_mult_82_n6017), .ZN(u5_mult_82_CARRYB_19__29_) );
  NAND2_X1 u5_mult_82_U11150 ( .A1(u5_mult_82_SUMB_18__30_), .A2(
        u5_mult_82_CARRYB_18__29_), .ZN(u5_mult_82_n6017) );
  NAND2_X1 u5_mult_82_U11149 ( .A1(u5_mult_82_ab_19__29_), .A2(
        u5_mult_82_CARRYB_18__29_), .ZN(u5_mult_82_n6015) );
  NAND3_X2 u5_mult_82_U11148 ( .A1(u5_mult_82_n6012), .A2(u5_mult_82_n6013), 
        .A3(u5_mult_82_n6014), .ZN(u5_mult_82_CARRYB_18__30_) );
  NAND2_X1 u5_mult_82_U11147 ( .A1(u5_mult_82_ab_18__30_), .A2(
        u5_mult_82_CARRYB_17__30_), .ZN(u5_mult_82_n6012) );
  NAND3_X2 u5_mult_82_U11146 ( .A1(u5_mult_82_n6009), .A2(u5_mult_82_n6010), 
        .A3(u5_mult_82_n6011), .ZN(u5_mult_82_CARRYB_31__17_) );
  NAND2_X1 u5_mult_82_U11145 ( .A1(u5_mult_82_SUMB_30__18_), .A2(
        u5_mult_82_CARRYB_30__17_), .ZN(u5_mult_82_n6011) );
  NAND2_X1 u5_mult_82_U11144 ( .A1(u5_mult_82_ab_31__17_), .A2(
        u5_mult_82_SUMB_30__18_), .ZN(u5_mult_82_n6010) );
  NAND2_X1 u5_mult_82_U11143 ( .A1(u5_mult_82_ab_31__17_), .A2(
        u5_mult_82_CARRYB_30__17_), .ZN(u5_mult_82_n6009) );
  NAND2_X1 u5_mult_82_U11142 ( .A1(u5_mult_82_ab_30__18_), .A2(
        u5_mult_82_CARRYB_29__18_), .ZN(u5_mult_82_net79263) );
  NAND2_X2 u5_mult_82_U11141 ( .A1(u5_mult_82_ab_41__7_), .A2(u5_mult_82_n1752), .ZN(u5_mult_82_n6004) );
  NAND2_X1 u5_mult_82_U11140 ( .A1(u5_mult_82_ab_41__7_), .A2(
        u5_mult_82_CARRYB_40__7_), .ZN(u5_mult_82_n6003) );
  NAND3_X2 u5_mult_82_U11139 ( .A1(u5_mult_82_n6000), .A2(u5_mult_82_n6001), 
        .A3(u5_mult_82_n6002), .ZN(u5_mult_82_CARRYB_23__38_) );
  NAND2_X2 u5_mult_82_U11138 ( .A1(u5_mult_82_ab_22__39_), .A2(
        u5_mult_82_SUMB_21__40_), .ZN(u5_mult_82_n5998) );
  NAND3_X2 u5_mult_82_U11137 ( .A1(u5_mult_82_n5994), .A2(u5_mult_82_n5995), 
        .A3(u5_mult_82_n5996), .ZN(u5_mult_82_CARRYB_35__26_) );
  NAND2_X1 u5_mult_82_U11136 ( .A1(u5_mult_82_ab_35__26_), .A2(
        u5_mult_82_CARRYB_34__26_), .ZN(u5_mult_82_n5996) );
  NAND2_X2 u5_mult_82_U11135 ( .A1(u5_mult_82_ab_35__26_), .A2(
        u5_mult_82_SUMB_34__27_), .ZN(u5_mult_82_n5995) );
  NAND2_X1 u5_mult_82_U11134 ( .A1(u5_mult_82_ab_50__11_), .A2(
        u5_mult_82_CARRYB_49__11_), .ZN(u5_mult_82_n5991) );
  NAND2_X1 u5_mult_82_U11133 ( .A1(u5_mult_82_ab_49__12_), .A2(
        u5_mult_82_CARRYB_48__12_), .ZN(u5_mult_82_n5988) );
  INV_X8 u5_mult_82_U11132 ( .A(n4785), .ZN(u5_mult_82_n7008) );
  NOR2_X2 u5_mult_82_U11131 ( .A1(u5_mult_82_n6818), .A2(u5_mult_82_net66019), 
        .ZN(u5_mult_82_ab_6__42_) );
  NOR2_X1 u5_mult_82_U11130 ( .A1(u5_mult_82_n6920), .A2(u5_mult_82_n6700), 
        .ZN(u5_mult_82_ab_33__18_) );
  NAND2_X1 u5_mult_82_U11129 ( .A1(u5_mult_82_ab_6__42_), .A2(
        u5_mult_82_CARRYB_5__42_), .ZN(u5_mult_82_n5987) );
  NAND3_X2 u5_mult_82_U11128 ( .A1(u5_mult_82_n5982), .A2(u5_mult_82_n5983), 
        .A3(u5_mult_82_n5984), .ZN(u5_mult_82_CARRYB_33__18_) );
  NAND2_X1 u5_mult_82_U11127 ( .A1(u5_mult_82_ab_33__18_), .A2(
        u5_mult_82_CARRYB_32__18_), .ZN(u5_mult_82_n5984) );
  NAND2_X1 u5_mult_82_U11126 ( .A1(u5_mult_82_CARRYB_32__18_), .A2(
        u5_mult_82_SUMB_32__19_), .ZN(u5_mult_82_n5982) );
  NAND2_X1 u5_mult_82_U11125 ( .A1(u5_mult_82_ab_8__41_), .A2(
        u5_mult_82_CARRYB_7__41_), .ZN(u5_mult_82_n5979) );
  NAND2_X2 u5_mult_82_U11124 ( .A1(u5_mult_82_CARRYB_6__42_), .A2(
        u5_mult_82_SUMB_6__43_), .ZN(u5_mult_82_n5978) );
  NAND2_X2 u5_mult_82_U11123 ( .A1(u5_mult_82_ab_7__42_), .A2(
        u5_mult_82_SUMB_6__43_), .ZN(u5_mult_82_n5977) );
  XOR2_X2 u5_mult_82_U11122 ( .A(u5_mult_82_n5975), .B(u5_mult_82_SUMB_7__42_), 
        .Z(u5_mult_82_SUMB_8__41_) );
  XOR2_X2 u5_mult_82_U11121 ( .A(u5_mult_82_ab_8__41_), .B(
        u5_mult_82_CARRYB_7__41_), .Z(u5_mult_82_n5975) );
  NAND2_X1 u5_mult_82_U11120 ( .A1(u5_mult_82_ab_25__25_), .A2(
        u5_mult_82_CARRYB_24__25_), .ZN(u5_mult_82_n5972) );
  NAND2_X2 u5_mult_82_U11119 ( .A1(u5_mult_82_ab_24__26_), .A2(
        u5_mult_82_n1395), .ZN(u5_mult_82_n5970) );
  NAND2_X1 u5_mult_82_U11118 ( .A1(u5_mult_82_ab_24__26_), .A2(
        u5_mult_82_CARRYB_23__26_), .ZN(u5_mult_82_n5969) );
  NAND3_X2 u5_mult_82_U11117 ( .A1(u5_mult_82_n5965), .A2(u5_mult_82_n5967), 
        .A3(u5_mult_82_n5966), .ZN(u5_mult_82_CARRYB_37__17_) );
  NAND2_X1 u5_mult_82_U11116 ( .A1(u5_mult_82_ab_37__17_), .A2(
        u5_mult_82_CARRYB_36__17_), .ZN(u5_mult_82_n5965) );
  NAND2_X2 u5_mult_82_U11115 ( .A1(u5_mult_82_CARRYB_35__18_), .A2(
        u5_mult_82_SUMB_35__19_), .ZN(u5_mult_82_n5964) );
  NAND2_X2 u5_mult_82_U11114 ( .A1(u5_mult_82_ab_36__18_), .A2(
        u5_mult_82_SUMB_35__19_), .ZN(u5_mult_82_n5963) );
  NAND2_X1 u5_mult_82_U11113 ( .A1(u5_mult_82_ab_44__10_), .A2(
        u5_mult_82_CARRYB_43__10_), .ZN(u5_mult_82_n5961) );
  XNOR2_X2 u5_mult_82_U11112 ( .A(u5_mult_82_ab_47__5_), .B(
        u5_mult_82_CARRYB_46__5_), .ZN(u5_mult_82_n5960) );
  XNOR2_X2 u5_mult_82_U11111 ( .A(u5_mult_82_SUMB_41__10_), .B(
        u5_mult_82_n5959), .ZN(u5_mult_82_SUMB_42__9_) );
  NOR2_X1 u5_mult_82_U11110 ( .A1(u5_mult_82_n6843), .A2(u5_mult_82_n6693), 
        .ZN(u5_mult_82_ab_32__32_) );
  NAND3_X2 u5_mult_82_U11109 ( .A1(u5_mult_82_n5956), .A2(u5_mult_82_n5957), 
        .A3(u5_mult_82_n5958), .ZN(u5_mult_82_CARRYB_18__46_) );
  NAND2_X2 u5_mult_82_U11108 ( .A1(u5_mult_82_ab_17__47_), .A2(
        u5_mult_82_SUMB_16__48_), .ZN(u5_mult_82_n5954) );
  XOR2_X2 u5_mult_82_U11107 ( .A(u5_mult_82_n5952), .B(u5_mult_82_SUMB_16__48_), .Z(u5_mult_82_SUMB_17__47_) );
  XOR2_X2 u5_mult_82_U11106 ( .A(u5_mult_82_ab_17__47_), .B(u5_mult_82_n1711), 
        .Z(u5_mult_82_n5952) );
  NAND2_X1 u5_mult_82_U11105 ( .A1(u5_mult_82_ab_34__30_), .A2(
        u5_mult_82_n3825), .ZN(u5_mult_82_n5949) );
  NAND3_X2 u5_mult_82_U11104 ( .A1(u5_mult_82_n5942), .A2(u5_mult_82_n5943), 
        .A3(u5_mult_82_n5944), .ZN(u5_mult_82_CARRYB_32__32_) );
  NAND2_X2 u5_mult_82_U11103 ( .A1(u5_mult_82_ab_32__32_), .A2(
        u5_mult_82_SUMB_31__33_), .ZN(u5_mult_82_n5943) );
  NAND2_X1 u5_mult_82_U11102 ( .A1(u5_mult_82_CARRYB_31__32_), .A2(
        u5_mult_82_SUMB_31__33_), .ZN(u5_mult_82_n5942) );
  NAND3_X2 u5_mult_82_U11101 ( .A1(u5_mult_82_n5939), .A2(u5_mult_82_n5940), 
        .A3(u5_mult_82_n5941), .ZN(u5_mult_82_CARRYB_50__14_) );
  NAND2_X1 u5_mult_82_U11100 ( .A1(u5_mult_82_ab_50__14_), .A2(
        u5_mult_82_SUMB_49__15_), .ZN(u5_mult_82_n5940) );
  NAND2_X1 u5_mult_82_U11099 ( .A1(u5_mult_82_ab_50__14_), .A2(
        u5_mult_82_CARRYB_49__14_), .ZN(u5_mult_82_n5939) );
  NAND2_X2 u5_mult_82_U11098 ( .A1(u5_mult_82_CARRYB_48__15_), .A2(
        u5_mult_82_SUMB_48__16_), .ZN(u5_mult_82_n5938) );
  NAND2_X2 u5_mult_82_U11097 ( .A1(u5_mult_82_ab_49__15_), .A2(
        u5_mult_82_SUMB_48__16_), .ZN(u5_mult_82_n5937) );
  NAND2_X1 u5_mult_82_U11096 ( .A1(u5_mult_82_ab_49__15_), .A2(
        u5_mult_82_CARRYB_48__15_), .ZN(u5_mult_82_n5936) );
  XOR2_X2 u5_mult_82_U11095 ( .A(u5_mult_82_ab_25__24_), .B(
        u5_mult_82_CARRYB_24__24_), .Z(u5_mult_82_n6051) );
  NAND2_X1 u5_mult_82_U11094 ( .A1(u5_mult_82_ab_43__8_), .A2(
        u5_mult_82_SUMB_42__9_), .ZN(u5_mult_82_n5935) );
  NAND2_X2 u5_mult_82_U11093 ( .A1(u5_mult_82_ab_43__8_), .A2(
        u5_mult_82_CARRYB_42__8_), .ZN(u5_mult_82_n5934) );
  NAND2_X1 u5_mult_82_U11092 ( .A1(u5_mult_82_ab_47__6_), .A2(
        u5_mult_82_CARRYB_46__6_), .ZN(u5_mult_82_n5932) );
  NAND2_X2 u5_mult_82_U11091 ( .A1(u5_mult_82_ab_47__6_), .A2(
        u5_mult_82_SUMB_46__7_), .ZN(u5_mult_82_n5931) );
  NAND3_X2 u5_mult_82_U11090 ( .A1(u5_mult_82_n5927), .A2(u5_mult_82_n5928), 
        .A3(u5_mult_82_n5929), .ZN(u5_mult_82_CARRYB_21__26_) );
  NAND2_X1 u5_mult_82_U11089 ( .A1(u5_mult_82_CARRYB_20__26_), .A2(
        u5_mult_82_SUMB_20__27_), .ZN(u5_mult_82_n5929) );
  NAND2_X1 u5_mult_82_U11088 ( .A1(u5_mult_82_ab_21__26_), .A2(
        u5_mult_82_SUMB_20__27_), .ZN(u5_mult_82_n5928) );
  NAND2_X1 u5_mult_82_U11087 ( .A1(u5_mult_82_ab_21__26_), .A2(
        u5_mult_82_CARRYB_20__26_), .ZN(u5_mult_82_n5927) );
  NAND3_X2 u5_mult_82_U11086 ( .A1(u5_mult_82_n5924), .A2(u5_mult_82_n5925), 
        .A3(u5_mult_82_n5926), .ZN(u5_mult_82_CARRYB_20__27_) );
  NAND2_X1 u5_mult_82_U11085 ( .A1(u5_mult_82_ab_20__27_), .A2(
        u5_mult_82_CARRYB_19__27_), .ZN(u5_mult_82_n5924) );
  NAND3_X2 u5_mult_82_U11084 ( .A1(u5_mult_82_n5920), .A2(u5_mult_82_n5919), 
        .A3(u5_mult_82_n5918), .ZN(u5_mult_82_CARRYB_33__14_) );
  XOR2_X2 u5_mult_82_U11083 ( .A(u5_mult_82_n5917), .B(u5_mult_82_SUMB_33__14_), .Z(u5_mult_82_SUMB_34__13_) );
  XOR2_X2 u5_mult_82_U11082 ( .A(u5_mult_82_ab_34__13_), .B(
        u5_mult_82_CARRYB_33__13_), .Z(u5_mult_82_n5917) );
  NOR2_X1 u5_mult_82_U11081 ( .A1(u5_mult_82_net64469), .A2(u5_mult_82_n6736), 
        .ZN(u5_mult_82_ab_44__11_) );
  NOR2_X1 u5_mult_82_U11080 ( .A1(u5_mult_82_net64959), .A2(u5_mult_82_n6544), 
        .ZN(u5_mult_82_ab_9__38_) );
  NAND3_X2 u5_mult_82_U11079 ( .A1(u5_mult_82_n5914), .A2(u5_mult_82_n5915), 
        .A3(u5_mult_82_n5916), .ZN(u5_mult_82_CARRYB_17__31_) );
  NAND2_X2 u5_mult_82_U11078 ( .A1(u5_mult_82_ab_17__31_), .A2(
        u5_mult_82_CARRYB_16__31_), .ZN(u5_mult_82_n5915) );
  NAND3_X2 u5_mult_82_U11077 ( .A1(u5_mult_82_n5911), .A2(u5_mult_82_n5912), 
        .A3(u5_mult_82_n5913), .ZN(u5_mult_82_CARRYB_16__31_) );
  NAND2_X1 u5_mult_82_U11076 ( .A1(u5_mult_82_CARRYB_15__31_), .A2(
        u5_mult_82_SUMB_15__32_), .ZN(u5_mult_82_n5913) );
  NAND2_X2 u5_mult_82_U11075 ( .A1(u5_mult_82_ab_16__31_), .A2(
        u5_mult_82_SUMB_15__32_), .ZN(u5_mult_82_n5912) );
  NAND3_X2 u5_mult_82_U11074 ( .A1(u5_mult_82_net79444), .A2(u5_mult_82_n5910), 
        .A3(u5_mult_82_net79446), .ZN(u5_mult_82_CARRYB_44__11_) );
  NAND2_X2 u5_mult_82_U11073 ( .A1(u5_mult_82_ab_44__11_), .A2(
        u5_mult_82_SUMB_43__12_), .ZN(u5_mult_82_n5910) );
  NAND3_X2 u5_mult_82_U11072 ( .A1(u5_mult_82_n5907), .A2(u5_mult_82_n5908), 
        .A3(u5_mult_82_n5909), .ZN(u5_mult_82_CARRYB_11__36_) );
  NAND2_X1 u5_mult_82_U11071 ( .A1(u5_mult_82_CARRYB_10__36_), .A2(
        u5_mult_82_SUMB_10__37_), .ZN(u5_mult_82_n5909) );
  NAND2_X1 u5_mult_82_U11070 ( .A1(u5_mult_82_ab_11__36_), .A2(
        u5_mult_82_SUMB_10__37_), .ZN(u5_mult_82_n5908) );
  NAND2_X1 u5_mult_82_U11069 ( .A1(u5_mult_82_ab_11__36_), .A2(
        u5_mult_82_CARRYB_10__36_), .ZN(u5_mult_82_n5907) );
  NAND2_X2 u5_mult_82_U11068 ( .A1(u5_mult_82_ab_10__37_), .A2(
        u5_mult_82_SUMB_9__38_), .ZN(u5_mult_82_n5905) );
  NAND2_X1 u5_mult_82_U11067 ( .A1(u5_mult_82_ab_10__37_), .A2(
        u5_mult_82_CARRYB_9__37_), .ZN(u5_mult_82_n5904) );
  XOR2_X2 u5_mult_82_U11066 ( .A(u5_mult_82_n5903), .B(u5_mult_82_SUMB_10__37_), .Z(u5_mult_82_SUMB_11__36_) );
  XOR2_X2 u5_mult_82_U11065 ( .A(u5_mult_82_n5902), .B(u5_mult_82_SUMB_9__38_), 
        .Z(u5_mult_82_SUMB_10__37_) );
  NAND2_X1 u5_mult_82_U11064 ( .A1(u5_mult_82_ab_9__38_), .A2(
        u5_mult_82_CARRYB_8__38_), .ZN(u5_mult_82_n5901) );
  NAND2_X2 u5_mult_82_U11063 ( .A1(u5_mult_82_ab_9__38_), .A2(u5_mult_82_n1452), .ZN(u5_mult_82_n5900) );
  NAND2_X1 u5_mult_82_U11062 ( .A1(u5_mult_82_CARRYB_34__20_), .A2(
        u5_mult_82_SUMB_34__21_), .ZN(u5_mult_82_n5898) );
  NAND2_X1 u5_mult_82_U11061 ( .A1(u5_mult_82_ab_35__20_), .A2(
        u5_mult_82_SUMB_34__21_), .ZN(u5_mult_82_n5897) );
  NAND2_X1 u5_mult_82_U11060 ( .A1(u5_mult_82_ab_35__20_), .A2(
        u5_mult_82_CARRYB_34__20_), .ZN(u5_mult_82_n5896) );
  NAND2_X1 u5_mult_82_U11059 ( .A1(u5_mult_82_ab_34__21_), .A2(
        u5_mult_82_SUMB_33__22_), .ZN(u5_mult_82_n5894) );
  NAND2_X1 u5_mult_82_U11058 ( .A1(u5_mult_82_ab_34__21_), .A2(
        u5_mult_82_CARRYB_33__21_), .ZN(u5_mult_82_n5893) );
  XOR2_X2 u5_mult_82_U11057 ( .A(u5_mult_82_n5892), .B(u5_mult_82_SUMB_34__21_), .Z(u5_mult_82_SUMB_35__20_) );
  XOR2_X2 u5_mult_82_U11056 ( .A(u5_mult_82_n5891), .B(u5_mult_82_SUMB_33__22_), .Z(u5_mult_82_SUMB_34__21_) );
  NAND3_X2 u5_mult_82_U11055 ( .A1(u5_mult_82_n5888), .A2(u5_mult_82_n5889), 
        .A3(u5_mult_82_n5890), .ZN(u5_mult_82_CARRYB_22__37_) );
  NAND2_X1 u5_mult_82_U11054 ( .A1(u5_mult_82_CARRYB_21__37_), .A2(
        u5_mult_82_SUMB_21__38_), .ZN(u5_mult_82_n5890) );
  NAND2_X1 u5_mult_82_U11053 ( .A1(u5_mult_82_ab_22__37_), .A2(
        u5_mult_82_SUMB_21__38_), .ZN(u5_mult_82_n5889) );
  NAND2_X1 u5_mult_82_U11052 ( .A1(u5_mult_82_ab_22__37_), .A2(
        u5_mult_82_CARRYB_21__37_), .ZN(u5_mult_82_n5888) );
  NAND3_X2 u5_mult_82_U11051 ( .A1(u5_mult_82_n5885), .A2(u5_mult_82_n5886), 
        .A3(u5_mult_82_n5887), .ZN(u5_mult_82_CARRYB_21__38_) );
  NAND2_X2 u5_mult_82_U11050 ( .A1(u5_mult_82_CARRYB_20__38_), .A2(
        u5_mult_82_n1788), .ZN(u5_mult_82_n5887) );
  NAND2_X2 u5_mult_82_U11049 ( .A1(u5_mult_82_ab_21__38_), .A2(
        u5_mult_82_n1788), .ZN(u5_mult_82_n5886) );
  NAND2_X1 u5_mult_82_U11048 ( .A1(u5_mult_82_ab_21__38_), .A2(
        u5_mult_82_CARRYB_20__38_), .ZN(u5_mult_82_n5885) );
  XOR2_X2 u5_mult_82_U11047 ( .A(u5_mult_82_n5884), .B(u5_mult_82_n1788), .Z(
        u5_mult_82_SUMB_21__38_) );
  XOR2_X2 u5_mult_82_U11046 ( .A(u5_mult_82_ab_21__38_), .B(
        u5_mult_82_CARRYB_20__38_), .Z(u5_mult_82_n5884) );
  NAND3_X2 u5_mult_82_U11045 ( .A1(u5_mult_82_n5881), .A2(u5_mult_82_n5882), 
        .A3(u5_mult_82_n5883), .ZN(u5_mult_82_CARRYB_43__16_) );
  NAND2_X1 u5_mult_82_U11044 ( .A1(u5_mult_82_ab_43__16_), .A2(
        u5_mult_82_SUMB_42__17_), .ZN(u5_mult_82_n5882) );
  NAND2_X1 u5_mult_82_U11043 ( .A1(u5_mult_82_n1837), .A2(
        u5_mult_82_SUMB_42__17_), .ZN(u5_mult_82_n5881) );
  XOR2_X2 u5_mult_82_U11042 ( .A(u5_mult_82_SUMB_42__17_), .B(u5_mult_82_n5880), .Z(u5_mult_82_SUMB_43__16_) );
  NOR2_X1 u5_mult_82_U11041 ( .A1(u5_mult_82_n6805), .A2(u5_mult_82_n6615), 
        .ZN(u5_mult_82_ab_19__44_) );
  NOR2_X1 u5_mult_82_U11040 ( .A1(u5_mult_82_n6798), .A2(u5_mult_82_n6607), 
        .ZN(u5_mult_82_ab_18__45_) );
  NOR2_X1 u5_mult_82_U11039 ( .A1(u5_mult_82_n6919), .A2(u5_mult_82_net65321), 
        .ZN(u5_mult_82_ab_45__18_) );
  NAND3_X2 u5_mult_82_U11038 ( .A1(u5_mult_82_n5877), .A2(u5_mult_82_n5878), 
        .A3(u5_mult_82_n5879), .ZN(u5_mult_82_CARRYB_19__44_) );
  NAND3_X2 u5_mult_82_U11037 ( .A1(u5_mult_82_n5874), .A2(u5_mult_82_n5875), 
        .A3(u5_mult_82_n5876), .ZN(u5_mult_82_CARRYB_18__45_) );
  NAND2_X2 u5_mult_82_U11036 ( .A1(u5_mult_82_n1800), .A2(
        u5_mult_82_ab_32__31_), .ZN(u5_mult_82_n5869) );
  NAND2_X1 u5_mult_82_U11035 ( .A1(u5_mult_82_ab_32__31_), .A2(
        u5_mult_82_CARRYB_31__31_), .ZN(u5_mult_82_n5868) );
  NAND3_X2 u5_mult_82_U11034 ( .A1(u5_mult_82_n5864), .A2(u5_mult_82_n5865), 
        .A3(u5_mult_82_n5866), .ZN(u5_mult_82_CARRYB_47__16_) );
  NAND2_X1 u5_mult_82_U11033 ( .A1(u5_mult_82_CARRYB_46__16_), .A2(
        u5_mult_82_SUMB_46__17_), .ZN(u5_mult_82_n5866) );
  NAND2_X1 u5_mult_82_U11032 ( .A1(u5_mult_82_ab_47__16_), .A2(
        u5_mult_82_SUMB_46__17_), .ZN(u5_mult_82_n5865) );
  NAND2_X2 u5_mult_82_U11031 ( .A1(u5_mult_82_ab_46__17_), .A2(
        u5_mult_82_SUMB_45__18_), .ZN(u5_mult_82_n5862) );
  NAND2_X2 u5_mult_82_U11030 ( .A1(u5_mult_82_ab_45__18_), .A2(
        u5_mult_82_SUMB_44__19_), .ZN(u5_mult_82_n5858) );
  NOR2_X1 u5_mult_82_U11029 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6642), 
        .ZN(u5_mult_82_ab_24__38_) );
  NAND2_X2 u5_mult_82_U11028 ( .A1(u5_mult_82_ab_33__30_), .A2(
        u5_mult_82_CARRYB_32__30_), .ZN(u5_mult_82_n5871) );
  NOR2_X2 u5_mult_82_U11027 ( .A1(u5_mult_82_n6857), .A2(u5_mult_82_n6693), 
        .ZN(u5_mult_82_ab_32__30_) );
  NAND2_X2 u5_mult_82_U11026 ( .A1(u5_mult_82_ab_48__15_), .A2(
        u5_mult_82_CARRYB_47__15_), .ZN(u5_mult_82_n5854) );
  NAND3_X2 u5_mult_82_U11025 ( .A1(u5_mult_82_n5849), .A2(u5_mult_82_n5850), 
        .A3(u5_mult_82_n5851), .ZN(u5_mult_82_CARRYB_47__15_) );
  NAND2_X2 u5_mult_82_U11024 ( .A1(u5_mult_82_ab_47__15_), .A2(
        u5_mult_82_SUMB_46__16_), .ZN(u5_mult_82_n5850) );
  NAND2_X1 u5_mult_82_U11023 ( .A1(u5_mult_82_ab_47__15_), .A2(
        u5_mult_82_CARRYB_46__15_), .ZN(u5_mult_82_n5849) );
  NAND2_X2 u5_mult_82_U11022 ( .A1(u5_mult_82_ab_24__38_), .A2(
        u5_mult_82_SUMB_23__39_), .ZN(u5_mult_82_n5847) );
  NAND3_X2 u5_mult_82_U11021 ( .A1(u5_mult_82_n5843), .A2(u5_mult_82_n5844), 
        .A3(u5_mult_82_n5845), .ZN(u5_mult_82_CARRYB_20__42_) );
  NAND2_X1 u5_mult_82_U11020 ( .A1(u5_mult_82_ab_20__42_), .A2(
        u5_mult_82_CARRYB_19__42_), .ZN(u5_mult_82_n5843) );
  NAND2_X1 u5_mult_82_U11019 ( .A1(u5_mult_82_ab_19__43_), .A2(
        u5_mult_82_CARRYB_18__43_), .ZN(u5_mult_82_n5840) );
  NAND3_X2 u5_mult_82_U11018 ( .A1(u5_mult_82_n5837), .A2(u5_mult_82_n5838), 
        .A3(u5_mult_82_n5839), .ZN(u5_mult_82_CARRYB_44__18_) );
  NAND2_X1 u5_mult_82_U11017 ( .A1(u5_mult_82_ab_44__18_), .A2(
        u5_mult_82_CARRYB_43__18_), .ZN(u5_mult_82_n5837) );
  NAND3_X2 u5_mult_82_U11016 ( .A1(u5_mult_82_n5834), .A2(u5_mult_82_n5835), 
        .A3(u5_mult_82_n5836), .ZN(u5_mult_82_CARRYB_43__19_) );
  NAND2_X1 u5_mult_82_U11015 ( .A1(u5_mult_82_CARRYB_42__19_), .A2(
        u5_mult_82_SUMB_42__20_), .ZN(u5_mult_82_n5836) );
  NAND2_X1 u5_mult_82_U11014 ( .A1(u5_mult_82_ab_43__19_), .A2(
        u5_mult_82_SUMB_42__20_), .ZN(u5_mult_82_n5835) );
  NAND2_X1 u5_mult_82_U11013 ( .A1(u5_mult_82_ab_43__19_), .A2(
        u5_mult_82_CARRYB_42__19_), .ZN(u5_mult_82_n5834) );
  XOR2_X2 u5_mult_82_U11012 ( .A(u5_mult_82_n5833), .B(u5_mult_82_SUMB_42__20_), .Z(u5_mult_82_SUMB_43__19_) );
  NAND2_X1 u5_mult_82_U11011 ( .A1(u5_mult_82_ab_32__30_), .A2(
        u5_mult_82_SUMB_31__31_), .ZN(u5_mult_82_n5831) );
  NAND2_X1 u5_mult_82_U11010 ( .A1(u5_mult_82_CARRYB_31__30_), .A2(
        u5_mult_82_SUMB_31__31_), .ZN(u5_mult_82_n5830) );
  NAND3_X2 u5_mult_82_U11009 ( .A1(u5_mult_82_n5827), .A2(u5_mult_82_n5828), 
        .A3(u5_mult_82_n5829), .ZN(u5_mult_82_CARRYB_50__13_) );
  NAND2_X1 u5_mult_82_U11008 ( .A1(u5_mult_82_n2112), .A2(
        u5_mult_82_ab_50__13_), .ZN(u5_mult_82_n5827) );
  NAND2_X2 u5_mult_82_U11007 ( .A1(u5_mult_82_ab_49__14_), .A2(
        u5_mult_82_n1661), .ZN(u5_mult_82_n5825) );
  NAND2_X1 u5_mult_82_U11006 ( .A1(u5_mult_82_ab_49__14_), .A2(
        u5_mult_82_CARRYB_48__14_), .ZN(u5_mult_82_n5824) );
  NOR2_X2 u5_mult_82_U11005 ( .A1(u5_mult_82_net64379), .A2(
        u5_mult_82_net65391), .ZN(u5_mult_82_ab_41__6_) );
  NOR2_X1 u5_mult_82_U11004 ( .A1(u5_mult_82_net64381), .A2(
        u5_mult_82_net65409), .ZN(u5_mult_82_ab_40__6_) );
  NAND2_X2 u5_mult_82_U11003 ( .A1(u5_mult_82_ab_16__31_), .A2(
        u5_mult_82_CARRYB_15__31_), .ZN(u5_mult_82_n5911) );
  NAND2_X1 u5_mult_82_U11002 ( .A1(u5_mult_82_ab_41__6_), .A2(
        u5_mult_82_CARRYB_40__6_), .ZN(u5_mult_82_n5823) );
  XOR2_X2 u5_mult_82_U11001 ( .A(u5_mult_82_n1755), .B(u5_mult_82_n5820), .Z(
        u5_mult_82_SUMB_41__6_) );
  NAND3_X2 u5_mult_82_U11000 ( .A1(u5_mult_82_n5817), .A2(u5_mult_82_n5818), 
        .A3(u5_mult_82_n5819), .ZN(u5_mult_82_CARRYB_40__6_) );
  NAND2_X2 u5_mult_82_U10999 ( .A1(u5_mult_82_ab_40__6_), .A2(
        u5_mult_82_SUMB_39__7_), .ZN(u5_mult_82_n5818) );
  NAND3_X2 u5_mult_82_U10998 ( .A1(u5_mult_82_n5816), .A2(u5_mult_82_n5815), 
        .A3(u5_mult_82_n5814), .ZN(u5_mult_82_CARRYB_48__1_) );
  NAND2_X2 u5_mult_82_U10997 ( .A1(u5_mult_82_CARRYB_47__1_), .A2(
        u5_mult_82_ab_48__1_), .ZN(u5_mult_82_n5815) );
  NAND3_X2 u5_mult_82_U10996 ( .A1(u5_mult_82_n5810), .A2(u5_mult_82_n5811), 
        .A3(u5_mult_82_n5812), .ZN(u5_mult_82_CARRYB_47__1_) );
  NAND2_X2 u5_mult_82_U10995 ( .A1(u5_mult_82_ab_47__1_), .A2(
        u5_mult_82_SUMB_46__2_), .ZN(u5_mult_82_n5811) );
  NAND3_X2 u5_mult_82_U10994 ( .A1(u5_mult_82_n5807), .A2(u5_mult_82_n5808), 
        .A3(u5_mult_82_n5809), .ZN(u5_mult_82_CARRYB_8__38_) );
  NAND2_X1 u5_mult_82_U10993 ( .A1(u5_mult_82_CARRYB_7__38_), .A2(
        u5_mult_82_SUMB_7__39_), .ZN(u5_mult_82_n5809) );
  NAND2_X1 u5_mult_82_U10992 ( .A1(u5_mult_82_ab_8__38_), .A2(
        u5_mult_82_SUMB_7__39_), .ZN(u5_mult_82_n5808) );
  NAND2_X1 u5_mult_82_U10991 ( .A1(u5_mult_82_ab_8__38_), .A2(
        u5_mult_82_CARRYB_7__38_), .ZN(u5_mult_82_n5807) );
  NAND3_X2 u5_mult_82_U10990 ( .A1(u5_mult_82_n5804), .A2(u5_mult_82_n5805), 
        .A3(u5_mult_82_n5806), .ZN(u5_mult_82_CARRYB_7__39_) );
  NAND2_X1 u5_mult_82_U10989 ( .A1(u5_mult_82_ab_7__39_), .A2(u5_mult_82_n1592), .ZN(u5_mult_82_n5805) );
  NAND2_X1 u5_mult_82_U10988 ( .A1(u5_mult_82_ab_7__39_), .A2(
        u5_mult_82_CARRYB_6__39_), .ZN(u5_mult_82_n5804) );
  XOR2_X2 u5_mult_82_U10987 ( .A(u5_mult_82_n5803), .B(u5_mult_82_SUMB_7__39_), 
        .Z(u5_mult_82_SUMB_8__38_) );
  XOR2_X2 u5_mult_82_U10986 ( .A(u5_mult_82_ab_8__38_), .B(
        u5_mult_82_CARRYB_7__38_), .Z(u5_mult_82_n5803) );
  NAND3_X2 u5_mult_82_U10985 ( .A1(u5_mult_82_n5800), .A2(u5_mult_82_n5801), 
        .A3(u5_mult_82_n5802), .ZN(u5_mult_82_CARRYB_19__27_) );
  NAND2_X1 u5_mult_82_U10984 ( .A1(u5_mult_82_ab_19__27_), .A2(
        u5_mult_82_CARRYB_18__27_), .ZN(u5_mult_82_n5800) );
  NAND3_X2 u5_mult_82_U10983 ( .A1(u5_mult_82_n5799), .A2(u5_mult_82_n5798), 
        .A3(u5_mult_82_n5797), .ZN(u5_mult_82_CARRYB_18__28_) );
  NAND2_X1 u5_mult_82_U10982 ( .A1(u5_mult_82_CARRYB_17__28_), .A2(
        u5_mult_82_n31), .ZN(u5_mult_82_n5799) );
  NAND2_X1 u5_mult_82_U10981 ( .A1(u5_mult_82_ab_18__28_), .A2(
        u5_mult_82_CARRYB_17__28_), .ZN(u5_mult_82_n5797) );
  NAND2_X2 u5_mult_82_U10980 ( .A1(u5_mult_82_ab_15__31_), .A2(
        u5_mult_82_SUMB_14__32_), .ZN(u5_mult_82_n5795) );
  NAND3_X4 u5_mult_82_U10979 ( .A1(u5_mult_82_n5788), .A2(u5_mult_82_n5789), 
        .A3(u5_mult_82_n5790), .ZN(u5_mult_82_CARRYB_44__4_) );
  XOR2_X2 u5_mult_82_U10978 ( .A(u5_mult_82_n6298), .B(u5_mult_82_SUMB_30__23_), .Z(u5_mult_82_SUMB_31__22_) );
  NOR2_X1 u5_mult_82_U10977 ( .A1(u5_mult_82_net64939), .A2(u5_mult_82_n6621), 
        .ZN(u5_mult_82_ab_20__37_) );
  NOR2_X1 u5_mult_82_U10976 ( .A1(u5_mult_82_n6813), .A2(u5_mult_82_n6564), 
        .ZN(u5_mult_82_ab_12__43_) );
  NOR2_X2 u5_mult_82_U10975 ( .A1(u5_mult_82_net64523), .A2(u5_mult_82_n6742), 
        .ZN(u5_mult_82_ab_46__14_) );
  NAND2_X1 u5_mult_82_U10974 ( .A1(u5_mult_82_ab_20__37_), .A2(
        u5_mult_82_CARRYB_19__37_), .ZN(u5_mult_82_n5786) );
  NAND2_X2 u5_mult_82_U10973 ( .A1(u5_mult_82_ab_20__37_), .A2(
        u5_mult_82_SUMB_19__38_), .ZN(u5_mult_82_n5785) );
  NAND2_X1 u5_mult_82_U10972 ( .A1(u5_mult_82_CARRYB_19__37_), .A2(
        u5_mult_82_SUMB_19__38_), .ZN(u5_mult_82_n5784) );
  NAND3_X2 u5_mult_82_U10971 ( .A1(u5_mult_82_n5780), .A2(u5_mult_82_n5781), 
        .A3(u5_mult_82_n5782), .ZN(u5_mult_82_CARRYB_12__43_) );
  NAND2_X1 u5_mult_82_U10970 ( .A1(u5_mult_82_ab_12__43_), .A2(
        u5_mult_82_CARRYB_11__43_), .ZN(u5_mult_82_n5782) );
  XOR2_X2 u5_mult_82_U10969 ( .A(u5_mult_82_SUMB_11__44_), .B(u5_mult_82_n5779), .Z(u5_mult_82_SUMB_12__43_) );
  XOR2_X2 u5_mult_82_U10968 ( .A(u5_mult_82_CARRYB_11__43_), .B(
        u5_mult_82_ab_12__43_), .Z(u5_mult_82_n5779) );
  NAND3_X2 u5_mult_82_U10967 ( .A1(u5_mult_82_n5773), .A2(u5_mult_82_n5774), 
        .A3(u5_mult_82_n5775), .ZN(u5_mult_82_CARRYB_48__14_) );
  NAND2_X2 u5_mult_82_U10966 ( .A1(u5_mult_82_ab_48__14_), .A2(
        u5_mult_82_CARRYB_47__14_), .ZN(u5_mult_82_n5774) );
  NAND2_X1 u5_mult_82_U10965 ( .A1(u5_mult_82_ab_26__33_), .A2(
        u5_mult_82_n4553), .ZN(u5_mult_82_n5767) );
  XOR2_X2 u5_mult_82_U10964 ( .A(u5_mult_82_n5763), .B(u5_mult_82_SUMB_25__34_), .Z(u5_mult_82_SUMB_26__33_) );
  XOR2_X2 u5_mult_82_U10963 ( .A(u5_mult_82_ab_26__33_), .B(u5_mult_82_n4553), 
        .Z(u5_mult_82_n5763) );
  NAND2_X1 u5_mult_82_U10962 ( .A1(u5_mult_82_SUMB_49__13_), .A2(
        u5_mult_82_CARRYB_49__12_), .ZN(u5_mult_82_n5761) );
  NAND2_X1 u5_mult_82_U10961 ( .A1(u5_mult_82_ab_50__12_), .A2(
        u5_mult_82_SUMB_49__13_), .ZN(u5_mult_82_n5760) );
  NAND2_X1 u5_mult_82_U10960 ( .A1(u5_mult_82_CARRYB_49__12_), .A2(
        u5_mult_82_ab_50__12_), .ZN(u5_mult_82_n5759) );
  NAND2_X2 u5_mult_82_U10959 ( .A1(u5_mult_82_n1388), .A2(
        u5_mult_82_SUMB_48__14_), .ZN(u5_mult_82_n5758) );
  NAND2_X2 u5_mult_82_U10958 ( .A1(u5_mult_82_ab_49__13_), .A2(
        u5_mult_82_SUMB_48__14_), .ZN(u5_mult_82_n5757) );
  NAND2_X1 u5_mult_82_U10957 ( .A1(u5_mult_82_ab_49__13_), .A2(
        u5_mult_82_CARRYB_48__13_), .ZN(u5_mult_82_n5756) );
  XOR2_X2 u5_mult_82_U10956 ( .A(u5_mult_82_n5755), .B(u5_mult_82_SUMB_48__14_), .Z(u5_mult_82_SUMB_49__13_) );
  NAND3_X4 u5_mult_82_U10955 ( .A1(u5_mult_82_n5969), .A2(u5_mult_82_n5970), 
        .A3(u5_mult_82_n5971), .ZN(u5_mult_82_CARRYB_24__26_) );
  NOR2_X1 u5_mult_82_U10954 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6693), 
        .ZN(u5_mult_82_ab_32__36_) );
  NOR2_X1 u5_mult_82_U10953 ( .A1(u5_mult_82_n6919), .A2(u5_mult_82_net65229), 
        .ZN(u5_mult_82_ab_50__18_) );
  NAND3_X2 u5_mult_82_U10952 ( .A1(u5_mult_82_n5752), .A2(u5_mult_82_n5753), 
        .A3(u5_mult_82_n5754), .ZN(u5_mult_82_CARRYB_32__36_) );
  NAND2_X1 u5_mult_82_U10951 ( .A1(u5_mult_82_ab_32__36_), .A2(
        u5_mult_82_CARRYB_31__36_), .ZN(u5_mult_82_n5754) );
  NAND2_X2 u5_mult_82_U10950 ( .A1(u5_mult_82_ab_32__36_), .A2(
        u5_mult_82_SUMB_31__37_), .ZN(u5_mult_82_n5753) );
  NAND2_X1 u5_mult_82_U10949 ( .A1(u5_mult_82_CARRYB_31__36_), .A2(
        u5_mult_82_SUMB_31__37_), .ZN(u5_mult_82_n5752) );
  XOR2_X2 u5_mult_82_U10948 ( .A(u5_mult_82_SUMB_31__37_), .B(u5_mult_82_n5751), .Z(u5_mult_82_SUMB_32__36_) );
  XOR2_X2 u5_mult_82_U10947 ( .A(u5_mult_82_CARRYB_31__36_), .B(
        u5_mult_82_ab_32__36_), .Z(u5_mult_82_n5751) );
  NAND3_X2 u5_mult_82_U10946 ( .A1(u5_mult_82_n5748), .A2(u5_mult_82_n5749), 
        .A3(u5_mult_82_n5750), .ZN(u5_mult_82_CARRYB_48__20_) );
  NAND2_X1 u5_mult_82_U10945 ( .A1(u5_mult_82_ab_48__20_), .A2(
        u5_mult_82_CARRYB_47__20_), .ZN(u5_mult_82_n5748) );
  NAND3_X2 u5_mult_82_U10944 ( .A1(u5_mult_82_n5745), .A2(u5_mult_82_n5746), 
        .A3(u5_mult_82_n5747), .ZN(u5_mult_82_CARRYB_47__21_) );
  NAND2_X2 u5_mult_82_U10943 ( .A1(u5_mult_82_ab_47__21_), .A2(
        u5_mult_82_SUMB_46__22_), .ZN(u5_mult_82_n5746) );
  NAND2_X1 u5_mult_82_U10942 ( .A1(u5_mult_82_ab_47__21_), .A2(u5_mult_82_n702), .ZN(u5_mult_82_n5745) );
  XOR2_X2 u5_mult_82_U10941 ( .A(u5_mult_82_n5744), .B(u5_mult_82_SUMB_46__22_), .Z(u5_mult_82_SUMB_47__21_) );
  NOR2_X2 u5_mult_82_U10940 ( .A1(u5_mult_82_net64921), .A2(
        u5_mult_82_net65711), .ZN(u5_mult_82_ab_23__36_) );
  NOR2_X1 u5_mult_82_U10939 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6642), 
        .ZN(u5_mult_82_ab_24__36_) );
  NOR2_X1 u5_mult_82_U10938 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6663), 
        .ZN(u5_mult_82_ab_28__36_) );
  NOR2_X1 u5_mult_82_U10937 ( .A1(u5_mult_82_n6780), .A2(u5_mult_82_n6536), 
        .ZN(u5_mult_82_ab_8__48_) );
  NAND3_X2 u5_mult_82_U10936 ( .A1(u5_mult_82_n5738), .A2(u5_mult_82_n5739), 
        .A3(u5_mult_82_n5740), .ZN(u5_mult_82_CARRYB_23__36_) );
  NAND2_X1 u5_mult_82_U10935 ( .A1(u5_mult_82_ab_23__36_), .A2(
        u5_mult_82_CARRYB_22__36_), .ZN(u5_mult_82_n5740) );
  NAND2_X2 u5_mult_82_U10934 ( .A1(u5_mult_82_ab_24__36_), .A2(
        u5_mult_82_SUMB_23__37_), .ZN(u5_mult_82_n5736) );
  NAND2_X1 u5_mult_82_U10933 ( .A1(u5_mult_82_ab_28__36_), .A2(
        u5_mult_82_CARRYB_27__36_), .ZN(u5_mult_82_n5734) );
  NAND2_X2 u5_mult_82_U10932 ( .A1(u5_mult_82_ab_28__36_), .A2(
        u5_mult_82_SUMB_27__37_), .ZN(u5_mult_82_n5733) );
  NAND2_X1 u5_mult_82_U10931 ( .A1(u5_mult_82_CARRYB_27__36_), .A2(
        u5_mult_82_SUMB_27__37_), .ZN(u5_mult_82_n5732) );
  NAND3_X2 u5_mult_82_U10930 ( .A1(u5_mult_82_n5729), .A2(u5_mult_82_n5730), 
        .A3(u5_mult_82_n5731), .ZN(u5_mult_82_CARRYB_10__46_) );
  NAND2_X1 u5_mult_82_U10929 ( .A1(u5_mult_82_ab_10__46_), .A2(
        u5_mult_82_CARRYB_9__46_), .ZN(u5_mult_82_n5729) );
  NAND2_X2 u5_mult_82_U10928 ( .A1(u5_mult_82_CARRYB_8__47_), .A2(
        u5_mult_82_SUMB_8__48_), .ZN(u5_mult_82_n5728) );
  NAND2_X2 u5_mult_82_U10927 ( .A1(u5_mult_82_ab_9__47_), .A2(
        u5_mult_82_SUMB_8__48_), .ZN(u5_mult_82_n5727) );
  XOR2_X2 u5_mult_82_U10926 ( .A(u5_mult_82_n5725), .B(u5_mult_82_SUMB_8__48_), 
        .Z(u5_mult_82_SUMB_9__47_) );
  NAND3_X2 u5_mult_82_U10925 ( .A1(u5_mult_82_n5722), .A2(u5_mult_82_n5723), 
        .A3(u5_mult_82_n5724), .ZN(u5_mult_82_CARRYB_8__48_) );
  NAND2_X2 u5_mult_82_U10924 ( .A1(u5_mult_82_ab_8__48_), .A2(
        u5_mult_82_CARRYB_7__48_), .ZN(u5_mult_82_n5724) );
  NAND2_X2 u5_mult_82_U10923 ( .A1(u5_mult_82_ab_8__48_), .A2(
        u5_mult_82_SUMB_7__49_), .ZN(u5_mult_82_n5723) );
  NAND3_X2 u5_mult_82_U10922 ( .A1(u5_mult_82_n5719), .A2(u5_mult_82_n5720), 
        .A3(u5_mult_82_n5721), .ZN(u5_mult_82_CARRYB_38__28_) );
  NAND2_X1 u5_mult_82_U10921 ( .A1(u5_mult_82_ab_38__28_), .A2(
        u5_mult_82_CARRYB_37__28_), .ZN(u5_mult_82_n5719) );
  NAND3_X2 u5_mult_82_U10920 ( .A1(u5_mult_82_n5716), .A2(u5_mult_82_n5717), 
        .A3(u5_mult_82_n5718), .ZN(u5_mult_82_CARRYB_37__29_) );
  NAND2_X2 u5_mult_82_U10919 ( .A1(u5_mult_82_CARRYB_36__29_), .A2(
        u5_mult_82_n1857), .ZN(u5_mult_82_n5718) );
  NAND2_X2 u5_mult_82_U10918 ( .A1(u5_mult_82_ab_37__29_), .A2(
        u5_mult_82_n1857), .ZN(u5_mult_82_n5717) );
  NAND2_X1 u5_mult_82_U10917 ( .A1(u5_mult_82_ab_37__29_), .A2(
        u5_mult_82_CARRYB_36__29_), .ZN(u5_mult_82_n5716) );
  XOR2_X2 u5_mult_82_U10916 ( .A(u5_mult_82_n5715), .B(u5_mult_82_n1857), .Z(
        u5_mult_82_SUMB_37__29_) );
  XOR2_X2 u5_mult_82_U10915 ( .A(u5_mult_82_ab_37__29_), .B(
        u5_mult_82_CARRYB_36__29_), .Z(u5_mult_82_n5715) );
  NAND3_X2 u5_mult_82_U10914 ( .A1(u5_mult_82_n5712), .A2(u5_mult_82_n5713), 
        .A3(u5_mult_82_n5714), .ZN(u5_mult_82_CARRYB_48__18_) );
  NAND2_X2 u5_mult_82_U10913 ( .A1(u5_mult_82_CARRYB_46__19_), .A2(
        u5_mult_82_n1608), .ZN(u5_mult_82_n5711) );
  NAND2_X2 u5_mult_82_U10912 ( .A1(u5_mult_82_ab_47__19_), .A2(
        u5_mult_82_n1608), .ZN(u5_mult_82_n5710) );
  NAND2_X1 u5_mult_82_U10911 ( .A1(u5_mult_82_ab_47__19_), .A2(
        u5_mult_82_CARRYB_46__19_), .ZN(u5_mult_82_n5709) );
  XOR2_X2 u5_mult_82_U10910 ( .A(u5_mult_82_ab_47__19_), .B(
        u5_mult_82_CARRYB_46__19_), .Z(u5_mult_82_n5708) );
  NAND2_X1 u5_mult_82_U10909 ( .A1(u5_mult_82_ab_32__30_), .A2(
        u5_mult_82_CARRYB_31__30_), .ZN(u5_mult_82_n5832) );
  NAND3_X2 u5_mult_82_U10908 ( .A1(u5_mult_82_n5705), .A2(u5_mult_82_n5706), 
        .A3(u5_mult_82_n5707), .ZN(u5_mult_82_CARRYB_13__32_) );
  NAND2_X1 u5_mult_82_U10907 ( .A1(u5_mult_82_CARRYB_12__32_), .A2(
        u5_mult_82_SUMB_12__33_), .ZN(u5_mult_82_n5707) );
  NAND2_X1 u5_mult_82_U10906 ( .A1(u5_mult_82_ab_13__32_), .A2(
        u5_mult_82_SUMB_12__33_), .ZN(u5_mult_82_n5706) );
  NAND2_X1 u5_mult_82_U10905 ( .A1(u5_mult_82_ab_13__32_), .A2(
        u5_mult_82_CARRYB_12__32_), .ZN(u5_mult_82_n5705) );
  NAND2_X2 u5_mult_82_U10904 ( .A1(u5_mult_82_ab_12__33_), .A2(
        u5_mult_82_SUMB_11__34_), .ZN(u5_mult_82_n5703) );
  NAND2_X1 u5_mult_82_U10903 ( .A1(u5_mult_82_ab_10__35_), .A2(
        u5_mult_82_CARRYB_9__35_), .ZN(u5_mult_82_n5699) );
  NAND3_X2 u5_mult_82_U10902 ( .A1(u5_mult_82_n5696), .A2(u5_mult_82_n5697), 
        .A3(u5_mult_82_n5698), .ZN(u5_mult_82_CARRYB_9__36_) );
  NAND2_X2 u5_mult_82_U10901 ( .A1(u5_mult_82_CARRYB_8__36_), .A2(
        u5_mult_82_n1763), .ZN(u5_mult_82_n5698) );
  NAND2_X2 u5_mult_82_U10900 ( .A1(u5_mult_82_ab_9__36_), .A2(u5_mult_82_n1763), .ZN(u5_mult_82_n5697) );
  NAND2_X1 u5_mult_82_U10899 ( .A1(u5_mult_82_ab_9__36_), .A2(
        u5_mult_82_CARRYB_8__36_), .ZN(u5_mult_82_n5696) );
  NAND3_X2 u5_mult_82_U10898 ( .A1(u5_mult_82_n5690), .A2(u5_mult_82_n5691), 
        .A3(u5_mult_82_n5692), .ZN(u5_mult_82_CARRYB_24__21_) );
  NAND2_X2 u5_mult_82_U10897 ( .A1(u5_mult_82_ab_24__21_), .A2(
        u5_mult_82_SUMB_23__22_), .ZN(u5_mult_82_n5691) );
  NAND2_X1 u5_mult_82_U10896 ( .A1(u5_mult_82_ab_24__21_), .A2(
        u5_mult_82_CARRYB_23__21_), .ZN(u5_mult_82_n5690) );
  XOR2_X2 u5_mult_82_U10895 ( .A(u5_mult_82_n5689), .B(u5_mult_82_SUMB_24__21_), .Z(u5_mult_82_SUMB_25__20_) );
  NAND3_X2 u5_mult_82_U10894 ( .A1(u5_mult_82_n5686), .A2(u5_mult_82_n5687), 
        .A3(u5_mult_82_n5688), .ZN(u5_mult_82_CARRYB_16__29_) );
  NAND2_X1 u5_mult_82_U10893 ( .A1(u5_mult_82_CARRYB_15__29_), .A2(
        u5_mult_82_SUMB_15__30_), .ZN(u5_mult_82_n5688) );
  NAND2_X1 u5_mult_82_U10892 ( .A1(u5_mult_82_ab_16__29_), .A2(
        u5_mult_82_SUMB_15__30_), .ZN(u5_mult_82_n5687) );
  NAND2_X2 u5_mult_82_U10891 ( .A1(u5_mult_82_n1527), .A2(
        u5_mult_82_SUMB_14__31_), .ZN(u5_mult_82_n5685) );
  NAND2_X2 u5_mult_82_U10890 ( .A1(u5_mult_82_ab_15__30_), .A2(
        u5_mult_82_SUMB_14__31_), .ZN(u5_mult_82_n5684) );
  XOR2_X2 u5_mult_82_U10889 ( .A(u5_mult_82_n5682), .B(u5_mult_82_n1673), .Z(
        u5_mult_82_SUMB_15__30_) );
  NAND2_X1 u5_mult_82_U10888 ( .A1(u5_mult_82_ab_46__11_), .A2(
        u5_mult_82_CARRYB_45__11_), .ZN(u5_mult_82_n5679) );
  NAND2_X2 u5_mult_82_U10887 ( .A1(u5_mult_82_ab_45__12_), .A2(
        u5_mult_82_n3709), .ZN(u5_mult_82_n5677) );
  NAND2_X1 u5_mult_82_U10886 ( .A1(u5_mult_82_ab_45__12_), .A2(
        u5_mult_82_CARRYB_44__12_), .ZN(u5_mult_82_n5676) );
  XOR2_X2 u5_mult_82_U10885 ( .A(u5_mult_82_n5675), .B(u5_mult_82_n3709), .Z(
        u5_mult_82_SUMB_45__12_) );
  XOR2_X2 u5_mult_82_U10884 ( .A(u5_mult_82_ab_45__12_), .B(
        u5_mult_82_CARRYB_44__12_), .Z(u5_mult_82_n5675) );
  XNOR2_X2 u5_mult_82_U10883 ( .A(u5_mult_82_ab_48__18_), .B(
        u5_mult_82_CARRYB_47__18_), .ZN(u5_mult_82_n5674) );
  XNOR2_X2 u5_mult_82_U10882 ( .A(u5_mult_82_CARRYB_49__18_), .B(
        u5_mult_82_ab_50__18_), .ZN(u5_mult_82_n5673) );
  XNOR2_X2 u5_mult_82_U10881 ( .A(u5_mult_82_SUMB_49__19_), .B(
        u5_mult_82_n5673), .ZN(u5_mult_82_SUMB_50__18_) );
  NOR2_X1 u5_mult_82_U10880 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6649), 
        .ZN(u5_mult_82_ab_26__38_) );
  NOR2_X1 u5_mult_82_U10879 ( .A1(u5_mult_82_net64683), .A2(
        u5_mult_82_net65371), .ZN(u5_mult_82_ab_42__23_) );
  NAND2_X2 u5_mult_82_U10878 ( .A1(u5_mult_82_CARRYB_47__18_), .A2(
        u5_mult_82_SUMB_47__19_), .ZN(u5_mult_82_n5714) );
  NOR2_X2 u5_mult_82_U10877 ( .A1(u5_mult_82_n6919), .A2(u5_mult_82_net65285), 
        .ZN(u5_mult_82_ab_47__18_) );
  NOR2_X1 u5_mult_82_U10876 ( .A1(u5_mult_82_net64665), .A2(
        u5_mult_82_net65353), .ZN(u5_mult_82_ab_43__22_) );
  NAND2_X1 u5_mult_82_U10875 ( .A1(u5_mult_82_ab_26__38_), .A2(
        u5_mult_82_CARRYB_25__38_), .ZN(u5_mult_82_n5672) );
  NAND2_X1 u5_mult_82_U10874 ( .A1(u5_mult_82_CARRYB_25__38_), .A2(
        u5_mult_82_SUMB_25__39_), .ZN(u5_mult_82_n5670) );
  NAND2_X1 u5_mult_82_U10873 ( .A1(u5_mult_82_ab_29__36_), .A2(
        u5_mult_82_CARRYB_28__36_), .ZN(u5_mult_82_n5667) );
  NAND2_X1 u5_mult_82_U10872 ( .A1(u5_mult_82_ab_28__37_), .A2(
        u5_mult_82_CARRYB_27__37_), .ZN(u5_mult_82_n5664) );
  NAND2_X1 u5_mult_82_U10871 ( .A1(u5_mult_82_ab_42__23_), .A2(
        u5_mult_82_CARRYB_41__23_), .ZN(u5_mult_82_n5663) );
  NAND2_X1 u5_mult_82_U10870 ( .A1(u5_mult_82_ab_47__18_), .A2(
        u5_mult_82_CARRYB_46__18_), .ZN(u5_mult_82_n5660) );
  NAND3_X2 u5_mult_82_U10869 ( .A1(u5_mult_82_n5655), .A2(u5_mult_82_n5656), 
        .A3(u5_mult_82_n5657), .ZN(u5_mult_82_CARRYB_43__22_) );
  NAND2_X2 u5_mult_82_U10868 ( .A1(u5_mult_82_ab_43__22_), .A2(
        u5_mult_82_SUMB_42__23_), .ZN(u5_mult_82_n5656) );
  XNOR2_X2 u5_mult_82_U10867 ( .A(u5_mult_82_CARRYB_22__38_), .B(
        u5_mult_82_ab_23__38_), .ZN(u5_mult_82_n5653) );
  XNOR2_X2 u5_mult_82_U10866 ( .A(u5_mult_82_SUMB_52__13_), .B(
        u5_mult_82_n5652), .ZN(u5_mult_82_n5651) );
  XNOR2_X2 u5_mult_82_U10865 ( .A(u5_mult_82_CARRYB_46__18_), .B(
        u5_mult_82_ab_47__18_), .ZN(u5_mult_82_n5650) );
  XNOR2_X2 u5_mult_82_U10864 ( .A(u5_mult_82_CARRYB_27__36_), .B(
        u5_mult_82_ab_28__36_), .ZN(u5_mult_82_n5648) );
  NOR2_X1 u5_mult_82_U10863 ( .A1(u5_mult_82_n6818), .A2(u5_mult_82_n6580), 
        .ZN(u5_mult_82_ab_14__42_) );
  NOR2_X1 u5_mult_82_U10862 ( .A1(u5_mult_82_n6806), .A2(u5_mult_82_n6559), 
        .ZN(u5_mult_82_ab_11__44_) );
  NAND3_X2 u5_mult_82_U10861 ( .A1(u5_mult_82_n5645), .A2(u5_mult_82_n5646), 
        .A3(u5_mult_82_n5647), .ZN(u5_mult_82_CARRYB_14__42_) );
  NAND2_X1 u5_mult_82_U10860 ( .A1(u5_mult_82_ab_14__42_), .A2(
        u5_mult_82_CARRYB_13__42_), .ZN(u5_mult_82_n5647) );
  NAND2_X2 u5_mult_82_U10859 ( .A1(u5_mult_82_ab_14__42_), .A2(
        u5_mult_82_n1794), .ZN(u5_mult_82_n5646) );
  INV_X4 u5_mult_82_U10858 ( .A(u5_mult_82_n5640), .ZN(u5_mult_82_n5641) );
  INV_X2 u5_mult_82_U10857 ( .A(u5_mult_82_CARRYB_42__22_), .ZN(
        u5_mult_82_n5640) );
  NAND2_X1 u5_mult_82_U10856 ( .A1(u5_mult_82_SUMB_47__16_), .A2(
        u5_mult_82_CARRYB_47__15_), .ZN(u5_mult_82_n5855) );
  NAND2_X1 u5_mult_82_U10855 ( .A1(u5_mult_82_ab_48__15_), .A2(
        u5_mult_82_SUMB_47__16_), .ZN(u5_mult_82_n5853) );
  INV_X4 u5_mult_82_U10854 ( .A(u5_mult_82_CARRYB_52__12_), .ZN(
        u5_mult_82_n5652) );
  XNOR2_X2 u5_mult_82_U10853 ( .A(u5_mult_82_SUMB_43__12_), .B(
        u5_mult_82_net79780), .ZN(u5_mult_82_SUMB_44__11_) );
  XNOR2_X2 u5_mult_82_U10852 ( .A(u5_mult_82_n5641), .B(u5_mult_82_ab_43__22_), 
        .ZN(u5_mult_82_n5639) );
  XNOR2_X2 u5_mult_82_U10851 ( .A(u5_mult_82_SUMB_42__23_), .B(
        u5_mult_82_n5639), .ZN(u5_mult_82_SUMB_43__22_) );
  XNOR2_X2 u5_mult_82_U10850 ( .A(u5_mult_82_ab_45__3_), .B(u5_mult_82_n1721), 
        .ZN(u5_mult_82_n5638) );
  NOR2_X1 u5_mult_82_U10849 ( .A1(u5_mult_82_n6960), .A2(u5_mult_82_net65355), 
        .ZN(u5_mult_82_ab_43__2_) );
  NOR2_X1 u5_mult_82_U10848 ( .A1(u5_mult_82_n6960), .A2(u5_mult_82_net65375), 
        .ZN(u5_mult_82_ab_42__2_) );
  NOR2_X1 u5_mult_82_U10847 ( .A1(u5_mult_82_net64959), .A2(
        u5_mult_82_net66017), .ZN(u5_mult_82_ab_6__38_) );
  NOR2_X1 u5_mult_82_U10846 ( .A1(u5_mult_82_n6876), .A2(u5_mult_82_n6602), 
        .ZN(u5_mult_82_ab_17__27_) );
  NAND3_X4 u5_mult_82_U10845 ( .A1(u5_mult_82_n5635), .A2(u5_mult_82_n5636), 
        .A3(u5_mult_82_n5637), .ZN(u5_mult_82_CARRYB_43__2_) );
  NAND2_X1 u5_mult_82_U10844 ( .A1(u5_mult_82_ab_43__2_), .A2(
        u5_mult_82_CARRYB_42__2_), .ZN(u5_mult_82_n5637) );
  NAND2_X2 u5_mult_82_U10843 ( .A1(u5_mult_82_ab_43__2_), .A2(
        u5_mult_82_SUMB_42__3_), .ZN(u5_mult_82_n5636) );
  XOR2_X2 u5_mult_82_U10842 ( .A(u5_mult_82_SUMB_42__3_), .B(u5_mult_82_n5634), 
        .Z(u5_mult_82_SUMB_43__2_) );
  XOR2_X2 u5_mult_82_U10841 ( .A(u5_mult_82_CARRYB_42__2_), .B(
        u5_mult_82_ab_43__2_), .Z(u5_mult_82_n5634) );
  NAND2_X2 u5_mult_82_U10840 ( .A1(u5_mult_82_ab_45__2_), .A2(
        u5_mult_82_CARRYB_44__2_), .ZN(u5_mult_82_n5629) );
  XOR2_X2 u5_mult_82_U10839 ( .A(u5_mult_82_n5627), .B(
        u5_mult_82_CARRYB_44__2_), .Z(u5_mult_82_SUMB_45__2_) );
  NAND3_X2 u5_mult_82_U10838 ( .A1(u5_mult_82_n5624), .A2(u5_mult_82_n5625), 
        .A3(u5_mult_82_n5626), .ZN(u5_mult_82_CARRYB_44__2_) );
  NAND2_X1 u5_mult_82_U10837 ( .A1(u5_mult_82_CARRYB_43__2_), .A2(
        u5_mult_82_SUMB_43__3_), .ZN(u5_mult_82_n5626) );
  NAND2_X2 u5_mult_82_U10836 ( .A1(u5_mult_82_ab_44__2_), .A2(
        u5_mult_82_SUMB_43__3_), .ZN(u5_mult_82_n5625) );
  NAND2_X2 u5_mult_82_U10835 ( .A1(u5_mult_82_ab_44__2_), .A2(
        u5_mult_82_CARRYB_43__2_), .ZN(u5_mult_82_n5624) );
  NAND3_X4 u5_mult_82_U10834 ( .A1(u5_mult_82_n5623), .A2(u5_mult_82_n5622), 
        .A3(u5_mult_82_n5621), .ZN(u5_mult_82_CARRYB_8__36_) );
  NAND3_X2 u5_mult_82_U10833 ( .A1(u5_mult_82_n5618), .A2(u5_mult_82_n5619), 
        .A3(u5_mult_82_n5620), .ZN(u5_mult_82_CARRYB_7__37_) );
  NAND2_X2 u5_mult_82_U10832 ( .A1(u5_mult_82_ab_7__37_), .A2(
        u5_mult_82_SUMB_6__38_), .ZN(u5_mult_82_n5619) );
  NAND2_X1 u5_mult_82_U10831 ( .A1(u5_mult_82_ab_7__37_), .A2(
        u5_mult_82_CARRYB_6__37_), .ZN(u5_mult_82_n5618) );
  NAND3_X2 u5_mult_82_U10830 ( .A1(u5_mult_82_n5615), .A2(u5_mult_82_n5616), 
        .A3(u5_mult_82_n5617), .ZN(u5_mult_82_CARRYB_6__38_) );
  NAND2_X1 u5_mult_82_U10829 ( .A1(u5_mult_82_ab_6__38_), .A2(
        u5_mult_82_CARRYB_5__38_), .ZN(u5_mult_82_n5617) );
  XOR2_X2 u5_mult_82_U10828 ( .A(u5_mult_82_CARRYB_5__38_), .B(
        u5_mult_82_ab_6__38_), .Z(u5_mult_82_n5614) );
  NAND2_X1 u5_mult_82_U10827 ( .A1(u5_mult_82_ab_20__24_), .A2(
        u5_mult_82_CARRYB_19__24_), .ZN(u5_mult_82_n5611) );
  NAND3_X2 u5_mult_82_U10826 ( .A1(u5_mult_82_n5608), .A2(u5_mult_82_n5609), 
        .A3(u5_mult_82_n5610), .ZN(u5_mult_82_CARRYB_19__25_) );
  NAND2_X2 u5_mult_82_U10825 ( .A1(u5_mult_82_n37), .A2(u5_mult_82_ab_19__25_), 
        .ZN(u5_mult_82_n5609) );
  NAND2_X1 u5_mult_82_U10824 ( .A1(u5_mult_82_ab_19__25_), .A2(
        u5_mult_82_CARRYB_18__25_), .ZN(u5_mult_82_n5608) );
  XNOR2_X2 u5_mult_82_U10823 ( .A(u5_mult_82_ab_46__11_), .B(
        u5_mult_82_CARRYB_45__11_), .ZN(u5_mult_82_n5605) );
  XNOR2_X2 u5_mult_82_U10822 ( .A(u5_mult_82_n5605), .B(
        u5_mult_82_SUMB_45__12_), .ZN(u5_mult_82_SUMB_46__11_) );
  NAND3_X4 u5_mult_82_U10821 ( .A1(u5_mult_82_n5602), .A2(u5_mult_82_n5603), 
        .A3(u5_mult_82_n5604), .ZN(u5_mult_82_CARRYB_34__31_) );
  NAND2_X2 u5_mult_82_U10820 ( .A1(u5_mult_82_CARRYB_33__31_), .A2(
        u5_mult_82_SUMB_33__32_), .ZN(u5_mult_82_n5604) );
  NAND2_X2 u5_mult_82_U10819 ( .A1(u5_mult_82_ab_34__31_), .A2(
        u5_mult_82_SUMB_33__32_), .ZN(u5_mult_82_n5603) );
  NAND2_X1 u5_mult_82_U10818 ( .A1(u5_mult_82_ab_34__31_), .A2(
        u5_mult_82_CARRYB_33__31_), .ZN(u5_mult_82_n5602) );
  NAND2_X2 u5_mult_82_U10817 ( .A1(u5_mult_82_n72), .A2(
        u5_mult_82_CARRYB_32__32_), .ZN(u5_mult_82_n5601) );
  NAND2_X2 u5_mult_82_U10816 ( .A1(u5_mult_82_n72), .A2(u5_mult_82_ab_33__32_), 
        .ZN(u5_mult_82_n5600) );
  NAND2_X1 u5_mult_82_U10815 ( .A1(u5_mult_82_ab_33__32_), .A2(
        u5_mult_82_CARRYB_32__32_), .ZN(u5_mult_82_n5599) );
  XOR2_X2 u5_mult_82_U10814 ( .A(u5_mult_82_n5598), .B(u5_mult_82_SUMB_33__32_), .Z(u5_mult_82_SUMB_34__31_) );
  XOR2_X2 u5_mult_82_U10813 ( .A(u5_mult_82_ab_34__31_), .B(
        u5_mult_82_CARRYB_33__31_), .Z(u5_mult_82_n5598) );
  NAND3_X2 u5_mult_82_U10812 ( .A1(u5_mult_82_n5595), .A2(u5_mult_82_n5596), 
        .A3(u5_mult_82_n5597), .ZN(u5_mult_82_CARRYB_35__29_) );
  NAND2_X1 u5_mult_82_U10811 ( .A1(u5_mult_82_ab_35__29_), .A2(
        u5_mult_82_SUMB_34__30_), .ZN(u5_mult_82_n5597) );
  NAND2_X1 u5_mult_82_U10810 ( .A1(u5_mult_82_ab_35__29_), .A2(
        u5_mult_82_CARRYB_34__29_), .ZN(u5_mult_82_n5596) );
  NAND2_X1 u5_mult_82_U10809 ( .A1(u5_mult_82_SUMB_34__30_), .A2(
        u5_mult_82_CARRYB_34__29_), .ZN(u5_mult_82_n5595) );
  NAND3_X4 u5_mult_82_U10808 ( .A1(u5_mult_82_n5830), .A2(u5_mult_82_n5831), 
        .A3(u5_mult_82_n5832), .ZN(u5_mult_82_CARRYB_32__30_) );
  NAND2_X1 u5_mult_82_U10807 ( .A1(u5_mult_82_ab_26__43_), .A2(
        u5_mult_82_CARRYB_25__43_), .ZN(u5_mult_82_n5592) );
  NAND2_X2 u5_mult_82_U10806 ( .A1(u5_mult_82_n1568), .A2(
        u5_mult_82_SUMB_24__45_), .ZN(u5_mult_82_n5591) );
  NAND2_X2 u5_mult_82_U10805 ( .A1(u5_mult_82_ab_25__44_), .A2(
        u5_mult_82_SUMB_24__45_), .ZN(u5_mult_82_n5590) );
  XOR2_X2 u5_mult_82_U10804 ( .A(u5_mult_82_n5588), .B(u5_mult_82_SUMB_24__45_), .Z(u5_mult_82_SUMB_25__44_) );
  XOR2_X2 u5_mult_82_U10803 ( .A(u5_mult_82_ab_25__44_), .B(u5_mult_82_n1568), 
        .Z(u5_mult_82_n5588) );
  NAND3_X2 u5_mult_82_U10802 ( .A1(u5_mult_82_n5585), .A2(u5_mult_82_n5586), 
        .A3(u5_mult_82_n5587), .ZN(u5_mult_82_CARRYB_42__27_) );
  NAND2_X1 u5_mult_82_U10801 ( .A1(u5_mult_82_SUMB_41__28_), .A2(
        u5_mult_82_CARRYB_41__27_), .ZN(u5_mult_82_n5587) );
  NAND2_X1 u5_mult_82_U10800 ( .A1(u5_mult_82_ab_42__27_), .A2(
        u5_mult_82_SUMB_41__28_), .ZN(u5_mult_82_n5586) );
  NAND2_X1 u5_mult_82_U10799 ( .A1(u5_mult_82_ab_42__27_), .A2(
        u5_mult_82_CARRYB_41__27_), .ZN(u5_mult_82_n5585) );
  NAND2_X1 u5_mult_82_U10798 ( .A1(u5_mult_82_ab_41__28_), .A2(
        u5_mult_82_CARRYB_40__28_), .ZN(u5_mult_82_n5582) );
  XOR2_X2 u5_mult_82_U10797 ( .A(u5_mult_82_n5581), .B(u5_mult_82_SUMB_41__28_), .Z(u5_mult_82_SUMB_42__27_) );
  XOR2_X2 u5_mult_82_U10796 ( .A(u5_mult_82_ab_41__28_), .B(
        u5_mult_82_CARRYB_40__28_), .Z(u5_mult_82_n5580) );
  NAND3_X2 u5_mult_82_U10795 ( .A1(u5_mult_82_n5577), .A2(u5_mult_82_n5578), 
        .A3(u5_mult_82_n5579), .ZN(u5_mult_82_CARRYB_36__33_) );
  NAND2_X1 u5_mult_82_U10794 ( .A1(u5_mult_82_CARRYB_35__33_), .A2(
        u5_mult_82_SUMB_35__34_), .ZN(u5_mult_82_n5579) );
  NAND2_X1 u5_mult_82_U10793 ( .A1(u5_mult_82_ab_36__33_), .A2(
        u5_mult_82_SUMB_35__34_), .ZN(u5_mult_82_n5578) );
  NAND3_X4 u5_mult_82_U10792 ( .A1(u5_mult_82_n5574), .A2(u5_mult_82_n5575), 
        .A3(u5_mult_82_n5576), .ZN(u5_mult_82_CARRYB_35__34_) );
  NAND2_X2 u5_mult_82_U10791 ( .A1(u5_mult_82_CARRYB_34__34_), .A2(
        u5_mult_82_n442), .ZN(u5_mult_82_n5576) );
  NAND2_X2 u5_mult_82_U10790 ( .A1(u5_mult_82_ab_35__34_), .A2(u5_mult_82_n442), .ZN(u5_mult_82_n5575) );
  NAND2_X2 u5_mult_82_U10789 ( .A1(u5_mult_82_ab_35__34_), .A2(
        u5_mult_82_CARRYB_34__34_), .ZN(u5_mult_82_n5574) );
  XOR2_X2 u5_mult_82_U10788 ( .A(u5_mult_82_n5573), .B(u5_mult_82_SUMB_35__34_), .Z(u5_mult_82_SUMB_36__33_) );
  XOR2_X2 u5_mult_82_U10787 ( .A(u5_mult_82_ab_36__33_), .B(
        u5_mult_82_CARRYB_35__33_), .Z(u5_mult_82_n5573) );
  XOR2_X2 u5_mult_82_U10786 ( .A(u5_mult_82_n5572), .B(u5_mult_82_n442), .Z(
        u5_mult_82_SUMB_35__34_) );
  XOR2_X2 u5_mult_82_U10785 ( .A(u5_mult_82_ab_35__34_), .B(
        u5_mult_82_CARRYB_34__34_), .Z(u5_mult_82_n5572) );
  NAND3_X2 u5_mult_82_U10784 ( .A1(u5_mult_82_n5569), .A2(u5_mult_82_n5570), 
        .A3(u5_mult_82_n5571), .ZN(u5_mult_82_CARRYB_51__18_) );
  NAND2_X1 u5_mult_82_U10783 ( .A1(u5_mult_82_CARRYB_50__18_), .A2(
        u5_mult_82_SUMB_50__19_), .ZN(u5_mult_82_n5571) );
  NAND2_X1 u5_mult_82_U10782 ( .A1(u5_mult_82_ab_51__18_), .A2(
        u5_mult_82_CARRYB_50__18_), .ZN(u5_mult_82_n5569) );
  NAND2_X2 u5_mult_82_U10781 ( .A1(u5_mult_82_ab_50__19_), .A2(
        u5_mult_82_n1841), .ZN(u5_mult_82_n5567) );
  XOR2_X2 u5_mult_82_U10780 ( .A(u5_mult_82_CARRYB_52__16_), .B(
        u5_mult_82_SUMB_52__17_), .Z(u5_mult_82_n5565) );
  NOR2_X1 u5_mult_82_U10779 ( .A1(u5_mult_82_net64939), .A2(u5_mult_82_n6642), 
        .ZN(u5_mult_82_ab_24__37_) );
  NAND3_X4 u5_mult_82_U10778 ( .A1(u5_mult_82_n5735), .A2(u5_mult_82_n5736), 
        .A3(u5_mult_82_n5737), .ZN(u5_mult_82_CARRYB_24__36_) );
  NOR2_X1 u5_mult_82_U10777 ( .A1(u5_mult_82_net64921), .A2(
        u5_mult_82_net65675), .ZN(u5_mult_82_ab_25__36_) );
  INV_X4 u5_mult_82_U10776 ( .A(u5_mult_82_n5649), .ZN(u5_mult_82_n5562) );
  NAND2_X1 u5_mult_82_U10775 ( .A1(u5_mult_82_SUMB_31__31_), .A2(
        u5_mult_82_n5649), .ZN(u5_mult_82_n5563) );
  NAND3_X2 u5_mult_82_U10774 ( .A1(u5_mult_82_n5555), .A2(u5_mult_82_n5556), 
        .A3(u5_mult_82_n5557), .ZN(u5_mult_82_CARRYB_25__36_) );
  NAND2_X2 u5_mult_82_U10773 ( .A1(u5_mult_82_CARRYB_24__36_), .A2(
        u5_mult_82_SUMB_24__37_), .ZN(u5_mult_82_n5555) );
  XNOR2_X2 u5_mult_82_U10772 ( .A(u5_mult_82_n5554), .B(
        u5_mult_82_SUMB_19__43_), .ZN(u5_mult_82_SUMB_20__42_) );
  XNOR2_X2 u5_mult_82_U10771 ( .A(u5_mult_82_CARRYB_12__44_), .B(
        u5_mult_82_ab_13__44_), .ZN(u5_mult_82_n5553) );
  XNOR2_X2 u5_mult_82_U10770 ( .A(u5_mult_82_n5553), .B(
        u5_mult_82_SUMB_12__45_), .ZN(u5_mult_82_SUMB_13__44_) );
  INV_X4 u5_mult_82_U10769 ( .A(u5_mult_82_n5551), .ZN(u5_mult_82_n5552) );
  XOR2_X2 u5_mult_82_U10768 ( .A(u5_mult_82_n5654), .B(
        u5_mult_82_CARRYB_17__46_), .Z(u5_mult_82_n5550) );
  NAND2_X2 u5_mult_82_U10767 ( .A1(u5_mult_82_CARRYB_23__36_), .A2(
        u5_mult_82_SUMB_23__37_), .ZN(u5_mult_82_n5735) );
  XNOR2_X2 u5_mult_82_U10766 ( .A(u5_mult_82_CARRYB_15__42_), .B(
        u5_mult_82_n5549), .ZN(u5_mult_82_n6219) );
  NOR2_X1 u5_mult_82_U10765 ( .A1(u5_mult_82_net64885), .A2(u5_mult_82_n6628), 
        .ZN(u5_mult_82_ab_21__34_) );
  NAND3_X2 u5_mult_82_U10764 ( .A1(u5_mult_82_n5545), .A2(u5_mult_82_n5546), 
        .A3(u5_mult_82_n5547), .ZN(u5_mult_82_CARRYB_26__29_) );
  NAND2_X1 u5_mult_82_U10763 ( .A1(u5_mult_82_ab_26__29_), .A2(
        u5_mult_82_CARRYB_25__29_), .ZN(u5_mult_82_n5547) );
  NAND2_X2 u5_mult_82_U10762 ( .A1(u5_mult_82_ab_26__29_), .A2(
        u5_mult_82_n1428), .ZN(u5_mult_82_n5546) );
  XNOR2_X2 u5_mult_82_U10761 ( .A(u5_mult_82_CARRYB_46__12_), .B(
        u5_mult_82_n5541), .ZN(u5_mult_82_n6230) );
  NOR2_X1 u5_mult_82_U10760 ( .A1(u5_mult_82_n6886), .A2(u5_mult_82_n6650), 
        .ZN(u5_mult_82_ab_26__25_) );
  NOR2_X1 u5_mult_82_U10759 ( .A1(u5_mult_82_net64559), .A2(u5_mult_82_n6721), 
        .ZN(u5_mult_82_ab_37__16_) );
  NAND2_X1 u5_mult_82_U10758 ( .A1(u5_mult_82_ab_28__23_), .A2(
        u5_mult_82_CARRYB_27__23_), .ZN(u5_mult_82_n5538) );
  NAND2_X2 u5_mult_82_U10757 ( .A1(u5_mult_82_ab_27__24_), .A2(
        u5_mult_82_SUMB_26__25_), .ZN(u5_mult_82_n5536) );
  NAND2_X1 u5_mult_82_U10756 ( .A1(u5_mult_82_ab_27__24_), .A2(
        u5_mult_82_CARRYB_26__24_), .ZN(u5_mult_82_n5535) );
  NAND3_X2 u5_mult_82_U10755 ( .A1(u5_mult_82_n5532), .A2(u5_mult_82_n5533), 
        .A3(u5_mult_82_n5534), .ZN(u5_mult_82_CARRYB_26__25_) );
  NAND2_X1 u5_mult_82_U10754 ( .A1(u5_mult_82_ab_26__25_), .A2(
        u5_mult_82_CARRYB_25__25_), .ZN(u5_mult_82_n5534) );
  NAND2_X2 u5_mult_82_U10753 ( .A1(u5_mult_82_ab_26__25_), .A2(
        u5_mult_82_SUMB_25__26_), .ZN(u5_mult_82_n5533) );
  NAND3_X2 u5_mult_82_U10752 ( .A1(u5_mult_82_n5529), .A2(u5_mult_82_n5530), 
        .A3(u5_mult_82_n5531), .ZN(u5_mult_82_CARRYB_40__14_) );
  NAND2_X1 u5_mult_82_U10751 ( .A1(u5_mult_82_CARRYB_39__14_), .A2(
        u5_mult_82_SUMB_39__15_), .ZN(u5_mult_82_n5531) );
  NAND2_X1 u5_mult_82_U10750 ( .A1(u5_mult_82_ab_40__14_), .A2(
        u5_mult_82_SUMB_39__15_), .ZN(u5_mult_82_n5530) );
  NAND2_X1 u5_mult_82_U10749 ( .A1(u5_mult_82_ab_40__14_), .A2(
        u5_mult_82_CARRYB_39__14_), .ZN(u5_mult_82_n5529) );
  NAND2_X1 u5_mult_82_U10748 ( .A1(u5_mult_82_ab_37__16_), .A2(
        u5_mult_82_CARRYB_36__16_), .ZN(u5_mult_82_n5525) );
  NAND2_X1 u5_mult_82_U10747 ( .A1(u5_mult_82_ab_21__34_), .A2(
        u5_mult_82_CARRYB_20__34_), .ZN(u5_mult_82_n5544) );
  XNOR2_X2 u5_mult_82_U10746 ( .A(u5_mult_82_n5522), .B(
        u5_mult_82_CARRYB_32__30_), .ZN(u5_mult_82_n5867) );
  XNOR2_X2 u5_mult_82_U10745 ( .A(u5_mult_82_n5520), .B(
        u5_mult_82_SUMB_42__14_), .ZN(u5_mult_82_SUMB_43__13_) );
  NAND2_X1 u5_mult_82_U10744 ( .A1(u5_mult_82_ab_21__37_), .A2(
        u5_mult_82_CARRYB_20__37_), .ZN(u5_mult_82_n5517) );
  NAND3_X4 u5_mult_82_U10743 ( .A1(u5_mult_82_n5514), .A2(u5_mult_82_n5515), 
        .A3(u5_mult_82_n5516), .ZN(u5_mult_82_CARRYB_20__38_) );
  NAND2_X2 u5_mult_82_U10742 ( .A1(u5_mult_82_CARRYB_19__38_), .A2(
        u5_mult_82_SUMB_19__39_), .ZN(u5_mult_82_n5516) );
  NAND2_X2 u5_mult_82_U10741 ( .A1(u5_mult_82_ab_20__38_), .A2(
        u5_mult_82_SUMB_19__39_), .ZN(u5_mult_82_n5515) );
  NAND2_X1 u5_mult_82_U10740 ( .A1(u5_mult_82_ab_20__38_), .A2(
        u5_mult_82_CARRYB_19__38_), .ZN(u5_mult_82_n5514) );
  XOR2_X2 u5_mult_82_U10739 ( .A(u5_mult_82_SUMB_19__39_), .B(u5_mult_82_n5513), .Z(u5_mult_82_SUMB_20__38_) );
  XOR2_X2 u5_mult_82_U10738 ( .A(u5_mult_82_ab_20__38_), .B(
        u5_mult_82_CARRYB_19__38_), .Z(u5_mult_82_n5513) );
  XNOR2_X2 u5_mult_82_U10737 ( .A(u5_mult_82_n5512), .B(
        u5_mult_82_CARRYB_34__20_), .ZN(u5_mult_82_n5892) );
  NAND2_X1 u5_mult_82_U10736 ( .A1(u5_mult_82_ab_24__32_), .A2(
        u5_mult_82_CARRYB_23__32_), .ZN(u5_mult_82_n5511) );
  NAND2_X2 u5_mult_82_U10735 ( .A1(u5_mult_82_ab_24__32_), .A2(u5_mult_82_n433), .ZN(u5_mult_82_n5510) );
  XNOR2_X2 u5_mult_82_U10734 ( .A(u5_mult_82_ab_49__10_), .B(
        u5_mult_82_CARRYB_48__10_), .ZN(u5_mult_82_n5508) );
  INV_X4 u5_mult_82_U10733 ( .A(u5_mult_82_CARRYB_22__34_), .ZN(
        u5_mult_82_n5506) );
  NAND3_X2 u5_mult_82_U10732 ( .A1(u5_mult_82_n5503), .A2(u5_mult_82_n5504), 
        .A3(u5_mult_82_n5505), .ZN(u5_mult_82_CARRYB_4__39_) );
  NAND2_X1 u5_mult_82_U10731 ( .A1(u5_mult_82_CARRYB_3__39_), .A2(
        u5_mult_82_SUMB_3__40_), .ZN(u5_mult_82_n5505) );
  NAND2_X1 u5_mult_82_U10730 ( .A1(u5_mult_82_ab_4__39_), .A2(
        u5_mult_82_SUMB_3__40_), .ZN(u5_mult_82_n5504) );
  NAND2_X1 u5_mult_82_U10729 ( .A1(u5_mult_82_ab_4__39_), .A2(
        u5_mult_82_CARRYB_3__39_), .ZN(u5_mult_82_n5503) );
  NAND3_X2 u5_mult_82_U10728 ( .A1(u5_mult_82_n5502), .A2(u5_mult_82_n5501), 
        .A3(u5_mult_82_n5500), .ZN(u5_mult_82_CARRYB_3__40_) );
  NAND2_X2 u5_mult_82_U10727 ( .A1(u5_mult_82_ab_3__40_), .A2(
        u5_mult_82_SUMB_2__41_), .ZN(u5_mult_82_n5501) );
  NAND2_X1 u5_mult_82_U10726 ( .A1(u5_mult_82_ab_3__40_), .A2(
        u5_mult_82_CARRYB_2__40_), .ZN(u5_mult_82_n5500) );
  XOR2_X2 u5_mult_82_U10725 ( .A(u5_mult_82_n5499), .B(u5_mult_82_n1778), .Z(
        u5_mult_82_SUMB_3__40_) );
  NAND3_X2 u5_mult_82_U10724 ( .A1(u5_mult_82_n970), .A2(u5_mult_82_n5497), 
        .A3(u5_mult_82_n5498), .ZN(u5_mult_82_CARRYB_21__22_) );
  NAND2_X1 u5_mult_82_U10723 ( .A1(u5_mult_82_ab_21__22_), .A2(
        u5_mult_82_SUMB_20__23_), .ZN(u5_mult_82_n5497) );
  NAND3_X2 u5_mult_82_U10722 ( .A1(u5_mult_82_n5494), .A2(u5_mult_82_n5495), 
        .A3(u5_mult_82_n5496), .ZN(u5_mult_82_CARRYB_20__23_) );
  NAND2_X2 u5_mult_82_U10721 ( .A1(u5_mult_82_ab_20__23_), .A2(
        u5_mult_82_SUMB_19__24_), .ZN(u5_mult_82_n5495) );
  NAND2_X1 u5_mult_82_U10720 ( .A1(u5_mult_82_ab_20__23_), .A2(
        u5_mult_82_CARRYB_19__23_), .ZN(u5_mult_82_n5494) );
  NAND2_X1 u5_mult_82_U10719 ( .A1(u5_mult_82_ab_44__8_), .A2(
        u5_mult_82_CARRYB_43__8_), .ZN(u5_mult_82_n5491) );
  NAND3_X2 u5_mult_82_U10718 ( .A1(u5_mult_82_n5488), .A2(u5_mult_82_n5489), 
        .A3(u5_mult_82_n5490), .ZN(u5_mult_82_CARRYB_43__9_) );
  NAND2_X2 u5_mult_82_U10717 ( .A1(u5_mult_82_CARRYB_42__9_), .A2(
        u5_mult_82_SUMB_42__10_), .ZN(u5_mult_82_n5490) );
  NOR2_X1 u5_mult_82_U10716 ( .A1(u5_mult_82_n6813), .A2(u5_mult_82_n6585), 
        .ZN(u5_mult_82_ab_15__43_) );
  NOR2_X1 u5_mult_82_U10715 ( .A1(u5_mult_82_n6813), .A2(u5_mult_82_n6580), 
        .ZN(u5_mult_82_ab_14__43_) );
  NAND3_X2 u5_mult_82_U10714 ( .A1(u5_mult_82_n5485), .A2(u5_mult_82_n5486), 
        .A3(u5_mult_82_n5487), .ZN(u5_mult_82_CARRYB_15__43_) );
  NAND2_X1 u5_mult_82_U10713 ( .A1(u5_mult_82_ab_15__43_), .A2(
        u5_mult_82_CARRYB_14__43_), .ZN(u5_mult_82_n5487) );
  NAND2_X2 u5_mult_82_U10712 ( .A1(u5_mult_82_ab_15__43_), .A2(
        u5_mult_82_SUMB_14__44_), .ZN(u5_mult_82_n5486) );
  NAND2_X1 u5_mult_82_U10711 ( .A1(u5_mult_82_CARRYB_14__43_), .A2(
        u5_mult_82_SUMB_14__44_), .ZN(u5_mult_82_n5485) );
  XOR2_X2 u5_mult_82_U10710 ( .A(u5_mult_82_SUMB_14__44_), .B(u5_mult_82_n5484), .Z(u5_mult_82_SUMB_15__43_) );
  XOR2_X2 u5_mult_82_U10709 ( .A(u5_mult_82_CARRYB_14__43_), .B(
        u5_mult_82_ab_15__43_), .Z(u5_mult_82_n5484) );
  NAND3_X2 u5_mult_82_U10708 ( .A1(u5_mult_82_n5481), .A2(u5_mult_82_n5482), 
        .A3(u5_mult_82_n5483), .ZN(u5_mult_82_CARRYB_14__43_) );
  NAND2_X1 u5_mult_82_U10707 ( .A1(u5_mult_82_ab_14__43_), .A2(
        u5_mult_82_SUMB_13__44_), .ZN(u5_mult_82_n5483) );
  NAND2_X2 u5_mult_82_U10706 ( .A1(u5_mult_82_ab_14__43_), .A2(
        u5_mult_82_CARRYB_13__43_), .ZN(u5_mult_82_n5482) );
  XOR2_X2 u5_mult_82_U10705 ( .A(u5_mult_82_CARRYB_13__43_), .B(
        u5_mult_82_n5480), .Z(u5_mult_82_SUMB_14__43_) );
  XOR2_X2 u5_mult_82_U10704 ( .A(u5_mult_82_SUMB_13__44_), .B(
        u5_mult_82_ab_14__43_), .Z(u5_mult_82_n5480) );
  NOR2_X1 u5_mult_82_U10703 ( .A1(u5_mult_82_n6862), .A2(u5_mult_82_n6663), 
        .ZN(u5_mult_82_ab_28__29_) );
  NAND2_X2 u5_mult_82_U10702 ( .A1(u5_mult_82_SUMB_27__30_), .A2(
        u5_mult_82_ab_28__29_), .ZN(u5_mult_82_n5478) );
  NAND3_X2 u5_mult_82_U10701 ( .A1(u5_mult_82_n5474), .A2(u5_mult_82_n5475), 
        .A3(u5_mult_82_n5476), .ZN(u5_mult_82_CARRYB_25__32_) );
  NAND2_X1 u5_mult_82_U10700 ( .A1(u5_mult_82_SUMB_24__33_), .A2(
        u5_mult_82_CARRYB_24__32_), .ZN(u5_mult_82_n5476) );
  NAND2_X1 u5_mult_82_U10699 ( .A1(u5_mult_82_ab_25__32_), .A2(
        u5_mult_82_CARRYB_24__32_), .ZN(u5_mult_82_n5474) );
  NAND2_X2 u5_mult_82_U10698 ( .A1(u5_mult_82_ab_24__33_), .A2(
        u5_mult_82_SUMB_23__34_), .ZN(u5_mult_82_n5472) );
  NAND2_X1 u5_mult_82_U10697 ( .A1(u5_mult_82_ab_24__33_), .A2(
        u5_mult_82_CARRYB_23__33_), .ZN(u5_mult_82_n5471) );
  NAND3_X4 u5_mult_82_U10696 ( .A1(u5_mult_82_n6358), .A2(u5_mult_82_n6359), 
        .A3(u5_mult_82_n6360), .ZN(u5_mult_82_CARRYB_42__15_) );
  NOR2_X1 u5_mult_82_U10695 ( .A1(u5_mult_82_n6933), .A2(u5_mult_82_net65355), 
        .ZN(u5_mult_82_ab_43__15_) );
  NOR2_X1 u5_mult_82_U10694 ( .A1(u5_mult_82_net64523), .A2(u5_mult_82_n6736), 
        .ZN(u5_mult_82_ab_44__14_) );
  NAND3_X2 u5_mult_82_U10693 ( .A1(u5_mult_82_n5468), .A2(u5_mult_82_n5470), 
        .A3(u5_mult_82_n5469), .ZN(u5_mult_82_CARRYB_43__15_) );
  NAND2_X1 u5_mult_82_U10692 ( .A1(u5_mult_82_ab_43__15_), .A2(
        u5_mult_82_CARRYB_42__15_), .ZN(u5_mult_82_n5470) );
  NAND2_X1 u5_mult_82_U10691 ( .A1(u5_mult_82_ab_43__15_), .A2(
        u5_mult_82_SUMB_42__16_), .ZN(u5_mult_82_n5469) );
  NAND2_X1 u5_mult_82_U10690 ( .A1(u5_mult_82_CARRYB_42__15_), .A2(
        u5_mult_82_SUMB_42__16_), .ZN(u5_mult_82_n5468) );
  XOR2_X2 u5_mult_82_U10689 ( .A(u5_mult_82_SUMB_42__16_), .B(u5_mult_82_n5467), .Z(u5_mult_82_SUMB_43__15_) );
  XOR2_X2 u5_mult_82_U10688 ( .A(u5_mult_82_CARRYB_42__15_), .B(
        u5_mult_82_ab_43__15_), .Z(u5_mult_82_n5467) );
  XOR2_X2 u5_mult_82_U10687 ( .A(u5_mult_82_SUMB_44__14_), .B(u5_mult_82_n5460), .Z(u5_mult_82_SUMB_45__13_) );
  NAND3_X2 u5_mult_82_U10686 ( .A1(u5_mult_82_n5457), .A2(u5_mult_82_n5458), 
        .A3(u5_mult_82_n5459), .ZN(u5_mult_82_CARRYB_44__14_) );
  NAND2_X1 u5_mult_82_U10685 ( .A1(u5_mult_82_CARRYB_43__14_), .A2(
        u5_mult_82_SUMB_43__15_), .ZN(u5_mult_82_n5457) );
  NOR2_X1 u5_mult_82_U10684 ( .A1(u5_mult_82_net64941), .A2(u5_mult_82_n6557), 
        .ZN(u5_mult_82_ab_11__37_) );
  NAND2_X1 u5_mult_82_U10683 ( .A1(u5_mult_82_CARRYB_10__37_), .A2(
        u5_mult_82_SUMB_10__38_), .ZN(u5_mult_82_n5454) );
  NAND3_X2 u5_mult_82_U10682 ( .A1(u5_mult_82_n5451), .A2(u5_mult_82_n5452), 
        .A3(u5_mult_82_n5453), .ZN(u5_mult_82_CARRYB_30__24_) );
  NAND2_X1 u5_mult_82_U10681 ( .A1(u5_mult_82_CARRYB_29__24_), .A2(
        u5_mult_82_SUMB_29__25_), .ZN(u5_mult_82_n5453) );
  NAND2_X1 u5_mult_82_U10680 ( .A1(u5_mult_82_ab_30__24_), .A2(
        u5_mult_82_SUMB_29__25_), .ZN(u5_mult_82_n5452) );
  NAND2_X1 u5_mult_82_U10679 ( .A1(u5_mult_82_ab_30__24_), .A2(
        u5_mult_82_CARRYB_29__24_), .ZN(u5_mult_82_n5451) );
  NAND3_X2 u5_mult_82_U10678 ( .A1(u5_mult_82_n5449), .A2(u5_mult_82_n5448), 
        .A3(u5_mult_82_n5450), .ZN(u5_mult_82_CARRYB_29__25_) );
  NAND2_X1 u5_mult_82_U10677 ( .A1(u5_mult_82_ab_29__25_), .A2(
        u5_mult_82_CARRYB_28__25_), .ZN(u5_mult_82_n5448) );
  XOR2_X2 u5_mult_82_U10676 ( .A(u5_mult_82_n5447), .B(u5_mult_82_SUMB_29__25_), .Z(u5_mult_82_SUMB_30__24_) );
  XOR2_X2 u5_mult_82_U10675 ( .A(u5_mult_82_ab_30__24_), .B(
        u5_mult_82_CARRYB_29__24_), .Z(u5_mult_82_n5447) );
  XOR2_X2 u5_mult_82_U10674 ( .A(u5_mult_82_n5446), .B(u5_mult_82_n1816), .Z(
        u5_mult_82_SUMB_29__25_) );
  XOR2_X2 u5_mult_82_U10673 ( .A(u5_mult_82_ab_29__25_), .B(
        u5_mult_82_CARRYB_28__25_), .Z(u5_mult_82_n5446) );
  NAND3_X2 u5_mult_82_U10672 ( .A1(u5_mult_82_n5443), .A2(u5_mult_82_n5444), 
        .A3(u5_mult_82_n5445), .ZN(u5_mult_82_CARRYB_26__28_) );
  NAND2_X1 u5_mult_82_U10671 ( .A1(u5_mult_82_CARRYB_25__28_), .A2(
        u5_mult_82_SUMB_25__29_), .ZN(u5_mult_82_n5445) );
  NAND2_X1 u5_mult_82_U10670 ( .A1(u5_mult_82_ab_26__28_), .A2(
        u5_mult_82_SUMB_25__29_), .ZN(u5_mult_82_n5444) );
  NAND2_X1 u5_mult_82_U10669 ( .A1(u5_mult_82_ab_26__28_), .A2(
        u5_mult_82_CARRYB_25__28_), .ZN(u5_mult_82_n5443) );
  NAND3_X2 u5_mult_82_U10668 ( .A1(u5_mult_82_n5440), .A2(u5_mult_82_n5441), 
        .A3(u5_mult_82_n5442), .ZN(u5_mult_82_CARRYB_25__29_) );
  NAND2_X1 u5_mult_82_U10667 ( .A1(u5_mult_82_ab_25__29_), .A2(
        u5_mult_82_CARRYB_24__29_), .ZN(u5_mult_82_n5440) );
  INV_X4 u5_mult_82_U10666 ( .A(u5_mult_82_n6782), .ZN(u5_mult_82_n6781) );
  XNOR2_X2 u5_mult_82_U10665 ( .A(u5_mult_82_ab_48__14_), .B(
        u5_mult_82_SUMB_47__15_), .ZN(u5_mult_82_n5438) );
  XNOR2_X2 u5_mult_82_U10664 ( .A(u5_mult_82_n5438), .B(
        u5_mult_82_CARRYB_47__14_), .ZN(u5_mult_82_SUMB_48__14_) );
  XNOR2_X2 u5_mult_82_U10663 ( .A(u5_mult_82_net80099), .B(
        u5_mult_82_CARRYB_42__10_), .ZN(u5_mult_82_net78853) );
  NAND2_X1 u5_mult_82_U10662 ( .A1(u5_mult_82_ab_42__9_), .A2(
        u5_mult_82_CARRYB_41__9_), .ZN(u5_mult_82_n6133) );
  NAND2_X1 u5_mult_82_U10661 ( .A1(u5_mult_82_ab_4__49_), .A2(u5_mult_82_n1468), .ZN(u5_mult_82_n6318) );
  NAND2_X1 u5_mult_82_U10660 ( .A1(u5_mult_82_SUMB_13__44_), .A2(
        u5_mult_82_CARRYB_13__43_), .ZN(u5_mult_82_n5481) );
  NOR2_X1 u5_mult_82_U10659 ( .A1(u5_mult_82_n6896), .A2(u5_mult_82_n6672), 
        .ZN(u5_mult_82_ab_29__21_) );
  NOR2_X1 u5_mult_82_U10658 ( .A1(u5_mult_82_net64559), .A2(
        u5_mult_82_net65443), .ZN(u5_mult_82_ab_38__16_) );
  NAND3_X2 u5_mult_82_U10657 ( .A1(u5_mult_82_n5435), .A2(u5_mult_82_n5436), 
        .A3(u5_mult_82_n5437), .ZN(u5_mult_82_CARRYB_29__21_) );
  NAND3_X2 u5_mult_82_U10656 ( .A1(u5_mult_82_n5432), .A2(u5_mult_82_n5433), 
        .A3(u5_mult_82_n5434), .ZN(u5_mult_82_CARRYB_38__16_) );
  NAND2_X1 u5_mult_82_U10655 ( .A1(u5_mult_82_ab_38__16_), .A2(
        u5_mult_82_CARRYB_37__16_), .ZN(u5_mult_82_n5434) );
  NAND2_X2 u5_mult_82_U10654 ( .A1(u5_mult_82_CARRYB_18__28_), .A2(
        u5_mult_82_SUMB_18__29_), .ZN(u5_mult_82_n5431) );
  NAND2_X2 u5_mult_82_U10653 ( .A1(u5_mult_82_ab_19__28_), .A2(
        u5_mult_82_SUMB_18__29_), .ZN(u5_mult_82_n5430) );
  NAND3_X4 u5_mult_82_U10652 ( .A1(u5_mult_82_n5426), .A2(u5_mult_82_n5427), 
        .A3(u5_mult_82_n5428), .ZN(u5_mult_82_CARRYB_18__29_) );
  NAND2_X2 u5_mult_82_U10651 ( .A1(u5_mult_82_n303), .A2(u5_mult_82_n1680), 
        .ZN(u5_mult_82_n5428) );
  NAND2_X2 u5_mult_82_U10650 ( .A1(u5_mult_82_ab_18__29_), .A2(
        u5_mult_82_n1680), .ZN(u5_mult_82_n5427) );
  NAND3_X2 u5_mult_82_U10649 ( .A1(u5_mult_82_n5423), .A2(u5_mult_82_n5424), 
        .A3(u5_mult_82_n5425), .ZN(u5_mult_82_CARRYB_5__40_) );
  NAND2_X1 u5_mult_82_U10648 ( .A1(u5_mult_82_CARRYB_4__40_), .A2(
        u5_mult_82_SUMB_4__41_), .ZN(u5_mult_82_n5425) );
  NAND2_X1 u5_mult_82_U10647 ( .A1(u5_mult_82_ab_5__40_), .A2(
        u5_mult_82_SUMB_4__41_), .ZN(u5_mult_82_n5424) );
  NAND2_X1 u5_mult_82_U10646 ( .A1(u5_mult_82_ab_5__40_), .A2(
        u5_mult_82_CARRYB_4__40_), .ZN(u5_mult_82_n5423) );
  NAND3_X2 u5_mult_82_U10645 ( .A1(u5_mult_82_n5420), .A2(u5_mult_82_n5421), 
        .A3(u5_mult_82_n5422), .ZN(u5_mult_82_CARRYB_4__41_) );
  NAND2_X2 u5_mult_82_U10644 ( .A1(u5_mult_82_CARRYB_3__41_), .A2(
        u5_mult_82_SUMB_3__42_), .ZN(u5_mult_82_n5422) );
  NAND2_X2 u5_mult_82_U10643 ( .A1(u5_mult_82_ab_4__41_), .A2(
        u5_mult_82_SUMB_3__42_), .ZN(u5_mult_82_n5421) );
  NAND2_X1 u5_mult_82_U10642 ( .A1(u5_mult_82_ab_4__41_), .A2(
        u5_mult_82_CARRYB_3__41_), .ZN(u5_mult_82_n5420) );
  XOR2_X2 u5_mult_82_U10641 ( .A(u5_mult_82_n5419), .B(u5_mult_82_SUMB_4__41_), 
        .Z(u5_mult_82_SUMB_5__40_) );
  XOR2_X2 u5_mult_82_U10640 ( .A(u5_mult_82_ab_5__40_), .B(
        u5_mult_82_CARRYB_4__40_), .Z(u5_mult_82_n5419) );
  XOR2_X2 u5_mult_82_U10639 ( .A(u5_mult_82_n5418), .B(u5_mult_82_SUMB_3__42_), 
        .Z(u5_mult_82_SUMB_4__41_) );
  XOR2_X2 u5_mult_82_U10638 ( .A(u5_mult_82_ab_4__41_), .B(
        u5_mult_82_CARRYB_3__41_), .Z(u5_mult_82_n5418) );
  NAND3_X2 u5_mult_82_U10637 ( .A1(u5_mult_82_n5415), .A2(u5_mult_82_n5416), 
        .A3(u5_mult_82_n5417), .ZN(u5_mult_82_CARRYB_33__19_) );
  NAND2_X1 u5_mult_82_U10636 ( .A1(u5_mult_82_SUMB_32__20_), .A2(
        u5_mult_82_CARRYB_32__19_), .ZN(u5_mult_82_n5417) );
  NAND2_X1 u5_mult_82_U10635 ( .A1(u5_mult_82_ab_33__19_), .A2(
        u5_mult_82_CARRYB_32__19_), .ZN(u5_mult_82_n5415) );
  NAND2_X2 u5_mult_82_U10634 ( .A1(u5_mult_82_CARRYB_31__20_), .A2(
        u5_mult_82_SUMB_31__21_), .ZN(u5_mult_82_n5414) );
  NAND2_X2 u5_mult_82_U10633 ( .A1(u5_mult_82_ab_32__20_), .A2(
        u5_mult_82_SUMB_31__21_), .ZN(u5_mult_82_n5413) );
  NAND2_X1 u5_mult_82_U10632 ( .A1(u5_mult_82_ab_32__20_), .A2(
        u5_mult_82_CARRYB_31__20_), .ZN(u5_mult_82_n5412) );
  XOR2_X2 u5_mult_82_U10631 ( .A(u5_mult_82_n5411), .B(u5_mult_82_SUMB_32__20_), .Z(u5_mult_82_SUMB_33__19_) );
  XOR2_X2 u5_mult_82_U10630 ( .A(u5_mult_82_n5410), .B(u5_mult_82_n86), .Z(
        u5_mult_82_SUMB_32__20_) );
  NAND3_X4 u5_mult_82_U10629 ( .A1(u5_mult_82_n5407), .A2(u5_mult_82_n5408), 
        .A3(u5_mult_82_n5409), .ZN(u5_mult_82_CARRYB_45__11_) );
  NAND2_X2 u5_mult_82_U10628 ( .A1(u5_mult_82_SUMB_44__12_), .A2(
        u5_mult_82_CARRYB_44__11_), .ZN(u5_mult_82_n5409) );
  NAND2_X2 u5_mult_82_U10627 ( .A1(u5_mult_82_ab_45__11_), .A2(
        u5_mult_82_SUMB_44__12_), .ZN(u5_mult_82_n5408) );
  NAND3_X4 u5_mult_82_U10626 ( .A1(u5_mult_82_n5404), .A2(u5_mult_82_n5405), 
        .A3(u5_mult_82_n5406), .ZN(u5_mult_82_CARRYB_44__12_) );
  NAND2_X2 u5_mult_82_U10625 ( .A1(u5_mult_82_ab_44__12_), .A2(
        u5_mult_82_SUMB_43__13_), .ZN(u5_mult_82_n5405) );
  XOR2_X2 u5_mult_82_U10624 ( .A(u5_mult_82_n5403), .B(u5_mult_82_n707), .Z(
        u5_mult_82_SUMB_45__11_) );
  XOR2_X2 u5_mult_82_U10623 ( .A(u5_mult_82_n5402), .B(u5_mult_82_SUMB_43__13_), .Z(u5_mult_82_SUMB_44__12_) );
  NOR2_X1 u5_mult_82_U10622 ( .A1(u5_mult_82_n6818), .A2(u5_mult_82_n6552), 
        .ZN(u5_mult_82_ab_10__42_) );
  NAND2_X1 u5_mult_82_U10621 ( .A1(u5_mult_82_ab_10__42_), .A2(
        u5_mult_82_CARRYB_9__42_), .ZN(u5_mult_82_n5401) );
  NAND2_X2 u5_mult_82_U10620 ( .A1(u5_mult_82_ab_10__42_), .A2(
        u5_mult_82_SUMB_9__43_), .ZN(u5_mult_82_n5400) );
  NAND2_X2 u5_mult_82_U10619 ( .A1(u5_mult_82_ab_11__43_), .A2(
        u5_mult_82_CARRYB_10__43_), .ZN(u5_mult_82_n5396) );
  NAND2_X2 u5_mult_82_U10618 ( .A1(u5_mult_82_ab_10__43_), .A2(
        u5_mult_82_SUMB_9__44_), .ZN(u5_mult_82_n5392) );
  NAND2_X1 u5_mult_82_U10617 ( .A1(u5_mult_82_ab_10__43_), .A2(
        u5_mult_82_CARRYB_9__43_), .ZN(u5_mult_82_n5391) );
  NAND3_X2 u5_mult_82_U10616 ( .A1(u5_mult_82_n5388), .A2(u5_mult_82_n5389), 
        .A3(u5_mult_82_n5390), .ZN(u5_mult_82_CARRYB_15__39_) );
  NAND2_X1 u5_mult_82_U10615 ( .A1(u5_mult_82_CARRYB_14__39_), .A2(
        u5_mult_82_SUMB_14__40_), .ZN(u5_mult_82_n5390) );
  NAND2_X1 u5_mult_82_U10614 ( .A1(u5_mult_82_ab_15__39_), .A2(
        u5_mult_82_SUMB_14__40_), .ZN(u5_mult_82_n5389) );
  NAND2_X1 u5_mult_82_U10613 ( .A1(u5_mult_82_ab_15__39_), .A2(
        u5_mult_82_CARRYB_14__39_), .ZN(u5_mult_82_n5388) );
  NAND2_X2 u5_mult_82_U10612 ( .A1(u5_mult_82_CARRYB_13__40_), .A2(
        u5_mult_82_SUMB_13__41_), .ZN(u5_mult_82_n5387) );
  XOR2_X2 u5_mult_82_U10611 ( .A(u5_mult_82_n5384), .B(u5_mult_82_SUMB_13__41_), .Z(u5_mult_82_SUMB_14__40_) );
  NAND2_X1 u5_mult_82_U10610 ( .A1(u5_mult_82_ab_8__34_), .A2(
        u5_mult_82_SUMB_7__35_), .ZN(u5_mult_82_n5383) );
  NAND3_X2 u5_mult_82_U10609 ( .A1(u5_mult_82_net80185), .A2(u5_mult_82_n5382), 
        .A3(u5_mult_82_net80187), .ZN(u5_mult_82_CARRYB_7__35_) );
  NAND2_X2 u5_mult_82_U10608 ( .A1(u5_mult_82_ab_7__35_), .A2(
        u5_mult_82_SUMB_6__36_), .ZN(u5_mult_82_n5382) );
  XOR2_X2 u5_mult_82_U10607 ( .A(u5_mult_82_net80183), .B(
        u5_mult_82_SUMB_6__36_), .Z(u5_mult_82_SUMB_7__35_) );
  NAND3_X2 u5_mult_82_U10606 ( .A1(u5_mult_82_n5379), .A2(u5_mult_82_n5380), 
        .A3(u5_mult_82_n5381), .ZN(u5_mult_82_CARRYB_25__17_) );
  NAND2_X1 u5_mult_82_U10605 ( .A1(u5_mult_82_ab_25__17_), .A2(
        u5_mult_82_CARRYB_24__17_), .ZN(u5_mult_82_n5379) );
  NAND3_X2 u5_mult_82_U10604 ( .A1(u5_mult_82_n5376), .A2(u5_mult_82_n5377), 
        .A3(u5_mult_82_n5378), .ZN(u5_mult_82_CARRYB_24__18_) );
  NAND2_X2 u5_mult_82_U10603 ( .A1(u5_mult_82_CARRYB_23__18_), .A2(
        u5_mult_82_SUMB_23__19_), .ZN(u5_mult_82_n5378) );
  NAND2_X2 u5_mult_82_U10602 ( .A1(u5_mult_82_ab_24__18_), .A2(
        u5_mult_82_SUMB_23__19_), .ZN(u5_mult_82_n5377) );
  NAND2_X1 u5_mult_82_U10601 ( .A1(u5_mult_82_ab_24__18_), .A2(
        u5_mult_82_CARRYB_23__18_), .ZN(u5_mult_82_n5376) );
  XOR2_X2 u5_mult_82_U10600 ( .A(u5_mult_82_n5375), .B(u5_mult_82_SUMB_24__18_), .Z(u5_mult_82_SUMB_25__17_) );
  XOR2_X2 u5_mult_82_U10599 ( .A(u5_mult_82_ab_25__17_), .B(
        u5_mult_82_CARRYB_24__17_), .Z(u5_mult_82_n5375) );
  XOR2_X2 u5_mult_82_U10598 ( .A(u5_mult_82_n5374), .B(u5_mult_82_SUMB_23__19_), .Z(u5_mult_82_SUMB_24__18_) );
  XOR2_X2 u5_mult_82_U10597 ( .A(u5_mult_82_ab_24__18_), .B(
        u5_mult_82_CARRYB_23__18_), .Z(u5_mult_82_n5374) );
  NAND2_X1 u5_mult_82_U10596 ( .A1(u5_mult_82_ab_43__16_), .A2(
        u5_mult_82_CARRYB_42__16_), .ZN(u5_mult_82_n5883) );
  NOR2_X2 u5_mult_82_U10595 ( .A1(u5_mult_82_n6980), .A2(u5_mult_82_n6568), 
        .ZN(u5_mult_82_ab_12__52_) );
  NOR2_X2 u5_mult_82_U10594 ( .A1(u5_mult_82_n6980), .A2(u5_mult_82_n6560), 
        .ZN(u5_mult_82_ab_11__52_) );
  NOR2_X2 u5_mult_82_U10593 ( .A1(u5_mult_82_n6980), .A2(u5_mult_82_n6553), 
        .ZN(u5_mult_82_ab_10__52_) );
  NOR2_X2 u5_mult_82_U10592 ( .A1(u5_mult_82_n6980), .A2(u5_mult_82_n6547), 
        .ZN(u5_mult_82_ab_9__52_) );
  NOR2_X2 u5_mult_82_U10591 ( .A1(u5_mult_82_n6980), .A2(u5_mult_82_n6538), 
        .ZN(u5_mult_82_ab_8__52_) );
  NOR2_X2 u5_mult_82_U10590 ( .A1(u5_mult_82_n6980), .A2(u5_mult_82_n6531), 
        .ZN(u5_mult_82_ab_7__52_) );
  NOR2_X2 u5_mult_82_U10589 ( .A1(u5_mult_82_n6980), .A2(u5_mult_82_net66023), 
        .ZN(u5_mult_82_ab_6__52_) );
  NOR2_X2 u5_mult_82_U10588 ( .A1(u5_mult_82_n6980), .A2(u5_mult_82_net66041), 
        .ZN(u5_mult_82_ab_5__52_) );
  NOR2_X2 u5_mult_82_U10587 ( .A1(u5_mult_82_n6980), .A2(u5_mult_82_n6515), 
        .ZN(u5_mult_82_ab_3__52_) );
  NOR2_X2 u5_mult_82_U10586 ( .A1(u5_mult_82_n6980), .A2(u5_mult_82_net66091), 
        .ZN(u5_mult_82_ab_2__52_) );
  NOR2_X2 u5_mult_82_U10585 ( .A1(u5_mult_82_n6981), .A2(u5_mult_82_net65681), 
        .ZN(u5_mult_82_ab_25__52_) );
  NOR2_X2 u5_mult_82_U10584 ( .A1(u5_mult_82_n6981), .A2(u5_mult_82_n6645), 
        .ZN(u5_mult_82_ab_24__52_) );
  NOR2_X2 u5_mult_82_U10583 ( .A1(u5_mult_82_n6981), .A2(u5_mult_82_net65717), 
        .ZN(u5_mult_82_ab_23__52_) );
  NOR2_X2 u5_mult_82_U10582 ( .A1(u5_mult_82_n6981), .A2(u5_mult_82_n6638), 
        .ZN(u5_mult_82_ab_22__52_) );
  NOR2_X2 u5_mult_82_U10581 ( .A1(u5_mult_82_n6981), .A2(u5_mult_82_n6631), 
        .ZN(u5_mult_82_ab_21__52_) );
  NOR2_X2 u5_mult_82_U10580 ( .A1(u5_mult_82_n6981), .A2(u5_mult_82_n6624), 
        .ZN(u5_mult_82_ab_20__52_) );
  NOR2_X2 u5_mult_82_U10579 ( .A1(u5_mult_82_n6981), .A2(u5_mult_82_n6617), 
        .ZN(u5_mult_82_ab_19__52_) );
  NOR2_X2 u5_mult_82_U10578 ( .A1(u5_mult_82_n6981), .A2(u5_mult_82_n6611), 
        .ZN(u5_mult_82_ab_18__52_) );
  NOR2_X2 u5_mult_82_U10577 ( .A1(u5_mult_82_n6981), .A2(u5_mult_82_n6604), 
        .ZN(u5_mult_82_ab_17__52_) );
  NOR2_X2 u5_mult_82_U10576 ( .A1(u5_mult_82_n6981), .A2(u5_mult_82_n6597), 
        .ZN(u5_mult_82_ab_16__52_) );
  NOR2_X2 u5_mult_82_U10575 ( .A1(u5_mult_82_n6981), .A2(u5_mult_82_n6589), 
        .ZN(u5_mult_82_ab_15__52_) );
  NOR2_X2 u5_mult_82_U10574 ( .A1(u5_mult_82_n6981), .A2(u5_mult_82_n6581), 
        .ZN(u5_mult_82_ab_14__52_) );
  NOR2_X2 u5_mult_82_U10573 ( .A1(u5_mult_82_n6981), .A2(u5_mult_82_n6574), 
        .ZN(u5_mult_82_ab_13__52_) );
  XNOR2_X2 u5_mult_82_U10572 ( .A(u5_mult_82_CARRYB_40__9_), .B(
        u5_mult_82_ab_41__9_), .ZN(u5_mult_82_n5373) );
  XNOR2_X2 u5_mult_82_U10571 ( .A(u5_mult_82_n1486), .B(u5_mult_82_n5373), 
        .ZN(u5_mult_82_SUMB_41__9_) );
  XNOR2_X2 u5_mult_82_U10570 ( .A(u5_mult_82_CARRYB_20__34_), .B(
        u5_mult_82_ab_21__34_), .ZN(u5_mult_82_n5372) );
  XNOR2_X2 u5_mult_82_U10569 ( .A(u5_mult_82_n1725), .B(u5_mult_82_n5372), 
        .ZN(u5_mult_82_SUMB_21__34_) );
  NOR2_X4 u5_mult_82_U10568 ( .A1(u5_mult_82_n6980), .A2(u5_mult_82_net66111), 
        .ZN(u5_mult_82_ab_1__52_) );
  XNOR2_X2 u5_mult_82_U10567 ( .A(u5_mult_82_ab_4__39_), .B(
        u5_mult_82_CARRYB_3__39_), .ZN(u5_mult_82_n5371) );
  XNOR2_X2 u5_mult_82_U10566 ( .A(u5_mult_82_n5371), .B(u5_mult_82_SUMB_3__40_), .ZN(u5_mult_82_SUMB_4__39_) );
  NOR2_X1 u5_mult_82_U10565 ( .A1(u5_mult_82_n6806), .A2(u5_mult_82_n6537), 
        .ZN(u5_mult_82_ab_8__44_) );
  NOR2_X1 u5_mult_82_U10564 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6594), 
        .ZN(u5_mult_82_ab_16__38_) );
  NOR2_X1 u5_mult_82_U10563 ( .A1(u5_mult_82_n6903), .A2(u5_mult_82_n6735), 
        .ZN(u5_mult_82_ab_44__20_) );
  NAND2_X1 u5_mult_82_U10562 ( .A1(u5_mult_82_ab_12__41_), .A2(
        u5_mult_82_CARRYB_11__41_), .ZN(u5_mult_82_n5368) );
  NAND3_X2 u5_mult_82_U10561 ( .A1(u5_mult_82_n5365), .A2(u5_mult_82_n5366), 
        .A3(u5_mult_82_n5367), .ZN(u5_mult_82_CARRYB_11__42_) );
  NAND2_X2 u5_mult_82_U10560 ( .A1(u5_mult_82_ab_11__42_), .A2(
        u5_mult_82_SUMB_10__43_), .ZN(u5_mult_82_n5366) );
  NAND2_X1 u5_mult_82_U10559 ( .A1(u5_mult_82_ab_11__42_), .A2(
        u5_mult_82_CARRYB_10__42_), .ZN(u5_mult_82_n5365) );
  XOR2_X2 u5_mult_82_U10558 ( .A(u5_mult_82_n5364), .B(u5_mult_82_SUMB_10__43_), .Z(u5_mult_82_SUMB_11__42_) );
  XOR2_X2 u5_mult_82_U10557 ( .A(u5_mult_82_ab_11__42_), .B(
        u5_mult_82_CARRYB_10__42_), .Z(u5_mult_82_n5364) );
  NAND3_X2 u5_mult_82_U10556 ( .A1(u5_mult_82_n5361), .A2(u5_mult_82_n5362), 
        .A3(u5_mult_82_n5363), .ZN(u5_mult_82_CARRYB_8__44_) );
  NAND2_X2 u5_mult_82_U10555 ( .A1(u5_mult_82_ab_8__44_), .A2(
        u5_mult_82_CARRYB_7__44_), .ZN(u5_mult_82_n5363) );
  NAND2_X2 u5_mult_82_U10554 ( .A1(u5_mult_82_ab_8__44_), .A2(
        u5_mult_82_SUMB_7__45_), .ZN(u5_mult_82_n5362) );
  NAND2_X2 u5_mult_82_U10553 ( .A1(u5_mult_82_CARRYB_7__44_), .A2(
        u5_mult_82_SUMB_7__45_), .ZN(u5_mult_82_n5361) );
  NAND3_X2 u5_mult_82_U10552 ( .A1(u5_mult_82_n5358), .A2(u5_mult_82_n5359), 
        .A3(u5_mult_82_n5360), .ZN(u5_mult_82_CARRYB_16__38_) );
  NAND2_X1 u5_mult_82_U10551 ( .A1(u5_mult_82_ab_16__38_), .A2(
        u5_mult_82_CARRYB_15__38_), .ZN(u5_mult_82_n5360) );
  NAND2_X2 u5_mult_82_U10550 ( .A1(u5_mult_82_ab_16__38_), .A2(
        u5_mult_82_SUMB_15__39_), .ZN(u5_mult_82_n5359) );
  NAND2_X1 u5_mult_82_U10549 ( .A1(u5_mult_82_CARRYB_15__38_), .A2(
        u5_mult_82_SUMB_15__39_), .ZN(u5_mult_82_n5358) );
  NAND2_X2 u5_mult_82_U10548 ( .A1(u5_mult_82_ab_15__38_), .A2(
        u5_mult_82_SUMB_14__39_), .ZN(u5_mult_82_n5356) );
  NAND2_X2 u5_mult_82_U10547 ( .A1(u5_mult_82_ab_14__39_), .A2(
        u5_mult_82_SUMB_13__40_), .ZN(u5_mult_82_n5353) );
  XOR2_X2 u5_mult_82_U10546 ( .A(u5_mult_82_n5351), .B(u5_mult_82_n634), .Z(
        u5_mult_82_SUMB_14__39_) );
  NAND2_X1 u5_mult_82_U10545 ( .A1(u5_mult_82_ab_47__17_), .A2(
        u5_mult_82_CARRYB_46__17_), .ZN(u5_mult_82_n5348) );
  NAND2_X2 u5_mult_82_U10544 ( .A1(u5_mult_82_CARRYB_45__18_), .A2(
        u5_mult_82_n1493), .ZN(u5_mult_82_n5347) );
  NAND2_X2 u5_mult_82_U10543 ( .A1(u5_mult_82_ab_46__18_), .A2(
        u5_mult_82_n1493), .ZN(u5_mult_82_n5346) );
  NAND2_X1 u5_mult_82_U10542 ( .A1(u5_mult_82_ab_46__18_), .A2(
        u5_mult_82_CARRYB_45__18_), .ZN(u5_mult_82_n5345) );
  NAND3_X2 u5_mult_82_U10541 ( .A1(u5_mult_82_n5341), .A2(u5_mult_82_n5342), 
        .A3(u5_mult_82_n5343), .ZN(u5_mult_82_CARRYB_44__20_) );
  NAND2_X1 u5_mult_82_U10540 ( .A1(u5_mult_82_ab_44__20_), .A2(
        u5_mult_82_CARRYB_43__20_), .ZN(u5_mult_82_n5343) );
  NAND2_X2 u5_mult_82_U10539 ( .A1(u5_mult_82_ab_44__20_), .A2(
        u5_mult_82_SUMB_43__21_), .ZN(u5_mult_82_n5342) );
  NAND2_X2 u5_mult_82_U10538 ( .A1(u5_mult_82_ab_16__29_), .A2(
        u5_mult_82_CARRYB_15__29_), .ZN(u5_mult_82_n5686) );
  NOR2_X2 u5_mult_82_U10537 ( .A1(u5_mult_82_n6864), .A2(u5_mult_82_n6586), 
        .ZN(u5_mult_82_ab_15__29_) );
  NOR2_X1 u5_mult_82_U10536 ( .A1(u5_mult_82_n6864), .A2(u5_mult_82_n6578), 
        .ZN(u5_mult_82_ab_14__29_) );
  NOR2_X1 u5_mult_82_U10535 ( .A1(u5_mult_82_net64669), .A2(
        u5_mult_82_net65713), .ZN(u5_mult_82_ab_23__22_) );
  NOR2_X1 u5_mult_82_U10534 ( .A1(u5_mult_82_net64433), .A2(u5_mult_82_n6722), 
        .ZN(u5_mult_82_ab_37__9_) );
  NAND2_X1 u5_mult_82_U10533 ( .A1(u5_mult_82_ab_15__29_), .A2(
        u5_mult_82_CARRYB_14__29_), .ZN(u5_mult_82_n5340) );
  NAND2_X2 u5_mult_82_U10532 ( .A1(u5_mult_82_ab_15__29_), .A2(
        u5_mult_82_SUMB_14__30_), .ZN(u5_mult_82_n5339) );
  NAND3_X2 u5_mult_82_U10531 ( .A1(u5_mult_82_net80252), .A2(u5_mult_82_n5337), 
        .A3(u5_mult_82_net80254), .ZN(u5_mult_82_CARRYB_14__29_) );
  NAND2_X2 u5_mult_82_U10530 ( .A1(u5_mult_82_ab_14__29_), .A2(
        u5_mult_82_net83274), .ZN(u5_mult_82_n5337) );
  NAND3_X2 u5_mult_82_U10529 ( .A1(u5_mult_82_n5335), .A2(u5_mult_82_n5334), 
        .A3(u5_mult_82_n5336), .ZN(u5_mult_82_CARRYB_23__22_) );
  NAND2_X1 u5_mult_82_U10528 ( .A1(u5_mult_82_ab_23__22_), .A2(
        u5_mult_82_CARRYB_22__22_), .ZN(u5_mult_82_n5336) );
  NAND2_X2 u5_mult_82_U10527 ( .A1(u5_mult_82_ab_23__22_), .A2(
        u5_mult_82_SUMB_22__23_), .ZN(u5_mult_82_n5335) );
  NAND3_X2 u5_mult_82_U10526 ( .A1(u5_mult_82_n5331), .A2(u5_mult_82_n5332), 
        .A3(u5_mult_82_n5333), .ZN(u5_mult_82_CARRYB_37__9_) );
  NAND2_X1 u5_mult_82_U10525 ( .A1(u5_mult_82_ab_37__9_), .A2(
        u5_mult_82_CARRYB_36__9_), .ZN(u5_mult_82_n5333) );
  NAND2_X2 u5_mult_82_U10524 ( .A1(u5_mult_82_ab_37__9_), .A2(
        u5_mult_82_SUMB_36__10_), .ZN(u5_mult_82_n5332) );
  NAND2_X1 u5_mult_82_U10523 ( .A1(u5_mult_82_CARRYB_36__9_), .A2(
        u5_mult_82_SUMB_36__10_), .ZN(u5_mult_82_n5331) );
  XOR2_X2 u5_mult_82_U10522 ( .A(u5_mult_82_n6205), .B(u5_mult_82_SUMB_47__11_), .Z(u5_mult_82_SUMB_48__10_) );
  NAND2_X1 u5_mult_82_U10521 ( .A1(u5_mult_82_ab_46__14_), .A2(
        u5_mult_82_CARRYB_45__14_), .ZN(u5_mult_82_n5778) );
  NAND2_X1 u5_mult_82_U10520 ( .A1(u5_mult_82_CARRYB_49__11_), .A2(
        u5_mult_82_SUMB_49__12_), .ZN(u5_mult_82_n5993) );
  NAND3_X2 u5_mult_82_U10519 ( .A1(u5_mult_82_n1366), .A2(u5_mult_82_n5328), 
        .A3(u5_mult_82_n5329), .ZN(u5_mult_82_CARRYB_5__36_) );
  NAND2_X1 u5_mult_82_U10518 ( .A1(u5_mult_82_CARRYB_4__36_), .A2(
        u5_mult_82_SUMB_4__37_), .ZN(u5_mult_82_n5329) );
  NAND2_X1 u5_mult_82_U10517 ( .A1(u5_mult_82_ab_5__36_), .A2(
        u5_mult_82_SUMB_4__37_), .ZN(u5_mult_82_n5328) );
  NAND3_X2 u5_mult_82_U10516 ( .A1(u5_mult_82_n5322), .A2(u5_mult_82_n5323), 
        .A3(u5_mult_82_n5324), .ZN(u5_mult_82_CARRYB_17__24_) );
  NAND3_X2 u5_mult_82_U10515 ( .A1(u5_mult_82_n5319), .A2(u5_mult_82_n5320), 
        .A3(u5_mult_82_n5321), .ZN(u5_mult_82_CARRYB_16__25_) );
  NAND2_X2 u5_mult_82_U10514 ( .A1(u5_mult_82_SUMB_15__26_), .A2(
        u5_mult_82_CARRYB_15__25_), .ZN(u5_mult_82_n5321) );
  NAND2_X2 u5_mult_82_U10513 ( .A1(u5_mult_82_ab_16__25_), .A2(
        u5_mult_82_SUMB_15__26_), .ZN(u5_mult_82_n5320) );
  NAND2_X1 u5_mult_82_U10512 ( .A1(u5_mult_82_ab_16__25_), .A2(
        u5_mult_82_CARRYB_15__25_), .ZN(u5_mult_82_n5319) );
  NAND3_X2 u5_mult_82_U10511 ( .A1(u5_mult_82_n5316), .A2(u5_mult_82_n5317), 
        .A3(u5_mult_82_n5318), .ZN(u5_mult_82_CARRYB_12__29_) );
  NAND2_X1 u5_mult_82_U10510 ( .A1(u5_mult_82_CARRYB_11__29_), .A2(
        u5_mult_82_SUMB_11__30_), .ZN(u5_mult_82_n5318) );
  NAND2_X1 u5_mult_82_U10509 ( .A1(u5_mult_82_ab_12__29_), .A2(
        u5_mult_82_SUMB_11__30_), .ZN(u5_mult_82_n5317) );
  NAND2_X1 u5_mult_82_U10508 ( .A1(u5_mult_82_ab_12__29_), .A2(
        u5_mult_82_CARRYB_11__29_), .ZN(u5_mult_82_n5316) );
  NAND2_X2 u5_mult_82_U10507 ( .A1(u5_mult_82_n448), .A2(
        u5_mult_82_CARRYB_10__30_), .ZN(u5_mult_82_n5315) );
  NAND2_X2 u5_mult_82_U10506 ( .A1(u5_mult_82_ab_11__30_), .A2(u5_mult_82_n448), .ZN(u5_mult_82_n5314) );
  NAND2_X1 u5_mult_82_U10505 ( .A1(u5_mult_82_ab_11__30_), .A2(
        u5_mult_82_CARRYB_10__30_), .ZN(u5_mult_82_n5313) );
  XOR2_X2 u5_mult_82_U10504 ( .A(u5_mult_82_n5312), .B(u5_mult_82_n448), .Z(
        u5_mult_82_SUMB_11__30_) );
  XOR2_X2 u5_mult_82_U10503 ( .A(u5_mult_82_ab_11__30_), .B(
        u5_mult_82_CARRYB_10__30_), .Z(u5_mult_82_n5312) );
  NAND3_X2 u5_mult_82_U10502 ( .A1(u5_mult_82_n5309), .A2(u5_mult_82_n5310), 
        .A3(u5_mult_82_n5311), .ZN(u5_mult_82_CARRYB_31__10_) );
  NAND2_X1 u5_mult_82_U10501 ( .A1(u5_mult_82_SUMB_30__11_), .A2(
        u5_mult_82_CARRYB_30__10_), .ZN(u5_mult_82_n5311) );
  NAND2_X1 u5_mult_82_U10500 ( .A1(u5_mult_82_ab_31__10_), .A2(
        u5_mult_82_SUMB_30__11_), .ZN(u5_mult_82_n5310) );
  NAND2_X2 u5_mult_82_U10499 ( .A1(u5_mult_82_CARRYB_29__11_), .A2(
        u5_mult_82_SUMB_29__12_), .ZN(u5_mult_82_n5308) );
  NAND2_X2 u5_mult_82_U10498 ( .A1(u5_mult_82_ab_30__11_), .A2(
        u5_mult_82_SUMB_29__12_), .ZN(u5_mult_82_n5307) );
  XOR2_X2 u5_mult_82_U10497 ( .A(u5_mult_82_n5305), .B(u5_mult_82_SUMB_30__11_), .Z(u5_mult_82_SUMB_31__10_) );
  XOR2_X2 u5_mult_82_U10496 ( .A(u5_mult_82_ab_31__10_), .B(
        u5_mult_82_CARRYB_30__10_), .Z(u5_mult_82_n5305) );
  NAND3_X4 u5_mult_82_U10495 ( .A1(u5_mult_82_n5299), .A2(u5_mult_82_n5300), 
        .A3(u5_mult_82_n5301), .ZN(u5_mult_82_CARRYB_23__18_) );
  NAND2_X2 u5_mult_82_U10494 ( .A1(u5_mult_82_CARRYB_22__18_), .A2(
        u5_mult_82_n743), .ZN(u5_mult_82_n5301) );
  NAND2_X2 u5_mult_82_U10493 ( .A1(u5_mult_82_ab_23__18_), .A2(u5_mult_82_n743), .ZN(u5_mult_82_n5300) );
  NAND2_X1 u5_mult_82_U10492 ( .A1(u5_mult_82_ab_23__18_), .A2(
        u5_mult_82_CARRYB_22__18_), .ZN(u5_mult_82_n5299) );
  XOR2_X2 u5_mult_82_U10491 ( .A(u5_mult_82_n5298), .B(u5_mult_82_n743), .Z(
        u5_mult_82_SUMB_23__18_) );
  XOR2_X2 u5_mult_82_U10490 ( .A(u5_mult_82_ab_23__18_), .B(
        u5_mult_82_CARRYB_22__18_), .Z(u5_mult_82_n5298) );
  XNOR2_X2 u5_mult_82_U10489 ( .A(u5_mult_82_ab_50__11_), .B(
        u5_mult_82_CARRYB_49__11_), .ZN(u5_mult_82_n5297) );
  NOR2_X1 u5_mult_82_U10488 ( .A1(u5_mult_82_net64559), .A2(
        u5_mult_82_net65389), .ZN(u5_mult_82_ab_41__16_) );
  NOR2_X1 u5_mult_82_U10487 ( .A1(u5_mult_82_net64667), .A2(u5_mult_82_n6700), 
        .ZN(u5_mult_82_ab_33__22_) );
  NOR2_X1 u5_mult_82_U10486 ( .A1(u5_mult_82_n6974), .A2(u5_mult_82_net64415), 
        .ZN(u5_mult_82_ab_52__8_) );
  NOR2_X4 u5_mult_82_U10485 ( .A1(u5_mult_82_net64559), .A2(
        u5_mult_82_net65353), .ZN(u5_mult_82_ab_43__16_) );
  NAND3_X2 u5_mult_82_U10484 ( .A1(u5_mult_82_n5294), .A2(u5_mult_82_n5295), 
        .A3(u5_mult_82_n5296), .ZN(u5_mult_82_CARRYB_41__16_) );
  NAND2_X1 u5_mult_82_U10483 ( .A1(u5_mult_82_ab_41__16_), .A2(
        u5_mult_82_CARRYB_40__16_), .ZN(u5_mult_82_n5296) );
  NAND2_X2 u5_mult_82_U10482 ( .A1(u5_mult_82_ab_41__16_), .A2(
        u5_mult_82_SUMB_40__17_), .ZN(u5_mult_82_n5295) );
  XOR2_X2 u5_mult_82_U10481 ( .A(u5_mult_82_SUMB_40__17_), .B(u5_mult_82_n5293), .Z(u5_mult_82_SUMB_41__16_) );
  NAND3_X2 u5_mult_82_U10480 ( .A1(u5_mult_82_n5290), .A2(u5_mult_82_n5291), 
        .A3(u5_mult_82_n5292), .ZN(u5_mult_82_CARRYB_33__22_) );
  NAND2_X1 u5_mult_82_U10479 ( .A1(u5_mult_82_ab_33__22_), .A2(
        u5_mult_82_CARRYB_32__22_), .ZN(u5_mult_82_n5292) );
  NAND2_X1 u5_mult_82_U10478 ( .A1(u5_mult_82_CARRYB_32__22_), .A2(
        u5_mult_82_SUMB_32__23_), .ZN(u5_mult_82_n5290) );
  NAND3_X2 u5_mult_82_U10477 ( .A1(u5_mult_82_n5287), .A2(u5_mult_82_n5288), 
        .A3(u5_mult_82_n5289), .ZN(u5_mult_82_CARRYB_52__8_) );
  NAND2_X2 u5_mult_82_U10476 ( .A1(u5_mult_82_ab_52__8_), .A2(
        u5_mult_82_CARRYB_51__8_), .ZN(u5_mult_82_n5289) );
  NAND2_X1 u5_mult_82_U10475 ( .A1(u5_mult_82_ab_52__8_), .A2(
        u5_mult_82_SUMB_51__9_), .ZN(u5_mult_82_n5288) );
  NAND2_X1 u5_mult_82_U10474 ( .A1(u5_mult_82_CARRYB_51__8_), .A2(
        u5_mult_82_SUMB_51__9_), .ZN(u5_mult_82_n5287) );
  XOR2_X2 u5_mult_82_U10473 ( .A(u5_mult_82_SUMB_51__9_), .B(u5_mult_82_n5286), 
        .Z(u5_mult_82_SUMB_52__8_) );
  XOR2_X2 u5_mult_82_U10472 ( .A(u5_mult_82_CARRYB_51__8_), .B(
        u5_mult_82_ab_52__8_), .Z(u5_mult_82_n5286) );
  INV_X1 u5_mult_82_U10471 ( .A(u5_mult_82_ab_43__16_), .ZN(u5_mult_82_n5283)
         );
  XNOR2_X2 u5_mult_82_U10470 ( .A(u5_mult_82_n5281), .B(
        u5_mult_82_CARRYB_44__11_), .ZN(u5_mult_82_n5403) );
  NOR2_X1 u5_mult_82_U10469 ( .A1(u5_mult_82_n6868), .A2(u5_mult_82_n6727), 
        .ZN(u5_mult_82_ab_39__28_) );
  NOR2_X1 u5_mult_82_U10468 ( .A1(u5_mult_82_n6862), .A2(u5_mult_82_net65441), 
        .ZN(u5_mult_82_ab_38__29_) );
  NAND3_X2 u5_mult_82_U10467 ( .A1(u5_mult_82_n5278), .A2(u5_mult_82_n5279), 
        .A3(u5_mult_82_n5280), .ZN(u5_mult_82_CARRYB_39__28_) );
  NAND2_X2 u5_mult_82_U10466 ( .A1(u5_mult_82_ab_39__28_), .A2(
        u5_mult_82_SUMB_38__29_), .ZN(u5_mult_82_n5279) );
  NAND3_X2 u5_mult_82_U10465 ( .A1(u5_mult_82_n5275), .A2(u5_mult_82_n5276), 
        .A3(u5_mult_82_n5277), .ZN(u5_mult_82_CARRYB_38__29_) );
  NAND2_X1 u5_mult_82_U10464 ( .A1(u5_mult_82_ab_38__29_), .A2(
        u5_mult_82_CARRYB_37__29_), .ZN(u5_mult_82_n5277) );
  NAND2_X1 u5_mult_82_U10463 ( .A1(u5_mult_82_CARRYB_37__29_), .A2(
        u5_mult_82_SUMB_37__30_), .ZN(u5_mult_82_n5275) );
  NAND2_X1 u5_mult_82_U10462 ( .A1(u5_mult_82_ab_44__12_), .A2(
        u5_mult_82_CARRYB_43__12_), .ZN(u5_mult_82_n5404) );
  NAND2_X1 u5_mult_82_U10461 ( .A1(u5_mult_82_ab_16__40_), .A2(
        u5_mult_82_CARRYB_15__40_), .ZN(u5_mult_82_n6287) );
  XNOR2_X2 u5_mult_82_U10460 ( .A(u5_mult_82_CARRYB_24__36_), .B(
        u5_mult_82_ab_25__36_), .ZN(u5_mult_82_n5274) );
  XNOR2_X2 u5_mult_82_U10459 ( .A(u5_mult_82_SUMB_24__37_), .B(
        u5_mult_82_n5274), .ZN(u5_mult_82_SUMB_25__36_) );
  XNOR2_X2 u5_mult_82_U10458 ( .A(u5_mult_82_ab_16__31_), .B(
        u5_mult_82_CARRYB_15__31_), .ZN(u5_mult_82_n5273) );
  XNOR2_X2 u5_mult_82_U10457 ( .A(u5_mult_82_SUMB_15__32_), .B(
        u5_mult_82_n5273), .ZN(u5_mult_82_SUMB_16__31_) );
  NAND3_X2 u5_mult_82_U10456 ( .A1(u5_mult_82_n5961), .A2(u5_mult_82_net79317), 
        .A3(u5_mult_82_net79318), .ZN(u5_mult_82_CARRYB_44__10_) );
  XNOR2_X2 u5_mult_82_U10455 ( .A(u5_mult_82_n5272), .B(
        u5_mult_82_SUMB_10__44_), .ZN(u5_mult_82_n5394) );
  NAND3_X2 u5_mult_82_U10454 ( .A1(u5_mult_82_n5269), .A2(u5_mult_82_n5270), 
        .A3(u5_mult_82_n5271), .ZN(u5_mult_82_CARRYB_23__30_) );
  NAND2_X1 u5_mult_82_U10453 ( .A1(u5_mult_82_CARRYB_22__30_), .A2(
        u5_mult_82_SUMB_22__31_), .ZN(u5_mult_82_n5271) );
  NAND2_X1 u5_mult_82_U10452 ( .A1(u5_mult_82_ab_23__30_), .A2(
        u5_mult_82_SUMB_22__31_), .ZN(u5_mult_82_n5270) );
  NAND2_X1 u5_mult_82_U10451 ( .A1(u5_mult_82_ab_23__30_), .A2(
        u5_mult_82_CARRYB_22__30_), .ZN(u5_mult_82_n5269) );
  NAND3_X2 u5_mult_82_U10450 ( .A1(u5_mult_82_n5267), .A2(u5_mult_82_n5266), 
        .A3(u5_mult_82_n5268), .ZN(u5_mult_82_CARRYB_22__31_) );
  NAND2_X1 u5_mult_82_U10449 ( .A1(u5_mult_82_SUMB_21__32_), .A2(
        u5_mult_82_ab_22__31_), .ZN(u5_mult_82_n5267) );
  NAND2_X1 u5_mult_82_U10448 ( .A1(u5_mult_82_ab_22__31_), .A2(
        u5_mult_82_CARRYB_21__31_), .ZN(u5_mult_82_n5266) );
  XOR2_X2 u5_mult_82_U10447 ( .A(u5_mult_82_n5265), .B(u5_mult_82_SUMB_21__32_), .Z(u5_mult_82_SUMB_22__31_) );
  NAND2_X1 u5_mult_82_U10446 ( .A1(u5_mult_82_ab_49__8_), .A2(
        u5_mult_82_CARRYB_48__8_), .ZN(u5_mult_82_n5262) );
  NAND2_X2 u5_mult_82_U10445 ( .A1(u5_mult_82_CARRYB_47__9_), .A2(
        u5_mult_82_SUMB_47__10_), .ZN(u5_mult_82_n5261) );
  NAND2_X2 u5_mult_82_U10444 ( .A1(u5_mult_82_ab_48__9_), .A2(
        u5_mult_82_SUMB_47__10_), .ZN(u5_mult_82_n5260) );
  XNOR2_X2 u5_mult_82_U10443 ( .A(u5_mult_82_CARRYB_23__36_), .B(
        u5_mult_82_ab_24__36_), .ZN(u5_mult_82_n5258) );
  XNOR2_X2 u5_mult_82_U10442 ( .A(u5_mult_82_SUMB_23__37_), .B(
        u5_mult_82_n5258), .ZN(u5_mult_82_SUMB_24__36_) );
  NAND2_X2 u5_mult_82_U10441 ( .A1(u5_mult_82_CARRYB_31__31_), .A2(
        u5_mult_82_n1800), .ZN(u5_mult_82_n5870) );
  XNOR2_X2 u5_mult_82_U10440 ( .A(u5_mult_82_ab_51__7_), .B(
        u5_mult_82_CARRYB_50__7_), .ZN(u5_mult_82_n5256) );
  INV_X1 u5_mult_82_U10439 ( .A(u5_mult_82_SUMB_17__47_), .ZN(u5_mult_82_n5253) );
  NAND2_X2 u5_mult_82_U10438 ( .A1(u5_mult_82_n5252), .A2(u5_mult_82_n5253), 
        .ZN(u5_mult_82_n5255) );
  NOR2_X1 u5_mult_82_U10437 ( .A1(u5_mult_82_n6868), .A2(u5_mult_82_n6693), 
        .ZN(u5_mult_82_ab_32__28_) );
  NAND3_X2 u5_mult_82_U10436 ( .A1(u5_mult_82_n5249), .A2(u5_mult_82_n5250), 
        .A3(u5_mult_82_n5251), .ZN(u5_mult_82_CARRYB_32__28_) );
  NAND2_X1 u5_mult_82_U10435 ( .A1(u5_mult_82_ab_32__28_), .A2(
        u5_mult_82_CARRYB_31__28_), .ZN(u5_mult_82_n5251) );
  NAND2_X1 u5_mult_82_U10434 ( .A1(u5_mult_82_CARRYB_31__28_), .A2(
        u5_mult_82_SUMB_31__29_), .ZN(u5_mult_82_n5249) );
  INV_X4 u5_mult_82_U10433 ( .A(u5_mult_82_n5247), .ZN(u5_mult_82_n5248) );
  XNOR2_X2 u5_mult_82_U10432 ( .A(u5_mult_82_n5246), .B(
        u5_mult_82_CARRYB_43__12_), .ZN(u5_mult_82_n5402) );
  NOR2_X2 u5_mult_82_U10431 ( .A1(u5_mult_82_net64361), .A2(
        u5_mult_82_net65355), .ZN(u5_mult_82_ab_43__5_) );
  NOR2_X1 u5_mult_82_U10430 ( .A1(u5_mult_82_n6952), .A2(u5_mult_82_net65189), 
        .ZN(u5_mult_82_ab_51__3_) );
  NAND3_X2 u5_mult_82_U10429 ( .A1(u5_mult_82_n5240), .A2(u5_mult_82_n5241), 
        .A3(u5_mult_82_n5242), .ZN(u5_mult_82_CARRYB_51__3_) );
  NAND2_X1 u5_mult_82_U10428 ( .A1(u5_mult_82_ab_51__3_), .A2(
        u5_mult_82_SUMB_50__4_), .ZN(u5_mult_82_n5242) );
  NAND3_X4 u5_mult_82_U10427 ( .A1(u5_mult_82_n5237), .A2(u5_mult_82_n5238), 
        .A3(u5_mult_82_n5239), .ZN(u5_mult_82_CARRYB_4__36_) );
  NAND2_X2 u5_mult_82_U10426 ( .A1(u5_mult_82_SUMB_3__37_), .A2(
        u5_mult_82_CARRYB_3__36_), .ZN(u5_mult_82_n5239) );
  NAND2_X2 u5_mult_82_U10425 ( .A1(u5_mult_82_SUMB_3__37_), .A2(
        u5_mult_82_ab_4__36_), .ZN(u5_mult_82_n5238) );
  NAND2_X1 u5_mult_82_U10424 ( .A1(u5_mult_82_ab_4__36_), .A2(
        u5_mult_82_CARRYB_3__36_), .ZN(u5_mult_82_n5237) );
  NAND3_X2 u5_mult_82_U10423 ( .A1(u5_mult_82_n5234), .A2(u5_mult_82_n5235), 
        .A3(u5_mult_82_n5236), .ZN(u5_mult_82_CARRYB_21__19_) );
  NAND2_X1 u5_mult_82_U10422 ( .A1(u5_mult_82_CARRYB_20__19_), .A2(
        u5_mult_82_SUMB_20__20_), .ZN(u5_mult_82_n5236) );
  NAND2_X1 u5_mult_82_U10421 ( .A1(u5_mult_82_ab_21__19_), .A2(
        u5_mult_82_SUMB_20__20_), .ZN(u5_mult_82_n5235) );
  NAND2_X1 u5_mult_82_U10420 ( .A1(u5_mult_82_ab_21__19_), .A2(
        u5_mult_82_CARRYB_20__19_), .ZN(u5_mult_82_n5234) );
  NAND2_X2 u5_mult_82_U10419 ( .A1(u5_mult_82_CARRYB_19__20_), .A2(
        u5_mult_82_SUMB_19__21_), .ZN(u5_mult_82_n5233) );
  NAND2_X2 u5_mult_82_U10418 ( .A1(u5_mult_82_ab_20__20_), .A2(
        u5_mult_82_SUMB_19__21_), .ZN(u5_mult_82_n5232) );
  NAND2_X1 u5_mult_82_U10417 ( .A1(u5_mult_82_ab_20__20_), .A2(
        u5_mult_82_CARRYB_19__20_), .ZN(u5_mult_82_n5231) );
  XOR2_X2 u5_mult_82_U10416 ( .A(u5_mult_82_n5230), .B(u5_mult_82_SUMB_20__20_), .Z(u5_mult_82_SUMB_21__19_) );
  XOR2_X2 u5_mult_82_U10415 ( .A(u5_mult_82_ab_21__19_), .B(
        u5_mult_82_CARRYB_20__19_), .Z(u5_mult_82_n5230) );
  XOR2_X2 u5_mult_82_U10414 ( .A(u5_mult_82_n5229), .B(u5_mult_82_SUMB_19__21_), .Z(u5_mult_82_SUMB_20__20_) );
  XOR2_X2 u5_mult_82_U10413 ( .A(u5_mult_82_ab_20__20_), .B(
        u5_mult_82_CARRYB_19__20_), .Z(u5_mult_82_n5229) );
  NAND3_X2 u5_mult_82_U10412 ( .A1(u5_mult_82_n5223), .A2(u5_mult_82_n5224), 
        .A3(u5_mult_82_n5225), .ZN(u5_mult_82_CARRYB_32__12_) );
  NAND2_X2 u5_mult_82_U10411 ( .A1(u5_mult_82_CARRYB_31__12_), .A2(
        u5_mult_82_SUMB_31__13_), .ZN(u5_mult_82_n5225) );
  NAND2_X2 u5_mult_82_U10410 ( .A1(u5_mult_82_ab_32__12_), .A2(
        u5_mult_82_SUMB_31__13_), .ZN(u5_mult_82_n5224) );
  NAND2_X1 u5_mult_82_U10409 ( .A1(u5_mult_82_ab_32__12_), .A2(
        u5_mult_82_CARRYB_31__12_), .ZN(u5_mult_82_n5223) );
  XNOR2_X2 u5_mult_82_U10408 ( .A(u5_mult_82_CARRYB_16__35_), .B(
        u5_mult_82_n5221), .ZN(u5_mult_82_n6186) );
  XNOR2_X2 u5_mult_82_U10407 ( .A(u5_mult_82_ab_13__37_), .B(
        u5_mult_82_CARRYB_12__37_), .ZN(u5_mult_82_n5220) );
  XNOR2_X2 u5_mult_82_U10406 ( .A(u5_mult_82_n5220), .B(
        u5_mult_82_SUMB_12__38_), .ZN(u5_mult_82_SUMB_13__37_) );
  INV_X8 u5_mult_82_U10405 ( .A(n4762), .ZN(u5_mult_82_n7010) );
  XNOR2_X2 u5_mult_82_U10404 ( .A(u5_mult_82_CARRYB_14__29_), .B(
        u5_mult_82_n5219), .ZN(u5_mult_82_net80255) );
  NOR2_X1 u5_mult_82_U10403 ( .A1(u5_mult_82_n6892), .A2(u5_mult_82_n6629), 
        .ZN(u5_mult_82_ab_21__24_) );
  NAND2_X2 u5_mult_82_U10402 ( .A1(u5_mult_82_ab_34__13_), .A2(
        u5_mult_82_CARRYB_33__13_), .ZN(u5_mult_82_n5921) );
  NOR2_X2 u5_mult_82_U10401 ( .A1(u5_mult_82_net64505), .A2(u5_mult_82_n6701), 
        .ZN(u5_mult_82_ab_33__13_) );
  NAND2_X1 u5_mult_82_U10400 ( .A1(u5_mult_82_ab_21__24_), .A2(
        u5_mult_82_CARRYB_20__24_), .ZN(u5_mult_82_n5218) );
  NAND2_X2 u5_mult_82_U10399 ( .A1(u5_mult_82_CARRYB_17__27_), .A2(
        u5_mult_82_SUMB_17__28_), .ZN(u5_mult_82_n5217) );
  NAND2_X2 u5_mult_82_U10398 ( .A1(u5_mult_82_ab_18__27_), .A2(
        u5_mult_82_SUMB_17__28_), .ZN(u5_mult_82_n5216) );
  NAND2_X1 u5_mult_82_U10397 ( .A1(u5_mult_82_ab_18__27_), .A2(
        u5_mult_82_CARRYB_17__27_), .ZN(u5_mult_82_n5215) );
  NAND3_X4 u5_mult_82_U10396 ( .A1(u5_mult_82_net80535), .A2(u5_mult_82_n5214), 
        .A3(u5_mult_82_net80537), .ZN(u5_mult_82_CARRYB_17__28_) );
  NAND2_X2 u5_mult_82_U10395 ( .A1(u5_mult_82_ab_17__28_), .A2(
        u5_mult_82_SUMB_16__29_), .ZN(u5_mult_82_n5214) );
  NAND3_X4 u5_mult_82_U10394 ( .A1(u5_mult_82_n5211), .A2(u5_mult_82_n5212), 
        .A3(u5_mult_82_n5213), .ZN(u5_mult_82_CARRYB_33__13_) );
  NAND2_X2 u5_mult_82_U10393 ( .A1(u5_mult_82_ab_33__13_), .A2(
        u5_mult_82_SUMB_32__14_), .ZN(u5_mult_82_n5212) );
  XOR2_X2 u5_mult_82_U10392 ( .A(u5_mult_82_SUMB_32__14_), .B(u5_mult_82_n5210), .Z(u5_mult_82_SUMB_33__13_) );
  NAND3_X2 u5_mult_82_U10391 ( .A1(u5_mult_82_n5207), .A2(u5_mult_82_n5208), 
        .A3(u5_mult_82_n5209), .ZN(u5_mult_82_CARRYB_39__8_) );
  NAND2_X1 u5_mult_82_U10390 ( .A1(u5_mult_82_CARRYB_38__8_), .A2(
        u5_mult_82_SUMB_38__9_), .ZN(u5_mult_82_n5209) );
  NAND2_X1 u5_mult_82_U10389 ( .A1(u5_mult_82_ab_39__8_), .A2(
        u5_mult_82_SUMB_38__9_), .ZN(u5_mult_82_n5208) );
  NAND2_X1 u5_mult_82_U10388 ( .A1(u5_mult_82_ab_39__8_), .A2(
        u5_mult_82_CARRYB_38__8_), .ZN(u5_mult_82_n5207) );
  NAND2_X2 u5_mult_82_U10387 ( .A1(u5_mult_82_CARRYB_37__9_), .A2(
        u5_mult_82_SUMB_37__10_), .ZN(u5_mult_82_n5206) );
  NAND2_X2 u5_mult_82_U10386 ( .A1(u5_mult_82_ab_38__9_), .A2(
        u5_mult_82_SUMB_37__10_), .ZN(u5_mult_82_n5205) );
  NAND2_X1 u5_mult_82_U10385 ( .A1(u5_mult_82_ab_38__9_), .A2(
        u5_mult_82_CARRYB_37__9_), .ZN(u5_mult_82_n5204) );
  XOR2_X2 u5_mult_82_U10384 ( .A(u5_mult_82_n5202), .B(u5_mult_82_n1854), .Z(
        u5_mult_82_SUMB_38__9_) );
  XOR2_X2 u5_mult_82_U10383 ( .A(u5_mult_82_ab_38__9_), .B(
        u5_mult_82_CARRYB_37__9_), .Z(u5_mult_82_n5202) );
  NAND3_X2 u5_mult_82_U10382 ( .A1(u5_mult_82_n6333), .A2(u5_mult_82_n6334), 
        .A3(u5_mult_82_n6335), .ZN(u5_mult_82_CARRYB_34__20_) );
  NOR2_X2 u5_mult_82_U10381 ( .A1(u5_mult_82_net64923), .A2(u5_mult_82_n6571), 
        .ZN(u5_mult_82_ab_13__36_) );
  NOR2_X1 u5_mult_82_U10380 ( .A1(u5_mult_82_net64923), .A2(u5_mult_82_n6578), 
        .ZN(u5_mult_82_ab_14__36_) );
  NOR2_X1 u5_mult_82_U10379 ( .A1(u5_mult_82_n6904), .A2(u5_mult_82_n6721), 
        .ZN(u5_mult_82_ab_37__20_) );
  NAND3_X2 u5_mult_82_U10378 ( .A1(u5_mult_82_n5198), .A2(u5_mult_82_n5199), 
        .A3(u5_mult_82_n5200), .ZN(u5_mult_82_CARRYB_13__36_) );
  NAND2_X1 u5_mult_82_U10377 ( .A1(u5_mult_82_ab_13__36_), .A2(
        u5_mult_82_SUMB_12__37_), .ZN(u5_mult_82_n5199) );
  NAND2_X1 u5_mult_82_U10376 ( .A1(u5_mult_82_CARRYB_12__36_), .A2(
        u5_mult_82_SUMB_12__37_), .ZN(u5_mult_82_n5198) );
  NAND3_X2 u5_mult_82_U10375 ( .A1(u5_mult_82_n5194), .A2(u5_mult_82_n5195), 
        .A3(u5_mult_82_n5196), .ZN(u5_mult_82_CARRYB_14__36_) );
  NAND2_X2 u5_mult_82_U10374 ( .A1(u5_mult_82_ab_14__36_), .A2(
        u5_mult_82_SUMB_13__37_), .ZN(u5_mult_82_n5196) );
  NAND2_X2 u5_mult_82_U10373 ( .A1(u5_mult_82_ab_14__36_), .A2(
        u5_mult_82_CARRYB_13__36_), .ZN(u5_mult_82_n5195) );
  NAND2_X1 u5_mult_82_U10372 ( .A1(u5_mult_82_SUMB_13__37_), .A2(
        u5_mult_82_CARRYB_13__36_), .ZN(u5_mult_82_n5194) );
  NAND3_X2 u5_mult_82_U10371 ( .A1(u5_mult_82_n5191), .A2(u5_mult_82_n5192), 
        .A3(u5_mult_82_n5193), .ZN(u5_mult_82_CARRYB_40__17_) );
  NAND2_X1 u5_mult_82_U10370 ( .A1(u5_mult_82_ab_40__17_), .A2(
        u5_mult_82_CARRYB_39__17_), .ZN(u5_mult_82_n5191) );
  NAND2_X2 u5_mult_82_U10369 ( .A1(u5_mult_82_ab_39__18_), .A2(u5_mult_82_n735), .ZN(u5_mult_82_n5189) );
  NAND2_X1 u5_mult_82_U10368 ( .A1(u5_mult_82_ab_39__18_), .A2(
        u5_mult_82_CARRYB_38__18_), .ZN(u5_mult_82_n5188) );
  NAND3_X2 u5_mult_82_U10367 ( .A1(u5_mult_82_n5185), .A2(u5_mult_82_n5186), 
        .A3(u5_mult_82_n5187), .ZN(u5_mult_82_CARRYB_37__20_) );
  NAND2_X1 u5_mult_82_U10366 ( .A1(u5_mult_82_ab_37__20_), .A2(
        u5_mult_82_CARRYB_36__20_), .ZN(u5_mult_82_n5187) );
  NAND2_X1 u5_mult_82_U10365 ( .A1(u5_mult_82_CARRYB_36__20_), .A2(
        u5_mult_82_SUMB_36__21_), .ZN(u5_mult_82_n5185) );
  INV_X2 u5_mult_82_U10364 ( .A(u5_mult_82_SUMB_11__39_), .ZN(u5_mult_82_n5183) );
  NAND2_X2 u5_mult_82_U10363 ( .A1(u5_mult_82_ab_9__45_), .A2(
        u5_mult_82_CARRYB_8__45_), .ZN(u5_mult_82_n6352) );
  NOR2_X2 u5_mult_82_U10362 ( .A1(u5_mult_82_n6799), .A2(u5_mult_82_n6537), 
        .ZN(u5_mult_82_ab_8__45_) );
  NOR2_X1 u5_mult_82_U10361 ( .A1(u5_mult_82_n6850), .A2(u5_mult_82_n6678), 
        .ZN(u5_mult_82_ab_30__31_) );
  NAND3_X2 u5_mult_82_U10360 ( .A1(u5_mult_82_n5180), .A2(u5_mult_82_n5181), 
        .A3(u5_mult_82_n5182), .ZN(u5_mult_82_CARRYB_44__21_) );
  NAND2_X1 u5_mult_82_U10359 ( .A1(u5_mult_82_ab_44__21_), .A2(
        u5_mult_82_CARRYB_43__21_), .ZN(u5_mult_82_n5181) );
  NAND3_X2 u5_mult_82_U10358 ( .A1(u5_mult_82_n5177), .A2(u5_mult_82_n5178), 
        .A3(u5_mult_82_n5179), .ZN(u5_mult_82_CARRYB_43__21_) );
  NAND2_X1 u5_mult_82_U10357 ( .A1(u5_mult_82_CARRYB_42__21_), .A2(
        u5_mult_82_SUMB_42__22_), .ZN(u5_mult_82_n5179) );
  NAND2_X1 u5_mult_82_U10356 ( .A1(u5_mult_82_ab_43__21_), .A2(
        u5_mult_82_SUMB_42__22_), .ZN(u5_mult_82_n5178) );
  NAND2_X1 u5_mult_82_U10355 ( .A1(u5_mult_82_ab_43__21_), .A2(
        u5_mult_82_CARRYB_42__21_), .ZN(u5_mult_82_n5177) );
  XOR2_X2 u5_mult_82_U10354 ( .A(u5_mult_82_n5176), .B(u5_mult_82_SUMB_42__22_), .Z(u5_mult_82_SUMB_43__21_) );
  NAND3_X4 u5_mult_82_U10353 ( .A1(u5_mult_82_n5173), .A2(u5_mult_82_n5174), 
        .A3(u5_mult_82_n5175), .ZN(u5_mult_82_CARRYB_13__41_) );
  NAND2_X1 u5_mult_82_U10352 ( .A1(u5_mult_82_ab_13__41_), .A2(
        u5_mult_82_CARRYB_12__41_), .ZN(u5_mult_82_n5173) );
  NAND2_X2 u5_mult_82_U10351 ( .A1(u5_mult_82_CARRYB_11__42_), .A2(
        u5_mult_82_n1505), .ZN(u5_mult_82_n5172) );
  NAND2_X2 u5_mult_82_U10350 ( .A1(u5_mult_82_ab_12__42_), .A2(
        u5_mult_82_n1505), .ZN(u5_mult_82_n5171) );
  NAND2_X2 u5_mult_82_U10349 ( .A1(u5_mult_82_ab_12__42_), .A2(
        u5_mult_82_CARRYB_11__42_), .ZN(u5_mult_82_n5170) );
  XOR2_X2 u5_mult_82_U10348 ( .A(u5_mult_82_n5169), .B(u5_mult_82_SUMB_12__42_), .Z(u5_mult_82_SUMB_13__41_) );
  XOR2_X2 u5_mult_82_U10347 ( .A(u5_mult_82_ab_13__41_), .B(
        u5_mult_82_CARRYB_12__41_), .Z(u5_mult_82_n5169) );
  XOR2_X2 u5_mult_82_U10346 ( .A(u5_mult_82_n5168), .B(u5_mult_82_n1505), .Z(
        u5_mult_82_SUMB_12__42_) );
  XOR2_X2 u5_mult_82_U10345 ( .A(u5_mult_82_ab_12__42_), .B(
        u5_mult_82_CARRYB_11__42_), .Z(u5_mult_82_n5168) );
  NAND2_X1 u5_mult_82_U10344 ( .A1(u5_mult_82_ab_8__45_), .A2(
        u5_mult_82_SUMB_7__46_), .ZN(u5_mult_82_n5167) );
  NAND2_X2 u5_mult_82_U10343 ( .A1(u5_mult_82_ab_8__45_), .A2(
        u5_mult_82_CARRYB_7__45_), .ZN(u5_mult_82_n5166) );
  NAND2_X1 u5_mult_82_U10342 ( .A1(u5_mult_82_SUMB_7__46_), .A2(
        u5_mult_82_CARRYB_7__45_), .ZN(u5_mult_82_n5165) );
  NAND3_X2 u5_mult_82_U10341 ( .A1(u5_mult_82_n5162), .A2(u5_mult_82_n5163), 
        .A3(u5_mult_82_n5164), .ZN(u5_mult_82_CARRYB_30__31_) );
  NAND2_X2 u5_mult_82_U10340 ( .A1(u5_mult_82_ab_30__31_), .A2(
        u5_mult_82_CARRYB_29__31_), .ZN(u5_mult_82_n5164) );
  NOR2_X1 u5_mult_82_U10339 ( .A1(u5_mult_82_n6953), .A2(u5_mult_82_net65393), 
        .ZN(u5_mult_82_ab_41__3_) );
  NOR2_X1 u5_mult_82_U10338 ( .A1(u5_mult_82_n6882), .A2(u5_mult_82_n6572), 
        .ZN(u5_mult_82_ab_13__26_) );
  NAND3_X2 u5_mult_82_U10337 ( .A1(u5_mult_82_n5158), .A2(u5_mult_82_n5159), 
        .A3(u5_mult_82_n5160), .ZN(u5_mult_82_CARRYB_41__3_) );
  NAND2_X1 u5_mult_82_U10336 ( .A1(u5_mult_82_ab_41__3_), .A2(
        u5_mult_82_CARRYB_40__3_), .ZN(u5_mult_82_n5160) );
  NAND2_X2 u5_mult_82_U10335 ( .A1(u5_mult_82_ab_41__3_), .A2(
        u5_mult_82_SUMB_40__4_), .ZN(u5_mult_82_n5159) );
  XOR2_X2 u5_mult_82_U10334 ( .A(u5_mult_82_CARRYB_40__3_), .B(
        u5_mult_82_ab_41__3_), .Z(u5_mult_82_n5157) );
  NAND3_X2 u5_mult_82_U10333 ( .A1(u5_mult_82_n5156), .A2(u5_mult_82_net80618), 
        .A3(u5_mult_82_net80619), .ZN(u5_mult_82_CARRYB_4__35_) );
  NAND3_X2 u5_mult_82_U10332 ( .A1(u5_mult_82_n5152), .A2(u5_mult_82_n5153), 
        .A3(u5_mult_82_n5154), .ZN(u5_mult_82_CARRYB_15__24_) );
  NAND2_X1 u5_mult_82_U10331 ( .A1(u5_mult_82_CARRYB_14__24_), .A2(
        u5_mult_82_SUMB_14__25_), .ZN(u5_mult_82_n5154) );
  NAND2_X1 u5_mult_82_U10330 ( .A1(u5_mult_82_ab_15__24_), .A2(
        u5_mult_82_SUMB_14__25_), .ZN(u5_mult_82_n5153) );
  NAND2_X1 u5_mult_82_U10329 ( .A1(u5_mult_82_ab_15__24_), .A2(
        u5_mult_82_CARRYB_14__24_), .ZN(u5_mult_82_n5152) );
  NAND3_X2 u5_mult_82_U10328 ( .A1(u5_mult_82_n5149), .A2(u5_mult_82_n5150), 
        .A3(u5_mult_82_n5151), .ZN(u5_mult_82_CARRYB_14__25_) );
  NAND2_X2 u5_mult_82_U10327 ( .A1(u5_mult_82_ab_14__25_), .A2(
        u5_mult_82_SUMB_13__26_), .ZN(u5_mult_82_n5150) );
  NAND2_X1 u5_mult_82_U10326 ( .A1(u5_mult_82_ab_14__25_), .A2(
        u5_mult_82_CARRYB_13__25_), .ZN(u5_mult_82_n5149) );
  XOR2_X2 u5_mult_82_U10325 ( .A(u5_mult_82_n5148), .B(u5_mult_82_SUMB_13__26_), .Z(u5_mult_82_SUMB_14__25_) );
  XOR2_X2 u5_mult_82_U10324 ( .A(u5_mult_82_ab_14__25_), .B(
        u5_mult_82_CARRYB_13__25_), .Z(u5_mult_82_n5148) );
  NAND3_X2 u5_mult_82_U10323 ( .A1(u5_mult_82_n5145), .A2(u5_mult_82_n5146), 
        .A3(u5_mult_82_n5147), .ZN(u5_mult_82_CARRYB_13__26_) );
  NAND2_X1 u5_mult_82_U10322 ( .A1(u5_mult_82_ab_13__26_), .A2(
        u5_mult_82_CARRYB_12__26_), .ZN(u5_mult_82_n5147) );
  NAND2_X2 u5_mult_82_U10321 ( .A1(u5_mult_82_ab_13__26_), .A2(
        u5_mult_82_n1530), .ZN(u5_mult_82_n5146) );
  NAND2_X2 u5_mult_82_U10320 ( .A1(u5_mult_82_CARRYB_12__26_), .A2(
        u5_mult_82_n1530), .ZN(u5_mult_82_n5145) );
  XOR2_X2 u5_mult_82_U10319 ( .A(u5_mult_82_n1530), .B(u5_mult_82_n5144), .Z(
        u5_mult_82_SUMB_13__26_) );
  XOR2_X2 u5_mult_82_U10318 ( .A(u5_mult_82_CARRYB_12__26_), .B(
        u5_mult_82_ab_13__26_), .Z(u5_mult_82_n5144) );
  XNOR2_X2 u5_mult_82_U10317 ( .A(u5_mult_82_n5143), .B(
        u5_mult_82_CARRYB_32__19_), .ZN(u5_mult_82_n5411) );
  XNOR2_X2 u5_mult_82_U10316 ( .A(u5_mult_82_ab_44__9_), .B(
        u5_mult_82_CARRYB_43__9_), .ZN(u5_mult_82_n5142) );
  NOR2_X1 u5_mult_82_U10315 ( .A1(u5_mult_82_n6897), .A2(u5_mult_82_n6657), 
        .ZN(u5_mult_82_ab_27__21_) );
  NAND3_X2 u5_mult_82_U10314 ( .A1(u5_mult_82_net80645), .A2(u5_mult_82_n5141), 
        .A3(u5_mult_82_net80647), .ZN(u5_mult_82_CARRYB_27__21_) );
  NAND2_X1 u5_mult_82_U10313 ( .A1(u5_mult_82_ab_27__21_), .A2(
        u5_mult_82_SUMB_26__22_), .ZN(u5_mult_82_n5141) );
  NAND2_X1 u5_mult_82_U10312 ( .A1(u5_mult_82_CARRYB_22__25_), .A2(
        u5_mult_82_SUMB_22__26_), .ZN(u5_mult_82_n5140) );
  NAND2_X1 u5_mult_82_U10311 ( .A1(u5_mult_82_ab_23__25_), .A2(
        u5_mult_82_SUMB_22__26_), .ZN(u5_mult_82_n5139) );
  NAND2_X1 u5_mult_82_U10310 ( .A1(u5_mult_82_ab_23__25_), .A2(
        u5_mult_82_CARRYB_22__25_), .ZN(u5_mult_82_n5138) );
  NAND3_X2 u5_mult_82_U10309 ( .A1(u5_mult_82_n5137), .A2(u5_mult_82_n5135), 
        .A3(u5_mult_82_n5136), .ZN(u5_mult_82_CARRYB_22__26_) );
  NAND2_X1 u5_mult_82_U10308 ( .A1(u5_mult_82_CARRYB_21__26_), .A2(
        u5_mult_82_SUMB_21__27_), .ZN(u5_mult_82_n5137) );
  NAND2_X1 u5_mult_82_U10307 ( .A1(u5_mult_82_ab_22__26_), .A2(
        u5_mult_82_SUMB_21__27_), .ZN(u5_mult_82_n5136) );
  NAND2_X1 u5_mult_82_U10306 ( .A1(u5_mult_82_ab_22__26_), .A2(
        u5_mult_82_CARRYB_21__26_), .ZN(u5_mult_82_n5135) );
  XOR2_X2 u5_mult_82_U10305 ( .A(u5_mult_82_n5134), .B(u5_mult_82_SUMB_21__27_), .Z(u5_mult_82_SUMB_22__26_) );
  XOR2_X2 u5_mult_82_U10304 ( .A(u5_mult_82_ab_22__26_), .B(
        u5_mult_82_CARRYB_21__26_), .Z(u5_mult_82_n5134) );
  NAND3_X2 u5_mult_82_U10303 ( .A1(u5_mult_82_n5128), .A2(u5_mult_82_n5129), 
        .A3(u5_mult_82_n5130), .ZN(u5_mult_82_CARRYB_38__12_) );
  NAND2_X1 u5_mult_82_U10302 ( .A1(u5_mult_82_ab_38__12_), .A2(
        u5_mult_82_CARRYB_37__12_), .ZN(u5_mult_82_n5128) );
  NAND3_X2 u5_mult_82_U10301 ( .A1(u5_mult_82_n5124), .A2(u5_mult_82_n5125), 
        .A3(u5_mult_82_n5126), .ZN(u5_mult_82_CARRYB_37__35_) );
  NAND2_X1 u5_mult_82_U10300 ( .A1(u5_mult_82_ab_37__35_), .A2(
        u5_mult_82_CARRYB_36__35_), .ZN(u5_mult_82_n5124) );
  NAND2_X2 u5_mult_82_U10299 ( .A1(u5_mult_82_CARRYB_35__36_), .A2(
        u5_mult_82_n710), .ZN(u5_mult_82_n5123) );
  NAND2_X2 u5_mult_82_U10298 ( .A1(u5_mult_82_ab_36__36_), .A2(u5_mult_82_n710), .ZN(u5_mult_82_n5122) );
  NAND2_X1 u5_mult_82_U10297 ( .A1(u5_mult_82_ab_36__36_), .A2(
        u5_mult_82_CARRYB_35__36_), .ZN(u5_mult_82_n5121) );
  NAND3_X2 u5_mult_82_U10296 ( .A1(u5_mult_82_n5118), .A2(u5_mult_82_n5119), 
        .A3(u5_mult_82_n5120), .ZN(u5_mult_82_CARRYB_46__26_) );
  NAND2_X1 u5_mult_82_U10295 ( .A1(u5_mult_82_CARRYB_45__26_), .A2(
        u5_mult_82_SUMB_45__27_), .ZN(u5_mult_82_n5120) );
  NAND2_X1 u5_mult_82_U10294 ( .A1(u5_mult_82_ab_46__26_), .A2(
        u5_mult_82_SUMB_45__27_), .ZN(u5_mult_82_n5119) );
  NAND2_X1 u5_mult_82_U10293 ( .A1(u5_mult_82_ab_46__26_), .A2(
        u5_mult_82_CARRYB_45__26_), .ZN(u5_mult_82_n5118) );
  NAND2_X2 u5_mult_82_U10292 ( .A1(u5_mult_82_n465), .A2(u5_mult_82_n1408), 
        .ZN(u5_mult_82_n5117) );
  NAND2_X2 u5_mult_82_U10291 ( .A1(u5_mult_82_ab_45__27_), .A2(
        u5_mult_82_n1408), .ZN(u5_mult_82_n5116) );
  NAND2_X1 u5_mult_82_U10290 ( .A1(u5_mult_82_ab_45__27_), .A2(
        u5_mult_82_CARRYB_44__27_), .ZN(u5_mult_82_n5115) );
  XOR2_X2 u5_mult_82_U10289 ( .A(u5_mult_82_n5114), .B(u5_mult_82_n1408), .Z(
        u5_mult_82_SUMB_45__27_) );
  XOR2_X2 u5_mult_82_U10288 ( .A(u5_mult_82_ab_45__27_), .B(
        u5_mult_82_CARRYB_44__27_), .Z(u5_mult_82_n5114) );
  NAND3_X2 u5_mult_82_U10287 ( .A1(u5_mult_82_n5111), .A2(u5_mult_82_n5112), 
        .A3(u5_mult_82_n5113), .ZN(u5_mult_82_CARRYB_40__32_) );
  NAND2_X1 u5_mult_82_U10286 ( .A1(u5_mult_82_SUMB_39__33_), .A2(
        u5_mult_82_CARRYB_39__32_), .ZN(u5_mult_82_n5113) );
  NAND2_X1 u5_mult_82_U10285 ( .A1(u5_mult_82_ab_40__32_), .A2(
        u5_mult_82_CARRYB_39__32_), .ZN(u5_mult_82_n5111) );
  NAND3_X2 u5_mult_82_U10284 ( .A1(u5_mult_82_n5108), .A2(u5_mult_82_n5109), 
        .A3(u5_mult_82_n5110), .ZN(u5_mult_82_CARRYB_39__33_) );
  NAND2_X2 u5_mult_82_U10283 ( .A1(u5_mult_82_CARRYB_38__33_), .A2(
        u5_mult_82_SUMB_38__34_), .ZN(u5_mult_82_n5110) );
  NAND2_X2 u5_mult_82_U10282 ( .A1(u5_mult_82_ab_39__33_), .A2(
        u5_mult_82_SUMB_38__34_), .ZN(u5_mult_82_n5109) );
  NAND2_X1 u5_mult_82_U10281 ( .A1(u5_mult_82_ab_39__33_), .A2(
        u5_mult_82_CARRYB_38__33_), .ZN(u5_mult_82_n5108) );
  XOR2_X2 u5_mult_82_U10280 ( .A(u5_mult_82_n5107), .B(u5_mult_82_n1560), .Z(
        u5_mult_82_SUMB_39__33_) );
  XOR2_X2 u5_mult_82_U10279 ( .A(u5_mult_82_ab_39__33_), .B(
        u5_mult_82_CARRYB_38__33_), .Z(u5_mult_82_n5107) );
  NAND3_X2 u5_mult_82_U10278 ( .A1(u5_mult_82_n5104), .A2(u5_mult_82_n5105), 
        .A3(u5_mult_82_n5106), .ZN(u5_mult_82_CARRYB_52__20_) );
  NAND2_X1 u5_mult_82_U10277 ( .A1(u5_mult_82_CARRYB_51__20_), .A2(
        u5_mult_82_SUMB_51__21_), .ZN(u5_mult_82_n5106) );
  NAND2_X1 u5_mult_82_U10276 ( .A1(u5_mult_82_ab_52__20_), .A2(
        u5_mult_82_SUMB_51__21_), .ZN(u5_mult_82_n5105) );
  NAND2_X1 u5_mult_82_U10275 ( .A1(u5_mult_82_ab_52__20_), .A2(
        u5_mult_82_CARRYB_51__20_), .ZN(u5_mult_82_n5104) );
  NAND2_X2 u5_mult_82_U10274 ( .A1(u5_mult_82_SUMB_50__22_), .A2(
        u5_mult_82_ab_51__21_), .ZN(u5_mult_82_n5102) );
  XOR2_X2 u5_mult_82_U10273 ( .A(u5_mult_82_n5100), .B(u5_mult_82_SUMB_51__21_), .Z(u5_mult_82_SUMB_52__20_) );
  NAND3_X2 u5_mult_82_U10272 ( .A1(u5_mult_82_n5097), .A2(u5_mult_82_n5098), 
        .A3(u5_mult_82_n5099), .ZN(u5_mult_82_CARRYB_50__22_) );
  NAND2_X2 u5_mult_82_U10271 ( .A1(u5_mult_82_ab_50__22_), .A2(
        u5_mult_82_SUMB_49__23_), .ZN(u5_mult_82_n5098) );
  NOR2_X2 u5_mult_82_U10270 ( .A1(u5_mult_82_n6775), .A2(u5_mult_82_n6531), 
        .ZN(u5_mult_82_ab_7__49_) );
  NOR2_X1 u5_mult_82_U10269 ( .A1(u5_mult_82_n6774), .A2(u5_mult_82_n6628), 
        .ZN(u5_mult_82_ab_21__49_) );
  NOR2_X1 u5_mult_82_U10268 ( .A1(u5_mult_82_n6832), .A2(u5_mult_82_n6693), 
        .ZN(u5_mult_82_ab_32__39_) );
  NOR2_X2 u5_mult_82_U10267 ( .A1(u5_mult_82_n6895), .A2(u5_mult_82_net65229), 
        .ZN(u5_mult_82_ab_50__21_) );
  NAND3_X2 u5_mult_82_U10266 ( .A1(u5_mult_82_n5094), .A2(u5_mult_82_n5095), 
        .A3(u5_mult_82_n5096), .ZN(u5_mult_82_CARRYB_7__49_) );
  NAND2_X2 u5_mult_82_U10265 ( .A1(u5_mult_82_ab_7__49_), .A2(
        u5_mult_82_CARRYB_6__49_), .ZN(u5_mult_82_n5095) );
  NAND3_X2 u5_mult_82_U10264 ( .A1(u5_mult_82_n5091), .A2(u5_mult_82_n5092), 
        .A3(u5_mult_82_n5093), .ZN(u5_mult_82_CARRYB_21__49_) );
  NAND2_X1 u5_mult_82_U10263 ( .A1(u5_mult_82_ab_21__49_), .A2(
        u5_mult_82_SUMB_20__50_), .ZN(u5_mult_82_n5093) );
  NAND2_X2 u5_mult_82_U10262 ( .A1(u5_mult_82_ab_21__49_), .A2(
        u5_mult_82_CARRYB_20__49_), .ZN(u5_mult_82_n5092) );
  NAND2_X1 u5_mult_82_U10261 ( .A1(u5_mult_82_SUMB_20__50_), .A2(
        u5_mult_82_CARRYB_20__49_), .ZN(u5_mult_82_n5091) );
  NAND3_X2 u5_mult_82_U10260 ( .A1(u5_mult_82_n5087), .A2(u5_mult_82_n5088), 
        .A3(u5_mult_82_n5089), .ZN(u5_mult_82_CARRYB_3__51_) );
  NAND2_X2 u5_mult_82_U10259 ( .A1(u5_mult_82_ab_2__52_), .A2(
        u5_mult_82_ab_3__51_), .ZN(u5_mult_82_n5089) );
  NAND2_X2 u5_mult_82_U10258 ( .A1(u5_mult_82_CARRYB_2__51_), .A2(
        u5_mult_82_ab_2__52_), .ZN(u5_mult_82_n5088) );
  NAND2_X2 u5_mult_82_U10257 ( .A1(u5_mult_82_CARRYB_2__51_), .A2(
        u5_mult_82_ab_3__51_), .ZN(u5_mult_82_n5087) );
  NAND2_X1 u5_mult_82_U10256 ( .A1(u5_mult_82_ab_36__35_), .A2(
        u5_mult_82_CARRYB_35__35_), .ZN(u5_mult_82_n5084) );
  NAND3_X4 u5_mult_82_U10255 ( .A1(u5_mult_82_n5081), .A2(u5_mult_82_n5082), 
        .A3(u5_mult_82_n5083), .ZN(u5_mult_82_CARRYB_35__36_) );
  NAND2_X2 u5_mult_82_U10254 ( .A1(u5_mult_82_ab_35__36_), .A2(
        u5_mult_82_SUMB_34__37_), .ZN(u5_mult_82_n5082) );
  NAND2_X1 u5_mult_82_U10253 ( .A1(u5_mult_82_ab_32__39_), .A2(
        u5_mult_82_CARRYB_31__39_), .ZN(u5_mult_82_n5080) );
  NAND2_X1 u5_mult_82_U10252 ( .A1(u5_mult_82_CARRYB_31__39_), .A2(
        u5_mult_82_SUMB_31__40_), .ZN(u5_mult_82_n5078) );
  NAND3_X2 u5_mult_82_U10251 ( .A1(u5_mult_82_n5075), .A2(u5_mult_82_n5076), 
        .A3(u5_mult_82_n5077), .ZN(u5_mult_82_CARRYB_52__19_) );
  NAND2_X1 u5_mult_82_U10250 ( .A1(u5_mult_82_CARRYB_51__19_), .A2(
        u5_mult_82_SUMB_51__20_), .ZN(u5_mult_82_n5077) );
  NAND2_X1 u5_mult_82_U10249 ( .A1(u5_mult_82_ab_52__19_), .A2(
        u5_mult_82_SUMB_51__20_), .ZN(u5_mult_82_n5076) );
  NAND2_X1 u5_mult_82_U10248 ( .A1(u5_mult_82_ab_52__19_), .A2(
        u5_mult_82_CARRYB_51__19_), .ZN(u5_mult_82_n5075) );
  NAND3_X4 u5_mult_82_U10247 ( .A1(u5_mult_82_n5073), .A2(u5_mult_82_n5074), 
        .A3(u5_mult_82_n5072), .ZN(u5_mult_82_CARRYB_51__20_) );
  NAND2_X2 u5_mult_82_U10246 ( .A1(u5_mult_82_CARRYB_50__20_), .A2(
        u5_mult_82_SUMB_50__21_), .ZN(u5_mult_82_n5074) );
  NAND2_X2 u5_mult_82_U10245 ( .A1(u5_mult_82_ab_51__20_), .A2(
        u5_mult_82_SUMB_50__21_), .ZN(u5_mult_82_n5073) );
  NAND2_X2 u5_mult_82_U10244 ( .A1(u5_mult_82_ab_51__20_), .A2(
        u5_mult_82_CARRYB_50__20_), .ZN(u5_mult_82_n5072) );
  XOR2_X2 u5_mult_82_U10243 ( .A(u5_mult_82_n5071), .B(u5_mult_82_SUMB_50__21_), .Z(u5_mult_82_SUMB_51__20_) );
  XOR2_X2 u5_mult_82_U10242 ( .A(u5_mult_82_ab_51__20_), .B(
        u5_mult_82_CARRYB_50__20_), .Z(u5_mult_82_n5071) );
  NAND3_X2 u5_mult_82_U10241 ( .A1(u5_mult_82_n5068), .A2(u5_mult_82_n5069), 
        .A3(u5_mult_82_n5070), .ZN(u5_mult_82_CARRYB_50__21_) );
  NAND2_X1 u5_mult_82_U10240 ( .A1(u5_mult_82_ab_50__21_), .A2(
        u5_mult_82_CARRYB_49__21_), .ZN(u5_mult_82_n5070) );
  XOR2_X2 u5_mult_82_U10239 ( .A(u5_mult_82_SUMB_49__22_), .B(u5_mult_82_n5067), .Z(u5_mult_82_SUMB_50__21_) );
  XOR2_X2 u5_mult_82_U10238 ( .A(u5_mult_82_CARRYB_49__21_), .B(
        u5_mult_82_ab_50__21_), .Z(u5_mult_82_n5067) );
  NOR2_X1 u5_mult_82_U10237 ( .A1(u5_mult_82_n6863), .A2(u5_mult_82_n6628), 
        .ZN(u5_mult_82_ab_21__29_) );
  NAND3_X2 u5_mult_82_U10236 ( .A1(u5_mult_82_n5064), .A2(u5_mult_82_n5065), 
        .A3(u5_mult_82_n5066), .ZN(u5_mult_82_CARRYB_42__17_) );
  NAND2_X2 u5_mult_82_U10235 ( .A1(u5_mult_82_ab_42__17_), .A2(
        u5_mult_82_CARRYB_41__17_), .ZN(u5_mult_82_n5065) );
  NAND2_X1 u5_mult_82_U10234 ( .A1(u5_mult_82_CARRYB_40__17_), .A2(
        u5_mult_82_SUMB_40__18_), .ZN(u5_mult_82_n5063) );
  NAND2_X1 u5_mult_82_U10233 ( .A1(u5_mult_82_ab_41__17_), .A2(
        u5_mult_82_SUMB_40__18_), .ZN(u5_mult_82_n5062) );
  NAND2_X1 u5_mult_82_U10232 ( .A1(u5_mult_82_ab_21__29_), .A2(
        u5_mult_82_CARRYB_20__29_), .ZN(u5_mult_82_n5060) );
  NAND2_X2 u5_mult_82_U10231 ( .A1(u5_mult_82_SUMB_20__30_), .A2(
        u5_mult_82_ab_21__29_), .ZN(u5_mult_82_n5059) );
  XOR2_X2 u5_mult_82_U10230 ( .A(u5_mult_82_SUMB_20__30_), .B(u5_mult_82_n5057), .Z(u5_mult_82_SUMB_21__29_) );
  NAND3_X2 u5_mult_82_U10229 ( .A1(u5_mult_82_n5054), .A2(u5_mult_82_n5055), 
        .A3(u5_mult_82_n5056), .ZN(u5_mult_82_CARRYB_16__34_) );
  NAND2_X1 u5_mult_82_U10228 ( .A1(u5_mult_82_CARRYB_15__34_), .A2(
        u5_mult_82_SUMB_15__35_), .ZN(u5_mult_82_n5056) );
  NAND2_X1 u5_mult_82_U10227 ( .A1(u5_mult_82_ab_16__34_), .A2(
        u5_mult_82_SUMB_15__35_), .ZN(u5_mult_82_n5055) );
  NAND3_X2 u5_mult_82_U10226 ( .A1(u5_mult_82_n5053), .A2(u5_mult_82_n5052), 
        .A3(u5_mult_82_n5051), .ZN(u5_mult_82_CARRYB_15__35_) );
  NAND2_X2 u5_mult_82_U10225 ( .A1(u5_mult_82_ab_15__35_), .A2(
        u5_mult_82_SUMB_14__36_), .ZN(u5_mult_82_n5052) );
  NAND2_X1 u5_mult_82_U10224 ( .A1(u5_mult_82_ab_15__35_), .A2(
        u5_mult_82_CARRYB_14__35_), .ZN(u5_mult_82_n5051) );
  XOR2_X2 u5_mult_82_U10223 ( .A(u5_mult_82_n5050), .B(u5_mult_82_SUMB_15__35_), .Z(u5_mult_82_SUMB_16__34_) );
  XOR2_X2 u5_mult_82_U10222 ( .A(u5_mult_82_n5049), .B(u5_mult_82_SUMB_14__36_), .Z(u5_mult_82_SUMB_15__35_) );
  NAND2_X2 u5_mult_82_U10221 ( .A1(u5_mult_82_ab_14__40_), .A2(
        u5_mult_82_CARRYB_13__40_), .ZN(u5_mult_82_n5385) );
  NAND3_X4 u5_mult_82_U10220 ( .A1(u5_mult_82_n5872), .A2(u5_mult_82_n5873), 
        .A3(u5_mult_82_n5871), .ZN(u5_mult_82_CARRYB_33__30_) );
  NAND3_X2 u5_mult_82_U10219 ( .A1(u5_mult_82_n5046), .A2(u5_mult_82_n5047), 
        .A3(u5_mult_82_n5048), .ZN(u5_mult_82_CARRYB_4__46_) );
  NAND2_X1 u5_mult_82_U10218 ( .A1(u5_mult_82_CARRYB_3__46_), .A2(
        u5_mult_82_SUMB_3__47_), .ZN(u5_mult_82_n5048) );
  NAND2_X1 u5_mult_82_U10217 ( .A1(u5_mult_82_ab_4__46_), .A2(
        u5_mult_82_SUMB_3__47_), .ZN(u5_mult_82_n5047) );
  NAND2_X1 u5_mult_82_U10216 ( .A1(u5_mult_82_ab_4__46_), .A2(
        u5_mult_82_CARRYB_3__46_), .ZN(u5_mult_82_n5046) );
  NAND3_X4 u5_mult_82_U10215 ( .A1(u5_mult_82_n5043), .A2(u5_mult_82_n5044), 
        .A3(u5_mult_82_n5045), .ZN(u5_mult_82_CARRYB_3__47_) );
  NAND2_X2 u5_mult_82_U10214 ( .A1(u5_mult_82_CARRYB_2__47_), .A2(
        u5_mult_82_SUMB_2__48_), .ZN(u5_mult_82_n5045) );
  NAND2_X2 u5_mult_82_U10213 ( .A1(u5_mult_82_ab_3__47_), .A2(
        u5_mult_82_SUMB_2__48_), .ZN(u5_mult_82_n5044) );
  NAND2_X2 u5_mult_82_U10212 ( .A1(u5_mult_82_ab_3__47_), .A2(
        u5_mult_82_CARRYB_2__47_), .ZN(u5_mult_82_n5043) );
  XOR2_X2 u5_mult_82_U10211 ( .A(u5_mult_82_n5042), .B(u5_mult_82_SUMB_3__47_), 
        .Z(u5_mult_82_SUMB_4__46_) );
  XOR2_X2 u5_mult_82_U10210 ( .A(u5_mult_82_ab_4__46_), .B(
        u5_mult_82_CARRYB_3__46_), .Z(u5_mult_82_n5042) );
  XOR2_X2 u5_mult_82_U10209 ( .A(u5_mult_82_n5041), .B(u5_mult_82_n1547), .Z(
        u5_mult_82_SUMB_3__47_) );
  XOR2_X2 u5_mult_82_U10208 ( .A(u5_mult_82_ab_3__47_), .B(
        u5_mult_82_CARRYB_2__47_), .Z(u5_mult_82_n5041) );
  NAND3_X2 u5_mult_82_U10207 ( .A1(u5_mult_82_n5035), .A2(u5_mult_82_n5036), 
        .A3(u5_mult_82_n5037), .ZN(u5_mult_82_CARRYB_17__37_) );
  NAND2_X2 u5_mult_82_U10206 ( .A1(u5_mult_82_CARRYB_16__37_), .A2(
        u5_mult_82_SUMB_16__38_), .ZN(u5_mult_82_n5037) );
  NAND2_X2 u5_mult_82_U10205 ( .A1(u5_mult_82_ab_17__37_), .A2(
        u5_mult_82_SUMB_16__38_), .ZN(u5_mult_82_n5036) );
  NAND3_X2 u5_mult_82_U10204 ( .A1(u5_mult_82_n5033), .A2(u5_mult_82_n5032), 
        .A3(u5_mult_82_n5034), .ZN(u5_mult_82_CARRYB_36__24_) );
  NAND2_X1 u5_mult_82_U10203 ( .A1(u5_mult_82_CARRYB_35__24_), .A2(
        u5_mult_82_SUMB_35__25_), .ZN(u5_mult_82_n5034) );
  NAND2_X1 u5_mult_82_U10202 ( .A1(u5_mult_82_ab_36__24_), .A2(
        u5_mult_82_SUMB_35__25_), .ZN(u5_mult_82_n5033) );
  NAND2_X2 u5_mult_82_U10201 ( .A1(u5_mult_82_CARRYB_34__25_), .A2(
        u5_mult_82_n1815), .ZN(u5_mult_82_n5031) );
  NAND2_X2 u5_mult_82_U10200 ( .A1(u5_mult_82_ab_35__25_), .A2(
        u5_mult_82_n1815), .ZN(u5_mult_82_n5030) );
  XOR2_X2 u5_mult_82_U10199 ( .A(u5_mult_82_n5028), .B(u5_mult_82_n1815), .Z(
        u5_mult_82_SUMB_35__25_) );
  XOR2_X2 u5_mult_82_U10198 ( .A(u5_mult_82_ab_35__25_), .B(
        u5_mult_82_CARRYB_34__25_), .Z(u5_mult_82_n5028) );
  XNOR2_X2 u5_mult_82_U10197 ( .A(u5_mult_82_net83274), .B(u5_mult_82_net80786), .ZN(u5_mult_82_SUMB_14__29_) );
  XOR2_X2 u5_mult_82_U10196 ( .A(u5_mult_82_n6261), .B(u5_mult_82_n1488), .Z(
        u5_mult_82_SUMB_46__10_) );
  NAND2_X1 u5_mult_82_U10195 ( .A1(u5_mult_82_CARRYB_20__37_), .A2(
        u5_mult_82_SUMB_20__38_), .ZN(u5_mult_82_n5519) );
  NAND2_X2 u5_mult_82_U10194 ( .A1(u5_mult_82_ab_13__37_), .A2(
        u5_mult_82_SUMB_12__38_), .ZN(u5_mult_82_n6093) );
  XNOR2_X2 u5_mult_82_U10193 ( .A(u5_mult_82_ab_44__8_), .B(
        u5_mult_82_CARRYB_43__8_), .ZN(u5_mult_82_n5027) );
  NOR2_X1 u5_mult_82_U10192 ( .A1(u5_mult_82_n6920), .A2(u5_mult_82_n6721), 
        .ZN(u5_mult_82_ab_37__18_) );
  NAND2_X1 u5_mult_82_U10191 ( .A1(u5_mult_82_CARRYB_15__35_), .A2(
        u5_mult_82_SUMB_15__36_), .ZN(u5_mult_82_n5026) );
  NAND2_X1 u5_mult_82_U10190 ( .A1(u5_mult_82_ab_16__35_), .A2(
        u5_mult_82_SUMB_15__36_), .ZN(u5_mult_82_n5025) );
  NAND2_X1 u5_mult_82_U10189 ( .A1(u5_mult_82_ab_16__35_), .A2(
        u5_mult_82_CARRYB_15__35_), .ZN(u5_mult_82_n5024) );
  NAND2_X2 u5_mult_82_U10188 ( .A1(u5_mult_82_n1859), .A2(
        u5_mult_82_CARRYB_14__36_), .ZN(u5_mult_82_n5023) );
  NAND2_X1 u5_mult_82_U10187 ( .A1(u5_mult_82_ab_15__36_), .A2(
        u5_mult_82_CARRYB_14__36_), .ZN(u5_mult_82_n5021) );
  XOR2_X2 u5_mult_82_U10186 ( .A(u5_mult_82_n5020), .B(u5_mult_82_SUMB_15__36_), .Z(u5_mult_82_SUMB_16__35_) );
  NAND3_X4 u5_mult_82_U10185 ( .A1(u5_mult_82_n5017), .A2(u5_mult_82_n5018), 
        .A3(u5_mult_82_n5019), .ZN(u5_mult_82_CARRYB_41__14_) );
  NAND2_X2 u5_mult_82_U10184 ( .A1(u5_mult_82_CARRYB_40__14_), .A2(
        u5_mult_82_SUMB_40__15_), .ZN(u5_mult_82_n5019) );
  NAND2_X2 u5_mult_82_U10183 ( .A1(u5_mult_82_ab_41__14_), .A2(
        u5_mult_82_SUMB_40__15_), .ZN(u5_mult_82_n5018) );
  NAND2_X1 u5_mult_82_U10182 ( .A1(u5_mult_82_ab_41__14_), .A2(
        u5_mult_82_CARRYB_40__14_), .ZN(u5_mult_82_n5017) );
  NAND2_X2 u5_mult_82_U10181 ( .A1(u5_mult_82_CARRYB_39__15_), .A2(
        u5_mult_82_SUMB_39__16_), .ZN(u5_mult_82_n5016) );
  NAND2_X2 u5_mult_82_U10180 ( .A1(u5_mult_82_ab_40__15_), .A2(
        u5_mult_82_SUMB_39__16_), .ZN(u5_mult_82_n5015) );
  NAND2_X1 u5_mult_82_U10179 ( .A1(u5_mult_82_ab_40__15_), .A2(
        u5_mult_82_CARRYB_39__15_), .ZN(u5_mult_82_n5014) );
  NAND3_X2 u5_mult_82_U10178 ( .A1(u5_mult_82_n5011), .A2(u5_mult_82_n5012), 
        .A3(u5_mult_82_n5013), .ZN(u5_mult_82_CARRYB_37__18_) );
  NAND2_X1 u5_mult_82_U10177 ( .A1(u5_mult_82_ab_37__18_), .A2(
        u5_mult_82_CARRYB_36__18_), .ZN(u5_mult_82_n5013) );
  NAND2_X2 u5_mult_82_U10176 ( .A1(u5_mult_82_ab_37__18_), .A2(
        u5_mult_82_SUMB_36__19_), .ZN(u5_mult_82_n5012) );
  XOR2_X2 u5_mult_82_U10175 ( .A(u5_mult_82_SUMB_36__19_), .B(u5_mult_82_n5010), .Z(u5_mult_82_SUMB_37__18_) );
  XOR2_X2 u5_mult_82_U10174 ( .A(u5_mult_82_CARRYB_36__18_), .B(
        u5_mult_82_ab_37__18_), .Z(u5_mult_82_n5010) );
  NAND3_X2 u5_mult_82_U10173 ( .A1(u5_mult_82_n5007), .A2(u5_mult_82_n5008), 
        .A3(u5_mult_82_n5009), .ZN(u5_mult_82_CARRYB_50__7_) );
  NAND2_X1 u5_mult_82_U10172 ( .A1(u5_mult_82_ab_50__7_), .A2(
        u5_mult_82_SUMB_49__8_), .ZN(u5_mult_82_n5008) );
  NAND2_X1 u5_mult_82_U10171 ( .A1(u5_mult_82_ab_50__7_), .A2(
        u5_mult_82_CARRYB_49__7_), .ZN(u5_mult_82_n5007) );
  NAND3_X4 u5_mult_82_U10170 ( .A1(u5_mult_82_n5004), .A2(u5_mult_82_n5005), 
        .A3(u5_mult_82_n5006), .ZN(u5_mult_82_CARRYB_43__12_) );
  NAND2_X2 u5_mult_82_U10169 ( .A1(u5_mult_82_ab_43__12_), .A2(
        u5_mult_82_SUMB_42__13_), .ZN(u5_mult_82_n5006) );
  NAND2_X2 u5_mult_82_U10168 ( .A1(u5_mult_82_CARRYB_42__12_), .A2(
        u5_mult_82_SUMB_42__13_), .ZN(u5_mult_82_n5005) );
  NAND3_X4 u5_mult_82_U10167 ( .A1(u5_mult_82_net80797), .A2(u5_mult_82_n5003), 
        .A3(u5_mult_82_net80795), .ZN(u5_mult_82_CARRYB_42__13_) );
  NAND2_X2 u5_mult_82_U10166 ( .A1(u5_mult_82_ab_42__13_), .A2(
        u5_mult_82_SUMB_41__14_), .ZN(u5_mult_82_n5003) );
  XOR2_X2 u5_mult_82_U10165 ( .A(u5_mult_82_net80793), .B(
        u5_mult_82_SUMB_41__14_), .Z(u5_mult_82_SUMB_42__13_) );
  NOR2_X1 u5_mult_82_U10164 ( .A1(u5_mult_82_n6904), .A2(u5_mult_82_n6728), 
        .ZN(u5_mult_82_ab_39__20_) );
  NAND3_X2 u5_mult_82_U10163 ( .A1(u5_mult_82_n4999), .A2(u5_mult_82_n5000), 
        .A3(u5_mult_82_n5001), .ZN(u5_mult_82_CARRYB_9__42_) );
  NAND2_X1 u5_mult_82_U10162 ( .A1(u5_mult_82_ab_9__42_), .A2(
        u5_mult_82_CARRYB_8__42_), .ZN(u5_mult_82_n5001) );
  NAND2_X2 u5_mult_82_U10161 ( .A1(u5_mult_82_CARRYB_5__44_), .A2(
        u5_mult_82_SUMB_5__45_), .ZN(u5_mult_82_n4998) );
  NAND2_X2 u5_mult_82_U10160 ( .A1(u5_mult_82_ab_6__44_), .A2(
        u5_mult_82_SUMB_5__45_), .ZN(u5_mult_82_n4997) );
  NAND2_X1 u5_mult_82_U10159 ( .A1(u5_mult_82_ab_6__44_), .A2(
        u5_mult_82_CARRYB_5__44_), .ZN(u5_mult_82_n4996) );
  NAND3_X2 u5_mult_82_U10158 ( .A1(u5_mult_82_n4993), .A2(u5_mult_82_n4994), 
        .A3(u5_mult_82_n4995), .ZN(u5_mult_82_CARRYB_5__45_) );
  NAND2_X1 u5_mult_82_U10157 ( .A1(u5_mult_82_ab_5__45_), .A2(
        u5_mult_82_CARRYB_4__45_), .ZN(u5_mult_82_n4993) );
  XOR2_X2 u5_mult_82_U10156 ( .A(u5_mult_82_n4992), .B(u5_mult_82_SUMB_4__46_), 
        .Z(u5_mult_82_SUMB_5__45_) );
  NAND3_X2 u5_mult_82_U10155 ( .A1(u5_mult_82_n4989), .A2(u5_mult_82_n4990), 
        .A3(u5_mult_82_n4991), .ZN(u5_mult_82_CARRYB_22__34_) );
  NAND2_X1 u5_mult_82_U10154 ( .A1(u5_mult_82_ab_22__34_), .A2(
        u5_mult_82_CARRYB_21__34_), .ZN(u5_mult_82_n4989) );
  NAND2_X2 u5_mult_82_U10153 ( .A1(u5_mult_82_ab_21__35_), .A2(
        u5_mult_82_SUMB_20__36_), .ZN(u5_mult_82_n4987) );
  NAND2_X1 u5_mult_82_U10152 ( .A1(u5_mult_82_CARRYB_40__18_), .A2(
        u5_mult_82_SUMB_40__19_), .ZN(u5_mult_82_n4985) );
  NAND2_X1 u5_mult_82_U10151 ( .A1(u5_mult_82_ab_41__18_), .A2(
        u5_mult_82_SUMB_40__19_), .ZN(u5_mult_82_n4984) );
  NAND2_X1 u5_mult_82_U10150 ( .A1(u5_mult_82_ab_41__18_), .A2(
        u5_mult_82_CARRYB_40__18_), .ZN(u5_mult_82_n4983) );
  NAND3_X4 u5_mult_82_U10149 ( .A1(u5_mult_82_n4980), .A2(u5_mult_82_n4981), 
        .A3(u5_mult_82_n4982), .ZN(u5_mult_82_CARRYB_40__19_) );
  NAND2_X2 u5_mult_82_U10148 ( .A1(u5_mult_82_CARRYB_39__19_), .A2(
        u5_mult_82_SUMB_39__20_), .ZN(u5_mult_82_n4982) );
  NAND2_X2 u5_mult_82_U10147 ( .A1(u5_mult_82_ab_40__19_), .A2(
        u5_mult_82_SUMB_39__20_), .ZN(u5_mult_82_n4981) );
  NAND2_X2 u5_mult_82_U10146 ( .A1(u5_mult_82_ab_40__19_), .A2(
        u5_mult_82_CARRYB_39__19_), .ZN(u5_mult_82_n4980) );
  NAND3_X2 u5_mult_82_U10145 ( .A1(u5_mult_82_n4977), .A2(u5_mult_82_n4978), 
        .A3(u5_mult_82_n4979), .ZN(u5_mult_82_CARRYB_39__20_) );
  NAND2_X1 u5_mult_82_U10144 ( .A1(u5_mult_82_ab_39__20_), .A2(
        u5_mult_82_CARRYB_38__20_), .ZN(u5_mult_82_n4979) );
  NAND2_X2 u5_mult_82_U10143 ( .A1(u5_mult_82_ab_39__20_), .A2(
        u5_mult_82_SUMB_38__21_), .ZN(u5_mult_82_n4978) );
  NOR2_X2 u5_mult_82_U10142 ( .A1(u5_mult_82_net64363), .A2(
        u5_mult_82_net65409), .ZN(u5_mult_82_ab_40__5_) );
  INV_X2 u5_mult_82_U10141 ( .A(u5_mult_82_ab_45__2_), .ZN(u5_mult_82_n5398)
         );
  NAND3_X2 u5_mult_82_U10140 ( .A1(u5_mult_82_n4974), .A2(u5_mult_82_n4975), 
        .A3(u5_mult_82_n4976), .ZN(u5_mult_82_CARRYB_27__11_) );
  NAND2_X1 u5_mult_82_U10139 ( .A1(u5_mult_82_SUMB_26__12_), .A2(
        u5_mult_82_CARRYB_26__11_), .ZN(u5_mult_82_n4976) );
  NAND2_X1 u5_mult_82_U10138 ( .A1(u5_mult_82_ab_27__11_), .A2(
        u5_mult_82_SUMB_26__12_), .ZN(u5_mult_82_n4975) );
  NAND2_X1 u5_mult_82_U10137 ( .A1(u5_mult_82_ab_27__11_), .A2(
        u5_mult_82_CARRYB_26__11_), .ZN(u5_mult_82_n4974) );
  NAND3_X2 u5_mult_82_U10136 ( .A1(u5_mult_82_n4971), .A2(u5_mult_82_n4972), 
        .A3(u5_mult_82_n4973), .ZN(u5_mult_82_CARRYB_26__12_) );
  NAND2_X1 u5_mult_82_U10135 ( .A1(u5_mult_82_CARRYB_25__12_), .A2(
        u5_mult_82_SUMB_25__13_), .ZN(u5_mult_82_n4973) );
  NAND2_X1 u5_mult_82_U10134 ( .A1(u5_mult_82_ab_26__12_), .A2(
        u5_mult_82_SUMB_25__13_), .ZN(u5_mult_82_n4972) );
  NAND2_X1 u5_mult_82_U10133 ( .A1(u5_mult_82_ab_26__12_), .A2(
        u5_mult_82_CARRYB_25__12_), .ZN(u5_mult_82_n4971) );
  XOR2_X2 u5_mult_82_U10132 ( .A(u5_mult_82_n4970), .B(u5_mult_82_SUMB_26__12_), .Z(u5_mult_82_SUMB_27__11_) );
  XOR2_X2 u5_mult_82_U10131 ( .A(u5_mult_82_n4969), .B(u5_mult_82_SUMB_25__13_), .Z(u5_mult_82_SUMB_26__12_) );
  XOR2_X2 u5_mult_82_U10130 ( .A(u5_mult_82_ab_26__12_), .B(
        u5_mult_82_CARRYB_25__12_), .Z(u5_mult_82_n4969) );
  NAND3_X2 u5_mult_82_U10129 ( .A1(u5_mult_82_n4966), .A2(u5_mult_82_n4967), 
        .A3(u5_mult_82_n4968), .ZN(u5_mult_82_CARRYB_40__5_) );
  NAND3_X2 u5_mult_82_U10128 ( .A1(u5_mult_82_n4965), .A2(u5_mult_82_n4964), 
        .A3(u5_mult_82_n4963), .ZN(u5_mult_82_CARRYB_42__3_) );
  NAND2_X2 u5_mult_82_U10127 ( .A1(u5_mult_82_CARRYB_41__3_), .A2(
        u5_mult_82_SUMB_41__4_), .ZN(u5_mult_82_n4965) );
  NAND2_X2 u5_mult_82_U10126 ( .A1(u5_mult_82_ab_42__3_), .A2(
        u5_mult_82_SUMB_41__4_), .ZN(u5_mult_82_n4964) );
  NAND3_X2 u5_mult_82_U10125 ( .A1(u5_mult_82_n4960), .A2(u5_mult_82_n4961), 
        .A3(u5_mult_82_n4962), .ZN(u5_mult_82_CARRYB_41__4_) );
  NAND2_X2 u5_mult_82_U10124 ( .A1(u5_mult_82_ab_41__4_), .A2(
        u5_mult_82_SUMB_40__5_), .ZN(u5_mult_82_n4961) );
  XOR2_X2 u5_mult_82_U10123 ( .A(u5_mult_82_CARRYB_41__3_), .B(
        u5_mult_82_ab_42__3_), .Z(u5_mult_82_n4959) );
  NAND2_X2 u5_mult_82_U10122 ( .A1(u5_mult_82_ab_45__2_), .A2(u5_mult_82_n1832), .ZN(u5_mult_82_n4958) );
  XNOR2_X2 u5_mult_82_U10121 ( .A(u5_mult_82_n5653), .B(
        u5_mult_82_SUMB_22__39_), .ZN(u5_mult_82_SUMB_23__38_) );
  NAND2_X1 u5_mult_82_U10120 ( .A1(u5_mult_82_ab_34__14_), .A2(
        u5_mult_82_CARRYB_33__14_), .ZN(u5_mult_82_n4951) );
  XOR2_X2 u5_mult_82_U10119 ( .A(u5_mult_82_n4950), .B(u5_mult_82_SUMB_34__14_), .Z(u5_mult_82_SUMB_35__13_) );
  XOR2_X2 u5_mult_82_U10118 ( .A(u5_mult_82_ab_35__13_), .B(
        u5_mult_82_CARRYB_34__13_), .Z(u5_mult_82_n4950) );
  NAND2_X1 u5_mult_82_U10117 ( .A1(u5_mult_82_ab_32__32_), .A2(
        u5_mult_82_CARRYB_31__32_), .ZN(u5_mult_82_n5944) );
  NAND2_X2 u5_mult_82_U10116 ( .A1(u5_mult_82_ab_41__6_), .A2(u5_mult_82_n1755), .ZN(u5_mult_82_n5822) );
  XOR2_X2 u5_mult_82_U10115 ( .A(u5_mult_82_n5203), .B(u5_mult_82_SUMB_38__9_), 
        .Z(u5_mult_82_SUMB_39__8_) );
  NOR2_X1 u5_mult_82_U10114 ( .A1(u5_mult_82_net64939), .A2(
        u5_mult_82_net65675), .ZN(u5_mult_82_ab_25__37_) );
  NAND3_X2 u5_mult_82_U10113 ( .A1(u5_mult_82_n4947), .A2(u5_mult_82_n4948), 
        .A3(u5_mult_82_n4949), .ZN(u5_mult_82_CARRYB_25__37_) );
  NAND2_X1 u5_mult_82_U10112 ( .A1(u5_mult_82_ab_25__37_), .A2(
        u5_mult_82_CARRYB_24__37_), .ZN(u5_mult_82_n4949) );
  NAND2_X2 u5_mult_82_U10111 ( .A1(u5_mult_82_ab_25__37_), .A2(
        u5_mult_82_SUMB_24__38_), .ZN(u5_mult_82_n4948) );
  NAND2_X1 u5_mult_82_U10110 ( .A1(u5_mult_82_CARRYB_24__37_), .A2(
        u5_mult_82_SUMB_24__38_), .ZN(u5_mult_82_n4947) );
  NAND2_X2 u5_mult_82_U10109 ( .A1(u5_mult_82_ab_21__39_), .A2(
        u5_mult_82_SUMB_20__40_), .ZN(u5_mult_82_n4945) );
  NAND3_X2 u5_mult_82_U10108 ( .A1(u5_mult_82_n4938), .A2(u5_mult_82_n4939), 
        .A3(u5_mult_82_n4940), .ZN(u5_mult_82_CARRYB_30__32_) );
  NAND2_X1 u5_mult_82_U10107 ( .A1(u5_mult_82_CARRYB_29__32_), .A2(
        u5_mult_82_SUMB_29__33_), .ZN(u5_mult_82_n4940) );
  NAND2_X1 u5_mult_82_U10106 ( .A1(u5_mult_82_ab_30__32_), .A2(
        u5_mult_82_SUMB_29__33_), .ZN(u5_mult_82_n4939) );
  NAND2_X1 u5_mult_82_U10105 ( .A1(u5_mult_82_ab_30__32_), .A2(
        u5_mult_82_CARRYB_29__32_), .ZN(u5_mult_82_n4938) );
  NAND2_X2 u5_mult_82_U10104 ( .A1(u5_mult_82_CARRYB_28__33_), .A2(
        u5_mult_82_n1550), .ZN(u5_mult_82_n4937) );
  NAND2_X2 u5_mult_82_U10103 ( .A1(u5_mult_82_ab_29__33_), .A2(
        u5_mult_82_n1550), .ZN(u5_mult_82_n4936) );
  NAND2_X2 u5_mult_82_U10102 ( .A1(u5_mult_82_ab_29__33_), .A2(
        u5_mult_82_CARRYB_28__33_), .ZN(u5_mult_82_n4935) );
  NAND2_X1 u5_mult_82_U10101 ( .A1(u5_mult_82_CARRYB_26__35_), .A2(
        u5_mult_82_SUMB_26__36_), .ZN(u5_mult_82_n4932) );
  NOR2_X1 u5_mult_82_U10100 ( .A1(u5_mult_82_n6822), .A2(u5_mult_82_n6630), 
        .ZN(u5_mult_82_ab_21__41_) );
  NOR2_X1 u5_mult_82_U10099 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6693), 
        .ZN(u5_mult_82_ab_32__38_) );
  NOR2_X1 u5_mult_82_U10098 ( .A1(u5_mult_82_n6879), .A2(u5_mult_82_n6735), 
        .ZN(u5_mult_82_ab_44__26_) );
  NAND3_X2 u5_mult_82_U10097 ( .A1(u5_mult_82_n4929), .A2(u5_mult_82_n4930), 
        .A3(u5_mult_82_n4931), .ZN(u5_mult_82_CARRYB_21__41_) );
  NAND2_X1 u5_mult_82_U10096 ( .A1(u5_mult_82_ab_21__41_), .A2(
        u5_mult_82_SUMB_20__42_), .ZN(u5_mult_82_n4931) );
  NAND2_X2 u5_mult_82_U10095 ( .A1(u5_mult_82_ab_21__41_), .A2(
        u5_mult_82_CARRYB_20__41_), .ZN(u5_mult_82_n4930) );
  NAND2_X1 u5_mult_82_U10094 ( .A1(u5_mult_82_SUMB_20__42_), .A2(
        u5_mult_82_CARRYB_20__41_), .ZN(u5_mult_82_n4929) );
  XOR2_X2 u5_mult_82_U10093 ( .A(u5_mult_82_CARRYB_20__41_), .B(
        u5_mult_82_n4928), .Z(u5_mult_82_SUMB_21__41_) );
  NAND3_X2 u5_mult_82_U10092 ( .A1(u5_mult_82_n4925), .A2(u5_mult_82_n4926), 
        .A3(u5_mult_82_n4927), .ZN(u5_mult_82_CARRYB_32__38_) );
  NAND3_X2 u5_mult_82_U10091 ( .A1(u5_mult_82_n4921), .A2(u5_mult_82_n4922), 
        .A3(u5_mult_82_n4923), .ZN(u5_mult_82_CARRYB_44__26_) );
  NAND2_X1 u5_mult_82_U10090 ( .A1(u5_mult_82_CARRYB_43__26_), .A2(
        u5_mult_82_SUMB_43__27_), .ZN(u5_mult_82_n4921) );
  XOR2_X2 u5_mult_82_U10089 ( .A(u5_mult_82_SUMB_43__27_), .B(u5_mult_82_n4920), .Z(u5_mult_82_SUMB_44__26_) );
  NAND2_X1 u5_mult_82_U10088 ( .A1(u5_mult_82_ab_40__30_), .A2(
        u5_mult_82_CARRYB_39__30_), .ZN(u5_mult_82_n4917) );
  NAND2_X2 u5_mult_82_U10087 ( .A1(u5_mult_82_CARRYB_38__31_), .A2(
        u5_mult_82_SUMB_38__32_), .ZN(u5_mult_82_n4916) );
  NAND2_X2 u5_mult_82_U10086 ( .A1(u5_mult_82_ab_39__31_), .A2(
        u5_mult_82_SUMB_38__32_), .ZN(u5_mult_82_n4915) );
  NAND2_X1 u5_mult_82_U10085 ( .A1(u5_mult_82_ab_39__31_), .A2(
        u5_mult_82_CARRYB_38__31_), .ZN(u5_mult_82_n4914) );
  NAND3_X4 u5_mult_82_U10084 ( .A1(u5_mult_82_n4908), .A2(u5_mult_82_n4909), 
        .A3(u5_mult_82_n4910), .ZN(u5_mult_82_CARRYB_50__20_) );
  NAND2_X2 u5_mult_82_U10083 ( .A1(u5_mult_82_CARRYB_49__20_), .A2(
        u5_mult_82_SUMB_49__21_), .ZN(u5_mult_82_n4910) );
  NAND2_X2 u5_mult_82_U10082 ( .A1(u5_mult_82_ab_50__20_), .A2(
        u5_mult_82_SUMB_49__21_), .ZN(u5_mult_82_n4909) );
  XNOR2_X2 u5_mult_82_U10081 ( .A(u5_mult_82_ab_23__30_), .B(
        u5_mult_82_CARRYB_22__30_), .ZN(u5_mult_82_n4907) );
  XNOR2_X2 u5_mult_82_U10080 ( .A(u5_mult_82_n4906), .B(
        u5_mult_82_CARRYB_15__35_), .ZN(u5_mult_82_n5020) );
  XNOR2_X2 u5_mult_82_U10079 ( .A(u5_mult_82_CARRYB_46__3_), .B(
        u5_mult_82_ab_47__3_), .ZN(u5_mult_82_n4905) );
  XNOR2_X2 u5_mult_82_U10078 ( .A(u5_mult_82_SUMB_46__4_), .B(u5_mult_82_n4905), .ZN(u5_mult_82_SUMB_47__3_) );
  NOR2_X1 u5_mult_82_U10077 ( .A1(u5_mult_82_n6897), .A2(u5_mult_82_n6629), 
        .ZN(u5_mult_82_ab_21__21_) );
  NAND3_X2 u5_mult_82_U10076 ( .A1(u5_mult_82_n4902), .A2(u5_mult_82_n4903), 
        .A3(u5_mult_82_n4904), .ZN(u5_mult_82_CARRYB_21__21_) );
  NAND2_X1 u5_mult_82_U10075 ( .A1(u5_mult_82_ab_21__21_), .A2(
        u5_mult_82_CARRYB_20__21_), .ZN(u5_mult_82_n4904) );
  NAND2_X2 u5_mult_82_U10074 ( .A1(u5_mult_82_ab_21__21_), .A2(
        u5_mult_82_SUMB_20__22_), .ZN(u5_mult_82_n4903) );
  NAND2_X1 u5_mult_82_U10073 ( .A1(u5_mult_82_CARRYB_20__21_), .A2(
        u5_mult_82_SUMB_20__22_), .ZN(u5_mult_82_n4902) );
  XOR2_X2 u5_mult_82_U10072 ( .A(u5_mult_82_SUMB_20__22_), .B(u5_mult_82_n4901), .Z(u5_mult_82_SUMB_21__21_) );
  XOR2_X2 u5_mult_82_U10071 ( .A(u5_mult_82_CARRYB_20__21_), .B(
        u5_mult_82_ab_21__21_), .Z(u5_mult_82_n4901) );
  NAND3_X2 u5_mult_82_U10070 ( .A1(u5_mult_82_n4898), .A2(u5_mult_82_n4899), 
        .A3(u5_mult_82_n4900), .ZN(u5_mult_82_CARRYB_28__15_) );
  NAND2_X1 u5_mult_82_U10069 ( .A1(u5_mult_82_CARRYB_27__15_), .A2(
        u5_mult_82_SUMB_27__16_), .ZN(u5_mult_82_n4899) );
  NAND2_X1 u5_mult_82_U10068 ( .A1(u5_mult_82_CARRYB_27__15_), .A2(
        u5_mult_82_ab_28__15_), .ZN(u5_mult_82_n4898) );
  NAND2_X2 u5_mult_82_U10067 ( .A1(u5_mult_82_CARRYB_26__16_), .A2(
        u5_mult_82_SUMB_26__17_), .ZN(u5_mult_82_n4897) );
  NAND2_X2 u5_mult_82_U10066 ( .A1(u5_mult_82_ab_27__16_), .A2(
        u5_mult_82_SUMB_26__17_), .ZN(u5_mult_82_n4896) );
  NAND2_X1 u5_mult_82_U10065 ( .A1(u5_mult_82_ab_27__16_), .A2(
        u5_mult_82_CARRYB_26__16_), .ZN(u5_mult_82_n4895) );
  XOR2_X2 u5_mult_82_U10064 ( .A(u5_mult_82_n4894), .B(u5_mult_82_SUMB_27__16_), .Z(u5_mult_82_SUMB_28__15_) );
  XOR2_X2 u5_mult_82_U10063 ( .A(u5_mult_82_CARRYB_27__15_), .B(
        u5_mult_82_ab_28__15_), .Z(u5_mult_82_n4894) );
  XOR2_X2 u5_mult_82_U10062 ( .A(u5_mult_82_n4893), .B(u5_mult_82_SUMB_26__17_), .Z(u5_mult_82_SUMB_27__16_) );
  XOR2_X2 u5_mult_82_U10061 ( .A(u5_mult_82_ab_27__16_), .B(
        u5_mult_82_CARRYB_26__16_), .Z(u5_mult_82_n4893) );
  NAND2_X2 u5_mult_82_U10060 ( .A1(u5_mult_82_SUMB_42__7_), .A2(
        u5_mult_82_ab_43__6_), .ZN(u5_mult_82_n6031) );
  NAND2_X1 u5_mult_82_U10059 ( .A1(u5_mult_82_ab_12__46_), .A2(
        u5_mult_82_n1866), .ZN(u5_mult_82_n4892) );
  NAND3_X4 u5_mult_82_U10058 ( .A1(u5_mult_82_n4884), .A2(u5_mult_82_n4885), 
        .A3(u5_mult_82_n4886), .ZN(u5_mult_82_CARRYB_17__44_) );
  NAND2_X2 u5_mult_82_U10057 ( .A1(u5_mult_82_CARRYB_16__44_), .A2(
        u5_mult_82_SUMB_16__45_), .ZN(u5_mult_82_n4886) );
  NAND2_X2 u5_mult_82_U10056 ( .A1(u5_mult_82_ab_17__44_), .A2(
        u5_mult_82_SUMB_16__45_), .ZN(u5_mult_82_n4885) );
  NAND2_X1 u5_mult_82_U10055 ( .A1(u5_mult_82_ab_17__44_), .A2(
        u5_mult_82_CARRYB_16__44_), .ZN(u5_mult_82_n4884) );
  XOR2_X2 u5_mult_82_U10054 ( .A(u5_mult_82_n4883), .B(u5_mult_82_SUMB_16__45_), .Z(u5_mult_82_SUMB_17__44_) );
  XOR2_X2 u5_mult_82_U10053 ( .A(u5_mult_82_ab_17__44_), .B(
        u5_mult_82_CARRYB_16__44_), .Z(u5_mult_82_n4883) );
  NAND3_X2 u5_mult_82_U10052 ( .A1(u5_mult_82_n4880), .A2(u5_mult_82_n4881), 
        .A3(u5_mult_82_n4882), .ZN(u5_mult_82_CARRYB_16__45_) );
  NAND2_X1 u5_mult_82_U10051 ( .A1(u5_mult_82_CARRYB_15__45_), .A2(
        u5_mult_82_SUMB_15__46_), .ZN(u5_mult_82_n4882) );
  NAND2_X1 u5_mult_82_U10050 ( .A1(u5_mult_82_ab_16__45_), .A2(
        u5_mult_82_SUMB_15__46_), .ZN(u5_mult_82_n4881) );
  NAND2_X1 u5_mult_82_U10049 ( .A1(u5_mult_82_ab_16__45_), .A2(
        u5_mult_82_CARRYB_15__45_), .ZN(u5_mult_82_n4880) );
  NAND3_X2 u5_mult_82_U10048 ( .A1(u5_mult_82_n4877), .A2(u5_mult_82_n4878), 
        .A3(u5_mult_82_n4879), .ZN(u5_mult_82_CARRYB_15__46_) );
  NAND2_X1 u5_mult_82_U10047 ( .A1(u5_mult_82_ab_15__46_), .A2(
        u5_mult_82_CARRYB_14__46_), .ZN(u5_mult_82_n4877) );
  NAND3_X4 u5_mult_82_U10046 ( .A1(u5_mult_82_n4874), .A2(u5_mult_82_n4875), 
        .A3(u5_mult_82_n4876), .ZN(u5_mult_82_CARRYB_36__29_) );
  NAND2_X1 u5_mult_82_U10045 ( .A1(u5_mult_82_ab_36__29_), .A2(
        u5_mult_82_CARRYB_35__29_), .ZN(u5_mult_82_n4874) );
  NAND3_X2 u5_mult_82_U10044 ( .A1(u5_mult_82_n4871), .A2(u5_mult_82_n4872), 
        .A3(u5_mult_82_n4873), .ZN(u5_mult_82_CARRYB_35__30_) );
  NAND2_X2 u5_mult_82_U10043 ( .A1(u5_mult_82_ab_35__30_), .A2(
        u5_mult_82_SUMB_34__31_), .ZN(u5_mult_82_n4872) );
  NAND2_X1 u5_mult_82_U10042 ( .A1(u5_mult_82_ab_35__30_), .A2(
        u5_mult_82_CARRYB_34__30_), .ZN(u5_mult_82_n4871) );
  XNOR2_X2 u5_mult_82_U10041 ( .A(u5_mult_82_SUMB_50__4_), .B(
        u5_mult_82_ab_51__3_), .ZN(u5_mult_82_n4870) );
  XNOR2_X2 u5_mult_82_U10040 ( .A(u5_mult_82_n4870), .B(
        u5_mult_82_CARRYB_50__3_), .ZN(u5_mult_82_SUMB_51__3_) );
  XNOR2_X2 u5_mult_82_U10039 ( .A(u5_mult_82_CARRYB_41__7_), .B(
        u5_mult_82_ab_42__7_), .ZN(u5_mult_82_n4869) );
  XNOR2_X2 u5_mult_82_U10038 ( .A(u5_mult_82_n4869), .B(u5_mult_82_n47), .ZN(
        u5_mult_82_SUMB_42__7_) );
  NAND2_X1 u5_mult_82_U10037 ( .A1(u5_mult_82_ab_39__28_), .A2(
        u5_mult_82_CARRYB_38__28_), .ZN(u5_mult_82_n5280) );
  XNOR2_X2 u5_mult_82_U10036 ( .A(u5_mult_82_ab_26__28_), .B(
        u5_mult_82_CARRYB_25__28_), .ZN(u5_mult_82_n4867) );
  XNOR2_X2 u5_mult_82_U10035 ( .A(u5_mult_82_n4866), .B(
        u5_mult_82_CARRYB_16__32_), .ZN(u5_mult_82_n6044) );
  NOR2_X1 u5_mult_82_U10034 ( .A1(u5_mult_82_net64887), .A2(u5_mult_82_n6578), 
        .ZN(u5_mult_82_ab_14__34_) );
  NAND2_X1 u5_mult_82_U10033 ( .A1(u5_mult_82_ab_16__32_), .A2(
        u5_mult_82_SUMB_15__33_), .ZN(u5_mult_82_n4863) );
  NAND2_X1 u5_mult_82_U10032 ( .A1(u5_mult_82_ab_16__32_), .A2(
        u5_mult_82_CARRYB_15__32_), .ZN(u5_mult_82_n4862) );
  XOR2_X2 u5_mult_82_U10031 ( .A(u5_mult_82_n4858), .B(u5_mult_82_SUMB_14__34_), .Z(u5_mult_82_SUMB_15__33_) );
  NAND3_X2 u5_mult_82_U10030 ( .A1(u5_mult_82_n4855), .A2(u5_mult_82_n4856), 
        .A3(u5_mult_82_n4857), .ZN(u5_mult_82_CARRYB_14__34_) );
  NAND2_X1 u5_mult_82_U10029 ( .A1(u5_mult_82_ab_14__34_), .A2(
        u5_mult_82_CARRYB_13__34_), .ZN(u5_mult_82_n4857) );
  NAND2_X1 u5_mult_82_U10028 ( .A1(u5_mult_82_CARRYB_13__34_), .A2(
        u5_mult_82_SUMB_13__35_), .ZN(u5_mult_82_n4855) );
  XOR2_X2 u5_mult_82_U10027 ( .A(u5_mult_82_SUMB_13__35_), .B(u5_mult_82_n4854), .Z(u5_mult_82_SUMB_14__34_) );
  XOR2_X2 u5_mult_82_U10026 ( .A(u5_mult_82_CARRYB_13__34_), .B(
        u5_mult_82_ab_14__34_), .Z(u5_mult_82_n4854) );
  XNOR2_X2 u5_mult_82_U10025 ( .A(u5_mult_82_ab_30__32_), .B(
        u5_mult_82_CARRYB_29__32_), .ZN(u5_mult_82_n4853) );
  NAND3_X2 u5_mult_82_U10024 ( .A1(u5_mult_82_n6006), .A2(u5_mult_82_n6007), 
        .A3(u5_mult_82_n6008), .ZN(u5_mult_82_CARRYB_42__6_) );
  XNOR2_X2 u5_mult_82_U10023 ( .A(u5_mult_82_n4852), .B(
        u5_mult_82_CARRYB_45__6_), .ZN(u5_mult_82_n6165) );
  NOR2_X1 u5_mult_82_U10022 ( .A1(u5_mult_82_n6987), .A2(u5_mult_82_net65411), 
        .ZN(u5_mult_82_ab_40__0_) );
  NOR2_X1 u5_mult_82_U10021 ( .A1(u5_mult_82_n6987), .A2(u5_mult_82_n6730), 
        .ZN(u5_mult_82_ab_39__0_) );
  NOR2_X1 u5_mult_82_U10020 ( .A1(u5_mult_82_n6986), .A2(u5_mult_82_n6737), 
        .ZN(u5_mult_82_ab_44__0_) );
  NOR2_X1 u5_mult_82_U10019 ( .A1(u5_mult_82_n6986), .A2(u5_mult_82_net65355), 
        .ZN(u5_mult_82_ab_43__0_) );
  NAND2_X2 u5_mult_82_U10018 ( .A1(u5_mult_82_ab_40__0_), .A2(
        u5_mult_82_SUMB_39__1_), .ZN(u5_mult_82_n4850) );
  XOR2_X2 u5_mult_82_U10017 ( .A(u5_mult_82_CARRYB_39__0_), .B(
        u5_mult_82_ab_40__0_), .Z(u5_mult_82_n4848) );
  NAND3_X2 u5_mult_82_U10016 ( .A1(u5_mult_82_n4845), .A2(u5_mult_82_n4846), 
        .A3(u5_mult_82_n4847), .ZN(u5_mult_82_CARRYB_39__0_) );
  NAND2_X2 u5_mult_82_U10015 ( .A1(u5_mult_82_ab_39__0_), .A2(
        u5_mult_82_SUMB_38__1_), .ZN(u5_mult_82_n4846) );
  NAND3_X2 u5_mult_82_U10014 ( .A1(u5_mult_82_n4841), .A2(u5_mult_82_n4842), 
        .A3(u5_mult_82_n4843), .ZN(u5_mult_82_CARRYB_44__0_) );
  NAND2_X2 u5_mult_82_U10013 ( .A1(u5_mult_82_ab_44__0_), .A2(
        u5_mult_82_SUMB_43__1_), .ZN(u5_mult_82_n4842) );
  XOR2_X2 u5_mult_82_U10012 ( .A(u5_mult_82_SUMB_43__1_), .B(u5_mult_82_n4840), 
        .Z(u5_N44) );
  NAND3_X2 u5_mult_82_U10011 ( .A1(u5_mult_82_n4837), .A2(u5_mult_82_n4838), 
        .A3(u5_mult_82_n4839), .ZN(u5_mult_82_CARRYB_43__0_) );
  NAND2_X2 u5_mult_82_U10010 ( .A1(u5_mult_82_ab_43__0_), .A2(
        u5_mult_82_SUMB_42__1_), .ZN(u5_mult_82_n4838) );
  XOR2_X2 u5_mult_82_U10009 ( .A(u5_mult_82_SUMB_42__1_), .B(u5_mult_82_n4836), 
        .Z(u5_N43) );
  NAND3_X2 u5_mult_82_U10008 ( .A1(u5_mult_82_n4833), .A2(u5_mult_82_n4834), 
        .A3(u5_mult_82_n4835), .ZN(u5_mult_82_CARRYB_26__13_) );
  NAND2_X2 u5_mult_82_U10007 ( .A1(u5_mult_82_CARRYB_24__14_), .A2(
        u5_mult_82_SUMB_24__15_), .ZN(u5_mult_82_n4832) );
  NAND2_X2 u5_mult_82_U10006 ( .A1(u5_mult_82_ab_25__14_), .A2(
        u5_mult_82_SUMB_24__15_), .ZN(u5_mult_82_n4831) );
  NAND2_X1 u5_mult_82_U10005 ( .A1(u5_mult_82_ab_25__14_), .A2(
        u5_mult_82_CARRYB_24__14_), .ZN(u5_mult_82_n4830) );
  XOR2_X2 u5_mult_82_U10004 ( .A(u5_mult_82_n4829), .B(u5_mult_82_n78), .Z(
        u5_mult_82_SUMB_26__13_) );
  XOR2_X2 u5_mult_82_U10003 ( .A(u5_mult_82_n4828), .B(u5_mult_82_n1795), .Z(
        u5_mult_82_SUMB_25__14_) );
  NOR2_X1 u5_mult_82_U10002 ( .A1(u5_mult_82_net64667), .A2(
        u5_mult_82_net65443), .ZN(u5_mult_82_ab_38__22_) );
  NAND3_X2 u5_mult_82_U10001 ( .A1(u5_mult_82_n4825), .A2(u5_mult_82_n4826), 
        .A3(u5_mult_82_n4827), .ZN(u5_mult_82_CARRYB_37__23_) );
  NAND2_X1 u5_mult_82_U10000 ( .A1(u5_mult_82_SUMB_36__24_), .A2(
        u5_mult_82_CARRYB_36__23_), .ZN(u5_mult_82_n4827) );
  NAND2_X2 u5_mult_82_U9999 ( .A1(u5_mult_82_ab_37__23_), .A2(
        u5_mult_82_CARRYB_36__23_), .ZN(u5_mult_82_n4826) );
  NAND2_X1 u5_mult_82_U9998 ( .A1(u5_mult_82_ab_37__23_), .A2(
        u5_mult_82_SUMB_36__24_), .ZN(u5_mult_82_n4825) );
  XOR2_X2 u5_mult_82_U9997 ( .A(u5_mult_82_n4824), .B(
        u5_mult_82_CARRYB_36__23_), .Z(u5_mult_82_SUMB_37__23_) );
  XOR2_X2 u5_mult_82_U9996 ( .A(u5_mult_82_ab_37__23_), .B(
        u5_mult_82_SUMB_36__24_), .Z(u5_mult_82_n4824) );
  NAND3_X2 u5_mult_82_U9995 ( .A1(u5_mult_82_n4821), .A2(u5_mult_82_n4822), 
        .A3(u5_mult_82_n4823), .ZN(u5_mult_82_CARRYB_36__23_) );
  NAND2_X1 u5_mult_82_U9994 ( .A1(u5_mult_82_CARRYB_35__23_), .A2(
        u5_mult_82_SUMB_35__24_), .ZN(u5_mult_82_n4823) );
  NAND2_X2 u5_mult_82_U9993 ( .A1(u5_mult_82_ab_36__23_), .A2(
        u5_mult_82_SUMB_35__24_), .ZN(u5_mult_82_n4822) );
  NAND2_X1 u5_mult_82_U9992 ( .A1(u5_mult_82_ab_36__23_), .A2(
        u5_mult_82_CARRYB_35__23_), .ZN(u5_mult_82_n4821) );
  NAND3_X2 u5_mult_82_U9991 ( .A1(u5_mult_82_n4818), .A2(u5_mult_82_n4820), 
        .A3(u5_mult_82_n4819), .ZN(u5_mult_82_CARRYB_21__33_) );
  NAND2_X2 u5_mult_82_U9990 ( .A1(u5_mult_82_ab_21__33_), .A2(
        u5_mult_82_CARRYB_20__33_), .ZN(u5_mult_82_n4819) );
  XOR2_X2 u5_mult_82_U9989 ( .A(u5_mult_82_n4817), .B(
        u5_mult_82_CARRYB_20__33_), .Z(u5_mult_82_SUMB_21__33_) );
  NAND3_X2 u5_mult_82_U9988 ( .A1(u5_mult_82_n4814), .A2(u5_mult_82_n4815), 
        .A3(u5_mult_82_n4816), .ZN(u5_mult_82_CARRYB_20__33_) );
  NAND2_X1 u5_mult_82_U9987 ( .A1(u5_mult_82_CARRYB_19__33_), .A2(
        u5_mult_82_SUMB_19__34_), .ZN(u5_mult_82_n4815) );
  NAND2_X1 u5_mult_82_U9986 ( .A1(u5_mult_82_CARRYB_19__33_), .A2(
        u5_mult_82_ab_20__33_), .ZN(u5_mult_82_n4814) );
  NAND2_X2 u5_mult_82_U9985 ( .A1(u5_mult_82_CARRYB_23__31_), .A2(
        u5_mult_82_SUMB_23__32_), .ZN(u5_mult_82_n4813) );
  NAND2_X2 u5_mult_82_U9984 ( .A1(u5_mult_82_ab_24__31_), .A2(
        u5_mult_82_SUMB_23__32_), .ZN(u5_mult_82_n4812) );
  NAND2_X1 u5_mult_82_U9983 ( .A1(u5_mult_82_ab_24__31_), .A2(
        u5_mult_82_CARRYB_23__31_), .ZN(u5_mult_82_n4811) );
  NAND2_X2 u5_mult_82_U9982 ( .A1(u5_mult_82_CARRYB_22__32_), .A2(
        u5_mult_82_SUMB_22__33_), .ZN(u5_mult_82_n4810) );
  NAND2_X2 u5_mult_82_U9981 ( .A1(u5_mult_82_ab_23__32_), .A2(
        u5_mult_82_SUMB_22__33_), .ZN(u5_mult_82_n4809) );
  NAND2_X1 u5_mult_82_U9980 ( .A1(u5_mult_82_ab_23__32_), .A2(
        u5_mult_82_CARRYB_22__32_), .ZN(u5_mult_82_n4808) );
  XOR2_X2 u5_mult_82_U9979 ( .A(u5_mult_82_n4807), .B(u5_mult_82_SUMB_23__32_), 
        .Z(u5_mult_82_SUMB_24__31_) );
  XOR2_X2 u5_mult_82_U9978 ( .A(u5_mult_82_ab_24__31_), .B(
        u5_mult_82_CARRYB_23__31_), .Z(u5_mult_82_n4807) );
  NAND3_X2 u5_mult_82_U9977 ( .A1(u5_mult_82_n4804), .A2(u5_mult_82_n4805), 
        .A3(u5_mult_82_n4806), .ZN(u5_mult_82_CARRYB_38__22_) );
  NAND2_X1 u5_mult_82_U9976 ( .A1(u5_mult_82_ab_38__22_), .A2(u5_mult_82_n1623), .ZN(u5_mult_82_n4806) );
  XOR2_X2 u5_mult_82_U9975 ( .A(u5_mult_82_SUMB_37__23_), .B(u5_mult_82_n4803), 
        .Z(u5_mult_82_SUMB_38__22_) );
  XOR2_X2 u5_mult_82_U9974 ( .A(u5_mult_82_CARRYB_37__22_), .B(
        u5_mult_82_ab_38__22_), .Z(u5_mult_82_n4803) );
  NAND3_X4 u5_mult_82_U9973 ( .A1(u5_mult_82_n6027), .A2(u5_mult_82_n6028), 
        .A3(u5_mult_82_n6029), .ZN(u5_mult_82_CARRYB_42__7_) );
  XOR2_X2 u5_mult_82_U9972 ( .A(u5_mult_82_ab_12__45_), .B(
        u5_mult_82_CARRYB_11__45_), .Z(u5_mult_82_n6378) );
  XOR2_X2 u5_mult_82_U9971 ( .A(u5_mult_82_n5439), .B(u5_mult_82_n54), .Z(
        u5_mult_82_SUMB_25__29_) );
  NAND2_X2 u5_mult_82_U9970 ( .A1(u5_mult_82_ab_9__46_), .A2(
        u5_mult_82_SUMB_8__47_), .ZN(u5_mult_82_n4797) );
  NAND3_X2 u5_mult_82_U9969 ( .A1(u5_mult_82_n4793), .A2(u5_mult_82_n4794), 
        .A3(u5_mult_82_n4795), .ZN(u5_mult_82_CARRYB_21__40_) );
  NAND2_X2 u5_mult_82_U9968 ( .A1(u5_mult_82_CARRYB_20__40_), .A2(
        u5_mult_82_SUMB_20__41_), .ZN(u5_mult_82_n4795) );
  NAND2_X2 u5_mult_82_U9967 ( .A1(u5_mult_82_ab_21__40_), .A2(
        u5_mult_82_SUMB_20__41_), .ZN(u5_mult_82_n4794) );
  NAND2_X1 u5_mult_82_U9966 ( .A1(u5_mult_82_ab_21__40_), .A2(
        u5_mult_82_CARRYB_20__40_), .ZN(u5_mult_82_n4793) );
  NAND3_X2 u5_mult_82_U9965 ( .A1(u5_mult_82_n4790), .A2(u5_mult_82_n4791), 
        .A3(u5_mult_82_n4792), .ZN(u5_mult_82_CARRYB_20__41_) );
  NAND2_X1 u5_mult_82_U9964 ( .A1(u5_mult_82_ab_20__41_), .A2(
        u5_mult_82_SUMB_19__42_), .ZN(u5_mult_82_n4792) );
  NAND2_X1 u5_mult_82_U9963 ( .A1(u5_mult_82_CARRYB_19__41_), .A2(
        u5_mult_82_SUMB_19__42_), .ZN(u5_mult_82_n4791) );
  NAND2_X1 u5_mult_82_U9962 ( .A1(u5_mult_82_CARRYB_19__41_), .A2(
        u5_mult_82_ab_20__41_), .ZN(u5_mult_82_n4790) );
  XNOR2_X2 u5_mult_82_U9961 ( .A(u5_mult_82_n1808), .B(u5_mult_82_ab_47__1_), 
        .ZN(u5_mult_82_n4789) );
  XNOR2_X2 u5_mult_82_U9960 ( .A(u5_mult_82_n4787), .B(u5_mult_82_n4101), .ZN(
        u5_mult_82_SUMB_12__46_) );
  NAND2_X2 u5_mult_82_U9959 ( .A1(u5_mult_82_CARRYB_32__13_), .A2(
        u5_mult_82_SUMB_32__14_), .ZN(u5_mult_82_n5211) );
  NOR2_X2 u5_mult_82_U9958 ( .A1(u5_mult_82_net64505), .A2(u5_mult_82_n6695), 
        .ZN(u5_mult_82_ab_32__13_) );
  NAND3_X2 u5_mult_82_U9957 ( .A1(u5_mult_82_n4784), .A2(u5_mult_82_n4785), 
        .A3(u5_mult_82_n4786), .ZN(u5_mult_82_CARRYB_25__19_) );
  NAND2_X1 u5_mult_82_U9956 ( .A1(u5_mult_82_ab_25__19_), .A2(
        u5_mult_82_SUMB_24__20_), .ZN(u5_mult_82_n4785) );
  NAND2_X1 u5_mult_82_U9955 ( .A1(u5_mult_82_ab_25__19_), .A2(
        u5_mult_82_CARRYB_24__19_), .ZN(u5_mult_82_n4784) );
  NAND3_X4 u5_mult_82_U9954 ( .A1(u5_mult_82_n4781), .A2(u5_mult_82_n4782), 
        .A3(u5_mult_82_n4783), .ZN(u5_mult_82_CARRYB_24__20_) );
  NAND2_X2 u5_mult_82_U9953 ( .A1(u5_mult_82_n457), .A2(
        u5_mult_82_SUMB_23__21_), .ZN(u5_mult_82_n4783) );
  NAND2_X2 u5_mult_82_U9952 ( .A1(u5_mult_82_ab_24__20_), .A2(
        u5_mult_82_SUMB_23__21_), .ZN(u5_mult_82_n4782) );
  NAND2_X1 u5_mult_82_U9951 ( .A1(u5_mult_82_CARRYB_23__20_), .A2(
        u5_mult_82_ab_24__20_), .ZN(u5_mult_82_n4781) );
  XOR2_X2 u5_mult_82_U9950 ( .A(u5_mult_82_n4780), .B(u5_mult_82_SUMB_23__21_), 
        .Z(u5_mult_82_SUMB_24__20_) );
  XOR2_X2 u5_mult_82_U9949 ( .A(u5_mult_82_ab_24__20_), .B(
        u5_mult_82_CARRYB_23__20_), .Z(u5_mult_82_n4780) );
  NAND2_X1 u5_mult_82_U9948 ( .A1(u5_mult_82_ab_18__25_), .A2(
        u5_mult_82_CARRYB_17__25_), .ZN(u5_mult_82_n4777) );
  NAND3_X2 u5_mult_82_U9947 ( .A1(u5_mult_82_n4775), .A2(u5_mult_82_n4774), 
        .A3(u5_mult_82_n4776), .ZN(u5_mult_82_CARRYB_17__26_) );
  NAND2_X1 u5_mult_82_U9946 ( .A1(u5_mult_82_ab_17__26_), .A2(
        u5_mult_82_CARRYB_16__26_), .ZN(u5_mult_82_n4774) );
  NAND3_X2 u5_mult_82_U9945 ( .A1(u5_mult_82_n4771), .A2(u5_mult_82_n4772), 
        .A3(u5_mult_82_n4773), .ZN(u5_mult_82_CARRYB_39__9_) );
  NAND2_X1 u5_mult_82_U9944 ( .A1(u5_mult_82_CARRYB_38__9_), .A2(
        u5_mult_82_SUMB_38__10_), .ZN(u5_mult_82_n4773) );
  NAND2_X1 u5_mult_82_U9943 ( .A1(u5_mult_82_ab_39__9_), .A2(
        u5_mult_82_SUMB_38__10_), .ZN(u5_mult_82_n4772) );
  NAND2_X2 u5_mult_82_U9942 ( .A1(u5_mult_82_ab_38__10_), .A2(
        u5_mult_82_SUMB_37__11_), .ZN(u5_mult_82_n4770) );
  NAND2_X2 u5_mult_82_U9941 ( .A1(u5_mult_82_CARRYB_37__10_), .A2(
        u5_mult_82_SUMB_37__11_), .ZN(u5_mult_82_n4769) );
  NAND2_X1 u5_mult_82_U9940 ( .A1(u5_mult_82_CARRYB_37__10_), .A2(
        u5_mult_82_ab_38__10_), .ZN(u5_mult_82_n4768) );
  XOR2_X2 u5_mult_82_U9939 ( .A(u5_mult_82_n4767), .B(u5_mult_82_SUMB_38__10_), 
        .Z(u5_mult_82_SUMB_39__9_) );
  XOR2_X2 u5_mult_82_U9938 ( .A(u5_mult_82_ab_39__9_), .B(
        u5_mult_82_CARRYB_38__9_), .Z(u5_mult_82_n4767) );
  XOR2_X2 u5_mult_82_U9937 ( .A(u5_mult_82_n4766), .B(u5_mult_82_SUMB_37__11_), 
        .Z(u5_mult_82_SUMB_38__10_) );
  XOR2_X2 u5_mult_82_U9936 ( .A(u5_mult_82_CARRYB_37__10_), .B(
        u5_mult_82_ab_38__10_), .Z(u5_mult_82_n4766) );
  NAND2_X1 u5_mult_82_U9935 ( .A1(u5_mult_82_ab_32__13_), .A2(
        u5_mult_82_CARRYB_31__13_), .ZN(u5_mult_82_n4765) );
  NAND2_X1 u5_mult_82_U9934 ( .A1(u5_mult_82_CARRYB_31__13_), .A2(
        u5_mult_82_SUMB_31__14_), .ZN(u5_mult_82_n4763) );
  NAND3_X2 u5_mult_82_U9933 ( .A1(u5_mult_82_n4760), .A2(u5_mult_82_n4761), 
        .A3(u5_mult_82_n4762), .ZN(u5_mult_82_CARRYB_39__17_) );
  NAND2_X1 u5_mult_82_U9932 ( .A1(u5_mult_82_CARRYB_38__17_), .A2(
        u5_mult_82_SUMB_38__18_), .ZN(u5_mult_82_n4762) );
  NAND2_X1 u5_mult_82_U9931 ( .A1(u5_mult_82_ab_39__17_), .A2(
        u5_mult_82_SUMB_38__18_), .ZN(u5_mult_82_n4761) );
  NAND2_X1 u5_mult_82_U9930 ( .A1(u5_mult_82_ab_39__17_), .A2(
        u5_mult_82_CARRYB_38__17_), .ZN(u5_mult_82_n4760) );
  NAND3_X4 u5_mult_82_U9929 ( .A1(u5_mult_82_n4757), .A2(u5_mult_82_n4758), 
        .A3(u5_mult_82_n4759), .ZN(u5_mult_82_CARRYB_38__18_) );
  NAND2_X2 u5_mult_82_U9928 ( .A1(u5_mult_82_ab_38__18_), .A2(u5_mult_82_n741), 
        .ZN(u5_mult_82_n4758) );
  NAND2_X1 u5_mult_82_U9927 ( .A1(u5_mult_82_ab_38__18_), .A2(
        u5_mult_82_CARRYB_37__18_), .ZN(u5_mult_82_n4757) );
  XOR2_X2 u5_mult_82_U9926 ( .A(u5_mult_82_n4756), .B(u5_mult_82_SUMB_38__18_), 
        .Z(u5_mult_82_SUMB_39__17_) );
  XOR2_X2 u5_mult_82_U9925 ( .A(u5_mult_82_ab_39__17_), .B(
        u5_mult_82_CARRYB_38__17_), .Z(u5_mult_82_n4756) );
  XOR2_X2 u5_mult_82_U9924 ( .A(u5_mult_82_n4755), .B(u5_mult_82_n741), .Z(
        u5_mult_82_SUMB_38__18_) );
  XOR2_X2 u5_mult_82_U9923 ( .A(u5_mult_82_ab_38__18_), .B(
        u5_mult_82_CARRYB_37__18_), .Z(u5_mult_82_n4755) );
  NAND3_X2 u5_mult_82_U9922 ( .A1(u5_mult_82_n4752), .A2(u5_mult_82_n4753), 
        .A3(u5_mult_82_n4754), .ZN(u5_mult_82_CARRYB_11__35_) );
  NAND2_X2 u5_mult_82_U9921 ( .A1(u5_mult_82_ab_11__35_), .A2(
        u5_mult_82_SUMB_10__36_), .ZN(u5_mult_82_n4753) );
  NAND2_X1 u5_mult_82_U9920 ( .A1(u5_mult_82_ab_11__35_), .A2(
        u5_mult_82_CARRYB_10__35_), .ZN(u5_mult_82_n4752) );
  NAND2_X2 u5_mult_82_U9919 ( .A1(u5_mult_82_CARRYB_9__36_), .A2(
        u5_mult_82_SUMB_9__37_), .ZN(u5_mult_82_n4751) );
  NAND2_X2 u5_mult_82_U9918 ( .A1(u5_mult_82_ab_10__36_), .A2(
        u5_mult_82_SUMB_9__37_), .ZN(u5_mult_82_n4750) );
  NAND2_X1 u5_mult_82_U9917 ( .A1(u5_mult_82_ab_10__36_), .A2(
        u5_mult_82_CARRYB_9__36_), .ZN(u5_mult_82_n4749) );
  XOR2_X2 u5_mult_82_U9916 ( .A(u5_mult_82_n4748), .B(u5_mult_82_SUMB_10__36_), 
        .Z(u5_mult_82_SUMB_11__35_) );
  XOR2_X2 u5_mult_82_U9915 ( .A(u5_mult_82_ab_11__35_), .B(
        u5_mult_82_CARRYB_10__35_), .Z(u5_mult_82_n4748) );
  XOR2_X2 u5_mult_82_U9914 ( .A(u5_mult_82_ab_10__36_), .B(
        u5_mult_82_CARRYB_9__36_), .Z(u5_mult_82_n4747) );
  NAND2_X1 u5_mult_82_U9913 ( .A1(u5_mult_82_ab_7__38_), .A2(
        u5_mult_82_CARRYB_6__38_), .ZN(u5_mult_82_n4744) );
  NAND2_X1 u5_mult_82_U9912 ( .A1(u5_mult_82_CARRYB_5__39_), .A2(
        u5_mult_82_SUMB_5__40_), .ZN(u5_mult_82_n4743) );
  NAND2_X1 u5_mult_82_U9911 ( .A1(u5_mult_82_ab_6__39_), .A2(
        u5_mult_82_SUMB_5__40_), .ZN(u5_mult_82_n4742) );
  NAND2_X1 u5_mult_82_U9910 ( .A1(u5_mult_82_ab_6__39_), .A2(
        u5_mult_82_CARRYB_5__39_), .ZN(u5_mult_82_n4741) );
  INV_X8 u5_mult_82_U9909 ( .A(u5_mult_82_n7007), .ZN(u5_mult_82_n6790) );
  NAND2_X2 u5_mult_82_U9908 ( .A1(u5_mult_82_ab_24__17_), .A2(
        u5_mult_82_CARRYB_23__17_), .ZN(u5_mult_82_n5302) );
  NOR2_X1 u5_mult_82_U9907 ( .A1(u5_mult_82_n6928), .A2(u5_mult_82_net65713), 
        .ZN(u5_mult_82_ab_23__17_) );
  NAND3_X4 u5_mult_82_U9906 ( .A1(u5_mult_82_n4738), .A2(u5_mult_82_n4739), 
        .A3(u5_mult_82_n4740), .ZN(u5_mult_82_CARRYB_22__18_) );
  NAND2_X2 u5_mult_82_U9905 ( .A1(u5_mult_82_ab_22__18_), .A2(
        u5_mult_82_CARRYB_21__18_), .ZN(u5_mult_82_n4739) );
  NAND3_X2 u5_mult_82_U9904 ( .A1(u5_mult_82_n4735), .A2(u5_mult_82_n4736), 
        .A3(u5_mult_82_n4737), .ZN(u5_mult_82_CARRYB_21__18_) );
  NAND2_X1 u5_mult_82_U9903 ( .A1(u5_mult_82_CARRYB_20__18_), .A2(
        u5_mult_82_SUMB_20__19_), .ZN(u5_mult_82_n4737) );
  NAND2_X2 u5_mult_82_U9902 ( .A1(u5_mult_82_ab_21__18_), .A2(
        u5_mult_82_SUMB_20__19_), .ZN(u5_mult_82_n4736) );
  NAND2_X1 u5_mult_82_U9901 ( .A1(u5_mult_82_ab_21__18_), .A2(
        u5_mult_82_CARRYB_20__18_), .ZN(u5_mult_82_n4735) );
  NAND3_X4 u5_mult_82_U9900 ( .A1(u5_mult_82_n4732), .A2(u5_mult_82_n4733), 
        .A3(u5_mult_82_n4734), .ZN(u5_mult_82_CARRYB_23__17_) );
  NAND2_X2 u5_mult_82_U9899 ( .A1(u5_mult_82_ab_23__17_), .A2(
        u5_mult_82_SUMB_22__18_), .ZN(u5_mult_82_n4733) );
  NAND2_X2 u5_mult_82_U9898 ( .A1(u5_mult_82_ab_42__4_), .A2(
        u5_mult_82_SUMB_41__5_), .ZN(u5_mult_82_n4731) );
  NAND2_X2 u5_mult_82_U9897 ( .A1(u5_mult_82_CARRYB_41__4_), .A2(
        u5_mult_82_SUMB_41__5_), .ZN(u5_mult_82_n4730) );
  NAND3_X2 u5_mult_82_U9896 ( .A1(u5_mult_82_n4726), .A2(u5_mult_82_n4727), 
        .A3(u5_mult_82_n4728), .ZN(u5_mult_82_CARRYB_41__5_) );
  NAND2_X1 u5_mult_82_U9895 ( .A1(u5_mult_82_ab_41__5_), .A2(
        u5_mult_82_CARRYB_40__5_), .ZN(u5_mult_82_n4726) );
  XNOR2_X2 u5_mult_82_U9894 ( .A(u5_mult_82_SUMB_20__42_), .B(u5_mult_82_n4725), .ZN(u5_mult_82_n4928) );
  XNOR2_X2 u5_mult_82_U9893 ( .A(u5_mult_82_CARRYB_31__39_), .B(
        u5_mult_82_ab_32__39_), .ZN(u5_mult_82_n4723) );
  XNOR2_X2 u5_mult_82_U9892 ( .A(u5_mult_82_n1670), .B(u5_mult_82_n4723), .ZN(
        u5_mult_82_SUMB_32__39_) );
  XNOR2_X2 u5_mult_82_U9891 ( .A(u5_mult_82_ab_44__18_), .B(
        u5_mult_82_CARRYB_43__18_), .ZN(u5_mult_82_n4722) );
  XNOR2_X2 u5_mult_82_U9890 ( .A(u5_mult_82_SUMB_43__19_), .B(u5_mult_82_n4722), .ZN(u5_mult_82_SUMB_44__18_) );
  XNOR2_X2 u5_mult_82_U9889 ( .A(u5_mult_82_SUMB_31__14_), .B(u5_mult_82_n4721), .ZN(u5_mult_82_SUMB_32__13_) );
  NAND2_X2 u5_mult_82_U9888 ( .A1(u5_mult_82_ab_9__47_), .A2(
        u5_mult_82_CARRYB_8__47_), .ZN(u5_mult_82_n5726) );
  NOR2_X1 u5_mult_82_U9887 ( .A1(u5_mult_82_n6775), .A2(u5_mult_82_n6585), 
        .ZN(u5_mult_82_ab_15__49_) );
  NAND3_X2 u5_mult_82_U9886 ( .A1(u5_mult_82_n4718), .A2(u5_mult_82_n4719), 
        .A3(u5_mult_82_n4720), .ZN(u5_mult_82_CARRYB_15__49_) );
  NAND2_X1 u5_mult_82_U9885 ( .A1(u5_mult_82_ab_15__49_), .A2(u5_mult_82_n1392), .ZN(u5_mult_82_n4720) );
  NAND2_X2 u5_mult_82_U9884 ( .A1(u5_mult_82_ab_15__49_), .A2(
        u5_mult_82_CARRYB_14__49_), .ZN(u5_mult_82_n4719) );
  NAND2_X1 u5_mult_82_U9883 ( .A1(u5_mult_82_n1392), .A2(
        u5_mult_82_CARRYB_14__49_), .ZN(u5_mult_82_n4718) );
  XOR2_X2 u5_mult_82_U9882 ( .A(u5_mult_82_CARRYB_14__49_), .B(
        u5_mult_82_n4717), .Z(u5_mult_82_SUMB_15__49_) );
  NAND2_X1 u5_mult_82_U9881 ( .A1(u5_mult_82_ab_39__29_), .A2(
        u5_mult_82_SUMB_38__30_), .ZN(u5_mult_82_n4715) );
  NAND2_X1 u5_mult_82_U9880 ( .A1(u5_mult_82_ab_39__29_), .A2(
        u5_mult_82_CARRYB_38__29_), .ZN(u5_mult_82_n4714) );
  NAND3_X4 u5_mult_82_U9879 ( .A1(u5_mult_82_n4711), .A2(u5_mult_82_n4712), 
        .A3(u5_mult_82_n4713), .ZN(u5_mult_82_CARRYB_38__30_) );
  NAND2_X2 u5_mult_82_U9878 ( .A1(u5_mult_82_ab_38__30_), .A2(
        u5_mult_82_SUMB_37__31_), .ZN(u5_mult_82_n4712) );
  XOR2_X2 u5_mult_82_U9877 ( .A(u5_mult_82_n4710), .B(u5_mult_82_SUMB_37__31_), 
        .Z(u5_mult_82_SUMB_38__30_) );
  XOR2_X2 u5_mult_82_U9876 ( .A(u5_mult_82_n1475), .B(u5_mult_82_ab_38__30_), 
        .Z(u5_mult_82_n4710) );
  NAND3_X2 u5_mult_82_U9875 ( .A1(u5_mult_82_n4707), .A2(u5_mult_82_n4708), 
        .A3(u5_mult_82_n4709), .ZN(u5_mult_82_CARRYB_46__23_) );
  NAND2_X1 u5_mult_82_U9874 ( .A1(u5_mult_82_n1595), .A2(
        u5_mult_82_SUMB_45__24_), .ZN(u5_mult_82_n4709) );
  NAND2_X1 u5_mult_82_U9873 ( .A1(u5_mult_82_ab_46__23_), .A2(
        u5_mult_82_SUMB_45__24_), .ZN(u5_mult_82_n4708) );
  NAND2_X1 u5_mult_82_U9872 ( .A1(u5_mult_82_ab_46__23_), .A2(u5_mult_82_n1595), .ZN(u5_mult_82_n4707) );
  NAND3_X2 u5_mult_82_U9871 ( .A1(u5_mult_82_n4704), .A2(u5_mult_82_n4705), 
        .A3(u5_mult_82_n4706), .ZN(u5_mult_82_CARRYB_45__24_) );
  NAND2_X2 u5_mult_82_U9870 ( .A1(u5_mult_82_CARRYB_44__24_), .A2(
        u5_mult_82_SUMB_44__25_), .ZN(u5_mult_82_n4706) );
  NAND2_X2 u5_mult_82_U9869 ( .A1(u5_mult_82_ab_45__24_), .A2(
        u5_mult_82_SUMB_44__25_), .ZN(u5_mult_82_n4705) );
  NAND2_X1 u5_mult_82_U9868 ( .A1(u5_mult_82_ab_45__24_), .A2(
        u5_mult_82_CARRYB_44__24_), .ZN(u5_mult_82_n4704) );
  XOR2_X2 u5_mult_82_U9867 ( .A(u5_mult_82_n4703), .B(u5_mult_82_SUMB_45__24_), 
        .Z(u5_mult_82_SUMB_46__23_) );
  XNOR2_X2 u5_mult_82_U9866 ( .A(u5_mult_82_n4702), .B(
        u5_mult_82_CARRYB_38__8_), .ZN(u5_mult_82_n5203) );
  NOR2_X1 u5_mult_82_U9865 ( .A1(u5_mult_82_n6974), .A2(u5_mult_82_net64469), 
        .ZN(u5_mult_82_ab_52__11_) );
  NOR2_X1 u5_mult_82_U9864 ( .A1(u5_mult_82_net64469), .A2(u5_mult_82_net65189), .ZN(u5_mult_82_ab_51__11_) );
  INV_X8 u5_mult_82_U9863 ( .A(u5_mult_82_n6397), .ZN(u5_mult_82_CLA_SUM[63])
         );
  NAND3_X2 u5_mult_82_U9862 ( .A1(u5_mult_82_n4699), .A2(u5_mult_82_n4700), 
        .A3(u5_mult_82_n4701), .ZN(u5_mult_82_CARRYB_52__11_) );
  NAND2_X1 u5_mult_82_U9861 ( .A1(u5_mult_82_ab_52__11_), .A2(u5_mult_82_n406), 
        .ZN(u5_mult_82_n4701) );
  NAND2_X2 u5_mult_82_U9860 ( .A1(u5_mult_82_ab_52__11_), .A2(
        u5_mult_82_SUMB_51__12_), .ZN(u5_mult_82_n4700) );
  NAND2_X1 u5_mult_82_U9859 ( .A1(u5_mult_82_CARRYB_51__11_), .A2(
        u5_mult_82_SUMB_51__12_), .ZN(u5_mult_82_n4699) );
  XOR2_X2 u5_mult_82_U9858 ( .A(u5_mult_82_SUMB_51__12_), .B(u5_mult_82_n4698), 
        .Z(u5_mult_82_SUMB_52__11_) );
  NAND3_X2 u5_mult_82_U9857 ( .A1(u5_mult_82_n4695), .A2(u5_mult_82_n4696), 
        .A3(u5_mult_82_n4697), .ZN(u5_mult_82_CARRYB_51__11_) );
  NAND2_X1 u5_mult_82_U9856 ( .A1(u5_mult_82_ab_51__11_), .A2(
        u5_mult_82_CARRYB_50__11_), .ZN(u5_mult_82_n4697) );
  XOR2_X2 u5_mult_82_U9855 ( .A(u5_mult_82_SUMB_50__12_), .B(u5_mult_82_n4694), 
        .Z(u5_mult_82_SUMB_51__11_) );
  XOR2_X2 u5_mult_82_U9854 ( .A(u5_mult_82_CARRYB_50__11_), .B(
        u5_mult_82_ab_51__11_), .Z(u5_mult_82_n4694) );
  INV_X1 u5_mult_82_U9853 ( .A(u5_mult_82_CARRYB_52__10_), .ZN(
        u5_mult_82_n4690) );
  XNOR2_X2 u5_mult_82_U9852 ( .A(u5_mult_82_net81335), .B(
        u5_mult_82_SUMB_16__29_), .ZN(u5_mult_82_SUMB_17__28_) );
  NAND2_X2 u5_mult_82_U9851 ( .A1(u5_mult_82_SUMB_5__51_), .A2(
        u5_mult_82_CARRYB_5__50_), .ZN(u5_mult_82_n6288) );
  INV_X1 u5_mult_82_U9850 ( .A(u5_mult_82_SUMB_46__2_), .ZN(u5_mult_82_n4687)
         );
  NAND3_X2 u5_mult_82_U9849 ( .A1(u5_mult_82_n4683), .A2(u5_mult_82_n4684), 
        .A3(u5_mult_82_n4685), .ZN(u5_mult_82_CARRYB_38__2_) );
  NAND2_X2 u5_mult_82_U9848 ( .A1(u5_mult_82_ab_37__3_), .A2(
        u5_mult_82_SUMB_36__4_), .ZN(u5_mult_82_n4681) );
  XOR2_X2 u5_mult_82_U9847 ( .A(u5_mult_82_n4679), .B(u5_mult_82_SUMB_36__4_), 
        .Z(u5_mult_82_SUMB_37__3_) );
  NOR2_X1 u5_mult_82_U9846 ( .A1(u5_mult_82_n6946), .A2(u5_mult_82_net65355), 
        .ZN(u5_mult_82_ab_43__4_) );
  NAND3_X4 u5_mult_82_U9845 ( .A1(u5_mult_82_n4676), .A2(u5_mult_82_n4677), 
        .A3(u5_mult_82_n4678), .ZN(u5_mult_82_CARRYB_43__4_) );
  NAND2_X2 u5_mult_82_U9844 ( .A1(u5_mult_82_ab_43__4_), .A2(
        u5_mult_82_CARRYB_42__4_), .ZN(u5_mult_82_n4678) );
  NAND2_X2 u5_mult_82_U9843 ( .A1(u5_mult_82_CARRYB_42__4_), .A2(
        u5_mult_82_n3707), .ZN(u5_mult_82_n4676) );
  NOR2_X1 u5_mult_82_U9842 ( .A1(u5_mult_82_n6914), .A2(u5_mult_82_net65713), 
        .ZN(u5_mult_82_ab_23__19_) );
  NOR2_X1 u5_mult_82_U9841 ( .A1(u5_mult_82_n6905), .A2(u5_mult_82_n6629), 
        .ZN(u5_mult_82_ab_21__20_) );
  NAND3_X4 u5_mult_82_U9840 ( .A1(u5_mult_82_n4673), .A2(u5_mult_82_n4674), 
        .A3(u5_mult_82_n4675), .ZN(u5_mult_82_CARRYB_20__21_) );
  NAND2_X2 u5_mult_82_U9839 ( .A1(u5_mult_82_SUMB_19__22_), .A2(
        u5_mult_82_CARRYB_19__21_), .ZN(u5_mult_82_n4675) );
  NAND2_X2 u5_mult_82_U9838 ( .A1(u5_mult_82_ab_20__21_), .A2(
        u5_mult_82_CARRYB_19__21_), .ZN(u5_mult_82_n4674) );
  NAND2_X2 u5_mult_82_U9837 ( .A1(u5_mult_82_ab_20__21_), .A2(
        u5_mult_82_SUMB_19__22_), .ZN(u5_mult_82_n4673) );
  NAND3_X2 u5_mult_82_U9836 ( .A1(u5_mult_82_n4670), .A2(u5_mult_82_n4671), 
        .A3(u5_mult_82_n4672), .ZN(u5_mult_82_CARRYB_19__21_) );
  NAND2_X1 u5_mult_82_U9835 ( .A1(u5_mult_82_CARRYB_18__21_), .A2(
        u5_mult_82_SUMB_18__22_), .ZN(u5_mult_82_n4672) );
  NAND2_X2 u5_mult_82_U9834 ( .A1(u5_mult_82_ab_19__21_), .A2(
        u5_mult_82_SUMB_18__22_), .ZN(u5_mult_82_n4671) );
  NAND2_X1 u5_mult_82_U9833 ( .A1(u5_mult_82_ab_19__21_), .A2(
        u5_mult_82_CARRYB_18__21_), .ZN(u5_mult_82_n4670) );
  XOR2_X2 u5_mult_82_U9832 ( .A(u5_mult_82_n4669), .B(u5_mult_82_SUMB_18__22_), 
        .Z(u5_mult_82_SUMB_19__21_) );
  NAND3_X2 u5_mult_82_U9831 ( .A1(u5_mult_82_n4666), .A2(u5_mult_82_n4667), 
        .A3(u5_mult_82_n4668), .ZN(u5_mult_82_CARRYB_23__19_) );
  NAND2_X1 u5_mult_82_U9830 ( .A1(u5_mult_82_ab_23__19_), .A2(
        u5_mult_82_CARRYB_22__19_), .ZN(u5_mult_82_n4668) );
  NAND2_X2 u5_mult_82_U9829 ( .A1(u5_mult_82_ab_23__19_), .A2(
        u5_mult_82_SUMB_22__20_), .ZN(u5_mult_82_n4667) );
  XOR2_X2 u5_mult_82_U9828 ( .A(u5_mult_82_SUMB_22__20_), .B(u5_mult_82_n4665), 
        .Z(u5_mult_82_SUMB_23__19_) );
  XOR2_X2 u5_mult_82_U9827 ( .A(u5_mult_82_CARRYB_22__19_), .B(
        u5_mult_82_ab_23__19_), .Z(u5_mult_82_n4665) );
  NAND3_X2 u5_mult_82_U9826 ( .A1(u5_mult_82_n4662), .A2(u5_mult_82_n4663), 
        .A3(u5_mult_82_n4664), .ZN(u5_mult_82_CARRYB_21__20_) );
  NAND2_X1 u5_mult_82_U9825 ( .A1(u5_mult_82_ab_21__20_), .A2(
        u5_mult_82_CARRYB_20__20_), .ZN(u5_mult_82_n4664) );
  NAND2_X1 u5_mult_82_U9824 ( .A1(u5_mult_82_ab_46__5_), .A2(
        u5_mult_82_CARRYB_45__5_), .ZN(u5_mult_82_n4659) );
  NAND2_X2 u5_mult_82_U9823 ( .A1(u5_mult_82_CARRYB_44__6_), .A2(
        u5_mult_82_n1610), .ZN(u5_mult_82_n4658) );
  NAND2_X2 u5_mult_82_U9822 ( .A1(u5_mult_82_ab_45__6_), .A2(u5_mult_82_n1610), 
        .ZN(u5_mult_82_n4657) );
  NAND2_X1 u5_mult_82_U9821 ( .A1(u5_mult_82_ab_23__17_), .A2(
        u5_mult_82_CARRYB_22__17_), .ZN(u5_mult_82_n4734) );
  NAND2_X2 u5_mult_82_U9820 ( .A1(u5_mult_82_CARRYB_43__0_), .A2(
        u5_mult_82_SUMB_43__1_), .ZN(u5_mult_82_n4841) );
  NAND2_X1 u5_mult_82_U9819 ( .A1(u5_mult_82_CARRYB_22__36_), .A2(
        u5_mult_82_SUMB_22__37_), .ZN(u5_mult_82_n5738) );
  NAND3_X2 u5_mult_82_U9818 ( .A1(u5_mult_82_n4653), .A2(u5_mult_82_n4654), 
        .A3(u5_mult_82_n4655), .ZN(u5_mult_82_CARRYB_12__51_) );
  NAND2_X2 u5_mult_82_U9817 ( .A1(u5_mult_82_ab_11__52_), .A2(
        u5_mult_82_CARRYB_11__51_), .ZN(u5_mult_82_n4655) );
  NAND2_X2 u5_mult_82_U9816 ( .A1(u5_mult_82_ab_12__51_), .A2(
        u5_mult_82_CARRYB_11__51_), .ZN(u5_mult_82_n4654) );
  NAND2_X2 u5_mult_82_U9815 ( .A1(u5_mult_82_ab_12__51_), .A2(
        u5_mult_82_ab_11__52_), .ZN(u5_mult_82_n4653) );
  XOR2_X1 u5_mult_82_U9814 ( .A(u5_mult_82_n4652), .B(
        u5_mult_82_CARRYB_11__51_), .Z(u5_mult_82_SUMB_12__51_) );
  XOR2_X2 u5_mult_82_U9813 ( .A(u5_mult_82_ab_12__51_), .B(
        u5_mult_82_ab_11__52_), .Z(u5_mult_82_n4652) );
  NAND3_X2 u5_mult_82_U9812 ( .A1(u5_mult_82_n4649), .A2(u5_mult_82_n4650), 
        .A3(u5_mult_82_n4651), .ZN(u5_mult_82_CARRYB_11__51_) );
  NAND2_X2 u5_mult_82_U9811 ( .A1(u5_mult_82_ab_11__51_), .A2(
        u5_mult_82_ab_10__52_), .ZN(u5_mult_82_n4650) );
  NAND2_X1 u5_mult_82_U9810 ( .A1(u5_mult_82_ab_30__36_), .A2(
        u5_mult_82_CARRYB_29__36_), .ZN(u5_mult_82_n4645) );
  NAND2_X2 u5_mult_82_U9809 ( .A1(u5_mult_82_ab_29__37_), .A2(u5_mult_82_n1702), .ZN(u5_mult_82_n4643) );
  NAND2_X1 u5_mult_82_U9808 ( .A1(u5_mult_82_ab_29__37_), .A2(
        u5_mult_82_CARRYB_28__37_), .ZN(u5_mult_82_n4642) );
  XOR2_X2 u5_mult_82_U9807 ( .A(u5_mult_82_n4641), .B(u5_mult_82_SUMB_29__37_), 
        .Z(u5_mult_82_SUMB_30__36_) );
  XOR2_X2 u5_mult_82_U9806 ( .A(u5_mult_82_ab_30__36_), .B(
        u5_mult_82_CARRYB_29__36_), .Z(u5_mult_82_n4641) );
  NAND2_X2 u5_mult_82_U9805 ( .A1(u5_mult_82_ab_10__46_), .A2(
        u5_mult_82_SUMB_9__47_), .ZN(u5_mult_82_n5730) );
  NAND2_X2 u5_mult_82_U9804 ( .A1(u5_mult_82_ab_21__20_), .A2(
        u5_mult_82_SUMB_20__21_), .ZN(u5_mult_82_n4663) );
  NAND2_X2 u5_mult_82_U9803 ( .A1(u5_mult_82_CARRYB_20__20_), .A2(
        u5_mult_82_SUMB_20__21_), .ZN(u5_mult_82_n4662) );
  INV_X16 u5_mult_82_U9802 ( .A(u5_mult_82_n6984), .ZN(u5_mult_82_n6980) );
  INV_X8 u5_mult_82_U9801 ( .A(u5_mult_82_n6979), .ZN(u5_mult_82_n6984) );
  NAND2_X2 u5_mult_82_U9800 ( .A1(u5_mult_82_n1776), .A2(u5_mult_82_n1635), 
        .ZN(u5_mult_82_n6381) );
  XNOR2_X2 u5_mult_82_U9799 ( .A(u5_mult_82_ab_31__17_), .B(
        u5_mult_82_CARRYB_30__17_), .ZN(u5_mult_82_n4639) );
  NAND2_X2 u5_mult_82_U9798 ( .A1(u5_mult_82_ab_49__11_), .A2(
        u5_mult_82_CARRYB_48__11_), .ZN(u5_mult_82_n6111) );
  NAND2_X2 u5_mult_82_U9797 ( .A1(u5_mult_82_CARRYB_19__22_), .A2(
        u5_mult_82_SUMB_19__23_), .ZN(u5_mult_82_n4638) );
  NAND2_X2 u5_mult_82_U9796 ( .A1(u5_mult_82_ab_20__22_), .A2(
        u5_mult_82_SUMB_19__23_), .ZN(u5_mult_82_n4637) );
  NAND2_X1 u5_mult_82_U9795 ( .A1(u5_mult_82_ab_20__22_), .A2(
        u5_mult_82_CARRYB_19__22_), .ZN(u5_mult_82_n4636) );
  NAND3_X2 u5_mult_82_U9794 ( .A1(u5_mult_82_n4633), .A2(u5_mult_82_n4634), 
        .A3(u5_mult_82_n4635), .ZN(u5_mult_82_CARRYB_19__23_) );
  NAND2_X1 u5_mult_82_U9793 ( .A1(u5_mult_82_CARRYB_18__23_), .A2(
        u5_mult_82_SUMB_18__24_), .ZN(u5_mult_82_n4635) );
  NAND2_X1 u5_mult_82_U9792 ( .A1(u5_mult_82_ab_19__23_), .A2(
        u5_mult_82_SUMB_18__24_), .ZN(u5_mult_82_n4634) );
  NAND2_X1 u5_mult_82_U9791 ( .A1(u5_mult_82_ab_19__23_), .A2(
        u5_mult_82_CARRYB_18__23_), .ZN(u5_mult_82_n4633) );
  XOR2_X2 u5_mult_82_U9790 ( .A(u5_mult_82_n4632), .B(u5_mult_82_SUMB_19__23_), 
        .Z(u5_mult_82_SUMB_20__22_) );
  XOR2_X2 u5_mult_82_U9789 ( .A(u5_mult_82_ab_20__22_), .B(
        u5_mult_82_CARRYB_19__22_), .Z(u5_mult_82_n4632) );
  NAND3_X2 u5_mult_82_U9788 ( .A1(u5_mult_82_n4631), .A2(u5_mult_82_n4630), 
        .A3(u5_mult_82_n4629), .ZN(u5_mult_82_CARRYB_17__25_) );
  NAND2_X2 u5_mult_82_U9787 ( .A1(u5_mult_82_ab_16__26_), .A2(
        u5_mult_82_net86785), .ZN(u5_mult_82_n4627) );
  NAND2_X1 u5_mult_82_U9786 ( .A1(u5_mult_82_ab_16__26_), .A2(
        u5_mult_82_CARRYB_15__26_), .ZN(u5_mult_82_n4626) );
  XOR2_X2 u5_mult_82_U9785 ( .A(u5_mult_82_n4624), .B(u5_mult_82_SUMB_38__13_), 
        .Z(u5_mult_82_SUMB_39__12_) );
  XOR2_X2 u5_mult_82_U9784 ( .A(u5_mult_82_ab_39__12_), .B(
        u5_mult_82_CARRYB_38__12_), .Z(u5_mult_82_n4624) );
  XNOR2_X2 u5_mult_82_U9783 ( .A(u5_mult_82_ab_49__12_), .B(
        u5_mult_82_CARRYB_48__12_), .ZN(u5_mult_82_n4622) );
  XNOR2_X2 u5_mult_82_U9782 ( .A(u5_mult_82_n1843), .B(u5_mult_82_n4622), .ZN(
        u5_mult_82_SUMB_49__12_) );
  NOR2_X1 u5_mult_82_U9781 ( .A1(u5_mult_82_net64665), .A2(u5_mult_82_n6735), 
        .ZN(u5_mult_82_ab_44__22_) );
  NAND3_X2 u5_mult_82_U9780 ( .A1(u5_mult_82_n4619), .A2(u5_mult_82_n4620), 
        .A3(u5_mult_82_n4621), .ZN(u5_mult_82_CARRYB_44__22_) );
  NAND2_X1 u5_mult_82_U9779 ( .A1(u5_mult_82_ab_44__22_), .A2(
        u5_mult_82_CARRYB_43__22_), .ZN(u5_mult_82_n4621) );
  NAND2_X1 u5_mult_82_U9778 ( .A1(u5_mult_82_ab_44__22_), .A2(
        u5_mult_82_SUMB_43__23_), .ZN(u5_mult_82_n4620) );
  NAND2_X1 u5_mult_82_U9777 ( .A1(u5_mult_82_CARRYB_43__22_), .A2(
        u5_mult_82_SUMB_43__23_), .ZN(u5_mult_82_n4619) );
  XOR2_X2 u5_mult_82_U9776 ( .A(u5_mult_82_SUMB_43__23_), .B(u5_mult_82_n4618), 
        .Z(u5_mult_82_SUMB_44__22_) );
  XOR2_X2 u5_mult_82_U9775 ( .A(u5_mult_82_CARRYB_43__22_), .B(
        u5_mult_82_ab_44__22_), .Z(u5_mult_82_n4618) );
  XNOR2_X2 u5_mult_82_U9774 ( .A(u5_mult_82_CARRYB_29__31_), .B(
        u5_mult_82_ab_30__31_), .ZN(u5_mult_82_n4617) );
  XNOR2_X2 u5_mult_82_U9773 ( .A(u5_mult_82_SUMB_29__32_), .B(u5_mult_82_n4617), .ZN(u5_mult_82_SUMB_30__31_) );
  XNOR2_X2 u5_mult_82_U9772 ( .A(u5_mult_82_ab_21__18_), .B(
        u5_mult_82_CARRYB_20__18_), .ZN(u5_mult_82_n4616) );
  XNOR2_X2 u5_mult_82_U9771 ( .A(u5_mult_82_n4616), .B(u5_mult_82_SUMB_20__19_), .ZN(u5_mult_82_SUMB_21__18_) );
  NOR2_X1 u5_mult_82_U9770 ( .A1(u5_mult_82_n6791), .A2(u5_mult_82_n6733), 
        .ZN(u5_mult_82_ab_44__46_) );
  NOR2_X1 u5_mult_82_U9769 ( .A1(u5_mult_82_n6791), .A2(u5_mult_82_net65313), 
        .ZN(u5_mult_82_ab_45__46_) );
  NOR2_X1 u5_mult_82_U9768 ( .A1(u5_mult_82_n6791), .A2(u5_mult_82_n6740), 
        .ZN(u5_mult_82_ab_46__46_) );
  NOR2_X1 u5_mult_82_U9767 ( .A1(u5_mult_82_n6791), .A2(u5_mult_82_net65277), 
        .ZN(u5_mult_82_ab_47__46_) );
  NOR2_X1 u5_mult_82_U9766 ( .A1(u5_mult_82_n6791), .A2(u5_mult_82_n6746), 
        .ZN(u5_mult_82_ab_48__46_) );
  NOR2_X1 u5_mult_82_U9765 ( .A1(u5_mult_82_n6791), .A2(u5_mult_82_n6752), 
        .ZN(u5_mult_82_ab_49__46_) );
  NOR2_X1 u5_mult_82_U9764 ( .A1(u5_mult_82_n6791), .A2(u5_mult_82_net65223), 
        .ZN(u5_mult_82_ab_50__46_) );
  NOR2_X1 u5_mult_82_U9763 ( .A1(u5_mult_82_n6791), .A2(u5_mult_82_net65193), 
        .ZN(u5_mult_82_ab_51__46_) );
  NOR2_X1 u5_mult_82_U9762 ( .A1(u5_mult_82_n6977), .A2(u5_mult_82_n6791), 
        .ZN(u5_mult_82_ab_52__46_) );
  NAND3_X2 u5_mult_82_U9761 ( .A1(u5_mult_82_n4612), .A2(u5_mult_82_n4613), 
        .A3(u5_mult_82_n4614), .ZN(u5_mult_82_CARRYB_16__46_) );
  NAND2_X1 u5_mult_82_U9760 ( .A1(u5_mult_82_ab_16__46_), .A2(
        u5_mult_82_CARRYB_15__46_), .ZN(u5_mult_82_n4612) );
  NAND2_X2 u5_mult_82_U9759 ( .A1(u5_mult_82_CARRYB_14__47_), .A2(
        u5_mult_82_SUMB_14__48_), .ZN(u5_mult_82_n4611) );
  NAND2_X2 u5_mult_82_U9758 ( .A1(u5_mult_82_ab_15__47_), .A2(
        u5_mult_82_SUMB_14__48_), .ZN(u5_mult_82_n4610) );
  XOR2_X2 u5_mult_82_U9757 ( .A(u5_mult_82_n4608), .B(u5_mult_82_SUMB_15__47_), 
        .Z(u5_mult_82_SUMB_16__46_) );
  XOR2_X2 u5_mult_82_U9756 ( .A(u5_mult_82_ab_16__46_), .B(
        u5_mult_82_CARRYB_15__46_), .Z(u5_mult_82_n4608) );
  NAND3_X2 u5_mult_82_U9755 ( .A1(u5_mult_82_n4605), .A2(u5_mult_82_n4606), 
        .A3(u5_mult_82_n4607), .ZN(u5_mult_82_CARRYB_21__42_) );
  NAND2_X1 u5_mult_82_U9754 ( .A1(u5_mult_82_CARRYB_20__42_), .A2(
        u5_mult_82_SUMB_20__43_), .ZN(u5_mult_82_n4607) );
  NAND2_X1 u5_mult_82_U9753 ( .A1(u5_mult_82_ab_21__42_), .A2(
        u5_mult_82_SUMB_20__43_), .ZN(u5_mult_82_n4606) );
  NAND2_X1 u5_mult_82_U9752 ( .A1(u5_mult_82_ab_21__42_), .A2(
        u5_mult_82_CARRYB_20__42_), .ZN(u5_mult_82_n4605) );
  NAND2_X2 u5_mult_82_U9751 ( .A1(u5_mult_82_ab_20__43_), .A2(
        u5_mult_82_SUMB_19__44_), .ZN(u5_mult_82_n4603) );
  XOR2_X2 u5_mult_82_U9750 ( .A(u5_mult_82_n4601), .B(u5_mult_82_SUMB_19__44_), 
        .Z(u5_mult_82_SUMB_20__43_) );
  XOR2_X2 u5_mult_82_U9749 ( .A(u5_mult_82_ab_20__43_), .B(
        u5_mult_82_CARRYB_19__43_), .Z(u5_mult_82_n4601) );
  NAND3_X4 u5_mult_82_U9748 ( .A1(u5_mult_82_n4598), .A2(u5_mult_82_n4599), 
        .A3(u5_mult_82_n4600), .ZN(u5_mult_82_CARRYB_46__4_) );
  NAND2_X2 u5_mult_82_U9747 ( .A1(u5_mult_82_CARRYB_45__4_), .A2(
        u5_mult_82_SUMB_45__5_), .ZN(u5_mult_82_n4600) );
  NAND2_X2 u5_mult_82_U9746 ( .A1(u5_mult_82_ab_46__4_), .A2(
        u5_mult_82_SUMB_45__5_), .ZN(u5_mult_82_n4599) );
  NAND2_X1 u5_mult_82_U9745 ( .A1(u5_mult_82_ab_45__5_), .A2(
        u5_mult_82_CARRYB_44__5_), .ZN(u5_mult_82_n4595) );
  INV_X16 u5_mult_82_U9744 ( .A(u5_mult_82_net64949), .ZN(u5_mult_82_net64947)
         );
  NAND3_X2 u5_mult_82_U9743 ( .A1(u5_mult_82_n4592), .A2(u5_mult_82_n4593), 
        .A3(u5_mult_82_n4594), .ZN(u5_mult_82_CARRYB_13__46_) );
  NAND2_X1 u5_mult_82_U9742 ( .A1(u5_mult_82_ab_13__46_), .A2(
        u5_mult_82_SUMB_12__47_), .ZN(u5_mult_82_n4593) );
  NAND3_X2 u5_mult_82_U9741 ( .A1(u5_mult_82_n4589), .A2(u5_mult_82_n4590), 
        .A3(u5_mult_82_n4591), .ZN(u5_mult_82_CARRYB_12__47_) );
  NAND2_X2 u5_mult_82_U9740 ( .A1(u5_mult_82_ab_12__47_), .A2(
        u5_mult_82_SUMB_11__48_), .ZN(u5_mult_82_n4590) );
  XOR2_X2 u5_mult_82_U9739 ( .A(u5_mult_82_n4588), .B(u5_mult_82_SUMB_12__47_), 
        .Z(u5_mult_82_SUMB_13__46_) );
  XOR2_X2 u5_mult_82_U9738 ( .A(u5_mult_82_n4587), .B(u5_mult_82_SUMB_11__48_), 
        .Z(u5_mult_82_SUMB_12__47_) );
  NOR2_X1 u5_mult_82_U9737 ( .A1(u5_mult_82_n6905), .A2(u5_mult_82_n6650), 
        .ZN(u5_mult_82_ab_26__20_) );
  NAND3_X2 u5_mult_82_U9736 ( .A1(u5_mult_82_n4584), .A2(u5_mult_82_n4585), 
        .A3(u5_mult_82_n4586), .ZN(u5_mult_82_CARRYB_26__20_) );
  NAND2_X1 u5_mult_82_U9735 ( .A1(u5_mult_82_CARRYB_25__20_), .A2(
        u5_mult_82_SUMB_25__21_), .ZN(u5_mult_82_n4584) );
  XOR2_X2 u5_mult_82_U9734 ( .A(u5_mult_82_SUMB_25__21_), .B(u5_mult_82_n4583), 
        .Z(u5_mult_82_SUMB_26__20_) );
  XOR2_X2 u5_mult_82_U9733 ( .A(u5_mult_82_CARRYB_25__20_), .B(
        u5_mult_82_ab_26__20_), .Z(u5_mult_82_n4583) );
  INV_X8 u5_mult_82_U9732 ( .A(n4284), .ZN(u5_mult_82_net57161) );
  NAND3_X2 u5_mult_82_U9731 ( .A1(u5_mult_82_n4580), .A2(u5_mult_82_n4581), 
        .A3(u5_mult_82_n4582), .ZN(u5_mult_82_CARRYB_49__24_) );
  NAND2_X1 u5_mult_82_U9730 ( .A1(u5_mult_82_ab_49__24_), .A2(
        u5_mult_82_SUMB_48__25_), .ZN(u5_mult_82_n4581) );
  NAND2_X1 u5_mult_82_U9729 ( .A1(u5_mult_82_ab_49__24_), .A2(
        u5_mult_82_CARRYB_48__24_), .ZN(u5_mult_82_n4580) );
  NAND3_X2 u5_mult_82_U9728 ( .A1(u5_mult_82_n4579), .A2(u5_mult_82_n4578), 
        .A3(u5_mult_82_n4577), .ZN(u5_mult_82_CARRYB_48__25_) );
  NAND2_X2 u5_mult_82_U9727 ( .A1(u5_mult_82_ab_48__25_), .A2(
        u5_mult_82_SUMB_47__26_), .ZN(u5_mult_82_n4578) );
  NAND2_X1 u5_mult_82_U9726 ( .A1(u5_mult_82_ab_48__25_), .A2(
        u5_mult_82_CARRYB_47__25_), .ZN(u5_mult_82_n4577) );
  NAND2_X2 u5_mult_82_U9725 ( .A1(u5_mult_82_ab_46__27_), .A2(
        u5_mult_82_SUMB_45__28_), .ZN(u5_mult_82_n4574) );
  NAND2_X1 u5_mult_82_U9724 ( .A1(u5_mult_82_ab_46__27_), .A2(
        u5_mult_82_CARRYB_45__27_), .ZN(u5_mult_82_n4573) );
  NAND2_X2 u5_mult_82_U9723 ( .A1(u5_mult_82_CARRYB_44__28_), .A2(
        u5_mult_82_SUMB_44__29_), .ZN(u5_mult_82_n4572) );
  NAND2_X2 u5_mult_82_U9722 ( .A1(u5_mult_82_ab_45__28_), .A2(
        u5_mult_82_SUMB_44__29_), .ZN(u5_mult_82_n4571) );
  XOR2_X2 u5_mult_82_U9721 ( .A(u5_mult_82_n4569), .B(u5_mult_82_SUMB_45__28_), 
        .Z(u5_mult_82_SUMB_46__27_) );
  NOR2_X1 u5_mult_82_U9720 ( .A1(u5_mult_82_n6876), .A2(u5_mult_82_n6595), 
        .ZN(u5_mult_82_ab_16__27_) );
  NAND3_X2 u5_mult_82_U9719 ( .A1(u5_mult_82_net81534), .A2(u5_mult_82_n4568), 
        .A3(u5_mult_82_net81536), .ZN(u5_mult_82_CARRYB_16__27_) );
  NAND2_X2 u5_mult_82_U9718 ( .A1(u5_mult_82_ab_16__27_), .A2(
        u5_mult_82_SUMB_15__28_), .ZN(u5_mult_82_n4568) );
  NAND3_X2 u5_mult_82_U9717 ( .A1(u5_mult_82_n4566), .A2(u5_mult_82_net81531), 
        .A3(u5_mult_82_n4567), .ZN(u5_mult_82_CARRYB_22__24_) );
  NAND2_X1 u5_mult_82_U9716 ( .A1(u5_mult_82_ab_22__24_), .A2(
        u5_mult_82_CARRYB_21__24_), .ZN(u5_mult_82_n4567) );
  NAND2_X1 u5_mult_82_U9715 ( .A1(u5_mult_82_CARRYB_21__24_), .A2(
        u5_mult_82_SUMB_21__25_), .ZN(u5_mult_82_n4566) );
  NAND3_X2 u5_mult_82_U9714 ( .A1(u5_mult_82_n4563), .A2(u5_mult_82_n4564), 
        .A3(u5_mult_82_n4565), .ZN(u5_mult_82_CARRYB_30__17_) );
  NAND2_X1 u5_mult_82_U9713 ( .A1(u5_mult_82_ab_30__17_), .A2(
        u5_mult_82_SUMB_29__18_), .ZN(u5_mult_82_n4564) );
  NAND2_X1 u5_mult_82_U9712 ( .A1(u5_mult_82_ab_30__17_), .A2(
        u5_mult_82_CARRYB_29__17_), .ZN(u5_mult_82_n4563) );
  NAND2_X2 u5_mult_82_U9711 ( .A1(u5_mult_82_ab_29__18_), .A2(
        u5_mult_82_SUMB_28__19_), .ZN(u5_mult_82_n4561) );
  NAND2_X1 u5_mult_82_U9710 ( .A1(u5_mult_82_ab_29__18_), .A2(
        u5_mult_82_CARRYB_28__18_), .ZN(u5_mult_82_n4560) );
  XOR2_X2 u5_mult_82_U9709 ( .A(u5_mult_82_n4559), .B(u5_mult_82_SUMB_29__18_), 
        .Z(u5_mult_82_SUMB_30__17_) );
  XOR2_X2 u5_mult_82_U9708 ( .A(u5_mult_82_n4558), .B(u5_mult_82_SUMB_28__19_), 
        .Z(u5_mult_82_SUMB_29__18_) );
  NAND2_X1 u5_mult_82_U9707 ( .A1(u5_mult_82_SUMB_25__34_), .A2(
        u5_mult_82_n4553), .ZN(u5_mult_82_n5769) );
  XNOR2_X2 u5_mult_82_U9706 ( .A(u5_mult_82_SUMB_26__36_), .B(u5_mult_82_n4557), .ZN(u5_mult_82_SUMB_27__35_) );
  NOR2_X1 u5_mult_82_U9705 ( .A1(u5_mult_82_n6885), .A2(u5_mult_82_n6715), 
        .ZN(u5_mult_82_ab_36__25_) );
  NAND3_X2 u5_mult_82_U9704 ( .A1(u5_mult_82_n4554), .A2(u5_mult_82_n4555), 
        .A3(u5_mult_82_n4556), .ZN(u5_mult_82_CARRYB_36__25_) );
  NAND2_X1 u5_mult_82_U9703 ( .A1(u5_mult_82_ab_36__25_), .A2(
        u5_mult_82_CARRYB_35__25_), .ZN(u5_mult_82_n4556) );
  NAND2_X2 u5_mult_82_U9702 ( .A1(u5_mult_82_ab_36__25_), .A2(
        u5_mult_82_SUMB_35__26_), .ZN(u5_mult_82_n4555) );
  NAND2_X1 u5_mult_82_U9701 ( .A1(u5_mult_82_ab_33__13_), .A2(
        u5_mult_82_CARRYB_32__13_), .ZN(u5_mult_82_n5213) );
  NAND3_X2 u5_mult_82_U9700 ( .A1(u5_mult_82_n4550), .A2(u5_mult_82_n4551), 
        .A3(u5_mult_82_n4552), .ZN(u5_mult_82_CARRYB_35__28_) );
  NAND2_X1 u5_mult_82_U9699 ( .A1(u5_mult_82_ab_35__28_), .A2(
        u5_mult_82_SUMB_34__29_), .ZN(u5_mult_82_n4552) );
  NAND2_X1 u5_mult_82_U9698 ( .A1(u5_mult_82_CARRYB_34__28_), .A2(
        u5_mult_82_SUMB_34__29_), .ZN(u5_mult_82_n4551) );
  NAND2_X1 u5_mult_82_U9697 ( .A1(u5_mult_82_CARRYB_34__28_), .A2(
        u5_mult_82_ab_35__28_), .ZN(u5_mult_82_n4550) );
  NAND3_X2 u5_mult_82_U9696 ( .A1(u5_mult_82_n4547), .A2(u5_mult_82_n4548), 
        .A3(u5_mult_82_n4549), .ZN(u5_mult_82_CARRYB_34__29_) );
  NAND2_X2 u5_mult_82_U9695 ( .A1(u5_mult_82_ab_34__29_), .A2(
        u5_mult_82_SUMB_33__30_), .ZN(u5_mult_82_n4548) );
  XOR2_X2 u5_mult_82_U9694 ( .A(u5_mult_82_n4546), .B(u5_mult_82_SUMB_33__30_), 
        .Z(u5_mult_82_SUMB_34__29_) );
  XOR2_X1 u5_mult_82_U9693 ( .A(u5_mult_82_ab_34__29_), .B(
        u5_mult_82_CARRYB_33__29_), .Z(u5_mult_82_n4546) );
  NAND3_X2 u5_mult_82_U9692 ( .A1(u5_mult_82_n4543), .A2(u5_mult_82_n4544), 
        .A3(u5_mult_82_n4545), .ZN(u5_mult_82_CARRYB_32__27_) );
  NAND2_X2 u5_mult_82_U9691 ( .A1(u5_mult_82_ab_31__28_), .A2(
        u5_mult_82_SUMB_30__29_), .ZN(u5_mult_82_n4541) );
  NAND2_X2 u5_mult_82_U9690 ( .A1(u5_mult_82_ab_31__28_), .A2(u5_mult_82_n1628), .ZN(u5_mult_82_n4540) );
  NAND3_X2 u5_mult_82_U9689 ( .A1(u5_mult_82_n4536), .A2(u5_mult_82_n4535), 
        .A3(u5_mult_82_n4534), .ZN(u5_mult_82_CARRYB_29__30_) );
  NAND2_X1 u5_mult_82_U9688 ( .A1(u5_mult_82_ab_29__30_), .A2(
        u5_mult_82_CARRYB_28__30_), .ZN(u5_mult_82_n4534) );
  XOR2_X2 u5_mult_82_U9687 ( .A(u5_mult_82_n4533), .B(u5_mult_82_SUMB_28__31_), 
        .Z(u5_mult_82_SUMB_29__30_) );
  NAND3_X2 u5_mult_82_U9686 ( .A1(u5_mult_82_n5784), .A2(u5_mult_82_n5785), 
        .A3(u5_mult_82_n5786), .ZN(u5_mult_82_CARRYB_20__37_) );
  INV_X2 u5_mult_82_U9685 ( .A(u5_mult_82_ab_21__37_), .ZN(u5_mult_82_n5002)
         );
  NAND2_X2 u5_mult_82_U9684 ( .A1(u5_mult_82_n4530), .A2(u5_mult_82_ab_21__37_), .ZN(u5_mult_82_n4532) );
  NOR2_X1 u5_mult_82_U9683 ( .A1(u5_mult_82_n6967), .A2(u5_mult_82_net65393), 
        .ZN(u5_mult_82_ab_41__1_) );
  NAND3_X2 u5_mult_82_U9682 ( .A1(u5_mult_82_n4527), .A2(u5_mult_82_n4528), 
        .A3(u5_mult_82_n4529), .ZN(u5_mult_82_CARRYB_41__1_) );
  NAND2_X2 u5_mult_82_U9681 ( .A1(u5_mult_82_ab_41__1_), .A2(
        u5_mult_82_SUMB_40__2_), .ZN(u5_mult_82_n4528) );
  NAND3_X2 u5_mult_82_U9680 ( .A1(u5_mult_82_n4524), .A2(u5_mult_82_n4525), 
        .A3(u5_mult_82_n4526), .ZN(u5_mult_82_CARRYB_34__8_) );
  NAND2_X1 u5_mult_82_U9679 ( .A1(u5_mult_82_CARRYB_33__8_), .A2(
        u5_mult_82_SUMB_33__9_), .ZN(u5_mult_82_n4526) );
  NAND2_X1 u5_mult_82_U9678 ( .A1(u5_mult_82_ab_34__8_), .A2(
        u5_mult_82_SUMB_33__9_), .ZN(u5_mult_82_n4525) );
  NAND2_X1 u5_mult_82_U9677 ( .A1(u5_mult_82_ab_34__8_), .A2(
        u5_mult_82_CARRYB_33__8_), .ZN(u5_mult_82_n4524) );
  NAND2_X2 u5_mult_82_U9676 ( .A1(u5_mult_82_n1688), .A2(u5_mult_82_n388), 
        .ZN(u5_mult_82_n4523) );
  NAND2_X2 u5_mult_82_U9675 ( .A1(u5_mult_82_ab_33__9_), .A2(u5_mult_82_n1688), 
        .ZN(u5_mult_82_n4522) );
  NAND2_X1 u5_mult_82_U9674 ( .A1(u5_mult_82_ab_33__9_), .A2(
        u5_mult_82_CARRYB_32__9_), .ZN(u5_mult_82_n4521) );
  XOR2_X2 u5_mult_82_U9673 ( .A(u5_mult_82_n4520), .B(u5_mult_82_SUMB_33__9_), 
        .Z(u5_mult_82_SUMB_34__8_) );
  XOR2_X2 u5_mult_82_U9672 ( .A(u5_mult_82_n4519), .B(u5_mult_82_n1688), .Z(
        u5_mult_82_SUMB_33__9_) );
  NAND2_X2 u5_mult_82_U9671 ( .A1(u5_mult_82_CARRYB_46__2_), .A2(
        u5_mult_82_SUMB_46__3_), .ZN(u5_mult_82_n4517) );
  NAND2_X2 u5_mult_82_U9670 ( .A1(u5_mult_82_ab_47__2_), .A2(
        u5_mult_82_SUMB_46__3_), .ZN(u5_mult_82_n4516) );
  NAND2_X2 u5_mult_82_U9669 ( .A1(u5_mult_82_CARRYB_45__3_), .A2(
        u5_mult_82_SUMB_45__4_), .ZN(u5_mult_82_n4514) );
  NAND2_X2 u5_mult_82_U9668 ( .A1(u5_mult_82_ab_46__3_), .A2(
        u5_mult_82_SUMB_45__4_), .ZN(u5_mult_82_n4513) );
  XOR2_X2 u5_mult_82_U9667 ( .A(u5_mult_82_n4511), .B(u5_mult_82_n412), .Z(
        u5_mult_82_SUMB_47__2_) );
  XNOR2_X2 u5_mult_82_U9666 ( .A(u5_mult_82_CARRYB_22__36_), .B(
        u5_mult_82_ab_23__36_), .ZN(u5_mult_82_n4509) );
  XNOR2_X2 u5_mult_82_U9665 ( .A(u5_mult_82_SUMB_22__37_), .B(u5_mult_82_n4509), .ZN(u5_mult_82_SUMB_23__36_) );
  NAND2_X2 u5_mult_82_U9664 ( .A1(u5_mult_82_n5002), .A2(
        u5_mult_82_CARRYB_20__37_), .ZN(u5_mult_82_n4531) );
  NOR2_X1 u5_mult_82_U9663 ( .A1(u5_mult_82_net64561), .A2(u5_mult_82_n6629), 
        .ZN(u5_mult_82_ab_21__16_) );
  NAND3_X2 u5_mult_82_U9662 ( .A1(u5_mult_82_n4506), .A2(u5_mult_82_n4507), 
        .A3(u5_mult_82_n4508), .ZN(u5_mult_82_CARRYB_21__16_) );
  NAND2_X1 u5_mult_82_U9661 ( .A1(u5_mult_82_ab_21__16_), .A2(
        u5_mult_82_CARRYB_20__16_), .ZN(u5_mult_82_n4508) );
  NAND2_X2 u5_mult_82_U9660 ( .A1(u5_mult_82_ab_21__16_), .A2(
        u5_mult_82_SUMB_20__17_), .ZN(u5_mult_82_n4507) );
  NAND2_X1 u5_mult_82_U9659 ( .A1(u5_mult_82_CARRYB_20__16_), .A2(
        u5_mult_82_SUMB_20__17_), .ZN(u5_mult_82_n4506) );
  NAND3_X2 u5_mult_82_U9658 ( .A1(u5_mult_82_n4503), .A2(u5_mult_82_n4504), 
        .A3(u5_mult_82_n4505), .ZN(u5_mult_82_CARRYB_4__33_) );
  NAND2_X1 u5_mult_82_U9657 ( .A1(u5_mult_82_ab_4__33_), .A2(
        u5_mult_82_SUMB_3__34_), .ZN(u5_mult_82_n4504) );
  NAND3_X2 u5_mult_82_U9656 ( .A1(u5_mult_82_n4500), .A2(u5_mult_82_n4501), 
        .A3(u5_mult_82_n4502), .ZN(u5_mult_82_CARRYB_3__34_) );
  NAND2_X2 u5_mult_82_U9655 ( .A1(u5_mult_82_CARRYB_2__34_), .A2(
        u5_mult_82_SUMB_2__35_), .ZN(u5_mult_82_n4502) );
  NAND2_X2 u5_mult_82_U9654 ( .A1(u5_mult_82_ab_3__34_), .A2(
        u5_mult_82_SUMB_2__35_), .ZN(u5_mult_82_n4501) );
  NAND2_X1 u5_mult_82_U9653 ( .A1(u5_mult_82_ab_3__34_), .A2(
        u5_mult_82_CARRYB_2__34_), .ZN(u5_mult_82_n4500) );
  XOR2_X2 u5_mult_82_U9652 ( .A(u5_mult_82_n4499), .B(u5_mult_82_SUMB_3__34_), 
        .Z(u5_mult_82_SUMB_4__33_) );
  XOR2_X2 u5_mult_82_U9651 ( .A(u5_mult_82_ab_4__33_), .B(
        u5_mult_82_CARRYB_3__33_), .Z(u5_mult_82_n4499) );
  XOR2_X2 u5_mult_82_U9650 ( .A(u5_mult_82_n4498), .B(u5_mult_82_SUMB_2__35_), 
        .Z(u5_mult_82_SUMB_3__34_) );
  XOR2_X2 u5_mult_82_U9649 ( .A(u5_mult_82_ab_3__34_), .B(
        u5_mult_82_CARRYB_2__34_), .Z(u5_mult_82_n4498) );
  NAND3_X2 u5_mult_82_U9648 ( .A1(u5_mult_82_n4495), .A2(u5_mult_82_n4496), 
        .A3(u5_mult_82_n4497), .ZN(u5_mult_82_CARRYB_2__35_) );
  NAND2_X2 u5_mult_82_U9647 ( .A1(u5_mult_82_ab_2__35_), .A2(u5_mult_82_n586), 
        .ZN(u5_mult_82_n4497) );
  NAND2_X2 u5_mult_82_U9646 ( .A1(u5_mult_82_ab_2__35_), .A2(
        u5_mult_82_SUMB_1__36_), .ZN(u5_mult_82_n4496) );
  NAND2_X2 u5_mult_82_U9645 ( .A1(u5_mult_82_n586), .A2(u5_mult_82_SUMB_1__36_), .ZN(u5_mult_82_n4495) );
  XOR2_X2 u5_mult_82_U9644 ( .A(u5_mult_82_SUMB_1__36_), .B(u5_mult_82_n4494), 
        .Z(u5_mult_82_SUMB_2__35_) );
  XOR2_X2 u5_mult_82_U9643 ( .A(u5_mult_82_n586), .B(u5_mult_82_ab_2__35_), 
        .Z(u5_mult_82_n4494) );
  NAND3_X2 u5_mult_82_U9642 ( .A1(u5_mult_82_n4491), .A2(u5_mult_82_n4492), 
        .A3(u5_mult_82_n4493), .ZN(u5_mult_82_CARRYB_13__24_) );
  NAND2_X1 u5_mult_82_U9641 ( .A1(u5_mult_82_CARRYB_12__24_), .A2(
        u5_mult_82_SUMB_12__25_), .ZN(u5_mult_82_n4493) );
  NAND2_X1 u5_mult_82_U9640 ( .A1(u5_mult_82_ab_13__24_), .A2(
        u5_mult_82_SUMB_12__25_), .ZN(u5_mult_82_n4492) );
  NAND2_X1 u5_mult_82_U9639 ( .A1(u5_mult_82_ab_13__24_), .A2(
        u5_mult_82_CARRYB_12__24_), .ZN(u5_mult_82_n4491) );
  NAND3_X2 u5_mult_82_U9638 ( .A1(u5_mult_82_n4490), .A2(u5_mult_82_n4489), 
        .A3(u5_mult_82_n4488), .ZN(u5_mult_82_CARRYB_12__25_) );
  NAND2_X2 u5_mult_82_U9637 ( .A1(u5_mult_82_CARRYB_11__25_), .A2(
        u5_mult_82_n1572), .ZN(u5_mult_82_n4490) );
  NAND2_X2 u5_mult_82_U9636 ( .A1(u5_mult_82_ab_12__25_), .A2(u5_mult_82_n1572), .ZN(u5_mult_82_n4489) );
  XOR2_X2 u5_mult_82_U9635 ( .A(u5_mult_82_n4487), .B(u5_mult_82_SUMB_12__25_), 
        .Z(u5_mult_82_SUMB_13__24_) );
  XOR2_X2 u5_mult_82_U9634 ( .A(u5_mult_82_n4486), .B(u5_mult_82_n1572), .Z(
        u5_mult_82_SUMB_12__25_) );
  XOR2_X2 u5_mult_82_U9633 ( .A(u5_mult_82_ab_12__25_), .B(
        u5_mult_82_CARRYB_11__25_), .Z(u5_mult_82_n4486) );
  XNOR2_X2 u5_mult_82_U9632 ( .A(u5_mult_82_n4485), .B(
        u5_mult_82_CARRYB_48__24_), .ZN(u5_mult_82_n4576) );
  NAND3_X4 u5_mult_82_U9631 ( .A1(u5_mult_82_n6319), .A2(u5_mult_82_n6320), 
        .A3(u5_mult_82_n6321), .ZN(u5_mult_82_CARRYB_6__47_) );
  NAND3_X2 u5_mult_82_U9630 ( .A1(u5_mult_82_n4482), .A2(u5_mult_82_n4483), 
        .A3(u5_mult_82_n4484), .ZN(u5_mult_82_CARRYB_33__42_) );
  NAND2_X1 u5_mult_82_U9629 ( .A1(u5_mult_82_CARRYB_32__42_), .A2(
        u5_mult_82_SUMB_32__43_), .ZN(u5_mult_82_n4484) );
  NAND2_X1 u5_mult_82_U9628 ( .A1(u5_mult_82_ab_33__42_), .A2(
        u5_mult_82_SUMB_32__43_), .ZN(u5_mult_82_n4483) );
  NAND2_X1 u5_mult_82_U9627 ( .A1(u5_mult_82_ab_33__42_), .A2(
        u5_mult_82_CARRYB_32__42_), .ZN(u5_mult_82_n4482) );
  NAND3_X2 u5_mult_82_U9626 ( .A1(u5_mult_82_n4479), .A2(u5_mult_82_n4480), 
        .A3(u5_mult_82_n4481), .ZN(u5_mult_82_CARRYB_32__43_) );
  NAND2_X2 u5_mult_82_U9625 ( .A1(u5_mult_82_CARRYB_31__43_), .A2(
        u5_mult_82_SUMB_31__44_), .ZN(u5_mult_82_n4481) );
  NAND2_X2 u5_mult_82_U9624 ( .A1(u5_mult_82_ab_32__43_), .A2(
        u5_mult_82_SUMB_31__44_), .ZN(u5_mult_82_n4480) );
  NAND2_X1 u5_mult_82_U9623 ( .A1(u5_mult_82_ab_32__43_), .A2(
        u5_mult_82_CARRYB_31__43_), .ZN(u5_mult_82_n4479) );
  XOR2_X2 u5_mult_82_U9622 ( .A(u5_mult_82_n4478), .B(u5_mult_82_SUMB_31__44_), 
        .Z(u5_mult_82_SUMB_32__43_) );
  XOR2_X2 u5_mult_82_U9621 ( .A(u5_mult_82_CARRYB_31__43_), .B(
        u5_mult_82_ab_32__43_), .Z(u5_mult_82_n4478) );
  NAND3_X2 u5_mult_82_U9620 ( .A1(u5_mult_82_n4475), .A2(u5_mult_82_n4476), 
        .A3(u5_mult_82_n4477), .ZN(u5_mult_82_CARRYB_39__36_) );
  NAND2_X1 u5_mult_82_U9619 ( .A1(u5_mult_82_CARRYB_38__36_), .A2(
        u5_mult_82_SUMB_38__37_), .ZN(u5_mult_82_n4477) );
  NAND2_X1 u5_mult_82_U9618 ( .A1(u5_mult_82_ab_39__36_), .A2(
        u5_mult_82_SUMB_38__37_), .ZN(u5_mult_82_n4476) );
  NAND2_X1 u5_mult_82_U9617 ( .A1(u5_mult_82_ab_39__36_), .A2(
        u5_mult_82_CARRYB_38__36_), .ZN(u5_mult_82_n4475) );
  NAND2_X2 u5_mult_82_U9616 ( .A1(u5_mult_82_CARRYB_37__37_), .A2(
        u5_mult_82_SUMB_37__38_), .ZN(u5_mult_82_n4474) );
  NAND2_X2 u5_mult_82_U9615 ( .A1(u5_mult_82_ab_38__37_), .A2(
        u5_mult_82_SUMB_37__38_), .ZN(u5_mult_82_n4473) );
  XOR2_X2 u5_mult_82_U9614 ( .A(u5_mult_82_n4470), .B(u5_mult_82_SUMB_37__38_), 
        .Z(u5_mult_82_SUMB_38__37_) );
  NAND3_X2 u5_mult_82_U9613 ( .A1(u5_mult_82_n4467), .A2(u5_mult_82_n4468), 
        .A3(u5_mult_82_n4469), .ZN(u5_mult_82_CARRYB_51__24_) );
  NAND2_X1 u5_mult_82_U9612 ( .A1(u5_mult_82_ab_51__24_), .A2(
        u5_mult_82_SUMB_50__25_), .ZN(u5_mult_82_n4468) );
  NAND2_X2 u5_mult_82_U9611 ( .A1(u5_mult_82_CARRYB_49__25_), .A2(
        u5_mult_82_SUMB_49__26_), .ZN(u5_mult_82_n4466) );
  NAND2_X2 u5_mult_82_U9610 ( .A1(u5_mult_82_ab_50__25_), .A2(
        u5_mult_82_SUMB_49__26_), .ZN(u5_mult_82_n4465) );
  NAND2_X1 u5_mult_82_U9609 ( .A1(u5_mult_82_ab_50__25_), .A2(
        u5_mult_82_CARRYB_49__25_), .ZN(u5_mult_82_n4464) );
  XOR2_X2 u5_mult_82_U9608 ( .A(u5_mult_82_n4463), .B(u5_mult_82_SUMB_50__25_), 
        .Z(u5_mult_82_SUMB_51__24_) );
  XOR2_X2 u5_mult_82_U9607 ( .A(u5_mult_82_n4462), .B(u5_mult_82_SUMB_49__26_), 
        .Z(u5_mult_82_SUMB_50__25_) );
  NOR2_X1 u5_mult_82_U9606 ( .A1(u5_mult_82_n6768), .A2(u5_mult_82_n6607), 
        .ZN(u5_mult_82_ab_18__50_) );
  NOR2_X1 u5_mult_82_U9605 ( .A1(u5_mult_82_net64683), .A2(u5_mult_82_net65191), .ZN(u5_mult_82_ab_51__23_) );
  NAND3_X2 u5_mult_82_U9604 ( .A1(u5_mult_82_n4459), .A2(u5_mult_82_n4460), 
        .A3(u5_mult_82_n4461), .ZN(u5_mult_82_CARRYB_18__50_) );
  NAND2_X2 u5_mult_82_U9603 ( .A1(u5_mult_82_ab_18__50_), .A2(
        u5_mult_82_SUMB_17__51_), .ZN(u5_mult_82_n4461) );
  NAND2_X2 u5_mult_82_U9602 ( .A1(u5_mult_82_ab_18__50_), .A2(
        u5_mult_82_CARRYB_17__50_), .ZN(u5_mult_82_n4460) );
  NAND3_X2 u5_mult_82_U9601 ( .A1(u5_mult_82_n4456), .A2(u5_mult_82_n4457), 
        .A3(u5_mult_82_n4458), .ZN(u5_mult_82_CARRYB_51__23_) );
  NAND2_X1 u5_mult_82_U9600 ( .A1(u5_mult_82_ab_51__23_), .A2(
        u5_mult_82_SUMB_50__24_), .ZN(u5_mult_82_n4458) );
  NAND2_X2 u5_mult_82_U9599 ( .A1(u5_mult_82_ab_51__23_), .A2(
        u5_mult_82_CARRYB_50__23_), .ZN(u5_mult_82_n4457) );
  NAND3_X2 u5_mult_82_U9598 ( .A1(u5_mult_82_n4453), .A2(u5_mult_82_n4454), 
        .A3(u5_mult_82_n4455), .ZN(u5_mult_82_CARRYB_40__34_) );
  NAND2_X1 u5_mult_82_U9597 ( .A1(u5_mult_82_CARRYB_39__34_), .A2(
        u5_mult_82_SUMB_39__35_), .ZN(u5_mult_82_n4455) );
  NAND2_X1 u5_mult_82_U9596 ( .A1(u5_mult_82_ab_40__34_), .A2(
        u5_mult_82_SUMB_39__35_), .ZN(u5_mult_82_n4454) );
  NAND2_X1 u5_mult_82_U9595 ( .A1(u5_mult_82_ab_40__34_), .A2(
        u5_mult_82_CARRYB_39__34_), .ZN(u5_mult_82_n4453) );
  NAND3_X2 u5_mult_82_U9594 ( .A1(u5_mult_82_n4450), .A2(u5_mult_82_n4451), 
        .A3(u5_mult_82_n4452), .ZN(u5_mult_82_CARRYB_39__35_) );
  NAND2_X2 u5_mult_82_U9593 ( .A1(u5_mult_82_CARRYB_38__35_), .A2(
        u5_mult_82_n3472), .ZN(u5_mult_82_n4452) );
  NAND2_X2 u5_mult_82_U9592 ( .A1(u5_mult_82_ab_39__35_), .A2(u5_mult_82_n3472), .ZN(u5_mult_82_n4451) );
  NAND2_X1 u5_mult_82_U9591 ( .A1(u5_mult_82_ab_39__35_), .A2(
        u5_mult_82_CARRYB_38__35_), .ZN(u5_mult_82_n4450) );
  XOR2_X2 u5_mult_82_U9590 ( .A(u5_mult_82_ab_40__34_), .B(
        u5_mult_82_CARRYB_39__34_), .Z(u5_mult_82_n4449) );
  XOR2_X2 u5_mult_82_U9589 ( .A(u5_mult_82_n4448), .B(u5_mult_82_n3472), .Z(
        u5_mult_82_SUMB_39__35_) );
  XOR2_X2 u5_mult_82_U9588 ( .A(u5_mult_82_ab_39__35_), .B(
        u5_mult_82_CARRYB_38__35_), .Z(u5_mult_82_n4448) );
  NAND2_X1 u5_mult_82_U9587 ( .A1(u5_mult_82_ab_50__24_), .A2(
        u5_mult_82_CARRYB_49__24_), .ZN(u5_mult_82_n4445) );
  NAND2_X2 u5_mult_82_U9586 ( .A1(u5_mult_82_CARRYB_48__25_), .A2(
        u5_mult_82_n1663), .ZN(u5_mult_82_n4444) );
  NAND2_X2 u5_mult_82_U9585 ( .A1(u5_mult_82_ab_49__25_), .A2(u5_mult_82_n1663), .ZN(u5_mult_82_n4443) );
  NAND2_X2 u5_mult_82_U9584 ( .A1(u5_mult_82_ab_49__25_), .A2(
        u5_mult_82_CARRYB_48__25_), .ZN(u5_mult_82_n4442) );
  INV_X4 u5_mult_82_U9583 ( .A(u5_mult_82_n6801), .ZN(u5_mult_82_n6800) );
  NAND2_X1 u5_mult_82_U9582 ( .A1(u5_mult_82_CARRYB_14__29_), .A2(
        u5_mult_82_SUMB_14__30_), .ZN(u5_mult_82_n5338) );
  INV_X16 u5_mult_82_U9581 ( .A(u5_mult_82_n7008), .ZN(u5_mult_82_n6801) );
  NAND3_X4 u5_mult_82_U9580 ( .A1(u5_mult_82_n5764), .A2(u5_mult_82_n5765), 
        .A3(u5_mult_82_n5766), .ZN(u5_mult_82_CARRYB_25__34_) );
  NOR2_X1 u5_mult_82_U9579 ( .A1(u5_mult_82_net64885), .A2(u5_mult_82_n6649), 
        .ZN(u5_mult_82_ab_26__34_) );
  NAND2_X1 u5_mult_82_U9578 ( .A1(u5_mult_82_ab_26__34_), .A2(
        u5_mult_82_CARRYB_25__34_), .ZN(u5_mult_82_n4441) );
  INV_X4 u5_mult_82_U9577 ( .A(u5_mult_82_n4853), .ZN(u5_mult_82_n4436) );
  NAND2_X4 u5_mult_82_U9576 ( .A1(u5_mult_82_n4437), .A2(u5_mult_82_n4438), 
        .ZN(u5_mult_82_SUMB_30__32_) );
  NAND2_X4 u5_mult_82_U9575 ( .A1(u5_mult_82_n4436), .A2(u5_mult_82_n79), .ZN(
        u5_mult_82_n4438) );
  NAND2_X2 u5_mult_82_U9574 ( .A1(u5_mult_82_n4853), .A2(
        u5_mult_82_SUMB_29__33_), .ZN(u5_mult_82_n4437) );
  NAND2_X2 u5_mult_82_U9573 ( .A1(u5_mult_82_ab_19__29_), .A2(
        u5_mult_82_SUMB_18__30_), .ZN(u5_mult_82_n6016) );
  NAND2_X1 u5_mult_82_U9572 ( .A1(u5_mult_82_CARRYB_40__5_), .A2(
        u5_mult_82_SUMB_40__6_), .ZN(u5_mult_82_n4728) );
  XNOR2_X2 u5_mult_82_U9571 ( .A(u5_mult_82_CARRYB_36__16_), .B(
        u5_mult_82_ab_37__16_), .ZN(u5_mult_82_n4435) );
  XNOR2_X2 u5_mult_82_U9570 ( .A(u5_mult_82_n738), .B(u5_mult_82_n4435), .ZN(
        u5_mult_82_SUMB_37__16_) );
  NOR2_X1 u5_mult_82_U9569 ( .A1(u5_mult_82_net64683), .A2(u5_mult_82_n6749), 
        .ZN(u5_mult_82_ab_48__23_) );
  NAND3_X2 u5_mult_82_U9568 ( .A1(u5_mult_82_n4432), .A2(u5_mult_82_n4433), 
        .A3(u5_mult_82_n4434), .ZN(u5_mult_82_CARRYB_48__23_) );
  NAND2_X1 u5_mult_82_U9567 ( .A1(u5_mult_82_ab_48__23_), .A2(
        u5_mult_82_CARRYB_47__23_), .ZN(u5_mult_82_n4434) );
  NAND2_X2 u5_mult_82_U9566 ( .A1(u5_mult_82_ab_48__23_), .A2(
        u5_mult_82_SUMB_47__24_), .ZN(u5_mult_82_n4433) );
  NAND2_X1 u5_mult_82_U9565 ( .A1(u5_mult_82_CARRYB_47__23_), .A2(
        u5_mult_82_SUMB_47__24_), .ZN(u5_mult_82_n4432) );
  NAND2_X1 u5_mult_82_U9564 ( .A1(u5_mult_82_CARRYB_17__47_), .A2(
        u5_mult_82_SUMB_17__48_), .ZN(u5_mult_82_n4431) );
  NAND2_X1 u5_mult_82_U9563 ( .A1(u5_mult_82_ab_18__47_), .A2(
        u5_mult_82_SUMB_17__48_), .ZN(u5_mult_82_n4430) );
  NAND2_X1 u5_mult_82_U9562 ( .A1(u5_mult_82_ab_18__47_), .A2(
        u5_mult_82_CARRYB_17__47_), .ZN(u5_mult_82_n4429) );
  NAND3_X2 u5_mult_82_U9561 ( .A1(u5_mult_82_n4426), .A2(u5_mult_82_n4427), 
        .A3(u5_mult_82_n4428), .ZN(u5_mult_82_CARRYB_17__48_) );
  NAND2_X2 u5_mult_82_U9560 ( .A1(u5_mult_82_ab_17__48_), .A2(
        u5_mult_82_SUMB_16__49_), .ZN(u5_mult_82_n4427) );
  XOR2_X2 u5_mult_82_U9559 ( .A(u5_mult_82_n4425), .B(u5_mult_82_SUMB_16__49_), 
        .Z(u5_mult_82_SUMB_17__48_) );
  NAND3_X2 u5_mult_82_U9558 ( .A1(u5_mult_82_n4422), .A2(u5_mult_82_n4423), 
        .A3(u5_mult_82_n4424), .ZN(u5_mult_82_CARRYB_42__29_) );
  NAND2_X1 u5_mult_82_U9557 ( .A1(u5_mult_82_CARRYB_41__29_), .A2(
        u5_mult_82_SUMB_41__30_), .ZN(u5_mult_82_n4424) );
  NAND2_X1 u5_mult_82_U9556 ( .A1(u5_mult_82_ab_42__29_), .A2(
        u5_mult_82_CARRYB_41__29_), .ZN(u5_mult_82_n4422) );
  NAND2_X2 u5_mult_82_U9555 ( .A1(u5_mult_82_CARRYB_40__30_), .A2(
        u5_mult_82_SUMB_40__31_), .ZN(u5_mult_82_n4421) );
  NAND2_X2 u5_mult_82_U9554 ( .A1(u5_mult_82_ab_41__30_), .A2(
        u5_mult_82_SUMB_40__31_), .ZN(u5_mult_82_n4420) );
  NAND2_X1 u5_mult_82_U9553 ( .A1(u5_mult_82_ab_41__30_), .A2(
        u5_mult_82_CARRYB_40__30_), .ZN(u5_mult_82_n4419) );
  NOR2_X1 u5_mult_82_U9552 ( .A1(u5_mult_82_n6813), .A2(u5_mult_82_n6513), 
        .ZN(u5_mult_82_ab_3__43_) );
  NAND3_X2 u5_mult_82_U9551 ( .A1(u5_mult_82_n4415), .A2(u5_mult_82_n4416), 
        .A3(u5_mult_82_n4417), .ZN(u5_mult_82_CARRYB_3__43_) );
  NAND2_X1 u5_mult_82_U9550 ( .A1(u5_mult_82_ab_3__43_), .A2(
        u5_mult_82_CARRYB_2__43_), .ZN(u5_mult_82_n4417) );
  NAND2_X2 u5_mult_82_U9549 ( .A1(u5_mult_82_ab_3__43_), .A2(
        u5_mult_82_SUMB_2__44_), .ZN(u5_mult_82_n4416) );
  NAND2_X1 u5_mult_82_U9548 ( .A1(u5_mult_82_CARRYB_2__43_), .A2(
        u5_mult_82_SUMB_2__44_), .ZN(u5_mult_82_n4415) );
  AND2_X2 u5_mult_82_U9547 ( .A1(u5_mult_82_net86084), .A2(n4783), .ZN(
        u5_mult_82_n4414) );
  NAND2_X2 u5_mult_82_U9546 ( .A1(u5_mult_82_CARRYB_18__38_), .A2(
        u5_mult_82_SUMB_18__39_), .ZN(u5_mult_82_n4413) );
  NAND2_X2 u5_mult_82_U9545 ( .A1(u5_mult_82_ab_19__38_), .A2(
        u5_mult_82_SUMB_18__39_), .ZN(u5_mult_82_n4412) );
  NAND2_X1 u5_mult_82_U9544 ( .A1(u5_mult_82_ab_19__38_), .A2(
        u5_mult_82_CARRYB_18__38_), .ZN(u5_mult_82_n4411) );
  NAND3_X2 u5_mult_82_U9543 ( .A1(u5_mult_82_n4408), .A2(u5_mult_82_n4409), 
        .A3(u5_mult_82_n4410), .ZN(u5_mult_82_CARRYB_18__39_) );
  NAND2_X2 u5_mult_82_U9542 ( .A1(u5_mult_82_ab_18__39_), .A2(
        u5_mult_82_CARRYB_17__39_), .ZN(u5_mult_82_n4408) );
  NAND3_X2 u5_mult_82_U9541 ( .A1(u5_mult_82_n4405), .A2(u5_mult_82_n4406), 
        .A3(u5_mult_82_n4407), .ZN(u5_mult_82_CARRYB_27__34_) );
  NAND2_X1 u5_mult_82_U9540 ( .A1(u5_mult_82_CARRYB_26__34_), .A2(
        u5_mult_82_SUMB_26__35_), .ZN(u5_mult_82_n4407) );
  NAND2_X1 u5_mult_82_U9539 ( .A1(u5_mult_82_ab_27__34_), .A2(
        u5_mult_82_SUMB_26__35_), .ZN(u5_mult_82_n4406) );
  NAND2_X1 u5_mult_82_U9538 ( .A1(u5_mult_82_ab_27__34_), .A2(
        u5_mult_82_CARRYB_26__34_), .ZN(u5_mult_82_n4405) );
  NAND3_X2 u5_mult_82_U9537 ( .A1(u5_mult_82_n4402), .A2(u5_mult_82_n4403), 
        .A3(u5_mult_82_n4404), .ZN(u5_mult_82_CARRYB_26__35_) );
  NAND2_X2 u5_mult_82_U9536 ( .A1(u5_mult_82_SUMB_25__36_), .A2(
        u5_mult_82_CARRYB_25__35_), .ZN(u5_mult_82_n4404) );
  NAND2_X2 u5_mult_82_U9535 ( .A1(u5_mult_82_ab_26__35_), .A2(
        u5_mult_82_SUMB_25__36_), .ZN(u5_mult_82_n4403) );
  XOR2_X2 u5_mult_82_U9534 ( .A(u5_mult_82_n4401), .B(u5_mult_82_n1672), .Z(
        u5_mult_82_SUMB_26__35_) );
  XOR2_X2 u5_mult_82_U9533 ( .A(u5_mult_82_CARRYB_25__35_), .B(
        u5_mult_82_ab_26__35_), .Z(u5_mult_82_n4401) );
  NAND3_X4 u5_mult_82_U9532 ( .A1(u5_mult_82_n4395), .A2(u5_mult_82_n4396), 
        .A3(u5_mult_82_n4397), .ZN(u5_mult_82_CARRYB_49__18_) );
  NAND2_X2 u5_mult_82_U9531 ( .A1(u5_mult_82_CARRYB_48__18_), .A2(
        u5_mult_82_SUMB_48__19_), .ZN(u5_mult_82_n4397) );
  NAND2_X2 u5_mult_82_U9530 ( .A1(u5_mult_82_ab_49__18_), .A2(
        u5_mult_82_SUMB_48__19_), .ZN(u5_mult_82_n4396) );
  XOR2_X2 u5_mult_82_U9529 ( .A(u5_mult_82_ab_50__17_), .B(
        u5_mult_82_CARRYB_49__17_), .Z(u5_mult_82_n4394) );
  NAND3_X2 u5_mult_82_U9528 ( .A1(u5_mult_82_n4391), .A2(u5_mult_82_n4392), 
        .A3(u5_mult_82_n4393), .ZN(u5_mult_82_CARRYB_48__19_) );
  NAND2_X1 u5_mult_82_U9527 ( .A1(u5_mult_82_ab_48__19_), .A2(
        u5_mult_82_CARRYB_47__19_), .ZN(u5_mult_82_n4391) );
  NAND2_X2 u5_mult_82_U9526 ( .A1(u5_mult_82_n1719), .A2(u5_mult_82_n1863), 
        .ZN(u5_mult_82_n4390) );
  NAND2_X2 u5_mult_82_U9525 ( .A1(u5_mult_82_ab_47__20_), .A2(u5_mult_82_n1863), .ZN(u5_mult_82_n4389) );
  NAND2_X1 u5_mult_82_U9524 ( .A1(u5_mult_82_ab_47__20_), .A2(
        u5_mult_82_CARRYB_46__20_), .ZN(u5_mult_82_n4388) );
  NOR2_X1 u5_mult_82_U9523 ( .A1(u5_mult_82_net64415), .A2(u5_mult_82_net65373), .ZN(u5_mult_82_ab_42__8_) );
  NOR2_X1 u5_mult_82_U9522 ( .A1(u5_mult_82_net64379), .A2(u5_mult_82_n6748), 
        .ZN(u5_mult_82_ab_48__6_) );
  NOR2_X2 u5_mult_82_U9521 ( .A1(u5_mult_82_n6882), .A2(u5_mult_82_n6551), 
        .ZN(u5_mult_82_ab_10__26_) );
  NAND2_X1 u5_mult_82_U9520 ( .A1(u5_mult_82_ab_42__8_), .A2(
        u5_mult_82_SUMB_41__9_), .ZN(u5_mult_82_n4387) );
  NAND2_X1 u5_mult_82_U9519 ( .A1(u5_mult_82_SUMB_41__9_), .A2(
        u5_mult_82_CARRYB_41__8_), .ZN(u5_mult_82_n4385) );
  NAND2_X1 u5_mult_82_U9518 ( .A1(u5_mult_82_ab_48__6_), .A2(
        u5_mult_82_CARRYB_47__6_), .ZN(u5_mult_82_n4383) );
  NAND2_X2 u5_mult_82_U9517 ( .A1(u5_mult_82_ab_48__6_), .A2(
        u5_mult_82_SUMB_47__7_), .ZN(u5_mult_82_n4382) );
  XOR2_X2 u5_mult_82_U9516 ( .A(u5_mult_82_SUMB_47__7_), .B(u5_mult_82_n4380), 
        .Z(u5_mult_82_SUMB_48__6_) );
  XOR2_X2 u5_mult_82_U9515 ( .A(u5_mult_82_CARRYB_47__6_), .B(
        u5_mult_82_ab_48__6_), .Z(u5_mult_82_n4380) );
  NAND3_X2 u5_mult_82_U9514 ( .A1(u5_mult_82_n4377), .A2(u5_mult_82_n4378), 
        .A3(u5_mult_82_n4379), .ZN(u5_mult_82_CARRYB_46__7_) );
  NAND2_X2 u5_mult_82_U9513 ( .A1(u5_mult_82_ab_46__7_), .A2(
        u5_mult_82_CARRYB_45__7_), .ZN(u5_mult_82_n4378) );
  NAND3_X2 u5_mult_82_U9512 ( .A1(u5_mult_82_n4374), .A2(u5_mult_82_n4375), 
        .A3(u5_mult_82_n4376), .ZN(u5_mult_82_CARRYB_45__7_) );
  NAND2_X1 u5_mult_82_U9511 ( .A1(u5_mult_82_CARRYB_44__7_), .A2(
        u5_mult_82_SUMB_44__8_), .ZN(u5_mult_82_n4376) );
  NAND2_X2 u5_mult_82_U9510 ( .A1(u5_mult_82_ab_45__7_), .A2(
        u5_mult_82_SUMB_44__8_), .ZN(u5_mult_82_n4375) );
  NAND2_X1 u5_mult_82_U9509 ( .A1(u5_mult_82_ab_45__7_), .A2(
        u5_mult_82_CARRYB_44__7_), .ZN(u5_mult_82_n4374) );
  NAND3_X2 u5_mult_82_U9508 ( .A1(u5_mult_82_n4371), .A2(u5_mult_82_n4372), 
        .A3(u5_mult_82_n4373), .ZN(u5_mult_82_CARRYB_10__26_) );
  NAND2_X1 u5_mult_82_U9507 ( .A1(u5_mult_82_ab_10__26_), .A2(
        u5_mult_82_CARRYB_9__26_), .ZN(u5_mult_82_n4373) );
  NAND2_X2 u5_mult_82_U9506 ( .A1(u5_mult_82_ab_10__26_), .A2(u5_mult_82_n382), 
        .ZN(u5_mult_82_n4372) );
  NAND3_X2 u5_mult_82_U9505 ( .A1(u5_mult_82_n4368), .A2(u5_mult_82_n4369), 
        .A3(u5_mult_82_n4370), .ZN(u5_mult_82_CARRYB_18__20_) );
  NAND2_X1 u5_mult_82_U9504 ( .A1(u5_mult_82_ab_18__20_), .A2(
        u5_mult_82_SUMB_17__21_), .ZN(u5_mult_82_n4369) );
  NAND3_X2 u5_mult_82_U9503 ( .A1(u5_mult_82_n4365), .A2(u5_mult_82_n4366), 
        .A3(u5_mult_82_n4367), .ZN(u5_mult_82_CARRYB_17__21_) );
  NAND2_X2 u5_mult_82_U9502 ( .A1(u5_mult_82_CARRYB_16__21_), .A2(
        u5_mult_82_SUMB_16__22_), .ZN(u5_mult_82_n4367) );
  NAND2_X2 u5_mult_82_U9501 ( .A1(u5_mult_82_ab_17__21_), .A2(
        u5_mult_82_SUMB_16__22_), .ZN(u5_mult_82_n4366) );
  NAND2_X1 u5_mult_82_U9500 ( .A1(u5_mult_82_ab_17__21_), .A2(
        u5_mult_82_CARRYB_16__21_), .ZN(u5_mult_82_n4365) );
  XOR2_X2 u5_mult_82_U9499 ( .A(u5_mult_82_n4364), .B(u5_mult_82_SUMB_16__22_), 
        .Z(u5_mult_82_SUMB_17__21_) );
  XOR2_X2 u5_mult_82_U9498 ( .A(u5_mult_82_ab_17__21_), .B(
        u5_mult_82_CARRYB_16__21_), .Z(u5_mult_82_n4364) );
  NAND3_X4 u5_mult_82_U9497 ( .A1(u5_mult_82_net79785), .A2(
        u5_mult_82_net79786), .A3(u5_mult_82_n5606), .ZN(
        u5_mult_82_CARRYB_17__27_) );
  XOR2_X2 u5_mult_82_U9496 ( .A(u5_mult_82_SUMB_14__50_), .B(
        u5_mult_82_ab_15__49_), .Z(u5_mult_82_n4717) );
  NAND2_X2 u5_mult_82_U9495 ( .A1(u5_mult_82_SUMB_36__18_), .A2(
        u5_mult_82_CARRYB_36__17_), .ZN(u5_mult_82_n5967) );
  NAND2_X2 u5_mult_82_U9494 ( .A1(u5_mult_82_CARRYB_22__17_), .A2(
        u5_mult_82_SUMB_22__18_), .ZN(u5_mult_82_n4732) );
  NAND2_X2 u5_mult_82_U9493 ( .A1(u5_mult_82_SUMB_6__50_), .A2(
        u5_mult_82_CARRYB_6__49_), .ZN(u5_mult_82_n5094) );
  XNOR2_X2 u5_mult_82_U9492 ( .A(u5_mult_82_CARRYB_45__14_), .B(
        u5_mult_82_ab_46__14_), .ZN(u5_mult_82_n4363) );
  XNOR2_X2 u5_mult_82_U9491 ( .A(u5_mult_82_SUMB_45__15_), .B(u5_mult_82_n4363), .ZN(u5_mult_82_SUMB_46__14_) );
  XOR2_X2 u5_mult_82_U9490 ( .A(u5_mult_82_ab_13__24_), .B(
        u5_mult_82_CARRYB_12__24_), .Z(u5_mult_82_n4487) );
  NAND3_X2 u5_mult_82_U9489 ( .A1(u5_mult_82_n5538), .A2(u5_mult_82_n5539), 
        .A3(u5_mult_82_n5540), .ZN(u5_mult_82_CARRYB_28__23_) );
  NAND2_X2 u5_mult_82_U9488 ( .A1(u5_mult_82_CARRYB_44__12_), .A2(
        u5_mult_82_n3709), .ZN(u5_mult_82_n5678) );
  XNOR2_X2 u5_mult_82_U9487 ( .A(u5_mult_82_ab_25__25_), .B(
        u5_mult_82_CARRYB_24__25_), .ZN(u5_mult_82_n4361) );
  XNOR2_X2 u5_mult_82_U9486 ( .A(u5_mult_82_n4361), .B(u5_mult_82_SUMB_24__26_), .ZN(u5_mult_82_SUMB_25__25_) );
  XNOR2_X2 u5_mult_82_U9485 ( .A(u5_mult_82_ab_50__14_), .B(
        u5_mult_82_CARRYB_49__14_), .ZN(u5_mult_82_n4362) );
  NOR2_X2 u5_mult_82_U9484 ( .A1(u5_mult_82_net64559), .A2(u5_mult_82_n6685), 
        .ZN(u5_mult_82_ab_31__16_) );
  NAND3_X2 u5_mult_82_U9483 ( .A1(u5_mult_82_n4357), .A2(u5_mult_82_n4359), 
        .A3(u5_mult_82_n4358), .ZN(u5_mult_82_CARRYB_31__16_) );
  NAND2_X1 u5_mult_82_U9482 ( .A1(u5_mult_82_SUMB_30__17_), .A2(
        u5_mult_82_CARRYB_30__16_), .ZN(u5_mult_82_n4357) );
  NAND3_X2 u5_mult_82_U9481 ( .A1(u5_mult_82_n4354), .A2(u5_mult_82_n4355), 
        .A3(u5_mult_82_n4356), .ZN(u5_mult_82_CARRYB_11__27_) );
  NAND2_X1 u5_mult_82_U9480 ( .A1(u5_mult_82_CARRYB_10__27_), .A2(
        u5_mult_82_SUMB_10__28_), .ZN(u5_mult_82_n4356) );
  NAND2_X1 u5_mult_82_U9479 ( .A1(u5_mult_82_ab_11__27_), .A2(
        u5_mult_82_SUMB_10__28_), .ZN(u5_mult_82_n4355) );
  NAND2_X1 u5_mult_82_U9478 ( .A1(u5_mult_82_ab_11__27_), .A2(
        u5_mult_82_CARRYB_10__27_), .ZN(u5_mult_82_n4354) );
  NAND3_X2 u5_mult_82_U9477 ( .A1(u5_mult_82_n4351), .A2(u5_mult_82_n4352), 
        .A3(u5_mult_82_n4353), .ZN(u5_mult_82_CARRYB_10__28_) );
  NAND2_X2 u5_mult_82_U9476 ( .A1(u5_mult_82_CARRYB_9__28_), .A2(
        u5_mult_82_SUMB_9__29_), .ZN(u5_mult_82_n4353) );
  NAND2_X2 u5_mult_82_U9475 ( .A1(u5_mult_82_ab_10__28_), .A2(
        u5_mult_82_SUMB_9__29_), .ZN(u5_mult_82_n4352) );
  NAND2_X1 u5_mult_82_U9474 ( .A1(u5_mult_82_ab_10__28_), .A2(
        u5_mult_82_CARRYB_9__28_), .ZN(u5_mult_82_n4351) );
  XOR2_X2 u5_mult_82_U9473 ( .A(u5_mult_82_n4350), .B(u5_mult_82_SUMB_10__28_), 
        .Z(u5_mult_82_SUMB_11__27_) );
  XOR2_X2 u5_mult_82_U9472 ( .A(u5_mult_82_ab_11__27_), .B(
        u5_mult_82_CARRYB_10__27_), .Z(u5_mult_82_n4350) );
  XOR2_X2 u5_mult_82_U9471 ( .A(u5_mult_82_n4349), .B(u5_mult_82_SUMB_9__29_), 
        .Z(u5_mult_82_SUMB_10__28_) );
  XOR2_X2 u5_mult_82_U9470 ( .A(u5_mult_82_ab_10__28_), .B(
        u5_mult_82_CARRYB_9__28_), .Z(u5_mult_82_n4349) );
  NAND3_X2 u5_mult_82_U9469 ( .A1(u5_mult_82_n4346), .A2(u5_mult_82_n4347), 
        .A3(u5_mult_82_n4348), .ZN(u5_mult_82_CARRYB_7__31_) );
  NAND2_X1 u5_mult_82_U9468 ( .A1(u5_mult_82_CARRYB_6__31_), .A2(
        u5_mult_82_SUMB_6__32_), .ZN(u5_mult_82_n4348) );
  NAND2_X1 u5_mult_82_U9467 ( .A1(u5_mult_82_ab_7__31_), .A2(
        u5_mult_82_SUMB_6__32_), .ZN(u5_mult_82_n4347) );
  NAND2_X1 u5_mult_82_U9466 ( .A1(u5_mult_82_ab_7__31_), .A2(
        u5_mult_82_CARRYB_6__31_), .ZN(u5_mult_82_n4346) );
  NAND3_X2 u5_mult_82_U9465 ( .A1(u5_mult_82_n4343), .A2(u5_mult_82_n4344), 
        .A3(u5_mult_82_n4345), .ZN(u5_mult_82_CARRYB_6__32_) );
  NAND2_X2 u5_mult_82_U9464 ( .A1(u5_mult_82_CARRYB_5__32_), .A2(
        u5_mult_82_SUMB_5__33_), .ZN(u5_mult_82_n4345) );
  NAND2_X2 u5_mult_82_U9463 ( .A1(u5_mult_82_ab_6__32_), .A2(
        u5_mult_82_SUMB_5__33_), .ZN(u5_mult_82_n4344) );
  NAND2_X1 u5_mult_82_U9462 ( .A1(u5_mult_82_ab_6__32_), .A2(
        u5_mult_82_CARRYB_5__32_), .ZN(u5_mult_82_n4343) );
  XOR2_X2 u5_mult_82_U9461 ( .A(u5_mult_82_n4342), .B(u5_mult_82_SUMB_5__33_), 
        .Z(u5_mult_82_SUMB_6__32_) );
  XOR2_X2 u5_mult_82_U9460 ( .A(u5_mult_82_ab_6__32_), .B(
        u5_mult_82_CARRYB_5__32_), .Z(u5_mult_82_n4342) );
  NAND2_X2 u5_mult_82_U9459 ( .A1(u5_mult_82_ab_48__8_), .A2(
        u5_mult_82_SUMB_47__9_), .ZN(u5_mult_82_n4341) );
  XNOR2_X2 u5_mult_82_U9458 ( .A(u5_mult_82_ab_50__24_), .B(
        u5_mult_82_CARRYB_49__24_), .ZN(u5_mult_82_n4340) );
  XNOR2_X2 u5_mult_82_U9457 ( .A(u5_mult_82_n4340), .B(u5_mult_82_SUMB_49__25_), .ZN(u5_mult_82_SUMB_50__24_) );
  XNOR2_X2 u5_mult_82_U9456 ( .A(u5_mult_82_ab_47__15_), .B(
        u5_mult_82_CARRYB_46__15_), .ZN(u5_mult_82_n4339) );
  XNOR2_X2 u5_mult_82_U9455 ( .A(u5_mult_82_n4339), .B(u5_mult_82_SUMB_46__16_), .ZN(u5_mult_82_SUMB_47__15_) );
  NOR2_X1 u5_mult_82_U9454 ( .A1(u5_mult_82_n6775), .A2(u5_mult_82_n6550), 
        .ZN(u5_mult_82_ab_10__49_) );
  NOR2_X2 u5_mult_82_U9453 ( .A1(u5_mult_82_n6775), .A2(u5_mult_82_n6543), 
        .ZN(u5_mult_82_ab_9__49_) );
  NOR2_X1 u5_mult_82_U9452 ( .A1(u5_mult_82_n6863), .A2(u5_mult_82_net65405), 
        .ZN(u5_mult_82_ab_40__29_) );
  NAND2_X1 u5_mult_82_U9451 ( .A1(u5_mult_82_ab_10__49_), .A2(
        u5_mult_82_CARRYB_9__49_), .ZN(u5_mult_82_n4338) );
  NAND2_X2 u5_mult_82_U9450 ( .A1(u5_mult_82_ab_10__49_), .A2(
        u5_mult_82_SUMB_9__50_), .ZN(u5_mult_82_n4337) );
  NAND2_X1 u5_mult_82_U9449 ( .A1(u5_mult_82_CARRYB_9__49_), .A2(
        u5_mult_82_SUMB_9__50_), .ZN(u5_mult_82_n4336) );
  XOR2_X2 u5_mult_82_U9448 ( .A(u5_mult_82_n1539), .B(u5_mult_82_n4335), .Z(
        u5_mult_82_SUMB_10__49_) );
  XOR2_X2 u5_mult_82_U9447 ( .A(u5_mult_82_CARRYB_9__49_), .B(
        u5_mult_82_ab_10__49_), .Z(u5_mult_82_n4335) );
  NAND3_X2 u5_mult_82_U9446 ( .A1(u5_mult_82_n4332), .A2(u5_mult_82_n4333), 
        .A3(u5_mult_82_n4334), .ZN(u5_mult_82_CARRYB_9__49_) );
  NAND2_X1 u5_mult_82_U9445 ( .A1(u5_mult_82_ab_9__49_), .A2(
        u5_mult_82_SUMB_8__50_), .ZN(u5_mult_82_n4334) );
  NAND2_X2 u5_mult_82_U9444 ( .A1(u5_mult_82_ab_9__49_), .A2(
        u5_mult_82_CARRYB_8__49_), .ZN(u5_mult_82_n4333) );
  NAND2_X1 u5_mult_82_U9443 ( .A1(u5_mult_82_SUMB_8__50_), .A2(
        u5_mult_82_CARRYB_8__49_), .ZN(u5_mult_82_n4332) );
  NAND2_X2 u5_mult_82_U9442 ( .A1(u5_mult_82_ab_40__29_), .A2(
        u5_mult_82_SUMB_39__30_), .ZN(u5_mult_82_n4330) );
  NAND3_X2 u5_mult_82_U9441 ( .A1(u5_mult_82_n4326), .A2(u5_mult_82_n4327), 
        .A3(u5_mult_82_n4328), .ZN(u5_mult_82_CARRYB_15__48_) );
  NAND3_X2 u5_mult_82_U9440 ( .A1(u5_mult_82_n4323), .A2(u5_mult_82_n4324), 
        .A3(u5_mult_82_n4325), .ZN(u5_mult_82_CARRYB_14__49_) );
  NAND2_X1 u5_mult_82_U9439 ( .A1(u5_mult_82_CARRYB_13__49_), .A2(
        u5_mult_82_SUMB_13__50_), .ZN(u5_mult_82_n4325) );
  NAND2_X2 u5_mult_82_U9438 ( .A1(u5_mult_82_ab_14__49_), .A2(
        u5_mult_82_SUMB_13__50_), .ZN(u5_mult_82_n4324) );
  NAND3_X4 u5_mult_82_U9437 ( .A1(u5_mult_82_n4319), .A2(u5_mult_82_n4320), 
        .A3(u5_mult_82_n4321), .ZN(u5_mult_82_CARRYB_31__36_) );
  NAND3_X2 u5_mult_82_U9436 ( .A1(u5_mult_82_n4316), .A2(u5_mult_82_n4317), 
        .A3(u5_mult_82_n4318), .ZN(u5_mult_82_CARRYB_30__37_) );
  NAND2_X2 u5_mult_82_U9435 ( .A1(u5_mult_82_CARRYB_29__37_), .A2(
        u5_mult_82_SUMB_29__38_), .ZN(u5_mult_82_n4318) );
  NAND2_X2 u5_mult_82_U9434 ( .A1(u5_mult_82_ab_30__37_), .A2(
        u5_mult_82_SUMB_29__38_), .ZN(u5_mult_82_n4317) );
  NAND2_X1 u5_mult_82_U9433 ( .A1(u5_mult_82_ab_30__37_), .A2(
        u5_mult_82_CARRYB_29__37_), .ZN(u5_mult_82_n4316) );
  XOR2_X2 u5_mult_82_U9432 ( .A(u5_mult_82_n4315), .B(u5_mult_82_SUMB_30__37_), 
        .Z(u5_mult_82_SUMB_31__36_) );
  XOR2_X2 u5_mult_82_U9431 ( .A(u5_mult_82_ab_31__36_), .B(
        u5_mult_82_CARRYB_30__36_), .Z(u5_mult_82_n4315) );
  NAND2_X1 u5_mult_82_U9430 ( .A1(u5_mult_82_CARRYB_51__21_), .A2(
        u5_mult_82_SUMB_51__22_), .ZN(u5_mult_82_n4314) );
  NAND2_X1 u5_mult_82_U9429 ( .A1(u5_mult_82_ab_52__21_), .A2(
        u5_mult_82_SUMB_51__22_), .ZN(u5_mult_82_n4313) );
  NAND2_X1 u5_mult_82_U9428 ( .A1(u5_mult_82_ab_52__21_), .A2(
        u5_mult_82_CARRYB_51__21_), .ZN(u5_mult_82_n4312) );
  NAND3_X2 u5_mult_82_U9427 ( .A1(u5_mult_82_n4309), .A2(u5_mult_82_n4310), 
        .A3(u5_mult_82_n4311), .ZN(u5_mult_82_CARRYB_51__22_) );
  NAND2_X2 u5_mult_82_U9426 ( .A1(u5_mult_82_CARRYB_50__22_), .A2(
        u5_mult_82_SUMB_50__23_), .ZN(u5_mult_82_n4311) );
  NAND2_X2 u5_mult_82_U9425 ( .A1(u5_mult_82_ab_51__22_), .A2(
        u5_mult_82_SUMB_50__23_), .ZN(u5_mult_82_n4310) );
  NAND2_X1 u5_mult_82_U9424 ( .A1(u5_mult_82_ab_51__22_), .A2(
        u5_mult_82_CARRYB_50__22_), .ZN(u5_mult_82_n4309) );
  XOR2_X2 u5_mult_82_U9423 ( .A(u5_mult_82_n4308), .B(u5_mult_82_SUMB_51__22_), 
        .Z(u5_mult_82_SUMB_52__21_) );
  XOR2_X2 u5_mult_82_U9422 ( .A(u5_mult_82_n4307), .B(u5_mult_82_n1434), .Z(
        u5_mult_82_SUMB_51__22_) );
  XOR2_X2 u5_mult_82_U9421 ( .A(u5_mult_82_ab_51__22_), .B(
        u5_mult_82_CARRYB_50__22_), .Z(u5_mult_82_n4307) );
  NAND3_X2 u5_mult_82_U9420 ( .A1(u5_mult_82_n4304), .A2(u5_mult_82_n4305), 
        .A3(u5_mult_82_n4306), .ZN(u5_mult_82_CARRYB_49__23_) );
  NAND2_X2 u5_mult_82_U9419 ( .A1(u5_mult_82_CARRYB_48__23_), .A2(
        u5_mult_82_SUMB_48__24_), .ZN(u5_mult_82_n4306) );
  NAND2_X2 u5_mult_82_U9418 ( .A1(u5_mult_82_ab_49__23_), .A2(
        u5_mult_82_SUMB_48__24_), .ZN(u5_mult_82_n4305) );
  NAND2_X1 u5_mult_82_U9417 ( .A1(u5_mult_82_ab_49__23_), .A2(
        u5_mult_82_CARRYB_48__23_), .ZN(u5_mult_82_n4304) );
  NAND3_X4 u5_mult_82_U9416 ( .A1(u5_mult_82_n4301), .A2(u5_mult_82_n4302), 
        .A3(u5_mult_82_n4303), .ZN(u5_mult_82_CARRYB_48__24_) );
  NAND2_X2 u5_mult_82_U9415 ( .A1(u5_mult_82_CARRYB_47__24_), .A2(
        u5_mult_82_SUMB_47__25_), .ZN(u5_mult_82_n4303) );
  NAND2_X2 u5_mult_82_U9414 ( .A1(u5_mult_82_ab_48__24_), .A2(
        u5_mult_82_SUMB_47__25_), .ZN(u5_mult_82_n4302) );
  NAND2_X2 u5_mult_82_U9413 ( .A1(u5_mult_82_ab_38__12_), .A2(
        u5_mult_82_SUMB_37__13_), .ZN(u5_mult_82_n5129) );
  NOR2_X1 u5_mult_82_U9412 ( .A1(u5_mult_82_n6927), .A2(u5_mult_82_net65353), 
        .ZN(u5_mult_82_ab_43__17_) );
  NAND3_X2 u5_mult_82_U9411 ( .A1(u5_mult_82_n4297), .A2(u5_mult_82_n4298), 
        .A3(u5_mult_82_n4299), .ZN(u5_mult_82_CARRYB_23__28_) );
  NAND2_X1 u5_mult_82_U9410 ( .A1(u5_mult_82_ab_22__29_), .A2(
        u5_mult_82_CARRYB_21__29_), .ZN(u5_mult_82_n4294) );
  XOR2_X2 u5_mult_82_U9409 ( .A(u5_mult_82_n4293), .B(u5_mult_82_SUMB_22__29_), 
        .Z(u5_mult_82_SUMB_23__28_) );
  NAND2_X1 u5_mult_82_U9408 ( .A1(u5_mult_82_CARRYB_44__15_), .A2(
        u5_mult_82_SUMB_44__16_), .ZN(u5_mult_82_n4291) );
  NAND2_X1 u5_mult_82_U9407 ( .A1(u5_mult_82_ab_45__15_), .A2(
        u5_mult_82_SUMB_44__16_), .ZN(u5_mult_82_n4290) );
  NAND2_X1 u5_mult_82_U9406 ( .A1(u5_mult_82_ab_45__15_), .A2(
        u5_mult_82_CARRYB_44__15_), .ZN(u5_mult_82_n4289) );
  NAND2_X2 u5_mult_82_U9405 ( .A1(u5_mult_82_CARRYB_43__16_), .A2(
        u5_mult_82_SUMB_43__17_), .ZN(u5_mult_82_n4288) );
  NAND2_X2 u5_mult_82_U9404 ( .A1(u5_mult_82_ab_44__16_), .A2(
        u5_mult_82_SUMB_43__17_), .ZN(u5_mult_82_n4287) );
  XOR2_X2 u5_mult_82_U9403 ( .A(u5_mult_82_n4285), .B(u5_mult_82_SUMB_43__17_), 
        .Z(u5_mult_82_SUMB_44__16_) );
  XOR2_X2 u5_mult_82_U9402 ( .A(u5_mult_82_ab_44__16_), .B(
        u5_mult_82_CARRYB_43__16_), .Z(u5_mult_82_n4285) );
  NAND3_X2 u5_mult_82_U9401 ( .A1(u5_mult_82_n4282), .A2(u5_mult_82_n4283), 
        .A3(u5_mult_82_n4284), .ZN(u5_mult_82_CARRYB_43__17_) );
  NAND2_X1 u5_mult_82_U9400 ( .A1(u5_mult_82_ab_43__17_), .A2(
        u5_mult_82_CARRYB_42__17_), .ZN(u5_mult_82_n4284) );
  XOR2_X2 u5_mult_82_U9399 ( .A(u5_mult_82_CARRYB_42__17_), .B(
        u5_mult_82_ab_43__17_), .Z(u5_mult_82_n4281) );
  XNOR2_X2 u5_mult_82_U9398 ( .A(u5_mult_82_CARRYB_20__16_), .B(
        u5_mult_82_ab_21__16_), .ZN(u5_mult_82_n4280) );
  XNOR2_X2 u5_mult_82_U9397 ( .A(u5_mult_82_SUMB_20__17_), .B(u5_mult_82_n4280), .ZN(u5_mult_82_SUMB_21__16_) );
  XNOR2_X2 u5_mult_82_U9396 ( .A(u5_mult_82_ab_48__7_), .B(
        u5_mult_82_CARRYB_47__7_), .ZN(u5_mult_82_net81962) );
  NOR2_X2 u5_mult_82_U9395 ( .A1(u5_mult_82_n6986), .A2(u5_mult_82_net65285), 
        .ZN(u5_mult_82_ab_47__0_) );
  NOR2_X1 u5_mult_82_U9394 ( .A1(u5_mult_82_n6852), .A2(u5_mult_82_n6521), 
        .ZN(u5_mult_82_ab_4__31_) );
  NAND3_X2 u5_mult_82_U9393 ( .A1(u5_mult_82_n4276), .A2(u5_mult_82_n4277), 
        .A3(u5_mult_82_n4278), .ZN(u5_mult_82_CARRYB_47__0_) );
  NAND2_X1 u5_mult_82_U9392 ( .A1(u5_mult_82_ab_47__0_), .A2(
        u5_mult_82_SUMB_46__1_), .ZN(u5_mult_82_n4277) );
  NAND3_X2 u5_mult_82_U9391 ( .A1(u5_mult_82_n4273), .A2(u5_mult_82_n4274), 
        .A3(u5_mult_82_n4275), .ZN(u5_mult_82_CARRYB_6__29_) );
  NAND2_X1 u5_mult_82_U9390 ( .A1(u5_mult_82_CARRYB_5__29_), .A2(
        u5_mult_82_SUMB_5__30_), .ZN(u5_mult_82_n4275) );
  NAND2_X1 u5_mult_82_U9389 ( .A1(u5_mult_82_ab_6__29_), .A2(
        u5_mult_82_SUMB_5__30_), .ZN(u5_mult_82_n4274) );
  NAND3_X2 u5_mult_82_U9388 ( .A1(u5_mult_82_n4270), .A2(u5_mult_82_n4271), 
        .A3(u5_mult_82_n4272), .ZN(u5_mult_82_CARRYB_5__30_) );
  NAND2_X2 u5_mult_82_U9387 ( .A1(u5_mult_82_CARRYB_4__30_), .A2(
        u5_mult_82_SUMB_4__31_), .ZN(u5_mult_82_n4272) );
  NAND2_X2 u5_mult_82_U9386 ( .A1(u5_mult_82_ab_5__30_), .A2(
        u5_mult_82_SUMB_4__31_), .ZN(u5_mult_82_n4271) );
  NAND2_X1 u5_mult_82_U9385 ( .A1(u5_mult_82_ab_5__30_), .A2(
        u5_mult_82_CARRYB_4__30_), .ZN(u5_mult_82_n4270) );
  XOR2_X2 u5_mult_82_U9384 ( .A(u5_mult_82_n4269), .B(u5_mult_82_SUMB_5__30_), 
        .Z(u5_mult_82_SUMB_6__29_) );
  XOR2_X2 u5_mult_82_U9383 ( .A(u5_mult_82_ab_6__29_), .B(
        u5_mult_82_CARRYB_5__29_), .Z(u5_mult_82_n4269) );
  XOR2_X2 u5_mult_82_U9382 ( .A(u5_mult_82_n4268), .B(u5_mult_82_SUMB_4__31_), 
        .Z(u5_mult_82_SUMB_5__30_) );
  XOR2_X2 u5_mult_82_U9381 ( .A(u5_mult_82_ab_5__30_), .B(
        u5_mult_82_CARRYB_4__30_), .Z(u5_mult_82_n4268) );
  NAND3_X2 u5_mult_82_U9380 ( .A1(u5_mult_82_n4265), .A2(u5_mult_82_n4266), 
        .A3(u5_mult_82_n4267), .ZN(u5_mult_82_CARRYB_4__31_) );
  NAND2_X1 u5_mult_82_U9379 ( .A1(u5_mult_82_ab_4__31_), .A2(
        u5_mult_82_CARRYB_3__31_), .ZN(u5_mult_82_n4267) );
  NAND2_X1 u5_mult_82_U9378 ( .A1(u5_mult_82_CARRYB_3__31_), .A2(
        u5_mult_82_SUMB_3__32_), .ZN(u5_mult_82_n4265) );
  XOR2_X2 u5_mult_82_U9377 ( .A(u5_mult_82_SUMB_3__32_), .B(u5_mult_82_n4264), 
        .Z(u5_mult_82_SUMB_4__31_) );
  XOR2_X2 u5_mult_82_U9376 ( .A(u5_mult_82_CARRYB_3__31_), .B(
        u5_mult_82_ab_4__31_), .Z(u5_mult_82_n4264) );
  NAND3_X2 u5_mult_82_U9375 ( .A1(u5_mult_82_n4261), .A2(u5_mult_82_n4262), 
        .A3(u5_mult_82_n4263), .ZN(u5_mult_82_CARRYB_11__24_) );
  NAND2_X1 u5_mult_82_U9374 ( .A1(u5_mult_82_CARRYB_10__24_), .A2(
        u5_mult_82_SUMB_10__25_), .ZN(u5_mult_82_n4263) );
  NAND2_X1 u5_mult_82_U9373 ( .A1(u5_mult_82_ab_11__24_), .A2(
        u5_mult_82_SUMB_10__25_), .ZN(u5_mult_82_n4262) );
  NAND2_X1 u5_mult_82_U9372 ( .A1(u5_mult_82_ab_11__24_), .A2(
        u5_mult_82_CARRYB_10__24_), .ZN(u5_mult_82_n4261) );
  NAND3_X2 u5_mult_82_U9371 ( .A1(u5_mult_82_n4258), .A2(u5_mult_82_n4259), 
        .A3(u5_mult_82_n4260), .ZN(u5_mult_82_CARRYB_10__25_) );
  NAND2_X2 u5_mult_82_U9370 ( .A1(u5_mult_82_CARRYB_9__25_), .A2(
        u5_mult_82_SUMB_9__26_), .ZN(u5_mult_82_n4260) );
  NAND2_X2 u5_mult_82_U9369 ( .A1(u5_mult_82_ab_10__25_), .A2(
        u5_mult_82_SUMB_9__26_), .ZN(u5_mult_82_n4259) );
  NAND2_X1 u5_mult_82_U9368 ( .A1(u5_mult_82_ab_10__25_), .A2(
        u5_mult_82_CARRYB_9__25_), .ZN(u5_mult_82_n4258) );
  XOR2_X2 u5_mult_82_U9367 ( .A(u5_mult_82_n4257), .B(u5_mult_82_SUMB_10__25_), 
        .Z(u5_mult_82_SUMB_11__24_) );
  NAND3_X2 u5_mult_82_U9366 ( .A1(u5_mult_82_n4254), .A2(u5_mult_82_n4255), 
        .A3(u5_mult_82_n4256), .ZN(u5_mult_82_CARRYB_9__26_) );
  NAND2_X1 u5_mult_82_U9365 ( .A1(u5_mult_82_CARRYB_8__26_), .A2(
        u5_mult_82_SUMB_8__27_), .ZN(u5_mult_82_n4256) );
  NAND2_X1 u5_mult_82_U9364 ( .A1(u5_mult_82_ab_9__26_), .A2(
        u5_mult_82_SUMB_8__27_), .ZN(u5_mult_82_n4255) );
  NAND2_X1 u5_mult_82_U9363 ( .A1(u5_mult_82_ab_9__26_), .A2(
        u5_mult_82_CARRYB_8__26_), .ZN(u5_mult_82_n4254) );
  NAND3_X2 u5_mult_82_U9362 ( .A1(u5_mult_82_n4251), .A2(u5_mult_82_n4252), 
        .A3(u5_mult_82_n4253), .ZN(u5_mult_82_CARRYB_8__27_) );
  NAND2_X1 u5_mult_82_U9361 ( .A1(u5_mult_82_CARRYB_7__27_), .A2(
        u5_mult_82_SUMB_7__28_), .ZN(u5_mult_82_n4253) );
  NAND2_X1 u5_mult_82_U9360 ( .A1(u5_mult_82_ab_8__27_), .A2(
        u5_mult_82_SUMB_7__28_), .ZN(u5_mult_82_n4252) );
  NAND2_X1 u5_mult_82_U9359 ( .A1(u5_mult_82_ab_8__27_), .A2(
        u5_mult_82_CARRYB_7__27_), .ZN(u5_mult_82_n4251) );
  XOR2_X2 u5_mult_82_U9358 ( .A(u5_mult_82_n4250), .B(u5_mult_82_SUMB_8__27_), 
        .Z(u5_mult_82_SUMB_9__26_) );
  XOR2_X2 u5_mult_82_U9357 ( .A(u5_mult_82_ab_9__26_), .B(
        u5_mult_82_CARRYB_8__26_), .Z(u5_mult_82_n4250) );
  XOR2_X2 u5_mult_82_U9356 ( .A(u5_mult_82_n4249), .B(u5_mult_82_SUMB_7__28_), 
        .Z(u5_mult_82_SUMB_8__27_) );
  XOR2_X2 u5_mult_82_U9355 ( .A(u5_mult_82_ab_8__27_), .B(
        u5_mult_82_CARRYB_7__27_), .Z(u5_mult_82_n4249) );
  NAND3_X4 u5_mult_82_U9354 ( .A1(u5_mult_82_n5658), .A2(u5_mult_82_n5659), 
        .A3(u5_mult_82_n5660), .ZN(u5_mult_82_CARRYB_47__18_) );
  XNOR2_X2 u5_mult_82_U9353 ( .A(u5_mult_82_ab_41__17_), .B(
        u5_mult_82_CARRYB_40__17_), .ZN(u5_mult_82_n4248) );
  XNOR2_X2 u5_mult_82_U9352 ( .A(u5_mult_82_n4248), .B(u5_mult_82_SUMB_40__18_), .ZN(u5_mult_82_SUMB_41__17_) );
  NAND2_X1 u5_mult_82_U9351 ( .A1(u5_mult_82_ab_35__21_), .A2(
        u5_mult_82_CARRYB_34__21_), .ZN(u5_mult_82_n4245) );
  NAND2_X2 u5_mult_82_U9350 ( .A1(u5_mult_82_CARRYB_33__22_), .A2(
        u5_mult_82_SUMB_33__23_), .ZN(u5_mult_82_n4244) );
  NAND2_X2 u5_mult_82_U9349 ( .A1(u5_mult_82_ab_34__22_), .A2(
        u5_mult_82_SUMB_33__23_), .ZN(u5_mult_82_n4243) );
  NAND2_X1 u5_mult_82_U9348 ( .A1(u5_mult_82_ab_34__22_), .A2(
        u5_mult_82_CARRYB_33__22_), .ZN(u5_mult_82_n4242) );
  NAND3_X2 u5_mult_82_U9347 ( .A1(u5_mult_82_n4239), .A2(u5_mult_82_n4240), 
        .A3(u5_mult_82_n4241), .ZN(u5_mult_82_CARRYB_32__24_) );
  NAND2_X1 u5_mult_82_U9346 ( .A1(u5_mult_82_ab_32__24_), .A2(
        u5_mult_82_CARRYB_31__24_), .ZN(u5_mult_82_n4239) );
  NAND3_X2 u5_mult_82_U9345 ( .A1(u5_mult_82_n4236), .A2(u5_mult_82_n4237), 
        .A3(u5_mult_82_n4238), .ZN(u5_mult_82_CARRYB_31__25_) );
  NAND2_X2 u5_mult_82_U9344 ( .A1(u5_mult_82_ab_31__25_), .A2(
        u5_mult_82_SUMB_30__26_), .ZN(u5_mult_82_n4237) );
  XOR2_X2 u5_mult_82_U9343 ( .A(u5_mult_82_n4235), .B(u5_mult_82_SUMB_30__26_), 
        .Z(u5_mult_82_SUMB_31__25_) );
  NAND3_X2 u5_mult_82_U9342 ( .A1(u5_mult_82_n4232), .A2(u5_mult_82_n4233), 
        .A3(u5_mult_82_n4234), .ZN(u5_mult_82_CARRYB_43__18_) );
  NAND3_X4 u5_mult_82_U9341 ( .A1(u5_mult_82_n4229), .A2(u5_mult_82_n4230), 
        .A3(u5_mult_82_n4231), .ZN(u5_mult_82_CARRYB_42__19_) );
  NAND2_X2 u5_mult_82_U9340 ( .A1(u5_mult_82_CARRYB_41__19_), .A2(
        u5_mult_82_n25), .ZN(u5_mult_82_n4231) );
  NAND2_X2 u5_mult_82_U9339 ( .A1(u5_mult_82_ab_42__19_), .A2(u5_mult_82_n25), 
        .ZN(u5_mult_82_n4230) );
  NAND2_X1 u5_mult_82_U9338 ( .A1(u5_mult_82_ab_42__19_), .A2(
        u5_mult_82_CARRYB_41__19_), .ZN(u5_mult_82_n4229) );
  XOR2_X2 u5_mult_82_U9337 ( .A(u5_mult_82_ab_42__19_), .B(
        u5_mult_82_CARRYB_41__19_), .Z(u5_mult_82_n4228) );
  NAND2_X2 u5_mult_82_U9336 ( .A1(u5_mult_82_n4226), .A2(u5_mult_82_n4227), 
        .ZN(u5_mult_82_n5852) );
  NAND2_X2 u5_mult_82_U9335 ( .A1(u5_mult_82_ab_48__15_), .A2(u5_mult_82_n1418), .ZN(u5_mult_82_n4227) );
  NAND2_X1 u5_mult_82_U9334 ( .A1(u5_mult_82_n5521), .A2(
        u5_mult_82_SUMB_47__16_), .ZN(u5_mult_82_n4226) );
  NAND2_X1 u5_mult_82_U9333 ( .A1(u5_mult_82_ab_32__38_), .A2(
        u5_mult_82_CARRYB_31__38_), .ZN(u5_mult_82_n4927) );
  NAND2_X2 u5_mult_82_U9332 ( .A1(u5_mult_82_SUMB_47__2_), .A2(
        u5_mult_82_CARRYB_47__1_), .ZN(u5_mult_82_n5816) );
  NOR2_X1 u5_mult_82_U9331 ( .A1(u5_mult_82_n6933), .A2(u5_mult_82_net65229), 
        .ZN(u5_mult_82_ab_50__15_) );
  NAND3_X2 u5_mult_82_U9330 ( .A1(u5_mult_82_n4223), .A2(u5_mult_82_n4224), 
        .A3(u5_mult_82_n4225), .ZN(u5_mult_82_CARRYB_50__15_) );
  NAND2_X1 u5_mult_82_U9329 ( .A1(u5_mult_82_ab_50__15_), .A2(
        u5_mult_82_CARRYB_49__15_), .ZN(u5_mult_82_n4225) );
  NAND2_X2 u5_mult_82_U9328 ( .A1(u5_mult_82_ab_50__15_), .A2(
        u5_mult_82_SUMB_49__16_), .ZN(u5_mult_82_n4224) );
  NAND2_X1 u5_mult_82_U9327 ( .A1(u5_mult_82_CARRYB_49__15_), .A2(
        u5_mult_82_SUMB_49__16_), .ZN(u5_mult_82_n4223) );
  XNOR2_X2 u5_mult_82_U9326 ( .A(u5_mult_82_n5222), .B(
        u5_mult_82_CARRYB_47__10_), .ZN(u5_mult_82_n6205) );
  NAND2_X2 u5_mult_82_U9325 ( .A1(u5_mult_82_CARRYB_42__7_), .A2(
        u5_mult_82_SUMB_42__8_), .ZN(u5_mult_82_n6073) );
  NAND2_X1 u5_mult_82_U9324 ( .A1(u5_mult_82_CARRYB_37__12_), .A2(
        u5_mult_82_SUMB_37__13_), .ZN(u5_mult_82_n5130) );
  NAND2_X2 u5_mult_82_U9323 ( .A1(u5_mult_82_ab_38__13_), .A2(
        u5_mult_82_CARRYB_37__13_), .ZN(u5_mult_82_n4625) );
  NOR2_X2 u5_mult_82_U9322 ( .A1(u5_mult_82_net64505), .A2(u5_mult_82_n6722), 
        .ZN(u5_mult_82_ab_37__13_) );
  NAND3_X2 u5_mult_82_U9321 ( .A1(u5_mult_82_n5491), .A2(u5_mult_82_n5492), 
        .A3(u5_mult_82_n5493), .ZN(u5_mult_82_CARRYB_44__8_) );
  NOR2_X1 u5_mult_82_U9320 ( .A1(u5_mult_82_net64415), .A2(u5_mult_82_net65319), .ZN(u5_mult_82_ab_45__8_) );
  NOR2_X1 u5_mult_82_U9319 ( .A1(u5_mult_82_n6913), .A2(u5_mult_82_n6664), 
        .ZN(u5_mult_82_ab_28__19_) );
  NAND3_X2 u5_mult_82_U9318 ( .A1(u5_mult_82_n4221), .A2(u5_mult_82_n4220), 
        .A3(u5_mult_82_n4219), .ZN(u5_mult_82_CARRYB_45__8_) );
  NAND2_X1 u5_mult_82_U9317 ( .A1(u5_mult_82_ab_45__8_), .A2(
        u5_mult_82_SUMB_44__9_), .ZN(u5_mult_82_n4221) );
  NAND2_X2 u5_mult_82_U9316 ( .A1(u5_mult_82_ab_45__8_), .A2(
        u5_mult_82_CARRYB_44__8_), .ZN(u5_mult_82_n4220) );
  NAND2_X1 u5_mult_82_U9315 ( .A1(u5_mult_82_ab_28__19_), .A2(
        u5_mult_82_CARRYB_27__19_), .ZN(u5_mult_82_n4217) );
  XOR2_X2 u5_mult_82_U9314 ( .A(u5_mult_82_CARRYB_27__19_), .B(
        u5_mult_82_ab_28__19_), .Z(u5_mult_82_net82046) );
  INV_X4 u5_mult_82_U9313 ( .A(u5_mult_82_net80255), .ZN(u5_mult_82_net82039)
         );
  NAND2_X1 u5_mult_82_U9312 ( .A1(u5_mult_82_SUMB_14__30_), .A2(
        u5_mult_82_net82039), .ZN(u5_mult_82_net82040) );
  NAND2_X2 u5_mult_82_U9311 ( .A1(u5_mult_82_ab_48__1_), .A2(
        u5_mult_82_SUMB_47__2_), .ZN(u5_mult_82_n5814) );
  NAND2_X2 u5_mult_82_U9310 ( .A1(u5_mult_82_ab_47__11_), .A2(
        u5_mult_82_SUMB_46__12_), .ZN(u5_mult_82_n6207) );
  NAND2_X1 u5_mult_82_U9309 ( .A1(u5_mult_82_CARRYB_38__19_), .A2(
        u5_mult_82_SUMB_38__20_), .ZN(u5_mult_82_n4216) );
  NAND2_X1 u5_mult_82_U9308 ( .A1(u5_mult_82_ab_39__19_), .A2(
        u5_mult_82_SUMB_38__20_), .ZN(u5_mult_82_n4215) );
  NAND2_X1 u5_mult_82_U9307 ( .A1(u5_mult_82_ab_39__19_), .A2(
        u5_mult_82_CARRYB_38__19_), .ZN(u5_mult_82_n4214) );
  NAND2_X2 u5_mult_82_U9306 ( .A1(u5_mult_82_CARRYB_37__20_), .A2(
        u5_mult_82_SUMB_37__21_), .ZN(u5_mult_82_n4213) );
  NAND2_X2 u5_mult_82_U9305 ( .A1(u5_mult_82_ab_38__20_), .A2(
        u5_mult_82_SUMB_37__21_), .ZN(u5_mult_82_n4212) );
  NAND2_X1 u5_mult_82_U9304 ( .A1(u5_mult_82_ab_38__20_), .A2(
        u5_mult_82_CARRYB_37__20_), .ZN(u5_mult_82_n4211) );
  NAND2_X2 u5_mult_82_U9303 ( .A1(u5_mult_82_CARRYB_45__13_), .A2(
        u5_mult_82_SUMB_45__14_), .ZN(u5_mult_82_n4210) );
  NAND2_X2 u5_mult_82_U9302 ( .A1(u5_mult_82_ab_46__13_), .A2(
        u5_mult_82_SUMB_45__14_), .ZN(u5_mult_82_n4209) );
  NAND2_X1 u5_mult_82_U9301 ( .A1(u5_mult_82_ab_46__13_), .A2(
        u5_mult_82_CARRYB_45__13_), .ZN(u5_mult_82_n4208) );
  NAND3_X2 u5_mult_82_U9300 ( .A1(u5_mult_82_n4207), .A2(u5_mult_82_n4206), 
        .A3(u5_mult_82_n4205), .ZN(u5_mult_82_CARRYB_45__14_) );
  NAND2_X2 u5_mult_82_U9299 ( .A1(u5_mult_82_ab_45__14_), .A2(
        u5_mult_82_CARRYB_44__14_), .ZN(u5_mult_82_n4205) );
  XNOR2_X2 u5_mult_82_U9298 ( .A(u5_mult_82_n4204), .B(u5_mult_82_SUMB_42__19_), .ZN(u5_mult_82_SUMB_43__18_) );
  NOR2_X1 u5_mult_82_U9297 ( .A1(u5_mult_82_n6867), .A2(u5_mult_82_n6747), 
        .ZN(u5_mult_82_ab_48__28_) );
  NOR2_X1 u5_mult_82_U9296 ( .A1(u5_mult_82_net64937), .A2(u5_mult_82_n6727), 
        .ZN(u5_mult_82_ab_39__37_) );
  NAND3_X2 u5_mult_82_U9295 ( .A1(u5_mult_82_n4201), .A2(u5_mult_82_n4202), 
        .A3(u5_mult_82_n4203), .ZN(u5_mult_82_CARRYB_35__41_) );
  NAND2_X1 u5_mult_82_U9294 ( .A1(u5_mult_82_CARRYB_34__41_), .A2(
        u5_mult_82_SUMB_34__42_), .ZN(u5_mult_82_n4203) );
  NAND2_X2 u5_mult_82_U9293 ( .A1(u5_mult_82_ab_35__41_), .A2(
        u5_mult_82_SUMB_34__42_), .ZN(u5_mult_82_n4202) );
  NAND2_X1 u5_mult_82_U9292 ( .A1(u5_mult_82_ab_35__41_), .A2(
        u5_mult_82_CARRYB_34__41_), .ZN(u5_mult_82_n4201) );
  NAND3_X2 u5_mult_82_U9291 ( .A1(u5_mult_82_n4198), .A2(u5_mult_82_n4199), 
        .A3(u5_mult_82_n4200), .ZN(u5_mult_82_CARRYB_34__42_) );
  NAND2_X2 u5_mult_82_U9290 ( .A1(u5_mult_82_CARRYB_33__42_), .A2(
        u5_mult_82_n1563), .ZN(u5_mult_82_n4200) );
  NAND2_X2 u5_mult_82_U9289 ( .A1(u5_mult_82_ab_34__42_), .A2(u5_mult_82_n1563), .ZN(u5_mult_82_n4199) );
  NAND2_X2 u5_mult_82_U9288 ( .A1(u5_mult_82_ab_34__42_), .A2(
        u5_mult_82_CARRYB_33__42_), .ZN(u5_mult_82_n4198) );
  XOR2_X2 u5_mult_82_U9287 ( .A(u5_mult_82_n4197), .B(u5_mult_82_n1563), .Z(
        u5_mult_82_SUMB_34__42_) );
  XOR2_X2 u5_mult_82_U9286 ( .A(u5_mult_82_ab_34__42_), .B(
        u5_mult_82_CARRYB_33__42_), .Z(u5_mult_82_n4197) );
  NAND3_X2 u5_mult_82_U9285 ( .A1(u5_mult_82_n4194), .A2(u5_mult_82_n4195), 
        .A3(u5_mult_82_n4196), .ZN(u5_mult_82_CARRYB_48__28_) );
  NAND2_X1 u5_mult_82_U9284 ( .A1(u5_mult_82_ab_48__28_), .A2(
        u5_mult_82_CARRYB_47__28_), .ZN(u5_mult_82_n4196) );
  NAND2_X1 u5_mult_82_U9283 ( .A1(u5_mult_82_ab_48__28_), .A2(
        u5_mult_82_SUMB_47__29_), .ZN(u5_mult_82_n4195) );
  NAND2_X1 u5_mult_82_U9282 ( .A1(u5_mult_82_CARRYB_47__28_), .A2(
        u5_mult_82_SUMB_47__29_), .ZN(u5_mult_82_n4194) );
  NAND3_X2 u5_mult_82_U9281 ( .A1(u5_mult_82_n4191), .A2(u5_mult_82_n4192), 
        .A3(u5_mult_82_n4193), .ZN(u5_mult_82_CARRYB_39__37_) );
  NAND2_X1 u5_mult_82_U9280 ( .A1(u5_mult_82_ab_39__37_), .A2(
        u5_mult_82_CARRYB_38__37_), .ZN(u5_mult_82_n4193) );
  NAND2_X1 u5_mult_82_U9279 ( .A1(u5_mult_82_ab_39__37_), .A2(
        u5_mult_82_SUMB_38__38_), .ZN(u5_mult_82_n4192) );
  NAND2_X1 u5_mult_82_U9278 ( .A1(u5_mult_82_CARRYB_38__37_), .A2(
        u5_mult_82_SUMB_38__38_), .ZN(u5_mult_82_n4191) );
  XOR2_X2 u5_mult_82_U9277 ( .A(u5_mult_82_SUMB_38__38_), .B(u5_mult_82_n4190), 
        .Z(u5_mult_82_SUMB_39__37_) );
  XOR2_X2 u5_mult_82_U9276 ( .A(u5_mult_82_CARRYB_38__37_), .B(
        u5_mult_82_ab_39__37_), .Z(u5_mult_82_n4190) );
  NAND3_X2 u5_mult_82_U9275 ( .A1(u5_mult_82_n4187), .A2(u5_mult_82_n4188), 
        .A3(u5_mult_82_n4189), .ZN(u5_mult_82_CARRYB_51__25_) );
  NAND2_X1 u5_mult_82_U9274 ( .A1(u5_mult_82_SUMB_50__26_), .A2(
        u5_mult_82_CARRYB_50__25_), .ZN(u5_mult_82_n4189) );
  NAND2_X1 u5_mult_82_U9273 ( .A1(u5_mult_82_ab_51__25_), .A2(
        u5_mult_82_CARRYB_50__25_), .ZN(u5_mult_82_n4187) );
  NAND3_X2 u5_mult_82_U9272 ( .A1(u5_mult_82_n4184), .A2(u5_mult_82_n4185), 
        .A3(u5_mult_82_n4186), .ZN(u5_mult_82_CARRYB_50__26_) );
  NAND2_X1 u5_mult_82_U9271 ( .A1(u5_mult_82_CARRYB_49__26_), .A2(
        u5_mult_82_SUMB_49__27_), .ZN(u5_mult_82_n4186) );
  NAND2_X1 u5_mult_82_U9270 ( .A1(u5_mult_82_ab_50__26_), .A2(
        u5_mult_82_SUMB_49__27_), .ZN(u5_mult_82_n4185) );
  XNOR2_X2 u5_mult_82_U9269 ( .A(u5_mult_82_n4182), .B(u5_mult_82_SUMB_49__9_), 
        .ZN(u5_mult_82_SUMB_50__8_) );
  NAND2_X2 u5_mult_82_U9268 ( .A1(u5_mult_82_ab_38__16_), .A2(
        u5_mult_82_SUMB_37__17_), .ZN(u5_mult_82_n5433) );
  NAND2_X2 u5_mult_82_U9267 ( .A1(u5_mult_82_ab_48__10_), .A2(
        u5_mult_82_CARRYB_47__10_), .ZN(u5_mult_82_n6209) );
  NOR2_X2 u5_mult_82_U9266 ( .A1(u5_mult_82_net64455), .A2(u5_mult_82_net65283), .ZN(u5_mult_82_ab_47__10_) );
  NAND3_X4 u5_mult_82_U9265 ( .A1(u5_mult_82_n4179), .A2(u5_mult_82_n4180), 
        .A3(u5_mult_82_n4181), .ZN(u5_mult_82_CARRYB_47__10_) );
  NAND2_X2 u5_mult_82_U9264 ( .A1(u5_mult_82_ab_47__10_), .A2(
        u5_mult_82_CARRYB_46__10_), .ZN(u5_mult_82_n4180) );
  NAND3_X2 u5_mult_82_U9263 ( .A1(u5_mult_82_n4176), .A2(u5_mult_82_n4177), 
        .A3(u5_mult_82_n4178), .ZN(u5_mult_82_CARRYB_4__38_) );
  NAND2_X1 u5_mult_82_U9262 ( .A1(u5_mult_82_CARRYB_3__38_), .A2(
        u5_mult_82_SUMB_3__39_), .ZN(u5_mult_82_n4178) );
  NAND2_X1 u5_mult_82_U9261 ( .A1(u5_mult_82_ab_4__38_), .A2(
        u5_mult_82_SUMB_3__39_), .ZN(u5_mult_82_n4177) );
  NAND2_X1 u5_mult_82_U9260 ( .A1(u5_mult_82_ab_4__38_), .A2(
        u5_mult_82_CARRYB_3__38_), .ZN(u5_mult_82_n4176) );
  NAND3_X2 u5_mult_82_U9259 ( .A1(u5_mult_82_n4173), .A2(u5_mult_82_n4174), 
        .A3(u5_mult_82_n4175), .ZN(u5_mult_82_CARRYB_3__39_) );
  NAND2_X1 u5_mult_82_U9258 ( .A1(u5_mult_82_ab_3__39_), .A2(
        u5_mult_82_CARRYB_2__39_), .ZN(u5_mult_82_n4173) );
  XOR2_X2 u5_mult_82_U9257 ( .A(u5_mult_82_n4172), .B(u5_mult_82_SUMB_2__40_), 
        .Z(u5_mult_82_SUMB_3__39_) );
  XOR2_X2 u5_mult_82_U9256 ( .A(u5_mult_82_ab_3__39_), .B(
        u5_mult_82_CARRYB_2__39_), .Z(u5_mult_82_n4172) );
  NAND2_X1 u5_mult_82_U9255 ( .A1(u5_mult_82_ab_51__8_), .A2(
        u5_mult_82_SUMB_50__9_), .ZN(u5_mult_82_n4170) );
  NAND2_X1 u5_mult_82_U9254 ( .A1(u5_mult_82_ab_51__8_), .A2(
        u5_mult_82_CARRYB_50__8_), .ZN(u5_mult_82_n4169) );
  NAND3_X2 u5_mult_82_U9253 ( .A1(u5_mult_82_n4166), .A2(u5_mult_82_n4167), 
        .A3(u5_mult_82_n4168), .ZN(u5_mult_82_CARRYB_50__9_) );
  NAND2_X1 u5_mult_82_U9252 ( .A1(u5_mult_82_CARRYB_49__9_), .A2(
        u5_mult_82_SUMB_49__10_), .ZN(u5_mult_82_n4168) );
  NAND2_X1 u5_mult_82_U9251 ( .A1(u5_mult_82_ab_50__9_), .A2(
        u5_mult_82_SUMB_49__10_), .ZN(u5_mult_82_n4167) );
  NAND2_X1 u5_mult_82_U9250 ( .A1(u5_mult_82_ab_50__9_), .A2(
        u5_mult_82_CARRYB_49__9_), .ZN(u5_mult_82_n4166) );
  XOR2_X2 u5_mult_82_U9249 ( .A(u5_mult_82_n4165), .B(u5_mult_82_SUMB_49__10_), 
        .Z(u5_mult_82_SUMB_50__9_) );
  XOR2_X2 u5_mult_82_U9248 ( .A(u5_mult_82_n6223), .B(u5_mult_82_SUMB_24__34_), 
        .Z(u5_mult_82_SUMB_25__33_) );
  NAND2_X2 u5_mult_82_U9247 ( .A1(u5_mult_82_CARRYB_46__18_), .A2(
        u5_mult_82_SUMB_46__19_), .ZN(u5_mult_82_n5658) );
  NAND2_X4 u5_mult_82_U9246 ( .A1(u5_mult_82_n4157), .A2(u5_mult_82_n1636), 
        .ZN(u5_mult_82_n4159) );
  NAND2_X4 u5_mult_82_U9245 ( .A1(u5_mult_82_n4686), .A2(u5_mult_82_n4687), 
        .ZN(u5_mult_82_n4689) );
  NOR2_X1 u5_mult_82_U9244 ( .A1(u5_mult_82_net64361), .A2(u5_mult_82_net65445), .ZN(u5_mult_82_ab_38__5_) );
  NAND3_X2 u5_mult_82_U9243 ( .A1(u5_mult_82_n4154), .A2(u5_mult_82_n4155), 
        .A3(u5_mult_82_n4156), .ZN(u5_mult_82_CARRYB_34__9_) );
  NAND2_X1 u5_mult_82_U9242 ( .A1(u5_mult_82_ab_34__9_), .A2(
        u5_mult_82_CARRYB_33__9_), .ZN(u5_mult_82_n4154) );
  NAND2_X2 u5_mult_82_U9241 ( .A1(u5_mult_82_SUMB_32__11_), .A2(
        u5_mult_82_n1514), .ZN(u5_mult_82_n4153) );
  NAND2_X2 u5_mult_82_U9240 ( .A1(u5_mult_82_ab_33__10_), .A2(
        u5_mult_82_SUMB_32__11_), .ZN(u5_mult_82_n4152) );
  NAND3_X2 u5_mult_82_U9239 ( .A1(u5_mult_82_n4148), .A2(u5_mult_82_n4149), 
        .A3(u5_mult_82_n4150), .ZN(u5_mult_82_CARRYB_38__5_) );
  NAND2_X2 u5_mult_82_U9238 ( .A1(u5_mult_82_ab_38__5_), .A2(
        u5_mult_82_SUMB_37__6_), .ZN(u5_mult_82_n4149) );
  NAND2_X1 u5_mult_82_U9237 ( .A1(u5_mult_82_CARRYB_37__5_), .A2(
        u5_mult_82_SUMB_37__6_), .ZN(u5_mult_82_n4148) );
  NAND2_X2 u5_mult_82_U9236 ( .A1(u5_mult_82_CARRYB_22__19_), .A2(
        u5_mult_82_SUMB_22__20_), .ZN(u5_mult_82_n4666) );
  XOR2_X2 u5_mult_82_U9235 ( .A(u5_mult_82_ab_11__24_), .B(
        u5_mult_82_CARRYB_10__24_), .Z(u5_mult_82_n4257) );
  XNOR2_X2 u5_mult_82_U9234 ( .A(u5_mult_82_n4146), .B(u5_mult_82_SUMB_46__7_), 
        .ZN(u5_mult_82_SUMB_47__6_) );
  XOR2_X2 u5_mult_82_U9233 ( .A(u5_mult_82_n4648), .B(u5_mult_82_ab_10__52_), 
        .Z(u5_mult_82_SUMB_11__51_) );
  XNOR2_X2 u5_mult_82_U9232 ( .A(u5_mult_82_CARRYB_22__17_), .B(
        u5_mult_82_ab_23__17_), .ZN(u5_mult_82_n4145) );
  XNOR2_X2 u5_mult_82_U9231 ( .A(u5_mult_82_SUMB_22__18_), .B(u5_mult_82_n4145), .ZN(u5_mult_82_SUMB_23__17_) );
  NAND2_X1 u5_mult_82_U9230 ( .A1(u5_mult_82_CARRYB_12__37_), .A2(
        u5_mult_82_SUMB_12__38_), .ZN(u5_mult_82_n6094) );
  XNOR2_X2 u5_mult_82_U9229 ( .A(u5_mult_82_ab_48__20_), .B(
        u5_mult_82_CARRYB_47__20_), .ZN(u5_mult_82_n4144) );
  XNOR2_X2 u5_mult_82_U9228 ( .A(u5_mult_82_n4144), .B(u5_mult_82_SUMB_47__21_), .ZN(u5_mult_82_SUMB_48__20_) );
  NOR2_X2 u5_mult_82_U9227 ( .A1(u5_mult_82_net64361), .A2(u5_mult_82_n6722), 
        .ZN(u5_mult_82_ab_37__5_) );
  NAND3_X2 u5_mult_82_U9226 ( .A1(u5_mult_82_n4141), .A2(u5_mult_82_n4142), 
        .A3(u5_mult_82_n4143), .ZN(u5_mult_82_CARRYB_3__31_) );
  NAND2_X1 u5_mult_82_U9225 ( .A1(u5_mult_82_CARRYB_2__31_), .A2(
        u5_mult_82_SUMB_2__32_), .ZN(u5_mult_82_n4143) );
  NAND2_X1 u5_mult_82_U9224 ( .A1(u5_mult_82_ab_3__31_), .A2(
        u5_mult_82_SUMB_2__32_), .ZN(u5_mult_82_n4142) );
  NAND2_X1 u5_mult_82_U9223 ( .A1(u5_mult_82_ab_3__31_), .A2(
        u5_mult_82_CARRYB_2__31_), .ZN(u5_mult_82_n4141) );
  NAND3_X2 u5_mult_82_U9222 ( .A1(u5_mult_82_n4138), .A2(u5_mult_82_n4139), 
        .A3(u5_mult_82_n4140), .ZN(u5_mult_82_CARRYB_2__32_) );
  NAND2_X2 u5_mult_82_U9221 ( .A1(u5_mult_82_CARRYB_1__32_), .A2(
        u5_mult_82_SUMB_1__33_), .ZN(u5_mult_82_n4140) );
  NAND2_X2 u5_mult_82_U9220 ( .A1(u5_mult_82_ab_2__32_), .A2(
        u5_mult_82_SUMB_1__33_), .ZN(u5_mult_82_n4139) );
  NAND2_X1 u5_mult_82_U9219 ( .A1(u5_mult_82_ab_2__32_), .A2(
        u5_mult_82_CARRYB_1__32_), .ZN(u5_mult_82_n4138) );
  XOR2_X2 u5_mult_82_U9218 ( .A(u5_mult_82_n4137), .B(u5_mult_82_SUMB_2__32_), 
        .Z(u5_mult_82_SUMB_3__31_) );
  XOR2_X2 u5_mult_82_U9217 ( .A(u5_mult_82_ab_3__31_), .B(
        u5_mult_82_CARRYB_2__31_), .Z(u5_mult_82_n4137) );
  XOR2_X2 u5_mult_82_U9216 ( .A(u5_mult_82_n4136), .B(u5_mult_82_SUMB_1__33_), 
        .Z(u5_mult_82_SUMB_2__32_) );
  XOR2_X2 u5_mult_82_U9215 ( .A(u5_mult_82_ab_2__32_), .B(
        u5_mult_82_CARRYB_1__32_), .Z(u5_mult_82_n4136) );
  NAND3_X2 u5_mult_82_U9214 ( .A1(u5_mult_82_n4133), .A2(u5_mult_82_n4134), 
        .A3(u5_mult_82_n4135), .ZN(u5_mult_82_CARRYB_14__20_) );
  NAND2_X1 u5_mult_82_U9213 ( .A1(u5_mult_82_CARRYB_13__20_), .A2(
        u5_mult_82_SUMB_13__21_), .ZN(u5_mult_82_n4135) );
  NAND2_X1 u5_mult_82_U9212 ( .A1(u5_mult_82_ab_14__20_), .A2(
        u5_mult_82_SUMB_13__21_), .ZN(u5_mult_82_n4134) );
  NAND2_X1 u5_mult_82_U9211 ( .A1(u5_mult_82_ab_14__20_), .A2(
        u5_mult_82_CARRYB_13__20_), .ZN(u5_mult_82_n4133) );
  NAND3_X2 u5_mult_82_U9210 ( .A1(u5_mult_82_n4130), .A2(u5_mult_82_n4131), 
        .A3(u5_mult_82_n4132), .ZN(u5_mult_82_CARRYB_13__21_) );
  NAND2_X2 u5_mult_82_U9209 ( .A1(u5_mult_82_CARRYB_12__21_), .A2(
        u5_mult_82_SUMB_12__22_), .ZN(u5_mult_82_n4132) );
  NAND2_X2 u5_mult_82_U9208 ( .A1(u5_mult_82_ab_13__21_), .A2(
        u5_mult_82_SUMB_12__22_), .ZN(u5_mult_82_n4131) );
  NAND2_X1 u5_mult_82_U9207 ( .A1(u5_mult_82_ab_13__21_), .A2(
        u5_mult_82_CARRYB_12__21_), .ZN(u5_mult_82_n4130) );
  XOR2_X2 u5_mult_82_U9206 ( .A(u5_mult_82_n4129), .B(u5_mult_82_SUMB_13__21_), 
        .Z(u5_mult_82_SUMB_14__20_) );
  XOR2_X2 u5_mult_82_U9205 ( .A(u5_mult_82_ab_14__20_), .B(
        u5_mult_82_CARRYB_13__20_), .Z(u5_mult_82_n4129) );
  XOR2_X2 u5_mult_82_U9204 ( .A(u5_mult_82_n4128), .B(u5_mult_82_SUMB_12__22_), 
        .Z(u5_mult_82_SUMB_13__21_) );
  XOR2_X2 u5_mult_82_U9203 ( .A(u5_mult_82_ab_13__21_), .B(
        u5_mult_82_CARRYB_12__21_), .Z(u5_mult_82_n4128) );
  NAND3_X4 u5_mult_82_U9202 ( .A1(u5_mult_82_n4125), .A2(u5_mult_82_n4126), 
        .A3(u5_mult_82_n4127), .ZN(u5_mult_82_CARRYB_7__27_) );
  NAND2_X1 u5_mult_82_U9201 ( .A1(u5_mult_82_CARRYB_6__27_), .A2(
        u5_mult_82_SUMB_6__28_), .ZN(u5_mult_82_n4127) );
  NAND2_X1 u5_mult_82_U9200 ( .A1(u5_mult_82_ab_7__27_), .A2(
        u5_mult_82_SUMB_6__28_), .ZN(u5_mult_82_n4126) );
  NAND2_X1 u5_mult_82_U9199 ( .A1(u5_mult_82_ab_7__27_), .A2(
        u5_mult_82_CARRYB_6__27_), .ZN(u5_mult_82_n4125) );
  NAND3_X2 u5_mult_82_U9198 ( .A1(u5_mult_82_n4122), .A2(u5_mult_82_n4123), 
        .A3(u5_mult_82_n4124), .ZN(u5_mult_82_CARRYB_6__28_) );
  NAND2_X1 u5_mult_82_U9197 ( .A1(u5_mult_82_CARRYB_5__28_), .A2(
        u5_mult_82_SUMB_5__29_), .ZN(u5_mult_82_n4124) );
  NAND2_X1 u5_mult_82_U9196 ( .A1(u5_mult_82_ab_6__28_), .A2(
        u5_mult_82_SUMB_5__29_), .ZN(u5_mult_82_n4123) );
  NAND2_X1 u5_mult_82_U9195 ( .A1(u5_mult_82_ab_6__28_), .A2(
        u5_mult_82_CARRYB_5__28_), .ZN(u5_mult_82_n4122) );
  NAND3_X2 u5_mult_82_U9194 ( .A1(u5_mult_82_n4119), .A2(u5_mult_82_n4120), 
        .A3(u5_mult_82_n4121), .ZN(u5_mult_82_CARRYB_24__10_) );
  NAND2_X1 u5_mult_82_U9193 ( .A1(u5_mult_82_CARRYB_23__10_), .A2(
        u5_mult_82_ab_24__10_), .ZN(u5_mult_82_n4119) );
  NAND3_X2 u5_mult_82_U9192 ( .A1(u5_mult_82_n4116), .A2(u5_mult_82_n4117), 
        .A3(u5_mult_82_n4118), .ZN(u5_mult_82_CARRYB_23__11_) );
  NAND2_X2 u5_mult_82_U9191 ( .A1(u5_mult_82_CARRYB_22__11_), .A2(
        u5_mult_82_SUMB_22__12_), .ZN(u5_mult_82_n4118) );
  NAND2_X2 u5_mult_82_U9190 ( .A1(u5_mult_82_ab_23__11_), .A2(
        u5_mult_82_SUMB_22__12_), .ZN(u5_mult_82_n4117) );
  XOR2_X2 u5_mult_82_U9189 ( .A(u5_mult_82_n4115), .B(u5_mult_82_SUMB_23__11_), 
        .Z(u5_mult_82_SUMB_24__10_) );
  NAND3_X2 u5_mult_82_U9188 ( .A1(u5_mult_82_n4112), .A2(u5_mult_82_n4113), 
        .A3(u5_mult_82_n4114), .ZN(u5_mult_82_CARRYB_18__16_) );
  NAND2_X1 u5_mult_82_U9187 ( .A1(u5_mult_82_CARRYB_17__16_), .A2(
        u5_mult_82_SUMB_17__17_), .ZN(u5_mult_82_n4114) );
  NAND2_X1 u5_mult_82_U9186 ( .A1(u5_mult_82_ab_18__16_), .A2(
        u5_mult_82_SUMB_17__17_), .ZN(u5_mult_82_n4113) );
  NAND3_X2 u5_mult_82_U9185 ( .A1(u5_mult_82_n4109), .A2(u5_mult_82_n4110), 
        .A3(u5_mult_82_n4111), .ZN(u5_mult_82_CARRYB_17__17_) );
  NAND2_X2 u5_mult_82_U9184 ( .A1(u5_mult_82_CARRYB_16__17_), .A2(
        u5_mult_82_SUMB_16__18_), .ZN(u5_mult_82_n4111) );
  NAND2_X2 u5_mult_82_U9183 ( .A1(u5_mult_82_ab_17__17_), .A2(
        u5_mult_82_SUMB_16__18_), .ZN(u5_mult_82_n4110) );
  NAND2_X1 u5_mult_82_U9182 ( .A1(u5_mult_82_ab_17__17_), .A2(
        u5_mult_82_CARRYB_16__17_), .ZN(u5_mult_82_n4109) );
  XOR2_X2 u5_mult_82_U9181 ( .A(u5_mult_82_n4108), .B(u5_mult_82_SUMB_17__17_), 
        .Z(u5_mult_82_SUMB_18__16_) );
  XOR2_X2 u5_mult_82_U9180 ( .A(u5_mult_82_n4107), .B(u5_mult_82_n1597), .Z(
        u5_mult_82_SUMB_17__17_) );
  NAND2_X1 u5_mult_82_U9179 ( .A1(u5_mult_82_ab_37__5_), .A2(
        u5_mult_82_CARRYB_36__5_), .ZN(u5_mult_82_n4106) );
  XNOR2_X2 u5_mult_82_U9178 ( .A(u5_mult_82_ab_44__21_), .B(
        u5_mult_82_SUMB_43__22_), .ZN(u5_mult_82_n4103) );
  XNOR2_X2 u5_mult_82_U9177 ( .A(u5_mult_82_n4103), .B(
        u5_mult_82_CARRYB_43__21_), .ZN(u5_mult_82_SUMB_44__21_) );
  NAND2_X2 u5_mult_82_U9176 ( .A1(u5_mult_82_ab_29__24_), .A2(
        u5_mult_82_SUMB_28__25_), .ZN(u5_mult_82_n6296) );
  NAND2_X2 u5_mult_82_U9175 ( .A1(u5_mult_82_ab_50__8_), .A2(
        u5_mult_82_SUMB_49__9_), .ZN(u5_mult_82_n6200) );
  NAND3_X4 u5_mult_82_U9174 ( .A1(u5_mult_82_n6131), .A2(u5_mult_82_n6132), 
        .A3(u5_mult_82_n6133), .ZN(u5_mult_82_CARRYB_42__9_) );
  INV_X1 u5_mult_82_U9173 ( .A(u5_mult_82_CARRYB_15__44_), .ZN(
        u5_mult_82_n5551) );
  XNOR2_X2 u5_mult_82_U9172 ( .A(u5_mult_82_n4102), .B(
        u5_mult_82_CARRYB_28__26_), .ZN(u5_mult_82_n6249) );
  INV_X8 u5_mult_82_U9171 ( .A(u5_mult_82_n4100), .ZN(u5_mult_82_n4101) );
  INV_X2 u5_mult_82_U9170 ( .A(u5_mult_82_SUMB_11__47_), .ZN(u5_mult_82_n4100)
         );
  XNOR2_X2 u5_mult_82_U9169 ( .A(u5_mult_82_CARRYB_41__4_), .B(
        u5_mult_82_ab_42__4_), .ZN(u5_mult_82_n4099) );
  NOR2_X1 u5_mult_82_U9168 ( .A1(u5_mult_82_net64665), .A2(u5_mult_82_n6741), 
        .ZN(u5_mult_82_ab_46__22_) );
  NAND3_X2 u5_mult_82_U9167 ( .A1(u5_mult_82_n4096), .A2(u5_mult_82_n4097), 
        .A3(u5_mult_82_n4098), .ZN(u5_mult_82_CARRYB_46__22_) );
  NAND2_X1 u5_mult_82_U9166 ( .A1(u5_mult_82_ab_46__22_), .A2(
        u5_mult_82_CARRYB_45__22_), .ZN(u5_mult_82_n4098) );
  NAND2_X2 u5_mult_82_U9165 ( .A1(u5_mult_82_ab_46__22_), .A2(
        u5_mult_82_SUMB_45__23_), .ZN(u5_mult_82_n4097) );
  NAND2_X1 u5_mult_82_U9164 ( .A1(u5_mult_82_CARRYB_45__22_), .A2(
        u5_mult_82_SUMB_45__23_), .ZN(u5_mult_82_n4096) );
  NAND3_X2 u5_mult_82_U9163 ( .A1(u5_mult_82_n4093), .A2(u5_mult_82_n4094), 
        .A3(u5_mult_82_n4095), .ZN(u5_mult_82_CARRYB_42__26_) );
  NAND2_X1 u5_mult_82_U9162 ( .A1(u5_mult_82_CARRYB_41__26_), .A2(
        u5_mult_82_SUMB_41__27_), .ZN(u5_mult_82_n4095) );
  NAND2_X1 u5_mult_82_U9161 ( .A1(u5_mult_82_ab_42__26_), .A2(
        u5_mult_82_SUMB_41__27_), .ZN(u5_mult_82_n4094) );
  NAND2_X1 u5_mult_82_U9160 ( .A1(u5_mult_82_ab_42__26_), .A2(
        u5_mult_82_CARRYB_41__26_), .ZN(u5_mult_82_n4093) );
  NAND2_X2 u5_mult_82_U9159 ( .A1(u5_mult_82_CARRYB_40__27_), .A2(
        u5_mult_82_n1730), .ZN(u5_mult_82_n4092) );
  NAND2_X2 u5_mult_82_U9158 ( .A1(u5_mult_82_ab_41__27_), .A2(u5_mult_82_n1730), .ZN(u5_mult_82_n4091) );
  NAND2_X1 u5_mult_82_U9157 ( .A1(u5_mult_82_ab_41__27_), .A2(
        u5_mult_82_CARRYB_40__27_), .ZN(u5_mult_82_n4090) );
  XOR2_X2 u5_mult_82_U9156 ( .A(u5_mult_82_n4089), .B(u5_mult_82_n1730), .Z(
        u5_mult_82_SUMB_41__27_) );
  XOR2_X2 u5_mult_82_U9155 ( .A(u5_mult_82_ab_41__27_), .B(
        u5_mult_82_CARRYB_40__27_), .Z(u5_mult_82_n4089) );
  NAND3_X2 u5_mult_82_U9154 ( .A1(u5_mult_82_n4086), .A2(u5_mult_82_n4087), 
        .A3(u5_mult_82_n4088), .ZN(u5_mult_82_CARRYB_36__31_) );
  NAND2_X1 u5_mult_82_U9153 ( .A1(u5_mult_82_CARRYB_35__31_), .A2(
        u5_mult_82_SUMB_35__32_), .ZN(u5_mult_82_n4088) );
  NAND2_X1 u5_mult_82_U9152 ( .A1(u5_mult_82_ab_36__31_), .A2(
        u5_mult_82_SUMB_35__32_), .ZN(u5_mult_82_n4087) );
  NAND2_X1 u5_mult_82_U9151 ( .A1(u5_mult_82_ab_36__31_), .A2(
        u5_mult_82_CARRYB_35__31_), .ZN(u5_mult_82_n4086) );
  NAND3_X2 u5_mult_82_U9150 ( .A1(u5_mult_82_n4083), .A2(u5_mult_82_n4084), 
        .A3(u5_mult_82_n4085), .ZN(u5_mult_82_CARRYB_35__32_) );
  NAND2_X2 u5_mult_82_U9149 ( .A1(u5_mult_82_CARRYB_34__32_), .A2(
        u5_mult_82_n1575), .ZN(u5_mult_82_n4085) );
  NAND2_X2 u5_mult_82_U9148 ( .A1(u5_mult_82_ab_35__32_), .A2(u5_mult_82_n1575), .ZN(u5_mult_82_n4084) );
  NAND2_X1 u5_mult_82_U9147 ( .A1(u5_mult_82_ab_35__32_), .A2(
        u5_mult_82_CARRYB_34__32_), .ZN(u5_mult_82_n4083) );
  XOR2_X2 u5_mult_82_U9146 ( .A(u5_mult_82_n4082), .B(u5_mult_82_SUMB_35__32_), 
        .Z(u5_mult_82_SUMB_36__31_) );
  XOR2_X2 u5_mult_82_U9145 ( .A(u5_mult_82_ab_36__31_), .B(
        u5_mult_82_CARRYB_35__31_), .Z(u5_mult_82_n4082) );
  XOR2_X2 u5_mult_82_U9144 ( .A(u5_mult_82_n4081), .B(u5_mult_82_n1575), .Z(
        u5_mult_82_SUMB_35__32_) );
  XOR2_X2 u5_mult_82_U9143 ( .A(u5_mult_82_ab_35__32_), .B(
        u5_mult_82_CARRYB_34__32_), .Z(u5_mult_82_n4081) );
  NAND2_X2 u5_mult_82_U9142 ( .A1(u5_mult_82_ab_43__9_), .A2(
        u5_mult_82_SUMB_42__10_), .ZN(u5_mult_82_n5489) );
  XOR2_X2 u5_mult_82_U9141 ( .A(u5_mult_82_n5127), .B(u5_mult_82_SUMB_37__13_), 
        .Z(u5_mult_82_SUMB_38__12_) );
  INV_X8 u5_mult_82_U9140 ( .A(n4746), .ZN(u5_mult_82_n7012) );
  XNOR2_X2 u5_mult_82_U9139 ( .A(u5_mult_82_ab_35__14_), .B(
        u5_mult_82_CARRYB_34__14_), .ZN(u5_mult_82_n4079) );
  NAND3_X4 u5_mult_82_U9138 ( .A1(u5_mult_82_n6375), .A2(u5_mult_82_n6376), 
        .A3(u5_mult_82_n6377), .ZN(u5_mult_82_CARRYB_23__34_) );
  NAND2_X2 u5_mult_82_U9137 ( .A1(u5_mult_82_CARRYB_24__33_), .A2(
        u5_mult_82_SUMB_24__34_), .ZN(u5_mult_82_n6229) );
  NOR2_X1 u5_mult_82_U9136 ( .A1(u5_mult_82_net64451), .A2(u5_mult_82_net65517), .ZN(u5_mult_82_ab_34__10_) );
  NAND2_X1 u5_mult_82_U9135 ( .A1(u5_mult_82_CARRYB_35__8_), .A2(
        u5_mult_82_SUMB_35__9_), .ZN(u5_mult_82_n4078) );
  NAND2_X1 u5_mult_82_U9134 ( .A1(u5_mult_82_ab_36__8_), .A2(
        u5_mult_82_SUMB_35__9_), .ZN(u5_mult_82_n4077) );
  NAND2_X1 u5_mult_82_U9133 ( .A1(u5_mult_82_ab_36__8_), .A2(
        u5_mult_82_CARRYB_35__8_), .ZN(u5_mult_82_n4076) );
  NAND3_X2 u5_mult_82_U9132 ( .A1(u5_mult_82_n4073), .A2(u5_mult_82_n4074), 
        .A3(u5_mult_82_n4075), .ZN(u5_mult_82_CARRYB_35__9_) );
  NAND2_X2 u5_mult_82_U9131 ( .A1(u5_mult_82_CARRYB_34__9_), .A2(
        u5_mult_82_SUMB_34__10_), .ZN(u5_mult_82_n4075) );
  NAND2_X2 u5_mult_82_U9130 ( .A1(u5_mult_82_ab_35__9_), .A2(
        u5_mult_82_SUMB_34__10_), .ZN(u5_mult_82_n4074) );
  NAND2_X1 u5_mult_82_U9129 ( .A1(u5_mult_82_ab_35__9_), .A2(
        u5_mult_82_CARRYB_34__9_), .ZN(u5_mult_82_n4073) );
  NAND3_X2 u5_mult_82_U9128 ( .A1(u5_mult_82_n4070), .A2(u5_mult_82_n4071), 
        .A3(u5_mult_82_n4072), .ZN(u5_mult_82_CARRYB_34__10_) );
  XOR2_X2 u5_mult_82_U9127 ( .A(u5_mult_82_n1442), .B(u5_mult_82_n5090), .Z(
        u5_mult_82_SUMB_21__49_) );
  NAND2_X1 u5_mult_82_U9126 ( .A1(u5_mult_82_ab_33__14_), .A2(
        u5_mult_82_SUMB_32__15_), .ZN(u5_mult_82_n5919) );
  XOR2_X2 u5_mult_82_U9125 ( .A(u5_mult_82_CARRYB_9__26_), .B(u5_mult_82_n4279), .Z(u5_mult_82_n4069) );
  XNOR2_X2 u5_mult_82_U9124 ( .A(u5_mult_82_n382), .B(u5_mult_82_n4069), .ZN(
        u5_mult_82_SUMB_10__26_) );
  XNOR2_X2 u5_mult_82_U9123 ( .A(u5_mult_82_ab_34__14_), .B(
        u5_mult_82_CARRYB_33__14_), .ZN(u5_mult_82_n4068) );
  XNOR2_X2 u5_mult_82_U9122 ( .A(u5_mult_82_n4068), .B(u5_mult_82_SUMB_33__15_), .ZN(u5_mult_82_SUMB_34__14_) );
  NAND3_X4 u5_mult_82_U9121 ( .A1(u5_mult_82_n4464), .A2(u5_mult_82_n4465), 
        .A3(u5_mult_82_n4466), .ZN(u5_mult_82_CARRYB_50__25_) );
  XOR2_X2 u5_mult_82_U9120 ( .A(u5_mult_82_CARRYB_46__4_), .B(
        u5_mult_82_ab_47__4_), .Z(u5_mult_82_n6134) );
  NOR2_X1 u5_mult_82_U9119 ( .A1(u5_mult_82_net64525), .A2(u5_mult_82_n6651), 
        .ZN(u5_mult_82_ab_26__14_) );
  NAND3_X2 u5_mult_82_U9118 ( .A1(u5_mult_82_n4065), .A2(u5_mult_82_n4066), 
        .A3(u5_mult_82_n4067), .ZN(u5_mult_82_CARRYB_26__14_) );
  NAND2_X1 u5_mult_82_U9117 ( .A1(u5_mult_82_ab_26__14_), .A2(
        u5_mult_82_CARRYB_25__14_), .ZN(u5_mult_82_n4067) );
  NAND3_X2 u5_mult_82_U9116 ( .A1(u5_mult_82_n4062), .A2(u5_mult_82_n4063), 
        .A3(u5_mult_82_n4064), .ZN(u5_mult_82_CARRYB_29__11_) );
  NAND2_X1 u5_mult_82_U9115 ( .A1(u5_mult_82_CARRYB_28__11_), .A2(
        u5_mult_82_SUMB_28__12_), .ZN(u5_mult_82_n4064) );
  NAND2_X1 u5_mult_82_U9114 ( .A1(u5_mult_82_ab_29__11_), .A2(
        u5_mult_82_SUMB_28__12_), .ZN(u5_mult_82_n4063) );
  NAND2_X1 u5_mult_82_U9113 ( .A1(u5_mult_82_ab_29__11_), .A2(
        u5_mult_82_CARRYB_28__11_), .ZN(u5_mult_82_n4062) );
  NAND3_X2 u5_mult_82_U9112 ( .A1(u5_mult_82_n4059), .A2(u5_mult_82_n4060), 
        .A3(u5_mult_82_n4061), .ZN(u5_mult_82_CARRYB_28__12_) );
  NAND2_X1 u5_mult_82_U9111 ( .A1(u5_mult_82_CARRYB_27__12_), .A2(
        u5_mult_82_SUMB_27__13_), .ZN(u5_mult_82_n4061) );
  NAND2_X1 u5_mult_82_U9110 ( .A1(u5_mult_82_ab_28__12_), .A2(
        u5_mult_82_SUMB_27__13_), .ZN(u5_mult_82_n4060) );
  NAND2_X1 u5_mult_82_U9109 ( .A1(u5_mult_82_ab_28__12_), .A2(
        u5_mult_82_CARRYB_27__12_), .ZN(u5_mult_82_n4059) );
  XOR2_X2 u5_mult_82_U9108 ( .A(u5_mult_82_n4058), .B(u5_mult_82_SUMB_27__13_), 
        .Z(u5_mult_82_SUMB_28__12_) );
  XOR2_X2 u5_mult_82_U9107 ( .A(u5_mult_82_CARRYB_27__12_), .B(
        u5_mult_82_ab_28__12_), .Z(u5_mult_82_n4058) );
  XNOR2_X2 u5_mult_82_U9106 ( .A(u5_mult_82_ab_43__14_), .B(
        u5_mult_82_CARRYB_42__14_), .ZN(u5_mult_82_n4057) );
  XNOR2_X2 u5_mult_82_U9105 ( .A(u5_mult_82_n4057), .B(u5_mult_82_SUMB_42__15_), .ZN(u5_mult_82_SUMB_43__14_) );
  NOR2_X1 u5_mult_82_U9104 ( .A1(u5_mult_82_net64361), .A2(u5_mult_82_n6665), 
        .ZN(u5_mult_82_ab_28__5_) );
  NOR2_X2 u5_mult_82_U9103 ( .A1(u5_mult_82_net64561), .A2(u5_mult_82_n6602), 
        .ZN(u5_mult_82_ab_17__16_) );
  NAND3_X2 u5_mult_82_U9102 ( .A1(u5_mult_82_n4054), .A2(u5_mult_82_n4055), 
        .A3(u5_mult_82_n4056), .ZN(u5_mult_82_CARRYB_28__5_) );
  NAND2_X2 u5_mult_82_U9101 ( .A1(u5_mult_82_ab_28__5_), .A2(
        u5_mult_82_SUMB_27__6_), .ZN(u5_mult_82_n4055) );
  NAND2_X1 u5_mult_82_U9100 ( .A1(u5_mult_82_CARRYB_27__5_), .A2(
        u5_mult_82_SUMB_27__6_), .ZN(u5_mult_82_n4054) );
  XOR2_X2 u5_mult_82_U9099 ( .A(u5_mult_82_n4053), .B(u5_mult_82_SUMB_27__6_), 
        .Z(u5_mult_82_SUMB_28__5_) );
  NAND3_X2 u5_mult_82_U9098 ( .A1(u5_mult_82_n4050), .A2(u5_mult_82_n4051), 
        .A3(u5_mult_82_n4052), .ZN(u5_mult_82_CARRYB_9__24_) );
  NAND2_X1 u5_mult_82_U9097 ( .A1(u5_mult_82_CARRYB_8__24_), .A2(
        u5_mult_82_SUMB_8__25_), .ZN(u5_mult_82_n4052) );
  NAND2_X1 u5_mult_82_U9096 ( .A1(u5_mult_82_ab_9__24_), .A2(
        u5_mult_82_SUMB_8__25_), .ZN(u5_mult_82_n4051) );
  NAND2_X1 u5_mult_82_U9095 ( .A1(u5_mult_82_ab_9__24_), .A2(
        u5_mult_82_CARRYB_8__24_), .ZN(u5_mult_82_n4050) );
  NAND3_X2 u5_mult_82_U9094 ( .A1(u5_mult_82_n4047), .A2(u5_mult_82_n4048), 
        .A3(u5_mult_82_n4049), .ZN(u5_mult_82_CARRYB_8__25_) );
  NAND2_X2 u5_mult_82_U9093 ( .A1(u5_mult_82_CARRYB_7__25_), .A2(
        u5_mult_82_SUMB_7__26_), .ZN(u5_mult_82_n4049) );
  NAND2_X2 u5_mult_82_U9092 ( .A1(u5_mult_82_ab_8__25_), .A2(
        u5_mult_82_SUMB_7__26_), .ZN(u5_mult_82_n4048) );
  NAND2_X1 u5_mult_82_U9091 ( .A1(u5_mult_82_ab_8__25_), .A2(
        u5_mult_82_CARRYB_7__25_), .ZN(u5_mult_82_n4047) );
  XOR2_X2 u5_mult_82_U9090 ( .A(u5_mult_82_ab_9__24_), .B(
        u5_mult_82_CARRYB_8__24_), .Z(u5_mult_82_n4046) );
  XOR2_X2 u5_mult_82_U9089 ( .A(u5_mult_82_n4045), .B(u5_mult_82_SUMB_7__26_), 
        .Z(u5_mult_82_SUMB_8__25_) );
  XOR2_X2 u5_mult_82_U9088 ( .A(u5_mult_82_ab_8__25_), .B(
        u5_mult_82_CARRYB_7__25_), .Z(u5_mult_82_n4045) );
  NAND3_X2 u5_mult_82_U9087 ( .A1(u5_mult_82_n4042), .A2(u5_mult_82_n4043), 
        .A3(u5_mult_82_n4044), .ZN(u5_mult_82_CARRYB_5__28_) );
  NAND2_X1 u5_mult_82_U9086 ( .A1(u5_mult_82_CARRYB_4__28_), .A2(
        u5_mult_82_SUMB_4__29_), .ZN(u5_mult_82_n4044) );
  NAND2_X1 u5_mult_82_U9085 ( .A1(u5_mult_82_ab_5__28_), .A2(
        u5_mult_82_SUMB_4__29_), .ZN(u5_mult_82_n4043) );
  NAND2_X1 u5_mult_82_U9084 ( .A1(u5_mult_82_ab_5__28_), .A2(
        u5_mult_82_CARRYB_4__28_), .ZN(u5_mult_82_n4042) );
  NAND3_X2 u5_mult_82_U9083 ( .A1(u5_mult_82_n4039), .A2(u5_mult_82_n4040), 
        .A3(u5_mult_82_n4041), .ZN(u5_mult_82_CARRYB_4__29_) );
  NAND2_X1 u5_mult_82_U9082 ( .A1(u5_mult_82_CARRYB_3__29_), .A2(
        u5_mult_82_SUMB_3__30_), .ZN(u5_mult_82_n4041) );
  NAND2_X1 u5_mult_82_U9081 ( .A1(u5_mult_82_ab_4__29_), .A2(
        u5_mult_82_SUMB_3__30_), .ZN(u5_mult_82_n4040) );
  NAND2_X1 u5_mult_82_U9080 ( .A1(u5_mult_82_ab_4__29_), .A2(
        u5_mult_82_CARRYB_3__29_), .ZN(u5_mult_82_n4039) );
  XOR2_X2 u5_mult_82_U9079 ( .A(u5_mult_82_n4038), .B(u5_mult_82_SUMB_4__29_), 
        .Z(u5_mult_82_SUMB_5__28_) );
  XOR2_X2 u5_mult_82_U9078 ( .A(u5_mult_82_n4037), .B(u5_mult_82_SUMB_3__30_), 
        .Z(u5_mult_82_SUMB_4__29_) );
  XOR2_X2 u5_mult_82_U9077 ( .A(u5_mult_82_ab_4__29_), .B(
        u5_mult_82_CARRYB_3__29_), .Z(u5_mult_82_n4037) );
  NAND3_X2 u5_mult_82_U9076 ( .A1(u5_mult_82_n4034), .A2(u5_mult_82_n4035), 
        .A3(u5_mult_82_n4036), .ZN(u5_mult_82_CARRYB_19__14_) );
  NAND2_X1 u5_mult_82_U9075 ( .A1(u5_mult_82_CARRYB_18__14_), .A2(
        u5_mult_82_SUMB_18__15_), .ZN(u5_mult_82_n4036) );
  NAND2_X1 u5_mult_82_U9074 ( .A1(u5_mult_82_ab_19__14_), .A2(
        u5_mult_82_SUMB_18__15_), .ZN(u5_mult_82_n4035) );
  NAND2_X1 u5_mult_82_U9073 ( .A1(u5_mult_82_ab_19__14_), .A2(
        u5_mult_82_CARRYB_18__14_), .ZN(u5_mult_82_n4034) );
  NAND3_X2 u5_mult_82_U9072 ( .A1(u5_mult_82_n4031), .A2(u5_mult_82_n4032), 
        .A3(u5_mult_82_n4033), .ZN(u5_mult_82_CARRYB_18__15_) );
  NAND2_X2 u5_mult_82_U9071 ( .A1(u5_mult_82_CARRYB_17__15_), .A2(
        u5_mult_82_SUMB_17__16_), .ZN(u5_mult_82_n4033) );
  NAND2_X2 u5_mult_82_U9070 ( .A1(u5_mult_82_ab_18__15_), .A2(
        u5_mult_82_SUMB_17__16_), .ZN(u5_mult_82_n4032) );
  NAND2_X1 u5_mult_82_U9069 ( .A1(u5_mult_82_ab_18__15_), .A2(
        u5_mult_82_CARRYB_17__15_), .ZN(u5_mult_82_n4031) );
  XOR2_X2 u5_mult_82_U9068 ( .A(u5_mult_82_n4030), .B(u5_mult_82_SUMB_18__15_), 
        .Z(u5_mult_82_SUMB_19__14_) );
  XOR2_X2 u5_mult_82_U9067 ( .A(u5_mult_82_ab_19__14_), .B(
        u5_mult_82_CARRYB_18__14_), .Z(u5_mult_82_n4030) );
  XOR2_X2 u5_mult_82_U9066 ( .A(u5_mult_82_n4029), .B(u5_mult_82_SUMB_17__16_), 
        .Z(u5_mult_82_SUMB_18__15_) );
  XOR2_X2 u5_mult_82_U9065 ( .A(u5_mult_82_ab_18__15_), .B(
        u5_mult_82_CARRYB_17__15_), .Z(u5_mult_82_n4029) );
  NAND2_X1 u5_mult_82_U9064 ( .A1(u5_mult_82_ab_17__16_), .A2(
        u5_mult_82_CARRYB_16__16_), .ZN(u5_mult_82_n4028) );
  XOR2_X2 u5_mult_82_U9063 ( .A(u5_mult_82_SUMB_16__17_), .B(u5_mult_82_n4025), 
        .Z(u5_mult_82_SUMB_17__16_) );
  XOR2_X2 u5_mult_82_U9062 ( .A(u5_mult_82_CARRYB_16__16_), .B(
        u5_mult_82_ab_17__16_), .Z(u5_mult_82_n4025) );
  NAND3_X4 u5_mult_82_U9061 ( .A1(u5_mult_82_n5368), .A2(u5_mult_82_n5369), 
        .A3(u5_mult_82_n5370), .ZN(u5_mult_82_CARRYB_12__41_) );
  NAND3_X4 u5_mult_82_U9060 ( .A1(u5_mult_82_n5471), .A2(u5_mult_82_n5472), 
        .A3(u5_mult_82_n5473), .ZN(u5_mult_82_CARRYB_24__33_) );
  XNOR2_X2 u5_mult_82_U9059 ( .A(u5_mult_82_ab_36__23_), .B(
        u5_mult_82_CARRYB_35__23_), .ZN(u5_mult_82_n4024) );
  XNOR2_X2 u5_mult_82_U9058 ( .A(u5_mult_82_n4024), .B(u5_mult_82_SUMB_35__24_), .ZN(u5_mult_82_SUMB_36__23_) );
  XNOR2_X2 u5_mult_82_U9057 ( .A(u5_mult_82_ab_17__24_), .B(
        u5_mult_82_CARRYB_16__24_), .ZN(u5_mult_82_n4023) );
  NOR2_X1 u5_mult_82_U9056 ( .A1(u5_mult_82_n6829), .A2(u5_mult_82_n6528), 
        .ZN(u5_mult_82_ab_7__40_) );
  NAND2_X2 u5_mult_82_U9055 ( .A1(u5_mult_82_ab_16__34_), .A2(
        u5_mult_82_CARRYB_15__34_), .ZN(u5_mult_82_n5054) );
  NOR2_X2 u5_mult_82_U9054 ( .A1(u5_mult_82_net64887), .A2(u5_mult_82_n6586), 
        .ZN(u5_mult_82_ab_15__34_) );
  NAND2_X2 u5_mult_82_U9053 ( .A1(u5_mult_82_CARRYB_45__17_), .A2(
        u5_mult_82_SUMB_45__18_), .ZN(u5_mult_82_n5863) );
  NOR2_X1 u5_mult_82_U9052 ( .A1(u5_mult_82_n6927), .A2(u5_mult_82_net65321), 
        .ZN(u5_mult_82_ab_45__17_) );
  NOR2_X1 u5_mult_82_U9051 ( .A1(u5_mult_82_net64959), .A2(u5_mult_82_n6550), 
        .ZN(u5_mult_82_ab_10__38_) );
  NOR2_X1 u5_mult_82_U9050 ( .A1(u5_mult_82_net64685), .A2(u5_mult_82_n6700), 
        .ZN(u5_mult_82_ab_33__23_) );
  NOR2_X1 u5_mult_82_U9049 ( .A1(u5_mult_82_n6858), .A2(u5_mult_82_n6621), 
        .ZN(u5_mult_82_ab_20__30_) );
  NOR2_X1 u5_mult_82_U9048 ( .A1(u5_mult_82_n6896), .A2(u5_mult_82_net65443), 
        .ZN(u5_mult_82_ab_38__21_) );
  NAND3_X2 u5_mult_82_U9047 ( .A1(u5_mult_82_n4020), .A2(u5_mult_82_n4021), 
        .A3(u5_mult_82_n4022), .ZN(u5_mult_82_CARRYB_7__40_) );
  NAND2_X1 u5_mult_82_U9046 ( .A1(u5_mult_82_ab_7__40_), .A2(
        u5_mult_82_CARRYB_6__40_), .ZN(u5_mult_82_n4022) );
  NAND3_X4 u5_mult_82_U9045 ( .A1(u5_mult_82_n4016), .A2(u5_mult_82_n4017), 
        .A3(u5_mult_82_n4018), .ZN(u5_mult_82_CARRYB_15__34_) );
  NAND2_X1 u5_mult_82_U9044 ( .A1(u5_mult_82_ab_15__34_), .A2(
        u5_mult_82_CARRYB_14__34_), .ZN(u5_mult_82_n4018) );
  NAND2_X2 u5_mult_82_U9043 ( .A1(u5_mult_82_CARRYB_14__34_), .A2(
        u5_mult_82_n1616), .ZN(u5_mult_82_n4016) );
  NAND3_X2 u5_mult_82_U9042 ( .A1(u5_mult_82_n4013), .A2(u5_mult_82_n4014), 
        .A3(u5_mult_82_n4015), .ZN(u5_mult_82_CARRYB_45__17_) );
  NAND2_X2 u5_mult_82_U9041 ( .A1(u5_mult_82_ab_45__17_), .A2(
        u5_mult_82_CARRYB_44__17_), .ZN(u5_mult_82_n4014) );
  NAND3_X2 u5_mult_82_U9040 ( .A1(u5_mult_82_n4010), .A2(u5_mult_82_n4011), 
        .A3(u5_mult_82_n4012), .ZN(u5_mult_82_CARRYB_10__38_) );
  NAND2_X1 u5_mult_82_U9039 ( .A1(u5_mult_82_ab_10__38_), .A2(
        u5_mult_82_CARRYB_9__38_), .ZN(u5_mult_82_n4012) );
  NAND2_X1 u5_mult_82_U9038 ( .A1(u5_mult_82_CARRYB_9__38_), .A2(
        u5_mult_82_SUMB_9__39_), .ZN(u5_mult_82_n4010) );
  NAND3_X2 u5_mult_82_U9037 ( .A1(u5_mult_82_n4007), .A2(u5_mult_82_n4008), 
        .A3(u5_mult_82_n4009), .ZN(u5_mult_82_CARRYB_33__23_) );
  NAND2_X1 u5_mult_82_U9036 ( .A1(u5_mult_82_SUMB_32__24_), .A2(
        u5_mult_82_CARRYB_32__23_), .ZN(u5_mult_82_n4007) );
  NAND3_X2 u5_mult_82_U9035 ( .A1(u5_mult_82_n4004), .A2(u5_mult_82_n4005), 
        .A3(u5_mult_82_n4006), .ZN(u5_mult_82_CARRYB_20__30_) );
  NAND2_X1 u5_mult_82_U9034 ( .A1(u5_mult_82_ab_20__30_), .A2(
        u5_mult_82_CARRYB_19__30_), .ZN(u5_mult_82_n4006) );
  NAND2_X2 u5_mult_82_U9033 ( .A1(u5_mult_82_ab_20__30_), .A2(
        u5_mult_82_SUMB_19__31_), .ZN(u5_mult_82_n4005) );
  NAND2_X1 u5_mult_82_U9032 ( .A1(u5_mult_82_CARRYB_19__30_), .A2(
        u5_mult_82_SUMB_19__31_), .ZN(u5_mult_82_n4004) );
  NAND3_X2 u5_mult_82_U9031 ( .A1(u5_mult_82_n4001), .A2(u5_mult_82_n4002), 
        .A3(u5_mult_82_n4003), .ZN(u5_mult_82_CARRYB_38__21_) );
  NAND2_X1 u5_mult_82_U9030 ( .A1(u5_mult_82_SUMB_37__22_), .A2(
        u5_mult_82_CARRYB_37__21_), .ZN(u5_mult_82_n4001) );
  XOR2_X2 u5_mult_82_U9029 ( .A(u5_mult_82_n4000), .B(u5_mult_82_n1444), .Z(
        u5_mult_82_SUMB_38__21_) );
  XOR2_X2 u5_mult_82_U9028 ( .A(u5_mult_82_SUMB_37__22_), .B(
        u5_mult_82_ab_38__21_), .Z(u5_mult_82_n4000) );
  XOR2_X2 u5_mult_82_U9027 ( .A(u5_mult_82_SUMB_20__50_), .B(
        u5_mult_82_ab_21__49_), .Z(u5_mult_82_n5090) );
  XNOR2_X2 u5_mult_82_U9026 ( .A(u5_mult_82_CARRYB_6__40_), .B(
        u5_mult_82_n3999), .ZN(u5_mult_82_n4019) );
  NAND2_X1 u5_mult_82_U9025 ( .A1(u5_mult_82_CARRYB_7__40_), .A2(
        u5_mult_82_SUMB_7__41_), .ZN(u5_mult_82_n6023) );
  NAND2_X1 u5_mult_82_U9024 ( .A1(u5_mult_82_CARRYB_32__14_), .A2(
        u5_mult_82_SUMB_32__15_), .ZN(u5_mult_82_n5920) );
  NAND2_X2 u5_mult_82_U9023 ( .A1(u5_mult_82_ab_33__14_), .A2(
        u5_mult_82_CARRYB_32__14_), .ZN(u5_mult_82_n5918) );
  NOR2_X2 u5_mult_82_U9022 ( .A1(u5_mult_82_net64523), .A2(u5_mult_82_n6695), 
        .ZN(u5_mult_82_ab_32__14_) );
  NOR2_X1 u5_mult_82_U9021 ( .A1(u5_mult_82_net64451), .A2(u5_mult_82_n6729), 
        .ZN(u5_mult_82_ab_39__10_) );
  NAND3_X4 u5_mult_82_U9020 ( .A1(u5_mult_82_n3996), .A2(u5_mult_82_n3997), 
        .A3(u5_mult_82_n3998), .ZN(u5_mult_82_CARRYB_32__14_) );
  NAND2_X2 u5_mult_82_U9019 ( .A1(u5_mult_82_ab_32__14_), .A2(
        u5_mult_82_SUMB_31__15_), .ZN(u5_mult_82_n3997) );
  NAND2_X2 u5_mult_82_U9018 ( .A1(u5_mult_82_CARRYB_31__14_), .A2(
        u5_mult_82_SUMB_31__15_), .ZN(u5_mult_82_n3996) );
  NAND3_X2 u5_mult_82_U9017 ( .A1(u5_mult_82_n3994), .A2(u5_mult_82_n3993), 
        .A3(u5_mult_82_n3995), .ZN(u5_mult_82_CARRYB_39__10_) );
  NAND2_X1 u5_mult_82_U9016 ( .A1(u5_mult_82_ab_39__10_), .A2(
        u5_mult_82_CARRYB_38__10_), .ZN(u5_mult_82_n3995) );
  NAND2_X2 u5_mult_82_U9015 ( .A1(u5_mult_82_ab_39__10_), .A2(
        u5_mult_82_SUMB_38__11_), .ZN(u5_mult_82_n3994) );
  NAND2_X2 u5_mult_82_U9014 ( .A1(u5_mult_82_ab_44__5_), .A2(
        u5_mult_82_CARRYB_43__5_), .ZN(u5_mult_82_n6035) );
  XOR2_X2 u5_mult_82_U9013 ( .A(u5_mult_82_n6308), .B(u5_mult_82_SUMB_16__37_), 
        .Z(u5_mult_82_SUMB_17__36_) );
  XOR2_X2 u5_mult_82_U9012 ( .A(u5_mult_82_CARRYB_20__29_), .B(
        u5_mult_82_ab_21__29_), .Z(u5_mult_82_n5057) );
  NAND3_X2 u5_mult_82_U9011 ( .A1(u5_mult_82_n6291), .A2(u5_mult_82_n6292), 
        .A3(u5_mult_82_n6293), .ZN(u5_mult_82_CARRYB_5__50_) );
  NAND3_X2 u5_mult_82_U9010 ( .A1(u5_mult_82_n3991), .A2(u5_mult_82_net82468), 
        .A3(u5_mult_82_net82469), .ZN(u5_mult_82_CARRYB_39__13_) );
  NAND2_X2 u5_mult_82_U9009 ( .A1(u5_mult_82_CARRYB_25__34_), .A2(
        u5_mult_82_SUMB_25__35_), .ZN(u5_mult_82_n4439) );
  NAND3_X2 u5_mult_82_U9008 ( .A1(u5_mult_82_n3988), .A2(u5_mult_82_n3989), 
        .A3(u5_mult_82_n3990), .ZN(u5_mult_82_CARRYB_8__24_) );
  NAND2_X1 u5_mult_82_U9007 ( .A1(u5_mult_82_ab_8__24_), .A2(
        u5_mult_82_SUMB_7__25_), .ZN(u5_mult_82_n3989) );
  NAND3_X4 u5_mult_82_U9006 ( .A1(u5_mult_82_n3985), .A2(u5_mult_82_n3986), 
        .A3(u5_mult_82_n3987), .ZN(u5_mult_82_CARRYB_7__25_) );
  NAND2_X2 u5_mult_82_U9005 ( .A1(u5_mult_82_CARRYB_6__25_), .A2(
        u5_mult_82_SUMB_6__26_), .ZN(u5_mult_82_n3987) );
  NAND2_X2 u5_mult_82_U9004 ( .A1(u5_mult_82_ab_7__25_), .A2(
        u5_mult_82_SUMB_6__26_), .ZN(u5_mult_82_n3986) );
  XOR2_X2 u5_mult_82_U9003 ( .A(u5_mult_82_n3984), .B(u5_mult_82_SUMB_7__25_), 
        .Z(u5_mult_82_SUMB_8__24_) );
  XOR2_X2 u5_mult_82_U9002 ( .A(u5_mult_82_ab_8__24_), .B(
        u5_mult_82_CARRYB_7__24_), .Z(u5_mult_82_n3984) );
  NAND3_X2 u5_mult_82_U9001 ( .A1(u5_mult_82_n3981), .A2(u5_mult_82_n3982), 
        .A3(u5_mult_82_n3983), .ZN(u5_mult_82_CARRYB_5__27_) );
  NAND3_X4 u5_mult_82_U9000 ( .A1(u5_mult_82_n3978), .A2(u5_mult_82_n3979), 
        .A3(u5_mult_82_n3980), .ZN(u5_mult_82_CARRYB_4__28_) );
  NAND2_X2 u5_mult_82_U8999 ( .A1(u5_mult_82_CARRYB_3__28_), .A2(
        u5_mult_82_SUMB_3__29_), .ZN(u5_mult_82_n3980) );
  NAND2_X2 u5_mult_82_U8998 ( .A1(u5_mult_82_ab_4__28_), .A2(
        u5_mult_82_SUMB_3__29_), .ZN(u5_mult_82_n3979) );
  NAND2_X1 u5_mult_82_U8997 ( .A1(u5_mult_82_ab_4__28_), .A2(
        u5_mult_82_CARRYB_3__28_), .ZN(u5_mult_82_n3978) );
  XOR2_X2 u5_mult_82_U8996 ( .A(u5_mult_82_n3977), .B(u5_mult_82_SUMB_3__29_), 
        .Z(u5_mult_82_SUMB_4__28_) );
  XOR2_X2 u5_mult_82_U8995 ( .A(u5_mult_82_ab_4__28_), .B(
        u5_mult_82_CARRYB_3__28_), .Z(u5_mult_82_n3977) );
  NAND3_X2 u5_mult_82_U8994 ( .A1(u5_mult_82_n3974), .A2(u5_mult_82_n3975), 
        .A3(u5_mult_82_n3976), .ZN(u5_mult_82_CARRYB_17__15_) );
  NAND2_X1 u5_mult_82_U8993 ( .A1(u5_mult_82_CARRYB_16__15_), .A2(
        u5_mult_82_SUMB_16__16_), .ZN(u5_mult_82_n3976) );
  NAND2_X1 u5_mult_82_U8992 ( .A1(u5_mult_82_ab_17__15_), .A2(
        u5_mult_82_SUMB_16__16_), .ZN(u5_mult_82_n3975) );
  NAND2_X1 u5_mult_82_U8991 ( .A1(u5_mult_82_ab_17__15_), .A2(
        u5_mult_82_CARRYB_16__15_), .ZN(u5_mult_82_n3974) );
  NAND3_X4 u5_mult_82_U8990 ( .A1(u5_mult_82_n3971), .A2(u5_mult_82_n3972), 
        .A3(u5_mult_82_n3973), .ZN(u5_mult_82_CARRYB_16__16_) );
  NAND2_X2 u5_mult_82_U8989 ( .A1(u5_mult_82_CARRYB_15__16_), .A2(
        u5_mult_82_n1651), .ZN(u5_mult_82_n3973) );
  NAND2_X2 u5_mult_82_U8988 ( .A1(u5_mult_82_ab_16__16_), .A2(u5_mult_82_n1651), .ZN(u5_mult_82_n3972) );
  NAND2_X1 u5_mult_82_U8987 ( .A1(u5_mult_82_ab_16__16_), .A2(
        u5_mult_82_CARRYB_15__16_), .ZN(u5_mult_82_n3971) );
  XOR2_X2 u5_mult_82_U8986 ( .A(u5_mult_82_n3970), .B(u5_mult_82_SUMB_16__16_), 
        .Z(u5_mult_82_SUMB_17__15_) );
  XNOR2_X2 u5_mult_82_U8985 ( .A(u5_mult_82_ab_15__48_), .B(
        u5_mult_82_CARRYB_14__48_), .ZN(u5_mult_82_n3969) );
  XNOR2_X2 u5_mult_82_U8984 ( .A(u5_mult_82_ab_4__38_), .B(
        u5_mult_82_CARRYB_3__38_), .ZN(u5_mult_82_n3968) );
  XNOR2_X2 u5_mult_82_U8983 ( .A(u5_mult_82_n3968), .B(u5_mult_82_SUMB_3__39_), 
        .ZN(u5_mult_82_SUMB_4__38_) );
  XNOR2_X2 u5_mult_82_U8982 ( .A(u5_mult_82_n3967), .B(u5_mult_82_SUMB_15__33_), .ZN(u5_mult_82_SUMB_16__32_) );
  NAND3_X2 u5_mult_82_U8981 ( .A1(u5_mult_82_n3964), .A2(u5_mult_82_n3965), 
        .A3(u5_mult_82_n3966), .ZN(u5_mult_82_CARRYB_39__6_) );
  NAND2_X1 u5_mult_82_U8980 ( .A1(u5_mult_82_CARRYB_38__6_), .A2(
        u5_mult_82_SUMB_38__7_), .ZN(u5_mult_82_n3966) );
  NAND2_X1 u5_mult_82_U8979 ( .A1(u5_mult_82_ab_39__6_), .A2(
        u5_mult_82_SUMB_38__7_), .ZN(u5_mult_82_n3965) );
  NAND2_X1 u5_mult_82_U8978 ( .A1(u5_mult_82_ab_39__6_), .A2(
        u5_mult_82_CARRYB_38__6_), .ZN(u5_mult_82_n3964) );
  NAND2_X1 u5_mult_82_U8977 ( .A1(u5_mult_82_ab_38__7_), .A2(
        u5_mult_82_SUMB_37__8_), .ZN(u5_mult_82_n3962) );
  NAND2_X1 u5_mult_82_U8976 ( .A1(u5_mult_82_CARRYB_37__7_), .A2(
        u5_mult_82_ab_38__7_), .ZN(u5_mult_82_n3961) );
  NAND2_X1 u5_mult_82_U8975 ( .A1(u5_mult_82_n702), .A2(
        u5_mult_82_SUMB_46__22_), .ZN(u5_mult_82_n5747) );
  NAND2_X2 u5_mult_82_U8974 ( .A1(u5_mult_82_SUMB_32__26_), .A2(
        u5_mult_82_n1432), .ZN(u5_mult_82_n3959) );
  NAND2_X2 u5_mult_82_U8973 ( .A1(u5_mult_82_ab_33__25_), .A2(
        u5_mult_82_SUMB_32__26_), .ZN(u5_mult_82_n3958) );
  NAND2_X1 u5_mult_82_U8972 ( .A1(u5_mult_82_ab_33__25_), .A2(
        u5_mult_82_CARRYB_32__25_), .ZN(u5_mult_82_n3957) );
  NAND2_X1 u5_mult_82_U8971 ( .A1(u5_mult_82_ab_32__26_), .A2(
        u5_mult_82_CARRYB_31__26_), .ZN(u5_mult_82_n3954) );
  XOR2_X2 u5_mult_82_U8970 ( .A(u5_mult_82_n3953), .B(u5_mult_82_SUMB_32__26_), 
        .Z(u5_mult_82_SUMB_33__25_) );
  XOR2_X2 u5_mult_82_U8969 ( .A(u5_mult_82_ab_33__25_), .B(
        u5_mult_82_CARRYB_32__25_), .Z(u5_mult_82_n3953) );
  XOR2_X2 u5_mult_82_U8968 ( .A(u5_mult_82_SUMB_6__41_), .B(u5_mult_82_n4019), 
        .Z(u5_mult_82_SUMB_7__40_) );
  NAND3_X2 u5_mult_82_U8967 ( .A1(u5_mult_82_n3950), .A2(u5_mult_82_n3951), 
        .A3(u5_mult_82_n3952), .ZN(u5_mult_82_CARRYB_23__43_) );
  NAND2_X1 u5_mult_82_U8966 ( .A1(u5_mult_82_CARRYB_22__43_), .A2(
        u5_mult_82_SUMB_22__44_), .ZN(u5_mult_82_n3952) );
  NAND2_X1 u5_mult_82_U8965 ( .A1(u5_mult_82_ab_23__43_), .A2(
        u5_mult_82_SUMB_22__44_), .ZN(u5_mult_82_n3951) );
  NAND2_X1 u5_mult_82_U8964 ( .A1(u5_mult_82_CARRYB_22__43_), .A2(
        u5_mult_82_ab_23__43_), .ZN(u5_mult_82_n3950) );
  NAND2_X2 u5_mult_82_U8963 ( .A1(u5_mult_82_CARRYB_21__44_), .A2(
        u5_mult_82_SUMB_21__45_), .ZN(u5_mult_82_n3949) );
  NAND2_X2 u5_mult_82_U8962 ( .A1(u5_mult_82_ab_22__44_), .A2(
        u5_mult_82_SUMB_21__45_), .ZN(u5_mult_82_n3948) );
  XOR2_X2 u5_mult_82_U8961 ( .A(u5_mult_82_n3945), .B(u5_mult_82_SUMB_21__45_), 
        .Z(u5_mult_82_SUMB_22__44_) );
  NAND3_X2 u5_mult_82_U8960 ( .A1(u5_mult_82_n3942), .A2(u5_mult_82_n3943), 
        .A3(u5_mult_82_n3944), .ZN(u5_mult_82_CARRYB_42__31_) );
  NAND2_X1 u5_mult_82_U8959 ( .A1(u5_mult_82_ab_42__31_), .A2(
        u5_mult_82_SUMB_41__32_), .ZN(u5_mult_82_n3943) );
  NAND3_X2 u5_mult_82_U8958 ( .A1(u5_mult_82_n3939), .A2(u5_mult_82_n3940), 
        .A3(u5_mult_82_n3941), .ZN(u5_mult_82_CARRYB_41__32_) );
  NAND2_X2 u5_mult_82_U8957 ( .A1(u5_mult_82_CARRYB_40__32_), .A2(
        u5_mult_82_SUMB_40__33_), .ZN(u5_mult_82_n3941) );
  NAND2_X2 u5_mult_82_U8956 ( .A1(u5_mult_82_ab_41__32_), .A2(
        u5_mult_82_SUMB_40__33_), .ZN(u5_mult_82_n3940) );
  NAND2_X1 u5_mult_82_U8955 ( .A1(u5_mult_82_ab_41__32_), .A2(
        u5_mult_82_CARRYB_40__32_), .ZN(u5_mult_82_n3939) );
  XOR2_X2 u5_mult_82_U8954 ( .A(u5_mult_82_n3938), .B(u5_mult_82_n1431), .Z(
        u5_mult_82_SUMB_41__32_) );
  XOR2_X2 u5_mult_82_U8953 ( .A(u5_mult_82_ab_41__32_), .B(
        u5_mult_82_CARRYB_40__32_), .Z(u5_mult_82_n3938) );
  NAND2_X1 u5_mult_82_U8952 ( .A1(u5_mult_82_ab_39__34_), .A2(
        u5_mult_82_CARRYB_38__34_), .ZN(u5_mult_82_n3935) );
  NAND2_X2 u5_mult_82_U8951 ( .A1(u5_mult_82_ab_38__35_), .A2(
        u5_mult_82_SUMB_37__36_), .ZN(u5_mult_82_n3933) );
  NAND2_X1 u5_mult_82_U8950 ( .A1(u5_mult_82_ab_38__35_), .A2(
        u5_mult_82_CARRYB_37__35_), .ZN(u5_mult_82_n3932) );
  NAND3_X2 u5_mult_82_U8949 ( .A1(u5_mult_82_n4810), .A2(u5_mult_82_n4809), 
        .A3(u5_mult_82_n4808), .ZN(u5_mult_82_CARRYB_23__32_) );
  NAND2_X1 u5_mult_82_U8948 ( .A1(u5_mult_82_ab_10__38_), .A2(
        u5_mult_82_SUMB_9__39_), .ZN(u5_mult_82_n4011) );
  XNOR2_X2 u5_mult_82_U8947 ( .A(u5_mult_82_CARRYB_38__36_), .B(
        u5_mult_82_n3931), .ZN(u5_mult_82_n4471) );
  NOR2_X1 u5_mult_82_U8946 ( .A1(u5_mult_82_n6856), .A2(u5_mult_82_net65369), 
        .ZN(u5_mult_82_ab_42__30_) );
  NAND2_X1 u5_mult_82_U8945 ( .A1(u5_mult_82_ab_36__34_), .A2(
        u5_mult_82_CARRYB_35__34_), .ZN(u5_mult_82_n3928) );
  NAND3_X4 u5_mult_82_U8944 ( .A1(u5_mult_82_n3925), .A2(u5_mult_82_n3926), 
        .A3(u5_mult_82_n3927), .ZN(u5_mult_82_CARRYB_35__35_) );
  NAND2_X2 u5_mult_82_U8943 ( .A1(u5_mult_82_n1631), .A2(
        u5_mult_82_SUMB_34__36_), .ZN(u5_mult_82_n3927) );
  NAND2_X2 u5_mult_82_U8942 ( .A1(u5_mult_82_ab_35__35_), .A2(
        u5_mult_82_SUMB_34__36_), .ZN(u5_mult_82_n3926) );
  NAND2_X1 u5_mult_82_U8941 ( .A1(u5_mult_82_ab_35__35_), .A2(
        u5_mult_82_CARRYB_34__35_), .ZN(u5_mult_82_n3925) );
  XOR2_X2 u5_mult_82_U8940 ( .A(u5_mult_82_n3923), .B(u5_mult_82_n3), .Z(
        u5_mult_82_SUMB_35__35_) );
  XOR2_X2 u5_mult_82_U8939 ( .A(u5_mult_82_ab_35__35_), .B(
        u5_mult_82_CARRYB_34__35_), .Z(u5_mult_82_n3923) );
  NAND3_X2 u5_mult_82_U8938 ( .A1(u5_mult_82_n3920), .A2(u5_mult_82_n3921), 
        .A3(u5_mult_82_n3922), .ZN(u5_mult_82_CARRYB_42__30_) );
  NAND2_X1 u5_mult_82_U8937 ( .A1(u5_mult_82_ab_42__30_), .A2(
        u5_mult_82_CARRYB_41__30_), .ZN(u5_mult_82_n3922) );
  NAND2_X2 u5_mult_82_U8936 ( .A1(u5_mult_82_ab_42__30_), .A2(
        u5_mult_82_SUMB_41__31_), .ZN(u5_mult_82_n3921) );
  NAND2_X1 u5_mult_82_U8935 ( .A1(u5_mult_82_CARRYB_41__30_), .A2(
        u5_mult_82_SUMB_41__31_), .ZN(u5_mult_82_n3920) );
  XOR2_X2 u5_mult_82_U8934 ( .A(u5_mult_82_SUMB_41__31_), .B(u5_mult_82_n3919), 
        .Z(u5_mult_82_SUMB_42__30_) );
  XOR2_X2 u5_mult_82_U8933 ( .A(u5_mult_82_CARRYB_41__30_), .B(
        u5_mult_82_ab_42__30_), .Z(u5_mult_82_n3919) );
  NAND3_X2 u5_mult_82_U8932 ( .A1(u5_mult_82_n4863), .A2(u5_mult_82_n4862), 
        .A3(u5_mult_82_n4864), .ZN(u5_mult_82_CARRYB_16__32_) );
  NOR2_X1 u5_mult_82_U8931 ( .A1(u5_mult_82_net64683), .A2(u5_mult_82_n6735), 
        .ZN(u5_mult_82_ab_44__23_) );
  NAND3_X2 u5_mult_82_U8930 ( .A1(u5_mult_82_n3916), .A2(u5_mult_82_n3917), 
        .A3(u5_mult_82_n3918), .ZN(u5_mult_82_CARRYB_44__23_) );
  NAND2_X1 u5_mult_82_U8929 ( .A1(u5_mult_82_ab_44__23_), .A2(
        u5_mult_82_CARRYB_43__23_), .ZN(u5_mult_82_n3918) );
  NAND2_X2 u5_mult_82_U8928 ( .A1(u5_mult_82_ab_44__23_), .A2(
        u5_mult_82_SUMB_43__24_), .ZN(u5_mult_82_n3917) );
  NAND2_X1 u5_mult_82_U8927 ( .A1(u5_mult_82_CARRYB_43__23_), .A2(
        u5_mult_82_SUMB_43__24_), .ZN(u5_mult_82_n3916) );
  NAND2_X2 u5_mult_82_U8926 ( .A1(u5_mult_82_n1425), .A2(
        u5_mult_82_SUMB_41__25_), .ZN(u5_mult_82_n3914) );
  NAND2_X2 u5_mult_82_U8925 ( .A1(u5_mult_82_ab_42__24_), .A2(
        u5_mult_82_SUMB_41__25_), .ZN(u5_mult_82_n3913) );
  NAND2_X1 u5_mult_82_U8924 ( .A1(u5_mult_82_ab_42__24_), .A2(
        u5_mult_82_CARRYB_41__24_), .ZN(u5_mult_82_n3912) );
  NAND3_X2 u5_mult_82_U8923 ( .A1(u5_mult_82_n3911), .A2(u5_mult_82_n3910), 
        .A3(u5_mult_82_n3909), .ZN(u5_mult_82_CARRYB_41__25_) );
  NAND2_X2 u5_mult_82_U8922 ( .A1(u5_mult_82_CARRYB_40__25_), .A2(
        u5_mult_82_SUMB_40__26_), .ZN(u5_mult_82_n3911) );
  NAND2_X2 u5_mult_82_U8921 ( .A1(u5_mult_82_ab_41__25_), .A2(
        u5_mult_82_SUMB_40__26_), .ZN(u5_mult_82_n3910) );
  NAND2_X1 u5_mult_82_U8920 ( .A1(u5_mult_82_ab_41__25_), .A2(
        u5_mult_82_CARRYB_40__25_), .ZN(u5_mult_82_n3909) );
  XOR2_X2 u5_mult_82_U8919 ( .A(u5_mult_82_n3908), .B(u5_mult_82_n1844), .Z(
        u5_mult_82_SUMB_41__25_) );
  XOR2_X2 u5_mult_82_U8918 ( .A(u5_mult_82_ab_41__25_), .B(
        u5_mult_82_CARRYB_40__25_), .Z(u5_mult_82_n3908) );
  XNOR2_X2 u5_mult_82_U8917 ( .A(u5_mult_82_CARRYB_43__20_), .B(
        u5_mult_82_ab_44__20_), .ZN(u5_mult_82_n3907) );
  XNOR2_X2 u5_mult_82_U8916 ( .A(u5_mult_82_SUMB_43__21_), .B(u5_mult_82_n3907), .ZN(u5_mult_82_SUMB_44__20_) );
  NOR2_X1 u5_mult_82_U8915 ( .A1(u5_mult_82_net64453), .A2(u5_mult_82_n6658), 
        .ZN(u5_mult_82_ab_27__10_) );
  NOR2_X1 u5_mult_82_U8914 ( .A1(u5_mult_82_net64453), .A2(u5_mult_82_n6651), 
        .ZN(u5_mult_82_ab_26__10_) );
  NAND2_X2 u5_mult_82_U8913 ( .A1(u5_mult_82_ab_12__25_), .A2(
        u5_mult_82_CARRYB_11__25_), .ZN(u5_mult_82_n4488) );
  NOR2_X2 u5_mult_82_U8912 ( .A1(u5_mult_82_n6887), .A2(u5_mult_82_n6558), 
        .ZN(u5_mult_82_ab_11__25_) );
  NAND3_X2 u5_mult_82_U8911 ( .A1(u5_mult_82_n3904), .A2(u5_mult_82_n3905), 
        .A3(u5_mult_82_n3906), .ZN(u5_mult_82_CARRYB_27__10_) );
  NAND2_X1 u5_mult_82_U8910 ( .A1(u5_mult_82_ab_27__10_), .A2(
        u5_mult_82_CARRYB_26__10_), .ZN(u5_mult_82_n3906) );
  NAND2_X1 u5_mult_82_U8909 ( .A1(u5_mult_82_CARRYB_26__10_), .A2(
        u5_mult_82_SUMB_26__11_), .ZN(u5_mult_82_n3904) );
  NAND3_X2 u5_mult_82_U8908 ( .A1(u5_mult_82_n3901), .A2(u5_mult_82_n3902), 
        .A3(u5_mult_82_n3903), .ZN(u5_mult_82_CARRYB_26__10_) );
  NAND2_X1 u5_mult_82_U8907 ( .A1(u5_mult_82_ab_26__10_), .A2(
        u5_mult_82_CARRYB_25__10_), .ZN(u5_mult_82_n3903) );
  NAND2_X2 u5_mult_82_U8906 ( .A1(u5_mult_82_ab_26__10_), .A2(
        u5_mult_82_SUMB_25__11_), .ZN(u5_mult_82_n3902) );
  NAND2_X1 u5_mult_82_U8905 ( .A1(u5_mult_82_SUMB_25__11_), .A2(
        u5_mult_82_CARRYB_25__10_), .ZN(u5_mult_82_n3901) );
  NAND3_X4 u5_mult_82_U8904 ( .A1(u5_mult_82_n3898), .A2(u5_mult_82_n3899), 
        .A3(u5_mult_82_n3900), .ZN(u5_mult_82_CARRYB_11__25_) );
  NAND2_X2 u5_mult_82_U8903 ( .A1(u5_mult_82_ab_11__25_), .A2(
        u5_mult_82_SUMB_10__26_), .ZN(u5_mult_82_n3899) );
  NAND3_X2 u5_mult_82_U8902 ( .A1(u5_mult_82_n3895), .A2(u5_mult_82_n3896), 
        .A3(u5_mult_82_n3897), .ZN(u5_mult_82_CARRYB_17__19_) );
  NAND2_X1 u5_mult_82_U8901 ( .A1(u5_mult_82_CARRYB_16__19_), .A2(
        u5_mult_82_SUMB_16__20_), .ZN(u5_mult_82_n3897) );
  NAND2_X1 u5_mult_82_U8900 ( .A1(u5_mult_82_ab_17__19_), .A2(
        u5_mult_82_SUMB_16__20_), .ZN(u5_mult_82_n3896) );
  NAND2_X1 u5_mult_82_U8899 ( .A1(u5_mult_82_ab_17__19_), .A2(
        u5_mult_82_CARRYB_16__19_), .ZN(u5_mult_82_n3895) );
  NAND2_X1 u5_mult_82_U8898 ( .A1(u5_mult_82_ab_16__20_), .A2(
        u5_mult_82_SUMB_15__21_), .ZN(u5_mult_82_n3893) );
  NAND2_X1 u5_mult_82_U8897 ( .A1(u5_mult_82_ab_16__20_), .A2(
        u5_mult_82_CARRYB_15__20_), .ZN(u5_mult_82_n3892) );
  NAND3_X2 u5_mult_82_U8896 ( .A1(u5_mult_82_n3888), .A2(u5_mult_82_n3889), 
        .A3(u5_mult_82_n3890), .ZN(u5_mult_82_CARRYB_14__22_) );
  NAND2_X1 u5_mult_82_U8895 ( .A1(u5_mult_82_CARRYB_13__22_), .A2(
        u5_mult_82_SUMB_13__23_), .ZN(u5_mult_82_n3890) );
  NAND2_X1 u5_mult_82_U8894 ( .A1(u5_mult_82_ab_14__22_), .A2(
        u5_mult_82_SUMB_13__23_), .ZN(u5_mult_82_n3889) );
  NAND2_X1 u5_mult_82_U8893 ( .A1(u5_mult_82_ab_14__22_), .A2(
        u5_mult_82_CARRYB_13__22_), .ZN(u5_mult_82_n3888) );
  NAND3_X2 u5_mult_82_U8892 ( .A1(u5_mult_82_n3885), .A2(u5_mult_82_n3886), 
        .A3(u5_mult_82_n3887), .ZN(u5_mult_82_CARRYB_13__23_) );
  NAND2_X2 u5_mult_82_U8891 ( .A1(u5_mult_82_ab_13__23_), .A2(
        u5_mult_82_SUMB_12__24_), .ZN(u5_mult_82_n3886) );
  XOR2_X2 u5_mult_82_U8890 ( .A(u5_mult_82_n3884), .B(u5_mult_82_SUMB_12__24_), 
        .Z(u5_mult_82_SUMB_13__23_) );
  NAND2_X1 u5_mult_82_U8889 ( .A1(u5_mult_82_ab_38__15_), .A2(
        u5_mult_82_CARRYB_37__15_), .ZN(u5_mult_82_n3880) );
  XNOR2_X2 u5_mult_82_U8888 ( .A(u5_mult_82_ab_27__34_), .B(
        u5_mult_82_CARRYB_26__34_), .ZN(u5_mult_82_n3879) );
  XNOR2_X2 u5_mult_82_U8887 ( .A(u5_mult_82_n3879), .B(u5_mult_82_SUMB_26__35_), .ZN(u5_mult_82_SUMB_27__34_) );
  NOR2_X1 u5_mult_82_U8886 ( .A1(u5_mult_82_n6891), .A2(u5_mult_82_net65353), 
        .ZN(u5_mult_82_ab_43__24_) );
  NAND3_X2 u5_mult_82_U8885 ( .A1(u5_mult_82_n3876), .A2(u5_mult_82_n3877), 
        .A3(u5_mult_82_n3878), .ZN(u5_mult_82_CARRYB_43__24_) );
  NAND2_X1 u5_mult_82_U8884 ( .A1(u5_mult_82_ab_43__24_), .A2(
        u5_mult_82_CARRYB_42__24_), .ZN(u5_mult_82_n3878) );
  NAND2_X2 u5_mult_82_U8883 ( .A1(u5_mult_82_ab_43__24_), .A2(
        u5_mult_82_SUMB_42__25_), .ZN(u5_mult_82_n3877) );
  XOR2_X2 u5_mult_82_U8882 ( .A(u5_mult_82_SUMB_42__25_), .B(u5_mult_82_n3875), 
        .Z(u5_mult_82_SUMB_43__24_) );
  XOR2_X2 u5_mult_82_U8881 ( .A(u5_mult_82_CARRYB_42__24_), .B(
        u5_mult_82_ab_43__24_), .Z(u5_mult_82_n3875) );
  NOR2_X1 u5_mult_82_U8880 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6628), 
        .ZN(u5_mult_82_ab_21__36_) );
  NOR2_X1 u5_mult_82_U8879 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6621), 
        .ZN(u5_mult_82_ab_20__36_) );
  NAND2_X2 u5_mult_82_U8878 ( .A1(u5_mult_82_ab_34__29_), .A2(
        u5_mult_82_CARRYB_33__29_), .ZN(u5_mult_82_n4547) );
  NAND2_X1 u5_mult_82_U8877 ( .A1(u5_mult_82_CARRYB_33__29_), .A2(
        u5_mult_82_SUMB_33__30_), .ZN(u5_mult_82_n4549) );
  NAND2_X4 u5_mult_82_U8876 ( .A1(u5_mult_82_n5563), .A2(u5_mult_82_n5564), 
        .ZN(u5_mult_82_SUMB_32__30_) );
  NOR2_X1 u5_mult_82_U8875 ( .A1(u5_mult_82_n6862), .A2(u5_mult_82_n6699), 
        .ZN(u5_mult_82_ab_33__29_) );
  NAND3_X2 u5_mult_82_U8874 ( .A1(u5_mult_82_n3872), .A2(u5_mult_82_n3873), 
        .A3(u5_mult_82_n3874), .ZN(u5_mult_82_CARRYB_21__36_) );
  NAND2_X1 u5_mult_82_U8873 ( .A1(u5_mult_82_ab_21__36_), .A2(
        u5_mult_82_CARRYB_20__36_), .ZN(u5_mult_82_n3874) );
  NAND2_X1 u5_mult_82_U8872 ( .A1(u5_mult_82_CARRYB_20__36_), .A2(
        u5_mult_82_SUMB_20__37_), .ZN(u5_mult_82_n3872) );
  XOR2_X2 u5_mult_82_U8871 ( .A(u5_mult_82_SUMB_20__37_), .B(u5_mult_82_n3871), 
        .Z(u5_mult_82_SUMB_21__36_) );
  XOR2_X2 u5_mult_82_U8870 ( .A(u5_mult_82_CARRYB_20__36_), .B(
        u5_mult_82_ab_21__36_), .Z(u5_mult_82_n3871) );
  NAND3_X2 u5_mult_82_U8869 ( .A1(u5_mult_82_n3868), .A2(u5_mult_82_n3869), 
        .A3(u5_mult_82_n3870), .ZN(u5_mult_82_CARRYB_20__36_) );
  NAND2_X1 u5_mult_82_U8868 ( .A1(u5_mult_82_ab_20__36_), .A2(
        u5_mult_82_CARRYB_19__36_), .ZN(u5_mult_82_n3870) );
  NAND2_X2 u5_mult_82_U8867 ( .A1(u5_mult_82_ab_20__36_), .A2(
        u5_mult_82_SUMB_19__37_), .ZN(u5_mult_82_n3869) );
  NAND2_X1 u5_mult_82_U8866 ( .A1(u5_mult_82_CARRYB_19__36_), .A2(
        u5_mult_82_SUMB_19__37_), .ZN(u5_mult_82_n3868) );
  XOR2_X2 u5_mult_82_U8865 ( .A(u5_mult_82_SUMB_19__37_), .B(u5_mult_82_n3867), 
        .Z(u5_mult_82_SUMB_20__36_) );
  XOR2_X2 u5_mult_82_U8864 ( .A(u5_mult_82_CARRYB_19__36_), .B(
        u5_mult_82_ab_20__36_), .Z(u5_mult_82_n3867) );
  NAND3_X2 u5_mult_82_U8863 ( .A1(u5_mult_82_n3864), .A2(u5_mult_82_n3865), 
        .A3(u5_mult_82_n3866), .ZN(u5_mult_82_CARRYB_33__29_) );
  NAND2_X1 u5_mult_82_U8862 ( .A1(u5_mult_82_ab_33__29_), .A2(
        u5_mult_82_SUMB_32__30_), .ZN(u5_mult_82_n3866) );
  NAND2_X2 u5_mult_82_U8861 ( .A1(u5_mult_82_CARRYB_32__29_), .A2(
        u5_mult_82_ab_33__29_), .ZN(u5_mult_82_n3865) );
  NAND2_X2 u5_mult_82_U8860 ( .A1(u5_mult_82_SUMB_32__30_), .A2(
        u5_mult_82_CARRYB_32__29_), .ZN(u5_mult_82_n3864) );
  XOR2_X2 u5_mult_82_U8859 ( .A(u5_mult_82_CARRYB_32__29_), .B(
        u5_mult_82_n3863), .Z(u5_mult_82_SUMB_33__29_) );
  XOR2_X2 u5_mult_82_U8858 ( .A(u5_mult_82_SUMB_32__30_), .B(
        u5_mult_82_ab_33__29_), .Z(u5_mult_82_n3863) );
  NOR2_X1 u5_mult_82_U8857 ( .A1(u5_mult_82_n6885), .A2(u5_mult_82_n6728), 
        .ZN(u5_mult_82_ab_39__25_) );
  NAND2_X1 u5_mult_82_U8856 ( .A1(u5_mult_82_ab_41__23_), .A2(
        u5_mult_82_SUMB_40__24_), .ZN(u5_mult_82_n3861) );
  NAND2_X1 u5_mult_82_U8855 ( .A1(u5_mult_82_ab_41__23_), .A2(
        u5_mult_82_CARRYB_40__23_), .ZN(u5_mult_82_n3860) );
  NAND3_X2 u5_mult_82_U8854 ( .A1(u5_mult_82_n3858), .A2(u5_mult_82_n3857), 
        .A3(u5_mult_82_n3859), .ZN(u5_mult_82_CARRYB_40__24_) );
  NAND2_X1 u5_mult_82_U8853 ( .A1(u5_mult_82_ab_40__24_), .A2(
        u5_mult_82_SUMB_39__25_), .ZN(u5_mult_82_n3858) );
  NAND2_X1 u5_mult_82_U8852 ( .A1(u5_mult_82_ab_40__24_), .A2(
        u5_mult_82_CARRYB_39__24_), .ZN(u5_mult_82_n3857) );
  XOR2_X2 u5_mult_82_U8851 ( .A(u5_mult_82_n3855), .B(u5_mult_82_SUMB_39__25_), 
        .Z(u5_mult_82_SUMB_40__24_) );
  XOR2_X2 u5_mult_82_U8850 ( .A(u5_mult_82_ab_40__24_), .B(
        u5_mult_82_CARRYB_39__24_), .Z(u5_mult_82_n3855) );
  NAND3_X2 u5_mult_82_U8849 ( .A1(u5_mult_82_n3852), .A2(u5_mult_82_n3853), 
        .A3(u5_mult_82_n3854), .ZN(u5_mult_82_CARRYB_39__25_) );
  NAND2_X1 u5_mult_82_U8848 ( .A1(u5_mult_82_ab_39__25_), .A2(
        u5_mult_82_CARRYB_38__25_), .ZN(u5_mult_82_n3854) );
  NAND2_X1 u5_mult_82_U8847 ( .A1(u5_mult_82_CARRYB_38__25_), .A2(
        u5_mult_82_SUMB_38__26_), .ZN(u5_mult_82_n3852) );
  XOR2_X2 u5_mult_82_U8846 ( .A(u5_mult_82_n1632), .B(u5_mult_82_n3851), .Z(
        u5_mult_82_SUMB_39__25_) );
  NAND3_X4 u5_mult_82_U8845 ( .A1(u5_mult_82_n3848), .A2(u5_mult_82_n3850), 
        .A3(u5_mult_82_n3849), .ZN(u5_mult_82_CARRYB_46__19_) );
  NAND3_X2 u5_mult_82_U8844 ( .A1(u5_mult_82_n3845), .A2(u5_mult_82_n3846), 
        .A3(u5_mult_82_n3847), .ZN(u5_mult_82_CARRYB_45__20_) );
  NAND2_X2 u5_mult_82_U8843 ( .A1(u5_mult_82_ab_45__20_), .A2(
        u5_mult_82_SUMB_44__21_), .ZN(u5_mult_82_n3846) );
  NAND2_X1 u5_mult_82_U8842 ( .A1(u5_mult_82_ab_45__20_), .A2(
        u5_mult_82_CARRYB_44__20_), .ZN(u5_mult_82_n3845) );
  XNOR2_X2 u5_mult_82_U8841 ( .A(u5_mult_82_CARRYB_32__42_), .B(
        u5_mult_82_ab_33__42_), .ZN(u5_mult_82_n3843) );
  XNOR2_X2 u5_mult_82_U8840 ( .A(u5_mult_82_n3843), .B(u5_mult_82_SUMB_32__43_), .ZN(u5_mult_82_SUMB_33__42_) );
  NAND3_X2 u5_mult_82_U8839 ( .A1(u5_mult_82_n3840), .A2(u5_mult_82_n3841), 
        .A3(u5_mult_82_n3842), .ZN(u5_mult_82_CARRYB_33__39_) );
  NAND2_X2 u5_mult_82_U8838 ( .A1(u5_mult_82_CARRYB_32__39_), .A2(
        u5_mult_82_SUMB_32__40_), .ZN(u5_mult_82_n3842) );
  NAND2_X2 u5_mult_82_U8837 ( .A1(u5_mult_82_ab_33__39_), .A2(
        u5_mult_82_SUMB_32__40_), .ZN(u5_mult_82_n3841) );
  NAND3_X2 u5_mult_82_U8836 ( .A1(u5_mult_82_n3839), .A2(u5_mult_82_n3838), 
        .A3(u5_mult_82_n3837), .ZN(u5_mult_82_CARRYB_32__40_) );
  XOR2_X2 u5_mult_82_U8835 ( .A(u5_mult_82_n3836), .B(u5_mult_82_SUMB_32__40_), 
        .Z(u5_mult_82_SUMB_33__39_) );
  XOR2_X2 u5_mult_82_U8834 ( .A(u5_mult_82_ab_33__39_), .B(
        u5_mult_82_CARRYB_32__39_), .Z(u5_mult_82_n3836) );
  NAND3_X2 u5_mult_82_U8833 ( .A1(u5_mult_82_n3833), .A2(u5_mult_82_n3834), 
        .A3(u5_mult_82_n3835), .ZN(u5_mult_82_CARRYB_46__31_) );
  NAND2_X1 u5_mult_82_U8832 ( .A1(u5_mult_82_ab_46__31_), .A2(
        u5_mult_82_SUMB_45__32_), .ZN(u5_mult_82_n3834) );
  NAND3_X4 u5_mult_82_U8831 ( .A1(u5_mult_82_n3830), .A2(u5_mult_82_n3831), 
        .A3(u5_mult_82_n3832), .ZN(u5_mult_82_CARRYB_45__32_) );
  NAND2_X2 u5_mult_82_U8830 ( .A1(u5_mult_82_CARRYB_44__32_), .A2(
        u5_mult_82_SUMB_44__33_), .ZN(u5_mult_82_n3832) );
  NAND2_X2 u5_mult_82_U8829 ( .A1(u5_mult_82_ab_45__32_), .A2(
        u5_mult_82_SUMB_44__33_), .ZN(u5_mult_82_n3831) );
  NAND2_X1 u5_mult_82_U8828 ( .A1(u5_mult_82_ab_45__32_), .A2(
        u5_mult_82_CARRYB_44__32_), .ZN(u5_mult_82_n3830) );
  XOR2_X2 u5_mult_82_U8827 ( .A(u5_mult_82_n3829), .B(u5_mult_82_SUMB_45__32_), 
        .Z(u5_mult_82_SUMB_46__31_) );
  XOR2_X2 u5_mult_82_U8826 ( .A(u5_mult_82_ab_46__31_), .B(
        u5_mult_82_CARRYB_45__31_), .Z(u5_mult_82_n3829) );
  XOR2_X2 u5_mult_82_U8825 ( .A(u5_mult_82_n3828), .B(u5_mult_82_n1577), .Z(
        u5_mult_82_SUMB_45__32_) );
  XOR2_X2 u5_mult_82_U8824 ( .A(u5_mult_82_ab_45__32_), .B(
        u5_mult_82_CARRYB_44__32_), .Z(u5_mult_82_n3828) );
  XNOR2_X2 u5_mult_82_U8823 ( .A(u5_mult_82_ab_40__30_), .B(
        u5_mult_82_CARRYB_39__30_), .ZN(u5_mult_82_n3827) );
  XNOR2_X2 u5_mult_82_U8822 ( .A(u5_mult_82_n3827), .B(u5_mult_82_SUMB_39__31_), .ZN(u5_mult_82_SUMB_40__30_) );
  XNOR2_X2 u5_mult_82_U8821 ( .A(u5_mult_82_ab_42__26_), .B(
        u5_mult_82_CARRYB_41__26_), .ZN(u5_mult_82_n3826) );
  XNOR2_X2 u5_mult_82_U8820 ( .A(u5_mult_82_n3826), .B(u5_mult_82_SUMB_41__27_), .ZN(u5_mult_82_SUMB_42__26_) );
  NAND2_X2 u5_mult_82_U8819 ( .A1(u5_mult_82_ab_28__29_), .A2(
        u5_mult_82_CARRYB_27__29_), .ZN(u5_mult_82_n5479) );
  XNOR2_X2 u5_mult_82_U8818 ( .A(u5_mult_82_CARRYB_38__10_), .B(
        u5_mult_82_ab_39__10_), .ZN(u5_mult_82_n3824) );
  XNOR2_X2 u5_mult_82_U8817 ( .A(u5_mult_82_n1426), .B(u5_mult_82_n3824), .ZN(
        u5_mult_82_SUMB_39__10_) );
  NAND2_X1 u5_mult_82_U8816 ( .A1(u5_mult_82_ab_7__24_), .A2(u5_mult_82_n104), 
        .ZN(u5_mult_82_n3820) );
  NAND3_X4 u5_mult_82_U8815 ( .A1(u5_mult_82_n3817), .A2(u5_mult_82_n3818), 
        .A3(u5_mult_82_n3819), .ZN(u5_mult_82_CARRYB_6__25_) );
  NAND2_X2 u5_mult_82_U8814 ( .A1(u5_mult_82_CARRYB_5__25_), .A2(
        u5_mult_82_n1824), .ZN(u5_mult_82_n3819) );
  NAND2_X2 u5_mult_82_U8813 ( .A1(u5_mult_82_ab_6__25_), .A2(u5_mult_82_n1824), 
        .ZN(u5_mult_82_n3818) );
  NAND2_X1 u5_mult_82_U8812 ( .A1(u5_mult_82_ab_6__25_), .A2(
        u5_mult_82_CARRYB_5__25_), .ZN(u5_mult_82_n3817) );
  XOR2_X2 u5_mult_82_U8811 ( .A(u5_mult_82_n3816), .B(u5_mult_82_n1667), .Z(
        u5_mult_82_SUMB_7__24_) );
  XOR2_X2 u5_mult_82_U8810 ( .A(u5_mult_82_ab_6__25_), .B(
        u5_mult_82_CARRYB_5__25_), .Z(u5_mult_82_n3815) );
  NAND3_X2 u5_mult_82_U8809 ( .A1(u5_mult_82_n3812), .A2(u5_mult_82_n3813), 
        .A3(u5_mult_82_n3814), .ZN(u5_mult_82_CARRYB_3__28_) );
  NAND2_X1 u5_mult_82_U8808 ( .A1(u5_mult_82_CARRYB_2__28_), .A2(
        u5_mult_82_SUMB_2__29_), .ZN(u5_mult_82_n3814) );
  NAND2_X1 u5_mult_82_U8807 ( .A1(u5_mult_82_ab_3__28_), .A2(
        u5_mult_82_SUMB_2__29_), .ZN(u5_mult_82_n3813) );
  NAND3_X2 u5_mult_82_U8806 ( .A1(u5_mult_82_n3809), .A2(u5_mult_82_n3810), 
        .A3(u5_mult_82_n3811), .ZN(u5_mult_82_CARRYB_2__29_) );
  NAND2_X2 u5_mult_82_U8805 ( .A1(u5_mult_82_CARRYB_1__29_), .A2(
        u5_mult_82_SUMB_1__30_), .ZN(u5_mult_82_n3811) );
  NAND2_X2 u5_mult_82_U8804 ( .A1(u5_mult_82_ab_2__29_), .A2(
        u5_mult_82_SUMB_1__30_), .ZN(u5_mult_82_n3810) );
  NAND2_X1 u5_mult_82_U8803 ( .A1(u5_mult_82_ab_2__29_), .A2(
        u5_mult_82_CARRYB_1__29_), .ZN(u5_mult_82_n3809) );
  XOR2_X2 u5_mult_82_U8802 ( .A(u5_mult_82_n3808), .B(u5_mult_82_SUMB_1__30_), 
        .Z(u5_mult_82_SUMB_2__29_) );
  XOR2_X2 u5_mult_82_U8801 ( .A(u5_mult_82_ab_2__29_), .B(
        u5_mult_82_CARRYB_1__29_), .Z(u5_mult_82_n3808) );
  NAND3_X2 u5_mult_82_U8800 ( .A1(u5_mult_82_n3805), .A2(u5_mult_82_n3806), 
        .A3(u5_mult_82_n3807), .ZN(u5_mult_82_CARRYB_17__14_) );
  NAND2_X1 u5_mult_82_U8799 ( .A1(u5_mult_82_CARRYB_16__14_), .A2(
        u5_mult_82_SUMB_16__15_), .ZN(u5_mult_82_n3807) );
  NAND2_X1 u5_mult_82_U8798 ( .A1(u5_mult_82_ab_17__14_), .A2(
        u5_mult_82_SUMB_16__15_), .ZN(u5_mult_82_n3806) );
  NAND2_X1 u5_mult_82_U8797 ( .A1(u5_mult_82_ab_17__14_), .A2(
        u5_mult_82_CARRYB_16__14_), .ZN(u5_mult_82_n3805) );
  NAND3_X4 u5_mult_82_U8796 ( .A1(u5_mult_82_n3802), .A2(u5_mult_82_n3803), 
        .A3(u5_mult_82_n3804), .ZN(u5_mult_82_CARRYB_16__15_) );
  NAND2_X2 u5_mult_82_U8795 ( .A1(u5_mult_82_CARRYB_15__15_), .A2(
        u5_mult_82_SUMB_15__16_), .ZN(u5_mult_82_n3804) );
  NAND2_X2 u5_mult_82_U8794 ( .A1(u5_mult_82_ab_16__15_), .A2(
        u5_mult_82_SUMB_15__16_), .ZN(u5_mult_82_n3803) );
  NAND3_X2 u5_mult_82_U8793 ( .A1(u5_mult_82_n3799), .A2(u5_mult_82_n3800), 
        .A3(u5_mult_82_n3801), .ZN(u5_mult_82_CARRYB_14__17_) );
  NAND2_X1 u5_mult_82_U8792 ( .A1(u5_mult_82_CARRYB_13__17_), .A2(
        u5_mult_82_SUMB_13__18_), .ZN(u5_mult_82_n3801) );
  NAND2_X1 u5_mult_82_U8791 ( .A1(u5_mult_82_ab_14__17_), .A2(
        u5_mult_82_SUMB_13__18_), .ZN(u5_mult_82_n3800) );
  NAND2_X1 u5_mult_82_U8790 ( .A1(u5_mult_82_ab_14__17_), .A2(
        u5_mult_82_CARRYB_13__17_), .ZN(u5_mult_82_n3799) );
  NAND3_X2 u5_mult_82_U8789 ( .A1(u5_mult_82_n3796), .A2(u5_mult_82_n3797), 
        .A3(u5_mult_82_n3798), .ZN(u5_mult_82_CARRYB_13__18_) );
  NAND2_X2 u5_mult_82_U8788 ( .A1(u5_mult_82_CARRYB_12__18_), .A2(
        u5_mult_82_SUMB_12__19_), .ZN(u5_mult_82_n3798) );
  NAND2_X2 u5_mult_82_U8787 ( .A1(u5_mult_82_ab_13__18_), .A2(
        u5_mult_82_SUMB_12__19_), .ZN(u5_mult_82_n3797) );
  NAND2_X1 u5_mult_82_U8786 ( .A1(u5_mult_82_ab_13__18_), .A2(
        u5_mult_82_CARRYB_12__18_), .ZN(u5_mult_82_n3796) );
  XOR2_X2 u5_mult_82_U8785 ( .A(u5_mult_82_n3795), .B(u5_mult_82_SUMB_12__19_), 
        .Z(u5_mult_82_SUMB_13__18_) );
  XOR2_X2 u5_mult_82_U8784 ( .A(u5_mult_82_ab_13__18_), .B(
        u5_mult_82_CARRYB_12__18_), .Z(u5_mult_82_n3795) );
  NAND3_X2 u5_mult_82_U8783 ( .A1(u5_mult_82_n3792), .A2(u5_mult_82_n3793), 
        .A3(u5_mult_82_n3794), .ZN(u5_mult_82_CARRYB_34__6_) );
  NAND2_X1 u5_mult_82_U8782 ( .A1(u5_mult_82_ab_34__6_), .A2(
        u5_mult_82_SUMB_33__7_), .ZN(u5_mult_82_n3794) );
  NAND2_X1 u5_mult_82_U8781 ( .A1(u5_mult_82_CARRYB_33__6_), .A2(
        u5_mult_82_SUMB_33__7_), .ZN(u5_mult_82_n3793) );
  NAND2_X1 u5_mult_82_U8780 ( .A1(u5_mult_82_CARRYB_33__6_), .A2(
        u5_mult_82_ab_34__6_), .ZN(u5_mult_82_n3792) );
  NAND2_X2 u5_mult_82_U8779 ( .A1(u5_mult_82_n3823), .A2(
        u5_mult_82_SUMB_32__8_), .ZN(u5_mult_82_n3791) );
  NAND2_X2 u5_mult_82_U8778 ( .A1(u5_mult_82_ab_33__7_), .A2(
        u5_mult_82_SUMB_32__8_), .ZN(u5_mult_82_n3790) );
  NAND2_X1 u5_mult_82_U8777 ( .A1(u5_mult_82_ab_33__7_), .A2(u5_mult_82_n3823), 
        .ZN(u5_mult_82_n3789) );
  XOR2_X2 u5_mult_82_U8776 ( .A(u5_mult_82_n3788), .B(u5_mult_82_SUMB_32__8_), 
        .Z(u5_mult_82_SUMB_33__7_) );
  XOR2_X2 u5_mult_82_U8775 ( .A(u5_mult_82_ab_38__12_), .B(
        u5_mult_82_CARRYB_37__12_), .Z(u5_mult_82_n5127) );
  XNOR2_X2 u5_mult_82_U8774 ( .A(u5_mult_82_ab_22__34_), .B(
        u5_mult_82_CARRYB_21__34_), .ZN(u5_mult_82_n3787) );
  XNOR2_X2 u5_mult_82_U8773 ( .A(u5_mult_82_n3787), .B(u5_mult_82_SUMB_21__35_), .ZN(u5_mult_82_SUMB_22__34_) );
  INV_X1 u5_mult_82_U8772 ( .A(u5_mult_82_SUMB_34__15_), .ZN(u5_mult_82_n3784)
         );
  NAND2_X2 u5_mult_82_U8771 ( .A1(u5_mult_82_n3783), .A2(u5_mult_82_n3784), 
        .ZN(u5_mult_82_n3786) );
  NOR2_X1 u5_mult_82_U8770 ( .A1(u5_mult_82_n6861), .A2(u5_mult_82_n6742), 
        .ZN(u5_mult_82_ab_46__29_) );
  NAND3_X2 u5_mult_82_U8769 ( .A1(u5_mult_82_n3780), .A2(u5_mult_82_n3781), 
        .A3(u5_mult_82_n3782), .ZN(u5_mult_82_CARRYB_46__29_) );
  NAND2_X1 u5_mult_82_U8768 ( .A1(u5_mult_82_ab_46__29_), .A2(
        u5_mult_82_CARRYB_45__29_), .ZN(u5_mult_82_n3782) );
  NAND2_X2 u5_mult_82_U8767 ( .A1(u5_mult_82_ab_46__29_), .A2(
        u5_mult_82_SUMB_45__30_), .ZN(u5_mult_82_n3781) );
  NAND2_X1 u5_mult_82_U8766 ( .A1(u5_mult_82_SUMB_45__30_), .A2(
        u5_mult_82_CARRYB_45__29_), .ZN(u5_mult_82_n3780) );
  NAND2_X2 u5_mult_82_U8765 ( .A1(u5_mult_82_CARRYB_32__40_), .A2(
        u5_mult_82_SUMB_32__41_), .ZN(u5_mult_82_n3779) );
  NAND2_X2 u5_mult_82_U8764 ( .A1(u5_mult_82_ab_33__40_), .A2(
        u5_mult_82_SUMB_32__41_), .ZN(u5_mult_82_n3778) );
  NAND2_X1 u5_mult_82_U8763 ( .A1(u5_mult_82_ab_33__40_), .A2(
        u5_mult_82_CARRYB_32__40_), .ZN(u5_mult_82_n3777) );
  NAND2_X2 u5_mult_82_U8762 ( .A1(u5_mult_82_CARRYB_31__41_), .A2(
        u5_mult_82_SUMB_31__42_), .ZN(u5_mult_82_n3776) );
  NAND2_X2 u5_mult_82_U8761 ( .A1(u5_mult_82_ab_32__41_), .A2(
        u5_mult_82_SUMB_31__42_), .ZN(u5_mult_82_n3775) );
  NAND2_X1 u5_mult_82_U8760 ( .A1(u5_mult_82_ab_32__41_), .A2(
        u5_mult_82_CARRYB_31__41_), .ZN(u5_mult_82_n3774) );
  XNOR2_X2 u5_mult_82_U8759 ( .A(u5_mult_82_CARRYB_36__9_), .B(
        u5_mult_82_ab_37__9_), .ZN(u5_mult_82_n3773) );
  XNOR2_X2 u5_mult_82_U8758 ( .A(u5_mult_82_SUMB_36__10_), .B(u5_mult_82_n3773), .ZN(u5_mult_82_SUMB_37__9_) );
  NAND3_X2 u5_mult_82_U8757 ( .A1(u5_mult_82_n4429), .A2(u5_mult_82_n4430), 
        .A3(u5_mult_82_n4431), .ZN(u5_mult_82_CARRYB_18__47_) );
  XNOR2_X2 u5_mult_82_U8756 ( .A(u5_mult_82_ab_34__30_), .B(
        u5_mult_82_CARRYB_33__30_), .ZN(u5_mult_82_n3771) );
  NAND2_X1 u5_mult_82_U8755 ( .A1(u5_mult_82_ab_38__22_), .A2(
        u5_mult_82_SUMB_37__23_), .ZN(u5_mult_82_n4805) );
  NAND2_X2 u5_mult_82_U8754 ( .A1(u5_mult_82_ab_25__33_), .A2(
        u5_mult_82_SUMB_24__34_), .ZN(u5_mult_82_n6228) );
  NAND2_X2 u5_mult_82_U8753 ( .A1(u5_mult_82_CARRYB_47__6_), .A2(
        u5_mult_82_SUMB_47__7_), .ZN(u5_mult_82_n4381) );
  NAND3_X4 u5_mult_82_U8752 ( .A1(u5_mult_82_n4381), .A2(u5_mult_82_n4382), 
        .A3(u5_mult_82_n4383), .ZN(u5_mult_82_CARRYB_48__6_) );
  XOR2_X2 u5_mult_82_U8751 ( .A(u5_mult_82_ab_11__51_), .B(
        u5_mult_82_CARRYB_10__51_), .Z(u5_mult_82_n4648) );
  NOR2_X1 u5_mult_82_U8750 ( .A1(u5_mult_82_n6779), .A2(u5_mult_82_n6642), 
        .ZN(u5_mult_82_ab_24__48_) );
  NOR2_X1 u5_mult_82_U8749 ( .A1(u5_mult_82_n6861), .A2(u5_mult_82_n6747), 
        .ZN(u5_mult_82_ab_48__29_) );
  NAND3_X2 u5_mult_82_U8748 ( .A1(u5_mult_82_n3768), .A2(u5_mult_82_n3769), 
        .A3(u5_mult_82_n3770), .ZN(u5_mult_82_CARRYB_24__48_) );
  NAND2_X1 u5_mult_82_U8747 ( .A1(u5_mult_82_ab_24__48_), .A2(
        u5_mult_82_SUMB_23__49_), .ZN(u5_mult_82_n3770) );
  NAND2_X2 u5_mult_82_U8746 ( .A1(u5_mult_82_ab_24__48_), .A2(
        u5_mult_82_CARRYB_23__48_), .ZN(u5_mult_82_n3769) );
  NAND2_X2 u5_mult_82_U8745 ( .A1(u5_mult_82_SUMB_23__49_), .A2(
        u5_mult_82_CARRYB_23__48_), .ZN(u5_mult_82_n3768) );
  XOR2_X2 u5_mult_82_U8744 ( .A(u5_mult_82_SUMB_23__49_), .B(
        u5_mult_82_ab_24__48_), .Z(u5_mult_82_n3767) );
  NAND2_X2 u5_mult_82_U8743 ( .A1(u5_mult_82_CARRYB_33__40_), .A2(
        u5_mult_82_SUMB_33__41_), .ZN(u5_mult_82_n3766) );
  NAND2_X2 u5_mult_82_U8742 ( .A1(u5_mult_82_ab_34__40_), .A2(
        u5_mult_82_SUMB_33__41_), .ZN(u5_mult_82_n3765) );
  NAND2_X1 u5_mult_82_U8741 ( .A1(u5_mult_82_ab_34__40_), .A2(
        u5_mult_82_CARRYB_33__40_), .ZN(u5_mult_82_n3764) );
  NAND3_X4 u5_mult_82_U8740 ( .A1(u5_mult_82_n3761), .A2(u5_mult_82_n3762), 
        .A3(u5_mult_82_n3763), .ZN(u5_mult_82_CARRYB_33__41_) );
  NAND2_X2 u5_mult_82_U8739 ( .A1(u5_mult_82_CARRYB_32__41_), .A2(
        u5_mult_82_SUMB_32__42_), .ZN(u5_mult_82_n3763) );
  NAND2_X2 u5_mult_82_U8738 ( .A1(u5_mult_82_ab_33__41_), .A2(
        u5_mult_82_SUMB_32__42_), .ZN(u5_mult_82_n3762) );
  NAND2_X1 u5_mult_82_U8737 ( .A1(u5_mult_82_ab_33__41_), .A2(
        u5_mult_82_CARRYB_32__41_), .ZN(u5_mult_82_n3761) );
  XOR2_X2 u5_mult_82_U8736 ( .A(u5_mult_82_n3760), .B(u5_mult_82_SUMB_33__41_), 
        .Z(u5_mult_82_SUMB_34__40_) );
  XOR2_X2 u5_mult_82_U8735 ( .A(u5_mult_82_ab_34__40_), .B(
        u5_mult_82_CARRYB_33__40_), .Z(u5_mult_82_n3760) );
  NAND2_X1 u5_mult_82_U8734 ( .A1(u5_mult_82_ab_48__29_), .A2(
        u5_mult_82_CARRYB_47__29_), .ZN(u5_mult_82_n3759) );
  NAND3_X2 u5_mult_82_U8733 ( .A1(u5_mult_82_n3754), .A2(u5_mult_82_n3755), 
        .A3(u5_mult_82_n3756), .ZN(u5_mult_82_CARRYB_51__26_) );
  NAND2_X1 u5_mult_82_U8732 ( .A1(u5_mult_82_CARRYB_50__26_), .A2(
        u5_mult_82_SUMB_50__27_), .ZN(u5_mult_82_n3756) );
  NAND2_X1 u5_mult_82_U8731 ( .A1(u5_mult_82_ab_51__26_), .A2(
        u5_mult_82_SUMB_50__27_), .ZN(u5_mult_82_n3755) );
  NAND2_X1 u5_mult_82_U8730 ( .A1(u5_mult_82_ab_51__26_), .A2(
        u5_mult_82_CARRYB_50__26_), .ZN(u5_mult_82_n3754) );
  NAND3_X2 u5_mult_82_U8729 ( .A1(u5_mult_82_n3751), .A2(u5_mult_82_n3752), 
        .A3(u5_mult_82_n3753), .ZN(u5_mult_82_CARRYB_50__27_) );
  NAND2_X2 u5_mult_82_U8728 ( .A1(u5_mult_82_ab_50__27_), .A2(
        u5_mult_82_SUMB_49__28_), .ZN(u5_mult_82_n3752) );
  NAND3_X4 u5_mult_82_U8727 ( .A1(u5_mult_82_n5509), .A2(u5_mult_82_n5510), 
        .A3(u5_mult_82_n5511), .ZN(u5_mult_82_CARRYB_24__32_) );
  NAND2_X2 u5_mult_82_U8726 ( .A1(u5_mult_82_ab_46__4_), .A2(
        u5_mult_82_CARRYB_45__4_), .ZN(u5_mult_82_n4598) );
  XNOR2_X2 u5_mult_82_U8725 ( .A(u5_mult_82_ab_24__17_), .B(
        u5_mult_82_CARRYB_23__17_), .ZN(u5_mult_82_n3750) );
  XNOR2_X2 u5_mult_82_U8724 ( .A(u5_mult_82_n3750), .B(u5_mult_82_SUMB_23__18_), .ZN(u5_mult_82_SUMB_24__17_) );
  XNOR2_X2 u5_mult_82_U8723 ( .A(u5_mult_82_n3749), .B(u5_mult_82_SUMB_44__6_), 
        .ZN(u5_mult_82_SUMB_45__5_) );
  NAND2_X2 u5_mult_82_U8722 ( .A1(u5_mult_82_ab_23__31_), .A2(
        u5_mult_82_SUMB_22__32_), .ZN(u5_mult_82_n6343) );
  XNOR2_X2 u5_mult_82_U8721 ( .A(u5_mult_82_n446), .B(u5_mult_82_ab_21__39_), 
        .ZN(u5_mult_82_n3748) );
  XNOR2_X2 u5_mult_82_U8720 ( .A(u5_mult_82_n3748), .B(u5_mult_82_SUMB_20__40_), .ZN(u5_mult_82_SUMB_21__39_) );
  XOR2_X2 u5_mult_82_U8719 ( .A(u5_mult_82_SUMB_42__6_), .B(u5_mult_82_n4802), 
        .Z(u5_mult_82_n3747) );
  XNOR2_X2 u5_mult_82_U8718 ( .A(u5_mult_82_n1835), .B(u5_mult_82_n3747), .ZN(
        u5_mult_82_SUMB_43__5_) );
  NAND2_X2 u5_mult_82_U8717 ( .A1(u5_mult_82_ab_49__5_), .A2(
        u5_mult_82_SUMB_48__6_), .ZN(u5_mult_82_n6326) );
  NAND2_X1 u5_mult_82_U8716 ( .A1(u5_mult_82_CARRYB_4__50_), .A2(
        u5_mult_82_ab_5__50_), .ZN(u5_mult_82_n6293) );
  NAND2_X2 u5_mult_82_U8715 ( .A1(u5_mult_82_SUMB_42__7_), .A2(
        u5_mult_82_CARRYB_42__6_), .ZN(u5_mult_82_n6032) );
  NAND2_X2 u5_mult_82_U8714 ( .A1(u5_mult_82_ab_42__6_), .A2(
        u5_mult_82_SUMB_41__7_), .ZN(u5_mult_82_n6007) );
  XNOR2_X2 u5_mult_82_U8713 ( .A(u5_mult_82_n3746), .B(
        u5_mult_82_CARRYB_24__34_), .ZN(u5_mult_82_n5762) );
  NAND2_X2 u5_mult_82_U8712 ( .A1(u5_mult_82_n1721), .A2(
        u5_mult_82_SUMB_44__4_), .ZN(u5_mult_82_n5793) );
  XNOR2_X2 u5_mult_82_U8711 ( .A(u5_mult_82_n3745), .B(u5_mult_82_SUMB_20__34_), .ZN(u5_mult_82_n4817) );
  NAND2_X2 u5_mult_82_U8710 ( .A1(u5_mult_82_ab_45__3_), .A2(
        u5_mult_82_SUMB_44__4_), .ZN(u5_mult_82_n5792) );
  NAND3_X2 u5_mult_82_U8709 ( .A1(u5_mult_82_n3741), .A2(u5_mult_82_n3742), 
        .A3(u5_mult_82_n3743), .ZN(u5_mult_82_CARRYB_34__7_) );
  NAND2_X1 u5_mult_82_U8708 ( .A1(u5_mult_82_ab_34__7_), .A2(
        u5_mult_82_SUMB_33__8_), .ZN(u5_mult_82_n3743) );
  NAND2_X1 u5_mult_82_U8707 ( .A1(u5_mult_82_CARRYB_33__7_), .A2(
        u5_mult_82_SUMB_33__8_), .ZN(u5_mult_82_n3742) );
  NAND2_X1 u5_mult_82_U8706 ( .A1(u5_mult_82_CARRYB_33__7_), .A2(
        u5_mult_82_ab_34__7_), .ZN(u5_mult_82_n3741) );
  NAND2_X2 u5_mult_82_U8705 ( .A1(u5_mult_82_ab_29__10_), .A2(
        u5_mult_82_SUMB_28__11_), .ZN(u5_mult_82_n3736) );
  NAND2_X1 u5_mult_82_U8704 ( .A1(u5_mult_82_ab_29__10_), .A2(
        u5_mult_82_CARRYB_28__10_), .ZN(u5_mult_82_n3735) );
  NAND3_X4 u5_mult_82_U8703 ( .A1(u5_mult_82_n3732), .A2(u5_mult_82_n3733), 
        .A3(u5_mult_82_n3734), .ZN(u5_mult_82_CARRYB_28__11_) );
  NAND2_X2 u5_mult_82_U8702 ( .A1(u5_mult_82_CARRYB_27__11_), .A2(
        u5_mult_82_SUMB_27__12_), .ZN(u5_mult_82_n3734) );
  NAND2_X2 u5_mult_82_U8701 ( .A1(u5_mult_82_ab_28__11_), .A2(
        u5_mult_82_SUMB_27__12_), .ZN(u5_mult_82_n3733) );
  NAND2_X2 u5_mult_82_U8700 ( .A1(u5_mult_82_ab_28__11_), .A2(
        u5_mult_82_CARRYB_27__11_), .ZN(u5_mult_82_n3732) );
  XNOR2_X2 u5_mult_82_U8699 ( .A(u5_mult_82_net82990), .B(
        u5_mult_82_SUMB_26__22_), .ZN(u5_mult_82_SUMB_27__21_) );
  XNOR2_X2 u5_mult_82_U8698 ( .A(u5_mult_82_ab_45__6_), .B(
        u5_mult_82_CARRYB_44__6_), .ZN(u5_mult_82_n3731) );
  XNOR2_X2 u5_mult_82_U8697 ( .A(u5_mult_82_n3731), .B(u5_mult_82_n1610), .ZN(
        u5_mult_82_SUMB_45__6_) );
  NOR2_X1 u5_mult_82_U8696 ( .A1(u5_mult_82_net64435), .A2(u5_mult_82_n6637), 
        .ZN(u5_mult_82_ab_22__9_) );
  NOR2_X1 u5_mult_82_U8695 ( .A1(u5_mult_82_net64435), .A2(u5_mult_82_n6630), 
        .ZN(u5_mult_82_ab_21__9_) );
  NOR2_X1 u5_mult_82_U8694 ( .A1(u5_mult_82_net64671), .A2(u5_mult_82_n6536), 
        .ZN(u5_mult_82_ab_8__22_) );
  NAND2_X1 u5_mult_82_U8693 ( .A1(u5_mult_82_ab_22__9_), .A2(
        u5_mult_82_CARRYB_21__9_), .ZN(u5_mult_82_n3730) );
  NAND2_X2 u5_mult_82_U8692 ( .A1(u5_mult_82_ab_22__9_), .A2(
        u5_mult_82_SUMB_21__10_), .ZN(u5_mult_82_n3729) );
  XOR2_X2 u5_mult_82_U8691 ( .A(u5_mult_82_SUMB_21__10_), .B(u5_mult_82_n3727), 
        .Z(u5_mult_82_SUMB_22__9_) );
  XOR2_X2 u5_mult_82_U8690 ( .A(u5_mult_82_CARRYB_21__9_), .B(
        u5_mult_82_ab_22__9_), .Z(u5_mult_82_n3727) );
  NAND3_X2 u5_mult_82_U8689 ( .A1(u5_mult_82_n3720), .A2(u5_mult_82_n3721), 
        .A3(u5_mult_82_n3722), .ZN(u5_mult_82_CARRYB_10__20_) );
  NAND2_X1 u5_mult_82_U8688 ( .A1(u5_mult_82_CARRYB_9__20_), .A2(
        u5_mult_82_SUMB_9__21_), .ZN(u5_mult_82_n3722) );
  NAND2_X1 u5_mult_82_U8687 ( .A1(u5_mult_82_ab_10__20_), .A2(
        u5_mult_82_SUMB_9__21_), .ZN(u5_mult_82_n3721) );
  NAND2_X1 u5_mult_82_U8686 ( .A1(u5_mult_82_ab_10__20_), .A2(
        u5_mult_82_CARRYB_9__20_), .ZN(u5_mult_82_n3720) );
  NAND3_X2 u5_mult_82_U8685 ( .A1(u5_mult_82_n3717), .A2(u5_mult_82_n3718), 
        .A3(u5_mult_82_n3719), .ZN(u5_mult_82_CARRYB_9__21_) );
  NAND2_X2 u5_mult_82_U8684 ( .A1(u5_mult_82_CARRYB_8__21_), .A2(
        u5_mult_82_SUMB_8__22_), .ZN(u5_mult_82_n3719) );
  NAND2_X2 u5_mult_82_U8683 ( .A1(u5_mult_82_ab_9__21_), .A2(
        u5_mult_82_SUMB_8__22_), .ZN(u5_mult_82_n3718) );
  NAND2_X1 u5_mult_82_U8682 ( .A1(u5_mult_82_ab_9__21_), .A2(
        u5_mult_82_CARRYB_8__21_), .ZN(u5_mult_82_n3717) );
  XOR2_X2 u5_mult_82_U8681 ( .A(u5_mult_82_n3716), .B(u5_mult_82_SUMB_9__21_), 
        .Z(u5_mult_82_SUMB_10__20_) );
  XOR2_X2 u5_mult_82_U8680 ( .A(u5_mult_82_n3715), .B(u5_mult_82_SUMB_8__22_), 
        .Z(u5_mult_82_SUMB_9__21_) );
  XOR2_X2 u5_mult_82_U8679 ( .A(u5_mult_82_ab_9__21_), .B(
        u5_mult_82_CARRYB_8__21_), .Z(u5_mult_82_n3715) );
  NAND3_X2 u5_mult_82_U8678 ( .A1(u5_mult_82_n3712), .A2(u5_mult_82_n3713), 
        .A3(u5_mult_82_n3714), .ZN(u5_mult_82_CARRYB_8__22_) );
  NAND2_X1 u5_mult_82_U8677 ( .A1(u5_mult_82_ab_8__22_), .A2(
        u5_mult_82_CARRYB_7__22_), .ZN(u5_mult_82_n3714) );
  NAND2_X1 u5_mult_82_U8676 ( .A1(u5_mult_82_CARRYB_7__22_), .A2(
        u5_mult_82_SUMB_7__23_), .ZN(u5_mult_82_n3712) );
  XOR2_X2 u5_mult_82_U8675 ( .A(u5_mult_82_SUMB_7__23_), .B(u5_mult_82_n3711), 
        .Z(u5_mult_82_SUMB_8__22_) );
  XOR2_X2 u5_mult_82_U8674 ( .A(u5_mult_82_CARRYB_7__22_), .B(
        u5_mult_82_ab_8__22_), .Z(u5_mult_82_n3711) );
  XNOR2_X2 u5_mult_82_U8673 ( .A(u5_mult_82_n3710), .B(
        u5_mult_82_CARRYB_24__29_), .ZN(u5_mult_82_n5439) );
  INV_X4 u5_mult_82_U8672 ( .A(u5_mult_82_n3708), .ZN(u5_mult_82_n3709) );
  INV_X2 u5_mult_82_U8671 ( .A(u5_mult_82_SUMB_44__13_), .ZN(u5_mult_82_n3708)
         );
  INV_X4 u5_mult_82_U8670 ( .A(u5_mult_82_n3706), .ZN(u5_mult_82_n3707) );
  INV_X2 u5_mult_82_U8669 ( .A(u5_mult_82_SUMB_42__5_), .ZN(u5_mult_82_n3706)
         );
  XNOR2_X2 u5_mult_82_U8668 ( .A(u5_mult_82_ab_45__7_), .B(
        u5_mult_82_CARRYB_44__7_), .ZN(u5_mult_82_n3705) );
  XNOR2_X2 u5_mult_82_U8667 ( .A(u5_mult_82_n3705), .B(u5_mult_82_SUMB_44__8_), 
        .ZN(u5_mult_82_SUMB_45__7_) );
  XNOR2_X2 u5_mult_82_U8666 ( .A(u5_mult_82_CARRYB_41__2_), .B(
        u5_mult_82_ab_42__2_), .ZN(u5_mult_82_n4623) );
  XNOR2_X2 u5_mult_82_U8665 ( .A(u5_mult_82_CARRYB_50__25_), .B(
        u5_mult_82_n3704), .ZN(u5_mult_82_n4183) );
  XNOR2_X2 u5_mult_82_U8664 ( .A(u5_mult_82_CARRYB_32__13_), .B(
        u5_mult_82_n3703), .ZN(u5_mult_82_n5210) );
  XOR2_X2 u5_mult_82_U8663 ( .A(u5_mult_82_CARRYB_45__10_), .B(
        u5_mult_82_ab_46__10_), .Z(u5_mult_82_n6261) );
  NAND2_X1 u5_mult_82_U8662 ( .A1(u5_mult_82_ab_46__10_), .A2(
        u5_mult_82_CARRYB_45__10_), .ZN(u5_mult_82_n6262) );
  XNOR2_X2 u5_mult_82_U8661 ( .A(u5_mult_82_CARRYB_36__13_), .B(
        u5_mult_82_ab_37__13_), .ZN(u5_mult_82_net83047) );
  NAND2_X2 u5_mult_82_U8660 ( .A1(u5_mult_82_ab_50__24_), .A2(
        u5_mult_82_SUMB_49__25_), .ZN(u5_mult_82_n4446) );
  XNOR2_X2 u5_mult_82_U8659 ( .A(u5_mult_82_n3701), .B(
        u5_mult_82_CARRYB_41__27_), .ZN(u5_mult_82_n5581) );
  XNOR2_X2 u5_mult_82_U8658 ( .A(u5_mult_82_ab_46__4_), .B(
        u5_mult_82_CARRYB_45__4_), .ZN(u5_mult_82_n3700) );
  XNOR2_X2 u5_mult_82_U8657 ( .A(u5_mult_82_n3700), .B(u5_mult_82_n1411), .ZN(
        u5_mult_82_SUMB_46__4_) );
  NAND2_X2 u5_mult_82_U8656 ( .A1(u5_mult_82_CARRYB_42__24_), .A2(
        u5_mult_82_SUMB_42__25_), .ZN(u5_mult_82_n3876) );
  NAND2_X2 u5_mult_82_U8655 ( .A1(u5_mult_82_CARRYB_11__41_), .A2(
        u5_mult_82_SUMB_11__42_), .ZN(u5_mult_82_n5370) );
  XNOR2_X2 u5_mult_82_U8654 ( .A(u5_mult_82_CARRYB_7__44_), .B(
        u5_mult_82_ab_8__44_), .ZN(u5_mult_82_n3699) );
  XNOR2_X2 u5_mult_82_U8653 ( .A(u5_mult_82_n33), .B(u5_mult_82_n3699), .ZN(
        u5_mult_82_SUMB_8__44_) );
  INV_X2 u5_mult_82_U8652 ( .A(u5_mult_82_ab_39__11_), .ZN(u5_mult_82_n3696)
         );
  NAND2_X2 u5_mult_82_U8651 ( .A1(u5_mult_82_n5131), .A2(u5_mult_82_n3698), 
        .ZN(u5_mult_82_n4164) );
  NAND2_X2 u5_mult_82_U8650 ( .A1(u5_mult_82_n3696), .A2(u5_mult_82_n3697), 
        .ZN(u5_mult_82_n3698) );
  NAND2_X1 u5_mult_82_U8649 ( .A1(u5_mult_82_CARRYB_48__24_), .A2(
        u5_mult_82_SUMB_48__25_), .ZN(u5_mult_82_n4582) );
  NAND2_X2 u5_mult_82_U8648 ( .A1(u5_mult_82_ab_47__4_), .A2(
        u5_mult_82_SUMB_46__5_), .ZN(u5_mult_82_n6136) );
  NAND2_X2 u5_mult_82_U8647 ( .A1(u5_mult_82_CARRYB_37__16_), .A2(
        u5_mult_82_SUMB_37__17_), .ZN(u5_mult_82_n5432) );
  NAND2_X2 u5_mult_82_U8646 ( .A1(u5_mult_82_CARRYB_45__12_), .A2(
        u5_mult_82_SUMB_45__13_), .ZN(u5_mult_82_n5466) );
  NAND2_X2 u5_mult_82_U8645 ( .A1(u5_mult_82_n1833), .A2(
        u5_mult_82_CARRYB_44__2_), .ZN(u5_mult_82_n5630) );
  NAND2_X1 u5_mult_82_U8644 ( .A1(u5_mult_82_ab_21__37_), .A2(
        u5_mult_82_SUMB_20__38_), .ZN(u5_mult_82_n5518) );
  XOR2_X2 u5_mult_82_U8643 ( .A(u5_mult_82_CARRYB_44__4_), .B(u5_mult_82_n5856), .Z(u5_mult_82_n3695) );
  XNOR2_X2 u5_mult_82_U8642 ( .A(u5_mult_82_SUMB_44__5_), .B(u5_mult_82_n3695), 
        .ZN(u5_mult_82_SUMB_45__4_) );
  XNOR2_X2 u5_mult_82_U8641 ( .A(u5_mult_82_n4724), .B(u5_mult_82_n3694), .ZN(
        u5_mult_82_n4721) );
  XOR2_X2 u5_mult_82_U8640 ( .A(u5_mult_82_SUMB_19__38_), .B(u5_mult_82_n5783), 
        .Z(u5_mult_82_SUMB_20__37_) );
  NAND2_X2 u5_mult_82_U8639 ( .A1(u5_mult_82_CARRYB_12__41_), .A2(
        u5_mult_82_SUMB_12__42_), .ZN(u5_mult_82_n5175) );
  XNOR2_X2 u5_mult_82_U8638 ( .A(u5_mult_82_n3692), .B(
        u5_mult_82_CARRYB_45__23_), .ZN(u5_mult_82_n4703) );
  XNOR2_X2 u5_mult_82_U8637 ( .A(u5_mult_82_n3691), .B(u5_mult_82_SUMB_20__38_), .ZN(u5_mult_82_SUMB_21__37_) );
  NAND2_X2 u5_mult_82_U8636 ( .A1(u5_mult_82_CARRYB_7__48_), .A2(
        u5_mult_82_SUMB_7__49_), .ZN(u5_mult_82_n5722) );
  XNOR2_X2 u5_mult_82_U8635 ( .A(u5_mult_82_net83139), .B(u5_mult_82_n9), .ZN(
        u5_mult_82_SUMB_16__27_) );
  XNOR2_X2 u5_mult_82_U8634 ( .A(u5_mult_82_ab_39__29_), .B(
        u5_mult_82_CARRYB_38__29_), .ZN(u5_mult_82_n3690) );
  XNOR2_X2 u5_mult_82_U8633 ( .A(u5_mult_82_n3690), .B(u5_mult_82_SUMB_38__30_), .ZN(u5_mult_82_SUMB_39__29_) );
  XNOR2_X2 u5_mult_82_U8632 ( .A(u5_mult_82_CARRYB_3__49_), .B(
        u5_mult_82_ab_4__49_), .ZN(u5_mult_82_n3689) );
  XNOR2_X2 u5_mult_82_U8631 ( .A(u5_mult_82_SUMB_3__50_), .B(u5_mult_82_n3689), 
        .ZN(u5_mult_82_SUMB_4__49_) );
  NAND2_X2 u5_mult_82_U8630 ( .A1(u5_mult_82_CARRYB_40__3_), .A2(
        u5_mult_82_SUMB_40__4_), .ZN(u5_mult_82_n5158) );
  NAND2_X1 u5_mult_82_U8629 ( .A1(u5_mult_82_CARRYB_42__20_), .A2(
        u5_mult_82_SUMB_42__21_), .ZN(u5_mult_82_n4160) );
  NAND2_X1 u5_mult_82_U8628 ( .A1(u5_mult_82_n1469), .A2(
        u5_mult_82_CARRYB_42__8_), .ZN(u5_mult_82_n5933) );
  XNOR2_X2 u5_mult_82_U8627 ( .A(u5_mult_82_CARRYB_33__9_), .B(
        u5_mult_82_ab_34__9_), .ZN(u5_mult_82_n3688) );
  XNOR2_X2 u5_mult_82_U8626 ( .A(u5_mult_82_n3688), .B(u5_mult_82_SUMB_33__10_), .ZN(u5_mult_82_SUMB_34__9_) );
  XOR2_X2 u5_mult_82_U8625 ( .A(u5_mult_82_n4576), .B(u5_mult_82_n45), .Z(
        u5_mult_82_SUMB_49__24_) );
  NAND2_X4 u5_mult_82_U8624 ( .A1(u5_mult_82_n4689), .A2(u5_mult_82_n4688), 
        .ZN(u5_mult_82_SUMB_47__1_) );
  NAND3_X4 u5_mult_82_U8623 ( .A1(u5_mult_82_n4442), .A2(u5_mult_82_n4443), 
        .A3(u5_mult_82_n4444), .ZN(u5_mult_82_CARRYB_49__25_) );
  XNOR2_X2 u5_mult_82_U8622 ( .A(u5_mult_82_ab_42__24_), .B(
        u5_mult_82_CARRYB_41__24_), .ZN(u5_mult_82_n3687) );
  XNOR2_X2 u5_mult_82_U8621 ( .A(u5_mult_82_n3687), .B(u5_mult_82_SUMB_41__25_), .ZN(u5_mult_82_SUMB_42__24_) );
  NAND2_X2 u5_mult_82_U8620 ( .A1(u5_mult_82_ab_39__30_), .A2(
        u5_mult_82_SUMB_38__31_), .ZN(u5_mult_82_n3685) );
  NAND2_X1 u5_mult_82_U8619 ( .A1(u5_mult_82_ab_39__30_), .A2(
        u5_mult_82_CARRYB_38__30_), .ZN(u5_mult_82_n3684) );
  NAND3_X4 u5_mult_82_U8618 ( .A1(u5_mult_82_n3681), .A2(u5_mult_82_n3682), 
        .A3(u5_mult_82_n3683), .ZN(u5_mult_82_CARRYB_38__31_) );
  NAND2_X2 u5_mult_82_U8617 ( .A1(u5_mult_82_CARRYB_37__31_), .A2(
        u5_mult_82_n1850), .ZN(u5_mult_82_n3683) );
  NAND2_X2 u5_mult_82_U8616 ( .A1(u5_mult_82_ab_38__31_), .A2(u5_mult_82_n1850), .ZN(u5_mult_82_n3682) );
  NAND2_X2 u5_mult_82_U8615 ( .A1(u5_mult_82_ab_38__31_), .A2(
        u5_mult_82_CARRYB_37__31_), .ZN(u5_mult_82_n3681) );
  NAND3_X4 u5_mult_82_U8614 ( .A1(u5_mult_82_n3678), .A2(u5_mult_82_n3679), 
        .A3(u5_mult_82_n3680), .ZN(u5_mult_82_CARRYB_37__31_) );
  NAND2_X2 u5_mult_82_U8613 ( .A1(u5_mult_82_CARRYB_36__31_), .A2(
        u5_mult_82_SUMB_36__32_), .ZN(u5_mult_82_n3680) );
  NAND2_X2 u5_mult_82_U8612 ( .A1(u5_mult_82_ab_37__31_), .A2(
        u5_mult_82_SUMB_36__32_), .ZN(u5_mult_82_n3679) );
  NAND2_X1 u5_mult_82_U8611 ( .A1(u5_mult_82_ab_37__31_), .A2(
        u5_mult_82_CARRYB_36__31_), .ZN(u5_mult_82_n3678) );
  NAND2_X2 u5_mult_82_U8610 ( .A1(u5_mult_82_CARRYB_35__32_), .A2(
        u5_mult_82_SUMB_35__33_), .ZN(u5_mult_82_n3677) );
  NAND2_X2 u5_mult_82_U8609 ( .A1(u5_mult_82_ab_36__32_), .A2(
        u5_mult_82_SUMB_35__33_), .ZN(u5_mult_82_n3676) );
  NAND2_X1 u5_mult_82_U8608 ( .A1(u5_mult_82_ab_36__32_), .A2(
        u5_mult_82_CARRYB_35__32_), .ZN(u5_mult_82_n3675) );
  NAND3_X2 u5_mult_82_U8607 ( .A1(u5_mult_82_n3672), .A2(u5_mult_82_n3673), 
        .A3(u5_mult_82_n3674), .ZN(u5_mult_82_CARRYB_49__21_) );
  NAND2_X2 u5_mult_82_U8606 ( .A1(u5_mult_82_CARRYB_48__21_), .A2(
        u5_mult_82_SUMB_48__22_), .ZN(u5_mult_82_n3674) );
  NAND2_X2 u5_mult_82_U8605 ( .A1(u5_mult_82_ab_49__21_), .A2(
        u5_mult_82_SUMB_48__22_), .ZN(u5_mult_82_n3673) );
  NAND2_X1 u5_mult_82_U8604 ( .A1(u5_mult_82_ab_49__21_), .A2(
        u5_mult_82_CARRYB_48__21_), .ZN(u5_mult_82_n3672) );
  NAND3_X2 u5_mult_82_U8603 ( .A1(u5_mult_82_n3669), .A2(u5_mult_82_n3670), 
        .A3(u5_mult_82_n3671), .ZN(u5_mult_82_CARRYB_48__22_) );
  NAND2_X2 u5_mult_82_U8602 ( .A1(u5_mult_82_CARRYB_47__22_), .A2(
        u5_mult_82_SUMB_47__23_), .ZN(u5_mult_82_n3671) );
  NAND2_X2 u5_mult_82_U8601 ( .A1(u5_mult_82_ab_48__22_), .A2(
        u5_mult_82_SUMB_47__23_), .ZN(u5_mult_82_n3670) );
  NAND2_X1 u5_mult_82_U8600 ( .A1(u5_mult_82_ab_48__22_), .A2(
        u5_mult_82_CARRYB_47__22_), .ZN(u5_mult_82_n3669) );
  XOR2_X2 u5_mult_82_U8599 ( .A(u5_mult_82_n3668), .B(u5_mult_82_SUMB_48__22_), 
        .Z(u5_mult_82_SUMB_49__21_) );
  XOR2_X2 u5_mult_82_U8598 ( .A(u5_mult_82_ab_49__21_), .B(
        u5_mult_82_CARRYB_48__21_), .Z(u5_mult_82_n3668) );
  XOR2_X2 u5_mult_82_U8597 ( .A(u5_mult_82_ab_48__22_), .B(
        u5_mult_82_CARRYB_47__22_), .Z(u5_mult_82_n3667) );
  XNOR2_X2 u5_mult_82_U8596 ( .A(u5_mult_82_n3666), .B(
        u5_mult_82_CARRYB_29__17_), .ZN(u5_mult_82_n4559) );
  NAND2_X2 u5_mult_82_U8595 ( .A1(u5_mult_82_CARRYB_42__14_), .A2(
        u5_mult_82_SUMB_42__15_), .ZN(u5_mult_82_n6363) );
  XNOR2_X2 u5_mult_82_U8594 ( .A(u5_mult_82_CARRYB_4__28_), .B(
        u5_mult_82_n3665), .ZN(u5_mult_82_n4038) );
  NOR2_X1 u5_mult_82_U8593 ( .A1(u5_mult_82_net64687), .A2(u5_mult_82_n6602), 
        .ZN(u5_mult_82_ab_17__23_) );
  NOR2_X1 u5_mult_82_U8592 ( .A1(u5_mult_82_net64559), .A2(u5_mult_82_n6672), 
        .ZN(u5_mult_82_ab_29__16_) );
  NOR2_X4 u5_mult_82_U8591 ( .A1(u5_mult_82_net64433), .A2(u5_mult_82_net65373), .ZN(u5_mult_82_ab_42__9_) );
  NAND3_X4 u5_mult_82_U8590 ( .A1(u5_mult_82_n3662), .A2(u5_mult_82_n3663), 
        .A3(u5_mult_82_n3664), .ZN(u5_mult_82_CARRYB_17__23_) );
  NAND2_X1 u5_mult_82_U8589 ( .A1(u5_mult_82_ab_17__23_), .A2(
        u5_mult_82_CARRYB_16__23_), .ZN(u5_mult_82_n3664) );
  NAND2_X2 u5_mult_82_U8588 ( .A1(u5_mult_82_ab_17__23_), .A2(
        u5_mult_82_SUMB_16__24_), .ZN(u5_mult_82_n3663) );
  NAND2_X2 u5_mult_82_U8587 ( .A1(u5_mult_82_CARRYB_16__23_), .A2(
        u5_mult_82_SUMB_16__24_), .ZN(u5_mult_82_n3662) );
  NAND3_X2 u5_mult_82_U8586 ( .A1(u5_mult_82_n3659), .A2(u5_mult_82_n3660), 
        .A3(u5_mult_82_n3661), .ZN(u5_mult_82_CARRYB_31__14_) );
  NAND2_X2 u5_mult_82_U8585 ( .A1(u5_mult_82_ab_31__14_), .A2(
        u5_mult_82_SUMB_30__15_), .ZN(u5_mult_82_n3661) );
  NAND2_X1 u5_mult_82_U8584 ( .A1(u5_mult_82_CARRYB_30__14_), .A2(
        u5_mult_82_ab_31__14_), .ZN(u5_mult_82_n3659) );
  NAND2_X1 u5_mult_82_U8583 ( .A1(u5_mult_82_ab_30__15_), .A2(
        u5_mult_82_CARRYB_29__15_), .ZN(u5_mult_82_n3656) );
  XOR2_X2 u5_mult_82_U8582 ( .A(u5_mult_82_ab_30__15_), .B(
        u5_mult_82_CARRYB_29__15_), .Z(u5_mult_82_n3655) );
  NAND3_X2 u5_mult_82_U8581 ( .A1(u5_mult_82_n3652), .A2(u5_mult_82_n3653), 
        .A3(u5_mult_82_n3654), .ZN(u5_mult_82_CARRYB_29__16_) );
  NAND2_X1 u5_mult_82_U8580 ( .A1(u5_mult_82_ab_29__16_), .A2(
        u5_mult_82_CARRYB_28__16_), .ZN(u5_mult_82_n3654) );
  NAND2_X2 u5_mult_82_U8579 ( .A1(u5_mult_82_ab_29__16_), .A2(
        u5_mult_82_SUMB_28__17_), .ZN(u5_mult_82_n3653) );
  INV_X1 u5_mult_82_U8578 ( .A(u5_mult_82_ab_42__9_), .ZN(u5_mult_82_n3649) );
  NOR2_X1 u5_mult_82_U8577 ( .A1(u5_mult_82_n6839), .A2(u5_mult_82_n6608), 
        .ZN(u5_mult_82_ab_18__33_) );
  NAND2_X4 u5_mult_82_U8576 ( .A1(u5_mult_82_n4158), .A2(u5_mult_82_n4159), 
        .ZN(u5_mult_82_SUMB_48__18_) );
  NOR2_X2 u5_mult_82_U8575 ( .A1(u5_mult_82_n6927), .A2(u5_mult_82_n6754), 
        .ZN(u5_mult_82_ab_49__17_) );
  NOR2_X1 u5_mult_82_U8574 ( .A1(u5_mult_82_n6891), .A2(u5_mult_82_net65443), 
        .ZN(u5_mult_82_ab_38__24_) );
  NAND3_X2 u5_mult_82_U8573 ( .A1(u5_mult_82_n3645), .A2(u5_mult_82_n3646), 
        .A3(u5_mult_82_n3647), .ZN(u5_mult_82_CARRYB_18__33_) );
  NAND2_X1 u5_mult_82_U8572 ( .A1(u5_mult_82_ab_18__33_), .A2(
        u5_mult_82_CARRYB_17__33_), .ZN(u5_mult_82_n3647) );
  NAND2_X2 u5_mult_82_U8571 ( .A1(u5_mult_82_ab_18__33_), .A2(
        u5_mult_82_SUMB_17__34_), .ZN(u5_mult_82_n3646) );
  NAND3_X4 u5_mult_82_U8570 ( .A1(u5_mult_82_n3644), .A2(u5_mult_82_n3643), 
        .A3(u5_mult_82_n3642), .ZN(u5_mult_82_CARRYB_12__37_) );
  NAND2_X2 u5_mult_82_U8569 ( .A1(u5_mult_82_CARRYB_11__37_), .A2(
        u5_mult_82_n1386), .ZN(u5_mult_82_n3644) );
  NAND2_X2 u5_mult_82_U8568 ( .A1(u5_mult_82_ab_12__37_), .A2(u5_mult_82_n1386), .ZN(u5_mult_82_n3643) );
  NAND2_X1 u5_mult_82_U8567 ( .A1(u5_mult_82_ab_12__37_), .A2(
        u5_mult_82_CARRYB_11__37_), .ZN(u5_mult_82_n3642) );
  NAND3_X4 u5_mult_82_U8566 ( .A1(u5_mult_82_n3639), .A2(u5_mult_82_n3640), 
        .A3(u5_mult_82_n3641), .ZN(u5_mult_82_CARRYB_11__38_) );
  NAND2_X2 u5_mult_82_U8565 ( .A1(u5_mult_82_ab_11__38_), .A2(
        u5_mult_82_SUMB_10__39_), .ZN(u5_mult_82_n3640) );
  NAND2_X1 u5_mult_82_U8564 ( .A1(u5_mult_82_ab_11__38_), .A2(
        u5_mult_82_CARRYB_10__38_), .ZN(u5_mult_82_n3639) );
  NAND2_X2 u5_mult_82_U8563 ( .A1(u5_mult_82_ab_49__17_), .A2(
        u5_mult_82_CARRYB_48__17_), .ZN(u5_mult_82_n3637) );
  NAND2_X2 u5_mult_82_U8562 ( .A1(u5_mult_82_SUMB_48__18_), .A2(
        u5_mult_82_CARRYB_48__17_), .ZN(u5_mult_82_n3636) );
  NAND3_X2 u5_mult_82_U8561 ( .A1(u5_mult_82_n3633), .A2(u5_mult_82_n3634), 
        .A3(u5_mult_82_n3635), .ZN(u5_mult_82_CARRYB_38__24_) );
  NAND2_X1 u5_mult_82_U8560 ( .A1(u5_mult_82_CARRYB_37__24_), .A2(
        u5_mult_82_ab_38__24_), .ZN(u5_mult_82_n3635) );
  NAND2_X1 u5_mult_82_U8559 ( .A1(u5_mult_82_CARRYB_37__24_), .A2(
        u5_mult_82_SUMB_37__25_), .ZN(u5_mult_82_n3633) );
  XOR2_X2 u5_mult_82_U8558 ( .A(u5_mult_82_n3632), .B(u5_mult_82_SUMB_37__25_), 
        .Z(u5_mult_82_SUMB_38__24_) );
  NAND2_X1 u5_mult_82_U8557 ( .A1(u5_mult_82_CARRYB_50__15_), .A2(
        u5_mult_82_SUMB_50__16_), .ZN(u5_mult_82_n3631) );
  NAND2_X1 u5_mult_82_U8556 ( .A1(u5_mult_82_ab_51__15_), .A2(
        u5_mult_82_SUMB_50__16_), .ZN(u5_mult_82_n3630) );
  NAND2_X1 u5_mult_82_U8555 ( .A1(u5_mult_82_ab_51__15_), .A2(
        u5_mult_82_CARRYB_50__15_), .ZN(u5_mult_82_n3629) );
  NAND2_X2 u5_mult_82_U8554 ( .A1(u5_mult_82_CARRYB_49__16_), .A2(
        u5_mult_82_SUMB_49__17_), .ZN(u5_mult_82_n3628) );
  NAND2_X2 u5_mult_82_U8553 ( .A1(u5_mult_82_ab_50__16_), .A2(
        u5_mult_82_SUMB_49__17_), .ZN(u5_mult_82_n3627) );
  NAND2_X2 u5_mult_82_U8552 ( .A1(u5_mult_82_ab_50__16_), .A2(
        u5_mult_82_CARRYB_49__16_), .ZN(u5_mult_82_n3626) );
  XOR2_X2 u5_mult_82_U8551 ( .A(u5_mult_82_n3625), .B(u5_mult_82_SUMB_50__16_), 
        .Z(u5_mult_82_SUMB_51__15_) );
  XOR2_X2 u5_mult_82_U8550 ( .A(u5_mult_82_ab_51__15_), .B(
        u5_mult_82_CARRYB_50__15_), .Z(u5_mult_82_n3625) );
  XOR2_X2 u5_mult_82_U8549 ( .A(u5_mult_82_n3624), .B(u5_mult_82_SUMB_49__17_), 
        .Z(u5_mult_82_SUMB_50__16_) );
  XOR2_X2 u5_mult_82_U8548 ( .A(u5_mult_82_ab_50__16_), .B(
        u5_mult_82_CARRYB_49__16_), .Z(u5_mult_82_n3624) );
  NAND3_X2 u5_mult_82_U8547 ( .A1(u5_mult_82_n3621), .A2(u5_mult_82_n3622), 
        .A3(u5_mult_82_n3623), .ZN(u5_mult_82_CARRYB_27__8_) );
  NAND2_X1 u5_mult_82_U8546 ( .A1(u5_mult_82_ab_27__8_), .A2(
        u5_mult_82_CARRYB_26__8_), .ZN(u5_mult_82_n3621) );
  NAND2_X2 u5_mult_82_U8545 ( .A1(u5_mult_82_CARRYB_25__9_), .A2(
        u5_mult_82_SUMB_25__10_), .ZN(u5_mult_82_n3620) );
  NAND2_X2 u5_mult_82_U8544 ( .A1(u5_mult_82_ab_26__9_), .A2(
        u5_mult_82_SUMB_25__10_), .ZN(u5_mult_82_n3619) );
  NAND2_X1 u5_mult_82_U8543 ( .A1(u5_mult_82_ab_26__9_), .A2(
        u5_mult_82_CARRYB_25__9_), .ZN(u5_mult_82_n3618) );
  INV_X8 u5_mult_82_U8542 ( .A(n4738), .ZN(u5_mult_82_n7014) );
  INV_X4 u5_mult_82_U8541 ( .A(u5_mult_82_net83273), .ZN(u5_mult_82_net83274)
         );
  INV_X2 u5_mult_82_U8540 ( .A(u5_mult_82_SUMB_13__30_), .ZN(
        u5_mult_82_net83273) );
  NOR2_X2 u5_mult_82_U8539 ( .A1(u5_mult_82_net64687), .A2(u5_mult_82_n6629), 
        .ZN(u5_mult_82_ab_21__23_) );
  NOR2_X2 u5_mult_82_U8538 ( .A1(u5_mult_82_net64687), .A2(u5_mult_82_n6636), 
        .ZN(u5_mult_82_ab_22__23_) );
  NOR2_X1 u5_mult_82_U8537 ( .A1(u5_mult_82_net64887), .A2(u5_mult_82_n6521), 
        .ZN(u5_mult_82_ab_4__34_) );
  NAND3_X2 u5_mult_82_U8536 ( .A1(u5_mult_82_n6138), .A2(u5_mult_82_net79084), 
        .A3(u5_mult_82_net79086), .ZN(u5_mult_82_CARRYB_36__15_) );
  XOR2_X2 u5_mult_82_U8535 ( .A(u5_mult_82_CARRYB_21__23_), .B(
        u5_mult_82_n3614), .Z(u5_mult_82_SUMB_22__23_) );
  NAND2_X1 u5_mult_82_U8534 ( .A1(u5_mult_82_ab_32__17_), .A2(
        u5_mult_82_CARRYB_31__17_), .ZN(u5_mult_82_n3613) );
  NAND3_X2 u5_mult_82_U8533 ( .A1(u5_mult_82_net83288), .A2(
        u5_mult_82_net83289), .A3(u5_mult_82_net83290), .ZN(
        u5_mult_82_CARRYB_31__18_) );
  NAND2_X2 u5_mult_82_U8532 ( .A1(u5_mult_82_SUMB_41__24_), .A2(
        u5_mult_82_CARRYB_41__23_), .ZN(u5_mult_82_n5661) );
  NAND2_X2 u5_mult_82_U8531 ( .A1(u5_mult_82_ab_36__33_), .A2(
        u5_mult_82_CARRYB_35__33_), .ZN(u5_mult_82_n5577) );
  NOR2_X2 u5_mult_82_U8530 ( .A1(u5_mult_82_n6838), .A2(u5_mult_82_n6707), 
        .ZN(u5_mult_82_ab_35__33_) );
  NAND2_X2 u5_mult_82_U8529 ( .A1(u5_mult_82_ab_35__33_), .A2(
        u5_mult_82_CARRYB_34__33_), .ZN(u5_mult_82_n3611) );
  INV_X4 u5_mult_82_U8528 ( .A(u5_mult_82_n4183), .ZN(u5_mult_82_n3606) );
  NAND2_X2 u5_mult_82_U8527 ( .A1(u5_mult_82_n4183), .A2(u5_mult_82_n3607), 
        .ZN(u5_mult_82_n3608) );
  NAND3_X4 u5_mult_82_U8526 ( .A1(u5_mult_82_n6361), .A2(u5_mult_82_n6362), 
        .A3(u5_mult_82_n6363), .ZN(u5_mult_82_CARRYB_43__14_) );
  NAND2_X1 u5_mult_82_U8525 ( .A1(u5_mult_82_ab_45__13_), .A2(
        u5_mult_82_CARRYB_44__13_), .ZN(u5_mult_82_n5461) );
  NAND3_X2 u5_mult_82_U8524 ( .A1(u5_mult_82_n3602), .A2(u5_mult_82_n3603), 
        .A3(u5_mult_82_n3604), .ZN(u5_mult_82_CARRYB_12__50_) );
  NAND2_X2 u5_mult_82_U8523 ( .A1(u5_mult_82_ab_12__50_), .A2(
        u5_mult_82_CARRYB_11__50_), .ZN(u5_mult_82_n3603) );
  NAND3_X2 u5_mult_82_U8522 ( .A1(u5_mult_82_n3599), .A2(u5_mult_82_n3600), 
        .A3(u5_mult_82_n3601), .ZN(u5_mult_82_CARRYB_11__50_) );
  NAND2_X2 u5_mult_82_U8521 ( .A1(u5_mult_82_ab_11__50_), .A2(
        u5_mult_82_SUMB_10__51_), .ZN(u5_mult_82_n3600) );
  NAND3_X2 u5_mult_82_U8520 ( .A1(u5_mult_82_n3597), .A2(u5_mult_82_n3596), 
        .A3(u5_mult_82_n3598), .ZN(u5_mult_82_CARRYB_26__45_) );
  NAND2_X1 u5_mult_82_U8519 ( .A1(u5_mult_82_CARRYB_25__45_), .A2(
        u5_mult_82_SUMB_25__46_), .ZN(u5_mult_82_n3598) );
  NAND2_X1 u5_mult_82_U8518 ( .A1(u5_mult_82_ab_26__45_), .A2(
        u5_mult_82_SUMB_25__46_), .ZN(u5_mult_82_n3597) );
  NAND2_X1 u5_mult_82_U8517 ( .A1(u5_mult_82_ab_26__45_), .A2(
        u5_mult_82_CARRYB_25__45_), .ZN(u5_mult_82_n3596) );
  NAND2_X2 u5_mult_82_U8516 ( .A1(u5_mult_82_CARRYB_24__46_), .A2(
        u5_mult_82_SUMB_24__47_), .ZN(u5_mult_82_n3595) );
  NAND2_X2 u5_mult_82_U8515 ( .A1(u5_mult_82_ab_25__46_), .A2(
        u5_mult_82_SUMB_24__47_), .ZN(u5_mult_82_n3594) );
  NAND2_X2 u5_mult_82_U8514 ( .A1(u5_mult_82_ab_25__46_), .A2(
        u5_mult_82_CARRYB_24__46_), .ZN(u5_mult_82_n3593) );
  XOR2_X2 u5_mult_82_U8513 ( .A(u5_mult_82_n3592), .B(u5_mult_82_n1584), .Z(
        u5_mult_82_SUMB_25__46_) );
  XOR2_X2 u5_mult_82_U8512 ( .A(u5_mult_82_ab_25__46_), .B(
        u5_mult_82_CARRYB_24__46_), .Z(u5_mult_82_n3592) );
  INV_X8 u5_mult_82_U8511 ( .A(n4780), .ZN(u5_mult_82_n7013) );
  NAND2_X2 u5_mult_82_U8510 ( .A1(u5_mult_82_ab_37__17_), .A2(
        u5_mult_82_SUMB_36__18_), .ZN(u5_mult_82_n5966) );
  NAND2_X2 u5_mult_82_U8509 ( .A1(u5_mult_82_ab_46__12_), .A2(
        u5_mult_82_SUMB_45__13_), .ZN(u5_mult_82_n5465) );
  XOR2_X2 u5_mult_82_U8508 ( .A(u5_mult_82_ab_10__20_), .B(
        u5_mult_82_CARRYB_9__20_), .Z(u5_mult_82_n3716) );
  INV_X8 u5_mult_82_U8507 ( .A(n4758), .ZN(u5_mult_82_n7016) );
  NAND2_X2 u5_mult_82_U8506 ( .A1(u5_mult_82_ab_35__25_), .A2(
        u5_mult_82_CARRYB_34__25_), .ZN(u5_mult_82_n5029) );
  NAND2_X1 u5_mult_82_U8505 ( .A1(u5_mult_82_ab_33__18_), .A2(
        u5_mult_82_SUMB_32__19_), .ZN(u5_mult_82_n5983) );
  NAND2_X2 u5_mult_82_U8504 ( .A1(u5_mult_82_n5398), .A2(u5_mult_82_n1833), 
        .ZN(u5_mult_82_n4957) );
  XNOR2_X2 u5_mult_82_U8503 ( .A(u5_mult_82_n3591), .B(u5_mult_82_n27), .ZN(
        u5_mult_82_SUMB_42__6_) );
  XNOR2_X2 u5_mult_82_U8502 ( .A(u5_mult_82_SUMB_16__25_), .B(u5_mult_82_n4023), .ZN(u5_mult_82_SUMB_17__24_) );
  XNOR2_X2 u5_mult_82_U8501 ( .A(u5_mult_82_CARRYB_26__11_), .B(
        u5_mult_82_n3590), .ZN(u5_mult_82_n4970) );
  XNOR2_X2 u5_mult_82_U8500 ( .A(u5_mult_82_SUMB_41__9_), .B(u5_mult_82_n3589), 
        .ZN(u5_mult_82_n4384) );
  NAND3_X4 u5_mult_82_U8499 ( .A1(u5_mult_82_n5962), .A2(u5_mult_82_n5963), 
        .A3(u5_mult_82_n5964), .ZN(u5_mult_82_CARRYB_36__18_) );
  XNOR2_X1 u5_mult_82_U8498 ( .A(u5_mult_82_n5508), .B(u5_mult_82_SUMB_48__11_), .ZN(u5_mult_82_SUMB_49__10_) );
  XNOR2_X2 u5_mult_82_U8497 ( .A(u5_mult_82_CARRYB_38__28_), .B(
        u5_mult_82_ab_39__28_), .ZN(u5_mult_82_n3587) );
  XNOR2_X2 u5_mult_82_U8496 ( .A(u5_mult_82_SUMB_38__29_), .B(u5_mult_82_n3587), .ZN(u5_mult_82_SUMB_39__28_) );
  INV_X4 u5_mult_82_U8495 ( .A(u5_mult_82_ab_33__31_), .ZN(u5_mult_82_n3605)
         );
  NAND2_X4 u5_mult_82_U8494 ( .A1(u5_mult_82_n3584), .A2(u5_mult_82_n3583), 
        .ZN(u5_mult_82_n3586) );
  XNOR2_X2 u5_mult_82_U8493 ( .A(u5_mult_82_n3582), .B(u5_mult_82_SUMB_30__20_), .ZN(u5_mult_82_SUMB_31__19_) );
  NAND2_X2 u5_mult_82_U8492 ( .A1(u5_mult_82_ab_37__16_), .A2(u5_mult_82_n738), 
        .ZN(u5_mult_82_n5524) );
  NAND2_X1 u5_mult_82_U8491 ( .A1(u5_mult_82_ab_3__36_), .A2(
        u5_mult_82_SUMB_2__37_), .ZN(u5_mult_82_n5155) );
  NAND2_X2 u5_mult_82_U8490 ( .A1(u5_mult_82_CARRYB_46__6_), .A2(
        u5_mult_82_SUMB_46__7_), .ZN(u5_mult_82_n5930) );
  NAND3_X4 u5_mult_82_U8489 ( .A1(u5_mult_82_n5932), .A2(u5_mult_82_n5931), 
        .A3(u5_mult_82_n5930), .ZN(u5_mult_82_CARRYB_47__6_) );
  NAND2_X1 u5_mult_82_U8488 ( .A1(u5_mult_82_ab_44__14_), .A2(
        u5_mult_82_CARRYB_43__14_), .ZN(u5_mult_82_n5459) );
  XNOR2_X2 u5_mult_82_U8487 ( .A(u5_mult_82_CARRYB_25__10_), .B(
        u5_mult_82_ab_26__10_), .ZN(u5_mult_82_n3581) );
  XNOR2_X2 u5_mult_82_U8486 ( .A(u5_mult_82_SUMB_25__11_), .B(u5_mult_82_n3581), .ZN(u5_mult_82_SUMB_26__10_) );
  NAND2_X1 u5_mult_82_U8485 ( .A1(u5_mult_82_ab_33__31_), .A2(
        u5_mult_82_CARRYB_32__31_), .ZN(u5_mult_82_n5946) );
  NAND3_X4 u5_mult_82_U8484 ( .A1(u5_mult_82_n5770), .A2(u5_mult_82_n5771), 
        .A3(u5_mult_82_n5772), .ZN(u5_mult_82_CARRYB_47__14_) );
  NOR2_X1 u5_mult_82_U8483 ( .A1(u5_mult_82_net64469), .A2(u5_mult_82_net65517), .ZN(u5_mult_82_ab_34__11_) );
  NAND3_X2 u5_mult_82_U8482 ( .A1(u5_mult_82_n3577), .A2(u5_mult_82_n3578), 
        .A3(u5_mult_82_n3579), .ZN(u5_mult_82_CARRYB_34__11_) );
  NAND2_X1 u5_mult_82_U8481 ( .A1(u5_mult_82_ab_34__11_), .A2(
        u5_mult_82_CARRYB_33__11_), .ZN(u5_mult_82_n3579) );
  NAND2_X1 u5_mult_82_U8480 ( .A1(u5_mult_82_CARRYB_33__11_), .A2(
        u5_mult_82_SUMB_33__12_), .ZN(u5_mult_82_n3577) );
  NAND2_X2 u5_mult_82_U8479 ( .A1(u5_mult_82_CARRYB_25__17_), .A2(
        u5_mult_82_SUMB_25__18_), .ZN(u5_mult_82_n3576) );
  NAND2_X2 u5_mult_82_U8478 ( .A1(u5_mult_82_ab_26__17_), .A2(
        u5_mult_82_SUMB_25__18_), .ZN(u5_mult_82_n3575) );
  NAND2_X1 u5_mult_82_U8477 ( .A1(u5_mult_82_ab_26__17_), .A2(
        u5_mult_82_CARRYB_25__17_), .ZN(u5_mult_82_n3574) );
  NAND3_X2 u5_mult_82_U8476 ( .A1(u5_mult_82_n3571), .A2(u5_mult_82_n3572), 
        .A3(u5_mult_82_n3573), .ZN(u5_mult_82_CARRYB_25__18_) );
  NAND2_X2 u5_mult_82_U8475 ( .A1(u5_mult_82_n85), .A2(
        u5_mult_82_CARRYB_24__18_), .ZN(u5_mult_82_n3573) );
  NAND2_X2 u5_mult_82_U8474 ( .A1(u5_mult_82_ab_25__18_), .A2(u5_mult_82_n85), 
        .ZN(u5_mult_82_n3572) );
  NAND2_X1 u5_mult_82_U8473 ( .A1(u5_mult_82_ab_25__18_), .A2(
        u5_mult_82_CARRYB_24__18_), .ZN(u5_mult_82_n3571) );
  XOR2_X2 u5_mult_82_U8472 ( .A(u5_mult_82_n3570), .B(u5_mult_82_SUMB_25__18_), 
        .Z(u5_mult_82_SUMB_26__17_) );
  XOR2_X2 u5_mult_82_U8471 ( .A(u5_mult_82_ab_26__17_), .B(
        u5_mult_82_CARRYB_25__17_), .Z(u5_mult_82_n3570) );
  XOR2_X2 u5_mult_82_U8470 ( .A(u5_mult_82_n3569), .B(u5_mult_82_n85), .Z(
        u5_mult_82_SUMB_25__18_) );
  XOR2_X2 u5_mult_82_U8469 ( .A(u5_mult_82_ab_25__18_), .B(
        u5_mult_82_CARRYB_24__18_), .Z(u5_mult_82_n3569) );
  NOR2_X1 u5_mult_82_U8468 ( .A1(u5_mult_82_n6947), .A2(u5_mult_82_net65679), 
        .ZN(u5_mult_82_ab_25__4_) );
  NOR2_X1 u5_mult_82_U8467 ( .A1(u5_mult_82_net64563), .A2(u5_mult_82_n6572), 
        .ZN(u5_mult_82_ab_13__16_) );
  NAND3_X2 u5_mult_82_U8466 ( .A1(u5_mult_82_n3566), .A2(u5_mult_82_n3567), 
        .A3(u5_mult_82_n3568), .ZN(u5_mult_82_CARRYB_25__4_) );
  NAND2_X1 u5_mult_82_U8465 ( .A1(u5_mult_82_ab_25__4_), .A2(
        u5_mult_82_CARRYB_24__4_), .ZN(u5_mult_82_n3568) );
  NAND2_X2 u5_mult_82_U8464 ( .A1(u5_mult_82_ab_25__4_), .A2(
        u5_mult_82_SUMB_24__5_), .ZN(u5_mult_82_n3567) );
  NAND2_X1 u5_mult_82_U8463 ( .A1(u5_mult_82_CARRYB_24__4_), .A2(
        u5_mult_82_SUMB_24__5_), .ZN(u5_mult_82_n3566) );
  XOR2_X2 u5_mult_82_U8462 ( .A(u5_mult_82_SUMB_24__5_), .B(u5_mult_82_n3565), 
        .Z(u5_mult_82_SUMB_25__4_) );
  XOR2_X2 u5_mult_82_U8461 ( .A(u5_mult_82_CARRYB_24__4_), .B(
        u5_mult_82_ab_25__4_), .Z(u5_mult_82_n3565) );
  NAND2_X2 u5_mult_82_U8460 ( .A1(u5_mult_82_n3562), .A2(u5_mult_82_n1781), 
        .ZN(u5_mult_82_n3564) );
  NAND3_X2 u5_mult_82_U8459 ( .A1(u5_mult_82_n3559), .A2(u5_mult_82_n3560), 
        .A3(u5_mult_82_n3561), .ZN(u5_mult_82_CARRYB_3__26_) );
  NAND2_X1 u5_mult_82_U8458 ( .A1(u5_mult_82_CARRYB_2__26_), .A2(
        u5_mult_82_SUMB_2__27_), .ZN(u5_mult_82_n3561) );
  NAND2_X1 u5_mult_82_U8457 ( .A1(u5_mult_82_ab_3__26_), .A2(
        u5_mult_82_SUMB_2__27_), .ZN(u5_mult_82_n3560) );
  NAND2_X1 u5_mult_82_U8456 ( .A1(u5_mult_82_ab_3__26_), .A2(
        u5_mult_82_CARRYB_2__26_), .ZN(u5_mult_82_n3559) );
  NAND3_X2 u5_mult_82_U8455 ( .A1(u5_mult_82_n3556), .A2(u5_mult_82_n3557), 
        .A3(u5_mult_82_n3558), .ZN(u5_mult_82_CARRYB_2__27_) );
  NAND2_X2 u5_mult_82_U8454 ( .A1(u5_mult_82_CARRYB_1__27_), .A2(
        u5_mult_82_n469), .ZN(u5_mult_82_n3558) );
  NAND2_X2 u5_mult_82_U8453 ( .A1(u5_mult_82_ab_2__27_), .A2(u5_mult_82_n469), 
        .ZN(u5_mult_82_n3557) );
  NAND2_X1 u5_mult_82_U8452 ( .A1(u5_mult_82_ab_2__27_), .A2(
        u5_mult_82_CARRYB_1__27_), .ZN(u5_mult_82_n3556) );
  XOR2_X2 u5_mult_82_U8451 ( .A(u5_mult_82_n3555), .B(u5_mult_82_n469), .Z(
        u5_mult_82_SUMB_2__27_) );
  XOR2_X2 u5_mult_82_U8450 ( .A(u5_mult_82_ab_2__27_), .B(
        u5_mult_82_CARRYB_1__27_), .Z(u5_mult_82_n3555) );
  NAND3_X2 u5_mult_82_U8449 ( .A1(u5_mult_82_n3552), .A2(u5_mult_82_n3553), 
        .A3(u5_mult_82_n3554), .ZN(u5_mult_82_CARRYB_15__14_) );
  NAND2_X1 u5_mult_82_U8448 ( .A1(u5_mult_82_CARRYB_14__14_), .A2(
        u5_mult_82_SUMB_14__15_), .ZN(u5_mult_82_n3554) );
  NAND2_X1 u5_mult_82_U8447 ( .A1(u5_mult_82_ab_15__14_), .A2(
        u5_mult_82_SUMB_14__15_), .ZN(u5_mult_82_n3553) );
  NAND3_X2 u5_mult_82_U8446 ( .A1(u5_mult_82_n3549), .A2(u5_mult_82_n3550), 
        .A3(u5_mult_82_n3551), .ZN(u5_mult_82_CARRYB_14__15_) );
  NAND2_X2 u5_mult_82_U8445 ( .A1(u5_mult_82_CARRYB_13__15_), .A2(
        u5_mult_82_SUMB_13__16_), .ZN(u5_mult_82_n3551) );
  NAND2_X2 u5_mult_82_U8444 ( .A1(u5_mult_82_ab_14__15_), .A2(
        u5_mult_82_SUMB_13__16_), .ZN(u5_mult_82_n3550) );
  NAND2_X1 u5_mult_82_U8443 ( .A1(u5_mult_82_ab_14__15_), .A2(
        u5_mult_82_CARRYB_13__15_), .ZN(u5_mult_82_n3549) );
  XOR2_X2 u5_mult_82_U8442 ( .A(u5_mult_82_n3548), .B(u5_mult_82_SUMB_14__15_), 
        .Z(u5_mult_82_SUMB_15__14_) );
  XOR2_X2 u5_mult_82_U8441 ( .A(u5_mult_82_ab_15__14_), .B(
        u5_mult_82_CARRYB_14__14_), .Z(u5_mult_82_n3548) );
  XOR2_X2 u5_mult_82_U8440 ( .A(u5_mult_82_n3547), .B(u5_mult_82_SUMB_13__16_), 
        .Z(u5_mult_82_SUMB_14__15_) );
  XOR2_X2 u5_mult_82_U8439 ( .A(u5_mult_82_ab_14__15_), .B(
        u5_mult_82_CARRYB_13__15_), .Z(u5_mult_82_n3547) );
  NAND3_X2 u5_mult_82_U8438 ( .A1(u5_mult_82_n3544), .A2(u5_mult_82_n3545), 
        .A3(u5_mult_82_n3546), .ZN(u5_mult_82_CARRYB_13__16_) );
  NAND2_X1 u5_mult_82_U8437 ( .A1(u5_mult_82_ab_13__16_), .A2(
        u5_mult_82_CARRYB_12__16_), .ZN(u5_mult_82_n3546) );
  NAND2_X2 u5_mult_82_U8436 ( .A1(u5_mult_82_ab_13__16_), .A2(
        u5_mult_82_SUMB_12__17_), .ZN(u5_mult_82_n3545) );
  XOR2_X2 u5_mult_82_U8435 ( .A(u5_mult_82_SUMB_12__17_), .B(u5_mult_82_n3543), 
        .Z(u5_mult_82_SUMB_13__16_) );
  XOR2_X2 u5_mult_82_U8434 ( .A(u5_mult_82_CARRYB_12__16_), .B(
        u5_mult_82_ab_13__16_), .Z(u5_mult_82_n3543) );
  INV_X4 u5_mult_82_U8433 ( .A(u5_mult_82_n5297), .ZN(u5_mult_82_n3539) );
  NAND3_X2 u5_mult_82_U8432 ( .A1(u5_mult_82_n3536), .A2(u5_mult_82_n3537), 
        .A3(u5_mult_82_n3538), .ZN(u5_mult_82_CARRYB_20__32_) );
  NAND2_X2 u5_mult_82_U8431 ( .A1(u5_mult_82_ab_20__32_), .A2(
        u5_mult_82_SUMB_19__33_), .ZN(u5_mult_82_n3537) );
  NAND2_X2 u5_mult_82_U8430 ( .A1(u5_mult_82_CARRYB_18__33_), .A2(
        u5_mult_82_SUMB_18__34_), .ZN(u5_mult_82_n3535) );
  NAND2_X2 u5_mult_82_U8429 ( .A1(u5_mult_82_ab_19__33_), .A2(
        u5_mult_82_SUMB_18__34_), .ZN(u5_mult_82_n3534) );
  NAND2_X1 u5_mult_82_U8428 ( .A1(u5_mult_82_ab_19__33_), .A2(
        u5_mult_82_CARRYB_18__33_), .ZN(u5_mult_82_n3533) );
  NAND3_X2 u5_mult_82_U8427 ( .A1(u5_mult_82_n3530), .A2(u5_mult_82_n3531), 
        .A3(u5_mult_82_n3532), .ZN(u5_mult_82_CARRYB_3__41_) );
  NAND2_X1 u5_mult_82_U8426 ( .A1(u5_mult_82_CARRYB_2__41_), .A2(
        u5_mult_82_SUMB_2__42_), .ZN(u5_mult_82_n3532) );
  NAND2_X1 u5_mult_82_U8425 ( .A1(u5_mult_82_ab_3__41_), .A2(
        u5_mult_82_SUMB_2__42_), .ZN(u5_mult_82_n3531) );
  NAND2_X1 u5_mult_82_U8424 ( .A1(u5_mult_82_ab_3__41_), .A2(
        u5_mult_82_CARRYB_2__41_), .ZN(u5_mult_82_n3530) );
  NAND2_X2 u5_mult_82_U8423 ( .A1(u5_mult_82_CARRYB_1__42_), .A2(
        u5_mult_82_n481), .ZN(u5_mult_82_n3529) );
  NAND2_X2 u5_mult_82_U8422 ( .A1(u5_mult_82_ab_2__42_), .A2(u5_mult_82_n481), 
        .ZN(u5_mult_82_n3528) );
  NAND2_X1 u5_mult_82_U8421 ( .A1(u5_mult_82_ab_2__42_), .A2(
        u5_mult_82_CARRYB_1__42_), .ZN(u5_mult_82_n3527) );
  XOR2_X2 u5_mult_82_U8420 ( .A(u5_mult_82_n3526), .B(u5_mult_82_n481), .Z(
        u5_mult_82_SUMB_2__42_) );
  XOR2_X2 u5_mult_82_U8419 ( .A(u5_mult_82_ab_2__42_), .B(
        u5_mult_82_CARRYB_1__42_), .Z(u5_mult_82_n3526) );
  NAND3_X4 u5_mult_82_U8418 ( .A1(u5_mult_82_n3523), .A2(u5_mult_82_n3524), 
        .A3(u5_mult_82_n3525), .ZN(u5_mult_82_CARRYB_32__22_) );
  NAND2_X2 u5_mult_82_U8417 ( .A1(u5_mult_82_ab_32__22_), .A2(
        u5_mult_82_SUMB_31__23_), .ZN(u5_mult_82_n3524) );
  NAND2_X1 u5_mult_82_U8416 ( .A1(u5_mult_82_ab_32__22_), .A2(
        u5_mult_82_CARRYB_31__22_), .ZN(u5_mult_82_n3523) );
  NAND3_X2 u5_mult_82_U8415 ( .A1(u5_mult_82_n3520), .A2(u5_mult_82_n3521), 
        .A3(u5_mult_82_n3522), .ZN(u5_mult_82_CARRYB_31__23_) );
  NAND2_X2 u5_mult_82_U8414 ( .A1(u5_mult_82_CARRYB_30__23_), .A2(
        u5_mult_82_SUMB_30__24_), .ZN(u5_mult_82_n3522) );
  NAND2_X2 u5_mult_82_U8413 ( .A1(u5_mult_82_ab_31__23_), .A2(
        u5_mult_82_SUMB_30__24_), .ZN(u5_mult_82_n3521) );
  NAND2_X1 u5_mult_82_U8412 ( .A1(u5_mult_82_ab_31__23_), .A2(
        u5_mult_82_CARRYB_30__23_), .ZN(u5_mult_82_n3520) );
  XOR2_X2 u5_mult_82_U8411 ( .A(u5_mult_82_n3519), .B(u5_mult_82_SUMB_31__23_), 
        .Z(u5_mult_82_SUMB_32__22_) );
  NAND3_X4 u5_mult_82_U8410 ( .A1(u5_mult_82_n3516), .A2(u5_mult_82_n3517), 
        .A3(u5_mult_82_n3518), .ZN(u5_mult_82_CARRYB_28__25_) );
  NAND2_X2 u5_mult_82_U8409 ( .A1(u5_mult_82_CARRYB_27__25_), .A2(
        u5_mult_82_SUMB_27__26_), .ZN(u5_mult_82_n3518) );
  NAND2_X2 u5_mult_82_U8408 ( .A1(u5_mult_82_ab_28__25_), .A2(
        u5_mult_82_SUMB_27__26_), .ZN(u5_mult_82_n3517) );
  NAND2_X1 u5_mult_82_U8407 ( .A1(u5_mult_82_ab_28__25_), .A2(
        u5_mult_82_CARRYB_27__25_), .ZN(u5_mult_82_n3516) );
  NAND3_X2 u5_mult_82_U8406 ( .A1(u5_mult_82_n3515), .A2(u5_mult_82_n3514), 
        .A3(u5_mult_82_n3513), .ZN(u5_mult_82_CARRYB_27__26_) );
  NAND2_X2 u5_mult_82_U8405 ( .A1(u5_mult_82_CARRYB_26__26_), .A2(
        u5_mult_82_SUMB_26__27_), .ZN(u5_mult_82_n3515) );
  NAND2_X2 u5_mult_82_U8404 ( .A1(u5_mult_82_ab_27__26_), .A2(
        u5_mult_82_SUMB_26__27_), .ZN(u5_mult_82_n3514) );
  NAND2_X1 u5_mult_82_U8403 ( .A1(u5_mult_82_ab_27__26_), .A2(
        u5_mult_82_CARRYB_26__26_), .ZN(u5_mult_82_n3513) );
  XOR2_X2 u5_mult_82_U8402 ( .A(u5_mult_82_ab_28__25_), .B(
        u5_mult_82_CARRYB_27__25_), .Z(u5_mult_82_n3512) );
  XOR2_X2 u5_mult_82_U8401 ( .A(u5_mult_82_n3511), .B(u5_mult_82_n1769), .Z(
        u5_mult_82_SUMB_27__26_) );
  XOR2_X2 u5_mult_82_U8400 ( .A(u5_mult_82_ab_27__26_), .B(
        u5_mult_82_CARRYB_26__26_), .Z(u5_mult_82_n3511) );
  XNOR2_X2 u5_mult_82_U8399 ( .A(u5_mult_82_ab_18__36_), .B(
        u5_mult_82_CARRYB_17__36_), .ZN(u5_mult_82_n3510) );
  NAND2_X1 u5_mult_82_U8398 ( .A1(u5_mult_82_CARRYB_47__10_), .A2(
        u5_mult_82_SUMB_47__11_), .ZN(u5_mult_82_n6211) );
  NAND2_X2 u5_mult_82_U8397 ( .A1(u5_mult_82_n1548), .A2(u5_mult_82_n1752), 
        .ZN(u5_mult_82_n6005) );
  XNOR2_X2 u5_mult_82_U8396 ( .A(u5_mult_82_ab_46__13_), .B(
        u5_mult_82_CARRYB_45__13_), .ZN(u5_mult_82_n3509) );
  XNOR2_X2 u5_mult_82_U8395 ( .A(u5_mult_82_n3509), .B(u5_mult_82_SUMB_45__14_), .ZN(u5_mult_82_SUMB_46__13_) );
  NAND2_X2 u5_mult_82_U8394 ( .A1(u5_mult_82_ab_14__40_), .A2(
        u5_mult_82_SUMB_13__41_), .ZN(u5_mult_82_n5386) );
  XOR2_X2 u5_mult_82_U8393 ( .A(u5_mult_82_n3856), .B(u5_mult_82_SUMB_40__24_), 
        .Z(u5_mult_82_SUMB_41__23_) );
  NAND2_X2 u5_mult_82_U8392 ( .A1(u5_mult_82_CARRYB_19__40_), .A2(
        u5_mult_82_n66), .ZN(u5_mult_82_n4943) );
  NAND2_X2 u5_mult_82_U8391 ( .A1(u5_mult_82_CARRYB_21__39_), .A2(
        u5_mult_82_SUMB_21__40_), .ZN(u5_mult_82_n5999) );
  NAND3_X4 u5_mult_82_U8390 ( .A1(u5_mult_82_n5259), .A2(u5_mult_82_n5260), 
        .A3(u5_mult_82_n5261), .ZN(u5_mult_82_CARRYB_48__9_) );
  NAND3_X2 u5_mult_82_U8389 ( .A1(u5_mult_82_n5466), .A2(u5_mult_82_n5465), 
        .A3(u5_mult_82_n5464), .ZN(u5_mult_82_CARRYB_46__12_) );
  XNOR2_X2 u5_mult_82_U8388 ( .A(u5_mult_82_n3508), .B(
        u5_mult_82_CARRYB_8__47_), .ZN(u5_mult_82_n5725) );
  XNOR2_X2 u5_mult_82_U8387 ( .A(u5_mult_82_ab_10__46_), .B(
        u5_mult_82_CARRYB_9__46_), .ZN(u5_mult_82_n3507) );
  NAND2_X2 u5_mult_82_U8386 ( .A1(u5_mult_82_ab_2__50_), .A2(
        u5_mult_82_CARRYB_1__50_), .ZN(u5_mult_82_n3506) );
  NAND2_X2 u5_mult_82_U8385 ( .A1(u5_mult_82_CARRYB_1__50_), .A2(
        u5_mult_82_SUMB_1__51_), .ZN(u5_mult_82_n3504) );
  XOR2_X2 u5_mult_82_U8384 ( .A(u5_mult_82_n3503), .B(u5_mult_82_SUMB_1__51_), 
        .Z(u5_mult_82_SUMB_2__50_) );
  XOR2_X2 u5_mult_82_U8383 ( .A(u5_mult_82_CARRYB_1__50_), .B(
        u5_mult_82_ab_2__50_), .Z(u5_mult_82_n3503) );
  XNOR2_X2 u5_mult_82_U8382 ( .A(u5_mult_82_ab_51__8_), .B(
        u5_mult_82_CARRYB_50__8_), .ZN(u5_mult_82_n3502) );
  XNOR2_X2 u5_mult_82_U8381 ( .A(u5_mult_82_n3502), .B(u5_mult_82_SUMB_50__9_), 
        .ZN(u5_mult_82_SUMB_51__8_) );
  XNOR2_X2 u5_mult_82_U8380 ( .A(u5_mult_82_n3501), .B(
        u5_mult_82_CARRYB_16__36_), .ZN(u5_mult_82_n6308) );
  XNOR2_X2 u5_mult_82_U8379 ( .A(u5_mult_82_SUMB_44__9_), .B(u5_mult_82_n3500), 
        .ZN(u5_mult_82_n4218) );
  XNOR2_X1 u5_mult_82_U8378 ( .A(u5_mult_82_ab_22__18_), .B(
        u5_mult_82_SUMB_21__19_), .ZN(u5_mult_82_n3499) );
  XNOR2_X2 u5_mult_82_U8377 ( .A(u5_mult_82_n3499), .B(
        u5_mult_82_CARRYB_21__18_), .ZN(u5_mult_82_SUMB_22__18_) );
  NAND2_X2 u5_mult_82_U8376 ( .A1(u5_mult_82_SUMB_38__11_), .A2(
        u5_mult_82_CARRYB_38__10_), .ZN(u5_mult_82_n3993) );
  XNOR2_X2 u5_mult_82_U8375 ( .A(u5_mult_82_n3498), .B(u5_mult_82_n1541), .ZN(
        u5_mult_82_SUMB_48__11_) );
  NAND2_X2 u5_mult_82_U8374 ( .A1(u5_mult_82_ab_43__7_), .A2(
        u5_mult_82_CARRYB_42__7_), .ZN(u5_mult_82_n6071) );
  NAND2_X2 u5_mult_82_U8373 ( .A1(u5_mult_82_ab_47__5_), .A2(
        u5_mult_82_SUMB_46__6_), .ZN(u5_mult_82_n6170) );
  XNOR2_X2 u5_mult_82_U8372 ( .A(u5_mult_82_ab_39__34_), .B(
        u5_mult_82_CARRYB_38__34_), .ZN(u5_mult_82_n3497) );
  XNOR2_X2 u5_mult_82_U8371 ( .A(u5_mult_82_n3497), .B(u5_mult_82_SUMB_38__35_), .ZN(u5_mult_82_SUMB_39__34_) );
  XNOR2_X2 u5_mult_82_U8370 ( .A(u5_mult_82_ab_26__45_), .B(
        u5_mult_82_CARRYB_25__45_), .ZN(u5_mult_82_n3496) );
  NAND2_X1 u5_mult_82_U8369 ( .A1(u5_mult_82_ab_42__23_), .A2(
        u5_mult_82_SUMB_41__24_), .ZN(u5_mult_82_n5662) );
  INV_X4 u5_mult_82_U8368 ( .A(u5_mult_82_n3494), .ZN(u5_mult_82_n3495) );
  NAND2_X2 u5_mult_82_U8367 ( .A1(u5_mult_82_n5663), .A2(u5_mult_82_n5661), 
        .ZN(u5_mult_82_n3494) );
  NAND3_X2 u5_mult_82_U8366 ( .A1(u5_mult_82_n3491), .A2(u5_mult_82_n3492), 
        .A3(u5_mult_82_n3493), .ZN(u5_mult_82_CARRYB_40__25_) );
  NAND2_X1 u5_mult_82_U8365 ( .A1(u5_mult_82_CARRYB_39__25_), .A2(
        u5_mult_82_SUMB_39__26_), .ZN(u5_mult_82_n3493) );
  NAND2_X1 u5_mult_82_U8364 ( .A1(u5_mult_82_ab_40__25_), .A2(
        u5_mult_82_SUMB_39__26_), .ZN(u5_mult_82_n3492) );
  NAND2_X1 u5_mult_82_U8363 ( .A1(u5_mult_82_ab_40__25_), .A2(
        u5_mult_82_CARRYB_39__25_), .ZN(u5_mult_82_n3491) );
  NAND3_X2 u5_mult_82_U8362 ( .A1(u5_mult_82_n3489), .A2(u5_mult_82_n3488), 
        .A3(u5_mult_82_n3490), .ZN(u5_mult_82_CARRYB_39__26_) );
  NAND2_X1 u5_mult_82_U8361 ( .A1(u5_mult_82_CARRYB_38__26_), .A2(
        u5_mult_82_SUMB_38__27_), .ZN(u5_mult_82_n3490) );
  NAND2_X1 u5_mult_82_U8360 ( .A1(u5_mult_82_ab_39__26_), .A2(
        u5_mult_82_SUMB_38__27_), .ZN(u5_mult_82_n3489) );
  NAND2_X1 u5_mult_82_U8359 ( .A1(u5_mult_82_ab_39__26_), .A2(
        u5_mult_82_CARRYB_38__26_), .ZN(u5_mult_82_n3488) );
  XOR2_X2 u5_mult_82_U8358 ( .A(u5_mult_82_n3487), .B(u5_mult_82_SUMB_39__26_), 
        .Z(u5_mult_82_SUMB_40__25_) );
  XOR2_X2 u5_mult_82_U8357 ( .A(u5_mult_82_ab_40__25_), .B(
        u5_mult_82_CARRYB_39__25_), .Z(u5_mult_82_n3487) );
  XOR2_X2 u5_mult_82_U8356 ( .A(u5_mult_82_n3486), .B(u5_mult_82_SUMB_38__27_), 
        .Z(u5_mult_82_SUMB_39__26_) );
  XOR2_X2 u5_mult_82_U8355 ( .A(u5_mult_82_ab_39__26_), .B(
        u5_mult_82_CARRYB_38__26_), .Z(u5_mult_82_n3486) );
  INV_X8 u5_mult_82_U8354 ( .A(u5_mult_82_net57161), .ZN(u5_mult_82_net64915)
         );
  NAND2_X2 u5_mult_82_U8353 ( .A1(u5_mult_82_CARRYB_15__26_), .A2(
        u5_mult_82_net86785), .ZN(u5_mult_82_n4628) );
  NOR2_X1 u5_mult_82_U8352 ( .A1(u5_mult_82_n6960), .A2(u5_mult_82_n6730), 
        .ZN(u5_mult_82_ab_39__2_) );
  NAND3_X2 u5_mult_82_U8351 ( .A1(u5_mult_82_n3483), .A2(u5_mult_82_n3484), 
        .A3(u5_mult_82_n3485), .ZN(u5_mult_82_CARRYB_39__2_) );
  NAND2_X1 u5_mult_82_U8350 ( .A1(u5_mult_82_CARRYB_38__2_), .A2(
        u5_mult_82_ab_39__2_), .ZN(u5_mult_82_n3485) );
  NAND2_X2 u5_mult_82_U8349 ( .A1(u5_mult_82_ab_39__2_), .A2(
        u5_mult_82_SUMB_38__3_), .ZN(u5_mult_82_n3484) );
  INV_X4 u5_mult_82_U8348 ( .A(u5_mult_82_n4623), .ZN(u5_mult_82_n3480) );
  NAND2_X2 u5_mult_82_U8347 ( .A1(u5_mult_82_n3480), .A2(u5_mult_82_n728), 
        .ZN(u5_mult_82_n3482) );
  NAND2_X2 u5_mult_82_U8346 ( .A1(u5_mult_82_n4623), .A2(
        u5_mult_82_SUMB_41__3_), .ZN(u5_mult_82_n3481) );
  NAND3_X2 u5_mult_82_U8345 ( .A1(u5_mult_82_n3477), .A2(u5_mult_82_n3478), 
        .A3(u5_mult_82_n3479), .ZN(u5_mult_82_CARRYB_17__18_) );
  NAND2_X1 u5_mult_82_U8344 ( .A1(u5_mult_82_CARRYB_16__18_), .A2(
        u5_mult_82_SUMB_16__19_), .ZN(u5_mult_82_n3479) );
  NAND2_X1 u5_mult_82_U8343 ( .A1(u5_mult_82_ab_17__18_), .A2(
        u5_mult_82_SUMB_16__19_), .ZN(u5_mult_82_n3478) );
  NAND2_X1 u5_mult_82_U8342 ( .A1(u5_mult_82_ab_17__18_), .A2(
        u5_mult_82_CARRYB_16__18_), .ZN(u5_mult_82_n3477) );
  NAND2_X2 u5_mult_82_U8341 ( .A1(u5_mult_82_CARRYB_15__19_), .A2(
        u5_mult_82_n1829), .ZN(u5_mult_82_n3476) );
  NAND2_X2 u5_mult_82_U8340 ( .A1(u5_mult_82_ab_16__19_), .A2(u5_mult_82_n1829), .ZN(u5_mult_82_n3475) );
  NAND2_X1 u5_mult_82_U8339 ( .A1(u5_mult_82_ab_16__19_), .A2(
        u5_mult_82_CARRYB_15__19_), .ZN(u5_mult_82_n3474) );
  XOR2_X2 u5_mult_82_U8338 ( .A(u5_mult_82_n3473), .B(u5_mult_82_SUMB_16__19_), 
        .Z(u5_mult_82_SUMB_17__18_) );
  INV_X4 u5_mult_82_U8337 ( .A(u5_mult_82_n3471), .ZN(u5_mult_82_n3472) );
  INV_X2 u5_mult_82_U8336 ( .A(u5_mult_82_SUMB_38__36_), .ZN(u5_mult_82_n3471)
         );
  NAND2_X2 u5_mult_82_U8335 ( .A1(u5_mult_82_ab_50__21_), .A2(u5_mult_82_n1669), .ZN(u5_mult_82_n5069) );
  XNOR2_X2 u5_mult_82_U8334 ( .A(u5_mult_82_ab_38__28_), .B(
        u5_mult_82_CARRYB_37__28_), .ZN(u5_mult_82_n3470) );
  XNOR2_X2 u5_mult_82_U8333 ( .A(u5_mult_82_n3470), .B(u5_mult_82_SUMB_37__29_), .ZN(u5_mult_82_SUMB_38__28_) );
  NOR2_X1 u5_mult_82_U8332 ( .A1(u5_mult_82_net64937), .A2(u5_mult_82_n6714), 
        .ZN(u5_mult_82_ab_36__37_) );
  NAND3_X2 u5_mult_82_U8331 ( .A1(u5_mult_82_n3467), .A2(u5_mult_82_n3468), 
        .A3(u5_mult_82_n3469), .ZN(u5_mult_82_CARRYB_36__37_) );
  NAND2_X1 u5_mult_82_U8330 ( .A1(u5_mult_82_ab_36__37_), .A2(
        u5_mult_82_SUMB_35__38_), .ZN(u5_mult_82_n3469) );
  NAND2_X2 u5_mult_82_U8329 ( .A1(u5_mult_82_ab_36__37_), .A2(
        u5_mult_82_CARRYB_35__37_), .ZN(u5_mult_82_n3468) );
  NAND2_X1 u5_mult_82_U8328 ( .A1(u5_mult_82_SUMB_35__38_), .A2(
        u5_mult_82_CARRYB_35__37_), .ZN(u5_mult_82_n3467) );
  NOR2_X1 u5_mult_82_U8327 ( .A1(u5_mult_82_n6859), .A2(u5_mult_82_net66017), 
        .ZN(u5_mult_82_ab_6__30_) );
  NOR2_X1 u5_mult_82_U8326 ( .A1(u5_mult_82_net64689), .A2(u5_mult_82_n6587), 
        .ZN(u5_mult_82_ab_15__23_) );
  NAND2_X2 u5_mult_82_U8325 ( .A1(u5_mult_82_ab_6__30_), .A2(
        u5_mult_82_CARRYB_5__30_), .ZN(u5_mult_82_n3466) );
  XOR2_X2 u5_mult_82_U8324 ( .A(u5_mult_82_SUMB_5__31_), .B(u5_mult_82_n3463), 
        .Z(u5_mult_82_SUMB_6__30_) );
  XOR2_X2 u5_mult_82_U8323 ( .A(u5_mult_82_CARRYB_5__30_), .B(
        u5_mult_82_ab_6__30_), .Z(u5_mult_82_n3463) );
  NAND3_X2 u5_mult_82_U8322 ( .A1(u5_mult_82_n3460), .A2(u5_mult_82_n3461), 
        .A3(u5_mult_82_n3462), .ZN(u5_mult_82_CARRYB_15__23_) );
  NAND2_X2 u5_mult_82_U8321 ( .A1(u5_mult_82_ab_15__23_), .A2(
        u5_mult_82_CARRYB_14__23_), .ZN(u5_mult_82_n3462) );
  NAND2_X1 u5_mult_82_U8320 ( .A1(u5_mult_82_CARRYB_14__23_), .A2(
        u5_mult_82_SUMB_14__24_), .ZN(u5_mult_82_n3460) );
  XOR2_X2 u5_mult_82_U8319 ( .A(u5_mult_82_SUMB_14__24_), .B(u5_mult_82_n3459), 
        .Z(u5_mult_82_SUMB_15__23_) );
  NAND3_X2 u5_mult_82_U8318 ( .A1(u5_mult_82_n3456), .A2(u5_mult_82_n3457), 
        .A3(u5_mult_82_n3458), .ZN(u5_mult_82_CARRYB_8__29_) );
  NAND2_X2 u5_mult_82_U8317 ( .A1(u5_mult_82_CARRYB_7__29_), .A2(
        u5_mult_82_SUMB_7__30_), .ZN(u5_mult_82_n3458) );
  NAND2_X2 u5_mult_82_U8316 ( .A1(u5_mult_82_ab_8__29_), .A2(
        u5_mult_82_SUMB_7__30_), .ZN(u5_mult_82_n3457) );
  NAND2_X1 u5_mult_82_U8315 ( .A1(u5_mult_82_ab_8__29_), .A2(
        u5_mult_82_CARRYB_7__29_), .ZN(u5_mult_82_n3456) );
  NAND3_X2 u5_mult_82_U8314 ( .A1(u5_mult_82_n3453), .A2(u5_mult_82_n3454), 
        .A3(u5_mult_82_n3455), .ZN(u5_mult_82_CARRYB_7__30_) );
  NAND2_X2 u5_mult_82_U8313 ( .A1(u5_mult_82_CARRYB_6__30_), .A2(
        u5_mult_82_n1534), .ZN(u5_mult_82_n3455) );
  NAND2_X2 u5_mult_82_U8312 ( .A1(u5_mult_82_ab_7__30_), .A2(u5_mult_82_n1534), 
        .ZN(u5_mult_82_n3454) );
  NAND2_X2 u5_mult_82_U8311 ( .A1(u5_mult_82_ab_7__30_), .A2(
        u5_mult_82_CARRYB_6__30_), .ZN(u5_mult_82_n3453) );
  XOR2_X2 u5_mult_82_U8310 ( .A(u5_mult_82_n3452), .B(u5_mult_82_SUMB_7__30_), 
        .Z(u5_mult_82_SUMB_8__29_) );
  XOR2_X2 u5_mult_82_U8309 ( .A(u5_mult_82_ab_8__29_), .B(
        u5_mult_82_CARRYB_7__29_), .Z(u5_mult_82_n3452) );
  NAND3_X4 u5_mult_82_U8308 ( .A1(u5_mult_82_n3449), .A2(u5_mult_82_n3450), 
        .A3(u5_mult_82_n3451), .ZN(u5_mult_82_CARRYB_10__27_) );
  NAND2_X1 u5_mult_82_U8307 ( .A1(u5_mult_82_ab_10__27_), .A2(u5_mult_82_n1390), .ZN(u5_mult_82_n3449) );
  NAND2_X2 u5_mult_82_U8306 ( .A1(u5_mult_82_ab_9__28_), .A2(
        u5_mult_82_SUMB_8__29_), .ZN(u5_mult_82_n3447) );
  XOR2_X2 u5_mult_82_U8305 ( .A(u5_mult_82_n3445), .B(u5_mult_82_SUMB_9__28_), 
        .Z(u5_mult_82_SUMB_10__27_) );
  XOR2_X2 u5_mult_82_U8304 ( .A(u5_mult_82_n3444), .B(u5_mult_82_SUMB_8__29_), 
        .Z(u5_mult_82_SUMB_9__28_) );
  XOR2_X2 u5_mult_82_U8303 ( .A(u5_mult_82_ab_9__28_), .B(
        u5_mult_82_CARRYB_8__28_), .Z(u5_mult_82_n3444) );
  NAND2_X1 u5_mult_82_U8302 ( .A1(u5_mult_82_CARRYB_27__23_), .A2(
        u5_mult_82_SUMB_27__24_), .ZN(u5_mult_82_n5540) );
  XOR2_X2 u5_mult_82_U8301 ( .A(u5_mult_82_CARRYB_19__37_), .B(
        u5_mult_82_ab_20__37_), .Z(u5_mult_82_n5783) );
  NAND3_X4 u5_mult_82_U8300 ( .A1(u5_mult_82_n4090), .A2(u5_mult_82_n4091), 
        .A3(u5_mult_82_n4092), .ZN(u5_mult_82_CARRYB_41__27_) );
  XNOR2_X2 u5_mult_82_U8299 ( .A(u5_mult_82_ab_30__30_), .B(
        u5_mult_82_CARRYB_29__30_), .ZN(u5_mult_82_n3443) );
  XNOR2_X2 u5_mult_82_U8298 ( .A(u5_mult_82_n3442), .B(
        u5_mult_82_CARRYB_13__40_), .ZN(u5_mult_82_n5384) );
  XNOR2_X2 u5_mult_82_U8297 ( .A(u5_mult_82_CARRYB_4__50_), .B(
        u5_mult_82_ab_5__50_), .ZN(u5_mult_82_n3441) );
  XNOR2_X2 u5_mult_82_U8296 ( .A(u5_mult_82_SUMB_4__51_), .B(u5_mult_82_n3441), 
        .ZN(u5_mult_82_SUMB_5__50_) );
  NAND2_X2 u5_mult_82_U8295 ( .A1(u5_mult_82_n421), .A2(
        u5_mult_82_SUMB_14__39_), .ZN(u5_mult_82_n5357) );
  NAND3_X4 u5_mult_82_U8294 ( .A1(u5_mult_82_n5355), .A2(u5_mult_82_n5356), 
        .A3(u5_mult_82_n5357), .ZN(u5_mult_82_CARRYB_15__38_) );
  NOR2_X1 u5_mult_82_U8293 ( .A1(u5_mult_82_n6967), .A2(u5_mult_82_net65321), 
        .ZN(u5_mult_82_ab_45__1_) );
  NOR2_X1 u5_mult_82_U8292 ( .A1(u5_mult_82_n6953), .A2(u5_mult_82_net65447), 
        .ZN(u5_mult_82_ab_38__3_) );
  NOR2_X1 u5_mult_82_U8291 ( .A1(u5_mult_82_n6986), .A2(u5_mult_82_net65229), 
        .ZN(u5_mult_82_ab_50__0_) );
  NAND2_X2 u5_mult_82_U8290 ( .A1(u5_mult_82_ab_15__14_), .A2(
        u5_mult_82_CARRYB_14__14_), .ZN(u5_mult_82_n3552) );
  NOR2_X2 u5_mult_82_U8289 ( .A1(u5_mult_82_net64527), .A2(u5_mult_82_n6580), 
        .ZN(u5_mult_82_ab_14__14_) );
  NAND3_X2 u5_mult_82_U8288 ( .A1(u5_mult_82_n3438), .A2(u5_mult_82_n3439), 
        .A3(u5_mult_82_n3440), .ZN(u5_mult_82_CARRYB_45__1_) );
  NAND2_X1 u5_mult_82_U8287 ( .A1(u5_mult_82_ab_45__1_), .A2(
        u5_mult_82_SUMB_44__2_), .ZN(u5_mult_82_n3440) );
  NAND2_X2 u5_mult_82_U8286 ( .A1(u5_mult_82_CARRYB_44__1_), .A2(
        u5_mult_82_ab_45__1_), .ZN(u5_mult_82_n3439) );
  NAND2_X2 u5_mult_82_U8285 ( .A1(u5_mult_82_ab_25__9_), .A2(
        u5_mult_82_CARRYB_24__9_), .ZN(u5_mult_82_n3436) );
  XOR2_X2 u5_mult_82_U8284 ( .A(u5_mult_82_n3434), .B(u5_mult_82_CARRYB_24__9_), .Z(u5_mult_82_SUMB_25__9_) );
  NAND3_X2 u5_mult_82_U8283 ( .A1(u5_mult_82_n3431), .A2(u5_mult_82_n3432), 
        .A3(u5_mult_82_n3433), .ZN(u5_mult_82_CARRYB_24__9_) );
  NAND2_X1 u5_mult_82_U8282 ( .A1(u5_mult_82_CARRYB_23__9_), .A2(
        u5_mult_82_SUMB_23__10_), .ZN(u5_mult_82_n3433) );
  NAND3_X2 u5_mult_82_U8281 ( .A1(u5_mult_82_n3428), .A2(u5_mult_82_n3429), 
        .A3(u5_mult_82_n3430), .ZN(u5_mult_82_CARRYB_38__3_) );
  NAND2_X1 u5_mult_82_U8280 ( .A1(u5_mult_82_ab_38__3_), .A2(
        u5_mult_82_SUMB_37__4_), .ZN(u5_mult_82_n3429) );
  NAND2_X1 u5_mult_82_U8279 ( .A1(u5_mult_82_CARRYB_37__3_), .A2(
        u5_mult_82_SUMB_37__4_), .ZN(u5_mult_82_n3428) );
  XOR2_X2 u5_mult_82_U8278 ( .A(u5_mult_82_SUMB_37__4_), .B(u5_mult_82_n3427), 
        .Z(u5_mult_82_SUMB_38__3_) );
  NAND3_X2 u5_mult_82_U8277 ( .A1(u5_mult_82_n3424), .A2(u5_mult_82_n3425), 
        .A3(u5_mult_82_n3426), .ZN(u5_mult_82_CARRYB_50__0_) );
  NAND2_X1 u5_mult_82_U8276 ( .A1(u5_mult_82_ab_50__0_), .A2(
        u5_mult_82_SUMB_49__1_), .ZN(u5_mult_82_n3426) );
  NAND2_X2 u5_mult_82_U8275 ( .A1(u5_mult_82_CARRYB_49__0_), .A2(
        u5_mult_82_ab_50__0_), .ZN(u5_mult_82_n3425) );
  XOR2_X2 u5_mult_82_U8274 ( .A(u5_mult_82_SUMB_49__1_), .B(
        u5_mult_82_ab_50__0_), .Z(u5_mult_82_n3423) );
  NAND2_X1 u5_mult_82_U8273 ( .A1(u5_mult_82_ab_14__14_), .A2(
        u5_mult_82_CARRYB_13__14_), .ZN(u5_mult_82_n3422) );
  NAND2_X1 u5_mult_82_U8272 ( .A1(u5_mult_82_ab_14__14_), .A2(
        u5_mult_82_SUMB_13__15_), .ZN(u5_mult_82_n3421) );
  NAND2_X1 u5_mult_82_U8271 ( .A1(u5_mult_82_CARRYB_13__14_), .A2(
        u5_mult_82_SUMB_13__15_), .ZN(u5_mult_82_n3420) );
  XOR2_X2 u5_mult_82_U8270 ( .A(u5_mult_82_SUMB_13__15_), .B(u5_mult_82_n3419), 
        .Z(u5_mult_82_SUMB_14__14_) );
  XOR2_X2 u5_mult_82_U8269 ( .A(u5_mult_82_CARRYB_13__14_), .B(
        u5_mult_82_ab_14__14_), .Z(u5_mult_82_n3419) );
  NAND3_X2 u5_mult_82_U8268 ( .A1(u5_mult_82_n3416), .A2(u5_mult_82_n3417), 
        .A3(u5_mult_82_n3418), .ZN(u5_mult_82_CARRYB_11__17_) );
  NAND2_X1 u5_mult_82_U8267 ( .A1(u5_mult_82_CARRYB_10__17_), .A2(
        u5_mult_82_SUMB_10__18_), .ZN(u5_mult_82_n3418) );
  NAND2_X1 u5_mult_82_U8266 ( .A1(u5_mult_82_ab_11__17_), .A2(
        u5_mult_82_SUMB_10__18_), .ZN(u5_mult_82_n3417) );
  NAND2_X1 u5_mult_82_U8265 ( .A1(u5_mult_82_ab_11__17_), .A2(
        u5_mult_82_CARRYB_10__17_), .ZN(u5_mult_82_n3416) );
  NAND3_X2 u5_mult_82_U8264 ( .A1(u5_mult_82_n3413), .A2(u5_mult_82_n3414), 
        .A3(u5_mult_82_n3415), .ZN(u5_mult_82_CARRYB_10__18_) );
  NAND2_X2 u5_mult_82_U8263 ( .A1(u5_mult_82_CARRYB_9__18_), .A2(
        u5_mult_82_SUMB_9__19_), .ZN(u5_mult_82_n3415) );
  NAND2_X2 u5_mult_82_U8262 ( .A1(u5_mult_82_ab_10__18_), .A2(
        u5_mult_82_SUMB_9__19_), .ZN(u5_mult_82_n3414) );
  NAND2_X1 u5_mult_82_U8261 ( .A1(u5_mult_82_ab_10__18_), .A2(
        u5_mult_82_CARRYB_9__18_), .ZN(u5_mult_82_n3413) );
  XOR2_X2 u5_mult_82_U8260 ( .A(u5_mult_82_n3412), .B(u5_mult_82_SUMB_10__18_), 
        .Z(u5_mult_82_SUMB_11__17_) );
  XOR2_X2 u5_mult_82_U8259 ( .A(u5_mult_82_ab_11__17_), .B(
        u5_mult_82_CARRYB_10__17_), .Z(u5_mult_82_n3412) );
  XOR2_X2 u5_mult_82_U8258 ( .A(u5_mult_82_n3411), .B(u5_mult_82_SUMB_9__19_), 
        .Z(u5_mult_82_SUMB_10__18_) );
  XOR2_X2 u5_mult_82_U8257 ( .A(u5_mult_82_ab_10__18_), .B(
        u5_mult_82_CARRYB_9__18_), .Z(u5_mult_82_n3411) );
  NAND3_X2 u5_mult_82_U8256 ( .A1(u5_mult_82_n3408), .A2(u5_mult_82_n3409), 
        .A3(u5_mult_82_n3410), .ZN(u5_mult_82_CARRYB_27__7_) );
  NAND2_X1 u5_mult_82_U8255 ( .A1(u5_mult_82_ab_27__7_), .A2(
        u5_mult_82_SUMB_26__8_), .ZN(u5_mult_82_n3410) );
  NAND2_X1 u5_mult_82_U8254 ( .A1(u5_mult_82_CARRYB_26__7_), .A2(
        u5_mult_82_SUMB_26__8_), .ZN(u5_mult_82_n3409) );
  NAND2_X1 u5_mult_82_U8253 ( .A1(u5_mult_82_CARRYB_26__7_), .A2(
        u5_mult_82_ab_27__7_), .ZN(u5_mult_82_n3408) );
  NAND3_X4 u5_mult_82_U8252 ( .A1(u5_mult_82_n3405), .A2(u5_mult_82_n3406), 
        .A3(u5_mult_82_n3407), .ZN(u5_mult_82_CARRYB_26__8_) );
  NAND2_X2 u5_mult_82_U8251 ( .A1(u5_mult_82_n1435), .A2(
        u5_mult_82_SUMB_25__9_), .ZN(u5_mult_82_n3407) );
  NAND2_X2 u5_mult_82_U8250 ( .A1(u5_mult_82_ab_26__8_), .A2(
        u5_mult_82_SUMB_25__9_), .ZN(u5_mult_82_n3406) );
  NAND2_X2 u5_mult_82_U8249 ( .A1(u5_mult_82_ab_26__8_), .A2(u5_mult_82_n1435), 
        .ZN(u5_mult_82_n3405) );
  XOR2_X2 u5_mult_82_U8248 ( .A(u5_mult_82_CARRYB_26__7_), .B(
        u5_mult_82_ab_27__7_), .Z(u5_mult_82_n3404) );
  XOR2_X2 u5_mult_82_U8247 ( .A(u5_mult_82_n3403), .B(u5_mult_82_SUMB_25__9_), 
        .Z(u5_mult_82_SUMB_26__8_) );
  XOR2_X2 u5_mult_82_U8246 ( .A(u5_mult_82_ab_26__8_), .B(
        u5_mult_82_CARRYB_25__8_), .Z(u5_mult_82_n3403) );
  NAND2_X1 u5_mult_82_U8245 ( .A1(u5_mult_82_n483), .A2(u5_mult_82_ab_36__15_), 
        .ZN(u5_mult_82_n6138) );
  NAND2_X2 u5_mult_82_U8244 ( .A1(u5_mult_82_ab_12__41_), .A2(
        u5_mult_82_SUMB_11__42_), .ZN(u5_mult_82_n5369) );
  NAND2_X1 u5_mult_82_U8243 ( .A1(u5_mult_82_ab_11__37_), .A2(
        u5_mult_82_CARRYB_10__37_), .ZN(u5_mult_82_n5456) );
  NAND2_X2 u5_mult_82_U8242 ( .A1(u5_mult_82_ab_43__14_), .A2(
        u5_mult_82_SUMB_42__15_), .ZN(u5_mult_82_n6362) );
  NAND2_X2 u5_mult_82_U8241 ( .A1(u5_mult_82_CARRYB_4__49_), .A2(
        u5_mult_82_SUMB_4__50_), .ZN(u5_mult_82_n6347) );
  XOR2_X1 u5_mult_82_U8240 ( .A(u5_mult_82_n3580), .B(
        u5_mult_82_CARRYB_33__15_), .Z(u5_mult_82_n3402) );
  XNOR2_X2 u5_mult_82_U8239 ( .A(u5_mult_82_n3402), .B(u5_mult_82_SUMB_33__16_), .ZN(u5_mult_82_SUMB_34__15_) );
  XNOR2_X2 u5_mult_82_U8238 ( .A(u5_mult_82_net83655), .B(
        u5_mult_82_SUMB_38__15_), .ZN(u5_mult_82_SUMB_39__14_) );
  NAND3_X4 u5_mult_82_U8237 ( .A1(u5_mult_82_n5904), .A2(u5_mult_82_n5905), 
        .A3(u5_mult_82_n5906), .ZN(u5_mult_82_CARRYB_10__37_) );
  NOR2_X1 u5_mult_82_U8236 ( .A1(u5_mult_82_n6829), .A2(u5_mult_82_n6559), 
        .ZN(u5_mult_82_ab_11__40_) );
  NAND2_X1 u5_mult_82_U8235 ( .A1(u5_mult_82_ab_11__40_), .A2(
        u5_mult_82_SUMB_10__41_), .ZN(u5_mult_82_n3401) );
  NAND2_X2 u5_mult_82_U8234 ( .A1(u5_mult_82_ab_11__40_), .A2(
        u5_mult_82_CARRYB_10__40_), .ZN(u5_mult_82_n3400) );
  NAND3_X2 u5_mult_82_U8233 ( .A1(u5_mult_82_n3396), .A2(u5_mult_82_n3397), 
        .A3(u5_mult_82_n3398), .ZN(u5_mult_82_CARRYB_18__37_) );
  NAND2_X1 u5_mult_82_U8232 ( .A1(u5_mult_82_CARRYB_17__37_), .A2(
        u5_mult_82_SUMB_17__38_), .ZN(u5_mult_82_n3398) );
  NAND2_X1 u5_mult_82_U8231 ( .A1(u5_mult_82_ab_18__37_), .A2(
        u5_mult_82_SUMB_17__38_), .ZN(u5_mult_82_n3397) );
  NAND2_X1 u5_mult_82_U8230 ( .A1(u5_mult_82_ab_18__37_), .A2(u5_mult_82_n350), 
        .ZN(u5_mult_82_n3396) );
  NAND3_X4 u5_mult_82_U8229 ( .A1(u5_mult_82_n3393), .A2(u5_mult_82_n3394), 
        .A3(u5_mult_82_n3395), .ZN(u5_mult_82_CARRYB_17__38_) );
  NAND2_X2 u5_mult_82_U8228 ( .A1(u5_mult_82_CARRYB_16__38_), .A2(
        u5_mult_82_n76), .ZN(u5_mult_82_n3395) );
  NAND2_X2 u5_mult_82_U8227 ( .A1(u5_mult_82_ab_17__38_), .A2(u5_mult_82_n76), 
        .ZN(u5_mult_82_n3394) );
  NAND2_X1 u5_mult_82_U8226 ( .A1(u5_mult_82_ab_17__38_), .A2(
        u5_mult_82_CARRYB_16__38_), .ZN(u5_mult_82_n3393) );
  XOR2_X2 u5_mult_82_U8225 ( .A(u5_mult_82_n3392), .B(u5_mult_82_SUMB_17__38_), 
        .Z(u5_mult_82_SUMB_18__37_) );
  XOR2_X2 u5_mult_82_U8224 ( .A(u5_mult_82_n3391), .B(u5_mult_82_n76), .Z(
        u5_mult_82_SUMB_17__38_) );
  XOR2_X2 u5_mult_82_U8223 ( .A(u5_mult_82_ab_17__38_), .B(
        u5_mult_82_CARRYB_16__38_), .Z(u5_mult_82_n3391) );
  NAND2_X2 u5_mult_82_U8222 ( .A1(u5_mult_82_ab_34__25_), .A2(
        u5_mult_82_SUMB_33__26_), .ZN(u5_mult_82_n3389) );
  NAND2_X1 u5_mult_82_U8221 ( .A1(u5_mult_82_ab_34__25_), .A2(
        u5_mult_82_CARRYB_33__25_), .ZN(u5_mult_82_n3388) );
  NAND2_X2 u5_mult_82_U8220 ( .A1(u5_mult_82_SUMB_32__27_), .A2(
        u5_mult_82_CARRYB_32__26_), .ZN(u5_mult_82_n3387) );
  NAND2_X2 u5_mult_82_U8219 ( .A1(u5_mult_82_ab_33__26_), .A2(
        u5_mult_82_SUMB_32__27_), .ZN(u5_mult_82_n3386) );
  XOR2_X2 u5_mult_82_U8218 ( .A(u5_mult_82_n3384), .B(u5_mult_82_SUMB_33__26_), 
        .Z(u5_mult_82_SUMB_34__25_) );
  XOR2_X2 u5_mult_82_U8217 ( .A(u5_mult_82_ab_34__25_), .B(
        u5_mult_82_CARRYB_33__25_), .Z(u5_mult_82_n3384) );
  NAND2_X4 u5_mult_82_U8216 ( .A1(u5_mult_82_n3383), .A2(u5_mult_82_n3382), 
        .ZN(u5_mult_82_n6223) );
  XNOR2_X2 u5_mult_82_U8215 ( .A(u5_mult_82_ab_27__25_), .B(
        u5_mult_82_CARRYB_26__25_), .ZN(u5_mult_82_n3380) );
  XNOR2_X2 u5_mult_82_U8214 ( .A(u5_mult_82_n3380), .B(u5_mult_82_SUMB_26__26_), .ZN(u5_mult_82_SUMB_27__25_) );
  NAND3_X4 u5_mult_82_U8213 ( .A1(u5_mult_82_n4890), .A2(u5_mult_82_n4891), 
        .A3(u5_mult_82_n4892), .ZN(u5_mult_82_CARRYB_12__46_) );
  NAND2_X2 u5_mult_82_U8212 ( .A1(u5_mult_82_ab_32__13_), .A2(
        u5_mult_82_SUMB_31__14_), .ZN(u5_mult_82_n4764) );
  NAND2_X2 u5_mult_82_U8211 ( .A1(u5_mult_82_CARRYB_46__5_), .A2(
        u5_mult_82_SUMB_46__6_), .ZN(u5_mult_82_n6171) );
  NAND2_X2 u5_mult_82_U8210 ( .A1(u5_mult_82_ab_15__48_), .A2(
        u5_mult_82_CARRYB_14__48_), .ZN(u5_mult_82_n4326) );
  NOR2_X2 u5_mult_82_U8209 ( .A1(u5_mult_82_n6780), .A2(u5_mult_82_n6580), 
        .ZN(u5_mult_82_ab_14__48_) );
  NOR2_X1 u5_mult_82_U8208 ( .A1(u5_mult_82_n6798), .A2(u5_mult_82_n6644), 
        .ZN(u5_mult_82_ab_24__45_) );
  NOR2_X1 u5_mult_82_U8207 ( .A1(u5_mult_82_n6831), .A2(u5_mult_82_net65405), 
        .ZN(u5_mult_82_ab_40__39_) );
  NOR2_X1 u5_mult_82_U8206 ( .A1(u5_mult_82_n6798), .A2(u5_mult_82_n6615), 
        .ZN(u5_mult_82_ab_19__45_) );
  NAND3_X2 u5_mult_82_U8205 ( .A1(u5_mult_82_n3377), .A2(u5_mult_82_n3378), 
        .A3(u5_mult_82_n3379), .ZN(u5_mult_82_CARRYB_14__48_) );
  NAND2_X1 u5_mult_82_U8204 ( .A1(u5_mult_82_ab_14__48_), .A2(
        u5_mult_82_SUMB_13__49_), .ZN(u5_mult_82_n3379) );
  NAND2_X2 u5_mult_82_U8203 ( .A1(u5_mult_82_ab_14__48_), .A2(
        u5_mult_82_CARRYB_13__48_), .ZN(u5_mult_82_n3378) );
  NAND3_X2 u5_mult_82_U8202 ( .A1(u5_mult_82_n3374), .A2(u5_mult_82_n3375), 
        .A3(u5_mult_82_n3376), .ZN(u5_mult_82_CARRYB_24__45_) );
  NAND2_X2 u5_mult_82_U8201 ( .A1(u5_mult_82_CARRYB_23__45_), .A2(
        u5_mult_82_ab_24__45_), .ZN(u5_mult_82_n3375) );
  NAND3_X2 u5_mult_82_U8200 ( .A1(u5_mult_82_n3371), .A2(u5_mult_82_n3372), 
        .A3(u5_mult_82_n3373), .ZN(u5_mult_82_CARRYB_40__39_) );
  NAND2_X2 u5_mult_82_U8199 ( .A1(u5_mult_82_ab_40__39_), .A2(
        u5_mult_82_SUMB_39__40_), .ZN(u5_mult_82_n3372) );
  XOR2_X2 u5_mult_82_U8198 ( .A(u5_mult_82_SUMB_39__40_), .B(u5_mult_82_n3370), 
        .Z(u5_mult_82_SUMB_40__39_) );
  XOR2_X2 u5_mult_82_U8197 ( .A(u5_mult_82_CARRYB_39__39_), .B(
        u5_mult_82_ab_40__39_), .Z(u5_mult_82_n3370) );
  NAND3_X2 u5_mult_82_U8196 ( .A1(u5_mult_82_n3367), .A2(u5_mult_82_n3368), 
        .A3(u5_mult_82_n3369), .ZN(u5_mult_82_CARRYB_19__45_) );
  NAND2_X1 u5_mult_82_U8195 ( .A1(u5_mult_82_ab_19__45_), .A2(
        u5_mult_82_CARRYB_18__45_), .ZN(u5_mult_82_n3369) );
  NAND2_X2 u5_mult_82_U8194 ( .A1(u5_mult_82_ab_19__45_), .A2(
        u5_mult_82_SUMB_18__46_), .ZN(u5_mult_82_n3368) );
  XOR2_X2 u5_mult_82_U8193 ( .A(u5_mult_82_SUMB_18__46_), .B(u5_mult_82_n3366), 
        .Z(u5_mult_82_SUMB_19__45_) );
  XOR2_X2 u5_mult_82_U8192 ( .A(u5_mult_82_CARRYB_18__45_), .B(
        u5_mult_82_ab_19__45_), .Z(u5_mult_82_n3366) );
  INV_X4 u5_mult_82_U8191 ( .A(u5_mult_82_n3969), .ZN(u5_mult_82_n3363) );
  NAND2_X4 u5_mult_82_U8190 ( .A1(u5_mult_82_n3363), .A2(u5_mult_82_n1438), 
        .ZN(u5_mult_82_n3365) );
  NAND2_X2 u5_mult_82_U8189 ( .A1(u5_mult_82_ab_5__49_), .A2(
        u5_mult_82_SUMB_4__50_), .ZN(u5_mult_82_n6346) );
  XNOR2_X2 u5_mult_82_U8188 ( .A(u5_mult_82_CARRYB_17__43_), .B(
        u5_mult_82_ab_18__43_), .ZN(u5_mult_82_n3362) );
  XNOR2_X2 u5_mult_82_U8187 ( .A(u5_mult_82_n3362), .B(u5_mult_82_SUMB_17__44_), .ZN(u5_mult_82_SUMB_18__43_) );
  NAND2_X2 u5_mult_82_U8186 ( .A1(u5_mult_82_ab_18__45_), .A2(
        u5_mult_82_SUMB_17__46_), .ZN(u5_mult_82_n5875) );
  XOR2_X1 u5_mult_82_U8185 ( .A(u5_mult_82_CARRYB_16__48_), .B(
        u5_mult_82_ab_17__48_), .Z(u5_mult_82_n4425) );
  NAND3_X4 u5_mult_82_U8184 ( .A1(u5_mult_82_n4887), .A2(u5_mult_82_n4888), 
        .A3(u5_mult_82_n4889), .ZN(u5_mult_82_CARRYB_18__43_) );
  NAND2_X2 u5_mult_82_U8183 ( .A1(u5_mult_82_CARRYB_33__13_), .A2(
        u5_mult_82_SUMB_33__14_), .ZN(u5_mult_82_n5923) );
  NAND2_X2 u5_mult_82_U8182 ( .A1(u5_mult_82_n1486), .A2(u5_mult_82_ab_41__9_), 
        .ZN(u5_mult_82_n6068) );
  XOR2_X2 u5_mult_82_U8181 ( .A(u5_mult_82_CARRYB_23__48_), .B(
        u5_mult_82_n3767), .Z(u5_mult_82_SUMB_24__48_) );
  NAND3_X2 u5_mult_82_U8180 ( .A1(u5_mult_82_n4211), .A2(u5_mult_82_n4212), 
        .A3(u5_mult_82_n4213), .ZN(u5_mult_82_CARRYB_38__20_) );
  NOR2_X1 u5_mult_82_U8179 ( .A1(u5_mult_82_n6784), .A2(u5_mult_82_n6670), 
        .ZN(u5_mult_82_ab_29__47_) );
  NOR2_X1 u5_mult_82_U8178 ( .A1(u5_mult_82_net64913), .A2(u5_mult_82_net65351), .ZN(u5_mult_82_ab_43__35_) );
  NAND3_X2 u5_mult_82_U8177 ( .A1(u5_mult_82_n3359), .A2(u5_mult_82_n3360), 
        .A3(u5_mult_82_n3361), .ZN(u5_mult_82_CARRYB_29__47_) );
  NAND2_X1 u5_mult_82_U8176 ( .A1(u5_mult_82_ab_29__47_), .A2(
        u5_mult_82_SUMB_28__48_), .ZN(u5_mult_82_n3361) );
  NAND2_X1 u5_mult_82_U8175 ( .A1(u5_mult_82_ab_29__47_), .A2(
        u5_mult_82_CARRYB_28__47_), .ZN(u5_mult_82_n3360) );
  NAND2_X1 u5_mult_82_U8174 ( .A1(u5_mult_82_SUMB_28__48_), .A2(
        u5_mult_82_CARRYB_28__47_), .ZN(u5_mult_82_n3359) );
  NAND3_X2 u5_mult_82_U8173 ( .A1(u5_mult_82_n3356), .A2(u5_mult_82_n3357), 
        .A3(u5_mult_82_n3358), .ZN(u5_mult_82_CARRYB_43__35_) );
  NAND2_X1 u5_mult_82_U8172 ( .A1(u5_mult_82_ab_43__35_), .A2(
        u5_mult_82_CARRYB_42__35_), .ZN(u5_mult_82_n3358) );
  NAND2_X2 u5_mult_82_U8171 ( .A1(u5_mult_82_ab_43__35_), .A2(
        u5_mult_82_SUMB_42__36_), .ZN(u5_mult_82_n3357) );
  NAND2_X1 u5_mult_82_U8170 ( .A1(u5_mult_82_CARRYB_42__35_), .A2(
        u5_mult_82_SUMB_42__36_), .ZN(u5_mult_82_n3356) );
  XOR2_X2 u5_mult_82_U8169 ( .A(u5_mult_82_SUMB_42__36_), .B(u5_mult_82_n3355), 
        .Z(u5_mult_82_SUMB_43__35_) );
  NAND3_X4 u5_mult_82_U8168 ( .A1(u5_mult_82_n3352), .A2(u5_mult_82_n3353), 
        .A3(u5_mult_82_n3354), .ZN(u5_mult_82_CARRYB_46__32_) );
  NAND2_X2 u5_mult_82_U8167 ( .A1(u5_mult_82_CARRYB_45__32_), .A2(
        u5_mult_82_SUMB_45__33_), .ZN(u5_mult_82_n3354) );
  NAND2_X2 u5_mult_82_U8166 ( .A1(u5_mult_82_ab_46__32_), .A2(
        u5_mult_82_SUMB_45__33_), .ZN(u5_mult_82_n3353) );
  NAND2_X1 u5_mult_82_U8165 ( .A1(u5_mult_82_ab_46__32_), .A2(
        u5_mult_82_CARRYB_45__32_), .ZN(u5_mult_82_n3352) );
  NAND3_X2 u5_mult_82_U8164 ( .A1(u5_mult_82_n3349), .A2(u5_mult_82_n3350), 
        .A3(u5_mult_82_n3351), .ZN(u5_mult_82_CARRYB_45__33_) );
  NAND2_X2 u5_mult_82_U8163 ( .A1(u5_mult_82_CARRYB_44__33_), .A2(
        u5_mult_82_SUMB_44__34_), .ZN(u5_mult_82_n3351) );
  NAND2_X2 u5_mult_82_U8162 ( .A1(u5_mult_82_ab_45__33_), .A2(
        u5_mult_82_SUMB_44__34_), .ZN(u5_mult_82_n3350) );
  NAND2_X1 u5_mult_82_U8161 ( .A1(u5_mult_82_ab_45__33_), .A2(
        u5_mult_82_CARRYB_44__33_), .ZN(u5_mult_82_n3349) );
  NAND3_X2 u5_mult_82_U8160 ( .A1(u5_mult_82_n6168), .A2(u5_mult_82_n6167), 
        .A3(u5_mult_82_n6166), .ZN(u5_mult_82_CARRYB_46__6_) );
  INV_X8 u5_mult_82_U8159 ( .A(n4756), .ZN(u5_mult_82_n7017) );
  NAND2_X2 u5_mult_82_U8158 ( .A1(u5_mult_82_CARRYB_36__15_), .A2(
        u5_mult_82_SUMB_36__16_), .ZN(u5_mult_82_n6178) );
  NOR2_X1 u5_mult_82_U8157 ( .A1(u5_mult_82_net64887), .A2(u5_mult_82_n6557), 
        .ZN(u5_mult_82_ab_11__34_) );
  NOR2_X1 u5_mult_82_U8156 ( .A1(u5_mult_82_net64887), .A2(u5_mult_82_n6544), 
        .ZN(u5_mult_82_ab_9__34_) );
  NAND3_X2 u5_mult_82_U8155 ( .A1(u5_mult_82_n3346), .A2(u5_mult_82_n3347), 
        .A3(u5_mult_82_n3348), .ZN(u5_mult_82_CARRYB_11__34_) );
  NAND2_X1 u5_mult_82_U8154 ( .A1(u5_mult_82_ab_11__34_), .A2(
        u5_mult_82_CARRYB_10__34_), .ZN(u5_mult_82_n3348) );
  NAND2_X2 u5_mult_82_U8153 ( .A1(u5_mult_82_ab_11__34_), .A2(
        u5_mult_82_SUMB_10__35_), .ZN(u5_mult_82_n3347) );
  NAND2_X1 u5_mult_82_U8152 ( .A1(u5_mult_82_CARRYB_10__34_), .A2(
        u5_mult_82_SUMB_10__35_), .ZN(u5_mult_82_n3346) );
  XOR2_X2 u5_mult_82_U8151 ( .A(u5_mult_82_SUMB_10__35_), .B(u5_mult_82_n3345), 
        .Z(u5_mult_82_SUMB_11__34_) );
  XOR2_X2 u5_mult_82_U8150 ( .A(u5_mult_82_CARRYB_10__34_), .B(
        u5_mult_82_ab_11__34_), .Z(u5_mult_82_n3345) );
  NAND3_X2 u5_mult_82_U8149 ( .A1(u5_mult_82_n3342), .A2(u5_mult_82_n3343), 
        .A3(u5_mult_82_n3344), .ZN(u5_mult_82_CARRYB_9__34_) );
  NAND2_X2 u5_mult_82_U8148 ( .A1(u5_mult_82_ab_9__34_), .A2(
        u5_mult_82_CARRYB_8__34_), .ZN(u5_mult_82_n3344) );
  NAND2_X1 u5_mult_82_U8147 ( .A1(u5_mult_82_ab_9__34_), .A2(
        u5_mult_82_SUMB_8__35_), .ZN(u5_mult_82_n3343) );
  NAND2_X1 u5_mult_82_U8146 ( .A1(u5_mult_82_CARRYB_8__34_), .A2(
        u5_mult_82_SUMB_8__35_), .ZN(u5_mult_82_n3342) );
  XOR2_X2 u5_mult_82_U8145 ( .A(u5_mult_82_SUMB_8__35_), .B(u5_mult_82_n3341), 
        .Z(u5_mult_82_SUMB_9__34_) );
  XOR2_X2 u5_mult_82_U8144 ( .A(u5_mult_82_CARRYB_8__34_), .B(
        u5_mult_82_ab_9__34_), .Z(u5_mult_82_n3341) );
  NAND3_X2 u5_mult_82_U8143 ( .A1(u5_mult_82_n3338), .A2(u5_mult_82_n3339), 
        .A3(u5_mult_82_n3340), .ZN(u5_mult_82_CARRYB_21__28_) );
  NAND2_X1 u5_mult_82_U8142 ( .A1(u5_mult_82_CARRYB_20__28_), .A2(
        u5_mult_82_SUMB_20__29_), .ZN(u5_mult_82_n3340) );
  NAND2_X1 u5_mult_82_U8141 ( .A1(u5_mult_82_ab_21__28_), .A2(
        u5_mult_82_SUMB_20__29_), .ZN(u5_mult_82_n3339) );
  NAND2_X1 u5_mult_82_U8140 ( .A1(u5_mult_82_ab_21__28_), .A2(
        u5_mult_82_CARRYB_20__28_), .ZN(u5_mult_82_n3338) );
  NAND3_X4 u5_mult_82_U8139 ( .A1(u5_mult_82_n3335), .A2(u5_mult_82_n3336), 
        .A3(u5_mult_82_n3337), .ZN(u5_mult_82_CARRYB_20__29_) );
  NAND2_X2 u5_mult_82_U8138 ( .A1(u5_mult_82_CARRYB_19__29_), .A2(
        u5_mult_82_SUMB_19__30_), .ZN(u5_mult_82_n3337) );
  NAND2_X2 u5_mult_82_U8137 ( .A1(u5_mult_82_ab_20__29_), .A2(
        u5_mult_82_SUMB_19__30_), .ZN(u5_mult_82_n3336) );
  NAND2_X1 u5_mult_82_U8136 ( .A1(u5_mult_82_ab_20__29_), .A2(
        u5_mult_82_CARRYB_19__29_), .ZN(u5_mult_82_n3335) );
  XOR2_X2 u5_mult_82_U8135 ( .A(u5_mult_82_n3334), .B(u5_mult_82_SUMB_20__29_), 
        .Z(u5_mult_82_SUMB_21__28_) );
  XOR2_X2 u5_mult_82_U8134 ( .A(u5_mult_82_n3333), .B(u5_mult_82_n1760), .Z(
        u5_mult_82_SUMB_20__29_) );
  XOR2_X2 u5_mult_82_U8133 ( .A(u5_mult_82_ab_20__29_), .B(
        u5_mult_82_CARRYB_19__29_), .Z(u5_mult_82_n3333) );
  NAND2_X2 u5_mult_82_U8132 ( .A1(u5_mult_82_ab_17__24_), .A2(
        u5_mult_82_CARRYB_16__24_), .ZN(u5_mult_82_n5322) );
  NOR2_X2 u5_mult_82_U8131 ( .A1(u5_mult_82_n6892), .A2(u5_mult_82_n6595), 
        .ZN(u5_mult_82_ab_16__24_) );
  NOR2_X1 u5_mult_82_U8130 ( .A1(u5_mult_82_n6864), .A2(u5_mult_82_n6550), 
        .ZN(u5_mult_82_ab_10__29_) );
  NAND2_X2 u5_mult_82_U8129 ( .A1(u5_mult_82_ab_16__24_), .A2(
        u5_mult_82_CARRYB_15__24_), .ZN(u5_mult_82_n3332) );
  NAND3_X2 u5_mult_82_U8128 ( .A1(u5_mult_82_n3327), .A2(u5_mult_82_n3328), 
        .A3(u5_mult_82_n3329), .ZN(u5_mult_82_CARRYB_10__29_) );
  NAND2_X1 u5_mult_82_U8127 ( .A1(u5_mult_82_ab_10__29_), .A2(
        u5_mult_82_CARRYB_9__29_), .ZN(u5_mult_82_n3329) );
  NAND2_X1 u5_mult_82_U8126 ( .A1(u5_mult_82_CARRYB_9__29_), .A2(
        u5_mult_82_SUMB_9__30_), .ZN(u5_mult_82_n3327) );
  XOR2_X2 u5_mult_82_U8125 ( .A(u5_mult_82_SUMB_9__30_), .B(u5_mult_82_n3326), 
        .Z(u5_mult_82_SUMB_10__29_) );
  XOR2_X2 u5_mult_82_U8124 ( .A(u5_mult_82_CARRYB_9__29_), .B(
        u5_mult_82_ab_10__29_), .Z(u5_mult_82_n3326) );
  NAND3_X2 u5_mult_82_U8123 ( .A1(u5_mult_82_n4160), .A2(u5_mult_82_n4161), 
        .A3(u5_mult_82_n4162), .ZN(u5_mult_82_CARRYB_43__20_) );
  NOR2_X1 u5_mult_82_U8122 ( .A1(u5_mult_82_net64471), .A2(u5_mult_82_n6616), 
        .ZN(u5_mult_82_ab_19__11_) );
  NAND3_X2 u5_mult_82_U8121 ( .A1(u5_mult_82_n3323), .A2(u5_mult_82_n3324), 
        .A3(u5_mult_82_n3325), .ZN(u5_mult_82_CARRYB_19__11_) );
  NAND2_X1 u5_mult_82_U8120 ( .A1(u5_mult_82_ab_19__11_), .A2(
        u5_mult_82_CARRYB_18__11_), .ZN(u5_mult_82_n3325) );
  NAND2_X2 u5_mult_82_U8119 ( .A1(u5_mult_82_ab_19__11_), .A2(
        u5_mult_82_SUMB_18__12_), .ZN(u5_mult_82_n3324) );
  NAND2_X1 u5_mult_82_U8118 ( .A1(u5_mult_82_CARRYB_18__11_), .A2(
        u5_mult_82_SUMB_18__12_), .ZN(u5_mult_82_n3323) );
  NAND3_X2 u5_mult_82_U8117 ( .A1(u5_mult_82_n3319), .A2(u5_mult_82_n3320), 
        .A3(u5_mult_82_n3321), .ZN(u5_mult_82_CARRYB_12__18_) );
  NAND2_X1 u5_mult_82_U8116 ( .A1(u5_mult_82_SUMB_11__19_), .A2(
        u5_mult_82_CARRYB_11__18_), .ZN(u5_mult_82_n3321) );
  NAND2_X1 u5_mult_82_U8115 ( .A1(u5_mult_82_ab_12__18_), .A2(
        u5_mult_82_SUMB_11__19_), .ZN(u5_mult_82_n3320) );
  NAND2_X1 u5_mult_82_U8114 ( .A1(u5_mult_82_ab_12__18_), .A2(
        u5_mult_82_CARRYB_11__18_), .ZN(u5_mult_82_n3319) );
  NAND3_X2 u5_mult_82_U8113 ( .A1(u5_mult_82_n3316), .A2(u5_mult_82_n3317), 
        .A3(u5_mult_82_n3318), .ZN(u5_mult_82_CARRYB_11__19_) );
  NAND2_X1 u5_mult_82_U8112 ( .A1(u5_mult_82_CARRYB_10__19_), .A2(
        u5_mult_82_SUMB_10__20_), .ZN(u5_mult_82_n3318) );
  NAND2_X1 u5_mult_82_U8111 ( .A1(u5_mult_82_ab_11__19_), .A2(
        u5_mult_82_SUMB_10__20_), .ZN(u5_mult_82_n3317) );
  NAND2_X1 u5_mult_82_U8110 ( .A1(u5_mult_82_ab_11__19_), .A2(
        u5_mult_82_CARRYB_10__19_), .ZN(u5_mult_82_n3316) );
  XOR2_X2 u5_mult_82_U8109 ( .A(u5_mult_82_n3315), .B(u5_mult_82_SUMB_11__19_), 
        .Z(u5_mult_82_SUMB_12__18_) );
  XOR2_X2 u5_mult_82_U8108 ( .A(u5_mult_82_n3314), .B(u5_mult_82_SUMB_10__20_), 
        .Z(u5_mult_82_SUMB_11__19_) );
  XOR2_X2 u5_mult_82_U8107 ( .A(u5_mult_82_ab_11__19_), .B(
        u5_mult_82_CARRYB_10__19_), .Z(u5_mult_82_n3314) );
  NAND3_X2 u5_mult_82_U8106 ( .A1(u5_mult_82_n3311), .A2(u5_mult_82_n3312), 
        .A3(u5_mult_82_n3313), .ZN(u5_mult_82_CARRYB_26__6_) );
  NAND2_X1 u5_mult_82_U8105 ( .A1(u5_mult_82_CARRYB_25__6_), .A2(
        u5_mult_82_SUMB_25__7_), .ZN(u5_mult_82_n3313) );
  NAND2_X1 u5_mult_82_U8104 ( .A1(u5_mult_82_ab_26__6_), .A2(
        u5_mult_82_SUMB_25__7_), .ZN(u5_mult_82_n3312) );
  NAND2_X1 u5_mult_82_U8103 ( .A1(u5_mult_82_ab_26__6_), .A2(
        u5_mult_82_CARRYB_25__6_), .ZN(u5_mult_82_n3311) );
  NAND3_X2 u5_mult_82_U8102 ( .A1(u5_mult_82_n3308), .A2(u5_mult_82_n3309), 
        .A3(u5_mult_82_n3310), .ZN(u5_mult_82_CARRYB_25__7_) );
  NAND2_X2 u5_mult_82_U8101 ( .A1(u5_mult_82_ab_25__7_), .A2(
        u5_mult_82_SUMB_24__8_), .ZN(u5_mult_82_n3309) );
  NAND2_X1 u5_mult_82_U8100 ( .A1(u5_mult_82_ab_25__7_), .A2(
        u5_mult_82_CARRYB_24__7_), .ZN(u5_mult_82_n3308) );
  XOR2_X2 u5_mult_82_U8099 ( .A(u5_mult_82_n3307), .B(u5_mult_82_SUMB_25__7_), 
        .Z(u5_mult_82_SUMB_26__6_) );
  XOR2_X2 u5_mult_82_U8098 ( .A(u5_mult_82_ab_26__6_), .B(
        u5_mult_82_CARRYB_25__6_), .Z(u5_mult_82_n3307) );
  XOR2_X2 u5_mult_82_U8097 ( .A(u5_mult_82_n3306), .B(u5_mult_82_SUMB_24__8_), 
        .Z(u5_mult_82_SUMB_25__7_) );
  XOR2_X2 u5_mult_82_U8096 ( .A(u5_mult_82_CARRYB_24__7_), .B(
        u5_mult_82_ab_25__7_), .Z(u5_mult_82_n3306) );
  XNOR2_X2 u5_mult_82_U8095 ( .A(u5_mult_82_ab_31__28_), .B(u5_mult_82_n1628), 
        .ZN(u5_mult_82_n3305) );
  XNOR2_X2 u5_mult_82_U8094 ( .A(u5_mult_82_n3305), .B(u5_mult_82_SUMB_30__29_), .ZN(u5_mult_82_SUMB_31__28_) );
  NAND2_X2 u5_mult_82_U8093 ( .A1(u5_mult_82_CARRYB_49__21_), .A2(
        u5_mult_82_n1669), .ZN(u5_mult_82_n5068) );
  NAND2_X2 u5_mult_82_U8092 ( .A1(u5_mult_82_n3074), .A2(
        u5_mult_82_SUMB_28__22_), .ZN(u5_mult_82_n5435) );
  NAND2_X2 u5_mult_82_U8091 ( .A1(u5_mult_82_n446), .A2(
        u5_mult_82_SUMB_20__40_), .ZN(u5_mult_82_n4946) );
  NAND3_X4 u5_mult_82_U8090 ( .A1(u5_mult_82_n4944), .A2(u5_mult_82_n4945), 
        .A3(u5_mult_82_n4946), .ZN(u5_mult_82_CARRYB_21__39_) );
  NAND3_X4 u5_mult_82_U8089 ( .A1(u5_mult_82_n6189), .A2(u5_mult_82_n6188), 
        .A3(u5_mult_82_n6187), .ZN(u5_mult_82_CARRYB_16__36_) );
  NAND2_X2 u5_mult_82_U8088 ( .A1(u5_mult_82_ab_39__25_), .A2(
        u5_mult_82_SUMB_38__26_), .ZN(u5_mult_82_n3853) );
  NAND2_X1 u5_mult_82_U8087 ( .A1(u5_mult_82_ab_28__23_), .A2(
        u5_mult_82_SUMB_27__24_), .ZN(u5_mult_82_n5539) );
  NOR2_X1 u5_mult_82_U8086 ( .A1(u5_mult_82_n6927), .A2(u5_mult_82_n6700), 
        .ZN(u5_mult_82_ab_33__17_) );
  NAND3_X2 u5_mult_82_U8085 ( .A1(u5_mult_82_n3302), .A2(u5_mult_82_n3303), 
        .A3(u5_mult_82_n3304), .ZN(u5_mult_82_CARRYB_33__17_) );
  NAND2_X2 u5_mult_82_U8084 ( .A1(u5_mult_82_ab_33__17_), .A2(
        u5_mult_82_SUMB_32__18_), .ZN(u5_mult_82_n3303) );
  NAND2_X2 u5_mult_82_U8083 ( .A1(u5_mult_82_CARRYB_17__43_), .A2(
        u5_mult_82_SUMB_17__44_), .ZN(u5_mult_82_n4889) );
  XNOR2_X2 u5_mult_82_U8082 ( .A(u5_mult_82_ab_51__21_), .B(
        u5_mult_82_CARRYB_50__21_), .ZN(u5_mult_82_n3301) );
  XNOR2_X2 u5_mult_82_U8081 ( .A(u5_mult_82_n3301), .B(u5_mult_82_SUMB_50__22_), .ZN(u5_mult_82_SUMB_51__21_) );
  XNOR2_X2 u5_mult_82_U8080 ( .A(u5_mult_82_CARRYB_41__31_), .B(
        u5_mult_82_ab_42__31_), .ZN(u5_mult_82_n3300) );
  XNOR2_X2 u5_mult_82_U8079 ( .A(u5_mult_82_n3300), .B(u5_mult_82_SUMB_41__32_), .ZN(u5_mult_82_SUMB_42__31_) );
  XOR2_X2 u5_mult_82_U8078 ( .A(u5_mult_82_ab_43__21_), .B(
        u5_mult_82_CARRYB_42__21_), .Z(u5_mult_82_n5176) );
  NAND3_X4 u5_mult_82_U8077 ( .A1(u5_mult_82_n5542), .A2(u5_mult_82_n5543), 
        .A3(u5_mult_82_n5544), .ZN(u5_mult_82_CARRYB_21__34_) );
  XNOR2_X2 u5_mult_82_U8076 ( .A(u5_mult_82_n4099), .B(u5_mult_82_SUMB_41__5_), 
        .ZN(u5_mult_82_SUMB_42__4_) );
  NAND2_X1 u5_mult_82_U8075 ( .A1(u5_mult_82_ab_3__39_), .A2(
        u5_mult_82_SUMB_2__40_), .ZN(u5_mult_82_n4174) );
  NAND2_X2 u5_mult_82_U8074 ( .A1(u5_mult_82_ab_18__43_), .A2(
        u5_mult_82_SUMB_17__44_), .ZN(u5_mult_82_n4888) );
  NAND2_X4 u5_mult_82_U8073 ( .A1(u5_mult_82_n3495), .A2(u5_mult_82_n5662), 
        .ZN(u5_mult_82_CARRYB_42__23_) );
  NAND2_X2 u5_mult_82_U8072 ( .A1(u5_mult_82_ab_18__43_), .A2(
        u5_mult_82_CARRYB_17__43_), .ZN(u5_mult_82_n4887) );
  NAND3_X2 u5_mult_82_U8071 ( .A1(u5_mult_82_n3297), .A2(u5_mult_82_n3298), 
        .A3(u5_mult_82_n3299), .ZN(u5_mult_82_CARRYB_14__44_) );
  NAND2_X2 u5_mult_82_U8070 ( .A1(u5_mult_82_CARRYB_13__44_), .A2(
        u5_mult_82_SUMB_13__45_), .ZN(u5_mult_82_n3299) );
  NAND2_X2 u5_mult_82_U8069 ( .A1(u5_mult_82_ab_14__44_), .A2(
        u5_mult_82_SUMB_13__45_), .ZN(u5_mult_82_n3298) );
  NAND2_X1 u5_mult_82_U8068 ( .A1(u5_mult_82_ab_14__44_), .A2(
        u5_mult_82_CARRYB_13__44_), .ZN(u5_mult_82_n3297) );
  NAND3_X2 u5_mult_82_U8067 ( .A1(u5_mult_82_n3294), .A2(u5_mult_82_n3295), 
        .A3(u5_mult_82_n3296), .ZN(u5_mult_82_CARRYB_13__45_) );
  NAND2_X2 u5_mult_82_U8066 ( .A1(u5_mult_82_CARRYB_12__45_), .A2(
        u5_mult_82_SUMB_12__46_), .ZN(u5_mult_82_n3296) );
  NAND2_X2 u5_mult_82_U8065 ( .A1(u5_mult_82_ab_13__45_), .A2(u5_mult_82_n1404), .ZN(u5_mult_82_n3295) );
  NAND2_X1 u5_mult_82_U8064 ( .A1(u5_mult_82_ab_13__45_), .A2(
        u5_mult_82_CARRYB_12__45_), .ZN(u5_mult_82_n3294) );
  XOR2_X2 u5_mult_82_U8063 ( .A(u5_mult_82_n3293), .B(u5_mult_82_SUMB_13__45_), 
        .Z(u5_mult_82_SUMB_14__44_) );
  XOR2_X2 u5_mult_82_U8062 ( .A(u5_mult_82_ab_14__44_), .B(
        u5_mult_82_CARRYB_13__44_), .Z(u5_mult_82_n3293) );
  NAND2_X1 u5_mult_82_U8061 ( .A1(u5_mult_82_CARRYB_5__37_), .A2(
        u5_mult_82_SUMB_5__38_), .ZN(u5_mult_82_n3292) );
  NAND2_X1 u5_mult_82_U8060 ( .A1(u5_mult_82_ab_6__37_), .A2(
        u5_mult_82_CARRYB_5__37_), .ZN(u5_mult_82_n3290) );
  NAND3_X2 u5_mult_82_U8059 ( .A1(u5_mult_82_n3287), .A2(u5_mult_82_n3288), 
        .A3(u5_mult_82_n3289), .ZN(u5_mult_82_CARRYB_5__38_) );
  NAND2_X2 u5_mult_82_U8058 ( .A1(u5_mult_82_CARRYB_4__38_), .A2(
        u5_mult_82_SUMB_4__39_), .ZN(u5_mult_82_n3289) );
  NAND2_X2 u5_mult_82_U8057 ( .A1(u5_mult_82_ab_5__38_), .A2(
        u5_mult_82_SUMB_4__39_), .ZN(u5_mult_82_n3288) );
  NAND2_X1 u5_mult_82_U8056 ( .A1(u5_mult_82_ab_5__38_), .A2(
        u5_mult_82_CARRYB_4__38_), .ZN(u5_mult_82_n3287) );
  XOR2_X2 u5_mult_82_U8055 ( .A(u5_mult_82_n3286), .B(u5_mult_82_SUMB_4__39_), 
        .Z(u5_mult_82_SUMB_5__38_) );
  XOR2_X2 u5_mult_82_U8054 ( .A(u5_mult_82_ab_5__38_), .B(
        u5_mult_82_CARRYB_4__38_), .Z(u5_mult_82_n3286) );
  INV_X4 u5_mult_82_U8053 ( .A(u5_mult_82_n2480), .ZN(u5_mult_82_n6824) );
  XNOR2_X2 u5_mult_82_U8052 ( .A(u5_mult_82_CARRYB_5__48_), .B(
        u5_mult_82_ab_6__48_), .ZN(u5_mult_82_n3285) );
  XNOR2_X2 u5_mult_82_U8051 ( .A(u5_mult_82_n3285), .B(u5_mult_82_SUMB_5__49_), 
        .ZN(u5_mult_82_SUMB_6__48_) );
  NAND2_X2 u5_mult_82_U8050 ( .A1(u5_mult_82_ab_34__13_), .A2(
        u5_mult_82_SUMB_33__14_), .ZN(u5_mult_82_n5922) );
  NAND3_X4 u5_mult_82_U8049 ( .A1(u5_mult_82_n5921), .A2(u5_mult_82_n5922), 
        .A3(u5_mult_82_n5923), .ZN(u5_mult_82_CARRYB_34__13_) );
  XNOR2_X2 u5_mult_82_U8048 ( .A(u5_mult_82_SUMB_30__17_), .B(
        u5_mult_82_ab_31__16_), .ZN(u5_mult_82_n3702) );
  XNOR2_X2 u5_mult_82_U8047 ( .A(u5_mult_82_ab_23__25_), .B(
        u5_mult_82_CARRYB_22__25_), .ZN(u5_mult_82_n3284) );
  XNOR2_X2 u5_mult_82_U8046 ( .A(u5_mult_82_n3284), .B(u5_mult_82_SUMB_22__26_), .ZN(u5_mult_82_SUMB_23__25_) );
  XNOR2_X2 u5_mult_82_U8045 ( .A(u5_mult_82_n3283), .B(
        u5_mult_82_CARRYB_24__20_), .ZN(u5_mult_82_n5689) );
  NAND2_X1 u5_mult_82_U8044 ( .A1(u5_mult_82_ab_13__46_), .A2(
        u5_mult_82_CARRYB_12__46_), .ZN(u5_mult_82_n4592) );
  NAND2_X1 u5_mult_82_U8043 ( .A1(u5_mult_82_CARRYB_12__46_), .A2(
        u5_mult_82_SUMB_12__47_), .ZN(u5_mult_82_n4594) );
  NAND2_X1 u5_mult_82_U8042 ( .A1(u5_mult_82_ab_26__20_), .A2(
        u5_mult_82_CARRYB_25__20_), .ZN(u5_mult_82_n4586) );
  NAND2_X2 u5_mult_82_U8041 ( .A1(u5_mult_82_CARRYB_5__47_), .A2(
        u5_mult_82_n1822), .ZN(u5_mult_82_n6321) );
  NAND3_X4 u5_mult_82_U8040 ( .A1(u5_mult_82_n5899), .A2(u5_mult_82_n5900), 
        .A3(u5_mult_82_n5901), .ZN(u5_mult_82_CARRYB_9__38_) );
  XNOR2_X2 u5_mult_82_U8039 ( .A(u5_mult_82_CARRYB_2__41_), .B(
        u5_mult_82_ab_3__41_), .ZN(u5_mult_82_n3282) );
  XNOR2_X2 u5_mult_82_U8038 ( .A(u5_mult_82_n3282), .B(u5_mult_82_SUMB_2__42_), 
        .ZN(u5_mult_82_SUMB_3__41_) );
  NAND2_X2 u5_mult_82_U8037 ( .A1(u5_mult_82_ab_6__48_), .A2(
        u5_mult_82_SUMB_5__49_), .ZN(u5_mult_82_n6349) );
  NAND2_X2 u5_mult_82_U8036 ( .A1(u5_mult_82_CARRYB_32__11_), .A2(
        u5_mult_82_SUMB_32__12_), .ZN(u5_mult_82_n5228) );
  NAND2_X2 u5_mult_82_U8035 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n1755), 
        .ZN(u5_mult_82_n5821) );
  NAND2_X2 u5_mult_82_U8034 ( .A1(u5_mult_82_ab_11__43_), .A2(
        u5_mult_82_SUMB_10__44_), .ZN(u5_mult_82_n5395) );
  INV_X2 u5_mult_82_U8033 ( .A(u5_mult_82_n5638), .ZN(u5_mult_82_n3562) );
  NAND2_X2 u5_mult_82_U8032 ( .A1(u5_mult_82_ab_37__15_), .A2(
        u5_mult_82_SUMB_36__16_), .ZN(u5_mult_82_n6177) );
  NAND3_X4 u5_mult_82_U8031 ( .A1(u5_mult_82_n6176), .A2(u5_mult_82_n6177), 
        .A3(u5_mult_82_n6178), .ZN(u5_mult_82_CARRYB_37__15_) );
  XNOR2_X2 u5_mult_82_U8030 ( .A(u5_mult_82_SUMB_5__47_), .B(u5_mult_82_n3279), 
        .ZN(u5_mult_82_SUMB_6__46_) );
  INV_X8 u5_mult_82_U8029 ( .A(u6_N52), .ZN(u5_mult_82_n6979) );
  XNOR2_X2 u5_mult_82_U8028 ( .A(u5_mult_82_SUMB_7__46_), .B(
        u5_mult_82_ab_8__45_), .ZN(u5_mult_82_n3278) );
  NAND2_X2 u5_mult_82_U8027 ( .A1(u5_mult_82_ab_13__38_), .A2(
        u5_mult_82_SUMB_12__39_), .ZN(u5_mult_82_n6160) );
  NAND3_X4 u5_mult_82_U8026 ( .A1(u5_mult_82_n5215), .A2(u5_mult_82_n5216), 
        .A3(u5_mult_82_n5217), .ZN(u5_mult_82_CARRYB_18__27_) );
  XNOR2_X2 u5_mult_82_U8025 ( .A(u5_mult_82_ab_8__36_), .B(
        u5_mult_82_CARRYB_7__36_), .ZN(u5_mult_82_n3277) );
  XNOR2_X2 u5_mult_82_U8024 ( .A(u5_mult_82_CARRYB_50__24_), .B(
        u5_mult_82_n3276), .ZN(u5_mult_82_n4463) );
  NAND2_X2 u5_mult_82_U8023 ( .A1(u5_mult_82_ab_33__11_), .A2(
        u5_mult_82_SUMB_32__12_), .ZN(u5_mult_82_n5227) );
  XNOR2_X2 u5_mult_82_U8022 ( .A(u5_mult_82_SUMB_7__49_), .B(u5_mult_82_n3275), 
        .ZN(u5_mult_82_SUMB_8__48_) );
  XNOR2_X2 u5_mult_82_U8021 ( .A(u5_mult_82_n3274), .B(
        u5_mult_82_CARRYB_49__25_), .ZN(u5_mult_82_n4462) );
  XNOR2_X1 u5_mult_82_U8020 ( .A(u5_mult_82_ab_16__25_), .B(
        u5_mult_82_CARRYB_15__25_), .ZN(u5_mult_82_n3273) );
  XNOR2_X2 u5_mult_82_U8019 ( .A(u5_mult_82_SUMB_9__47_), .B(u5_mult_82_n3507), 
        .ZN(u5_mult_82_SUMB_10__46_) );
  NAND3_X2 u5_mult_82_U8018 ( .A1(u5_mult_82_n3738), .A2(u5_mult_82_n3739), 
        .A3(u5_mult_82_n3740), .ZN(u5_mult_82_CARRYB_33__8_) );
  NOR2_X1 u5_mult_82_U8017 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_net65441), .ZN(u5_mult_82_ab_38__38_) );
  NOR2_X1 u5_mult_82_U8016 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6720), 
        .ZN(u5_mult_82_ab_37__38_) );
  NOR2_X1 u5_mult_82_U8015 ( .A1(u5_mult_82_n6849), .A2(u5_mult_82_net65279), 
        .ZN(u5_mult_82_ab_47__31_) );
  NAND3_X2 u5_mult_82_U8014 ( .A1(u5_mult_82_n3270), .A2(u5_mult_82_n3271), 
        .A3(u5_mult_82_n3272), .ZN(u5_mult_82_CARRYB_38__38_) );
  NAND2_X1 u5_mult_82_U8013 ( .A1(u5_mult_82_ab_38__38_), .A2(
        u5_mult_82_CARRYB_37__38_), .ZN(u5_mult_82_n3272) );
  NAND2_X2 u5_mult_82_U8012 ( .A1(u5_mult_82_ab_38__38_), .A2(
        u5_mult_82_SUMB_37__39_), .ZN(u5_mult_82_n3271) );
  NAND2_X1 u5_mult_82_U8011 ( .A1(u5_mult_82_CARRYB_37__38_), .A2(
        u5_mult_82_SUMB_37__39_), .ZN(u5_mult_82_n3270) );
  XOR2_X2 u5_mult_82_U8010 ( .A(u5_mult_82_SUMB_37__39_), .B(u5_mult_82_n3269), 
        .Z(u5_mult_82_SUMB_38__38_) );
  XOR2_X2 u5_mult_82_U8009 ( .A(u5_mult_82_CARRYB_37__38_), .B(
        u5_mult_82_ab_38__38_), .Z(u5_mult_82_n3269) );
  NAND3_X2 u5_mult_82_U8008 ( .A1(u5_mult_82_n3266), .A2(u5_mult_82_n3267), 
        .A3(u5_mult_82_n3268), .ZN(u5_mult_82_CARRYB_37__38_) );
  NAND2_X1 u5_mult_82_U8007 ( .A1(u5_mult_82_ab_37__38_), .A2(
        u5_mult_82_SUMB_36__39_), .ZN(u5_mult_82_n3268) );
  NAND2_X2 u5_mult_82_U8006 ( .A1(u5_mult_82_ab_37__38_), .A2(
        u5_mult_82_CARRYB_36__38_), .ZN(u5_mult_82_n3267) );
  NAND2_X1 u5_mult_82_U8005 ( .A1(u5_mult_82_SUMB_36__39_), .A2(
        u5_mult_82_CARRYB_36__38_), .ZN(u5_mult_82_n3266) );
  NAND3_X2 u5_mult_82_U8004 ( .A1(u5_mult_82_n3263), .A2(u5_mult_82_n3264), 
        .A3(u5_mult_82_n3265), .ZN(u5_mult_82_CARRYB_49__29_) );
  NAND2_X1 u5_mult_82_U8003 ( .A1(u5_mult_82_CARRYB_48__29_), .A2(
        u5_mult_82_SUMB_48__30_), .ZN(u5_mult_82_n3265) );
  NAND2_X1 u5_mult_82_U8002 ( .A1(u5_mult_82_ab_49__29_), .A2(
        u5_mult_82_SUMB_48__30_), .ZN(u5_mult_82_n3264) );
  NAND2_X1 u5_mult_82_U8001 ( .A1(u5_mult_82_ab_49__29_), .A2(
        u5_mult_82_CARRYB_48__29_), .ZN(u5_mult_82_n3263) );
  NAND2_X2 u5_mult_82_U8000 ( .A1(u5_mult_82_n1602), .A2(
        u5_mult_82_SUMB_47__31_), .ZN(u5_mult_82_n3262) );
  NAND2_X2 u5_mult_82_U7999 ( .A1(u5_mult_82_ab_48__30_), .A2(
        u5_mult_82_SUMB_47__31_), .ZN(u5_mult_82_n3261) );
  NAND2_X2 u5_mult_82_U7998 ( .A1(u5_mult_82_n1602), .A2(u5_mult_82_ab_48__30_), .ZN(u5_mult_82_n3260) );
  XOR2_X2 u5_mult_82_U7997 ( .A(u5_mult_82_n3259), .B(u5_mult_82_SUMB_47__31_), 
        .Z(u5_mult_82_SUMB_48__30_) );
  NAND3_X2 u5_mult_82_U7996 ( .A1(u5_mult_82_n3256), .A2(u5_mult_82_n3257), 
        .A3(u5_mult_82_n3258), .ZN(u5_mult_82_CARRYB_47__31_) );
  NAND2_X2 u5_mult_82_U7995 ( .A1(u5_mult_82_ab_47__31_), .A2(
        u5_mult_82_CARRYB_46__31_), .ZN(u5_mult_82_n3258) );
  NAND2_X2 u5_mult_82_U7994 ( .A1(u5_mult_82_ab_47__31_), .A2(
        u5_mult_82_SUMB_46__32_), .ZN(u5_mult_82_n3257) );
  NAND2_X2 u5_mult_82_U7993 ( .A1(u5_mult_82_CARRYB_46__31_), .A2(
        u5_mult_82_SUMB_46__32_), .ZN(u5_mult_82_n3256) );
  XNOR2_X2 u5_mult_82_U7992 ( .A(u5_mult_82_ab_32__24_), .B(
        u5_mult_82_CARRYB_31__24_), .ZN(u5_mult_82_n3255) );
  XOR2_X2 u5_mult_82_U7991 ( .A(u5_mult_82_n5607), .B(u5_mult_82_SUMB_19__25_), 
        .Z(u5_mult_82_SUMB_20__24_) );
  XNOR2_X2 u5_mult_82_U7990 ( .A(u5_mult_82_ab_46__5_), .B(
        u5_mult_82_CARRYB_45__5_), .ZN(u5_mult_82_n3254) );
  XNOR2_X2 u5_mult_82_U7989 ( .A(u5_mult_82_n3254), .B(u5_mult_82_SUMB_45__6_), 
        .ZN(u5_mult_82_SUMB_46__5_) );
  NAND2_X2 u5_mult_82_U7988 ( .A1(u5_mult_82_ab_33__11_), .A2(
        u5_mult_82_CARRYB_32__11_), .ZN(u5_mult_82_n5226) );
  NAND2_X2 u5_mult_82_U7987 ( .A1(u5_mult_82_ab_34__10_), .A2(
        u5_mult_82_SUMB_33__11_), .ZN(u5_mult_82_n4071) );
  XNOR2_X2 u5_mult_82_U7986 ( .A(u5_mult_82_CARRYB_16__25_), .B(
        u5_mult_82_ab_17__25_), .ZN(u5_mult_82_n3253) );
  XNOR2_X2 u5_mult_82_U7985 ( .A(u5_mult_82_n3253), .B(u5_mult_82_SUMB_16__26_), .ZN(u5_mult_82_SUMB_17__25_) );
  XNOR2_X2 u5_mult_82_U7984 ( .A(u5_mult_82_CARRYB_10__37_), .B(
        u5_mult_82_ab_11__37_), .ZN(u5_mult_82_n3252) );
  XNOR2_X2 u5_mult_82_U7983 ( .A(u5_mult_82_SUMB_10__38_), .B(u5_mult_82_n3252), .ZN(u5_mult_82_SUMB_11__37_) );
  XNOR2_X2 u5_mult_82_U7982 ( .A(u5_mult_82_ab_24__9_), .B(
        u5_mult_82_CARRYB_23__9_), .ZN(u5_mult_82_n3251) );
  XNOR2_X2 u5_mult_82_U7981 ( .A(u5_mult_82_CARRYB_9__42_), .B(
        u5_mult_82_ab_10__42_), .ZN(u5_mult_82_n3250) );
  XNOR2_X2 u5_mult_82_U7980 ( .A(u5_mult_82_SUMB_9__43_), .B(u5_mult_82_n3250), 
        .ZN(u5_mult_82_SUMB_10__42_) );
  NAND2_X2 u5_mult_82_U7979 ( .A1(u5_mult_82_ab_51__3_), .A2(
        u5_mult_82_CARRYB_50__3_), .ZN(u5_mult_82_n5241) );
  NOR2_X1 u5_mult_82_U7978 ( .A1(u5_mult_82_n6952), .A2(u5_mult_82_net65229), 
        .ZN(u5_mult_82_ab_50__3_) );
  NAND2_X1 u5_mult_82_U7977 ( .A1(u5_mult_82_ab_50__3_), .A2(
        u5_mult_82_CARRYB_49__3_), .ZN(u5_mult_82_n3249) );
  NAND2_X2 u5_mult_82_U7976 ( .A1(u5_mult_82_ab_50__3_), .A2(
        u5_mult_82_SUMB_49__4_), .ZN(u5_mult_82_n3248) );
  NAND2_X1 u5_mult_82_U7975 ( .A1(u5_mult_82_CARRYB_49__3_), .A2(
        u5_mult_82_SUMB_49__4_), .ZN(u5_mult_82_n3247) );
  NAND2_X1 u5_mult_82_U7974 ( .A1(u5_mult_82_ab_19__22_), .A2(
        u5_mult_82_SUMB_18__23_), .ZN(u5_mult_82_n3245) );
  NAND2_X1 u5_mult_82_U7973 ( .A1(u5_mult_82_ab_19__22_), .A2(
        u5_mult_82_CARRYB_18__22_), .ZN(u5_mult_82_n3244) );
  NAND3_X4 u5_mult_82_U7972 ( .A1(u5_mult_82_n3241), .A2(u5_mult_82_n3242), 
        .A3(u5_mult_82_n3243), .ZN(u5_mult_82_CARRYB_18__23_) );
  NAND2_X2 u5_mult_82_U7971 ( .A1(u5_mult_82_ab_18__23_), .A2(
        u5_mult_82_SUMB_17__24_), .ZN(u5_mult_82_n3243) );
  NAND2_X2 u5_mult_82_U7970 ( .A1(u5_mult_82_CARRYB_17__23_), .A2(
        u5_mult_82_SUMB_17__24_), .ZN(u5_mult_82_n3242) );
  NAND2_X1 u5_mult_82_U7969 ( .A1(u5_mult_82_CARRYB_17__23_), .A2(
        u5_mult_82_ab_18__23_), .ZN(u5_mult_82_n3241) );
  XOR2_X2 u5_mult_82_U7968 ( .A(u5_mult_82_n3240), .B(u5_mult_82_SUMB_17__24_), 
        .Z(u5_mult_82_SUMB_18__23_) );
  XOR2_X2 u5_mult_82_U7967 ( .A(u5_mult_82_CARRYB_17__23_), .B(
        u5_mult_82_ab_18__23_), .Z(u5_mult_82_n3240) );
  NAND3_X4 u5_mult_82_U7966 ( .A1(u5_mult_82_n4540), .A2(u5_mult_82_n4541), 
        .A3(u5_mult_82_n4542), .ZN(u5_mult_82_CARRYB_31__28_) );
  XNOR2_X2 u5_mult_82_U7965 ( .A(u5_mult_82_ab_19__43_), .B(
        u5_mult_82_CARRYB_18__43_), .ZN(u5_mult_82_n3239) );
  XNOR2_X2 u5_mult_82_U7964 ( .A(u5_mult_82_n1559), .B(u5_mult_82_n3239), .ZN(
        u5_mult_82_SUMB_19__43_) );
  XNOR2_X2 u5_mult_82_U7963 ( .A(u5_mult_82_n3238), .B(u5_mult_82_n104), .ZN(
        u5_mult_82_n3816) );
  NAND2_X1 u5_mult_82_U7962 ( .A1(u5_mult_82_CARRYB_44__17_), .A2(
        u5_mult_82_SUMB_44__18_), .ZN(u5_mult_82_n4013) );
  NOR2_X1 u5_mult_82_U7961 ( .A1(u5_mult_82_n6912), .A2(u5_mult_82_n6735), 
        .ZN(u5_mult_82_ab_44__19_) );
  NAND3_X2 u5_mult_82_U7960 ( .A1(u5_mult_82_n3235), .A2(u5_mult_82_n3236), 
        .A3(u5_mult_82_n3237), .ZN(u5_mult_82_CARRYB_44__19_) );
  NAND2_X1 u5_mult_82_U7959 ( .A1(u5_mult_82_ab_44__19_), .A2(
        u5_mult_82_CARRYB_43__19_), .ZN(u5_mult_82_n3237) );
  NAND2_X2 u5_mult_82_U7958 ( .A1(u5_mult_82_ab_44__19_), .A2(
        u5_mult_82_SUMB_43__20_), .ZN(u5_mult_82_n3236) );
  INV_X4 u5_mult_82_U7957 ( .A(u5_mult_82_n3510), .ZN(u5_mult_82_n3231) );
  NAND2_X4 u5_mult_82_U7956 ( .A1(u5_mult_82_n3233), .A2(u5_mult_82_n3234), 
        .ZN(u5_mult_82_SUMB_18__36_) );
  NAND2_X2 u5_mult_82_U7955 ( .A1(u5_mult_82_n3231), .A2(u5_mult_82_n3232), 
        .ZN(u5_mult_82_n3234) );
  NAND3_X2 u5_mult_82_U7954 ( .A1(u5_mult_82_n3228), .A2(u5_mult_82_n3229), 
        .A3(u5_mult_82_n3230), .ZN(u5_mult_82_CARRYB_29__29_) );
  NAND2_X1 u5_mult_82_U7953 ( .A1(u5_mult_82_SUMB_28__30_), .A2(
        u5_mult_82_CARRYB_28__29_), .ZN(u5_mult_82_n3230) );
  NAND2_X1 u5_mult_82_U7952 ( .A1(u5_mult_82_ab_29__29_), .A2(
        u5_mult_82_SUMB_28__30_), .ZN(u5_mult_82_n3229) );
  NAND2_X1 u5_mult_82_U7951 ( .A1(u5_mult_82_ab_29__29_), .A2(
        u5_mult_82_CARRYB_28__29_), .ZN(u5_mult_82_n3228) );
  NAND3_X2 u5_mult_82_U7950 ( .A1(u5_mult_82_n3225), .A2(u5_mult_82_n3226), 
        .A3(u5_mult_82_n3227), .ZN(u5_mult_82_CARRYB_28__30_) );
  NAND2_X1 u5_mult_82_U7949 ( .A1(u5_mult_82_ab_28__30_), .A2(
        u5_mult_82_CARRYB_27__30_), .ZN(u5_mult_82_n3225) );
  XOR2_X2 u5_mult_82_U7948 ( .A(u5_mult_82_n3224), .B(u5_mult_82_SUMB_28__30_), 
        .Z(u5_mult_82_SUMB_29__29_) );
  XOR2_X2 u5_mult_82_U7947 ( .A(u5_mult_82_ab_29__29_), .B(
        u5_mult_82_CARRYB_28__29_), .Z(u5_mult_82_n3224) );
  XOR2_X2 u5_mult_82_U7946 ( .A(u5_mult_82_n3223), .B(u5_mult_82_n1851), .Z(
        u5_mult_82_SUMB_28__30_) );
  NAND3_X2 u5_mult_82_U7945 ( .A1(u5_mult_82_n3220), .A2(u5_mult_82_n3221), 
        .A3(u5_mult_82_n3222), .ZN(u5_mult_82_CARRYB_49__16_) );
  NAND2_X1 u5_mult_82_U7944 ( .A1(u5_mult_82_ab_49__16_), .A2(
        u5_mult_82_SUMB_48__17_), .ZN(u5_mult_82_n3222) );
  NAND2_X1 u5_mult_82_U7943 ( .A1(u5_mult_82_CARRYB_48__16_), .A2(
        u5_mult_82_SUMB_48__17_), .ZN(u5_mult_82_n3221) );
  NAND2_X1 u5_mult_82_U7942 ( .A1(u5_mult_82_CARRYB_48__16_), .A2(
        u5_mult_82_ab_49__16_), .ZN(u5_mult_82_n3220) );
  NAND2_X2 u5_mult_82_U7941 ( .A1(u5_mult_82_CARRYB_47__17_), .A2(
        u5_mult_82_SUMB_47__18_), .ZN(u5_mult_82_n3219) );
  NAND2_X2 u5_mult_82_U7940 ( .A1(u5_mult_82_ab_48__17_), .A2(
        u5_mult_82_SUMB_47__18_), .ZN(u5_mult_82_n3218) );
  NAND2_X1 u5_mult_82_U7939 ( .A1(u5_mult_82_ab_48__17_), .A2(
        u5_mult_82_CARRYB_47__17_), .ZN(u5_mult_82_n3217) );
  XOR2_X2 u5_mult_82_U7938 ( .A(u5_mult_82_n3216), .B(u5_mult_82_SUMB_48__17_), 
        .Z(u5_mult_82_SUMB_49__16_) );
  XOR2_X2 u5_mult_82_U7937 ( .A(u5_mult_82_CARRYB_48__16_), .B(
        u5_mult_82_ab_49__16_), .Z(u5_mult_82_n3216) );
  NAND2_X2 u5_mult_82_U7936 ( .A1(u5_mult_82_ab_31__10_), .A2(
        u5_mult_82_CARRYB_30__10_), .ZN(u5_mult_82_n5309) );
  NAND3_X4 u5_mult_82_U7935 ( .A1(u5_mult_82_n3735), .A2(u5_mult_82_n3736), 
        .A3(u5_mult_82_n3737), .ZN(u5_mult_82_CARRYB_29__10_) );
  NOR2_X2 u5_mult_82_U7934 ( .A1(u5_mult_82_net64451), .A2(u5_mult_82_n6680), 
        .ZN(u5_mult_82_ab_30__10_) );
  NOR2_X1 u5_mult_82_U7933 ( .A1(u5_mult_82_n6905), .A2(u5_mult_82_n6602), 
        .ZN(u5_mult_82_ab_17__20_) );
  NAND2_X2 u5_mult_82_U7932 ( .A1(u5_mult_82_ab_26__13_), .A2(
        u5_mult_82_CARRYB_25__13_), .ZN(u5_mult_82_n4833) );
  NAND2_X2 u5_mult_82_U7931 ( .A1(u5_mult_82_CARRYB_25__13_), .A2(
        u5_mult_82_SUMB_25__14_), .ZN(u5_mult_82_n4835) );
  NOR2_X2 u5_mult_82_U7930 ( .A1(u5_mult_82_net64507), .A2(u5_mult_82_net65679), .ZN(u5_mult_82_ab_25__13_) );
  NAND2_X2 u5_mult_82_U7929 ( .A1(u5_mult_82_ab_47__2_), .A2(
        u5_mult_82_CARRYB_46__2_), .ZN(u5_mult_82_n4515) );
  NAND2_X4 u5_mult_82_U7928 ( .A1(u5_mult_82_n3563), .A2(u5_mult_82_n3564), 
        .ZN(u5_mult_82_SUMB_45__3_) );
  NOR2_X2 u5_mult_82_U7927 ( .A1(u5_mult_82_n6960), .A2(u5_mult_82_n6743), 
        .ZN(u5_mult_82_ab_46__2_) );
  NOR2_X2 u5_mult_82_U7926 ( .A1(u5_mult_82_net64361), .A2(u5_mult_82_n6729), 
        .ZN(u5_mult_82_ab_39__5_) );
  NOR2_X1 u5_mult_82_U7925 ( .A1(u5_mult_82_net64379), .A2(u5_mult_82_n6722), 
        .ZN(u5_mult_82_ab_37__6_) );
  NAND2_X1 u5_mult_82_U7924 ( .A1(u5_mult_82_ab_30__10_), .A2(
        u5_mult_82_CARRYB_29__10_), .ZN(u5_mult_82_n3215) );
  NAND2_X2 u5_mult_82_U7923 ( .A1(u5_mult_82_CARRYB_29__10_), .A2(
        u5_mult_82_SUMB_29__11_), .ZN(u5_mult_82_n3213) );
  XOR2_X2 u5_mult_82_U7922 ( .A(u5_mult_82_SUMB_29__11_), .B(u5_mult_82_n3212), 
        .Z(u5_mult_82_SUMB_30__10_) );
  NAND3_X4 u5_mult_82_U7921 ( .A1(u5_mult_82_n3209), .A2(u5_mult_82_n3210), 
        .A3(u5_mult_82_n3211), .ZN(u5_mult_82_CARRYB_17__20_) );
  NAND2_X1 u5_mult_82_U7920 ( .A1(u5_mult_82_ab_17__20_), .A2(
        u5_mult_82_CARRYB_16__20_), .ZN(u5_mult_82_n3211) );
  NAND2_X2 u5_mult_82_U7919 ( .A1(u5_mult_82_ab_17__20_), .A2(u5_mult_82_n1642), .ZN(u5_mult_82_n3210) );
  NAND3_X4 u5_mult_82_U7918 ( .A1(u5_mult_82_n3206), .A2(u5_mult_82_n3207), 
        .A3(u5_mult_82_n3208), .ZN(u5_mult_82_CARRYB_25__13_) );
  NAND2_X1 u5_mult_82_U7917 ( .A1(u5_mult_82_ab_25__13_), .A2(
        u5_mult_82_CARRYB_24__13_), .ZN(u5_mult_82_n3208) );
  NAND2_X2 u5_mult_82_U7916 ( .A1(u5_mult_82_ab_25__13_), .A2(u5_mult_82_n1797), .ZN(u5_mult_82_n3207) );
  NAND2_X2 u5_mult_82_U7915 ( .A1(u5_mult_82_CARRYB_24__13_), .A2(
        u5_mult_82_n1797), .ZN(u5_mult_82_n3206) );
  XOR2_X2 u5_mult_82_U7914 ( .A(u5_mult_82_n1797), .B(u5_mult_82_n3205), .Z(
        u5_mult_82_SUMB_25__13_) );
  XOR2_X2 u5_mult_82_U7913 ( .A(u5_mult_82_CARRYB_24__13_), .B(
        u5_mult_82_ab_25__13_), .Z(u5_mult_82_n3205) );
  NAND3_X4 u5_mult_82_U7912 ( .A1(u5_mult_82_n3202), .A2(u5_mult_82_n3203), 
        .A3(u5_mult_82_n3204), .ZN(u5_mult_82_CARRYB_46__2_) );
  NAND2_X2 u5_mult_82_U7911 ( .A1(u5_mult_82_ab_46__2_), .A2(
        u5_mult_82_CARRYB_45__2_), .ZN(u5_mult_82_n3204) );
  NAND2_X4 u5_mult_82_U7910 ( .A1(u5_mult_82_ab_46__2_), .A2(
        u5_mult_82_SUMB_45__3_), .ZN(u5_mult_82_n3203) );
  NAND2_X2 u5_mult_82_U7909 ( .A1(u5_mult_82_CARRYB_45__2_), .A2(
        u5_mult_82_SUMB_45__3_), .ZN(u5_mult_82_n3202) );
  NAND2_X1 u5_mult_82_U7908 ( .A1(u5_mult_82_ab_39__5_), .A2(
        u5_mult_82_CARRYB_38__5_), .ZN(u5_mult_82_n3201) );
  NAND2_X2 u5_mult_82_U7907 ( .A1(u5_mult_82_SUMB_38__6_), .A2(
        u5_mult_82_ab_39__5_), .ZN(u5_mult_82_n3200) );
  NAND2_X2 u5_mult_82_U7906 ( .A1(u5_mult_82_CARRYB_38__5_), .A2(
        u5_mult_82_SUMB_38__6_), .ZN(u5_mult_82_n3199) );
  NAND3_X2 u5_mult_82_U7905 ( .A1(u5_mult_82_n3196), .A2(u5_mult_82_n3197), 
        .A3(u5_mult_82_n3198), .ZN(u5_mult_82_CARRYB_37__6_) );
  NAND2_X2 u5_mult_82_U7904 ( .A1(u5_mult_82_ab_37__6_), .A2(
        u5_mult_82_CARRYB_36__6_), .ZN(u5_mult_82_n3197) );
  NAND2_X1 u5_mult_82_U7903 ( .A1(u5_mult_82_SUMB_36__7_), .A2(
        u5_mult_82_CARRYB_36__6_), .ZN(u5_mult_82_n3196) );
  XNOR2_X2 u5_mult_82_U7902 ( .A(u5_mult_82_ab_12__29_), .B(
        u5_mult_82_CARRYB_11__29_), .ZN(u5_mult_82_n3195) );
  XNOR2_X2 u5_mult_82_U7901 ( .A(u5_mult_82_n3195), .B(u5_mult_82_SUMB_11__30_), .ZN(u5_mult_82_SUMB_12__29_) );
  XNOR2_X2 u5_mult_82_U7900 ( .A(u5_mult_82_CARRYB_8__46_), .B(
        u5_mult_82_ab_9__46_), .ZN(u5_mult_82_n3194) );
  XNOR2_X2 u5_mult_82_U7899 ( .A(u5_mult_82_n3194), .B(u5_mult_82_n1681), .ZN(
        u5_mult_82_SUMB_9__46_) );
  NAND2_X2 u5_mult_82_U7898 ( .A1(u5_mult_82_CARRYB_49__0_), .A2(
        u5_mult_82_SUMB_49__1_), .ZN(u5_mult_82_n3424) );
  XNOR2_X2 u5_mult_82_U7897 ( .A(u5_mult_82_n3193), .B(
        u5_mult_82_CARRYB_45__3_), .ZN(u5_mult_82_n4510) );
  NAND2_X1 u5_mult_82_U7896 ( .A1(u5_mult_82_ab_34__15_), .A2(
        u5_mult_82_CARRYB_33__15_), .ZN(u5_mult_82_n6037) );
  NAND2_X2 u5_mult_82_U7895 ( .A1(u5_mult_82_ab_25__20_), .A2(
        u5_mult_82_SUMB_24__21_), .ZN(u5_mult_82_n5694) );
  NAND2_X2 u5_mult_82_U7894 ( .A1(u5_mult_82_CARRYB_24__20_), .A2(
        u5_mult_82_SUMB_24__21_), .ZN(u5_mult_82_n5695) );
  NOR2_X1 u5_mult_82_U7893 ( .A1(u5_mult_82_net64489), .A2(u5_mult_82_n6610), 
        .ZN(u5_mult_82_ab_18__12_) );
  NAND3_X2 u5_mult_82_U7892 ( .A1(u5_mult_82_n3190), .A2(u5_mult_82_n3191), 
        .A3(u5_mult_82_n3192), .ZN(u5_mult_82_CARRYB_18__12_) );
  NAND2_X1 u5_mult_82_U7891 ( .A1(u5_mult_82_ab_18__12_), .A2(
        u5_mult_82_CARRYB_17__12_), .ZN(u5_mult_82_n3192) );
  NAND2_X2 u5_mult_82_U7890 ( .A1(u5_mult_82_ab_18__12_), .A2(
        u5_mult_82_SUMB_17__13_), .ZN(u5_mult_82_n3191) );
  NAND2_X1 u5_mult_82_U7889 ( .A1(u5_mult_82_CARRYB_17__12_), .A2(
        u5_mult_82_SUMB_17__13_), .ZN(u5_mult_82_n3190) );
  XOR2_X2 u5_mult_82_U7888 ( .A(u5_mult_82_SUMB_17__13_), .B(u5_mult_82_n3189), 
        .Z(u5_mult_82_SUMB_18__12_) );
  XOR2_X2 u5_mult_82_U7887 ( .A(u5_mult_82_CARRYB_17__12_), .B(
        u5_mult_82_ab_18__12_), .Z(u5_mult_82_n3189) );
  NAND3_X2 u5_mult_82_U7886 ( .A1(u5_mult_82_n3186), .A2(u5_mult_82_n3187), 
        .A3(u5_mult_82_n3188), .ZN(u5_mult_82_CARRYB_3__25_) );
  NAND2_X1 u5_mult_82_U7885 ( .A1(u5_mult_82_CARRYB_2__25_), .A2(
        u5_mult_82_SUMB_2__26_), .ZN(u5_mult_82_n3188) );
  NAND2_X1 u5_mult_82_U7884 ( .A1(u5_mult_82_ab_3__25_), .A2(
        u5_mult_82_SUMB_2__26_), .ZN(u5_mult_82_n3187) );
  NAND2_X1 u5_mult_82_U7883 ( .A1(u5_mult_82_CARRYB_2__25_), .A2(
        u5_mult_82_ab_3__25_), .ZN(u5_mult_82_n3186) );
  NAND3_X4 u5_mult_82_U7882 ( .A1(u5_mult_82_n3183), .A2(u5_mult_82_n3184), 
        .A3(u5_mult_82_n3185), .ZN(u5_mult_82_CARRYB_2__26_) );
  NAND2_X2 u5_mult_82_U7881 ( .A1(u5_mult_82_CARRYB_1__26_), .A2(
        u5_mult_82_SUMB_1__27_), .ZN(u5_mult_82_n3185) );
  NAND2_X2 u5_mult_82_U7880 ( .A1(u5_mult_82_ab_2__26_), .A2(
        u5_mult_82_SUMB_1__27_), .ZN(u5_mult_82_n3184) );
  NAND2_X1 u5_mult_82_U7879 ( .A1(u5_mult_82_ab_2__26_), .A2(
        u5_mult_82_CARRYB_1__26_), .ZN(u5_mult_82_n3183) );
  XOR2_X2 u5_mult_82_U7878 ( .A(u5_mult_82_n3182), .B(u5_mult_82_SUMB_1__27_), 
        .Z(u5_mult_82_SUMB_2__26_) );
  NAND3_X2 u5_mult_82_U7877 ( .A1(u5_mult_82_n3179), .A2(u5_mult_82_n3180), 
        .A3(u5_mult_82_n3181), .ZN(u5_mult_82_CARRYB_35__4_) );
  NAND2_X1 u5_mult_82_U7876 ( .A1(u5_mult_82_CARRYB_34__4_), .A2(
        u5_mult_82_SUMB_34__5_), .ZN(u5_mult_82_n3181) );
  NAND2_X1 u5_mult_82_U7875 ( .A1(u5_mult_82_ab_35__4_), .A2(
        u5_mult_82_CARRYB_34__4_), .ZN(u5_mult_82_n3179) );
  NAND3_X2 u5_mult_82_U7874 ( .A1(u5_mult_82_n3176), .A2(u5_mult_82_n3177), 
        .A3(u5_mult_82_n3178), .ZN(u5_mult_82_CARRYB_34__5_) );
  NAND2_X2 u5_mult_82_U7873 ( .A1(u5_mult_82_CARRYB_33__5_), .A2(
        u5_mult_82_SUMB_33__6_), .ZN(u5_mult_82_n3178) );
  NAND2_X2 u5_mult_82_U7872 ( .A1(u5_mult_82_ab_34__5_), .A2(
        u5_mult_82_SUMB_33__6_), .ZN(u5_mult_82_n3177) );
  XOR2_X1 u5_mult_82_U7871 ( .A(u5_mult_82_ab_35__4_), .B(
        u5_mult_82_CARRYB_34__4_), .Z(u5_mult_82_n3175) );
  XNOR2_X2 u5_mult_82_U7870 ( .A(u5_mult_82_n3174), .B(u5_mult_82_SUMB_42__10_), .ZN(u5_mult_82_SUMB_43__9_) );
  INV_X2 u5_mult_82_U7869 ( .A(u5_mult_82_SUMB_50__26_), .ZN(u5_mult_82_n3607)
         );
  XNOR2_X2 u5_mult_82_U7868 ( .A(u5_mult_82_ab_36__35_), .B(
        u5_mult_82_CARRYB_35__35_), .ZN(u5_mult_82_n3173) );
  XNOR2_X2 u5_mult_82_U7867 ( .A(u5_mult_82_n3173), .B(u5_mult_82_SUMB_35__36_), .ZN(u5_mult_82_SUMB_36__35_) );
  XNOR2_X2 u5_mult_82_U7866 ( .A(u5_mult_82_ab_19__27_), .B(
        u5_mult_82_CARRYB_18__27_), .ZN(u5_mult_82_n3172) );
  XNOR2_X2 u5_mult_82_U7865 ( .A(u5_mult_82_n3172), .B(u5_mult_82_SUMB_18__28_), .ZN(u5_mult_82_SUMB_19__27_) );
  NOR2_X1 u5_mult_82_U7864 ( .A1(u5_mult_82_n6882), .A2(u5_mult_82_n6579), 
        .ZN(u5_mult_82_ab_14__26_) );
  NAND3_X2 u5_mult_82_U7863 ( .A1(u5_mult_82_n3169), .A2(u5_mult_82_n3170), 
        .A3(u5_mult_82_n3171), .ZN(u5_mult_82_CARRYB_14__26_) );
  NAND2_X1 u5_mult_82_U7862 ( .A1(u5_mult_82_ab_14__26_), .A2(
        u5_mult_82_CARRYB_13__26_), .ZN(u5_mult_82_n3171) );
  NAND2_X2 u5_mult_82_U7861 ( .A1(u5_mult_82_ab_14__26_), .A2(
        u5_mult_82_SUMB_13__27_), .ZN(u5_mult_82_n3170) );
  NAND2_X1 u5_mult_82_U7860 ( .A1(u5_mult_82_CARRYB_13__26_), .A2(
        u5_mult_82_SUMB_13__27_), .ZN(u5_mult_82_n3169) );
  NAND3_X4 u5_mult_82_U7859 ( .A1(u5_mult_82_n3166), .A2(u5_mult_82_n3167), 
        .A3(u5_mult_82_n3168), .ZN(u5_mult_82_CARRYB_23__21_) );
  NAND2_X2 u5_mult_82_U7858 ( .A1(u5_mult_82_CARRYB_22__21_), .A2(
        u5_mult_82_SUMB_22__22_), .ZN(u5_mult_82_n3168) );
  NAND2_X2 u5_mult_82_U7857 ( .A1(u5_mult_82_ab_23__21_), .A2(
        u5_mult_82_SUMB_22__22_), .ZN(u5_mult_82_n3167) );
  NAND2_X1 u5_mult_82_U7856 ( .A1(u5_mult_82_ab_23__21_), .A2(
        u5_mult_82_CARRYB_22__21_), .ZN(u5_mult_82_n3166) );
  NAND3_X4 u5_mult_82_U7855 ( .A1(u5_mult_82_n3163), .A2(u5_mult_82_n3164), 
        .A3(u5_mult_82_n3165), .ZN(u5_mult_82_CARRYB_22__22_) );
  NAND2_X2 u5_mult_82_U7854 ( .A1(u5_mult_82_CARRYB_21__22_), .A2(
        u5_mult_82_SUMB_21__23_), .ZN(u5_mult_82_n3165) );
  NAND2_X2 u5_mult_82_U7853 ( .A1(u5_mult_82_ab_22__22_), .A2(
        u5_mult_82_SUMB_21__23_), .ZN(u5_mult_82_n3164) );
  NAND2_X1 u5_mult_82_U7852 ( .A1(u5_mult_82_ab_22__22_), .A2(
        u5_mult_82_CARRYB_21__22_), .ZN(u5_mult_82_n3163) );
  XOR2_X2 u5_mult_82_U7851 ( .A(u5_mult_82_n3162), .B(u5_mult_82_SUMB_22__22_), 
        .Z(u5_mult_82_SUMB_23__21_) );
  NAND2_X1 u5_mult_82_U7850 ( .A1(u5_mult_82_CARRYB_26__18_), .A2(
        u5_mult_82_SUMB_26__19_), .ZN(u5_mult_82_n3161) );
  NAND2_X1 u5_mult_82_U7849 ( .A1(u5_mult_82_ab_27__18_), .A2(
        u5_mult_82_SUMB_26__19_), .ZN(u5_mult_82_n3160) );
  NAND2_X1 u5_mult_82_U7848 ( .A1(u5_mult_82_ab_27__18_), .A2(
        u5_mult_82_CARRYB_26__18_), .ZN(u5_mult_82_n3159) );
  NAND3_X2 u5_mult_82_U7847 ( .A1(u5_mult_82_n3156), .A2(u5_mult_82_n3157), 
        .A3(u5_mult_82_n3158), .ZN(u5_mult_82_CARRYB_26__19_) );
  NAND2_X2 u5_mult_82_U7846 ( .A1(u5_mult_82_ab_26__19_), .A2(
        u5_mult_82_SUMB_25__20_), .ZN(u5_mult_82_n3157) );
  NAND2_X1 u5_mult_82_U7845 ( .A1(u5_mult_82_ab_26__19_), .A2(
        u5_mult_82_CARRYB_25__19_), .ZN(u5_mult_82_n3156) );
  XOR2_X2 u5_mult_82_U7844 ( .A(u5_mult_82_n3155), .B(u5_mult_82_SUMB_25__20_), 
        .Z(u5_mult_82_SUMB_26__19_) );
  XOR2_X2 u5_mult_82_U7843 ( .A(u5_mult_82_ab_26__19_), .B(
        u5_mult_82_CARRYB_25__19_), .Z(u5_mult_82_n3155) );
  INV_X4 u5_mult_82_U7842 ( .A(u5_mult_82_SUMB_12__37_), .ZN(u5_mult_82_n4868)
         );
  NAND3_X2 u5_mult_82_U7841 ( .A1(u5_mult_82_n5991), .A2(u5_mult_82_n5992), 
        .A3(u5_mult_82_n5993), .ZN(u5_mult_82_CARRYB_50__11_) );
  NAND2_X1 u5_mult_82_U7840 ( .A1(u5_mult_82_n3969), .A2(
        u5_mult_82_SUMB_14__49_), .ZN(u5_mult_82_n3364) );
  NAND2_X2 u5_mult_82_U7839 ( .A1(u5_mult_82_CARRYB_17__25_), .A2(
        u5_mult_82_SUMB_17__26_), .ZN(u5_mult_82_n4779) );
  XNOR2_X2 u5_mult_82_U7838 ( .A(u5_mult_82_n3154), .B(u5_mult_82_SUMB_27__24_), .ZN(u5_mult_82_SUMB_28__23_) );
  NAND2_X1 u5_mult_82_U7837 ( .A1(u5_mult_82_n633), .A2(u5_mult_82_SUMB_36__6_), .ZN(u5_mult_82_n4104) );
  XNOR2_X2 u5_mult_82_U7836 ( .A(u5_mult_82_n3152), .B(
        u5_mult_82_CARRYB_12__46_), .ZN(u5_mult_82_n4588) );
  NAND2_X2 u5_mult_82_U7835 ( .A1(u5_mult_82_CARRYB_44__1_), .A2(
        u5_mult_82_SUMB_44__2_), .ZN(u5_mult_82_n3438) );
  XNOR2_X2 u5_mult_82_U7834 ( .A(u5_mult_82_n3151), .B(u5_mult_82_SUMB_19__33_), .ZN(u5_mult_82_SUMB_20__32_) );
  INV_X2 u5_mult_82_U7833 ( .A(u5_mult_82_ab_16__34_), .ZN(u5_mult_82_n4865)
         );
  NAND3_X2 u5_mult_82_U7832 ( .A1(u5_mult_82_n3148), .A2(u5_mult_82_n3149), 
        .A3(u5_mult_82_n3150), .ZN(u5_mult_82_CARRYB_23__29_) );
  NAND2_X1 u5_mult_82_U7831 ( .A1(u5_mult_82_CARRYB_22__29_), .A2(
        u5_mult_82_SUMB_22__30_), .ZN(u5_mult_82_n3150) );
  NAND2_X1 u5_mult_82_U7830 ( .A1(u5_mult_82_ab_23__29_), .A2(
        u5_mult_82_SUMB_22__30_), .ZN(u5_mult_82_n3149) );
  NAND2_X1 u5_mult_82_U7829 ( .A1(u5_mult_82_ab_23__29_), .A2(
        u5_mult_82_CARRYB_22__29_), .ZN(u5_mult_82_n3148) );
  NAND2_X2 u5_mult_82_U7828 ( .A1(u5_mult_82_ab_22__30_), .A2(u5_mult_82_n1791), .ZN(u5_mult_82_n3146) );
  NAND2_X1 u5_mult_82_U7827 ( .A1(u5_mult_82_ab_22__30_), .A2(
        u5_mult_82_CARRYB_21__30_), .ZN(u5_mult_82_n3145) );
  XOR2_X2 u5_mult_82_U7826 ( .A(u5_mult_82_n3144), .B(u5_mult_82_SUMB_22__30_), 
        .Z(u5_mult_82_SUMB_23__29_) );
  XOR2_X2 u5_mult_82_U7825 ( .A(u5_mult_82_n3143), .B(u5_mult_82_n1791), .Z(
        u5_mult_82_SUMB_22__30_) );
  INV_X4 u5_mult_82_U7824 ( .A(u5_mult_82_CARRYB_15__34_), .ZN(
        u5_mult_82_n3140) );
  NAND2_X2 u5_mult_82_U7823 ( .A1(u5_mult_82_n4865), .A2(
        u5_mult_82_CARRYB_15__34_), .ZN(u5_mult_82_n3141) );
  INV_X2 u5_mult_82_U7822 ( .A(u5_mult_82_ab_43__18_), .ZN(u5_mult_82_n3137)
         );
  NAND2_X2 u5_mult_82_U7821 ( .A1(u5_mult_82_n3138), .A2(u5_mult_82_n3137), 
        .ZN(u5_mult_82_n3139) );
  NAND2_X2 u5_mult_82_U7820 ( .A1(u5_mult_82_CARRYB_8__45_), .A2(
        u5_mult_82_n1853), .ZN(u5_mult_82_n6354) );
  NAND2_X1 u5_mult_82_U7819 ( .A1(u5_mult_82_CARRYB_15__41_), .A2(
        u5_mult_82_SUMB_15__42_), .ZN(u5_mult_82_n3136) );
  NAND2_X1 u5_mult_82_U7818 ( .A1(u5_mult_82_ab_16__41_), .A2(
        u5_mult_82_SUMB_15__42_), .ZN(u5_mult_82_n3135) );
  NAND2_X1 u5_mult_82_U7817 ( .A1(u5_mult_82_ab_16__41_), .A2(
        u5_mult_82_CARRYB_15__41_), .ZN(u5_mult_82_n3134) );
  NAND3_X2 u5_mult_82_U7816 ( .A1(u5_mult_82_n3131), .A2(u5_mult_82_n3132), 
        .A3(u5_mult_82_n3133), .ZN(u5_mult_82_CARRYB_15__42_) );
  NAND2_X1 u5_mult_82_U7815 ( .A1(u5_mult_82_ab_15__42_), .A2(
        u5_mult_82_CARRYB_14__42_), .ZN(u5_mult_82_n3131) );
  NAND2_X1 u5_mult_82_U7814 ( .A1(u5_mult_82_CARRYB_7__47_), .A2(
        u5_mult_82_SUMB_7__48_), .ZN(u5_mult_82_n3130) );
  NAND2_X1 u5_mult_82_U7813 ( .A1(u5_mult_82_ab_8__47_), .A2(
        u5_mult_82_CARRYB_7__47_), .ZN(u5_mult_82_n3128) );
  NAND3_X2 u5_mult_82_U7812 ( .A1(u5_mult_82_n3125), .A2(u5_mult_82_n3126), 
        .A3(u5_mult_82_n3127), .ZN(u5_mult_82_CARRYB_7__48_) );
  NAND2_X2 u5_mult_82_U7811 ( .A1(u5_mult_82_CARRYB_6__48_), .A2(
        u5_mult_82_SUMB_6__49_), .ZN(u5_mult_82_n3127) );
  NAND2_X2 u5_mult_82_U7810 ( .A1(u5_mult_82_ab_7__48_), .A2(
        u5_mult_82_SUMB_6__49_), .ZN(u5_mult_82_n3126) );
  NAND2_X1 u5_mult_82_U7809 ( .A1(u5_mult_82_ab_7__48_), .A2(
        u5_mult_82_CARRYB_6__48_), .ZN(u5_mult_82_n3125) );
  XOR2_X2 u5_mult_82_U7808 ( .A(u5_mult_82_n3124), .B(u5_mult_82_SUMB_7__48_), 
        .Z(u5_mult_82_SUMB_8__47_) );
  XOR2_X2 u5_mult_82_U7807 ( .A(u5_mult_82_n3123), .B(u5_mult_82_SUMB_6__49_), 
        .Z(u5_mult_82_SUMB_7__48_) );
  XOR2_X2 u5_mult_82_U7806 ( .A(u5_mult_82_ab_7__48_), .B(
        u5_mult_82_CARRYB_6__48_), .Z(u5_mult_82_n3123) );
  NAND3_X2 u5_mult_82_U7805 ( .A1(u5_mult_82_n3120), .A2(u5_mult_82_n3121), 
        .A3(u5_mult_82_n3122), .ZN(u5_mult_82_CARRYB_29__34_) );
  NAND2_X1 u5_mult_82_U7804 ( .A1(u5_mult_82_n1665), .A2(
        u5_mult_82_SUMB_28__35_), .ZN(u5_mult_82_n3122) );
  NAND2_X1 u5_mult_82_U7803 ( .A1(u5_mult_82_ab_29__34_), .A2(
        u5_mult_82_SUMB_28__35_), .ZN(u5_mult_82_n3121) );
  NAND2_X1 u5_mult_82_U7802 ( .A1(u5_mult_82_ab_29__34_), .A2(u5_mult_82_n1665), .ZN(u5_mult_82_n3120) );
  NAND2_X2 u5_mult_82_U7801 ( .A1(u5_mult_82_ab_28__35_), .A2(u5_mult_82_n2320), .ZN(u5_mult_82_n3119) );
  NAND2_X1 u5_mult_82_U7800 ( .A1(u5_mult_82_CARRYB_27__35_), .A2(
        u5_mult_82_ab_28__35_), .ZN(u5_mult_82_n3117) );
  XOR2_X2 u5_mult_82_U7799 ( .A(u5_mult_82_n3116), .B(u5_mult_82_n2320), .Z(
        u5_mult_82_SUMB_28__35_) );
  XOR2_X2 u5_mult_82_U7798 ( .A(u5_mult_82_CARRYB_27__35_), .B(
        u5_mult_82_ab_28__35_), .Z(u5_mult_82_n3116) );
  XNOR2_X2 u5_mult_82_U7797 ( .A(u5_mult_82_CARRYB_46__16_), .B(
        u5_mult_82_n3115), .ZN(u5_mult_82_n5860) );
  NAND3_X2 u5_mult_82_U7796 ( .A1(u5_mult_82_n3114), .A2(u5_mult_82_n3113), 
        .A3(u5_mult_82_n3112), .ZN(u5_mult_82_CARRYB_20__34_) );
  NAND2_X1 u5_mult_82_U7795 ( .A1(u5_mult_82_CARRYB_19__34_), .A2(
        u5_mult_82_SUMB_19__35_), .ZN(u5_mult_82_n3114) );
  NAND3_X2 u5_mult_82_U7794 ( .A1(u5_mult_82_n3109), .A2(u5_mult_82_n3110), 
        .A3(u5_mult_82_n3111), .ZN(u5_mult_82_CARRYB_19__35_) );
  NAND2_X2 u5_mult_82_U7793 ( .A1(u5_mult_82_CARRYB_18__35_), .A2(
        u5_mult_82_SUMB_18__36_), .ZN(u5_mult_82_n3111) );
  NAND2_X2 u5_mult_82_U7792 ( .A1(u5_mult_82_ab_19__35_), .A2(
        u5_mult_82_SUMB_18__36_), .ZN(u5_mult_82_n3110) );
  XNOR2_X2 u5_mult_82_U7791 ( .A(u5_mult_82_CARRYB_33__6_), .B(
        u5_mult_82_ab_34__6_), .ZN(u5_mult_82_n3108) );
  NOR2_X1 u5_mult_82_U7790 ( .A1(u5_mult_82_n6785), .A2(u5_mult_82_n6615), 
        .ZN(u5_mult_82_ab_19__47_) );
  NOR2_X1 u5_mult_82_U7789 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_net65279), .ZN(u5_mult_82_ab_47__36_) );
  NOR2_X1 u5_mult_82_U7788 ( .A1(u5_mult_82_net64913), .A2(u5_mult_82_n6747), 
        .ZN(u5_mult_82_ab_48__35_) );
  NAND3_X2 u5_mult_82_U7787 ( .A1(u5_mult_82_n3105), .A2(u5_mult_82_n3106), 
        .A3(u5_mult_82_n3107), .ZN(u5_mult_82_CARRYB_19__47_) );
  NAND2_X2 u5_mult_82_U7786 ( .A1(u5_mult_82_ab_19__47_), .A2(
        u5_mult_82_CARRYB_18__47_), .ZN(u5_mult_82_n3106) );
  NAND3_X2 u5_mult_82_U7785 ( .A1(u5_mult_82_n3102), .A2(u5_mult_82_n3103), 
        .A3(u5_mult_82_n3104), .ZN(u5_mult_82_CARRYB_47__36_) );
  NAND2_X1 u5_mult_82_U7784 ( .A1(u5_mult_82_ab_47__36_), .A2(u5_mult_82_n5), 
        .ZN(u5_mult_82_n3104) );
  NAND2_X2 u5_mult_82_U7783 ( .A1(u5_mult_82_ab_47__36_), .A2(
        u5_mult_82_CARRYB_46__36_), .ZN(u5_mult_82_n3103) );
  NAND2_X1 u5_mult_82_U7782 ( .A1(u5_mult_82_n5), .A2(
        u5_mult_82_CARRYB_46__36_), .ZN(u5_mult_82_n3102) );
  NAND3_X2 u5_mult_82_U7781 ( .A1(u5_mult_82_n3099), .A2(u5_mult_82_n3100), 
        .A3(u5_mult_82_n3101), .ZN(u5_mult_82_CARRYB_52__31_) );
  NAND2_X1 u5_mult_82_U7780 ( .A1(u5_mult_82_CARRYB_51__31_), .A2(
        u5_mult_82_SUMB_51__32_), .ZN(u5_mult_82_n3101) );
  NAND2_X1 u5_mult_82_U7779 ( .A1(u5_mult_82_ab_52__31_), .A2(
        u5_mult_82_SUMB_51__32_), .ZN(u5_mult_82_n3100) );
  NAND2_X1 u5_mult_82_U7778 ( .A1(u5_mult_82_ab_52__31_), .A2(
        u5_mult_82_CARRYB_51__31_), .ZN(u5_mult_82_n3099) );
  NAND3_X2 u5_mult_82_U7777 ( .A1(u5_mult_82_n3096), .A2(u5_mult_82_n3097), 
        .A3(u5_mult_82_n3098), .ZN(u5_mult_82_CARRYB_51__32_) );
  NAND2_X2 u5_mult_82_U7776 ( .A1(u5_mult_82_CARRYB_50__32_), .A2(
        u5_mult_82_n1749), .ZN(u5_mult_82_n3098) );
  NAND2_X2 u5_mult_82_U7775 ( .A1(u5_mult_82_ab_51__32_), .A2(u5_mult_82_n1749), .ZN(u5_mult_82_n3097) );
  NAND2_X1 u5_mult_82_U7774 ( .A1(u5_mult_82_ab_51__32_), .A2(
        u5_mult_82_CARRYB_50__32_), .ZN(u5_mult_82_n3096) );
  XOR2_X2 u5_mult_82_U7773 ( .A(u5_mult_82_n3095), .B(u5_mult_82_SUMB_51__32_), 
        .Z(u5_mult_82_SUMB_52__31_) );
  XOR2_X2 u5_mult_82_U7772 ( .A(u5_mult_82_ab_52__31_), .B(
        u5_mult_82_CARRYB_51__31_), .Z(u5_mult_82_n3095) );
  XOR2_X2 u5_mult_82_U7771 ( .A(u5_mult_82_n3094), .B(u5_mult_82_n1749), .Z(
        u5_mult_82_SUMB_51__32_) );
  XOR2_X2 u5_mult_82_U7770 ( .A(u5_mult_82_ab_51__32_), .B(
        u5_mult_82_CARRYB_50__32_), .Z(u5_mult_82_n3094) );
  NAND2_X1 u5_mult_82_U7769 ( .A1(u5_mult_82_ab_48__35_), .A2(
        u5_mult_82_CARRYB_47__35_), .ZN(u5_mult_82_n3093) );
  NOR2_X1 u5_mult_82_U7768 ( .A1(u5_mult_82_n6850), .A2(u5_mult_82_net65387), 
        .ZN(u5_mult_82_ab_41__31_) );
  NOR2_X1 u5_mult_82_U7767 ( .A1(u5_mult_82_n6851), .A2(u5_mult_82_net65405), 
        .ZN(u5_mult_82_ab_40__31_) );
  NOR2_X1 u5_mult_82_U7766 ( .A1(u5_mult_82_n6817), .A2(u5_mult_82_n6644), 
        .ZN(u5_mult_82_ab_24__42_) );
  NAND2_X1 u5_mult_82_U7765 ( .A1(u5_mult_82_ab_41__31_), .A2(
        u5_mult_82_CARRYB_40__31_), .ZN(u5_mult_82_n3090) );
  NAND3_X2 u5_mult_82_U7764 ( .A1(u5_mult_82_n3085), .A2(u5_mult_82_n3086), 
        .A3(u5_mult_82_n3087), .ZN(u5_mult_82_CARRYB_40__31_) );
  NAND2_X1 u5_mult_82_U7763 ( .A1(u5_mult_82_ab_40__31_), .A2(
        u5_mult_82_CARRYB_39__31_), .ZN(u5_mult_82_n3087) );
  NAND3_X2 u5_mult_82_U7762 ( .A1(u5_mult_82_n3082), .A2(u5_mult_82_n3083), 
        .A3(u5_mult_82_n3084), .ZN(u5_mult_82_CARRYB_26__40_) );
  NAND2_X1 u5_mult_82_U7761 ( .A1(u5_mult_82_n2174), .A2(
        u5_mult_82_SUMB_25__41_), .ZN(u5_mult_82_n3084) );
  NAND2_X1 u5_mult_82_U7760 ( .A1(u5_mult_82_ab_26__40_), .A2(
        u5_mult_82_SUMB_25__41_), .ZN(u5_mult_82_n3083) );
  NAND2_X1 u5_mult_82_U7759 ( .A1(u5_mult_82_ab_26__40_), .A2(u5_mult_82_n2174), .ZN(u5_mult_82_n3082) );
  NAND3_X2 u5_mult_82_U7758 ( .A1(u5_mult_82_n3079), .A2(u5_mult_82_n3080), 
        .A3(u5_mult_82_n3081), .ZN(u5_mult_82_CARRYB_25__41_) );
  NAND2_X2 u5_mult_82_U7757 ( .A1(u5_mult_82_CARRYB_24__41_), .A2(
        u5_mult_82_SUMB_24__42_), .ZN(u5_mult_82_n3081) );
  NAND2_X2 u5_mult_82_U7756 ( .A1(u5_mult_82_ab_25__41_), .A2(
        u5_mult_82_SUMB_24__42_), .ZN(u5_mult_82_n3080) );
  NAND3_X2 u5_mult_82_U7755 ( .A1(u5_mult_82_n3076), .A2(u5_mult_82_n3077), 
        .A3(u5_mult_82_n3078), .ZN(u5_mult_82_CARRYB_24__42_) );
  NAND2_X2 u5_mult_82_U7754 ( .A1(u5_mult_82_ab_24__42_), .A2(
        u5_mult_82_CARRYB_23__42_), .ZN(u5_mult_82_n3078) );
  NAND2_X2 u5_mult_82_U7753 ( .A1(u5_mult_82_ab_24__42_), .A2(
        u5_mult_82_SUMB_23__43_), .ZN(u5_mult_82_n3077) );
  XNOR2_X2 u5_mult_82_U7752 ( .A(u5_mult_82_CARRYB_37__16_), .B(
        u5_mult_82_ab_38__16_), .ZN(u5_mult_82_n3075) );
  XNOR2_X2 u5_mult_82_U7751 ( .A(u5_mult_82_SUMB_37__17_), .B(u5_mult_82_n3075), .ZN(u5_mult_82_SUMB_38__16_) );
  XOR2_X2 u5_mult_82_U7750 ( .A(u5_mult_82_ab_41__23_), .B(
        u5_mult_82_CARRYB_40__23_), .Z(u5_mult_82_n3856) );
  INV_X4 u5_mult_82_U7749 ( .A(u5_mult_82_n3073), .ZN(u5_mult_82_n3074) );
  INV_X2 u5_mult_82_U7748 ( .A(u5_mult_82_CARRYB_28__21_), .ZN(
        u5_mult_82_n3073) );
  NOR2_X1 u5_mult_82_U7747 ( .A1(u5_mult_82_n6842), .A2(u5_mult_82_net65369), 
        .ZN(u5_mult_82_ab_42__32_) );
  NAND3_X2 u5_mult_82_U7746 ( .A1(u5_mult_82_n3070), .A2(u5_mult_82_n3071), 
        .A3(u5_mult_82_n3072), .ZN(u5_mult_82_CARRYB_46__28_) );
  NAND2_X1 u5_mult_82_U7745 ( .A1(u5_mult_82_CARRYB_45__28_), .A2(
        u5_mult_82_SUMB_45__29_), .ZN(u5_mult_82_n3072) );
  NAND2_X1 u5_mult_82_U7744 ( .A1(u5_mult_82_ab_46__28_), .A2(
        u5_mult_82_SUMB_45__29_), .ZN(u5_mult_82_n3071) );
  NAND2_X1 u5_mult_82_U7743 ( .A1(u5_mult_82_ab_46__28_), .A2(
        u5_mult_82_CARRYB_45__28_), .ZN(u5_mult_82_n3070) );
  NAND3_X4 u5_mult_82_U7742 ( .A1(u5_mult_82_n3069), .A2(u5_mult_82_n3068), 
        .A3(u5_mult_82_n3067), .ZN(u5_mult_82_CARRYB_45__29_) );
  NAND2_X2 u5_mult_82_U7741 ( .A1(u5_mult_82_n1700), .A2(u5_mult_82_n1594), 
        .ZN(u5_mult_82_n3069) );
  NAND2_X2 u5_mult_82_U7740 ( .A1(u5_mult_82_ab_45__29_), .A2(u5_mult_82_n1594), .ZN(u5_mult_82_n3068) );
  NAND2_X1 u5_mult_82_U7739 ( .A1(u5_mult_82_ab_45__29_), .A2(
        u5_mult_82_CARRYB_44__29_), .ZN(u5_mult_82_n3067) );
  XOR2_X2 u5_mult_82_U7738 ( .A(u5_mult_82_n3066), .B(u5_mult_82_SUMB_45__29_), 
        .Z(u5_mult_82_SUMB_46__28_) );
  NAND3_X2 u5_mult_82_U7737 ( .A1(u5_mult_82_n3063), .A2(u5_mult_82_n3064), 
        .A3(u5_mult_82_n3065), .ZN(u5_mult_82_CARRYB_42__32_) );
  NAND2_X1 u5_mult_82_U7736 ( .A1(u5_mult_82_ab_42__32_), .A2(
        u5_mult_82_CARRYB_41__32_), .ZN(u5_mult_82_n3065) );
  NAND2_X2 u5_mult_82_U7735 ( .A1(u5_mult_82_ab_42__32_), .A2(
        u5_mult_82_SUMB_41__33_), .ZN(u5_mult_82_n3064) );
  NAND2_X1 u5_mult_82_U7734 ( .A1(u5_mult_82_CARRYB_41__32_), .A2(
        u5_mult_82_SUMB_41__33_), .ZN(u5_mult_82_n3063) );
  XOR2_X2 u5_mult_82_U7733 ( .A(u5_mult_82_SUMB_41__33_), .B(u5_mult_82_n3062), 
        .Z(u5_mult_82_SUMB_42__32_) );
  XOR2_X2 u5_mult_82_U7732 ( .A(u5_mult_82_CARRYB_41__32_), .B(
        u5_mult_82_ab_42__32_), .Z(u5_mult_82_n3062) );
  NAND2_X2 u5_mult_82_U7731 ( .A1(u5_mult_82_ab_18__25_), .A2(
        u5_mult_82_SUMB_17__26_), .ZN(u5_mult_82_n4778) );
  NAND3_X2 u5_mult_82_U7730 ( .A1(u5_mult_82_n5243), .A2(u5_mult_82_n5245), 
        .A3(u5_mult_82_n5244), .ZN(u5_mult_82_CARRYB_43__5_) );
  XOR2_X2 u5_mult_82_U7729 ( .A(u5_mult_82_ab_10__27_), .B(
        u5_mult_82_CARRYB_9__27_), .Z(u5_mult_82_n3445) );
  XNOR2_X2 u5_mult_82_U7728 ( .A(u5_mult_82_n3061), .B(
        u5_mult_82_CARRYB_48__11_), .ZN(u5_mult_82_n6107) );
  XNOR2_X2 u5_mult_82_U7727 ( .A(u5_mult_82_n3443), .B(u5_mult_82_SUMB_29__31_), .ZN(u5_mult_82_SUMB_30__30_) );
  NAND2_X1 u5_mult_82_U7726 ( .A1(u5_mult_82_ab_42__6_), .A2(
        u5_mult_82_CARRYB_41__6_), .ZN(u5_mult_82_n6006) );
  XNOR2_X2 u5_mult_82_U7725 ( .A(u5_mult_82_ab_28__23_), .B(
        u5_mult_82_CARRYB_27__23_), .ZN(u5_mult_82_n3154) );
  XNOR2_X2 u5_mult_82_U7724 ( .A(u5_mult_82_ab_27__23_), .B(
        u5_mult_82_CARRYB_26__23_), .ZN(u5_mult_82_n3060) );
  XNOR2_X2 u5_mult_82_U7723 ( .A(u5_mult_82_ab_42__6_), .B(
        u5_mult_82_CARRYB_41__6_), .ZN(u5_mult_82_n3591) );
  NOR2_X1 u5_mult_82_U7722 ( .A1(u5_mult_82_net64687), .A2(u5_mult_82_n6643), 
        .ZN(u5_mult_82_ab_24__23_) );
  NOR2_X1 u5_mult_82_U7721 ( .A1(u5_mult_82_n6886), .A2(u5_mult_82_n6622), 
        .ZN(u5_mult_82_ab_20__25_) );
  NAND2_X1 u5_mult_82_U7720 ( .A1(u5_mult_82_ab_20__25_), .A2(
        u5_mult_82_CARRYB_19__25_), .ZN(u5_mult_82_n3057) );
  XNOR2_X2 u5_mult_82_U7719 ( .A(u5_mult_82_CARRYB_33__7_), .B(
        u5_mult_82_ab_34__7_), .ZN(u5_mult_82_n3056) );
  XNOR2_X2 u5_mult_82_U7718 ( .A(u5_mult_82_ab_48__11_), .B(
        u5_mult_82_CARRYB_47__11_), .ZN(u5_mult_82_n3498) );
  NAND3_X4 u5_mult_82_U7717 ( .A1(u5_mult_82_n3757), .A2(u5_mult_82_n3758), 
        .A3(u5_mult_82_n3759), .ZN(u5_mult_82_CARRYB_48__29_) );
  XNOR2_X2 u5_mult_82_U7716 ( .A(u5_mult_82_SUMB_18__48_), .B(
        u5_mult_82_ab_19__47_), .ZN(u5_mult_82_n3055) );
  XNOR2_X2 u5_mult_82_U7715 ( .A(u5_mult_82_CARRYB_18__47_), .B(
        u5_mult_82_n3055), .ZN(u5_mult_82_SUMB_19__47_) );
  NAND2_X2 u5_mult_82_U7714 ( .A1(u5_mult_82_ab_46__19_), .A2(
        u5_mult_82_SUMB_45__20_), .ZN(u5_mult_82_n3849) );
  NAND2_X2 u5_mult_82_U7713 ( .A1(u5_mult_82_ab_48__18_), .A2(
        u5_mult_82_SUMB_47__19_), .ZN(u5_mult_82_n5713) );
  NOR2_X2 u5_mult_82_U7712 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6714), 
        .ZN(u5_mult_82_ab_36__38_) );
  NAND2_X4 u5_mult_82_U7711 ( .A1(u5_mult_82_ab_38__37_), .A2(
        u5_mult_82_CARRYB_37__37_), .ZN(u5_mult_82_n4472) );
  NOR2_X2 u5_mult_82_U7710 ( .A1(u5_mult_82_net64937), .A2(u5_mult_82_n6720), 
        .ZN(u5_mult_82_ab_37__37_) );
  NAND2_X2 u5_mult_82_U7709 ( .A1(u5_mult_82_ab_36__38_), .A2(
        u5_mult_82_SUMB_35__39_), .ZN(u5_mult_82_n3054) );
  NAND2_X2 u5_mult_82_U7708 ( .A1(u5_mult_82_ab_36__38_), .A2(
        u5_mult_82_CARRYB_35__38_), .ZN(u5_mult_82_n3053) );
  NAND2_X2 u5_mult_82_U7707 ( .A1(u5_mult_82_SUMB_35__39_), .A2(
        u5_mult_82_CARRYB_35__38_), .ZN(u5_mult_82_n3052) );
  XOR2_X2 u5_mult_82_U7706 ( .A(u5_mult_82_CARRYB_35__38_), .B(
        u5_mult_82_n3051), .Z(u5_mult_82_SUMB_36__38_) );
  XOR2_X2 u5_mult_82_U7705 ( .A(u5_mult_82_SUMB_35__39_), .B(
        u5_mult_82_ab_36__38_), .Z(u5_mult_82_n3051) );
  NAND3_X4 u5_mult_82_U7704 ( .A1(u5_mult_82_n3048), .A2(u5_mult_82_n3049), 
        .A3(u5_mult_82_n3050), .ZN(u5_mult_82_CARRYB_37__37_) );
  NAND2_X2 u5_mult_82_U7703 ( .A1(u5_mult_82_ab_37__37_), .A2(
        u5_mult_82_CARRYB_36__37_), .ZN(u5_mult_82_n3050) );
  NAND2_X2 u5_mult_82_U7702 ( .A1(u5_mult_82_ab_37__37_), .A2(
        u5_mult_82_SUMB_36__38_), .ZN(u5_mult_82_n3049) );
  NAND2_X2 u5_mult_82_U7701 ( .A1(u5_mult_82_CARRYB_36__37_), .A2(
        u5_mult_82_SUMB_36__38_), .ZN(u5_mult_82_n3048) );
  XOR2_X2 u5_mult_82_U7700 ( .A(u5_mult_82_CARRYB_40__16_), .B(
        u5_mult_82_ab_41__16_), .Z(u5_mult_82_n5293) );
  NOR2_X1 u5_mult_82_U7699 ( .A1(u5_mult_82_net64881), .A2(u5_mult_82_net65369), .ZN(u5_mult_82_ab_42__34_) );
  NAND3_X2 u5_mult_82_U7698 ( .A1(u5_mult_82_n3045), .A2(u5_mult_82_n3046), 
        .A3(u5_mult_82_n3047), .ZN(u5_mult_82_CARRYB_42__34_) );
  NAND2_X1 u5_mult_82_U7697 ( .A1(u5_mult_82_ab_42__34_), .A2(
        u5_mult_82_SUMB_41__35_), .ZN(u5_mult_82_n3047) );
  NAND2_X2 u5_mult_82_U7696 ( .A1(u5_mult_82_ab_42__34_), .A2(
        u5_mult_82_CARRYB_41__34_), .ZN(u5_mult_82_n3046) );
  NAND2_X1 u5_mult_82_U7695 ( .A1(u5_mult_82_SUMB_41__35_), .A2(
        u5_mult_82_CARRYB_41__34_), .ZN(u5_mult_82_n3045) );
  XOR2_X2 u5_mult_82_U7694 ( .A(u5_mult_82_CARRYB_41__34_), .B(
        u5_mult_82_n3044), .Z(u5_mult_82_SUMB_42__34_) );
  XOR2_X2 u5_mult_82_U7693 ( .A(u5_mult_82_SUMB_41__35_), .B(
        u5_mult_82_ab_42__34_), .Z(u5_mult_82_n3044) );
  NAND3_X4 u5_mult_82_U7692 ( .A1(u5_mult_82_n3041), .A2(u5_mult_82_n3042), 
        .A3(u5_mult_82_n3043), .ZN(u5_mult_82_CARRYB_44__32_) );
  NAND2_X1 u5_mult_82_U7691 ( .A1(u5_mult_82_CARRYB_43__32_), .A2(
        u5_mult_82_SUMB_43__33_), .ZN(u5_mult_82_n3043) );
  NAND2_X1 u5_mult_82_U7690 ( .A1(u5_mult_82_ab_44__32_), .A2(
        u5_mult_82_SUMB_43__33_), .ZN(u5_mult_82_n3042) );
  NAND2_X1 u5_mult_82_U7689 ( .A1(u5_mult_82_ab_44__32_), .A2(
        u5_mult_82_CARRYB_43__32_), .ZN(u5_mult_82_n3041) );
  NAND2_X1 u5_mult_82_U7688 ( .A1(u5_mult_82_ab_43__33_), .A2(
        u5_mult_82_CARRYB_42__33_), .ZN(u5_mult_82_n3038) );
  XOR2_X2 u5_mult_82_U7687 ( .A(u5_mult_82_n3037), .B(u5_mult_82_SUMB_42__34_), 
        .Z(u5_mult_82_SUMB_43__33_) );
  XOR2_X2 u5_mult_82_U7686 ( .A(u5_mult_82_ab_43__33_), .B(
        u5_mult_82_CARRYB_42__33_), .Z(u5_mult_82_n3037) );
  NOR2_X1 u5_mult_82_U7685 ( .A1(u5_mult_82_n6822), .A2(u5_mult_82_net65717), 
        .ZN(u5_mult_82_ab_23__41_) );
  NAND3_X2 u5_mult_82_U7684 ( .A1(u5_mult_82_n3034), .A2(u5_mult_82_n3035), 
        .A3(u5_mult_82_n3036), .ZN(u5_mult_82_CARRYB_25__39_) );
  NAND2_X1 u5_mult_82_U7683 ( .A1(u5_mult_82_ab_25__39_), .A2(
        u5_mult_82_SUMB_24__40_), .ZN(u5_mult_82_n3035) );
  NAND2_X1 u5_mult_82_U7682 ( .A1(u5_mult_82_ab_25__39_), .A2(
        u5_mult_82_CARRYB_24__39_), .ZN(u5_mult_82_n3034) );
  NAND2_X2 u5_mult_82_U7681 ( .A1(u5_mult_82_ab_24__40_), .A2(
        u5_mult_82_SUMB_23__41_), .ZN(u5_mult_82_n3033) );
  NAND2_X1 u5_mult_82_U7680 ( .A1(u5_mult_82_CARRYB_23__40_), .A2(
        u5_mult_82_ab_24__40_), .ZN(u5_mult_82_n3031) );
  XOR2_X2 u5_mult_82_U7679 ( .A(u5_mult_82_n3030), .B(u5_mult_82_SUMB_23__41_), 
        .Z(u5_mult_82_SUMB_24__40_) );
  XOR2_X2 u5_mult_82_U7678 ( .A(u5_mult_82_CARRYB_23__40_), .B(
        u5_mult_82_ab_24__40_), .Z(u5_mult_82_n3030) );
  NAND2_X1 u5_mult_82_U7677 ( .A1(u5_mult_82_ab_23__41_), .A2(
        u5_mult_82_CARRYB_22__41_), .ZN(u5_mult_82_n3029) );
  NAND2_X2 u5_mult_82_U7676 ( .A1(u5_mult_82_ab_23__41_), .A2(
        u5_mult_82_SUMB_22__42_), .ZN(u5_mult_82_n3028) );
  NAND3_X4 u5_mult_82_U7675 ( .A1(u5_mult_82_n3024), .A2(u5_mult_82_n3025), 
        .A3(u5_mult_82_n3026), .ZN(u5_mult_82_CARRYB_45__30_) );
  NAND2_X1 u5_mult_82_U7674 ( .A1(u5_mult_82_CARRYB_44__30_), .A2(
        u5_mult_82_SUMB_44__31_), .ZN(u5_mult_82_n3026) );
  NAND2_X1 u5_mult_82_U7673 ( .A1(u5_mult_82_ab_45__30_), .A2(
        u5_mult_82_SUMB_44__31_), .ZN(u5_mult_82_n3025) );
  NAND2_X1 u5_mult_82_U7672 ( .A1(u5_mult_82_ab_45__30_), .A2(
        u5_mult_82_CARRYB_44__30_), .ZN(u5_mult_82_n3024) );
  NAND3_X2 u5_mult_82_U7671 ( .A1(u5_mult_82_n3023), .A2(u5_mult_82_n3022), 
        .A3(u5_mult_82_n3021), .ZN(u5_mult_82_CARRYB_44__31_) );
  NAND2_X2 u5_mult_82_U7670 ( .A1(u5_mult_82_SUMB_43__32_), .A2(
        u5_mult_82_ab_44__31_), .ZN(u5_mult_82_n3022) );
  NAND2_X1 u5_mult_82_U7669 ( .A1(u5_mult_82_ab_44__31_), .A2(
        u5_mult_82_CARRYB_43__31_), .ZN(u5_mult_82_n3021) );
  XOR2_X2 u5_mult_82_U7668 ( .A(u5_mult_82_n3020), .B(u5_mult_82_SUMB_44__31_), 
        .Z(u5_mult_82_SUMB_45__30_) );
  XOR2_X2 u5_mult_82_U7667 ( .A(u5_mult_82_SUMB_43__32_), .B(u5_mult_82_n3019), 
        .Z(u5_mult_82_SUMB_44__31_) );
  XNOR2_X2 u5_mult_82_U7666 ( .A(u5_mult_82_CARRYB_5__46_), .B(
        u5_mult_82_ab_6__46_), .ZN(u5_mult_82_n3279) );
  NAND2_X1 u5_mult_82_U7665 ( .A1(u5_mult_82_CARRYB_40__23_), .A2(
        u5_mult_82_SUMB_40__24_), .ZN(u5_mult_82_n3862) );
  NAND2_X2 u5_mult_82_U7664 ( .A1(u5_mult_82_n407), .A2(
        u5_mult_82_SUMB_49__19_), .ZN(u5_mult_82_n5741) );
  NOR2_X1 u5_mult_82_U7663 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6742), 
        .ZN(u5_mult_82_ab_46__36_) );
  NOR2_X1 u5_mult_82_U7662 ( .A1(u5_mult_82_n6831), .A2(u5_mult_82_net65351), 
        .ZN(u5_mult_82_ab_43__39_) );
  NAND3_X2 u5_mult_82_U7661 ( .A1(u5_mult_82_n3016), .A2(u5_mult_82_n3017), 
        .A3(u5_mult_82_n3018), .ZN(u5_mult_82_CARRYB_46__36_) );
  NAND2_X1 u5_mult_82_U7660 ( .A1(u5_mult_82_ab_46__36_), .A2(
        u5_mult_82_CARRYB_45__36_), .ZN(u5_mult_82_n3018) );
  NAND2_X2 u5_mult_82_U7659 ( .A1(u5_mult_82_ab_46__36_), .A2(
        u5_mult_82_SUMB_45__37_), .ZN(u5_mult_82_n3017) );
  NAND2_X1 u5_mult_82_U7658 ( .A1(u5_mult_82_CARRYB_45__36_), .A2(
        u5_mult_82_SUMB_45__37_), .ZN(u5_mult_82_n3016) );
  NAND3_X2 u5_mult_82_U7657 ( .A1(u5_mult_82_n3013), .A2(u5_mult_82_n3014), 
        .A3(u5_mult_82_n3015), .ZN(u5_mult_82_CARRYB_43__39_) );
  NAND2_X1 u5_mult_82_U7656 ( .A1(u5_mult_82_ab_43__39_), .A2(u5_mult_82_n1412), .ZN(u5_mult_82_n3015) );
  NAND2_X2 u5_mult_82_U7655 ( .A1(u5_mult_82_ab_43__39_), .A2(
        u5_mult_82_SUMB_42__40_), .ZN(u5_mult_82_n3014) );
  NAND2_X1 u5_mult_82_U7654 ( .A1(u5_mult_82_n1412), .A2(
        u5_mult_82_SUMB_42__40_), .ZN(u5_mult_82_n3013) );
  XOR2_X2 u5_mult_82_U7653 ( .A(u5_mult_82_SUMB_42__40_), .B(u5_mult_82_n3012), 
        .Z(u5_mult_82_SUMB_43__39_) );
  XOR2_X2 u5_mult_82_U7652 ( .A(u5_mult_82_CARRYB_42__39_), .B(
        u5_mult_82_ab_43__39_), .Z(u5_mult_82_n3012) );
  NAND3_X2 u5_mult_82_U7651 ( .A1(u5_mult_82_n3009), .A2(u5_mult_82_n3010), 
        .A3(u5_mult_82_n3011), .ZN(u5_mult_82_CARRYB_49__33_) );
  NAND2_X1 u5_mult_82_U7650 ( .A1(u5_mult_82_CARRYB_48__33_), .A2(
        u5_mult_82_SUMB_48__34_), .ZN(u5_mult_82_n3011) );
  NAND2_X1 u5_mult_82_U7649 ( .A1(u5_mult_82_ab_49__33_), .A2(
        u5_mult_82_SUMB_48__34_), .ZN(u5_mult_82_n3010) );
  NAND2_X1 u5_mult_82_U7648 ( .A1(u5_mult_82_ab_49__33_), .A2(
        u5_mult_82_CARRYB_48__33_), .ZN(u5_mult_82_n3009) );
  NAND2_X2 u5_mult_82_U7647 ( .A1(u5_mult_82_CARRYB_47__34_), .A2(
        u5_mult_82_n1581), .ZN(u5_mult_82_n3008) );
  NAND2_X2 u5_mult_82_U7646 ( .A1(u5_mult_82_ab_48__34_), .A2(u5_mult_82_n1581), .ZN(u5_mult_82_n3007) );
  NAND2_X1 u5_mult_82_U7645 ( .A1(u5_mult_82_ab_48__34_), .A2(
        u5_mult_82_CARRYB_47__34_), .ZN(u5_mult_82_n3006) );
  XOR2_X2 u5_mult_82_U7644 ( .A(u5_mult_82_n3005), .B(u5_mult_82_n1581), .Z(
        u5_mult_82_SUMB_48__34_) );
  XOR2_X2 u5_mult_82_U7643 ( .A(u5_mult_82_ab_48__34_), .B(
        u5_mult_82_CARRYB_47__34_), .Z(u5_mult_82_n3005) );
  NAND2_X1 u5_mult_82_U7642 ( .A1(u5_mult_82_ab_42__29_), .A2(
        u5_mult_82_SUMB_41__30_), .ZN(u5_mult_82_n4423) );
  XNOR2_X2 u5_mult_82_U7641 ( .A(u5_mult_82_ab_45__5_), .B(
        u5_mult_82_CARRYB_44__5_), .ZN(u5_mult_82_n3749) );
  NAND3_X2 u5_mult_82_U7640 ( .A1(u5_mult_82_n3002), .A2(u5_mult_82_n3003), 
        .A3(u5_mult_82_n3004), .ZN(u5_mult_82_CARRYB_48__36_) );
  NAND2_X1 u5_mult_82_U7639 ( .A1(u5_mult_82_ab_48__36_), .A2(
        u5_mult_82_SUMB_47__37_), .ZN(u5_mult_82_n3003) );
  NAND2_X1 u5_mult_82_U7638 ( .A1(u5_mult_82_ab_48__36_), .A2(
        u5_mult_82_CARRYB_47__36_), .ZN(u5_mult_82_n3002) );
  NAND2_X2 u5_mult_82_U7637 ( .A1(u5_mult_82_CARRYB_46__37_), .A2(
        u5_mult_82_SUMB_46__38_), .ZN(u5_mult_82_n3001) );
  NAND2_X1 u5_mult_82_U7636 ( .A1(u5_mult_82_ab_47__37_), .A2(
        u5_mult_82_CARRYB_46__37_), .ZN(u5_mult_82_n2999) );
  XOR2_X2 u5_mult_82_U7635 ( .A(u5_mult_82_n2998), .B(u5_mult_82_SUMB_46__38_), 
        .Z(u5_mult_82_SUMB_47__37_) );
  XOR2_X2 u5_mult_82_U7634 ( .A(u5_mult_82_ab_47__37_), .B(
        u5_mult_82_CARRYB_46__37_), .Z(u5_mult_82_n2998) );
  XNOR2_X2 u5_mult_82_U7633 ( .A(u5_mult_82_ab_44__32_), .B(
        u5_mult_82_CARRYB_43__32_), .ZN(u5_mult_82_n2997) );
  XNOR2_X2 u5_mult_82_U7632 ( .A(u5_mult_82_n2997), .B(u5_mult_82_SUMB_43__33_), .ZN(u5_mult_82_SUMB_44__32_) );
  NAND2_X2 u5_mult_82_U7631 ( .A1(u5_mult_82_CARRYB_21__29_), .A2(
        u5_mult_82_SUMB_21__30_), .ZN(u5_mult_82_n4296) );
  NAND3_X4 u5_mult_82_U7630 ( .A1(u5_mult_82_n4777), .A2(u5_mult_82_n4778), 
        .A3(u5_mult_82_n4779), .ZN(u5_mult_82_CARRYB_18__25_) );
  NAND3_X4 u5_mult_82_U7629 ( .A1(u5_mult_82_n4296), .A2(u5_mult_82_n4295), 
        .A3(u5_mult_82_n4294), .ZN(u5_mult_82_CARRYB_22__29_) );
  NAND3_X2 u5_mult_82_U7628 ( .A1(u5_mult_82_n2994), .A2(u5_mult_82_n2995), 
        .A3(u5_mult_82_n2996), .ZN(u5_mult_82_CARRYB_26__15_) );
  NAND2_X1 u5_mult_82_U7627 ( .A1(u5_mult_82_CARRYB_25__15_), .A2(
        u5_mult_82_SUMB_25__16_), .ZN(u5_mult_82_n2995) );
  NAND2_X2 u5_mult_82_U7626 ( .A1(u5_mult_82_CARRYB_24__16_), .A2(
        u5_mult_82_SUMB_24__17_), .ZN(u5_mult_82_n2993) );
  NAND2_X2 u5_mult_82_U7625 ( .A1(u5_mult_82_ab_25__16_), .A2(
        u5_mult_82_SUMB_24__17_), .ZN(u5_mult_82_n2992) );
  NAND2_X2 u5_mult_82_U7624 ( .A1(u5_mult_82_ab_25__16_), .A2(
        u5_mult_82_CARRYB_24__16_), .ZN(u5_mult_82_n2991) );
  XOR2_X2 u5_mult_82_U7623 ( .A(u5_mult_82_n2990), .B(u5_mult_82_SUMB_24__17_), 
        .Z(u5_mult_82_SUMB_25__16_) );
  NAND2_X1 u5_mult_82_U7622 ( .A1(u5_mult_82_ab_39__7_), .A2(
        u5_mult_82_CARRYB_38__7_), .ZN(u5_mult_82_n2987) );
  NAND3_X2 u5_mult_82_U7621 ( .A1(u5_mult_82_n2984), .A2(u5_mult_82_n2985), 
        .A3(u5_mult_82_n2986), .ZN(u5_mult_82_CARRYB_38__8_) );
  NAND2_X2 u5_mult_82_U7620 ( .A1(u5_mult_82_ab_38__8_), .A2(
        u5_mult_82_SUMB_37__9_), .ZN(u5_mult_82_n2985) );
  NAND2_X4 u5_mult_82_U7619 ( .A1(u5_mult_82_n2981), .A2(u5_mult_82_ab_41__6_), 
        .ZN(u5_mult_82_n2983) );
  NAND2_X2 u5_mult_82_U7618 ( .A1(u5_mult_82_CARRYB_40__6_), .A2(
        u5_mult_82_n4788), .ZN(u5_mult_82_n2982) );
  NAND2_X4 u5_mult_82_U7617 ( .A1(u5_mult_82_ab_44__4_), .A2(u5_mult_82_n2978), 
        .ZN(u5_mult_82_n2980) );
  NAND2_X1 u5_mult_82_U7616 ( .A1(u5_mult_82_n3992), .A2(
        u5_mult_82_CARRYB_43__4_), .ZN(u5_mult_82_n2979) );
  NAND2_X1 u5_mult_82_U7615 ( .A1(u5_mult_82_ab_20__27_), .A2(
        u5_mult_82_SUMB_19__28_), .ZN(u5_mult_82_n5925) );
  NAND2_X1 u5_mult_82_U7614 ( .A1(u5_mult_82_CARRYB_19__27_), .A2(
        u5_mult_82_SUMB_19__28_), .ZN(u5_mult_82_n5926) );
  NAND3_X2 u5_mult_82_U7613 ( .A1(u5_mult_82_n6206), .A2(u5_mult_82_n6207), 
        .A3(u5_mult_82_n6208), .ZN(u5_mult_82_CARRYB_47__11_) );
  XOR2_X2 u5_mult_82_U7612 ( .A(u5_mult_82_CARRYB_38__25_), .B(
        u5_mult_82_ab_39__25_), .Z(u5_mult_82_n3851) );
  XOR2_X2 u5_mult_82_U7611 ( .A(u5_mult_82_SUMB_43__24_), .B(u5_mult_82_n3915), 
        .Z(u5_mult_82_SUMB_44__23_) );
  XNOR2_X2 u5_mult_82_U7610 ( .A(u5_mult_82_ab_49__33_), .B(
        u5_mult_82_CARRYB_48__33_), .ZN(u5_mult_82_n2977) );
  XNOR2_X2 u5_mult_82_U7609 ( .A(u5_mult_82_n2977), .B(u5_mult_82_SUMB_48__34_), .ZN(u5_mult_82_SUMB_49__33_) );
  NOR2_X1 u5_mult_82_U7608 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_net65387), .ZN(u5_mult_82_ab_41__36_) );
  NAND3_X2 u5_mult_82_U7607 ( .A1(u5_mult_82_n2974), .A2(u5_mult_82_n2976), 
        .A3(u5_mult_82_n2975), .ZN(u5_mult_82_CARRYB_41__36_) );
  NAND2_X1 u5_mult_82_U7606 ( .A1(u5_mult_82_ab_41__36_), .A2(
        u5_mult_82_CARRYB_40__36_), .ZN(u5_mult_82_n2976) );
  NAND2_X1 u5_mult_82_U7605 ( .A1(u5_mult_82_CARRYB_40__36_), .A2(
        u5_mult_82_SUMB_40__37_), .ZN(u5_mult_82_n2974) );
  XOR2_X2 u5_mult_82_U7604 ( .A(u5_mult_82_SUMB_40__37_), .B(u5_mult_82_n2973), 
        .Z(u5_mult_82_SUMB_41__36_) );
  XOR2_X2 u5_mult_82_U7603 ( .A(u5_mult_82_CARRYB_40__36_), .B(
        u5_mult_82_ab_41__36_), .Z(u5_mult_82_n2973) );
  NAND3_X2 u5_mult_82_U7602 ( .A1(u5_mult_82_n2970), .A2(u5_mult_82_n2971), 
        .A3(u5_mult_82_n2972), .ZN(u5_mult_82_CARRYB_38__39_) );
  NAND2_X1 u5_mult_82_U7601 ( .A1(u5_mult_82_SUMB_37__40_), .A2(
        u5_mult_82_CARRYB_37__39_), .ZN(u5_mult_82_n2972) );
  NAND2_X1 u5_mult_82_U7600 ( .A1(u5_mult_82_ab_38__39_), .A2(
        u5_mult_82_SUMB_37__40_), .ZN(u5_mult_82_n2971) );
  NAND2_X1 u5_mult_82_U7599 ( .A1(u5_mult_82_ab_38__39_), .A2(
        u5_mult_82_CARRYB_37__39_), .ZN(u5_mult_82_n2970) );
  NAND3_X2 u5_mult_82_U7598 ( .A1(u5_mult_82_n2967), .A2(u5_mult_82_n2968), 
        .A3(u5_mult_82_n2969), .ZN(u5_mult_82_CARRYB_37__40_) );
  NAND2_X2 u5_mult_82_U7597 ( .A1(u5_mult_82_CARRYB_36__40_), .A2(
        u5_mult_82_SUMB_36__41_), .ZN(u5_mult_82_n2969) );
  NAND2_X2 u5_mult_82_U7596 ( .A1(u5_mult_82_ab_37__40_), .A2(
        u5_mult_82_SUMB_36__41_), .ZN(u5_mult_82_n2968) );
  NAND2_X1 u5_mult_82_U7595 ( .A1(u5_mult_82_ab_37__40_), .A2(
        u5_mult_82_CARRYB_36__40_), .ZN(u5_mult_82_n2967) );
  XOR2_X2 u5_mult_82_U7594 ( .A(u5_mult_82_n2966), .B(u5_mult_82_SUMB_37__40_), 
        .Z(u5_mult_82_SUMB_38__39_) );
  XOR2_X2 u5_mult_82_U7593 ( .A(u5_mult_82_ab_38__39_), .B(
        u5_mult_82_CARRYB_37__39_), .Z(u5_mult_82_n2966) );
  XOR2_X2 u5_mult_82_U7592 ( .A(u5_mult_82_n2965), .B(u5_mult_82_SUMB_36__41_), 
        .Z(u5_mult_82_SUMB_37__40_) );
  XOR2_X2 u5_mult_82_U7591 ( .A(u5_mult_82_ab_37__40_), .B(
        u5_mult_82_CARRYB_36__40_), .Z(u5_mult_82_n2965) );
  NAND3_X2 u5_mult_82_U7590 ( .A1(u5_mult_82_n2962), .A2(u5_mult_82_n2963), 
        .A3(u5_mult_82_n2964), .ZN(u5_mult_82_CARRYB_48__31_) );
  NAND2_X1 u5_mult_82_U7589 ( .A1(u5_mult_82_CARRYB_47__31_), .A2(
        u5_mult_82_SUMB_47__32_), .ZN(u5_mult_82_n2964) );
  NAND2_X1 u5_mult_82_U7588 ( .A1(u5_mult_82_ab_48__31_), .A2(
        u5_mult_82_SUMB_47__32_), .ZN(u5_mult_82_n2963) );
  NAND2_X1 u5_mult_82_U7587 ( .A1(u5_mult_82_ab_48__31_), .A2(
        u5_mult_82_CARRYB_47__31_), .ZN(u5_mult_82_n2962) );
  NAND2_X2 u5_mult_82_U7586 ( .A1(u5_mult_82_CARRYB_46__32_), .A2(
        u5_mult_82_SUMB_46__33_), .ZN(u5_mult_82_n2961) );
  NAND2_X2 u5_mult_82_U7585 ( .A1(u5_mult_82_ab_47__32_), .A2(
        u5_mult_82_SUMB_46__33_), .ZN(u5_mult_82_n2960) );
  NAND2_X2 u5_mult_82_U7584 ( .A1(u5_mult_82_ab_47__32_), .A2(
        u5_mult_82_CARRYB_46__32_), .ZN(u5_mult_82_n2959) );
  NAND3_X2 u5_mult_82_U7583 ( .A1(u5_mult_82_n2955), .A2(u5_mult_82_n2956), 
        .A3(u5_mult_82_n2957), .ZN(u5_mult_82_CARRYB_52__27_) );
  NAND2_X1 u5_mult_82_U7582 ( .A1(u5_mult_82_CARRYB_51__27_), .A2(
        u5_mult_82_SUMB_51__28_), .ZN(u5_mult_82_n2957) );
  NAND2_X1 u5_mult_82_U7581 ( .A1(u5_mult_82_ab_52__27_), .A2(
        u5_mult_82_SUMB_51__28_), .ZN(u5_mult_82_n2956) );
  NAND2_X1 u5_mult_82_U7580 ( .A1(u5_mult_82_ab_52__27_), .A2(
        u5_mult_82_CARRYB_51__27_), .ZN(u5_mult_82_n2955) );
  NAND3_X2 u5_mult_82_U7579 ( .A1(u5_mult_82_n2952), .A2(u5_mult_82_n2953), 
        .A3(u5_mult_82_n2954), .ZN(u5_mult_82_CARRYB_51__28_) );
  NAND2_X2 u5_mult_82_U7578 ( .A1(u5_mult_82_CARRYB_50__28_), .A2(
        u5_mult_82_SUMB_50__29_), .ZN(u5_mult_82_n2954) );
  NAND2_X2 u5_mult_82_U7577 ( .A1(u5_mult_82_ab_51__28_), .A2(
        u5_mult_82_SUMB_50__29_), .ZN(u5_mult_82_n2953) );
  NAND2_X2 u5_mult_82_U7576 ( .A1(u5_mult_82_ab_51__28_), .A2(
        u5_mult_82_CARRYB_50__28_), .ZN(u5_mult_82_n2952) );
  XOR2_X2 u5_mult_82_U7575 ( .A(u5_mult_82_n2951), .B(u5_mult_82_SUMB_51__28_), 
        .Z(u5_mult_82_SUMB_52__27_) );
  XOR2_X2 u5_mult_82_U7574 ( .A(u5_mult_82_ab_52__27_), .B(
        u5_mult_82_CARRYB_51__27_), .Z(u5_mult_82_n2951) );
  XOR2_X1 u5_mult_82_U7573 ( .A(u5_mult_82_n2950), .B(u5_mult_82_SUMB_50__29_), 
        .Z(u5_mult_82_SUMB_51__28_) );
  XOR2_X2 u5_mult_82_U7572 ( .A(u5_mult_82_ab_51__28_), .B(
        u5_mult_82_CARRYB_50__28_), .Z(u5_mult_82_n2950) );
  NAND3_X2 u5_mult_82_U7571 ( .A1(u5_mult_82_n2947), .A2(u5_mult_82_n2948), 
        .A3(u5_mult_82_n2949), .ZN(u5_mult_82_CARRYB_25__45_) );
  NAND2_X1 u5_mult_82_U7570 ( .A1(u5_mult_82_CARRYB_24__45_), .A2(
        u5_mult_82_SUMB_24__46_), .ZN(u5_mult_82_n2949) );
  NAND2_X1 u5_mult_82_U7569 ( .A1(u5_mult_82_ab_25__45_), .A2(
        u5_mult_82_SUMB_24__46_), .ZN(u5_mult_82_n2948) );
  NAND2_X1 u5_mult_82_U7568 ( .A1(u5_mult_82_ab_25__45_), .A2(
        u5_mult_82_CARRYB_24__45_), .ZN(u5_mult_82_n2947) );
  NAND3_X2 u5_mult_82_U7567 ( .A1(u5_mult_82_n2944), .A2(u5_mult_82_n2945), 
        .A3(u5_mult_82_n2946), .ZN(u5_mult_82_CARRYB_24__46_) );
  NAND2_X2 u5_mult_82_U7566 ( .A1(u5_mult_82_ab_24__46_), .A2(
        u5_mult_82_SUMB_23__47_), .ZN(u5_mult_82_n2946) );
  NAND2_X2 u5_mult_82_U7565 ( .A1(u5_mult_82_CARRYB_23__46_), .A2(
        u5_mult_82_SUMB_23__47_), .ZN(u5_mult_82_n2945) );
  NAND2_X1 u5_mult_82_U7564 ( .A1(u5_mult_82_CARRYB_23__46_), .A2(
        u5_mult_82_ab_24__46_), .ZN(u5_mult_82_n2944) );
  XOR2_X2 u5_mult_82_U7563 ( .A(u5_mult_82_n2943), .B(u5_mult_82_n1598), .Z(
        u5_mult_82_SUMB_24__46_) );
  XOR2_X1 u5_mult_82_U7562 ( .A(u5_mult_82_CARRYB_23__46_), .B(
        u5_mult_82_ab_24__46_), .Z(u5_mult_82_n2943) );
  NAND3_X2 u5_mult_82_U7561 ( .A1(u5_mult_82_n2940), .A2(u5_mult_82_n2941), 
        .A3(u5_mult_82_n2942), .ZN(u5_mult_82_CARRYB_49__31_) );
  NAND2_X2 u5_mult_82_U7560 ( .A1(u5_mult_82_ab_49__31_), .A2(
        u5_mult_82_SUMB_48__32_), .ZN(u5_mult_82_n2941) );
  NAND2_X1 u5_mult_82_U7559 ( .A1(u5_mult_82_ab_49__31_), .A2(
        u5_mult_82_CARRYB_48__31_), .ZN(u5_mult_82_n2940) );
  NAND3_X2 u5_mult_82_U7558 ( .A1(u5_mult_82_n2937), .A2(u5_mult_82_n2938), 
        .A3(u5_mult_82_n2939), .ZN(u5_mult_82_CARRYB_48__32_) );
  NAND2_X2 u5_mult_82_U7557 ( .A1(u5_mult_82_CARRYB_47__32_), .A2(
        u5_mult_82_n2710), .ZN(u5_mult_82_n2939) );
  NAND2_X2 u5_mult_82_U7556 ( .A1(u5_mult_82_ab_48__32_), .A2(u5_mult_82_n2710), .ZN(u5_mult_82_n2938) );
  NAND2_X1 u5_mult_82_U7555 ( .A1(u5_mult_82_ab_48__32_), .A2(
        u5_mult_82_CARRYB_47__32_), .ZN(u5_mult_82_n2937) );
  XOR2_X2 u5_mult_82_U7554 ( .A(u5_mult_82_n2936), .B(u5_mult_82_SUMB_48__32_), 
        .Z(u5_mult_82_SUMB_49__31_) );
  XOR2_X2 u5_mult_82_U7553 ( .A(u5_mult_82_n2935), .B(u5_mult_82_n2710), .Z(
        u5_mult_82_SUMB_48__32_) );
  XOR2_X2 u5_mult_82_U7552 ( .A(u5_mult_82_ab_48__32_), .B(
        u5_mult_82_CARRYB_47__32_), .Z(u5_mult_82_n2935) );
  NOR2_X1 u5_mult_82_U7551 ( .A1(u5_mult_82_n6805), .A2(u5_mult_82_net65713), 
        .ZN(u5_mult_82_ab_23__44_) );
  NOR2_X1 u5_mult_82_U7550 ( .A1(u5_mult_82_n6792), .A2(u5_mult_82_n6628), 
        .ZN(u5_mult_82_ab_21__46_) );
  NOR2_X1 u5_mult_82_U7549 ( .A1(u5_mult_82_net64913), .A2(u5_mult_82_n6742), 
        .ZN(u5_mult_82_ab_46__35_) );
  NAND3_X2 u5_mult_82_U7548 ( .A1(u5_mult_82_n2932), .A2(u5_mult_82_n2933), 
        .A3(u5_mult_82_n2934), .ZN(u5_mult_82_CARRYB_23__44_) );
  NAND2_X1 u5_mult_82_U7547 ( .A1(u5_mult_82_ab_23__44_), .A2(
        u5_mult_82_CARRYB_22__44_), .ZN(u5_mult_82_n2934) );
  NAND2_X2 u5_mult_82_U7546 ( .A1(u5_mult_82_ab_23__44_), .A2(
        u5_mult_82_SUMB_22__45_), .ZN(u5_mult_82_n2933) );
  NAND2_X1 u5_mult_82_U7545 ( .A1(u5_mult_82_CARRYB_22__44_), .A2(
        u5_mult_82_SUMB_22__45_), .ZN(u5_mult_82_n2932) );
  XOR2_X2 u5_mult_82_U7544 ( .A(u5_mult_82_SUMB_22__45_), .B(u5_mult_82_n2931), 
        .Z(u5_mult_82_SUMB_23__44_) );
  XOR2_X2 u5_mult_82_U7543 ( .A(u5_mult_82_CARRYB_22__44_), .B(
        u5_mult_82_ab_23__44_), .Z(u5_mult_82_n2931) );
  NAND2_X2 u5_mult_82_U7542 ( .A1(u5_mult_82_ab_21__46_), .A2(
        u5_mult_82_CARRYB_20__46_), .ZN(u5_mult_82_n2929) );
  NAND2_X1 u5_mult_82_U7541 ( .A1(u5_mult_82_SUMB_20__47_), .A2(
        u5_mult_82_CARRYB_20__46_), .ZN(u5_mult_82_n2928) );
  XOR2_X2 u5_mult_82_U7540 ( .A(u5_mult_82_CARRYB_20__46_), .B(
        u5_mult_82_n2927), .Z(u5_mult_82_SUMB_21__46_) );
  NAND3_X2 u5_mult_82_U7539 ( .A1(u5_mult_82_n2924), .A2(u5_mult_82_n2925), 
        .A3(u5_mult_82_n2926), .ZN(u5_mult_82_CARRYB_48__33_) );
  NAND2_X1 u5_mult_82_U7538 ( .A1(u5_mult_82_CARRYB_47__33_), .A2(
        u5_mult_82_SUMB_47__34_), .ZN(u5_mult_82_n2926) );
  NAND2_X1 u5_mult_82_U7537 ( .A1(u5_mult_82_ab_48__33_), .A2(
        u5_mult_82_SUMB_47__34_), .ZN(u5_mult_82_n2925) );
  NAND2_X1 u5_mult_82_U7536 ( .A1(u5_mult_82_ab_48__33_), .A2(
        u5_mult_82_CARRYB_47__33_), .ZN(u5_mult_82_n2924) );
  NAND3_X2 u5_mult_82_U7535 ( .A1(u5_mult_82_n2921), .A2(u5_mult_82_n2922), 
        .A3(u5_mult_82_n2923), .ZN(u5_mult_82_CARRYB_47__34_) );
  NAND2_X2 u5_mult_82_U7534 ( .A1(u5_mult_82_CARRYB_46__34_), .A2(
        u5_mult_82_SUMB_46__35_), .ZN(u5_mult_82_n2923) );
  NAND2_X2 u5_mult_82_U7533 ( .A1(u5_mult_82_ab_47__34_), .A2(
        u5_mult_82_SUMB_46__35_), .ZN(u5_mult_82_n2922) );
  NAND2_X2 u5_mult_82_U7532 ( .A1(u5_mult_82_ab_47__34_), .A2(
        u5_mult_82_CARRYB_46__34_), .ZN(u5_mult_82_n2921) );
  XOR2_X2 u5_mult_82_U7531 ( .A(u5_mult_82_n2920), .B(u5_mult_82_SUMB_46__35_), 
        .Z(u5_mult_82_SUMB_47__34_) );
  NAND3_X2 u5_mult_82_U7530 ( .A1(u5_mult_82_n2917), .A2(u5_mult_82_n2918), 
        .A3(u5_mult_82_n2919), .ZN(u5_mult_82_CARRYB_46__35_) );
  NAND2_X1 u5_mult_82_U7529 ( .A1(u5_mult_82_ab_46__35_), .A2(
        u5_mult_82_CARRYB_45__35_), .ZN(u5_mult_82_n2919) );
  XOR2_X2 u5_mult_82_U7528 ( .A(u5_mult_82_n1570), .B(u5_mult_82_n2916), .Z(
        u5_mult_82_SUMB_46__35_) );
  XOR2_X2 u5_mult_82_U7527 ( .A(u5_mult_82_CARRYB_45__35_), .B(
        u5_mult_82_ab_46__35_), .Z(u5_mult_82_n2916) );
  XNOR2_X2 u5_mult_82_U7526 ( .A(u5_mult_82_ab_27__24_), .B(
        u5_mult_82_CARRYB_26__24_), .ZN(u5_mult_82_n2915) );
  XNOR2_X2 u5_mult_82_U7525 ( .A(u5_mult_82_n2915), .B(u5_mult_82_SUMB_26__25_), .ZN(u5_mult_82_SUMB_27__24_) );
  NAND3_X4 u5_mult_82_U7524 ( .A1(u5_mult_82_n5204), .A2(u5_mult_82_n5205), 
        .A3(u5_mult_82_n5206), .ZN(u5_mult_82_CARRYB_38__9_) );
  NAND3_X2 u5_mult_82_U7523 ( .A1(u5_mult_82_n2912), .A2(u5_mult_82_n2913), 
        .A3(u5_mult_82_n2914), .ZN(u5_mult_82_CARRYB_38__32_) );
  NAND2_X1 u5_mult_82_U7522 ( .A1(u5_mult_82_CARRYB_37__32_), .A2(
        u5_mult_82_SUMB_37__33_), .ZN(u5_mult_82_n2914) );
  NAND2_X1 u5_mult_82_U7521 ( .A1(u5_mult_82_ab_38__32_), .A2(
        u5_mult_82_SUMB_37__33_), .ZN(u5_mult_82_n2913) );
  NAND2_X1 u5_mult_82_U7520 ( .A1(u5_mult_82_ab_38__32_), .A2(
        u5_mult_82_CARRYB_37__32_), .ZN(u5_mult_82_n2912) );
  NAND3_X4 u5_mult_82_U7519 ( .A1(u5_mult_82_n2911), .A2(u5_mult_82_n2910), 
        .A3(u5_mult_82_n2909), .ZN(u5_mult_82_CARRYB_37__33_) );
  NAND2_X2 u5_mult_82_U7518 ( .A1(u5_mult_82_CARRYB_36__33_), .A2(
        u5_mult_82_SUMB_36__34_), .ZN(u5_mult_82_n2911) );
  NAND2_X2 u5_mult_82_U7517 ( .A1(u5_mult_82_ab_37__33_), .A2(
        u5_mult_82_SUMB_36__34_), .ZN(u5_mult_82_n2910) );
  NAND2_X1 u5_mult_82_U7516 ( .A1(u5_mult_82_ab_37__33_), .A2(
        u5_mult_82_CARRYB_36__33_), .ZN(u5_mult_82_n2909) );
  XOR2_X2 u5_mult_82_U7515 ( .A(u5_mult_82_n2908), .B(u5_mult_82_SUMB_37__33_), 
        .Z(u5_mult_82_SUMB_38__32_) );
  XOR2_X2 u5_mult_82_U7514 ( .A(u5_mult_82_ab_38__32_), .B(
        u5_mult_82_CARRYB_37__32_), .Z(u5_mult_82_n2908) );
  XOR2_X2 u5_mult_82_U7513 ( .A(u5_mult_82_n2907), .B(u5_mult_82_n443), .Z(
        u5_mult_82_SUMB_37__33_) );
  XOR2_X2 u5_mult_82_U7512 ( .A(u5_mult_82_ab_37__33_), .B(
        u5_mult_82_CARRYB_36__33_), .Z(u5_mult_82_n2907) );
  NAND2_X2 u5_mult_82_U7511 ( .A1(u5_mult_82_CARRYB_24__40_), .A2(
        u5_mult_82_SUMB_24__41_), .ZN(u5_mult_82_n2906) );
  NAND2_X2 u5_mult_82_U7510 ( .A1(u5_mult_82_ab_25__40_), .A2(
        u5_mult_82_SUMB_24__41_), .ZN(u5_mult_82_n2905) );
  NAND2_X1 u5_mult_82_U7509 ( .A1(u5_mult_82_ab_25__40_), .A2(
        u5_mult_82_CARRYB_24__40_), .ZN(u5_mult_82_n2904) );
  NAND2_X2 u5_mult_82_U7508 ( .A1(u5_mult_82_ab_24__41_), .A2(u5_mult_82_n1691), .ZN(u5_mult_82_n2902) );
  NAND2_X1 u5_mult_82_U7507 ( .A1(u5_mult_82_ab_24__41_), .A2(
        u5_mult_82_CARRYB_23__41_), .ZN(u5_mult_82_n2901) );
  XOR2_X2 u5_mult_82_U7506 ( .A(u5_mult_82_n2900), .B(u5_mult_82_SUMB_24__41_), 
        .Z(u5_mult_82_SUMB_25__40_) );
  XOR2_X2 u5_mult_82_U7505 ( .A(u5_mult_82_ab_25__40_), .B(
        u5_mult_82_CARRYB_24__40_), .Z(u5_mult_82_n2900) );
  NAND3_X4 u5_mult_82_U7504 ( .A1(u5_mult_82_n2897), .A2(u5_mult_82_n2898), 
        .A3(u5_mult_82_n2899), .ZN(u5_mult_82_CARRYB_30__22_) );
  NAND2_X1 u5_mult_82_U7503 ( .A1(u5_mult_82_ab_30__22_), .A2(
        u5_mult_82_CARRYB_29__22_), .ZN(u5_mult_82_n2897) );
  NAND2_X2 u5_mult_82_U7502 ( .A1(u5_mult_82_CARRYB_28__23_), .A2(
        u5_mult_82_n1522), .ZN(u5_mult_82_n2896) );
  NAND2_X2 u5_mult_82_U7501 ( .A1(u5_mult_82_ab_29__23_), .A2(u5_mult_82_n1522), .ZN(u5_mult_82_n2895) );
  NAND2_X1 u5_mult_82_U7500 ( .A1(u5_mult_82_ab_29__23_), .A2(
        u5_mult_82_CARRYB_28__23_), .ZN(u5_mult_82_n2894) );
  NAND2_X1 u5_mult_82_U7499 ( .A1(u5_mult_82_CARRYB_40__15_), .A2(
        u5_mult_82_SUMB_40__16_), .ZN(u5_mult_82_n2893) );
  NAND2_X1 u5_mult_82_U7498 ( .A1(u5_mult_82_ab_41__15_), .A2(
        u5_mult_82_SUMB_40__16_), .ZN(u5_mult_82_n2892) );
  NAND2_X1 u5_mult_82_U7497 ( .A1(u5_mult_82_ab_41__15_), .A2(
        u5_mult_82_CARRYB_40__15_), .ZN(u5_mult_82_n2891) );
  NAND2_X2 u5_mult_82_U7496 ( .A1(u5_mult_82_CARRYB_39__16_), .A2(
        u5_mult_82_SUMB_39__17_), .ZN(u5_mult_82_n2890) );
  NAND2_X2 u5_mult_82_U7495 ( .A1(u5_mult_82_ab_40__16_), .A2(
        u5_mult_82_SUMB_39__17_), .ZN(u5_mult_82_n2889) );
  NAND2_X2 u5_mult_82_U7494 ( .A1(u5_mult_82_ab_40__16_), .A2(
        u5_mult_82_CARRYB_39__16_), .ZN(u5_mult_82_n2888) );
  XOR2_X2 u5_mult_82_U7493 ( .A(u5_mult_82_n2887), .B(u5_mult_82_SUMB_39__17_), 
        .Z(u5_mult_82_SUMB_40__16_) );
  XOR2_X2 u5_mult_82_U7492 ( .A(u5_mult_82_ab_40__16_), .B(
        u5_mult_82_CARRYB_39__16_), .Z(u5_mult_82_n2887) );
  NAND3_X4 u5_mult_82_U7491 ( .A1(u5_mult_82_n2886), .A2(u5_mult_82_n2885), 
        .A3(u5_mult_82_n2884), .ZN(u5_mult_82_CARRYB_39__16_) );
  NAND2_X2 u5_mult_82_U7490 ( .A1(u5_mult_82_CARRYB_38__16_), .A2(
        u5_mult_82_SUMB_38__17_), .ZN(u5_mult_82_n2886) );
  NAND2_X2 u5_mult_82_U7489 ( .A1(u5_mult_82_ab_39__16_), .A2(
        u5_mult_82_SUMB_38__17_), .ZN(u5_mult_82_n2885) );
  NAND2_X2 u5_mult_82_U7488 ( .A1(u5_mult_82_CARRYB_37__17_), .A2(
        u5_mult_82_SUMB_37__18_), .ZN(u5_mult_82_n2883) );
  NAND2_X2 u5_mult_82_U7487 ( .A1(u5_mult_82_ab_38__17_), .A2(
        u5_mult_82_SUMB_37__18_), .ZN(u5_mult_82_n2882) );
  NAND2_X1 u5_mult_82_U7486 ( .A1(u5_mult_82_ab_38__17_), .A2(
        u5_mult_82_CARRYB_37__17_), .ZN(u5_mult_82_n2881) );
  XOR2_X2 u5_mult_82_U7485 ( .A(u5_mult_82_n2880), .B(u5_mult_82_SUMB_37__18_), 
        .Z(u5_mult_82_SUMB_38__17_) );
  XOR2_X2 u5_mult_82_U7484 ( .A(u5_mult_82_ab_38__17_), .B(
        u5_mult_82_CARRYB_37__17_), .Z(u5_mult_82_n2880) );
  NAND2_X2 u5_mult_82_U7483 ( .A1(u5_mult_82_CARRYB_40__9_), .A2(
        u5_mult_82_n1486), .ZN(u5_mult_82_n6067) );
  XNOR2_X2 u5_mult_82_U7482 ( .A(u5_mult_82_ab_24__25_), .B(
        u5_mult_82_CARRYB_23__25_), .ZN(u5_mult_82_n2879) );
  NAND2_X2 u5_mult_82_U7481 ( .A1(u5_mult_82_ab_29__21_), .A2(
        u5_mult_82_SUMB_28__22_), .ZN(u5_mult_82_n5436) );
  NOR2_X1 u5_mult_82_U7480 ( .A1(u5_mult_82_n6946), .A2(u5_mult_82_n6748), 
        .ZN(u5_mult_82_ab_48__4_) );
  NAND3_X4 u5_mult_82_U7479 ( .A1(u5_mult_82_n2876), .A2(u5_mult_82_n2877), 
        .A3(u5_mult_82_n2878), .ZN(u5_mult_82_CARRYB_41__8_) );
  NAND2_X1 u5_mult_82_U7478 ( .A1(u5_mult_82_ab_41__8_), .A2(
        u5_mult_82_SUMB_40__9_), .ZN(u5_mult_82_n2877) );
  NAND2_X1 u5_mult_82_U7477 ( .A1(u5_mult_82_ab_41__8_), .A2(
        u5_mult_82_CARRYB_40__8_), .ZN(u5_mult_82_n2876) );
  NAND3_X2 u5_mult_82_U7476 ( .A1(u5_mult_82_n2873), .A2(u5_mult_82_n2874), 
        .A3(u5_mult_82_n2875), .ZN(u5_mult_82_CARRYB_40__9_) );
  NAND2_X2 u5_mult_82_U7475 ( .A1(u5_mult_82_CARRYB_39__9_), .A2(
        u5_mult_82_SUMB_39__10_), .ZN(u5_mult_82_n2875) );
  NAND2_X2 u5_mult_82_U7474 ( .A1(u5_mult_82_ab_40__9_), .A2(
        u5_mult_82_SUMB_39__10_), .ZN(u5_mult_82_n2874) );
  NAND2_X1 u5_mult_82_U7473 ( .A1(u5_mult_82_ab_40__9_), .A2(
        u5_mult_82_CARRYB_39__9_), .ZN(u5_mult_82_n2873) );
  XOR2_X2 u5_mult_82_U7472 ( .A(u5_mult_82_n2872), .B(u5_mult_82_SUMB_39__10_), 
        .Z(u5_mult_82_SUMB_40__9_) );
  XOR2_X2 u5_mult_82_U7471 ( .A(u5_mult_82_ab_40__9_), .B(
        u5_mult_82_CARRYB_39__9_), .Z(u5_mult_82_n2872) );
  NAND3_X2 u5_mult_82_U7470 ( .A1(u5_mult_82_n2869), .A2(u5_mult_82_n2870), 
        .A3(u5_mult_82_n2871), .ZN(u5_mult_82_CARRYB_48__4_) );
  NAND2_X1 u5_mult_82_U7469 ( .A1(u5_mult_82_ab_48__4_), .A2(
        u5_mult_82_CARRYB_47__4_), .ZN(u5_mult_82_n2871) );
  NAND2_X2 u5_mult_82_U7468 ( .A1(u5_mult_82_ab_48__4_), .A2(
        u5_mult_82_SUMB_47__5_), .ZN(u5_mult_82_n2870) );
  NAND2_X1 u5_mult_82_U7467 ( .A1(u5_mult_82_CARRYB_47__4_), .A2(
        u5_mult_82_SUMB_47__5_), .ZN(u5_mult_82_n2869) );
  XOR2_X2 u5_mult_82_U7466 ( .A(u5_mult_82_SUMB_47__5_), .B(u5_mult_82_n2868), 
        .Z(u5_mult_82_SUMB_48__4_) );
  XOR2_X2 u5_mult_82_U7465 ( .A(u5_mult_82_CARRYB_47__4_), .B(
        u5_mult_82_ab_48__4_), .Z(u5_mult_82_n2868) );
  NAND2_X2 u5_mult_82_U7464 ( .A1(u5_mult_82_ab_13__41_), .A2(
        u5_mult_82_SUMB_12__42_), .ZN(u5_mult_82_n5174) );
  NAND2_X2 u5_mult_82_U7463 ( .A1(u5_mult_82_ab_21__36_), .A2(
        u5_mult_82_SUMB_20__37_), .ZN(u5_mult_82_n3873) );
  INV_X4 u5_mult_82_U7462 ( .A(u5_mult_82_net78853), .ZN(u5_mult_82_net84440)
         );
  NAND3_X4 u5_mult_82_U7461 ( .A1(u5_mult_82_n6339), .A2(u5_mult_82_n6340), 
        .A3(u5_mult_82_n6341), .ZN(u5_mult_82_CARRYB_22__32_) );
  INV_X2 u5_mult_82_U7460 ( .A(u5_mult_82_CARRYB_20__28_), .ZN(
        u5_mult_82_n2864) );
  INV_X2 u5_mult_82_U7459 ( .A(u5_mult_82_ab_21__28_), .ZN(u5_mult_82_n2863)
         );
  NAND2_X2 u5_mult_82_U7458 ( .A1(u5_mult_82_n2865), .A2(u5_mult_82_n2866), 
        .ZN(u5_mult_82_n3334) );
  NAND2_X1 u5_mult_82_U7457 ( .A1(u5_mult_82_n2863), .A2(
        u5_mult_82_CARRYB_20__28_), .ZN(u5_mult_82_n2866) );
  NAND2_X2 u5_mult_82_U7456 ( .A1(u5_mult_82_ab_21__28_), .A2(u5_mult_82_n2864), .ZN(u5_mult_82_n2865) );
  CLKBUF_X3 u5_mult_82_U7455 ( .A(u5_mult_82_CARRYB_32__7_), .Z(
        u5_mult_82_n3823) );
  NAND3_X2 u5_mult_82_U7454 ( .A1(u5_mult_82_n2860), .A2(u5_mult_82_n2861), 
        .A3(u5_mult_82_n2862), .ZN(u5_mult_82_CARRYB_22__13_) );
  NAND2_X1 u5_mult_82_U7453 ( .A1(u5_mult_82_CARRYB_21__13_), .A2(
        u5_mult_82_SUMB_21__14_), .ZN(u5_mult_82_n2862) );
  NAND2_X1 u5_mult_82_U7452 ( .A1(u5_mult_82_ab_22__13_), .A2(
        u5_mult_82_SUMB_21__14_), .ZN(u5_mult_82_n2861) );
  NAND2_X1 u5_mult_82_U7451 ( .A1(u5_mult_82_ab_22__13_), .A2(
        u5_mult_82_CARRYB_21__13_), .ZN(u5_mult_82_n2860) );
  NAND3_X2 u5_mult_82_U7450 ( .A1(u5_mult_82_n2857), .A2(u5_mult_82_n2858), 
        .A3(u5_mult_82_n2859), .ZN(u5_mult_82_CARRYB_21__14_) );
  NAND2_X2 u5_mult_82_U7449 ( .A1(u5_mult_82_CARRYB_20__14_), .A2(
        u5_mult_82_n1717), .ZN(u5_mult_82_n2859) );
  NAND2_X2 u5_mult_82_U7448 ( .A1(u5_mult_82_ab_21__14_), .A2(u5_mult_82_n1717), .ZN(u5_mult_82_n2858) );
  XOR2_X2 u5_mult_82_U7447 ( .A(u5_mult_82_n2856), .B(u5_mult_82_SUMB_21__14_), 
        .Z(u5_mult_82_SUMB_22__13_) );
  NAND3_X4 u5_mult_82_U7446 ( .A1(u5_mult_82_n2853), .A2(u5_mult_82_n2854), 
        .A3(u5_mult_82_n2855), .ZN(u5_mult_82_CARRYB_32__7_) );
  NAND2_X2 u5_mult_82_U7445 ( .A1(u5_mult_82_CARRYB_31__7_), .A2(
        u5_mult_82_SUMB_31__8_), .ZN(u5_mult_82_n2855) );
  NAND2_X2 u5_mult_82_U7444 ( .A1(u5_mult_82_ab_32__7_), .A2(
        u5_mult_82_SUMB_31__8_), .ZN(u5_mult_82_n2854) );
  NAND3_X2 u5_mult_82_U7443 ( .A1(u5_mult_82_n2850), .A2(u5_mult_82_n2851), 
        .A3(u5_mult_82_n2852), .ZN(u5_mult_82_CARRYB_31__8_) );
  NAND2_X2 u5_mult_82_U7442 ( .A1(u5_mult_82_CARRYB_30__8_), .A2(
        u5_mult_82_SUMB_30__9_), .ZN(u5_mult_82_n2852) );
  NAND2_X1 u5_mult_82_U7441 ( .A1(u5_mult_82_ab_31__8_), .A2(
        u5_mult_82_SUMB_30__9_), .ZN(u5_mult_82_n2851) );
  NAND2_X1 u5_mult_82_U7440 ( .A1(u5_mult_82_ab_31__8_), .A2(
        u5_mult_82_CARRYB_30__8_), .ZN(u5_mult_82_n2850) );
  XOR2_X2 u5_mult_82_U7439 ( .A(u5_mult_82_n2849), .B(u5_mult_82_SUMB_30__9_), 
        .Z(u5_mult_82_SUMB_31__8_) );
  XOR2_X2 u5_mult_82_U7438 ( .A(u5_mult_82_ab_31__8_), .B(
        u5_mult_82_CARRYB_30__8_), .Z(u5_mult_82_n2849) );
  XOR2_X2 u5_mult_82_U7437 ( .A(u5_mult_82_ab_22__29_), .B(
        u5_mult_82_CARRYB_21__29_), .Z(u5_mult_82_n4292) );
  NAND2_X2 u5_mult_82_U7436 ( .A1(u5_mult_82_ab_22__29_), .A2(
        u5_mult_82_SUMB_21__30_), .ZN(u5_mult_82_n4295) );
  NAND3_X4 u5_mult_82_U7435 ( .A1(u5_mult_82_n4286), .A2(u5_mult_82_n4287), 
        .A3(u5_mult_82_n4288), .ZN(u5_mult_82_CARRYB_44__16_) );
  NAND2_X1 u5_mult_82_U7434 ( .A1(u5_mult_82_ab_42__10_), .A2(
        u5_mult_82_CARRYB_41__10_), .ZN(u5_mult_82_n6164) );
  XNOR2_X2 u5_mult_82_U7433 ( .A(u5_mult_82_CARRYB_25__15_), .B(
        u5_mult_82_ab_26__15_), .ZN(u5_mult_82_n2848) );
  XNOR2_X2 u5_mult_82_U7432 ( .A(u5_mult_82_n2848), .B(u5_mult_82_n723), .ZN(
        u5_mult_82_SUMB_26__15_) );
  XNOR2_X2 u5_mult_82_U7431 ( .A(u5_mult_82_CARRYB_16__23_), .B(
        u5_mult_82_ab_17__23_), .ZN(u5_mult_82_n2847) );
  NAND2_X2 u5_mult_82_U7430 ( .A1(u5_mult_82_ab_39__7_), .A2(
        u5_mult_82_SUMB_38__8_), .ZN(u5_mult_82_n2988) );
  NAND2_X2 u5_mult_82_U7429 ( .A1(u5_mult_82_ab_16__37_), .A2(
        u5_mult_82_SUMB_15__38_), .ZN(u5_mult_82_n6306) );
  XNOR2_X2 u5_mult_82_U7428 ( .A(u5_mult_82_CARRYB_26__10_), .B(
        u5_mult_82_ab_27__10_), .ZN(u5_mult_82_n2846) );
  XNOR2_X2 u5_mult_82_U7427 ( .A(u5_mult_82_SUMB_26__11_), .B(u5_mult_82_n2846), .ZN(u5_mult_82_SUMB_27__10_) );
  NAND3_X2 u5_mult_82_U7426 ( .A1(u5_mult_82_n2843), .A2(u5_mult_82_n2844), 
        .A3(u5_mult_82_n2845), .ZN(u5_mult_82_CARRYB_21__15_) );
  NAND2_X1 u5_mult_82_U7425 ( .A1(u5_mult_82_CARRYB_20__15_), .A2(
        u5_mult_82_SUMB_20__16_), .ZN(u5_mult_82_n2845) );
  NAND2_X1 u5_mult_82_U7424 ( .A1(u5_mult_82_ab_21__15_), .A2(
        u5_mult_82_SUMB_20__16_), .ZN(u5_mult_82_n2844) );
  NAND2_X1 u5_mult_82_U7423 ( .A1(u5_mult_82_ab_21__15_), .A2(
        u5_mult_82_CARRYB_20__15_), .ZN(u5_mult_82_n2843) );
  NAND3_X4 u5_mult_82_U7422 ( .A1(u5_mult_82_n2840), .A2(u5_mult_82_n2841), 
        .A3(u5_mult_82_n2842), .ZN(u5_mult_82_CARRYB_20__16_) );
  NAND2_X2 u5_mult_82_U7421 ( .A1(u5_mult_82_ab_20__16_), .A2(
        u5_mult_82_SUMB_19__17_), .ZN(u5_mult_82_n2841) );
  NAND2_X2 u5_mult_82_U7420 ( .A1(u5_mult_82_CARRYB_19__16_), .A2(
        u5_mult_82_ab_20__16_), .ZN(u5_mult_82_n2840) );
  XOR2_X2 u5_mult_82_U7419 ( .A(u5_mult_82_n2839), .B(u5_mult_82_SUMB_19__17_), 
        .Z(u5_mult_82_SUMB_20__16_) );
  XOR2_X2 u5_mult_82_U7418 ( .A(u5_mult_82_ab_20__16_), .B(
        u5_mult_82_CARRYB_19__16_), .Z(u5_mult_82_n2839) );
  NAND3_X2 u5_mult_82_U7417 ( .A1(u5_mult_82_n2836), .A2(u5_mult_82_n2837), 
        .A3(u5_mult_82_n2838), .ZN(u5_mult_82_CARRYB_13__20_) );
  NAND2_X1 u5_mult_82_U7416 ( .A1(u5_mult_82_n1606), .A2(
        u5_mult_82_SUMB_12__21_), .ZN(u5_mult_82_n2838) );
  NAND2_X1 u5_mult_82_U7415 ( .A1(u5_mult_82_ab_13__20_), .A2(
        u5_mult_82_SUMB_12__21_), .ZN(u5_mult_82_n2837) );
  NAND2_X1 u5_mult_82_U7414 ( .A1(u5_mult_82_ab_13__20_), .A2(u5_mult_82_n1606), .ZN(u5_mult_82_n2836) );
  NAND3_X2 u5_mult_82_U7413 ( .A1(u5_mult_82_n2833), .A2(u5_mult_82_n2834), 
        .A3(u5_mult_82_n2835), .ZN(u5_mult_82_CARRYB_12__21_) );
  NAND2_X2 u5_mult_82_U7412 ( .A1(u5_mult_82_CARRYB_11__21_), .A2(
        u5_mult_82_SUMB_11__22_), .ZN(u5_mult_82_n2835) );
  NAND2_X2 u5_mult_82_U7411 ( .A1(u5_mult_82_ab_12__21_), .A2(
        u5_mult_82_SUMB_11__22_), .ZN(u5_mult_82_n2834) );
  NAND2_X1 u5_mult_82_U7410 ( .A1(u5_mult_82_ab_12__21_), .A2(
        u5_mult_82_CARRYB_11__21_), .ZN(u5_mult_82_n2833) );
  XOR2_X2 u5_mult_82_U7409 ( .A(u5_mult_82_n2832), .B(u5_mult_82_SUMB_12__21_), 
        .Z(u5_mult_82_SUMB_13__20_) );
  XOR2_X2 u5_mult_82_U7408 ( .A(u5_mult_82_ab_13__20_), .B(u5_mult_82_n1606), 
        .Z(u5_mult_82_n2832) );
  XOR2_X2 u5_mult_82_U7407 ( .A(u5_mult_82_n2831), .B(u5_mult_82_SUMB_11__22_), 
        .Z(u5_mult_82_SUMB_12__21_) );
  XOR2_X2 u5_mult_82_U7406 ( .A(u5_mult_82_ab_12__21_), .B(
        u5_mult_82_CARRYB_11__21_), .Z(u5_mult_82_n2831) );
  NAND3_X2 u5_mult_82_U7405 ( .A1(u5_mult_82_n2828), .A2(u5_mult_82_n2829), 
        .A3(u5_mult_82_n2830), .ZN(u5_mult_82_CARRYB_30__8_) );
  NAND2_X1 u5_mult_82_U7404 ( .A1(u5_mult_82_CARRYB_29__8_), .A2(
        u5_mult_82_SUMB_29__9_), .ZN(u5_mult_82_n2830) );
  NAND2_X1 u5_mult_82_U7403 ( .A1(u5_mult_82_ab_30__8_), .A2(
        u5_mult_82_SUMB_29__9_), .ZN(u5_mult_82_n2829) );
  NAND2_X1 u5_mult_82_U7402 ( .A1(u5_mult_82_ab_30__8_), .A2(
        u5_mult_82_CARRYB_29__8_), .ZN(u5_mult_82_n2828) );
  NAND3_X2 u5_mult_82_U7401 ( .A1(u5_mult_82_n2825), .A2(u5_mult_82_n2826), 
        .A3(u5_mult_82_n2827), .ZN(u5_mult_82_CARRYB_29__9_) );
  NAND2_X1 u5_mult_82_U7400 ( .A1(u5_mult_82_ab_29__9_), .A2(
        u5_mult_82_CARRYB_28__9_), .ZN(u5_mult_82_n2825) );
  XOR2_X2 u5_mult_82_U7399 ( .A(u5_mult_82_n399), .B(u5_mult_82_n2824), .Z(
        u5_mult_82_SUMB_29__9_) );
  XOR2_X2 u5_mult_82_U7398 ( .A(u5_mult_82_ab_29__9_), .B(
        u5_mult_82_CARRYB_28__9_), .Z(u5_mult_82_n2824) );
  NAND3_X2 u5_mult_82_U7397 ( .A1(u5_mult_82_n2821), .A2(u5_mult_82_n2822), 
        .A3(u5_mult_82_n2823), .ZN(u5_mult_82_CARRYB_25__11_) );
  NAND2_X1 u5_mult_82_U7396 ( .A1(u5_mult_82_ab_25__11_), .A2(
        u5_mult_82_CARRYB_24__11_), .ZN(u5_mult_82_n2821) );
  NAND2_X2 u5_mult_82_U7395 ( .A1(u5_mult_82_n397), .A2(
        u5_mult_82_CARRYB_23__12_), .ZN(u5_mult_82_n2820) );
  NAND2_X2 u5_mult_82_U7394 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_ab_24__12_), 
        .ZN(u5_mult_82_n2819) );
  NAND2_X1 u5_mult_82_U7393 ( .A1(u5_mult_82_ab_24__12_), .A2(
        u5_mult_82_CARRYB_23__12_), .ZN(u5_mult_82_n2818) );
  XOR2_X2 u5_mult_82_U7392 ( .A(u5_mult_82_n2817), .B(u5_mult_82_SUMB_24__12_), 
        .Z(u5_mult_82_SUMB_25__11_) );
  XOR2_X2 u5_mult_82_U7391 ( .A(u5_mult_82_ab_25__11_), .B(
        u5_mult_82_CARRYB_24__11_), .Z(u5_mult_82_n2817) );
  XOR2_X1 u5_mult_82_U7390 ( .A(u5_mult_82_ab_24__12_), .B(
        u5_mult_82_CARRYB_23__12_), .Z(u5_mult_82_n2816) );
  NAND3_X2 u5_mult_82_U7389 ( .A1(u5_mult_82_n2813), .A2(u5_mult_82_n2814), 
        .A3(u5_mult_82_n2815), .ZN(u5_mult_82_CARRYB_28__31_) );
  NAND2_X2 u5_mult_82_U7388 ( .A1(u5_mult_82_ab_28__31_), .A2(
        u5_mult_82_SUMB_27__32_), .ZN(u5_mult_82_n2814) );
  NAND3_X2 u5_mult_82_U7387 ( .A1(u5_mult_82_n2810), .A2(u5_mult_82_n2811), 
        .A3(u5_mult_82_n2812), .ZN(u5_mult_82_CARRYB_27__32_) );
  NAND2_X1 u5_mult_82_U7386 ( .A1(u5_mult_82_CARRYB_26__32_), .A2(
        u5_mult_82_SUMB_26__33_), .ZN(u5_mult_82_n2812) );
  NAND2_X1 u5_mult_82_U7385 ( .A1(u5_mult_82_ab_27__32_), .A2(
        u5_mult_82_SUMB_26__33_), .ZN(u5_mult_82_n2811) );
  NAND2_X1 u5_mult_82_U7384 ( .A1(u5_mult_82_ab_27__32_), .A2(
        u5_mult_82_CARRYB_26__32_), .ZN(u5_mult_82_n2810) );
  NAND3_X2 u5_mult_82_U7383 ( .A1(u5_mult_82_n2807), .A2(u5_mult_82_n2808), 
        .A3(u5_mult_82_n2809), .ZN(u5_mult_82_CARRYB_36__26_) );
  NAND2_X1 u5_mult_82_U7382 ( .A1(u5_mult_82_CARRYB_35__26_), .A2(
        u5_mult_82_SUMB_35__27_), .ZN(u5_mult_82_n2809) );
  NAND2_X1 u5_mult_82_U7381 ( .A1(u5_mult_82_ab_36__26_), .A2(
        u5_mult_82_SUMB_35__27_), .ZN(u5_mult_82_n2808) );
  NAND2_X1 u5_mult_82_U7380 ( .A1(u5_mult_82_ab_36__26_), .A2(
        u5_mult_82_CARRYB_35__26_), .ZN(u5_mult_82_n2807) );
  NAND3_X2 u5_mult_82_U7379 ( .A1(u5_mult_82_n2804), .A2(u5_mult_82_n2805), 
        .A3(u5_mult_82_n2806), .ZN(u5_mult_82_CARRYB_35__27_) );
  NAND2_X2 u5_mult_82_U7378 ( .A1(u5_mult_82_ab_35__27_), .A2(
        u5_mult_82_SUMB_34__28_), .ZN(u5_mult_82_n2805) );
  NAND2_X1 u5_mult_82_U7377 ( .A1(u5_mult_82_ab_35__27_), .A2(
        u5_mult_82_CARRYB_34__27_), .ZN(u5_mult_82_n2804) );
  XOR2_X2 u5_mult_82_U7376 ( .A(u5_mult_82_n2803), .B(u5_mult_82_n1479), .Z(
        u5_mult_82_SUMB_35__27_) );
  XOR2_X2 u5_mult_82_U7375 ( .A(u5_mult_82_CARRYB_34__27_), .B(
        u5_mult_82_ab_35__27_), .Z(u5_mult_82_n2803) );
  NAND2_X1 u5_mult_82_U7374 ( .A1(u5_mult_82_ab_20__43_), .A2(
        u5_mult_82_CARRYB_19__43_), .ZN(u5_mult_82_n4602) );
  XOR2_X2 u5_mult_82_U7373 ( .A(u5_mult_82_n3322), .B(u5_mult_82_SUMB_18__12_), 
        .Z(u5_mult_82_SUMB_19__11_) );
  NAND3_X4 u5_mult_82_U7372 ( .A1(u5_mult_82_n2799), .A2(u5_mult_82_n2800), 
        .A3(u5_mult_82_n2801), .ZN(u5_mult_82_CARRYB_20__19_) );
  NAND2_X2 u5_mult_82_U7371 ( .A1(u5_mult_82_CARRYB_19__19_), .A2(
        u5_mult_82_SUMB_19__20_), .ZN(u5_mult_82_n2801) );
  NAND2_X2 u5_mult_82_U7370 ( .A1(u5_mult_82_ab_20__19_), .A2(
        u5_mult_82_SUMB_19__20_), .ZN(u5_mult_82_n2800) );
  NAND2_X1 u5_mult_82_U7369 ( .A1(u5_mult_82_ab_20__19_), .A2(
        u5_mult_82_CARRYB_19__19_), .ZN(u5_mult_82_n2799) );
  NAND2_X2 u5_mult_82_U7368 ( .A1(u5_mult_82_CARRYB_18__20_), .A2(
        u5_mult_82_n692), .ZN(u5_mult_82_n2798) );
  NAND2_X2 u5_mult_82_U7367 ( .A1(u5_mult_82_ab_19__20_), .A2(u5_mult_82_n692), 
        .ZN(u5_mult_82_n2797) );
  NAND2_X1 u5_mult_82_U7366 ( .A1(u5_mult_82_ab_19__20_), .A2(
        u5_mult_82_CARRYB_18__20_), .ZN(u5_mult_82_n2796) );
  XOR2_X2 u5_mult_82_U7365 ( .A(u5_mult_82_n2795), .B(u5_mult_82_SUMB_19__20_), 
        .Z(u5_mult_82_SUMB_20__19_) );
  XOR2_X1 u5_mult_82_U7364 ( .A(u5_mult_82_ab_20__19_), .B(
        u5_mult_82_CARRYB_19__19_), .Z(u5_mult_82_n2795) );
  XOR2_X2 u5_mult_82_U7363 ( .A(u5_mult_82_n2794), .B(u5_mult_82_n692), .Z(
        u5_mult_82_SUMB_19__20_) );
  NAND3_X2 u5_mult_82_U7362 ( .A1(u5_mult_82_n2791), .A2(u5_mult_82_n2792), 
        .A3(u5_mult_82_n2793), .ZN(u5_mult_82_CARRYB_29__13_) );
  NAND2_X1 u5_mult_82_U7361 ( .A1(u5_mult_82_ab_29__13_), .A2(
        u5_mult_82_CARRYB_28__13_), .ZN(u5_mult_82_n2791) );
  NAND2_X2 u5_mult_82_U7360 ( .A1(u5_mult_82_n1657), .A2(
        u5_mult_82_SUMB_27__15_), .ZN(u5_mult_82_n2790) );
  NAND2_X2 u5_mult_82_U7359 ( .A1(u5_mult_82_ab_28__14_), .A2(
        u5_mult_82_SUMB_27__15_), .ZN(u5_mult_82_n2789) );
  NAND2_X2 u5_mult_82_U7358 ( .A1(u5_mult_82_ab_28__14_), .A2(u5_mult_82_n1657), .ZN(u5_mult_82_n2788) );
  XOR2_X2 u5_mult_82_U7357 ( .A(u5_mult_82_n2787), .B(u5_mult_82_SUMB_27__15_), 
        .Z(u5_mult_82_SUMB_28__14_) );
  NAND2_X2 u5_mult_82_U7356 ( .A1(u5_mult_82_ab_27__15_), .A2(
        u5_mult_82_SUMB_26__16_), .ZN(u5_mult_82_n2786) );
  NAND2_X1 u5_mult_82_U7355 ( .A1(u5_mult_82_CARRYB_26__15_), .A2(
        u5_mult_82_ab_27__15_), .ZN(u5_mult_82_n2784) );
  NAND2_X1 u5_mult_82_U7354 ( .A1(u5_mult_82_ab_26__16_), .A2(
        u5_mult_82_CARRYB_25__16_), .ZN(u5_mult_82_n2781) );
  NAND2_X1 u5_mult_82_U7353 ( .A1(u5_mult_82_SUMB_22__9_), .A2(
        u5_mult_82_CARRYB_22__8_), .ZN(u5_mult_82_n2780) );
  NAND2_X2 u5_mult_82_U7352 ( .A1(u5_mult_82_ab_23__8_), .A2(
        u5_mult_82_CARRYB_22__8_), .ZN(u5_mult_82_n2779) );
  NAND2_X1 u5_mult_82_U7351 ( .A1(u5_mult_82_ab_23__8_), .A2(
        u5_mult_82_SUMB_22__9_), .ZN(u5_mult_82_n2778) );
  NAND3_X2 u5_mult_82_U7350 ( .A1(u5_mult_82_n2775), .A2(u5_mult_82_n2776), 
        .A3(u5_mult_82_n2777), .ZN(u5_mult_82_CARRYB_22__8_) );
  NAND2_X1 u5_mult_82_U7349 ( .A1(u5_mult_82_CARRYB_21__8_), .A2(
        u5_mult_82_SUMB_21__9_), .ZN(u5_mult_82_n2777) );
  NAND2_X2 u5_mult_82_U7348 ( .A1(u5_mult_82_ab_22__8_), .A2(
        u5_mult_82_SUMB_21__9_), .ZN(u5_mult_82_n2776) );
  NAND2_X1 u5_mult_82_U7347 ( .A1(u5_mult_82_ab_22__8_), .A2(
        u5_mult_82_CARRYB_21__8_), .ZN(u5_mult_82_n2775) );
  XOR2_X2 u5_mult_82_U7346 ( .A(u5_mult_82_n2774), .B(u5_mult_82_SUMB_21__9_), 
        .Z(u5_mult_82_SUMB_22__8_) );
  XOR2_X2 u5_mult_82_U7345 ( .A(u5_mult_82_ab_22__8_), .B(
        u5_mult_82_CARRYB_21__8_), .Z(u5_mult_82_n2774) );
  NAND3_X2 u5_mult_82_U7344 ( .A1(u5_mult_82_n2771), .A2(u5_mult_82_n2772), 
        .A3(u5_mult_82_n2773), .ZN(u5_mult_82_CARRYB_11__16_) );
  NAND2_X1 u5_mult_82_U7343 ( .A1(u5_mult_82_CARRYB_10__16_), .A2(
        u5_mult_82_SUMB_10__17_), .ZN(u5_mult_82_n2773) );
  NAND2_X1 u5_mult_82_U7342 ( .A1(u5_mult_82_ab_11__16_), .A2(
        u5_mult_82_SUMB_10__17_), .ZN(u5_mult_82_n2772) );
  NAND2_X1 u5_mult_82_U7341 ( .A1(u5_mult_82_ab_11__16_), .A2(
        u5_mult_82_CARRYB_10__16_), .ZN(u5_mult_82_n2771) );
  NAND3_X4 u5_mult_82_U7340 ( .A1(u5_mult_82_n2768), .A2(u5_mult_82_n2769), 
        .A3(u5_mult_82_n2770), .ZN(u5_mult_82_CARRYB_10__17_) );
  NAND2_X2 u5_mult_82_U7339 ( .A1(u5_mult_82_CARRYB_9__17_), .A2(
        u5_mult_82_SUMB_9__18_), .ZN(u5_mult_82_n2770) );
  NAND2_X2 u5_mult_82_U7338 ( .A1(u5_mult_82_ab_10__17_), .A2(
        u5_mult_82_SUMB_9__18_), .ZN(u5_mult_82_n2769) );
  NAND2_X1 u5_mult_82_U7337 ( .A1(u5_mult_82_ab_10__17_), .A2(
        u5_mult_82_CARRYB_9__17_), .ZN(u5_mult_82_n2768) );
  XOR2_X2 u5_mult_82_U7336 ( .A(u5_mult_82_n2767), .B(u5_mult_82_SUMB_9__18_), 
        .Z(u5_mult_82_SUMB_10__17_) );
  XOR2_X2 u5_mult_82_U7335 ( .A(u5_mult_82_ab_10__17_), .B(
        u5_mult_82_CARRYB_9__17_), .Z(u5_mult_82_n2767) );
  NAND3_X2 u5_mult_82_U7334 ( .A1(u5_mult_82_n2764), .A2(u5_mult_82_n2765), 
        .A3(u5_mult_82_n2766), .ZN(u5_mult_82_CARRYB_9__18_) );
  NAND2_X1 u5_mult_82_U7333 ( .A1(u5_mult_82_CARRYB_8__18_), .A2(
        u5_mult_82_SUMB_8__19_), .ZN(u5_mult_82_n2766) );
  NAND2_X1 u5_mult_82_U7332 ( .A1(u5_mult_82_ab_9__18_), .A2(
        u5_mult_82_SUMB_8__19_), .ZN(u5_mult_82_n2765) );
  NAND2_X1 u5_mult_82_U7331 ( .A1(u5_mult_82_ab_9__18_), .A2(
        u5_mult_82_CARRYB_8__18_), .ZN(u5_mult_82_n2764) );
  NAND3_X2 u5_mult_82_U7330 ( .A1(u5_mult_82_n2761), .A2(u5_mult_82_n2762), 
        .A3(u5_mult_82_n2763), .ZN(u5_mult_82_CARRYB_8__19_) );
  NAND2_X1 u5_mult_82_U7329 ( .A1(u5_mult_82_CARRYB_7__19_), .A2(
        u5_mult_82_SUMB_7__20_), .ZN(u5_mult_82_n2763) );
  NAND2_X1 u5_mult_82_U7328 ( .A1(u5_mult_82_ab_8__19_), .A2(
        u5_mult_82_SUMB_7__20_), .ZN(u5_mult_82_n2762) );
  XOR2_X2 u5_mult_82_U7327 ( .A(u5_mult_82_n2760), .B(u5_mult_82_SUMB_8__19_), 
        .Z(u5_mult_82_SUMB_9__18_) );
  XOR2_X2 u5_mult_82_U7326 ( .A(u5_mult_82_ab_9__18_), .B(
        u5_mult_82_CARRYB_8__18_), .Z(u5_mult_82_n2760) );
  XOR2_X2 u5_mult_82_U7325 ( .A(u5_mult_82_n2759), .B(u5_mult_82_SUMB_7__20_), 
        .Z(u5_mult_82_SUMB_8__19_) );
  XOR2_X2 u5_mult_82_U7324 ( .A(u5_mult_82_ab_8__19_), .B(
        u5_mult_82_CARRYB_7__19_), .Z(u5_mult_82_n2759) );
  XNOR2_X2 u5_mult_82_U7323 ( .A(u5_mult_82_CARRYB_47__35_), .B(
        u5_mult_82_ab_48__35_), .ZN(u5_mult_82_n2758) );
  XNOR2_X2 u5_mult_82_U7322 ( .A(u5_mult_82_n1503), .B(u5_mult_82_n2758), .ZN(
        u5_mult_82_SUMB_48__35_) );
  XNOR2_X2 u5_mult_82_U7321 ( .A(u5_mult_82_n3056), .B(u5_mult_82_SUMB_33__8_), 
        .ZN(u5_mult_82_SUMB_34__7_) );
  INV_X4 u5_mult_82_U7320 ( .A(u5_mult_82_CARRYB_30__19_), .ZN(
        u5_mult_82_n2755) );
  INV_X8 u5_mult_82_U7319 ( .A(u5_mult_82_ab_31__19_), .ZN(u5_mult_82_n2754)
         );
  NAND2_X4 u5_mult_82_U7318 ( .A1(u5_mult_82_n2756), .A2(u5_mult_82_n2757), 
        .ZN(u5_mult_82_n3582) );
  NAND2_X4 u5_mult_82_U7317 ( .A1(u5_mult_82_n2754), .A2(u5_mult_82_n2755), 
        .ZN(u5_mult_82_n2757) );
  XNOR2_X2 u5_mult_82_U7316 ( .A(u5_mult_82_SUMB_28__22_), .B(u5_mult_82_n2753), .ZN(u5_mult_82_SUMB_29__21_) );
  XNOR2_X2 u5_mult_82_U7315 ( .A(u5_mult_82_n2752), .B(u5_mult_82_SUMB_10__51_), .ZN(u5_mult_82_SUMB_11__50_) );
  XNOR2_X2 u5_mult_82_U7314 ( .A(u5_mult_82_n2751), .B(u5_mult_82_SUMB_26__19_), .ZN(u5_mult_82_SUMB_27__18_) );
  XNOR2_X2 u5_mult_82_U7313 ( .A(u5_mult_82_ab_32__17_), .B(
        u5_mult_82_CARRYB_31__17_), .ZN(u5_mult_82_net84580) );
  NAND3_X2 u5_mult_82_U7312 ( .A1(u5_mult_82_net80614), .A2(u5_mult_82_n5155), 
        .A3(u5_mult_82_net80616), .ZN(u5_mult_82_CARRYB_3__36_) );
  XNOR2_X2 u5_mult_82_U7311 ( .A(u5_mult_82_n1428), .B(u5_mult_82_n2749), .ZN(
        u5_mult_82_SUMB_26__29_) );
  NAND2_X2 u5_mult_82_U7310 ( .A1(u5_mult_82_ab_17__16_), .A2(
        u5_mult_82_SUMB_16__17_), .ZN(u5_mult_82_n4027) );
  NAND2_X1 u5_mult_82_U7309 ( .A1(u5_mult_82_ab_18__16_), .A2(
        u5_mult_82_CARRYB_17__16_), .ZN(u5_mult_82_n4112) );
  NAND2_X2 u5_mult_82_U7308 ( .A1(u5_mult_82_ab_46__7_), .A2(
        u5_mult_82_SUMB_45__8_), .ZN(u5_mult_82_n4377) );
  NAND2_X2 u5_mult_82_U7307 ( .A1(u5_mult_82_ab_43__9_), .A2(
        u5_mult_82_CARRYB_42__9_), .ZN(u5_mult_82_n5488) );
  INV_X4 u5_mult_82_U7306 ( .A(u5_mult_82_n4218), .ZN(u5_mult_82_n2745) );
  INV_X1 u5_mult_82_U7305 ( .A(u5_mult_82_CARRYB_44__8_), .ZN(u5_mult_82_n2744) );
  INV_X1 u5_mult_82_U7304 ( .A(u5_mult_82_SUMB_43__10_), .ZN(
        u5_mult_82_net84601) );
  INV_X4 u5_mult_82_U7303 ( .A(u5_mult_82_n5142), .ZN(u5_mult_82_n2741) );
  NAND2_X2 u5_mult_82_U7302 ( .A1(u5_mult_82_n2741), .A2(u5_mult_82_net84601), 
        .ZN(u5_mult_82_n2743) );
  NAND3_X2 u5_mult_82_U7301 ( .A1(u5_mult_82_n5488), .A2(u5_mult_82_n5489), 
        .A3(u5_mult_82_n5490), .ZN(u5_mult_82_net84599) );
  XNOR2_X2 u5_mult_82_U7300 ( .A(u5_mult_82_ab_13__32_), .B(
        u5_mult_82_CARRYB_12__32_), .ZN(u5_mult_82_n2740) );
  XNOR2_X2 u5_mult_82_U7299 ( .A(u5_mult_82_ab_18__47_), .B(
        u5_mult_82_CARRYB_17__47_), .ZN(u5_mult_82_n2739) );
  XNOR2_X2 u5_mult_82_U7298 ( .A(u5_mult_82_n2739), .B(u5_mult_82_SUMB_17__48_), .ZN(u5_mult_82_SUMB_18__47_) );
  INV_X1 u5_mult_82_U7297 ( .A(u5_mult_82_SUMB_7__37_), .ZN(u5_mult_82_n2736)
         );
  INV_X4 u5_mult_82_U7296 ( .A(u5_mult_82_n3277), .ZN(u5_mult_82_n2735) );
  NAND2_X2 u5_mult_82_U7295 ( .A1(u5_mult_82_n2737), .A2(u5_mult_82_n2738), 
        .ZN(u5_mult_82_SUMB_8__36_) );
  NAND2_X2 u5_mult_82_U7294 ( .A1(u5_mult_82_n2735), .A2(u5_mult_82_n2736), 
        .ZN(u5_mult_82_n2738) );
  XNOR2_X2 u5_mult_82_U7293 ( .A(u5_mult_82_ab_29__36_), .B(
        u5_mult_82_CARRYB_28__36_), .ZN(u5_mult_82_n2734) );
  XNOR2_X2 u5_mult_82_U7292 ( .A(u5_mult_82_n2734), .B(u5_mult_82_SUMB_28__37_), .ZN(u5_mult_82_SUMB_29__36_) );
  XNOR2_X2 u5_mult_82_U7291 ( .A(u5_mult_82_ab_6__37_), .B(
        u5_mult_82_CARRYB_5__37_), .ZN(u5_mult_82_n2733) );
  NAND2_X2 u5_mult_82_U7290 ( .A1(u5_mult_82_net78853), .A2(
        u5_mult_82_net84441), .ZN(u5_mult_82_n2867) );
  NAND2_X4 u5_mult_82_U7289 ( .A1(u5_mult_82_n2867), .A2(u5_mult_82_net84443), 
        .ZN(u5_mult_82_SUMB_43__10_) );
  NAND2_X2 u5_mult_82_U7288 ( .A1(u5_mult_82_ab_15__45_), .A2(
        u5_mult_82_CARRYB_14__45_), .ZN(u5_mult_82_n6125) );
  NAND2_X1 u5_mult_82_U7287 ( .A1(u5_mult_82_CARRYB_14__45_), .A2(
        u5_mult_82_n1639), .ZN(u5_mult_82_n6127) );
  NOR2_X2 u5_mult_82_U7286 ( .A1(u5_mult_82_n6799), .A2(u5_mult_82_n6580), 
        .ZN(u5_mult_82_ab_14__45_) );
  NAND3_X2 u5_mult_82_U7285 ( .A1(u5_mult_82_n2731), .A2(u5_mult_82_n2730), 
        .A3(u5_mult_82_n2732), .ZN(u5_mult_82_CARRYB_17__42_) );
  NAND2_X1 u5_mult_82_U7284 ( .A1(u5_mult_82_ab_17__42_), .A2(
        u5_mult_82_SUMB_16__43_), .ZN(u5_mult_82_n2731) );
  NAND2_X1 u5_mult_82_U7283 ( .A1(u5_mult_82_ab_17__42_), .A2(
        u5_mult_82_CARRYB_16__42_), .ZN(u5_mult_82_n2730) );
  NAND2_X2 u5_mult_82_U7282 ( .A1(u5_mult_82_CARRYB_15__43_), .A2(
        u5_mult_82_SUMB_15__44_), .ZN(u5_mult_82_n2729) );
  NAND2_X2 u5_mult_82_U7281 ( .A1(u5_mult_82_ab_16__43_), .A2(
        u5_mult_82_SUMB_15__44_), .ZN(u5_mult_82_n2728) );
  NAND3_X4 u5_mult_82_U7280 ( .A1(u5_mult_82_n2724), .A2(u5_mult_82_n2725), 
        .A3(u5_mult_82_n2726), .ZN(u5_mult_82_CARRYB_14__45_) );
  NAND2_X1 u5_mult_82_U7279 ( .A1(u5_mult_82_ab_14__45_), .A2(
        u5_mult_82_CARRYB_13__45_), .ZN(u5_mult_82_n2726) );
  NAND2_X2 u5_mult_82_U7278 ( .A1(u5_mult_82_ab_14__45_), .A2(
        u5_mult_82_SUMB_13__46_), .ZN(u5_mult_82_n2725) );
  XOR2_X2 u5_mult_82_U7277 ( .A(u5_mult_82_SUMB_13__46_), .B(u5_mult_82_n2723), 
        .Z(u5_mult_82_SUMB_14__45_) );
  XOR2_X2 u5_mult_82_U7276 ( .A(u5_mult_82_CARRYB_13__45_), .B(
        u5_mult_82_ab_14__45_), .Z(u5_mult_82_n2723) );
  NAND3_X4 u5_mult_82_U7275 ( .A1(u5_mult_82_n2720), .A2(u5_mult_82_n2721), 
        .A3(u5_mult_82_n2722), .ZN(u5_mult_82_CARRYB_35__31_) );
  NAND2_X2 u5_mult_82_U7274 ( .A1(u5_mult_82_CARRYB_34__31_), .A2(
        u5_mult_82_SUMB_34__32_), .ZN(u5_mult_82_n2722) );
  NAND2_X2 u5_mult_82_U7273 ( .A1(u5_mult_82_ab_35__31_), .A2(
        u5_mult_82_SUMB_34__32_), .ZN(u5_mult_82_n2721) );
  NAND2_X1 u5_mult_82_U7272 ( .A1(u5_mult_82_ab_35__31_), .A2(
        u5_mult_82_CARRYB_34__31_), .ZN(u5_mult_82_n2720) );
  NAND3_X4 u5_mult_82_U7271 ( .A1(u5_mult_82_n2719), .A2(u5_mult_82_n2718), 
        .A3(u5_mult_82_n2717), .ZN(u5_mult_82_CARRYB_34__32_) );
  NAND2_X1 u5_mult_82_U7270 ( .A1(u5_mult_82_ab_34__32_), .A2(
        u5_mult_82_CARRYB_33__32_), .ZN(u5_mult_82_n2717) );
  XOR2_X2 u5_mult_82_U7269 ( .A(u5_mult_82_n4292), .B(u5_mult_82_SUMB_21__30_), 
        .Z(u5_mult_82_SUMB_22__29_) );
  NAND2_X2 u5_mult_82_U7268 ( .A1(u5_mult_82_SUMB_16__27_), .A2(
        u5_mult_82_CARRYB_16__26_), .ZN(u5_mult_82_n4776) );
  NAND3_X4 u5_mult_82_U7267 ( .A1(u5_mult_82_n4026), .A2(u5_mult_82_n4027), 
        .A3(u5_mult_82_n4028), .ZN(u5_mult_82_CARRYB_17__16_) );
  INV_X1 u5_mult_82_U7266 ( .A(u5_mult_82_net64911), .ZN(u5_mult_82_net64899)
         );
  NAND2_X1 u5_mult_82_U7265 ( .A1(u5_mult_82_ab_0__30_), .A2(
        u5_mult_82_ab_1__29_), .ZN(u5_mult_82_n6482) );
  NAND2_X2 u5_mult_82_U7264 ( .A1(u5_mult_82_CARRYB_20__34_), .A2(
        u5_mult_82_n1725), .ZN(u5_mult_82_n5542) );
  XNOR2_X2 u5_mult_82_U7263 ( .A(u5_mult_82_ab_48__36_), .B(
        u5_mult_82_CARRYB_47__36_), .ZN(u5_mult_82_n2714) );
  INV_X16 u5_mult_82_U7262 ( .A(u5_mult_82_n7014), .ZN(u5_mult_82_n6866) );
  XNOR2_X2 u5_mult_82_U7261 ( .A(u5_mult_82_CARRYB_34__28_), .B(
        u5_mult_82_ab_35__28_), .ZN(u5_mult_82_n2713) );
  XNOR2_X2 u5_mult_82_U7260 ( .A(u5_mult_82_n2713), .B(u5_mult_82_SUMB_34__29_), .ZN(u5_mult_82_SUMB_35__28_) );
  XNOR2_X2 u5_mult_82_U7259 ( .A(u5_mult_82_SUMB_20__47_), .B(u5_mult_82_n2711), .ZN(u5_mult_82_n2927) );
  NAND2_X2 u5_mult_82_U7258 ( .A1(u5_mult_82_ab_11__51_), .A2(
        u5_mult_82_CARRYB_10__51_), .ZN(u5_mult_82_n4649) );
  NAND2_X4 u5_mult_82_U7257 ( .A1(u5_mult_82_ab_1__34_), .A2(
        u5_mult_82_ab_0__35_), .ZN(u5_mult_82_n6489) );
  XNOR2_X2 u5_mult_82_U7256 ( .A(u5_mult_82_n5), .B(u5_mult_82_ab_47__36_), 
        .ZN(u5_mult_82_n2802) );
  NAND2_X2 u5_mult_82_U7255 ( .A1(u5_mult_82_CARRYB_16__16_), .A2(
        u5_mult_82_SUMB_16__17_), .ZN(u5_mult_82_n4026) );
  XNOR2_X2 u5_mult_82_U7254 ( .A(u5_mult_82_ab_48__33_), .B(
        u5_mult_82_CARRYB_47__33_), .ZN(u5_mult_82_n2712) );
  NAND3_X2 u5_mult_82_U7253 ( .A1(u5_mult_82_net80542), .A2(
        u5_mult_82_net80543), .A3(u5_mult_82_n5218), .ZN(
        u5_mult_82_CARRYB_21__24_) );
  INV_X2 u5_mult_82_U7252 ( .A(u5_mult_82_SUMB_47__33_), .ZN(u5_mult_82_n2709)
         );
  NAND2_X2 u5_mult_82_U7251 ( .A1(u5_mult_82_ab_32__39_), .A2(
        u5_mult_82_SUMB_31__40_), .ZN(u5_mult_82_n5079) );
  XNOR2_X2 u5_mult_82_U7250 ( .A(u5_mult_82_CARRYB_16__20_), .B(
        u5_mult_82_ab_17__20_), .ZN(u5_mult_82_n2708) );
  XNOR2_X2 u5_mult_82_U7249 ( .A(u5_mult_82_n1642), .B(u5_mult_82_n2708), .ZN(
        u5_mult_82_SUMB_17__20_) );
  XNOR2_X2 u5_mult_82_U7248 ( .A(u5_mult_82_ab_17__14_), .B(
        u5_mult_82_CARRYB_16__14_), .ZN(u5_mult_82_n2707) );
  XNOR2_X2 u5_mult_82_U7247 ( .A(u5_mult_82_n2707), .B(u5_mult_82_SUMB_16__15_), .ZN(u5_mult_82_SUMB_17__14_) );
  INV_X8 u5_mult_82_U7246 ( .A(n4752), .ZN(u5_mult_82_n7018) );
  NOR2_X1 u5_mult_82_U7245 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6753), 
        .ZN(u5_mult_82_ab_49__36_) );
  NOR2_X1 u5_mult_82_U7244 ( .A1(u5_mult_82_net64935), .A2(u5_mult_82_n6747), 
        .ZN(u5_mult_82_ab_48__37_) );
  NAND3_X2 u5_mult_82_U7243 ( .A1(u5_mult_82_n2705), .A2(u5_mult_82_n2704), 
        .A3(u5_mult_82_n2706), .ZN(u5_mult_82_CARRYB_49__36_) );
  NAND2_X1 u5_mult_82_U7242 ( .A1(u5_mult_82_ab_49__36_), .A2(
        u5_mult_82_CARRYB_48__36_), .ZN(u5_mult_82_n2706) );
  NAND2_X2 u5_mult_82_U7241 ( .A1(u5_mult_82_ab_49__36_), .A2(
        u5_mult_82_SUMB_48__37_), .ZN(u5_mult_82_n2705) );
  XOR2_X2 u5_mult_82_U7240 ( .A(u5_mult_82_SUMB_48__37_), .B(u5_mult_82_n2703), 
        .Z(u5_mult_82_SUMB_49__36_) );
  XOR2_X2 u5_mult_82_U7239 ( .A(u5_mult_82_CARRYB_48__36_), .B(
        u5_mult_82_ab_49__36_), .Z(u5_mult_82_n2703) );
  NAND3_X2 u5_mult_82_U7238 ( .A1(u5_mult_82_n2700), .A2(u5_mult_82_n2701), 
        .A3(u5_mult_82_n2702), .ZN(u5_mult_82_CARRYB_48__37_) );
  NAND2_X1 u5_mult_82_U7237 ( .A1(u5_mult_82_ab_48__37_), .A2(
        u5_mult_82_CARRYB_47__37_), .ZN(u5_mult_82_n2702) );
  NAND2_X1 u5_mult_82_U7236 ( .A1(u5_mult_82_ab_48__37_), .A2(
        u5_mult_82_SUMB_47__38_), .ZN(u5_mult_82_n2701) );
  NAND2_X1 u5_mult_82_U7235 ( .A1(u5_mult_82_CARRYB_47__37_), .A2(
        u5_mult_82_SUMB_47__38_), .ZN(u5_mult_82_n2700) );
  XOR2_X1 u5_mult_82_U7234 ( .A(u5_mult_82_SUMB_47__38_), .B(u5_mult_82_n2699), 
        .Z(u5_mult_82_SUMB_48__37_) );
  XOR2_X2 u5_mult_82_U7233 ( .A(u5_mult_82_CARRYB_47__37_), .B(
        u5_mult_82_ab_48__37_), .Z(u5_mult_82_n2699) );
  NAND3_X2 u5_mult_82_U7232 ( .A1(u5_mult_82_n2696), .A2(u5_mult_82_n2697), 
        .A3(u5_mult_82_n2698), .ZN(u5_mult_82_CARRYB_51__34_) );
  NAND2_X1 u5_mult_82_U7231 ( .A1(u5_mult_82_CARRYB_50__34_), .A2(
        u5_mult_82_SUMB_50__35_), .ZN(u5_mult_82_n2698) );
  NAND2_X1 u5_mult_82_U7230 ( .A1(u5_mult_82_ab_51__34_), .A2(
        u5_mult_82_SUMB_50__35_), .ZN(u5_mult_82_n2697) );
  NAND3_X2 u5_mult_82_U7229 ( .A1(u5_mult_82_n2693), .A2(u5_mult_82_n2694), 
        .A3(u5_mult_82_n2695), .ZN(u5_mult_82_CARRYB_50__35_) );
  NAND2_X1 u5_mult_82_U7228 ( .A1(u5_mult_82_ab_50__35_), .A2(
        u5_mult_82_SUMB_49__36_), .ZN(u5_mult_82_n2694) );
  XOR2_X2 u5_mult_82_U7227 ( .A(u5_mult_82_n2692), .B(u5_mult_82_SUMB_49__36_), 
        .Z(u5_mult_82_SUMB_50__35_) );
  XOR2_X2 u5_mult_82_U7226 ( .A(u5_mult_82_ab_50__35_), .B(
        u5_mult_82_CARRYB_49__35_), .Z(u5_mult_82_n2692) );
  INV_X32 u5_mult_82_U7225 ( .A(u5_mult_82_n6789), .ZN(u5_mult_82_n6795) );
  XNOR2_X2 u5_mult_82_U7224 ( .A(u5_mult_82_n2691), .B(u5_mult_82_SUMB_31__41_), .ZN(u5_mult_82_SUMB_32__40_) );
  NAND2_X2 u5_mult_82_U7223 ( .A1(u5_mult_82_ab_21__9_), .A2(
        u5_mult_82_SUMB_20__10_), .ZN(u5_mult_82_n3725) );
  NAND2_X2 u5_mult_82_U7222 ( .A1(u5_mult_82_CARRYB_40__1_), .A2(
        u5_mult_82_ab_41__1_), .ZN(u5_mult_82_n4529) );
  NAND3_X2 u5_mult_82_U7221 ( .A1(u5_mult_82_n2687), .A2(u5_mult_82_n2688), 
        .A3(u5_mult_82_n2689), .ZN(u5_mult_82_CARRYB_2__45_) );
  NAND2_X2 u5_mult_82_U7220 ( .A1(u5_mult_82_ab_2__45_), .A2(
        u5_mult_82_SUMB_1__46_), .ZN(u5_mult_82_n2688) );
  NAND2_X1 u5_mult_82_U7219 ( .A1(u5_mult_82_CARRYB_1__45_), .A2(
        u5_mult_82_SUMB_1__46_), .ZN(u5_mult_82_n2687) );
  XOR2_X2 u5_mult_82_U7218 ( .A(u5_mult_82_SUMB_1__46_), .B(u5_mult_82_n2686), 
        .Z(u5_mult_82_SUMB_2__45_) );
  XOR2_X2 u5_mult_82_U7217 ( .A(u5_mult_82_CARRYB_1__45_), .B(
        u5_mult_82_ab_2__45_), .Z(u5_mult_82_n2686) );
  NAND3_X4 u5_mult_82_U7216 ( .A1(u5_mult_82_n2683), .A2(u5_mult_82_n2684), 
        .A3(u5_mult_82_n2685), .ZN(u5_mult_82_CARRYB_28__39_) );
  NAND2_X2 u5_mult_82_U7215 ( .A1(u5_mult_82_CARRYB_27__39_), .A2(
        u5_mult_82_SUMB_27__40_), .ZN(u5_mult_82_n2685) );
  NAND2_X2 u5_mult_82_U7214 ( .A1(u5_mult_82_ab_28__39_), .A2(
        u5_mult_82_SUMB_27__40_), .ZN(u5_mult_82_n2684) );
  NAND2_X2 u5_mult_82_U7213 ( .A1(u5_mult_82_ab_28__39_), .A2(
        u5_mult_82_CARRYB_27__39_), .ZN(u5_mult_82_n2683) );
  NAND2_X2 u5_mult_82_U7212 ( .A1(u5_mult_82_CARRYB_26__40_), .A2(
        u5_mult_82_SUMB_26__41_), .ZN(u5_mult_82_n2682) );
  NAND2_X2 u5_mult_82_U7211 ( .A1(u5_mult_82_ab_27__40_), .A2(
        u5_mult_82_SUMB_26__41_), .ZN(u5_mult_82_n2681) );
  NAND2_X1 u5_mult_82_U7210 ( .A1(u5_mult_82_ab_27__40_), .A2(
        u5_mult_82_CARRYB_26__40_), .ZN(u5_mult_82_n2680) );
  XOR2_X2 u5_mult_82_U7209 ( .A(u5_mult_82_n2679), .B(u5_mult_82_SUMB_26__41_), 
        .Z(u5_mult_82_SUMB_27__40_) );
  XOR2_X2 u5_mult_82_U7208 ( .A(u5_mult_82_ab_27__40_), .B(
        u5_mult_82_CARRYB_26__40_), .Z(u5_mult_82_n2679) );
  NAND2_X2 u5_mult_82_U7207 ( .A1(u5_mult_82_ab_40__5_), .A2(
        u5_mult_82_SUMB_39__6_), .ZN(u5_mult_82_n4967) );
  XOR2_X2 u5_mult_82_U7206 ( .A(u5_mult_82_n3946), .B(u5_mult_82_SUMB_22__44_), 
        .Z(u5_mult_82_SUMB_23__43_) );
  NAND3_X4 u5_mult_82_U7205 ( .A1(u5_mult_82_n4572), .A2(u5_mult_82_n4571), 
        .A3(u5_mult_82_n4570), .ZN(u5_mult_82_CARRYB_45__28_) );
  XNOR2_X2 u5_mult_82_U7204 ( .A(u5_mult_82_ab_36__8_), .B(
        u5_mult_82_CARRYB_35__8_), .ZN(u5_mult_82_n2678) );
  XNOR2_X2 u5_mult_82_U7203 ( .A(u5_mult_82_n2678), .B(u5_mult_82_SUMB_35__9_), 
        .ZN(u5_mult_82_SUMB_36__8_) );
  XNOR2_X2 u5_mult_82_U7202 ( .A(u5_mult_82_n5648), .B(u5_mult_82_SUMB_27__37_), .ZN(u5_mult_82_SUMB_28__36_) );
  NAND2_X1 u5_mult_82_U7201 ( .A1(u5_mult_82_CARRYB_8__42_), .A2(
        u5_mult_82_SUMB_8__43_), .ZN(u5_mult_82_n4999) );
  XNOR2_X2 u5_mult_82_U7200 ( .A(u5_mult_82_n4867), .B(u5_mult_82_SUMB_25__29_), .ZN(u5_mult_82_SUMB_26__28_) );
  XOR2_X2 u5_mult_82_U7199 ( .A(u5_mult_82_ab_22__30_), .B(
        u5_mult_82_CARRYB_21__30_), .Z(u5_mult_82_n3143) );
  NAND3_X2 u5_mult_82_U7198 ( .A1(u5_mult_82_n4388), .A2(u5_mult_82_n4389), 
        .A3(u5_mult_82_n4390), .ZN(u5_mult_82_CARRYB_47__20_) );
  XNOR2_X2 u5_mult_82_U7197 ( .A(u5_mult_82_CARRYB_45__36_), .B(
        u5_mult_82_ab_46__36_), .ZN(u5_mult_82_n2677) );
  XNOR2_X2 u5_mult_82_U7196 ( .A(u5_mult_82_SUMB_45__37_), .B(u5_mult_82_n2677), .ZN(u5_mult_82_SUMB_46__36_) );
  XNOR2_X2 u5_mult_82_U7195 ( .A(u5_mult_82_CARRYB_29__10_), .B(
        u5_mult_82_n2676), .ZN(u5_mult_82_n3212) );
  NOR2_X2 u5_mult_82_U7194 ( .A1(u5_mult_82_n7007), .A2(u5_mult_82_net66107), 
        .ZN(u5_mult_82_ab_1__46_) );
  NAND2_X2 u5_mult_82_U7193 ( .A1(u5_mult_82_ab_33__8_), .A2(
        u5_mult_82_CARRYB_32__8_), .ZN(u5_mult_82_n3738) );
  NOR2_X1 u5_mult_82_U7192 ( .A1(u5_mult_82_net64415), .A2(u5_mult_82_n6695), 
        .ZN(u5_mult_82_ab_32__8_) );
  NAND2_X1 u5_mult_82_U7191 ( .A1(u5_mult_82_ab_32__8_), .A2(
        u5_mult_82_CARRYB_31__8_), .ZN(u5_mult_82_n2675) );
  NAND2_X2 u5_mult_82_U7190 ( .A1(u5_mult_82_ab_32__8_), .A2(
        u5_mult_82_SUMB_31__9_), .ZN(u5_mult_82_n2674) );
  NAND2_X2 u5_mult_82_U7189 ( .A1(u5_mult_82_CARRYB_31__8_), .A2(
        u5_mult_82_SUMB_31__9_), .ZN(u5_mult_82_n2673) );
  NAND3_X2 u5_mult_82_U7188 ( .A1(u5_mult_82_n2668), .A2(u5_mult_82_n2669), 
        .A3(u5_mult_82_n2670), .ZN(u5_mult_82_CARRYB_40__3_) );
  XOR2_X2 u5_mult_82_U7187 ( .A(u5_mult_82_CARRYB_39__3_), .B(
        u5_mult_82_ab_40__3_), .Z(u5_mult_82_n2667) );
  NAND3_X2 u5_mult_82_U7186 ( .A1(u5_mult_82_n2664), .A2(u5_mult_82_n2665), 
        .A3(u5_mult_82_n2666), .ZN(u5_mult_82_CARRYB_41__39_) );
  NAND2_X1 u5_mult_82_U7185 ( .A1(u5_mult_82_CARRYB_40__39_), .A2(
        u5_mult_82_SUMB_40__40_), .ZN(u5_mult_82_n2666) );
  NAND2_X1 u5_mult_82_U7184 ( .A1(u5_mult_82_ab_41__39_), .A2(
        u5_mult_82_SUMB_40__40_), .ZN(u5_mult_82_n2665) );
  NAND2_X1 u5_mult_82_U7183 ( .A1(u5_mult_82_ab_41__39_), .A2(
        u5_mult_82_CARRYB_40__39_), .ZN(u5_mult_82_n2664) );
  NAND3_X2 u5_mult_82_U7182 ( .A1(u5_mult_82_n2661), .A2(u5_mult_82_n2662), 
        .A3(u5_mult_82_n2663), .ZN(u5_mult_82_CARRYB_40__40_) );
  NAND2_X2 u5_mult_82_U7181 ( .A1(u5_mult_82_CARRYB_39__40_), .A2(
        u5_mult_82_SUMB_39__41_), .ZN(u5_mult_82_n2663) );
  NAND2_X2 u5_mult_82_U7180 ( .A1(u5_mult_82_ab_40__40_), .A2(
        u5_mult_82_SUMB_39__41_), .ZN(u5_mult_82_n2662) );
  NAND2_X1 u5_mult_82_U7179 ( .A1(u5_mult_82_ab_40__40_), .A2(
        u5_mult_82_CARRYB_39__40_), .ZN(u5_mult_82_n2661) );
  XOR2_X2 u5_mult_82_U7178 ( .A(u5_mult_82_n2660), .B(u5_mult_82_SUMB_40__40_), 
        .Z(u5_mult_82_SUMB_41__39_) );
  XOR2_X2 u5_mult_82_U7177 ( .A(u5_mult_82_ab_41__39_), .B(
        u5_mult_82_CARRYB_40__39_), .Z(u5_mult_82_n2660) );
  XOR2_X2 u5_mult_82_U7176 ( .A(u5_mult_82_n2659), .B(u5_mult_82_SUMB_39__41_), 
        .Z(u5_mult_82_SUMB_40__40_) );
  XOR2_X2 u5_mult_82_U7175 ( .A(u5_mult_82_ab_40__40_), .B(
        u5_mult_82_CARRYB_39__40_), .Z(u5_mult_82_n2659) );
  NAND3_X4 u5_mult_82_U7174 ( .A1(u5_mult_82_n2656), .A2(u5_mult_82_n2657), 
        .A3(u5_mult_82_n2658), .ZN(u5_mult_82_CARRYB_46__34_) );
  NAND2_X1 u5_mult_82_U7173 ( .A1(u5_mult_82_ab_46__34_), .A2(
        u5_mult_82_SUMB_45__35_), .ZN(u5_mult_82_n2657) );
  NAND2_X1 u5_mult_82_U7172 ( .A1(u5_mult_82_ab_46__34_), .A2(
        u5_mult_82_CARRYB_45__34_), .ZN(u5_mult_82_n2656) );
  NAND3_X4 u5_mult_82_U7171 ( .A1(u5_mult_82_n2653), .A2(u5_mult_82_n2654), 
        .A3(u5_mult_82_n2655), .ZN(u5_mult_82_CARRYB_45__35_) );
  NAND2_X2 u5_mult_82_U7170 ( .A1(u5_mult_82_CARRYB_44__35_), .A2(
        u5_mult_82_SUMB_44__36_), .ZN(u5_mult_82_n2655) );
  NAND2_X2 u5_mult_82_U7169 ( .A1(u5_mult_82_ab_45__35_), .A2(
        u5_mult_82_SUMB_44__36_), .ZN(u5_mult_82_n2654) );
  XOR2_X2 u5_mult_82_U7168 ( .A(u5_mult_82_n2652), .B(u5_mult_82_SUMB_44__36_), 
        .Z(u5_mult_82_SUMB_45__35_) );
  XOR2_X2 u5_mult_82_U7167 ( .A(u5_mult_82_ab_45__35_), .B(
        u5_mult_82_CARRYB_44__35_), .Z(u5_mult_82_n2652) );
  NAND3_X2 u5_mult_82_U7166 ( .A1(u5_mult_82_n2649), .A2(u5_mult_82_n2650), 
        .A3(u5_mult_82_n2651), .ZN(u5_mult_82_CARRYB_12__14_) );
  NAND2_X1 u5_mult_82_U7165 ( .A1(u5_mult_82_CARRYB_11__14_), .A2(
        u5_mult_82_SUMB_11__15_), .ZN(u5_mult_82_n2651) );
  NAND2_X1 u5_mult_82_U7164 ( .A1(u5_mult_82_ab_12__14_), .A2(
        u5_mult_82_SUMB_11__15_), .ZN(u5_mult_82_n2650) );
  NAND2_X1 u5_mult_82_U7163 ( .A1(u5_mult_82_ab_12__14_), .A2(
        u5_mult_82_CARRYB_11__14_), .ZN(u5_mult_82_n2649) );
  NAND3_X2 u5_mult_82_U7162 ( .A1(u5_mult_82_n2646), .A2(u5_mult_82_n2647), 
        .A3(u5_mult_82_n2648), .ZN(u5_mult_82_CARRYB_11__15_) );
  NAND2_X2 u5_mult_82_U7161 ( .A1(u5_mult_82_CARRYB_10__15_), .A2(
        u5_mult_82_n1660), .ZN(u5_mult_82_n2648) );
  NAND2_X2 u5_mult_82_U7160 ( .A1(u5_mult_82_ab_11__15_), .A2(u5_mult_82_n1660), .ZN(u5_mult_82_n2647) );
  NAND2_X1 u5_mult_82_U7159 ( .A1(u5_mult_82_ab_11__15_), .A2(
        u5_mult_82_CARRYB_10__15_), .ZN(u5_mult_82_n2646) );
  XOR2_X2 u5_mult_82_U7158 ( .A(u5_mult_82_n2645), .B(u5_mult_82_SUMB_11__15_), 
        .Z(u5_mult_82_SUMB_12__14_) );
  XOR2_X2 u5_mult_82_U7157 ( .A(u5_mult_82_ab_12__14_), .B(
        u5_mult_82_CARRYB_11__14_), .Z(u5_mult_82_n2645) );
  XOR2_X2 u5_mult_82_U7156 ( .A(u5_mult_82_ab_11__15_), .B(
        u5_mult_82_CARRYB_10__15_), .Z(u5_mult_82_n2644) );
  XNOR2_X2 u5_mult_82_U7155 ( .A(u5_mult_82_CARRYB_13__42_), .B(
        u5_mult_82_ab_14__42_), .ZN(u5_mult_82_n2643) );
  NOR2_X1 u5_mult_82_U7154 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_net65193), .ZN(u5_mult_82_ab_51__36_) );
  NAND3_X2 u5_mult_82_U7153 ( .A1(u5_mult_82_n2640), .A2(u5_mult_82_n2641), 
        .A3(u5_mult_82_n2642), .ZN(u5_mult_82_CARRYB_35__43_) );
  NAND2_X1 u5_mult_82_U7152 ( .A1(u5_mult_82_SUMB_34__44_), .A2(
        u5_mult_82_CARRYB_34__43_), .ZN(u5_mult_82_n2642) );
  NAND2_X1 u5_mult_82_U7151 ( .A1(u5_mult_82_ab_35__43_), .A2(
        u5_mult_82_SUMB_34__44_), .ZN(u5_mult_82_n2641) );
  NAND2_X1 u5_mult_82_U7150 ( .A1(u5_mult_82_ab_35__43_), .A2(
        u5_mult_82_CARRYB_34__43_), .ZN(u5_mult_82_n2640) );
  NAND3_X2 u5_mult_82_U7149 ( .A1(u5_mult_82_n2637), .A2(u5_mult_82_n2638), 
        .A3(u5_mult_82_n2639), .ZN(u5_mult_82_CARRYB_34__44_) );
  NAND2_X2 u5_mult_82_U7148 ( .A1(u5_mult_82_ab_34__44_), .A2(
        u5_mult_82_SUMB_33__45_), .ZN(u5_mult_82_n2638) );
  NAND2_X1 u5_mult_82_U7147 ( .A1(u5_mult_82_ab_34__44_), .A2(
        u5_mult_82_CARRYB_33__44_), .ZN(u5_mult_82_n2637) );
  XOR2_X2 u5_mult_82_U7146 ( .A(u5_mult_82_n2636), .B(u5_mult_82_SUMB_34__44_), 
        .Z(u5_mult_82_SUMB_35__43_) );
  XOR2_X2 u5_mult_82_U7145 ( .A(u5_mult_82_ab_35__43_), .B(
        u5_mult_82_CARRYB_34__43_), .Z(u5_mult_82_n2636) );
  XOR2_X2 u5_mult_82_U7144 ( .A(u5_mult_82_n2635), .B(u5_mult_82_SUMB_33__45_), 
        .Z(u5_mult_82_SUMB_34__44_) );
  NAND3_X2 u5_mult_82_U7143 ( .A1(u5_mult_82_n2632), .A2(u5_mult_82_n2633), 
        .A3(u5_mult_82_n2634), .ZN(u5_mult_82_CARRYB_51__36_) );
  NAND2_X1 u5_mult_82_U7142 ( .A1(u5_mult_82_ab_51__36_), .A2(
        u5_mult_82_CARRYB_50__36_), .ZN(u5_mult_82_n2634) );
  NAND2_X2 u5_mult_82_U7141 ( .A1(u5_mult_82_ab_51__36_), .A2(
        u5_mult_82_SUMB_50__37_), .ZN(u5_mult_82_n2633) );
  NAND2_X1 u5_mult_82_U7140 ( .A1(u5_mult_82_CARRYB_50__36_), .A2(
        u5_mult_82_SUMB_50__37_), .ZN(u5_mult_82_n2632) );
  XNOR2_X2 u5_mult_82_U7139 ( .A(u5_mult_82_n4164), .B(u5_mult_82_SUMB_38__12_), .ZN(u5_mult_82_SUMB_39__11_) );
  NAND3_X4 u5_mult_82_U7138 ( .A1(u5_mult_82_n6067), .A2(u5_mult_82_n6068), 
        .A3(u5_mult_82_n6069), .ZN(u5_mult_82_CARRYB_41__9_) );
  NAND2_X2 u5_mult_82_U7137 ( .A1(u5_mult_82_CARRYB_38__30_), .A2(
        u5_mult_82_SUMB_38__31_), .ZN(u5_mult_82_n3686) );
  XNOR2_X2 u5_mult_82_U7136 ( .A(u5_mult_82_ab_29__13_), .B(
        u5_mult_82_CARRYB_28__13_), .ZN(u5_mult_82_n2630) );
  XNOR2_X2 u5_mult_82_U7135 ( .A(u5_mult_82_ab_46__34_), .B(
        u5_mult_82_CARRYB_45__34_), .ZN(u5_mult_82_n2629) );
  XNOR2_X2 u5_mult_82_U7134 ( .A(u5_mult_82_n2629), .B(u5_mult_82_SUMB_45__35_), .ZN(u5_mult_82_SUMB_46__34_) );
  NAND2_X2 u5_mult_82_U7133 ( .A1(u5_mult_82_ab_6__29_), .A2(
        u5_mult_82_CARRYB_5__29_), .ZN(u5_mult_82_n4273) );
  NOR2_X1 u5_mult_82_U7132 ( .A1(u5_mult_82_n6864), .A2(u5_mult_82_net66035), 
        .ZN(u5_mult_82_ab_5__29_) );
  NOR2_X1 u5_mult_82_U7131 ( .A1(u5_mult_82_n6870), .A2(u5_mult_82_n6528), 
        .ZN(u5_mult_82_ab_7__28_) );
  NAND3_X4 u5_mult_82_U7130 ( .A1(u5_mult_82_n2626), .A2(u5_mult_82_n2627), 
        .A3(u5_mult_82_n2628), .ZN(u5_mult_82_CARRYB_5__29_) );
  NAND2_X1 u5_mult_82_U7129 ( .A1(u5_mult_82_ab_5__29_), .A2(
        u5_mult_82_CARRYB_4__29_), .ZN(u5_mult_82_n2628) );
  NAND2_X2 u5_mult_82_U7128 ( .A1(u5_mult_82_ab_5__29_), .A2(u5_mult_82_n380), 
        .ZN(u5_mult_82_n2627) );
  NAND2_X2 u5_mult_82_U7127 ( .A1(u5_mult_82_CARRYB_4__29_), .A2(
        u5_mult_82_n380), .ZN(u5_mult_82_n2626) );
  NAND3_X2 u5_mult_82_U7126 ( .A1(u5_mult_82_n2623), .A2(u5_mult_82_n2624), 
        .A3(u5_mult_82_n2625), .ZN(u5_mult_82_CARRYB_7__28_) );
  NAND2_X1 u5_mult_82_U7125 ( .A1(u5_mult_82_ab_7__28_), .A2(
        u5_mult_82_CARRYB_6__28_), .ZN(u5_mult_82_n2625) );
  NAND2_X2 u5_mult_82_U7124 ( .A1(u5_mult_82_ab_7__28_), .A2(
        u5_mult_82_SUMB_6__29_), .ZN(u5_mult_82_n2624) );
  XOR2_X2 u5_mult_82_U7123 ( .A(u5_mult_82_SUMB_6__29_), .B(u5_mult_82_n2622), 
        .Z(u5_mult_82_SUMB_7__28_) );
  XOR2_X2 u5_mult_82_U7122 ( .A(u5_mult_82_CARRYB_6__28_), .B(
        u5_mult_82_ab_7__28_), .Z(u5_mult_82_n2622) );
  NOR2_X1 u5_mult_82_U7121 ( .A1(u5_mult_82_n6779), .A2(u5_mult_82_n6648), 
        .ZN(u5_mult_82_ab_26__48_) );
  NOR2_X1 u5_mult_82_U7120 ( .A1(u5_mult_82_n6779), .A2(u5_mult_82_n1381), 
        .ZN(u5_mult_82_ab_25__48_) );
  NAND3_X2 u5_mult_82_U7119 ( .A1(u5_mult_82_n2619), .A2(u5_mult_82_n2620), 
        .A3(u5_mult_82_n2621), .ZN(u5_mult_82_CARRYB_26__48_) );
  NAND2_X1 u5_mult_82_U7118 ( .A1(u5_mult_82_ab_26__48_), .A2(
        u5_mult_82_CARRYB_25__48_), .ZN(u5_mult_82_n2621) );
  NAND2_X2 u5_mult_82_U7117 ( .A1(u5_mult_82_ab_26__48_), .A2(
        u5_mult_82_SUMB_25__49_), .ZN(u5_mult_82_n2620) );
  NAND2_X1 u5_mult_82_U7116 ( .A1(u5_mult_82_CARRYB_25__48_), .A2(
        u5_mult_82_SUMB_25__49_), .ZN(u5_mult_82_n2619) );
  XOR2_X2 u5_mult_82_U7115 ( .A(u5_mult_82_SUMB_25__49_), .B(u5_mult_82_n2618), 
        .Z(u5_mult_82_SUMB_26__48_) );
  XOR2_X2 u5_mult_82_U7114 ( .A(u5_mult_82_CARRYB_25__48_), .B(
        u5_mult_82_ab_26__48_), .Z(u5_mult_82_n2618) );
  NAND3_X2 u5_mult_82_U7113 ( .A1(u5_mult_82_n2615), .A2(u5_mult_82_n2616), 
        .A3(u5_mult_82_n2617), .ZN(u5_mult_82_CARRYB_25__48_) );
  NAND2_X1 u5_mult_82_U7112 ( .A1(u5_mult_82_ab_25__48_), .A2(
        u5_mult_82_CARRYB_24__48_), .ZN(u5_mult_82_n2617) );
  NAND2_X2 u5_mult_82_U7111 ( .A1(u5_mult_82_ab_25__48_), .A2(
        u5_mult_82_SUMB_24__49_), .ZN(u5_mult_82_n2616) );
  NAND2_X1 u5_mult_82_U7110 ( .A1(u5_mult_82_CARRYB_24__48_), .A2(
        u5_mult_82_SUMB_24__49_), .ZN(u5_mult_82_n2615) );
  XOR2_X2 u5_mult_82_U7109 ( .A(u5_mult_82_SUMB_24__49_), .B(u5_mult_82_n2614), 
        .Z(u5_mult_82_SUMB_25__48_) );
  XOR2_X2 u5_mult_82_U7108 ( .A(u5_mult_82_CARRYB_24__48_), .B(
        u5_mult_82_ab_25__48_), .Z(u5_mult_82_n2614) );
  NAND3_X2 u5_mult_82_U7107 ( .A1(u5_mult_82_n2611), .A2(u5_mult_82_n2612), 
        .A3(u5_mult_82_n2613), .ZN(u5_mult_82_CARRYB_46__33_) );
  NAND2_X2 u5_mult_82_U7106 ( .A1(u5_mult_82_CARRYB_45__33_), .A2(
        u5_mult_82_SUMB_45__34_), .ZN(u5_mult_82_n2613) );
  NAND2_X2 u5_mult_82_U7105 ( .A1(u5_mult_82_ab_46__33_), .A2(
        u5_mult_82_SUMB_45__34_), .ZN(u5_mult_82_n2612) );
  NAND2_X1 u5_mult_82_U7104 ( .A1(u5_mult_82_ab_46__33_), .A2(
        u5_mult_82_CARRYB_45__33_), .ZN(u5_mult_82_n2611) );
  NAND3_X4 u5_mult_82_U7103 ( .A1(u5_mult_82_n2608), .A2(u5_mult_82_n2609), 
        .A3(u5_mult_82_n2610), .ZN(u5_mult_82_CARRYB_45__34_) );
  NAND2_X2 u5_mult_82_U7102 ( .A1(u5_mult_82_ab_45__34_), .A2(
        u5_mult_82_SUMB_44__35_), .ZN(u5_mult_82_n2609) );
  NAND2_X2 u5_mult_82_U7101 ( .A1(u5_mult_82_CARRYB_44__5_), .A2(
        u5_mult_82_SUMB_44__6_), .ZN(u5_mult_82_n4597) );
  NAND3_X2 u5_mult_82_U7100 ( .A1(u5_mult_82_n2605), .A2(u5_mult_82_n2606), 
        .A3(u5_mult_82_n2607), .ZN(u5_mult_82_CARRYB_32__11_) );
  NAND2_X2 u5_mult_82_U7099 ( .A1(u5_mult_82_CARRYB_31__11_), .A2(
        u5_mult_82_SUMB_31__12_), .ZN(u5_mult_82_n2607) );
  NAND2_X2 u5_mult_82_U7098 ( .A1(u5_mult_82_ab_32__11_), .A2(
        u5_mult_82_SUMB_31__12_), .ZN(u5_mult_82_n2606) );
  NAND2_X1 u5_mult_82_U7097 ( .A1(u5_mult_82_ab_32__11_), .A2(
        u5_mult_82_CARRYB_31__11_), .ZN(u5_mult_82_n2605) );
  NAND2_X2 u5_mult_82_U7096 ( .A1(u5_mult_82_n1839), .A2(
        u5_mult_82_CARRYB_30__12_), .ZN(u5_mult_82_n2604) );
  NAND2_X2 u5_mult_82_U7095 ( .A1(u5_mult_82_ab_31__12_), .A2(u5_mult_82_n1839), .ZN(u5_mult_82_n2603) );
  NAND2_X1 u5_mult_82_U7094 ( .A1(u5_mult_82_ab_31__12_), .A2(
        u5_mult_82_CARRYB_30__12_), .ZN(u5_mult_82_n2602) );
  NAND2_X2 u5_mult_82_U7093 ( .A1(u5_mult_82_CARRYB_28__12_), .A2(
        u5_mult_82_SUMB_28__13_), .ZN(u5_mult_82_n2601) );
  NAND2_X2 u5_mult_82_U7092 ( .A1(u5_mult_82_ab_29__12_), .A2(
        u5_mult_82_SUMB_28__13_), .ZN(u5_mult_82_n2600) );
  NAND2_X1 u5_mult_82_U7091 ( .A1(u5_mult_82_ab_29__12_), .A2(
        u5_mult_82_CARRYB_28__12_), .ZN(u5_mult_82_n2599) );
  NAND3_X4 u5_mult_82_U7090 ( .A1(u5_mult_82_n2596), .A2(u5_mult_82_n2597), 
        .A3(u5_mult_82_n2598), .ZN(u5_mult_82_CARRYB_28__13_) );
  NAND2_X2 u5_mult_82_U7089 ( .A1(u5_mult_82_n1848), .A2(u5_mult_82_n394), 
        .ZN(u5_mult_82_n2598) );
  NOR2_X2 u5_mult_82_U7088 ( .A1(u5_mult_82_net64469), .A2(u5_mult_82_net65391), .ZN(u5_mult_82_ab_41__11_) );
  NAND2_X1 u5_mult_82_U7087 ( .A1(u5_mult_82_CARRYB_40__31_), .A2(
        u5_mult_82_SUMB_40__32_), .ZN(u5_mult_82_n3088) );
  NAND2_X1 u5_mult_82_U7086 ( .A1(u5_mult_82_ab_51__24_), .A2(
        u5_mult_82_CARRYB_50__24_), .ZN(u5_mult_82_n4467) );
  NAND2_X1 u5_mult_82_U7085 ( .A1(u5_mult_82_CARRYB_50__24_), .A2(
        u5_mult_82_SUMB_50__25_), .ZN(u5_mult_82_n4469) );
  NAND2_X2 u5_mult_82_U7084 ( .A1(u5_mult_82_SUMB_10__44_), .A2(
        u5_mult_82_CARRYB_10__43_), .ZN(u5_mult_82_n5397) );
  NAND2_X2 u5_mult_82_U7083 ( .A1(u5_mult_82_ab_15__40_), .A2(
        u5_mult_82_SUMB_14__41_), .ZN(u5_mult_82_n6245) );
  NAND2_X2 u5_mult_82_U7082 ( .A1(u5_mult_82_CARRYB_14__40_), .A2(
        u5_mult_82_SUMB_14__41_), .ZN(u5_mult_82_n6246) );
  NAND3_X4 u5_mult_82_U7081 ( .A1(u5_mult_82_n6244), .A2(u5_mult_82_n6245), 
        .A3(u5_mult_82_n6246), .ZN(u5_mult_82_CARRYB_15__40_) );
  NAND2_X2 u5_mult_82_U7080 ( .A1(u5_mult_82_ab_45__5_), .A2(
        u5_mult_82_SUMB_44__6_), .ZN(u5_mult_82_n4596) );
  XNOR2_X2 u5_mult_82_U7079 ( .A(u5_mult_82_ab_43__9_), .B(
        u5_mult_82_CARRYB_42__9_), .ZN(u5_mult_82_n3174) );
  XNOR2_X2 u5_mult_82_U7078 ( .A(u5_mult_82_n5027), .B(u5_mult_82_SUMB_43__9_), 
        .ZN(u5_mult_82_SUMB_44__8_) );
  NAND2_X2 u5_mult_82_U7077 ( .A1(u5_mult_82_n5142), .A2(
        u5_mult_82_SUMB_43__10_), .ZN(u5_mult_82_n2742) );
  NAND2_X4 u5_mult_82_U7076 ( .A1(u5_mult_82_n2742), .A2(u5_mult_82_n2743), 
        .ZN(u5_mult_82_SUMB_44__9_) );
  NAND2_X2 u5_mult_82_U7075 ( .A1(u5_mult_82_ab_17__26_), .A2(
        u5_mult_82_SUMB_16__27_), .ZN(u5_mult_82_n4775) );
  XNOR2_X2 u5_mult_82_U7074 ( .A(u5_mult_82_ab_4__36_), .B(
        u5_mult_82_CARRYB_3__36_), .ZN(u5_mult_82_n2594) );
  NAND2_X2 u5_mult_82_U7073 ( .A1(u5_mult_82_ab_4__37_), .A2(
        u5_mult_82_CARRYB_3__37_), .ZN(u5_mult_82_n5325) );
  NAND3_X2 u5_mult_82_U7072 ( .A1(u5_mult_82_n4104), .A2(u5_mult_82_n4105), 
        .A3(u5_mult_82_n4106), .ZN(u5_mult_82_CARRYB_37__5_) );
  NAND2_X1 u5_mult_82_U7071 ( .A1(u5_mult_82_ab_31__25_), .A2(
        u5_mult_82_CARRYB_30__25_), .ZN(u5_mult_82_n4236) );
  NAND2_X1 u5_mult_82_U7070 ( .A1(u5_mult_82_CARRYB_30__25_), .A2(
        u5_mult_82_SUMB_30__26_), .ZN(u5_mult_82_n4238) );
  INV_X4 u5_mult_82_U7069 ( .A(u5_mult_82_SUMB_52__11_), .ZN(u5_mult_82_n4691)
         );
  XNOR2_X2 u5_mult_82_U7068 ( .A(u5_mult_82_n5256), .B(u5_mult_82_SUMB_50__8_), 
        .ZN(u5_mult_82_SUMB_51__7_) );
  INV_X2 u5_mult_82_U7067 ( .A(u5_mult_82_SUMB_49__12_), .ZN(u5_mult_82_n3540)
         );
  XNOR2_X2 u5_mult_82_U7066 ( .A(u5_mult_82_CARRYB_11__18_), .B(
        u5_mult_82_n2593), .ZN(u5_mult_82_n3315) );
  XNOR2_X2 u5_mult_82_U7065 ( .A(u5_mult_82_n2592), .B(
        u5_mult_82_CARRYB_17__16_), .ZN(u5_mult_82_n4108) );
  XNOR2_X2 u5_mult_82_U7064 ( .A(u5_mult_82_CARRYB_16__18_), .B(
        u5_mult_82_n2591), .ZN(u5_mult_82_n3473) );
  XNOR2_X2 u5_mult_82_U7063 ( .A(u5_mult_82_ab_27__8_), .B(
        u5_mult_82_CARRYB_26__8_), .ZN(u5_mult_82_n2590) );
  XNOR2_X2 u5_mult_82_U7062 ( .A(u5_mult_82_n2590), .B(u5_mult_82_SUMB_26__9_), 
        .ZN(u5_mult_82_SUMB_27__8_) );
  NAND2_X2 u5_mult_82_U7061 ( .A1(u5_mult_82_ab_18__46_), .A2(
        u5_mult_82_SUMB_17__47_), .ZN(u5_mult_82_n5957) );
  NAND2_X2 u5_mult_82_U7060 ( .A1(u5_mult_82_CARRYB_41__6_), .A2(
        u5_mult_82_SUMB_41__7_), .ZN(u5_mult_82_n6008) );
  XNOR2_X2 u5_mult_82_U7059 ( .A(u5_mult_82_CARRYB_15__40_), .B(
        u5_mult_82_ab_16__40_), .ZN(u5_mult_82_n2589) );
  XNOR2_X2 u5_mult_82_U7058 ( .A(u5_mult_82_SUMB_15__41_), .B(u5_mult_82_n2589), .ZN(u5_mult_82_SUMB_16__40_) );
  NOR2_X1 u5_mult_82_U7057 ( .A1(u5_mult_82_n6769), .A2(u5_mult_82_n6585), 
        .ZN(u5_mult_82_ab_15__50_) );
  NAND2_X1 u5_mult_82_U7056 ( .A1(u5_mult_82_SUMB_17__51_), .A2(
        u5_mult_82_CARRYB_17__50_), .ZN(u5_mult_82_n4459) );
  NOR2_X1 u5_mult_82_U7055 ( .A1(u5_mult_82_n6768), .A2(u5_mult_82_n6600), 
        .ZN(u5_mult_82_ab_17__50_) );
  NAND3_X2 u5_mult_82_U7054 ( .A1(u5_mult_82_n2586), .A2(u5_mult_82_n2587), 
        .A3(u5_mult_82_n2588), .ZN(u5_mult_82_CARRYB_15__50_) );
  NAND2_X1 u5_mult_82_U7053 ( .A1(u5_mult_82_ab_15__50_), .A2(
        u5_mult_82_SUMB_14__51_), .ZN(u5_mult_82_n2588) );
  NAND2_X2 u5_mult_82_U7052 ( .A1(u5_mult_82_ab_15__50_), .A2(u5_mult_82_n416), 
        .ZN(u5_mult_82_n2587) );
  NAND2_X2 u5_mult_82_U7051 ( .A1(u5_mult_82_SUMB_14__51_), .A2(
        u5_mult_82_n416), .ZN(u5_mult_82_n2586) );
  XOR2_X2 u5_mult_82_U7050 ( .A(u5_mult_82_n416), .B(u5_mult_82_n2585), .Z(
        u5_mult_82_SUMB_15__50_) );
  XOR2_X2 u5_mult_82_U7049 ( .A(u5_mult_82_SUMB_14__51_), .B(
        u5_mult_82_ab_15__50_), .Z(u5_mult_82_n2585) );
  NAND3_X2 u5_mult_82_U7048 ( .A1(u5_mult_82_n2582), .A2(u5_mult_82_n2583), 
        .A3(u5_mult_82_n2584), .ZN(u5_mult_82_CARRYB_17__50_) );
  NAND2_X1 u5_mult_82_U7047 ( .A1(u5_mult_82_ab_17__50_), .A2(
        u5_mult_82_SUMB_16__51_), .ZN(u5_mult_82_n2584) );
  NAND2_X2 u5_mult_82_U7046 ( .A1(u5_mult_82_CARRYB_16__50_), .A2(
        u5_mult_82_ab_17__50_), .ZN(u5_mult_82_n2583) );
  NAND2_X2 u5_mult_82_U7045 ( .A1(u5_mult_82_SUMB_16__51_), .A2(
        u5_mult_82_CARRYB_16__50_), .ZN(u5_mult_82_n2582) );
  XOR2_X2 u5_mult_82_U7044 ( .A(u5_mult_82_SUMB_16__51_), .B(
        u5_mult_82_ab_17__50_), .Z(u5_mult_82_n2581) );
  NAND3_X2 u5_mult_82_U7043 ( .A1(u5_mult_82_n2578), .A2(u5_mult_82_n2579), 
        .A3(u5_mult_82_n2580), .ZN(u5_mult_82_CARRYB_26__42_) );
  NAND2_X1 u5_mult_82_U7042 ( .A1(u5_mult_82_ab_26__42_), .A2(
        u5_mult_82_SUMB_25__43_), .ZN(u5_mult_82_n2580) );
  NAND2_X1 u5_mult_82_U7041 ( .A1(u5_mult_82_CARRYB_25__42_), .A2(
        u5_mult_82_SUMB_25__43_), .ZN(u5_mult_82_n2579) );
  NAND2_X1 u5_mult_82_U7040 ( .A1(u5_mult_82_CARRYB_25__42_), .A2(
        u5_mult_82_ab_26__42_), .ZN(u5_mult_82_n2578) );
  NAND3_X2 u5_mult_82_U7039 ( .A1(u5_mult_82_n2575), .A2(u5_mult_82_n2576), 
        .A3(u5_mult_82_n2577), .ZN(u5_mult_82_CARRYB_25__43_) );
  NAND2_X2 u5_mult_82_U7038 ( .A1(u5_mult_82_ab_25__43_), .A2(
        u5_mult_82_SUMB_24__44_), .ZN(u5_mult_82_n2576) );
  NAND2_X1 u5_mult_82_U7037 ( .A1(u5_mult_82_ab_25__43_), .A2(
        u5_mult_82_CARRYB_24__43_), .ZN(u5_mult_82_n2575) );
  XOR2_X2 u5_mult_82_U7036 ( .A(u5_mult_82_n2574), .B(u5_mult_82_SUMB_25__43_), 
        .Z(u5_mult_82_SUMB_26__42_) );
  XOR2_X2 u5_mult_82_U7035 ( .A(u5_mult_82_CARRYB_25__42_), .B(
        u5_mult_82_ab_26__42_), .Z(u5_mult_82_n2574) );
  NAND2_X2 u5_mult_82_U7034 ( .A1(u5_mult_82_CARRYB_10__51_), .A2(
        u5_mult_82_ab_10__52_), .ZN(u5_mult_82_n4651) );
  NAND2_X1 u5_mult_82_U7033 ( .A1(u5_mult_82_n1623), .A2(
        u5_mult_82_SUMB_37__23_), .ZN(u5_mult_82_n4804) );
  XNOR2_X2 u5_mult_82_U7032 ( .A(u5_mult_82_ab_11__16_), .B(
        u5_mult_82_CARRYB_10__16_), .ZN(u5_mult_82_n2572) );
  XNOR2_X2 u5_mult_82_U7031 ( .A(u5_mult_82_n2572), .B(u5_mult_82_SUMB_10__17_), .ZN(u5_mult_82_SUMB_11__16_) );
  XNOR2_X2 u5_mult_82_U7030 ( .A(u5_mult_82_n2571), .B(u5_mult_82_SUMB_31__8_), 
        .ZN(u5_mult_82_SUMB_32__7_) );
  NAND3_X4 u5_mult_82_U7029 ( .A1(u5_mult_82_net84888), .A2(u5_mult_82_n2570), 
        .A3(u5_mult_82_net84890), .ZN(u5_mult_82_CARRYB_46__9_) );
  NAND2_X2 u5_mult_82_U7028 ( .A1(u5_mult_82_ab_46__9_), .A2(
        u5_mult_82_SUMB_45__10_), .ZN(u5_mult_82_n2570) );
  NAND3_X4 u5_mult_82_U7027 ( .A1(u5_mult_82_n2567), .A2(u5_mult_82_n2568), 
        .A3(u5_mult_82_n2569), .ZN(u5_mult_82_CARRYB_45__10_) );
  NAND2_X2 u5_mult_82_U7026 ( .A1(u5_mult_82_CARRYB_44__10_), .A2(
        u5_mult_82_SUMB_44__11_), .ZN(u5_mult_82_n2569) );
  NAND2_X2 u5_mult_82_U7025 ( .A1(u5_mult_82_ab_45__10_), .A2(
        u5_mult_82_SUMB_44__11_), .ZN(u5_mult_82_n2568) );
  NAND3_X2 u5_mult_82_U7024 ( .A1(u5_mult_82_n6326), .A2(u5_mult_82_n6325), 
        .A3(u5_mult_82_n6327), .ZN(u5_mult_82_CARRYB_49__5_) );
  XNOR2_X1 u5_mult_82_U7023 ( .A(u5_mult_82_ab_34__5_), .B(
        u5_mult_82_CARRYB_33__5_), .ZN(u5_mult_82_n2566) );
  XNOR2_X2 u5_mult_82_U7022 ( .A(u5_mult_82_CARRYB_34__29_), .B(
        u5_mult_82_n2565), .ZN(u5_mult_82_SUMB_35__29_) );
  XNOR2_X2 u5_mult_82_U7021 ( .A(u5_mult_82_n2564), .B(u5_mult_82_SUMB_20__23_), .ZN(u5_mult_82_SUMB_21__22_) );
  XNOR2_X2 u5_mult_82_U7020 ( .A(u5_mult_82_n3255), .B(u5_mult_82_SUMB_31__25_), .ZN(u5_mult_82_SUMB_32__24_) );
  NAND2_X2 u5_mult_82_U7019 ( .A1(u5_mult_82_n2979), .A2(u5_mult_82_n2980), 
        .ZN(u5_mult_82_n5787) );
  NAND3_X4 u5_mult_82_U7018 ( .A1(u5_mult_82_n5226), .A2(u5_mult_82_n5227), 
        .A3(u5_mult_82_n5228), .ZN(u5_mult_82_CARRYB_33__11_) );
  XNOR2_X2 u5_mult_82_U7017 ( .A(u5_mult_82_n2566), .B(u5_mult_82_n1600), .ZN(
        u5_mult_82_SUMB_34__5_) );
  NAND2_X2 u5_mult_82_U7016 ( .A1(u5_mult_82_ab_35__4_), .A2(
        u5_mult_82_SUMB_34__5_), .ZN(u5_mult_82_n3180) );
  INV_X4 u5_mult_82_U7015 ( .A(u5_mult_82_n4079), .ZN(u5_mult_82_n3783) );
  NAND2_X2 u5_mult_82_U7014 ( .A1(u5_mult_82_n1413), .A2(
        u5_mult_82_SUMB_38__12_), .ZN(u5_mult_82_n5133) );
  NAND2_X1 u5_mult_82_U7013 ( .A1(u5_mult_82_ab_27__29_), .A2(
        u5_mult_82_CARRYB_26__29_), .ZN(u5_mult_82_n6282) );
  NAND2_X2 u5_mult_82_U7012 ( .A1(u5_mult_82_ab_24__9_), .A2(
        u5_mult_82_CARRYB_23__9_), .ZN(u5_mult_82_n3431) );
  NOR2_X1 u5_mult_82_U7011 ( .A1(u5_mult_82_net64435), .A2(u5_mult_82_net65713), .ZN(u5_mult_82_ab_23__9_) );
  NAND2_X1 u5_mult_82_U7010 ( .A1(u5_mult_82_ab_23__9_), .A2(
        u5_mult_82_CARRYB_22__9_), .ZN(u5_mult_82_n2563) );
  NAND2_X1 u5_mult_82_U7009 ( .A1(u5_mult_82_ab_23__9_), .A2(
        u5_mult_82_SUMB_22__10_), .ZN(u5_mult_82_n2562) );
  NAND2_X1 u5_mult_82_U7008 ( .A1(u5_mult_82_CARRYB_22__9_), .A2(
        u5_mult_82_SUMB_22__10_), .ZN(u5_mult_82_n2561) );
  INV_X4 u5_mult_82_U7007 ( .A(u5_mult_82_n3251), .ZN(u5_mult_82_n2557) );
  NAND2_X2 u5_mult_82_U7006 ( .A1(u5_mult_82_n2557), .A2(u5_mult_82_n2558), 
        .ZN(u5_mult_82_n2560) );
  NAND2_X2 u5_mult_82_U7005 ( .A1(u5_mult_82_n3251), .A2(
        u5_mult_82_SUMB_23__10_), .ZN(u5_mult_82_n2559) );
  NAND3_X2 u5_mult_82_U7004 ( .A1(u5_mult_82_n3626), .A2(u5_mult_82_n3627), 
        .A3(u5_mult_82_n3628), .ZN(u5_mult_82_CARRYB_50__16_) );
  XNOR2_X2 u5_mult_82_U7003 ( .A(u5_mult_82_CARRYB_6__44_), .B(
        u5_mult_82_n2556), .ZN(u5_mult_82_n6148) );
  XNOR2_X2 u5_mult_82_U7002 ( .A(u5_mult_82_CARRYB_20__15_), .B(
        u5_mult_82_ab_21__15_), .ZN(u5_mult_82_n2555) );
  XNOR2_X2 u5_mult_82_U7001 ( .A(u5_mult_82_n2555), .B(u5_mult_82_SUMB_20__16_), .ZN(u5_mult_82_SUMB_21__15_) );
  XNOR2_X2 u5_mult_82_U7000 ( .A(u5_mult_82_CARRYB_30__14_), .B(
        u5_mult_82_ab_31__14_), .ZN(u5_mult_82_n2554) );
  XNOR2_X2 u5_mult_82_U6999 ( .A(u5_mult_82_n2554), .B(u5_mult_82_SUMB_30__15_), .ZN(u5_mult_82_SUMB_31__14_) );
  NAND2_X2 u5_mult_82_U6998 ( .A1(u5_mult_82_ab_32__24_), .A2(
        u5_mult_82_SUMB_31__25_), .ZN(u5_mult_82_n4240) );
  NAND2_X2 u5_mult_82_U6997 ( .A1(u5_mult_82_SUMB_44__9_), .A2(
        u5_mult_82_CARRYB_44__8_), .ZN(u5_mult_82_n4219) );
  NAND3_X2 u5_mult_82_U6996 ( .A1(u5_mult_82_n6045), .A2(u5_mult_82_n6046), 
        .A3(u5_mult_82_n6047), .ZN(u5_mult_82_CARRYB_16__33_) );
  NAND2_X2 u5_mult_82_U6995 ( .A1(u5_mult_82_n3481), .A2(u5_mult_82_n3482), 
        .ZN(u5_mult_82_SUMB_42__2_) );
  NOR2_X2 u5_mult_82_U6994 ( .A1(u5_mult_82_n6967), .A2(u5_mult_82_net65355), 
        .ZN(u5_mult_82_ab_43__1_) );
  NOR2_X1 u5_mult_82_U6993 ( .A1(u5_mult_82_n6929), .A2(u5_mult_82_n6536), 
        .ZN(u5_mult_82_ab_8__17_) );
  NAND3_X2 u5_mult_82_U6992 ( .A1(u5_mult_82_n2551), .A2(u5_mult_82_n2552), 
        .A3(u5_mult_82_n2553), .ZN(u5_mult_82_CARRYB_39__1_) );
  NAND2_X2 u5_mult_82_U6991 ( .A1(u5_mult_82_SUMB_38__2_), .A2(
        u5_mult_82_CARRYB_38__1_), .ZN(u5_mult_82_n2553) );
  NAND2_X2 u5_mult_82_U6990 ( .A1(u5_mult_82_ab_39__1_), .A2(
        u5_mult_82_CARRYB_38__1_), .ZN(u5_mult_82_n2552) );
  NAND2_X2 u5_mult_82_U6989 ( .A1(u5_mult_82_ab_39__1_), .A2(
        u5_mult_82_SUMB_38__2_), .ZN(u5_mult_82_n2551) );
  NAND3_X2 u5_mult_82_U6988 ( .A1(u5_mult_82_n2548), .A2(u5_mult_82_n2549), 
        .A3(u5_mult_82_n2550), .ZN(u5_mult_82_CARRYB_38__1_) );
  NAND2_X2 u5_mult_82_U6987 ( .A1(u5_mult_82_ab_38__1_), .A2(
        u5_mult_82_SUMB_37__2_), .ZN(u5_mult_82_n2549) );
  XOR2_X2 u5_mult_82_U6986 ( .A(u5_mult_82_n2547), .B(u5_mult_82_SUMB_37__2_), 
        .Z(u5_mult_82_SUMB_38__1_) );
  NAND3_X2 u5_mult_82_U6985 ( .A1(u5_mult_82_n2544), .A2(u5_mult_82_n2545), 
        .A3(u5_mult_82_n2546), .ZN(u5_mult_82_CARRYB_43__1_) );
  NAND2_X2 u5_mult_82_U6984 ( .A1(u5_mult_82_ab_43__1_), .A2(
        u5_mult_82_CARRYB_42__1_), .ZN(u5_mult_82_n2545) );
  NAND3_X2 u5_mult_82_U6983 ( .A1(u5_mult_82_n2541), .A2(u5_mult_82_n2542), 
        .A3(u5_mult_82_n2543), .ZN(u5_mult_82_CARRYB_10__15_) );
  NAND2_X1 u5_mult_82_U6982 ( .A1(u5_mult_82_CARRYB_9__15_), .A2(
        u5_mult_82_SUMB_9__16_), .ZN(u5_mult_82_n2543) );
  NAND2_X1 u5_mult_82_U6981 ( .A1(u5_mult_82_ab_10__15_), .A2(
        u5_mult_82_SUMB_9__16_), .ZN(u5_mult_82_n2542) );
  NAND2_X1 u5_mult_82_U6980 ( .A1(u5_mult_82_ab_10__15_), .A2(
        u5_mult_82_CARRYB_9__15_), .ZN(u5_mult_82_n2541) );
  NAND3_X2 u5_mult_82_U6979 ( .A1(u5_mult_82_n2538), .A2(u5_mult_82_n2539), 
        .A3(u5_mult_82_n2540), .ZN(u5_mult_82_CARRYB_9__16_) );
  NAND2_X1 u5_mult_82_U6978 ( .A1(u5_mult_82_CARRYB_8__16_), .A2(
        u5_mult_82_SUMB_8__17_), .ZN(u5_mult_82_n2540) );
  NAND2_X1 u5_mult_82_U6977 ( .A1(u5_mult_82_ab_9__16_), .A2(
        u5_mult_82_SUMB_8__17_), .ZN(u5_mult_82_n2539) );
  NAND2_X1 u5_mult_82_U6976 ( .A1(u5_mult_82_ab_9__16_), .A2(
        u5_mult_82_CARRYB_8__16_), .ZN(u5_mult_82_n2538) );
  XOR2_X2 u5_mult_82_U6975 ( .A(u5_mult_82_n2537), .B(u5_mult_82_SUMB_9__16_), 
        .Z(u5_mult_82_SUMB_10__15_) );
  XOR2_X2 u5_mult_82_U6974 ( .A(u5_mult_82_ab_10__15_), .B(
        u5_mult_82_CARRYB_9__15_), .Z(u5_mult_82_n2537) );
  XOR2_X2 u5_mult_82_U6973 ( .A(u5_mult_82_n2536), .B(u5_mult_82_SUMB_8__17_), 
        .Z(u5_mult_82_SUMB_9__16_) );
  XOR2_X2 u5_mult_82_U6972 ( .A(u5_mult_82_ab_9__16_), .B(
        u5_mult_82_CARRYB_8__16_), .Z(u5_mult_82_n2536) );
  NAND3_X2 u5_mult_82_U6971 ( .A1(u5_mult_82_n2533), .A2(u5_mult_82_n2534), 
        .A3(u5_mult_82_n2535), .ZN(u5_mult_82_CARRYB_8__17_) );
  NAND2_X1 u5_mult_82_U6970 ( .A1(u5_mult_82_ab_8__17_), .A2(
        u5_mult_82_CARRYB_7__17_), .ZN(u5_mult_82_n2535) );
  NAND2_X2 u5_mult_82_U6969 ( .A1(u5_mult_82_ab_8__17_), .A2(
        u5_mult_82_SUMB_7__18_), .ZN(u5_mult_82_n2534) );
  NAND2_X1 u5_mult_82_U6968 ( .A1(u5_mult_82_CARRYB_7__17_), .A2(
        u5_mult_82_SUMB_7__18_), .ZN(u5_mult_82_n2533) );
  XOR2_X2 u5_mult_82_U6967 ( .A(u5_mult_82_SUMB_7__18_), .B(u5_mult_82_n2532), 
        .Z(u5_mult_82_SUMB_8__17_) );
  XOR2_X2 u5_mult_82_U6966 ( .A(u5_mult_82_CARRYB_7__17_), .B(
        u5_mult_82_ab_8__17_), .Z(u5_mult_82_n2532) );
  NAND2_X2 u5_mult_82_U6965 ( .A1(u5_mult_82_ab_21__30_), .A2(
        u5_mult_82_SUMB_20__31_), .ZN(u5_mult_82_n2530) );
  NAND2_X1 u5_mult_82_U6964 ( .A1(u5_mult_82_ab_21__30_), .A2(
        u5_mult_82_CARRYB_20__30_), .ZN(u5_mult_82_n2529) );
  NAND3_X2 u5_mult_82_U6963 ( .A1(u5_mult_82_n2526), .A2(u5_mult_82_n2527), 
        .A3(u5_mult_82_n2528), .ZN(u5_mult_82_CARRYB_20__31_) );
  NAND2_X1 u5_mult_82_U6962 ( .A1(u5_mult_82_CARRYB_19__31_), .A2(
        u5_mult_82_SUMB_19__32_), .ZN(u5_mult_82_n2528) );
  NAND2_X1 u5_mult_82_U6961 ( .A1(u5_mult_82_ab_20__31_), .A2(
        u5_mult_82_SUMB_19__32_), .ZN(u5_mult_82_n2527) );
  NAND2_X1 u5_mult_82_U6960 ( .A1(u5_mult_82_ab_20__31_), .A2(
        u5_mult_82_CARRYB_19__31_), .ZN(u5_mult_82_n2526) );
  NAND2_X2 u5_mult_82_U6959 ( .A1(u5_mult_82_ab_22__44_), .A2(
        u5_mult_82_CARRYB_21__44_), .ZN(u5_mult_82_n3947) );
  NAND2_X2 u5_mult_82_U6958 ( .A1(u5_mult_82_SUMB_49__25_), .A2(
        u5_mult_82_CARRYB_49__24_), .ZN(u5_mult_82_n4447) );
  NAND3_X2 u5_mult_82_U6957 ( .A1(u5_mult_82_n3088), .A2(u5_mult_82_n3089), 
        .A3(u5_mult_82_n3090), .ZN(u5_mult_82_CARRYB_41__31_) );
  XOR2_X2 u5_mult_82_U6956 ( .A(u5_mult_82_CARRYB_43__26_), .B(
        u5_mult_82_ab_44__26_), .Z(u5_mult_82_n4920) );
  NAND2_X2 u5_mult_82_U6955 ( .A1(u5_mult_82_CARRYB_17__36_), .A2(
        u5_mult_82_SUMB_17__37_), .ZN(u5_mult_82_n5040) );
  INV_X4 u5_mult_82_U6954 ( .A(u5_mult_82_n3278), .ZN(u5_mult_82_n2523) );
  INV_X1 u5_mult_82_U6953 ( .A(u5_mult_82_CARRYB_7__45_), .ZN(u5_mult_82_n2522) );
  INV_X1 u5_mult_82_U6952 ( .A(u5_mult_82_n1794), .ZN(u5_mult_82_n2518) );
  NAND2_X2 u5_mult_82_U6951 ( .A1(u5_mult_82_n2520), .A2(u5_mult_82_n2521), 
        .ZN(u5_mult_82_SUMB_14__42_) );
  NAND2_X2 u5_mult_82_U6950 ( .A1(u5_mult_82_n2518), .A2(u5_mult_82_n2519), 
        .ZN(u5_mult_82_n2521) );
  NAND2_X1 u5_mult_82_U6949 ( .A1(u5_mult_82_n1794), .A2(u5_mult_82_n2643), 
        .ZN(u5_mult_82_n2520) );
  NAND3_X2 u5_mult_82_U6948 ( .A1(u5_mult_82_n2515), .A2(u5_mult_82_n2516), 
        .A3(u5_mult_82_n2517), .ZN(u5_mult_82_CARRYB_41__26_) );
  NAND2_X1 u5_mult_82_U6947 ( .A1(u5_mult_82_ab_41__26_), .A2(
        u5_mult_82_SUMB_40__27_), .ZN(u5_mult_82_n2517) );
  NAND2_X1 u5_mult_82_U6946 ( .A1(u5_mult_82_n1450), .A2(
        u5_mult_82_SUMB_40__27_), .ZN(u5_mult_82_n2516) );
  NAND2_X1 u5_mult_82_U6945 ( .A1(u5_mult_82_n1450), .A2(u5_mult_82_ab_41__26_), .ZN(u5_mult_82_n2515) );
  NAND3_X4 u5_mult_82_U6944 ( .A1(u5_mult_82_n2512), .A2(u5_mult_82_n2513), 
        .A3(u5_mult_82_n2514), .ZN(u5_mult_82_CARRYB_40__27_) );
  NAND2_X2 u5_mult_82_U6943 ( .A1(u5_mult_82_n706), .A2(
        u5_mult_82_SUMB_39__28_), .ZN(u5_mult_82_n2514) );
  NAND2_X2 u5_mult_82_U6942 ( .A1(u5_mult_82_ab_40__27_), .A2(
        u5_mult_82_SUMB_39__28_), .ZN(u5_mult_82_n2513) );
  NAND2_X2 u5_mult_82_U6941 ( .A1(u5_mult_82_ab_40__27_), .A2(u5_mult_82_n706), 
        .ZN(u5_mult_82_n2512) );
  XOR2_X2 u5_mult_82_U6940 ( .A(u5_mult_82_n2511), .B(u5_mult_82_SUMB_40__27_), 
        .Z(u5_mult_82_SUMB_41__26_) );
  XOR2_X2 u5_mult_82_U6939 ( .A(u5_mult_82_CARRYB_40__26_), .B(
        u5_mult_82_ab_41__26_), .Z(u5_mult_82_n2511) );
  XOR2_X2 u5_mult_82_U6938 ( .A(u5_mult_82_n2510), .B(u5_mult_82_SUMB_39__28_), 
        .Z(u5_mult_82_SUMB_40__27_) );
  XOR2_X2 u5_mult_82_U6937 ( .A(u5_mult_82_n706), .B(u5_mult_82_ab_40__27_), 
        .Z(u5_mult_82_n2510) );
  XNOR2_X2 u5_mult_82_U6936 ( .A(u5_mult_82_ab_49__6_), .B(
        u5_mult_82_CARRYB_48__6_), .ZN(u5_mult_82_net84845) );
  NOR2_X2 u5_mult_82_U6935 ( .A1(u5_mult_82_n6824), .A2(u5_mult_82_net66087), 
        .ZN(u5_mult_82_ab_2__41_) );
  NAND2_X2 u5_mult_82_U6934 ( .A1(u5_mult_82_ab_9__28_), .A2(
        u5_mult_82_CARRYB_8__28_), .ZN(u5_mult_82_n3446) );
  NOR2_X1 u5_mult_82_U6933 ( .A1(u5_mult_82_n6870), .A2(u5_mult_82_n6535), 
        .ZN(u5_mult_82_ab_8__28_) );
  NOR2_X4 u5_mult_82_U6932 ( .A1(u5_mult_82_net64415), .A2(u5_mult_82_net65355), .ZN(u5_mult_82_ab_43__8_) );
  NAND2_X1 u5_mult_82_U6931 ( .A1(u5_mult_82_ab_8__28_), .A2(
        u5_mult_82_CARRYB_7__28_), .ZN(u5_mult_82_n2509) );
  XOR2_X2 u5_mult_82_U6930 ( .A(u5_mult_82_SUMB_7__29_), .B(u5_mult_82_n2506), 
        .Z(u5_mult_82_SUMB_8__28_) );
  XOR2_X2 u5_mult_82_U6929 ( .A(u5_mult_82_CARRYB_7__28_), .B(
        u5_mult_82_ab_8__28_), .Z(u5_mult_82_n2506) );
  INV_X2 u5_mult_82_U6928 ( .A(u5_mult_82_ab_43__8_), .ZN(u5_mult_82_n2503) );
  INV_X4 u5_mult_82_U6927 ( .A(u5_mult_82_SUMB_42__9_), .ZN(u5_mult_82_n2502)
         );
  NAND2_X4 u5_mult_82_U6926 ( .A1(u5_mult_82_n2504), .A2(u5_mult_82_n2505), 
        .ZN(u5_mult_82_n5257) );
  NAND2_X4 u5_mult_82_U6925 ( .A1(u5_mult_82_n2502), .A2(u5_mult_82_n2503), 
        .ZN(u5_mult_82_n2505) );
  NAND2_X2 u5_mult_82_U6924 ( .A1(u5_mult_82_n1469), .A2(u5_mult_82_ab_43__8_), 
        .ZN(u5_mult_82_n2504) );
  NAND2_X2 u5_mult_82_U6923 ( .A1(u5_mult_82_ab_0__42_), .A2(
        u5_mult_82_ab_1__41_), .ZN(u5_mult_82_n6494) );
  XOR2_X2 u5_mult_82_U6922 ( .A(u5_mult_82_ab_41__30_), .B(
        u5_mult_82_CARRYB_40__30_), .Z(u5_mult_82_n4418) );
  XNOR2_X2 u5_mult_82_U6921 ( .A(u5_mult_82_n2501), .B(
        u5_mult_82_CARRYB_21__13_), .ZN(u5_mult_82_n2856) );
  XNOR2_X2 u5_mult_82_U6920 ( .A(u5_mult_82_ab_16__36_), .B(
        u5_mult_82_CARRYB_15__36_), .ZN(u5_mult_82_n2500) );
  XNOR2_X2 u5_mult_82_U6919 ( .A(u5_mult_82_n2500), .B(u5_mult_82_n1827), .ZN(
        u5_mult_82_SUMB_16__36_) );
  NAND2_X2 u5_mult_82_U6918 ( .A1(u5_mult_82_CARRYB_21__9_), .A2(
        u5_mult_82_SUMB_21__10_), .ZN(u5_mult_82_n3728) );
  NAND2_X2 u5_mult_82_U6917 ( .A1(u5_mult_82_CARRYB_23__40_), .A2(
        u5_mult_82_SUMB_23__41_), .ZN(u5_mult_82_n3032) );
  XNOR2_X1 u5_mult_82_U6916 ( .A(u5_mult_82_ab_12__41_), .B(
        u5_mult_82_CARRYB_11__41_), .ZN(u5_mult_82_n2499) );
  XNOR2_X2 u5_mult_82_U6915 ( .A(u5_mult_82_n2499), .B(u5_mult_82_SUMB_11__42_), .ZN(u5_mult_82_SUMB_12__41_) );
  XNOR2_X2 u5_mult_82_U6914 ( .A(u5_mult_82_CARRYB_22__43_), .B(
        u5_mult_82_n2498), .ZN(u5_mult_82_n3946) );
  XOR2_X2 u5_mult_82_U6913 ( .A(u5_mult_82_n5580), .B(u5_mult_82_SUMB_40__29_), 
        .Z(u5_mult_82_SUMB_41__28_) );
  NAND3_X4 u5_mult_82_U6912 ( .A1(u5_mult_82_n4439), .A2(u5_mult_82_n4440), 
        .A3(u5_mult_82_n4441), .ZN(u5_mult_82_CARRYB_26__34_) );
  NAND3_X4 u5_mult_82_U6911 ( .A1(u5_mult_82_n5741), .A2(u5_mult_82_n5742), 
        .A3(u5_mult_82_n5743), .ZN(u5_mult_82_CARRYB_50__18_) );
  XNOR2_X2 u5_mult_82_U6910 ( .A(u5_mult_82_ab_18__25_), .B(
        u5_mult_82_CARRYB_17__25_), .ZN(u5_mult_82_n2497) );
  XNOR2_X2 u5_mult_82_U6909 ( .A(u5_mult_82_n2497), .B(u5_mult_82_SUMB_17__26_), .ZN(u5_mult_82_SUMB_18__25_) );
  NAND2_X2 u5_mult_82_U6908 ( .A1(u5_mult_82_SUMB_37__31_), .A2(
        u5_mult_82_n1475), .ZN(u5_mult_82_n4713) );
  NAND3_X4 u5_mult_82_U6907 ( .A1(u5_mult_82_n2494), .A2(u5_mult_82_n2495), 
        .A3(u5_mult_82_n2496), .ZN(u5_mult_82_CARRYB_35__42_) );
  NAND2_X2 u5_mult_82_U6906 ( .A1(u5_mult_82_CARRYB_34__42_), .A2(
        u5_mult_82_SUMB_34__43_), .ZN(u5_mult_82_n2496) );
  NAND2_X2 u5_mult_82_U6905 ( .A1(u5_mult_82_ab_35__42_), .A2(
        u5_mult_82_SUMB_34__43_), .ZN(u5_mult_82_n2495) );
  NAND2_X1 u5_mult_82_U6904 ( .A1(u5_mult_82_ab_35__42_), .A2(
        u5_mult_82_CARRYB_34__42_), .ZN(u5_mult_82_n2494) );
  NAND3_X4 u5_mult_82_U6903 ( .A1(u5_mult_82_n2493), .A2(u5_mult_82_n2492), 
        .A3(u5_mult_82_n2491), .ZN(u5_mult_82_CARRYB_34__43_) );
  NAND2_X2 u5_mult_82_U6902 ( .A1(u5_mult_82_CARRYB_33__43_), .A2(
        u5_mult_82_SUMB_33__44_), .ZN(u5_mult_82_n2493) );
  NAND2_X2 u5_mult_82_U6901 ( .A1(u5_mult_82_ab_34__43_), .A2(
        u5_mult_82_SUMB_33__44_), .ZN(u5_mult_82_n2492) );
  NAND2_X1 u5_mult_82_U6900 ( .A1(u5_mult_82_ab_34__43_), .A2(
        u5_mult_82_CARRYB_33__43_), .ZN(u5_mult_82_n2491) );
  XOR2_X2 u5_mult_82_U6899 ( .A(u5_mult_82_n2490), .B(u5_mult_82_SUMB_34__43_), 
        .Z(u5_mult_82_SUMB_35__42_) );
  XOR2_X2 u5_mult_82_U6898 ( .A(u5_mult_82_ab_35__42_), .B(
        u5_mult_82_CARRYB_34__42_), .Z(u5_mult_82_n2490) );
  XOR2_X2 u5_mult_82_U6897 ( .A(u5_mult_82_n2489), .B(u5_mult_82_n1508), .Z(
        u5_mult_82_SUMB_34__43_) );
  XOR2_X1 u5_mult_82_U6896 ( .A(u5_mult_82_ab_34__43_), .B(
        u5_mult_82_CARRYB_33__43_), .Z(u5_mult_82_n2489) );
  NAND3_X2 u5_mult_82_U6895 ( .A1(u5_mult_82_n2486), .A2(u5_mult_82_n2487), 
        .A3(u5_mult_82_n2488), .ZN(u5_mult_82_CARRYB_26__46_) );
  NAND2_X1 u5_mult_82_U6894 ( .A1(u5_mult_82_CARRYB_25__46_), .A2(
        u5_mult_82_SUMB_25__47_), .ZN(u5_mult_82_n2488) );
  NAND2_X1 u5_mult_82_U6893 ( .A1(u5_mult_82_ab_26__46_), .A2(
        u5_mult_82_SUMB_25__47_), .ZN(u5_mult_82_n2487) );
  NAND2_X1 u5_mult_82_U6892 ( .A1(u5_mult_82_ab_26__46_), .A2(
        u5_mult_82_CARRYB_25__46_), .ZN(u5_mult_82_n2486) );
  NAND3_X2 u5_mult_82_U6891 ( .A1(u5_mult_82_n2483), .A2(u5_mult_82_n2484), 
        .A3(u5_mult_82_n2485), .ZN(u5_mult_82_CARRYB_25__47_) );
  NAND2_X2 u5_mult_82_U6890 ( .A1(u5_mult_82_ab_25__47_), .A2(
        u5_mult_82_SUMB_24__48_), .ZN(u5_mult_82_n2485) );
  NAND2_X1 u5_mult_82_U6889 ( .A1(u5_mult_82_CARRYB_24__47_), .A2(
        u5_mult_82_SUMB_24__48_), .ZN(u5_mult_82_n2484) );
  NAND2_X1 u5_mult_82_U6888 ( .A1(u5_mult_82_CARRYB_24__47_), .A2(
        u5_mult_82_ab_25__47_), .ZN(u5_mult_82_n2483) );
  XOR2_X2 u5_mult_82_U6887 ( .A(u5_mult_82_n2482), .B(u5_mult_82_SUMB_25__47_), 
        .Z(u5_mult_82_SUMB_26__46_) );
  XOR2_X2 u5_mult_82_U6886 ( .A(u5_mult_82_ab_26__46_), .B(
        u5_mult_82_CARRYB_25__46_), .Z(u5_mult_82_n2482) );
  XOR2_X2 u5_mult_82_U6885 ( .A(u5_mult_82_n2481), .B(u5_mult_82_SUMB_24__48_), 
        .Z(u5_mult_82_SUMB_25__47_) );
  XOR2_X2 u5_mult_82_U6884 ( .A(u5_mult_82_CARRYB_24__47_), .B(
        u5_mult_82_ab_25__47_), .Z(u5_mult_82_n2481) );
  INV_X16 u5_mult_82_U6883 ( .A(u5_mult_82_n6820), .ZN(u5_mult_82_n2480) );
  NAND3_X4 u5_mult_82_U6882 ( .A1(u5_mult_82_n5599), .A2(u5_mult_82_n5600), 
        .A3(u5_mult_82_n5601), .ZN(u5_mult_82_CARRYB_33__32_) );
  NAND3_X2 u5_mult_82_U6881 ( .A1(u5_mult_82_n5976), .A2(u5_mult_82_n5977), 
        .A3(u5_mult_82_n5978), .ZN(u5_mult_82_CARRYB_7__42_) );
  NAND2_X2 u5_mult_82_U6880 ( .A1(u5_mult_82_ab_21__14_), .A2(
        u5_mult_82_CARRYB_20__14_), .ZN(u5_mult_82_n2857) );
  NOR2_X2 u5_mult_82_U6879 ( .A1(u5_mult_82_net64525), .A2(u5_mult_82_n6623), 
        .ZN(u5_mult_82_ab_20__14_) );
  NAND3_X4 u5_mult_82_U6878 ( .A1(u5_mult_82_n2479), .A2(u5_mult_82_n2478), 
        .A3(u5_mult_82_n2477), .ZN(u5_mult_82_CARRYB_5__25_) );
  NAND2_X2 u5_mult_82_U6877 ( .A1(u5_mult_82_ab_5__25_), .A2(
        u5_mult_82_SUMB_4__26_), .ZN(u5_mult_82_n2478) );
  NAND2_X1 u5_mult_82_U6876 ( .A1(u5_mult_82_ab_5__25_), .A2(
        u5_mult_82_CARRYB_4__25_), .ZN(u5_mult_82_n2477) );
  NAND3_X2 u5_mult_82_U6875 ( .A1(u5_mult_82_n2474), .A2(u5_mult_82_n2475), 
        .A3(u5_mult_82_n2476), .ZN(u5_mult_82_CARRYB_4__26_) );
  NAND2_X2 u5_mult_82_U6874 ( .A1(u5_mult_82_ab_4__26_), .A2(
        u5_mult_82_CARRYB_3__26_), .ZN(u5_mult_82_n2474) );
  XOR2_X2 u5_mult_82_U6873 ( .A(u5_mult_82_n2473), .B(u5_mult_82_SUMB_4__26_), 
        .Z(u5_mult_82_SUMB_5__25_) );
  XOR2_X2 u5_mult_82_U6872 ( .A(u5_mult_82_ab_5__25_), .B(
        u5_mult_82_CARRYB_4__25_), .Z(u5_mult_82_n2473) );
  NAND3_X2 u5_mult_82_U6871 ( .A1(u5_mult_82_n2472), .A2(u5_mult_82_n2471), 
        .A3(u5_mult_82_n2470), .ZN(u5_mult_82_CARRYB_22__12_) );
  NAND2_X2 u5_mult_82_U6870 ( .A1(u5_mult_82_CARRYB_21__12_), .A2(
        u5_mult_82_SUMB_21__13_), .ZN(u5_mult_82_n2472) );
  NAND2_X2 u5_mult_82_U6869 ( .A1(u5_mult_82_ab_22__12_), .A2(
        u5_mult_82_SUMB_21__13_), .ZN(u5_mult_82_n2471) );
  NAND2_X1 u5_mult_82_U6868 ( .A1(u5_mult_82_CARRYB_20__13_), .A2(
        u5_mult_82_SUMB_20__14_), .ZN(u5_mult_82_n2469) );
  NAND2_X1 u5_mult_82_U6867 ( .A1(u5_mult_82_ab_21__13_), .A2(
        u5_mult_82_CARRYB_20__13_), .ZN(u5_mult_82_n2467) );
  NAND3_X2 u5_mult_82_U6866 ( .A1(u5_mult_82_n2464), .A2(u5_mult_82_n2465), 
        .A3(u5_mult_82_n2466), .ZN(u5_mult_82_CARRYB_20__14_) );
  NAND2_X2 u5_mult_82_U6865 ( .A1(u5_mult_82_ab_20__14_), .A2(
        u5_mult_82_CARRYB_19__14_), .ZN(u5_mult_82_n2466) );
  NAND2_X2 u5_mult_82_U6864 ( .A1(u5_mult_82_ab_20__14_), .A2(
        u5_mult_82_SUMB_19__15_), .ZN(u5_mult_82_n2465) );
  NAND2_X2 u5_mult_82_U6863 ( .A1(u5_mult_82_CARRYB_19__14_), .A2(
        u5_mult_82_SUMB_19__15_), .ZN(u5_mult_82_n2464) );
  NAND3_X4 u5_mult_82_U6862 ( .A1(u5_mult_82_n3677), .A2(u5_mult_82_n3676), 
        .A3(u5_mult_82_n3675), .ZN(u5_mult_82_CARRYB_36__32_) );
  NOR2_X1 u5_mult_82_U6861 ( .A1(u5_mult_82_n6792), .A2(u5_mult_82_n6615), 
        .ZN(u5_mult_82_ab_19__46_) );
  NAND3_X2 u5_mult_82_U6860 ( .A1(u5_mult_82_n2461), .A2(u5_mult_82_n2462), 
        .A3(u5_mult_82_n2463), .ZN(u5_mult_82_CARRYB_31__39_) );
  NAND2_X1 u5_mult_82_U6859 ( .A1(u5_mult_82_SUMB_30__40_), .A2(
        u5_mult_82_CARRYB_30__39_), .ZN(u5_mult_82_n2463) );
  NAND2_X2 u5_mult_82_U6858 ( .A1(u5_mult_82_ab_31__39_), .A2(
        u5_mult_82_CARRYB_30__39_), .ZN(u5_mult_82_n2462) );
  NAND2_X1 u5_mult_82_U6857 ( .A1(u5_mult_82_ab_31__39_), .A2(
        u5_mult_82_SUMB_30__40_), .ZN(u5_mult_82_n2461) );
  NAND3_X2 u5_mult_82_U6856 ( .A1(u5_mult_82_n2458), .A2(u5_mult_82_n2459), 
        .A3(u5_mult_82_n2460), .ZN(u5_mult_82_CARRYB_30__39_) );
  NAND2_X1 u5_mult_82_U6855 ( .A1(u5_mult_82_CARRYB_29__39_), .A2(
        u5_mult_82_SUMB_29__40_), .ZN(u5_mult_82_n2460) );
  NAND2_X2 u5_mult_82_U6854 ( .A1(u5_mult_82_ab_30__39_), .A2(
        u5_mult_82_SUMB_29__40_), .ZN(u5_mult_82_n2459) );
  NAND2_X1 u5_mult_82_U6853 ( .A1(u5_mult_82_ab_30__39_), .A2(
        u5_mult_82_CARRYB_29__39_), .ZN(u5_mult_82_n2458) );
  XOR2_X2 u5_mult_82_U6852 ( .A(u5_mult_82_n2457), .B(u5_mult_82_SUMB_29__40_), 
        .Z(u5_mult_82_SUMB_30__39_) );
  NAND3_X2 u5_mult_82_U6851 ( .A1(u5_mult_82_n2454), .A2(u5_mult_82_n2455), 
        .A3(u5_mult_82_n2456), .ZN(u5_mult_82_CARRYB_19__46_) );
  NAND2_X1 u5_mult_82_U6850 ( .A1(u5_mult_82_ab_19__46_), .A2(
        u5_mult_82_SUMB_18__47_), .ZN(u5_mult_82_n2456) );
  NAND2_X1 u5_mult_82_U6849 ( .A1(u5_mult_82_SUMB_18__47_), .A2(
        u5_mult_82_CARRYB_18__46_), .ZN(u5_mult_82_n2454) );
  XOR2_X2 u5_mult_82_U6848 ( .A(u5_mult_82_CARRYB_18__46_), .B(
        u5_mult_82_n2453), .Z(u5_mult_82_SUMB_19__46_) );
  XOR2_X2 u5_mult_82_U6847 ( .A(u5_mult_82_SUMB_18__47_), .B(
        u5_mult_82_ab_19__46_), .Z(u5_mult_82_n2453) );
  NAND3_X2 u5_mult_82_U6846 ( .A1(u5_mult_82_n2450), .A2(u5_mult_82_n2451), 
        .A3(u5_mult_82_n2452), .ZN(u5_mult_82_CARRYB_29__40_) );
  NAND2_X1 u5_mult_82_U6845 ( .A1(u5_mult_82_CARRYB_28__40_), .A2(
        u5_mult_82_SUMB_28__41_), .ZN(u5_mult_82_n2452) );
  NAND2_X1 u5_mult_82_U6844 ( .A1(u5_mult_82_ab_29__40_), .A2(
        u5_mult_82_SUMB_28__41_), .ZN(u5_mult_82_n2451) );
  NAND3_X2 u5_mult_82_U6843 ( .A1(u5_mult_82_n2447), .A2(u5_mult_82_n2448), 
        .A3(u5_mult_82_n2449), .ZN(u5_mult_82_CARRYB_28__41_) );
  NAND2_X2 u5_mult_82_U6842 ( .A1(u5_mult_82_ab_28__41_), .A2(
        u5_mult_82_SUMB_27__42_), .ZN(u5_mult_82_n2448) );
  XOR2_X2 u5_mult_82_U6841 ( .A(u5_mult_82_n2446), .B(u5_mult_82_SUMB_28__41_), 
        .Z(u5_mult_82_SUMB_29__40_) );
  XOR2_X2 u5_mult_82_U6840 ( .A(u5_mult_82_ab_29__40_), .B(
        u5_mult_82_CARRYB_28__40_), .Z(u5_mult_82_n2446) );
  XOR2_X2 u5_mult_82_U6839 ( .A(u5_mult_82_n2445), .B(u5_mult_82_n1836), .Z(
        u5_mult_82_SUMB_28__41_) );
  XOR2_X2 u5_mult_82_U6838 ( .A(u5_mult_82_CARRYB_27__41_), .B(
        u5_mult_82_ab_28__41_), .Z(u5_mult_82_n2445) );
  NAND2_X2 u5_mult_82_U6837 ( .A1(u5_mult_82_CARRYB_46__29_), .A2(
        u5_mult_82_SUMB_46__30_), .ZN(u5_mult_82_n2444) );
  NAND2_X2 u5_mult_82_U6836 ( .A1(u5_mult_82_ab_47__29_), .A2(
        u5_mult_82_SUMB_46__30_), .ZN(u5_mult_82_n2443) );
  NAND2_X1 u5_mult_82_U6835 ( .A1(u5_mult_82_ab_47__29_), .A2(
        u5_mult_82_CARRYB_46__29_), .ZN(u5_mult_82_n2442) );
  NAND3_X2 u5_mult_82_U6834 ( .A1(u5_mult_82_n2441), .A2(u5_mult_82_n2440), 
        .A3(u5_mult_82_n2439), .ZN(u5_mult_82_CARRYB_46__30_) );
  NAND2_X1 u5_mult_82_U6833 ( .A1(u5_mult_82_CARRYB_45__30_), .A2(
        u5_mult_82_SUMB_45__31_), .ZN(u5_mult_82_n2441) );
  NAND2_X1 u5_mult_82_U6832 ( .A1(u5_mult_82_ab_46__30_), .A2(
        u5_mult_82_SUMB_45__31_), .ZN(u5_mult_82_n2440) );
  NAND2_X1 u5_mult_82_U6831 ( .A1(u5_mult_82_ab_46__30_), .A2(
        u5_mult_82_CARRYB_45__30_), .ZN(u5_mult_82_n2439) );
  XOR2_X2 u5_mult_82_U6830 ( .A(u5_mult_82_n2437), .B(u5_mult_82_SUMB_45__31_), 
        .Z(u5_mult_82_SUMB_46__30_) );
  XOR2_X2 u5_mult_82_U6829 ( .A(u5_mult_82_ab_46__30_), .B(
        u5_mult_82_CARRYB_45__30_), .Z(u5_mult_82_n2437) );
  NAND2_X2 u5_mult_82_U6828 ( .A1(u5_mult_82_ab_5__47_), .A2(
        u5_mult_82_CARRYB_4__47_), .ZN(u5_mult_82_n6195) );
  NOR2_X2 u5_mult_82_U6827 ( .A1(u5_mult_82_n6786), .A2(u5_mult_82_n6520), 
        .ZN(u5_mult_82_ab_4__47_) );
  NAND3_X2 u5_mult_82_U6826 ( .A1(u5_mult_82_n2434), .A2(u5_mult_82_n2435), 
        .A3(u5_mult_82_n2436), .ZN(u5_mult_82_CARRYB_19__37_) );
  NAND2_X2 u5_mult_82_U6825 ( .A1(u5_mult_82_CARRYB_18__37_), .A2(
        u5_mult_82_SUMB_18__38_), .ZN(u5_mult_82_n2436) );
  NAND2_X2 u5_mult_82_U6824 ( .A1(u5_mult_82_ab_19__37_), .A2(
        u5_mult_82_SUMB_18__38_), .ZN(u5_mult_82_n2435) );
  NAND2_X1 u5_mult_82_U6823 ( .A1(u5_mult_82_ab_19__37_), .A2(
        u5_mult_82_CARRYB_18__37_), .ZN(u5_mult_82_n2434) );
  NAND3_X4 u5_mult_82_U6822 ( .A1(u5_mult_82_n2431), .A2(u5_mult_82_n2432), 
        .A3(u5_mult_82_n2433), .ZN(u5_mult_82_CARRYB_18__38_) );
  NAND2_X2 u5_mult_82_U6821 ( .A1(u5_mult_82_CARRYB_17__38_), .A2(
        u5_mult_82_n1512), .ZN(u5_mult_82_n2433) );
  NAND2_X2 u5_mult_82_U6820 ( .A1(u5_mult_82_ab_18__38_), .A2(u5_mult_82_n1512), .ZN(u5_mult_82_n2432) );
  NAND2_X1 u5_mult_82_U6819 ( .A1(u5_mult_82_ab_18__38_), .A2(
        u5_mult_82_CARRYB_17__38_), .ZN(u5_mult_82_n2431) );
  XOR2_X2 u5_mult_82_U6818 ( .A(u5_mult_82_n2430), .B(u5_mult_82_SUMB_18__38_), 
        .Z(u5_mult_82_SUMB_19__37_) );
  XOR2_X2 u5_mult_82_U6817 ( .A(u5_mult_82_ab_19__37_), .B(
        u5_mult_82_CARRYB_18__37_), .Z(u5_mult_82_n2430) );
  NAND2_X1 u5_mult_82_U6816 ( .A1(u5_mult_82_ab_29__32_), .A2(
        u5_mult_82_CARRYB_28__32_), .ZN(u5_mult_82_n2427) );
  NAND3_X4 u5_mult_82_U6815 ( .A1(u5_mult_82_n2424), .A2(u5_mult_82_n2425), 
        .A3(u5_mult_82_n2426), .ZN(u5_mult_82_CARRYB_28__33_) );
  NAND2_X2 u5_mult_82_U6814 ( .A1(u5_mult_82_ab_28__33_), .A2(
        u5_mult_82_SUMB_27__34_), .ZN(u5_mult_82_n2425) );
  NAND2_X1 u5_mult_82_U6813 ( .A1(u5_mult_82_ab_28__33_), .A2(u5_mult_82_n1614), .ZN(u5_mult_82_n2424) );
  XOR2_X2 u5_mult_82_U6812 ( .A(u5_mult_82_n2423), .B(u5_mult_82_SUMB_28__33_), 
        .Z(u5_mult_82_SUMB_29__32_) );
  NAND3_X4 u5_mult_82_U6811 ( .A1(u5_mult_82_n2420), .A2(u5_mult_82_n2421), 
        .A3(u5_mult_82_n2422), .ZN(u5_mult_82_CARRYB_4__47_) );
  NAND2_X1 u5_mult_82_U6810 ( .A1(u5_mult_82_ab_4__47_), .A2(
        u5_mult_82_CARRYB_3__47_), .ZN(u5_mult_82_n2422) );
  XOR2_X2 u5_mult_82_U6809 ( .A(u5_mult_82_CARRYB_3__47_), .B(
        u5_mult_82_ab_4__47_), .Z(u5_mult_82_n2419) );
  NAND3_X4 u5_mult_82_U6808 ( .A1(u5_mult_82_n3684), .A2(u5_mult_82_n3685), 
        .A3(u5_mult_82_n3686), .ZN(u5_mult_82_CARRYB_39__30_) );
  XNOR2_X2 u5_mult_82_U6807 ( .A(u5_mult_82_CARRYB_22__9_), .B(
        u5_mult_82_ab_23__9_), .ZN(u5_mult_82_n2417) );
  NAND2_X2 u5_mult_82_U6806 ( .A1(u5_mult_82_ab_42__10_), .A2(
        u5_mult_82_SUMB_41__11_), .ZN(u5_mult_82_n6163) );
  NOR2_X1 u5_mult_82_U6805 ( .A1(u5_mult_82_n6977), .A2(u5_mult_82_n6820), 
        .ZN(u5_mult_82_ab_52__41_) );
  NOR2_X1 u5_mult_82_U6804 ( .A1(u5_mult_82_n6820), .A2(u5_mult_82_net65193), 
        .ZN(u5_mult_82_ab_51__41_) );
  NOR2_X1 u5_mult_82_U6803 ( .A1(u5_mult_82_n6820), .A2(u5_mult_82_net65223), 
        .ZN(u5_mult_82_ab_50__41_) );
  NOR2_X1 u5_mult_82_U6802 ( .A1(u5_mult_82_n6820), .A2(u5_mult_82_n6752), 
        .ZN(u5_mult_82_ab_49__41_) );
  NOR2_X1 u5_mult_82_U6801 ( .A1(u5_mult_82_n6820), .A2(u5_mult_82_n6746), 
        .ZN(u5_mult_82_ab_48__41_) );
  NOR2_X1 u5_mult_82_U6800 ( .A1(u5_mult_82_n6820), .A2(u5_mult_82_net65277), 
        .ZN(u5_mult_82_ab_47__41_) );
  NOR2_X1 u5_mult_82_U6799 ( .A1(u5_mult_82_n6820), .A2(u5_mult_82_n6742), 
        .ZN(u5_mult_82_ab_46__41_) );
  NOR2_X1 u5_mult_82_U6798 ( .A1(u5_mult_82_n6820), .A2(u5_mult_82_net65313), 
        .ZN(u5_mult_82_ab_45__41_) );
  NOR2_X1 u5_mult_82_U6797 ( .A1(u5_mult_82_n6820), .A2(u5_mult_82_n6735), 
        .ZN(u5_mult_82_ab_44__41_) );
  NOR2_X1 u5_mult_82_U6796 ( .A1(u5_mult_82_n6820), .A2(u5_mult_82_net65349), 
        .ZN(u5_mult_82_ab_43__41_) );
  NOR2_X1 u5_mult_82_U6795 ( .A1(u5_mult_82_n6820), .A2(u5_mult_82_net65371), 
        .ZN(u5_mult_82_ab_42__41_) );
  NAND2_X2 u5_mult_82_U6794 ( .A1(u5_mult_82_n1711), .A2(
        u5_mult_82_SUMB_16__48_), .ZN(u5_mult_82_n5955) );
  NAND2_X2 u5_mult_82_U6793 ( .A1(u5_mult_82_SUMB_43__5_), .A2(
        u5_mult_82_CARRYB_43__4_), .ZN(u5_mult_82_n5790) );
  NAND2_X2 u5_mult_82_U6792 ( .A1(u5_mult_82_n1625), .A2(u5_mult_82_n1642), 
        .ZN(u5_mult_82_n3209) );
  XNOR2_X2 u5_mult_82_U6791 ( .A(u5_mult_82_n2415), .B(
        u5_mult_82_CARRYB_12__38_), .ZN(u5_mult_82_n6155) );
  NAND2_X2 u5_mult_82_U6790 ( .A1(u5_mult_82_CARRYB_31__26_), .A2(
        u5_mult_82_n1500), .ZN(u5_mult_82_n3956) );
  NAND2_X2 u5_mult_82_U6789 ( .A1(u5_mult_82_CARRYB_29__29_), .A2(
        u5_mult_82_SUMB_29__30_), .ZN(u5_mult_82_n4539) );
  NAND3_X2 u5_mult_82_U6788 ( .A1(u5_mult_82_n4076), .A2(u5_mult_82_n4077), 
        .A3(u5_mult_82_n4078), .ZN(u5_mult_82_CARRYB_36__8_) );
  NAND2_X2 u5_mult_82_U6787 ( .A1(u5_mult_82_SUMB_43__5_), .A2(
        u5_mult_82_ab_44__4_), .ZN(u5_mult_82_n5789) );
  XOR2_X1 u5_mult_82_U6786 ( .A(u5_mult_82_n2644), .B(u5_mult_82_n1660), .Z(
        u5_mult_82_SUMB_11__15_) );
  XNOR2_X2 u5_mult_82_U6785 ( .A(u5_mult_82_n2414), .B(
        u5_mult_82_CARRYB_27__30_), .ZN(u5_mult_82_n3223) );
  NAND3_X4 u5_mult_82_U6784 ( .A1(u5_mult_82_n5936), .A2(u5_mult_82_n5937), 
        .A3(u5_mult_82_n5938), .ZN(u5_mult_82_CARRYB_49__15_) );
  XNOR2_X2 u5_mult_82_U6783 ( .A(u5_mult_82_ab_23__34_), .B(u5_mult_82_n5506), 
        .ZN(u5_mult_82_n6371) );
  INV_X16 u5_mult_82_U6782 ( .A(n4760), .ZN(u5_mult_82_n7019) );
  NAND3_X4 u5_mult_82_U6781 ( .A1(u5_mult_82_n3724), .A2(u5_mult_82_n3725), 
        .A3(u5_mult_82_n3726), .ZN(u5_mult_82_CARRYB_21__9_) );
  XNOR2_X2 u5_mult_82_U6780 ( .A(u5_mult_82_CARRYB_44__17_), .B(
        u5_mult_82_n2412), .ZN(u5_mult_82_SUMB_45__17_) );
  XNOR2_X2 u5_mult_82_U6779 ( .A(u5_mult_82_ab_41__8_), .B(
        u5_mult_82_CARRYB_40__8_), .ZN(u5_mult_82_n2411) );
  XNOR2_X2 u5_mult_82_U6778 ( .A(u5_mult_82_n2411), .B(u5_mult_82_SUMB_40__9_), 
        .ZN(u5_mult_82_SUMB_41__8_) );
  NAND3_X2 u5_mult_82_U6777 ( .A1(u5_mult_82_n5896), .A2(u5_mult_82_n5897), 
        .A3(u5_mult_82_n5898), .ZN(u5_mult_82_CARRYB_35__20_) );
  XNOR2_X2 u5_mult_82_U6776 ( .A(u5_mult_82_CARRYB_38__5_), .B(
        u5_mult_82_ab_39__5_), .ZN(u5_mult_82_n2690) );
  XNOR2_X2 u5_mult_82_U6775 ( .A(u5_mult_82_n2410), .B(u5_mult_82_n1387), .ZN(
        u5_mult_82_SUMB_36__22_) );
  XOR2_X2 u5_mult_82_U6774 ( .A(u5_mult_82_n4360), .B(
        u5_mult_82_CARRYB_45__17_), .Z(u5_mult_82_n2409) );
  NAND2_X2 u5_mult_82_U6773 ( .A1(u5_mult_82_n4957), .A2(u5_mult_82_n4958), 
        .ZN(u5_mult_82_n5627) );
  XNOR2_X2 u5_mult_82_U6772 ( .A(u5_mult_82_n2630), .B(u5_mult_82_SUMB_28__14_), .ZN(u5_mult_82_SUMB_29__13_) );
  NAND3_X2 u5_mult_82_U6771 ( .A1(u5_mult_82_n2599), .A2(u5_mult_82_n2600), 
        .A3(u5_mult_82_n2601), .ZN(u5_mult_82_CARRYB_29__12_) );
  NAND2_X2 u5_mult_82_U6770 ( .A1(u5_mult_82_ab_17__47_), .A2(u5_mult_82_n1711), .ZN(u5_mult_82_n5953) );
  XNOR2_X2 u5_mult_82_U6769 ( .A(u5_mult_82_CARRYB_32__18_), .B(
        u5_mult_82_ab_33__18_), .ZN(u5_mult_82_n2408) );
  XNOR2_X2 u5_mult_82_U6768 ( .A(u5_mult_82_n2408), .B(u5_mult_82_SUMB_32__19_), .ZN(u5_mult_82_SUMB_33__18_) );
  NAND3_X4 u5_mult_82_U6767 ( .A1(u5_mult_82_n5863), .A2(u5_mult_82_n5862), 
        .A3(u5_mult_82_n5861), .ZN(u5_mult_82_CARRYB_46__17_) );
  NAND2_X1 u5_mult_82_U6766 ( .A1(u5_mult_82_ab_9__42_), .A2(
        u5_mult_82_SUMB_8__43_), .ZN(u5_mult_82_n5000) );
  NAND2_X2 u5_mult_82_U6765 ( .A1(u5_mult_82_ab_20__42_), .A2(
        u5_mult_82_SUMB_19__43_), .ZN(u5_mult_82_n5844) );
  NAND2_X2 u5_mult_82_U6764 ( .A1(u5_mult_82_ab_35__33_), .A2(
        u5_mult_82_SUMB_34__34_), .ZN(u5_mult_82_n3612) );
  NAND2_X2 u5_mult_82_U6763 ( .A1(u5_mult_82_CARRYB_39__30_), .A2(
        u5_mult_82_SUMB_39__31_), .ZN(u5_mult_82_n4919) );
  NAND2_X2 u5_mult_82_U6762 ( .A1(u5_mult_82_ab_39__11_), .A2(
        u5_mult_82_SUMB_38__12_), .ZN(u5_mult_82_n5132) );
  NAND3_X4 u5_mult_82_U6761 ( .A1(u5_mult_82_n4917), .A2(u5_mult_82_n4918), 
        .A3(u5_mult_82_n4919), .ZN(u5_mult_82_CARRYB_40__30_) );
  XNOR2_X2 u5_mult_82_U6760 ( .A(u5_mult_82_ab_6__44_), .B(
        u5_mult_82_CARRYB_5__44_), .ZN(u5_mult_82_n2407) );
  XNOR2_X2 u5_mult_82_U6759 ( .A(u5_mult_82_n2407), .B(u5_mult_82_SUMB_5__45_), 
        .ZN(u5_mult_82_SUMB_6__44_) );
  NAND2_X1 u5_mult_82_U6758 ( .A1(u5_mult_82_CARRYB_50__3_), .A2(
        u5_mult_82_SUMB_50__4_), .ZN(u5_mult_82_n5240) );
  NAND2_X1 u5_mult_82_U6757 ( .A1(u5_mult_82_ab_13__36_), .A2(
        u5_mult_82_CARRYB_12__36_), .ZN(u5_mult_82_n5200) );
  XNOR2_X2 u5_mult_82_U6756 ( .A(u5_mult_82_SUMB_28__48_), .B(
        u5_mult_82_ab_29__47_), .ZN(u5_mult_82_n2406) );
  XNOR2_X2 u5_mult_82_U6755 ( .A(u5_mult_82_CARRYB_28__47_), .B(
        u5_mult_82_n2406), .ZN(u5_mult_82_SUMB_29__47_) );
  XNOR2_X2 u5_mult_82_U6754 ( .A(u5_mult_82_ab_51__26_), .B(
        u5_mult_82_CARRYB_50__26_), .ZN(u5_mult_82_n2405) );
  XNOR2_X2 u5_mult_82_U6753 ( .A(u5_mult_82_n2405), .B(u5_mult_82_SUMB_50__27_), .ZN(u5_mult_82_SUMB_51__26_) );
  NAND2_X2 u5_mult_82_U6752 ( .A1(u5_mult_82_SUMB_20__10_), .A2(
        u5_mult_82_CARRYB_20__9_), .ZN(u5_mult_82_n3724) );
  NAND3_X2 u5_mult_82_U6751 ( .A1(u5_mult_82_n2402), .A2(u5_mult_82_n2403), 
        .A3(u5_mult_82_n2404), .ZN(u5_mult_82_CARRYB_30__38_) );
  NAND2_X1 u5_mult_82_U6750 ( .A1(u5_mult_82_CARRYB_29__38_), .A2(
        u5_mult_82_SUMB_29__39_), .ZN(u5_mult_82_n2404) );
  NAND2_X1 u5_mult_82_U6749 ( .A1(u5_mult_82_ab_30__38_), .A2(
        u5_mult_82_SUMB_29__39_), .ZN(u5_mult_82_n2403) );
  NAND3_X4 u5_mult_82_U6748 ( .A1(u5_mult_82_n2399), .A2(u5_mult_82_n2400), 
        .A3(u5_mult_82_n2401), .ZN(u5_mult_82_CARRYB_29__39_) );
  NAND2_X2 u5_mult_82_U6747 ( .A1(u5_mult_82_n1810), .A2(
        u5_mult_82_CARRYB_28__39_), .ZN(u5_mult_82_n2401) );
  NAND2_X2 u5_mult_82_U6746 ( .A1(u5_mult_82_ab_29__39_), .A2(
        u5_mult_82_CARRYB_28__39_), .ZN(u5_mult_82_n2399) );
  XOR2_X2 u5_mult_82_U6745 ( .A(u5_mult_82_n2398), .B(u5_mult_82_n1810), .Z(
        u5_mult_82_SUMB_29__39_) );
  XOR2_X2 u5_mult_82_U6744 ( .A(u5_mult_82_ab_29__39_), .B(
        u5_mult_82_CARRYB_28__39_), .Z(u5_mult_82_n2398) );
  XNOR2_X2 u5_mult_82_U6743 ( .A(u5_mult_82_ab_15__24_), .B(
        u5_mult_82_CARRYB_14__24_), .ZN(u5_mult_82_n2397) );
  XNOR2_X2 u5_mult_82_U6742 ( .A(u5_mult_82_n2397), .B(u5_mult_82_SUMB_14__25_), .ZN(u5_mult_82_SUMB_15__24_) );
  NAND2_X2 u5_mult_82_U6741 ( .A1(u5_mult_82_CARRYB_49__35_), .A2(
        u5_mult_82_SUMB_49__36_), .ZN(u5_mult_82_n2695) );
  NAND2_X2 u5_mult_82_U6740 ( .A1(u5_mult_82_ab_50__35_), .A2(
        u5_mult_82_CARRYB_49__35_), .ZN(u5_mult_82_n2693) );
  NAND3_X4 u5_mult_82_U6739 ( .A1(u5_mult_82_n3091), .A2(u5_mult_82_n3092), 
        .A3(u5_mult_82_n3093), .ZN(u5_mult_82_CARRYB_48__35_) );
  NOR2_X1 u5_mult_82_U6738 ( .A1(u5_mult_82_net64913), .A2(u5_mult_82_n6753), 
        .ZN(u5_mult_82_ab_49__35_) );
  NAND3_X2 u5_mult_82_U6737 ( .A1(u5_mult_82_n2394), .A2(u5_mult_82_n2395), 
        .A3(u5_mult_82_n2396), .ZN(u5_mult_82_CARRYB_43__40_) );
  NAND2_X1 u5_mult_82_U6736 ( .A1(u5_mult_82_CARRYB_42__40_), .A2(
        u5_mult_82_SUMB_42__41_), .ZN(u5_mult_82_n2396) );
  NAND2_X1 u5_mult_82_U6735 ( .A1(u5_mult_82_ab_43__40_), .A2(
        u5_mult_82_SUMB_42__41_), .ZN(u5_mult_82_n2395) );
  NAND2_X1 u5_mult_82_U6734 ( .A1(u5_mult_82_ab_43__40_), .A2(
        u5_mult_82_CARRYB_42__40_), .ZN(u5_mult_82_n2394) );
  NAND3_X2 u5_mult_82_U6733 ( .A1(u5_mult_82_n2391), .A2(u5_mult_82_n2392), 
        .A3(u5_mult_82_n2393), .ZN(u5_mult_82_CARRYB_42__41_) );
  NAND2_X2 u5_mult_82_U6732 ( .A1(u5_mult_82_CARRYB_41__41_), .A2(
        u5_mult_82_SUMB_41__42_), .ZN(u5_mult_82_n2393) );
  NAND2_X2 u5_mult_82_U6731 ( .A1(u5_mult_82_ab_42__41_), .A2(
        u5_mult_82_SUMB_41__42_), .ZN(u5_mult_82_n2392) );
  NAND2_X1 u5_mult_82_U6730 ( .A1(u5_mult_82_ab_42__41_), .A2(
        u5_mult_82_CARRYB_41__41_), .ZN(u5_mult_82_n2391) );
  XOR2_X2 u5_mult_82_U6729 ( .A(u5_mult_82_n2390), .B(u5_mult_82_SUMB_42__41_), 
        .Z(u5_mult_82_SUMB_43__40_) );
  XOR2_X2 u5_mult_82_U6728 ( .A(u5_mult_82_ab_43__40_), .B(
        u5_mult_82_CARRYB_42__40_), .Z(u5_mult_82_n2390) );
  XOR2_X2 u5_mult_82_U6727 ( .A(u5_mult_82_n2389), .B(u5_mult_82_SUMB_41__42_), 
        .Z(u5_mult_82_SUMB_42__41_) );
  XOR2_X2 u5_mult_82_U6726 ( .A(u5_mult_82_CARRYB_41__41_), .B(
        u5_mult_82_ab_42__41_), .Z(u5_mult_82_n2389) );
  NAND3_X2 u5_mult_82_U6725 ( .A1(u5_mult_82_n2386), .A2(u5_mult_82_n2387), 
        .A3(u5_mult_82_n2388), .ZN(u5_mult_82_CARRYB_24__47_) );
  NAND2_X1 u5_mult_82_U6724 ( .A1(u5_mult_82_CARRYB_23__47_), .A2(
        u5_mult_82_SUMB_23__48_), .ZN(u5_mult_82_n2388) );
  NAND2_X1 u5_mult_82_U6723 ( .A1(u5_mult_82_ab_24__47_), .A2(
        u5_mult_82_SUMB_23__48_), .ZN(u5_mult_82_n2387) );
  NAND2_X1 u5_mult_82_U6722 ( .A1(u5_mult_82_ab_24__47_), .A2(
        u5_mult_82_CARRYB_23__47_), .ZN(u5_mult_82_n2386) );
  NAND3_X2 u5_mult_82_U6721 ( .A1(u5_mult_82_n2383), .A2(u5_mult_82_n2384), 
        .A3(u5_mult_82_n2385), .ZN(u5_mult_82_CARRYB_23__48_) );
  NAND2_X1 u5_mult_82_U6720 ( .A1(u5_mult_82_CARRYB_22__48_), .A2(
        u5_mult_82_SUMB_22__49_), .ZN(u5_mult_82_n2385) );
  NAND2_X1 u5_mult_82_U6719 ( .A1(u5_mult_82_ab_23__48_), .A2(
        u5_mult_82_SUMB_22__49_), .ZN(u5_mult_82_n2384) );
  NAND2_X1 u5_mult_82_U6718 ( .A1(u5_mult_82_ab_23__48_), .A2(
        u5_mult_82_CARRYB_22__48_), .ZN(u5_mult_82_n2383) );
  XOR2_X2 u5_mult_82_U6717 ( .A(u5_mult_82_n2382), .B(u5_mult_82_SUMB_23__48_), 
        .Z(u5_mult_82_SUMB_24__47_) );
  XOR2_X2 u5_mult_82_U6716 ( .A(u5_mult_82_n2381), .B(u5_mult_82_SUMB_22__49_), 
        .Z(u5_mult_82_SUMB_23__48_) );
  XOR2_X2 u5_mult_82_U6715 ( .A(u5_mult_82_CARRYB_22__48_), .B(
        u5_mult_82_ab_23__48_), .Z(u5_mult_82_n2381) );
  NAND3_X2 u5_mult_82_U6714 ( .A1(u5_mult_82_n2378), .A2(u5_mult_82_n2379), 
        .A3(u5_mult_82_n2380), .ZN(u5_mult_82_CARRYB_36__44_) );
  NAND2_X1 u5_mult_82_U6713 ( .A1(u5_mult_82_ab_36__44_), .A2(
        u5_mult_82_SUMB_35__45_), .ZN(u5_mult_82_n2380) );
  NAND2_X1 u5_mult_82_U6712 ( .A1(u5_mult_82_CARRYB_35__44_), .A2(
        u5_mult_82_SUMB_35__45_), .ZN(u5_mult_82_n2379) );
  NAND2_X1 u5_mult_82_U6711 ( .A1(u5_mult_82_CARRYB_35__44_), .A2(
        u5_mult_82_ab_36__44_), .ZN(u5_mult_82_n2378) );
  NAND3_X2 u5_mult_82_U6710 ( .A1(u5_mult_82_n2375), .A2(u5_mult_82_n2376), 
        .A3(u5_mult_82_n2377), .ZN(u5_mult_82_CARRYB_35__45_) );
  NAND2_X2 u5_mult_82_U6709 ( .A1(u5_mult_82_CARRYB_34__45_), .A2(
        u5_mult_82_SUMB_34__46_), .ZN(u5_mult_82_n2377) );
  NAND2_X2 u5_mult_82_U6708 ( .A1(u5_mult_82_ab_35__45_), .A2(
        u5_mult_82_SUMB_34__46_), .ZN(u5_mult_82_n2376) );
  NAND2_X1 u5_mult_82_U6707 ( .A1(u5_mult_82_ab_35__45_), .A2(
        u5_mult_82_CARRYB_34__45_), .ZN(u5_mult_82_n2375) );
  XOR2_X2 u5_mult_82_U6706 ( .A(u5_mult_82_n2374), .B(u5_mult_82_SUMB_35__45_), 
        .Z(u5_mult_82_SUMB_36__44_) );
  XOR2_X2 u5_mult_82_U6705 ( .A(u5_mult_82_CARRYB_35__44_), .B(
        u5_mult_82_ab_36__44_), .Z(u5_mult_82_n2374) );
  XOR2_X2 u5_mult_82_U6704 ( .A(u5_mult_82_n2373), .B(u5_mult_82_SUMB_34__46_), 
        .Z(u5_mult_82_SUMB_35__45_) );
  XOR2_X2 u5_mult_82_U6703 ( .A(u5_mult_82_ab_35__45_), .B(
        u5_mult_82_CARRYB_34__45_), .Z(u5_mult_82_n2373) );
  NAND3_X2 u5_mult_82_U6702 ( .A1(u5_mult_82_n2370), .A2(u5_mult_82_n2371), 
        .A3(u5_mult_82_n2372), .ZN(u5_mult_82_CARRYB_52__32_) );
  NAND2_X1 u5_mult_82_U6701 ( .A1(u5_mult_82_CARRYB_51__32_), .A2(
        u5_mult_82_SUMB_51__33_), .ZN(u5_mult_82_n2372) );
  NAND2_X1 u5_mult_82_U6700 ( .A1(u5_mult_82_ab_52__32_), .A2(
        u5_mult_82_SUMB_51__33_), .ZN(u5_mult_82_n2371) );
  NAND2_X1 u5_mult_82_U6699 ( .A1(u5_mult_82_ab_52__32_), .A2(
        u5_mult_82_CARRYB_51__32_), .ZN(u5_mult_82_n2370) );
  NAND3_X2 u5_mult_82_U6698 ( .A1(u5_mult_82_n2367), .A2(u5_mult_82_n2368), 
        .A3(u5_mult_82_n2369), .ZN(u5_mult_82_CARRYB_51__33_) );
  NAND2_X1 u5_mult_82_U6697 ( .A1(u5_mult_82_CARRYB_50__33_), .A2(
        u5_mult_82_SUMB_50__34_), .ZN(u5_mult_82_n2369) );
  NAND2_X1 u5_mult_82_U6696 ( .A1(u5_mult_82_ab_51__33_), .A2(
        u5_mult_82_SUMB_50__34_), .ZN(u5_mult_82_n2368) );
  NAND2_X1 u5_mult_82_U6695 ( .A1(u5_mult_82_ab_51__33_), .A2(
        u5_mult_82_CARRYB_50__33_), .ZN(u5_mult_82_n2367) );
  XOR2_X2 u5_mult_82_U6694 ( .A(u5_mult_82_n2366), .B(u5_mult_82_n1416), .Z(
        u5_mult_82_SUMB_51__33_) );
  XOR2_X2 u5_mult_82_U6693 ( .A(u5_mult_82_ab_51__33_), .B(
        u5_mult_82_CARRYB_50__33_), .Z(u5_mult_82_n2366) );
  NAND3_X2 u5_mult_82_U6692 ( .A1(u5_mult_82_n2363), .A2(u5_mult_82_n2364), 
        .A3(u5_mult_82_n2365), .ZN(u5_mult_82_CARRYB_49__35_) );
  NAND2_X1 u5_mult_82_U6691 ( .A1(u5_mult_82_ab_49__35_), .A2(
        u5_mult_82_CARRYB_48__35_), .ZN(u5_mult_82_n2365) );
  NAND2_X2 u5_mult_82_U6690 ( .A1(u5_mult_82_ab_49__35_), .A2(
        u5_mult_82_SUMB_48__36_), .ZN(u5_mult_82_n2364) );
  NAND2_X1 u5_mult_82_U6689 ( .A1(u5_mult_82_CARRYB_48__35_), .A2(
        u5_mult_82_SUMB_48__36_), .ZN(u5_mult_82_n2363) );
  XOR2_X2 u5_mult_82_U6688 ( .A(u5_mult_82_n7), .B(u5_mult_82_n2362), .Z(
        u5_mult_82_SUMB_49__35_) );
  XOR2_X2 u5_mult_82_U6687 ( .A(u5_mult_82_CARRYB_48__35_), .B(
        u5_mult_82_ab_49__35_), .Z(u5_mult_82_n2362) );
  NAND2_X2 u5_mult_82_U6686 ( .A1(u5_mult_82_ab_36__22_), .A2(u5_mult_82_n718), 
        .ZN(u5_mult_82_n6216) );
  NAND2_X2 u5_mult_82_U6685 ( .A1(u5_mult_82_n2359), .A2(u5_mult_82_n2360), 
        .ZN(u5_mult_82_SUMB_17__35_) );
  NAND2_X1 u5_mult_82_U6684 ( .A1(u5_mult_82_n6186), .A2(u5_mult_82_n2358), 
        .ZN(u5_mult_82_n2359) );
  NAND3_X2 u5_mult_82_U6683 ( .A1(u5_mult_82_n2355), .A2(u5_mult_82_n2356), 
        .A3(u5_mult_82_n2357), .ZN(u5_mult_82_CARRYB_30__27_) );
  NAND2_X1 u5_mult_82_U6682 ( .A1(u5_mult_82_CARRYB_29__27_), .A2(
        u5_mult_82_SUMB_29__28_), .ZN(u5_mult_82_n2357) );
  NAND2_X1 u5_mult_82_U6681 ( .A1(u5_mult_82_ab_30__27_), .A2(
        u5_mult_82_SUMB_29__28_), .ZN(u5_mult_82_n2356) );
  NAND2_X1 u5_mult_82_U6680 ( .A1(u5_mult_82_ab_30__27_), .A2(
        u5_mult_82_CARRYB_29__27_), .ZN(u5_mult_82_n2355) );
  NAND2_X2 u5_mult_82_U6679 ( .A1(u5_mult_82_ab_29__28_), .A2(
        u5_mult_82_SUMB_28__29_), .ZN(u5_mult_82_n2353) );
  NAND2_X1 u5_mult_82_U6678 ( .A1(u5_mult_82_ab_29__28_), .A2(
        u5_mult_82_CARRYB_28__28_), .ZN(u5_mult_82_n2352) );
  XOR2_X2 u5_mult_82_U6677 ( .A(u5_mult_82_n2351), .B(u5_mult_82_SUMB_28__29_), 
        .Z(u5_mult_82_SUMB_29__28_) );
  NAND2_X2 u5_mult_82_U6676 ( .A1(u5_mult_82_n718), .A2(
        u5_mult_82_SUMB_35__23_), .ZN(u5_mult_82_n6218) );
  XNOR2_X2 u5_mult_82_U6675 ( .A(u5_mult_82_ab_30__27_), .B(
        u5_mult_82_CARRYB_29__27_), .ZN(u5_mult_82_n2350) );
  XNOR2_X2 u5_mult_82_U6674 ( .A(u5_mult_82_n2350), .B(u5_mult_82_SUMB_29__28_), .ZN(u5_mult_82_SUMB_30__27_) );
  NAND2_X2 u5_mult_82_U6673 ( .A1(u5_mult_82_CARRYB_41__10_), .A2(
        u5_mult_82_SUMB_41__11_), .ZN(u5_mult_82_n6162) );
  NOR2_X1 u5_mult_82_U6672 ( .A1(u5_mult_82_n6946), .A2(u5_mult_82_n6722), 
        .ZN(u5_mult_82_ab_37__4_) );
  NAND3_X2 u5_mult_82_U6671 ( .A1(u5_mult_82_n2347), .A2(u5_mult_82_n2348), 
        .A3(u5_mult_82_n2349), .ZN(u5_mult_82_CARRYB_34__4_) );
  NAND2_X1 u5_mult_82_U6670 ( .A1(u5_mult_82_SUMB_33__5_), .A2(
        u5_mult_82_CARRYB_33__4_), .ZN(u5_mult_82_n2349) );
  NAND2_X2 u5_mult_82_U6669 ( .A1(u5_mult_82_ab_34__4_), .A2(
        u5_mult_82_CARRYB_33__4_), .ZN(u5_mult_82_n2348) );
  NAND2_X1 u5_mult_82_U6668 ( .A1(u5_mult_82_ab_34__4_), .A2(
        u5_mult_82_SUMB_33__5_), .ZN(u5_mult_82_n2347) );
  XOR2_X2 u5_mult_82_U6667 ( .A(u5_mult_82_n2346), .B(u5_mult_82_CARRYB_33__4_), .Z(u5_mult_82_SUMB_34__4_) );
  XOR2_X2 u5_mult_82_U6666 ( .A(u5_mult_82_ab_34__4_), .B(
        u5_mult_82_SUMB_33__5_), .Z(u5_mult_82_n2346) );
  NAND3_X2 u5_mult_82_U6665 ( .A1(u5_mult_82_n2343), .A2(u5_mult_82_n2344), 
        .A3(u5_mult_82_n2345), .ZN(u5_mult_82_CARRYB_33__4_) );
  NAND2_X1 u5_mult_82_U6664 ( .A1(u5_mult_82_CARRYB_32__4_), .A2(
        u5_mult_82_SUMB_32__5_), .ZN(u5_mult_82_n2345) );
  NAND2_X2 u5_mult_82_U6663 ( .A1(u5_mult_82_ab_33__4_), .A2(
        u5_mult_82_SUMB_32__5_), .ZN(u5_mult_82_n2344) );
  NAND2_X1 u5_mult_82_U6662 ( .A1(u5_mult_82_ab_33__4_), .A2(
        u5_mult_82_CARRYB_32__4_), .ZN(u5_mult_82_n2343) );
  NAND3_X2 u5_mult_82_U6661 ( .A1(u5_mult_82_n2340), .A2(u5_mult_82_n2341), 
        .A3(u5_mult_82_n2342), .ZN(u5_mult_82_CARRYB_37__4_) );
  NAND2_X2 u5_mult_82_U6660 ( .A1(u5_mult_82_ab_37__4_), .A2(
        u5_mult_82_CARRYB_36__4_), .ZN(u5_mult_82_n2341) );
  XOR2_X2 u5_mult_82_U6659 ( .A(u5_mult_82_CARRYB_36__4_), .B(u5_mult_82_n2339), .Z(u5_mult_82_SUMB_37__4_) );
  XOR2_X2 u5_mult_82_U6658 ( .A(u5_mult_82_n390), .B(u5_mult_82_ab_37__4_), 
        .Z(u5_mult_82_n2339) );
  NAND3_X2 u5_mult_82_U6657 ( .A1(u5_mult_82_n2336), .A2(u5_mult_82_n2337), 
        .A3(u5_mult_82_n2338), .ZN(u5_mult_82_CARRYB_13__11_) );
  NAND2_X1 u5_mult_82_U6656 ( .A1(u5_mult_82_CARRYB_12__11_), .A2(
        u5_mult_82_SUMB_12__12_), .ZN(u5_mult_82_n2338) );
  NAND2_X1 u5_mult_82_U6655 ( .A1(u5_mult_82_ab_13__11_), .A2(
        u5_mult_82_SUMB_12__12_), .ZN(u5_mult_82_n2337) );
  NAND2_X1 u5_mult_82_U6654 ( .A1(u5_mult_82_ab_13__11_), .A2(
        u5_mult_82_CARRYB_12__11_), .ZN(u5_mult_82_n2336) );
  NAND3_X2 u5_mult_82_U6653 ( .A1(u5_mult_82_n2333), .A2(u5_mult_82_n2334), 
        .A3(u5_mult_82_n2335), .ZN(u5_mult_82_CARRYB_12__12_) );
  NAND2_X2 u5_mult_82_U6652 ( .A1(u5_mult_82_CARRYB_11__12_), .A2(
        u5_mult_82_SUMB_11__13_), .ZN(u5_mult_82_n2335) );
  NAND2_X2 u5_mult_82_U6651 ( .A1(u5_mult_82_ab_12__12_), .A2(
        u5_mult_82_SUMB_11__13_), .ZN(u5_mult_82_n2334) );
  NAND2_X1 u5_mult_82_U6650 ( .A1(u5_mult_82_ab_12__12_), .A2(
        u5_mult_82_CARRYB_11__12_), .ZN(u5_mult_82_n2333) );
  XOR2_X2 u5_mult_82_U6649 ( .A(u5_mult_82_n2332), .B(u5_mult_82_SUMB_12__12_), 
        .Z(u5_mult_82_SUMB_13__11_) );
  XOR2_X2 u5_mult_82_U6648 ( .A(u5_mult_82_ab_13__11_), .B(
        u5_mult_82_CARRYB_12__11_), .Z(u5_mult_82_n2332) );
  XOR2_X2 u5_mult_82_U6647 ( .A(u5_mult_82_n2331), .B(u5_mult_82_SUMB_11__13_), 
        .Z(u5_mult_82_SUMB_12__12_) );
  XOR2_X2 u5_mult_82_U6646 ( .A(u5_mult_82_ab_12__12_), .B(
        u5_mult_82_CARRYB_11__12_), .Z(u5_mult_82_n2331) );
  XNOR2_X2 u5_mult_82_U6645 ( .A(u5_mult_82_ab_46__26_), .B(
        u5_mult_82_CARRYB_45__26_), .ZN(u5_mult_82_n2330) );
  INV_X2 u5_mult_82_U6644 ( .A(u5_mult_82_n5550), .ZN(u5_mult_82_n5252) );
  NAND2_X1 u5_mult_82_U6643 ( .A1(u5_mult_82_n1422), .A2(
        u5_mult_82_SUMB_17__47_), .ZN(u5_mult_82_n5958) );
  NAND2_X1 u5_mult_82_U6642 ( .A1(u5_mult_82_ab_18__46_), .A2(u5_mult_82_n1422), .ZN(u5_mult_82_n5956) );
  XOR2_X2 u5_mult_82_U6641 ( .A(u5_mult_82_n4449), .B(u5_mult_82_SUMB_39__35_), 
        .Z(u5_mult_82_SUMB_40__34_) );
  NAND2_X2 u5_mult_82_U6640 ( .A1(u5_mult_82_ab_20__24_), .A2(
        u5_mult_82_SUMB_19__25_), .ZN(u5_mult_82_n5612) );
  NAND3_X4 u5_mult_82_U6639 ( .A1(u5_mult_82_n4445), .A2(u5_mult_82_n4446), 
        .A3(u5_mult_82_n4447), .ZN(u5_mult_82_CARRYB_50__24_) );
  XNOR2_X2 u5_mult_82_U6638 ( .A(u5_mult_82_n2329), .B(
        u5_mult_82_CARRYB_45__18_), .ZN(u5_mult_82_n5344) );
  XNOR2_X2 u5_mult_82_U6637 ( .A(u5_mult_82_CARRYB_36__5_), .B(
        u5_mult_82_ab_37__5_), .ZN(u5_mult_82_n2328) );
  XNOR2_X2 u5_mult_82_U6636 ( .A(u5_mult_82_n2328), .B(u5_mult_82_SUMB_36__6_), 
        .ZN(u5_mult_82_SUMB_37__5_) );
  NAND2_X2 u5_mult_82_U6635 ( .A1(u5_mult_82_CARRYB_30__36_), .A2(
        u5_mult_82_SUMB_30__37_), .ZN(u5_mult_82_n4321) );
  NAND3_X4 u5_mult_82_U6634 ( .A1(u5_mult_82_n4645), .A2(u5_mult_82_n4646), 
        .A3(u5_mult_82_n4647), .ZN(u5_mult_82_CARRYB_30__36_) );
  XNOR2_X2 u5_mult_82_U6633 ( .A(u5_mult_82_ab_42__29_), .B(
        u5_mult_82_CARRYB_41__29_), .ZN(u5_mult_82_n2327) );
  XNOR2_X2 u5_mult_82_U6632 ( .A(u5_mult_82_n2327), .B(u5_mult_82_SUMB_41__30_), .ZN(u5_mult_82_SUMB_42__29_) );
  XNOR2_X2 u5_mult_82_U6631 ( .A(u5_mult_82_n2326), .B(u5_mult_82_SUMB_48__30_), .ZN(u5_mult_82_SUMB_49__29_) );
  XNOR2_X2 u5_mult_82_U6630 ( .A(u5_mult_82_n2325), .B(
        u5_mult_82_CARRYB_34__23_), .ZN(u5_mult_82_n6212) );
  NAND2_X2 u5_mult_82_U6629 ( .A1(u5_mult_82_ab_29__36_), .A2(
        u5_mult_82_SUMB_28__37_), .ZN(u5_mult_82_n5668) );
  XNOR2_X2 u5_mult_82_U6628 ( .A(u5_mult_82_CARRYB_32__9_), .B(
        u5_mult_82_n2324), .ZN(u5_mult_82_n4519) );
  NAND2_X1 u5_mult_82_U6627 ( .A1(u5_mult_82_CARRYB_13__45_), .A2(
        u5_mult_82_SUMB_13__46_), .ZN(u5_mult_82_n2724) );
  XNOR2_X2 u5_mult_82_U6626 ( .A(u5_mult_82_ab_28__39_), .B(
        u5_mult_82_CARRYB_27__39_), .ZN(u5_mult_82_n2323) );
  XNOR2_X2 u5_mult_82_U6625 ( .A(u5_mult_82_n2323), .B(u5_mult_82_SUMB_27__40_), .ZN(u5_mult_82_SUMB_28__39_) );
  NAND2_X2 u5_mult_82_U6624 ( .A1(u5_mult_82_CARRYB_30__22_), .A2(
        u5_mult_82_SUMB_30__23_), .ZN(u5_mult_82_n6304) );
  NAND2_X2 u5_mult_82_U6623 ( .A1(u5_mult_82_ab_31__22_), .A2(
        u5_mult_82_SUMB_30__23_), .ZN(u5_mult_82_n6303) );
  XNOR2_X2 u5_mult_82_U6622 ( .A(u5_mult_82_CARRYB_20__24_), .B(
        u5_mult_82_ab_21__24_), .ZN(u5_mult_82_n2322) );
  XNOR2_X2 u5_mult_82_U6621 ( .A(u5_mult_82_ab_33__24_), .B(
        u5_mult_82_CARRYB_32__24_), .ZN(u5_mult_82_n2321) );
  XNOR2_X2 u5_mult_82_U6620 ( .A(u5_mult_82_n2321), .B(u5_mult_82_SUMB_32__25_), .ZN(u5_mult_82_SUMB_33__24_) );
  NAND2_X2 u5_mult_82_U6619 ( .A1(u5_mult_82_SUMB_8__42_), .A2(
        u5_mult_82_CARRYB_8__41_), .ZN(u5_mult_82_n6105) );
  NAND2_X1 u5_mult_82_U6618 ( .A1(u5_mult_82_CARRYB_12__23_), .A2(
        u5_mult_82_SUMB_12__24_), .ZN(u5_mult_82_n3887) );
  NAND2_X2 u5_mult_82_U6617 ( .A1(u5_mult_82_ab_11__44_), .A2(
        u5_mult_82_SUMB_10__45_), .ZN(u5_mult_82_n5643) );
  NAND3_X4 u5_mult_82_U6616 ( .A1(u5_mult_82_n6236), .A2(u5_mult_82_n6235), 
        .A3(u5_mult_82_n6234), .ZN(u5_mult_82_CARRYB_48__11_) );
  NAND3_X4 u5_mult_82_U6615 ( .A1(u5_mult_82_n2894), .A2(u5_mult_82_n2895), 
        .A3(u5_mult_82_n2896), .ZN(u5_mult_82_CARRYB_29__23_) );
  NAND2_X2 u5_mult_82_U6614 ( .A1(u5_mult_82_CARRYB_29__36_), .A2(
        u5_mult_82_SUMB_29__37_), .ZN(u5_mult_82_n4647) );
  XOR2_X2 u5_mult_82_U6613 ( .A(u5_mult_82_n3512), .B(u5_mult_82_SUMB_27__26_), 
        .Z(u5_mult_82_SUMB_28__25_) );
  NAND2_X2 u5_mult_82_U6612 ( .A1(u5_mult_82_ab_30__36_), .A2(
        u5_mult_82_SUMB_29__37_), .ZN(u5_mult_82_n4646) );
  NAND2_X1 u5_mult_82_U6611 ( .A1(u5_mult_82_ab_11__25_), .A2(
        u5_mult_82_CARRYB_10__25_), .ZN(u5_mult_82_n3900) );
  NAND2_X1 u5_mult_82_U6610 ( .A1(u5_mult_82_CARRYB_10__25_), .A2(
        u5_mult_82_SUMB_10__26_), .ZN(u5_mult_82_n3898) );
  XOR2_X1 u5_mult_82_U6609 ( .A(u5_mult_82_CARRYB_14__23_), .B(
        u5_mult_82_ab_15__23_), .Z(u5_mult_82_n3459) );
  XNOR2_X2 u5_mult_82_U6608 ( .A(u5_mult_82_n2413), .B(u5_mult_82_SUMB_31__28_), .ZN(u5_mult_82_SUMB_32__27_) );
  NAND2_X1 u5_mult_82_U6607 ( .A1(u5_mult_82_ab_45__18_), .A2(u5_mult_82_n721), 
        .ZN(u5_mult_82_n5859) );
  XNOR2_X1 u5_mult_82_U6606 ( .A(u5_mult_82_ab_10__25_), .B(
        u5_mult_82_CARRYB_9__25_), .ZN(u5_mult_82_n2318) );
  XNOR2_X2 u5_mult_82_U6605 ( .A(u5_mult_82_n2318), .B(u5_mult_82_SUMB_9__26_), 
        .ZN(u5_mult_82_SUMB_10__25_) );
  NAND3_X2 u5_mult_82_U6604 ( .A1(u5_mult_82_n2315), .A2(u5_mult_82_n2316), 
        .A3(u5_mult_82_n2317), .ZN(u5_mult_82_CARRYB_24__39_) );
  NAND2_X1 u5_mult_82_U6603 ( .A1(u5_mult_82_CARRYB_23__39_), .A2(
        u5_mult_82_SUMB_23__40_), .ZN(u5_mult_82_n2317) );
  NAND2_X1 u5_mult_82_U6602 ( .A1(u5_mult_82_ab_24__39_), .A2(
        u5_mult_82_SUMB_23__40_), .ZN(u5_mult_82_n2316) );
  NAND2_X1 u5_mult_82_U6601 ( .A1(u5_mult_82_ab_24__39_), .A2(
        u5_mult_82_CARRYB_23__39_), .ZN(u5_mult_82_n2315) );
  NAND2_X2 u5_mult_82_U6600 ( .A1(u5_mult_82_ab_23__40_), .A2(
        u5_mult_82_CARRYB_22__40_), .ZN(u5_mult_82_n2314) );
  NAND2_X2 u5_mult_82_U6599 ( .A1(u5_mult_82_n1708), .A2(
        u5_mult_82_CARRYB_22__40_), .ZN(u5_mult_82_n2313) );
  NAND2_X2 u5_mult_82_U6598 ( .A1(u5_mult_82_n1708), .A2(u5_mult_82_ab_23__40_), .ZN(u5_mult_82_n2312) );
  NAND3_X2 u5_mult_82_U6597 ( .A1(u5_mult_82_n4242), .A2(u5_mult_82_n4243), 
        .A3(u5_mult_82_n4244), .ZN(u5_mult_82_CARRYB_34__22_) );
  XNOR2_X2 u5_mult_82_U6596 ( .A(u5_mult_82_n2309), .B(
        u5_mult_82_CARRYB_12__23_), .ZN(u5_mult_82_n3884) );
  NOR2_X1 u5_mult_82_U6595 ( .A1(u5_mult_82_n6840), .A2(u5_mult_82_n6528), 
        .ZN(u5_mult_82_ab_7__33_) );
  NAND3_X2 u5_mult_82_U6594 ( .A1(u5_mult_82_net85372), .A2(
        u5_mult_82_net85373), .A3(u5_mult_82_n2308), .ZN(
        u5_mult_82_CARRYB_7__33_) );
  NAND2_X1 u5_mult_82_U6593 ( .A1(u5_mult_82_ab_7__33_), .A2(
        u5_mult_82_CARRYB_6__33_), .ZN(u5_mult_82_n2308) );
  XOR2_X2 u5_mult_82_U6592 ( .A(u5_mult_82_CARRYB_6__33_), .B(
        u5_mult_82_ab_7__33_), .Z(u5_mult_82_net85371) );
  NAND2_X1 u5_mult_82_U6591 ( .A1(u5_mult_82_ab_11__29_), .A2(
        u5_mult_82_CARRYB_10__29_), .ZN(u5_mult_82_n2305) );
  NAND3_X4 u5_mult_82_U6590 ( .A1(u5_mult_82_n2302), .A2(u5_mult_82_n2303), 
        .A3(u5_mult_82_n2304), .ZN(u5_mult_82_CARRYB_10__30_) );
  NAND2_X2 u5_mult_82_U6589 ( .A1(u5_mult_82_CARRYB_9__30_), .A2(
        u5_mult_82_SUMB_9__31_), .ZN(u5_mult_82_n2304) );
  NAND2_X2 u5_mult_82_U6588 ( .A1(u5_mult_82_ab_10__30_), .A2(
        u5_mult_82_SUMB_9__31_), .ZN(u5_mult_82_n2303) );
  XOR2_X2 u5_mult_82_U6587 ( .A(u5_mult_82_n2301), .B(u5_mult_82_SUMB_9__31_), 
        .Z(u5_mult_82_SUMB_10__30_) );
  XOR2_X2 u5_mult_82_U6586 ( .A(u5_mult_82_ab_10__30_), .B(
        u5_mult_82_CARRYB_9__30_), .Z(u5_mult_82_n2301) );
  NAND3_X4 u5_mult_82_U6585 ( .A1(u5_mult_82_n2298), .A2(u5_mult_82_n2299), 
        .A3(u5_mult_82_n2300), .ZN(u5_mult_82_CARRYB_29__15_) );
  NAND2_X2 u5_mult_82_U6584 ( .A1(u5_mult_82_CARRYB_28__15_), .A2(
        u5_mult_82_SUMB_28__16_), .ZN(u5_mult_82_n2300) );
  NAND2_X2 u5_mult_82_U6583 ( .A1(u5_mult_82_ab_29__15_), .A2(
        u5_mult_82_SUMB_28__16_), .ZN(u5_mult_82_n2299) );
  NAND2_X1 u5_mult_82_U6582 ( .A1(u5_mult_82_ab_29__15_), .A2(
        u5_mult_82_CARRYB_28__15_), .ZN(u5_mult_82_n2298) );
  NAND3_X4 u5_mult_82_U6581 ( .A1(u5_mult_82_n2295), .A2(u5_mult_82_n2296), 
        .A3(u5_mult_82_n2297), .ZN(u5_mult_82_CARRYB_28__16_) );
  NAND2_X2 u5_mult_82_U6580 ( .A1(u5_mult_82_CARRYB_27__16_), .A2(
        u5_mult_82_n1498), .ZN(u5_mult_82_n2297) );
  NAND2_X2 u5_mult_82_U6579 ( .A1(u5_mult_82_ab_28__16_), .A2(u5_mult_82_n1498), .ZN(u5_mult_82_n2296) );
  NAND2_X2 u5_mult_82_U6578 ( .A1(u5_mult_82_ab_28__16_), .A2(
        u5_mult_82_CARRYB_27__16_), .ZN(u5_mult_82_n2295) );
  XOR2_X2 u5_mult_82_U6577 ( .A(u5_mult_82_n2294), .B(u5_mult_82_n1498), .Z(
        u5_mult_82_SUMB_28__16_) );
  XOR2_X2 u5_mult_82_U6576 ( .A(u5_mult_82_ab_28__16_), .B(
        u5_mult_82_CARRYB_27__16_), .Z(u5_mult_82_n2294) );
  NAND2_X2 u5_mult_82_U6575 ( .A1(u5_mult_82_ab_31__36_), .A2(
        u5_mult_82_SUMB_30__37_), .ZN(u5_mult_82_n4320) );
  XNOR2_X2 u5_mult_82_U6574 ( .A(u5_mult_82_n2293), .B(
        u5_mult_82_CARRYB_33__8_), .ZN(u5_mult_82_n4520) );
  XOR2_X2 u5_mult_82_U6573 ( .A(u5_mult_82_ab_5__45_), .B(
        u5_mult_82_CARRYB_4__45_), .Z(u5_mult_82_n4992) );
  NAND3_X4 u5_mult_82_U6572 ( .A1(u5_mult_82_n5857), .A2(u5_mult_82_n5858), 
        .A3(u5_mult_82_n5859), .ZN(u5_mult_82_CARRYB_45__18_) );
  NAND2_X2 u5_mult_82_U6571 ( .A1(u5_mult_82_ab_47__0_), .A2(
        u5_mult_82_CARRYB_46__0_), .ZN(u5_mult_82_n4278) );
  NAND2_X2 u5_mult_82_U6570 ( .A1(u5_mult_82_CARRYB_23__41_), .A2(
        u5_mult_82_n1691), .ZN(u5_mult_82_n2903) );
  NAND2_X2 u5_mult_82_U6569 ( .A1(u5_mult_82_CARRYB_28__13_), .A2(
        u5_mult_82_SUMB_28__14_), .ZN(u5_mult_82_n2793) );
  NAND2_X2 u5_mult_82_U6568 ( .A1(u5_mult_82_ab_29__13_), .A2(
        u5_mult_82_SUMB_28__14_), .ZN(u5_mult_82_n2792) );
  XNOR2_X2 u5_mult_82_U6567 ( .A(u5_mult_82_n2292), .B(
        u5_mult_82_CARRYB_42__19_), .ZN(u5_mult_82_n5833) );
  NAND2_X2 u5_mult_82_U6566 ( .A1(u5_mult_82_ab_30__29_), .A2(
        u5_mult_82_SUMB_29__30_), .ZN(u5_mult_82_n4538) );
  XNOR2_X2 u5_mult_82_U6565 ( .A(u5_mult_82_ab_24__39_), .B(
        u5_mult_82_CARRYB_23__39_), .ZN(u5_mult_82_n2291) );
  XNOR2_X2 u5_mult_82_U6564 ( .A(u5_mult_82_n2291), .B(u5_mult_82_SUMB_23__40_), .ZN(u5_mult_82_SUMB_24__39_) );
  NAND3_X4 u5_mult_82_U6563 ( .A1(u5_mult_82_n3027), .A2(u5_mult_82_n3028), 
        .A3(u5_mult_82_n3029), .ZN(u5_mult_82_CARRYB_23__41_) );
  XNOR2_X2 u5_mult_82_U6562 ( .A(u5_mult_82_CARRYB_25__14_), .B(
        u5_mult_82_ab_26__14_), .ZN(u5_mult_82_n2290) );
  NAND2_X2 u5_mult_82_U6561 ( .A1(u5_mult_82_n5297), .A2(u5_mult_82_n1419), 
        .ZN(u5_mult_82_n3541) );
  NAND2_X1 u5_mult_82_U6560 ( .A1(u5_mult_82_CARRYB_14__42_), .A2(
        u5_mult_82_SUMB_14__43_), .ZN(u5_mult_82_n3133) );
  NAND2_X1 u5_mult_82_U6559 ( .A1(u5_mult_82_CARRYB_44__20_), .A2(
        u5_mult_82_SUMB_44__21_), .ZN(u5_mult_82_n3847) );
  XNOR2_X2 u5_mult_82_U6558 ( .A(u5_mult_82_CARRYB_10__25_), .B(
        u5_mult_82_ab_11__25_), .ZN(u5_mult_82_n2289) );
  XNOR2_X2 u5_mult_82_U6557 ( .A(u5_mult_82_SUMB_10__26_), .B(u5_mult_82_n2289), .ZN(u5_mult_82_SUMB_11__25_) );
  NAND2_X2 u5_mult_82_U6556 ( .A1(u5_mult_82_CARRYB_52__10_), .A2(
        u5_mult_82_SUMB_52__11_), .ZN(u5_mult_82_n4692) );
  XNOR2_X2 u5_mult_82_U6555 ( .A(u5_mult_82_ab_6__47_), .B(
        u5_mult_82_CARRYB_5__47_), .ZN(u5_mult_82_n2287) );
  XNOR2_X2 u5_mult_82_U6554 ( .A(u5_mult_82_n2287), .B(u5_mult_82_n1822), .ZN(
        u5_mult_82_SUMB_6__47_) );
  NAND2_X1 u5_mult_82_U6553 ( .A1(u5_mult_82_ab_35__36_), .A2(
        u5_mult_82_CARRYB_34__36_), .ZN(u5_mult_82_n5081) );
  NAND2_X2 u5_mult_82_U6552 ( .A1(u5_mult_82_ab_9__41_), .A2(
        u5_mult_82_SUMB_8__42_), .ZN(u5_mult_82_n6104) );
  NAND2_X1 u5_mult_82_U6551 ( .A1(u5_mult_82_CARRYB_24__12_), .A2(
        u5_mult_82_SUMB_24__13_), .ZN(u5_mult_82_n2286) );
  NAND2_X1 u5_mult_82_U6550 ( .A1(u5_mult_82_ab_25__12_), .A2(
        u5_mult_82_SUMB_24__13_), .ZN(u5_mult_82_n2285) );
  NAND2_X1 u5_mult_82_U6549 ( .A1(u5_mult_82_ab_25__12_), .A2(
        u5_mult_82_CARRYB_24__12_), .ZN(u5_mult_82_n2284) );
  NAND3_X4 u5_mult_82_U6548 ( .A1(u5_mult_82_n2281), .A2(u5_mult_82_n2282), 
        .A3(u5_mult_82_n2283), .ZN(u5_mult_82_CARRYB_24__13_) );
  NAND2_X2 u5_mult_82_U6547 ( .A1(u5_mult_82_n1596), .A2(
        u5_mult_82_SUMB_23__14_), .ZN(u5_mult_82_n2283) );
  NAND2_X2 u5_mult_82_U6546 ( .A1(u5_mult_82_ab_24__13_), .A2(
        u5_mult_82_SUMB_23__14_), .ZN(u5_mult_82_n2282) );
  NAND2_X1 u5_mult_82_U6545 ( .A1(u5_mult_82_ab_24__13_), .A2(
        u5_mult_82_CARRYB_23__13_), .ZN(u5_mult_82_n2281) );
  XOR2_X2 u5_mult_82_U6544 ( .A(u5_mult_82_n2280), .B(u5_mult_82_SUMB_24__13_), 
        .Z(u5_mult_82_SUMB_25__12_) );
  XOR2_X2 u5_mult_82_U6543 ( .A(u5_mult_82_n2279), .B(u5_mult_82_SUMB_23__14_), 
        .Z(u5_mult_82_SUMB_24__13_) );
  XOR2_X2 u5_mult_82_U6542 ( .A(u5_mult_82_ab_24__13_), .B(
        u5_mult_82_CARRYB_23__13_), .Z(u5_mult_82_n2279) );
  NAND2_X2 u5_mult_82_U6541 ( .A1(u5_mult_82_SUMB_50__12_), .A2(
        u5_mult_82_ab_51__11_), .ZN(u5_mult_82_n4696) );
  NAND2_X2 u5_mult_82_U6540 ( .A1(u5_mult_82_n721), .A2(
        u5_mult_82_SUMB_44__19_), .ZN(u5_mult_82_n5857) );
  XNOR2_X2 u5_mult_82_U6539 ( .A(u5_mult_82_SUMB_44__18_), .B(
        u5_mult_82_ab_45__17_), .ZN(u5_mult_82_n2412) );
  NAND2_X2 u5_mult_82_U6538 ( .A1(u5_mult_82_SUMB_27__30_), .A2(
        u5_mult_82_CARRYB_27__29_), .ZN(u5_mult_82_n5477) );
  NAND2_X4 u5_mult_82_U6537 ( .A1(u5_mult_82_ab_43__4_), .A2(u5_mult_82_n3707), 
        .ZN(u5_mult_82_n4677) );
  NAND2_X2 u5_mult_82_U6536 ( .A1(u5_mult_82_CARRYB_50__11_), .A2(
        u5_mult_82_SUMB_50__12_), .ZN(u5_mult_82_n4695) );
  NAND3_X4 u5_mult_82_U6535 ( .A1(u5_mult_82_n2901), .A2(u5_mult_82_n2902), 
        .A3(u5_mult_82_n2903), .ZN(u5_mult_82_CARRYB_24__41_) );
  NAND2_X2 u5_mult_82_U6534 ( .A1(u5_mult_82_ab_25__41_), .A2(
        u5_mult_82_CARRYB_24__41_), .ZN(u5_mult_82_n3079) );
  XOR2_X1 u5_mult_82_U6533 ( .A(u5_mult_82_n14), .B(u5_mult_82_ab_43__0_), .Z(
        u5_mult_82_n4836) );
  CLKBUF_X3 u5_mult_82_U6532 ( .A(u5_mult_82_CARRYB_33__30_), .Z(
        u5_mult_82_n3825) );
  NAND2_X2 u5_mult_82_U6531 ( .A1(u5_mult_82_n37), .A2(
        u5_mult_82_CARRYB_18__25_), .ZN(u5_mult_82_n5610) );
  NAND3_X2 u5_mult_82_U6530 ( .A1(u5_mult_82_n2276), .A2(u5_mult_82_n2277), 
        .A3(u5_mult_82_n2278), .ZN(u5_mult_82_CARRYB_33__51_) );
  NAND2_X2 u5_mult_82_U6529 ( .A1(u5_mult_82_ab_32__52_), .A2(
        u5_mult_82_CARRYB_32__51_), .ZN(u5_mult_82_n2278) );
  NAND2_X2 u5_mult_82_U6528 ( .A1(u5_mult_82_ab_33__51_), .A2(
        u5_mult_82_CARRYB_32__51_), .ZN(u5_mult_82_n2277) );
  NAND2_X2 u5_mult_82_U6527 ( .A1(u5_mult_82_ab_33__51_), .A2(
        u5_mult_82_ab_32__52_), .ZN(u5_mult_82_n2276) );
  XOR2_X1 u5_mult_82_U6526 ( .A(u5_mult_82_n2275), .B(
        u5_mult_82_CARRYB_32__51_), .Z(u5_mult_82_SUMB_33__51_) );
  XOR2_X2 u5_mult_82_U6525 ( .A(u5_mult_82_ab_33__51_), .B(
        u5_mult_82_ab_32__52_), .Z(u5_mult_82_n2275) );
  NAND3_X2 u5_mult_82_U6524 ( .A1(u5_mult_82_n2272), .A2(u5_mult_82_n2273), 
        .A3(u5_mult_82_n2274), .ZN(u5_mult_82_CARRYB_32__51_) );
  NAND2_X1 u5_mult_82_U6523 ( .A1(u5_mult_82_CARRYB_31__51_), .A2(
        u5_mult_82_ab_31__52_), .ZN(u5_mult_82_n2274) );
  NAND2_X2 u5_mult_82_U6522 ( .A1(u5_mult_82_ab_32__51_), .A2(
        u5_mult_82_ab_31__52_), .ZN(u5_mult_82_n2273) );
  NAND2_X1 u5_mult_82_U6521 ( .A1(u5_mult_82_ab_32__51_), .A2(
        u5_mult_82_CARRYB_31__51_), .ZN(u5_mult_82_n2272) );
  XOR2_X2 u5_mult_82_U6520 ( .A(u5_mult_82_n2271), .B(u5_mult_82_ab_31__52_), 
        .Z(u5_mult_82_SUMB_32__51_) );
  XOR2_X2 u5_mult_82_U6519 ( .A(u5_mult_82_ab_32__51_), .B(
        u5_mult_82_CARRYB_31__51_), .Z(u5_mult_82_n2271) );
  NAND3_X2 u5_mult_82_U6518 ( .A1(u5_mult_82_n2268), .A2(u5_mult_82_n2269), 
        .A3(u5_mult_82_n2270), .ZN(u5_mult_82_CARRYB_45__43_) );
  NAND2_X1 u5_mult_82_U6517 ( .A1(u5_mult_82_CARRYB_44__43_), .A2(
        u5_mult_82_SUMB_44__44_), .ZN(u5_mult_82_n2270) );
  NAND2_X1 u5_mult_82_U6516 ( .A1(u5_mult_82_ab_45__43_), .A2(
        u5_mult_82_SUMB_44__44_), .ZN(u5_mult_82_n2269) );
  NAND2_X1 u5_mult_82_U6515 ( .A1(u5_mult_82_ab_45__43_), .A2(
        u5_mult_82_CARRYB_44__43_), .ZN(u5_mult_82_n2268) );
  NAND2_X2 u5_mult_82_U6514 ( .A1(u5_mult_82_CARRYB_43__44_), .A2(
        u5_mult_82_SUMB_43__45_), .ZN(u5_mult_82_n2267) );
  NAND2_X2 u5_mult_82_U6513 ( .A1(u5_mult_82_ab_44__44_), .A2(
        u5_mult_82_SUMB_43__45_), .ZN(u5_mult_82_n2266) );
  NAND2_X1 u5_mult_82_U6512 ( .A1(u5_mult_82_ab_44__44_), .A2(
        u5_mult_82_CARRYB_43__44_), .ZN(u5_mult_82_n2265) );
  XOR2_X2 u5_mult_82_U6511 ( .A(u5_mult_82_n2264), .B(u5_mult_82_SUMB_44__44_), 
        .Z(u5_mult_82_SUMB_45__43_) );
  XOR2_X2 u5_mult_82_U6510 ( .A(u5_mult_82_ab_45__43_), .B(
        u5_mult_82_CARRYB_44__43_), .Z(u5_mult_82_n2264) );
  XOR2_X2 u5_mult_82_U6509 ( .A(u5_mult_82_n2263), .B(u5_mult_82_SUMB_43__45_), 
        .Z(u5_mult_82_SUMB_44__44_) );
  XOR2_X2 u5_mult_82_U6508 ( .A(u5_mult_82_ab_44__44_), .B(
        u5_mult_82_CARRYB_43__44_), .Z(u5_mult_82_n2263) );
  NAND2_X2 u5_mult_82_U6507 ( .A1(u5_mult_82_ab_26__13_), .A2(
        u5_mult_82_SUMB_25__14_), .ZN(u5_mult_82_n4834) );
  NAND3_X2 u5_mult_82_U6506 ( .A1(u5_mult_82_n2987), .A2(u5_mult_82_n2988), 
        .A3(u5_mult_82_n2989), .ZN(u5_mult_82_CARRYB_39__7_) );
  NAND2_X2 u5_mult_82_U6505 ( .A1(u5_mult_82_CARRYB_43__5_), .A2(
        u5_mult_82_SUMB_43__6_), .ZN(u5_mult_82_n6033) );
  NAND3_X4 u5_mult_82_U6504 ( .A1(u5_mult_82_n6033), .A2(u5_mult_82_n6034), 
        .A3(u5_mult_82_n6035), .ZN(u5_mult_82_CARRYB_44__5_) );
  XNOR2_X2 u5_mult_82_U6503 ( .A(u5_mult_82_n2261), .B(
        u5_mult_82_CARRYB_29__39_), .ZN(u5_mult_82_n2457) );
  NAND2_X2 u5_mult_82_U6502 ( .A1(u5_mult_82_CARRYB_33__25_), .A2(
        u5_mult_82_SUMB_33__26_), .ZN(u5_mult_82_n3390) );
  NAND2_X1 u5_mult_82_U6501 ( .A1(u5_mult_82_ab_36__20_), .A2(
        u5_mult_82_CARRYB_35__20_), .ZN(u5_mult_82_n6277) );
  BUF_X8 u5_mult_82_U6500 ( .A(u5_mult_82_SUMB_21__39_), .Z(u5_mult_82_n2260)
         );
  NAND2_X2 u5_mult_82_U6499 ( .A1(u5_mult_82_ab_23__37_), .A2(
        u5_mult_82_SUMB_22__38_), .ZN(u5_mult_82_n2258) );
  NAND2_X1 u5_mult_82_U6498 ( .A1(u5_mult_82_ab_23__37_), .A2(
        u5_mult_82_CARRYB_22__37_), .ZN(u5_mult_82_n2257) );
  NAND3_X4 u5_mult_82_U6497 ( .A1(u5_mult_82_n2251), .A2(u5_mult_82_n2252), 
        .A3(u5_mult_82_n2253), .ZN(u5_mult_82_CARRYB_42__21_) );
  NAND2_X1 u5_mult_82_U6496 ( .A1(u5_mult_82_ab_42__21_), .A2(
        u5_mult_82_CARRYB_41__21_), .ZN(u5_mult_82_n2251) );
  NAND3_X2 u5_mult_82_U6495 ( .A1(u5_mult_82_n2248), .A2(u5_mult_82_n2249), 
        .A3(u5_mult_82_n2250), .ZN(u5_mult_82_CARRYB_41__22_) );
  NAND2_X1 u5_mult_82_U6494 ( .A1(u5_mult_82_CARRYB_40__22_), .A2(
        u5_mult_82_SUMB_40__23_), .ZN(u5_mult_82_n2249) );
  XOR2_X2 u5_mult_82_U6493 ( .A(u5_mult_82_n2247), .B(u5_mult_82_SUMB_41__22_), 
        .Z(u5_mult_82_SUMB_42__21_) );
  XOR2_X2 u5_mult_82_U6492 ( .A(u5_mult_82_n2246), .B(u5_mult_82_SUMB_40__23_), 
        .Z(u5_mult_82_SUMB_41__22_) );
  XOR2_X2 u5_mult_82_U6491 ( .A(u5_mult_82_CARRYB_40__22_), .B(
        u5_mult_82_ab_41__22_), .Z(u5_mult_82_n2246) );
  NAND2_X1 u5_mult_82_U6490 ( .A1(u5_mult_82_CARRYB_39__23_), .A2(
        u5_mult_82_SUMB_39__24_), .ZN(u5_mult_82_n2245) );
  NAND2_X1 u5_mult_82_U6489 ( .A1(u5_mult_82_ab_40__23_), .A2(
        u5_mult_82_SUMB_39__24_), .ZN(u5_mult_82_n2244) );
  NAND2_X1 u5_mult_82_U6488 ( .A1(u5_mult_82_ab_40__23_), .A2(
        u5_mult_82_CARRYB_39__23_), .ZN(u5_mult_82_n2243) );
  NAND3_X4 u5_mult_82_U6487 ( .A1(u5_mult_82_n2240), .A2(u5_mult_82_n2241), 
        .A3(u5_mult_82_n2242), .ZN(u5_mult_82_CARRYB_39__24_) );
  NAND2_X2 u5_mult_82_U6486 ( .A1(u5_mult_82_ab_39__24_), .A2(u5_mult_82_n1812), .ZN(u5_mult_82_n2242) );
  NAND2_X2 u5_mult_82_U6485 ( .A1(u5_mult_82_CARRYB_38__24_), .A2(
        u5_mult_82_n1812), .ZN(u5_mult_82_n2241) );
  NAND2_X1 u5_mult_82_U6484 ( .A1(u5_mult_82_CARRYB_38__24_), .A2(
        u5_mult_82_ab_39__24_), .ZN(u5_mult_82_n2240) );
  XOR2_X2 u5_mult_82_U6483 ( .A(u5_mult_82_n2239), .B(u5_mult_82_SUMB_39__24_), 
        .Z(u5_mult_82_SUMB_40__23_) );
  NAND2_X2 u5_mult_82_U6482 ( .A1(u5_mult_82_CARRYB_29__22_), .A2(
        u5_mult_82_SUMB_29__23_), .ZN(u5_mult_82_n2899) );
  NAND3_X4 u5_mult_82_U6481 ( .A1(u5_mult_82_n5014), .A2(u5_mult_82_n5015), 
        .A3(u5_mult_82_n5016), .ZN(u5_mult_82_CARRYB_40__15_) );
  NAND3_X4 u5_mult_82_U6480 ( .A1(u5_mult_82_n6201), .A2(u5_mult_82_n6200), 
        .A3(u5_mult_82_n6199), .ZN(u5_mult_82_CARRYB_50__8_) );
  NAND2_X2 u5_mult_82_U6479 ( .A1(u5_mult_82_ab_15__23_), .A2(
        u5_mult_82_SUMB_14__24_), .ZN(u5_mult_82_n3461) );
  NAND3_X2 u5_mult_82_U6478 ( .A1(u5_mult_82_n2507), .A2(u5_mult_82_n2508), 
        .A3(u5_mult_82_n2509), .ZN(u5_mult_82_CARRYB_8__28_) );
  XOR2_X2 u5_mult_82_U6477 ( .A(u5_mult_82_n2750), .B(
        u5_mult_82_CARRYB_20__26_), .Z(u5_mult_82_n2238) );
  XNOR2_X2 u5_mult_82_U6476 ( .A(u5_mult_82_n2238), .B(u5_mult_82_SUMB_20__27_), .ZN(u5_mult_82_SUMB_21__26_) );
  NAND2_X1 u5_mult_82_U6475 ( .A1(u5_mult_82_CARRYB_43__43_), .A2(
        u5_mult_82_SUMB_43__44_), .ZN(u5_mult_82_n2237) );
  NAND2_X1 u5_mult_82_U6474 ( .A1(u5_mult_82_ab_44__43_), .A2(
        u5_mult_82_SUMB_43__44_), .ZN(u5_mult_82_n2236) );
  NAND2_X1 u5_mult_82_U6473 ( .A1(u5_mult_82_ab_44__43_), .A2(
        u5_mult_82_CARRYB_43__43_), .ZN(u5_mult_82_n2235) );
  NAND3_X4 u5_mult_82_U6472 ( .A1(u5_mult_82_n2232), .A2(u5_mult_82_n2233), 
        .A3(u5_mult_82_n2234), .ZN(u5_mult_82_CARRYB_43__44_) );
  NAND2_X2 u5_mult_82_U6471 ( .A1(u5_mult_82_CARRYB_42__44_), .A2(
        u5_mult_82_SUMB_42__45_), .ZN(u5_mult_82_n2234) );
  NAND2_X2 u5_mult_82_U6470 ( .A1(u5_mult_82_ab_43__44_), .A2(
        u5_mult_82_SUMB_42__45_), .ZN(u5_mult_82_n2233) );
  NAND2_X1 u5_mult_82_U6469 ( .A1(u5_mult_82_ab_43__44_), .A2(
        u5_mult_82_CARRYB_42__44_), .ZN(u5_mult_82_n2232) );
  XOR2_X2 u5_mult_82_U6468 ( .A(u5_mult_82_n2231), .B(u5_mult_82_SUMB_43__44_), 
        .Z(u5_mult_82_SUMB_44__43_) );
  XOR2_X2 u5_mult_82_U6467 ( .A(u5_mult_82_ab_44__43_), .B(
        u5_mult_82_CARRYB_43__43_), .Z(u5_mult_82_n2231) );
  XOR2_X2 u5_mult_82_U6466 ( .A(u5_mult_82_n2230), .B(u5_mult_82_SUMB_42__45_), 
        .Z(u5_mult_82_SUMB_43__44_) );
  XOR2_X2 u5_mult_82_U6465 ( .A(u5_mult_82_ab_43__44_), .B(
        u5_mult_82_CARRYB_42__44_), .Z(u5_mult_82_n2230) );
  NAND3_X2 u5_mult_82_U6464 ( .A1(u5_mult_82_n2227), .A2(u5_mult_82_n2228), 
        .A3(u5_mult_82_n2229), .ZN(u5_mult_82_CARRYB_50__37_) );
  NAND2_X2 u5_mult_82_U6463 ( .A1(u5_mult_82_CARRYB_49__37_), .A2(
        u5_mult_82_SUMB_49__38_), .ZN(u5_mult_82_n2229) );
  NAND2_X2 u5_mult_82_U6462 ( .A1(u5_mult_82_ab_50__37_), .A2(
        u5_mult_82_SUMB_49__38_), .ZN(u5_mult_82_n2228) );
  NAND2_X1 u5_mult_82_U6461 ( .A1(u5_mult_82_ab_50__37_), .A2(
        u5_mult_82_CARRYB_49__37_), .ZN(u5_mult_82_n2227) );
  NAND3_X4 u5_mult_82_U6460 ( .A1(u5_mult_82_n2224), .A2(u5_mult_82_n2225), 
        .A3(u5_mult_82_n2226), .ZN(u5_mult_82_CARRYB_49__38_) );
  NAND2_X2 u5_mult_82_U6459 ( .A1(u5_mult_82_CARRYB_48__38_), .A2(
        u5_mult_82_SUMB_48__39_), .ZN(u5_mult_82_n2226) );
  NAND2_X2 u5_mult_82_U6458 ( .A1(u5_mult_82_ab_49__38_), .A2(
        u5_mult_82_SUMB_48__39_), .ZN(u5_mult_82_n2225) );
  NAND2_X1 u5_mult_82_U6457 ( .A1(u5_mult_82_ab_49__38_), .A2(
        u5_mult_82_CARRYB_48__38_), .ZN(u5_mult_82_n2224) );
  XOR2_X2 u5_mult_82_U6456 ( .A(u5_mult_82_n2223), .B(u5_mult_82_SUMB_49__38_), 
        .Z(u5_mult_82_SUMB_50__37_) );
  XOR2_X2 u5_mult_82_U6455 ( .A(u5_mult_82_ab_50__37_), .B(
        u5_mult_82_CARRYB_49__37_), .Z(u5_mult_82_n2223) );
  XOR2_X2 u5_mult_82_U6454 ( .A(u5_mult_82_n2222), .B(u5_mult_82_SUMB_48__39_), 
        .Z(u5_mult_82_SUMB_49__38_) );
  XOR2_X2 u5_mult_82_U6453 ( .A(u5_mult_82_ab_49__38_), .B(
        u5_mult_82_CARRYB_48__38_), .Z(u5_mult_82_n2222) );
  NAND3_X4 u5_mult_82_U6452 ( .A1(u5_mult_82_n3006), .A2(u5_mult_82_n3007), 
        .A3(u5_mult_82_n3008), .ZN(u5_mult_82_CARRYB_48__34_) );
  INV_X8 u5_mult_82_U6451 ( .A(u5_mult_82_n6789), .ZN(u5_mult_82_n6796) );
  NAND3_X4 u5_mult_82_U6450 ( .A1(u5_mult_82_n3040), .A2(u5_mult_82_n3039), 
        .A3(u5_mult_82_n3038), .ZN(u5_mult_82_CARRYB_43__33_) );
  NOR2_X1 u5_mult_82_U6449 ( .A1(u5_mult_82_n6831), .A2(u5_mult_82_n6742), 
        .ZN(u5_mult_82_ab_46__39_) );
  NOR2_X1 u5_mult_82_U6448 ( .A1(u5_mult_82_n6831), .A2(u5_mult_82_net65315), 
        .ZN(u5_mult_82_ab_45__39_) );
  NAND2_X1 u5_mult_82_U6447 ( .A1(u5_mult_82_ab_46__39_), .A2(
        u5_mult_82_CARRYB_45__39_), .ZN(u5_mult_82_n2221) );
  NAND2_X2 u5_mult_82_U6446 ( .A1(u5_mult_82_ab_46__39_), .A2(
        u5_mult_82_SUMB_45__40_), .ZN(u5_mult_82_n2220) );
  NAND2_X1 u5_mult_82_U6445 ( .A1(u5_mult_82_CARRYB_45__39_), .A2(
        u5_mult_82_SUMB_45__40_), .ZN(u5_mult_82_n2219) );
  XOR2_X2 u5_mult_82_U6444 ( .A(u5_mult_82_SUMB_45__40_), .B(u5_mult_82_n2218), 
        .Z(u5_mult_82_SUMB_46__39_) );
  XOR2_X2 u5_mult_82_U6443 ( .A(u5_mult_82_CARRYB_45__39_), .B(
        u5_mult_82_ab_46__39_), .Z(u5_mult_82_n2218) );
  NAND3_X2 u5_mult_82_U6442 ( .A1(u5_mult_82_n2215), .A2(u5_mult_82_n2216), 
        .A3(u5_mult_82_n2217), .ZN(u5_mult_82_CARRYB_45__39_) );
  NAND2_X1 u5_mult_82_U6441 ( .A1(u5_mult_82_ab_45__39_), .A2(
        u5_mult_82_CARRYB_44__39_), .ZN(u5_mult_82_n2217) );
  NAND2_X2 u5_mult_82_U6440 ( .A1(u5_mult_82_ab_45__39_), .A2(
        u5_mult_82_SUMB_44__40_), .ZN(u5_mult_82_n2216) );
  NAND2_X1 u5_mult_82_U6439 ( .A1(u5_mult_82_CARRYB_44__39_), .A2(
        u5_mult_82_SUMB_44__40_), .ZN(u5_mult_82_n2215) );
  XOR2_X2 u5_mult_82_U6438 ( .A(u5_mult_82_SUMB_44__40_), .B(u5_mult_82_n2214), 
        .Z(u5_mult_82_SUMB_45__39_) );
  XOR2_X2 u5_mult_82_U6437 ( .A(u5_mult_82_CARRYB_44__39_), .B(
        u5_mult_82_ab_45__39_), .Z(u5_mult_82_n2214) );
  INV_X2 u5_mult_82_U6436 ( .A(u5_mult_82_ab_26__40_), .ZN(u5_mult_82_n2288)
         );
  INV_X4 u5_mult_82_U6435 ( .A(u5_mult_82_n2174), .ZN(u5_mult_82_n2211) );
  NAND2_X1 u5_mult_82_U6434 ( .A1(u5_mult_82_n2288), .A2(u5_mult_82_n2174), 
        .ZN(u5_mult_82_n2212) );
  NAND2_X2 u5_mult_82_U6433 ( .A1(u5_mult_82_CARRYB_8__29_), .A2(
        u5_mult_82_SUMB_8__30_), .ZN(u5_mult_82_n2210) );
  NAND2_X2 u5_mult_82_U6432 ( .A1(u5_mult_82_ab_9__29_), .A2(
        u5_mult_82_SUMB_8__30_), .ZN(u5_mult_82_n2209) );
  NAND2_X1 u5_mult_82_U6431 ( .A1(u5_mult_82_ab_9__29_), .A2(
        u5_mult_82_CARRYB_8__29_), .ZN(u5_mult_82_n2208) );
  NAND2_X2 u5_mult_82_U6430 ( .A1(u5_mult_82_ab_8__30_), .A2(
        u5_mult_82_SUMB_7__31_), .ZN(u5_mult_82_n2206) );
  NAND2_X1 u5_mult_82_U6429 ( .A1(u5_mult_82_ab_8__30_), .A2(
        u5_mult_82_CARRYB_7__30_), .ZN(u5_mult_82_n2205) );
  NAND3_X4 u5_mult_82_U6428 ( .A1(u5_mult_82_n2202), .A2(u5_mult_82_n2203), 
        .A3(u5_mult_82_n2204), .ZN(u5_mult_82_CARRYB_13__25_) );
  NAND2_X1 u5_mult_82_U6427 ( .A1(u5_mult_82_ab_13__25_), .A2(
        u5_mult_82_CARRYB_12__25_), .ZN(u5_mult_82_n2202) );
  NAND3_X4 u5_mult_82_U6426 ( .A1(u5_mult_82_n2199), .A2(u5_mult_82_n2200), 
        .A3(u5_mult_82_n2201), .ZN(u5_mult_82_CARRYB_12__26_) );
  NAND2_X2 u5_mult_82_U6425 ( .A1(u5_mult_82_ab_12__26_), .A2(
        u5_mult_82_SUMB_11__27_), .ZN(u5_mult_82_n2201) );
  NAND2_X1 u5_mult_82_U6424 ( .A1(u5_mult_82_CARRYB_11__26_), .A2(
        u5_mult_82_ab_12__26_), .ZN(u5_mult_82_n2199) );
  NAND2_X1 u5_mult_82_U6423 ( .A1(u5_mult_82_ab_4__37_), .A2(
        u5_mult_82_SUMB_3__38_), .ZN(u5_mult_82_n5326) );
  NAND2_X1 u5_mult_82_U6422 ( .A1(u5_mult_82_CARRYB_3__37_), .A2(
        u5_mult_82_SUMB_3__38_), .ZN(u5_mult_82_n5327) );
  NAND3_X2 u5_mult_82_U6421 ( .A1(u5_mult_82_n5327), .A2(u5_mult_82_n5326), 
        .A3(u5_mult_82_n5325), .ZN(u5_mult_82_CARRYB_4__37_) );
  XNOR2_X2 u5_mult_82_U6420 ( .A(u5_mult_82_n2198), .B(u5_mult_82_SUMB_24__10_), .ZN(u5_mult_82_n3434) );
  NAND3_X4 u5_mult_82_U6419 ( .A1(u5_mult_82_n2529), .A2(u5_mult_82_n2530), 
        .A3(u5_mult_82_n2531), .ZN(u5_mult_82_CARRYB_21__30_) );
  NAND2_X2 u5_mult_82_U6418 ( .A1(u5_mult_82_ab_48__14_), .A2(
        u5_mult_82_SUMB_47__15_), .ZN(u5_mult_82_n5773) );
  NAND2_X2 u5_mult_82_U6417 ( .A1(u5_mult_82_ab_50__13_), .A2(
        u5_mult_82_SUMB_49__14_), .ZN(u5_mult_82_n5829) );
  NAND3_X2 u5_mult_82_U6416 ( .A1(u5_mult_82_n2197), .A2(u5_mult_82_n2196), 
        .A3(u5_mult_82_n2195), .ZN(u5_mult_82_CARRYB_23__24_) );
  NAND2_X1 u5_mult_82_U6415 ( .A1(u5_mult_82_ab_23__24_), .A2(
        u5_mult_82_SUMB_22__25_), .ZN(u5_mult_82_n2197) );
  NAND2_X1 u5_mult_82_U6414 ( .A1(u5_mult_82_CARRYB_22__24_), .A2(
        u5_mult_82_ab_23__24_), .ZN(u5_mult_82_n2195) );
  NAND2_X2 u5_mult_82_U6413 ( .A1(u5_mult_82_ab_22__25_), .A2(
        u5_mult_82_SUMB_21__26_), .ZN(u5_mult_82_n2193) );
  NAND2_X2 u5_mult_82_U6412 ( .A1(u5_mult_82_CARRYB_20__25_), .A2(
        u5_mult_82_SUMB_20__26_), .ZN(u5_mult_82_n2191) );
  NAND2_X2 u5_mult_82_U6411 ( .A1(u5_mult_82_ab_21__25_), .A2(
        u5_mult_82_SUMB_20__26_), .ZN(u5_mult_82_n2190) );
  NAND3_X2 u5_mult_82_U6410 ( .A1(u5_mult_82_net85540), .A2(
        u5_mult_82_net85541), .A3(u5_mult_82_n2188), .ZN(
        u5_mult_82_CARRYB_20__26_) );
  NAND2_X2 u5_mult_82_U6409 ( .A1(u5_mult_82_ab_20__26_), .A2(
        u5_mult_82_SUMB_19__27_), .ZN(u5_mult_82_n2188) );
  INV_X8 u5_mult_82_U6408 ( .A(u5_mult_82_n6795), .ZN(u5_mult_82_n6794) );
  NOR2_X1 u5_mult_82_U6407 ( .A1(u5_mult_82_n6774), .A2(u5_mult_82_n6593), 
        .ZN(u5_mult_82_ab_16__49_) );
  NAND3_X2 u5_mult_82_U6406 ( .A1(u5_mult_82_n2185), .A2(u5_mult_82_n2186), 
        .A3(u5_mult_82_n2187), .ZN(u5_mult_82_CARRYB_16__49_) );
  NAND2_X1 u5_mult_82_U6405 ( .A1(u5_mult_82_ab_16__49_), .A2(
        u5_mult_82_SUMB_15__50_), .ZN(u5_mult_82_n2187) );
  NAND2_X2 u5_mult_82_U6404 ( .A1(u5_mult_82_ab_16__49_), .A2(
        u5_mult_82_CARRYB_15__49_), .ZN(u5_mult_82_n2186) );
  NAND2_X1 u5_mult_82_U6403 ( .A1(u5_mult_82_SUMB_15__50_), .A2(
        u5_mult_82_CARRYB_15__49_), .ZN(u5_mult_82_n2185) );
  XOR2_X2 u5_mult_82_U6402 ( .A(u5_mult_82_CARRYB_15__49_), .B(
        u5_mult_82_n2184), .Z(u5_mult_82_SUMB_16__49_) );
  XOR2_X2 u5_mult_82_U6401 ( .A(u5_mult_82_SUMB_15__50_), .B(
        u5_mult_82_ab_16__49_), .Z(u5_mult_82_n2184) );
  NAND2_X1 u5_mult_82_U6400 ( .A1(u5_mult_82_CARRYB_28__41_), .A2(
        u5_mult_82_SUMB_28__42_), .ZN(u5_mult_82_n2183) );
  NAND2_X1 u5_mult_82_U6399 ( .A1(u5_mult_82_ab_29__41_), .A2(
        u5_mult_82_SUMB_28__42_), .ZN(u5_mult_82_n2182) );
  NAND2_X1 u5_mult_82_U6398 ( .A1(u5_mult_82_ab_29__41_), .A2(
        u5_mult_82_CARRYB_28__41_), .ZN(u5_mult_82_n2181) );
  NAND3_X2 u5_mult_82_U6397 ( .A1(u5_mult_82_n2178), .A2(u5_mult_82_n2179), 
        .A3(u5_mult_82_n2180), .ZN(u5_mult_82_CARRYB_28__42_) );
  NAND2_X2 u5_mult_82_U6396 ( .A1(u5_mult_82_ab_28__42_), .A2(
        u5_mult_82_SUMB_27__43_), .ZN(u5_mult_82_n2180) );
  NAND2_X1 u5_mult_82_U6395 ( .A1(u5_mult_82_CARRYB_27__42_), .A2(
        u5_mult_82_ab_28__42_), .ZN(u5_mult_82_n2178) );
  XOR2_X2 u5_mult_82_U6394 ( .A(u5_mult_82_n2177), .B(u5_mult_82_SUMB_28__42_), 
        .Z(u5_mult_82_SUMB_29__41_) );
  XOR2_X2 u5_mult_82_U6393 ( .A(u5_mult_82_ab_29__41_), .B(
        u5_mult_82_CARRYB_28__41_), .Z(u5_mult_82_n2177) );
  XOR2_X2 u5_mult_82_U6392 ( .A(u5_mult_82_n2176), .B(u5_mult_82_SUMB_27__43_), 
        .Z(u5_mult_82_SUMB_28__42_) );
  XNOR2_X2 u5_mult_82_U6391 ( .A(u5_mult_82_n2175), .B(
        u5_mult_82_CARRYB_23__26_), .ZN(u5_mult_82_n5968) );
  NAND3_X2 u5_mult_82_U6390 ( .A1(u5_mult_82_n2906), .A2(u5_mult_82_n2905), 
        .A3(u5_mult_82_n2904), .ZN(u5_mult_82_n2174) );
  NAND2_X2 u5_mult_82_U6389 ( .A1(u5_mult_82_ab_23__11_), .A2(
        u5_mult_82_CARRYB_22__11_), .ZN(u5_mult_82_n4116) );
  NAND2_X2 u5_mult_82_U6388 ( .A1(u5_mult_82_ab_37__4_), .A2(u5_mult_82_n390), 
        .ZN(u5_mult_82_n2342) );
  NAND2_X2 u5_mult_82_U6387 ( .A1(u5_mult_82_ab_32__7_), .A2(
        u5_mult_82_CARRYB_31__7_), .ZN(u5_mult_82_n2853) );
  XNOR2_X2 u5_mult_82_U6386 ( .A(u5_mult_82_n2173), .B(
        u5_mult_82_CARRYB_48__13_), .ZN(u5_mult_82_n5755) );
  XNOR2_X2 u5_mult_82_U6385 ( .A(u5_mult_82_n2171), .B(u5_mult_82_SUMB_21__13_), .ZN(u5_mult_82_SUMB_22__12_) );
  NAND2_X1 u5_mult_82_U6384 ( .A1(u5_mult_82_ab_24__9_), .A2(
        u5_mult_82_SUMB_23__10_), .ZN(u5_mult_82_n3432) );
  NAND3_X2 u5_mult_82_U6383 ( .A1(u5_mult_82_n3435), .A2(u5_mult_82_n3436), 
        .A3(u5_mult_82_n3437), .ZN(u5_mult_82_CARRYB_25__9_) );
  NAND2_X2 u5_mult_82_U6382 ( .A1(u5_mult_82_n2112), .A2(
        u5_mult_82_SUMB_49__14_), .ZN(u5_mult_82_n5828) );
  NOR2_X1 u5_mult_82_U6381 ( .A1(u5_mult_82_net64453), .A2(u5_mult_82_n6630), 
        .ZN(u5_mult_82_ab_21__10_) );
  NOR2_X1 u5_mult_82_U6380 ( .A1(u5_mult_82_net64417), .A2(u5_mult_82_n6644), 
        .ZN(u5_mult_82_ab_24__8_) );
  NOR2_X1 u5_mult_82_U6379 ( .A1(u5_mult_82_net64381), .A2(u5_mult_82_n6658), 
        .ZN(u5_mult_82_ab_27__6_) );
  NOR2_X1 u5_mult_82_U6378 ( .A1(u5_mult_82_net64507), .A2(u5_mult_82_n6610), 
        .ZN(u5_mult_82_ab_18__13_) );
  NAND3_X2 u5_mult_82_U6377 ( .A1(u5_mult_82_n2168), .A2(u5_mult_82_n2169), 
        .A3(u5_mult_82_n2170), .ZN(u5_mult_82_CARRYB_21__10_) );
  NAND2_X1 u5_mult_82_U6376 ( .A1(u5_mult_82_ab_21__10_), .A2(
        u5_mult_82_CARRYB_20__10_), .ZN(u5_mult_82_n2170) );
  NAND2_X2 u5_mult_82_U6375 ( .A1(u5_mult_82_ab_21__10_), .A2(
        u5_mult_82_SUMB_20__11_), .ZN(u5_mult_82_n2169) );
  NAND2_X1 u5_mult_82_U6374 ( .A1(u5_mult_82_CARRYB_20__10_), .A2(
        u5_mult_82_SUMB_20__11_), .ZN(u5_mult_82_n2168) );
  XOR2_X2 u5_mult_82_U6373 ( .A(u5_mult_82_SUMB_20__11_), .B(u5_mult_82_n2167), 
        .Z(u5_mult_82_SUMB_21__10_) );
  XOR2_X2 u5_mult_82_U6372 ( .A(u5_mult_82_CARRYB_20__10_), .B(
        u5_mult_82_ab_21__10_), .Z(u5_mult_82_n2167) );
  NAND3_X2 u5_mult_82_U6371 ( .A1(u5_mult_82_n2164), .A2(u5_mult_82_n2165), 
        .A3(u5_mult_82_n2166), .ZN(u5_mult_82_CARRYB_24__8_) );
  NAND2_X1 u5_mult_82_U6370 ( .A1(u5_mult_82_ab_24__8_), .A2(
        u5_mult_82_CARRYB_23__8_), .ZN(u5_mult_82_n2166) );
  NAND2_X2 u5_mult_82_U6369 ( .A1(u5_mult_82_ab_24__8_), .A2(
        u5_mult_82_SUMB_23__9_), .ZN(u5_mult_82_n2165) );
  NAND2_X1 u5_mult_82_U6368 ( .A1(u5_mult_82_CARRYB_23__8_), .A2(
        u5_mult_82_SUMB_23__9_), .ZN(u5_mult_82_n2164) );
  XOR2_X2 u5_mult_82_U6367 ( .A(u5_mult_82_SUMB_23__9_), .B(u5_mult_82_n2163), 
        .Z(u5_mult_82_SUMB_24__8_) );
  XOR2_X2 u5_mult_82_U6366 ( .A(u5_mult_82_CARRYB_23__8_), .B(
        u5_mult_82_ab_24__8_), .Z(u5_mult_82_n2163) );
  NAND3_X2 u5_mult_82_U6365 ( .A1(u5_mult_82_n2160), .A2(u5_mult_82_n2161), 
        .A3(u5_mult_82_n2162), .ZN(u5_mult_82_CARRYB_27__6_) );
  NAND2_X1 u5_mult_82_U6364 ( .A1(u5_mult_82_ab_27__6_), .A2(
        u5_mult_82_CARRYB_26__6_), .ZN(u5_mult_82_n2162) );
  NAND2_X2 u5_mult_82_U6363 ( .A1(u5_mult_82_ab_27__6_), .A2(
        u5_mult_82_SUMB_26__7_), .ZN(u5_mult_82_n2161) );
  NAND2_X1 u5_mult_82_U6362 ( .A1(u5_mult_82_CARRYB_26__6_), .A2(
        u5_mult_82_SUMB_26__7_), .ZN(u5_mult_82_n2160) );
  XOR2_X2 u5_mult_82_U6361 ( .A(u5_mult_82_SUMB_26__7_), .B(u5_mult_82_n2159), 
        .Z(u5_mult_82_SUMB_27__6_) );
  XOR2_X2 u5_mult_82_U6360 ( .A(u5_mult_82_CARRYB_26__6_), .B(
        u5_mult_82_ab_27__6_), .Z(u5_mult_82_n2159) );
  NAND3_X2 u5_mult_82_U6359 ( .A1(u5_mult_82_n2156), .A2(u5_mult_82_n2157), 
        .A3(u5_mult_82_n2158), .ZN(u5_mult_82_CARRYB_18__13_) );
  NAND2_X1 u5_mult_82_U6358 ( .A1(u5_mult_82_ab_18__13_), .A2(
        u5_mult_82_SUMB_17__14_), .ZN(u5_mult_82_n2158) );
  NAND2_X1 u5_mult_82_U6357 ( .A1(u5_mult_82_ab_18__13_), .A2(
        u5_mult_82_CARRYB_17__13_), .ZN(u5_mult_82_n2157) );
  NAND2_X1 u5_mult_82_U6356 ( .A1(u5_mult_82_SUMB_17__14_), .A2(
        u5_mult_82_CARRYB_17__13_), .ZN(u5_mult_82_n2156) );
  NAND3_X4 u5_mult_82_U6355 ( .A1(u5_mult_82_n2959), .A2(u5_mult_82_n2960), 
        .A3(u5_mult_82_n2961), .ZN(u5_mult_82_CARRYB_47__32_) );
  NAND2_X1 u5_mult_82_U6354 ( .A1(u5_mult_82_SUMB_32__23_), .A2(
        u5_mult_82_ab_33__22_), .ZN(u5_mult_82_n5291) );
  NAND2_X4 u5_mult_82_U6353 ( .A1(u5_mult_82_n4690), .A2(u5_mult_82_n4691), 
        .ZN(u5_mult_82_n4693) );
  NAND2_X4 u5_mult_82_U6352 ( .A1(u5_mult_82_n4692), .A2(u5_mult_82_n4693), 
        .ZN(u5_mult_82_n6397) );
  NAND2_X2 u5_mult_82_U6351 ( .A1(u5_mult_82_CARRYB_23__26_), .A2(
        u5_mult_82_n1395), .ZN(u5_mult_82_n5971) );
  NAND2_X2 u5_mult_82_U6350 ( .A1(u5_mult_82_ab_30__22_), .A2(
        u5_mult_82_SUMB_29__23_), .ZN(u5_mult_82_n2898) );
  NOR2_X1 u5_mult_82_U6349 ( .A1(u5_mult_82_n6831), .A2(u5_mult_82_net65279), 
        .ZN(u5_mult_82_ab_47__39_) );
  NAND3_X2 u5_mult_82_U6348 ( .A1(u5_mult_82_n2153), .A2(u5_mult_82_n2154), 
        .A3(u5_mult_82_n2155), .ZN(u5_mult_82_CARRYB_47__39_) );
  NAND2_X1 u5_mult_82_U6347 ( .A1(u5_mult_82_ab_47__39_), .A2(
        u5_mult_82_CARRYB_46__39_), .ZN(u5_mult_82_n2155) );
  NAND2_X1 u5_mult_82_U6346 ( .A1(u5_mult_82_ab_47__39_), .A2(
        u5_mult_82_SUMB_46__40_), .ZN(u5_mult_82_n2154) );
  NAND2_X1 u5_mult_82_U6345 ( .A1(u5_mult_82_CARRYB_46__39_), .A2(
        u5_mult_82_SUMB_46__40_), .ZN(u5_mult_82_n2153) );
  XOR2_X2 u5_mult_82_U6344 ( .A(u5_mult_82_SUMB_46__40_), .B(u5_mult_82_n2152), 
        .Z(u5_mult_82_SUMB_47__39_) );
  XOR2_X2 u5_mult_82_U6343 ( .A(u5_mult_82_CARRYB_46__39_), .B(
        u5_mult_82_ab_47__39_), .Z(u5_mult_82_n2152) );
  NAND3_X2 u5_mult_82_U6342 ( .A1(u5_mult_82_n2149), .A2(u5_mult_82_n2150), 
        .A3(u5_mult_82_n2151), .ZN(u5_mult_82_CARRYB_49__37_) );
  NAND2_X1 u5_mult_82_U6341 ( .A1(u5_mult_82_CARRYB_48__37_), .A2(
        u5_mult_82_SUMB_48__38_), .ZN(u5_mult_82_n2151) );
  NAND2_X1 u5_mult_82_U6340 ( .A1(u5_mult_82_ab_49__37_), .A2(
        u5_mult_82_SUMB_48__38_), .ZN(u5_mult_82_n2150) );
  NAND2_X1 u5_mult_82_U6339 ( .A1(u5_mult_82_ab_49__37_), .A2(
        u5_mult_82_CARRYB_48__37_), .ZN(u5_mult_82_n2149) );
  NAND3_X2 u5_mult_82_U6338 ( .A1(u5_mult_82_n2146), .A2(u5_mult_82_n2147), 
        .A3(u5_mult_82_n2148), .ZN(u5_mult_82_CARRYB_48__38_) );
  NAND2_X1 u5_mult_82_U6337 ( .A1(u5_mult_82_CARRYB_47__38_), .A2(
        u5_mult_82_SUMB_47__39_), .ZN(u5_mult_82_n2148) );
  NAND2_X1 u5_mult_82_U6336 ( .A1(u5_mult_82_ab_48__38_), .A2(
        u5_mult_82_SUMB_47__39_), .ZN(u5_mult_82_n2147) );
  NAND2_X1 u5_mult_82_U6335 ( .A1(u5_mult_82_ab_48__38_), .A2(
        u5_mult_82_CARRYB_47__38_), .ZN(u5_mult_82_n2146) );
  XOR2_X2 u5_mult_82_U6334 ( .A(u5_mult_82_n2145), .B(u5_mult_82_SUMB_48__38_), 
        .Z(u5_mult_82_SUMB_49__37_) );
  XOR2_X2 u5_mult_82_U6333 ( .A(u5_mult_82_ab_49__37_), .B(
        u5_mult_82_CARRYB_48__37_), .Z(u5_mult_82_n2145) );
  XOR2_X2 u5_mult_82_U6332 ( .A(u5_mult_82_n2144), .B(u5_mult_82_SUMB_47__39_), 
        .Z(u5_mult_82_SUMB_48__38_) );
  XOR2_X2 u5_mult_82_U6331 ( .A(u5_mult_82_ab_48__38_), .B(
        u5_mult_82_CARRYB_47__38_), .Z(u5_mult_82_n2144) );
  NAND2_X2 u5_mult_82_U6330 ( .A1(u5_mult_82_ab_48__29_), .A2(u5_mult_82_n1826), .ZN(u5_mult_82_n3758) );
  XNOR2_X2 u5_mult_82_U6329 ( .A(u5_mult_82_ab_47__14_), .B(
        u5_mult_82_CARRYB_46__14_), .ZN(u5_mult_82_n2143) );
  XNOR2_X2 u5_mult_82_U6328 ( .A(u5_mult_82_n2143), .B(u5_mult_82_n1693), .ZN(
        u5_mult_82_SUMB_47__14_) );
  XNOR2_X2 u5_mult_82_U6327 ( .A(u5_mult_82_CARRYB_45__29_), .B(
        u5_mult_82_ab_46__29_), .ZN(u5_mult_82_n2142) );
  XNOR2_X2 u5_mult_82_U6326 ( .A(u5_mult_82_SUMB_45__30_), .B(u5_mult_82_n2142), .ZN(u5_mult_82_SUMB_46__29_) );
  XNOR2_X2 u5_mult_82_U6325 ( .A(u5_mult_82_CARRYB_18__22_), .B(
        u5_mult_82_ab_19__22_), .ZN(u5_mult_82_n2141) );
  XNOR2_X2 u5_mult_82_U6324 ( .A(u5_mult_82_n2141), .B(u5_mult_82_SUMB_18__23_), .ZN(u5_mult_82_SUMB_19__22_) );
  XNOR2_X2 u5_mult_82_U6323 ( .A(u5_mult_82_SUMB_17__51_), .B(
        u5_mult_82_ab_18__50_), .ZN(u5_mult_82_n2140) );
  XNOR2_X2 u5_mult_82_U6322 ( .A(u5_mult_82_CARRYB_17__50_), .B(
        u5_mult_82_n2140), .ZN(u5_mult_82_SUMB_18__50_) );
  NAND2_X2 u5_mult_82_U6321 ( .A1(u5_mult_82_CARRYB_23__27_), .A2(
        u5_mult_82_ab_24__27_), .ZN(u5_mult_82_n6141) );
  NAND2_X1 u5_mult_82_U6320 ( .A1(u5_mult_82_ab_33__23_), .A2(
        u5_mult_82_CARRYB_32__23_), .ZN(u5_mult_82_n4008) );
  NAND2_X1 u5_mult_82_U6319 ( .A1(u5_mult_82_ab_38__21_), .A2(
        u5_mult_82_CARRYB_37__21_), .ZN(u5_mult_82_n4002) );
  NAND2_X2 u5_mult_82_U6318 ( .A1(u5_mult_82_n455), .A2(
        u5_mult_82_CARRYB_42__17_), .ZN(u5_mult_82_n4282) );
  XNOR2_X2 u5_mult_82_U6317 ( .A(u5_mult_82_ab_19__29_), .B(
        u5_mult_82_CARRYB_18__29_), .ZN(u5_mult_82_n2139) );
  XNOR2_X2 u5_mult_82_U6316 ( .A(u5_mult_82_n2139), .B(u5_mult_82_SUMB_18__30_), .ZN(u5_mult_82_SUMB_19__29_) );
  NAND2_X2 u5_mult_82_U6315 ( .A1(u5_mult_82_ab_48__35_), .A2(u5_mult_82_n1503), .ZN(u5_mult_82_n3092) );
  XNOR2_X1 u5_mult_82_U6314 ( .A(u5_mult_82_ab_12__50_), .B(
        u5_mult_82_SUMB_11__51_), .ZN(u5_mult_82_n2138) );
  XNOR2_X2 u5_mult_82_U6313 ( .A(u5_mult_82_CARRYB_48__5_), .B(
        u5_mult_82_ab_49__5_), .ZN(u5_mult_82_n2137) );
  XNOR2_X2 u5_mult_82_U6312 ( .A(u5_mult_82_n2137), .B(u5_mult_82_SUMB_48__6_), 
        .ZN(u5_mult_82_SUMB_49__5_) );
  NAND2_X2 u5_mult_82_U6311 ( .A1(u5_mult_82_CARRYB_44__4_), .A2(
        u5_mult_82_SUMB_44__5_), .ZN(u5_mult_82_n6024) );
  XNOR2_X2 u5_mult_82_U6310 ( .A(u5_mult_82_n2136), .B(
        u5_mult_82_CARRYB_45__7_), .ZN(u5_mult_82_SUMB_46__7_) );
  NAND2_X1 u5_mult_82_U6309 ( .A1(u5_mult_82_n1866), .A2(u5_mult_82_n4101), 
        .ZN(u5_mult_82_n4890) );
  NAND3_X4 u5_mult_82_U6308 ( .A1(u5_mult_82_n4658), .A2(u5_mult_82_n4657), 
        .A3(u5_mult_82_n4656), .ZN(u5_mult_82_CARRYB_45__6_) );
  XNOR2_X2 u5_mult_82_U6307 ( .A(u5_mult_82_ab_51__34_), .B(
        u5_mult_82_CARRYB_50__34_), .ZN(u5_mult_82_n2135) );
  NAND2_X1 u5_mult_82_U6306 ( .A1(u5_mult_82_CARRYB_27__37_), .A2(
        u5_mult_82_SUMB_27__38_), .ZN(u5_mult_82_n5666) );
  NAND3_X4 u5_mult_82_U6305 ( .A1(u5_mult_82_n3613), .A2(u5_mult_82_net83292), 
        .A3(u5_mult_82_net83293), .ZN(u5_mult_82_CARRYB_32__17_) );
  NAND2_X2 u5_mult_82_U6304 ( .A1(u5_mult_82_n5248), .A2(
        u5_mult_82_SUMB_18__45_), .ZN(u5_mult_82_n5877) );
  NAND2_X2 u5_mult_82_U6303 ( .A1(u5_mult_82_CARRYB_39__0_), .A2(
        u5_mult_82_SUMB_39__1_), .ZN(u5_mult_82_n4849) );
  XOR2_X1 u5_mult_82_U6302 ( .A(u5_mult_82_SUMB_39__1_), .B(u5_mult_82_n4848), 
        .Z(u5_N40) );
  XNOR2_X2 u5_mult_82_U6301 ( .A(u5_mult_82_CARRYB_24__32_), .B(
        u5_mult_82_ab_25__32_), .ZN(u5_mult_82_n2134) );
  XNOR2_X2 u5_mult_82_U6300 ( .A(u5_mult_82_n2134), .B(u5_mult_82_SUMB_24__33_), .ZN(u5_mult_82_SUMB_25__32_) );
  NAND3_X2 u5_mult_82_U6299 ( .A1(u5_mult_82_n6365), .A2(u5_mult_82_n6366), 
        .A3(u5_mult_82_n6367), .ZN(u5_mult_82_CARRYB_32__25_) );
  NAND3_X2 u5_mult_82_U6298 ( .A1(u5_mult_82_n6171), .A2(u5_mult_82_n6170), 
        .A3(u5_mult_82_n6169), .ZN(u5_mult_82_CARRYB_47__5_) );
  NAND3_X2 u5_mult_82_U6297 ( .A1(u5_mult_82_n4986), .A2(u5_mult_82_n4987), 
        .A3(u5_mult_82_n4988), .ZN(u5_mult_82_CARRYB_21__35_) );
  NAND2_X2 u5_mult_82_U6296 ( .A1(u5_mult_82_ab_37__6_), .A2(
        u5_mult_82_SUMB_36__7_), .ZN(u5_mult_82_n3198) );
  XNOR2_X2 u5_mult_82_U6295 ( .A(u5_mult_82_n2131), .B(
        u5_mult_82_CARRYB_24__14_), .ZN(u5_mult_82_n4828) );
  NAND3_X4 u5_mult_82_U6294 ( .A1(u5_mult_82_n4941), .A2(u5_mult_82_n4942), 
        .A3(u5_mult_82_n4943), .ZN(u5_mult_82_CARRYB_20__40_) );
  XNOR2_X2 u5_mult_82_U6293 ( .A(u5_mult_82_n433), .B(u5_mult_82_n3693), .ZN(
        u5_mult_82_SUMB_24__32_) );
  NAND2_X1 u5_mult_82_U6292 ( .A1(u5_mult_82_CARRYB_36__3_), .A2(
        u5_mult_82_SUMB_36__4_), .ZN(u5_mult_82_n4682) );
  NAND2_X1 u5_mult_82_U6291 ( .A1(u5_mult_82_ab_37__3_), .A2(
        u5_mult_82_CARRYB_36__3_), .ZN(u5_mult_82_n4680) );
  XOR2_X2 u5_mult_82_U6290 ( .A(u5_mult_82_ab_37__3_), .B(
        u5_mult_82_CARRYB_36__3_), .Z(u5_mult_82_n4679) );
  XNOR2_X2 u5_mult_82_U6289 ( .A(u5_mult_82_ab_11__29_), .B(
        u5_mult_82_CARRYB_10__29_), .ZN(u5_mult_82_n2130) );
  XNOR2_X2 u5_mult_82_U6288 ( .A(u5_mult_82_n2130), .B(u5_mult_82_SUMB_10__30_), .ZN(u5_mult_82_SUMB_11__29_) );
  XNOR2_X2 u5_mult_82_U6287 ( .A(u5_mult_82_n2129), .B(u5_mult_82_SUMB_15__21_), .ZN(u5_mult_82_SUMB_16__20_) );
  NAND3_X4 u5_mult_82_U6286 ( .A1(u5_mult_82_n4597), .A2(u5_mult_82_n4596), 
        .A3(u5_mult_82_n4595), .ZN(u5_mult_82_CARRYB_45__5_) );
  NAND3_X4 u5_mult_82_U6285 ( .A1(u5_mult_82_n6003), .A2(u5_mult_82_n6004), 
        .A3(u5_mult_82_n6005), .ZN(u5_mult_82_CARRYB_41__7_) );
  XNOR2_X2 u5_mult_82_U6284 ( .A(u5_mult_82_CARRYB_35__25_), .B(
        u5_mult_82_ab_36__25_), .ZN(u5_mult_82_n2128) );
  XNOR2_X2 u5_mult_82_U6283 ( .A(u5_mult_82_SUMB_35__26_), .B(u5_mult_82_n2128), .ZN(u5_mult_82_SUMB_36__25_) );
  INV_X2 u5_mult_82_U6282 ( .A(u5_mult_82_CARRYB_42__18_), .ZN(
        u5_mult_82_n3138) );
  NAND2_X1 u5_mult_82_U6281 ( .A1(u5_mult_82_CARRYB_37__8_), .A2(
        u5_mult_82_SUMB_37__9_), .ZN(u5_mult_82_n2986) );
  NAND2_X1 u5_mult_82_U6280 ( .A1(u5_mult_82_ab_38__8_), .A2(
        u5_mult_82_CARRYB_37__8_), .ZN(u5_mult_82_n2984) );
  XNOR2_X2 u5_mult_82_U6279 ( .A(u5_mult_82_n2127), .B(
        u5_mult_82_CARRYB_47__31_), .ZN(u5_mult_82_n2958) );
  NAND2_X2 u5_mult_82_U6278 ( .A1(u5_mult_82_CARRYB_45__35_), .A2(
        u5_mult_82_n1570), .ZN(u5_mult_82_n2917) );
  NAND2_X2 u5_mult_82_U6277 ( .A1(u5_mult_82_SUMB_42__2_), .A2(
        u5_mult_82_n1652), .ZN(u5_mult_82_n2544) );
  XOR2_X2 u5_mult_82_U6276 ( .A(u5_mult_82_ab_47__21_), .B(u5_mult_82_n702), 
        .Z(u5_mult_82_n5744) );
  XNOR2_X2 u5_mult_82_U6275 ( .A(u5_mult_82_ab_41__5_), .B(
        u5_mult_82_CARRYB_40__5_), .ZN(u5_mult_82_n2126) );
  XNOR2_X2 u5_mult_82_U6274 ( .A(u5_mult_82_n2126), .B(u5_mult_82_SUMB_40__6_), 
        .ZN(u5_mult_82_SUMB_41__5_) );
  NAND2_X2 u5_mult_82_U6273 ( .A1(u5_mult_82_ab_19__28_), .A2(
        u5_mult_82_CARRYB_18__28_), .ZN(u5_mult_82_n5429) );
  XNOR2_X1 u5_mult_82_U6272 ( .A(u5_mult_82_SUMB_8__50_), .B(
        u5_mult_82_ab_9__49_), .ZN(u5_mult_82_n2125) );
  XNOR2_X2 u5_mult_82_U6271 ( .A(u5_mult_82_CARRYB_8__49_), .B(
        u5_mult_82_n2125), .ZN(u5_mult_82_SUMB_9__49_) );
  XNOR2_X2 u5_mult_82_U6270 ( .A(u5_mult_82_CARRYB_36__6_), .B(
        u5_mult_82_n2123), .ZN(u5_mult_82_SUMB_37__6_) );
  XNOR2_X2 u5_mult_82_U6269 ( .A(u5_mult_82_n2122), .B(u5_mult_82_SUMB_16__27_), .ZN(u5_mult_82_SUMB_17__26_) );
  XNOR2_X2 u5_mult_82_U6268 ( .A(u5_mult_82_ab_24__41_), .B(
        u5_mult_82_CARRYB_23__41_), .ZN(u5_mult_82_n2121) );
  XNOR2_X2 u5_mult_82_U6267 ( .A(u5_mult_82_n2121), .B(u5_mult_82_n1691), .ZN(
        u5_mult_82_SUMB_24__41_) );
  XNOR2_X2 u5_mult_82_U6266 ( .A(u5_mult_82_SUMB_17__14_), .B(
        u5_mult_82_ab_18__13_), .ZN(u5_mult_82_n2120) );
  XNOR2_X2 u5_mult_82_U6265 ( .A(u5_mult_82_n630), .B(u5_mult_82_n2120), .ZN(
        u5_mult_82_SUMB_18__13_) );
  XNOR2_X2 u5_mult_82_U6264 ( .A(u5_mult_82_n303), .B(u5_mult_82_ab_18__29_), 
        .ZN(u5_mult_82_n2119) );
  XNOR2_X2 u5_mult_82_U6263 ( .A(u5_mult_82_n2119), .B(u5_mult_82_n1680), .ZN(
        u5_mult_82_SUMB_18__29_) );
  NAND2_X2 u5_mult_82_U6262 ( .A1(u5_mult_82_ab_42__2_), .A2(
        u5_mult_82_CARRYB_41__2_), .ZN(u5_mult_82_n5633) );
  XNOR2_X2 u5_mult_82_U6261 ( .A(u5_mult_82_CARRYB_33__11_), .B(
        u5_mult_82_ab_34__11_), .ZN(u5_mult_82_n2118) );
  NAND2_X1 u5_mult_82_U6260 ( .A1(u5_mult_82_SUMB_41__18_), .A2(
        u5_mult_82_CARRYB_41__17_), .ZN(u5_mult_82_n5066) );
  XNOR2_X2 u5_mult_82_U6259 ( .A(u5_mult_82_ab_16__44_), .B(
        u5_mult_82_CARRYB_15__44_), .ZN(u5_mult_82_n2117) );
  XNOR2_X2 u5_mult_82_U6258 ( .A(u5_mult_82_n2117), .B(u5_mult_82_SUMB_15__45_), .ZN(u5_mult_82_SUMB_16__44_) );
  NAND3_X4 u5_mult_82_U6257 ( .A1(u5_mult_82_n5759), .A2(u5_mult_82_n5760), 
        .A3(u5_mult_82_n5761), .ZN(u5_mult_82_CARRYB_50__12_) );
  NOR2_X1 u5_mult_82_U6256 ( .A1(u5_mult_82_net64487), .A2(u5_mult_82_net65189), .ZN(u5_mult_82_ab_51__12_) );
  NAND3_X2 u5_mult_82_U6255 ( .A1(u5_mult_82_n2114), .A2(u5_mult_82_n2115), 
        .A3(u5_mult_82_n2116), .ZN(u5_mult_82_CARRYB_51__12_) );
  NAND2_X1 u5_mult_82_U6254 ( .A1(u5_mult_82_ab_51__12_), .A2(
        u5_mult_82_CARRYB_50__12_), .ZN(u5_mult_82_n2116) );
  NAND2_X2 u5_mult_82_U6253 ( .A1(u5_mult_82_ab_51__12_), .A2(
        u5_mult_82_SUMB_50__13_), .ZN(u5_mult_82_n2115) );
  NAND2_X1 u5_mult_82_U6252 ( .A1(u5_mult_82_SUMB_50__13_), .A2(
        u5_mult_82_CARRYB_50__12_), .ZN(u5_mult_82_n2114) );
  XOR2_X2 u5_mult_82_U6251 ( .A(u5_mult_82_SUMB_50__13_), .B(u5_mult_82_n2113), 
        .Z(u5_mult_82_SUMB_51__12_) );
  XOR2_X2 u5_mult_82_U6250 ( .A(u5_mult_82_CARRYB_50__12_), .B(
        u5_mult_82_ab_51__12_), .Z(u5_mult_82_n2113) );
  NAND3_X2 u5_mult_82_U6249 ( .A1(u5_mult_82_n3199), .A2(u5_mult_82_n3200), 
        .A3(u5_mult_82_n3201), .ZN(u5_mult_82_CARRYB_39__5_) );
  NAND2_X2 u5_mult_82_U6248 ( .A1(u5_mult_82_n5507), .A2(
        u5_mult_82_SUMB_22__35_), .ZN(u5_mult_82_n6377) );
  NAND2_X2 u5_mult_82_U6247 ( .A1(u5_mult_82_CARRYB_13__42_), .A2(
        u5_mult_82_n1794), .ZN(u5_mult_82_n5645) );
  NAND2_X2 u5_mult_82_U6246 ( .A1(u5_mult_82_ab_42__3_), .A2(
        u5_mult_82_CARRYB_41__3_), .ZN(u5_mult_82_n4963) );
  NAND2_X2 u5_mult_82_U6245 ( .A1(u5_mult_82_CARRYB_47__29_), .A2(
        u5_mult_82_n1826), .ZN(u5_mult_82_n3757) );
  NAND2_X2 u5_mult_82_U6244 ( .A1(u5_mult_82_CARRYB_42__0_), .A2(
        u5_mult_82_ab_43__0_), .ZN(u5_mult_82_n4839) );
  NAND2_X2 u5_mult_82_U6243 ( .A1(u5_mult_82_ab_20__40_), .A2(
        u5_mult_82_CARRYB_19__40_), .ZN(u5_mult_82_n4941) );
  NAND3_X2 u5_mult_82_U6242 ( .A1(u5_mult_82_n3260), .A2(u5_mult_82_n3261), 
        .A3(u5_mult_82_n3262), .ZN(u5_mult_82_CARRYB_48__30_) );
  XNOR2_X1 u5_mult_82_U6241 ( .A(u5_mult_82_n3496), .B(u5_mult_82_SUMB_25__46_), .ZN(u5_mult_82_SUMB_26__45_) );
  NAND3_X2 u5_mult_82_U6240 ( .A1(u5_mult_82_n4602), .A2(u5_mult_82_n4603), 
        .A3(u5_mult_82_n4604), .ZN(u5_mult_82_CARRYB_20__43_) );
  XNOR2_X2 u5_mult_82_U6239 ( .A(u5_mult_82_n2111), .B(u5_mult_82_SUMB_5__44_), 
        .ZN(u5_mult_82_SUMB_6__43_) );
  NAND2_X1 u5_mult_82_U6238 ( .A1(u5_mult_82_CARRYB_48__31_), .A2(
        u5_mult_82_SUMB_48__32_), .ZN(u5_mult_82_n2942) );
  NOR2_X1 u5_mult_82_U6237 ( .A1(u5_mult_82_net64913), .A2(u5_mult_82_n6734), 
        .ZN(u5_mult_82_ab_44__35_) );
  NOR2_X1 u5_mult_82_U6236 ( .A1(u5_mult_82_n6811), .A2(u5_mult_82_n6664), 
        .ZN(u5_mult_82_ab_28__43_) );
  NAND3_X4 u5_mult_82_U6235 ( .A1(u5_mult_82_n5592), .A2(u5_mult_82_n5593), 
        .A3(u5_mult_82_n5594), .ZN(u5_mult_82_CARRYB_26__43_) );
  NOR2_X1 u5_mult_82_U6234 ( .A1(u5_mult_82_n6812), .A2(u5_mult_82_n6655), 
        .ZN(u5_mult_82_ab_27__43_) );
  NOR2_X1 u5_mult_82_U6233 ( .A1(u5_mult_82_n6792), .A2(u5_mult_82_n6636), 
        .ZN(u5_mult_82_ab_22__46_) );
  NAND3_X4 u5_mult_82_U6232 ( .A1(u5_mult_82_n2108), .A2(u5_mult_82_n2109), 
        .A3(u5_mult_82_n2110), .ZN(u5_mult_82_CARRYB_44__35_) );
  NAND2_X1 u5_mult_82_U6231 ( .A1(u5_mult_82_ab_44__35_), .A2(
        u5_mult_82_CARRYB_43__35_), .ZN(u5_mult_82_n2110) );
  NAND2_X2 u5_mult_82_U6230 ( .A1(u5_mult_82_SUMB_43__36_), .A2(
        u5_mult_82_ab_44__35_), .ZN(u5_mult_82_n2109) );
  NAND2_X2 u5_mult_82_U6229 ( .A1(u5_mult_82_CARRYB_43__35_), .A2(
        u5_mult_82_SUMB_43__36_), .ZN(u5_mult_82_n2108) );
  XOR2_X2 u5_mult_82_U6228 ( .A(u5_mult_82_SUMB_43__36_), .B(u5_mult_82_n2107), 
        .Z(u5_mult_82_SUMB_44__35_) );
  XOR2_X2 u5_mult_82_U6227 ( .A(u5_mult_82_CARRYB_43__35_), .B(
        u5_mult_82_ab_44__35_), .Z(u5_mult_82_n2107) );
  NAND3_X2 u5_mult_82_U6226 ( .A1(u5_mult_82_n2104), .A2(u5_mult_82_n2105), 
        .A3(u5_mult_82_n2106), .ZN(u5_mult_82_CARRYB_28__43_) );
  NAND2_X1 u5_mult_82_U6225 ( .A1(u5_mult_82_ab_28__43_), .A2(
        u5_mult_82_CARRYB_27__43_), .ZN(u5_mult_82_n2106) );
  NAND2_X2 u5_mult_82_U6224 ( .A1(u5_mult_82_ab_28__43_), .A2(
        u5_mult_82_SUMB_27__44_), .ZN(u5_mult_82_n2105) );
  NAND2_X2 u5_mult_82_U6223 ( .A1(u5_mult_82_CARRYB_27__43_), .A2(
        u5_mult_82_SUMB_27__44_), .ZN(u5_mult_82_n2104) );
  XOR2_X2 u5_mult_82_U6222 ( .A(u5_mult_82_SUMB_27__44_), .B(u5_mult_82_n2103), 
        .Z(u5_mult_82_SUMB_28__43_) );
  XOR2_X2 u5_mult_82_U6221 ( .A(u5_mult_82_CARRYB_27__43_), .B(
        u5_mult_82_ab_28__43_), .Z(u5_mult_82_n2103) );
  NAND3_X2 u5_mult_82_U6220 ( .A1(u5_mult_82_n2100), .A2(u5_mult_82_n2101), 
        .A3(u5_mult_82_n2102), .ZN(u5_mult_82_CARRYB_27__43_) );
  NAND2_X1 u5_mult_82_U6219 ( .A1(u5_mult_82_ab_27__43_), .A2(
        u5_mult_82_CARRYB_26__43_), .ZN(u5_mult_82_n2102) );
  NAND2_X2 u5_mult_82_U6218 ( .A1(u5_mult_82_ab_27__43_), .A2(
        u5_mult_82_SUMB_26__44_), .ZN(u5_mult_82_n2101) );
  NAND2_X1 u5_mult_82_U6217 ( .A1(u5_mult_82_CARRYB_26__43_), .A2(
        u5_mult_82_SUMB_26__44_), .ZN(u5_mult_82_n2100) );
  XOR2_X2 u5_mult_82_U6216 ( .A(u5_mult_82_SUMB_26__44_), .B(u5_mult_82_n2099), 
        .Z(u5_mult_82_SUMB_27__43_) );
  XOR2_X2 u5_mult_82_U6215 ( .A(u5_mult_82_CARRYB_26__43_), .B(
        u5_mult_82_ab_27__43_), .Z(u5_mult_82_n2099) );
  NAND3_X2 u5_mult_82_U6214 ( .A1(u5_mult_82_n2096), .A2(u5_mult_82_n2097), 
        .A3(u5_mult_82_n2098), .ZN(u5_mult_82_CARRYB_14__51_) );
  NAND2_X2 u5_mult_82_U6213 ( .A1(u5_mult_82_ab_13__52_), .A2(
        u5_mult_82_CARRYB_13__51_), .ZN(u5_mult_82_n2098) );
  NAND2_X2 u5_mult_82_U6212 ( .A1(u5_mult_82_ab_14__51_), .A2(
        u5_mult_82_CARRYB_13__51_), .ZN(u5_mult_82_n2097) );
  NAND2_X2 u5_mult_82_U6211 ( .A1(u5_mult_82_ab_14__51_), .A2(
        u5_mult_82_ab_13__52_), .ZN(u5_mult_82_n2096) );
  XOR2_X2 u5_mult_82_U6210 ( .A(u5_mult_82_ab_14__51_), .B(
        u5_mult_82_ab_13__52_), .Z(u5_mult_82_n2095) );
  NAND3_X2 u5_mult_82_U6209 ( .A1(u5_mult_82_n2092), .A2(u5_mult_82_n2093), 
        .A3(u5_mult_82_n2094), .ZN(u5_mult_82_CARRYB_13__51_) );
  NAND2_X1 u5_mult_82_U6208 ( .A1(u5_mult_82_CARRYB_12__51_), .A2(
        u5_mult_82_ab_12__52_), .ZN(u5_mult_82_n2094) );
  NAND2_X2 u5_mult_82_U6207 ( .A1(u5_mult_82_ab_13__51_), .A2(
        u5_mult_82_ab_12__52_), .ZN(u5_mult_82_n2093) );
  NAND2_X1 u5_mult_82_U6206 ( .A1(u5_mult_82_ab_13__51_), .A2(
        u5_mult_82_CARRYB_12__51_), .ZN(u5_mult_82_n2092) );
  XOR2_X2 u5_mult_82_U6205 ( .A(u5_mult_82_n2091), .B(u5_mult_82_ab_12__52_), 
        .Z(u5_mult_82_SUMB_13__51_) );
  XOR2_X2 u5_mult_82_U6204 ( .A(u5_mult_82_ab_13__51_), .B(
        u5_mult_82_CARRYB_12__51_), .Z(u5_mult_82_n2091) );
  NAND3_X2 u5_mult_82_U6203 ( .A1(u5_mult_82_n2088), .A2(u5_mult_82_n2089), 
        .A3(u5_mult_82_n2090), .ZN(u5_mult_82_CARRYB_10__51_) );
  NAND2_X2 u5_mult_82_U6202 ( .A1(u5_mult_82_ab_9__52_), .A2(
        u5_mult_82_CARRYB_9__51_), .ZN(u5_mult_82_n2090) );
  NAND2_X2 u5_mult_82_U6201 ( .A1(u5_mult_82_ab_10__51_), .A2(
        u5_mult_82_CARRYB_9__51_), .ZN(u5_mult_82_n2089) );
  NAND2_X2 u5_mult_82_U6200 ( .A1(u5_mult_82_ab_10__51_), .A2(
        u5_mult_82_ab_9__52_), .ZN(u5_mult_82_n2088) );
  XOR2_X2 u5_mult_82_U6199 ( .A(u5_mult_82_ab_10__51_), .B(
        u5_mult_82_ab_9__52_), .Z(u5_mult_82_n2087) );
  NAND3_X2 u5_mult_82_U6198 ( .A1(u5_mult_82_n2084), .A2(u5_mult_82_n2085), 
        .A3(u5_mult_82_n2086), .ZN(u5_mult_82_CARRYB_9__51_) );
  NAND2_X2 u5_mult_82_U6197 ( .A1(u5_mult_82_ab_9__51_), .A2(
        u5_mult_82_ab_8__52_), .ZN(u5_mult_82_n2085) );
  XOR2_X2 u5_mult_82_U6196 ( .A(u5_mult_82_n2083), .B(u5_mult_82_ab_8__52_), 
        .Z(u5_mult_82_SUMB_9__51_) );
  NAND3_X2 u5_mult_82_U6195 ( .A1(u5_mult_82_n2080), .A2(u5_mult_82_n2081), 
        .A3(u5_mult_82_n2082), .ZN(u5_mult_82_CARRYB_22__46_) );
  NAND2_X1 u5_mult_82_U6194 ( .A1(u5_mult_82_ab_22__46_), .A2(
        u5_mult_82_CARRYB_21__46_), .ZN(u5_mult_82_n2082) );
  NAND2_X2 u5_mult_82_U6193 ( .A1(u5_mult_82_ab_22__46_), .A2(
        u5_mult_82_SUMB_21__47_), .ZN(u5_mult_82_n2081) );
  NAND2_X1 u5_mult_82_U6192 ( .A1(u5_mult_82_CARRYB_21__46_), .A2(
        u5_mult_82_SUMB_21__47_), .ZN(u5_mult_82_n2080) );
  XOR2_X2 u5_mult_82_U6191 ( .A(u5_mult_82_SUMB_21__47_), .B(u5_mult_82_n2079), 
        .Z(u5_mult_82_SUMB_22__46_) );
  XOR2_X2 u5_mult_82_U6190 ( .A(u5_mult_82_CARRYB_21__46_), .B(
        u5_mult_82_ab_22__46_), .Z(u5_mult_82_n2079) );
  INV_X1 u5_mult_82_U6189 ( .A(u5_mult_82_SUMB_47__34_), .ZN(u5_mult_82_n2076)
         );
  NAND2_X2 u5_mult_82_U6188 ( .A1(u5_mult_82_n2077), .A2(u5_mult_82_n2078), 
        .ZN(u5_mult_82_SUMB_48__33_) );
  NAND2_X2 u5_mult_82_U6187 ( .A1(u5_mult_82_n2075), .A2(u5_mult_82_n2076), 
        .ZN(u5_mult_82_n2078) );
  NAND2_X2 u5_mult_82_U6186 ( .A1(u5_mult_82_SUMB_47__15_), .A2(
        u5_mult_82_CARRYB_47__14_), .ZN(u5_mult_82_n5775) );
  NAND2_X2 u5_mult_82_U6185 ( .A1(u5_mult_82_CARRYB_33__9_), .A2(
        u5_mult_82_SUMB_33__10_), .ZN(u5_mult_82_n4156) );
  XOR2_X2 u5_mult_82_U6184 ( .A(u5_mult_82_n1834), .B(u5_mult_82_n6385), .Z(
        u5_mult_82_SUMB_5__51_) );
  NAND3_X2 u5_mult_82_U6183 ( .A1(u5_mult_82_n5840), .A2(u5_mult_82_n5841), 
        .A3(u5_mult_82_n5842), .ZN(u5_mult_82_CARRYB_19__43_) );
  XNOR2_X2 u5_mult_82_U6182 ( .A(u5_mult_82_n5960), .B(u5_mult_82_n35), .ZN(
        u5_mult_82_SUMB_47__5_) );
  NAND2_X2 u5_mult_82_U6181 ( .A1(u5_mult_82_ab_34__9_), .A2(
        u5_mult_82_SUMB_33__10_), .ZN(u5_mult_82_n4155) );
  XNOR2_X2 u5_mult_82_U6180 ( .A(u5_mult_82_n2074), .B(u5_mult_82_SUMB_22__12_), .ZN(u5_mult_82_SUMB_23__11_) );
  XNOR2_X2 u5_mult_82_U6179 ( .A(u5_mult_82_ab_27__29_), .B(
        u5_mult_82_CARRYB_26__29_), .ZN(u5_mult_82_n2073) );
  XNOR2_X2 u5_mult_82_U6178 ( .A(u5_mult_82_n2073), .B(u5_mult_82_SUMB_26__30_), .ZN(u5_mult_82_SUMB_27__29_) );
  NAND2_X1 u5_mult_82_U6177 ( .A1(u5_mult_82_CARRYB_24__39_), .A2(
        u5_mult_82_SUMB_24__40_), .ZN(u5_mult_82_n3036) );
  NAND2_X2 u5_mult_82_U6176 ( .A1(u5_mult_82_ab_26__38_), .A2(
        u5_mult_82_SUMB_25__39_), .ZN(u5_mult_82_n5671) );
  NAND2_X1 u5_mult_82_U6175 ( .A1(u5_mult_82_ab_28__37_), .A2(
        u5_mult_82_SUMB_27__38_), .ZN(u5_mult_82_n5665) );
  XNOR2_X2 u5_mult_82_U6174 ( .A(u5_mult_82_ab_20__23_), .B(
        u5_mult_82_CARRYB_19__23_), .ZN(u5_mult_82_n2072) );
  XNOR2_X2 u5_mult_82_U6173 ( .A(u5_mult_82_n2072), .B(u5_mult_82_SUMB_19__24_), .ZN(u5_mult_82_SUMB_20__23_) );
  XNOR2_X2 u5_mult_82_U6172 ( .A(u5_mult_82_CARRYB_6__27_), .B(
        u5_mult_82_ab_7__27_), .ZN(u5_mult_82_n2071) );
  XNOR2_X2 u5_mult_82_U6171 ( .A(u5_mult_82_n2071), .B(u5_mult_82_SUMB_6__28_), 
        .ZN(u5_mult_82_SUMB_7__27_) );
  NAND3_X4 u5_mult_82_U6170 ( .A1(u5_mult_82_n4537), .A2(u5_mult_82_n4538), 
        .A3(u5_mult_82_n4539), .ZN(u5_mult_82_CARRYB_30__29_) );
  XOR2_X2 u5_mult_82_U6169 ( .A(u5_mult_82_CARRYB_43__23_), .B(
        u5_mult_82_ab_44__23_), .Z(u5_mult_82_n3915) );
  NAND2_X2 u5_mult_82_U6168 ( .A1(u5_mult_82_n14), .A2(u5_mult_82_SUMB_42__1_), 
        .ZN(u5_mult_82_n4837) );
  NAND3_X4 u5_mult_82_U6167 ( .A1(u5_mult_82_net84193), .A2(
        u5_mult_82_net84194), .A3(u5_mult_82_n3057), .ZN(
        u5_mult_82_CARRYB_20__25_) );
  NAND2_X1 u5_mult_82_U6166 ( .A1(u5_mult_82_SUMB_34__28_), .A2(
        u5_mult_82_CARRYB_34__27_), .ZN(u5_mult_82_n2806) );
  XNOR2_X2 u5_mult_82_U6165 ( .A(u5_mult_82_ab_19__28_), .B(
        u5_mult_82_CARRYB_18__28_), .ZN(u5_mult_82_n2070) );
  XNOR2_X2 u5_mult_82_U6164 ( .A(u5_mult_82_n2070), .B(u5_mult_82_n32), .ZN(
        u5_mult_82_SUMB_19__28_) );
  NAND2_X2 u5_mult_82_U6163 ( .A1(u5_mult_82_ab_24__37_), .A2(
        u5_mult_82_SUMB_23__38_), .ZN(u5_mult_82_n5560) );
  XNOR2_X2 u5_mult_82_U6162 ( .A(u5_mult_82_n2124), .B(u5_mult_82_ab_1__51_), 
        .ZN(u5_mult_82_n6512) );
  XOR2_X2 u5_mult_82_U6161 ( .A(u5_mult_82_n2667), .B(u5_mult_82_n1637), .Z(
        u5_mult_82_SUMB_40__3_) );
  NAND3_X2 u5_mult_82_U6160 ( .A1(u5_mult_82_n1033), .A2(u5_mult_82_n2671), 
        .A3(u5_mult_82_n2672), .ZN(u5_mult_82_CARRYB_41__2_) );
  NAND2_X1 u5_mult_82_U6159 ( .A1(u5_mult_82_CARRYB_24__7_), .A2(
        u5_mult_82_SUMB_24__8_), .ZN(u5_mult_82_n3310) );
  XNOR2_X2 u5_mult_82_U6158 ( .A(u5_mult_82_ab_30__38_), .B(
        u5_mult_82_CARRYB_29__38_), .ZN(u5_mult_82_n2069) );
  XNOR2_X2 u5_mult_82_U6157 ( .A(u5_mult_82_n2069), .B(u5_mult_82_SUMB_29__39_), .ZN(u5_mult_82_SUMB_30__38_) );
  NAND3_X4 u5_mult_82_U6156 ( .A1(u5_mult_82_n6183), .A2(u5_mult_82_n6184), 
        .A3(u5_mult_82_n6185), .ZN(u5_mult_82_CARRYB_27__25_) );
  NAND2_X2 u5_mult_82_U6155 ( .A1(u5_mult_82_CARRYB_20__29_), .A2(
        u5_mult_82_SUMB_20__30_), .ZN(u5_mult_82_n5058) );
  NAND2_X2 u5_mult_82_U6154 ( .A1(u5_mult_82_CARRYB_28__37_), .A2(
        u5_mult_82_n1702), .ZN(u5_mult_82_n4644) );
  NAND2_X2 u5_mult_82_U6153 ( .A1(u5_mult_82_CARRYB_6__39_), .A2(
        u5_mult_82_n1592), .ZN(u5_mult_82_n5806) );
  NAND3_X2 u5_mult_82_U6152 ( .A1(u5_mult_82_n5454), .A2(u5_mult_82_n5455), 
        .A3(u5_mult_82_n5456), .ZN(u5_mult_82_CARRYB_11__37_) );
  XNOR2_X2 u5_mult_82_U6151 ( .A(u5_mult_82_ab_12__37_), .B(
        u5_mult_82_CARRYB_11__37_), .ZN(u5_mult_82_n2068) );
  XNOR2_X2 u5_mult_82_U6150 ( .A(u5_mult_82_SUMB_11__38_), .B(u5_mult_82_n2068), .ZN(u5_mult_82_SUMB_12__37_) );
  NAND2_X1 u5_mult_82_U6149 ( .A1(u5_mult_82_CARRYB_16__35_), .A2(
        u5_mult_82_SUMB_16__36_), .ZN(u5_mult_82_n6192) );
  NAND3_X4 u5_mult_82_U6148 ( .A1(u5_mult_82_n2729), .A2(u5_mult_82_n2728), 
        .A3(u5_mult_82_n2727), .ZN(u5_mult_82_CARRYB_16__43_) );
  NAND2_X2 u5_mult_82_U6147 ( .A1(u5_mult_82_ab_24__10_), .A2(
        u5_mult_82_SUMB_23__11_), .ZN(u5_mult_82_n4120) );
  NAND2_X2 u5_mult_82_U6146 ( .A1(u5_mult_82_SUMB_23__11_), .A2(
        u5_mult_82_CARRYB_23__10_), .ZN(u5_mult_82_n4121) );
  XNOR2_X2 u5_mult_82_U6145 ( .A(u5_mult_82_ab_5__44_), .B(
        u5_mult_82_CARRYB_4__44_), .ZN(u5_mult_82_n2067) );
  XNOR2_X2 u5_mult_82_U6144 ( .A(u5_mult_82_n2067), .B(u5_mult_82_SUMB_4__45_), 
        .ZN(u5_mult_82_SUMB_5__44_) );
  NAND2_X1 u5_mult_82_U6143 ( .A1(u5_mult_82_SUMB_15__33_), .A2(
        u5_mult_82_CARRYB_15__32_), .ZN(u5_mult_82_n4864) );
  NAND3_X2 u5_mult_82_U6142 ( .A1(u5_mult_82_n4680), .A2(u5_mult_82_n4681), 
        .A3(u5_mult_82_n4682), .ZN(u5_mult_82_CARRYB_37__3_) );
  NAND2_X1 u5_mult_82_U6141 ( .A1(u5_mult_82_CARRYB_25__29_), .A2(
        u5_mult_82_n1428), .ZN(u5_mult_82_n5545) );
  NAND2_X2 u5_mult_82_U6140 ( .A1(u5_mult_82_ab_34__5_), .A2(
        u5_mult_82_CARRYB_33__5_), .ZN(u5_mult_82_n3176) );
  INV_X2 u5_mult_82_U6139 ( .A(u5_mult_82_SUMB_23__10_), .ZN(u5_mult_82_n2558)
         );
  XOR2_X1 u5_mult_82_U6138 ( .A(u5_mult_82_CARRYB_43__0_), .B(
        u5_mult_82_ab_44__0_), .Z(u5_mult_82_n4840) );
  NAND2_X2 u5_mult_82_U6137 ( .A1(u5_mult_82_CARRYB_26__8_), .A2(
        u5_mult_82_SUMB_26__9_), .ZN(u5_mult_82_n3623) );
  XNOR2_X2 u5_mult_82_U6136 ( .A(u5_mult_82_CARRYB_31__7_), .B(
        u5_mult_82_ab_32__7_), .ZN(u5_mult_82_n2571) );
  XNOR2_X2 u5_mult_82_U6135 ( .A(u5_mult_82_n2066), .B(
        u5_mult_82_CARRYB_16__15_), .ZN(u5_mult_82_n3970) );
  NAND2_X1 u5_mult_82_U6134 ( .A1(u5_mult_82_ab_41__17_), .A2(
        u5_mult_82_CARRYB_40__17_), .ZN(u5_mult_82_n5061) );
  NAND2_X1 u5_mult_82_U6133 ( .A1(u5_mult_82_ab_38__5_), .A2(
        u5_mult_82_CARRYB_37__5_), .ZN(u5_mult_82_n4150) );
  NOR2_X2 u5_mult_82_U6132 ( .A1(u5_mult_82_net64379), .A2(u5_mult_82_n6665), 
        .ZN(u5_mult_82_ab_28__6_) );
  NAND3_X4 u5_mult_82_U6131 ( .A1(u5_mult_82_n2063), .A2(u5_mult_82_n2064), 
        .A3(u5_mult_82_n2065), .ZN(u5_mult_82_CARRYB_28__6_) );
  NAND2_X1 u5_mult_82_U6130 ( .A1(u5_mult_82_ab_28__6_), .A2(
        u5_mult_82_CARRYB_27__6_), .ZN(u5_mult_82_n2065) );
  NAND2_X2 u5_mult_82_U6129 ( .A1(u5_mult_82_ab_28__6_), .A2(
        u5_mult_82_SUMB_27__7_), .ZN(u5_mult_82_n2064) );
  NAND2_X2 u5_mult_82_U6128 ( .A1(u5_mult_82_CARRYB_27__6_), .A2(
        u5_mult_82_SUMB_27__7_), .ZN(u5_mult_82_n2063) );
  XOR2_X2 u5_mult_82_U6127 ( .A(u5_mult_82_CARRYB_27__6_), .B(
        u5_mult_82_ab_28__6_), .Z(u5_mult_82_n2062) );
  NAND3_X2 u5_mult_82_U6126 ( .A1(u5_mult_82_n2059), .A2(u5_mult_82_n2060), 
        .A3(u5_mult_82_n2061), .ZN(u5_mult_82_CARRYB_30__6_) );
  NAND2_X1 u5_mult_82_U6125 ( .A1(u5_mult_82_SUMB_29__7_), .A2(
        u5_mult_82_CARRYB_29__6_), .ZN(u5_mult_82_n2061) );
  NAND2_X2 u5_mult_82_U6124 ( .A1(u5_mult_82_ab_30__6_), .A2(
        u5_mult_82_CARRYB_29__6_), .ZN(u5_mult_82_n2060) );
  NAND2_X1 u5_mult_82_U6123 ( .A1(u5_mult_82_ab_30__6_), .A2(
        u5_mult_82_SUMB_29__7_), .ZN(u5_mult_82_n2059) );
  XOR2_X2 u5_mult_82_U6122 ( .A(u5_mult_82_n2058), .B(u5_mult_82_CARRYB_29__6_), .Z(u5_mult_82_SUMB_30__6_) );
  XOR2_X1 u5_mult_82_U6121 ( .A(u5_mult_82_ab_30__6_), .B(
        u5_mult_82_SUMB_29__7_), .Z(u5_mult_82_n2058) );
  NAND3_X2 u5_mult_82_U6120 ( .A1(u5_mult_82_n2055), .A2(u5_mult_82_n2056), 
        .A3(u5_mult_82_n2057), .ZN(u5_mult_82_CARRYB_29__6_) );
  NAND2_X2 u5_mult_82_U6119 ( .A1(u5_mult_82_ab_29__6_), .A2(
        u5_mult_82_SUMB_28__7_), .ZN(u5_mult_82_n2057) );
  NAND2_X1 u5_mult_82_U6118 ( .A1(u5_mult_82_CARRYB_28__6_), .A2(
        u5_mult_82_SUMB_28__7_), .ZN(u5_mult_82_n2056) );
  NAND2_X2 u5_mult_82_U6117 ( .A1(u5_mult_82_CARRYB_28__6_), .A2(
        u5_mult_82_ab_29__6_), .ZN(u5_mult_82_n2055) );
  XOR2_X1 u5_mult_82_U6116 ( .A(u5_mult_82_n2054), .B(u5_mult_82_SUMB_28__7_), 
        .Z(u5_mult_82_SUMB_29__6_) );
  XOR2_X2 u5_mult_82_U6115 ( .A(u5_mult_82_CARRYB_28__6_), .B(
        u5_mult_82_ab_29__6_), .Z(u5_mult_82_n2054) );
  NAND2_X1 u5_mult_82_U6114 ( .A1(u5_mult_82_CARRYB_35__29_), .A2(
        u5_mult_82_SUMB_35__30_), .ZN(u5_mult_82_n4876) );
  NAND2_X1 u5_mult_82_U6113 ( .A1(u5_mult_82_ab_15__42_), .A2(
        u5_mult_82_SUMB_14__43_), .ZN(u5_mult_82_n3132) );
  XNOR2_X2 u5_mult_82_U6112 ( .A(u5_mult_82_n2053), .B(u5_mult_82_n66), .ZN(
        u5_mult_82_SUMB_20__40_) );
  XNOR2_X2 u5_mult_82_U6111 ( .A(u5_mult_82_ab_30__22_), .B(
        u5_mult_82_CARRYB_29__22_), .ZN(u5_mult_82_n2052) );
  NAND2_X1 u5_mult_82_U6110 ( .A1(u5_mult_82_ab_31__36_), .A2(
        u5_mult_82_CARRYB_30__36_), .ZN(u5_mult_82_n4319) );
  NAND2_X1 u5_mult_82_U6109 ( .A1(u5_mult_82_SUMB_11__40_), .A2(
        u5_mult_82_CARRYB_11__39_), .ZN(u5_mult_82_n6158) );
  NAND2_X2 u5_mult_82_U6108 ( .A1(u5_mult_82_CARRYB_28__27_), .A2(
        u5_mult_82_n20), .ZN(u5_mult_82_n6270) );
  NAND3_X2 u5_mult_82_U6107 ( .A1(u5_mult_82_n2048), .A2(u5_mult_82_n2049), 
        .A3(u5_mult_82_n2050), .ZN(u5_mult_82_CARRYB_22__10_) );
  NAND2_X2 u5_mult_82_U6106 ( .A1(u5_mult_82_ab_22__10_), .A2(
        u5_mult_82_SUMB_21__11_), .ZN(u5_mult_82_n2050) );
  NAND2_X2 u5_mult_82_U6105 ( .A1(u5_mult_82_CARRYB_21__10_), .A2(
        u5_mult_82_SUMB_21__11_), .ZN(u5_mult_82_n2049) );
  NAND2_X1 u5_mult_82_U6104 ( .A1(u5_mult_82_CARRYB_21__10_), .A2(
        u5_mult_82_ab_22__10_), .ZN(u5_mult_82_n2048) );
  NAND2_X2 u5_mult_82_U6103 ( .A1(u5_mult_82_CARRYB_20__11_), .A2(
        u5_mult_82_SUMB_20__12_), .ZN(u5_mult_82_n2047) );
  NAND2_X2 u5_mult_82_U6102 ( .A1(u5_mult_82_ab_21__11_), .A2(
        u5_mult_82_SUMB_20__12_), .ZN(u5_mult_82_n2046) );
  NAND2_X2 u5_mult_82_U6101 ( .A1(u5_mult_82_ab_21__11_), .A2(
        u5_mult_82_CARRYB_20__11_), .ZN(u5_mult_82_n2045) );
  XOR2_X2 u5_mult_82_U6100 ( .A(u5_mult_82_n2044), .B(u5_mult_82_SUMB_21__11_), 
        .Z(u5_mult_82_SUMB_22__10_) );
  XOR2_X2 u5_mult_82_U6099 ( .A(u5_mult_82_CARRYB_21__10_), .B(
        u5_mult_82_ab_22__10_), .Z(u5_mult_82_n2044) );
  XOR2_X2 u5_mult_82_U6098 ( .A(u5_mult_82_n2043), .B(u5_mult_82_SUMB_20__12_), 
        .Z(u5_mult_82_SUMB_21__11_) );
  XOR2_X2 u5_mult_82_U6097 ( .A(u5_mult_82_ab_21__11_), .B(
        u5_mult_82_CARRYB_20__11_), .Z(u5_mult_82_n2043) );
  NAND2_X1 u5_mult_82_U6096 ( .A1(u5_mult_82_ab_40__5_), .A2(
        u5_mult_82_CARRYB_39__5_), .ZN(u5_mult_82_n4968) );
  XNOR2_X2 u5_mult_82_U6095 ( .A(u5_mult_82_CARRYB_25__13_), .B(
        u5_mult_82_n2042), .ZN(u5_mult_82_n4829) );
  NAND2_X2 u5_mult_82_U6094 ( .A1(u5_mult_82_ab_30__26_), .A2(
        u5_mult_82_SUMB_29__27_), .ZN(u5_mult_82_n6272) );
  NAND2_X2 u5_mult_82_U6093 ( .A1(u5_mult_82_CARRYB_29__26_), .A2(
        u5_mult_82_SUMB_29__27_), .ZN(u5_mult_82_n6273) );
  NAND2_X2 u5_mult_82_U6092 ( .A1(u5_mult_82_SUMB_7__42_), .A2(
        u5_mult_82_CARRYB_7__41_), .ZN(u5_mult_82_n5981) );
  NAND2_X2 u5_mult_82_U6091 ( .A1(u5_mult_82_ab_44__8_), .A2(
        u5_mult_82_SUMB_43__9_), .ZN(u5_mult_82_n5492) );
  NAND2_X2 u5_mult_82_U6090 ( .A1(u5_mult_82_CARRYB_43__8_), .A2(
        u5_mult_82_SUMB_43__9_), .ZN(u5_mult_82_n5493) );
  NAND3_X2 u5_mult_82_U6089 ( .A1(u5_mult_82_n3962), .A2(u5_mult_82_n3961), 
        .A3(u5_mult_82_n3963), .ZN(u5_mult_82_CARRYB_38__7_) );
  XNOR2_X2 u5_mult_82_U6088 ( .A(u5_mult_82_CARRYB_9__38_), .B(
        u5_mult_82_ab_10__38_), .ZN(u5_mult_82_n2041) );
  XNOR2_X2 u5_mult_82_U6087 ( .A(u5_mult_82_SUMB_9__39_), .B(u5_mult_82_n2041), 
        .ZN(u5_mult_82_SUMB_10__38_) );
  NAND2_X1 u5_mult_82_U6086 ( .A1(u5_mult_82_CARRYB_14__33_), .A2(
        u5_mult_82_ab_15__33_), .ZN(u5_mult_82_n4859) );
  NAND2_X1 u5_mult_82_U6085 ( .A1(u5_mult_82_SUMB_45__15_), .A2(
        u5_mult_82_CARRYB_45__14_), .ZN(u5_mult_82_n5776) );
  NAND2_X2 u5_mult_82_U6084 ( .A1(u5_mult_82_ab_38__2_), .A2(
        u5_mult_82_SUMB_37__3_), .ZN(u5_mult_82_n4684) );
  NAND2_X1 u5_mult_82_U6083 ( .A1(u5_mult_82_SUMB_26__11_), .A2(
        u5_mult_82_ab_27__10_), .ZN(u5_mult_82_n3905) );
  XNOR2_X2 u5_mult_82_U6082 ( .A(u5_mult_82_CARRYB_25__38_), .B(
        u5_mult_82_ab_26__38_), .ZN(u5_mult_82_n2040) );
  XNOR2_X2 u5_mult_82_U6081 ( .A(u5_mult_82_SUMB_25__39_), .B(u5_mult_82_n2040), .ZN(u5_mult_82_SUMB_26__38_) );
  NOR2_X1 u5_mult_82_U6080 ( .A1(u5_mult_82_n6953), .A2(u5_mult_82_n6687), 
        .ZN(u5_mult_82_ab_31__3_) );
  NOR2_X1 u5_mult_82_U6079 ( .A1(u5_mult_82_n6986), .A2(u5_mult_82_net65393), 
        .ZN(u5_mult_82_ab_41__0_) );
  NOR2_X1 u5_mult_82_U6078 ( .A1(u5_mult_82_n6986), .A2(u5_mult_82_n6749), 
        .ZN(u5_mult_82_ab_48__0_) );
  NAND3_X2 u5_mult_82_U6077 ( .A1(u5_mult_82_n2037), .A2(u5_mult_82_n2038), 
        .A3(u5_mult_82_n2039), .ZN(u5_mult_82_CARRYB_31__3_) );
  NAND2_X1 u5_mult_82_U6076 ( .A1(u5_mult_82_ab_31__3_), .A2(
        u5_mult_82_SUMB_30__4_), .ZN(u5_mult_82_n2039) );
  NAND2_X2 u5_mult_82_U6075 ( .A1(u5_mult_82_ab_31__3_), .A2(
        u5_mult_82_CARRYB_30__3_), .ZN(u5_mult_82_n2038) );
  XOR2_X2 u5_mult_82_U6074 ( .A(u5_mult_82_SUMB_30__4_), .B(
        u5_mult_82_ab_31__3_), .Z(u5_mult_82_n2036) );
  NAND3_X2 u5_mult_82_U6073 ( .A1(u5_mult_82_n2033), .A2(u5_mult_82_n2034), 
        .A3(u5_mult_82_n2035), .ZN(u5_mult_82_CARRYB_41__0_) );
  NAND2_X1 u5_mult_82_U6072 ( .A1(u5_mult_82_ab_41__0_), .A2(
        u5_mult_82_CARRYB_40__0_), .ZN(u5_mult_82_n2035) );
  NAND2_X2 u5_mult_82_U6071 ( .A1(u5_mult_82_ab_41__0_), .A2(
        u5_mult_82_SUMB_40__1_), .ZN(u5_mult_82_n2034) );
  XOR2_X2 u5_mult_82_U6070 ( .A(u5_mult_82_SUMB_40__1_), .B(u5_mult_82_n2032), 
        .Z(u5_N41) );
  XOR2_X2 u5_mult_82_U6069 ( .A(u5_mult_82_CARRYB_40__0_), .B(
        u5_mult_82_ab_41__0_), .Z(u5_mult_82_n2032) );
  NAND3_X2 u5_mult_82_U6068 ( .A1(u5_mult_82_n2031), .A2(u5_mult_82_n2030), 
        .A3(u5_mult_82_n2029), .ZN(u5_mult_82_CARRYB_48__0_) );
  XOR2_X2 u5_mult_82_U6067 ( .A(u5_mult_82_SUMB_47__1_), .B(
        u5_mult_82_ab_48__0_), .Z(u5_mult_82_n2028) );
  NAND3_X2 u5_mult_82_U6066 ( .A1(u5_mult_82_n2025), .A2(u5_mult_82_n2026), 
        .A3(u5_mult_82_n2027), .ZN(u5_mult_82_CARRYB_16__9_) );
  NAND2_X1 u5_mult_82_U6065 ( .A1(u5_mult_82_CARRYB_15__9_), .A2(
        u5_mult_82_SUMB_15__10_), .ZN(u5_mult_82_n2027) );
  NAND2_X1 u5_mult_82_U6064 ( .A1(u5_mult_82_ab_16__9_), .A2(
        u5_mult_82_SUMB_15__10_), .ZN(u5_mult_82_n2026) );
  NAND2_X1 u5_mult_82_U6063 ( .A1(u5_mult_82_ab_16__9_), .A2(
        u5_mult_82_CARRYB_15__9_), .ZN(u5_mult_82_n2025) );
  NAND3_X2 u5_mult_82_U6062 ( .A1(u5_mult_82_n2022), .A2(u5_mult_82_n2023), 
        .A3(u5_mult_82_n2024), .ZN(u5_mult_82_CARRYB_15__10_) );
  NAND2_X2 u5_mult_82_U6061 ( .A1(u5_mult_82_CARRYB_14__10_), .A2(
        u5_mult_82_SUMB_14__11_), .ZN(u5_mult_82_n2024) );
  NAND2_X2 u5_mult_82_U6060 ( .A1(u5_mult_82_ab_15__10_), .A2(
        u5_mult_82_SUMB_14__11_), .ZN(u5_mult_82_n2023) );
  NAND2_X1 u5_mult_82_U6059 ( .A1(u5_mult_82_ab_15__10_), .A2(
        u5_mult_82_CARRYB_14__10_), .ZN(u5_mult_82_n2022) );
  XOR2_X2 u5_mult_82_U6058 ( .A(u5_mult_82_n2021), .B(u5_mult_82_SUMB_15__10_), 
        .Z(u5_mult_82_SUMB_16__9_) );
  XOR2_X2 u5_mult_82_U6057 ( .A(u5_mult_82_ab_16__9_), .B(
        u5_mult_82_CARRYB_15__9_), .Z(u5_mult_82_n2021) );
  XOR2_X2 u5_mult_82_U6056 ( .A(u5_mult_82_n2020), .B(u5_mult_82_SUMB_14__11_), 
        .Z(u5_mult_82_SUMB_15__10_) );
  XOR2_X2 u5_mult_82_U6055 ( .A(u5_mult_82_ab_15__10_), .B(
        u5_mult_82_CARRYB_14__10_), .Z(u5_mult_82_n2020) );
  NAND2_X2 u5_mult_82_U6054 ( .A1(u5_mult_82_SUMB_7__42_), .A2(
        u5_mult_82_ab_8__41_), .ZN(u5_mult_82_n5980) );
  NAND3_X4 u5_mult_82_U6053 ( .A1(u5_mult_82_n5979), .A2(u5_mult_82_n5980), 
        .A3(u5_mult_82_n5981), .ZN(u5_mult_82_CARRYB_8__41_) );
  NAND3_X2 u5_mult_82_U6052 ( .A1(u5_mult_82_n3892), .A2(u5_mult_82_n3893), 
        .A3(u5_mult_82_n3894), .ZN(u5_mult_82_CARRYB_16__20_) );
  NAND2_X2 u5_mult_82_U6051 ( .A1(u5_mult_82_CARRYB_39__5_), .A2(
        u5_mult_82_SUMB_39__6_), .ZN(u5_mult_82_n4966) );
  NAND2_X2 u5_mult_82_U6050 ( .A1(u5_mult_82_ab_45__2_), .A2(u5_mult_82_n1833), 
        .ZN(u5_mult_82_n5628) );
  NAND2_X2 u5_mult_82_U6049 ( .A1(u5_mult_82_CARRYB_9__37_), .A2(
        u5_mult_82_SUMB_9__38_), .ZN(u5_mult_82_n5906) );
  NAND2_X2 u5_mult_82_U6048 ( .A1(u5_mult_82_CARRYB_38__28_), .A2(
        u5_mult_82_SUMB_38__29_), .ZN(u5_mult_82_n5278) );
  XNOR2_X2 u5_mult_82_U6047 ( .A(u5_mult_82_n2019), .B(
        u5_mult_82_CARRYB_51__20_), .ZN(u5_mult_82_n5100) );
  NAND3_X4 u5_mult_82_U6046 ( .A1(u5_mult_82_n5664), .A2(u5_mult_82_n5665), 
        .A3(u5_mult_82_n5666), .ZN(u5_mult_82_CARRYB_28__37_) );
  NAND2_X2 u5_mult_82_U6045 ( .A1(u5_mult_82_ab_24__37_), .A2(
        u5_mult_82_CARRYB_23__37_), .ZN(u5_mult_82_n5559) );
  XNOR2_X2 u5_mult_82_U6044 ( .A(u5_mult_82_ab_21__42_), .B(
        u5_mult_82_CARRYB_20__42_), .ZN(u5_mult_82_n2018) );
  XNOR2_X2 u5_mult_82_U6043 ( .A(u5_mult_82_n2018), .B(u5_mult_82_SUMB_20__43_), .ZN(u5_mult_82_SUMB_21__42_) );
  XNOR2_X2 u5_mult_82_U6042 ( .A(u5_mult_82_SUMB_14__32_), .B(u5_mult_82_n2017), .ZN(u5_mult_82_SUMB_15__31_) );
  INV_X4 u5_mult_82_U6041 ( .A(u5_mult_82_n6835), .ZN(u5_mult_82_n6831) );
  XNOR2_X2 u5_mult_82_U6040 ( .A(u5_mult_82_net86085), .B(
        u5_mult_82_SUMB_19__27_), .ZN(u5_mult_82_SUMB_20__26_) );
  NAND2_X4 u5_mult_82_U6039 ( .A1(u5_mult_82_net64225), .A2(n4762), .ZN(
        u5_mult_82_n2016) );
  XOR2_X2 u5_mult_82_U6038 ( .A(u5_mult_82_n5867), .B(u5_mult_82_SUMB_32__31_), 
        .Z(u5_mult_82_SUMB_33__30_) );
  NAND3_X2 u5_mult_82_U6037 ( .A1(u5_mult_82_n6030), .A2(u5_mult_82_n6031), 
        .A3(u5_mult_82_n6032), .ZN(u5_mult_82_CARRYB_43__6_) );
  NAND2_X1 u5_mult_82_U6036 ( .A1(u5_mult_82_CARRYB_34__30_), .A2(
        u5_mult_82_SUMB_34__31_), .ZN(u5_mult_82_n4873) );
  NAND3_X4 u5_mult_82_U6035 ( .A1(u5_mult_82_n5582), .A2(u5_mult_82_n5583), 
        .A3(u5_mult_82_n5584), .ZN(u5_mult_82_CARRYB_41__28_) );
  NAND2_X1 u5_mult_82_U6034 ( .A1(u5_mult_82_CARRYB_39__6_), .A2(
        u5_mult_82_SUMB_39__7_), .ZN(u5_mult_82_n5817) );
  INV_X4 u5_mult_82_U6033 ( .A(u5_mult_82_CARRYB_40__6_), .ZN(u5_mult_82_n2981) );
  NAND2_X2 u5_mult_82_U6032 ( .A1(u5_mult_82_ab_23__34_), .A2(
        u5_mult_82_SUMB_22__35_), .ZN(u5_mult_82_n6376) );
  NAND2_X2 u5_mult_82_U6031 ( .A1(u5_mult_82_ab_17__25_), .A2(
        u5_mult_82_SUMB_16__26_), .ZN(u5_mult_82_n4630) );
  NOR2_X4 u5_mult_82_U6030 ( .A1(u5_mult_82_n6793), .A2(u5_mult_82_n6564), 
        .ZN(u5_mult_82_ab_12__46_) );
  INV_X2 u5_mult_82_U6029 ( .A(u5_mult_82_ab_12__46_), .ZN(u5_mult_82_n2013)
         );
  INV_X4 u5_mult_82_U6028 ( .A(u5_mult_82_CARRYB_11__46_), .ZN(
        u5_mult_82_n2012) );
  NAND2_X4 u5_mult_82_U6027 ( .A1(u5_mult_82_n2014), .A2(u5_mult_82_n2015), 
        .ZN(u5_mult_82_n4787) );
  NAND2_X4 u5_mult_82_U6026 ( .A1(u5_mult_82_n2012), .A2(u5_mult_82_n2013), 
        .ZN(u5_mult_82_n2015) );
  NAND2_X2 u5_mult_82_U6025 ( .A1(u5_mult_82_CARRYB_11__46_), .A2(
        u5_mult_82_ab_12__46_), .ZN(u5_mult_82_n2014) );
  NAND2_X1 u5_mult_82_U6024 ( .A1(u5_mult_82_CARRYB_27__31_), .A2(
        u5_mult_82_SUMB_27__32_), .ZN(u5_mult_82_n2815) );
  INV_X8 u5_mult_82_U6023 ( .A(u5_mult_82_n7011), .ZN(u5_mult_82_n6847) );
  INV_X16 u5_mult_82_U6022 ( .A(u5_mult_82_n7011), .ZN(u5_mult_82_n6848) );
  INV_X8 u5_mult_82_U6021 ( .A(n4744), .ZN(u5_mult_82_n7011) );
  XOR2_X2 u5_mult_82_U6020 ( .A(u5_mult_82_n2573), .B(u5_mult_82_SUMB_24__44_), 
        .Z(u5_mult_82_SUMB_25__43_) );
  NAND3_X4 u5_mult_82_U6019 ( .A1(u5_mult_82_n2820), .A2(u5_mult_82_n2819), 
        .A3(u5_mult_82_n2818), .ZN(u5_mult_82_CARRYB_24__12_) );
  NAND2_X2 u5_mult_82_U6018 ( .A1(u5_mult_82_ab_27__8_), .A2(
        u5_mult_82_SUMB_26__9_), .ZN(u5_mult_82_n3622) );
  NAND2_X1 u5_mult_82_U6017 ( .A1(u5_mult_82_CARRYB_17__20_), .A2(
        u5_mult_82_SUMB_17__21_), .ZN(u5_mult_82_n4370) );
  NAND2_X1 u5_mult_82_U6016 ( .A1(u5_mult_82_ab_18__20_), .A2(
        u5_mult_82_CARRYB_17__20_), .ZN(u5_mult_82_n4368) );
  NAND2_X2 u5_mult_82_U6015 ( .A1(u5_mult_82_ab_18__30_), .A2(
        u5_mult_82_SUMB_17__31_), .ZN(u5_mult_82_n6013) );
  NAND2_X1 u5_mult_82_U6014 ( .A1(u5_mult_82_ab_23__28_), .A2(
        u5_mult_82_SUMB_22__29_), .ZN(u5_mult_82_n4298) );
  INV_X8 u5_mult_82_U6013 ( .A(u5_mult_82_n7010), .ZN(u5_mult_82_n6834) );
  XNOR2_X2 u5_mult_82_U6012 ( .A(u5_mult_82_ab_17__26_), .B(
        u5_mult_82_CARRYB_16__26_), .ZN(u5_mult_82_n2122) );
  NAND2_X1 u5_mult_82_U6011 ( .A1(u5_mult_82_ab_9__46_), .A2(
        u5_mult_82_CARRYB_8__46_), .ZN(u5_mult_82_n4796) );
  XNOR2_X2 u5_mult_82_U6010 ( .A(u5_mult_82_CARRYB_31__30_), .B(
        u5_mult_82_ab_32__30_), .ZN(u5_mult_82_n5649) );
  NAND2_X2 u5_mult_82_U6009 ( .A1(u5_mult_82_ab_24__27_), .A2(
        u5_mult_82_SUMB_23__28_), .ZN(u5_mult_82_n6142) );
  NAND2_X2 u5_mult_82_U6008 ( .A1(u5_mult_82_CARRYB_35__34_), .A2(
        u5_mult_82_SUMB_35__35_), .ZN(u5_mult_82_n3930) );
  XNOR2_X2 u5_mult_82_U6007 ( .A(u5_mult_82_CARRYB_14__33_), .B(
        u5_mult_82_n2011), .ZN(u5_mult_82_n4858) );
  XNOR2_X1 u5_mult_82_U6006 ( .A(u5_mult_82_ab_20__21_), .B(
        u5_mult_82_SUMB_19__22_), .ZN(u5_mult_82_n2010) );
  XNOR2_X2 u5_mult_82_U6005 ( .A(u5_mult_82_n2010), .B(
        u5_mult_82_CARRYB_19__21_), .ZN(u5_mult_82_SUMB_20__21_) );
  XNOR2_X2 u5_mult_82_U6004 ( .A(u5_mult_82_ab_12__38_), .B(
        u5_mult_82_CARRYB_11__38_), .ZN(u5_mult_82_n2009) );
  XNOR2_X2 u5_mult_82_U6003 ( .A(u5_mult_82_n2009), .B(u5_mult_82_n5184), .ZN(
        u5_mult_82_SUMB_12__38_) );
  NAND2_X2 u5_mult_82_U6002 ( .A1(u5_mult_82_CARRYB_12__16_), .A2(
        u5_mult_82_SUMB_12__17_), .ZN(u5_mult_82_n3544) );
  XNOR2_X2 u5_mult_82_U6001 ( .A(u5_mult_82_ab_23__31_), .B(
        u5_mult_82_CARRYB_22__31_), .ZN(u5_mult_82_n2008) );
  XNOR2_X2 u5_mult_82_U6000 ( .A(u5_mult_82_n2008), .B(u5_mult_82_SUMB_22__32_), .ZN(u5_mult_82_SUMB_23__31_) );
  XNOR2_X2 u5_mult_82_U5999 ( .A(u5_mult_82_CARRYB_9__37_), .B(
        u5_mult_82_n2007), .ZN(u5_mult_82_n5902) );
  NAND2_X2 u5_mult_82_U5998 ( .A1(u5_mult_82_CARRYB_23__27_), .A2(
        u5_mult_82_SUMB_23__28_), .ZN(u5_mult_82_n6143) );
  NAND2_X2 u5_mult_82_U5997 ( .A1(u5_mult_82_ab_0__45_), .A2(
        u5_mult_82_ab_1__44_), .ZN(u5_mult_82_n6498) );
  NAND2_X1 u5_mult_82_U5996 ( .A1(u5_mult_82_ab_17__27_), .A2(
        u5_mult_82_CARRYB_16__27_), .ZN(u5_mult_82_n5606) );
  NAND2_X1 u5_mult_82_U5995 ( .A1(u5_mult_82_CARRYB_29__31_), .A2(
        u5_mult_82_SUMB_29__32_), .ZN(u5_mult_82_n5162) );
  NAND3_X4 u5_mult_82_U5994 ( .A1(u5_mult_82_n3610), .A2(u5_mult_82_n3611), 
        .A3(u5_mult_82_n3612), .ZN(u5_mult_82_CARRYB_35__33_) );
  XOR2_X2 u5_mult_82_U5993 ( .A(u5_mult_82_n11), .B(u5_mult_82_n2036), .Z(
        u5_mult_82_SUMB_31__3_) );
  NAND2_X2 u5_mult_82_U5992 ( .A1(u5_mult_82_CARRYB_40__1_), .A2(
        u5_mult_82_SUMB_40__2_), .ZN(u5_mult_82_n4527) );
  NOR2_X2 u5_mult_82_U5991 ( .A1(u5_mult_82_n6927), .A2(u5_mult_82_n6664), 
        .ZN(u5_mult_82_ab_28__17_) );
  NOR2_X1 u5_mult_82_U5990 ( .A1(u5_mult_82_n6933), .A2(u5_mult_82_n6686), 
        .ZN(u5_mult_82_ab_31__15_) );
  NAND2_X4 u5_mult_82_U5989 ( .A1(u5_mult_82_n3785), .A2(u5_mult_82_n3786), 
        .ZN(u5_mult_82_SUMB_35__14_) );
  NOR2_X1 u5_mult_82_U5988 ( .A1(u5_mult_82_net64505), .A2(u5_mult_82_n6716), 
        .ZN(u5_mult_82_ab_36__13_) );
  NAND3_X4 u5_mult_82_U5987 ( .A1(u5_mult_82_n2003), .A2(u5_mult_82_n2004), 
        .A3(u5_mult_82_n2005), .ZN(u5_mult_82_CARRYB_28__17_) );
  NAND2_X2 u5_mult_82_U5986 ( .A1(u5_mult_82_ab_28__17_), .A2(
        u5_mult_82_SUMB_27__18_), .ZN(u5_mult_82_n2005) );
  NAND2_X2 u5_mult_82_U5985 ( .A1(u5_mult_82_ab_28__17_), .A2(
        u5_mult_82_CARRYB_27__17_), .ZN(u5_mult_82_n2004) );
  NAND2_X2 u5_mult_82_U5984 ( .A1(u5_mult_82_SUMB_27__18_), .A2(
        u5_mult_82_CARRYB_27__17_), .ZN(u5_mult_82_n2003) );
  NAND3_X2 u5_mult_82_U5983 ( .A1(u5_mult_82_n2000), .A2(u5_mult_82_n2001), 
        .A3(u5_mult_82_n2002), .ZN(u5_mult_82_CARRYB_31__15_) );
  NAND2_X1 u5_mult_82_U5982 ( .A1(u5_mult_82_ab_31__15_), .A2(
        u5_mult_82_CARRYB_30__15_), .ZN(u5_mult_82_n2002) );
  NAND2_X2 u5_mult_82_U5981 ( .A1(u5_mult_82_ab_31__15_), .A2(
        u5_mult_82_SUMB_30__16_), .ZN(u5_mult_82_n2001) );
  XOR2_X2 u5_mult_82_U5980 ( .A(u5_mult_82_SUMB_30__16_), .B(u5_mult_82_n1999), 
        .Z(u5_mult_82_SUMB_31__15_) );
  XOR2_X2 u5_mult_82_U5979 ( .A(u5_mult_82_CARRYB_30__15_), .B(
        u5_mult_82_ab_31__15_), .Z(u5_mult_82_n1999) );
  NAND2_X1 u5_mult_82_U5978 ( .A1(u5_mult_82_ab_36__13_), .A2(
        u5_mult_82_CARRYB_35__13_), .ZN(u5_mult_82_n1998) );
  NAND3_X2 u5_mult_82_U5977 ( .A1(u5_mult_82_n1993), .A2(u5_mult_82_n1994), 
        .A3(u5_mult_82_n1995), .ZN(u5_mult_82_CARRYB_30__16_) );
  NAND2_X2 u5_mult_82_U5976 ( .A1(u5_mult_82_CARRYB_29__16_), .A2(
        u5_mult_82_SUMB_29__17_), .ZN(u5_mult_82_n1995) );
  NAND2_X2 u5_mult_82_U5975 ( .A1(u5_mult_82_ab_30__16_), .A2(
        u5_mult_82_SUMB_29__17_), .ZN(u5_mult_82_n1994) );
  NAND2_X1 u5_mult_82_U5974 ( .A1(u5_mult_82_ab_30__16_), .A2(
        u5_mult_82_CARRYB_29__16_), .ZN(u5_mult_82_n1993) );
  NAND3_X4 u5_mult_82_U5973 ( .A1(u5_mult_82_n1992), .A2(u5_mult_82_n1991), 
        .A3(u5_mult_82_n1990), .ZN(u5_mult_82_CARRYB_29__17_) );
  NAND2_X2 u5_mult_82_U5972 ( .A1(u5_mult_82_CARRYB_28__17_), .A2(
        u5_mult_82_n431), .ZN(u5_mult_82_n1992) );
  NAND2_X2 u5_mult_82_U5971 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_ab_29__17_), 
        .ZN(u5_mult_82_n1991) );
  XOR2_X2 u5_mult_82_U5970 ( .A(u5_mult_82_n1989), .B(u5_mult_82_SUMB_29__17_), 
        .Z(u5_mult_82_SUMB_30__16_) );
  XOR2_X2 u5_mult_82_U5969 ( .A(u5_mult_82_ab_30__16_), .B(
        u5_mult_82_CARRYB_29__16_), .Z(u5_mult_82_n1989) );
  XOR2_X1 u5_mult_82_U5968 ( .A(u5_mult_82_n431), .B(u5_mult_82_n1988), .Z(
        u5_mult_82_SUMB_29__17_) );
  XOR2_X1 u5_mult_82_U5967 ( .A(u5_mult_82_ab_29__17_), .B(
        u5_mult_82_CARRYB_28__17_), .Z(u5_mult_82_n1988) );
  NAND3_X4 u5_mult_82_U5966 ( .A1(u5_mult_82_n1985), .A2(u5_mult_82_n1986), 
        .A3(u5_mult_82_n1987), .ZN(u5_mult_82_CARRYB_47__7_) );
  NAND2_X1 u5_mult_82_U5965 ( .A1(u5_mult_82_CARRYB_46__7_), .A2(
        u5_mult_82_SUMB_46__8_), .ZN(u5_mult_82_n1987) );
  NAND2_X1 u5_mult_82_U5964 ( .A1(u5_mult_82_ab_47__7_), .A2(
        u5_mult_82_SUMB_46__8_), .ZN(u5_mult_82_n1986) );
  NAND2_X1 u5_mult_82_U5963 ( .A1(u5_mult_82_ab_47__7_), .A2(
        u5_mult_82_CARRYB_46__7_), .ZN(u5_mult_82_n1985) );
  XOR2_X2 u5_mult_82_U5962 ( .A(u5_mult_82_n1984), .B(u5_mult_82_SUMB_46__8_), 
        .Z(u5_mult_82_SUMB_47__7_) );
  XOR2_X2 u5_mult_82_U5961 ( .A(u5_mult_82_ab_47__7_), .B(
        u5_mult_82_CARRYB_46__7_), .Z(u5_mult_82_n1984) );
  XOR2_X2 u5_mult_82_U5960 ( .A(u5_mult_82_n1983), .B(u5_mult_82_SUMB_45__9_), 
        .Z(u5_mult_82_SUMB_46__8_) );
  XOR2_X2 u5_mult_82_U5959 ( .A(u5_mult_82_ab_46__8_), .B(
        u5_mult_82_CARRYB_45__8_), .Z(u5_mult_82_n1983) );
  NAND2_X2 u5_mult_82_U5958 ( .A1(u5_mult_82_CARRYB_40__10_), .A2(
        u5_mult_82_SUMB_40__11_), .ZN(u5_mult_82_n1982) );
  NAND2_X2 u5_mult_82_U5957 ( .A1(u5_mult_82_ab_41__10_), .A2(
        u5_mult_82_SUMB_40__11_), .ZN(u5_mult_82_n1981) );
  NAND2_X1 u5_mult_82_U5956 ( .A1(u5_mult_82_ab_41__10_), .A2(
        u5_mult_82_CARRYB_40__10_), .ZN(u5_mult_82_n1980) );
  NAND3_X2 u5_mult_82_U5955 ( .A1(u5_mult_82_n1977), .A2(u5_mult_82_n1978), 
        .A3(u5_mult_82_n1979), .ZN(u5_mult_82_CARRYB_40__11_) );
  NAND2_X1 u5_mult_82_U5954 ( .A1(u5_mult_82_CARRYB_39__11_), .A2(
        u5_mult_82_SUMB_39__12_), .ZN(u5_mult_82_n1979) );
  NAND2_X1 u5_mult_82_U5953 ( .A1(u5_mult_82_ab_40__11_), .A2(
        u5_mult_82_SUMB_39__12_), .ZN(u5_mult_82_n1978) );
  NAND2_X1 u5_mult_82_U5952 ( .A1(u5_mult_82_ab_40__11_), .A2(
        u5_mult_82_CARRYB_39__11_), .ZN(u5_mult_82_n1977) );
  NAND2_X2 u5_mult_82_U5951 ( .A1(u5_mult_82_n733), .A2(
        u5_mult_82_SUMB_26__26_), .ZN(u5_mult_82_n6185) );
  NAND2_X2 u5_mult_82_U5950 ( .A1(u5_mult_82_CARRYB_31__22_), .A2(
        u5_mult_82_SUMB_31__23_), .ZN(u5_mult_82_n3525) );
  NAND2_X2 u5_mult_82_U5949 ( .A1(u5_mult_82_ab_25__26_), .A2(
        u5_mult_82_SUMB_24__27_), .ZN(u5_mult_82_n6145) );
  NAND2_X2 u5_mult_82_U5948 ( .A1(u5_mult_82_SUMB_24__27_), .A2(
        u5_mult_82_CARRYB_24__26_), .ZN(u5_mult_82_n6146) );
  NAND3_X4 u5_mult_82_U5947 ( .A1(u5_mult_82_n6144), .A2(u5_mult_82_n6145), 
        .A3(u5_mult_82_n6146), .ZN(u5_mult_82_CARRYB_25__26_) );
  XNOR2_X2 u5_mult_82_U5946 ( .A(u5_mult_82_ab_6__43_), .B(u5_mult_82_n1865), 
        .ZN(u5_mult_82_n2111) );
  NOR2_X1 u5_mult_82_U5945 ( .A1(u5_mult_82_net64489), .A2(u5_mult_82_n6616), 
        .ZN(u5_mult_82_ab_19__12_) );
  NOR2_X1 u5_mult_82_U5944 ( .A1(u5_mult_82_n6929), .A2(u5_mult_82_n6566), 
        .ZN(u5_mult_82_ab_12__17_) );
  NOR2_X1 u5_mult_82_U5943 ( .A1(u5_mult_82_net64379), .A2(u5_mult_82_n6686), 
        .ZN(u5_mult_82_ab_31__6_) );
  NOR2_X1 u5_mult_82_U5942 ( .A1(u5_mult_82_n6893), .A2(u5_mult_82_n6515), 
        .ZN(u5_mult_82_ab_3__24_) );
  NAND3_X2 u5_mult_82_U5941 ( .A1(u5_mult_82_n1974), .A2(u5_mult_82_n1975), 
        .A3(u5_mult_82_n1976), .ZN(u5_mult_82_CARRYB_19__12_) );
  NAND2_X1 u5_mult_82_U5940 ( .A1(u5_mult_82_SUMB_18__13_), .A2(
        u5_mult_82_ab_19__12_), .ZN(u5_mult_82_n1976) );
  NAND2_X2 u5_mult_82_U5939 ( .A1(u5_mult_82_ab_19__12_), .A2(
        u5_mult_82_CARRYB_18__12_), .ZN(u5_mult_82_n1975) );
  NAND2_X1 u5_mult_82_U5938 ( .A1(u5_mult_82_SUMB_18__13_), .A2(
        u5_mult_82_CARRYB_18__12_), .ZN(u5_mult_82_n1974) );
  XOR2_X2 u5_mult_82_U5937 ( .A(u5_mult_82_CARRYB_18__12_), .B(
        u5_mult_82_n1973), .Z(u5_mult_82_SUMB_19__12_) );
  XOR2_X2 u5_mult_82_U5936 ( .A(u5_mult_82_SUMB_18__13_), .B(
        u5_mult_82_ab_19__12_), .Z(u5_mult_82_n1973) );
  NAND3_X2 u5_mult_82_U5935 ( .A1(u5_mult_82_n1970), .A2(u5_mult_82_n1971), 
        .A3(u5_mult_82_n1972), .ZN(u5_mult_82_CARRYB_12__17_) );
  NAND2_X2 u5_mult_82_U5934 ( .A1(u5_mult_82_ab_12__17_), .A2(
        u5_mult_82_CARRYB_11__17_), .ZN(u5_mult_82_n1972) );
  NAND2_X1 u5_mult_82_U5933 ( .A1(u5_mult_82_CARRYB_11__17_), .A2(
        u5_mult_82_SUMB_11__18_), .ZN(u5_mult_82_n1970) );
  XOR2_X2 u5_mult_82_U5932 ( .A(u5_mult_82_CARRYB_11__17_), .B(
        u5_mult_82_ab_12__17_), .Z(u5_mult_82_n1969) );
  NAND3_X2 u5_mult_82_U5931 ( .A1(u5_mult_82_n1966), .A2(u5_mult_82_n1967), 
        .A3(u5_mult_82_n1968), .ZN(u5_mult_82_CARRYB_31__6_) );
  NAND2_X1 u5_mult_82_U5930 ( .A1(u5_mult_82_ab_31__6_), .A2(
        u5_mult_82_CARRYB_30__6_), .ZN(u5_mult_82_n1968) );
  NAND2_X2 u5_mult_82_U5929 ( .A1(u5_mult_82_ab_31__6_), .A2(
        u5_mult_82_SUMB_30__7_), .ZN(u5_mult_82_n1967) );
  NAND2_X1 u5_mult_82_U5928 ( .A1(u5_mult_82_CARRYB_30__6_), .A2(
        u5_mult_82_SUMB_30__7_), .ZN(u5_mult_82_n1966) );
  XOR2_X2 u5_mult_82_U5927 ( .A(u5_mult_82_n729), .B(u5_mult_82_n1965), .Z(
        u5_mult_82_SUMB_31__6_) );
  XOR2_X2 u5_mult_82_U5926 ( .A(u5_mult_82_CARRYB_30__6_), .B(
        u5_mult_82_ab_31__6_), .Z(u5_mult_82_n1965) );
  INV_X1 u5_mult_82_U5925 ( .A(u5_mult_82_SUMB_33__7_), .ZN(u5_mult_82_n1962)
         );
  NAND2_X2 u5_mult_82_U5924 ( .A1(u5_mult_82_n1963), .A2(u5_mult_82_n1964), 
        .ZN(u5_mult_82_SUMB_34__6_) );
  NAND2_X2 u5_mult_82_U5923 ( .A1(u5_mult_82_n1961), .A2(u5_mult_82_n1962), 
        .ZN(u5_mult_82_n1964) );
  NAND2_X2 u5_mult_82_U5922 ( .A1(u5_mult_82_n3108), .A2(
        u5_mult_82_SUMB_33__7_), .ZN(u5_mult_82_n1963) );
  NAND3_X2 u5_mult_82_U5921 ( .A1(u5_mult_82_n1958), .A2(u5_mult_82_n1959), 
        .A3(u5_mult_82_n1960), .ZN(u5_mult_82_CARRYB_5__22_) );
  NAND2_X1 u5_mult_82_U5920 ( .A1(u5_mult_82_ab_5__22_), .A2(
        u5_mult_82_SUMB_4__23_), .ZN(u5_mult_82_n1959) );
  NAND3_X2 u5_mult_82_U5919 ( .A1(u5_mult_82_n1955), .A2(u5_mult_82_n1956), 
        .A3(u5_mult_82_n1957), .ZN(u5_mult_82_CARRYB_4__23_) );
  NAND2_X2 u5_mult_82_U5918 ( .A1(u5_mult_82_CARRYB_3__23_), .A2(
        u5_mult_82_SUMB_3__24_), .ZN(u5_mult_82_n1957) );
  NAND2_X2 u5_mult_82_U5917 ( .A1(u5_mult_82_ab_4__23_), .A2(
        u5_mult_82_SUMB_3__24_), .ZN(u5_mult_82_n1956) );
  NAND2_X1 u5_mult_82_U5916 ( .A1(u5_mult_82_ab_4__23_), .A2(
        u5_mult_82_CARRYB_3__23_), .ZN(u5_mult_82_n1955) );
  XOR2_X2 u5_mult_82_U5915 ( .A(u5_mult_82_n1954), .B(u5_mult_82_SUMB_4__23_), 
        .Z(u5_mult_82_SUMB_5__22_) );
  XOR2_X2 u5_mult_82_U5914 ( .A(u5_mult_82_ab_5__22_), .B(
        u5_mult_82_CARRYB_4__22_), .Z(u5_mult_82_n1954) );
  XOR2_X2 u5_mult_82_U5913 ( .A(u5_mult_82_n1953), .B(u5_mult_82_SUMB_3__24_), 
        .Z(u5_mult_82_SUMB_4__23_) );
  XOR2_X2 u5_mult_82_U5912 ( .A(u5_mult_82_ab_4__23_), .B(
        u5_mult_82_CARRYB_3__23_), .Z(u5_mult_82_n1953) );
  NAND3_X2 u5_mult_82_U5911 ( .A1(u5_mult_82_n1950), .A2(u5_mult_82_n1951), 
        .A3(u5_mult_82_n1952), .ZN(u5_mult_82_CARRYB_3__24_) );
  NAND2_X1 u5_mult_82_U5910 ( .A1(u5_mult_82_ab_3__24_), .A2(
        u5_mult_82_CARRYB_2__24_), .ZN(u5_mult_82_n1952) );
  NAND2_X2 u5_mult_82_U5909 ( .A1(u5_mult_82_ab_3__24_), .A2(
        u5_mult_82_SUMB_2__25_), .ZN(u5_mult_82_n1951) );
  NAND2_X2 u5_mult_82_U5908 ( .A1(u5_mult_82_CARRYB_2__24_), .A2(
        u5_mult_82_SUMB_2__25_), .ZN(u5_mult_82_n1950) );
  XOR2_X2 u5_mult_82_U5907 ( .A(u5_mult_82_SUMB_2__25_), .B(u5_mult_82_n1949), 
        .Z(u5_mult_82_SUMB_3__24_) );
  XOR2_X2 u5_mult_82_U5906 ( .A(u5_mult_82_CARRYB_2__24_), .B(
        u5_mult_82_ab_3__24_), .Z(u5_mult_82_n1949) );
  XOR2_X2 u5_mult_82_U5905 ( .A(u5_mult_82_n4046), .B(u5_mult_82_SUMB_8__25_), 
        .Z(u5_mult_82_SUMB_9__24_) );
  NAND3_X2 u5_mult_82_U5904 ( .A1(u5_mult_82_n4914), .A2(u5_mult_82_n4915), 
        .A3(u5_mult_82_n4916), .ZN(u5_mult_82_CARRYB_39__31_) );
  XNOR2_X2 u5_mult_82_U5903 ( .A(u5_mult_82_n1948), .B(
        u5_mult_82_CARRYB_22__29_), .ZN(u5_mult_82_n3144) );
  NAND2_X1 u5_mult_82_U5902 ( .A1(u5_mult_82_ab_16__42_), .A2(
        u5_mult_82_CARRYB_15__42_), .ZN(u5_mult_82_n6222) );
  XNOR2_X2 u5_mult_82_U5901 ( .A(u5_mult_82_n1947), .B(
        u5_mult_82_CARRYB_33__32_), .ZN(u5_mult_82_n2716) );
  XNOR2_X2 u5_mult_82_U5900 ( .A(u5_mult_82_ab_17__42_), .B(
        u5_mult_82_CARRYB_16__42_), .ZN(u5_mult_82_n1946) );
  XNOR2_X1 u5_mult_82_U5899 ( .A(u5_mult_82_n1946), .B(u5_mult_82_SUMB_16__43_), .ZN(u5_mult_82_SUMB_17__42_) );
  XNOR2_X2 u5_mult_82_U5898 ( .A(u5_mult_82_CARRYB_24__37_), .B(
        u5_mult_82_ab_25__37_), .ZN(u5_mult_82_n1945) );
  XNOR2_X2 u5_mult_82_U5897 ( .A(u5_mult_82_SUMB_24__38_), .B(u5_mult_82_n1945), .ZN(u5_mult_82_SUMB_25__37_) );
  INV_X4 u5_mult_82_U5896 ( .A(u5_mult_82_SUMB_27__36_), .ZN(u5_mult_82_n2319)
         );
  INV_X4 u5_mult_82_U5895 ( .A(u5_mult_82_n2319), .ZN(u5_mult_82_n2320) );
  NAND2_X2 u5_mult_82_U5894 ( .A1(u5_mult_82_ab_5__27_), .A2(
        u5_mult_82_CARRYB_4__27_), .ZN(u5_mult_82_n3981) );
  NOR2_X1 u5_mult_82_U5893 ( .A1(u5_mult_82_n6882), .A2(u5_mult_82_net66019), 
        .ZN(u5_mult_82_ab_6__26_) );
  NOR2_X1 u5_mult_82_U5892 ( .A1(u5_mult_82_net64469), .A2(u5_mult_82_n6709), 
        .ZN(u5_mult_82_ab_35__11_) );
  NAND3_X2 u5_mult_82_U5891 ( .A1(u5_mult_82_n1942), .A2(u5_mult_82_n1943), 
        .A3(u5_mult_82_n1944), .ZN(u5_mult_82_CARRYB_6__26_) );
  NAND2_X1 u5_mult_82_U5890 ( .A1(u5_mult_82_ab_6__26_), .A2(
        u5_mult_82_CARRYB_5__26_), .ZN(u5_mult_82_n1944) );
  NAND2_X2 u5_mult_82_U5889 ( .A1(u5_mult_82_ab_6__26_), .A2(
        u5_mult_82_SUMB_5__27_), .ZN(u5_mult_82_n1943) );
  NAND2_X1 u5_mult_82_U5888 ( .A1(u5_mult_82_CARRYB_5__26_), .A2(
        u5_mult_82_SUMB_5__27_), .ZN(u5_mult_82_n1942) );
  NAND3_X2 u5_mult_82_U5887 ( .A1(u5_mult_82_n1939), .A2(u5_mult_82_n1940), 
        .A3(u5_mult_82_n1941), .ZN(u5_mult_82_CARRYB_35__11_) );
  NAND2_X1 u5_mult_82_U5886 ( .A1(u5_mult_82_ab_35__11_), .A2(
        u5_mult_82_CARRYB_34__11_), .ZN(u5_mult_82_n1941) );
  NAND2_X2 u5_mult_82_U5885 ( .A1(u5_mult_82_ab_35__11_), .A2(
        u5_mult_82_SUMB_34__12_), .ZN(u5_mult_82_n1940) );
  XNOR2_X2 u5_mult_82_U5884 ( .A(u5_mult_82_CARRYB_39__5_), .B(
        u5_mult_82_ab_40__5_), .ZN(u5_mult_82_n1938) );
  XNOR2_X2 u5_mult_82_U5883 ( .A(u5_mult_82_SUMB_39__6_), .B(u5_mult_82_n1938), 
        .ZN(u5_mult_82_SUMB_40__5_) );
  NAND3_X2 u5_mult_82_U5882 ( .A1(u5_mult_82_n5429), .A2(u5_mult_82_n5430), 
        .A3(u5_mult_82_n5431), .ZN(u5_mult_82_CARRYB_19__28_) );
  NAND2_X2 u5_mult_82_U5881 ( .A1(u5_mult_82_ab_15__30_), .A2(u5_mult_82_n1527), .ZN(u5_mult_82_n5683) );
  XNOR2_X2 u5_mult_82_U5880 ( .A(u5_mult_82_n1937), .B(u5_mult_82_SUMB_14__39_), .ZN(u5_mult_82_SUMB_15__38_) );
  XNOR2_X2 u5_mult_82_U5879 ( .A(u5_mult_82_ab_26__43_), .B(
        u5_mult_82_CARRYB_25__43_), .ZN(u5_mult_82_n1936) );
  XNOR2_X2 u5_mult_82_U5878 ( .A(u5_mult_82_n1936), .B(u5_mult_82_SUMB_25__44_), .ZN(u5_mult_82_SUMB_26__43_) );
  NAND3_X4 u5_mult_82_U5877 ( .A1(u5_mult_82_n5728), .A2(u5_mult_82_n5727), 
        .A3(u5_mult_82_n5726), .ZN(u5_mult_82_CARRYB_9__47_) );
  XNOR2_X2 u5_mult_82_U5876 ( .A(u5_mult_82_n3060), .B(u5_mult_82_n1622), .ZN(
        u5_mult_82_SUMB_27__23_) );
  NAND2_X2 u5_mult_82_U5875 ( .A1(u5_mult_82_ab_6__43_), .A2(u5_mult_82_n1865), 
        .ZN(u5_mult_82_n6061) );
  NAND2_X2 u5_mult_82_U5874 ( .A1(u5_mult_82_n1865), .A2(
        u5_mult_82_SUMB_5__44_), .ZN(u5_mult_82_n6063) );
  XNOR2_X2 u5_mult_82_U5873 ( .A(u5_mult_82_ab_33__4_), .B(
        u5_mult_82_CARRYB_32__4_), .ZN(u5_mult_82_n1935) );
  XNOR2_X2 u5_mult_82_U5872 ( .A(u5_mult_82_n1935), .B(u5_mult_82_SUMB_32__5_), 
        .ZN(u5_mult_82_SUMB_33__4_) );
  NAND3_X4 u5_mult_82_U5871 ( .A1(u5_mult_82_n4729), .A2(u5_mult_82_n4730), 
        .A3(u5_mult_82_n4731), .ZN(u5_mult_82_CARRYB_42__4_) );
  NAND2_X2 u5_mult_82_U5870 ( .A1(u5_mult_82_ab_24__23_), .A2(
        u5_mult_82_SUMB_23__24_), .ZN(u5_mult_82_n3059) );
  NAND2_X1 u5_mult_82_U5869 ( .A1(u5_mult_82_ab_3__46_), .A2(
        u5_mult_82_SUMB_2__47_), .ZN(u5_mult_82_n1933) );
  NAND2_X2 u5_mult_82_U5868 ( .A1(u5_mult_82_CARRYB_1__47_), .A2(
        u5_mult_82_SUMB_1__48_), .ZN(u5_mult_82_n1931) );
  NAND2_X2 u5_mult_82_U5867 ( .A1(u5_mult_82_ab_2__47_), .A2(
        u5_mult_82_SUMB_1__48_), .ZN(u5_mult_82_n1930) );
  NAND2_X1 u5_mult_82_U5866 ( .A1(u5_mult_82_ab_2__47_), .A2(
        u5_mult_82_CARRYB_1__47_), .ZN(u5_mult_82_n1929) );
  XOR2_X2 u5_mult_82_U5865 ( .A(u5_mult_82_ab_3__46_), .B(
        u5_mult_82_CARRYB_2__46_), .Z(u5_mult_82_n1928) );
  XOR2_X2 u5_mult_82_U5864 ( .A(u5_mult_82_n1927), .B(u5_mult_82_SUMB_1__48_), 
        .Z(u5_mult_82_SUMB_2__47_) );
  XOR2_X2 u5_mult_82_U5863 ( .A(u5_mult_82_ab_2__47_), .B(
        u5_mult_82_CARRYB_1__47_), .Z(u5_mult_82_n1927) );
  NAND3_X2 u5_mult_82_U5862 ( .A1(u5_mult_82_n1924), .A2(u5_mult_82_n1925), 
        .A3(u5_mult_82_n1926), .ZN(u5_mult_82_CARRYB_12__40_) );
  NAND2_X1 u5_mult_82_U5861 ( .A1(u5_mult_82_CARRYB_11__40_), .A2(
        u5_mult_82_SUMB_11__41_), .ZN(u5_mult_82_n1926) );
  NAND2_X1 u5_mult_82_U5860 ( .A1(u5_mult_82_ab_12__40_), .A2(
        u5_mult_82_SUMB_11__41_), .ZN(u5_mult_82_n1925) );
  NAND2_X1 u5_mult_82_U5859 ( .A1(u5_mult_82_ab_12__40_), .A2(
        u5_mult_82_CARRYB_11__40_), .ZN(u5_mult_82_n1924) );
  NAND3_X2 u5_mult_82_U5858 ( .A1(u5_mult_82_n1921), .A2(u5_mult_82_n1922), 
        .A3(u5_mult_82_n1923), .ZN(u5_mult_82_CARRYB_11__41_) );
  NAND2_X2 u5_mult_82_U5857 ( .A1(u5_mult_82_CARRYB_10__41_), .A2(
        u5_mult_82_SUMB_10__42_), .ZN(u5_mult_82_n1923) );
  NAND2_X2 u5_mult_82_U5856 ( .A1(u5_mult_82_ab_11__41_), .A2(
        u5_mult_82_SUMB_10__42_), .ZN(u5_mult_82_n1922) );
  NAND2_X1 u5_mult_82_U5855 ( .A1(u5_mult_82_ab_11__41_), .A2(
        u5_mult_82_CARRYB_10__41_), .ZN(u5_mult_82_n1921) );
  XOR2_X2 u5_mult_82_U5854 ( .A(u5_mult_82_n1920), .B(u5_mult_82_SUMB_11__41_), 
        .Z(u5_mult_82_SUMB_12__40_) );
  XOR2_X2 u5_mult_82_U5853 ( .A(u5_mult_82_ab_12__40_), .B(
        u5_mult_82_CARRYB_11__40_), .Z(u5_mult_82_n1920) );
  XOR2_X2 u5_mult_82_U5852 ( .A(u5_mult_82_n1919), .B(u5_mult_82_SUMB_10__42_), 
        .Z(u5_mult_82_SUMB_11__41_) );
  XOR2_X2 u5_mult_82_U5851 ( .A(u5_mult_82_ab_11__41_), .B(
        u5_mult_82_CARRYB_10__41_), .Z(u5_mult_82_n1919) );
  INV_X4 u5_mult_82_U5850 ( .A(u5_mult_82_CARRYB_17__35_), .ZN(
        u5_mult_82_n1916) );
  NAND2_X2 u5_mult_82_U5849 ( .A1(u5_mult_82_n1917), .A2(u5_mult_82_n1918), 
        .ZN(u5_mult_82_n6309) );
  NAND2_X2 u5_mult_82_U5848 ( .A1(u5_mult_82_ab_18__35_), .A2(u5_mult_82_n1916), .ZN(u5_mult_82_n1918) );
  NAND2_X1 u5_mult_82_U5847 ( .A1(u5_mult_82_n3153), .A2(
        u5_mult_82_CARRYB_17__35_), .ZN(u5_mult_82_n1917) );
  NAND2_X2 u5_mult_82_U5846 ( .A1(u5_mult_82_ab_28__5_), .A2(
        u5_mult_82_CARRYB_27__5_), .ZN(u5_mult_82_n4056) );
  XNOR2_X2 u5_mult_82_U5845 ( .A(u5_mult_82_CARRYB_28__10_), .B(
        u5_mult_82_ab_29__10_), .ZN(u5_mult_82_n1915) );
  XNOR2_X2 u5_mult_82_U5844 ( .A(u5_mult_82_n1915), .B(u5_mult_82_SUMB_28__11_), .ZN(u5_mult_82_SUMB_29__10_) );
  NAND2_X2 u5_mult_82_U5843 ( .A1(u5_mult_82_n1496), .A2(u5_mult_82_n3825), 
        .ZN(u5_mult_82_n5951) );
  NAND2_X2 u5_mult_82_U5842 ( .A1(u5_mult_82_ab_21__25_), .A2(
        u5_mult_82_CARRYB_20__25_), .ZN(u5_mult_82_n2189) );
  NAND3_X2 u5_mult_82_U5841 ( .A1(u5_mult_82_n2189), .A2(u5_mult_82_n2190), 
        .A3(u5_mult_82_n2191), .ZN(u5_mult_82_CARRYB_21__25_) );
  XNOR2_X2 u5_mult_82_U5840 ( .A(u5_mult_82_n1914), .B(
        u5_mult_82_CARRYB_45__27_), .ZN(u5_mult_82_n4569) );
  XNOR2_X2 u5_mult_82_U5839 ( .A(u5_mult_82_n1913), .B(u5_mult_82_n1782), .ZN(
        u5_mult_82_SUMB_15__46_) );
  XNOR2_X2 u5_mult_82_U5838 ( .A(u5_mult_82_n1912), .B(u5_mult_82_n1657), .ZN(
        u5_mult_82_n2787) );
  NAND2_X1 u5_mult_82_U5837 ( .A1(u5_mult_82_ab_7__42_), .A2(
        u5_mult_82_CARRYB_6__42_), .ZN(u5_mult_82_n5976) );
  NAND2_X2 u5_mult_82_U5836 ( .A1(u5_mult_82_ab_25__32_), .A2(
        u5_mult_82_SUMB_24__33_), .ZN(u5_mult_82_n5475) );
  NAND3_X2 u5_mult_82_U5835 ( .A1(u5_mult_82_n4573), .A2(u5_mult_82_n4574), 
        .A3(u5_mult_82_n4575), .ZN(u5_mult_82_CARRYB_46__27_) );
  NAND3_X4 u5_mult_82_U5834 ( .A1(u5_mult_82_net86288), .A2(
        u5_mult_82_net86289), .A3(u5_mult_82_net86290), .ZN(
        u5_mult_82_CARRYB_41__12_) );
  NAND3_X2 u5_mult_82_U5833 ( .A1(u5_mult_82_n1910), .A2(u5_mult_82_n1909), 
        .A3(u5_mult_82_n1911), .ZN(u5_mult_82_CARRYB_40__13_) );
  NAND2_X1 u5_mult_82_U5832 ( .A1(u5_mult_82_ab_40__13_), .A2(
        u5_mult_82_CARRYB_39__13_), .ZN(u5_mult_82_n1909) );
  INV_X4 u5_mult_82_U5831 ( .A(u5_mult_82_CARRYB_20__37_), .ZN(
        u5_mult_82_n4530) );
  XNOR2_X2 u5_mult_82_U5830 ( .A(u5_mult_82_n1908), .B(u5_mult_82_SUMB_37__3_), 
        .ZN(u5_mult_82_SUMB_38__2_) );
  XNOR2_X2 u5_mult_82_U5829 ( .A(u5_mult_82_n1907), .B(
        u5_mult_82_CARRYB_28__32_), .ZN(u5_mult_82_n2423) );
  NAND2_X2 u5_mult_82_U5828 ( .A1(u5_mult_82_net88030), .A2(
        u5_mult_82_SUMB_23__24_), .ZN(u5_mult_82_n3058) );
  NAND2_X2 u5_mult_82_U5827 ( .A1(u5_mult_82_ab_41__5_), .A2(
        u5_mult_82_SUMB_40__6_), .ZN(u5_mult_82_n4727) );
  XNOR2_X2 u5_mult_82_U5826 ( .A(u5_mult_82_n5161), .B(u5_mult_82_n374), .ZN(
        u5_mult_82_SUMB_40__6_) );
  NAND2_X2 u5_mult_82_U5825 ( .A1(u5_mult_82_ab_16__46_), .A2(
        u5_mult_82_SUMB_15__47_), .ZN(u5_mult_82_n4613) );
  NAND2_X1 u5_mult_82_U5824 ( .A1(u5_mult_82_ab_50__22_), .A2(
        u5_mult_82_CARRYB_49__22_), .ZN(u5_mult_82_n5099) );
  NAND3_X2 u5_mult_82_U5823 ( .A1(u5_mult_82_n2788), .A2(u5_mult_82_n2789), 
        .A3(u5_mult_82_n2790), .ZN(u5_mult_82_CARRYB_28__14_) );
  NAND2_X2 u5_mult_82_U5822 ( .A1(u5_mult_82_ab_23__36_), .A2(
        u5_mult_82_SUMB_22__37_), .ZN(u5_mult_82_n5739) );
  NOR2_X4 u5_mult_82_U5821 ( .A1(u5_mult_82_n6852), .A2(u5_mult_82_n6586), 
        .ZN(u5_mult_82_ab_15__31_) );
  NAND2_X1 u5_mult_82_U5820 ( .A1(u5_mult_82_ab_23__26_), .A2(
        u5_mult_82_CARRYB_22__26_), .ZN(u5_mult_82_n1903) );
  NAND3_X2 u5_mult_82_U5819 ( .A1(u5_mult_82_n1900), .A2(u5_mult_82_n1901), 
        .A3(u5_mult_82_n1902), .ZN(u5_mult_82_CARRYB_22__27_) );
  NAND2_X1 u5_mult_82_U5818 ( .A1(u5_mult_82_CARRYB_21__27_), .A2(
        u5_mult_82_SUMB_21__28_), .ZN(u5_mult_82_n1902) );
  NAND2_X1 u5_mult_82_U5817 ( .A1(u5_mult_82_ab_22__27_), .A2(
        u5_mult_82_SUMB_21__28_), .ZN(u5_mult_82_n1901) );
  NAND2_X1 u5_mult_82_U5816 ( .A1(u5_mult_82_ab_22__27_), .A2(
        u5_mult_82_CARRYB_21__27_), .ZN(u5_mult_82_n1900) );
  INV_X1 u5_mult_82_U5815 ( .A(u5_mult_82_ab_15__31_), .ZN(u5_mult_82_n1897)
         );
  INV_X4 u5_mult_82_U5814 ( .A(u5_mult_82_CARRYB_14__31_), .ZN(
        u5_mult_82_n1896) );
  NAND2_X4 u5_mult_82_U5813 ( .A1(u5_mult_82_n1898), .A2(u5_mult_82_n1899), 
        .ZN(u5_mult_82_n2017) );
  NAND2_X2 u5_mult_82_U5812 ( .A1(u5_mult_82_n1896), .A2(u5_mult_82_n1897), 
        .ZN(u5_mult_82_n1899) );
  NAND2_X2 u5_mult_82_U5811 ( .A1(u5_mult_82_CARRYB_14__31_), .A2(
        u5_mult_82_ab_15__31_), .ZN(u5_mult_82_n1898) );
  NOR2_X1 u5_mult_82_U5810 ( .A1(u5_mult_82_net64363), .A2(u5_mult_82_n6637), 
        .ZN(u5_mult_82_ab_22__5_) );
  NOR2_X1 u5_mult_82_U5809 ( .A1(u5_mult_82_net64363), .A2(u5_mult_82_n6630), 
        .ZN(u5_mult_82_ab_21__5_) );
  NOR2_X1 u5_mult_82_U5808 ( .A1(u5_mult_82_n6906), .A2(u5_mult_82_n6522), 
        .ZN(u5_mult_82_ab_4__20_) );
  NAND3_X2 u5_mult_82_U5807 ( .A1(u5_mult_82_n1893), .A2(u5_mult_82_n1894), 
        .A3(u5_mult_82_n1895), .ZN(u5_mult_82_CARRYB_33__5_) );
  NAND2_X1 u5_mult_82_U5806 ( .A1(u5_mult_82_SUMB_32__6_), .A2(
        u5_mult_82_CARRYB_32__5_), .ZN(u5_mult_82_n1895) );
  NAND2_X2 u5_mult_82_U5805 ( .A1(u5_mult_82_ab_33__5_), .A2(
        u5_mult_82_CARRYB_32__5_), .ZN(u5_mult_82_n1894) );
  NAND2_X1 u5_mult_82_U5804 ( .A1(u5_mult_82_ab_33__5_), .A2(
        u5_mult_82_SUMB_32__6_), .ZN(u5_mult_82_n1893) );
  XOR2_X2 u5_mult_82_U5803 ( .A(u5_mult_82_n1892), .B(u5_mult_82_CARRYB_32__5_), .Z(u5_mult_82_SUMB_33__5_) );
  XOR2_X2 u5_mult_82_U5802 ( .A(u5_mult_82_ab_33__5_), .B(
        u5_mult_82_SUMB_32__6_), .Z(u5_mult_82_n1892) );
  NAND3_X2 u5_mult_82_U5801 ( .A1(u5_mult_82_n1889), .A2(u5_mult_82_n1890), 
        .A3(u5_mult_82_n1891), .ZN(u5_mult_82_CARRYB_32__5_) );
  NAND2_X1 u5_mult_82_U5800 ( .A1(u5_mult_82_SUMB_31__6_), .A2(
        u5_mult_82_CARRYB_31__5_), .ZN(u5_mult_82_n1891) );
  NAND2_X2 u5_mult_82_U5799 ( .A1(u5_mult_82_ab_32__5_), .A2(
        u5_mult_82_CARRYB_31__5_), .ZN(u5_mult_82_n1890) );
  NAND2_X1 u5_mult_82_U5798 ( .A1(u5_mult_82_ab_32__5_), .A2(
        u5_mult_82_SUMB_31__6_), .ZN(u5_mult_82_n1889) );
  XOR2_X2 u5_mult_82_U5797 ( .A(u5_mult_82_n1888), .B(u5_mult_82_CARRYB_31__5_), .Z(u5_mult_82_SUMB_32__5_) );
  XOR2_X2 u5_mult_82_U5796 ( .A(u5_mult_82_ab_32__5_), .B(
        u5_mult_82_SUMB_31__6_), .Z(u5_mult_82_n1888) );
  NAND3_X2 u5_mult_82_U5795 ( .A1(u5_mult_82_n1885), .A2(u5_mult_82_n1886), 
        .A3(u5_mult_82_n1887), .ZN(u5_mult_82_CARRYB_22__5_) );
  NAND2_X1 u5_mult_82_U5794 ( .A1(u5_mult_82_ab_22__5_), .A2(
        u5_mult_82_CARRYB_21__5_), .ZN(u5_mult_82_n1887) );
  NAND2_X2 u5_mult_82_U5793 ( .A1(u5_mult_82_ab_22__5_), .A2(
        u5_mult_82_SUMB_21__6_), .ZN(u5_mult_82_n1886) );
  NAND2_X1 u5_mult_82_U5792 ( .A1(u5_mult_82_CARRYB_21__5_), .A2(
        u5_mult_82_SUMB_21__6_), .ZN(u5_mult_82_n1885) );
  XOR2_X2 u5_mult_82_U5791 ( .A(u5_mult_82_SUMB_21__6_), .B(u5_mult_82_n1884), 
        .Z(u5_mult_82_SUMB_22__5_) );
  XOR2_X2 u5_mult_82_U5790 ( .A(u5_mult_82_CARRYB_21__5_), .B(
        u5_mult_82_ab_22__5_), .Z(u5_mult_82_n1884) );
  NAND3_X2 u5_mult_82_U5789 ( .A1(u5_mult_82_n1881), .A2(u5_mult_82_n1882), 
        .A3(u5_mult_82_n1883), .ZN(u5_mult_82_CARRYB_21__5_) );
  NAND2_X1 u5_mult_82_U5788 ( .A1(u5_mult_82_ab_21__5_), .A2(
        u5_mult_82_CARRYB_20__5_), .ZN(u5_mult_82_n1883) );
  NAND2_X2 u5_mult_82_U5787 ( .A1(u5_mult_82_ab_21__5_), .A2(
        u5_mult_82_SUMB_20__6_), .ZN(u5_mult_82_n1882) );
  NAND2_X1 u5_mult_82_U5786 ( .A1(u5_mult_82_CARRYB_20__5_), .A2(
        u5_mult_82_SUMB_20__6_), .ZN(u5_mult_82_n1881) );
  NAND3_X2 u5_mult_82_U5785 ( .A1(u5_mult_82_n1878), .A2(u5_mult_82_n1879), 
        .A3(u5_mult_82_n1880), .ZN(u5_mult_82_CARRYB_6__18_) );
  NAND2_X1 u5_mult_82_U5784 ( .A1(u5_mult_82_CARRYB_5__18_), .A2(
        u5_mult_82_SUMB_5__19_), .ZN(u5_mult_82_n1880) );
  NAND2_X1 u5_mult_82_U5783 ( .A1(u5_mult_82_ab_6__18_), .A2(
        u5_mult_82_SUMB_5__19_), .ZN(u5_mult_82_n1879) );
  NAND2_X1 u5_mult_82_U5782 ( .A1(u5_mult_82_ab_6__18_), .A2(
        u5_mult_82_CARRYB_5__18_), .ZN(u5_mult_82_n1878) );
  NAND3_X2 u5_mult_82_U5781 ( .A1(u5_mult_82_n1875), .A2(u5_mult_82_n1876), 
        .A3(u5_mult_82_n1877), .ZN(u5_mult_82_CARRYB_5__19_) );
  NAND2_X2 u5_mult_82_U5780 ( .A1(u5_mult_82_CARRYB_4__19_), .A2(
        u5_mult_82_SUMB_4__20_), .ZN(u5_mult_82_n1877) );
  NAND2_X2 u5_mult_82_U5779 ( .A1(u5_mult_82_ab_5__19_), .A2(
        u5_mult_82_SUMB_4__20_), .ZN(u5_mult_82_n1876) );
  NAND2_X1 u5_mult_82_U5778 ( .A1(u5_mult_82_ab_5__19_), .A2(
        u5_mult_82_CARRYB_4__19_), .ZN(u5_mult_82_n1875) );
  XOR2_X2 u5_mult_82_U5777 ( .A(u5_mult_82_n1874), .B(u5_mult_82_SUMB_5__19_), 
        .Z(u5_mult_82_SUMB_6__18_) );
  XOR2_X2 u5_mult_82_U5776 ( .A(u5_mult_82_ab_6__18_), .B(
        u5_mult_82_CARRYB_5__18_), .Z(u5_mult_82_n1874) );
  XOR2_X2 u5_mult_82_U5775 ( .A(u5_mult_82_n1873), .B(u5_mult_82_SUMB_4__20_), 
        .Z(u5_mult_82_SUMB_5__19_) );
  XOR2_X2 u5_mult_82_U5774 ( .A(u5_mult_82_ab_5__19_), .B(
        u5_mult_82_CARRYB_4__19_), .Z(u5_mult_82_n1873) );
  NAND3_X2 u5_mult_82_U5773 ( .A1(u5_mult_82_n1870), .A2(u5_mult_82_n1871), 
        .A3(u5_mult_82_n1872), .ZN(u5_mult_82_CARRYB_4__20_) );
  NAND2_X1 u5_mult_82_U5772 ( .A1(u5_mult_82_ab_4__20_), .A2(
        u5_mult_82_CARRYB_3__20_), .ZN(u5_mult_82_n1872) );
  NAND2_X2 u5_mult_82_U5771 ( .A1(u5_mult_82_ab_4__20_), .A2(
        u5_mult_82_SUMB_3__21_), .ZN(u5_mult_82_n1871) );
  NAND2_X1 u5_mult_82_U5770 ( .A1(u5_mult_82_CARRYB_3__20_), .A2(
        u5_mult_82_SUMB_3__21_), .ZN(u5_mult_82_n1870) );
  XOR2_X2 u5_mult_82_U5769 ( .A(u5_mult_82_SUMB_3__21_), .B(u5_mult_82_n1869), 
        .Z(u5_mult_82_SUMB_4__20_) );
  XOR2_X2 u5_mult_82_U5768 ( .A(u5_mult_82_CARRYB_3__20_), .B(
        u5_mult_82_ab_4__20_), .Z(u5_mult_82_n1869) );
  XNOR2_X2 u5_mult_82_U5767 ( .A(u5_mult_82_n1728), .B(u5_mult_82_n1867), .ZN(
        u5_mult_82_SUMB_18__45_) );
  INV_X2 u5_mult_82_U5766 ( .A(u5_mult_82_n2012), .ZN(u5_mult_82_n1866) );
  INV_X8 u5_mult_82_U5765 ( .A(u5_mult_82_n1864), .ZN(u5_mult_82_n1865) );
  INV_X4 u5_mult_82_U5764 ( .A(u5_mult_82_CARRYB_5__43_), .ZN(u5_mult_82_n1864) );
  INV_X4 u5_mult_82_U5763 ( .A(u5_mult_82_n1862), .ZN(u5_mult_82_n1863) );
  INV_X2 u5_mult_82_U5762 ( .A(u5_mult_82_SUMB_46__21_), .ZN(u5_mult_82_n1862)
         );
  CLKBUF_X2 u5_mult_82_U5761 ( .A(u5_mult_82_SUMB_4__50_), .Z(u5_mult_82_n1861) );
  INV_X4 u5_mult_82_U5760 ( .A(u5_mult_82_n1858), .ZN(u5_mult_82_n1859) );
  INV_X2 u5_mult_82_U5759 ( .A(u5_mult_82_SUMB_14__37_), .ZN(u5_mult_82_n1858)
         );
  INV_X2 u5_mult_82_U5758 ( .A(u5_mult_82_SUMB_36__30_), .ZN(u5_mult_82_n1856)
         );
  XNOR2_X2 u5_mult_82_U5757 ( .A(u5_mult_82_SUMB_38__3_), .B(u5_mult_82_n1855), 
        .ZN(u5_mult_82_SUMB_39__2_) );
  CLKBUF_X3 u5_mult_82_U5756 ( .A(u5_mult_82_SUMB_37__10_), .Z(
        u5_mult_82_n1854) );
  INV_X4 u5_mult_82_U5755 ( .A(u5_mult_82_n1852), .ZN(u5_mult_82_n1853) );
  INV_X2 u5_mult_82_U5754 ( .A(u5_mult_82_SUMB_8__46_), .ZN(u5_mult_82_n1852)
         );
  INV_X4 u5_mult_82_U5753 ( .A(u5_mult_82_n1849), .ZN(u5_mult_82_n1850) );
  INV_X2 u5_mult_82_U5752 ( .A(u5_mult_82_SUMB_37__32_), .ZN(u5_mult_82_n1849)
         );
  INV_X4 u5_mult_82_U5751 ( .A(u5_mult_82_n1847), .ZN(u5_mult_82_n1848) );
  INV_X2 u5_mult_82_U5750 ( .A(u5_mult_82_SUMB_27__14_), .ZN(u5_mult_82_n1847)
         );
  CLKBUF_X2 u5_mult_82_U5749 ( .A(u5_mult_82_SUMB_32__42_), .Z(
        u5_mult_82_n1846) );
  NAND3_X2 u5_mult_82_U5748 ( .A1(u5_mult_82_n2442), .A2(u5_mult_82_n2443), 
        .A3(u5_mult_82_n2444), .ZN(u5_mult_82_CARRYB_47__29_) );
  CLKBUF_X2 u5_mult_82_U5747 ( .A(u5_mult_82_SUMB_48__16_), .Z(
        u5_mult_82_n1845) );
  CLKBUF_X2 u5_mult_82_U5746 ( .A(u5_mult_82_SUMB_40__26_), .Z(
        u5_mult_82_n1844) );
  INV_X4 u5_mult_82_U5745 ( .A(u5_mult_82_n1838), .ZN(u5_mult_82_n1839) );
  INV_X2 u5_mult_82_U5744 ( .A(u5_mult_82_SUMB_30__13_), .ZN(u5_mult_82_n1838)
         );
  INV_X1 u5_mult_82_U5743 ( .A(u5_mult_82_n5282), .ZN(u5_mult_82_n1837) );
  FA_X1 u5_mult_82_U5742 ( .A(u5_mult_82_ab_4__51_), .B(u5_mult_82_ab_3__52_), 
        .CI(u5_mult_82_n1495), .CO(u5_mult_82_n1834) );
  INV_X4 u5_mult_82_U5741 ( .A(u5_mult_82_SUMB_44__3_), .ZN(u5_mult_82_n1832)
         );
  XNOR2_X2 u5_mult_82_U5740 ( .A(u5_mult_82_ab_32__26_), .B(
        u5_mult_82_CARRYB_31__26_), .ZN(u5_mult_82_n1831) );
  XNOR2_X2 u5_mult_82_U5739 ( .A(u5_mult_82_n1500), .B(u5_mult_82_n1831), .ZN(
        u5_mult_82_SUMB_32__26_) );
  XNOR2_X2 u5_mult_82_U5738 ( .A(u5_mult_82_CARRYB_34__11_), .B(
        u5_mult_82_ab_35__11_), .ZN(u5_mult_82_n1830) );
  XNOR2_X2 u5_mult_82_U5737 ( .A(u5_mult_82_SUMB_34__12_), .B(u5_mult_82_n1830), .ZN(u5_mult_82_SUMB_35__11_) );
  INV_X8 u5_mult_82_U5736 ( .A(u5_mult_82_n1828), .ZN(u5_mult_82_n1829) );
  INV_X4 u5_mult_82_U5735 ( .A(u5_mult_82_SUMB_15__20_), .ZN(u5_mult_82_n1828)
         );
  NAND2_X1 u5_mult_82_U5734 ( .A1(u5_mult_82_CARRYB_47__12_), .A2(
        u5_mult_82_n1655), .ZN(u5_mult_82_n6110) );
  NAND2_X1 u5_mult_82_U5733 ( .A1(u5_mult_82_ab_48__12_), .A2(u5_mult_82_n1655), .ZN(u5_mult_82_n6109) );
  INV_X2 u5_mult_82_U5732 ( .A(u5_mult_82_SUMB_47__30_), .ZN(u5_mult_82_n1825)
         );
  XOR2_X2 u5_mult_82_U5731 ( .A(u5_mult_82_ab_49__31_), .B(
        u5_mult_82_CARRYB_48__31_), .Z(u5_mult_82_n2936) );
  INV_X2 u5_mult_82_U5730 ( .A(u5_mult_82_SUMB_5__48_), .ZN(u5_mult_82_n1821)
         );
  XNOR2_X2 u5_mult_82_U5729 ( .A(u5_mult_82_ab_41__15_), .B(
        u5_mult_82_CARRYB_40__15_), .ZN(u5_mult_82_n1819) );
  NAND3_X2 u5_mult_82_U5728 ( .A1(u5_mult_82_n6271), .A2(u5_mult_82_n6272), 
        .A3(u5_mult_82_n6273), .ZN(u5_mult_82_CARRYB_30__26_) );
  CLKBUF_X2 u5_mult_82_U5727 ( .A(u5_mult_82_SUMB_28__26_), .Z(
        u5_mult_82_n1816) );
  INV_X4 u5_mult_82_U5726 ( .A(u5_mult_82_n1814), .ZN(u5_mult_82_n1815) );
  XNOR2_X2 u5_mult_82_U5725 ( .A(u5_mult_82_ab_37__31_), .B(
        u5_mult_82_CARRYB_36__31_), .ZN(u5_mult_82_n1813) );
  XNOR2_X2 u5_mult_82_U5724 ( .A(u5_mult_82_n1813), .B(u5_mult_82_SUMB_36__32_), .ZN(u5_mult_82_SUMB_37__31_) );
  INV_X4 u5_mult_82_U5723 ( .A(u5_mult_82_n1811), .ZN(u5_mult_82_n1812) );
  INV_X2 u5_mult_82_U5722 ( .A(u5_mult_82_SUMB_38__25_), .ZN(u5_mult_82_n1811)
         );
  XOR2_X2 u5_mult_82_U5721 ( .A(u5_mult_82_n2958), .B(u5_mult_82_SUMB_47__32_), 
        .Z(u5_mult_82_SUMB_48__31_) );
  INV_X4 u5_mult_82_U5720 ( .A(u5_mult_82_n482), .ZN(u5_mult_82_n1810) );
  INV_X2 u5_mult_82_U5719 ( .A(u5_mult_82_n1807), .ZN(u5_mult_82_n1808) );
  XNOR2_X2 u5_mult_82_U5718 ( .A(u5_mult_82_ab_23__32_), .B(
        u5_mult_82_CARRYB_22__32_), .ZN(u5_mult_82_n1806) );
  XNOR2_X2 u5_mult_82_U5717 ( .A(u5_mult_82_n1806), .B(u5_mult_82_n1553), .ZN(
        u5_mult_82_SUMB_23__32_) );
  XNOR2_X2 u5_mult_82_U5716 ( .A(u5_mult_82_n1805), .B(u5_mult_82_n1462), .ZN(
        u5_mult_82_SUMB_7__42_) );
  XNOR2_X2 u5_mult_82_U5715 ( .A(u5_mult_82_n1804), .B(
        u5_mult_82_CARRYB_16__31_), .ZN(u5_mult_82_SUMB_17__31_) );
  XNOR2_X2 u5_mult_82_U5714 ( .A(u5_mult_82_ab_33__32_), .B(
        u5_mult_82_CARRYB_32__32_), .ZN(u5_mult_82_n1803) );
  XNOR2_X2 u5_mult_82_U5713 ( .A(u5_mult_82_n1803), .B(u5_mult_82_n72), .ZN(
        u5_mult_82_SUMB_33__32_) );
  XNOR2_X2 u5_mult_82_U5712 ( .A(u5_mult_82_CARRYB_19__41_), .B(
        u5_mult_82_ab_20__41_), .ZN(u5_mult_82_n1802) );
  XNOR2_X2 u5_mult_82_U5711 ( .A(u5_mult_82_n1802), .B(u5_mult_82_SUMB_19__42_), .ZN(u5_mult_82_SUMB_20__41_) );
  XNOR2_X2 u5_mult_82_U5710 ( .A(u5_mult_82_n1801), .B(u5_mult_82_SUMB_4__28_), 
        .ZN(u5_mult_82_SUMB_5__27_) );
  INV_X4 u5_mult_82_U5709 ( .A(u5_mult_82_n1799), .ZN(u5_mult_82_n1800) );
  XNOR2_X2 u5_mult_82_U5708 ( .A(u5_mult_82_n1798), .B(
        u5_mult_82_CARRYB_24__16_), .ZN(u5_mult_82_n2990) );
  INV_X8 u5_mult_82_U5707 ( .A(u5_mult_82_n1796), .ZN(u5_mult_82_n1797) );
  INV_X4 u5_mult_82_U5706 ( .A(u5_mult_82_SUMB_24__14_), .ZN(u5_mult_82_n1796)
         );
  INV_X4 u5_mult_82_U5705 ( .A(u5_mult_82_n1793), .ZN(u5_mult_82_n1794) );
  INV_X2 u5_mult_82_U5704 ( .A(u5_mult_82_SUMB_13__43_), .ZN(u5_mult_82_n1793)
         );
  XNOR2_X2 u5_mult_82_U5703 ( .A(u5_mult_82_ab_47__11_), .B(
        u5_mult_82_CARRYB_46__11_), .ZN(u5_mult_82_n1792) );
  XNOR2_X2 u5_mult_82_U5702 ( .A(u5_mult_82_n1792), .B(u5_mult_82_SUMB_46__12_), .ZN(u5_mult_82_SUMB_47__11_) );
  INV_X4 u5_mult_82_U5701 ( .A(u5_mult_82_n1790), .ZN(u5_mult_82_n1791) );
  INV_X2 u5_mult_82_U5700 ( .A(u5_mult_82_SUMB_21__31_), .ZN(u5_mult_82_n1790)
         );
  XOR2_X2 u5_mult_82_U5699 ( .A(u5_mult_82_n5201), .B(
        u5_mult_82_CARRYB_47__12_), .Z(u5_mult_82_n1789) );
  XNOR2_X2 u5_mult_82_U5698 ( .A(u5_mult_82_n1789), .B(u5_mult_82_SUMB_47__13_), .ZN(u5_mult_82_SUMB_48__12_) );
  INV_X4 u5_mult_82_U5697 ( .A(u5_mult_82_n1787), .ZN(u5_mult_82_n1788) );
  INV_X2 u5_mult_82_U5696 ( .A(u5_mult_82_SUMB_20__39_), .ZN(u5_mult_82_n1787)
         );
  NAND3_X2 u5_mult_82_U5695 ( .A1(u5_mult_82_n6175), .A2(u5_mult_82_n6174), 
        .A3(u5_mult_82_n6173), .ZN(u5_mult_82_CARRYB_36__16_) );
  NAND2_X1 u5_mult_82_U5694 ( .A1(u5_mult_82_CARRYB_35__16_), .A2(
        u5_mult_82_SUMB_35__17_), .ZN(u5_mult_82_n6175) );
  NAND2_X1 u5_mult_82_U5693 ( .A1(u5_mult_82_ab_36__16_), .A2(
        u5_mult_82_SUMB_35__17_), .ZN(u5_mult_82_n6174) );
  XNOR2_X2 u5_mult_82_U5692 ( .A(u5_mult_82_n1786), .B(u5_mult_82_SUMB_20__41_), .ZN(u5_mult_82_SUMB_21__40_) );
  XNOR2_X2 u5_mult_82_U5691 ( .A(u5_mult_82_CARRYB_6__43_), .B(
        u5_mult_82_n1785), .ZN(u5_mult_82_n6095) );
  XNOR2_X2 u5_mult_82_U5690 ( .A(u5_mult_82_n1784), .B(
        u5_mult_82_CARRYB_14__35_), .ZN(u5_mult_82_n5049) );
  XNOR2_X2 u5_mult_82_U5689 ( .A(u5_mult_82_n1783), .B(u5_mult_82_SUMB_14__48_), .ZN(u5_mult_82_SUMB_15__47_) );
  INV_X4 u5_mult_82_U5688 ( .A(u5_mult_82_n1781), .ZN(u5_mult_82_SUMB_44__4_)
         );
  XNOR2_X2 u5_mult_82_U5687 ( .A(u5_mult_82_n5787), .B(u5_mult_82_n417), .ZN(
        u5_mult_82_n1781) );
  XNOR2_X2 u5_mult_82_U5686 ( .A(u5_mult_82_CARRYB_14__34_), .B(
        u5_mult_82_ab_15__34_), .ZN(u5_mult_82_n1780) );
  XNOR2_X2 u5_mult_82_U5685 ( .A(u5_mult_82_n1616), .B(u5_mult_82_n1780), .ZN(
        u5_mult_82_SUMB_15__34_) );
  XNOR2_X2 u5_mult_82_U5684 ( .A(u5_mult_82_CARRYB_27__32_), .B(
        u5_mult_82_ab_28__32_), .ZN(u5_mult_82_n1779) );
  XNOR2_X2 u5_mult_82_U5683 ( .A(u5_mult_82_n1415), .B(u5_mult_82_n1779), .ZN(
        u5_mult_82_SUMB_28__32_) );
  CLKBUF_X2 u5_mult_82_U5682 ( .A(u5_mult_82_SUMB_2__41_), .Z(u5_mult_82_n1778) );
  NAND2_X2 u5_mult_82_U5681 ( .A1(u5_mult_82_ab_25__36_), .A2(
        u5_mult_82_SUMB_24__37_), .ZN(u5_mult_82_n5556) );
  XNOR2_X2 u5_mult_82_U5680 ( .A(u5_mult_82_ab_16__29_), .B(
        u5_mult_82_CARRYB_15__29_), .ZN(u5_mult_82_n1777) );
  XNOR2_X2 u5_mult_82_U5679 ( .A(u5_mult_82_n1777), .B(u5_mult_82_SUMB_15__30_), .ZN(u5_mult_82_SUMB_16__29_) );
  CLKBUF_X2 u5_mult_82_U5678 ( .A(u5_mult_82_CARRYB_11__45_), .Z(
        u5_mult_82_n1776) );
  XNOR2_X2 u5_mult_82_U5677 ( .A(u5_mult_82_CARRYB_34__33_), .B(
        u5_mult_82_n1775), .ZN(u5_mult_82_SUMB_35__33_) );
  XNOR2_X1 u5_mult_82_U5676 ( .A(u5_mult_82_ab_8__42_), .B(
        u5_mult_82_CARRYB_7__42_), .ZN(u5_mult_82_n1774) );
  XNOR2_X2 u5_mult_82_U5675 ( .A(u5_mult_82_n1774), .B(u5_mult_82_SUMB_7__43_), 
        .ZN(u5_mult_82_SUMB_8__42_) );
  XNOR2_X2 u5_mult_82_U5674 ( .A(u5_mult_82_n1773), .B(u5_mult_82_SUMB_20__31_), .ZN(u5_mult_82_SUMB_21__30_) );
  XNOR2_X2 u5_mult_82_U5673 ( .A(u5_mult_82_CARRYB_13__36_), .B(
        u5_mult_82_n1770), .ZN(u5_mult_82_SUMB_14__36_) );
  XNOR2_X2 u5_mult_82_U5672 ( .A(u5_mult_82_n1768), .B(u5_mult_82_n1752), .ZN(
        u5_mult_82_SUMB_41__7_) );
  XNOR2_X2 u5_mult_82_U5671 ( .A(u5_mult_82_CARRYB_8__38_), .B(
        u5_mult_82_ab_9__38_), .ZN(u5_mult_82_n1767) );
  XNOR2_X2 u5_mult_82_U5670 ( .A(u5_mult_82_n1452), .B(u5_mult_82_n1767), .ZN(
        u5_mult_82_SUMB_9__38_) );
  XNOR2_X2 u5_mult_82_U5669 ( .A(u5_mult_82_CARRYB_13__49_), .B(
        u5_mult_82_n1766), .ZN(u5_mult_82_n4322) );
  XNOR2_X2 u5_mult_82_U5668 ( .A(u5_mult_82_CARRYB_7__47_), .B(
        u5_mult_82_n1764), .ZN(u5_mult_82_n3124) );
  INV_X4 u5_mult_82_U5667 ( .A(u5_mult_82_net86784), .ZN(u5_mult_82_net86785)
         );
  INV_X2 u5_mult_82_U5666 ( .A(u5_mult_82_SUMB_8__37_), .ZN(u5_mult_82_n1762)
         );
  XNOR2_X2 u5_mult_82_U5665 ( .A(u5_mult_82_n1759), .B(u5_mult_82_n39), .ZN(
        u5_mult_82_SUMB_39__7_) );
  XNOR2_X2 u5_mult_82_U5664 ( .A(u5_mult_82_ab_20__31_), .B(
        u5_mult_82_CARRYB_19__31_), .ZN(u5_mult_82_n1758) );
  XNOR2_X2 u5_mult_82_U5663 ( .A(u5_mult_82_CARRYB_27__22_), .B(
        u5_mult_82_ab_28__22_), .ZN(u5_mult_82_n1757) );
  XNOR2_X2 u5_mult_82_U5662 ( .A(u5_mult_82_n1757), .B(u5_mult_82_SUMB_27__23_), .ZN(u5_mult_82_SUMB_28__22_) );
  XNOR2_X2 u5_mult_82_U5661 ( .A(u5_mult_82_SUMB_15__38_), .B(u5_mult_82_n1756), .ZN(u5_mult_82_SUMB_16__37_) );
  INV_X2 u5_mult_82_U5660 ( .A(u5_mult_82_SUMB_40__7_), .ZN(u5_mult_82_n1754)
         );
  XNOR2_X2 u5_mult_82_U5659 ( .A(u5_mult_82_ab_38__31_), .B(
        u5_mult_82_CARRYB_37__31_), .ZN(u5_mult_82_n1753) );
  XNOR2_X2 u5_mult_82_U5658 ( .A(u5_mult_82_n1753), .B(u5_mult_82_n1850), .ZN(
        u5_mult_82_SUMB_38__31_) );
  INV_X4 u5_mult_82_U5657 ( .A(u5_mult_82_n1751), .ZN(u5_mult_82_n1752) );
  INV_X2 u5_mult_82_U5656 ( .A(u5_mult_82_SUMB_40__8_), .ZN(u5_mult_82_n1751)
         );
  INV_X4 u5_mult_82_U5655 ( .A(u5_mult_82_SUMB_50__33_), .ZN(u5_mult_82_n1748)
         );
  XNOR2_X2 u5_mult_82_U5654 ( .A(u5_mult_82_n1746), .B(
        u5_mult_82_CARRYB_28__30_), .ZN(u5_mult_82_n4533) );
  INV_X8 u5_mult_82_U5653 ( .A(u5_mult_82_net64913), .ZN(u5_mult_82_net64911)
         );
  AND2_X2 u5_mult_82_U5652 ( .A1(u5_mult_82_net64911), .A2(u5_mult_82_net86863), .ZN(u5_mult_82_ab_2__35_) );
  XNOR2_X2 u5_mult_82_U5651 ( .A(u5_mult_82_n1745), .B(u5_mult_82_SUMB_27__32_), .ZN(u5_mult_82_SUMB_28__31_) );
  XNOR2_X2 u5_mult_82_U5650 ( .A(u5_mult_82_n1744), .B(u5_mult_82_SUMB_42__7_), 
        .ZN(u5_mult_82_SUMB_43__6_) );
  XNOR2_X2 u5_mult_82_U5649 ( .A(u5_mult_82_CARRYB_15__38_), .B(
        u5_mult_82_ab_16__38_), .ZN(u5_mult_82_n1743) );
  XNOR2_X2 u5_mult_82_U5648 ( .A(u5_mult_82_SUMB_15__39_), .B(u5_mult_82_n1743), .ZN(u5_mult_82_SUMB_16__38_) );
  XNOR2_X2 u5_mult_82_U5647 ( .A(u5_mult_82_ab_46__33_), .B(
        u5_mult_82_CARRYB_45__33_), .ZN(u5_mult_82_n1742) );
  XNOR2_X2 u5_mult_82_U5646 ( .A(u5_mult_82_n1742), .B(u5_mult_82_n1501), .ZN(
        u5_mult_82_SUMB_46__33_) );
  NAND2_X1 u5_mult_82_U5645 ( .A1(u5_mult_82_CARRYB_33__21_), .A2(
        u5_mult_82_SUMB_33__22_), .ZN(u5_mult_82_n5895) );
  XNOR2_X2 u5_mult_82_U5644 ( .A(u5_mult_82_n1741), .B(u5_mult_82_n1860), .ZN(
        u5_mult_82_SUMB_45__28_) );
  NAND2_X1 u5_mult_82_U5643 ( .A1(u5_mult_82_CARRYB_32__17_), .A2(
        u5_mult_82_SUMB_32__18_), .ZN(u5_mult_82_n3302) );
  XNOR2_X2 u5_mult_82_U5642 ( .A(u5_mult_82_CARRYB_19__30_), .B(
        u5_mult_82_ab_20__30_), .ZN(u5_mult_82_n1740) );
  XNOR2_X2 u5_mult_82_U5641 ( .A(u5_mult_82_SUMB_19__31_), .B(u5_mult_82_n1740), .ZN(u5_mult_82_SUMB_20__30_) );
  XNOR2_X2 u5_mult_82_U5640 ( .A(u5_mult_82_ab_45__33_), .B(
        u5_mult_82_CARRYB_44__33_), .ZN(u5_mult_82_n1739) );
  XNOR2_X2 u5_mult_82_U5639 ( .A(u5_mult_82_n1739), .B(u5_mult_82_SUMB_44__34_), .ZN(u5_mult_82_SUMB_45__33_) );
  NAND2_X2 u5_mult_82_U5638 ( .A1(u5_mult_82_n1721), .A2(u5_mult_82_ab_45__3_), 
        .ZN(u5_mult_82_n5791) );
  XNOR2_X2 u5_mult_82_U5637 ( .A(u5_mult_82_ab_50__26_), .B(
        u5_mult_82_CARRYB_49__26_), .ZN(u5_mult_82_n1738) );
  XNOR2_X2 u5_mult_82_U5636 ( .A(u5_mult_82_n1738), .B(u5_mult_82_n694), .ZN(
        u5_mult_82_SUMB_50__26_) );
  XOR2_X2 u5_mult_82_U5635 ( .A(u5_mult_82_n4615), .B(u5_mult_82_CARRYB_43__6_), .Z(u5_mult_82_n1737) );
  XNOR2_X2 u5_mult_82_U5634 ( .A(u5_mult_82_n1737), .B(u5_mult_82_SUMB_43__7_), 
        .ZN(u5_mult_82_SUMB_44__6_) );
  XNOR2_X2 u5_mult_82_U5633 ( .A(u5_mult_82_ab_10__44_), .B(
        u5_mult_82_CARRYB_9__44_), .ZN(u5_mult_82_n1736) );
  XNOR2_X2 u5_mult_82_U5632 ( .A(u5_mult_82_n1736), .B(u5_mult_82_SUMB_9__45_), 
        .ZN(u5_mult_82_SUMB_10__44_) );
  XNOR2_X2 u5_mult_82_U5631 ( .A(u5_mult_82_n1735), .B(u5_mult_82_SUMB_44__35_), .ZN(u5_mult_82_SUMB_45__34_) );
  XNOR2_X2 u5_mult_82_U5630 ( .A(u5_mult_82_n1734), .B(u5_mult_82_n410), .ZN(
        u5_mult_82_SUMB_30__29_) );
  XNOR2_X2 u5_mult_82_U5629 ( .A(u5_mult_82_CARRYB_33__21_), .B(
        u5_mult_82_n1733), .ZN(u5_mult_82_n5891) );
  XNOR2_X2 u5_mult_82_U5628 ( .A(u5_mult_82_ab_38__8_), .B(
        u5_mult_82_CARRYB_37__8_), .ZN(u5_mult_82_n1732) );
  XNOR2_X2 u5_mult_82_U5627 ( .A(u5_mult_82_n1732), .B(u5_mult_82_SUMB_37__9_), 
        .ZN(u5_mult_82_SUMB_38__8_) );
  XNOR2_X2 u5_mult_82_U5626 ( .A(u5_mult_82_SUMB_31__33_), .B(u5_mult_82_n1731), .ZN(u5_mult_82_SUMB_32__32_) );
  INV_X4 u5_mult_82_U5625 ( .A(u5_mult_82_n1729), .ZN(u5_mult_82_n1730) );
  INV_X2 u5_mult_82_U5624 ( .A(u5_mult_82_SUMB_40__28_), .ZN(u5_mult_82_n1729)
         );
  CLKBUF_X2 u5_mult_82_U5623 ( .A(u5_mult_82_SUMB_17__46_), .Z(
        u5_mult_82_n1728) );
  NAND3_X2 u5_mult_82_U5622 ( .A1(u5_mult_82_n4214), .A2(u5_mult_82_n4215), 
        .A3(u5_mult_82_n4216), .ZN(u5_mult_82_CARRYB_39__19_) );
  INV_X4 u5_mult_82_U5621 ( .A(u5_mult_82_n1724), .ZN(u5_mult_82_n1725) );
  XNOR2_X2 u5_mult_82_U5620 ( .A(u5_mult_82_n1723), .B(u5_mult_82_SUMB_21__40_), .ZN(u5_mult_82_SUMB_22__39_) );
  XNOR2_X2 u5_mult_82_U5619 ( .A(u5_mult_82_ab_45__14_), .B(
        u5_mult_82_CARRYB_44__14_), .ZN(u5_mult_82_n1722) );
  INV_X4 u5_mult_82_U5618 ( .A(u5_mult_82_n1720), .ZN(u5_mult_82_n1721) );
  INV_X2 u5_mult_82_U5617 ( .A(u5_mult_82_CARRYB_44__3_), .ZN(u5_mult_82_n1720) );
  XNOR2_X2 u5_mult_82_U5616 ( .A(u5_mult_82_n2879), .B(u5_mult_82_n70), .ZN(
        u5_mult_82_SUMB_24__25_) );
  XNOR2_X2 u5_mult_82_U5615 ( .A(u5_mult_82_net79208), .B(u5_mult_82_net87436), 
        .ZN(u5_mult_82_net86976) );
  BUF_X8 u5_mult_82_U5614 ( .A(u5_mult_82_CARRYB_46__20_), .Z(u5_mult_82_n1719) );
  XNOR2_X2 u5_mult_82_U5613 ( .A(u5_mult_82_ab_34__22_), .B(
        u5_mult_82_CARRYB_33__22_), .ZN(u5_mult_82_n1718) );
  INV_X2 u5_mult_82_U5612 ( .A(u5_mult_82_SUMB_20__15_), .ZN(u5_mult_82_n1716)
         );
  NAND2_X1 u5_mult_82_U5611 ( .A1(u5_mult_82_CARRYB_17__30_), .A2(
        u5_mult_82_SUMB_17__31_), .ZN(u5_mult_82_n6014) );
  CLKBUF_X2 u5_mult_82_U5610 ( .A(u5_mult_82_CARRYB_27__27_), .Z(
        u5_mult_82_n1715) );
  XNOR2_X2 u5_mult_82_U5609 ( .A(u5_mult_82_CARRYB_37__15_), .B(
        u5_mult_82_ab_38__15_), .ZN(u5_mult_82_n1714) );
  XNOR2_X2 u5_mult_82_U5608 ( .A(u5_mult_82_SUMB_37__16_), .B(u5_mult_82_n1714), .ZN(u5_mult_82_SUMB_38__15_) );
  NAND2_X2 u5_mult_82_U5607 ( .A1(u5_mult_82_SUMB_18__46_), .A2(
        u5_mult_82_CARRYB_18__45_), .ZN(u5_mult_82_n3367) );
  XNOR2_X2 u5_mult_82_U5606 ( .A(u5_mult_82_ab_33__26_), .B(
        u5_mult_82_CARRYB_32__26_), .ZN(u5_mult_82_n1713) );
  XNOR2_X2 u5_mult_82_U5605 ( .A(u5_mult_82_n1713), .B(u5_mult_82_SUMB_32__27_), .ZN(u5_mult_82_SUMB_33__26_) );
  XOR2_X2 u5_mult_82_U5604 ( .A(u5_mult_82_n4959), .B(u5_mult_82_n1531), .Z(
        u5_mult_82_SUMB_42__3_) );
  NAND2_X1 u5_mult_82_U5603 ( .A1(u5_mult_82_CARRYB_42__2_), .A2(
        u5_mult_82_SUMB_42__3_), .ZN(u5_mult_82_n5635) );
  INV_X4 u5_mult_82_U5602 ( .A(u5_mult_82_n1710), .ZN(u5_mult_82_n1711) );
  INV_X2 u5_mult_82_U5601 ( .A(u5_mult_82_CARRYB_16__47_), .ZN(
        u5_mult_82_n1710) );
  XNOR2_X2 u5_mult_82_U5600 ( .A(u5_mult_82_n1709), .B(u5_mult_82_n1449), .ZN(
        u5_mult_82_SUMB_10__45_) );
  INV_X4 u5_mult_82_U5599 ( .A(u5_mult_82_n1707), .ZN(u5_mult_82_n1708) );
  INV_X2 u5_mult_82_U5598 ( .A(u5_mult_82_SUMB_22__41_), .ZN(u5_mult_82_n1707)
         );
  NAND2_X1 u5_mult_82_U5597 ( .A1(u5_mult_82_CARRYB_27__41_), .A2(
        u5_mult_82_SUMB_27__42_), .ZN(u5_mult_82_n2449) );
  XNOR2_X1 u5_mult_82_U5596 ( .A(u5_mult_82_ab_49__15_), .B(
        u5_mult_82_CARRYB_48__15_), .ZN(u5_mult_82_n1706) );
  XNOR2_X2 u5_mult_82_U5595 ( .A(u5_mult_82_n1706), .B(u5_mult_82_n1845), .ZN(
        u5_mult_82_SUMB_49__15_) );
  CLKBUF_X2 u5_mult_82_U5594 ( .A(u5_mult_82_CARRYB_23__33_), .Z(
        u5_mult_82_n1705) );
  XNOR2_X2 u5_mult_82_U5593 ( .A(u5_mult_82_ab_35__36_), .B(
        u5_mult_82_CARRYB_34__36_), .ZN(u5_mult_82_n1704) );
  XNOR2_X2 u5_mult_82_U5592 ( .A(u5_mult_82_n1704), .B(u5_mult_82_SUMB_34__37_), .ZN(u5_mult_82_SUMB_35__36_) );
  NAND2_X1 u5_mult_82_U5591 ( .A1(u5_mult_82_ab_21__46_), .A2(
        u5_mult_82_SUMB_20__47_), .ZN(u5_mult_82_n2930) );
  XNOR2_X2 u5_mult_82_U5590 ( .A(u5_mult_82_ab_29__11_), .B(
        u5_mult_82_CARRYB_28__11_), .ZN(u5_mult_82_n1703) );
  XNOR2_X2 u5_mult_82_U5589 ( .A(u5_mult_82_n1703), .B(u5_mult_82_SUMB_28__12_), .ZN(u5_mult_82_SUMB_29__11_) );
  NAND3_X2 u5_mult_82_U5588 ( .A1(u5_mult_82_n4796), .A2(u5_mult_82_n4797), 
        .A3(u5_mult_82_n4798), .ZN(u5_mult_82_CARRYB_9__46_) );
  INV_X4 u5_mult_82_U5587 ( .A(u5_mult_82_n1701), .ZN(u5_mult_82_n1702) );
  INV_X2 u5_mult_82_U5586 ( .A(u5_mult_82_SUMB_28__38_), .ZN(u5_mult_82_n1701)
         );
  BUF_X2 u5_mult_82_U5585 ( .A(u5_mult_82_CARRYB_44__29_), .Z(u5_mult_82_n1700) );
  NAND3_X2 u5_mult_82_U5584 ( .A1(u5_mult_82_n5853), .A2(u5_mult_82_n5855), 
        .A3(u5_mult_82_n5854), .ZN(u5_mult_82_CARRYB_48__15_) );
  XNOR2_X2 u5_mult_82_U5583 ( .A(u5_mult_82_n1602), .B(u5_mult_82_n1699), .ZN(
        u5_mult_82_n3259) );
  XOR2_X2 u5_mult_82_U5582 ( .A(u5_mult_82_CARRYB_40__18_), .B(
        u5_mult_82_n4518), .Z(u5_mult_82_n1698) );
  XNOR2_X2 u5_mult_82_U5581 ( .A(u5_mult_82_n1698), .B(u5_mult_82_SUMB_40__19_), .ZN(u5_mult_82_SUMB_41__18_) );
  XNOR2_X2 u5_mult_82_U5580 ( .A(u5_mult_82_ab_36__18_), .B(
        u5_mult_82_CARRYB_35__18_), .ZN(u5_mult_82_n1697) );
  XNOR2_X2 u5_mult_82_U5579 ( .A(u5_mult_82_n1697), .B(u5_mult_82_SUMB_35__19_), .ZN(u5_mult_82_SUMB_36__18_) );
  XNOR2_X2 u5_mult_82_U5578 ( .A(u5_mult_82_CARRYB_46__10_), .B(
        u5_mult_82_n1696), .ZN(u5_mult_82_SUMB_47__10_) );
  XNOR2_X2 u5_mult_82_U5577 ( .A(u5_mult_82_n1460), .B(u5_mult_82_n1695), .ZN(
        u5_mult_82_SUMB_11__40_) );
  BUF_X8 u5_mult_82_U5576 ( .A(u5_mult_82_SUMB_25__10_), .Z(u5_mult_82_n1694)
         );
  INV_X4 u5_mult_82_U5575 ( .A(u5_mult_82_n1692), .ZN(u5_mult_82_n1693) );
  INV_X2 u5_mult_82_U5574 ( .A(u5_mult_82_SUMB_46__15_), .ZN(u5_mult_82_n1692)
         );
  INV_X4 u5_mult_82_U5573 ( .A(u5_mult_82_n1690), .ZN(u5_mult_82_n1691) );
  INV_X2 u5_mult_82_U5572 ( .A(u5_mult_82_SUMB_23__42_), .ZN(u5_mult_82_n1690)
         );
  XNOR2_X2 u5_mult_82_U5571 ( .A(u5_mult_82_ab_49__14_), .B(
        u5_mult_82_CARRYB_48__14_), .ZN(u5_mult_82_n1689) );
  XNOR2_X2 u5_mult_82_U5570 ( .A(u5_mult_82_n1689), .B(u5_mult_82_n1661), .ZN(
        u5_mult_82_SUMB_49__14_) );
  INV_X4 u5_mult_82_U5569 ( .A(u5_mult_82_SUMB_32__10_), .ZN(u5_mult_82_n1687)
         );
  XNOR2_X2 u5_mult_82_U5568 ( .A(u5_mult_82_CARRYB_19__34_), .B(
        u5_mult_82_ab_20__34_), .ZN(u5_mult_82_n1686) );
  XNOR2_X2 u5_mult_82_U5567 ( .A(u5_mult_82_n1686), .B(u5_mult_82_SUMB_19__35_), .ZN(u5_mult_82_SUMB_20__34_) );
  XNOR2_X2 u5_mult_82_U5566 ( .A(u5_mult_82_ab_30__37_), .B(
        u5_mult_82_CARRYB_29__37_), .ZN(u5_mult_82_n1685) );
  XNOR2_X2 u5_mult_82_U5565 ( .A(u5_mult_82_n1685), .B(u5_mult_82_SUMB_29__38_), .ZN(u5_mult_82_SUMB_30__37_) );
  XNOR2_X2 u5_mult_82_U5564 ( .A(u5_mult_82_ab_29__37_), .B(
        u5_mult_82_CARRYB_28__37_), .ZN(u5_mult_82_n1684) );
  XNOR2_X2 u5_mult_82_U5563 ( .A(u5_mult_82_n1684), .B(u5_mult_82_n1702), .ZN(
        u5_mult_82_SUMB_29__37_) );
  CLKBUF_X3 u5_mult_82_U5562 ( .A(u5_mult_82_SUMB_31__9_), .Z(u5_mult_82_n1683) );
  XNOR2_X2 u5_mult_82_U5561 ( .A(u5_mult_82_CARRYB_43__14_), .B(
        u5_mult_82_ab_44__14_), .ZN(u5_mult_82_n1682) );
  XNOR2_X2 u5_mult_82_U5560 ( .A(u5_mult_82_SUMB_43__15_), .B(u5_mult_82_n1682), .ZN(u5_mult_82_SUMB_44__14_) );
  CLKBUF_X2 u5_mult_82_U5559 ( .A(u5_mult_82_SUMB_8__47_), .Z(u5_mult_82_n1681) );
  NAND2_X1 u5_mult_82_U5558 ( .A1(u5_mult_82_CARRYB_2__39_), .A2(
        u5_mult_82_SUMB_2__40_), .ZN(u5_mult_82_n4175) );
  NAND3_X2 u5_mult_82_U5557 ( .A1(u5_mult_82_n2784), .A2(u5_mult_82_n2785), 
        .A3(u5_mult_82_n2786), .ZN(u5_mult_82_CARRYB_27__15_) );
  INV_X8 u5_mult_82_U5556 ( .A(u5_mult_82_n1679), .ZN(u5_mult_82_n1680) );
  INV_X2 u5_mult_82_U5555 ( .A(u5_mult_82_SUMB_17__30_), .ZN(u5_mult_82_n1679)
         );
  NAND2_X2 u5_mult_82_U5554 ( .A1(u5_mult_82_ab_15__31_), .A2(u5_mult_82_n1761), .ZN(u5_mult_82_n5796) );
  XNOR2_X1 u5_mult_82_U5553 ( .A(u5_mult_82_ab_10__35_), .B(
        u5_mult_82_CARRYB_9__35_), .ZN(u5_mult_82_n1678) );
  XNOR2_X2 u5_mult_82_U5552 ( .A(u5_mult_82_SUMB_23__43_), .B(u5_mult_82_n1677), .ZN(u5_mult_82_SUMB_24__42_) );
  XNOR2_X2 u5_mult_82_U5551 ( .A(u5_mult_82_CARRYB_49__22_), .B(
        u5_mult_82_ab_50__22_), .ZN(u5_mult_82_n1676) );
  XNOR2_X2 u5_mult_82_U5550 ( .A(u5_mult_82_SUMB_49__23_), .B(u5_mult_82_n1676), .ZN(u5_mult_82_SUMB_50__22_) );
  XNOR2_X2 u5_mult_82_U5549 ( .A(u5_mult_82_n1629), .B(u5_mult_82_n5157), .ZN(
        u5_mult_82_n1675) );
  XNOR2_X2 u5_mult_82_U5548 ( .A(u5_mult_82_ab_18__30_), .B(
        u5_mult_82_CARRYB_17__30_), .ZN(u5_mult_82_n1674) );
  XNOR2_X2 u5_mult_82_U5547 ( .A(u5_mult_82_n1674), .B(u5_mult_82_SUMB_17__31_), .ZN(u5_mult_82_SUMB_18__30_) );
  CLKBUF_X3 u5_mult_82_U5546 ( .A(u5_mult_82_SUMB_14__31_), .Z(
        u5_mult_82_n1673) );
  CLKBUF_X2 u5_mult_82_U5545 ( .A(u5_mult_82_SUMB_25__36_), .Z(
        u5_mult_82_n1672) );
  XNOR2_X2 u5_mult_82_U5544 ( .A(u5_mult_82_ab_31__39_), .B(
        u5_mult_82_SUMB_30__40_), .ZN(u5_mult_82_n1671) );
  XNOR2_X2 u5_mult_82_U5543 ( .A(u5_mult_82_n1671), .B(
        u5_mult_82_CARRYB_30__39_), .ZN(u5_mult_82_SUMB_31__39_) );
  CLKBUF_X2 u5_mult_82_U5542 ( .A(u5_mult_82_SUMB_31__40_), .Z(
        u5_mult_82_n1670) );
  FA_X1 u5_mult_82_U5541 ( .A(u5_mult_82_ab_49__22_), .B(
        u5_mult_82_CARRYB_48__22_), .CI(u5_mult_82_SUMB_48__23_), .S(
        u5_mult_82_n1669) );
  XNOR2_X2 u5_mult_82_U5540 ( .A(u5_mult_82_SUMB_23__46_), .B(
        u5_mult_82_ab_24__45_), .ZN(u5_mult_82_n1668) );
  XNOR2_X2 u5_mult_82_U5539 ( .A(u5_mult_82_CARRYB_23__45_), .B(
        u5_mult_82_n1668), .ZN(u5_mult_82_SUMB_24__45_) );
  XNOR2_X2 u5_mult_82_U5538 ( .A(u5_mult_82_CARRYB_39__31_), .B(
        u5_mult_82_ab_40__31_), .ZN(u5_mult_82_n1666) );
  XNOR2_X2 u5_mult_82_U5537 ( .A(u5_mult_82_SUMB_39__32_), .B(u5_mult_82_n1666), .ZN(u5_mult_82_SUMB_40__31_) );
  INV_X2 u5_mult_82_U5536 ( .A(u5_mult_82_n1664), .ZN(u5_mult_82_n1665) );
  INV_X4 u5_mult_82_U5535 ( .A(u5_mult_82_n1662), .ZN(u5_mult_82_n1663) );
  INV_X2 u5_mult_82_U5534 ( .A(u5_mult_82_SUMB_48__26_), .ZN(u5_mult_82_n1662)
         );
  XOR2_X2 u5_mult_82_U5533 ( .A(u5_mult_82_n5852), .B(
        u5_mult_82_CARRYB_47__15_), .Z(u5_mult_82_n1661) );
  NAND2_X2 u5_mult_82_U5532 ( .A1(u5_mult_82_ab_39__11_), .A2(
        u5_mult_82_CARRYB_38__11_), .ZN(u5_mult_82_n5131) );
  INV_X4 u5_mult_82_U5531 ( .A(u5_mult_82_n1659), .ZN(u5_mult_82_n1660) );
  INV_X2 u5_mult_82_U5530 ( .A(u5_mult_82_SUMB_10__16_), .ZN(u5_mult_82_n1659)
         );
  XNOR2_X2 u5_mult_82_U5529 ( .A(u5_mult_82_CARRYB_13__48_), .B(
        u5_mult_82_n1658), .ZN(u5_mult_82_SUMB_14__48_) );
  INV_X4 u5_mult_82_U5528 ( .A(u5_mult_82_n1656), .ZN(u5_mult_82_n1657) );
  INV_X2 u5_mult_82_U5527 ( .A(u5_mult_82_CARRYB_27__14_), .ZN(
        u5_mult_82_n1656) );
  FA_X1 u5_mult_82_U5526 ( .A(u5_mult_82_ab_47__13_), .B(
        u5_mult_82_CARRYB_46__13_), .CI(u5_mult_82_n1537), .S(u5_mult_82_n1655) );
  XNOR2_X2 u5_mult_82_U5525 ( .A(u5_mult_82_n1819), .B(u5_mult_82_SUMB_40__16_), .ZN(u5_mult_82_SUMB_41__15_) );
  XNOR2_X2 u5_mult_82_U5524 ( .A(u5_mult_82_ab_40__15_), .B(
        u5_mult_82_CARRYB_39__15_), .ZN(u5_mult_82_n1654) );
  XNOR2_X2 u5_mult_82_U5523 ( .A(u5_mult_82_n1654), .B(u5_mult_82_SUMB_39__16_), .ZN(u5_mult_82_SUMB_40__15_) );
  FA_X1 u5_mult_82_U5522 ( .A(u5_mult_82_ab_42__1_), .B(u5_mult_82_n1587), 
        .CI(u5_mult_82_n1484), .CO(u5_mult_82_n1653) );
  FA_X1 u5_mult_82_U5521 ( .A(u5_mult_82_ab_42__1_), .B(u5_mult_82_n1481), 
        .CI(u5_mult_82_n49), .CO(u5_mult_82_n1652) );
  INV_X2 u5_mult_82_U5520 ( .A(u5_mult_82_SUMB_15__17_), .ZN(u5_mult_82_n1650)
         );
  CLKBUF_X2 u5_mult_82_U5519 ( .A(u5_mult_82_SUMB_45__13_), .Z(
        u5_mult_82_n1649) );
  NAND2_X2 u5_mult_82_U5518 ( .A1(u5_mult_82_ab_25__44_), .A2(u5_mult_82_n1568), .ZN(u5_mult_82_n5589) );
  XNOR2_X2 u5_mult_82_U5517 ( .A(u5_mult_82_SUMB_39__30_), .B(u5_mult_82_n1648), .ZN(u5_mult_82_SUMB_40__29_) );
  INV_X4 u5_mult_82_U5516 ( .A(u5_mult_82_n1646), .ZN(u5_mult_82_n1647) );
  INV_X2 u5_mult_82_U5515 ( .A(u5_mult_82_SUMB_34__27_), .ZN(u5_mult_82_n1646)
         );
  NAND3_X2 u5_mult_82_U5514 ( .A1(u5_mult_82_n3860), .A2(u5_mult_82_n3861), 
        .A3(u5_mult_82_n3862), .ZN(u5_mult_82_CARRYB_41__23_) );
  NAND2_X1 u5_mult_82_U5513 ( .A1(u5_mult_82_ab_26__34_), .A2(
        u5_mult_82_SUMB_25__35_), .ZN(u5_mult_82_n4440) );
  XNOR2_X2 u5_mult_82_U5512 ( .A(u5_mult_82_n1645), .B(
        u5_mult_82_CARRYB_46__2_), .ZN(u5_mult_82_n4511) );
  XNOR2_X2 u5_mult_82_U5511 ( .A(u5_mult_82_ab_29__15_), .B(
        u5_mult_82_CARRYB_28__15_), .ZN(u5_mult_82_n1644) );
  XNOR2_X2 u5_mult_82_U5510 ( .A(u5_mult_82_n1643), .B(u5_mult_82_n1546), .ZN(
        u5_mult_82_SUMB_45__10_) );
  INV_X8 u5_mult_82_U5509 ( .A(u5_mult_82_n1641), .ZN(u5_mult_82_n1642) );
  INV_X2 u5_mult_82_U5508 ( .A(u5_mult_82_SUMB_16__21_), .ZN(u5_mult_82_n1641)
         );
  XNOR2_X2 u5_mult_82_U5507 ( .A(u5_mult_82_n4747), .B(u5_mult_82_n1868), .ZN(
        u5_mult_82_SUMB_10__36_) );
  XNOR2_X2 u5_mult_82_U5506 ( .A(u5_mult_82_ab_20__27_), .B(
        u5_mult_82_CARRYB_19__27_), .ZN(u5_mult_82_n1640) );
  XNOR2_X2 u5_mult_82_U5505 ( .A(u5_mult_82_n1640), .B(u5_mult_82_SUMB_19__28_), .ZN(u5_mult_82_SUMB_20__27_) );
  INV_X4 u5_mult_82_U5504 ( .A(u5_mult_82_n1638), .ZN(u5_mult_82_n1639) );
  INV_X2 u5_mult_82_U5503 ( .A(u5_mult_82_SUMB_14__46_), .ZN(u5_mult_82_n1638)
         );
  CLKBUF_X2 u5_mult_82_U5502 ( .A(u5_mult_82_SUMB_39__4_), .Z(u5_mult_82_n1637) );
  INV_X4 u5_mult_82_U5501 ( .A(u5_mult_82_n1636), .ZN(u5_mult_82_SUMB_47__19_)
         );
  XNOR2_X2 u5_mult_82_U5500 ( .A(u5_mult_82_n1608), .B(u5_mult_82_n5708), .ZN(
        u5_mult_82_n1636) );
  INV_X4 u5_mult_82_U5499 ( .A(u5_mult_82_n1634), .ZN(u5_mult_82_n1635) );
  INV_X2 u5_mult_82_U5498 ( .A(u5_mult_82_SUMB_11__46_), .ZN(u5_mult_82_n1634)
         );
  XNOR2_X1 u5_mult_82_U5497 ( .A(u5_mult_82_SUMB_3__37_), .B(u5_mult_82_n2594), 
        .ZN(u5_mult_82_SUMB_4__36_) );
  XNOR2_X2 u5_mult_82_U5496 ( .A(u5_mult_82_CARRYB_23__47_), .B(
        u5_mult_82_n1633), .ZN(u5_mult_82_n2382) );
  BUF_X4 u5_mult_82_U5495 ( .A(u5_mult_82_SUMB_38__26_), .Z(u5_mult_82_n1632)
         );
  CLKBUF_X2 u5_mult_82_U5494 ( .A(u5_mult_82_CARRYB_34__35_), .Z(
        u5_mult_82_n1631) );
  XNOR2_X2 u5_mult_82_U5493 ( .A(u5_mult_82_ab_39__31_), .B(
        u5_mult_82_CARRYB_38__31_), .ZN(u5_mult_82_n1630) );
  XNOR2_X2 u5_mult_82_U5492 ( .A(u5_mult_82_n1630), .B(u5_mult_82_SUMB_38__32_), .ZN(u5_mult_82_SUMB_39__31_) );
  BUF_X2 u5_mult_82_U5491 ( .A(u5_mult_82_SUMB_40__4_), .Z(u5_mult_82_n1629)
         );
  INV_X4 u5_mult_82_U5490 ( .A(u5_mult_82_n1627), .ZN(u5_mult_82_n1628) );
  CLKBUF_X2 u5_mult_82_U5489 ( .A(u5_mult_82_CARRYB_37__22_), .Z(
        u5_mult_82_n1623) );
  NAND2_X1 u5_mult_82_U5488 ( .A1(u5_mult_82_ab_38__24_), .A2(
        u5_mult_82_SUMB_37__25_), .ZN(u5_mult_82_n3634) );
  CLKBUF_X2 u5_mult_82_U5487 ( .A(u5_mult_82_SUMB_26__24_), .Z(
        u5_mult_82_n1622) );
  XNOR2_X2 u5_mult_82_U5486 ( .A(u5_mult_82_ab_35__30_), .B(
        u5_mult_82_CARRYB_34__30_), .ZN(u5_mult_82_n1621) );
  XNOR2_X2 u5_mult_82_U5485 ( .A(u5_mult_82_n1621), .B(u5_mult_82_SUMB_34__31_), .ZN(u5_mult_82_SUMB_35__30_) );
  INV_X1 u5_mult_82_U5484 ( .A(u5_mult_82_SUMB_45__4_), .ZN(u5_mult_82_n1624)
         );
  XNOR2_X2 u5_mult_82_U5483 ( .A(u5_mult_82_n4510), .B(u5_mult_82_n1624), .ZN(
        u5_mult_82_SUMB_46__3_) );
  XNOR2_X2 u5_mult_82_U5482 ( .A(u5_mult_82_SUMB_43__6_), .B(u5_mult_82_n1620), 
        .ZN(u5_mult_82_SUMB_44__5_) );
  XNOR2_X2 u5_mult_82_U5481 ( .A(u5_mult_82_ab_7__25_), .B(
        u5_mult_82_CARRYB_6__25_), .ZN(u5_mult_82_n1619) );
  XNOR2_X2 u5_mult_82_U5480 ( .A(u5_mult_82_n1619), .B(u5_mult_82_SUMB_6__26_), 
        .ZN(u5_mult_82_SUMB_7__25_) );
  XNOR2_X2 u5_mult_82_U5479 ( .A(u5_mult_82_ab_15__47_), .B(
        u5_mult_82_CARRYB_14__47_), .ZN(u5_mult_82_n1783) );
  NAND2_X2 u5_mult_82_U5478 ( .A1(u5_mult_82_ab_15__47_), .A2(
        u5_mult_82_CARRYB_14__47_), .ZN(u5_mult_82_n4609) );
  XNOR2_X2 u5_mult_82_U5477 ( .A(u5_mult_82_CARRYB_20__20_), .B(
        u5_mult_82_ab_21__20_), .ZN(u5_mult_82_n4163) );
  XNOR2_X2 u5_mult_82_U5476 ( .A(u5_mult_82_CARRYB_40__31_), .B(
        u5_mult_82_ab_41__31_), .ZN(u5_mult_82_n1618) );
  XNOR2_X2 u5_mult_82_U5475 ( .A(u5_mult_82_n1617), .B(u5_mult_82_SUMB_40__3_), 
        .ZN(u5_mult_82_SUMB_41__2_) );
  INV_X2 u5_mult_82_U5474 ( .A(u5_mult_82_SUMB_14__35_), .ZN(u5_mult_82_n1615)
         );
  XNOR2_X2 u5_mult_82_U5473 ( .A(u5_mult_82_SUMB_52__2_), .B(
        u5_mult_82_CARRYB_52__1_), .ZN(u5_mult_82_n6390) );
  INV_X8 u5_mult_82_U5472 ( .A(u5_mult_82_n1613), .ZN(u5_mult_82_n1614) );
  INV_X4 u5_mult_82_U5471 ( .A(u5_mult_82_CARRYB_27__33_), .ZN(
        u5_mult_82_n1613) );
  XNOR2_X2 u5_mult_82_U5470 ( .A(u5_mult_82_n394), .B(u5_mult_82_ab_28__13_), 
        .ZN(u5_mult_82_n1612) );
  XNOR2_X2 u5_mult_82_U5469 ( .A(u5_mult_82_n1612), .B(u5_mult_82_n1848), .ZN(
        u5_mult_82_SUMB_28__13_) );
  INV_X8 u5_mult_82_U5468 ( .A(u5_mult_82_n609), .ZN(u5_mult_82_n1827) );
  NAND2_X4 u5_mult_82_U5467 ( .A1(u5_mult_82_ab_16__36_), .A2(u5_mult_82_n1827), .ZN(u5_mult_82_n6188) );
  NAND2_X2 u5_mult_82_U5466 ( .A1(u5_mult_82_SUMB_50__20_), .A2(
        u5_mult_82_n2715), .ZN(u5_mult_82_n4913) );
  NAND2_X2 u5_mult_82_U5465 ( .A1(u5_mult_82_ab_51__19_), .A2(
        u5_mult_82_SUMB_50__20_), .ZN(u5_mult_82_n4912) );
  INV_X2 u5_mult_82_U5464 ( .A(u5_mult_82_SUMB_44__7_), .ZN(u5_mult_82_n1609)
         );
  INV_X4 u5_mult_82_U5463 ( .A(u5_mult_82_n1607), .ZN(u5_mult_82_n1608) );
  INV_X2 u5_mult_82_U5462 ( .A(u5_mult_82_SUMB_46__20_), .ZN(u5_mult_82_n1607)
         );
  INV_X4 u5_mult_82_U5461 ( .A(u5_mult_82_n1605), .ZN(u5_mult_82_n1606) );
  INV_X2 u5_mult_82_U5460 ( .A(u5_mult_82_CARRYB_12__20_), .ZN(
        u5_mult_82_n1605) );
  AND2_X4 u5_mult_82_U5459 ( .A1(u5_mult_82_SUMB_52__2_), .A2(
        u5_mult_82_CARRYB_52__1_), .ZN(u5_mult_82_n1604) );
  INV_X4 u5_mult_82_U5458 ( .A(u5_mult_82_n1601), .ZN(u5_mult_82_n1602) );
  INV_X2 u5_mult_82_U5457 ( .A(u5_mult_82_CARRYB_47__30_), .ZN(
        u5_mult_82_n1601) );
  CLKBUF_X2 u5_mult_82_U5456 ( .A(u5_mult_82_SUMB_33__6_), .Z(u5_mult_82_n1600) );
  NAND3_X2 u5_mult_82_U5455 ( .A1(u5_mult_82_n2245), .A2(u5_mult_82_n2244), 
        .A3(u5_mult_82_n2243), .ZN(u5_mult_82_CARRYB_40__23_) );
  XNOR2_X2 u5_mult_82_U5454 ( .A(u5_mult_82_CARRYB_46__31_), .B(
        u5_mult_82_ab_47__31_), .ZN(u5_mult_82_n1599) );
  XNOR2_X2 u5_mult_82_U5453 ( .A(u5_mult_82_SUMB_46__32_), .B(u5_mult_82_n1599), .ZN(u5_mult_82_SUMB_47__31_) );
  CLKBUF_X2 u5_mult_82_U5452 ( .A(u5_mult_82_SUMB_23__47_), .Z(
        u5_mult_82_n1598) );
  INV_X4 u5_mult_82_U5451 ( .A(u5_mult_82_net87429), .ZN(u5_mult_82_net87430)
         );
  CLKBUF_X2 u5_mult_82_U5450 ( .A(u5_mult_82_SUMB_16__18_), .Z(
        u5_mult_82_n1597) );
  NAND3_X2 u5_mult_82_U5449 ( .A1(u5_mult_82_n2181), .A2(u5_mult_82_n2182), 
        .A3(u5_mult_82_n2183), .ZN(u5_mult_82_CARRYB_29__41_) );
  XNOR2_X2 u5_mult_82_U5448 ( .A(u5_mult_82_ab_21__25_), .B(
        u5_mult_82_CARRYB_20__25_), .ZN(u5_mult_82_net87435) );
  CLKBUF_X2 u5_mult_82_U5447 ( .A(u5_mult_82_SUMB_28__21_), .Z(
        u5_mult_82_net87436) );
  NAND2_X1 u5_mult_82_U5446 ( .A1(u5_mult_82_ab_10__29_), .A2(
        u5_mult_82_SUMB_9__30_), .ZN(u5_mult_82_n3328) );
  INV_X4 u5_mult_82_U5445 ( .A(u5_mult_82_n1593), .ZN(u5_mult_82_n1594) );
  INV_X2 u5_mult_82_U5444 ( .A(u5_mult_82_SUMB_44__30_), .ZN(u5_mult_82_n1593)
         );
  INV_X4 u5_mult_82_U5443 ( .A(u5_mult_82_n1591), .ZN(u5_mult_82_n1592) );
  INV_X2 u5_mult_82_U5442 ( .A(u5_mult_82_SUMB_6__40_), .ZN(u5_mult_82_n1591)
         );
  XNOR2_X2 u5_mult_82_U5441 ( .A(u5_mult_82_n1590), .B(
        u5_mult_82_CARRYB_2__40_), .ZN(u5_mult_82_n5499) );
  XNOR2_X1 u5_mult_82_U5440 ( .A(u5_mult_82_ab_45__29_), .B(
        u5_mult_82_CARRYB_44__29_), .ZN(u5_mult_82_n1589) );
  XNOR2_X2 u5_mult_82_U5439 ( .A(u5_mult_82_n1589), .B(u5_mult_82_n1594), .ZN(
        u5_mult_82_SUMB_45__29_) );
  XNOR2_X2 u5_mult_82_U5438 ( .A(u5_mult_82_CARRYB_43__19_), .B(
        u5_mult_82_ab_44__19_), .ZN(u5_mult_82_n1588) );
  XNOR2_X2 u5_mult_82_U5437 ( .A(u5_mult_82_SUMB_43__20_), .B(u5_mult_82_n1588), .ZN(u5_mult_82_SUMB_44__19_) );
  XNOR2_X2 u5_mult_82_U5436 ( .A(u5_mult_82_n4639), .B(u5_mult_82_SUMB_30__18_), .ZN(u5_mult_82_SUMB_31__17_) );
  XNOR2_X2 u5_mult_82_U5435 ( .A(u5_mult_82_ab_6__39_), .B(
        u5_mult_82_CARRYB_5__39_), .ZN(u5_mult_82_n1586) );
  XNOR2_X2 u5_mult_82_U5434 ( .A(u5_mult_82_n1586), .B(u5_mult_82_SUMB_5__40_), 
        .ZN(u5_mult_82_SUMB_6__39_) );
  XNOR2_X2 u5_mult_82_U5433 ( .A(u5_mult_82_n1585), .B(
        u5_mult_82_CARRYB_41__21_), .ZN(u5_mult_82_n2247) );
  INV_X2 u5_mult_82_U5432 ( .A(u5_mult_82_n1583), .ZN(u5_mult_82_n1584) );
  INV_X1 u5_mult_82_U5431 ( .A(u5_mult_82_SUMB_24__47_), .ZN(u5_mult_82_n1583)
         );
  INV_X4 u5_mult_82_U5430 ( .A(u5_mult_82_n1580), .ZN(u5_mult_82_n1581) );
  INV_X2 u5_mult_82_U5429 ( .A(u5_mult_82_SUMB_47__35_), .ZN(u5_mult_82_n1580)
         );
  XNOR2_X2 u5_mult_82_U5428 ( .A(u5_mult_82_ab_48__19_), .B(
        u5_mult_82_CARRYB_47__19_), .ZN(u5_mult_82_n1579) );
  XNOR2_X2 u5_mult_82_U5427 ( .A(u5_mult_82_ab_23__26_), .B(
        u5_mult_82_CARRYB_22__26_), .ZN(u5_mult_82_n1578) );
  XNOR2_X2 u5_mult_82_U5426 ( .A(u5_mult_82_n1578), .B(u5_mult_82_SUMB_22__27_), .ZN(u5_mult_82_SUMB_23__26_) );
  INV_X1 u5_mult_82_U5425 ( .A(u5_mult_82_SUMB_44__33_), .ZN(u5_mult_82_n1576)
         );
  INV_X2 u5_mult_82_U5424 ( .A(u5_mult_82_SUMB_34__33_), .ZN(u5_mult_82_n1574)
         );
  NAND2_X2 u5_mult_82_U5423 ( .A1(u5_mult_82_ab_33__10_), .A2(u5_mult_82_n1514), .ZN(u5_mult_82_n4151) );
  XNOR2_X1 u5_mult_82_U5422 ( .A(u5_mult_82_ab_32__11_), .B(
        u5_mult_82_CARRYB_31__11_), .ZN(u5_mult_82_n1573) );
  XNOR2_X2 u5_mult_82_U5421 ( .A(u5_mult_82_n1573), .B(u5_mult_82_SUMB_31__12_), .ZN(u5_mult_82_SUMB_32__11_) );
  NAND2_X2 u5_mult_82_U5420 ( .A1(u5_mult_82_n42), .A2(u5_mult_82_SUMB_44__35_), .ZN(u5_mult_82_n2610) );
  INV_X4 u5_mult_82_U5419 ( .A(u5_mult_82_n1571), .ZN(u5_mult_82_n1572) );
  INV_X2 u5_mult_82_U5418 ( .A(u5_mult_82_SUMB_11__26_), .ZN(u5_mult_82_n1571)
         );
  INV_X4 u5_mult_82_U5417 ( .A(u5_mult_82_n1569), .ZN(u5_mult_82_n1570) );
  INV_X2 u5_mult_82_U5416 ( .A(u5_mult_82_SUMB_45__36_), .ZN(u5_mult_82_n1569)
         );
  XOR2_X1 u5_mult_82_U5415 ( .A(u5_mult_82_CARRYB_33__44_), .B(
        u5_mult_82_ab_34__44_), .Z(u5_mult_82_n2635) );
  NAND2_X1 u5_mult_82_U5414 ( .A1(u5_mult_82_CARRYB_33__44_), .A2(
        u5_mult_82_SUMB_33__45_), .ZN(u5_mult_82_n2639) );
  INV_X4 u5_mult_82_U5413 ( .A(u5_mult_82_n1567), .ZN(u5_mult_82_n1568) );
  INV_X2 u5_mult_82_U5412 ( .A(u5_mult_82_CARRYB_24__44_), .ZN(
        u5_mult_82_n1567) );
  XNOR2_X1 u5_mult_82_U5411 ( .A(u5_mult_82_ab_31__12_), .B(
        u5_mult_82_CARRYB_30__12_), .ZN(u5_mult_82_n1565) );
  XNOR2_X2 u5_mult_82_U5410 ( .A(u5_mult_82_n1565), .B(u5_mult_82_n1839), .ZN(
        u5_mult_82_SUMB_31__12_) );
  CLKBUF_X2 u5_mult_82_U5409 ( .A(u5_mult_82_SUMB_31__26_), .Z(
        u5_mult_82_n1564) );
  INV_X4 u5_mult_82_U5408 ( .A(u5_mult_82_n1562), .ZN(u5_mult_82_n1563) );
  INV_X2 u5_mult_82_U5407 ( .A(u5_mult_82_SUMB_33__43_), .ZN(u5_mult_82_n1562)
         );
  XNOR2_X2 u5_mult_82_U5406 ( .A(u5_mult_82_n1561), .B(u5_mult_82_n4384), .ZN(
        u5_mult_82_SUMB_42__8_) );
  CLKBUF_X3 u5_mult_82_U5405 ( .A(u5_mult_82_SUMB_38__34_), .Z(
        u5_mult_82_n1560) );
  INV_X4 u5_mult_82_U5404 ( .A(u5_mult_82_n1558), .ZN(u5_mult_82_n1559) );
  INV_X2 u5_mult_82_U5403 ( .A(u5_mult_82_SUMB_18__44_), .ZN(u5_mult_82_n1558)
         );
  XNOR2_X2 u5_mult_82_U5402 ( .A(u5_mult_82_ab_13__45_), .B(
        u5_mult_82_CARRYB_12__45_), .ZN(u5_mult_82_n1557) );
  XNOR2_X2 u5_mult_82_U5401 ( .A(u5_mult_82_n1557), .B(u5_mult_82_SUMB_12__46_), .ZN(u5_mult_82_SUMB_13__45_) );
  XNOR2_X2 u5_mult_82_U5400 ( .A(u5_mult_82_CARRYB_5__42_), .B(
        u5_mult_82_ab_6__42_), .ZN(u5_mult_82_n1556) );
  XNOR2_X2 u5_mult_82_U5399 ( .A(u5_mult_82_SUMB_5__43_), .B(u5_mult_82_n1556), 
        .ZN(u5_mult_82_SUMB_6__42_) );
  NAND2_X1 u5_mult_82_U5398 ( .A1(u5_mult_82_CARRYB_22__28_), .A2(
        u5_mult_82_SUMB_22__29_), .ZN(u5_mult_82_n4299) );
  XNOR2_X1 u5_mult_82_U5397 ( .A(u5_mult_82_ab_39__6_), .B(
        u5_mult_82_CARRYB_38__6_), .ZN(u5_mult_82_n1555) );
  XNOR2_X2 u5_mult_82_U5396 ( .A(u5_mult_82_n1555), .B(u5_mult_82_SUMB_38__7_), 
        .ZN(u5_mult_82_SUMB_39__6_) );
  XNOR2_X2 u5_mult_82_U5395 ( .A(u5_mult_82_ab_27__32_), .B(
        u5_mult_82_CARRYB_26__32_), .ZN(u5_mult_82_n1554) );
  XNOR2_X2 u5_mult_82_U5394 ( .A(u5_mult_82_n1554), .B(u5_mult_82_SUMB_26__33_), .ZN(u5_mult_82_SUMB_27__32_) );
  INV_X2 u5_mult_82_U5393 ( .A(u5_mult_82_SUMB_22__33_), .ZN(u5_mult_82_n1552)
         );
  XNOR2_X2 u5_mult_82_U5392 ( .A(u5_mult_82_CARRYB_44__18_), .B(
        u5_mult_82_ab_45__18_), .ZN(u5_mult_82_n1551) );
  XNOR2_X2 u5_mult_82_U5391 ( .A(u5_mult_82_SUMB_44__19_), .B(u5_mult_82_n1551), .ZN(u5_mult_82_SUMB_45__18_) );
  INV_X4 u5_mult_82_U5390 ( .A(u5_mult_82_n1549), .ZN(u5_mult_82_n1550) );
  INV_X2 u5_mult_82_U5389 ( .A(u5_mult_82_SUMB_28__34_), .ZN(u5_mult_82_n1549)
         );
  INV_X8 u5_mult_82_U5388 ( .A(u5_mult_82_n6390), .ZN(u5_mult_82_CLA_SUM[54])
         );
  CLKBUF_X2 u5_mult_82_U5387 ( .A(u5_mult_82_CARRYB_40__7_), .Z(
        u5_mult_82_n1548) );
  FA_X1 u5_mult_82_U5386 ( .A(u5_mult_82_ab_2__48_), .B(
        u5_mult_82_CARRYB_1__48_), .CI(u5_mult_82_SUMB_1__49_), .S(
        u5_mult_82_n1547) );
  NAND2_X1 u5_mult_82_U5385 ( .A1(u5_mult_82_ab_47__16_), .A2(
        u5_mult_82_CARRYB_46__16_), .ZN(u5_mult_82_n5864) );
  BUF_X2 u5_mult_82_U5384 ( .A(u5_mult_82_SUMB_44__11_), .Z(u5_mult_82_n1546)
         );
  XNOR2_X2 u5_mult_82_U5383 ( .A(u5_mult_82_ab_50__12_), .B(
        u5_mult_82_CARRYB_49__12_), .ZN(u5_mult_82_n1545) );
  XNOR2_X2 u5_mult_82_U5382 ( .A(u5_mult_82_n1545), .B(u5_mult_82_SUMB_49__13_), .ZN(u5_mult_82_SUMB_50__12_) );
  XNOR2_X2 u5_mult_82_U5381 ( .A(u5_mult_82_ab_49__23_), .B(
        u5_mult_82_CARRYB_48__23_), .ZN(u5_mult_82_n1544) );
  XNOR2_X2 u5_mult_82_U5380 ( .A(u5_mult_82_n1544), .B(u5_mult_82_SUMB_48__24_), .ZN(u5_mult_82_SUMB_49__23_) );
  XNOR2_X2 u5_mult_82_U5379 ( .A(u5_mult_82_ab_24__34_), .B(
        u5_mult_82_CARRYB_23__34_), .ZN(u5_mult_82_n1543) );
  XNOR2_X2 u5_mult_82_U5378 ( .A(u5_mult_82_n1543), .B(u5_mult_82_SUMB_23__35_), .ZN(u5_mult_82_SUMB_24__34_) );
  XNOR2_X1 u5_mult_82_U5377 ( .A(u5_mult_82_ab_24__33_), .B(
        u5_mult_82_CARRYB_23__33_), .ZN(u5_mult_82_n1542) );
  XNOR2_X2 u5_mult_82_U5376 ( .A(u5_mult_82_n1542), .B(u5_mult_82_n704), .ZN(
        u5_mult_82_SUMB_24__33_) );
  NAND2_X1 u5_mult_82_U5375 ( .A1(u5_mult_82_CARRYB_7__28_), .A2(
        u5_mult_82_SUMB_7__29_), .ZN(u5_mult_82_n2507) );
  XNOR2_X2 u5_mult_82_U5374 ( .A(u5_mult_82_ab_48__9_), .B(
        u5_mult_82_CARRYB_47__9_), .ZN(u5_mult_82_n1540) );
  XNOR2_X2 u5_mult_82_U5373 ( .A(u5_mult_82_n1540), .B(u5_mult_82_SUMB_47__10_), .ZN(u5_mult_82_SUMB_48__9_) );
  CLKBUF_X3 u5_mult_82_U5372 ( .A(u5_mult_82_SUMB_9__50_), .Z(u5_mult_82_n1539) );
  BUF_X2 u5_mult_82_U5371 ( .A(u5_mult_82_SUMB_23__28_), .Z(u5_mult_82_n1538)
         );
  XNOR2_X1 u5_mult_82_U5370 ( .A(u5_mult_82_SUMB_48__18_), .B(
        u5_mult_82_ab_49__17_), .ZN(u5_mult_82_n1536) );
  XNOR2_X2 u5_mult_82_U5369 ( .A(u5_mult_82_CARRYB_48__17_), .B(
        u5_mult_82_n1536), .ZN(u5_mult_82_SUMB_49__17_) );
  XNOR2_X2 u5_mult_82_U5368 ( .A(u5_mult_82_ab_22__25_), .B(
        u5_mult_82_CARRYB_21__25_), .ZN(u5_mult_82_n1535) );
  XNOR2_X2 u5_mult_82_U5367 ( .A(u5_mult_82_n1535), .B(u5_mult_82_SUMB_21__26_), .ZN(u5_mult_82_SUMB_22__25_) );
  INV_X8 u5_mult_82_U5366 ( .A(u5_mult_82_n1533), .ZN(u5_mult_82_n1534) );
  INV_X2 u5_mult_82_U5365 ( .A(u5_mult_82_SUMB_6__31_), .ZN(u5_mult_82_n1533)
         );
  NAND2_X1 u5_mult_82_U5364 ( .A1(u5_mult_82_ab_31__16_), .A2(
        u5_mult_82_SUMB_30__17_), .ZN(u5_mult_82_n4359) );
  NAND2_X1 u5_mult_82_U5363 ( .A1(u5_mult_82_CARRYB_40__4_), .A2(
        u5_mult_82_SUMB_40__5_), .ZN(u5_mult_82_n4962) );
  NAND2_X1 u5_mult_82_U5362 ( .A1(u5_mult_82_CARRYB_38__29_), .A2(
        u5_mult_82_SUMB_38__30_), .ZN(u5_mult_82_n4716) );
  XNOR2_X2 u5_mult_82_U5361 ( .A(u5_mult_82_ab_44__2_), .B(
        u5_mult_82_CARRYB_43__2_), .ZN(u5_mult_82_n1532) );
  XNOR2_X2 u5_mult_82_U5360 ( .A(u5_mult_82_n1532), .B(u5_mult_82_SUMB_43__3_), 
        .ZN(u5_mult_82_SUMB_44__2_) );
  INV_X8 u5_mult_82_U5359 ( .A(u5_mult_82_n1529), .ZN(u5_mult_82_n1530) );
  INV_X2 u5_mult_82_U5358 ( .A(u5_mult_82_SUMB_12__27_), .ZN(u5_mult_82_n1529)
         );
  NAND2_X1 u5_mult_82_U5357 ( .A1(u5_mult_82_CARRYB_17__39_), .A2(
        u5_mult_82_SUMB_17__40_), .ZN(u5_mult_82_n4410) );
  NAND2_X1 u5_mult_82_U5356 ( .A1(u5_mult_82_ab_18__39_), .A2(
        u5_mult_82_SUMB_17__40_), .ZN(u5_mult_82_n4409) );
  NAND3_X2 u5_mult_82_U5355 ( .A1(u5_mult_82_n4714), .A2(u5_mult_82_n4715), 
        .A3(u5_mult_82_n4716), .ZN(u5_mult_82_CARRYB_39__29_) );
  XNOR2_X2 u5_mult_82_U5354 ( .A(u5_mult_82_ab_3__51_), .B(
        u5_mult_82_ab_2__52_), .ZN(u5_mult_82_n1528) );
  INV_X4 u5_mult_82_U5353 ( .A(u5_mult_82_n1526), .ZN(u5_mult_82_n1527) );
  INV_X2 u5_mult_82_U5352 ( .A(u5_mult_82_CARRYB_14__30_), .ZN(
        u5_mult_82_n1526) );
  XNOR2_X2 u5_mult_82_U5351 ( .A(u5_mult_82_n2112), .B(u5_mult_82_ab_50__13_), 
        .ZN(u5_mult_82_n1525) );
  XNOR2_X2 u5_mult_82_U5350 ( .A(u5_mult_82_n1525), .B(u5_mult_82_SUMB_49__14_), .ZN(u5_mult_82_SUMB_50__13_) );
  XNOR2_X2 u5_mult_82_U5349 ( .A(u5_mult_82_ab_38__13_), .B(
        u5_mult_82_CARRYB_37__13_), .ZN(u5_mult_82_n1524) );
  XNOR2_X2 u5_mult_82_U5348 ( .A(u5_mult_82_n1524), .B(u5_mult_82_net87325), 
        .ZN(u5_mult_82_SUMB_38__13_) );
  XNOR2_X2 u5_mult_82_U5347 ( .A(u5_mult_82_ab_47__9_), .B(
        u5_mult_82_CARRYB_46__9_), .ZN(u5_mult_82_n1523) );
  XNOR2_X2 u5_mult_82_U5346 ( .A(u5_mult_82_n1523), .B(u5_mult_82_SUMB_46__10_), .ZN(u5_mult_82_SUMB_47__9_) );
  XNOR2_X2 u5_mult_82_U5345 ( .A(u5_mult_82_ab_48__25_), .B(
        u5_mult_82_CARRYB_47__25_), .ZN(u5_mult_82_n1520) );
  XNOR2_X2 u5_mult_82_U5344 ( .A(u5_mult_82_n1520), .B(u5_mult_82_n727), .ZN(
        u5_mult_82_SUMB_48__25_) );
  XNOR2_X2 u5_mult_82_U5343 ( .A(u5_mult_82_SUMB_32__23_), .B(u5_mult_82_n1519), .ZN(u5_mult_82_SUMB_33__22_) );
  XNOR2_X2 u5_mult_82_U5342 ( .A(u5_mult_82_ab_46__12_), .B(
        u5_mult_82_CARRYB_45__12_), .ZN(u5_mult_82_n1518) );
  XNOR2_X2 u5_mult_82_U5341 ( .A(u5_mult_82_n1518), .B(u5_mult_82_n1649), .ZN(
        u5_mult_82_SUMB_46__12_) );
  XNOR2_X2 u5_mult_82_U5340 ( .A(u5_mult_82_ab_5__49_), .B(
        u5_mult_82_CARRYB_4__49_), .ZN(u5_mult_82_n1517) );
  XNOR2_X2 u5_mult_82_U5339 ( .A(u5_mult_82_n1517), .B(u5_mult_82_n1861), .ZN(
        u5_mult_82_SUMB_5__49_) );
  XNOR2_X2 u5_mult_82_U5338 ( .A(u5_mult_82_n3702), .B(
        u5_mult_82_CARRYB_30__16_), .ZN(u5_mult_82_SUMB_31__16_) );
  XNOR2_X2 u5_mult_82_U5337 ( .A(u5_mult_82_ab_30__26_), .B(
        u5_mult_82_CARRYB_29__26_), .ZN(u5_mult_82_n1516) );
  XNOR2_X2 u5_mult_82_U5336 ( .A(u5_mult_82_n1516), .B(u5_mult_82_SUMB_29__27_), .ZN(u5_mult_82_SUMB_30__26_) );
  INV_X4 u5_mult_82_U5335 ( .A(u5_mult_82_n1513), .ZN(u5_mult_82_n1514) );
  INV_X2 u5_mult_82_U5334 ( .A(u5_mult_82_CARRYB_32__10_), .ZN(
        u5_mult_82_n1513) );
  INV_X4 u5_mult_82_U5333 ( .A(u5_mult_82_n1511), .ZN(u5_mult_82_n1512) );
  INV_X2 u5_mult_82_U5332 ( .A(u5_mult_82_SUMB_17__39_), .ZN(u5_mult_82_n1511)
         );
  NAND2_X2 u5_mult_82_U5331 ( .A1(u5_mult_82_ab_18__29_), .A2(u5_mult_82_n303), 
        .ZN(u5_mult_82_n5426) );
  INV_X4 u5_mult_82_U5330 ( .A(u5_mult_82_n1509), .ZN(u5_mult_82_n1510) );
  INV_X2 u5_mult_82_U5329 ( .A(u5_mult_82_CARRYB_6__41_), .ZN(u5_mult_82_n1509) );
  CLKBUF_X3 u5_mult_82_U5328 ( .A(u5_mult_82_SUMB_33__44_), .Z(
        u5_mult_82_n1508) );
  NAND2_X1 u5_mult_82_U5327 ( .A1(u5_mult_82_CARRYB_5__30_), .A2(
        u5_mult_82_SUMB_5__31_), .ZN(u5_mult_82_n3464) );
  NAND2_X1 u5_mult_82_U5326 ( .A1(u5_mult_82_ab_6__30_), .A2(
        u5_mult_82_SUMB_5__31_), .ZN(u5_mult_82_n3465) );
  XNOR2_X2 u5_mult_82_U5325 ( .A(u5_mult_82_ab_22__37_), .B(
        u5_mult_82_CARRYB_21__37_), .ZN(u5_mult_82_n1507) );
  XNOR2_X2 u5_mult_82_U5324 ( .A(u5_mult_82_n1507), .B(u5_mult_82_SUMB_21__38_), .ZN(u5_mult_82_SUMB_22__37_) );
  XNOR2_X2 u5_mult_82_U5323 ( .A(u5_mult_82_n1506), .B(u5_mult_82_SUMB_32__11_), .ZN(u5_mult_82_SUMB_33__10_) );
  NAND2_X1 u5_mult_82_U5322 ( .A1(u5_mult_82_CARRYB_27__30_), .A2(
        u5_mult_82_SUMB_27__31_), .ZN(u5_mult_82_n3227) );
  FA_X1 u5_mult_82_U5321 ( .A(u5_mult_82_ab_40__1_), .B(u5_mult_82_n208), .CI(
        u5_mult_82_SUMB_39__2_), .CO(u5_mult_82_n1504) );
  XNOR2_X2 u5_mult_82_U5320 ( .A(u5_mult_82_CARRYB_46__36_), .B(
        u5_mult_82_n2802), .ZN(u5_mult_82_n1503) );
  XNOR2_X2 u5_mult_82_U5319 ( .A(u5_mult_82_ab_22__32_), .B(
        u5_mult_82_CARRYB_21__32_), .ZN(u5_mult_82_n1502) );
  XNOR2_X2 u5_mult_82_U5318 ( .A(u5_mult_82_n17), .B(u5_mult_82_n1502), .ZN(
        u5_mult_82_SUMB_22__32_) );
  INV_X4 u5_mult_82_U5317 ( .A(u5_mult_82_n1499), .ZN(u5_mult_82_n1500) );
  INV_X2 u5_mult_82_U5316 ( .A(u5_mult_82_SUMB_31__27_), .ZN(u5_mult_82_n1499)
         );
  INV_X2 u5_mult_82_U5315 ( .A(u5_mult_82_SUMB_27__17_), .ZN(u5_mult_82_n1497)
         );
  NAND2_X2 u5_mult_82_U5314 ( .A1(u5_mult_82_CARRYB_28__10_), .A2(
        u5_mult_82_SUMB_28__11_), .ZN(u5_mult_82_n3737) );
  XOR2_X1 u5_mult_82_U5313 ( .A(u5_mult_82_n5945), .B(u5_mult_82_SUMB_32__32_), 
        .Z(u5_mult_82_n1496) );
  XNOR2_X2 u5_mult_82_U5312 ( .A(u5_mult_82_CARRYB_40__4_), .B(
        u5_mult_82_ab_41__4_), .ZN(u5_mult_82_n4640) );
  NAND3_X2 u5_mult_82_U5311 ( .A1(u5_mult_82_n5526), .A2(u5_mult_82_n5527), 
        .A3(u5_mult_82_n5528), .ZN(u5_mult_82_CARRYB_39__15_) );
  XNOR2_X2 u5_mult_82_U5310 ( .A(u5_mult_82_n1494), .B(u5_mult_82_SUMB_41__16_), .ZN(u5_mult_82_SUMB_42__15_) );
  NAND3_X2 u5_mult_82_U5309 ( .A1(u5_mult_82_n5990), .A2(u5_mult_82_n5989), 
        .A3(u5_mult_82_n5988), .ZN(u5_mult_82_CARRYB_49__12_) );
  NAND3_X1 u5_mult_82_U5308 ( .A1(u5_mult_82_n5087), .A2(u5_mult_82_n5088), 
        .A3(u5_mult_82_n5089), .ZN(u5_mult_82_n1495) );
  INV_X2 u5_mult_82_U5307 ( .A(u5_mult_82_SUMB_45__19_), .ZN(u5_mult_82_n1492)
         );
  CLKBUF_X2 u5_mult_82_U5306 ( .A(u5_mult_82_SUMB_32__9_), .Z(u5_mult_82_n1490) );
  XNOR2_X2 u5_mult_82_U5305 ( .A(u5_mult_82_ab_32__12_), .B(
        u5_mult_82_CARRYB_31__12_), .ZN(u5_mult_82_n1489) );
  XNOR2_X2 u5_mult_82_U5304 ( .A(u5_mult_82_n1489), .B(u5_mult_82_SUMB_31__13_), .ZN(u5_mult_82_SUMB_32__12_) );
  XNOR2_X2 u5_mult_82_U5303 ( .A(u5_mult_82_n1758), .B(u5_mult_82_n1582), .ZN(
        u5_mult_82_SUMB_20__31_) );
  XNOR2_X1 u5_mult_82_U5302 ( .A(u5_mult_82_SUMB_32__24_), .B(
        u5_mult_82_ab_33__23_), .ZN(u5_mult_82_n1487) );
  XNOR2_X2 u5_mult_82_U5301 ( .A(u5_mult_82_n1727), .B(u5_mult_82_n1487), .ZN(
        u5_mult_82_SUMB_33__23_) );
  NAND3_X2 u5_mult_82_U5300 ( .A1(u5_mult_82_n6344), .A2(u5_mult_82_n6343), 
        .A3(u5_mult_82_n6342), .ZN(u5_mult_82_CARRYB_23__31_) );
  INV_X4 u5_mult_82_U5299 ( .A(u5_mult_82_n1485), .ZN(u5_mult_82_n1486) );
  INV_X2 u5_mult_82_U5298 ( .A(u5_mult_82_SUMB_40__10_), .ZN(u5_mult_82_n1485)
         );
  XNOR2_X2 u5_mult_82_U5297 ( .A(u5_mult_82_CARRYB_27__29_), .B(
        u5_mult_82_ab_28__29_), .ZN(u5_mult_82_n1483) );
  XNOR2_X2 u5_mult_82_U5296 ( .A(u5_mult_82_n1809), .B(u5_mult_82_n1483), .ZN(
        u5_mult_82_SUMB_28__29_) );
  XNOR2_X2 u5_mult_82_U5295 ( .A(u5_mult_82_n1647), .B(u5_mult_82_n1482), .ZN(
        u5_mult_82_SUMB_35__26_) );
  NAND2_X4 u5_mult_82_U5294 ( .A1(u5_mult_82_n3651), .A2(u5_mult_82_n3650), 
        .ZN(u5_mult_82_n5959) );
  NAND3_X2 u5_mult_82_U5293 ( .A1(u5_mult_82_n4527), .A2(u5_mult_82_n4528), 
        .A3(u5_mult_82_n4529), .ZN(u5_mult_82_n1481) );
  INV_X4 u5_mult_82_U5292 ( .A(u5_mult_82_n1480), .ZN(u5_mult_82_SUMB_14__49_)
         );
  XNOR2_X2 u5_mult_82_U5291 ( .A(u5_mult_82_n4322), .B(u5_mult_82_SUMB_13__50_), .ZN(u5_mult_82_n1480) );
  CLKBUF_X3 u5_mult_82_U5290 ( .A(u5_mult_82_SUMB_34__28_), .Z(
        u5_mult_82_n1479) );
  XNOR2_X2 u5_mult_82_U5289 ( .A(u5_mult_82_ab_19__25_), .B(
        u5_mult_82_CARRYB_18__25_), .ZN(u5_mult_82_n1478) );
  XNOR2_X2 u5_mult_82_U5288 ( .A(u5_mult_82_n37), .B(u5_mult_82_n1478), .ZN(
        u5_mult_82_SUMB_19__25_) );
  XNOR2_X1 u5_mult_82_U5287 ( .A(u5_mult_82_ab_26__9_), .B(
        u5_mult_82_CARRYB_25__9_), .ZN(u5_mult_82_n1476) );
  XNOR2_X2 u5_mult_82_U5286 ( .A(u5_mult_82_n1476), .B(u5_mult_82_n1694), .ZN(
        u5_mult_82_SUMB_26__9_) );
  INV_X2 u5_mult_82_U5285 ( .A(u5_mult_82_CARRYB_37__30_), .ZN(
        u5_mult_82_n1474) );
  XNOR2_X1 u5_mult_82_U5284 ( .A(u5_mult_82_ab_21__13_), .B(
        u5_mult_82_CARRYB_20__13_), .ZN(u5_mult_82_n1473) );
  XNOR2_X2 u5_mult_82_U5283 ( .A(u5_mult_82_n1473), .B(u5_mult_82_SUMB_20__14_), .ZN(u5_mult_82_SUMB_21__13_) );
  XNOR2_X2 u5_mult_82_U5282 ( .A(u5_mult_82_ab_7__37_), .B(
        u5_mult_82_CARRYB_6__37_), .ZN(u5_mult_82_n1472) );
  XNOR2_X2 u5_mult_82_U5281 ( .A(u5_mult_82_n1472), .B(u5_mult_82_SUMB_6__38_), 
        .ZN(u5_mult_82_SUMB_7__37_) );
  XNOR2_X2 u5_mult_82_U5280 ( .A(u5_mult_82_n1471), .B(u5_mult_82_SUMB_40__11_), .ZN(u5_mult_82_SUMB_41__10_) );
  XNOR2_X2 u5_mult_82_U5279 ( .A(u5_mult_82_n1470), .B(u5_mult_82_SUMB_38__17_), .ZN(u5_mult_82_SUMB_39__16_) );
  XNOR2_X2 u5_mult_82_U5278 ( .A(u5_mult_82_SUMB_41__10_), .B(u5_mult_82_n5959), .ZN(u5_mult_82_n1469) );
  XNOR2_X2 u5_mult_82_U5277 ( .A(u5_mult_82_CARRYB_4__47_), .B(
        u5_mult_82_ab_5__47_), .ZN(u5_mult_82_n1467) );
  XNOR2_X2 u5_mult_82_U5276 ( .A(u5_mult_82_SUMB_4__48_), .B(u5_mult_82_n1467), 
        .ZN(u5_mult_82_SUMB_5__47_) );
  INV_X32 u5_mult_82_U5275 ( .A(n4772), .ZN(u5_mult_82_n6820) );
  NOR2_X4 u5_mult_82_U5274 ( .A1(u5_mult_82_net64219), .A2(u5_mult_82_n6820), 
        .ZN(u5_mult_82_ab_0__41_) );
  XNOR2_X2 u5_mult_82_U5273 ( .A(u5_mult_82_CARRYB_20__23_), .B(
        u5_mult_82_ab_21__23_), .ZN(u5_mult_82_n1466) );
  XNOR2_X1 u5_mult_82_U5272 ( .A(u5_mult_82_ab_12__39_), .B(
        u5_mult_82_CARRYB_11__39_), .ZN(u5_mult_82_n1465) );
  XNOR2_X2 u5_mult_82_U5271 ( .A(u5_mult_82_n1465), .B(u5_mult_82_SUMB_11__40_), .ZN(u5_mult_82_SUMB_12__39_) );
  NAND3_X2 u5_mult_82_U5270 ( .A1(u5_mult_82_n2673), .A2(u5_mult_82_n2674), 
        .A3(u5_mult_82_n2675), .ZN(u5_mult_82_CARRYB_32__8_) );
  XNOR2_X2 u5_mult_82_U5269 ( .A(u5_mult_82_ab_29__12_), .B(
        u5_mult_82_CARRYB_28__12_), .ZN(u5_mult_82_n1464) );
  XNOR2_X2 u5_mult_82_U5268 ( .A(u5_mult_82_n1464), .B(u5_mult_82_SUMB_28__13_), .ZN(u5_mult_82_SUMB_29__12_) );
  NAND2_X1 u5_mult_82_U5267 ( .A1(u5_mult_82_CARRYB_17__33_), .A2(
        u5_mult_82_SUMB_17__34_), .ZN(u5_mult_82_n3645) );
  XNOR2_X2 u5_mult_82_U5266 ( .A(u5_mult_82_n1463), .B(u5_mult_82_n1626), .ZN(
        u5_mult_82_SUMB_19__33_) );
  CLKBUF_X2 u5_mult_82_U5265 ( .A(u5_mult_82_SUMB_6__43_), .Z(u5_mult_82_n1462) );
  XNOR2_X2 u5_mult_82_U5264 ( .A(u5_mult_82_ab_33__8_), .B(
        u5_mult_82_CARRYB_32__8_), .ZN(u5_mult_82_n1461) );
  XNOR2_X2 u5_mult_82_U5263 ( .A(u5_mult_82_n1461), .B(u5_mult_82_n1490), .ZN(
        u5_mult_82_SUMB_33__8_) );
  CLKBUF_X2 u5_mult_82_U5262 ( .A(u5_mult_82_CARRYB_10__40_), .Z(
        u5_mult_82_n1460) );
  XNOR2_X2 u5_mult_82_U5261 ( .A(u5_mult_82_CARRYB_31__8_), .B(
        u5_mult_82_ab_32__8_), .ZN(u5_mult_82_n1459) );
  XNOR2_X2 u5_mult_82_U5260 ( .A(u5_mult_82_n1683), .B(u5_mult_82_n1459), .ZN(
        u5_mult_82_SUMB_32__8_) );
  NAND2_X2 u5_mult_82_U5259 ( .A1(u5_mult_82_ab_21__13_), .A2(
        u5_mult_82_SUMB_20__14_), .ZN(u5_mult_82_n2468) );
  XNOR2_X2 u5_mult_82_U5258 ( .A(u5_mult_82_ab_50__20_), .B(
        u5_mult_82_CARRYB_49__20_), .ZN(u5_mult_82_n1457) );
  XNOR2_X2 u5_mult_82_U5257 ( .A(u5_mult_82_n1457), .B(u5_mult_82_SUMB_49__21_), .ZN(u5_mult_82_SUMB_50__20_) );
  XNOR2_X2 u5_mult_82_U5256 ( .A(u5_mult_82_n1614), .B(u5_mult_82_ab_28__33_), 
        .ZN(u5_mult_82_n1456) );
  XNOR2_X2 u5_mult_82_U5255 ( .A(u5_mult_82_n1456), .B(u5_mult_82_SUMB_27__34_), .ZN(u5_mult_82_SUMB_28__33_) );
  NAND2_X1 u5_mult_82_U5254 ( .A1(u5_mult_82_CARRYB_24__43_), .A2(
        u5_mult_82_SUMB_24__44_), .ZN(u5_mult_82_n2577) );
  XOR2_X2 u5_mult_82_U5253 ( .A(u5_mult_82_CARRYB_35__24_), .B(
        u5_mult_82_n3744), .Z(u5_mult_82_n1455) );
  XNOR2_X2 u5_mult_82_U5252 ( .A(u5_mult_82_n1455), .B(u5_mult_82_SUMB_35__25_), .ZN(u5_mult_82_SUMB_36__24_) );
  XNOR2_X2 u5_mult_82_U5251 ( .A(u5_mult_82_CARRYB_19__14_), .B(
        u5_mult_82_ab_20__14_), .ZN(u5_mult_82_n1453) );
  XNOR2_X2 u5_mult_82_U5250 ( .A(u5_mult_82_SUMB_19__15_), .B(u5_mult_82_n1453), .ZN(u5_mult_82_SUMB_20__14_) );
  INV_X4 u5_mult_82_U5249 ( .A(u5_mult_82_n1451), .ZN(u5_mult_82_n1452) );
  INV_X2 u5_mult_82_U5248 ( .A(u5_mult_82_SUMB_8__39_), .ZN(u5_mult_82_n1451)
         );
  NAND2_X1 u5_mult_82_U5247 ( .A1(u5_mult_82_CARRYB_33__14_), .A2(
        u5_mult_82_SUMB_33__15_), .ZN(u5_mult_82_n4953) );
  NAND2_X1 u5_mult_82_U5246 ( .A1(u5_mult_82_ab_20__33_), .A2(
        u5_mult_82_SUMB_19__34_), .ZN(u5_mult_82_n4816) );
  XNOR2_X1 u5_mult_82_U5245 ( .A(u5_mult_82_CARRYB_45__22_), .B(
        u5_mult_82_ab_46__22_), .ZN(u5_mult_82_n1448) );
  XNOR2_X2 u5_mult_82_U5244 ( .A(u5_mult_82_n3772), .B(u5_mult_82_n1448), .ZN(
        u5_mult_82_SUMB_46__22_) );
  CLKBUF_X2 u5_mult_82_U5243 ( .A(u5_mult_82_SUMB_41__24_), .Z(
        u5_mult_82_n1447) );
  NAND2_X1 u5_mult_82_U5242 ( .A1(u5_mult_82_CARRYB_15__33_), .A2(
        u5_mult_82_SUMB_15__34_), .ZN(u5_mult_82_n6047) );
  XNOR2_X2 u5_mult_82_U5241 ( .A(u5_mult_82_ab_7__39_), .B(
        u5_mult_82_CARRYB_6__39_), .ZN(u5_mult_82_n1446) );
  XNOR2_X2 u5_mult_82_U5240 ( .A(u5_mult_82_n1446), .B(u5_mult_82_n1592), .ZN(
        u5_mult_82_SUMB_7__39_) );
  XNOR2_X2 u5_mult_82_U5239 ( .A(u5_mult_82_ab_17__37_), .B(
        u5_mult_82_CARRYB_16__37_), .ZN(u5_mult_82_n1445) );
  XNOR2_X2 u5_mult_82_U5238 ( .A(u5_mult_82_n1445), .B(u5_mult_82_SUMB_16__38_), .ZN(u5_mult_82_SUMB_17__37_) );
  CLKBUF_X2 u5_mult_82_U5237 ( .A(u5_mult_82_CARRYB_37__21_), .Z(
        u5_mult_82_n1444) );
  XNOR2_X2 u5_mult_82_U5236 ( .A(u5_mult_82_CARRYB_31__28_), .B(
        u5_mult_82_ab_32__28_), .ZN(u5_mult_82_n1443) );
  NAND2_X2 u5_mult_82_U5235 ( .A1(u5_mult_82_ab_4__35_), .A2(
        u5_mult_82_net86966), .ZN(u5_mult_82_n5156) );
  NAND3_X2 u5_mult_82_U5234 ( .A1(u5_mult_82_n2469), .A2(u5_mult_82_n2468), 
        .A3(u5_mult_82_n2467), .ZN(u5_mult_82_CARRYB_21__13_) );
  NAND2_X1 u5_mult_82_U5233 ( .A1(u5_mult_82_ab_12__17_), .A2(
        u5_mult_82_SUMB_11__18_), .ZN(u5_mult_82_n1971) );
  NAND3_X2 u5_mult_82_U5232 ( .A1(u5_mult_82_n5767), .A2(u5_mult_82_n5768), 
        .A3(u5_mult_82_n5769), .ZN(u5_mult_82_CARRYB_26__33_) );
  NAND2_X2 u5_mult_82_U5231 ( .A1(u5_mult_82_n1415), .A2(
        u5_mult_82_CARRYB_27__32_), .ZN(u5_mult_82_n6114) );
  XNOR2_X2 u5_mult_82_U5230 ( .A(u5_mult_82_CARRYB_3__34_), .B(
        u5_mult_82_ab_4__34_), .ZN(u5_mult_82_net88132) );
  BUF_X16 u5_mult_82_U5229 ( .A(u5_mult_82_CARRYB_20__49_), .Z(
        u5_mult_82_n1442) );
  XNOR2_X2 u5_mult_82_U5228 ( .A(u5_mult_82_ab_52__32_), .B(
        u5_mult_82_CARRYB_51__32_), .ZN(u5_mult_82_n1440) );
  XNOR2_X2 u5_mult_82_U5227 ( .A(u5_mult_82_n1440), .B(u5_mult_82_SUMB_51__33_), .ZN(u5_mult_82_SUMB_52__32_) );
  XNOR2_X2 u5_mult_82_U5226 ( .A(u5_mult_82_CARRYB_13__26_), .B(
        u5_mult_82_ab_14__26_), .ZN(u5_mult_82_n1439) );
  XNOR2_X2 u5_mult_82_U5225 ( .A(u5_mult_82_SUMB_13__27_), .B(u5_mult_82_n1439), .ZN(u5_mult_82_SUMB_14__26_) );
  INV_X1 u5_mult_82_U5224 ( .A(u5_mult_82_SUMB_14__49_), .ZN(u5_mult_82_n1438)
         );
  XNOR2_X2 u5_mult_82_U5223 ( .A(u5_mult_82_SUMB_47__24_), .B(u5_mult_82_n1437), .ZN(u5_mult_82_SUMB_48__23_) );
  XNOR2_X2 u5_mult_82_U5222 ( .A(u5_mult_82_CARRYB_41__23_), .B(
        u5_mult_82_ab_42__23_), .ZN(u5_mult_82_n1436) );
  XNOR2_X2 u5_mult_82_U5221 ( .A(u5_mult_82_n1447), .B(u5_mult_82_n1436), .ZN(
        u5_mult_82_SUMB_42__23_) );
  XNOR2_X2 u5_mult_82_U5220 ( .A(u5_mult_82_SUMB_13__49_), .B(
        u5_mult_82_ab_14__48_), .ZN(u5_mult_82_n1658) );
  NAND2_X4 u5_mult_82_U5219 ( .A1(u5_mult_82_n2559), .A2(u5_mult_82_n2560), 
        .ZN(u5_mult_82_SUMB_24__9_) );
  FA_X1 u5_mult_82_U5218 ( .A(u5_mult_82_ab_25__8_), .B(
        u5_mult_82_CARRYB_24__8_), .CI(u5_mult_82_SUMB_24__9_), .CO(
        u5_mult_82_n1435) );
  XNOR2_X2 u5_mult_82_U5217 ( .A(u5_mult_82_n2409), .B(u5_mult_82_n438), .ZN(
        u5_mult_82_SUMB_46__17_) );
  CLKBUF_X3 u5_mult_82_U5216 ( .A(u5_mult_82_SUMB_46__17_), .Z(
        u5_mult_82_n1433) );
  NAND2_X2 u5_mult_82_U5215 ( .A1(u5_mult_82_ab_36__22_), .A2(
        u5_mult_82_SUMB_35__23_), .ZN(u5_mult_82_n6217) );
  CLKBUF_X2 u5_mult_82_U5214 ( .A(u5_mult_82_SUMB_40__33_), .Z(
        u5_mult_82_n1431) );
  XNOR2_X2 u5_mult_82_U5213 ( .A(u5_mult_82_n1430), .B(
        u5_mult_82_CARRYB_24__43_), .ZN(u5_mult_82_n2573) );
  XNOR2_X2 u5_mult_82_U5212 ( .A(u5_mult_82_n1718), .B(u5_mult_82_SUMB_33__23_), .ZN(u5_mult_82_SUMB_34__22_) );
  XNOR2_X2 u5_mult_82_U5211 ( .A(u5_mult_82_CARRYB_47__23_), .B(
        u5_mult_82_ab_48__23_), .ZN(u5_mult_82_n1437) );
  XNOR2_X2 u5_mult_82_U5210 ( .A(u5_mult_82_ab_40__11_), .B(
        u5_mult_82_CARRYB_39__11_), .ZN(u5_mult_82_n1429) );
  XNOR2_X2 u5_mult_82_U5209 ( .A(u5_mult_82_n1429), .B(u5_mult_82_SUMB_39__12_), .ZN(u5_mult_82_SUMB_40__11_) );
  XNOR2_X1 u5_mult_82_U5208 ( .A(u5_mult_82_SUMB_15__26_), .B(u5_mult_82_n3273), .ZN(u5_mult_82_SUMB_16__25_) );
  INV_X4 u5_mult_82_U5207 ( .A(u5_mult_82_n1427), .ZN(u5_mult_82_n1428) );
  INV_X2 u5_mult_82_U5206 ( .A(u5_mult_82_SUMB_25__30_), .ZN(u5_mult_82_n1427)
         );
  CLKBUF_X3 u5_mult_82_U5205 ( .A(u5_mult_82_SUMB_38__11_), .Z(
        u5_mult_82_n1426) );
  NAND2_X2 u5_mult_82_U5204 ( .A1(u5_mult_82_CARRYB_16__24_), .A2(
        u5_mult_82_SUMB_16__25_), .ZN(u5_mult_82_n5324) );
  NAND2_X2 u5_mult_82_U5203 ( .A1(u5_mult_82_ab_17__24_), .A2(
        u5_mult_82_SUMB_16__25_), .ZN(u5_mult_82_n5323) );
  INV_X2 u5_mult_82_U5202 ( .A(u5_mult_82_n1424), .ZN(u5_mult_82_n1425) );
  INV_X1 u5_mult_82_U5201 ( .A(u5_mult_82_CARRYB_41__24_), .ZN(
        u5_mult_82_n1424) );
  XNOR2_X2 u5_mult_82_U5200 ( .A(u5_mult_82_ab_38__20_), .B(
        u5_mult_82_CARRYB_37__20_), .ZN(u5_mult_82_n1423) );
  XNOR2_X2 u5_mult_82_U5199 ( .A(u5_mult_82_n1423), .B(u5_mult_82_SUMB_37__21_), .ZN(u5_mult_82_SUMB_38__20_) );
  XNOR2_X2 u5_mult_82_U5198 ( .A(u5_mult_82_SUMB_20__21_), .B(u5_mult_82_n4163), .ZN(u5_mult_82_SUMB_21__20_) );
  XNOR2_X2 u5_mult_82_U5197 ( .A(u5_mult_82_CARRYB_31__14_), .B(
        u5_mult_82_ab_32__14_), .ZN(u5_mult_82_n1421) );
  XNOR2_X2 u5_mult_82_U5196 ( .A(u5_mult_82_SUMB_31__15_), .B(u5_mult_82_n1421), .ZN(u5_mult_82_SUMB_32__14_) );
  XNOR2_X2 u5_mult_82_U5195 ( .A(u5_mult_82_n1843), .B(u5_mult_82_n4622), .ZN(
        u5_mult_82_n1419) );
  INV_X4 u5_mult_82_U5194 ( .A(u5_mult_82_n1418), .ZN(u5_mult_82_SUMB_47__16_)
         );
  XNOR2_X2 u5_mult_82_U5193 ( .A(u5_mult_82_n5860), .B(u5_mult_82_n1433), .ZN(
        u5_mult_82_n1418) );
  XNOR2_X2 u5_mult_82_U5192 ( .A(u5_mult_82_CARRYB_37__7_), .B(
        u5_mult_82_ab_38__7_), .ZN(u5_mult_82_n1417) );
  XNOR2_X2 u5_mult_82_U5191 ( .A(u5_mult_82_n1417), .B(u5_mult_82_n55), .ZN(
        u5_mult_82_SUMB_38__7_) );
  CLKBUF_X2 u5_mult_82_U5190 ( .A(u5_mult_82_SUMB_50__34_), .Z(
        u5_mult_82_n1416) );
  XNOR2_X2 u5_mult_82_U5189 ( .A(u5_mult_82_ab_39__7_), .B(
        u5_mult_82_CARRYB_38__7_), .ZN(u5_mult_82_n1759) );
  INV_X2 u5_mult_82_U5188 ( .A(u5_mult_82_SUMB_27__33_), .ZN(u5_mult_82_n1414)
         );
  INV_X4 u5_mult_82_U5187 ( .A(u5_mult_82_CARRYB_38__11_), .ZN(
        u5_mult_82_n3697) );
  INV_X1 u5_mult_82_U5186 ( .A(u5_mult_82_n3697), .ZN(u5_mult_82_n1413) );
  CLKBUF_X2 u5_mult_82_U5185 ( .A(u5_mult_82_CARRYB_42__39_), .Z(
        u5_mult_82_n1412) );
  BUF_X2 u5_mult_82_U5184 ( .A(u5_mult_82_SUMB_45__5_), .Z(u5_mult_82_n1411)
         );
  XNOR2_X2 u5_mult_82_U5183 ( .A(u5_mult_82_ab_23__37_), .B(
        u5_mult_82_CARRYB_22__37_), .ZN(u5_mult_82_n1410) );
  NAND2_X2 u5_mult_82_U5182 ( .A1(u5_mult_82_CARRYB_28__9_), .A2(
        u5_mult_82_n399), .ZN(u5_mult_82_n2827) );
  NAND2_X2 u5_mult_82_U5181 ( .A1(u5_mult_82_ab_29__9_), .A2(u5_mult_82_n399), 
        .ZN(u5_mult_82_n2826) );
  XNOR2_X2 u5_mult_82_U5180 ( .A(u5_mult_82_n3667), .B(u5_mult_82_n1611), .ZN(
        u5_mult_82_SUMB_48__22_) );
  XNOR2_X2 u5_mult_82_U5179 ( .A(u5_mult_82_n1409), .B(u5_mult_82_SUMB_47__25_), .ZN(u5_mult_82_SUMB_48__24_) );
  INV_X4 u5_mult_82_U5178 ( .A(u5_mult_82_n1407), .ZN(u5_mult_82_n1408) );
  INV_X2 u5_mult_82_U5177 ( .A(u5_mult_82_SUMB_44__28_), .ZN(u5_mult_82_n1407)
         );
  NAND2_X1 u5_mult_82_U5176 ( .A1(u5_mult_82_ab_37__20_), .A2(
        u5_mult_82_SUMB_36__21_), .ZN(u5_mult_82_n5186) );
  XNOR2_X2 u5_mult_82_U5175 ( .A(u5_mult_82_CARRYB_23__37_), .B(
        u5_mult_82_n1406), .ZN(u5_mult_82_SUMB_24__37_) );
  XNOR2_X2 u5_mult_82_U5174 ( .A(u5_mult_82_CARRYB_49__3_), .B(
        u5_mult_82_ab_50__3_), .ZN(u5_mult_82_n1405) );
  XNOR2_X2 u5_mult_82_U5173 ( .A(u5_mult_82_SUMB_49__4_), .B(u5_mult_82_n1405), 
        .ZN(u5_mult_82_SUMB_50__3_) );
  NAND2_X1 u5_mult_82_U5172 ( .A1(u5_mult_82_ab_27__35_), .A2(
        u5_mult_82_SUMB_26__36_), .ZN(u5_mult_82_n4933) );
  XNOR2_X2 u5_mult_82_U5171 ( .A(u5_mult_82_n4787), .B(u5_mult_82_n4101), .ZN(
        u5_mult_82_n1404) );
  XNOR2_X2 u5_mult_82_U5170 ( .A(u5_mult_82_SUMB_18__45_), .B(u5_mult_82_n1403), .ZN(u5_mult_82_SUMB_19__44_) );
  INV_X2 u5_mult_82_U5169 ( .A(u5_mult_82_n1401), .ZN(u5_mult_82_n1402) );
  INV_X1 u5_mult_82_U5168 ( .A(u5_mult_82_CARRYB_49__0_), .ZN(u5_mult_82_n1401) );
  XNOR2_X2 u5_mult_82_U5167 ( .A(u5_mult_82_n1400), .B(u5_mult_82_SUMB_6__42_), 
        .ZN(u5_mult_82_SUMB_7__41_) );
  INV_X4 u5_mult_82_U5166 ( .A(u5_mult_82_n1398), .ZN(u5_mult_82_n1399) );
  INV_X2 u5_mult_82_U5165 ( .A(u5_mult_82_SUMB_33__21_), .ZN(u5_mult_82_n1398)
         );
  XNOR2_X1 u5_mult_82_U5164 ( .A(u5_mult_82_ab_25__39_), .B(
        u5_mult_82_CARRYB_24__39_), .ZN(u5_mult_82_n1397) );
  XNOR2_X2 u5_mult_82_U5163 ( .A(u5_mult_82_n1397), .B(u5_mult_82_SUMB_24__40_), .ZN(u5_mult_82_SUMB_25__39_) );
  XNOR2_X2 u5_mult_82_U5162 ( .A(u5_mult_82_ab_15__42_), .B(
        u5_mult_82_CARRYB_14__42_), .ZN(u5_mult_82_n1396) );
  XNOR2_X2 u5_mult_82_U5161 ( .A(u5_mult_82_n1396), .B(u5_mult_82_SUMB_14__43_), .ZN(u5_mult_82_SUMB_15__42_) );
  INV_X4 u5_mult_82_U5160 ( .A(u5_mult_82_n1394), .ZN(u5_mult_82_n1395) );
  NAND2_X2 u5_mult_82_U5159 ( .A1(u5_mult_82_SUMB_24__10_), .A2(
        u5_mult_82_CARRYB_24__9_), .ZN(u5_mult_82_n3437) );
  NAND2_X2 u5_mult_82_U5158 ( .A1(u5_mult_82_ab_25__9_), .A2(
        u5_mult_82_SUMB_24__10_), .ZN(u5_mult_82_n3435) );
  XNOR2_X2 u5_mult_82_U5157 ( .A(u5_mult_82_CARRYB_38__24_), .B(
        u5_mult_82_ab_39__24_), .ZN(u5_mult_82_n1393) );
  XNOR2_X2 u5_mult_82_U5156 ( .A(u5_mult_82_n1393), .B(u5_mult_82_n1812), .ZN(
        u5_mult_82_SUMB_39__24_) );
  CLKBUF_X2 u5_mult_82_U5155 ( .A(u5_mult_82_SUMB_14__50_), .Z(
        u5_mult_82_n1392) );
  XNOR2_X2 u5_mult_82_U5154 ( .A(u5_mult_82_SUMB_38__21_), .B(u5_mult_82_n1391), .ZN(u5_mult_82_SUMB_39__20_) );
  XNOR2_X2 u5_mult_82_U5153 ( .A(u5_mult_82_ab_29__27_), .B(
        u5_mult_82_CARRYB_28__27_), .ZN(u5_mult_82_n1389) );
  XNOR2_X1 u5_mult_82_U5152 ( .A(u5_mult_82_n1389), .B(u5_mult_82_n20), .ZN(
        u5_mult_82_SUMB_29__27_) );
  CLKBUF_X2 u5_mult_82_U5151 ( .A(u5_mult_82_CARRYB_48__13_), .Z(
        u5_mult_82_n1388) );
  XNOR2_X2 u5_mult_82_U5150 ( .A(u5_mult_82_n1603), .B(u5_mult_82_n1384), .ZN(
        u5_mult_82_n1386) );
  XNOR2_X2 u5_mult_82_U5149 ( .A(u5_mult_82_ab_30__23_), .B(
        u5_mult_82_CARRYB_29__23_), .ZN(u5_mult_82_n1385) );
  XNOR2_X2 u5_mult_82_U5148 ( .A(u5_mult_82_n1385), .B(u5_mult_82_SUMB_29__24_), .ZN(u5_mult_82_SUMB_30__23_) );
  NAND3_X2 u5_mult_82_U5147 ( .A1(u5_mult_82_n3618), .A2(u5_mult_82_n3619), 
        .A3(u5_mult_82_n3620), .ZN(u5_mult_82_CARRYB_26__9_) );
  INV_X4 u5_mult_82_U5146 ( .A(u5_mult_82_n1383), .ZN(u5_mult_82_n1384) );
  INV_X2 u5_mult_82_U5145 ( .A(u5_mult_82_SUMB_10__39_), .ZN(u5_mult_82_n1383)
         );
  NAND2_X2 u5_mult_82_U5144 ( .A1(u5_mult_82_ab_16__15_), .A2(
        u5_mult_82_CARRYB_15__15_), .ZN(u5_mult_82_n3802) );
  XOR2_X2 u5_mult_82_U5143 ( .A(u5_mult_82_n4300), .B(u5_mult_82_SUMB_41__18_), 
        .Z(u5_mult_82_n1382) );
  XNOR2_X2 u5_mult_82_U5142 ( .A(u5_mult_82_n1382), .B(
        u5_mult_82_CARRYB_41__17_), .ZN(u5_mult_82_SUMB_42__17_) );
  INV_X16 u5_mult_82_U5141 ( .A(n4764), .ZN(u5_mult_82_n7015) );
  FA_X1 u5_mult_82_U5140 ( .A(u5_mult_82_ab_2__37_), .B(
        u5_mult_82_CARRYB_1__37_), .CI(u5_mult_82_SUMB_1__38_), .S(
        u5_mult_82_net88595) );
  INV_X32 u5_mult_82_U5139 ( .A(u5_mult_82_n1379), .ZN(u5_mult_82_net64677) );
  INV_X32 u5_mult_82_U5138 ( .A(n4750), .ZN(u5_mult_82_n1379) );
  INV_X32 u5_mult_82_U5137 ( .A(u5_mult_82_n1378), .ZN(u5_mult_82_net64671) );
  INV_X32 u5_mult_82_U5136 ( .A(u5_mult_82_n1379), .ZN(u5_mult_82_n1378) );
  INV_X32 u5_mult_82_U5135 ( .A(u5_mult_82_n1378), .ZN(u5_mult_82_net64669) );
  INV_X32 u5_mult_82_U5134 ( .A(u5_mult_82_n1380), .ZN(u5_mult_82_net65679) );
  INV_X32 u5_mult_82_U5133 ( .A(u5_mult_82_net64569), .ZN(u5_mult_82_net64559)
         );
  INV_X32 u5_mult_82_U5132 ( .A(u5_mult_82_net64497), .ZN(u5_mult_82_net64487)
         );
  NOR2_X4 u5_mult_82_U5131 ( .A1(u5_mult_82_net64487), .A2(u5_mult_82_net65391), .ZN(u5_mult_82_ab_41__12_) );
  NAND2_X2 u5_mult_82_U5130 ( .A1(u5_mult_82_ab_41__12_), .A2(
        u5_mult_82_SUMB_40__13_), .ZN(u5_mult_82_net86289) );
  XNOR2_X2 u5_mult_82_U5129 ( .A(u5_mult_82_n1377), .B(u5_mult_82_SUMB_39__14_), .ZN(u5_mult_82_SUMB_40__13_) );
  INV_X32 u5_mult_82_U5128 ( .A(u5_mult_82_n1374), .ZN(u5_mult_82_net65353) );
  INV_X32 u5_mult_82_U5127 ( .A(u5_mult_82_n1374), .ZN(u5_mult_82_net65355) );
  NAND2_X1 u5_mult_82_U5126 ( .A1(u5_mult_82_ab_43__10_), .A2(
        u5_mult_82_CARRYB_42__10_), .ZN(u5_mult_82_n1376) );
  NOR2_X4 u5_mult_82_U5125 ( .A1(u5_mult_82_net64455), .A2(u5_mult_82_net65355), .ZN(u5_mult_82_ab_43__10_) );
  NAND3_X4 u5_mult_82_U5124 ( .A1(u5_mult_82_net78857), .A2(
        u5_mult_82_net78856), .A3(u5_mult_82_n1376), .ZN(
        u5_mult_82_CARRYB_43__10_) );
  NAND2_X1 u5_mult_82_U5123 ( .A1(u5_mult_82_net79209), .A2(
        u5_mult_82_net86976), .ZN(u5_mult_82_n1368) );
  INV_X4 u5_mult_82_U5122 ( .A(u5_mult_82_net79209), .ZN(u5_mult_82_net82042)
         );
  NAND2_X2 u5_mult_82_U5121 ( .A1(u5_mult_82_net87269), .A2(
        u5_mult_82_SUMB_29__20_), .ZN(u5_mult_82_net79215) );
  NAND2_X2 u5_mult_82_U5120 ( .A1(u5_mult_82_ab_30__19_), .A2(
        u5_mult_82_SUMB_29__20_), .ZN(u5_mult_82_net79214) );
  INV_X4 u5_mult_82_U5119 ( .A(u5_mult_82_net86976), .ZN(
        u5_mult_82_SUMB_29__20_) );
  NAND2_X2 u5_mult_82_U5118 ( .A1(u5_mult_82_net82042), .A2(
        u5_mult_82_SUMB_29__20_), .ZN(u5_mult_82_n1369) );
  NAND2_X4 u5_mult_82_U5117 ( .A1(u5_mult_82_n1368), .A2(u5_mult_82_n1369), 
        .ZN(u5_mult_82_SUMB_30__19_) );
  INV_X2 u5_mult_82_U5116 ( .A(u5_mult_82_ab_31__18_), .ZN(u5_mult_82_net86279) );
  NAND2_X4 u5_mult_82_U5115 ( .A1(u5_mult_82_net86279), .A2(
        u5_mult_82_net86280), .ZN(u5_mult_82_n1371) );
  NAND2_X2 u5_mult_82_U5114 ( .A1(u5_mult_82_net86281), .A2(u5_mult_82_n1371), 
        .ZN(u5_mult_82_n1370) );
  NAND2_X2 u5_mult_82_U5113 ( .A1(u5_mult_82_ab_32__17_), .A2(
        u5_mult_82_SUMB_31__18_), .ZN(u5_mult_82_net83292) );
  NAND2_X2 u5_mult_82_U5112 ( .A1(u5_mult_82_CARRYB_31__17_), .A2(
        u5_mult_82_SUMB_31__18_), .ZN(u5_mult_82_net83293) );
  XNOR2_X2 u5_mult_82_U5111 ( .A(u5_mult_82_n1370), .B(u5_mult_82_SUMB_30__19_), .ZN(u5_mult_82_SUMB_31__18_) );
  INV_X32 u5_mult_82_U5110 ( .A(u5_mult_82_n1357), .ZN(u5_mult_82_net64903) );
  INV_X16 u5_mult_82_U5109 ( .A(u5_mult_82_net64913), .ZN(u5_mult_82_n1357) );
  INV_X32 u5_mult_82_U5108 ( .A(u5_mult_82_n1357), .ZN(u5_mult_82_net64905) );
  INV_X32 u5_mult_82_U5107 ( .A(u5_mult_82_n1358), .ZN(u5_mult_82_net66017) );
  NAND2_X1 u5_mult_82_U5106 ( .A1(u5_mult_82_ab_5__35_), .A2(
        u5_mult_82_CARRYB_4__35_), .ZN(u5_mult_82_n1360) );
  NAND2_X2 u5_mult_82_U5105 ( .A1(u5_mult_82_n288), .A2(u5_mult_82_ab_5__35_), 
        .ZN(u5_mult_82_n1361) );
  NAND2_X2 u5_mult_82_U5104 ( .A1(u5_mult_82_n288), .A2(
        u5_mult_82_CARRYB_4__35_), .ZN(u5_mult_82_n1362) );
  NAND3_X4 u5_mult_82_U5103 ( .A1(u5_mult_82_n1360), .A2(u5_mult_82_n1361), 
        .A3(u5_mult_82_n1362), .ZN(u5_mult_82_CARRYB_5__35_) );
  INV_X4 u5_mult_82_U5102 ( .A(u5_mult_82_CARRYB_4__36_), .ZN(u5_mult_82_n1365) );
  NAND2_X4 u5_mult_82_U5101 ( .A1(u5_mult_82_n1367), .A2(u5_mult_82_n1366), 
        .ZN(u5_mult_82_n1363) );
  XNOR2_X2 u5_mult_82_U5100 ( .A(u5_mult_82_n1363), .B(u5_mult_82_SUMB_4__37_), 
        .ZN(u5_mult_82_SUMB_5__36_) );
  INV_X32 u5_mult_82_U5099 ( .A(u5_mult_82_n1351), .ZN(u5_mult_82_net65443) );
  NAND3_X2 u5_mult_82_U5098 ( .A1(u5_mult_82_net79087), .A2(
        u5_mult_82_net79088), .A3(u5_mult_82_net79089), .ZN(
        u5_mult_82_CARRYB_37__14_) );
  INV_X1 u5_mult_82_U5097 ( .A(u5_mult_82_ab_37__15_), .ZN(u5_mult_82_n1354)
         );
  NAND2_X4 u5_mult_82_U5096 ( .A1(u5_mult_82_n1355), .A2(u5_mult_82_n1354), 
        .ZN(u5_mult_82_n1356) );
  XNOR2_X2 u5_mult_82_U5095 ( .A(u5_mult_82_n1353), .B(u5_mult_82_SUMB_36__16_), .ZN(u5_mult_82_SUMB_37__15_) );
  XNOR2_X2 u5_mult_82_U5094 ( .A(u5_mult_82_CARRYB_38__14_), .B(
        u5_mult_82_ab_39__14_), .ZN(u5_mult_82_net83655) );
  INV_X4 u5_mult_82_U5093 ( .A(fracta_mul[51]), .ZN(u5_mult_82_n1349) );
  XNOR2_X2 u5_mult_82_U5092 ( .A(u5_mult_82_ab_50__7_), .B(
        u5_mult_82_CARRYB_49__7_), .ZN(u5_mult_82_n1350) );
  NAND2_X2 u5_mult_82_U5091 ( .A1(u5_mult_82_ab_51__6_), .A2(
        u5_mult_82_SUMB_50__7_), .ZN(u5_mult_82_net80807) );
  XNOR2_X2 u5_mult_82_U5090 ( .A(u5_mult_82_n1350), .B(u5_mult_82_SUMB_49__8_), 
        .ZN(u5_mult_82_SUMB_50__7_) );
  NAND2_X1 u5_mult_82_U5089 ( .A1(u5_mult_82_ab_22__24_), .A2(
        u5_mult_82_SUMB_21__25_), .ZN(u5_mult_82_net81531) );
  XNOR2_X2 u5_mult_82_U5088 ( .A(u5_mult_82_net87435), .B(
        u5_mult_82_SUMB_20__26_), .ZN(u5_mult_82_SUMB_21__25_) );
  INV_X8 u5_mult_82_U5087 ( .A(n4754), .ZN(u5_mult_82_n1342) );
  INV_X32 u5_mult_82_U5086 ( .A(u5_mult_82_n1342), .ZN(u5_mult_82_net64695) );
  INV_X32 u5_mult_82_U5085 ( .A(u5_mult_82_net64695), .ZN(u5_mult_82_net64689)
         );
  INV_X32 u5_mult_82_U5084 ( .A(u5_mult_82_net64695), .ZN(u5_mult_82_net64687)
         );
  NOR2_X4 u5_mult_82_U5083 ( .A1(u5_mult_82_net64687), .A2(u5_mult_82_net65713), .ZN(u5_mult_82_ab_23__23_) );
  NAND3_X2 u5_mult_82_U5082 ( .A1(u5_mult_82_n1345), .A2(u5_mult_82_n1346), 
        .A3(u5_mult_82_n1347), .ZN(u5_mult_82_CARRYB_22__23_) );
  XNOR2_X2 u5_mult_82_U5081 ( .A(u5_mult_82_SUMB_21__25_), .B(u5_mult_82_n1348), .ZN(u5_mult_82_SUMB_22__24_) );
  NAND2_X1 u5_mult_82_U5080 ( .A1(u5_mult_82_ab_24__23_), .A2(
        u5_mult_82_CARRYB_23__23_), .ZN(u5_mult_82_net84199) );
  INV_X32 u5_mult_82_U5079 ( .A(u5_mult_82_net65287), .ZN(u5_mult_82_net65283)
         );
  NAND2_X1 u5_mult_82_U5078 ( .A1(u5_mult_82_ab_46__8_), .A2(
        u5_mult_82_CARRYB_45__8_), .ZN(u5_mult_82_n1336) );
  NAND2_X2 u5_mult_82_U5077 ( .A1(u5_mult_82_ab_46__8_), .A2(
        u5_mult_82_SUMB_45__9_), .ZN(u5_mult_82_n1337) );
  NAND2_X2 u5_mult_82_U5076 ( .A1(u5_mult_82_CARRYB_45__8_), .A2(
        u5_mult_82_SUMB_45__9_), .ZN(u5_mult_82_n1338) );
  NAND3_X2 u5_mult_82_U5075 ( .A1(u5_mult_82_n1336), .A2(u5_mult_82_n1337), 
        .A3(u5_mult_82_n1338), .ZN(u5_mult_82_CARRYB_46__8_) );
  NAND2_X2 u5_mult_82_U5074 ( .A1(u5_mult_82_CARRYB_47__8_), .A2(
        u5_mult_82_SUMB_47__9_), .ZN(u5_mult_82_net81827) );
  XNOR2_X2 u5_mult_82_U5073 ( .A(u5_mult_82_n1341), .B(u5_mult_82_net81962), 
        .ZN(u5_mult_82_SUMB_48__7_) );
  NAND2_X2 u5_mult_82_U5072 ( .A1(u5_mult_82_ab_48__7_), .A2(u5_mult_82_n1341), 
        .ZN(u5_mult_82_n1333) );
  INV_X4 u5_mult_82_U5071 ( .A(u5_mult_82_n1340), .ZN(u5_mult_82_n1341) );
  NAND2_X2 u5_mult_82_U5070 ( .A1(u5_mult_82_CARRYB_47__7_), .A2(
        u5_mult_82_n1341), .ZN(u5_mult_82_n1334) );
  NAND2_X1 u5_mult_82_U5069 ( .A1(u5_mult_82_ab_49__7_), .A2(
        u5_mult_82_CARRYB_48__7_), .ZN(u5_mult_82_net81828) );
  NAND3_X4 u5_mult_82_U5068 ( .A1(u5_mult_82_n1334), .A2(u5_mult_82_n1333), 
        .A3(u5_mult_82_net78954), .ZN(u5_mult_82_CARRYB_48__7_) );
  XNOR2_X1 u5_mult_82_U5067 ( .A(u5_mult_82_ab_48__8_), .B(
        u5_mult_82_CARRYB_47__8_), .ZN(u5_mult_82_n1339) );
  NAND2_X2 u5_mult_82_U5066 ( .A1(u5_mult_82_ab_49__7_), .A2(
        u5_mult_82_SUMB_48__8_), .ZN(u5_mult_82_net81829) );
  XNOR2_X2 u5_mult_82_U5065 ( .A(u5_mult_82_n1339), .B(u5_mult_82_SUMB_47__9_), 
        .ZN(u5_mult_82_SUMB_48__8_) );
  XNOR2_X2 u5_mult_82_U5064 ( .A(u5_mult_82_CARRYB_48__7_), .B(
        u5_mult_82_n1335), .ZN(u5_mult_82_net81824) );
  INV_X32 u5_mult_82_U5063 ( .A(u5_mult_82_net65521), .ZN(u5_mult_82_net65515)
         );
  XOR2_X2 u5_mult_82_U5062 ( .A(u5_mult_82_CARRYB_32__17_), .B(
        u5_mult_82_ab_33__17_), .Z(u5_mult_82_n1332) );
  XOR2_X2 u5_mult_82_U5061 ( .A(u5_mult_82_SUMB_32__18_), .B(u5_mult_82_n1332), 
        .Z(u5_mult_82_SUMB_33__17_) );
  NAND2_X1 u5_mult_82_U5060 ( .A1(u5_mult_82_ab_36__15_), .A2(
        u5_mult_82_CARRYB_35__15_), .ZN(u5_mult_82_net79084) );
  NAND2_X2 u5_mult_82_U5059 ( .A1(u5_mult_82_n716), .A2(u5_mult_82_n483), .ZN(
        u5_mult_82_net79086) );
  NAND2_X2 u5_mult_82_U5058 ( .A1(u5_mult_82_ab_37__13_), .A2(
        u5_mult_82_SUMB_36__14_), .ZN(u5_mult_82_net82056) );
  NAND2_X2 u5_mult_82_U5057 ( .A1(u5_mult_82_CARRYB_36__13_), .A2(
        u5_mult_82_SUMB_36__14_), .ZN(u5_mult_82_net82055) );
  XNOR2_X2 u5_mult_82_U5056 ( .A(u5_mult_82_SUMB_36__14_), .B(
        u5_mult_82_net83047), .ZN(u5_mult_82_SUMB_37__13_) );
  NAND2_X1 u5_mult_82_U5055 ( .A1(u5_mult_82_ab_37__14_), .A2(
        u5_mult_82_CARRYB_36__14_), .ZN(u5_mult_82_net79087) );
  XNOR2_X2 u5_mult_82_U5054 ( .A(u5_mult_82_CARRYB_35__15_), .B(
        u5_mult_82_net83710), .ZN(u5_mult_82_net79082) );
  NAND2_X1 u5_mult_82_U5053 ( .A1(u5_mult_82_ab_37__14_), .A2(
        u5_mult_82_SUMB_36__15_), .ZN(u5_mult_82_net79088) );
  NAND2_X1 u5_mult_82_U5052 ( .A1(u5_mult_82_CARRYB_36__14_), .A2(
        u5_mult_82_SUMB_36__15_), .ZN(u5_mult_82_net79089) );
  XOR2_X2 u5_mult_82_U5051 ( .A(u5_mult_82_net79082), .B(u5_mult_82_n483), .Z(
        u5_mult_82_SUMB_36__15_) );
  NAND2_X1 u5_mult_82_U5050 ( .A1(u5_mult_82_net81198), .A2(
        u5_mult_82_CARRYB_36__14_), .ZN(u5_mult_82_net81422) );
  INV_X2 u5_mult_82_U5049 ( .A(u5_mult_82_ab_37__14_), .ZN(u5_mult_82_net81198) );
  NAND2_X2 u5_mult_82_U5048 ( .A1(u5_mult_82_ab_37__14_), .A2(
        u5_mult_82_net81421), .ZN(u5_mult_82_n1331) );
  NAND2_X4 u5_mult_82_U5047 ( .A1(u5_mult_82_net81422), .A2(u5_mult_82_n1331), 
        .ZN(u5_mult_82_n1330) );
  NAND2_X2 u5_mult_82_U5046 ( .A1(u5_mult_82_ab_38__13_), .A2(
        u5_mult_82_SUMB_37__14_), .ZN(u5_mult_82_net81427) );
  NAND2_X2 u5_mult_82_U5045 ( .A1(u5_mult_82_CARRYB_37__13_), .A2(
        u5_mult_82_SUMB_37__14_), .ZN(u5_mult_82_net81428) );
  CLKBUF_X3 u5_mult_82_U5044 ( .A(u5_mult_82_SUMB_37__14_), .Z(
        u5_mult_82_net87325) );
  XOR2_X2 u5_mult_82_U5043 ( .A(u5_mult_82_n1330), .B(u5_mult_82_SUMB_36__15_), 
        .Z(u5_mult_82_SUMB_37__14_) );
  XOR2_X2 u5_mult_82_U5042 ( .A(u5_mult_82_ab_7__35_), .B(
        u5_mult_82_CARRYB_6__35_), .Z(u5_mult_82_net80183) );
  NAND2_X1 u5_mult_82_U5041 ( .A1(u5_mult_82_ab_7__35_), .A2(
        u5_mult_82_CARRYB_6__35_), .ZN(u5_mult_82_net80185) );
  NAND2_X2 u5_mult_82_U5040 ( .A1(u5_mult_82_n34), .A2(u5_mult_82_SUMB_6__36_), 
        .ZN(u5_mult_82_net80187) );
  NAND2_X1 u5_mult_82_U5039 ( .A1(u5_mult_82_ab_8__34_), .A2(
        u5_mult_82_CARRYB_7__34_), .ZN(u5_mult_82_net80188) );
  NAND2_X1 u5_mult_82_U5038 ( .A1(u5_mult_82_CARRYB_7__34_), .A2(
        u5_mult_82_SUMB_7__35_), .ZN(u5_mult_82_net80190) );
  NAND2_X1 u5_mult_82_U5037 ( .A1(u5_mult_82_ab_14__29_), .A2(
        u5_mult_82_CARRYB_13__29_), .ZN(u5_mult_82_net80254) );
  XNOR2_X2 u5_mult_82_U5036 ( .A(u5_mult_82_CARRYB_13__29_), .B(
        u5_mult_82_ab_14__29_), .ZN(u5_mult_82_net80786) );
  INV_X2 u5_mult_82_U5035 ( .A(u5_mult_82_SUMB_15__27_), .ZN(
        u5_mult_82_net86784) );
  NAND2_X1 u5_mult_82_U5034 ( .A1(u5_mult_82_CARRYB_15__27_), .A2(
        u5_mult_82_SUMB_15__28_), .ZN(u5_mult_82_net81534) );
  NAND2_X1 u5_mult_82_U5033 ( .A1(u5_mult_82_ab_16__27_), .A2(
        u5_mult_82_CARRYB_15__27_), .ZN(u5_mult_82_net81536) );
  INV_X32 u5_mult_82_U5032 ( .A(u5_mult_82_net64515), .ZN(u5_mult_82_net64505)
         );
  INV_X4 u5_mult_82_U5031 ( .A(fracta_mul[41]), .ZN(u5_mult_82_n1325) );
  INV_X32 u5_mult_82_U5030 ( .A(u5_mult_82_n1326), .ZN(u5_mult_82_net65389) );
  INV_X32 u5_mult_82_U5029 ( .A(u5_mult_82_n1326), .ZN(u5_mult_82_net65391) );
  XNOR2_X2 u5_mult_82_U5028 ( .A(u5_mult_82_ab_40__14_), .B(
        u5_mult_82_CARRYB_39__14_), .ZN(u5_mult_82_n1329) );
  XNOR2_X2 u5_mult_82_U5027 ( .A(u5_mult_82_n1329), .B(u5_mult_82_SUMB_39__15_), .ZN(u5_mult_82_SUMB_40__14_) );
  XOR2_X2 u5_mult_82_U5026 ( .A(u5_mult_82_ab_42__13_), .B(
        u5_mult_82_CARRYB_41__13_), .Z(u5_mult_82_net80793) );
  NAND2_X1 u5_mult_82_U5025 ( .A1(u5_mult_82_ab_42__13_), .A2(
        u5_mult_82_CARRYB_41__13_), .ZN(u5_mult_82_net80795) );
  NAND2_X2 u5_mult_82_U5024 ( .A1(u5_mult_82_CARRYB_41__13_), .A2(
        u5_mult_82_SUMB_41__14_), .ZN(u5_mult_82_net80797) );
  NAND2_X1 u5_mult_82_U5023 ( .A1(u5_mult_82_ab_44__11_), .A2(
        u5_mult_82_CARRYB_43__11_), .ZN(u5_mult_82_net79446) );
  NAND2_X1 u5_mult_82_U5022 ( .A1(u5_mult_82_SUMB_43__12_), .A2(
        u5_mult_82_CARRYB_43__11_), .ZN(u5_mult_82_net79444) );
  INV_X32 u5_mult_82_U5021 ( .A(u5_mult_82_n1318), .ZN(u5_mult_82_net64469) );
  INV_X32 u5_mult_82_U5020 ( .A(u5_mult_82_n1320), .ZN(u5_mult_82_net65371) );
  INV_X32 u5_mult_82_U5019 ( .A(u5_mult_82_n1321), .ZN(u5_mult_82_n1320) );
  INV_X32 u5_mult_82_U5018 ( .A(u5_mult_82_n1320), .ZN(u5_mult_82_net65373) );
  NOR2_X1 u5_mult_82_U5017 ( .A1(u5_mult_82_net64469), .A2(u5_mult_82_net65373), .ZN(u5_mult_82_ab_42__11_) );
  NAND2_X2 u5_mult_82_U5016 ( .A1(u5_mult_82_SUMB_40__12_), .A2(
        u5_mult_82_CARRYB_40__11_), .ZN(u5_mult_82_n1322) );
  NAND2_X2 u5_mult_82_U5015 ( .A1(u5_mult_82_ab_41__11_), .A2(
        u5_mult_82_CARRYB_40__11_), .ZN(u5_mult_82_n1323) );
  NAND2_X1 u5_mult_82_U5014 ( .A1(u5_mult_82_ab_41__11_), .A2(
        u5_mult_82_SUMB_40__12_), .ZN(u5_mult_82_n1324) );
  NAND2_X2 u5_mult_82_U5013 ( .A1(u5_mult_82_ab_42__11_), .A2(
        u5_mult_82_CARRYB_41__11_), .ZN(u5_mult_82_net78852) );
  NAND3_X2 u5_mult_82_U5012 ( .A1(u5_mult_82_n1322), .A2(u5_mult_82_n1323), 
        .A3(u5_mult_82_n1324), .ZN(u5_mult_82_CARRYB_41__11_) );
  NAND2_X1 u5_mult_82_U5011 ( .A1(u5_mult_82_CARRYB_41__11_), .A2(
        u5_mult_82_SUMB_41__12_), .ZN(u5_mult_82_net78850) );
  NAND2_X2 u5_mult_82_U5010 ( .A1(u5_mult_82_ab_42__11_), .A2(
        u5_mult_82_SUMB_41__12_), .ZN(u5_mult_82_net78851) );
  XOR2_X2 u5_mult_82_U5009 ( .A(u5_mult_82_net86284), .B(
        u5_mult_82_SUMB_40__13_), .Z(u5_mult_82_SUMB_41__12_) );
  XNOR2_X2 u5_mult_82_U5008 ( .A(u5_mult_82_CARRYB_41__11_), .B(
        u5_mult_82_ab_42__11_), .ZN(u5_mult_82_net83870) );
  NAND2_X1 u5_mult_82_U5007 ( .A1(u5_mult_82_CARRYB_42__10_), .A2(
        u5_mult_82_SUMB_42__11_), .ZN(u5_mult_82_net78857) );
  INV_X1 u5_mult_82_U5006 ( .A(u5_mult_82_SUMB_42__11_), .ZN(
        u5_mult_82_net84441) );
  NAND2_X2 u5_mult_82_U5005 ( .A1(u5_mult_82_net84440), .A2(
        u5_mult_82_SUMB_42__11_), .ZN(u5_mult_82_net84443) );
  XNOR2_X2 u5_mult_82_U5004 ( .A(u5_mult_82_SUMB_41__12_), .B(
        u5_mult_82_net83870), .ZN(u5_mult_82_SUMB_42__11_) );
  INV_X1 u5_mult_82_U5003 ( .A(u5_mult_82_SUMB_14__30_), .ZN(u5_mult_82_n1311)
         );
  NAND2_X1 u5_mult_82_U5002 ( .A1(u5_mult_82_n1311), .A2(u5_mult_82_net80255), 
        .ZN(u5_mult_82_n1312) );
  NAND2_X2 u5_mult_82_U5001 ( .A1(u5_mult_82_net82040), .A2(u5_mult_82_n1312), 
        .ZN(u5_mult_82_SUMB_15__29_) );
  NAND2_X2 u5_mult_82_U5000 ( .A1(u5_mult_82_CARRYB_16__28_), .A2(
        u5_mult_82_SUMB_16__29_), .ZN(u5_mult_82_net80537) );
  NAND2_X2 u5_mult_82_U4999 ( .A1(u5_mult_82_ab_17__28_), .A2(
        u5_mult_82_CARRYB_16__28_), .ZN(u5_mult_82_net80535) );
  INV_X2 u5_mult_82_U4998 ( .A(u5_mult_82_SUMB_16__28_), .ZN(u5_mult_82_n1313)
         );
  NAND2_X4 u5_mult_82_U4997 ( .A1(u5_mult_82_ab_17__27_), .A2(u5_mult_82_n1314), .ZN(u5_mult_82_net79786) );
  NAND2_X2 u5_mult_82_U4996 ( .A1(u5_mult_82_CARRYB_16__27_), .A2(
        u5_mult_82_n1314), .ZN(u5_mult_82_net79785) );
  XNOR2_X2 u5_mult_82_U4995 ( .A(u5_mult_82_CARRYB_16__27_), .B(
        u5_mult_82_ab_17__27_), .ZN(u5_mult_82_n1309) );
  XNOR2_X2 u5_mult_82_U4994 ( .A(u5_mult_82_n1314), .B(u5_mult_82_n1309), .ZN(
        u5_mult_82_SUMB_17__27_) );
  XNOR2_X2 u5_mult_82_U4993 ( .A(u5_mult_82_ab_18__27_), .B(
        u5_mult_82_CARRYB_17__27_), .ZN(u5_mult_82_n1310) );
  XNOR2_X2 u5_mult_82_U4992 ( .A(u5_mult_82_n1310), .B(u5_mult_82_SUMB_17__28_), .ZN(u5_mult_82_SUMB_18__27_) );
  NAND2_X1 u5_mult_82_U4991 ( .A1(u5_mult_82_CARRYB_19__26_), .A2(
        u5_mult_82_ab_20__26_), .ZN(u5_mult_82_net85540) );
  XNOR2_X2 u5_mult_82_U4990 ( .A(u5_mult_82_CARRYB_19__26_), .B(
        u5_mult_82_ab_20__26_), .ZN(u5_mult_82_net86085) );
  INV_X2 u5_mult_82_U4989 ( .A(u5_mult_82_SUMB_19__26_), .ZN(u5_mult_82_n1316)
         );
  NAND2_X2 u5_mult_82_U4988 ( .A1(u5_mult_82_ab_20__25_), .A2(u5_mult_82_n1317), .ZN(u5_mult_82_net84194) );
  NAND2_X2 u5_mult_82_U4987 ( .A1(u5_mult_82_CARRYB_19__25_), .A2(
        u5_mult_82_n1317), .ZN(u5_mult_82_net84193) );
  INV_X8 u5_mult_82_U4986 ( .A(u5_mult_82_n1316), .ZN(u5_mult_82_n1317) );
  XNOR2_X2 u5_mult_82_U4985 ( .A(u5_mult_82_CARRYB_19__25_), .B(
        u5_mult_82_ab_20__25_), .ZN(u5_mult_82_n1315) );
  NAND2_X2 u5_mult_82_U4984 ( .A1(u5_mult_82_SUMB_20__25_), .A2(
        u5_mult_82_ab_21__24_), .ZN(u5_mult_82_net80543) );
  NAND2_X1 u5_mult_82_U4983 ( .A1(u5_mult_82_CARRYB_26__21_), .A2(
        u5_mult_82_SUMB_26__22_), .ZN(u5_mult_82_net80645) );
  NAND2_X1 u5_mult_82_U4982 ( .A1(u5_mult_82_ab_27__21_), .A2(
        u5_mult_82_CARRYB_26__21_), .ZN(u5_mult_82_net80647) );
  XNOR2_X2 u5_mult_82_U4981 ( .A(u5_mult_82_CARRYB_26__21_), .B(
        u5_mult_82_ab_27__21_), .ZN(u5_mult_82_net82990) );
  NAND2_X2 u5_mult_82_U4980 ( .A1(u5_mult_82_CARRYB_27__19_), .A2(
        u5_mult_82_n715), .ZN(u5_mult_82_net82047) );
  XOR2_X2 u5_mult_82_U4979 ( .A(u5_mult_82_n715), .B(u5_mult_82_net82046), .Z(
        u5_mult_82_SUMB_28__19_) );
  NAND2_X2 u5_mult_82_U4978 ( .A1(u5_mult_82_n715), .A2(u5_mult_82_ab_28__19_), 
        .ZN(u5_mult_82_net82048) );
  XOR2_X2 u5_mult_82_U4977 ( .A(u5_mult_82_ab_29__20_), .B(
        u5_mult_82_CARRYB_28__20_), .Z(u5_mult_82_net79208) );
  NAND2_X1 u5_mult_82_U4976 ( .A1(u5_mult_82_ab_29__20_), .A2(
        u5_mult_82_CARRYB_28__20_), .ZN(u5_mult_82_net79210) );
  NAND2_X2 u5_mult_82_U4975 ( .A1(u5_mult_82_CARRYB_28__20_), .A2(
        u5_mult_82_SUMB_28__21_), .ZN(u5_mult_82_net79212) );
  NAND2_X1 u5_mult_82_U4974 ( .A1(u5_mult_82_ab_30__19_), .A2(
        u5_mult_82_CARRYB_29__19_), .ZN(u5_mult_82_net79213) );
  XNOR2_X2 u5_mult_82_U4973 ( .A(u5_mult_82_net80364), .B(
        u5_mult_82_CARRYB_29__19_), .ZN(u5_mult_82_net79209) );
  CLKBUF_X3 u5_mult_82_U4972 ( .A(u5_mult_82_CARRYB_29__19_), .Z(
        u5_mult_82_net87269) );
  NAND2_X2 u5_mult_82_U4971 ( .A1(u5_mult_82_ab_30__18_), .A2(
        u5_mult_82_SUMB_29__19_), .ZN(u5_mult_82_n1307) );
  NAND2_X2 u5_mult_82_U4970 ( .A1(u5_mult_82_SUMB_29__19_), .A2(
        u5_mult_82_CARRYB_29__18_), .ZN(u5_mult_82_n1308) );
  NAND2_X1 u5_mult_82_U4969 ( .A1(u5_mult_82_ab_31__18_), .A2(
        u5_mult_82_CARRYB_30__18_), .ZN(u5_mult_82_net83288) );
  INV_X4 u5_mult_82_U4968 ( .A(u5_mult_82_CARRYB_30__18_), .ZN(
        u5_mult_82_net86280) );
  NAND2_X1 u5_mult_82_U4967 ( .A1(u5_mult_82_CARRYB_30__18_), .A2(
        u5_mult_82_SUMB_30__19_), .ZN(u5_mult_82_net83290) );
  NAND2_X2 u5_mult_82_U4966 ( .A1(u5_mult_82_CARRYB_30__18_), .A2(
        u5_mult_82_ab_31__18_), .ZN(u5_mult_82_net86281) );
  NAND3_X2 u5_mult_82_U4965 ( .A1(u5_mult_82_net79263), .A2(u5_mult_82_n1307), 
        .A3(u5_mult_82_n1308), .ZN(u5_mult_82_CARRYB_30__18_) );
  XOR2_X2 u5_mult_82_U4964 ( .A(u5_mult_82_ab_5__35_), .B(
        u5_mult_82_CARRYB_4__35_), .Z(u5_mult_82_n1306) );
  XOR2_X2 u5_mult_82_U4963 ( .A(u5_mult_82_n1306), .B(u5_mult_82_n288), .Z(
        u5_mult_82_SUMB_5__35_) );
  XOR2_X2 u5_mult_82_U4962 ( .A(u5_mult_82_SUMB_6__34_), .B(
        u5_mult_82_net85371), .Z(u5_mult_82_SUMB_7__33_) );
  NAND2_X1 u5_mult_82_U4961 ( .A1(u5_mult_82_CARRYB_6__33_), .A2(
        u5_mult_82_SUMB_6__34_), .ZN(u5_mult_82_net85372) );
  NAND2_X2 u5_mult_82_U4960 ( .A1(u5_mult_82_ab_7__33_), .A2(
        u5_mult_82_SUMB_6__34_), .ZN(u5_mult_82_net85373) );
  NAND2_X1 u5_mult_82_U4959 ( .A1(u5_mult_82_ab_4__35_), .A2(
        u5_mult_82_SUMB_3__36_), .ZN(u5_mult_82_net80618) );
  NAND2_X2 u5_mult_82_U4958 ( .A1(u5_mult_82_net86966), .A2(
        u5_mult_82_SUMB_3__36_), .ZN(u5_mult_82_net80619) );
  XNOR2_X2 u5_mult_82_U4957 ( .A(u5_mult_82_net85323), .B(
        u5_mult_82_SUMB_2__37_), .ZN(u5_mult_82_SUMB_3__36_) );
  INV_X16 u5_mult_82_U4956 ( .A(n4786), .ZN(u5_mult_82_net57160) );
  INV_X32 u5_mult_82_U4955 ( .A(u5_mult_82_net57160), .ZN(u5_mult_82_net64893)
         );
  INV_X32 u5_mult_82_U4954 ( .A(u5_mult_82_net64893), .ZN(u5_mult_82_net64885)
         );
  INV_X32 u5_mult_82_U4953 ( .A(u5_mult_82_net64893), .ZN(u5_mult_82_net64887)
         );
  INV_X4 u5_mult_82_U4952 ( .A(fracta_mul[5]), .ZN(u5_mult_82_n1301) );
  INV_X32 u5_mult_82_U4951 ( .A(u5_mult_82_n1303), .ZN(u5_mult_82_net66043) );
  INV_X32 u5_mult_82_U4950 ( .A(u5_mult_82_n1304), .ZN(u5_mult_82_n1303) );
  INV_X32 u5_mult_82_U4949 ( .A(u5_mult_82_n1302), .ZN(u5_mult_82_net66033) );
  INV_X32 u5_mult_82_U4948 ( .A(u5_mult_82_n1303), .ZN(u5_mult_82_n1302) );
  INV_X32 u5_mult_82_U4947 ( .A(u5_mult_82_n1302), .ZN(u5_mult_82_net66035) );
  NAND2_X2 u5_mult_82_U4946 ( .A1(u5_mult_82_ab_4__34_), .A2(
        u5_mult_82_CARRYB_3__34_), .ZN(u5_mult_82_n1305) );
  NAND3_X2 u5_mult_82_U4945 ( .A1(u5_mult_82_net83295), .A2(
        u5_mult_82_net83296), .A3(u5_mult_82_n1305), .ZN(
        u5_mult_82_CARRYB_4__34_) );
  XOR2_X2 u5_mult_82_U4944 ( .A(u5_mult_82_net80613), .B(
        u5_mult_82_SUMB_3__36_), .Z(u5_mult_82_SUMB_4__35_) );
  NAND2_X2 u5_mult_82_U4943 ( .A1(u5_mult_82_SUMB_48__7_), .A2(
        u5_mult_82_net84845), .ZN(u5_mult_82_n1299) );
  INV_X2 u5_mult_82_U4942 ( .A(u5_mult_82_SUMB_48__7_), .ZN(
        u5_mult_82_net86159) );
  INV_X4 u5_mult_82_U4941 ( .A(u5_mult_82_net84845), .ZN(u5_mult_82_n1298) );
  NAND2_X1 u5_mult_82_U4940 ( .A1(u5_mult_82_ab_52__5_), .A2(
        u5_mult_82_CARRYB_51__5_), .ZN(u5_mult_82_net78792) );
  INV_X1 u5_mult_82_U4939 ( .A(u5_mult_82_SUMB_50__7_), .ZN(
        u5_mult_82_net87846) );
  INV_X2 u5_mult_82_U4938 ( .A(u5_mult_82_net87846), .ZN(u5_mult_82_net87847)
         );
  NAND2_X1 u5_mult_82_U4937 ( .A1(u5_mult_82_CARRYB_51__5_), .A2(
        u5_mult_82_SUMB_51__6_), .ZN(u5_mult_82_net78790) );
  NAND2_X1 u5_mult_82_U4936 ( .A1(u5_mult_82_ab_52__5_), .A2(
        u5_mult_82_SUMB_51__6_), .ZN(u5_mult_82_net78791) );
  XOR2_X2 u5_mult_82_U4935 ( .A(u5_mult_82_net80802), .B(u5_mult_82_net87847), 
        .Z(u5_mult_82_SUMB_51__6_) );
  XNOR2_X2 u5_mult_82_U4934 ( .A(u5_mult_82_CARRYB_51__5_), .B(
        u5_mult_82_net87687), .ZN(u5_mult_82_net78789) );
  XNOR2_X2 u5_mult_82_U4933 ( .A(u5_mult_82_CARRYB_52__4_), .B(
        u5_mult_82_SUMB_52__5_), .ZN(u5_mult_82__UDW__89408_net70938) );
  XOR2_X2 u5_mult_82_U4932 ( .A(u5_mult_82_SUMB_51__6_), .B(
        u5_mult_82_net78789), .Z(u5_mult_82_SUMB_52__5_) );
  INV_X32 u5_mult_82_U4931 ( .A(u5_mult_82_n1289), .ZN(u5_mult_82_net64441) );
  INV_X32 u5_mult_82_U4930 ( .A(u5_mult_82_n1288), .ZN(u5_mult_82_net64433) );
  INV_X4 u5_mult_82_U4929 ( .A(fracta_mul[45]), .ZN(u5_mult_82_n1287) );
  INV_X32 u5_mult_82_U4928 ( .A(u5_mult_82_n1290), .ZN(u5_mult_82_net65321) );
  INV_X32 u5_mult_82_U4927 ( .A(u5_mult_82_n1290), .ZN(u5_mult_82_net65319) );
  NOR2_X4 u5_mult_82_U4926 ( .A1(u5_mult_82_net64433), .A2(u5_mult_82_net65319), .ZN(u5_mult_82_ab_45__9_) );
  XOR2_X2 u5_mult_82_U4925 ( .A(u5_mult_82_ab_44__10_), .B(
        u5_mult_82_CARRYB_43__10_), .Z(u5_mult_82_n1296) );
  XOR2_X2 u5_mult_82_U4924 ( .A(u5_mult_82_SUMB_43__11_), .B(u5_mult_82_n1296), 
        .Z(u5_mult_82_SUMB_44__10_) );
  NAND2_X2 u5_mult_82_U4923 ( .A1(u5_mult_82_net84599), .A2(
        u5_mult_82_SUMB_43__10_), .ZN(u5_mult_82_n1295) );
  NAND2_X2 u5_mult_82_U4922 ( .A1(u5_mult_82_ab_44__9_), .A2(
        u5_mult_82_SUMB_43__10_), .ZN(u5_mult_82_n1294) );
  NAND2_X2 u5_mult_82_U4921 ( .A1(u5_mult_82_ab_44__9_), .A2(
        u5_mult_82_net84599), .ZN(u5_mult_82_n1293) );
  XNOR2_X2 u5_mult_82_U4920 ( .A(u5_mult_82_CARRYB_44__9_), .B(
        u5_mult_82_ab_45__9_), .ZN(u5_mult_82_net83142) );
  NAND3_X4 u5_mult_82_U4919 ( .A1(u5_mult_82_n1295), .A2(u5_mult_82_n1294), 
        .A3(u5_mult_82_n1293), .ZN(u5_mult_82_CARRYB_44__9_) );
  NAND2_X1 u5_mult_82_U4918 ( .A1(u5_mult_82_ab_45__9_), .A2(
        u5_mult_82_CARRYB_44__9_), .ZN(u5_mult_82_n1297) );
  NAND2_X1 u5_mult_82_U4917 ( .A1(u5_mult_82_ab_46__9_), .A2(
        u5_mult_82_CARRYB_45__9_), .ZN(u5_mult_82_net84888) );
  NAND2_X2 u5_mult_82_U4916 ( .A1(u5_mult_82_CARRYB_45__9_), .A2(
        u5_mult_82_SUMB_45__10_), .ZN(u5_mult_82_net84890) );
  INV_X32 u5_mult_82_U4915 ( .A(u5_mult_82_net64495), .ZN(u5_mult_82_net64491)
         );
  INV_X32 u5_mult_82_U4914 ( .A(u5_mult_82_net64495), .ZN(u5_mult_82_net64489)
         );
  INV_X4 u5_mult_82_U4913 ( .A(fracta_mul[40]), .ZN(u5_mult_82_n1277) );
  INV_X32 u5_mult_82_U4912 ( .A(u5_mult_82_n1278), .ZN(u5_mult_82_net65411) );
  INV_X32 u5_mult_82_U4911 ( .A(u5_mult_82_n1278), .ZN(u5_mult_82_net65407) );
  INV_X32 u5_mult_82_U4910 ( .A(u5_mult_82_n1279), .ZN(u5_mult_82_n1278) );
  INV_X32 u5_mult_82_U4909 ( .A(u5_mult_82_n1278), .ZN(u5_mult_82_net65409) );
  NOR2_X4 u5_mult_82_U4908 ( .A1(u5_mult_82_net64489), .A2(u5_mult_82_net65409), .ZN(u5_mult_82_ab_40__12_) );
  XNOR2_X2 u5_mult_82_U4907 ( .A(u5_mult_82_net85894), .B(
        u5_mult_82_SUMB_39__13_), .ZN(u5_mult_82_SUMB_40__12_) );
  XOR2_X2 u5_mult_82_U4906 ( .A(u5_mult_82_n1284), .B(u5_mult_82_n1286), .Z(
        u5_mult_82_SUMB_39__13_) );
  NAND2_X1 u5_mult_82_U4905 ( .A1(u5_mult_82_ab_39__12_), .A2(
        u5_mult_82_CARRYB_38__12_), .ZN(u5_mult_82_n1281) );
  NAND2_X2 u5_mult_82_U4904 ( .A1(u5_mult_82_ab_39__12_), .A2(
        u5_mult_82_SUMB_38__13_), .ZN(u5_mult_82_n1282) );
  NAND2_X2 u5_mult_82_U4903 ( .A1(u5_mult_82_SUMB_38__13_), .A2(
        u5_mult_82_CARRYB_38__12_), .ZN(u5_mult_82_n1283) );
  XNOR2_X2 u5_mult_82_U4902 ( .A(u5_mult_82_ab_40__12_), .B(
        u5_mult_82_CARRYB_39__12_), .ZN(u5_mult_82_net85894) );
  NAND3_X4 u5_mult_82_U4901 ( .A1(u5_mult_82_n1281), .A2(u5_mult_82_n1282), 
        .A3(u5_mult_82_n1283), .ZN(u5_mult_82_CARRYB_39__12_) );
  NAND2_X1 u5_mult_82_U4900 ( .A1(u5_mult_82_ab_40__12_), .A2(
        u5_mult_82_CARRYB_39__12_), .ZN(u5_mult_82_n1285) );
  XOR2_X2 u5_mult_82_U4899 ( .A(u5_mult_82_ab_41__12_), .B(
        u5_mult_82_CARRYB_40__12_), .Z(u5_mult_82_net86284) );
  NAND2_X2 u5_mult_82_U4898 ( .A1(u5_mult_82_CARRYB_40__12_), .A2(
        u5_mult_82_SUMB_40__13_), .ZN(u5_mult_82_net86290) );
  NAND3_X2 u5_mult_82_U4897 ( .A1(u5_mult_82_n1285), .A2(u5_mult_82_net82471), 
        .A3(u5_mult_82_net82472), .ZN(u5_mult_82_CARRYB_40__12_) );
  XNOR2_X2 u5_mult_82_U4896 ( .A(u5_mult_82_SUMB_49__7_), .B(
        u5_mult_82_net84846), .ZN(u5_mult_82_SUMB_50__6_) );
  XOR2_X2 u5_mult_82_U4895 ( .A(u5_mult_82_net81824), .B(
        u5_mult_82_SUMB_48__8_), .Z(u5_mult_82_SUMB_49__7_) );
  NAND2_X1 u5_mult_82_U4894 ( .A1(u5_mult_82_ab_49__6_), .A2(
        u5_mult_82_CARRYB_48__6_), .ZN(u5_mult_82_n1274) );
  NAND2_X2 u5_mult_82_U4893 ( .A1(u5_mult_82_ab_49__6_), .A2(
        u5_mult_82_SUMB_48__7_), .ZN(u5_mult_82_n1275) );
  NAND2_X2 u5_mult_82_U4892 ( .A1(u5_mult_82_CARRYB_48__6_), .A2(
        u5_mult_82_SUMB_48__7_), .ZN(u5_mult_82_n1276) );
  NAND3_X4 u5_mult_82_U4891 ( .A1(u5_mult_82_n1274), .A2(u5_mult_82_n1275), 
        .A3(u5_mult_82_n1276), .ZN(u5_mult_82_CARRYB_49__6_) );
  INV_X32 u5_mult_82_U4890 ( .A(u5_mult_82_n1271), .ZN(u5_mult_82_net64387) );
  INV_X32 u5_mult_82_U4889 ( .A(u5_mult_82_n1270), .ZN(u5_mult_82_net64379) );
  INV_X4 u5_mult_82_U4888 ( .A(fracta_mul[50]), .ZN(u5_mult_82_net57179) );
  XNOR2_X2 u5_mult_82_U4887 ( .A(u5_mult_82_CARRYB_49__6_), .B(
        u5_mult_82_ab_50__6_), .ZN(u5_mult_82_net84846) );
  NOR2_X1 u5_mult_82_U4886 ( .A1(u5_mult_82_net64379), .A2(u5_mult_82_net65229), .ZN(u5_mult_82_ab_50__6_) );
  NAND2_X1 u5_mult_82_U4885 ( .A1(u5_mult_82_CARRYB_49__6_), .A2(
        u5_mult_82_SUMB_49__7_), .ZN(u5_mult_82_net78900) );
  NAND2_X1 u5_mult_82_U4884 ( .A1(u5_mult_82_ab_50__6_), .A2(
        u5_mult_82_CARRYB_49__6_), .ZN(u5_mult_82_n1273) );
  XOR2_X2 u5_mult_82_U4883 ( .A(u5_mult_82_ab_51__6_), .B(
        u5_mult_82_CARRYB_50__6_), .Z(u5_mult_82_net80802) );
  NAND2_X1 u5_mult_82_U4882 ( .A1(u5_mult_82_ab_51__6_), .A2(
        u5_mult_82_CARRYB_50__6_), .ZN(u5_mult_82_net80806) );
  NAND2_X2 u5_mult_82_U4881 ( .A1(u5_mult_82_CARRYB_50__6_), .A2(
        u5_mult_82_SUMB_50__7_), .ZN(u5_mult_82_net80808) );
  NAND3_X2 u5_mult_82_U4880 ( .A1(u5_mult_82_net78900), .A2(
        u5_mult_82_net78901), .A3(u5_mult_82_n1273), .ZN(
        u5_mult_82_CARRYB_50__6_) );
  AND2_X2 u5_mult_82_U4879 ( .A1(u5_mult_82_net64225), .A2(n4783), .ZN(
        u5_mult_82_ab_0__37_) );
  NAND2_X2 u5_mult_82_U4878 ( .A1(u5_mult_82_ab_1__36_), .A2(
        u5_mult_82_ab_0__37_), .ZN(u5_mult_82__UDW__88988_net69760) );
  INV_X4 u5_mult_82_U4877 ( .A(u5_mult_82__UDW__88988_net69760), .ZN(
        u5_mult_82_CARRYB_1__36_) );
  NOR2_X1 u5_mult_82_U4876 ( .A1(u5_mult_82_n1263), .A2(u5_mult_82_net66107), 
        .ZN(u5_mult_82_ab_1__36_) );
  INV_X8 u5_mult_82_U4875 ( .A(n4733), .ZN(u5_mult_82_n1263) );
  INV_X4 u5_mult_82_U4874 ( .A(u5_mult_82_n1263), .ZN(u5_mult_82_n1266) );
  INV_X4 u5_mult_82_U4873 ( .A(u5_mult_82_n1266), .ZN(u5_mult_82_n1269) );
  INV_X32 u5_mult_82_U4872 ( .A(u5_mult_82_n1265), .ZN(u5_mult_82_net64923) );
  INV_X32 u5_mult_82_U4871 ( .A(u5_mult_82_n1265), .ZN(u5_mult_82_net64921) );
  INV_X32 u5_mult_82_U4870 ( .A(u5_mult_82_n1268), .ZN(u5_mult_82_net66097) );
  INV_X32 u5_mult_82_U4869 ( .A(u5_mult_82_n1267), .ZN(u5_mult_82_net66087) );
  INV_X32 u5_mult_82_U4868 ( .A(u5_mult_82_n1267), .ZN(u5_mult_82_net66089) );
  XNOR2_X2 u5_mult_82_U4867 ( .A(u5_mult_82_ab_3__36_), .B(
        u5_mult_82_CARRYB_2__36_), .ZN(u5_mult_82_net85323) );
  NAND2_X1 u5_mult_82_U4866 ( .A1(u5_mult_82_ab_3__36_), .A2(
        u5_mult_82_CARRYB_2__36_), .ZN(u5_mult_82_net80614) );
  NAND2_X1 u5_mult_82_U4865 ( .A1(u5_mult_82_CARRYB_2__36_), .A2(
        u5_mult_82_net88595), .ZN(u5_mult_82_net80616) );
  NAND2_X2 u5_mult_82_U4864 ( .A1(u5_mult_82_ab_4__34_), .A2(
        u5_mult_82_SUMB_3__35_), .ZN(u5_mult_82_net83296) );
  XNOR2_X2 u5_mult_82_U4863 ( .A(u5_mult_82_SUMB_3__35_), .B(
        u5_mult_82_net88132), .ZN(u5_mult_82_SUMB_4__34_) );
  XNOR2_X2 u5_mult_82_U4862 ( .A(u5_mult_82_net85316), .B(
        u5_mult_82_CARRYB_3__35_), .ZN(u5_mult_82_net80613) );
  CLKBUF_X2 u5_mult_82_U4861 ( .A(u5_mult_82_CARRYB_3__35_), .Z(
        u5_mult_82_net86966) );
  INV_X16 u5_mult_82_U4860 ( .A(n4815), .ZN(u5_mult_82_net64217) );
  INV_X8 u5_mult_82_U4859 ( .A(n4815), .ZN(u5_mult_82_n1261) );
  NOR2_X1 u5_mult_82_U4858 ( .A1(u5_mult_82_net64219), .A2(u5_mult_82_net64961), .ZN(u5_mult_82_n1251) );
  INV_X32 u5_mult_82_U4857 ( .A(n4822), .ZN(u5_mult_82_net66107) );
  INV_X4 u5_mult_82_U4856 ( .A(u5_mult_82_n1255), .ZN(u5_mult_82_n1258) );
  INV_X4 u5_mult_82_U4855 ( .A(u5_mult_82_n1259), .ZN(u5_mult_82_CARRYB_2__36_) );
  INV_X4 u5_mult_82_U4854 ( .A(u5_mult_82_n1253), .ZN(u5_mult_82_n1252) );
  XNOR2_X2 u5_mult_82_U4853 ( .A(u5_mult_82_n1258), .B(u5_mult_82_n613), .ZN(
        u5_mult_82_n1257) );
  XNOR2_X2 u5_mult_82_U4852 ( .A(u5_mult_82_n1257), .B(u5_mult_82_n1254), .ZN(
        u5_mult_82_SUMB_2__36_) );
  XNOR2_X2 u5_mult_82_U4851 ( .A(u5_mult_82_n1256), .B(u5_mult_82_n1253), .ZN(
        u5_mult_82_n1255) );
  INV_X4 u5_mult_82_U4850 ( .A(u5_mult_82_CARRYB_1__36_), .ZN(u5_mult_82_n1254) );
  NAND2_X2 u5_mult_82_U4849 ( .A1(u5_mult_82_n1251), .A2(u5_mult_82_n1252), 
        .ZN(u5_mult_82__UDW__88983_net69746) );
  NAND2_X2 u5_mult_82_U4848 ( .A1(u5_mult_82_CARRYB_17__35_), .A2(
        u5_mult_82_SUMB_17__36_), .ZN(u5_mult_82_n6315) );
  XNOR2_X2 u5_mult_82_U4847 ( .A(u5_mult_82_SUMB_40__32_), .B(u5_mult_82_n1618), .ZN(u5_mult_82_SUMB_41__31_) );
  XNOR2_X2 u5_mult_82_U4846 ( .A(u5_mult_82_ab_39__15_), .B(
        u5_mult_82_CARRYB_38__15_), .ZN(u5_mult_82_n1250) );
  XNOR2_X2 u5_mult_82_U4845 ( .A(u5_mult_82_n1250), .B(u5_mult_82_SUMB_38__16_), .ZN(u5_mult_82_SUMB_39__15_) );
  INV_X8 u5_mult_82_U4844 ( .A(u5_mult_82_n6403), .ZN(u5_mult_82_CLA_SUM[70])
         );
  NAND2_X2 u5_mult_82_U4843 ( .A1(u5_mult_82_ab_18__35_), .A2(
        u5_mult_82_SUMB_17__36_), .ZN(u5_mult_82_n6314) );
  NAND3_X2 u5_mult_82_U4842 ( .A1(u5_mult_82_n5117), .A2(u5_mult_82_n5116), 
        .A3(u5_mult_82_n5115), .ZN(u5_mult_82_CARRYB_45__27_) );
  NAND2_X2 u5_mult_82_U4841 ( .A1(u5_mult_82_ab_18__45_), .A2(
        u5_mult_82_CARRYB_17__45_), .ZN(u5_mult_82_n5876) );
  NAND2_X1 u5_mult_82_U4840 ( .A1(u5_mult_82_ab_42__31_), .A2(
        u5_mult_82_CARRYB_41__31_), .ZN(u5_mult_82_n3942) );
  NAND2_X1 u5_mult_82_U4839 ( .A1(u5_mult_82_CARRYB_41__31_), .A2(
        u5_mult_82_SUMB_41__32_), .ZN(u5_mult_82_n3944) );
  NAND3_X2 u5_mult_82_U4838 ( .A1(u5_mult_82_n5138), .A2(u5_mult_82_n5139), 
        .A3(u5_mult_82_n5140), .ZN(u5_mult_82_CARRYB_23__25_) );
  NAND2_X2 u5_mult_82_U4837 ( .A1(u5_mult_82_SUMB_13__49_), .A2(
        u5_mult_82_CARRYB_13__48_), .ZN(u5_mult_82_n3377) );
  NAND2_X1 u5_mult_82_U4836 ( .A1(u5_mult_82_ab_44__26_), .A2(
        u5_mult_82_CARRYB_43__26_), .ZN(u5_mult_82_n4923) );
  NAND2_X1 u5_mult_82_U4835 ( .A1(u5_mult_82_CARRYB_49__22_), .A2(
        u5_mult_82_SUMB_49__23_), .ZN(u5_mult_82_n5097) );
  NAND2_X1 u5_mult_82_U4834 ( .A1(u5_mult_82_ab_42__17_), .A2(
        u5_mult_82_SUMB_41__18_), .ZN(u5_mult_82_n5064) );
  NAND2_X2 u5_mult_82_U4833 ( .A1(u5_mult_82_ab_36__34_), .A2(
        u5_mult_82_SUMB_35__35_), .ZN(u5_mult_82_n3929) );
  INV_X8 u5_mult_82_U4832 ( .A(u5_mult_82_n6407), .ZN(u5_mult_82_CLA_SUM[73])
         );
  NAND3_X2 u5_mult_82_U4831 ( .A1(u5_mult_82_n5953), .A2(u5_mult_82_n5954), 
        .A3(u5_mult_82_n5955), .ZN(u5_mult_82_CARRYB_17__47_) );
  NAND2_X1 u5_mult_82_U4830 ( .A1(u5_mult_82_ab_11__37_), .A2(
        u5_mult_82_SUMB_10__38_), .ZN(u5_mult_82_n5455) );
  NAND2_X2 u5_mult_82_U4829 ( .A1(u5_mult_82_SUMB_20__34_), .A2(
        u5_mult_82_CARRYB_20__33_), .ZN(u5_mult_82_n4820) );
  NAND2_X2 u5_mult_82_U4828 ( .A1(u5_mult_82_ab_7__41_), .A2(u5_mult_82_n1510), 
        .ZN(u5_mult_82_n6018) );
  XNOR2_X2 u5_mult_82_U4827 ( .A(u5_mult_82_ab_3__28_), .B(
        u5_mult_82_CARRYB_2__28_), .ZN(u5_mult_82_n1249) );
  XNOR2_X2 u5_mult_82_U4826 ( .A(u5_mult_82_n1249), .B(u5_mult_82_SUMB_2__29_), 
        .ZN(u5_mult_82_SUMB_3__28_) );
  NAND2_X2 u5_mult_82_U4825 ( .A1(u5_mult_82_ab_43__10_), .A2(
        u5_mult_82_SUMB_42__11_), .ZN(u5_mult_82_net78856) );
  NAND2_X2 u5_mult_82_U4824 ( .A1(u5_mult_82_CARRYB_41__4_), .A2(
        u5_mult_82_ab_42__4_), .ZN(u5_mult_82_n4729) );
  NAND2_X2 u5_mult_82_U4823 ( .A1(u5_mult_82_CARRYB_43__19_), .A2(
        u5_mult_82_SUMB_43__20_), .ZN(u5_mult_82_n3235) );
  NAND2_X2 u5_mult_82_U4822 ( .A1(u5_mult_82_CARRYB_13__39_), .A2(
        u5_mult_82_SUMB_13__40_), .ZN(u5_mult_82_n5354) );
  XNOR2_X2 u5_mult_82_U4821 ( .A(u5_mult_82_CARRYB_7__34_), .B(
        u5_mult_82_ab_8__34_), .ZN(u5_mult_82_n1248) );
  XNOR2_X2 u5_mult_82_U4820 ( .A(u5_mult_82_n1248), .B(u5_mult_82_SUMB_7__35_), 
        .ZN(u5_mult_82_SUMB_8__34_) );
  NAND2_X2 u5_mult_82_U4819 ( .A1(u5_mult_82_CARRYB_39__29_), .A2(
        u5_mult_82_SUMB_39__30_), .ZN(u5_mult_82_n4329) );
  NAND2_X1 u5_mult_82_U4818 ( .A1(u5_mult_82_CARRYB_37__28_), .A2(
        u5_mult_82_SUMB_37__29_), .ZN(u5_mult_82_n5721) );
  NAND2_X1 u5_mult_82_U4817 ( .A1(u5_mult_82_ab_38__28_), .A2(
        u5_mult_82_SUMB_37__29_), .ZN(u5_mult_82_n5720) );
  NAND2_X2 u5_mult_82_U4816 ( .A1(u5_mult_82_ab_21__23_), .A2(
        u5_mult_82_SUMB_20__24_), .ZN(u5_mult_82_n3616) );
  NAND2_X2 u5_mult_82_U4815 ( .A1(u5_mult_82_CARRYB_33__15_), .A2(
        u5_mult_82_SUMB_33__16_), .ZN(u5_mult_82_n6039) );
  NAND2_X1 u5_mult_82_U4814 ( .A1(u5_mult_82_CARRYB_48__7_), .A2(
        u5_mult_82_SUMB_48__8_), .ZN(u5_mult_82_net81830) );
  NAND2_X2 u5_mult_82_U4813 ( .A1(u5_mult_82_ab_32__38_), .A2(
        u5_mult_82_SUMB_31__39_), .ZN(u5_mult_82_n4926) );
  NAND2_X2 u5_mult_82_U4812 ( .A1(u5_mult_82_ab_25__34_), .A2(
        u5_mult_82_CARRYB_24__34_), .ZN(u5_mult_82_n5764) );
  XNOR2_X2 u5_mult_82_U4811 ( .A(u5_mult_82_SUMB_50__24_), .B(
        u5_mult_82_ab_51__23_), .ZN(u5_mult_82_n1247) );
  XNOR2_X2 u5_mult_82_U4810 ( .A(u5_mult_82_ab_7__42_), .B(
        u5_mult_82_CARRYB_6__42_), .ZN(u5_mult_82_n1805) );
  INV_X4 u5_mult_82_U4809 ( .A(u5_mult_82_SUMB_47__8_), .ZN(u5_mult_82_n1340)
         );
  INV_X2 u5_mult_82_U4808 ( .A(u5_mult_82_n1896), .ZN(u5_mult_82_n1761) );
  NAND2_X2 u5_mult_82_U4807 ( .A1(u5_mult_82_n1761), .A2(
        u5_mult_82_SUMB_14__32_), .ZN(u5_mult_82_n5794) );
  NAND3_X2 u5_mult_82_U4806 ( .A1(u5_mult_82_n2891), .A2(u5_mult_82_n2892), 
        .A3(u5_mult_82_n2893), .ZN(u5_mult_82_CARRYB_41__15_) );
  NAND2_X2 u5_mult_82_U4805 ( .A1(u5_mult_82_ab_42__15_), .A2(
        u5_mult_82_CARRYB_41__15_), .ZN(u5_mult_82_n6358) );
  NAND2_X2 u5_mult_82_U4804 ( .A1(u5_mult_82_ab_39__16_), .A2(
        u5_mult_82_CARRYB_38__16_), .ZN(u5_mult_82_n2884) );
  XNOR2_X2 u5_mult_82_U4803 ( .A(u5_mult_82_n2052), .B(u5_mult_82_SUMB_29__23_), .ZN(u5_mult_82_SUMB_30__22_) );
  NAND2_X2 u5_mult_82_U4802 ( .A1(u5_mult_82_CARRYB_44__9_), .A2(
        u5_mult_82_SUMB_44__10_), .ZN(u5_mult_82_net79321) );
  NAND2_X2 u5_mult_82_U4801 ( .A1(u5_mult_82_n82), .A2(u5_mult_82_ab_35__23_), 
        .ZN(u5_mult_82_n6214) );
  NAND2_X1 u5_mult_82_U4800 ( .A1(u5_mult_82_CARRYB_46__14_), .A2(
        u5_mult_82_n1693), .ZN(u5_mult_82_n5772) );
  NAND2_X1 u5_mult_82_U4799 ( .A1(u5_mult_82_ab_47__14_), .A2(u5_mult_82_n1693), .ZN(u5_mult_82_n5771) );
  XNOR2_X2 u5_mult_82_U4798 ( .A(u5_mult_82_n1246), .B(u5_mult_82_SUMB_6__39_), 
        .ZN(u5_mult_82_SUMB_7__38_) );
  XNOR2_X2 u5_mult_82_U4797 ( .A(u5_mult_82_n1245), .B(
        u5_mult_82_CARRYB_10__36_), .ZN(u5_mult_82_n5903) );
  NAND2_X4 u5_mult_82_U4796 ( .A1(u5_mult_82_n3586), .A2(u5_mult_82_n3585), 
        .ZN(u5_mult_82_n5945) );
  NAND3_X2 u5_mult_82_U4795 ( .A1(u5_mult_82_n4935), .A2(u5_mult_82_n4936), 
        .A3(u5_mult_82_n4937), .ZN(u5_mult_82_CARRYB_29__33_) );
  XOR2_X2 u5_mult_82_U4794 ( .A(u5_mult_82_SUMB_31__39_), .B(u5_mult_82_n4924), 
        .Z(u5_mult_82_SUMB_32__38_) );
  INV_X4 u5_mult_82_U4793 ( .A(u5_mult_82_n6419), .ZN(u5_mult_82_CLA_SUM[83])
         );
  NAND2_X2 u5_mult_82_U4792 ( .A1(u5_mult_82_ab_45__9_), .A2(
        u5_mult_82_SUMB_44__10_), .ZN(u5_mult_82_net79320) );
  NAND3_X2 u5_mult_82_U4791 ( .A1(u5_mult_82_n2259), .A2(u5_mult_82_n2258), 
        .A3(u5_mult_82_n2257), .ZN(u5_mult_82_CARRYB_23__37_) );
  NAND2_X2 u5_mult_82_U4790 ( .A1(u5_mult_82_ab_10__45_), .A2(
        u5_mult_82_CARRYB_9__45_), .ZN(u5_mult_82_n4799) );
  NAND2_X2 u5_mult_82_U4789 ( .A1(u5_mult_82_CARRYB_22__37_), .A2(
        u5_mult_82_SUMB_22__38_), .ZN(u5_mult_82_n2259) );
  BUF_X4 u5_mult_82_U4788 ( .A(u5_mult_82_SUMB_19__32_), .Z(u5_mult_82_n1582)
         );
  XNOR2_X2 u5_mult_82_U4787 ( .A(u5_mult_82_CARRYB_36__37_), .B(
        u5_mult_82_ab_37__37_), .ZN(u5_mult_82_n1244) );
  XNOR2_X2 u5_mult_82_U4786 ( .A(u5_mult_82_SUMB_36__38_), .B(u5_mult_82_n1244), .ZN(u5_mult_82_SUMB_37__37_) );
  XNOR2_X2 u5_mult_82_U4785 ( .A(u5_mult_82_CARRYB_19__33_), .B(
        u5_mult_82_ab_20__33_), .ZN(u5_mult_82_n1243) );
  XNOR2_X2 u5_mult_82_U4784 ( .A(u5_mult_82_n1243), .B(u5_mult_82_SUMB_19__34_), .ZN(u5_mult_82_SUMB_20__33_) );
  XNOR2_X2 u5_mult_82_U4783 ( .A(u5_mult_82_CARRYB_39__29_), .B(
        u5_mult_82_ab_40__29_), .ZN(u5_mult_82_n1648) );
  XNOR2_X2 u5_mult_82_U4782 ( .A(u5_mult_82_CARRYB_2__26_), .B(
        u5_mult_82_ab_3__26_), .ZN(u5_mult_82_n1242) );
  XNOR2_X2 u5_mult_82_U4781 ( .A(u5_mult_82_n1242), .B(u5_mult_82_SUMB_2__27_), 
        .ZN(u5_mult_82_SUMB_3__26_) );
  NAND2_X1 u5_mult_82_U4780 ( .A1(u5_mult_82_ab_38__29_), .A2(
        u5_mult_82_SUMB_37__30_), .ZN(u5_mult_82_n5276) );
  NAND2_X2 u5_mult_82_U4779 ( .A1(u5_mult_82_CARRYB_18__27_), .A2(
        u5_mult_82_SUMB_18__28_), .ZN(u5_mult_82_n5802) );
  XNOR2_X2 u5_mult_82_U4778 ( .A(u5_mult_82_ab_35__31_), .B(
        u5_mult_82_CARRYB_34__31_), .ZN(u5_mult_82_n1241) );
  XNOR2_X2 u5_mult_82_U4777 ( .A(u5_mult_82_n1241), .B(u5_mult_82_SUMB_34__32_), .ZN(u5_mult_82_SUMB_35__31_) );
  NAND2_X4 u5_mult_82_U4776 ( .A1(u5_mult_82_n2746), .A2(u5_mult_82_n2747), 
        .ZN(u5_mult_82_SUMB_45__8_) );
  XNOR2_X2 u5_mult_82_U4775 ( .A(u5_mult_82_ab_46__7_), .B(
        u5_mult_82_SUMB_45__8_), .ZN(u5_mult_82_n2136) );
  INV_X4 u5_mult_82_U4774 ( .A(u5_mult_82_n2016), .ZN(u5_mult_82_ab_0__39_) );
  XNOR2_X2 u5_mult_82_U4773 ( .A(u5_mult_82_ab_25__45_), .B(
        u5_mult_82_CARRYB_24__45_), .ZN(u5_mult_82_n1240) );
  XNOR2_X2 u5_mult_82_U4772 ( .A(u5_mult_82_CARRYB_16__28_), .B(
        u5_mult_82_ab_17__28_), .ZN(u5_mult_82_net81335) );
  NOR2_X1 u5_mult_82_U4771 ( .A1(u5_mult_82_n6876), .A2(u5_mult_82_n6650), 
        .ZN(u5_mult_82_ab_26__27_) );
  NAND3_X4 u5_mult_82_U4770 ( .A1(u5_mult_82_n4247), .A2(u5_mult_82_n4246), 
        .A3(u5_mult_82_n4245), .ZN(u5_mult_82_CARRYB_35__21_) );
  NOR2_X2 u5_mult_82_U4769 ( .A1(u5_mult_82_n6896), .A2(u5_mult_82_n6715), 
        .ZN(u5_mult_82_ab_36__21_) );
  NOR2_X2 u5_mult_82_U4768 ( .A1(u5_mult_82_n6896), .A2(u5_mult_82_n6721), 
        .ZN(u5_mult_82_ab_37__21_) );
  NAND2_X1 u5_mult_82_U4767 ( .A1(u5_mult_82_ab_26__27_), .A2(
        u5_mult_82_CARRYB_25__27_), .ZN(u5_mult_82_n1239) );
  NAND2_X2 u5_mult_82_U4766 ( .A1(u5_mult_82_ab_26__27_), .A2(
        u5_mult_82_SUMB_25__28_), .ZN(u5_mult_82_n1238) );
  NAND2_X1 u5_mult_82_U4765 ( .A1(u5_mult_82_CARRYB_25__27_), .A2(
        u5_mult_82_SUMB_25__28_), .ZN(u5_mult_82_n1237) );
  XOR2_X2 u5_mult_82_U4764 ( .A(u5_mult_82_n1236), .B(u5_mult_82_SUMB_25__28_), 
        .Z(u5_mult_82_SUMB_26__27_) );
  NAND3_X4 u5_mult_82_U4763 ( .A1(u5_mult_82_n1233), .A2(u5_mult_82_n1234), 
        .A3(u5_mult_82_n1235), .ZN(u5_mult_82_CARRYB_36__21_) );
  NAND2_X1 u5_mult_82_U4762 ( .A1(u5_mult_82_ab_36__21_), .A2(
        u5_mult_82_CARRYB_35__21_), .ZN(u5_mult_82_n1235) );
  NAND2_X2 u5_mult_82_U4761 ( .A1(u5_mult_82_ab_36__21_), .A2(
        u5_mult_82_SUMB_35__22_), .ZN(u5_mult_82_n1234) );
  NAND2_X2 u5_mult_82_U4760 ( .A1(u5_mult_82_CARRYB_35__21_), .A2(
        u5_mult_82_SUMB_35__22_), .ZN(u5_mult_82_n1233) );
  XOR2_X2 u5_mult_82_U4759 ( .A(u5_mult_82_SUMB_35__22_), .B(u5_mult_82_n1232), 
        .Z(u5_mult_82_SUMB_36__21_) );
  XOR2_X2 u5_mult_82_U4758 ( .A(u5_mult_82_CARRYB_35__21_), .B(
        u5_mult_82_ab_36__21_), .Z(u5_mult_82_n1232) );
  NAND3_X2 u5_mult_82_U4757 ( .A1(u5_mult_82_n1229), .A2(u5_mult_82_n1230), 
        .A3(u5_mult_82_n1231), .ZN(u5_mult_82_CARRYB_37__21_) );
  NAND2_X2 u5_mult_82_U4756 ( .A1(u5_mult_82_ab_37__21_), .A2(
        u5_mult_82_SUMB_36__22_), .ZN(u5_mult_82_n1231) );
  NAND2_X2 u5_mult_82_U4755 ( .A1(u5_mult_82_ab_37__21_), .A2(
        u5_mult_82_CARRYB_36__21_), .ZN(u5_mult_82_n1230) );
  NAND2_X1 u5_mult_82_U4754 ( .A1(u5_mult_82_SUMB_36__22_), .A2(
        u5_mult_82_CARRYB_36__21_), .ZN(u5_mult_82_n1229) );
  INV_X1 u5_mult_82_U4753 ( .A(u5_mult_82_n1384), .ZN(u5_mult_82_n1226) );
  NAND2_X2 u5_mult_82_U4752 ( .A1(u5_mult_82_n1225), .A2(u5_mult_82_n1226), 
        .ZN(u5_mult_82_n1228) );
  NAND2_X1 u5_mult_82_U4751 ( .A1(u5_mult_82_n1603), .A2(u5_mult_82_n1384), 
        .ZN(u5_mult_82_n1227) );
  NAND3_X4 u5_mult_82_U4750 ( .A1(u5_mult_82_n1297), .A2(u5_mult_82_net79320), 
        .A3(u5_mult_82_net79321), .ZN(u5_mult_82_CARRYB_45__9_) );
  NAND2_X1 u5_mult_82_U4749 ( .A1(u5_mult_82_ab_23__38_), .A2(
        u5_mult_82_SUMB_22__39_), .ZN(u5_mult_82_n6001) );
  NAND2_X4 u5_mult_82_U4748 ( .A1(u5_mult_82_CARRYB_15__36_), .A2(
        u5_mult_82_n1827), .ZN(u5_mult_82_n6189) );
  CLKBUF_X3 u5_mult_82_U4747 ( .A(u5_mult_82_CARRYB_40__26_), .Z(
        u5_mult_82_n1450) );
  NAND3_X4 u5_mult_82_U4746 ( .A1(u5_mult_82_n5558), .A2(u5_mult_82_n5559), 
        .A3(u5_mult_82_n5560), .ZN(u5_mult_82_CARRYB_24__37_) );
  NAND2_X2 u5_mult_82_U4745 ( .A1(u5_mult_82_ab_25__24_), .A2(
        u5_mult_82_CARRYB_24__24_), .ZN(u5_mult_82_n6055) );
  NOR2_X1 u5_mult_82_U4744 ( .A1(u5_mult_82_n6892), .A2(u5_mult_82_n6643), 
        .ZN(u5_mult_82_ab_24__24_) );
  NAND2_X2 u5_mult_82_U4743 ( .A1(u5_mult_82_ab_34__20_), .A2(
        u5_mult_82_CARRYB_33__20_), .ZN(u5_mult_82_n6333) );
  NOR2_X1 u5_mult_82_U4742 ( .A1(u5_mult_82_n6904), .A2(u5_mult_82_n6700), 
        .ZN(u5_mult_82_ab_33__20_) );
  NAND3_X2 u5_mult_82_U4741 ( .A1(u5_mult_82_n1222), .A2(u5_mult_82_n1223), 
        .A3(u5_mult_82_n1224), .ZN(u5_mult_82_CARRYB_13__31_) );
  NAND2_X1 u5_mult_82_U4740 ( .A1(u5_mult_82_CARRYB_12__31_), .A2(
        u5_mult_82_SUMB_12__32_), .ZN(u5_mult_82_n1224) );
  NAND2_X1 u5_mult_82_U4739 ( .A1(u5_mult_82_ab_13__31_), .A2(
        u5_mult_82_SUMB_12__32_), .ZN(u5_mult_82_n1223) );
  NAND2_X1 u5_mult_82_U4738 ( .A1(u5_mult_82_ab_13__31_), .A2(
        u5_mult_82_CARRYB_12__31_), .ZN(u5_mult_82_n1222) );
  NAND3_X4 u5_mult_82_U4737 ( .A1(u5_mult_82_n1219), .A2(u5_mult_82_n1220), 
        .A3(u5_mult_82_n1221), .ZN(u5_mult_82_CARRYB_12__32_) );
  NAND2_X2 u5_mult_82_U4736 ( .A1(u5_mult_82_CARRYB_11__32_), .A2(
        u5_mult_82_SUMB_11__33_), .ZN(u5_mult_82_n1221) );
  NAND2_X2 u5_mult_82_U4735 ( .A1(u5_mult_82_ab_12__32_), .A2(
        u5_mult_82_SUMB_11__33_), .ZN(u5_mult_82_n1220) );
  NAND2_X1 u5_mult_82_U4734 ( .A1(u5_mult_82_ab_12__32_), .A2(
        u5_mult_82_CARRYB_11__32_), .ZN(u5_mult_82_n1219) );
  NAND3_X2 u5_mult_82_U4733 ( .A1(u5_mult_82_n1216), .A2(u5_mult_82_n1217), 
        .A3(u5_mult_82_n1218), .ZN(u5_mult_82_CARRYB_24__24_) );
  NAND2_X1 u5_mult_82_U4732 ( .A1(u5_mult_82_ab_24__24_), .A2(
        u5_mult_82_CARRYB_23__24_), .ZN(u5_mult_82_n1218) );
  NAND2_X2 u5_mult_82_U4731 ( .A1(u5_mult_82_ab_24__24_), .A2(
        u5_mult_82_SUMB_23__25_), .ZN(u5_mult_82_n1217) );
  NAND2_X1 u5_mult_82_U4730 ( .A1(u5_mult_82_CARRYB_23__24_), .A2(
        u5_mult_82_SUMB_23__25_), .ZN(u5_mult_82_n1216) );
  XOR2_X2 u5_mult_82_U4729 ( .A(u5_mult_82_SUMB_23__25_), .B(u5_mult_82_n1215), 
        .Z(u5_mult_82_SUMB_24__24_) );
  NAND3_X2 u5_mult_82_U4728 ( .A1(u5_mult_82_n1212), .A2(u5_mult_82_n1213), 
        .A3(u5_mult_82_n1214), .ZN(u5_mult_82_CARRYB_33__20_) );
  NAND2_X1 u5_mult_82_U4727 ( .A1(u5_mult_82_ab_33__20_), .A2(
        u5_mult_82_CARRYB_32__20_), .ZN(u5_mult_82_n1214) );
  NAND2_X2 u5_mult_82_U4726 ( .A1(u5_mult_82_ab_33__20_), .A2(
        u5_mult_82_SUMB_32__21_), .ZN(u5_mult_82_n1213) );
  XOR2_X2 u5_mult_82_U4725 ( .A(u5_mult_82_SUMB_32__21_), .B(u5_mult_82_n1211), 
        .Z(u5_mult_82_SUMB_33__20_) );
  XOR2_X2 u5_mult_82_U4724 ( .A(u5_mult_82_CARRYB_32__20_), .B(
        u5_mult_82_ab_33__20_), .Z(u5_mult_82_n1211) );
  NAND2_X2 u5_mult_82_U4723 ( .A1(u5_mult_82_ab_3__46_), .A2(
        u5_mult_82_CARRYB_2__46_), .ZN(u5_mult_82_n1932) );
  NOR2_X2 u5_mult_82_U4722 ( .A1(u5_mult_82_n6794), .A2(u5_mult_82_net66087), 
        .ZN(u5_mult_82_ab_2__46_) );
  NOR2_X4 u5_mult_82_U4721 ( .A1(u5_mult_82_n6862), .A2(u5_mult_82_n6707), 
        .ZN(u5_mult_82_ab_35__29_) );
  NAND3_X4 u5_mult_82_U4720 ( .A1(u5_mult_82_n1208), .A2(u5_mult_82_n1209), 
        .A3(u5_mult_82_n1210), .ZN(u5_mult_82_CARRYB_2__46_) );
  NAND2_X2 u5_mult_82_U4719 ( .A1(u5_mult_82_ab_2__46_), .A2(
        u5_mult_82_CARRYB_1__46_), .ZN(u5_mult_82_n1210) );
  XOR2_X2 u5_mult_82_U4718 ( .A(u5_mult_82_SUMB_1__47_), .B(u5_mult_82_n1207), 
        .Z(u5_mult_82_SUMB_2__46_) );
  INV_X1 u5_mult_82_U4717 ( .A(u5_mult_82_ab_35__29_), .ZN(u5_mult_82_n1204)
         );
  NAND2_X2 u5_mult_82_U4716 ( .A1(u5_mult_82_n640), .A2(u5_mult_82_n1204), 
        .ZN(u5_mult_82_n1206) );
  XNOR2_X2 u5_mult_82_U4715 ( .A(u5_mult_82_CARRYB_12__36_), .B(
        u5_mult_82_n1203), .ZN(u5_mult_82_n5197) );
  NAND2_X2 u5_mult_82_U4714 ( .A1(u5_mult_82_ab_22__39_), .A2(
        u5_mult_82_CARRYB_21__39_), .ZN(u5_mult_82_n5997) );
  NAND3_X2 u5_mult_82_U4713 ( .A1(u5_mult_82_n5101), .A2(u5_mult_82_n5102), 
        .A3(u5_mult_82_n5103), .ZN(u5_mult_82_CARRYB_51__21_) );
  NAND2_X2 u5_mult_82_U4712 ( .A1(u5_mult_82_CARRYB_28__16_), .A2(
        u5_mult_82_SUMB_28__17_), .ZN(u5_mult_82_n3652) );
  NAND3_X2 u5_mult_82_U4711 ( .A1(u5_mult_82_n3244), .A2(u5_mult_82_n3245), 
        .A3(u5_mult_82_n3246), .ZN(u5_mult_82_CARRYB_19__22_) );
  XNOR2_X2 u5_mult_82_U4710 ( .A(u5_mult_82_ab_27__18_), .B(
        u5_mult_82_CARRYB_26__18_), .ZN(u5_mult_82_n2751) );
  NAND2_X2 u5_mult_82_U4709 ( .A1(u5_mult_82_CARRYB_14__48_), .A2(
        u5_mult_82_SUMB_14__49_), .ZN(u5_mult_82_n4328) );
  NAND2_X2 u5_mult_82_U4708 ( .A1(u5_mult_82_CARRYB_23__42_), .A2(
        u5_mult_82_SUMB_23__43_), .ZN(u5_mult_82_n3076) );
  NAND2_X4 u5_mult_82_U4707 ( .A1(u5_mult_82_CARRYB_43__0_), .A2(
        u5_mult_82_ab_44__0_), .ZN(u5_mult_82_n4843) );
  NAND2_X2 u5_mult_82_U4706 ( .A1(u5_mult_82_ab_14__49_), .A2(
        u5_mult_82_CARRYB_13__49_), .ZN(u5_mult_82_n4323) );
  XNOR2_X1 u5_mult_82_U4705 ( .A(u5_mult_82_n2138), .B(
        u5_mult_82_CARRYB_11__50_), .ZN(u5_mult_82_SUMB_12__50_) );
  NOR2_X2 u5_mult_82_U4704 ( .A1(u5_mult_82_n6775), .A2(u5_mult_82_n6572), 
        .ZN(u5_mult_82_ab_13__49_) );
  NOR2_X2 u5_mult_82_U4703 ( .A1(u5_mult_82_n6774), .A2(u5_mult_82_n6607), 
        .ZN(u5_mult_82_ab_18__49_) );
  NOR2_X1 u5_mult_82_U4702 ( .A1(u5_mult_82_n6791), .A2(u5_mult_82_n6720), 
        .ZN(u5_mult_82_ab_37__46_) );
  NAND3_X2 u5_mult_82_U4701 ( .A1(u5_mult_82_n1200), .A2(u5_mult_82_n1201), 
        .A3(u5_mult_82_n1202), .ZN(u5_mult_82_CARRYB_13__49_) );
  NAND2_X1 u5_mult_82_U4700 ( .A1(u5_mult_82_ab_13__49_), .A2(
        u5_mult_82_SUMB_12__50_), .ZN(u5_mult_82_n1202) );
  XOR2_X2 u5_mult_82_U4699 ( .A(u5_mult_82_CARRYB_12__49_), .B(
        u5_mult_82_n1199), .Z(u5_mult_82_SUMB_13__49_) );
  XOR2_X2 u5_mult_82_U4698 ( .A(u5_mult_82_SUMB_12__50_), .B(
        u5_mult_82_ab_13__49_), .Z(u5_mult_82_n1199) );
  NAND3_X4 u5_mult_82_U4697 ( .A1(u5_mult_82_n1196), .A2(u5_mult_82_n1197), 
        .A3(u5_mult_82_n1198), .ZN(u5_mult_82_CARRYB_18__49_) );
  NAND2_X2 u5_mult_82_U4696 ( .A1(u5_mult_82_ab_18__49_), .A2(
        u5_mult_82_CARRYB_17__49_), .ZN(u5_mult_82_n1197) );
  XOR2_X2 u5_mult_82_U4695 ( .A(u5_mult_82_CARRYB_17__49_), .B(
        u5_mult_82_n1195), .Z(u5_mult_82_SUMB_18__49_) );
  XOR2_X2 u5_mult_82_U4694 ( .A(u5_mult_82_SUMB_17__50_), .B(
        u5_mult_82_ab_18__49_), .Z(u5_mult_82_n1195) );
  NAND3_X2 u5_mult_82_U4693 ( .A1(u5_mult_82_n1192), .A2(u5_mult_82_n1193), 
        .A3(u5_mult_82_n1194), .ZN(u5_mult_82_CARRYB_20__49_) );
  NAND2_X1 u5_mult_82_U4692 ( .A1(u5_mult_82_SUMB_19__50_), .A2(
        u5_mult_82_CARRYB_19__49_), .ZN(u5_mult_82_n1194) );
  NAND2_X1 u5_mult_82_U4691 ( .A1(u5_mult_82_ab_20__49_), .A2(
        u5_mult_82_CARRYB_19__49_), .ZN(u5_mult_82_n1193) );
  NAND2_X1 u5_mult_82_U4690 ( .A1(u5_mult_82_ab_20__49_), .A2(
        u5_mult_82_SUMB_19__50_), .ZN(u5_mult_82_n1192) );
  XOR2_X2 u5_mult_82_U4689 ( .A(u5_mult_82_n1191), .B(
        u5_mult_82_CARRYB_19__49_), .Z(u5_mult_82_SUMB_20__49_) );
  XOR2_X2 u5_mult_82_U4688 ( .A(u5_mult_82_ab_20__49_), .B(
        u5_mult_82_SUMB_19__50_), .Z(u5_mult_82_n1191) );
  NAND3_X2 u5_mult_82_U4687 ( .A1(u5_mult_82_n1188), .A2(u5_mult_82_n1189), 
        .A3(u5_mult_82_n1190), .ZN(u5_mult_82_CARRYB_19__49_) );
  NAND2_X2 u5_mult_82_U4686 ( .A1(u5_mult_82_CARRYB_18__49_), .A2(
        u5_mult_82_SUMB_18__50_), .ZN(u5_mult_82_n1190) );
  NAND2_X2 u5_mult_82_U4685 ( .A1(u5_mult_82_ab_19__49_), .A2(
        u5_mult_82_SUMB_18__50_), .ZN(u5_mult_82_n1189) );
  NAND2_X2 u5_mult_82_U4684 ( .A1(u5_mult_82_ab_19__49_), .A2(
        u5_mult_82_CARRYB_18__49_), .ZN(u5_mult_82_n1188) );
  XOR2_X2 u5_mult_82_U4683 ( .A(u5_mult_82_n1187), .B(u5_mult_82_SUMB_18__50_), 
        .Z(u5_mult_82_SUMB_19__49_) );
  XOR2_X2 u5_mult_82_U4682 ( .A(u5_mult_82_ab_19__49_), .B(
        u5_mult_82_CARRYB_18__49_), .Z(u5_mult_82_n1187) );
  NAND3_X2 u5_mult_82_U4681 ( .A1(u5_mult_82_n1184), .A2(u5_mult_82_n1185), 
        .A3(u5_mult_82_n1186), .ZN(u5_mult_82_CARRYB_37__46_) );
  NAND2_X1 u5_mult_82_U4680 ( .A1(u5_mult_82_ab_37__46_), .A2(
        u5_mult_82_CARRYB_36__46_), .ZN(u5_mult_82_n1186) );
  NAND2_X1 u5_mult_82_U4679 ( .A1(u5_mult_82_ab_37__46_), .A2(
        u5_mult_82_SUMB_36__47_), .ZN(u5_mult_82_n1185) );
  NAND2_X1 u5_mult_82_U4678 ( .A1(u5_mult_82_CARRYB_36__46_), .A2(
        u5_mult_82_SUMB_36__47_), .ZN(u5_mult_82_n1184) );
  XOR2_X2 u5_mult_82_U4677 ( .A(u5_mult_82_SUMB_36__47_), .B(u5_mult_82_n1183), 
        .Z(u5_mult_82_SUMB_37__46_) );
  XOR2_X2 u5_mult_82_U4676 ( .A(u5_mult_82_CARRYB_36__46_), .B(
        u5_mult_82_ab_37__46_), .Z(u5_mult_82_n1183) );
  XNOR2_X2 u5_mult_82_U4675 ( .A(u5_mult_82_n5762), .B(u5_mult_82_n1817), .ZN(
        u5_mult_82_SUMB_25__34_) );
  NAND2_X2 u5_mult_82_U4674 ( .A1(u5_mult_82_ab_38__21_), .A2(
        u5_mult_82_SUMB_37__22_), .ZN(u5_mult_82_n4003) );
  NAND2_X2 u5_mult_82_U4673 ( .A1(u5_mult_82_CARRYB_31__24_), .A2(
        u5_mult_82_SUMB_31__25_), .ZN(u5_mult_82_n4241) );
  XNOR2_X2 u5_mult_82_U4672 ( .A(u5_mult_82_n1410), .B(u5_mult_82_SUMB_22__38_), .ZN(u5_mult_82_SUMB_23__37_) );
  NAND2_X2 u5_mult_82_U4671 ( .A1(u5_mult_82_ab_34__32_), .A2(u5_mult_82_n74), 
        .ZN(u5_mult_82_n2718) );
  XNOR2_X2 u5_mult_82_U4670 ( .A(u5_mult_82_ab_22__39_), .B(
        u5_mult_82_CARRYB_21__39_), .ZN(u5_mult_82_n1723) );
  INV_X4 u5_mult_82_U4669 ( .A(n4791), .ZN(u5_mult_82_net64959) );
  INV_X4 u5_mult_82_U4668 ( .A(n4791), .ZN(u5_mult_82_net64957) );
  CLKBUF_X3 u5_mult_82_U4667 ( .A(u5_mult_82_CARRYB_23__23_), .Z(
        u5_mult_82_net88030) );
  NAND2_X2 u5_mult_82_U4666 ( .A1(u5_mult_82_ab_51__7_), .A2(
        u5_mult_82_CARRYB_50__7_), .ZN(u5_mult_82_n6202) );
  NAND2_X2 u5_mult_82_U4665 ( .A1(u5_mult_82_n3605), .A2(
        u5_mult_82_CARRYB_32__31_), .ZN(u5_mult_82_n3585) );
  BUF_X8 u5_mult_82_U4664 ( .A(u5_mult_82_n49), .Z(u5_mult_82_n1484) );
  NAND2_X1 u5_mult_82_U4663 ( .A1(u5_mult_82_CARRYB_45__27_), .A2(
        u5_mult_82_SUMB_45__28_), .ZN(u5_mult_82_n4575) );
  NOR2_X1 u5_mult_82_U4662 ( .A1(u5_mult_82_net64453), .A2(u5_mult_82_n6603), 
        .ZN(u5_mult_82_ab_17__10_) );
  NAND2_X2 u5_mult_82_U4661 ( .A1(u5_mult_82_ab_5__22_), .A2(
        u5_mult_82_CARRYB_4__22_), .ZN(u5_mult_82_n1958) );
  NAND2_X2 u5_mult_82_U4660 ( .A1(u5_mult_82_CARRYB_4__22_), .A2(
        u5_mult_82_SUMB_4__23_), .ZN(u5_mult_82_n1960) );
  NOR2_X2 u5_mult_82_U4659 ( .A1(u5_mult_82_net64671), .A2(u5_mult_82_n6522), 
        .ZN(u5_mult_82_ab_4__22_) );
  NAND2_X2 u5_mult_82_U4658 ( .A1(u5_mult_82_ab_8__19_), .A2(
        u5_mult_82_CARRYB_7__19_), .ZN(u5_mult_82_n2761) );
  NOR2_X2 u5_mult_82_U4657 ( .A1(u5_mult_82_n6915), .A2(u5_mult_82_n6529), 
        .ZN(u5_mult_82_ab_7__19_) );
  NAND3_X2 u5_mult_82_U4656 ( .A1(u5_mult_82_n1180), .A2(u5_mult_82_n1181), 
        .A3(u5_mult_82_n1182), .ZN(u5_mult_82_CARRYB_17__10_) );
  NAND2_X1 u5_mult_82_U4655 ( .A1(u5_mult_82_ab_17__10_), .A2(
        u5_mult_82_CARRYB_16__10_), .ZN(u5_mult_82_n1182) );
  NAND2_X2 u5_mult_82_U4654 ( .A1(u5_mult_82_ab_17__10_), .A2(
        u5_mult_82_SUMB_16__11_), .ZN(u5_mult_82_n1181) );
  NAND2_X1 u5_mult_82_U4653 ( .A1(u5_mult_82_CARRYB_16__10_), .A2(
        u5_mult_82_SUMB_16__11_), .ZN(u5_mult_82_n1180) );
  XOR2_X2 u5_mult_82_U4652 ( .A(u5_mult_82_SUMB_16__11_), .B(u5_mult_82_n1179), 
        .Z(u5_mult_82_SUMB_17__10_) );
  XOR2_X2 u5_mult_82_U4651 ( .A(u5_mult_82_CARRYB_16__10_), .B(
        u5_mult_82_ab_17__10_), .Z(u5_mult_82_n1179) );
  NAND3_X2 u5_mult_82_U4650 ( .A1(u5_mult_82_n1176), .A2(u5_mult_82_n1177), 
        .A3(u5_mult_82_n1178), .ZN(u5_mult_82_CARRYB_6__20_) );
  NAND2_X1 u5_mult_82_U4649 ( .A1(u5_mult_82_CARRYB_5__20_), .A2(
        u5_mult_82_SUMB_5__21_), .ZN(u5_mult_82_n1178) );
  NAND2_X1 u5_mult_82_U4648 ( .A1(u5_mult_82_ab_6__20_), .A2(
        u5_mult_82_SUMB_5__21_), .ZN(u5_mult_82_n1177) );
  NAND2_X1 u5_mult_82_U4647 ( .A1(u5_mult_82_ab_6__20_), .A2(
        u5_mult_82_CARRYB_5__20_), .ZN(u5_mult_82_n1176) );
  NAND3_X2 u5_mult_82_U4646 ( .A1(u5_mult_82_n1173), .A2(u5_mult_82_n1174), 
        .A3(u5_mult_82_n1175), .ZN(u5_mult_82_CARRYB_5__21_) );
  NAND2_X1 u5_mult_82_U4645 ( .A1(u5_mult_82_CARRYB_4__21_), .A2(
        u5_mult_82_SUMB_4__22_), .ZN(u5_mult_82_n1175) );
  NAND2_X1 u5_mult_82_U4644 ( .A1(u5_mult_82_ab_5__21_), .A2(
        u5_mult_82_SUMB_4__22_), .ZN(u5_mult_82_n1174) );
  NAND2_X1 u5_mult_82_U4643 ( .A1(u5_mult_82_ab_5__21_), .A2(
        u5_mult_82_CARRYB_4__21_), .ZN(u5_mult_82_n1173) );
  XOR2_X2 u5_mult_82_U4642 ( .A(u5_mult_82_n1172), .B(u5_mult_82_SUMB_5__21_), 
        .Z(u5_mult_82_SUMB_6__20_) );
  XOR2_X2 u5_mult_82_U4641 ( .A(u5_mult_82_ab_6__20_), .B(
        u5_mult_82_CARRYB_5__20_), .Z(u5_mult_82_n1172) );
  XOR2_X2 u5_mult_82_U4640 ( .A(u5_mult_82_n1171), .B(u5_mult_82_SUMB_4__22_), 
        .Z(u5_mult_82_SUMB_5__21_) );
  XOR2_X2 u5_mult_82_U4639 ( .A(u5_mult_82_ab_5__21_), .B(
        u5_mult_82_CARRYB_4__21_), .Z(u5_mult_82_n1171) );
  NAND2_X1 u5_mult_82_U4638 ( .A1(u5_mult_82_ab_4__22_), .A2(
        u5_mult_82_CARRYB_3__22_), .ZN(u5_mult_82_n1170) );
  NAND2_X2 u5_mult_82_U4637 ( .A1(u5_mult_82_ab_4__22_), .A2(
        u5_mult_82_SUMB_3__23_), .ZN(u5_mult_82_n1169) );
  NAND2_X2 u5_mult_82_U4636 ( .A1(u5_mult_82_CARRYB_3__22_), .A2(
        u5_mult_82_SUMB_3__23_), .ZN(u5_mult_82_n1168) );
  XOR2_X2 u5_mult_82_U4635 ( .A(u5_mult_82_SUMB_3__23_), .B(u5_mult_82_n1167), 
        .Z(u5_mult_82_SUMB_4__22_) );
  XOR2_X2 u5_mult_82_U4634 ( .A(u5_mult_82_CARRYB_3__22_), .B(
        u5_mult_82_ab_4__22_), .Z(u5_mult_82_n1167) );
  NAND3_X2 u5_mult_82_U4633 ( .A1(u5_mult_82_n1164), .A2(u5_mult_82_n1165), 
        .A3(u5_mult_82_n1166), .ZN(u5_mult_82_CARRYB_7__19_) );
  NAND2_X1 u5_mult_82_U4632 ( .A1(u5_mult_82_ab_7__19_), .A2(
        u5_mult_82_CARRYB_6__19_), .ZN(u5_mult_82_n1166) );
  NAND2_X1 u5_mult_82_U4631 ( .A1(u5_mult_82_ab_7__19_), .A2(
        u5_mult_82_SUMB_6__20_), .ZN(u5_mult_82_n1165) );
  NAND2_X1 u5_mult_82_U4630 ( .A1(u5_mult_82_CARRYB_6__19_), .A2(
        u5_mult_82_SUMB_6__20_), .ZN(u5_mult_82_n1164) );
  XOR2_X2 u5_mult_82_U4629 ( .A(u5_mult_82_SUMB_6__20_), .B(u5_mult_82_n1163), 
        .Z(u5_mult_82_SUMB_7__19_) );
  XOR2_X2 u5_mult_82_U4628 ( .A(u5_mult_82_CARRYB_6__19_), .B(
        u5_mult_82_ab_7__19_), .Z(u5_mult_82_n1163) );
  NAND2_X2 u5_mult_82_U4627 ( .A1(u5_mult_82_ab_30__29_), .A2(
        u5_mult_82_CARRYB_29__29_), .ZN(u5_mult_82_n4537) );
  NAND2_X2 u5_mult_82_U4626 ( .A1(u5_mult_82_SUMB_22__32_), .A2(
        u5_mult_82_CARRYB_22__31_), .ZN(u5_mult_82_n6344) );
  NAND2_X1 u5_mult_82_U4625 ( .A1(u5_mult_82_CARRYB_26__29_), .A2(
        u5_mult_82_SUMB_26__30_), .ZN(u5_mult_82_n6284) );
  NAND2_X2 u5_mult_82_U4624 ( .A1(u5_mult_82_CARRYB_34__23_), .A2(
        u5_mult_82_n82), .ZN(u5_mult_82_n6215) );
  NOR2_X2 u5_mult_82_U4623 ( .A1(u5_mult_82_net64939), .A2(u5_mult_82_n6649), 
        .ZN(u5_mult_82_ab_26__37_) );
  NAND3_X2 u5_mult_82_U4622 ( .A1(u5_mult_82_n1160), .A2(u5_mult_82_n1161), 
        .A3(u5_mult_82_n1162), .ZN(u5_mult_82_CARRYB_26__37_) );
  NAND2_X1 u5_mult_82_U4621 ( .A1(u5_mult_82_ab_26__37_), .A2(
        u5_mult_82_CARRYB_25__37_), .ZN(u5_mult_82_n1162) );
  NAND2_X1 u5_mult_82_U4620 ( .A1(u5_mult_82_ab_26__37_), .A2(
        u5_mult_82_SUMB_25__38_), .ZN(u5_mult_82_n1161) );
  NAND2_X1 u5_mult_82_U4619 ( .A1(u5_mult_82_CARRYB_25__37_), .A2(
        u5_mult_82_SUMB_25__38_), .ZN(u5_mult_82_n1160) );
  XOR2_X2 u5_mult_82_U4618 ( .A(u5_mult_82_SUMB_25__38_), .B(u5_mult_82_n1159), 
        .Z(u5_mult_82_SUMB_26__37_) );
  XOR2_X2 u5_mult_82_U4617 ( .A(u5_mult_82_CARRYB_25__37_), .B(
        u5_mult_82_ab_26__37_), .Z(u5_mult_82_n1159) );
  NAND3_X4 u5_mult_82_U4616 ( .A1(u5_mult_82_n1156), .A2(u5_mult_82_n1157), 
        .A3(u5_mult_82_n1158), .ZN(u5_mult_82_CARRYB_23__39_) );
  NAND2_X2 u5_mult_82_U4615 ( .A1(u5_mult_82_CARRYB_22__39_), .A2(
        u5_mult_82_SUMB_22__40_), .ZN(u5_mult_82_n1158) );
  NAND2_X2 u5_mult_82_U4614 ( .A1(u5_mult_82_ab_23__39_), .A2(
        u5_mult_82_SUMB_22__40_), .ZN(u5_mult_82_n1157) );
  NAND2_X1 u5_mult_82_U4613 ( .A1(u5_mult_82_ab_23__39_), .A2(
        u5_mult_82_CARRYB_22__39_), .ZN(u5_mult_82_n1156) );
  NAND3_X4 u5_mult_82_U4612 ( .A1(u5_mult_82_n1153), .A2(u5_mult_82_n1154), 
        .A3(u5_mult_82_n1155), .ZN(u5_mult_82_CARRYB_22__40_) );
  NAND2_X2 u5_mult_82_U4611 ( .A1(u5_mult_82_CARRYB_21__40_), .A2(
        u5_mult_82_SUMB_21__41_), .ZN(u5_mult_82_n1155) );
  NAND2_X2 u5_mult_82_U4610 ( .A1(u5_mult_82_ab_22__40_), .A2(
        u5_mult_82_SUMB_21__41_), .ZN(u5_mult_82_n1154) );
  NAND2_X1 u5_mult_82_U4609 ( .A1(u5_mult_82_ab_22__40_), .A2(
        u5_mult_82_CARRYB_21__40_), .ZN(u5_mult_82_n1153) );
  XOR2_X2 u5_mult_82_U4608 ( .A(u5_mult_82_n1152), .B(u5_mult_82_SUMB_22__40_), 
        .Z(u5_mult_82_SUMB_23__39_) );
  XOR2_X2 u5_mult_82_U4607 ( .A(u5_mult_82_ab_23__39_), .B(
        u5_mult_82_CARRYB_22__39_), .Z(u5_mult_82_n1152) );
  XOR2_X2 u5_mult_82_U4606 ( .A(u5_mult_82_n1151), .B(u5_mult_82_SUMB_21__41_), 
        .Z(u5_mult_82_SUMB_22__40_) );
  XOR2_X2 u5_mult_82_U4605 ( .A(u5_mult_82_ab_22__40_), .B(
        u5_mult_82_CARRYB_21__40_), .Z(u5_mult_82_n1151) );
  NAND3_X2 u5_mult_82_U4604 ( .A1(u5_mult_82_n1148), .A2(u5_mult_82_n1149), 
        .A3(u5_mult_82_n1150), .ZN(u5_mult_82_CARRYB_46__25_) );
  NAND2_X1 u5_mult_82_U4603 ( .A1(u5_mult_82_CARRYB_45__25_), .A2(
        u5_mult_82_SUMB_45__26_), .ZN(u5_mult_82_n1150) );
  NAND2_X1 u5_mult_82_U4602 ( .A1(u5_mult_82_ab_46__25_), .A2(
        u5_mult_82_SUMB_45__26_), .ZN(u5_mult_82_n1149) );
  NAND2_X1 u5_mult_82_U4601 ( .A1(u5_mult_82_ab_46__25_), .A2(
        u5_mult_82_CARRYB_45__25_), .ZN(u5_mult_82_n1148) );
  NAND3_X2 u5_mult_82_U4600 ( .A1(u5_mult_82_n1145), .A2(u5_mult_82_n1146), 
        .A3(u5_mult_82_n1147), .ZN(u5_mult_82_CARRYB_45__26_) );
  NAND2_X2 u5_mult_82_U4599 ( .A1(u5_mult_82_CARRYB_44__26_), .A2(
        u5_mult_82_SUMB_44__27_), .ZN(u5_mult_82_n1147) );
  NAND2_X2 u5_mult_82_U4598 ( .A1(u5_mult_82_ab_45__26_), .A2(
        u5_mult_82_SUMB_44__27_), .ZN(u5_mult_82_n1146) );
  NAND2_X1 u5_mult_82_U4597 ( .A1(u5_mult_82_ab_45__26_), .A2(
        u5_mult_82_CARRYB_44__26_), .ZN(u5_mult_82_n1145) );
  XOR2_X2 u5_mult_82_U4596 ( .A(u5_mult_82_n1144), .B(u5_mult_82_SUMB_45__26_), 
        .Z(u5_mult_82_SUMB_46__25_) );
  NAND2_X2 u5_mult_82_U4595 ( .A1(u5_mult_82_SUMB_19__44_), .A2(
        u5_mult_82_CARRYB_19__43_), .ZN(u5_mult_82_n4604) );
  NAND2_X2 u5_mult_82_U4594 ( .A1(u5_mult_82_CARRYB_29__15_), .A2(
        u5_mult_82_SUMB_29__16_), .ZN(u5_mult_82_n3658) );
  NAND3_X2 u5_mult_82_U4593 ( .A1(u5_mult_82_n3385), .A2(u5_mult_82_n3386), 
        .A3(u5_mult_82_n3387), .ZN(u5_mult_82_CARRYB_33__26_) );
  NAND2_X2 u5_mult_82_U4592 ( .A1(u5_mult_82_ab_12__47_), .A2(
        u5_mult_82_CARRYB_11__47_), .ZN(u5_mult_82_n4589) );
  NAND2_X2 u5_mult_82_U4591 ( .A1(u5_mult_82_ab_44__18_), .A2(
        u5_mult_82_SUMB_43__19_), .ZN(u5_mult_82_n5838) );
  NAND2_X2 u5_mult_82_U4590 ( .A1(u5_mult_82_CARRYB_43__18_), .A2(
        u5_mult_82_SUMB_43__19_), .ZN(u5_mult_82_n5839) );
  NAND3_X2 u5_mult_82_U4589 ( .A1(u5_mult_82_n3932), .A2(u5_mult_82_n3933), 
        .A3(u5_mult_82_n3934), .ZN(u5_mult_82_CARRYB_38__35_) );
  NAND2_X2 u5_mult_82_U4588 ( .A1(u5_mult_82_CARRYB_11__47_), .A2(
        u5_mult_82_SUMB_11__48_), .ZN(u5_mult_82_n4591) );
  XOR2_X2 u5_mult_82_U4587 ( .A(u5_mult_82_n2595), .B(
        u5_mult_82_CARRYB_46__17_), .Z(u5_mult_82_n1143) );
  XNOR2_X2 u5_mult_82_U4586 ( .A(u5_mult_82_n1143), .B(u5_mult_82_SUMB_46__18_), .ZN(u5_mult_82_SUMB_47__17_) );
  NAND3_X2 u5_mult_82_U4585 ( .A1(u5_mult_82_n1237), .A2(u5_mult_82_n1238), 
        .A3(u5_mult_82_n1239), .ZN(u5_mult_82_CARRYB_26__27_) );
  XNOR2_X2 u5_mult_82_U4584 ( .A(u5_mult_82_ab_36__26_), .B(
        u5_mult_82_CARRYB_35__26_), .ZN(u5_mult_82_n1142) );
  XNOR2_X2 u5_mult_82_U4583 ( .A(u5_mult_82_n1142), .B(u5_mult_82_SUMB_35__27_), .ZN(u5_mult_82_SUMB_36__26_) );
  NAND2_X2 u5_mult_82_U4582 ( .A1(u5_mult_82_CARRYB_9__42_), .A2(
        u5_mult_82_SUMB_9__43_), .ZN(u5_mult_82_n5399) );
  AND2_X2 u5_mult_82_U4581 ( .A1(u5_mult_82_n4531), .A2(u5_mult_82_n4532), 
        .ZN(u5_mult_82_n3691) );
  NAND2_X2 u5_mult_82_U4580 ( .A1(u5_mult_82_ab_30__15_), .A2(
        u5_mult_82_SUMB_29__16_), .ZN(u5_mult_82_n3657) );
  NAND3_X4 u5_mult_82_U4579 ( .A1(u5_mult_82_n1139), .A2(u5_mult_82_n1140), 
        .A3(u5_mult_82_n1141), .ZN(u5_mult_82_CARRYB_25__28_) );
  NAND2_X2 u5_mult_82_U4578 ( .A1(u5_mult_82_CARRYB_24__28_), .A2(
        u5_mult_82_SUMB_24__29_), .ZN(u5_mult_82_n1141) );
  NAND2_X2 u5_mult_82_U4577 ( .A1(u5_mult_82_ab_25__28_), .A2(
        u5_mult_82_SUMB_24__29_), .ZN(u5_mult_82_n1140) );
  NAND3_X2 u5_mult_82_U4576 ( .A1(u5_mult_82_n1136), .A2(u5_mult_82_n1137), 
        .A3(u5_mult_82_n1138), .ZN(u5_mult_82_CARRYB_24__29_) );
  NAND2_X2 u5_mult_82_U4575 ( .A1(u5_mult_82_CARRYB_23__29_), .A2(
        u5_mult_82_ab_24__29_), .ZN(u5_mult_82_n1138) );
  NAND2_X1 u5_mult_82_U4574 ( .A1(u5_mult_82_SUMB_23__30_), .A2(
        u5_mult_82_ab_24__29_), .ZN(u5_mult_82_n1137) );
  NAND2_X1 u5_mult_82_U4573 ( .A1(u5_mult_82_SUMB_23__30_), .A2(
        u5_mult_82_CARRYB_23__29_), .ZN(u5_mult_82_n1136) );
  XOR2_X2 u5_mult_82_U4572 ( .A(u5_mult_82_n1135), .B(u5_mult_82_SUMB_24__29_), 
        .Z(u5_mult_82_SUMB_25__28_) );
  NAND3_X4 u5_mult_82_U4571 ( .A1(u5_mult_82_n1132), .A2(u5_mult_82_n1133), 
        .A3(u5_mult_82_n1134), .ZN(u5_mult_82_CARRYB_41__19_) );
  NAND2_X1 u5_mult_82_U4570 ( .A1(u5_mult_82_ab_41__19_), .A2(
        u5_mult_82_CARRYB_40__19_), .ZN(u5_mult_82_n1132) );
  NAND3_X2 u5_mult_82_U4569 ( .A1(u5_mult_82_n1129), .A2(u5_mult_82_n1130), 
        .A3(u5_mult_82_n1131), .ZN(u5_mult_82_CARRYB_40__20_) );
  NAND2_X1 u5_mult_82_U4568 ( .A1(u5_mult_82_CARRYB_39__20_), .A2(
        u5_mult_82_SUMB_39__21_), .ZN(u5_mult_82_n1131) );
  NAND2_X1 u5_mult_82_U4567 ( .A1(u5_mult_82_ab_40__20_), .A2(
        u5_mult_82_SUMB_39__21_), .ZN(u5_mult_82_n1130) );
  NAND2_X1 u5_mult_82_U4566 ( .A1(u5_mult_82_ab_40__20_), .A2(
        u5_mult_82_CARRYB_39__20_), .ZN(u5_mult_82_n1129) );
  XOR2_X2 u5_mult_82_U4565 ( .A(u5_mult_82_n1128), .B(u5_mult_82_SUMB_40__20_), 
        .Z(u5_mult_82_SUMB_41__19_) );
  XOR2_X2 u5_mult_82_U4564 ( .A(u5_mult_82_ab_41__19_), .B(
        u5_mult_82_CARRYB_40__19_), .Z(u5_mult_82_n1128) );
  INV_X4 u5_mult_82_U4563 ( .A(u5_mult_82_ab_20__32_), .ZN(u5_mult_82_n1125)
         );
  NAND2_X2 u5_mult_82_U4562 ( .A1(u5_mult_82_n1125), .A2(u5_mult_82_n1126), 
        .ZN(u5_mult_82_n1127) );
  NOR2_X1 u5_mult_82_U4561 ( .A1(u5_mult_82_n6862), .A2(u5_mult_82_n6684), 
        .ZN(u5_mult_82_ab_31__29_) );
  NAND2_X2 u5_mult_82_U4560 ( .A1(u5_mult_82_ab_50__19_), .A2(
        u5_mult_82_CARRYB_49__19_), .ZN(u5_mult_82_n5566) );
  NOR2_X2 u5_mult_82_U4559 ( .A1(u5_mult_82_n6912), .A2(u5_mult_82_n6754), 
        .ZN(u5_mult_82_ab_49__19_) );
  NAND3_X2 u5_mult_82_U4558 ( .A1(u5_mult_82_n1122), .A2(u5_mult_82_n1123), 
        .A3(u5_mult_82_n1124), .ZN(u5_mult_82_CARRYB_31__29_) );
  NAND2_X1 u5_mult_82_U4557 ( .A1(u5_mult_82_ab_31__29_), .A2(
        u5_mult_82_CARRYB_30__29_), .ZN(u5_mult_82_n1124) );
  NAND2_X2 u5_mult_82_U4556 ( .A1(u5_mult_82_ab_31__29_), .A2(
        u5_mult_82_SUMB_30__30_), .ZN(u5_mult_82_n1123) );
  NAND2_X1 u5_mult_82_U4555 ( .A1(u5_mult_82_CARRYB_30__29_), .A2(
        u5_mult_82_SUMB_30__30_), .ZN(u5_mult_82_n1122) );
  XOR2_X2 u5_mult_82_U4554 ( .A(u5_mult_82_SUMB_30__30_), .B(u5_mult_82_n1121), 
        .Z(u5_mult_82_SUMB_31__29_) );
  XOR2_X2 u5_mult_82_U4553 ( .A(u5_mult_82_CARRYB_30__29_), .B(
        u5_mult_82_ab_31__29_), .Z(u5_mult_82_n1121) );
  NAND3_X2 u5_mult_82_U4552 ( .A1(u5_mult_82_n1118), .A2(u5_mult_82_n1119), 
        .A3(u5_mult_82_n1120), .ZN(u5_mult_82_CARRYB_49__19_) );
  NAND2_X1 u5_mult_82_U4551 ( .A1(u5_mult_82_ab_49__19_), .A2(
        u5_mult_82_CARRYB_48__19_), .ZN(u5_mult_82_n1120) );
  NAND2_X2 u5_mult_82_U4550 ( .A1(u5_mult_82_ab_49__19_), .A2(
        u5_mult_82_SUMB_48__20_), .ZN(u5_mult_82_n1119) );
  NAND2_X1 u5_mult_82_U4549 ( .A1(u5_mult_82_CARRYB_48__19_), .A2(
        u5_mult_82_SUMB_48__20_), .ZN(u5_mult_82_n1118) );
  XNOR2_X2 u5_mult_82_U4548 ( .A(u5_mult_82_n1117), .B(
        u5_mult_82_CARRYB_45__28_), .ZN(u5_mult_82_n3066) );
  NAND2_X2 u5_mult_82_U4547 ( .A1(u5_mult_82_ab_28__31_), .A2(
        u5_mult_82_CARRYB_27__31_), .ZN(u5_mult_82_n2813) );
  NAND2_X1 u5_mult_82_U4546 ( .A1(u5_mult_82_ab_41__22_), .A2(
        u5_mult_82_SUMB_40__23_), .ZN(u5_mult_82_n2250) );
  XNOR2_X2 u5_mult_82_U4545 ( .A(u5_mult_82_ab_50__8_), .B(
        u5_mult_82_CARRYB_49__8_), .ZN(u5_mult_82_n4182) );
  NAND2_X2 u5_mult_82_U4544 ( .A1(u5_mult_82_CARRYB_32__30_), .A2(
        u5_mult_82_SUMB_32__31_), .ZN(u5_mult_82_n5873) );
  NAND2_X2 u5_mult_82_U4543 ( .A1(u5_mult_82_ab_33__30_), .A2(
        u5_mult_82_SUMB_32__31_), .ZN(u5_mult_82_n5872) );
  NAND3_X2 u5_mult_82_U4542 ( .A1(u5_mult_82_net81828), .A2(
        u5_mult_82_net81829), .A3(u5_mult_82_net81830), .ZN(
        u5_mult_82_CARRYB_49__7_) );
  NOR2_X2 u5_mult_82_U4541 ( .A1(u5_mult_82_n6827), .A2(u5_mult_82_n6664), 
        .ZN(u5_mult_82_ab_28__40_) );
  NAND3_X4 u5_mult_82_U4540 ( .A1(u5_mult_82_n2680), .A2(u5_mult_82_n2681), 
        .A3(u5_mult_82_n2682), .ZN(u5_mult_82_CARRYB_27__40_) );
  NAND2_X2 u5_mult_82_U4539 ( .A1(u5_mult_82_ab_50__26_), .A2(
        u5_mult_82_CARRYB_49__26_), .ZN(u5_mult_82_n4184) );
  NOR2_X2 u5_mult_82_U4538 ( .A1(u5_mult_82_n6879), .A2(u5_mult_82_n6754), 
        .ZN(u5_mult_82_ab_49__26_) );
  NAND3_X4 u5_mult_82_U4537 ( .A1(u5_mult_82_n1114), .A2(u5_mult_82_n1115), 
        .A3(u5_mult_82_n1116), .ZN(u5_mult_82_CARRYB_38__33_) );
  NAND2_X2 u5_mult_82_U4536 ( .A1(u5_mult_82_CARRYB_37__33_), .A2(
        u5_mult_82_SUMB_37__34_), .ZN(u5_mult_82_n1116) );
  NAND2_X2 u5_mult_82_U4535 ( .A1(u5_mult_82_ab_38__33_), .A2(
        u5_mult_82_SUMB_37__34_), .ZN(u5_mult_82_n1115) );
  NAND2_X1 u5_mult_82_U4534 ( .A1(u5_mult_82_ab_38__33_), .A2(
        u5_mult_82_CARRYB_37__33_), .ZN(u5_mult_82_n1114) );
  NAND3_X2 u5_mult_82_U4533 ( .A1(u5_mult_82_n1111), .A2(u5_mult_82_n1112), 
        .A3(u5_mult_82_n1113), .ZN(u5_mult_82_CARRYB_37__34_) );
  NAND2_X2 u5_mult_82_U4532 ( .A1(u5_mult_82_CARRYB_36__34_), .A2(
        u5_mult_82_SUMB_36__35_), .ZN(u5_mult_82_n1113) );
  NAND2_X2 u5_mult_82_U4531 ( .A1(u5_mult_82_ab_37__34_), .A2(
        u5_mult_82_SUMB_36__35_), .ZN(u5_mult_82_n1112) );
  NAND2_X1 u5_mult_82_U4530 ( .A1(u5_mult_82_ab_37__34_), .A2(
        u5_mult_82_CARRYB_36__34_), .ZN(u5_mult_82_n1111) );
  XOR2_X2 u5_mult_82_U4529 ( .A(u5_mult_82_n1110), .B(u5_mult_82_SUMB_37__34_), 
        .Z(u5_mult_82_SUMB_38__33_) );
  XOR2_X2 u5_mult_82_U4528 ( .A(u5_mult_82_ab_38__33_), .B(
        u5_mult_82_CARRYB_37__33_), .Z(u5_mult_82_n1110) );
  NAND3_X2 u5_mult_82_U4527 ( .A1(u5_mult_82_n1107), .A2(u5_mult_82_n1108), 
        .A3(u5_mult_82_n1109), .ZN(u5_mult_82_CARRYB_28__40_) );
  NAND2_X1 u5_mult_82_U4526 ( .A1(u5_mult_82_CARRYB_27__40_), .A2(
        u5_mult_82_ab_28__40_), .ZN(u5_mult_82_n1109) );
  NAND2_X1 u5_mult_82_U4525 ( .A1(u5_mult_82_CARRYB_27__40_), .A2(
        u5_mult_82_SUMB_27__41_), .ZN(u5_mult_82_n1107) );
  XOR2_X2 u5_mult_82_U4524 ( .A(u5_mult_82_CARRYB_27__40_), .B(
        u5_mult_82_ab_28__40_), .Z(u5_mult_82_n1106) );
  NAND3_X2 u5_mult_82_U4523 ( .A1(u5_mult_82_n1103), .A2(u5_mult_82_n1104), 
        .A3(u5_mult_82_n1105), .ZN(u5_mult_82_CARRYB_49__26_) );
  NAND2_X1 u5_mult_82_U4522 ( .A1(u5_mult_82_ab_49__26_), .A2(
        u5_mult_82_CARRYB_48__26_), .ZN(u5_mult_82_n1105) );
  NAND2_X1 u5_mult_82_U4521 ( .A1(u5_mult_82_ab_49__26_), .A2(
        u5_mult_82_SUMB_48__27_), .ZN(u5_mult_82_n1104) );
  NAND2_X1 u5_mult_82_U4520 ( .A1(u5_mult_82_CARRYB_48__26_), .A2(
        u5_mult_82_SUMB_48__27_), .ZN(u5_mult_82_n1103) );
  NAND2_X2 u5_mult_82_U4519 ( .A1(u5_mult_82_ab_48__8_), .A2(
        u5_mult_82_CARRYB_47__8_), .ZN(u5_mult_82_net81825) );
  NAND2_X2 u5_mult_82_U4518 ( .A1(u5_mult_82_CARRYB_39__12_), .A2(
        u5_mult_82_SUMB_39__13_), .ZN(u5_mult_82_net82472) );
  NAND2_X2 u5_mult_82_U4517 ( .A1(u5_mult_82_CARRYB_42__18_), .A2(
        u5_mult_82_SUMB_42__19_), .ZN(u5_mult_82_n4234) );
  NAND2_X2 u5_mult_82_U4516 ( .A1(u5_mult_82_ab_32__40_), .A2(
        u5_mult_82_CARRYB_31__40_), .ZN(u5_mult_82_n3837) );
  NAND2_X2 u5_mult_82_U4515 ( .A1(u5_mult_82_ab_32__40_), .A2(
        u5_mult_82_SUMB_31__41_), .ZN(u5_mult_82_n3838) );
  NAND2_X2 u5_mult_82_U4514 ( .A1(u5_mult_82_n1299), .A2(u5_mult_82_n1300), 
        .ZN(u5_mult_82_SUMB_49__6_) );
  NAND2_X2 u5_mult_82_U4513 ( .A1(u5_mult_82_CARRYB_44__8_), .A2(
        u5_mult_82_n2745), .ZN(u5_mult_82_n2746) );
  XNOR2_X2 u5_mult_82_U4512 ( .A(u5_mult_82_CARRYB_21__44_), .B(
        u5_mult_82_n1102), .ZN(u5_mult_82_n3945) );
  NAND2_X1 u5_mult_82_U4511 ( .A1(u5_mult_82_CARRYB_28__18_), .A2(
        u5_mult_82_SUMB_28__19_), .ZN(u5_mult_82_n4562) );
  XNOR2_X1 u5_mult_82_U4510 ( .A(u5_mult_82_CARRYB_15__27_), .B(
        u5_mult_82_ab_16__27_), .ZN(u5_mult_82_net83139) );
  NAND2_X2 u5_mult_82_U4509 ( .A1(u5_mult_82_CARRYB_40__0_), .A2(
        u5_mult_82_SUMB_40__1_), .ZN(u5_mult_82_n2033) );
  NAND2_X2 u5_mult_82_U4508 ( .A1(u5_mult_82_ab_48__19_), .A2(
        u5_mult_82_SUMB_47__20_), .ZN(u5_mult_82_n4392) );
  NAND2_X2 u5_mult_82_U4507 ( .A1(u5_mult_82_CARRYB_43__20_), .A2(
        u5_mult_82_SUMB_43__21_), .ZN(u5_mult_82_n5341) );
  INV_X4 u5_mult_82_U4506 ( .A(u5_mult_82_n1771), .ZN(u5_mult_82_n1772) );
  INV_X8 u5_mult_82_U4505 ( .A(u5_mult_82_n7021), .ZN(u5_mult_82_n6918) );
  NAND2_X2 u5_mult_82_U4504 ( .A1(u5_mult_82_ab_19__47_), .A2(
        u5_mult_82_SUMB_18__48_), .ZN(u5_mult_82_n3107) );
  NAND2_X2 u5_mult_82_U4503 ( .A1(u5_mult_82_ab_20__40_), .A2(u5_mult_82_n66), 
        .ZN(u5_mult_82_n4942) );
  XNOR2_X2 u5_mult_82_U4502 ( .A(u5_mult_82_ab_21__40_), .B(
        u5_mult_82_CARRYB_20__40_), .ZN(u5_mult_82_n1786) );
  NAND2_X2 u5_mult_82_U4501 ( .A1(u5_mult_82_CARRYB_47__25_), .A2(
        u5_mult_82_SUMB_47__26_), .ZN(u5_mult_82_n4579) );
  INV_X4 u5_mult_82_U4500 ( .A(u5_mult_82_SUMB_24__35_), .ZN(u5_mult_82_n1817)
         );
  NAND2_X2 u5_mult_82_U4499 ( .A1(u5_mult_82_ab_34__30_), .A2(u5_mult_82_n1496), .ZN(u5_mult_82_n5950) );
  NAND3_X4 u5_mult_82_U4498 ( .A1(u5_mult_82_n5949), .A2(u5_mult_82_n5950), 
        .A3(u5_mult_82_n5951), .ZN(u5_mult_82_CARRYB_34__30_) );
  NAND2_X2 u5_mult_82_U4497 ( .A1(u5_mult_82_n2631), .A2(
        u5_mult_82_SUMB_16__26_), .ZN(u5_mult_82_n4631) );
  NAND2_X2 u5_mult_82_U4496 ( .A1(u5_mult_82_SUMB_21__24_), .A2(
        u5_mult_82_CARRYB_21__23_), .ZN(u5_mult_82_n1345) );
  INV_X4 u5_mult_82_U4495 ( .A(u5_mult_82_n2322), .ZN(u5_mult_82_n1098) );
  INV_X4 u5_mult_82_U4494 ( .A(u5_mult_82_net87430), .ZN(u5_mult_82_n1097) );
  NAND2_X4 u5_mult_82_U4493 ( .A1(u5_mult_82_n1099), .A2(u5_mult_82_n1100), 
        .ZN(u5_mult_82_SUMB_21__24_) );
  NAND2_X4 u5_mult_82_U4492 ( .A1(u5_mult_82_n1097), .A2(u5_mult_82_n1098), 
        .ZN(u5_mult_82_n1100) );
  NAND2_X2 u5_mult_82_U4491 ( .A1(u5_mult_82_net87430), .A2(u5_mult_82_n2322), 
        .ZN(u5_mult_82_n1099) );
  NAND3_X2 u5_mult_82_U4490 ( .A1(u5_mult_82_n1094), .A2(u5_mult_82_n1095), 
        .A3(u5_mult_82_n1096), .ZN(u5_mult_82_CARRYB_12__30_) );
  NAND2_X1 u5_mult_82_U4489 ( .A1(u5_mult_82_CARRYB_11__30_), .A2(
        u5_mult_82_SUMB_11__31_), .ZN(u5_mult_82_n1096) );
  NAND2_X1 u5_mult_82_U4488 ( .A1(u5_mult_82_ab_12__30_), .A2(
        u5_mult_82_SUMB_11__31_), .ZN(u5_mult_82_n1095) );
  NAND2_X1 u5_mult_82_U4487 ( .A1(u5_mult_82_ab_12__30_), .A2(
        u5_mult_82_CARRYB_11__30_), .ZN(u5_mult_82_n1094) );
  NAND3_X2 u5_mult_82_U4486 ( .A1(u5_mult_82_n1091), .A2(u5_mult_82_n1092), 
        .A3(u5_mult_82_n1093), .ZN(u5_mult_82_CARRYB_11__31_) );
  NAND2_X2 u5_mult_82_U4485 ( .A1(u5_mult_82_ab_11__31_), .A2(
        u5_mult_82_SUMB_10__32_), .ZN(u5_mult_82_n1093) );
  NAND2_X2 u5_mult_82_U4484 ( .A1(u5_mult_82_CARRYB_10__31_), .A2(
        u5_mult_82_SUMB_10__32_), .ZN(u5_mult_82_n1092) );
  NAND2_X1 u5_mult_82_U4483 ( .A1(u5_mult_82_CARRYB_10__31_), .A2(
        u5_mult_82_ab_11__31_), .ZN(u5_mult_82_n1091) );
  XOR2_X2 u5_mult_82_U4482 ( .A(u5_mult_82_n1090), .B(u5_mult_82_SUMB_10__32_), 
        .Z(u5_mult_82_SUMB_11__31_) );
  XOR2_X2 u5_mult_82_U4481 ( .A(u5_mult_82_CARRYB_10__31_), .B(
        u5_mult_82_ab_11__31_), .Z(u5_mult_82_n1090) );
  XNOR2_X2 u5_mult_82_U4480 ( .A(u5_mult_82_ab_45__24_), .B(
        u5_mult_82_CARRYB_44__24_), .ZN(u5_mult_82_n1089) );
  XNOR2_X2 u5_mult_82_U4479 ( .A(u5_mult_82_n1089), .B(u5_mult_82_SUMB_44__25_), .ZN(u5_mult_82_SUMB_45__24_) );
  NAND3_X2 u5_mult_82_U4478 ( .A1(u5_mult_82_n3947), .A2(u5_mult_82_n3948), 
        .A3(u5_mult_82_n3949), .ZN(u5_mult_82_CARRYB_22__44_) );
  INV_X4 u5_mult_82_U4477 ( .A(u5_mult_82_n1825), .ZN(u5_mult_82_n1826) );
  XNOR2_X2 u5_mult_82_U4476 ( .A(u5_mult_82_ab_48__17_), .B(
        u5_mult_82_CARRYB_47__17_), .ZN(u5_mult_82_n1088) );
  XNOR2_X2 u5_mult_82_U4475 ( .A(u5_mult_82_n1088), .B(u5_mult_82_SUMB_47__18_), .ZN(u5_mult_82_SUMB_48__17_) );
  INV_X8 u5_mult_82_U4474 ( .A(u5_mult_82_n6418), .ZN(u5_mult_82_CLA_SUM[82])
         );
  NAND2_X2 u5_mult_82_U4473 ( .A1(u5_mult_82_ab_48__0_), .A2(
        u5_mult_82_CARRYB_47__0_), .ZN(u5_mult_82_n2030) );
  NAND2_X2 u5_mult_82_U4472 ( .A1(u5_mult_82_ab_25__17_), .A2(
        u5_mult_82_SUMB_24__18_), .ZN(u5_mult_82_n5380) );
  NAND2_X2 u5_mult_82_U4471 ( .A1(u5_mult_82_CARRYB_24__17_), .A2(
        u5_mult_82_SUMB_24__18_), .ZN(u5_mult_82_n5381) );
  NAND3_X4 u5_mult_82_U4470 ( .A1(u5_mult_82_n4895), .A2(u5_mult_82_n4896), 
        .A3(u5_mult_82_n4897), .ZN(u5_mult_82_CARRYB_27__16_) );
  NAND2_X1 u5_mult_82_U4469 ( .A1(u5_mult_82_ab_50__17_), .A2(
        u5_mult_82_CARRYB_49__17_), .ZN(u5_mult_82_n4398) );
  NAND2_X2 u5_mult_82_U4468 ( .A1(u5_mult_82_SUMB_47__1_), .A2(
        u5_mult_82_CARRYB_47__0_), .ZN(u5_mult_82_n2029) );
  NAND2_X1 u5_mult_82_U4467 ( .A1(u5_mult_82_ab_17__36_), .A2(
        u5_mult_82_CARRYB_16__36_), .ZN(u5_mult_82_n6310) );
  XNOR2_X2 u5_mult_82_U4466 ( .A(u5_mult_82_n695), .B(u5_mult_82_n1466), .ZN(
        u5_mult_82_SUMB_21__23_) );
  NAND3_X4 u5_mult_82_U4465 ( .A1(u5_mult_82_n6071), .A2(u5_mult_82_n6072), 
        .A3(u5_mult_82_n6073), .ZN(u5_mult_82_CARRYB_43__7_) );
  NAND2_X2 u5_mult_82_U4464 ( .A1(u5_mult_82_ab_43__33_), .A2(
        u5_mult_82_SUMB_42__34_), .ZN(u5_mult_82_n3039) );
  NAND2_X2 u5_mult_82_U4463 ( .A1(u5_mult_82_CARRYB_42__33_), .A2(
        u5_mult_82_SUMB_42__34_), .ZN(u5_mult_82_n3040) );
  NAND2_X2 u5_mult_82_U4462 ( .A1(u5_mult_82_CARRYB_41__2_), .A2(
        u5_mult_82_SUMB_41__3_), .ZN(u5_mult_82_n5631) );
  NAND2_X2 u5_mult_82_U4461 ( .A1(u5_mult_82_SUMB_30__4_), .A2(
        u5_mult_82_CARRYB_30__3_), .ZN(u5_mult_82_n2037) );
  INV_X4 u5_mult_82_U4460 ( .A(u5_mult_82_CARRYB_24__33_), .ZN(
        u5_mult_82_n3381) );
  NAND2_X4 u5_mult_82_U4459 ( .A1(u5_mult_82_n1705), .A2(u5_mult_82_n704), 
        .ZN(u5_mult_82_n5473) );
  XNOR2_X2 u5_mult_82_U4458 ( .A(u5_mult_82_CARRYB_50__36_), .B(
        u5_mult_82_ab_51__36_), .ZN(u5_mult_82_n1087) );
  XNOR2_X2 u5_mult_82_U4457 ( .A(u5_mult_82_SUMB_50__37_), .B(u5_mult_82_n1087), .ZN(u5_mult_82_SUMB_51__36_) );
  NAND3_X2 u5_mult_82_U4456 ( .A1(u5_mult_82_n6310), .A2(u5_mult_82_n6311), 
        .A3(u5_mult_82_n6312), .ZN(u5_mult_82_CARRYB_17__36_) );
  XNOR2_X2 u5_mult_82_U4455 ( .A(u5_mult_82_ab_25__41_), .B(
        u5_mult_82_CARRYB_24__41_), .ZN(u5_mult_82_n1086) );
  XNOR2_X2 u5_mult_82_U4454 ( .A(u5_mult_82_n1086), .B(u5_mult_82_SUMB_24__42_), .ZN(u5_mult_82_SUMB_25__41_) );
  NAND2_X2 u5_mult_82_U4453 ( .A1(u5_mult_82_SUMB_11__51_), .A2(
        u5_mult_82_CARRYB_11__50_), .ZN(u5_mult_82_n3604) );
  NAND2_X2 u5_mult_82_U4452 ( .A1(u5_mult_82_SUMB_34__34_), .A2(
        u5_mult_82_CARRYB_34__33_), .ZN(u5_mult_82_n3610) );
  NAND2_X2 u5_mult_82_U4451 ( .A1(u5_mult_82_ab_40__30_), .A2(
        u5_mult_82_SUMB_39__31_), .ZN(u5_mult_82_n4918) );
  NAND3_X2 u5_mult_82_U4450 ( .A1(u5_mult_82_n5170), .A2(u5_mult_82_n5171), 
        .A3(u5_mult_82_n5172), .ZN(u5_mult_82_CARRYB_12__42_) );
  CLKBUF_X3 u5_mult_82_U4449 ( .A(u5_mult_82_SUMB_45__11_), .Z(
        u5_mult_82_n1488) );
  XOR2_X2 u5_mult_82_U4448 ( .A(u5_mult_82_SUMB_52__7_), .B(
        u5_mult_82_CARRYB_52__6_), .Z(u5_mult_82_n5330) );
  NAND3_X2 u5_mult_82_U4447 ( .A1(u5_mult_82_n5589), .A2(u5_mult_82_n5590), 
        .A3(u5_mult_82_n5591), .ZN(u5_mult_82_CARRYB_25__44_) );
  XNOR2_X2 u5_mult_82_U4446 ( .A(u5_mult_82_ab_18__20_), .B(
        u5_mult_82_CARRYB_17__20_), .ZN(u5_mult_82_n1085) );
  XNOR2_X2 u5_mult_82_U4445 ( .A(u5_mult_82_n1085), .B(u5_mult_82_SUMB_17__21_), .ZN(u5_mult_82_SUMB_18__20_) );
  NAND3_X2 u5_mult_82_U4444 ( .A1(u5_mult_82_n1082), .A2(u5_mult_82_n1083), 
        .A3(u5_mult_82_n1084), .ZN(u5_mult_82_CARRYB_44__42_) );
  NAND2_X1 u5_mult_82_U4443 ( .A1(u5_mult_82_CARRYB_43__42_), .A2(
        u5_mult_82_SUMB_43__43_), .ZN(u5_mult_82_n1084) );
  NAND2_X1 u5_mult_82_U4442 ( .A1(u5_mult_82_ab_44__42_), .A2(
        u5_mult_82_SUMB_43__43_), .ZN(u5_mult_82_n1083) );
  NAND2_X1 u5_mult_82_U4441 ( .A1(u5_mult_82_ab_44__42_), .A2(
        u5_mult_82_CARRYB_43__42_), .ZN(u5_mult_82_n1082) );
  NAND3_X4 u5_mult_82_U4440 ( .A1(u5_mult_82_n1079), .A2(u5_mult_82_n1080), 
        .A3(u5_mult_82_n1081), .ZN(u5_mult_82_CARRYB_43__43_) );
  NAND2_X2 u5_mult_82_U4439 ( .A1(u5_mult_82_CARRYB_42__43_), .A2(
        u5_mult_82_SUMB_42__44_), .ZN(u5_mult_82_n1081) );
  NAND2_X2 u5_mult_82_U4438 ( .A1(u5_mult_82_ab_43__43_), .A2(
        u5_mult_82_SUMB_42__44_), .ZN(u5_mult_82_n1080) );
  NAND2_X2 u5_mult_82_U4437 ( .A1(u5_mult_82_ab_43__43_), .A2(
        u5_mult_82_CARRYB_42__43_), .ZN(u5_mult_82_n1079) );
  XOR2_X2 u5_mult_82_U4436 ( .A(u5_mult_82_n1078), .B(u5_mult_82_SUMB_43__43_), 
        .Z(u5_mult_82_SUMB_44__42_) );
  XOR2_X2 u5_mult_82_U4435 ( .A(u5_mult_82_ab_44__42_), .B(
        u5_mult_82_CARRYB_43__42_), .Z(u5_mult_82_n1078) );
  XOR2_X2 u5_mult_82_U4434 ( .A(u5_mult_82_n1077), .B(u5_mult_82_SUMB_42__44_), 
        .Z(u5_mult_82_SUMB_43__43_) );
  XOR2_X2 u5_mult_82_U4433 ( .A(u5_mult_82_ab_43__43_), .B(
        u5_mult_82_CARRYB_42__43_), .Z(u5_mult_82_n1077) );
  XNOR2_X2 u5_mult_82_U4432 ( .A(u5_mult_82_n383), .B(u5_mult_82_n2690), .ZN(
        u5_mult_82_SUMB_39__5_) );
  NAND3_X2 u5_mult_82_U4431 ( .A1(u5_mult_82_n5791), .A2(u5_mult_82_n5793), 
        .A3(u5_mult_82_n5792), .ZN(u5_mult_82_CARRYB_45__3_) );
  NAND2_X1 u5_mult_82_U4430 ( .A1(u5_mult_82_ab_43__5_), .A2(
        u5_mult_82_SUMB_42__6_), .ZN(u5_mult_82_n5245) );
  NAND2_X1 u5_mult_82_U4429 ( .A1(u5_mult_82_SUMB_42__6_), .A2(
        u5_mult_82_CARRYB_42__5_), .ZN(u5_mult_82_n5243) );
  XOR2_X2 u5_mult_82_U4428 ( .A(u5_mult_82_ab_44__31_), .B(
        u5_mult_82_CARRYB_43__31_), .Z(u5_mult_82_n3019) );
  NAND2_X1 u5_mult_82_U4427 ( .A1(u5_mult_82_n5550), .A2(
        u5_mult_82_SUMB_17__47_), .ZN(u5_mult_82_n5254) );
  NAND2_X1 u5_mult_82_U4426 ( .A1(u5_mult_82_ab_39__9_), .A2(
        u5_mult_82_CARRYB_38__9_), .ZN(u5_mult_82_n4771) );
  INV_X16 u5_mult_82_U4425 ( .A(n4813), .ZN(u5_mult_82_n6758) );
  NAND3_X4 u5_mult_82_U4424 ( .A1(u5_mult_82_n5933), .A2(u5_mult_82_n5934), 
        .A3(u5_mult_82_n5935), .ZN(u5_mult_82_CARRYB_43__8_) );
  INV_X2 u5_mult_82_U4423 ( .A(u5_mult_82_CARRYB_41__8_), .ZN(u5_mult_82_n1561) );
  NAND2_X2 u5_mult_82_U4422 ( .A1(u5_mult_82_ab_42__8_), .A2(
        u5_mult_82_CARRYB_41__8_), .ZN(u5_mult_82_n4386) );
  NAND2_X1 u5_mult_82_U4421 ( .A1(u5_mult_82_ab_49__18_), .A2(
        u5_mult_82_CARRYB_48__18_), .ZN(u5_mult_82_n4395) );
  XNOR2_X2 u5_mult_82_U4420 ( .A(u5_mult_82_CARRYB_43__5_), .B(
        u5_mult_82_ab_44__5_), .ZN(u5_mult_82_n1620) );
  XOR2_X1 u5_mult_82_U4419 ( .A(u5_mult_82_CARRYB_42__35_), .B(
        u5_mult_82_ab_43__35_), .Z(u5_mult_82_n3355) );
  INV_X2 u5_mult_82_U4418 ( .A(u5_mult_82_n2712), .ZN(u5_mult_82_n2075) );
  NAND2_X2 u5_mult_82_U4417 ( .A1(u5_mult_82_n2712), .A2(
        u5_mult_82_SUMB_47__34_), .ZN(u5_mult_82_n2077) );
  XNOR2_X2 u5_mult_82_U4416 ( .A(u5_mult_82_ab_12__30_), .B(
        u5_mult_82_CARRYB_11__30_), .ZN(u5_mult_82_n1076) );
  XNOR2_X2 u5_mult_82_U4415 ( .A(u5_mult_82_n1076), .B(u5_mult_82_SUMB_11__31_), .ZN(u5_mult_82_SUMB_12__30_) );
  NAND2_X2 u5_mult_82_U4414 ( .A1(u5_mult_82_n402), .A2(
        u5_mult_82_SUMB_22__27_), .ZN(u5_mult_82_n1905) );
  NAND3_X2 u5_mult_82_U4413 ( .A1(u5_mult_82_n5523), .A2(u5_mult_82_n5524), 
        .A3(u5_mult_82_n5525), .ZN(u5_mult_82_CARRYB_37__16_) );
  NAND2_X2 u5_mult_82_U4412 ( .A1(u5_mult_82_n738), .A2(
        u5_mult_82_CARRYB_36__16_), .ZN(u5_mult_82_n5523) );
  NAND3_X2 u5_mult_82_U4411 ( .A1(u5_mult_82_n4744), .A2(u5_mult_82_n4745), 
        .A3(u5_mult_82_n4746), .ZN(u5_mult_82_CARRYB_7__38_) );
  XOR2_X2 u5_mult_82_U4410 ( .A(u5_mult_82_SUMB_52__34_), .B(
        u5_mult_82_CARRYB_52__33_), .Z(u5_mult_82_n1075) );
  NAND2_X2 u5_mult_82_U4409 ( .A1(u5_mult_82_ab_43__18_), .A2(
        u5_mult_82_SUMB_42__19_), .ZN(u5_mult_82_n4233) );
  NAND2_X2 u5_mult_82_U4408 ( .A1(u5_mult_82_CARRYB_20__23_), .A2(
        u5_mult_82_SUMB_20__24_), .ZN(u5_mult_82_n3615) );
  NAND2_X2 u5_mult_82_U4407 ( .A1(u5_mult_82_ab_19__35_), .A2(
        u5_mult_82_CARRYB_18__35_), .ZN(u5_mult_82_n3109) );
  NAND2_X2 u5_mult_82_U4406 ( .A1(u5_mult_82_CARRYB_22__41_), .A2(
        u5_mult_82_SUMB_22__42_), .ZN(u5_mult_82_n3027) );
  NAND2_X2 u5_mult_82_U4405 ( .A1(u5_mult_82_ab_31__16_), .A2(
        u5_mult_82_CARRYB_30__16_), .ZN(u5_mult_82_n4358) );
  NAND2_X4 u5_mult_82_U4404 ( .A1(u5_mult_82_CARRYB_41__9_), .A2(
        u5_mult_82_ab_42__9_), .ZN(u5_mult_82_n3650) );
  NAND3_X4 u5_mult_82_U4403 ( .A1(u5_mult_82_n4636), .A2(u5_mult_82_n4637), 
        .A3(u5_mult_82_n4638), .ZN(u5_mult_82_CARRYB_20__22_) );
  XNOR2_X2 u5_mult_82_U4402 ( .A(u5_mult_82_ab_45__34_), .B(u5_mult_82_n42), 
        .ZN(u5_mult_82_n1735) );
  BUF_X2 u5_mult_82_U4401 ( .A(u5_mult_82_SUMB_45__34_), .Z(u5_mult_82_n1501)
         );
  NAND2_X2 u5_mult_82_U4400 ( .A1(u5_mult_82_CARRYB_21__34_), .A2(
        u5_mult_82_SUMB_21__35_), .ZN(u5_mult_82_n4991) );
  NAND2_X2 u5_mult_82_U4399 ( .A1(u5_mult_82_ab_22__34_), .A2(
        u5_mult_82_SUMB_21__35_), .ZN(u5_mult_82_n4990) );
  NAND3_X4 u5_mult_82_U4398 ( .A1(u5_mult_82_n1072), .A2(u5_mult_82_n1073), 
        .A3(u5_mult_82_n1074), .ZN(u5_mult_82_CARRYB_42__33_) );
  NAND2_X1 u5_mult_82_U4397 ( .A1(u5_mult_82_CARRYB_41__33_), .A2(
        u5_mult_82_SUMB_41__34_), .ZN(u5_mult_82_n1074) );
  NAND2_X1 u5_mult_82_U4396 ( .A1(u5_mult_82_ab_42__33_), .A2(
        u5_mult_82_SUMB_41__34_), .ZN(u5_mult_82_n1073) );
  NAND2_X1 u5_mult_82_U4395 ( .A1(u5_mult_82_ab_42__33_), .A2(
        u5_mult_82_CARRYB_41__33_), .ZN(u5_mult_82_n1072) );
  NAND2_X2 u5_mult_82_U4394 ( .A1(u5_mult_82_CARRYB_40__34_), .A2(
        u5_mult_82_SUMB_40__35_), .ZN(u5_mult_82_n1071) );
  NAND2_X2 u5_mult_82_U4393 ( .A1(u5_mult_82_ab_41__34_), .A2(
        u5_mult_82_SUMB_40__35_), .ZN(u5_mult_82_n1070) );
  NAND2_X1 u5_mult_82_U4392 ( .A1(u5_mult_82_ab_41__34_), .A2(
        u5_mult_82_CARRYB_40__34_), .ZN(u5_mult_82_n1069) );
  XOR2_X2 u5_mult_82_U4391 ( .A(u5_mult_82_n1068), .B(u5_mult_82_SUMB_41__34_), 
        .Z(u5_mult_82_SUMB_42__33_) );
  XOR2_X2 u5_mult_82_U4390 ( .A(u5_mult_82_ab_42__33_), .B(
        u5_mult_82_CARRYB_41__33_), .Z(u5_mult_82_n1068) );
  XOR2_X2 u5_mult_82_U4389 ( .A(u5_mult_82_n1067), .B(u5_mult_82_SUMB_40__35_), 
        .Z(u5_mult_82_SUMB_41__34_) );
  XOR2_X2 u5_mult_82_U4388 ( .A(u5_mult_82_ab_41__34_), .B(
        u5_mult_82_CARRYB_40__34_), .Z(u5_mult_82_n1067) );
  NOR2_X1 u5_mult_82_U4387 ( .A1(u5_mult_82_n6766), .A2(u5_mult_82_n6733), 
        .ZN(u5_mult_82_ab_44__50_) );
  NOR2_X1 u5_mult_82_U4386 ( .A1(u5_mult_82_n6766), .A2(u5_mult_82_net65313), 
        .ZN(u5_mult_82_ab_45__50_) );
  NOR2_X1 u5_mult_82_U4385 ( .A1(u5_mult_82_n6766), .A2(u5_mult_82_n6740), 
        .ZN(u5_mult_82_ab_46__50_) );
  NOR2_X1 u5_mult_82_U4384 ( .A1(u5_mult_82_n6766), .A2(u5_mult_82_net65277), 
        .ZN(u5_mult_82_ab_47__50_) );
  NOR2_X1 u5_mult_82_U4383 ( .A1(u5_mult_82_n6766), .A2(u5_mult_82_n6746), 
        .ZN(u5_mult_82_ab_48__50_) );
  NOR2_X1 u5_mult_82_U4382 ( .A1(u5_mult_82_n6766), .A2(u5_mult_82_n6752), 
        .ZN(u5_mult_82_ab_49__50_) );
  NOR2_X1 u5_mult_82_U4381 ( .A1(u5_mult_82_n6766), .A2(u5_mult_82_net65223), 
        .ZN(u5_mult_82_ab_50__50_) );
  NOR2_X1 u5_mult_82_U4380 ( .A1(u5_mult_82_n6766), .A2(u5_mult_82_net65191), 
        .ZN(u5_mult_82_ab_51__50_) );
  NOR2_X1 u5_mult_82_U4379 ( .A1(u5_mult_82_n6977), .A2(u5_mult_82_n6766), 
        .ZN(u5_mult_82_ab_52__50_) );
  NAND2_X2 u5_mult_82_U4378 ( .A1(u5_mult_82_ab_17__25_), .A2(u5_mult_82_n2631), .ZN(u5_mult_82_n4629) );
  XNOR2_X1 u5_mult_82_U4377 ( .A(u5_mult_82_CARRYB_22__41_), .B(
        u5_mult_82_ab_23__41_), .ZN(u5_mult_82_n1441) );
  NAND3_X4 u5_mult_82_U4376 ( .A1(u5_mult_82_n5670), .A2(u5_mult_82_n5671), 
        .A3(u5_mult_82_n5672), .ZN(u5_mult_82_CARRYB_26__38_) );
  NOR2_X1 u5_mult_82_U4375 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6656), 
        .ZN(u5_mult_82_ab_27__38_) );
  INV_X2 u5_mult_82_U4374 ( .A(u5_mult_82_n1441), .ZN(u5_mult_82_n1064) );
  INV_X2 u5_mult_82_U4373 ( .A(u5_mult_82_SUMB_22__42_), .ZN(u5_mult_82_n1063)
         );
  NAND2_X4 u5_mult_82_U4372 ( .A1(u5_mult_82_n1065), .A2(u5_mult_82_n1066), 
        .ZN(u5_mult_82_SUMB_23__41_) );
  NAND2_X4 u5_mult_82_U4371 ( .A1(u5_mult_82_n1063), .A2(u5_mult_82_n1064), 
        .ZN(u5_mult_82_n1066) );
  NAND2_X1 u5_mult_82_U4370 ( .A1(u5_mult_82_SUMB_22__42_), .A2(
        u5_mult_82_n1441), .ZN(u5_mult_82_n1065) );
  NAND3_X2 u5_mult_82_U4369 ( .A1(u5_mult_82_n1060), .A2(u5_mult_82_n1061), 
        .A3(u5_mult_82_n1062), .ZN(u5_mult_82_CARRYB_27__38_) );
  NAND2_X1 u5_mult_82_U4368 ( .A1(u5_mult_82_ab_27__38_), .A2(
        u5_mult_82_CARRYB_26__38_), .ZN(u5_mult_82_n1062) );
  NAND2_X2 u5_mult_82_U4367 ( .A1(u5_mult_82_ab_27__38_), .A2(
        u5_mult_82_SUMB_26__39_), .ZN(u5_mult_82_n1061) );
  XOR2_X2 u5_mult_82_U4366 ( .A(u5_mult_82_SUMB_26__39_), .B(u5_mult_82_n1059), 
        .Z(u5_mult_82_SUMB_27__38_) );
  XOR2_X2 u5_mult_82_U4365 ( .A(u5_mult_82_CARRYB_26__38_), .B(
        u5_mult_82_ab_27__38_), .Z(u5_mult_82_n1059) );
  NAND2_X4 u5_mult_82_U4364 ( .A1(u5_mult_82_n1818), .A2(u5_mult_82_ab_25__34_), .ZN(u5_mult_82_n5765) );
  NAND2_X4 u5_mult_82_U4363 ( .A1(u5_mult_82_n1818), .A2(
        u5_mult_82_CARRYB_24__34_), .ZN(u5_mult_82_n5766) );
  INV_X2 u5_mult_82_U4362 ( .A(u5_mult_82_n1552), .ZN(u5_mult_82_n1553) );
  NAND3_X2 u5_mult_82_U4361 ( .A1(u5_mult_82_n5702), .A2(u5_mult_82_n5703), 
        .A3(u5_mult_82_n5704), .ZN(u5_mult_82_CARRYB_12__33_) );
  BUF_X4 u5_mult_82_U4360 ( .A(u5_mult_82_SUMB_19__30_), .Z(u5_mult_82_n1760)
         );
  NAND2_X2 u5_mult_82_U4359 ( .A1(u5_mult_82_ab_51__34_), .A2(
        u5_mult_82_CARRYB_50__34_), .ZN(u5_mult_82_n2696) );
  NOR2_X2 u5_mult_82_U4358 ( .A1(u5_mult_82_net64881), .A2(u5_mult_82_net65225), .ZN(u5_mult_82_ab_50__34_) );
  NAND3_X4 u5_mult_82_U4357 ( .A1(u5_mult_82_n1056), .A2(u5_mult_82_n1057), 
        .A3(u5_mult_82_n1058), .ZN(u5_mult_82_CARRYB_50__34_) );
  NAND2_X1 u5_mult_82_U4356 ( .A1(u5_mult_82_ab_50__34_), .A2(
        u5_mult_82_CARRYB_49__34_), .ZN(u5_mult_82_n1058) );
  NAND2_X2 u5_mult_82_U4355 ( .A1(u5_mult_82_ab_50__34_), .A2(
        u5_mult_82_SUMB_49__35_), .ZN(u5_mult_82_n1057) );
  NAND2_X2 u5_mult_82_U4354 ( .A1(u5_mult_82_CARRYB_49__34_), .A2(
        u5_mult_82_SUMB_49__35_), .ZN(u5_mult_82_n1056) );
  XOR2_X2 u5_mult_82_U4353 ( .A(u5_mult_82_SUMB_49__35_), .B(u5_mult_82_n1055), 
        .Z(u5_mult_82_SUMB_50__34_) );
  XOR2_X1 u5_mult_82_U4352 ( .A(u5_mult_82_CARRYB_49__34_), .B(
        u5_mult_82_ab_50__34_), .Z(u5_mult_82_n1055) );
  INV_X1 u5_mult_82_U4351 ( .A(u5_mult_82_SUMB_50__35_), .ZN(u5_mult_82_n1052)
         );
  INV_X4 u5_mult_82_U4350 ( .A(u5_mult_82_n2135), .ZN(u5_mult_82_n1051) );
  NAND2_X2 u5_mult_82_U4349 ( .A1(u5_mult_82_n1051), .A2(u5_mult_82_n1052), 
        .ZN(u5_mult_82_n1054) );
  NAND2_X2 u5_mult_82_U4348 ( .A1(u5_mult_82_n2135), .A2(
        u5_mult_82_SUMB_50__35_), .ZN(u5_mult_82_n1053) );
  XNOR2_X1 u5_mult_82_U4347 ( .A(u5_mult_82_ab_1__30_), .B(
        u5_mult_82_ab_0__31_), .ZN(u5_mult_82_n6485) );
  NAND2_X2 u5_mult_82_U4346 ( .A1(u5_mult_82_ab_43__1_), .A2(
        u5_mult_82_SUMB_42__2_), .ZN(u5_mult_82_n2546) );
  NAND3_X2 u5_mult_82_U4345 ( .A1(u5_mult_82_n1048), .A2(u5_mult_82_n1049), 
        .A3(u5_mult_82_n1050), .ZN(u5_mult_82_CARRYB_43__41_) );
  NAND2_X1 u5_mult_82_U4344 ( .A1(u5_mult_82_ab_43__41_), .A2(
        u5_mult_82_CARRYB_42__41_), .ZN(u5_mult_82_n1050) );
  NAND2_X2 u5_mult_82_U4343 ( .A1(u5_mult_82_ab_43__41_), .A2(
        u5_mult_82_SUMB_42__42_), .ZN(u5_mult_82_n1049) );
  NAND2_X1 u5_mult_82_U4342 ( .A1(u5_mult_82_CARRYB_42__41_), .A2(
        u5_mult_82_SUMB_42__42_), .ZN(u5_mult_82_n1048) );
  XOR2_X2 u5_mult_82_U4341 ( .A(u5_mult_82_SUMB_42__42_), .B(u5_mult_82_n1047), 
        .Z(u5_mult_82_SUMB_43__41_) );
  XOR2_X2 u5_mult_82_U4340 ( .A(u5_mult_82_CARRYB_42__41_), .B(
        u5_mult_82_ab_43__41_), .Z(u5_mult_82_n1047) );
  NAND3_X2 u5_mult_82_U4339 ( .A1(u5_mult_82_n1044), .A2(u5_mult_82_n1045), 
        .A3(u5_mult_82_n1046), .ZN(u5_mult_82_CARRYB_11__49_) );
  NAND2_X2 u5_mult_82_U4338 ( .A1(u5_mult_82_CARRYB_10__49_), .A2(
        u5_mult_82_SUMB_10__50_), .ZN(u5_mult_82_n1046) );
  NAND2_X2 u5_mult_82_U4337 ( .A1(u5_mult_82_ab_11__49_), .A2(
        u5_mult_82_SUMB_10__50_), .ZN(u5_mult_82_n1045) );
  NAND2_X1 u5_mult_82_U4336 ( .A1(u5_mult_82_ab_11__49_), .A2(
        u5_mult_82_CARRYB_10__49_), .ZN(u5_mult_82_n1044) );
  NAND3_X2 u5_mult_82_U4335 ( .A1(u5_mult_82_n1041), .A2(u5_mult_82_n1042), 
        .A3(u5_mult_82_n1043), .ZN(u5_mult_82_CARRYB_10__50_) );
  NAND2_X2 u5_mult_82_U4334 ( .A1(u5_mult_82_ab_10__50_), .A2(
        u5_mult_82_SUMB_9__51_), .ZN(u5_mult_82_n1042) );
  XOR2_X2 u5_mult_82_U4333 ( .A(u5_mult_82_n1040), .B(u5_mult_82_SUMB_10__50_), 
        .Z(u5_mult_82_SUMB_11__49_) );
  XOR2_X2 u5_mult_82_U4332 ( .A(u5_mult_82_ab_11__49_), .B(
        u5_mult_82_CARRYB_10__49_), .Z(u5_mult_82_n1040) );
  XOR2_X2 u5_mult_82_U4331 ( .A(u5_mult_82_n1039), .B(u5_mult_82_SUMB_9__51_), 
        .Z(u5_mult_82_SUMB_10__50_) );
  NOR2_X1 u5_mult_82_U4330 ( .A1(u5_mult_82_net64455), .A2(u5_mult_82_n6567), 
        .ZN(u5_mult_82_ab_12__10_) );
  NAND3_X2 u5_mult_82_U4329 ( .A1(u5_mult_82_n1036), .A2(u5_mult_82_n1037), 
        .A3(u5_mult_82_n1038), .ZN(u5_mult_82_CARRYB_12__10_) );
  NAND2_X2 u5_mult_82_U4328 ( .A1(u5_mult_82_ab_12__10_), .A2(
        u5_mult_82_CARRYB_11__10_), .ZN(u5_mult_82_n1038) );
  NAND2_X2 u5_mult_82_U4327 ( .A1(u5_mult_82_ab_12__10_), .A2(
        u5_mult_82_SUMB_11__11_), .ZN(u5_mult_82_n1037) );
  NAND2_X1 u5_mult_82_U4326 ( .A1(u5_mult_82_CARRYB_11__10_), .A2(
        u5_mult_82_SUMB_11__11_), .ZN(u5_mult_82_n1036) );
  XOR2_X2 u5_mult_82_U4325 ( .A(u5_mult_82_SUMB_11__11_), .B(u5_mult_82_n1035), 
        .Z(u5_mult_82_SUMB_12__10_) );
  XOR2_X2 u5_mult_82_U4324 ( .A(u5_mult_82_CARRYB_11__10_), .B(
        u5_mult_82_ab_12__10_), .Z(u5_mult_82_n1035) );
  INV_X1 u5_mult_82_U4323 ( .A(u5_mult_82_CARRYB_40__2_), .ZN(u5_mult_82_n1032) );
  INV_X1 u5_mult_82_U4322 ( .A(u5_mult_82_ab_41__2_), .ZN(u5_mult_82_n1031) );
  NAND2_X2 u5_mult_82_U4321 ( .A1(u5_mult_82_n1031), .A2(u5_mult_82_n1032), 
        .ZN(u5_mult_82_n1034) );
  NAND2_X2 u5_mult_82_U4320 ( .A1(u5_mult_82_ab_41__2_), .A2(
        u5_mult_82_CARRYB_40__2_), .ZN(u5_mult_82_n1033) );
  NAND2_X1 u5_mult_82_U4319 ( .A1(u5_mult_82_ab_8__22_), .A2(
        u5_mult_82_SUMB_7__23_), .ZN(u5_mult_82_n3713) );
  NAND2_X2 u5_mult_82_U4318 ( .A1(u5_mult_82_n104), .A2(u5_mult_82_SUMB_6__25_), .ZN(u5_mult_82_n3822) );
  CLKBUF_X2 u5_mult_82_U4317 ( .A(u5_mult_82_SUMB_41__4_), .Z(u5_mult_82_n1531) );
  INV_X4 u5_mult_82_U4316 ( .A(u5_mult_82_n4640), .ZN(u5_mult_82_n1027) );
  NAND2_X4 u5_mult_82_U4315 ( .A1(u5_mult_82_n1029), .A2(u5_mult_82_n1030), 
        .ZN(u5_mult_82_SUMB_41__4_) );
  NAND2_X4 u5_mult_82_U4314 ( .A1(u5_mult_82_n1027), .A2(u5_mult_82_n1028), 
        .ZN(u5_mult_82_n1030) );
  NAND2_X2 u5_mult_82_U4313 ( .A1(u5_mult_82_n4640), .A2(
        u5_mult_82_SUMB_40__5_), .ZN(u5_mult_82_n1029) );
  NAND3_X2 u5_mult_82_U4312 ( .A1(u5_mult_82_n1024), .A2(u5_mult_82_n1025), 
        .A3(u5_mult_82_n1026), .ZN(u5_mult_82_CARRYB_16__12_) );
  NAND2_X1 u5_mult_82_U4311 ( .A1(u5_mult_82_CARRYB_15__12_), .A2(
        u5_mult_82_SUMB_15__13_), .ZN(u5_mult_82_n1026) );
  NAND2_X1 u5_mult_82_U4310 ( .A1(u5_mult_82_ab_16__12_), .A2(
        u5_mult_82_SUMB_15__13_), .ZN(u5_mult_82_n1025) );
  NAND2_X1 u5_mult_82_U4309 ( .A1(u5_mult_82_ab_16__12_), .A2(
        u5_mult_82_CARRYB_15__12_), .ZN(u5_mult_82_n1024) );
  NAND3_X2 u5_mult_82_U4308 ( .A1(u5_mult_82_n1021), .A2(u5_mult_82_n1022), 
        .A3(u5_mult_82_n1023), .ZN(u5_mult_82_CARRYB_15__13_) );
  NAND2_X2 u5_mult_82_U4307 ( .A1(u5_mult_82_CARRYB_14__13_), .A2(
        u5_mult_82_SUMB_14__14_), .ZN(u5_mult_82_n1023) );
  NAND2_X2 u5_mult_82_U4306 ( .A1(u5_mult_82_ab_15__13_), .A2(
        u5_mult_82_SUMB_14__14_), .ZN(u5_mult_82_n1022) );
  NAND2_X2 u5_mult_82_U4305 ( .A1(u5_mult_82_ab_15__13_), .A2(
        u5_mult_82_CARRYB_14__13_), .ZN(u5_mult_82_n1021) );
  XOR2_X2 u5_mult_82_U4304 ( .A(u5_mult_82_n1020), .B(u5_mult_82_SUMB_15__13_), 
        .Z(u5_mult_82_SUMB_16__12_) );
  XOR2_X2 u5_mult_82_U4303 ( .A(u5_mult_82_ab_16__12_), .B(
        u5_mult_82_CARRYB_15__12_), .Z(u5_mult_82_n1020) );
  XOR2_X2 u5_mult_82_U4302 ( .A(u5_mult_82_n1019), .B(u5_mult_82_SUMB_14__14_), 
        .Z(u5_mult_82_SUMB_15__13_) );
  XOR2_X1 u5_mult_82_U4301 ( .A(u5_mult_82_ab_15__13_), .B(
        u5_mult_82_CARRYB_14__13_), .Z(u5_mult_82_n1019) );
  NOR2_X2 u5_mult_82_U4300 ( .A1(u5_mult_82_net64961), .A2(u5_mult_82_net66107), .ZN(u5_mult_82_ab_1__38_) );
  XNOR2_X2 u5_mult_82_U4299 ( .A(u5_mult_82_ab_47__32_), .B(
        u5_mult_82_CARRYB_46__32_), .ZN(u5_mult_82_n1018) );
  XNOR2_X2 u5_mult_82_U4298 ( .A(u5_mult_82_n1018), .B(u5_mult_82_SUMB_46__33_), .ZN(u5_mult_82_SUMB_47__32_) );
  NAND2_X2 u5_mult_82_U4297 ( .A1(u5_mult_82_ab_27__25_), .A2(
        u5_mult_82_SUMB_26__26_), .ZN(u5_mult_82_n6184) );
  XNOR2_X2 u5_mult_82_U4296 ( .A(u5_mult_82_ab_17__31_), .B(
        u5_mult_82_SUMB_16__32_), .ZN(u5_mult_82_n1804) );
  XNOR2_X2 u5_mult_82_U4295 ( .A(u5_mult_82_ab_16__32_), .B(
        u5_mult_82_CARRYB_15__32_), .ZN(u5_mult_82_n3967) );
  XNOR2_X2 u5_mult_82_U4294 ( .A(u5_mult_82_CARRYB_23__27_), .B(
        u5_mult_82_n1491), .ZN(u5_mult_82_n6139) );
  CLKBUF_X3 u5_mult_82_U4293 ( .A(u5_mult_82_SUMB_44__29_), .Z(
        u5_mult_82_n1860) );
  NAND2_X4 u5_mult_82_U4292 ( .A1(u5_mult_82_ab_19__44_), .A2(u5_mult_82_n5248), .ZN(u5_mult_82_n5879) );
  CLKBUF_X2 u5_mult_82_U4291 ( .A(u5_mult_82_CARRYB_6__49_), .Z(
        u5_mult_82_n1765) );
  XOR2_X2 u5_mult_82_U4290 ( .A(u5_mult_82_n3924), .B(u5_mult_82_SUMB_35__35_), 
        .Z(u5_mult_82_SUMB_36__34_) );
  NAND2_X2 u5_mult_82_U4289 ( .A1(u5_mult_82_ab_7__24_), .A2(
        u5_mult_82_SUMB_6__25_), .ZN(u5_mult_82_n3821) );
  XOR2_X2 u5_mult_82_U4288 ( .A(u5_mult_82_ab_47__29_), .B(
        u5_mult_82_CARRYB_46__29_), .Z(u5_mult_82_n2438) );
  XNOR2_X2 u5_mult_82_U4287 ( .A(u5_mult_82_CARRYB_23__42_), .B(
        u5_mult_82_ab_24__42_), .ZN(u5_mult_82_n1677) );
  XOR2_X2 u5_mult_82_U4286 ( .A(u5_mult_82_ab_45__30_), .B(
        u5_mult_82_CARRYB_44__30_), .Z(u5_mult_82_n3020) );
  NAND2_X2 u5_mult_82_U4285 ( .A1(u5_mult_82_ab_18__36_), .A2(
        u5_mult_82_CARRYB_17__36_), .ZN(u5_mult_82_n5038) );
  NAND2_X2 u5_mult_82_U4284 ( .A1(u5_mult_82_CARRYB_25__15_), .A2(
        u5_mult_82_ab_26__15_), .ZN(u5_mult_82_n2994) );
  NOR2_X2 u5_mult_82_U4283 ( .A1(u5_mult_82_n6934), .A2(u5_mult_82_net65679), 
        .ZN(u5_mult_82_ab_25__15_) );
  NOR2_X1 u5_mult_82_U4282 ( .A1(u5_mult_82_n6882), .A2(u5_mult_82_n6529), 
        .ZN(u5_mult_82_ab_7__26_) );
  NAND2_X2 u5_mult_82_U4281 ( .A1(u5_mult_82_ab_13__23_), .A2(
        u5_mult_82_CARRYB_12__23_), .ZN(u5_mult_82_n3885) );
  NOR2_X1 u5_mult_82_U4280 ( .A1(u5_mult_82_net64689), .A2(u5_mult_82_n6566), 
        .ZN(u5_mult_82_ab_12__23_) );
  NAND2_X1 u5_mult_82_U4279 ( .A1(u5_mult_82_ab_25__15_), .A2(
        u5_mult_82_SUMB_24__16_), .ZN(u5_mult_82_n1016) );
  NAND2_X1 u5_mult_82_U4278 ( .A1(u5_mult_82_CARRYB_24__15_), .A2(
        u5_mult_82_SUMB_24__16_), .ZN(u5_mult_82_n1015) );
  NAND2_X1 u5_mult_82_U4277 ( .A1(u5_mult_82_ab_7__26_), .A2(
        u5_mult_82_CARRYB_6__26_), .ZN(u5_mult_82_n1014) );
  NAND2_X2 u5_mult_82_U4276 ( .A1(u5_mult_82_ab_7__26_), .A2(
        u5_mult_82_SUMB_6__27_), .ZN(u5_mult_82_n1013) );
  NAND2_X2 u5_mult_82_U4275 ( .A1(u5_mult_82_CARRYB_6__26_), .A2(
        u5_mult_82_SUMB_6__27_), .ZN(u5_mult_82_n1012) );
  XOR2_X2 u5_mult_82_U4274 ( .A(u5_mult_82_SUMB_6__27_), .B(u5_mult_82_n1011), 
        .Z(u5_mult_82_SUMB_7__26_) );
  XOR2_X2 u5_mult_82_U4273 ( .A(u5_mult_82_CARRYB_6__26_), .B(
        u5_mult_82_ab_7__26_), .Z(u5_mult_82_n1011) );
  INV_X1 u5_mult_82_U4272 ( .A(u5_mult_82_SUMB_16__20_), .ZN(u5_mult_82_n1008)
         );
  NAND2_X2 u5_mult_82_U4271 ( .A1(u5_mult_82_n1009), .A2(u5_mult_82_n1010), 
        .ZN(u5_mult_82_SUMB_17__19_) );
  NAND2_X1 u5_mult_82_U4270 ( .A1(u5_mult_82_n684), .A2(
        u5_mult_82_SUMB_16__20_), .ZN(u5_mult_82_n1010) );
  NAND3_X2 u5_mult_82_U4269 ( .A1(u5_mult_82_n1005), .A2(u5_mult_82_n1006), 
        .A3(u5_mult_82_n1007), .ZN(u5_mult_82_CARRYB_3__29_) );
  NAND2_X1 u5_mult_82_U4268 ( .A1(u5_mult_82_CARRYB_2__29_), .A2(
        u5_mult_82_SUMB_2__30_), .ZN(u5_mult_82_n1007) );
  NAND2_X1 u5_mult_82_U4267 ( .A1(u5_mult_82_ab_3__29_), .A2(
        u5_mult_82_SUMB_2__30_), .ZN(u5_mult_82_n1006) );
  NAND2_X1 u5_mult_82_U4266 ( .A1(u5_mult_82_ab_3__29_), .A2(
        u5_mult_82_CARRYB_2__29_), .ZN(u5_mult_82_n1005) );
  NAND3_X2 u5_mult_82_U4265 ( .A1(u5_mult_82_n1002), .A2(u5_mult_82_n1003), 
        .A3(u5_mult_82_n1004), .ZN(u5_mult_82_CARRYB_2__30_) );
  NAND2_X2 u5_mult_82_U4264 ( .A1(u5_mult_82_CARRYB_1__30_), .A2(
        u5_mult_82_SUMB_1__31_), .ZN(u5_mult_82_n1004) );
  NAND2_X2 u5_mult_82_U4263 ( .A1(u5_mult_82_ab_2__30_), .A2(
        u5_mult_82_SUMB_1__31_), .ZN(u5_mult_82_n1003) );
  NAND2_X1 u5_mult_82_U4262 ( .A1(u5_mult_82_ab_2__30_), .A2(
        u5_mult_82_CARRYB_1__30_), .ZN(u5_mult_82_n1002) );
  XOR2_X2 u5_mult_82_U4261 ( .A(u5_mult_82_n1001), .B(u5_mult_82_SUMB_2__30_), 
        .Z(u5_mult_82_SUMB_3__29_) );
  XOR2_X2 u5_mult_82_U4260 ( .A(u5_mult_82_ab_3__29_), .B(
        u5_mult_82_CARRYB_2__29_), .Z(u5_mult_82_n1001) );
  XOR2_X2 u5_mult_82_U4259 ( .A(u5_mult_82_n1000), .B(u5_mult_82_SUMB_1__31_), 
        .Z(u5_mult_82_SUMB_2__30_) );
  XOR2_X2 u5_mult_82_U4258 ( .A(u5_mult_82_ab_2__30_), .B(
        u5_mult_82_CARRYB_1__30_), .Z(u5_mult_82_n1000) );
  NAND3_X2 u5_mult_82_U4257 ( .A1(u5_mult_82_n997), .A2(u5_mult_82_n998), .A3(
        u5_mult_82_n999), .ZN(u5_mult_82_CARRYB_12__23_) );
  NAND2_X2 u5_mult_82_U4256 ( .A1(u5_mult_82_ab_12__23_), .A2(
        u5_mult_82_CARRYB_11__23_), .ZN(u5_mult_82_n999) );
  NAND2_X2 u5_mult_82_U4255 ( .A1(u5_mult_82_ab_12__23_), .A2(
        u5_mult_82_SUMB_11__24_), .ZN(u5_mult_82_n998) );
  NAND2_X1 u5_mult_82_U4254 ( .A1(u5_mult_82_CARRYB_11__23_), .A2(
        u5_mult_82_SUMB_11__24_), .ZN(u5_mult_82_n997) );
  XOR2_X2 u5_mult_82_U4253 ( .A(u5_mult_82_SUMB_11__24_), .B(u5_mult_82_n996), 
        .Z(u5_mult_82_SUMB_12__23_) );
  NAND3_X2 u5_mult_82_U4252 ( .A1(u5_mult_82_n993), .A2(u5_mult_82_n994), .A3(
        u5_mult_82_n995), .ZN(u5_mult_82_CARRYB_51__1_) );
  NAND2_X2 u5_mult_82_U4251 ( .A1(u5_mult_82_ab_51__1_), .A2(
        u5_mult_82_SUMB_50__2_), .ZN(u5_mult_82_n995) );
  NAND2_X1 u5_mult_82_U4250 ( .A1(u5_mult_82_CARRYB_50__1_), .A2(
        u5_mult_82_ab_51__1_), .ZN(u5_mult_82_n993) );
  NAND3_X2 u5_mult_82_U4249 ( .A1(u5_mult_82_n990), .A2(u5_mult_82_n991), .A3(
        u5_mult_82_n992), .ZN(u5_mult_82_CARRYB_50__2_) );
  NAND2_X2 u5_mult_82_U4248 ( .A1(u5_mult_82_ab_50__2_), .A2(
        u5_mult_82_SUMB_49__3_), .ZN(u5_mult_82_n992) );
  NAND2_X2 u5_mult_82_U4247 ( .A1(u5_mult_82_CARRYB_49__2_), .A2(
        u5_mult_82_SUMB_49__3_), .ZN(u5_mult_82_n991) );
  NAND2_X1 u5_mult_82_U4246 ( .A1(u5_mult_82_CARRYB_49__2_), .A2(
        u5_mult_82_ab_50__2_), .ZN(u5_mult_82_n990) );
  XOR2_X2 u5_mult_82_U4245 ( .A(u5_mult_82_n989), .B(u5_mult_82_n713), .Z(
        u5_mult_82_SUMB_50__2_) );
  NAND2_X1 u5_mult_82_U4244 ( .A1(u5_mult_82_ab_37__10_), .A2(
        u5_mult_82_SUMB_36__11_), .ZN(u5_mult_82_n987) );
  NAND2_X1 u5_mult_82_U4243 ( .A1(u5_mult_82_ab_37__10_), .A2(
        u5_mult_82_CARRYB_36__10_), .ZN(u5_mult_82_n986) );
  NAND3_X2 u5_mult_82_U4242 ( .A1(u5_mult_82_n983), .A2(u5_mult_82_n984), .A3(
        u5_mult_82_n985), .ZN(u5_mult_82_CARRYB_36__11_) );
  NAND2_X2 u5_mult_82_U4241 ( .A1(u5_mult_82_ab_36__11_), .A2(
        u5_mult_82_SUMB_35__12_), .ZN(u5_mult_82_n985) );
  NAND2_X2 u5_mult_82_U4240 ( .A1(u5_mult_82_CARRYB_35__11_), .A2(
        u5_mult_82_SUMB_35__12_), .ZN(u5_mult_82_n984) );
  NAND2_X1 u5_mult_82_U4239 ( .A1(u5_mult_82_CARRYB_35__11_), .A2(
        u5_mult_82_ab_36__11_), .ZN(u5_mult_82_n983) );
  XOR2_X2 u5_mult_82_U4238 ( .A(u5_mult_82_n982), .B(u5_mult_82_SUMB_36__11_), 
        .Z(u5_mult_82_SUMB_37__10_) );
  XOR2_X2 u5_mult_82_U4237 ( .A(u5_mult_82_n981), .B(u5_mult_82_SUMB_35__12_), 
        .Z(u5_mult_82_SUMB_36__11_) );
  XOR2_X2 u5_mult_82_U4236 ( .A(u5_mult_82_CARRYB_35__11_), .B(
        u5_mult_82_ab_36__11_), .Z(u5_mult_82_n981) );
  NAND3_X4 u5_mult_82_U4235 ( .A1(u5_mult_82_n6224), .A2(u5_mult_82_n6225), 
        .A3(u5_mult_82_n6226), .ZN(u5_mult_82_CARRYB_24__34_) );
  NAND2_X2 u5_mult_82_U4234 ( .A1(u5_mult_82_CARRYB_23__34_), .A2(
        u5_mult_82_SUMB_23__35_), .ZN(u5_mult_82_n6226) );
  NAND2_X2 u5_mult_82_U4233 ( .A1(u5_mult_82_ab_24__34_), .A2(
        u5_mult_82_SUMB_23__35_), .ZN(u5_mult_82_n6225) );
  NAND2_X1 u5_mult_82_U4232 ( .A1(u5_mult_82_ab_24__38_), .A2(
        u5_mult_82_CARRYB_23__38_), .ZN(u5_mult_82_n5848) );
  NAND2_X2 u5_mult_82_U4231 ( .A1(u5_mult_82_CARRYB_40__28_), .A2(
        u5_mult_82_SUMB_40__29_), .ZN(u5_mult_82_n5584) );
  NAND2_X2 u5_mult_82_U4230 ( .A1(u5_mult_82_ab_21__33_), .A2(
        u5_mult_82_SUMB_20__34_), .ZN(u5_mult_82_n4818) );
  NAND2_X2 u5_mult_82_U4229 ( .A1(u5_mult_82_ab_8__36_), .A2(
        u5_mult_82_CARRYB_7__36_), .ZN(u5_mult_82_n5621) );
  NAND3_X4 u5_mult_82_U4228 ( .A1(u5_mult_82_n6299), .A2(u5_mult_82_n6300), 
        .A3(u5_mult_82_n6301), .ZN(u5_mult_82_CARRYB_30__23_) );
  NAND2_X1 u5_mult_82_U4227 ( .A1(u5_mult_82_CARRYB_2__46_), .A2(
        u5_mult_82_SUMB_2__47_), .ZN(u5_mult_82_n1934) );
  NAND3_X2 u5_mult_82_U4226 ( .A1(u5_mult_82_n1932), .A2(u5_mult_82_n1933), 
        .A3(u5_mult_82_n1934), .ZN(u5_mult_82_CARRYB_3__46_) );
  NAND2_X1 u5_mult_82_U4225 ( .A1(u5_mult_82_SUMB_28__32_), .A2(
        u5_mult_82_CARRYB_28__31_), .ZN(u5_mult_82_n6120) );
  NAND2_X2 u5_mult_82_U4224 ( .A1(u5_mult_82_CARRYB_23__32_), .A2(
        u5_mult_82_n433), .ZN(u5_mult_82_n5509) );
  NAND2_X4 u5_mult_82_U4223 ( .A1(u5_mult_82_n3648), .A2(u5_mult_82_n3649), 
        .ZN(u5_mult_82_n3651) );
  NAND3_X2 u5_mult_82_U4222 ( .A1(u5_mult_82_n5084), .A2(u5_mult_82_n5085), 
        .A3(u5_mult_82_n5086), .ZN(u5_mult_82_CARRYB_36__35_) );
  BUF_X4 u5_mult_82_U4221 ( .A(u5_mult_82_CARRYB_17__46_), .Z(u5_mult_82_n1422) );
  NAND2_X2 u5_mult_82_U4220 ( .A1(u5_mult_82_CARRYB_25__43_), .A2(
        u5_mult_82_SUMB_25__44_), .ZN(u5_mult_82_n5594) );
  NAND2_X2 u5_mult_82_U4219 ( .A1(u5_mult_82_ab_33__31_), .A2(
        u5_mult_82_SUMB_32__32_), .ZN(u5_mult_82_n5947) );
  INV_X2 u5_mult_82_U4218 ( .A(u5_mult_82_CARRYB_19__32_), .ZN(
        u5_mult_82_n1126) );
  NAND3_X2 u5_mult_82_U4217 ( .A1(u5_mult_82_n5061), .A2(u5_mult_82_n5062), 
        .A3(u5_mult_82_n5063), .ZN(u5_mult_82_CARRYB_41__17_) );
  XNOR2_X2 u5_mult_82_U4216 ( .A(u5_mult_82_n4228), .B(u5_mult_82_n1750), .ZN(
        u5_mult_82_SUMB_42__19_) );
  XNOR2_X2 u5_mult_82_U4215 ( .A(u5_mult_82_CARRYB_25__34_), .B(
        u5_mult_82_ab_26__34_), .ZN(u5_mult_82_n980) );
  XNOR2_X2 u5_mult_82_U4214 ( .A(u5_mult_82_SUMB_25__35_), .B(u5_mult_82_n980), 
        .ZN(u5_mult_82_SUMB_26__34_) );
  NAND2_X2 u5_mult_82_U4213 ( .A1(u5_mult_82_CARRYB_9__45_), .A2(
        u5_mult_82_SUMB_9__46_), .ZN(u5_mult_82_n4801) );
  NAND3_X2 u5_mult_82_U4212 ( .A1(u5_mult_82_n4811), .A2(u5_mult_82_n4812), 
        .A3(u5_mult_82_n4813), .ZN(u5_mult_82_CARRYB_24__31_) );
  NAND2_X2 u5_mult_82_U4211 ( .A1(u5_mult_82_ab_26__43_), .A2(
        u5_mult_82_SUMB_25__44_), .ZN(u5_mult_82_n5593) );
  XOR2_X2 u5_mult_82_U4210 ( .A(u5_mult_82_n2438), .B(u5_mult_82_SUMB_46__30_), 
        .Z(u5_mult_82_SUMB_47__29_) );
  NAND2_X2 u5_mult_82_U4209 ( .A1(u5_mult_82_SUMB_8__47_), .A2(
        u5_mult_82_CARRYB_8__46_), .ZN(u5_mult_82_n4798) );
  XNOR2_X2 u5_mult_82_U4208 ( .A(u5_mult_82_n718), .B(u5_mult_82_ab_36__22_), 
        .ZN(u5_mult_82_n2410) );
  NAND2_X4 u5_mult_82_U4207 ( .A1(u5_mult_82_CARRYB_21__30_), .A2(
        u5_mult_82_n1791), .ZN(u5_mult_82_n3147) );
  NAND3_X4 u5_mult_82_U4206 ( .A1(u5_mult_82_n3145), .A2(u5_mult_82_n3146), 
        .A3(u5_mult_82_n3147), .ZN(u5_mult_82_CARRYB_22__30_) );
  NOR2_X4 u5_mult_82_U4205 ( .A1(u5_mult_82_n6844), .A2(u5_mult_82_n6642), 
        .ZN(u5_mult_82_ab_24__32_) );
  INV_X1 u5_mult_82_U4204 ( .A(u5_mult_82_ab_24__32_), .ZN(u5_mult_82_n977) );
  INV_X2 u5_mult_82_U4203 ( .A(u5_mult_82_CARRYB_23__32_), .ZN(u5_mult_82_n976) );
  NAND2_X2 u5_mult_82_U4202 ( .A1(u5_mult_82_n979), .A2(u5_mult_82_n978), .ZN(
        u5_mult_82_n3693) );
  NAND2_X2 u5_mult_82_U4201 ( .A1(u5_mult_82_n976), .A2(u5_mult_82_n977), .ZN(
        u5_mult_82_n979) );
  NAND2_X1 u5_mult_82_U4200 ( .A1(u5_mult_82_CARRYB_23__32_), .A2(
        u5_mult_82_ab_24__32_), .ZN(u5_mult_82_n978) );
  INV_X4 u5_mult_82_U4199 ( .A(u5_mult_82_n1521), .ZN(u5_mult_82_n1522) );
  NAND2_X2 u5_mult_82_U4198 ( .A1(u5_mult_82_ab_10__45_), .A2(
        u5_mult_82_SUMB_9__46_), .ZN(u5_mult_82_n4800) );
  NAND2_X1 u5_mult_82_U4197 ( .A1(u5_mult_82_ab_47__1_), .A2(
        u5_mult_82_CARRYB_46__1_), .ZN(u5_mult_82_n5810) );
  NAND2_X1 u5_mult_82_U4196 ( .A1(u5_mult_82_CARRYB_46__1_), .A2(
        u5_mult_82_SUMB_46__2_), .ZN(u5_mult_82_n5812) );
  NAND2_X2 u5_mult_82_U4195 ( .A1(u5_mult_82_n4789), .A2(
        u5_mult_82_SUMB_46__2_), .ZN(u5_mult_82_n4688) );
  NOR2_X2 u5_mult_82_U4194 ( .A1(u5_mult_82_n6840), .A2(u5_mult_82_n6514), 
        .ZN(u5_mult_82_ab_3__33_) );
  NAND2_X1 u5_mult_82_U4193 ( .A1(u5_mult_82_ab_3__33_), .A2(
        u5_mult_82_CARRYB_2__33_), .ZN(u5_mult_82_n975) );
  NAND2_X1 u5_mult_82_U4192 ( .A1(u5_mult_82_CARRYB_2__33_), .A2(
        u5_mult_82_SUMB_2__34_), .ZN(u5_mult_82_n973) );
  XOR2_X2 u5_mult_82_U4191 ( .A(u5_mult_82_SUMB_2__34_), .B(u5_mult_82_n972), 
        .Z(u5_mult_82_SUMB_3__33_) );
  XOR2_X2 u5_mult_82_U4190 ( .A(u5_mult_82_CARRYB_2__33_), .B(
        u5_mult_82_ab_3__33_), .Z(u5_mult_82_n972) );
  INV_X4 u5_mult_82_U4189 ( .A(u5_mult_82_CARRYB_20__22_), .ZN(u5_mult_82_n969) );
  INV_X2 u5_mult_82_U4188 ( .A(u5_mult_82_ab_21__22_), .ZN(u5_mult_82_n968) );
  NAND2_X2 u5_mult_82_U4187 ( .A1(u5_mult_82_n970), .A2(u5_mult_82_n971), .ZN(
        u5_mult_82_n2564) );
  NAND2_X2 u5_mult_82_U4186 ( .A1(u5_mult_82_n968), .A2(u5_mult_82_n969), .ZN(
        u5_mult_82_n971) );
  NAND2_X2 u5_mult_82_U4185 ( .A1(u5_mult_82_ab_17__48_), .A2(
        u5_mult_82_CARRYB_16__48_), .ZN(u5_mult_82_n4426) );
  NAND3_X2 u5_mult_82_U4184 ( .A1(u5_mult_82_n2999), .A2(u5_mult_82_n3000), 
        .A3(u5_mult_82_n3001), .ZN(u5_mult_82_CARRYB_47__37_) );
  NAND3_X4 u5_mult_82_U4183 ( .A1(u5_mult_82_n4336), .A2(u5_mult_82_n4337), 
        .A3(u5_mult_82_n4338), .ZN(u5_mult_82_CARRYB_10__49_) );
  XNOR2_X2 u5_mult_82_U4182 ( .A(u5_mult_82_CARRYB_20__5_), .B(
        u5_mult_82_ab_21__5_), .ZN(u5_mult_82_n967) );
  XNOR2_X2 u5_mult_82_U4181 ( .A(u5_mult_82_SUMB_20__6_), .B(u5_mult_82_n967), 
        .ZN(u5_mult_82_SUMB_21__5_) );
  NAND2_X2 u5_mult_82_U4180 ( .A1(u5_mult_82_CARRYB_41__21_), .A2(
        u5_mult_82_SUMB_41__22_), .ZN(u5_mult_82_n2253) );
  NAND3_X4 u5_mult_82_U4179 ( .A1(u5_mult_82_n5478), .A2(u5_mult_82_n5477), 
        .A3(u5_mult_82_n5479), .ZN(u5_mult_82_CARRYB_28__29_) );
  NAND2_X2 u5_mult_82_U4178 ( .A1(u5_mult_82_ab_20__34_), .A2(
        u5_mult_82_SUMB_19__35_), .ZN(u5_mult_82_n3113) );
  NAND2_X1 u5_mult_82_U4177 ( .A1(u5_mult_82_ab_36__29_), .A2(
        u5_mult_82_SUMB_35__30_), .ZN(u5_mult_82_n4875) );
  NOR2_X2 u5_mult_82_U4176 ( .A1(u5_mult_82_net64217), .A2(u5_mult_82_n6772), 
        .ZN(u5_mult_82_ab_0__49_) );
  NAND2_X2 u5_mult_82_U4175 ( .A1(u5_mult_82_ab_0__49_), .A2(
        u5_mult_82_ab_1__48_), .ZN(u5_mult_82_n6506) );
  XNOR2_X2 u5_mult_82_U4174 ( .A(u5_mult_82_ab_10__45_), .B(
        u5_mult_82_CARRYB_9__45_), .ZN(u5_mult_82_n1709) );
  NAND2_X2 u5_mult_82_U4173 ( .A1(u5_mult_82_n3510), .A2(
        u5_mult_82_SUMB_17__37_), .ZN(u5_mult_82_n3233) );
  INV_X2 u5_mult_82_U4172 ( .A(u5_mult_82_SUMB_17__37_), .ZN(u5_mult_82_n3232)
         );
  NAND2_X2 u5_mult_82_U4171 ( .A1(u5_mult_82_ab_18__36_), .A2(
        u5_mult_82_SUMB_17__37_), .ZN(u5_mult_82_n5039) );
  NAND2_X2 u5_mult_82_U4170 ( .A1(u5_mult_82_ab_42__2_), .A2(
        u5_mult_82_SUMB_41__3_), .ZN(u5_mult_82_n5632) );
  NAND3_X4 u5_mult_82_U4169 ( .A1(u5_mult_82_n5165), .A2(u5_mult_82_n5166), 
        .A3(u5_mult_82_n5167), .ZN(u5_mult_82_CARRYB_8__45_) );
  NAND2_X1 u5_mult_82_U4168 ( .A1(u5_mult_82_CARRYB_22__38_), .A2(
        u5_mult_82_SUMB_22__39_), .ZN(u5_mult_82_n6002) );
  NAND2_X1 u5_mult_82_U4167 ( .A1(u5_mult_82_ab_23__38_), .A2(
        u5_mult_82_CARRYB_22__38_), .ZN(u5_mult_82_n6000) );
  NOR2_X2 u5_mult_82_U4166 ( .A1(u5_mult_82_n966), .A2(u5_mult_82_n6979), .ZN(
        u5_mult_82_n965) );
  INV_X1 u5_mult_82_U4165 ( .A(u5_mult_82_n5506), .ZN(u5_mult_82_n5507) );
  INV_X8 u5_mult_82_U4164 ( .A(u5_mult_82_n6984), .ZN(u5_mult_82_n6981) );
  NOR2_X4 u5_mult_82_U4163 ( .A1(u5_mult_82_n7010), .A2(u5_mult_82_n2133), 
        .ZN(u5_mult_82_n2132) );
  XNOR2_X2 u5_mult_82_U4162 ( .A(u5_mult_82_n1420), .B(u5_mult_82_n730), .ZN(
        u5_mult_82_n3844) );
  NAND2_X2 u5_mult_82_U4161 ( .A1(u5_mult_82_ab_20__34_), .A2(
        u5_mult_82_CARRYB_19__34_), .ZN(u5_mult_82_n3112) );
  NAND2_X1 u5_mult_82_U4160 ( .A1(u5_mult_82_ab_16__37_), .A2(
        u5_mult_82_CARRYB_15__37_), .ZN(u5_mult_82_n6307) );
  NOR2_X2 u5_mult_82_U4159 ( .A1(u5_mult_82_net64941), .A2(u5_mult_82_n6586), 
        .ZN(u5_mult_82_ab_15__37_) );
  NAND3_X2 u5_mult_82_U4158 ( .A1(u5_mult_82_n962), .A2(u5_mult_82_n964), .A3(
        u5_mult_82_n963), .ZN(u5_mult_82_CARRYB_15__37_) );
  NAND2_X1 u5_mult_82_U4157 ( .A1(u5_mult_82_ab_15__37_), .A2(
        u5_mult_82_CARRYB_14__37_), .ZN(u5_mult_82_n964) );
  NAND2_X1 u5_mult_82_U4156 ( .A1(u5_mult_82_CARRYB_14__37_), .A2(
        u5_mult_82_SUMB_14__38_), .ZN(u5_mult_82_n962) );
  XOR2_X2 u5_mult_82_U4155 ( .A(u5_mult_82_CARRYB_14__37_), .B(
        u5_mult_82_ab_15__37_), .Z(u5_mult_82_n961) );
  XNOR2_X2 u5_mult_82_U4154 ( .A(u5_mult_82_CARRYB_13__39_), .B(
        u5_mult_82_n960), .ZN(u5_mult_82_n5351) );
  NAND2_X1 u5_mult_82_U4153 ( .A1(u5_mult_82_CARRYB_35__13_), .A2(
        u5_mult_82_SUMB_35__14_), .ZN(u5_mult_82_n1996) );
  INV_X8 u5_mult_82_U4152 ( .A(u5_mult_82_n5183), .ZN(u5_mult_82_n5184) );
  NAND2_X1 u5_mult_82_U4151 ( .A1(u5_mult_82_CARRYB_5__42_), .A2(
        u5_mult_82_SUMB_5__43_), .ZN(u5_mult_82_n5985) );
  NAND2_X2 u5_mult_82_U4150 ( .A1(u5_mult_82_SUMB_6__42_), .A2(
        u5_mult_82_n1510), .ZN(u5_mult_82_n6020) );
  NAND2_X1 u5_mult_82_U4149 ( .A1(u5_mult_82_ab_16__36_), .A2(
        u5_mult_82_CARRYB_15__36_), .ZN(u5_mult_82_n6187) );
  NAND3_X2 u5_mult_82_U4148 ( .A1(u5_mult_82_n5985), .A2(u5_mult_82_n5986), 
        .A3(u5_mult_82_n5987), .ZN(u5_mult_82_CARRYB_6__42_) );
  NAND2_X1 u5_mult_82_U4147 ( .A1(u5_mult_82_ab_6__42_), .A2(
        u5_mult_82_SUMB_5__43_), .ZN(u5_mult_82_n5986) );
  NAND2_X2 u5_mult_82_U4146 ( .A1(u5_mult_82_ab_17__31_), .A2(
        u5_mult_82_SUMB_16__32_), .ZN(u5_mult_82_n5914) );
  NAND2_X2 u5_mult_82_U4145 ( .A1(u5_mult_82_ab_1__51_), .A2(
        u5_mult_82_net64225), .ZN(u5_mult_82_n966) );
  NAND2_X2 u5_mult_82_U4144 ( .A1(u5_mult_82_CARRYB_41__9_), .A2(
        u5_mult_82_SUMB_41__10_), .ZN(u5_mult_82_n6131) );
  NAND2_X2 u5_mult_82_U4143 ( .A1(u5_mult_82_n2744), .A2(u5_mult_82_n4218), 
        .ZN(u5_mult_82_n2747) );
  OAI21_X2 u5_mult_82_U4142 ( .B1(u5_mult_82_n1255), .B2(u5_mult_82_n1254), 
        .A(u5_mult_82_n613), .ZN(u5_mult_82_n1260) );
  NAND3_X4 u5_mult_82_U4141 ( .A1(u5_mult_82_net79215), .A2(
        u5_mult_82_net79214), .A3(u5_mult_82_net79213), .ZN(
        u5_mult_82_CARRYB_30__19_) );
  NAND2_X2 u5_mult_82_U4140 ( .A1(u5_mult_82_n5254), .A2(u5_mult_82_n5255), 
        .ZN(u5_mult_82_SUMB_18__46_) );
  NAND2_X1 u5_mult_82_U4139 ( .A1(u5_mult_82_ab_47__37_), .A2(
        u5_mult_82_SUMB_46__38_), .ZN(u5_mult_82_n3000) );
  NAND2_X2 u5_mult_82_U4138 ( .A1(u5_mult_82_ab_40__0_), .A2(
        u5_mult_82_CARRYB_39__0_), .ZN(u5_mult_82_n4851) );
  NAND2_X2 u5_mult_82_U4137 ( .A1(u5_mult_82_CARRYB_27__35_), .A2(
        u5_mult_82_n2320), .ZN(u5_mult_82_n3118) );
  NAND3_X2 u5_mult_82_U4136 ( .A1(u5_mult_82_n5395), .A2(u5_mult_82_n5396), 
        .A3(u5_mult_82_n5397), .ZN(u5_mult_82_CARRYB_11__43_) );
  NAND3_X4 u5_mult_82_U4135 ( .A1(u5_mult_82_n5391), .A2(u5_mult_82_n5392), 
        .A3(u5_mult_82_n5393), .ZN(u5_mult_82_CARRYB_10__43_) );
  NAND2_X2 u5_mult_82_U4134 ( .A1(u5_mult_82_CARRYB_9__43_), .A2(
        u5_mult_82_SUMB_9__44_), .ZN(u5_mult_82_n5393) );
  NAND2_X4 u5_mult_82_U4133 ( .A1(u5_mult_82_n5184), .A2(
        u5_mult_82_CARRYB_11__38_), .ZN(u5_mult_82_n6091) );
  XNOR2_X2 u5_mult_82_U4132 ( .A(u5_mult_82_n1771), .B(u5_mult_82_n2419), .ZN(
        u5_mult_82_SUMB_4__47_) );
  NAND2_X2 u5_mult_82_U4131 ( .A1(u5_mult_82_ab_33__39_), .A2(
        u5_mult_82_CARRYB_32__39_), .ZN(u5_mult_82_n3840) );
  NAND2_X2 u5_mult_82_U4130 ( .A1(u5_mult_82_CARRYB_34__13_), .A2(
        u5_mult_82_SUMB_34__14_), .ZN(u5_mult_82_n4956) );
  NAND2_X1 u5_mult_82_U4129 ( .A1(u5_mult_82_CARRYB_37__35_), .A2(
        u5_mult_82_SUMB_37__36_), .ZN(u5_mult_82_n3934) );
  NAND2_X2 u5_mult_82_U4128 ( .A1(u5_mult_82_CARRYB_39__39_), .A2(
        u5_mult_82_SUMB_39__40_), .ZN(u5_mult_82_n3371) );
  NAND2_X2 u5_mult_82_U4127 ( .A1(u5_mult_82_ab_40__39_), .A2(
        u5_mult_82_CARRYB_39__39_), .ZN(u5_mult_82_n3373) );
  NOR2_X1 u5_mult_82_U4126 ( .A1(u5_mult_82_n6832), .A2(u5_mult_82_n6727), 
        .ZN(u5_mult_82_ab_39__39_) );
  NAND2_X1 u5_mult_82_U4125 ( .A1(u5_mult_82_ab_39__39_), .A2(
        u5_mult_82_CARRYB_38__39_), .ZN(u5_mult_82_n959) );
  NAND2_X2 u5_mult_82_U4124 ( .A1(u5_mult_82_ab_39__39_), .A2(
        u5_mult_82_SUMB_38__40_), .ZN(u5_mult_82_n958) );
  NAND2_X2 u5_mult_82_U4123 ( .A1(u5_mult_82_CARRYB_38__39_), .A2(
        u5_mult_82_SUMB_38__40_), .ZN(u5_mult_82_n957) );
  XOR2_X2 u5_mult_82_U4122 ( .A(u5_mult_82_SUMB_38__40_), .B(u5_mult_82_n956), 
        .Z(u5_mult_82_SUMB_39__39_) );
  XOR2_X2 u5_mult_82_U4121 ( .A(u5_mult_82_CARRYB_38__39_), .B(
        u5_mult_82_ab_39__39_), .Z(u5_mult_82_n956) );
  NAND3_X2 u5_mult_82_U4120 ( .A1(u5_mult_82_n953), .A2(u5_mult_82_n954), .A3(
        u5_mult_82_n955), .ZN(u5_mult_82_CARRYB_41__37_) );
  NAND2_X2 u5_mult_82_U4119 ( .A1(u5_mult_82_ab_41__37_), .A2(
        u5_mult_82_SUMB_40__38_), .ZN(u5_mult_82_n954) );
  NAND2_X1 u5_mult_82_U4118 ( .A1(u5_mult_82_ab_41__37_), .A2(
        u5_mult_82_CARRYB_40__37_), .ZN(u5_mult_82_n953) );
  NAND3_X4 u5_mult_82_U4117 ( .A1(u5_mult_82_n950), .A2(u5_mult_82_n951), .A3(
        u5_mult_82_n952), .ZN(u5_mult_82_CARRYB_40__38_) );
  NAND2_X1 u5_mult_82_U4116 ( .A1(u5_mult_82_CARRYB_39__38_), .A2(
        u5_mult_82_SUMB_39__39_), .ZN(u5_mult_82_n952) );
  NAND2_X2 u5_mult_82_U4115 ( .A1(u5_mult_82_ab_40__38_), .A2(
        u5_mult_82_SUMB_39__39_), .ZN(u5_mult_82_n951) );
  NAND2_X2 u5_mult_82_U4114 ( .A1(u5_mult_82_ab_40__38_), .A2(
        u5_mult_82_CARRYB_39__38_), .ZN(u5_mult_82_n950) );
  XOR2_X2 u5_mult_82_U4113 ( .A(u5_mult_82_n949), .B(u5_mult_82_SUMB_40__38_), 
        .Z(u5_mult_82_SUMB_41__37_) );
  XOR2_X2 u5_mult_82_U4112 ( .A(u5_mult_82_ab_41__37_), .B(
        u5_mult_82_CARRYB_40__37_), .Z(u5_mult_82_n949) );
  XOR2_X2 u5_mult_82_U4111 ( .A(u5_mult_82_n948), .B(u5_mult_82_SUMB_39__39_), 
        .Z(u5_mult_82_SUMB_40__38_) );
  XOR2_X2 u5_mult_82_U4110 ( .A(u5_mult_82_ab_40__38_), .B(
        u5_mult_82_CARRYB_39__38_), .Z(u5_mult_82_n948) );
  NAND2_X2 u5_mult_82_U4109 ( .A1(u5_mult_82_CARRYB_19__23_), .A2(
        u5_mult_82_SUMB_19__24_), .ZN(u5_mult_82_n5496) );
  NAND2_X2 u5_mult_82_U4108 ( .A1(u5_mult_82_ab_30__30_), .A2(
        u5_mult_82_CARRYB_29__30_), .ZN(u5_mult_82_n6121) );
  XNOR2_X2 u5_mult_82_U4107 ( .A(u5_mult_82_ab_13__31_), .B(
        u5_mult_82_CARRYB_12__31_), .ZN(u5_mult_82_n947) );
  XNOR2_X2 u5_mult_82_U4106 ( .A(u5_mult_82_n947), .B(u5_mult_82_SUMB_12__32_), 
        .ZN(u5_mult_82_SUMB_13__31_) );
  NAND3_X4 u5_mult_82_U4105 ( .A1(u5_mult_82_net80188), .A2(u5_mult_82_n5383), 
        .A3(u5_mult_82_net80190), .ZN(u5_mult_82_CARRYB_8__34_) );
  NAND2_X2 u5_mult_82_U4104 ( .A1(u5_mult_82_ab_40__32_), .A2(
        u5_mult_82_SUMB_39__33_), .ZN(u5_mult_82_n5112) );
  NAND2_X2 u5_mult_82_U4103 ( .A1(u5_mult_82_CARRYB_35__35_), .A2(
        u5_mult_82_SUMB_35__36_), .ZN(u5_mult_82_n5086) );
  NAND2_X2 u5_mult_82_U4102 ( .A1(u5_mult_82_CARRYB_2__40_), .A2(
        u5_mult_82_SUMB_2__41_), .ZN(u5_mult_82_n5502) );
  NAND2_X2 u5_mult_82_U4101 ( .A1(u5_mult_82_CARRYB_10__38_), .A2(
        u5_mult_82_SUMB_10__39_), .ZN(u5_mult_82_n3641) );
  NAND2_X2 u5_mult_82_U4100 ( .A1(u5_mult_82_ab_42__21_), .A2(
        u5_mult_82_SUMB_41__22_), .ZN(u5_mult_82_n2252) );
  XOR2_X2 u5_mult_82_U4099 ( .A(u5_mult_82_SUMB_27__7_), .B(u5_mult_82_n2062), 
        .Z(u5_mult_82_SUMB_28__6_) );
  NAND3_X2 u5_mult_82_U4098 ( .A1(u5_mult_82_n6079), .A2(u5_mult_82_n6078), 
        .A3(u5_mult_82_n6077), .ZN(u5_mult_82_CARRYB_27__23_) );
  NAND2_X2 u5_mult_82_U4097 ( .A1(u5_mult_82_ab_40__12_), .A2(
        u5_mult_82_SUMB_39__13_), .ZN(u5_mult_82_net82471) );
  INV_X4 u5_mult_82_U4096 ( .A(u5_mult_82_n1576), .ZN(u5_mult_82_n1577) );
  XNOR2_X2 u5_mult_82_U4095 ( .A(u5_mult_82_SUMB_23__38_), .B(
        u5_mult_82_ab_24__37_), .ZN(u5_mult_82_n1406) );
  NAND2_X2 u5_mult_82_U4094 ( .A1(u5_mult_82_ab_35__13_), .A2(
        u5_mult_82_SUMB_34__14_), .ZN(u5_mult_82_n4955) );
  INV_X4 u5_mult_82_U4093 ( .A(u5_mult_82_n6391), .ZN(u5_mult_82_CLA_SUM[55])
         );
  XOR2_X2 u5_mult_82_U4092 ( .A(u5_mult_82_CARRYB_8__42_), .B(u5_mult_82_n2361), .Z(u5_mult_82_n946) );
  XNOR2_X2 u5_mult_82_U4091 ( .A(u5_mult_82_SUMB_8__43_), .B(u5_mult_82_n946), 
        .ZN(u5_mult_82_SUMB_9__42_) );
  NAND2_X1 u5_mult_82_U4090 ( .A1(u5_mult_82_ab_29__31_), .A2(
        u5_mult_82_SUMB_28__32_), .ZN(u5_mult_82_n6119) );
  BUF_X8 u5_mult_82_U4089 ( .A(u5_mult_82_CARRYB_45__31_), .Z(u5_mult_82_n1566) );
  XNOR2_X2 u5_mult_82_U4088 ( .A(u5_mult_82_CARRYB_47__29_), .B(
        u5_mult_82_ab_48__29_), .ZN(u5_mult_82_n945) );
  XNOR2_X2 u5_mult_82_U4087 ( .A(u5_mult_82_n1826), .B(u5_mult_82_n945), .ZN(
        u5_mult_82_SUMB_48__29_) );
  NAND2_X1 u5_mult_82_U4086 ( .A1(u5_mult_82_ab_25__33_), .A2(
        u5_mult_82_CARRYB_24__33_), .ZN(u5_mult_82_n6227) );
  NAND2_X2 u5_mult_82_U4085 ( .A1(u5_mult_82_CARRYB_38__34_), .A2(
        u5_mult_82_SUMB_38__35_), .ZN(u5_mult_82_n3937) );
  XNOR2_X1 u5_mult_82_U4084 ( .A(u5_mult_82_CARRYB_11__33_), .B(
        u5_mult_82_ab_12__33_), .ZN(u5_mult_82_n944) );
  NAND3_X2 u5_mult_82_U4083 ( .A1(u5_mult_82_n2427), .A2(u5_mult_82_n2428), 
        .A3(u5_mult_82_n2429), .ZN(u5_mult_82_CARRYB_29__32_) );
  NAND2_X2 u5_mult_82_U4082 ( .A1(u5_mult_82_CARRYB_10__42_), .A2(
        u5_mult_82_SUMB_10__43_), .ZN(u5_mult_82_n5367) );
  NAND2_X2 u5_mult_82_U4081 ( .A1(u5_mult_82_CARRYB_4__45_), .A2(
        u5_mult_82_SUMB_4__46_), .ZN(u5_mult_82_n4995) );
  INV_X2 u5_mult_82_U4080 ( .A(u5_mult_82_SUMB_31__31_), .ZN(u5_mult_82_n5561)
         );
  NAND2_X2 u5_mult_82_U4079 ( .A1(u5_mult_82_ab_26__33_), .A2(
        u5_mult_82_SUMB_25__34_), .ZN(u5_mult_82_n5768) );
  NAND2_X1 u5_mult_82_U4078 ( .A1(u5_mult_82_CARRYB_31__40_), .A2(
        u5_mult_82_SUMB_31__41_), .ZN(u5_mult_82_n3839) );
  INV_X4 u5_mult_82_U4077 ( .A(u5_mult_82_n6389), .ZN(u5_mult_82_CLA_CARRY[53]) );
  NAND2_X2 u5_mult_82_U4076 ( .A1(u5_mult_82_ab_50__6_), .A2(
        u5_mult_82_SUMB_49__7_), .ZN(u5_mult_82_net78901) );
  NOR2_X2 u5_mult_82_U4075 ( .A1(u5_mult_82_n6797), .A2(u5_mult_82_net65349), 
        .ZN(u5_mult_82_ab_43__45_) );
  NOR2_X2 u5_mult_82_U4074 ( .A1(u5_mult_82_n6797), .A2(u5_mult_82_net65375), 
        .ZN(u5_mult_82_ab_42__45_) );
  NAND3_X4 u5_mult_82_U4073 ( .A1(u5_mult_82_n4799), .A2(u5_mult_82_n4801), 
        .A3(u5_mult_82_n4800), .ZN(u5_mult_82_CARRYB_10__45_) );
  NAND3_X4 u5_mult_82_U4072 ( .A1(u5_mult_82_n3134), .A2(u5_mult_82_n3135), 
        .A3(u5_mult_82_n3136), .ZN(u5_mult_82_CARRYB_16__41_) );
  NOR2_X1 u5_mult_82_U4071 ( .A1(u5_mult_82_n6822), .A2(u5_mult_82_n6600), 
        .ZN(u5_mult_82_ab_17__41_) );
  NAND3_X2 u5_mult_82_U4070 ( .A1(u5_mult_82_n941), .A2(u5_mult_82_n942), .A3(
        u5_mult_82_n943), .ZN(u5_mult_82_CARRYB_17__41_) );
  NAND2_X1 u5_mult_82_U4069 ( .A1(u5_mult_82_ab_17__41_), .A2(
        u5_mult_82_CARRYB_16__41_), .ZN(u5_mult_82_n943) );
  NAND2_X2 u5_mult_82_U4068 ( .A1(u5_mult_82_ab_17__41_), .A2(
        u5_mult_82_SUMB_16__42_), .ZN(u5_mult_82_n942) );
  NAND2_X2 u5_mult_82_U4067 ( .A1(u5_mult_82_CARRYB_16__41_), .A2(
        u5_mult_82_SUMB_16__42_), .ZN(u5_mult_82_n941) );
  XOR2_X2 u5_mult_82_U4066 ( .A(u5_mult_82_SUMB_16__42_), .B(u5_mult_82_n940), 
        .Z(u5_mult_82_SUMB_17__41_) );
  NAND3_X4 u5_mult_82_U4065 ( .A1(u5_mult_82_n937), .A2(u5_mult_82_n938), .A3(
        u5_mult_82_n939), .ZN(u5_mult_82_CARRYB_12__44_) );
  NAND2_X2 u5_mult_82_U4064 ( .A1(u5_mult_82_ab_12__44_), .A2(
        u5_mult_82_SUMB_11__45_), .ZN(u5_mult_82_n938) );
  NAND2_X1 u5_mult_82_U4063 ( .A1(u5_mult_82_ab_12__44_), .A2(u5_mult_82_n762), 
        .ZN(u5_mult_82_n937) );
  NAND3_X2 u5_mult_82_U4062 ( .A1(u5_mult_82_n934), .A2(u5_mult_82_n935), .A3(
        u5_mult_82_n936), .ZN(u5_mult_82_CARRYB_11__45_) );
  NAND2_X1 u5_mult_82_U4061 ( .A1(u5_mult_82_CARRYB_10__45_), .A2(
        u5_mult_82_SUMB_10__46_), .ZN(u5_mult_82_n936) );
  NAND2_X1 u5_mult_82_U4060 ( .A1(u5_mult_82_ab_11__45_), .A2(
        u5_mult_82_SUMB_10__46_), .ZN(u5_mult_82_n935) );
  NAND2_X1 u5_mult_82_U4059 ( .A1(u5_mult_82_ab_11__45_), .A2(
        u5_mult_82_CARRYB_10__45_), .ZN(u5_mult_82_n934) );
  XOR2_X2 u5_mult_82_U4058 ( .A(u5_mult_82_n933), .B(u5_mult_82_SUMB_10__46_), 
        .Z(u5_mult_82_SUMB_11__45_) );
  XOR2_X2 u5_mult_82_U4057 ( .A(u5_mult_82_ab_11__45_), .B(
        u5_mult_82_CARRYB_10__45_), .Z(u5_mult_82_n933) );
  NAND2_X2 u5_mult_82_U4056 ( .A1(u5_mult_82_ab_39__14_), .A2(
        u5_mult_82_SUMB_38__15_), .ZN(u5_mult_82_n3883) );
  XNOR2_X2 u5_mult_82_U4055 ( .A(u5_mult_82_ab_41__10_), .B(
        u5_mult_82_CARRYB_40__10_), .ZN(u5_mult_82_n1471) );
  XNOR2_X2 u5_mult_82_U4054 ( .A(u5_mult_82_n5394), .B(
        u5_mult_82_CARRYB_10__43_), .ZN(u5_mult_82_n932) );
  NAND2_X2 u5_mult_82_U4053 ( .A1(u5_mult_82_SUMB_32__32_), .A2(
        u5_mult_82_CARRYB_32__31_), .ZN(u5_mult_82_n5948) );
  NAND2_X2 u5_mult_82_U4052 ( .A1(u5_mult_82_SUMB_23__38_), .A2(
        u5_mult_82_CARRYB_23__37_), .ZN(u5_mult_82_n5558) );
  XNOR2_X1 u5_mult_82_U4051 ( .A(u5_mult_82_CARRYB_31__32_), .B(
        u5_mult_82_ab_32__32_), .ZN(u5_mult_82_n1731) );
  NOR2_X4 u5_mult_82_U4050 ( .A1(u5_mult_82_n6979), .A2(u5_mult_82_net64223), 
        .ZN(u5_mult_82_n2124) );
  INV_X16 u5_mult_82_U4049 ( .A(u5_mult_82_n6802), .ZN(u5_mult_82_n6797) );
  INV_X1 u5_mult_82_U4048 ( .A(u5_mult_82_n7008), .ZN(u5_mult_82_n6802) );
  XNOR2_X2 u5_mult_82_U4047 ( .A(u5_mult_82_ab_1__46_), .B(
        u5_mult_82_ab_0__47_), .ZN(u5_mult_82_n6503) );
  XNOR2_X2 u5_mult_82_U4046 ( .A(u5_mult_82_ab_37__35_), .B(
        u5_mult_82_CARRYB_36__35_), .ZN(u5_mult_82_n931) );
  XNOR2_X2 u5_mult_82_U4045 ( .A(u5_mult_82_ab_25__19_), .B(
        u5_mult_82_CARRYB_24__19_), .ZN(u5_mult_82_n930) );
  XNOR2_X1 u5_mult_82_U4044 ( .A(u5_mult_82_CARRYB_15__19_), .B(
        u5_mult_82_ab_16__19_), .ZN(u5_mult_82_n929) );
  XNOR2_X2 u5_mult_82_U4043 ( .A(u5_mult_82_n929), .B(u5_mult_82_n1829), .ZN(
        u5_mult_82_SUMB_16__19_) );
  NOR2_X1 u5_mult_82_U4042 ( .A1(u5_mult_82_n6822), .A2(u5_mult_82_n6655), 
        .ZN(u5_mult_82_ab_27__41_) );
  NOR2_X1 u5_mult_82_U4041 ( .A1(u5_mult_82_net64903), .A2(u5_mult_82_net65405), .ZN(u5_mult_82_ab_40__35_) );
  NAND3_X4 u5_mult_82_U4040 ( .A1(u5_mult_82_n5121), .A2(u5_mult_82_n5122), 
        .A3(u5_mult_82_n5123), .ZN(u5_mult_82_CARRYB_36__36_) );
  NOR2_X1 u5_mult_82_U4039 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6720), 
        .ZN(u5_mult_82_ab_37__36_) );
  NAND2_X2 u5_mult_82_U4038 ( .A1(u5_mult_82_ab_27__41_), .A2(
        u5_mult_82_SUMB_26__42_), .ZN(u5_mult_82_n927) );
  XOR2_X2 u5_mult_82_U4037 ( .A(u5_mult_82_SUMB_26__42_), .B(u5_mult_82_n925), 
        .Z(u5_mult_82_SUMB_27__41_) );
  XOR2_X2 u5_mult_82_U4036 ( .A(u5_mult_82_CARRYB_26__41_), .B(
        u5_mult_82_ab_27__41_), .Z(u5_mult_82_n925) );
  NAND3_X2 u5_mult_82_U4035 ( .A1(u5_mult_82_n922), .A2(u5_mult_82_n923), .A3(
        u5_mult_82_n924), .ZN(u5_mult_82_CARRYB_40__35_) );
  NAND2_X1 u5_mult_82_U4034 ( .A1(u5_mult_82_ab_40__35_), .A2(
        u5_mult_82_SUMB_39__36_), .ZN(u5_mult_82_n924) );
  NAND2_X2 u5_mult_82_U4033 ( .A1(u5_mult_82_ab_40__35_), .A2(
        u5_mult_82_CARRYB_39__35_), .ZN(u5_mult_82_n923) );
  NAND2_X1 u5_mult_82_U4032 ( .A1(u5_mult_82_SUMB_39__36_), .A2(
        u5_mult_82_CARRYB_39__35_), .ZN(u5_mult_82_n922) );
  XOR2_X2 u5_mult_82_U4031 ( .A(u5_mult_82_CARRYB_39__35_), .B(u5_mult_82_n921), .Z(u5_mult_82_SUMB_40__35_) );
  XOR2_X2 u5_mult_82_U4030 ( .A(u5_mult_82_SUMB_39__36_), .B(
        u5_mult_82_ab_40__35_), .Z(u5_mult_82_n921) );
  NAND3_X2 u5_mult_82_U4029 ( .A1(u5_mult_82_n918), .A2(u5_mult_82_n919), .A3(
        u5_mult_82_n920), .ZN(u5_mult_82_CARRYB_37__36_) );
  NAND2_X1 u5_mult_82_U4028 ( .A1(u5_mult_82_ab_37__36_), .A2(
        u5_mult_82_CARRYB_36__36_), .ZN(u5_mult_82_n920) );
  NAND2_X2 u5_mult_82_U4027 ( .A1(u5_mult_82_ab_37__36_), .A2(
        u5_mult_82_SUMB_36__37_), .ZN(u5_mult_82_n919) );
  NAND2_X1 u5_mult_82_U4026 ( .A1(u5_mult_82_CARRYB_36__36_), .A2(
        u5_mult_82_SUMB_36__37_), .ZN(u5_mult_82_n918) );
  XOR2_X2 u5_mult_82_U4025 ( .A(u5_mult_82_SUMB_36__37_), .B(u5_mult_82_n917), 
        .Z(u5_mult_82_SUMB_37__36_) );
  XOR2_X2 u5_mult_82_U4024 ( .A(u5_mult_82_CARRYB_36__36_), .B(
        u5_mult_82_ab_37__36_), .Z(u5_mult_82_n917) );
  INV_X1 u5_mult_82_U4023 ( .A(u5_mult_82_SUMB_38__37_), .ZN(u5_mult_82_n914)
         );
  INV_X4 u5_mult_82_U4022 ( .A(u5_mult_82_n4471), .ZN(u5_mult_82_n913) );
  NAND2_X2 u5_mult_82_U4021 ( .A1(u5_mult_82_n913), .A2(
        u5_mult_82_SUMB_38__37_), .ZN(u5_mult_82_n916) );
  NAND2_X2 u5_mult_82_U4020 ( .A1(u5_mult_82_n4471), .A2(u5_mult_82_n914), 
        .ZN(u5_mult_82_n915) );
  NAND3_X2 u5_mult_82_U4019 ( .A1(u5_mult_82_n910), .A2(u5_mult_82_n911), .A3(
        u5_mult_82_n912), .ZN(u5_mult_82_CARRYB_14__47_) );
  NAND2_X1 u5_mult_82_U4018 ( .A1(u5_mult_82_n424), .A2(
        u5_mult_82_SUMB_13__48_), .ZN(u5_mult_82_n912) );
  NAND2_X1 u5_mult_82_U4017 ( .A1(u5_mult_82_ab_14__47_), .A2(
        u5_mult_82_SUMB_13__48_), .ZN(u5_mult_82_n911) );
  NAND2_X1 u5_mult_82_U4016 ( .A1(u5_mult_82_ab_14__47_), .A2(u5_mult_82_n424), 
        .ZN(u5_mult_82_n910) );
  NAND3_X2 u5_mult_82_U4015 ( .A1(u5_mult_82_n907), .A2(u5_mult_82_n908), .A3(
        u5_mult_82_n909), .ZN(u5_mult_82_CARRYB_13__48_) );
  NAND2_X2 u5_mult_82_U4014 ( .A1(u5_mult_82_ab_13__48_), .A2(
        u5_mult_82_SUMB_12__49_), .ZN(u5_mult_82_n908) );
  XOR2_X2 u5_mult_82_U4013 ( .A(u5_mult_82_n906), .B(u5_mult_82_SUMB_13__48_), 
        .Z(u5_mult_82_SUMB_14__47_) );
  XOR2_X2 u5_mult_82_U4012 ( .A(u5_mult_82_ab_14__47_), .B(u5_mult_82_n424), 
        .Z(u5_mult_82_n906) );
  XOR2_X2 u5_mult_82_U4011 ( .A(u5_mult_82_n905), .B(u5_mult_82_SUMB_12__49_), 
        .Z(u5_mult_82_SUMB_13__48_) );
  XOR2_X2 u5_mult_82_U4010 ( .A(u5_mult_82_ab_13__48_), .B(
        u5_mult_82_CARRYB_12__48_), .Z(u5_mult_82_n905) );
  NAND3_X2 u5_mult_82_U4009 ( .A1(u5_mult_82_n902), .A2(u5_mult_82_n903), .A3(
        u5_mult_82_n904), .ZN(u5_mult_82_CARRYB_3__50_) );
  NAND2_X2 u5_mult_82_U4008 ( .A1(u5_mult_82_ab_3__50_), .A2(
        u5_mult_82_SUMB_2__51_), .ZN(u5_mult_82_n904) );
  NAND2_X2 u5_mult_82_U4007 ( .A1(u5_mult_82_CARRYB_2__50_), .A2(
        u5_mult_82_SUMB_2__51_), .ZN(u5_mult_82_n903) );
  NAND2_X1 u5_mult_82_U4006 ( .A1(u5_mult_82_CARRYB_2__50_), .A2(
        u5_mult_82_ab_3__50_), .ZN(u5_mult_82_n902) );
  NAND3_X2 u5_mult_82_U4005 ( .A1(u5_mult_82_n899), .A2(u5_mult_82_n900), .A3(
        u5_mult_82_n901), .ZN(u5_mult_82_CARRYB_2__51_) );
  NAND2_X1 u5_mult_82_U4004 ( .A1(u5_mult_82_ab_2__51_), .A2(u5_mult_82_n965), 
        .ZN(u5_mult_82_n899) );
  NAND2_X2 u5_mult_82_U4003 ( .A1(u5_mult_82_ab_48__0_), .A2(
        u5_mult_82_SUMB_47__1_), .ZN(u5_mult_82_n2031) );
  NAND3_X4 u5_mult_82_U4002 ( .A1(u5_mult_82_n5631), .A2(u5_mult_82_n5632), 
        .A3(u5_mult_82_n5633), .ZN(u5_mult_82_CARRYB_42__2_) );
  NAND2_X2 u5_mult_82_U4001 ( .A1(n4783), .A2(n4822), .ZN(u5_mult_82_n1253) );
  INV_X2 u5_mult_82_U4000 ( .A(u5_mult_82_SUMB_28__24_), .ZN(u5_mult_82_n1521)
         );
  NAND3_X2 u5_mult_82_U3999 ( .A1(u5_mult_82_n6018), .A2(u5_mult_82_n6019), 
        .A3(u5_mult_82_n6020), .ZN(u5_mult_82_CARRYB_7__41_) );
  NAND2_X2 u5_mult_82_U3998 ( .A1(u5_mult_82_CARRYB_37__1_), .A2(
        u5_mult_82_ab_38__1_), .ZN(u5_mult_82_n2548) );
  INV_X1 u5_mult_82_U3997 ( .A(u5_mult_82_CARRYB_36__14_), .ZN(
        u5_mult_82_net81421) );
  INV_X4 u5_mult_82_U3996 ( .A(u5_mult_82_n6502), .ZN(u5_mult_82_CARRYB_1__46_) );
  XNOR2_X2 u5_mult_82_U3995 ( .A(u5_mult_82_n6502), .B(u5_mult_82_ab_2__46_), 
        .ZN(u5_mult_82_n1207) );
  XNOR2_X2 u5_mult_82_U3994 ( .A(u5_mult_82_ab_30__18_), .B(
        u5_mult_82_CARRYB_29__18_), .ZN(u5_mult_82_n898) );
  XNOR2_X2 u5_mult_82_U3993 ( .A(u5_mult_82_SUMB_29__19_), .B(u5_mult_82_n898), 
        .ZN(u5_mult_82_SUMB_30__18_) );
  XNOR2_X1 u5_mult_82_U3992 ( .A(u5_mult_82_CARRYB_5__26_), .B(
        u5_mult_82_ab_6__26_), .ZN(u5_mult_82_n897) );
  XNOR2_X2 u5_mult_82_U3991 ( .A(u5_mult_82_SUMB_5__27_), .B(u5_mult_82_n897), 
        .ZN(u5_mult_82_SUMB_6__26_) );
  XNOR2_X2 u5_mult_82_U3990 ( .A(u5_mult_82_ab_15__40_), .B(
        u5_mult_82_CARRYB_14__40_), .ZN(u5_mult_82_n896) );
  XNOR2_X2 u5_mult_82_U3989 ( .A(u5_mult_82_n896), .B(u5_mult_82_SUMB_14__41_), 
        .ZN(u5_mult_82_SUMB_15__40_) );
  XNOR2_X2 u5_mult_82_U3988 ( .A(u5_mult_82_ab_3__25_), .B(
        u5_mult_82_CARRYB_2__25_), .ZN(u5_mult_82_n895) );
  XNOR2_X2 u5_mult_82_U3987 ( .A(u5_mult_82_n895), .B(u5_mult_82_SUMB_2__26_), 
        .ZN(u5_mult_82_SUMB_3__25_) );
  NAND2_X2 u5_mult_82_U3986 ( .A1(u5_mult_82_CARRYB_26__15_), .A2(
        u5_mult_82_SUMB_26__16_), .ZN(u5_mult_82_n2785) );
  NAND3_X4 u5_mult_82_U3985 ( .A1(u5_mult_82_n2796), .A2(u5_mult_82_n2797), 
        .A3(u5_mult_82_n2798), .ZN(u5_mult_82_CARRYB_19__20_) );
  NAND2_X2 u5_mult_82_U3984 ( .A1(u5_mult_82_ab_23__26_), .A2(
        u5_mult_82_SUMB_22__27_), .ZN(u5_mult_82_n1904) );
  NAND2_X2 u5_mult_82_U3983 ( .A1(u5_mult_82_ab_6__38_), .A2(
        u5_mult_82_SUMB_5__39_), .ZN(u5_mult_82_n5616) );
  NAND2_X2 u5_mult_82_U3982 ( .A1(u5_mult_82_CARRYB_26__24_), .A2(
        u5_mult_82_SUMB_26__25_), .ZN(u5_mult_82_n5537) );
  NAND2_X1 u5_mult_82_U3981 ( .A1(u5_mult_82_CARRYB_21__31_), .A2(
        u5_mult_82_SUMB_21__32_), .ZN(u5_mult_82_n5268) );
  NAND2_X2 u5_mult_82_U3980 ( .A1(u5_mult_82_ab_7__44_), .A2(
        u5_mult_82_CARRYB_6__44_), .ZN(u5_mult_82_n6152) );
  NAND3_X4 u5_mult_82_U3979 ( .A1(u5_mult_82_n4996), .A2(u5_mult_82_n4997), 
        .A3(u5_mult_82_n4998), .ZN(u5_mult_82_CARRYB_6__44_) );
  NAND3_X2 u5_mult_82_U3978 ( .A1(u5_mult_82_n6054), .A2(u5_mult_82_n6053), 
        .A3(u5_mult_82_n6052), .ZN(u5_mult_82_CARRYB_24__25_) );
  NAND2_X2 u5_mult_82_U3977 ( .A1(u5_mult_82_CARRYB_38__2_), .A2(
        u5_mult_82_SUMB_38__3_), .ZN(u5_mult_82_n3483) );
  INV_X4 u5_mult_82_U3976 ( .A(u5_mult_82_SUMB_5__26_), .ZN(u5_mult_82_n1823)
         );
  XNOR2_X2 u5_mult_82_U3975 ( .A(u5_mult_82_n3815), .B(u5_mult_82_n1823), .ZN(
        u5_mult_82_SUMB_6__25_) );
  XNOR2_X2 u5_mult_82_U3974 ( .A(u5_mult_82_SUMB_13__37_), .B(
        u5_mult_82_ab_14__36_), .ZN(u5_mult_82_n1770) );
  NAND2_X2 u5_mult_82_U3973 ( .A1(u5_mult_82_CARRYB_6__38_), .A2(
        u5_mult_82_SUMB_6__39_), .ZN(u5_mult_82_n4746) );
  NAND2_X1 u5_mult_82_U3972 ( .A1(u5_mult_82_SUMB_14__34_), .A2(
        u5_mult_82_CARRYB_14__33_), .ZN(u5_mult_82_n4861) );
  NAND3_X2 u5_mult_82_U3971 ( .A1(u5_mult_82_n892), .A2(u5_mult_82_n893), .A3(
        u5_mult_82_n894), .ZN(u5_mult_82_CARRYB_8__35_) );
  NAND2_X1 u5_mult_82_U3970 ( .A1(u5_mult_82_CARRYB_7__35_), .A2(
        u5_mult_82_SUMB_7__36_), .ZN(u5_mult_82_n894) );
  NAND2_X1 u5_mult_82_U3969 ( .A1(u5_mult_82_ab_8__35_), .A2(
        u5_mult_82_SUMB_7__36_), .ZN(u5_mult_82_n893) );
  NAND2_X1 u5_mult_82_U3968 ( .A1(u5_mult_82_ab_8__35_), .A2(
        u5_mult_82_CARRYB_7__35_), .ZN(u5_mult_82_n892) );
  NAND3_X4 u5_mult_82_U3967 ( .A1(u5_mult_82_n889), .A2(u5_mult_82_n890), .A3(
        u5_mult_82_n891), .ZN(u5_mult_82_CARRYB_7__36_) );
  NAND2_X2 u5_mult_82_U3966 ( .A1(u5_mult_82_ab_7__36_), .A2(
        u5_mult_82_CARRYB_6__36_), .ZN(u5_mult_82_n889) );
  XOR2_X2 u5_mult_82_U3965 ( .A(u5_mult_82_n888), .B(u5_mult_82_SUMB_7__36_), 
        .Z(u5_mult_82_SUMB_8__35_) );
  XOR2_X2 u5_mult_82_U3964 ( .A(u5_mult_82_ab_8__35_), .B(
        u5_mult_82_CARRYB_7__35_), .Z(u5_mult_82_n888) );
  XOR2_X2 u5_mult_82_U3963 ( .A(u5_mult_82_n887), .B(u5_mult_82_SUMB_6__37_), 
        .Z(u5_mult_82_SUMB_7__36_) );
  XOR2_X2 u5_mult_82_U3962 ( .A(u5_mult_82_ab_7__36_), .B(
        u5_mult_82_CARRYB_6__36_), .Z(u5_mult_82_n887) );
  NAND3_X4 u5_mult_82_U3961 ( .A1(u5_mult_82_n884), .A2(u5_mult_82_n885), .A3(
        u5_mult_82_n886), .ZN(u5_mult_82_CARRYB_6__36_) );
  NAND2_X2 u5_mult_82_U3960 ( .A1(u5_mult_82_ab_6__36_), .A2(
        u5_mult_82_SUMB_5__37_), .ZN(u5_mult_82_n886) );
  NAND2_X2 u5_mult_82_U3959 ( .A1(u5_mult_82_CARRYB_5__36_), .A2(
        u5_mult_82_SUMB_5__37_), .ZN(u5_mult_82_n885) );
  NAND2_X1 u5_mult_82_U3958 ( .A1(u5_mult_82_CARRYB_5__36_), .A2(
        u5_mult_82_ab_6__36_), .ZN(u5_mult_82_n884) );
  NAND3_X2 u5_mult_82_U3957 ( .A1(u5_mult_82_n881), .A2(u5_mult_82_n882), .A3(
        u5_mult_82_n883), .ZN(u5_mult_82_CARRYB_5__37_) );
  NAND2_X2 u5_mult_82_U3956 ( .A1(u5_mult_82_ab_5__37_), .A2(
        u5_mult_82_SUMB_4__38_), .ZN(u5_mult_82_n883) );
  NAND2_X1 u5_mult_82_U3955 ( .A1(u5_mult_82_CARRYB_4__37_), .A2(
        u5_mult_82_SUMB_4__38_), .ZN(u5_mult_82_n882) );
  NAND2_X1 u5_mult_82_U3954 ( .A1(u5_mult_82_CARRYB_4__37_), .A2(
        u5_mult_82_ab_5__37_), .ZN(u5_mult_82_n881) );
  XOR2_X2 u5_mult_82_U3953 ( .A(u5_mult_82_n880), .B(u5_mult_82_SUMB_5__37_), 
        .Z(u5_mult_82_SUMB_6__36_) );
  XOR2_X2 u5_mult_82_U3952 ( .A(u5_mult_82_CARRYB_5__36_), .B(
        u5_mult_82_ab_6__36_), .Z(u5_mult_82_n880) );
  XNOR2_X2 u5_mult_82_U3951 ( .A(u5_mult_82_n4868), .B(u5_mult_82_n5197), .ZN(
        u5_mult_82_SUMB_13__36_) );
  NOR2_X1 u5_mult_82_U3950 ( .A1(u5_mult_82_n6960), .A2(u5_mult_82_n6717), 
        .ZN(u5_mult_82_ab_36__2_) );
  NAND3_X2 u5_mult_82_U3949 ( .A1(u5_mult_82_n876), .A2(u5_mult_82_n877), .A3(
        u5_mult_82_n878), .ZN(u5_mult_82_CARRYB_36__2_) );
  NAND2_X1 u5_mult_82_U3948 ( .A1(u5_mult_82_ab_36__2_), .A2(
        u5_mult_82_SUMB_35__3_), .ZN(u5_mult_82_n878) );
  NAND2_X2 u5_mult_82_U3947 ( .A1(u5_mult_82_ab_36__2_), .A2(
        u5_mult_82_CARRYB_35__2_), .ZN(u5_mult_82_n877) );
  XOR2_X2 u5_mult_82_U3946 ( .A(u5_mult_82_n13), .B(u5_mult_82_n875), .Z(
        u5_mult_82_SUMB_36__2_) );
  XOR2_X2 u5_mult_82_U3945 ( .A(u5_mult_82_SUMB_35__3_), .B(
        u5_mult_82_ab_36__2_), .Z(u5_mult_82_n875) );
  NAND3_X2 u5_mult_82_U3944 ( .A1(u5_mult_82_n872), .A2(u5_mult_82_n873), .A3(
        u5_mult_82_n874), .ZN(u5_mult_82_CARRYB_11__11_) );
  NAND2_X1 u5_mult_82_U3943 ( .A1(u5_mult_82_CARRYB_10__11_), .A2(
        u5_mult_82_SUMB_10__12_), .ZN(u5_mult_82_n874) );
  NAND2_X1 u5_mult_82_U3942 ( .A1(u5_mult_82_ab_11__11_), .A2(
        u5_mult_82_SUMB_10__12_), .ZN(u5_mult_82_n873) );
  NAND2_X1 u5_mult_82_U3941 ( .A1(u5_mult_82_ab_11__11_), .A2(
        u5_mult_82_CARRYB_10__11_), .ZN(u5_mult_82_n872) );
  NAND3_X2 u5_mult_82_U3940 ( .A1(u5_mult_82_n869), .A2(u5_mult_82_n870), .A3(
        u5_mult_82_n871), .ZN(u5_mult_82_CARRYB_10__12_) );
  NAND2_X2 u5_mult_82_U3939 ( .A1(u5_mult_82_CARRYB_9__12_), .A2(
        u5_mult_82_SUMB_9__13_), .ZN(u5_mult_82_n871) );
  NAND2_X2 u5_mult_82_U3938 ( .A1(u5_mult_82_ab_10__12_), .A2(
        u5_mult_82_SUMB_9__13_), .ZN(u5_mult_82_n870) );
  NAND2_X1 u5_mult_82_U3937 ( .A1(u5_mult_82_ab_10__12_), .A2(
        u5_mult_82_CARRYB_9__12_), .ZN(u5_mult_82_n869) );
  XOR2_X2 u5_mult_82_U3936 ( .A(u5_mult_82_n868), .B(u5_mult_82_SUMB_10__12_), 
        .Z(u5_mult_82_SUMB_11__11_) );
  XOR2_X1 u5_mult_82_U3935 ( .A(u5_mult_82_ab_11__11_), .B(
        u5_mult_82_CARRYB_10__11_), .Z(u5_mult_82_n868) );
  XOR2_X2 u5_mult_82_U3934 ( .A(u5_mult_82_n867), .B(u5_mult_82_SUMB_9__13_), 
        .Z(u5_mult_82_SUMB_10__12_) );
  XOR2_X2 u5_mult_82_U3933 ( .A(u5_mult_82_ab_10__12_), .B(
        u5_mult_82_CARRYB_9__12_), .Z(u5_mult_82_n867) );
  NAND3_X2 u5_mult_82_U3932 ( .A1(u5_mult_82_n864), .A2(u5_mult_82_n865), .A3(
        u5_mult_82_n866), .ZN(u5_mult_82_CARRYB_7__15_) );
  NAND2_X1 u5_mult_82_U3931 ( .A1(u5_mult_82_CARRYB_6__15_), .A2(
        u5_mult_82_SUMB_6__16_), .ZN(u5_mult_82_n866) );
  NAND2_X1 u5_mult_82_U3930 ( .A1(u5_mult_82_ab_7__15_), .A2(
        u5_mult_82_SUMB_6__16_), .ZN(u5_mult_82_n865) );
  NAND2_X1 u5_mult_82_U3929 ( .A1(u5_mult_82_ab_7__15_), .A2(
        u5_mult_82_CARRYB_6__15_), .ZN(u5_mult_82_n864) );
  NAND3_X2 u5_mult_82_U3928 ( .A1(u5_mult_82_n861), .A2(u5_mult_82_n862), .A3(
        u5_mult_82_n863), .ZN(u5_mult_82_CARRYB_6__16_) );
  NAND2_X1 u5_mult_82_U3927 ( .A1(u5_mult_82_CARRYB_5__16_), .A2(
        u5_mult_82_SUMB_5__17_), .ZN(u5_mult_82_n863) );
  NAND2_X1 u5_mult_82_U3926 ( .A1(u5_mult_82_ab_6__16_), .A2(
        u5_mult_82_SUMB_5__17_), .ZN(u5_mult_82_n862) );
  NAND2_X1 u5_mult_82_U3925 ( .A1(u5_mult_82_ab_6__16_), .A2(
        u5_mult_82_CARRYB_5__16_), .ZN(u5_mult_82_n861) );
  XOR2_X2 u5_mult_82_U3924 ( .A(u5_mult_82_n860), .B(u5_mult_82_SUMB_6__16_), 
        .Z(u5_mult_82_SUMB_7__15_) );
  XOR2_X1 u5_mult_82_U3923 ( .A(u5_mult_82_ab_7__15_), .B(
        u5_mult_82_CARRYB_6__15_), .Z(u5_mult_82_n860) );
  XOR2_X2 u5_mult_82_U3922 ( .A(u5_mult_82_n859), .B(u5_mult_82_SUMB_5__17_), 
        .Z(u5_mult_82_SUMB_6__16_) );
  XOR2_X2 u5_mult_82_U3921 ( .A(u5_mult_82_ab_6__16_), .B(
        u5_mult_82_CARRYB_5__16_), .Z(u5_mult_82_n859) );
  XNOR2_X2 u5_mult_82_U3920 ( .A(u5_mult_82_ab_7__38_), .B(
        u5_mult_82_CARRYB_6__38_), .ZN(u5_mult_82_n1246) );
  XNOR2_X1 u5_mult_82_U3919 ( .A(u5_mult_82_CARRYB_32__22_), .B(
        u5_mult_82_ab_33__22_), .ZN(u5_mult_82_n1519) );
  NAND3_X4 u5_mult_82_U3918 ( .A1(u5_mult_82_n5893), .A2(u5_mult_82_n5894), 
        .A3(u5_mult_82_n5895), .ZN(u5_mult_82_CARRYB_34__21_) );
  NAND2_X2 u5_mult_82_U3917 ( .A1(u5_mult_82_CARRYB_8__38_), .A2(
        u5_mult_82_n1452), .ZN(u5_mult_82_n5899) );
  XOR2_X2 u5_mult_82_U3916 ( .A(u5_mult_82_ab_25__28_), .B(
        u5_mult_82_CARRYB_24__28_), .Z(u5_mult_82_n1135) );
  NAND2_X2 u5_mult_82_U3915 ( .A1(u5_mult_82_ab_38__3_), .A2(
        u5_mult_82_CARRYB_37__3_), .ZN(u5_mult_82_n3430) );
  NAND2_X2 u5_mult_82_U3914 ( .A1(u5_mult_82_CARRYB_48__8_), .A2(
        u5_mult_82_SUMB_48__9_), .ZN(u5_mult_82_n5264) );
  NAND3_X2 u5_mult_82_U3913 ( .A1(u5_mult_82_n5611), .A2(u5_mult_82_n5612), 
        .A3(u5_mult_82_n5613), .ZN(u5_mult_82_CARRYB_20__24_) );
  XOR2_X2 u5_mult_82_U3912 ( .A(u5_mult_82_n3815), .B(u5_mult_82_n1824), .Z(
        u5_mult_82_n1667) );
  INV_X4 u5_mult_82_U3911 ( .A(u5_mult_82_n1823), .ZN(u5_mult_82_n1824) );
  INV_X8 u5_mult_82_U3910 ( .A(u5_mult_82_CARRYB_41__9_), .ZN(u5_mult_82_n3648) );
  NAND3_X4 u5_mult_82_U3909 ( .A1(u5_mult_82_n5021), .A2(u5_mult_82_n5022), 
        .A3(u5_mult_82_n5023), .ZN(u5_mult_82_CARRYB_15__36_) );
  NAND2_X2 u5_mult_82_U3908 ( .A1(u5_mult_82_ab_7__38_), .A2(
        u5_mult_82_SUMB_6__39_), .ZN(u5_mult_82_n4745) );
  NAND2_X2 u5_mult_82_U3907 ( .A1(u5_mult_82_SUMB_16__32_), .A2(
        u5_mult_82_CARRYB_16__31_), .ZN(u5_mult_82_n5916) );
  XNOR2_X2 u5_mult_82_U3906 ( .A(u5_mult_82_ab_20__40_), .B(
        u5_mult_82_CARRYB_19__40_), .ZN(u5_mult_82_n2053) );
  NAND2_X4 u5_mult_82_U3905 ( .A1(u5_mult_82_ab_4__47_), .A2(u5_mult_82_n1772), 
        .ZN(u5_mult_82_n2421) );
  NAND2_X2 u5_mult_82_U3904 ( .A1(u5_mult_82_CARRYB_23__21_), .A2(
        u5_mult_82_SUMB_23__22_), .ZN(u5_mult_82_n5692) );
  XNOR2_X2 u5_mult_82_U3903 ( .A(u5_mult_82_CARRYB_38__2_), .B(
        u5_mult_82_ab_39__2_), .ZN(u5_mult_82_n1855) );
  NAND3_X2 u5_mult_82_U3902 ( .A1(u5_mult_82_n3159), .A2(u5_mult_82_n3160), 
        .A3(u5_mult_82_n3161), .ZN(u5_mult_82_CARRYB_27__18_) );
  NAND3_X4 u5_mult_82_U3901 ( .A1(u5_mult_82_n5693), .A2(u5_mult_82_n5694), 
        .A3(u5_mult_82_n5695), .ZN(u5_mult_82_CARRYB_25__20_) );
  XNOR2_X2 u5_mult_82_U3900 ( .A(u5_mult_82_ab_14__22_), .B(
        u5_mult_82_CARRYB_13__22_), .ZN(u5_mult_82_n856) );
  XNOR2_X2 u5_mult_82_U3899 ( .A(u5_mult_82_n856), .B(u5_mult_82_SUMB_13__23_), 
        .ZN(u5_mult_82_SUMB_14__22_) );
  NAND2_X2 u5_mult_82_U3898 ( .A1(u5_mult_82_ab_21__23_), .A2(
        u5_mult_82_CARRYB_20__23_), .ZN(u5_mult_82_n3617) );
  NAND3_X2 u5_mult_82_U3897 ( .A1(u5_mult_82_n4515), .A2(u5_mult_82_n4516), 
        .A3(u5_mult_82_n4517), .ZN(u5_mult_82_CARRYB_47__2_) );
  NAND2_X2 u5_mult_82_U3896 ( .A1(u5_mult_82_n5638), .A2(
        u5_mult_82_SUMB_44__4_), .ZN(u5_mult_82_n3563) );
  NAND3_X2 u5_mult_82_U3895 ( .A1(u5_mult_82_n853), .A2(u5_mult_82_n854), .A3(
        u5_mult_82_n855), .ZN(u5_mult_82_CARRYB_20__3_) );
  NAND2_X1 u5_mult_82_U3894 ( .A1(u5_mult_82_CARRYB_19__3_), .A2(
        u5_mult_82_SUMB_19__4_), .ZN(u5_mult_82_n855) );
  NAND2_X1 u5_mult_82_U3893 ( .A1(u5_mult_82_ab_20__3_), .A2(
        u5_mult_82_SUMB_19__4_), .ZN(u5_mult_82_n854) );
  NAND2_X1 u5_mult_82_U3892 ( .A1(u5_mult_82_ab_20__3_), .A2(
        u5_mult_82_CARRYB_19__3_), .ZN(u5_mult_82_n853) );
  NAND3_X2 u5_mult_82_U3891 ( .A1(u5_mult_82_n850), .A2(u5_mult_82_n851), .A3(
        u5_mult_82_n852), .ZN(u5_mult_82_CARRYB_19__4_) );
  NAND2_X2 u5_mult_82_U3890 ( .A1(u5_mult_82_CARRYB_18__4_), .A2(
        u5_mult_82_SUMB_18__5_), .ZN(u5_mult_82_n852) );
  NAND2_X2 u5_mult_82_U3889 ( .A1(u5_mult_82_ab_19__4_), .A2(
        u5_mult_82_SUMB_18__5_), .ZN(u5_mult_82_n851) );
  NAND2_X1 u5_mult_82_U3888 ( .A1(u5_mult_82_ab_19__4_), .A2(
        u5_mult_82_CARRYB_18__4_), .ZN(u5_mult_82_n850) );
  XOR2_X2 u5_mult_82_U3887 ( .A(u5_mult_82_n849), .B(u5_mult_82_SUMB_19__4_), 
        .Z(u5_mult_82_SUMB_20__3_) );
  XOR2_X2 u5_mult_82_U3886 ( .A(u5_mult_82_ab_20__3_), .B(
        u5_mult_82_CARRYB_19__3_), .Z(u5_mult_82_n849) );
  XOR2_X2 u5_mult_82_U3885 ( .A(u5_mult_82_n848), .B(u5_mult_82_SUMB_18__5_), 
        .Z(u5_mult_82_SUMB_19__4_) );
  XOR2_X1 u5_mult_82_U3884 ( .A(u5_mult_82_ab_19__4_), .B(
        u5_mult_82_CARRYB_18__4_), .Z(u5_mult_82_n848) );
  XNOR2_X2 u5_mult_82_U3883 ( .A(u5_mult_82_ab_15__36_), .B(
        u5_mult_82_CARRYB_14__36_), .ZN(u5_mult_82_n847) );
  XNOR2_X2 u5_mult_82_U3882 ( .A(u5_mult_82_n1859), .B(u5_mult_82_n847), .ZN(
        u5_mult_82_SUMB_15__36_) );
  NAND2_X2 u5_mult_82_U3881 ( .A1(u5_mult_82_SUMB_25__15_), .A2(
        u5_mult_82_CARRYB_25__14_), .ZN(u5_mult_82_n4065) );
  NAND3_X4 u5_mult_82_U3880 ( .A1(u5_mult_82_n1903), .A2(u5_mult_82_n1904), 
        .A3(u5_mult_82_n1905), .ZN(u5_mult_82_CARRYB_23__26_) );
  NAND2_X2 u5_mult_82_U3879 ( .A1(u5_mult_82_CARRYB_24__19_), .A2(
        u5_mult_82_SUMB_24__20_), .ZN(u5_mult_82_n4786) );
  NAND2_X2 u5_mult_82_U3878 ( .A1(u5_mult_82_ab_1__47_), .A2(
        u5_mult_82_ab_0__48_), .ZN(u5_mult_82_n6504) );
  NAND2_X2 u5_mult_82_U3877 ( .A1(u5_mult_82_ab_7__25_), .A2(
        u5_mult_82_CARRYB_6__25_), .ZN(u5_mult_82_n3985) );
  NAND2_X2 u5_mult_82_U3876 ( .A1(u5_mult_82_ab_26__15_), .A2(
        u5_mult_82_SUMB_25__16_), .ZN(u5_mult_82_n2996) );
  NAND2_X2 u5_mult_82_U3875 ( .A1(u5_mult_82_ab_22__23_), .A2(
        u5_mult_82_SUMB_21__24_), .ZN(u5_mult_82_n1347) );
  NAND2_X2 u5_mult_82_U3874 ( .A1(u5_mult_82_ab_22__23_), .A2(
        u5_mult_82_CARRYB_21__23_), .ZN(u5_mult_82_n1346) );
  XNOR2_X2 u5_mult_82_U3873 ( .A(u5_mult_82_n1644), .B(u5_mult_82_SUMB_28__16_), .ZN(u5_mult_82_SUMB_29__15_) );
  XOR2_X2 u5_mult_82_U3872 ( .A(u5_mult_82_CARRYB_49__2_), .B(
        u5_mult_82_ab_50__2_), .Z(u5_mult_82_n989) );
  NAND2_X1 u5_mult_82_U3871 ( .A1(u5_mult_82_ab_15__46_), .A2(
        u5_mult_82_SUMB_14__47_), .ZN(u5_mult_82_n4878) );
  CLKBUF_X3 u5_mult_82_U3870 ( .A(u5_mult_82_SUMB_14__47_), .Z(
        u5_mult_82_n1782) );
  CLKBUF_X3 u5_mult_82_U3869 ( .A(u5_mult_82_SUMB_37__30_), .Z(
        u5_mult_82_n1820) );
  NAND3_X2 u5_mult_82_U3868 ( .A1(u5_mult_82_n844), .A2(u5_mult_82_n845), .A3(
        u5_mult_82_n846), .ZN(u5_mult_82_CARRYB_20__4_) );
  NAND2_X2 u5_mult_82_U3867 ( .A1(u5_mult_82_CARRYB_19__4_), .A2(
        u5_mult_82_SUMB_19__5_), .ZN(u5_mult_82_n846) );
  NAND2_X2 u5_mult_82_U3866 ( .A1(u5_mult_82_ab_20__4_), .A2(
        u5_mult_82_SUMB_19__5_), .ZN(u5_mult_82_n845) );
  NAND2_X1 u5_mult_82_U3865 ( .A1(u5_mult_82_ab_20__4_), .A2(
        u5_mult_82_CARRYB_19__4_), .ZN(u5_mult_82_n844) );
  NAND3_X2 u5_mult_82_U3864 ( .A1(u5_mult_82_n841), .A2(u5_mult_82_n842), .A3(
        u5_mult_82_n843), .ZN(u5_mult_82_CARRYB_19__5_) );
  NAND2_X2 u5_mult_82_U3863 ( .A1(u5_mult_82_CARRYB_18__5_), .A2(
        u5_mult_82_SUMB_18__6_), .ZN(u5_mult_82_n843) );
  NAND2_X2 u5_mult_82_U3862 ( .A1(u5_mult_82_ab_19__5_), .A2(
        u5_mult_82_SUMB_18__6_), .ZN(u5_mult_82_n842) );
  NAND2_X1 u5_mult_82_U3861 ( .A1(u5_mult_82_ab_19__5_), .A2(
        u5_mult_82_CARRYB_18__5_), .ZN(u5_mult_82_n841) );
  XOR2_X2 u5_mult_82_U3860 ( .A(u5_mult_82_n840), .B(u5_mult_82_SUMB_19__5_), 
        .Z(u5_mult_82_SUMB_20__4_) );
  XOR2_X2 u5_mult_82_U3859 ( .A(u5_mult_82_ab_20__4_), .B(
        u5_mult_82_CARRYB_19__4_), .Z(u5_mult_82_n840) );
  XOR2_X2 u5_mult_82_U3858 ( .A(u5_mult_82_n839), .B(u5_mult_82_SUMB_18__6_), 
        .Z(u5_mult_82_SUMB_19__5_) );
  XOR2_X2 u5_mult_82_U3857 ( .A(u5_mult_82_ab_19__5_), .B(
        u5_mult_82_CARRYB_18__5_), .Z(u5_mult_82_n839) );
  XNOR2_X2 u5_mult_82_U3856 ( .A(u5_mult_82_n1527), .B(u5_mult_82_n838), .ZN(
        u5_mult_82_n5682) );
  NOR2_X4 u5_mult_82_U3855 ( .A1(u5_mult_82_net64217), .A2(u5_mult_82_n7007), 
        .ZN(u5_mult_82_ab_0__46_) );
  NAND2_X2 u5_mult_82_U3854 ( .A1(u5_mult_82_CARRYB_6__37_), .A2(
        u5_mult_82_SUMB_6__38_), .ZN(u5_mult_82_n5620) );
  NOR2_X1 u5_mult_82_U3853 ( .A1(u5_mult_82_n6941), .A2(u5_mult_82_n6630), 
        .ZN(u5_mult_82_ab_21__7_) );
  NAND3_X2 u5_mult_82_U3852 ( .A1(u5_mult_82_n835), .A2(u5_mult_82_n836), .A3(
        u5_mult_82_n837), .ZN(u5_mult_82_CARRYB_21__7_) );
  NAND2_X1 u5_mult_82_U3851 ( .A1(u5_mult_82_ab_21__7_), .A2(
        u5_mult_82_CARRYB_20__7_), .ZN(u5_mult_82_n837) );
  NAND2_X2 u5_mult_82_U3850 ( .A1(u5_mult_82_ab_21__7_), .A2(
        u5_mult_82_SUMB_20__8_), .ZN(u5_mult_82_n836) );
  NAND2_X1 u5_mult_82_U3849 ( .A1(u5_mult_82_CARRYB_20__7_), .A2(
        u5_mult_82_SUMB_20__8_), .ZN(u5_mult_82_n835) );
  XOR2_X2 u5_mult_82_U3848 ( .A(u5_mult_82_SUMB_20__8_), .B(u5_mult_82_n834), 
        .Z(u5_mult_82_SUMB_21__7_) );
  XOR2_X2 u5_mult_82_U3847 ( .A(u5_mult_82_CARRYB_20__7_), .B(
        u5_mult_82_ab_21__7_), .Z(u5_mult_82_n834) );
  NAND3_X2 u5_mult_82_U3846 ( .A1(u5_mult_82_n831), .A2(u5_mult_82_n832), .A3(
        u5_mult_82_n833), .ZN(u5_mult_82_CARRYB_25__3_) );
  NAND2_X1 u5_mult_82_U3845 ( .A1(u5_mult_82_CARRYB_24__3_), .A2(
        u5_mult_82_SUMB_24__4_), .ZN(u5_mult_82_n833) );
  NAND2_X1 u5_mult_82_U3844 ( .A1(u5_mult_82_ab_25__3_), .A2(
        u5_mult_82_SUMB_24__4_), .ZN(u5_mult_82_n832) );
  NAND2_X1 u5_mult_82_U3843 ( .A1(u5_mult_82_ab_25__3_), .A2(
        u5_mult_82_CARRYB_24__3_), .ZN(u5_mult_82_n831) );
  NAND3_X2 u5_mult_82_U3842 ( .A1(u5_mult_82_n828), .A2(u5_mult_82_n829), .A3(
        u5_mult_82_n830), .ZN(u5_mult_82_CARRYB_24__4_) );
  NAND2_X2 u5_mult_82_U3841 ( .A1(u5_mult_82_CARRYB_23__4_), .A2(
        u5_mult_82_SUMB_23__5_), .ZN(u5_mult_82_n830) );
  NAND2_X2 u5_mult_82_U3840 ( .A1(u5_mult_82_ab_24__4_), .A2(
        u5_mult_82_SUMB_23__5_), .ZN(u5_mult_82_n829) );
  NAND2_X1 u5_mult_82_U3839 ( .A1(u5_mult_82_ab_24__4_), .A2(
        u5_mult_82_CARRYB_23__4_), .ZN(u5_mult_82_n828) );
  XOR2_X2 u5_mult_82_U3838 ( .A(u5_mult_82_n827), .B(u5_mult_82_SUMB_24__4_), 
        .Z(u5_mult_82_SUMB_25__3_) );
  XOR2_X2 u5_mult_82_U3837 ( .A(u5_mult_82_ab_25__3_), .B(
        u5_mult_82_CARRYB_24__3_), .Z(u5_mult_82_n827) );
  XOR2_X2 u5_mult_82_U3836 ( .A(u5_mult_82_n826), .B(u5_mult_82_n51), .Z(
        u5_mult_82_SUMB_24__4_) );
  XOR2_X2 u5_mult_82_U3835 ( .A(u5_mult_82_ab_24__4_), .B(
        u5_mult_82_CARRYB_23__4_), .Z(u5_mult_82_n826) );
  XNOR2_X2 u5_mult_82_U3834 ( .A(u5_mult_82_ab_5__27_), .B(
        u5_mult_82_CARRYB_4__27_), .ZN(u5_mult_82_n1801) );
  NAND2_X2 u5_mult_82_U3833 ( .A1(u5_mult_82_CARRYB_4__27_), .A2(
        u5_mult_82_SUMB_4__28_), .ZN(u5_mult_82_n3983) );
  INV_X2 u5_mult_82_U3832 ( .A(u5_mult_82_SUMB_47__23_), .ZN(u5_mult_82_n1611)
         );
  NAND2_X2 u5_mult_82_U3831 ( .A1(u5_mult_82_ab_35__13_), .A2(
        u5_mult_82_CARRYB_34__13_), .ZN(u5_mult_82_n4954) );
  NAND3_X4 u5_mult_82_U3830 ( .A1(u5_mult_82_n4956), .A2(u5_mult_82_n4955), 
        .A3(u5_mult_82_n4954), .ZN(u5_mult_82_CARRYB_35__13_) );
  NAND2_X2 u5_mult_82_U3829 ( .A1(u5_mult_82_SUMB_3__50_), .A2(
        u5_mult_82_n1468), .ZN(u5_mult_82_n6316) );
  NAND2_X2 u5_mult_82_U3828 ( .A1(u5_mult_82_SUMB_9__47_), .A2(
        u5_mult_82_CARRYB_9__46_), .ZN(u5_mult_82_n5731) );
  NAND3_X4 u5_mult_82_U3827 ( .A1(u5_mult_82_n5313), .A2(u5_mult_82_n5314), 
        .A3(u5_mult_82_n5315), .ZN(u5_mult_82_CARRYB_11__30_) );
  NAND3_X2 u5_mult_82_U3826 ( .A1(u5_mult_82_n6096), .A2(u5_mult_82_n6097), 
        .A3(u5_mult_82_n6098), .ZN(u5_mult_82_CARRYB_7__43_) );
  NAND3_X4 u5_mult_82_U3825 ( .A1(u5_mult_82_n5399), .A2(u5_mult_82_n5400), 
        .A3(u5_mult_82_n5401), .ZN(u5_mult_82_CARRYB_10__42_) );
  NAND3_X2 u5_mult_82_U3824 ( .A1(u5_mult_82_n4849), .A2(u5_mult_82_n4850), 
        .A3(u5_mult_82_n4851), .ZN(u5_mult_82_CARRYB_40__0_) );
  NAND2_X2 u5_mult_82_U3823 ( .A1(u5_mult_82_ab_5__27_), .A2(
        u5_mult_82_SUMB_4__28_), .ZN(u5_mult_82_n3982) );
  NAND3_X2 u5_mult_82_U3822 ( .A1(u5_mult_82_n823), .A2(u5_mult_82_n824), .A3(
        u5_mult_82_n825), .ZN(u5_mult_82_CARRYB_24__6_) );
  NAND2_X2 u5_mult_82_U3821 ( .A1(u5_mult_82_ab_24__6_), .A2(
        u5_mult_82_SUMB_23__7_), .ZN(u5_mult_82_n825) );
  NAND2_X2 u5_mult_82_U3820 ( .A1(u5_mult_82_CARRYB_23__6_), .A2(
        u5_mult_82_SUMB_23__7_), .ZN(u5_mult_82_n824) );
  NAND2_X1 u5_mult_82_U3819 ( .A1(u5_mult_82_CARRYB_23__6_), .A2(
        u5_mult_82_ab_24__6_), .ZN(u5_mult_82_n823) );
  NAND3_X2 u5_mult_82_U3818 ( .A1(u5_mult_82_n820), .A2(u5_mult_82_n821), .A3(
        u5_mult_82_n822), .ZN(u5_mult_82_CARRYB_23__7_) );
  NAND2_X2 u5_mult_82_U3817 ( .A1(u5_mult_82_CARRYB_22__7_), .A2(
        u5_mult_82_SUMB_22__8_), .ZN(u5_mult_82_n822) );
  NAND2_X2 u5_mult_82_U3816 ( .A1(u5_mult_82_ab_23__7_), .A2(
        u5_mult_82_SUMB_22__8_), .ZN(u5_mult_82_n821) );
  NAND2_X2 u5_mult_82_U3815 ( .A1(u5_mult_82_ab_23__7_), .A2(
        u5_mult_82_CARRYB_22__7_), .ZN(u5_mult_82_n820) );
  XOR2_X2 u5_mult_82_U3814 ( .A(u5_mult_82_n819), .B(u5_mult_82_SUMB_23__7_), 
        .Z(u5_mult_82_SUMB_24__6_) );
  XOR2_X2 u5_mult_82_U3813 ( .A(u5_mult_82_CARRYB_23__6_), .B(
        u5_mult_82_ab_24__6_), .Z(u5_mult_82_n819) );
  XOR2_X2 u5_mult_82_U3812 ( .A(u5_mult_82_n818), .B(u5_mult_82_SUMB_22__8_), 
        .Z(u5_mult_82_SUMB_23__7_) );
  XOR2_X2 u5_mult_82_U3811 ( .A(u5_mult_82_ab_23__7_), .B(
        u5_mult_82_CARRYB_22__7_), .Z(u5_mult_82_n818) );
  NAND3_X2 u5_mult_82_U3810 ( .A1(u5_mult_82_n815), .A2(u5_mult_82_n816), .A3(
        u5_mult_82_n817), .ZN(u5_mult_82_CARRYB_26__4_) );
  NAND2_X2 u5_mult_82_U3809 ( .A1(u5_mult_82_CARRYB_25__4_), .A2(
        u5_mult_82_SUMB_25__5_), .ZN(u5_mult_82_n817) );
  NAND2_X2 u5_mult_82_U3808 ( .A1(u5_mult_82_ab_26__4_), .A2(
        u5_mult_82_SUMB_25__5_), .ZN(u5_mult_82_n816) );
  NAND2_X1 u5_mult_82_U3807 ( .A1(u5_mult_82_ab_26__4_), .A2(
        u5_mult_82_CARRYB_25__4_), .ZN(u5_mult_82_n815) );
  NAND3_X2 u5_mult_82_U3806 ( .A1(u5_mult_82_n812), .A2(u5_mult_82_n813), .A3(
        u5_mult_82_n814), .ZN(u5_mult_82_CARRYB_25__5_) );
  NAND2_X2 u5_mult_82_U3805 ( .A1(u5_mult_82_CARRYB_24__5_), .A2(
        u5_mult_82_SUMB_24__6_), .ZN(u5_mult_82_n814) );
  NAND2_X2 u5_mult_82_U3804 ( .A1(u5_mult_82_ab_25__5_), .A2(
        u5_mult_82_SUMB_24__6_), .ZN(u5_mult_82_n813) );
  NAND2_X1 u5_mult_82_U3803 ( .A1(u5_mult_82_ab_25__5_), .A2(
        u5_mult_82_CARRYB_24__5_), .ZN(u5_mult_82_n812) );
  XOR2_X2 u5_mult_82_U3802 ( .A(u5_mult_82_n811), .B(u5_mult_82_SUMB_25__5_), 
        .Z(u5_mult_82_SUMB_26__4_) );
  XOR2_X2 u5_mult_82_U3801 ( .A(u5_mult_82_ab_26__4_), .B(
        u5_mult_82_CARRYB_25__4_), .Z(u5_mult_82_n811) );
  XOR2_X2 u5_mult_82_U3800 ( .A(u5_mult_82_n810), .B(u5_mult_82_SUMB_24__6_), 
        .Z(u5_mult_82_SUMB_25__5_) );
  XOR2_X2 u5_mult_82_U3799 ( .A(u5_mult_82_ab_25__5_), .B(
        u5_mult_82_CARRYB_24__5_), .Z(u5_mult_82_n810) );
  NAND2_X4 u5_mult_82_U3798 ( .A1(u5_mult_82_CARRYB_3__47_), .A2(
        u5_mult_82_n1772), .ZN(u5_mult_82_n2420) );
  NAND2_X2 u5_mult_82_U3797 ( .A1(u5_mult_82_ab_10__30_), .A2(
        u5_mult_82_CARRYB_9__30_), .ZN(u5_mult_82_n2302) );
  NAND3_X4 u5_mult_82_U3796 ( .A1(u5_mult_82_n2205), .A2(u5_mult_82_n2206), 
        .A3(u5_mult_82_n2207), .ZN(u5_mult_82_CARRYB_8__30_) );
  NOR2_X1 u5_mult_82_U3795 ( .A1(u5_mult_82_n6859), .A2(u5_mult_82_n6544), 
        .ZN(u5_mult_82_ab_9__30_) );
  NAND3_X2 u5_mult_82_U3794 ( .A1(u5_mult_82_n807), .A2(u5_mult_82_n808), .A3(
        u5_mult_82_n809), .ZN(u5_mult_82_CARRYB_9__30_) );
  NAND2_X1 u5_mult_82_U3793 ( .A1(u5_mult_82_ab_9__30_), .A2(
        u5_mult_82_CARRYB_8__30_), .ZN(u5_mult_82_n809) );
  NAND2_X2 u5_mult_82_U3792 ( .A1(u5_mult_82_ab_9__30_), .A2(
        u5_mult_82_SUMB_8__31_), .ZN(u5_mult_82_n808) );
  NAND2_X1 u5_mult_82_U3791 ( .A1(u5_mult_82_CARRYB_8__30_), .A2(
        u5_mult_82_SUMB_8__31_), .ZN(u5_mult_82_n807) );
  XOR2_X2 u5_mult_82_U3790 ( .A(u5_mult_82_SUMB_8__31_), .B(u5_mult_82_n806), 
        .Z(u5_mult_82_SUMB_9__30_) );
  XOR2_X2 u5_mult_82_U3789 ( .A(u5_mult_82_CARRYB_8__30_), .B(
        u5_mult_82_ab_9__30_), .Z(u5_mult_82_n806) );
  INV_X16 u5_mult_82_U3788 ( .A(u5_mult_82_n6807), .ZN(u5_mult_82_n6805) );
  INV_X16 u5_mult_82_U3787 ( .A(u5_mult_82_n6807), .ZN(u5_mult_82_n6806) );
  INV_X4 u5_mult_82_U3786 ( .A(u5_mult_82_n7009), .ZN(u5_mult_82_n6807) );
  NAND2_X4 u5_mult_82_U3785 ( .A1(u5_mult_82_n5184), .A2(u5_mult_82_ab_12__38_), .ZN(u5_mult_82_n6090) );
  NAND2_X1 u5_mult_82_U3784 ( .A1(u5_mult_82_CARRYB_3__33_), .A2(
        u5_mult_82_SUMB_3__34_), .ZN(u5_mult_82_n4505) );
  XNOR2_X2 u5_mult_82_U3783 ( .A(u5_mult_82_CARRYB_11__23_), .B(
        u5_mult_82_n805), .ZN(u5_mult_82_n996) );
  NAND2_X1 u5_mult_82_U3782 ( .A1(u5_mult_82_ab_33__17_), .A2(
        u5_mult_82_CARRYB_32__17_), .ZN(u5_mult_82_n3304) );
  NAND2_X1 u5_mult_82_U3781 ( .A1(u5_mult_82_ab_11__44_), .A2(
        u5_mult_82_CARRYB_10__44_), .ZN(u5_mult_82_n5644) );
  NAND3_X4 u5_mult_82_U3780 ( .A1(u5_mult_82_n2991), .A2(u5_mult_82_n2992), 
        .A3(u5_mult_82_n2993), .ZN(u5_mult_82_CARRYB_25__16_) );
  NAND2_X1 u5_mult_82_U3779 ( .A1(u5_mult_82_ab_31__18_), .A2(
        u5_mult_82_SUMB_30__19_), .ZN(u5_mult_82_net83289) );
  NAND3_X4 u5_mult_82_U3778 ( .A1(u5_mult_82_n801), .A2(u5_mult_82_n802), .A3(
        u5_mult_82_n803), .ZN(u5_mult_82_CARRYB_13__34_) );
  NAND2_X1 u5_mult_82_U3777 ( .A1(u5_mult_82_CARRYB_12__34_), .A2(
        u5_mult_82_SUMB_12__35_), .ZN(u5_mult_82_n803) );
  NAND2_X1 u5_mult_82_U3776 ( .A1(u5_mult_82_ab_13__34_), .A2(
        u5_mult_82_SUMB_12__35_), .ZN(u5_mult_82_n802) );
  NAND2_X1 u5_mult_82_U3775 ( .A1(u5_mult_82_ab_13__34_), .A2(
        u5_mult_82_CARRYB_12__34_), .ZN(u5_mult_82_n801) );
  NAND3_X2 u5_mult_82_U3774 ( .A1(u5_mult_82_n798), .A2(u5_mult_82_n799), .A3(
        u5_mult_82_n800), .ZN(u5_mult_82_CARRYB_12__35_) );
  NAND2_X2 u5_mult_82_U3773 ( .A1(u5_mult_82_CARRYB_11__35_), .A2(
        u5_mult_82_SUMB_11__36_), .ZN(u5_mult_82_n800) );
  NAND2_X2 u5_mult_82_U3772 ( .A1(u5_mult_82_ab_12__35_), .A2(
        u5_mult_82_SUMB_11__36_), .ZN(u5_mult_82_n799) );
  NAND2_X1 u5_mult_82_U3771 ( .A1(u5_mult_82_ab_12__35_), .A2(
        u5_mult_82_CARRYB_11__35_), .ZN(u5_mult_82_n798) );
  XOR2_X2 u5_mult_82_U3770 ( .A(u5_mult_82_n797), .B(u5_mult_82_SUMB_12__35_), 
        .Z(u5_mult_82_SUMB_13__34_) );
  XOR2_X2 u5_mult_82_U3769 ( .A(u5_mult_82_CARRYB_12__34_), .B(
        u5_mult_82_ab_13__34_), .Z(u5_mult_82_n797) );
  XOR2_X2 u5_mult_82_U3768 ( .A(u5_mult_82_n796), .B(u5_mult_82_SUMB_11__36_), 
        .Z(u5_mult_82_SUMB_12__35_) );
  XOR2_X2 u5_mult_82_U3767 ( .A(u5_mult_82_ab_12__35_), .B(
        u5_mult_82_CARRYB_11__35_), .Z(u5_mult_82_n796) );
  NAND2_X2 u5_mult_82_U3766 ( .A1(u5_mult_82_ab_14__39_), .A2(
        u5_mult_82_CARRYB_13__39_), .ZN(u5_mult_82_n5352) );
  XOR2_X2 u5_mult_82_U3765 ( .A(u5_mult_82_CARRYB_37__3_), .B(
        u5_mult_82_ab_38__3_), .Z(u5_mult_82_n3427) );
  NAND2_X2 u5_mult_82_U3764 ( .A1(u5_mult_82_n1033), .A2(u5_mult_82_n1034), 
        .ZN(u5_mult_82_n1617) );
  BUF_X4 u5_mult_82_U3763 ( .A(u5_mult_82_SUMB_9__46_), .Z(u5_mult_82_n1449)
         );
  NOR2_X4 u5_mult_82_U3762 ( .A1(u5_mult_82_n6769), .A2(u5_mult_82_net66087), 
        .ZN(u5_mult_82_ab_2__50_) );
  XNOR2_X2 u5_mult_82_U3761 ( .A(u5_mult_82_ab_46__9_), .B(
        u5_mult_82_CARRYB_45__9_), .ZN(u5_mult_82_n795) );
  XNOR2_X2 u5_mult_82_U3760 ( .A(u5_mult_82_n795), .B(u5_mult_82_SUMB_45__10_), 
        .ZN(u5_mult_82_SUMB_46__9_) );
  NAND2_X2 u5_mult_82_U3759 ( .A1(u5_mult_82_CARRYB_10__44_), .A2(
        u5_mult_82_SUMB_10__45_), .ZN(u5_mult_82_n5642) );
  NAND2_X2 u5_mult_82_U3758 ( .A1(u5_mult_82_ab_15__38_), .A2(u5_mult_82_n421), 
        .ZN(u5_mult_82_n5355) );
  XNOR2_X2 u5_mult_82_U3757 ( .A(u5_mult_82_ab_15__38_), .B(u5_mult_82_n421), 
        .ZN(u5_mult_82_n1937) );
  NAND3_X2 u5_mult_82_U3756 ( .A1(u5_mult_82_n5642), .A2(u5_mult_82_n5643), 
        .A3(u5_mult_82_n5644), .ZN(u5_mult_82_CARRYB_11__44_) );
  NAND2_X2 u5_mult_82_U3755 ( .A1(u5_mult_82_ab_49__8_), .A2(
        u5_mult_82_SUMB_48__9_), .ZN(u5_mult_82_n5263) );
  NAND3_X4 u5_mult_82_U3754 ( .A1(u5_mult_82_n5262), .A2(u5_mult_82_n5263), 
        .A3(u5_mult_82_n5264), .ZN(u5_mult_82_CARRYB_49__8_) );
  NAND2_X2 u5_mult_82_U3753 ( .A1(u5_mult_82_SUMB_38__15_), .A2(
        u5_mult_82_CARRYB_38__14_), .ZN(u5_mult_82_net82678) );
  NAND2_X2 u5_mult_82_U3752 ( .A1(u5_mult_82_ab_50__17_), .A2(
        u5_mult_82_SUMB_49__18_), .ZN(u5_mult_82_n4399) );
  NAND3_X2 u5_mult_82_U3751 ( .A1(u5_mult_82_n792), .A2(u5_mult_82_n793), .A3(
        u5_mult_82_n794), .ZN(u5_mult_82_CARRYB_52__12_) );
  NAND2_X1 u5_mult_82_U3750 ( .A1(u5_mult_82_CARRYB_51__12_), .A2(
        u5_mult_82_SUMB_51__13_), .ZN(u5_mult_82_n794) );
  NAND2_X1 u5_mult_82_U3749 ( .A1(u5_mult_82_ab_52__12_), .A2(
        u5_mult_82_SUMB_51__13_), .ZN(u5_mult_82_n793) );
  NAND2_X1 u5_mult_82_U3748 ( .A1(u5_mult_82_ab_52__12_), .A2(
        u5_mult_82_CARRYB_51__12_), .ZN(u5_mult_82_n792) );
  NAND3_X2 u5_mult_82_U3747 ( .A1(u5_mult_82_n789), .A2(u5_mult_82_n790), .A3(
        u5_mult_82_n791), .ZN(u5_mult_82_CARRYB_51__13_) );
  NAND2_X2 u5_mult_82_U3746 ( .A1(u5_mult_82_CARRYB_50__13_), .A2(
        u5_mult_82_SUMB_50__14_), .ZN(u5_mult_82_n791) );
  NAND2_X2 u5_mult_82_U3745 ( .A1(u5_mult_82_ab_51__13_), .A2(
        u5_mult_82_SUMB_50__14_), .ZN(u5_mult_82_n790) );
  NAND2_X1 u5_mult_82_U3744 ( .A1(u5_mult_82_ab_51__13_), .A2(
        u5_mult_82_CARRYB_50__13_), .ZN(u5_mult_82_n789) );
  XOR2_X2 u5_mult_82_U3743 ( .A(u5_mult_82_n788), .B(u5_mult_82_SUMB_51__13_), 
        .Z(u5_mult_82_SUMB_52__12_) );
  XOR2_X2 u5_mult_82_U3742 ( .A(u5_mult_82_ab_52__12_), .B(
        u5_mult_82_CARRYB_51__12_), .Z(u5_mult_82_n788) );
  XOR2_X2 u5_mult_82_U3741 ( .A(u5_mult_82_n787), .B(u5_mult_82_SUMB_50__14_), 
        .Z(u5_mult_82_SUMB_51__13_) );
  XOR2_X2 u5_mult_82_U3740 ( .A(u5_mult_82_ab_51__13_), .B(
        u5_mult_82_CARRYB_50__13_), .Z(u5_mult_82_n787) );
  INV_X4 u5_mult_82_U3739 ( .A(u5_mult_82_n4362), .ZN(u5_mult_82_n783) );
  NAND2_X4 u5_mult_82_U3738 ( .A1(u5_mult_82_n785), .A2(u5_mult_82_n786), .ZN(
        u5_mult_82_SUMB_50__14_) );
  NAND2_X4 u5_mult_82_U3737 ( .A1(u5_mult_82_n783), .A2(u5_mult_82_n784), .ZN(
        u5_mult_82_n786) );
  NAND3_X2 u5_mult_82_U3736 ( .A1(u5_mult_82_n3058), .A2(u5_mult_82_n3059), 
        .A3(u5_mult_82_net84199), .ZN(u5_mult_82_CARRYB_24__23_) );
  XNOR2_X2 u5_mult_82_U3735 ( .A(u5_mult_82_SUMB_24__16_), .B(u5_mult_82_n782), 
        .ZN(u5_mult_82_SUMB_25__15_) );
  INV_X4 u5_mult_82_U3734 ( .A(u5_mult_82_SUMB_31__32_), .ZN(u5_mult_82_n1799)
         );
  NOR2_X2 u5_mult_82_U3733 ( .A1(u5_mult_82_net64683), .A2(u5_mult_82_net65285), .ZN(u5_mult_82_ab_47__23_) );
  NAND3_X2 u5_mult_82_U3732 ( .A1(u5_mult_82_n779), .A2(u5_mult_82_n780), .A3(
        u5_mult_82_n781), .ZN(u5_mult_82_CARRYB_47__23_) );
  NAND2_X2 u5_mult_82_U3731 ( .A1(u5_mult_82_ab_47__23_), .A2(
        u5_mult_82_CARRYB_46__23_), .ZN(u5_mult_82_n781) );
  NAND2_X1 u5_mult_82_U3730 ( .A1(u5_mult_82_ab_47__23_), .A2(
        u5_mult_82_SUMB_46__24_), .ZN(u5_mult_82_n780) );
  NAND2_X1 u5_mult_82_U3729 ( .A1(u5_mult_82_CARRYB_46__23_), .A2(
        u5_mult_82_SUMB_46__24_), .ZN(u5_mult_82_n779) );
  XOR2_X2 u5_mult_82_U3728 ( .A(u5_mult_82_CARRYB_46__23_), .B(
        u5_mult_82_ab_47__23_), .Z(u5_mult_82_n778) );
  NAND3_X2 u5_mult_82_U3727 ( .A1(u5_mult_82_n3292), .A2(u5_mult_82_n3291), 
        .A3(u5_mult_82_n3290), .ZN(u5_mult_82_CARRYB_6__37_) );
  XNOR2_X2 u5_mult_82_U3726 ( .A(u5_mult_82_SUMB_46__19_), .B(u5_mult_82_n5650), .ZN(u5_mult_82_SUMB_47__18_) );
  NAND3_X4 u5_mult_82_U3725 ( .A1(u5_mult_82_n3629), .A2(u5_mult_82_n3630), 
        .A3(u5_mult_82_n3631), .ZN(u5_mult_82_CARRYB_51__15_) );
  NOR2_X1 u5_mult_82_U3724 ( .A1(u5_mult_82_n6975), .A2(u5_mult_82_n6933), 
        .ZN(u5_mult_82_ab_52__15_) );
  INV_X1 u5_mult_82_U3723 ( .A(u5_mult_82_SUMB_45__20_), .ZN(u5_mult_82_n775)
         );
  INV_X4 u5_mult_82_U3722 ( .A(u5_mult_82_n3844), .ZN(u5_mult_82_n774) );
  NAND2_X4 u5_mult_82_U3721 ( .A1(u5_mult_82_n776), .A2(u5_mult_82_n777), .ZN(
        u5_mult_82_SUMB_46__19_) );
  NAND2_X2 u5_mult_82_U3720 ( .A1(u5_mult_82_n774), .A2(
        u5_mult_82_SUMB_45__20_), .ZN(u5_mult_82_n777) );
  NAND2_X2 u5_mult_82_U3719 ( .A1(u5_mult_82_n3844), .A2(u5_mult_82_n775), 
        .ZN(u5_mult_82_n776) );
  NAND3_X2 u5_mult_82_U3718 ( .A1(u5_mult_82_n771), .A2(u5_mult_82_n772), .A3(
        u5_mult_82_n773), .ZN(u5_mult_82_CARRYB_52__15_) );
  NAND2_X1 u5_mult_82_U3717 ( .A1(u5_mult_82_ab_52__15_), .A2(
        u5_mult_82_CARRYB_51__15_), .ZN(u5_mult_82_n773) );
  NAND2_X2 u5_mult_82_U3716 ( .A1(u5_mult_82_ab_52__15_), .A2(
        u5_mult_82_SUMB_51__16_), .ZN(u5_mult_82_n772) );
  NAND2_X1 u5_mult_82_U3715 ( .A1(u5_mult_82_CARRYB_51__15_), .A2(
        u5_mult_82_SUMB_51__16_), .ZN(u5_mult_82_n771) );
  XOR2_X2 u5_mult_82_U3714 ( .A(u5_mult_82_SUMB_51__16_), .B(u5_mult_82_n770), 
        .Z(u5_mult_82_SUMB_52__15_) );
  XOR2_X2 u5_mult_82_U3713 ( .A(u5_mult_82_CARRYB_51__15_), .B(
        u5_mult_82_ab_52__15_), .Z(u5_mult_82_n770) );
  NAND2_X4 u5_mult_82_U3712 ( .A1(u5_mult_82_ab_0__28_), .A2(
        u5_mult_82_ab_1__27_), .ZN(u5_mult_82_n6480) );
  NAND2_X1 u5_mult_82_U3711 ( .A1(u5_mult_82_CARRYB_8__28_), .A2(
        u5_mult_82_SUMB_8__29_), .ZN(u5_mult_82_n3448) );
  XNOR2_X2 u5_mult_82_U3710 ( .A(u5_mult_82_n1504), .B(u5_mult_82_ab_41__1_), 
        .ZN(u5_mult_82_n769) );
  XNOR2_X2 u5_mult_82_U3709 ( .A(u5_mult_82_SUMB_40__2_), .B(u5_mult_82_n769), 
        .ZN(u5_mult_82_SUMB_41__1_) );
  XNOR2_X2 u5_mult_82_U3708 ( .A(u5_mult_82_CARRYB_28__16_), .B(
        u5_mult_82_ab_29__16_), .ZN(u5_mult_82_n768) );
  XNOR2_X2 u5_mult_82_U3707 ( .A(u5_mult_82_SUMB_28__17_), .B(u5_mult_82_n768), 
        .ZN(u5_mult_82_SUMB_29__16_) );
  XNOR2_X2 u5_mult_82_U3706 ( .A(u5_mult_82_n1510), .B(u5_mult_82_ab_7__41_), 
        .ZN(u5_mult_82_n1400) );
  NOR2_X4 u5_mult_82_U3705 ( .A1(u5_mult_82_n6800), .A2(u5_mult_82_net66087), 
        .ZN(u5_mult_82_ab_2__45_) );
  XNOR2_X2 u5_mult_82_U3704 ( .A(u5_mult_82_CARRYB_38__19_), .B(
        u5_mult_82_ab_39__19_), .ZN(u5_mult_82_n767) );
  NAND2_X1 u5_mult_82_U3703 ( .A1(u5_mult_82_ab_26__35_), .A2(
        u5_mult_82_CARRYB_25__35_), .ZN(u5_mult_82_n4402) );
  NAND2_X2 u5_mult_82_U3702 ( .A1(u5_mult_82_CARRYB_21__38_), .A2(
        u5_mult_82_SUMB_21__39_), .ZN(u5_mult_82_n2256) );
  INV_X4 u5_mult_82_U3701 ( .A(u5_mult_82_SUMB_3__48_), .ZN(u5_mult_82_n1771)
         );
  INV_X2 u5_mult_82_U3700 ( .A(u5_mult_82_n2643), .ZN(u5_mult_82_n2519) );
  NAND2_X2 u5_mult_82_U3699 ( .A1(u5_mult_82_ab_48__9_), .A2(
        u5_mult_82_CARRYB_47__9_), .ZN(u5_mult_82_n5259) );
  INV_X4 u5_mult_82_U3698 ( .A(u5_mult_82_n6409), .ZN(u5_mult_82_CLA_SUM[75])
         );
  NAND3_X4 u5_mult_82_U3697 ( .A1(u5_mult_82_n4419), .A2(u5_mult_82_n4420), 
        .A3(u5_mult_82_n4421), .ZN(u5_mult_82_CARRYB_41__30_) );
  NAND3_X4 u5_mult_82_U3696 ( .A1(u5_mult_82_n6372), .A2(u5_mult_82_n6373), 
        .A3(u5_mult_82_n6374), .ZN(u5_mult_82_CARRYB_22__35_) );
  NOR2_X1 u5_mult_82_U3695 ( .A1(u5_mult_82_net64903), .A2(u5_mult_82_net65711), .ZN(u5_mult_82_ab_23__35_) );
  NAND3_X2 u5_mult_82_U3694 ( .A1(u5_mult_82_n764), .A2(u5_mult_82_n765), .A3(
        u5_mult_82_n766), .ZN(u5_mult_82_CARRYB_23__35_) );
  NAND2_X1 u5_mult_82_U3693 ( .A1(u5_mult_82_ab_23__35_), .A2(
        u5_mult_82_CARRYB_22__35_), .ZN(u5_mult_82_n766) );
  NAND2_X2 u5_mult_82_U3692 ( .A1(u5_mult_82_ab_23__35_), .A2(
        u5_mult_82_SUMB_22__36_), .ZN(u5_mult_82_n765) );
  NAND2_X1 u5_mult_82_U3691 ( .A1(u5_mult_82_CARRYB_22__35_), .A2(
        u5_mult_82_SUMB_22__36_), .ZN(u5_mult_82_n764) );
  XOR2_X2 u5_mult_82_U3690 ( .A(u5_mult_82_SUMB_22__36_), .B(u5_mult_82_n763), 
        .Z(u5_mult_82_SUMB_23__35_) );
  XOR2_X2 u5_mult_82_U3689 ( .A(u5_mult_82_CARRYB_22__35_), .B(
        u5_mult_82_ab_23__35_), .Z(u5_mult_82_n763) );
  NAND3_X4 u5_mult_82_U3688 ( .A1(u5_mult_82_n759), .A2(u5_mult_82_n760), .A3(
        u5_mult_82_n761), .ZN(u5_mult_82_CARRYB_32__29_) );
  NAND2_X1 u5_mult_82_U3687 ( .A1(u5_mult_82_CARRYB_31__29_), .A2(
        u5_mult_82_SUMB_31__30_), .ZN(u5_mult_82_n761) );
  NAND2_X1 u5_mult_82_U3686 ( .A1(u5_mult_82_ab_32__29_), .A2(
        u5_mult_82_SUMB_31__30_), .ZN(u5_mult_82_n760) );
  NAND2_X1 u5_mult_82_U3685 ( .A1(u5_mult_82_ab_32__29_), .A2(
        u5_mult_82_CARRYB_31__29_), .ZN(u5_mult_82_n759) );
  NAND3_X4 u5_mult_82_U3684 ( .A1(u5_mult_82_n756), .A2(u5_mult_82_n757), .A3(
        u5_mult_82_n758), .ZN(u5_mult_82_CARRYB_31__30_) );
  NAND2_X2 u5_mult_82_U3683 ( .A1(u5_mult_82_CARRYB_30__30_), .A2(
        u5_mult_82_SUMB_30__31_), .ZN(u5_mult_82_n758) );
  NAND2_X2 u5_mult_82_U3682 ( .A1(u5_mult_82_ab_31__30_), .A2(
        u5_mult_82_SUMB_30__31_), .ZN(u5_mult_82_n757) );
  NAND2_X1 u5_mult_82_U3681 ( .A1(u5_mult_82_ab_31__30_), .A2(
        u5_mult_82_CARRYB_30__30_), .ZN(u5_mult_82_n756) );
  XOR2_X2 u5_mult_82_U3680 ( .A(u5_mult_82_n755), .B(u5_mult_82_SUMB_31__30_), 
        .Z(u5_mult_82_SUMB_32__29_) );
  XOR2_X2 u5_mult_82_U3679 ( .A(u5_mult_82_ab_32__29_), .B(
        u5_mult_82_CARRYB_31__29_), .Z(u5_mult_82_n755) );
  XOR2_X2 u5_mult_82_U3678 ( .A(u5_mult_82_n754), .B(u5_mult_82_SUMB_30__31_), 
        .Z(u5_mult_82_SUMB_31__30_) );
  XOR2_X2 u5_mult_82_U3677 ( .A(u5_mult_82_ab_31__30_), .B(
        u5_mult_82_CARRYB_30__30_), .Z(u5_mult_82_n754) );
  XNOR2_X1 u5_mult_82_U3676 ( .A(u5_mult_82_CARRYB_26__15_), .B(
        u5_mult_82_ab_27__15_), .ZN(u5_mult_82_n753) );
  XNOR2_X2 u5_mult_82_U3675 ( .A(u5_mult_82_n753), .B(u5_mult_82_SUMB_26__16_), 
        .ZN(u5_mult_82_SUMB_27__15_) );
  NAND2_X2 u5_mult_82_U3674 ( .A1(u5_mult_82_ab_27__35_), .A2(
        u5_mult_82_CARRYB_26__35_), .ZN(u5_mult_82_n4934) );
  NOR2_X4 u5_mult_82_U3673 ( .A1(u5_mult_82_net64903), .A2(u5_mult_82_n6656), 
        .ZN(u5_mult_82_ab_27__35_) );
  INV_X1 u5_mult_82_U3672 ( .A(u5_mult_82_ab_27__35_), .ZN(u5_mult_82_n750) );
  INV_X2 u5_mult_82_U3671 ( .A(u5_mult_82_CARRYB_26__35_), .ZN(u5_mult_82_n749) );
  NAND2_X2 u5_mult_82_U3670 ( .A1(u5_mult_82_n751), .A2(u5_mult_82_n752), .ZN(
        u5_mult_82_n4557) );
  NAND2_X2 u5_mult_82_U3669 ( .A1(u5_mult_82_n749), .A2(u5_mult_82_n750), .ZN(
        u5_mult_82_n752) );
  NAND2_X2 u5_mult_82_U3668 ( .A1(u5_mult_82_CARRYB_26__35_), .A2(
        u5_mult_82_ab_27__35_), .ZN(u5_mult_82_n751) );
  XNOR2_X2 u5_mult_82_U3667 ( .A(u5_mult_82_CARRYB_7__48_), .B(
        u5_mult_82_ab_8__48_), .ZN(u5_mult_82_n3275) );
  NAND2_X2 u5_mult_82_U3666 ( .A1(u5_mult_82_n1475), .A2(u5_mult_82_ab_38__30_), .ZN(u5_mult_82_n4711) );
  NAND2_X2 u5_mult_82_U3665 ( .A1(u5_mult_82_ab_32__14_), .A2(
        u5_mult_82_CARRYB_31__14_), .ZN(u5_mult_82_n3998) );
  XOR2_X2 u5_mult_82_U3664 ( .A(u5_mult_82_n3655), .B(u5_mult_82_SUMB_29__16_), 
        .Z(u5_mult_82_SUMB_30__15_) );
  INV_X16 u5_mult_82_U3663 ( .A(n4818), .ZN(u5_mult_82_n6765) );
  NAND2_X2 u5_mult_82_U3662 ( .A1(u5_mult_82_CARRYB_49__7_), .A2(
        u5_mult_82_SUMB_49__8_), .ZN(u5_mult_82_n5009) );
  NAND2_X2 u5_mult_82_U3661 ( .A1(u5_mult_82_CARRYB_39__13_), .A2(
        u5_mult_82_SUMB_39__14_), .ZN(u5_mult_82_n1911) );
  NAND2_X2 u5_mult_82_U3660 ( .A1(u5_mult_82_CARRYB_40__16_), .A2(
        u5_mult_82_SUMB_40__17_), .ZN(u5_mult_82_n5294) );
  INV_X2 u5_mult_82_U3659 ( .A(u5_mult_82_CARRYB_42__16_), .ZN(
        u5_mult_82_n5282) );
  NAND2_X2 u5_mult_82_U3658 ( .A1(u5_mult_82_SUMB_45__8_), .A2(
        u5_mult_82_CARRYB_45__7_), .ZN(u5_mult_82_n4379) );
  NAND3_X4 u5_mult_82_U3657 ( .A1(u5_mult_82_n6090), .A2(u5_mult_82_n6091), 
        .A3(u5_mult_82_n6089), .ZN(u5_mult_82_CARRYB_12__38_) );
  NOR2_X1 u5_mult_82_U3656 ( .A1(u5_mult_82_n6810), .A2(u5_mult_82_net65313), 
        .ZN(u5_mult_82_ab_45__43_) );
  NOR2_X1 u5_mult_82_U3655 ( .A1(u5_mult_82_n6810), .A2(u5_mult_82_n6740), 
        .ZN(u5_mult_82_ab_46__43_) );
  NOR2_X1 u5_mult_82_U3654 ( .A1(u5_mult_82_n6810), .A2(u5_mult_82_net65277), 
        .ZN(u5_mult_82_ab_47__43_) );
  NOR2_X1 u5_mult_82_U3653 ( .A1(u5_mult_82_n6810), .A2(u5_mult_82_n6746), 
        .ZN(u5_mult_82_ab_48__43_) );
  NOR2_X1 u5_mult_82_U3652 ( .A1(u5_mult_82_n6810), .A2(u5_mult_82_n6752), 
        .ZN(u5_mult_82_ab_49__43_) );
  NOR2_X1 u5_mult_82_U3651 ( .A1(u5_mult_82_n6810), .A2(u5_mult_82_net65223), 
        .ZN(u5_mult_82_ab_50__43_) );
  NOR2_X1 u5_mult_82_U3650 ( .A1(u5_mult_82_n6810), .A2(u5_mult_82_net65193), 
        .ZN(u5_mult_82_ab_51__43_) );
  NOR2_X1 u5_mult_82_U3649 ( .A1(u5_mult_82_n6977), .A2(u5_mult_82_n6810), 
        .ZN(u5_mult_82_ab_52__43_) );
  NAND2_X2 u5_mult_82_U3648 ( .A1(u5_mult_82_CARRYB_32__20_), .A2(
        u5_mult_82_SUMB_32__21_), .ZN(u5_mult_82_n1212) );
  NAND2_X2 u5_mult_82_U3647 ( .A1(u5_mult_82_CARRYB_25__25_), .A2(
        u5_mult_82_SUMB_25__26_), .ZN(u5_mult_82_n5532) );
  NAND2_X2 u5_mult_82_U3646 ( .A1(u5_mult_82_ab_35__19_), .A2(
        u5_mult_82_SUMB_34__20_), .ZN(u5_mult_82_n6337) );
  NAND2_X1 u5_mult_82_U3645 ( .A1(u5_mult_82_CARRYB_31__38_), .A2(
        u5_mult_82_SUMB_31__39_), .ZN(u5_mult_82_n4925) );
  NAND2_X2 u5_mult_82_U3644 ( .A1(u5_mult_82_CARRYB_36__35_), .A2(
        u5_mult_82_SUMB_36__36_), .ZN(u5_mult_82_n5126) );
  NAND2_X2 u5_mult_82_U3643 ( .A1(u5_mult_82_ab_5__47_), .A2(
        u5_mult_82_SUMB_4__48_), .ZN(u5_mult_82_n6194) );
  NAND2_X4 u5_mult_82_U3642 ( .A1(u5_mult_82_n2522), .A2(u5_mult_82_n2523), 
        .ZN(u5_mult_82_n2525) );
  NAND2_X4 u5_mult_82_U3641 ( .A1(u5_mult_82_n2524), .A2(u5_mult_82_n2525), 
        .ZN(u5_mult_82_SUMB_8__45_) );
  NAND2_X2 u5_mult_82_U3640 ( .A1(u5_mult_82_ab_30__11_), .A2(
        u5_mult_82_CARRYB_29__11_), .ZN(u5_mult_82_n5306) );
  NAND2_X2 u5_mult_82_U3639 ( .A1(u5_mult_82_ab_45__6_), .A2(
        u5_mult_82_CARRYB_44__6_), .ZN(u5_mult_82_n4656) );
  NAND2_X2 u5_mult_82_U3638 ( .A1(u5_mult_82_ab_47__12_), .A2(
        u5_mult_82_SUMB_46__13_), .ZN(u5_mult_82_n6232) );
  XOR2_X2 u5_mult_82_U3637 ( .A(u5_mult_82_ab_35__19_), .B(
        u5_mult_82_CARRYB_34__19_), .Z(u5_mult_82_n6332) );
  XNOR2_X2 u5_mult_82_U3636 ( .A(u5_mult_82_ab_8__30_), .B(
        u5_mult_82_CARRYB_7__30_), .ZN(u5_mult_82_n748) );
  XNOR2_X2 u5_mult_82_U3635 ( .A(u5_mult_82_n748), .B(u5_mult_82_SUMB_7__31_), 
        .ZN(u5_mult_82_SUMB_8__30_) );
  XNOR2_X2 u5_mult_82_U3634 ( .A(u5_mult_82_ab_41__14_), .B(
        u5_mult_82_CARRYB_40__14_), .ZN(u5_mult_82_n747) );
  XNOR2_X2 u5_mult_82_U3633 ( .A(u5_mult_82_n747), .B(u5_mult_82_n720), .ZN(
        u5_mult_82_SUMB_41__14_) );
  XNOR2_X2 u5_mult_82_U3632 ( .A(u5_mult_82_SUMB_45__3_), .B(u5_mult_82_n746), 
        .ZN(u5_mult_82_SUMB_46__2_) );
  CLKBUF_X2 u5_mult_82_U3631 ( .A(u5_mult_82_SUMB_13__42_), .Z(u5_mult_82_n745) );
  XNOR2_X1 u5_mult_82_U3630 ( .A(u5_mult_82_ab_37__17_), .B(
        u5_mult_82_CARRYB_36__17_), .ZN(u5_mult_82_n744) );
  XNOR2_X2 u5_mult_82_U3629 ( .A(u5_mult_82_n744), .B(u5_mult_82_n304), .ZN(
        u5_mult_82_SUMB_37__17_) );
  INV_X8 u5_mult_82_U3628 ( .A(u5_mult_82_n742), .ZN(u5_mult_82_n743) );
  INV_X4 u5_mult_82_U3627 ( .A(u5_mult_82_SUMB_22__19_), .ZN(u5_mult_82_n742)
         );
  INV_X4 u5_mult_82_U3626 ( .A(u5_mult_82_n740), .ZN(u5_mult_82_n741) );
  INV_X2 u5_mult_82_U3625 ( .A(u5_mult_82_SUMB_37__19_), .ZN(u5_mult_82_n740)
         );
  XNOR2_X2 u5_mult_82_U3624 ( .A(u5_mult_82_ab_10__43_), .B(
        u5_mult_82_CARRYB_9__43_), .ZN(u5_mult_82_n739) );
  XNOR2_X2 u5_mult_82_U3623 ( .A(u5_mult_82_n739), .B(u5_mult_82_SUMB_9__44_), 
        .ZN(u5_mult_82_SUMB_10__43_) );
  INV_X2 u5_mult_82_U3622 ( .A(u5_mult_82_SUMB_36__17_), .ZN(u5_mult_82_n737)
         );
  INV_X8 u5_mult_82_U3621 ( .A(u5_mult_82_n734), .ZN(u5_mult_82_n735) );
  INV_X4 u5_mult_82_U3620 ( .A(u5_mult_82_SUMB_23__27_), .ZN(u5_mult_82_n1394)
         );
  XNOR2_X2 u5_mult_82_U3619 ( .A(u5_mult_82_n5968), .B(u5_mult_82_n1394), .ZN(
        u5_mult_82_SUMB_24__26_) );
  XNOR2_X2 u5_mult_82_U3618 ( .A(u5_mult_82_ab_40__17_), .B(
        u5_mult_82_CARRYB_39__17_), .ZN(u5_mult_82_n732) );
  XNOR2_X2 u5_mult_82_U3617 ( .A(u5_mult_82_n732), .B(u5_mult_82_SUMB_39__18_), 
        .ZN(u5_mult_82_SUMB_40__17_) );
  XNOR2_X2 u5_mult_82_U3616 ( .A(u5_mult_82_SUMB_25__15_), .B(u5_mult_82_n2290), .ZN(u5_mult_82_SUMB_26__14_) );
  NAND2_X1 u5_mult_82_U3615 ( .A1(u5_mult_82_CARRYB_40__4_), .A2(
        u5_mult_82_ab_41__4_), .ZN(u5_mult_82_n4960) );
  XNOR2_X2 u5_mult_82_U3614 ( .A(u5_mult_82_n731), .B(u5_mult_82_CARRYB_49__9_), .ZN(u5_mult_82_n4165) );
  CLKBUF_X3 u5_mult_82_U3613 ( .A(u5_mult_82_SUMB_30__7_), .Z(u5_mult_82_n729)
         );
  INV_X1 u5_mult_82_U3612 ( .A(u5_mult_82_SUMB_41__3_), .ZN(u5_mult_82_n728)
         );
  XNOR2_X2 u5_mult_82_U3611 ( .A(u5_mult_82_ab_49__8_), .B(
        u5_mult_82_CARRYB_48__8_), .ZN(u5_mult_82_n726) );
  XNOR2_X2 u5_mult_82_U3610 ( .A(u5_mult_82_n726), .B(u5_mult_82_SUMB_48__9_), 
        .ZN(u5_mult_82_SUMB_49__8_) );
  INV_X2 u5_mult_82_U3609 ( .A(u5_mult_82_n724), .ZN(u5_mult_82_n725) );
  INV_X1 u5_mult_82_U3608 ( .A(u5_mult_82_SUMB_52__7_), .ZN(u5_mult_82_n724)
         );
  CLKBUF_X2 u5_mult_82_U3607 ( .A(u5_mult_82_SUMB_25__16_), .Z(u5_mult_82_n723) );
  XNOR2_X2 u5_mult_82_U3606 ( .A(u5_mult_82_ab_26__16_), .B(
        u5_mult_82_CARRYB_25__16_), .ZN(u5_mult_82_n722) );
  XNOR2_X2 u5_mult_82_U3605 ( .A(u5_mult_82_n722), .B(u5_mult_82_SUMB_25__17_), 
        .ZN(u5_mult_82_SUMB_26__16_) );
  CLKBUF_X2 u5_mult_82_U3604 ( .A(u5_mult_82_CARRYB_44__18_), .Z(
        u5_mult_82_n721) );
  INV_X2 u5_mult_82_U3603 ( .A(u5_mult_82_n719), .ZN(u5_mult_82_n720) );
  INV_X1 u5_mult_82_U3602 ( .A(u5_mult_82_SUMB_40__15_), .ZN(u5_mult_82_n719)
         );
  INV_X8 u5_mult_82_U3601 ( .A(u5_mult_82_n717), .ZN(u5_mult_82_n718) );
  CLKBUF_X2 u5_mult_82_U3600 ( .A(u5_mult_82_CARRYB_35__15_), .Z(
        u5_mult_82_n716) );
  INV_X4 u5_mult_82_U3599 ( .A(u5_mult_82_n714), .ZN(u5_mult_82_n715) );
  INV_X2 u5_mult_82_U3598 ( .A(u5_mult_82_SUMB_27__20_), .ZN(u5_mult_82_n714)
         );
  CLKBUF_X2 u5_mult_82_U3597 ( .A(u5_mult_82_SUMB_49__3_), .Z(u5_mult_82_n713)
         );
  XNOR2_X2 u5_mult_82_U3596 ( .A(u5_mult_82_n712), .B(u5_mult_82_SUMB_42__13_), 
        .ZN(u5_mult_82_SUMB_43__12_) );
  XNOR2_X2 u5_mult_82_U3595 ( .A(u5_mult_82_SUMB_40__12_), .B(
        u5_mult_82_ab_41__11_), .ZN(u5_mult_82_n711) );
  XNOR2_X2 u5_mult_82_U3594 ( .A(u5_mult_82_CARRYB_40__11_), .B(
        u5_mult_82_n711), .ZN(u5_mult_82_SUMB_41__11_) );
  INV_X8 u5_mult_82_U3593 ( .A(u5_mult_82_n709), .ZN(u5_mult_82_n710) );
  INV_X2 u5_mult_82_U3592 ( .A(u5_mult_82_SUMB_35__37_), .ZN(u5_mult_82_n709)
         );
  XNOR2_X2 u5_mult_82_U3591 ( .A(u5_mult_82_ab_2__51_), .B(u5_mult_82_n965), 
        .ZN(u5_mult_82_n708) );
  XNOR2_X2 u5_mult_82_U3590 ( .A(u5_mult_82_n708), .B(u5_mult_82_n215), .ZN(
        u5_mult_82_SUMB_2__51_) );
  CLKBUF_X2 u5_mult_82_U3589 ( .A(u5_mult_82_SUMB_44__12_), .Z(u5_mult_82_n707) );
  INV_X4 u5_mult_82_U3588 ( .A(u5_mult_82_n705), .ZN(u5_mult_82_n706) );
  INV_X2 u5_mult_82_U3587 ( .A(u5_mult_82_CARRYB_39__27_), .ZN(u5_mult_82_n705) );
  XOR2_X1 u5_mult_82_U3586 ( .A(u5_mult_82_n6371), .B(u5_mult_82_SUMB_22__35_), 
        .Z(u5_mult_82_SUMB_23__34_) );
  XOR2_X2 u5_mult_82_U3585 ( .A(u5_mult_82_n6371), .B(u5_mult_82_SUMB_22__35_), 
        .Z(u5_mult_82_n704) );
  XNOR2_X1 u5_mult_82_U3584 ( .A(u5_mult_82_ab_19__35_), .B(
        u5_mult_82_CARRYB_18__35_), .ZN(u5_mult_82_n703) );
  XNOR2_X2 u5_mult_82_U3583 ( .A(u5_mult_82_n703), .B(u5_mult_82_SUMB_18__36_), 
        .ZN(u5_mult_82_SUMB_19__35_) );
  NAND2_X2 u5_mult_82_U3582 ( .A1(u5_mult_82_ab_20__32_), .A2(
        u5_mult_82_CARRYB_19__32_), .ZN(u5_mult_82_n3536) );
  INV_X2 u5_mult_82_U3581 ( .A(u5_mult_82_CARRYB_46__21_), .ZN(u5_mult_82_n701) );
  NAND2_X1 u5_mult_82_U3580 ( .A1(u5_mult_82_CARRYB_25__30_), .A2(
        u5_mult_82_SUMB_25__31_), .ZN(u5_mult_82_n6281) );
  NAND2_X1 u5_mult_82_U3579 ( .A1(u5_mult_82_CARRYB_24__25_), .A2(
        u5_mult_82_SUMB_24__26_), .ZN(u5_mult_82_n5974) );
  XNOR2_X2 u5_mult_82_U3578 ( .A(u5_mult_82_n700), .B(
        u5_mult_82_CARRYB_18__21_), .ZN(u5_mult_82_n4669) );
  XNOR2_X2 u5_mult_82_U3577 ( .A(u5_mult_82_ab_33__14_), .B(
        u5_mult_82_CARRYB_32__14_), .ZN(u5_mult_82_n699) );
  XNOR2_X2 u5_mult_82_U3576 ( .A(u5_mult_82_n699), .B(u5_mult_82_SUMB_32__15_), 
        .ZN(u5_mult_82_SUMB_33__14_) );
  XNOR2_X2 u5_mult_82_U3575 ( .A(u5_mult_82_ab_40__20_), .B(
        u5_mult_82_CARRYB_39__20_), .ZN(u5_mult_82_n698) );
  XNOR2_X2 u5_mult_82_U3574 ( .A(u5_mult_82_n698), .B(u5_mult_82_SUMB_39__21_), 
        .ZN(u5_mult_82_SUMB_40__20_) );
  XNOR2_X1 u5_mult_82_U3573 ( .A(u5_mult_82_CARRYB_17__45_), .B(
        u5_mult_82_ab_18__45_), .ZN(u5_mult_82_n1867) );
  NAND2_X1 u5_mult_82_U3572 ( .A1(u5_mult_82_CARRYB_17__45_), .A2(
        u5_mult_82_SUMB_17__46_), .ZN(u5_mult_82_n5874) );
  INV_X4 u5_mult_82_U3571 ( .A(u5_mult_82_n696), .ZN(u5_mult_82_n697) );
  INV_X2 u5_mult_82_U3570 ( .A(u5_mult_82_SUMB_44__15_), .ZN(u5_mult_82_n696)
         );
  CLKBUF_X2 u5_mult_82_U3569 ( .A(u5_mult_82_SUMB_20__24_), .Z(u5_mult_82_n695) );
  XNOR2_X2 u5_mult_82_U3568 ( .A(u5_mult_82_ab_28__37_), .B(
        u5_mult_82_CARRYB_27__37_), .ZN(u5_mult_82_n693) );
  XNOR2_X2 u5_mult_82_U3567 ( .A(u5_mult_82_n693), .B(u5_mult_82_SUMB_27__38_), 
        .ZN(u5_mult_82_SUMB_28__37_) );
  INV_X4 u5_mult_82_U3566 ( .A(u5_mult_82_n691), .ZN(u5_mult_82_n692) );
  INV_X2 u5_mult_82_U3565 ( .A(u5_mult_82_SUMB_18__21_), .ZN(u5_mult_82_n691)
         );
  XNOR2_X2 u5_mult_82_U3564 ( .A(u5_mult_82_CARRYB_15__15_), .B(
        u5_mult_82_ab_16__15_), .ZN(u5_mult_82_n690) );
  XNOR2_X2 u5_mult_82_U3563 ( .A(u5_mult_82_n690), .B(u5_mult_82_n1454), .ZN(
        u5_mult_82_SUMB_16__15_) );
  XNOR2_X2 u5_mult_82_U3562 ( .A(u5_mult_82_CARRYB_37__29_), .B(
        u5_mult_82_ab_38__29_), .ZN(u5_mult_82_n689) );
  XNOR2_X2 u5_mult_82_U3561 ( .A(u5_mult_82_n1820), .B(u5_mult_82_n689), .ZN(
        u5_mult_82_SUMB_38__29_) );
  XNOR2_X2 u5_mult_82_U3560 ( .A(u5_mult_82_ab_47__20_), .B(
        u5_mult_82_CARRYB_46__20_), .ZN(u5_mult_82_n688) );
  XNOR2_X2 u5_mult_82_U3559 ( .A(u5_mult_82_n688), .B(u5_mult_82_n1863), .ZN(
        u5_mult_82_SUMB_47__20_) );
  INV_X16 u5_mult_82_U3558 ( .A(u5_mult_82_n7009), .ZN(u5_mult_82_n6808) );
  INV_X2 u5_mult_82_U3557 ( .A(u5_mult_82_n6808), .ZN(u5_mult_82_n6804) );
  INV_X2 u5_mult_82_U3556 ( .A(u5_mult_82_n6835), .ZN(u5_mult_82_n6832) );
  NAND2_X2 u5_mult_82_U3555 ( .A1(u5_mult_82_CARRYB_13__29_), .A2(
        u5_mult_82_net83274), .ZN(u5_mult_82_net80252) );
  INV_X4 u5_mult_82_U3554 ( .A(u5_mult_82_n1492), .ZN(u5_mult_82_n1493) );
  NAND3_X4 u5_mult_82_U3553 ( .A1(u5_mult_82_n6100), .A2(u5_mult_82_n6101), 
        .A3(u5_mult_82_n6102), .ZN(u5_mult_82_CARRYB_8__42_) );
  XNOR2_X2 u5_mult_82_U3552 ( .A(u5_mult_82_CARRYB_39__6_), .B(
        u5_mult_82_ab_40__6_), .ZN(u5_mult_82_n5161) );
  XNOR2_X2 u5_mult_82_U3551 ( .A(u5_mult_82_ab_43__6_), .B(
        u5_mult_82_CARRYB_42__6_), .ZN(u5_mult_82_n1744) );
  NAND2_X2 u5_mult_82_U3550 ( .A1(u5_mult_82_CARRYB_5__38_), .A2(
        u5_mult_82_SUMB_5__39_), .ZN(u5_mult_82_n5615) );
  NAND2_X2 u5_mult_82_U3549 ( .A1(u5_mult_82_CARRYB_9__35_), .A2(
        u5_mult_82_SUMB_9__36_), .ZN(u5_mult_82_n5701) );
  XNOR2_X1 u5_mult_82_U3548 ( .A(u5_mult_82_n1678), .B(u5_mult_82_SUMB_9__36_), 
        .ZN(u5_mult_82_SUMB_10__35_) );
  NAND3_X2 u5_mult_82_U3547 ( .A1(u5_mult_82_n4859), .A2(u5_mult_82_n4860), 
        .A3(u5_mult_82_n4861), .ZN(u5_mult_82_CARRYB_15__33_) );
  NAND2_X1 u5_mult_82_U3546 ( .A1(u5_mult_82_ab_27__29_), .A2(
        u5_mult_82_SUMB_26__30_), .ZN(u5_mult_82_n6283) );
  NAND3_X2 u5_mult_82_U3545 ( .A1(u5_mult_82_n6282), .A2(u5_mult_82_n6283), 
        .A3(u5_mult_82_n6284), .ZN(u5_mult_82_CARRYB_27__29_) );
  NAND2_X2 u5_mult_82_U3544 ( .A1(u5_mult_82_ab_12__43_), .A2(
        u5_mult_82_SUMB_11__44_), .ZN(u5_mult_82_n5781) );
  NAND2_X2 u5_mult_82_U3543 ( .A1(u5_mult_82_ab_51__19_), .A2(u5_mult_82_n2715), .ZN(u5_mult_82_n4911) );
  XNOR2_X2 u5_mult_82_U3542 ( .A(u5_mult_82_CARRYB_42__4_), .B(
        u5_mult_82_ab_43__4_), .ZN(u5_mult_82_n687) );
  XNOR2_X2 u5_mult_82_U3541 ( .A(u5_mult_82_n3707), .B(u5_mult_82_n687), .ZN(
        u5_mult_82_SUMB_43__4_) );
  XNOR2_X2 u5_mult_82_U3540 ( .A(u5_mult_82_ab_12__32_), .B(
        u5_mult_82_CARRYB_11__32_), .ZN(u5_mult_82_n686) );
  XNOR2_X2 u5_mult_82_U3539 ( .A(u5_mult_82_n686), .B(u5_mult_82_SUMB_11__33_), 
        .ZN(u5_mult_82_SUMB_12__32_) );
  INV_X8 u5_mult_82_U3538 ( .A(u5_mult_82_n6512), .ZN(u5_mult_82_SUMB_1__51_)
         );
  NAND2_X2 u5_mult_82_U3537 ( .A1(u5_mult_82_ab_25__20_), .A2(
        u5_mult_82_CARRYB_24__20_), .ZN(u5_mult_82_n5693) );
  NAND2_X2 u5_mult_82_U3536 ( .A1(u5_mult_82_CARRYB_39__17_), .A2(
        u5_mult_82_SUMB_39__18_), .ZN(u5_mult_82_n5193) );
  XNOR2_X2 u5_mult_82_U3535 ( .A(u5_mult_82_n685), .B(u5_mult_82_SUMB_50__20_), 
        .ZN(u5_mult_82_SUMB_51__19_) );
  NAND2_X2 u5_mult_82_U3534 ( .A1(u5_mult_82_ab_40__13_), .A2(
        u5_mult_82_SUMB_39__14_), .ZN(u5_mult_82_n1910) );
  NAND2_X2 u5_mult_82_U3533 ( .A1(u5_mult_82_CARRYB_7__30_), .A2(
        u5_mult_82_SUMB_7__31_), .ZN(u5_mult_82_n2207) );
  NAND2_X2 u5_mult_82_U3532 ( .A1(u5_mult_82_ab_21__9_), .A2(
        u5_mult_82_CARRYB_20__9_), .ZN(u5_mult_82_n3726) );
  INV_X1 u5_mult_82_U3531 ( .A(u5_mult_82_n1603), .ZN(u5_mult_82_n1225) );
  NAND2_X1 u5_mult_82_U3530 ( .A1(u5_mult_82_n1390), .A2(
        u5_mult_82_SUMB_9__28_), .ZN(u5_mult_82_n3451) );
  NAND2_X1 u5_mult_82_U3529 ( .A1(u5_mult_82_ab_10__27_), .A2(
        u5_mult_82_SUMB_9__28_), .ZN(u5_mult_82_n3450) );
  NAND2_X2 u5_mult_82_U3528 ( .A1(u5_mult_82_ab_33__8_), .A2(
        u5_mult_82_SUMB_32__9_), .ZN(u5_mult_82_n3739) );
  NAND2_X2 u5_mult_82_U3527 ( .A1(u5_mult_82_CARRYB_32__8_), .A2(
        u5_mult_82_SUMB_32__9_), .ZN(u5_mult_82_n3740) );
  NAND2_X2 u5_mult_82_U3526 ( .A1(u5_mult_82_ab_37__5_), .A2(
        u5_mult_82_SUMB_36__6_), .ZN(u5_mult_82_n4105) );
  NAND2_X2 u5_mult_82_U3525 ( .A1(u5_mult_82_ab_40__3_), .A2(
        u5_mult_82_SUMB_39__4_), .ZN(u5_mult_82_n2669) );
  NAND2_X2 u5_mult_82_U3524 ( .A1(u5_mult_82_ab_39__34_), .A2(
        u5_mult_82_SUMB_38__35_), .ZN(u5_mult_82_n3936) );
  NAND3_X2 u5_mult_82_U3523 ( .A1(u5_mult_82_n2208), .A2(u5_mult_82_n2209), 
        .A3(u5_mult_82_n2210), .ZN(u5_mult_82_CARRYB_9__29_) );
  NAND2_X2 u5_mult_82_U3522 ( .A1(u5_mult_82_ab_45__4_), .A2(
        u5_mult_82_CARRYB_44__4_), .ZN(u5_mult_82_n6026) );
  NAND3_X4 u5_mult_82_U3521 ( .A1(u5_mult_82_n5821), .A2(u5_mult_82_n5822), 
        .A3(u5_mult_82_n5823), .ZN(u5_mult_82_CARRYB_41__6_) );
  XNOR2_X2 u5_mult_82_U3520 ( .A(u5_mult_82_SUMB_34__34_), .B(
        u5_mult_82_ab_35__33_), .ZN(u5_mult_82_n1775) );
  NAND2_X2 u5_mult_82_U3519 ( .A1(u5_mult_82_ab_25__15_), .A2(
        u5_mult_82_CARRYB_24__15_), .ZN(u5_mult_82_n1017) );
  INV_X4 u5_mult_82_U3518 ( .A(u5_mult_82_n684), .ZN(u5_mult_82_n3891) );
  XNOR2_X2 u5_mult_82_U3517 ( .A(u5_mult_82_ab_17__19_), .B(
        u5_mult_82_CARRYB_16__19_), .ZN(u5_mult_82_n684) );
  NAND2_X2 u5_mult_82_U3516 ( .A1(u5_mult_82_ab_2__50_), .A2(
        u5_mult_82_SUMB_1__51_), .ZN(u5_mult_82_n3505) );
  NAND2_X2 u5_mult_82_U3515 ( .A1(u5_mult_82_ab_37__35_), .A2(
        u5_mult_82_SUMB_36__36_), .ZN(u5_mult_82_n5125) );
  NAND3_X4 u5_mult_82_U3514 ( .A1(u5_mult_82_n3504), .A2(u5_mult_82_n3505), 
        .A3(u5_mult_82_n3506), .ZN(u5_mult_82_CARRYB_2__50_) );
  NAND2_X2 u5_mult_82_U3513 ( .A1(u5_mult_82_CARRYB_43__31_), .A2(
        u5_mult_82_SUMB_43__32_), .ZN(u5_mult_82_n3023) );
  XOR2_X2 u5_mult_82_U3512 ( .A(u5_mult_82_CARRYB_7__40_), .B(u5_mult_82_n857), 
        .Z(u5_mult_82_n683) );
  XNOR2_X2 u5_mult_82_U3511 ( .A(u5_mult_82_n683), .B(u5_mult_82_SUMB_7__41_), 
        .ZN(u5_mult_82_SUMB_8__40_) );
  NAND2_X2 u5_mult_82_U3510 ( .A1(u5_mult_82_ab_10__35_), .A2(
        u5_mult_82_SUMB_9__36_), .ZN(u5_mult_82_n5700) );
  INV_X4 u5_mult_82_U3509 ( .A(u5_mult_82_n6395), .ZN(u5_mult_82_CLA_SUM[61])
         );
  NAND2_X2 u5_mult_82_U3508 ( .A1(u5_mult_82_ab_40__17_), .A2(
        u5_mult_82_SUMB_39__18_), .ZN(u5_mult_82_n5192) );
  XNOR2_X2 u5_mult_82_U3507 ( .A(u5_mult_82_n5344), .B(u5_mult_82_n1492), .ZN(
        u5_mult_82_SUMB_46__18_) );
  NAND2_X2 u5_mult_82_U3506 ( .A1(u5_mult_82_CARRYB_40__2_), .A2(
        u5_mult_82_SUMB_40__3_), .ZN(u5_mult_82_n2672) );
  NAND2_X2 u5_mult_82_U3505 ( .A1(u5_mult_82_ab_3__28_), .A2(
        u5_mult_82_CARRYB_2__28_), .ZN(u5_mult_82_n3812) );
  NOR2_X1 u5_mult_82_U3504 ( .A1(u5_mult_82_net64487), .A2(u5_mult_82_net65517), .ZN(u5_mult_82_ab_34__12_) );
  NOR2_X1 u5_mult_82_U3503 ( .A1(u5_mult_82_net64561), .A2(u5_mult_82_n6636), 
        .ZN(u5_mult_82_ab_22__16_) );
  NOR2_X2 u5_mult_82_U3502 ( .A1(u5_mult_82_net64561), .A2(u5_mult_82_n6643), 
        .ZN(u5_mult_82_ab_24__16_) );
  NAND3_X2 u5_mult_82_U3501 ( .A1(u5_mult_82_n680), .A2(u5_mult_82_n681), .A3(
        u5_mult_82_n682), .ZN(u5_mult_82_CARRYB_2__28_) );
  NAND2_X1 u5_mult_82_U3500 ( .A1(u5_mult_82_ab_2__28_), .A2(
        u5_mult_82_SUMB_1__29_), .ZN(u5_mult_82_n682) );
  NAND2_X2 u5_mult_82_U3499 ( .A1(u5_mult_82_ab_2__28_), .A2(u5_mult_82_n470), 
        .ZN(u5_mult_82_n681) );
  NAND2_X1 u5_mult_82_U3498 ( .A1(u5_mult_82_SUMB_1__29_), .A2(u5_mult_82_n470), .ZN(u5_mult_82_n680) );
  XOR2_X2 u5_mult_82_U3497 ( .A(u5_mult_82_n470), .B(u5_mult_82_n679), .Z(
        u5_mult_82_SUMB_2__28_) );
  XOR2_X2 u5_mult_82_U3496 ( .A(u5_mult_82_SUMB_1__29_), .B(
        u5_mult_82_ab_2__28_), .Z(u5_mult_82_n679) );
  NAND3_X2 u5_mult_82_U3495 ( .A1(u5_mult_82_n676), .A2(u5_mult_82_n677), .A3(
        u5_mult_82_n678), .ZN(u5_mult_82_CARRYB_34__12_) );
  NAND2_X1 u5_mult_82_U3494 ( .A1(u5_mult_82_ab_34__12_), .A2(
        u5_mult_82_SUMB_33__13_), .ZN(u5_mult_82_n678) );
  NAND2_X2 u5_mult_82_U3493 ( .A1(u5_mult_82_ab_34__12_), .A2(
        u5_mult_82_CARRYB_33__12_), .ZN(u5_mult_82_n677) );
  NAND2_X1 u5_mult_82_U3492 ( .A1(u5_mult_82_SUMB_33__13_), .A2(
        u5_mult_82_CARRYB_33__12_), .ZN(u5_mult_82_n676) );
  XOR2_X2 u5_mult_82_U3491 ( .A(u5_mult_82_CARRYB_33__12_), .B(u5_mult_82_n675), .Z(u5_mult_82_SUMB_34__12_) );
  XOR2_X2 u5_mult_82_U3490 ( .A(u5_mult_82_SUMB_33__13_), .B(
        u5_mult_82_ab_34__12_), .Z(u5_mult_82_n675) );
  NAND3_X2 u5_mult_82_U3489 ( .A1(u5_mult_82_n672), .A2(u5_mult_82_n673), .A3(
        u5_mult_82_n674), .ZN(u5_mult_82_CARRYB_22__16_) );
  NAND2_X1 u5_mult_82_U3488 ( .A1(u5_mult_82_ab_22__16_), .A2(
        u5_mult_82_CARRYB_21__16_), .ZN(u5_mult_82_n674) );
  NAND2_X2 u5_mult_82_U3487 ( .A1(u5_mult_82_ab_22__16_), .A2(
        u5_mult_82_SUMB_21__17_), .ZN(u5_mult_82_n673) );
  NAND2_X1 u5_mult_82_U3486 ( .A1(u5_mult_82_CARRYB_21__16_), .A2(
        u5_mult_82_SUMB_21__17_), .ZN(u5_mult_82_n672) );
  XOR2_X2 u5_mult_82_U3485 ( .A(u5_mult_82_SUMB_21__17_), .B(u5_mult_82_n671), 
        .Z(u5_mult_82_SUMB_22__16_) );
  XOR2_X2 u5_mult_82_U3484 ( .A(u5_mult_82_CARRYB_21__16_), .B(
        u5_mult_82_ab_22__16_), .Z(u5_mult_82_n671) );
  INV_X4 u5_mult_82_U3483 ( .A(u5_mult_82_n5257), .ZN(u5_mult_82_n668) );
  INV_X1 u5_mult_82_U3482 ( .A(u5_mult_82_CARRYB_42__8_), .ZN(u5_mult_82_n667)
         );
  NAND2_X4 u5_mult_82_U3481 ( .A1(u5_mult_82_n669), .A2(u5_mult_82_n670), .ZN(
        u5_mult_82_SUMB_43__8_) );
  NAND2_X4 u5_mult_82_U3480 ( .A1(u5_mult_82_n668), .A2(u5_mult_82_n667), .ZN(
        u5_mult_82_n670) );
  NAND2_X2 u5_mult_82_U3479 ( .A1(u5_mult_82_CARRYB_42__8_), .A2(
        u5_mult_82_n5257), .ZN(u5_mult_82_n669) );
  NAND3_X2 u5_mult_82_U3478 ( .A1(u5_mult_82_n664), .A2(u5_mult_82_n665), .A3(
        u5_mult_82_n666), .ZN(u5_mult_82_CARRYB_14__21_) );
  NAND2_X1 u5_mult_82_U3477 ( .A1(u5_mult_82_CARRYB_13__21_), .A2(
        u5_mult_82_SUMB_13__22_), .ZN(u5_mult_82_n666) );
  NAND2_X1 u5_mult_82_U3476 ( .A1(u5_mult_82_ab_14__21_), .A2(
        u5_mult_82_SUMB_13__22_), .ZN(u5_mult_82_n665) );
  NAND2_X1 u5_mult_82_U3475 ( .A1(u5_mult_82_ab_14__21_), .A2(
        u5_mult_82_CARRYB_13__21_), .ZN(u5_mult_82_n664) );
  NAND3_X2 u5_mult_82_U3474 ( .A1(u5_mult_82_n661), .A2(u5_mult_82_n662), .A3(
        u5_mult_82_n663), .ZN(u5_mult_82_CARRYB_13__22_) );
  NAND2_X2 u5_mult_82_U3473 ( .A1(u5_mult_82_CARRYB_12__22_), .A2(
        u5_mult_82_SUMB_12__23_), .ZN(u5_mult_82_n663) );
  NAND2_X2 u5_mult_82_U3472 ( .A1(u5_mult_82_ab_13__22_), .A2(
        u5_mult_82_SUMB_12__23_), .ZN(u5_mult_82_n662) );
  NAND2_X2 u5_mult_82_U3471 ( .A1(u5_mult_82_ab_13__22_), .A2(
        u5_mult_82_CARRYB_12__22_), .ZN(u5_mult_82_n661) );
  XOR2_X2 u5_mult_82_U3470 ( .A(u5_mult_82_n660), .B(u5_mult_82_n392), .Z(
        u5_mult_82_SUMB_14__21_) );
  XOR2_X2 u5_mult_82_U3469 ( .A(u5_mult_82_ab_14__21_), .B(
        u5_mult_82_CARRYB_13__21_), .Z(u5_mult_82_n660) );
  XOR2_X2 u5_mult_82_U3468 ( .A(u5_mult_82_n659), .B(u5_mult_82_SUMB_12__23_), 
        .Z(u5_mult_82_SUMB_13__22_) );
  XOR2_X2 u5_mult_82_U3467 ( .A(u5_mult_82_CARRYB_12__22_), .B(
        u5_mult_82_ab_13__22_), .Z(u5_mult_82_n659) );
  NAND3_X2 u5_mult_82_U3466 ( .A1(u5_mult_82_n656), .A2(u5_mult_82_n657), .A3(
        u5_mult_82_n658), .ZN(u5_mult_82_CARRYB_24__16_) );
  NAND2_X1 u5_mult_82_U3465 ( .A1(u5_mult_82_ab_24__16_), .A2(
        u5_mult_82_SUMB_23__17_), .ZN(u5_mult_82_n658) );
  NAND2_X2 u5_mult_82_U3464 ( .A1(u5_mult_82_ab_24__16_), .A2(
        u5_mult_82_CARRYB_23__16_), .ZN(u5_mult_82_n657) );
  NAND2_X1 u5_mult_82_U3463 ( .A1(u5_mult_82_SUMB_23__17_), .A2(
        u5_mult_82_CARRYB_23__16_), .ZN(u5_mult_82_n656) );
  XOR2_X2 u5_mult_82_U3462 ( .A(u5_mult_82_CARRYB_23__16_), .B(u5_mult_82_n655), .Z(u5_mult_82_SUMB_24__16_) );
  XOR2_X2 u5_mult_82_U3461 ( .A(u5_mult_82_SUMB_23__17_), .B(
        u5_mult_82_ab_24__16_), .Z(u5_mult_82_n655) );
  NAND2_X2 u5_mult_82_U3460 ( .A1(u5_mult_82_ab_31__13_), .A2(
        u5_mult_82_SUMB_30__14_), .ZN(u5_mult_82_n653) );
  XOR2_X2 u5_mult_82_U3459 ( .A(u5_mult_82_SUMB_30__14_), .B(u5_mult_82_n651), 
        .Z(u5_mult_82_SUMB_31__13_) );
  XNOR2_X2 u5_mult_82_U3458 ( .A(u5_mult_82_ab_36__29_), .B(
        u5_mult_82_CARRYB_35__29_), .ZN(u5_mult_82_n650) );
  XNOR2_X2 u5_mult_82_U3457 ( .A(u5_mult_82_n650), .B(u5_mult_82_SUMB_35__30_), 
        .ZN(u5_mult_82_SUMB_36__29_) );
  XOR2_X2 u5_mult_82_U3456 ( .A(u5_mult_82_n3175), .B(u5_mult_82_SUMB_34__5_), 
        .Z(u5_mult_82_SUMB_35__4_) );
  XOR2_X2 u5_mult_82_U3455 ( .A(u5_mult_82_CARRYB_27__5_), .B(
        u5_mult_82_ab_28__5_), .Z(u5_mult_82_n4053) );
  XOR2_X2 u5_mult_82_U3454 ( .A(u5_mult_82_CARRYB_18__11_), .B(
        u5_mult_82_ab_19__11_), .Z(u5_mult_82_n3322) );
  NAND2_X2 u5_mult_82_U3453 ( .A1(u5_mult_82_ab_41__2_), .A2(
        u5_mult_82_SUMB_40__3_), .ZN(u5_mult_82_n2671) );
  XNOR2_X2 u5_mult_82_U3452 ( .A(u5_mult_82_n649), .B(
        u5_mult_82_CARRYB_16__17_), .ZN(u5_mult_82_n4107) );
  XNOR2_X2 u5_mult_82_U3451 ( .A(u5_mult_82_n2740), .B(u5_mult_82_SUMB_12__33_), .ZN(u5_mult_82_SUMB_13__32_) );
  NAND2_X2 u5_mult_82_U3450 ( .A1(u5_mult_82_SUMB_46__11_), .A2(
        u5_mult_82_CARRYB_46__10_), .ZN(u5_mult_82_n4179) );
  CLKBUF_X3 u5_mult_82_U3449 ( .A(u5_mult_82_SUMB_27__31_), .Z(
        u5_mult_82_n1851) );
  XNOR2_X2 u5_mult_82_U3448 ( .A(u5_mult_82_ab_30__29_), .B(
        u5_mult_82_CARRYB_29__29_), .ZN(u5_mult_82_n1734) );
  NAND2_X2 u5_mult_82_U3447 ( .A1(u5_mult_82_ab_43__20_), .A2(
        u5_mult_82_CARRYB_42__20_), .ZN(u5_mult_82_n4162) );
  NAND2_X2 u5_mult_82_U3446 ( .A1(u5_mult_82_ab_43__20_), .A2(
        u5_mult_82_SUMB_42__21_), .ZN(u5_mult_82_n4161) );
  XOR2_X2 u5_mult_82_U3445 ( .A(u5_mult_82_n1928), .B(u5_mult_82_SUMB_2__47_), 
        .Z(u5_mult_82_SUMB_3__46_) );
  NAND2_X2 u5_mult_82_U3444 ( .A1(u5_mult_82_n5674), .A2(
        u5_mult_82_SUMB_47__19_), .ZN(u5_mult_82_n4158) );
  NAND2_X2 u5_mult_82_U3443 ( .A1(u5_mult_82_CARRYB_43__10_), .A2(
        u5_mult_82_SUMB_43__11_), .ZN(u5_mult_82_net79318) );
  NAND2_X2 u5_mult_82_U3442 ( .A1(u5_mult_82_ab_39__14_), .A2(
        u5_mult_82_CARRYB_38__14_), .ZN(u5_mult_82_net82676) );
  XNOR2_X2 u5_mult_82_U3441 ( .A(u5_mult_82_ab_16__16_), .B(
        u5_mult_82_CARRYB_15__16_), .ZN(u5_mult_82_n648) );
  XNOR2_X2 u5_mult_82_U3440 ( .A(u5_mult_82_n648), .B(u5_mult_82_n1651), .ZN(
        u5_mult_82_SUMB_16__16_) );
  XOR2_X2 u5_mult_82_U3439 ( .A(u5_mult_82_n3960), .B(
        u5_mult_82_CARRYB_50__18_), .Z(u5_mult_82_n647) );
  XNOR2_X2 u5_mult_82_U3438 ( .A(u5_mult_82_SUMB_50__19_), .B(u5_mult_82_n647), 
        .ZN(u5_mult_82_SUMB_51__18_) );
  XNOR2_X2 u5_mult_82_U3437 ( .A(u5_mult_82_CARRYB_23__10_), .B(
        u5_mult_82_n2416), .ZN(u5_mult_82_n4115) );
  XNOR2_X2 u5_mult_82_U3436 ( .A(u5_mult_82_ab_30__8_), .B(
        u5_mult_82_CARRYB_29__8_), .ZN(u5_mult_82_n646) );
  XNOR2_X2 u5_mult_82_U3435 ( .A(u5_mult_82_n646), .B(u5_mult_82_SUMB_29__9_), 
        .ZN(u5_mult_82_SUMB_30__8_) );
  XNOR2_X2 u5_mult_82_U3434 ( .A(u5_mult_82_CARRYB_37__5_), .B(
        u5_mult_82_ab_38__5_), .ZN(u5_mult_82_n645) );
  XNOR2_X2 u5_mult_82_U3433 ( .A(u5_mult_82_SUMB_37__6_), .B(u5_mult_82_n645), 
        .ZN(u5_mult_82_SUMB_38__5_) );
  NAND3_X4 u5_mult_82_U3432 ( .A1(u5_mult_82_n3420), .A2(u5_mult_82_n3421), 
        .A3(u5_mult_82_n3422), .ZN(u5_mult_82_CARRYB_14__14_) );
  NAND2_X2 u5_mult_82_U3431 ( .A1(u5_mult_82_ab_39__13_), .A2(
        u5_mult_82_CARRYB_38__13_), .ZN(u5_mult_82_n3991) );
  NAND2_X2 u5_mult_82_U3430 ( .A1(u5_mult_82_ab_44__10_), .A2(
        u5_mult_82_SUMB_43__11_), .ZN(u5_mult_82_net79317) );
  NAND2_X4 u5_mult_82_U3429 ( .A1(u5_mult_82_SUMB_48__18_), .A2(
        u5_mult_82_ab_49__17_), .ZN(u5_mult_82_n3638) );
  NAND2_X4 u5_mult_82_U3428 ( .A1(u5_mult_82_ab_47__18_), .A2(
        u5_mult_82_SUMB_46__19_), .ZN(u5_mult_82_n5659) );
  XNOR2_X2 u5_mult_82_U3427 ( .A(u5_mult_82_n1579), .B(u5_mult_82_SUMB_47__20_), .ZN(u5_mult_82_SUMB_48__19_) );
  XNOR2_X2 u5_mult_82_U3426 ( .A(u5_mult_82_CARRYB_23__38_), .B(
        u5_mult_82_ab_24__38_), .ZN(u5_mult_82_n644) );
  XNOR2_X2 u5_mult_82_U3425 ( .A(u5_mult_82_SUMB_23__39_), .B(u5_mult_82_n644), 
        .ZN(u5_mult_82_SUMB_24__38_) );
  NAND3_X4 u5_mult_82_U3424 ( .A1(u5_mult_82_n5058), .A2(u5_mult_82_n5059), 
        .A3(u5_mult_82_n5060), .ZN(u5_mult_82_CARRYB_21__29_) );
  NAND2_X4 u5_mult_82_U3423 ( .A1(u5_mult_82_ab_15__34_), .A2(u5_mult_82_n1616), .ZN(u5_mult_82_n4017) );
  XNOR2_X2 u5_mult_82_U3422 ( .A(u5_mult_82_CARRYB_21__12_), .B(
        u5_mult_82_ab_22__12_), .ZN(u5_mult_82_n2171) );
  XNOR2_X2 u5_mult_82_U3421 ( .A(u5_mult_82_CARRYB_23__23_), .B(
        u5_mult_82_ab_24__23_), .ZN(u5_mult_82_n643) );
  NAND2_X2 u5_mult_82_U3420 ( .A1(u5_mult_82_CARRYB_49__17_), .A2(
        u5_mult_82_SUMB_49__18_), .ZN(u5_mult_82_n4400) );
  XNOR2_X2 u5_mult_82_U3419 ( .A(u5_mult_82_ab_23__8_), .B(
        u5_mult_82_SUMB_22__9_), .ZN(u5_mult_82_n642) );
  XNOR2_X2 u5_mult_82_U3418 ( .A(u5_mult_82_n642), .B(u5_mult_82_CARRYB_22__8_), .ZN(u5_mult_82_SUMB_23__8_) );
  NAND2_X2 u5_mult_82_U3417 ( .A1(u5_mult_82_ab_27__25_), .A2(u5_mult_82_n733), 
        .ZN(u5_mult_82_n6183) );
  NAND2_X2 u5_mult_82_U3416 ( .A1(u5_mult_82_CARRYB_28__24_), .A2(
        u5_mult_82_SUMB_28__25_), .ZN(u5_mult_82_n6295) );
  XNOR2_X2 u5_mult_82_U3415 ( .A(u5_mult_82_n944), .B(u5_mult_82_SUMB_11__34_), 
        .ZN(u5_mult_82_SUMB_12__33_) );
  NAND2_X2 u5_mult_82_U3414 ( .A1(u5_mult_82_CARRYB_9__26_), .A2(
        u5_mult_82_n382), .ZN(u5_mult_82_n4371) );
  NAND2_X2 u5_mult_82_U3413 ( .A1(u5_mult_82_ab_22__18_), .A2(
        u5_mult_82_SUMB_21__19_), .ZN(u5_mult_82_n4738) );
  NAND2_X2 u5_mult_82_U3412 ( .A1(u5_mult_82_CARRYB_16__42_), .A2(
        u5_mult_82_SUMB_16__43_), .ZN(u5_mult_82_n2732) );
  XNOR2_X1 u5_mult_82_U3411 ( .A(u5_mult_82_ab_20__42_), .B(
        u5_mult_82_CARRYB_19__42_), .ZN(u5_mult_82_n5554) );
  NAND2_X1 u5_mult_82_U3410 ( .A1(u5_mult_82_CARRYB_28__36_), .A2(
        u5_mult_82_SUMB_28__37_), .ZN(u5_mult_82_n5669) );
  XNOR2_X2 u5_mult_82_U3409 ( .A(u5_mult_82_n1722), .B(u5_mult_82_n697), .ZN(
        u5_mult_82_SUMB_45__14_) );
  XNOR2_X2 u5_mult_82_U3408 ( .A(u5_mult_82_n5945), .B(u5_mult_82_SUMB_32__32_), .ZN(u5_mult_82_n641) );
  INV_X4 u5_mult_82_U3407 ( .A(u5_mult_82_n640), .ZN(u5_mult_82_SUMB_34__30_)
         );
  XNOR2_X2 u5_mult_82_U3406 ( .A(u5_mult_82_n3771), .B(u5_mult_82_n641), .ZN(
        u5_mult_82_n640) );
  XNOR2_X2 u5_mult_82_U3405 ( .A(u5_mult_82_ab_40__32_), .B(
        u5_mult_82_CARRYB_39__32_), .ZN(u5_mult_82_n639) );
  XNOR2_X2 u5_mult_82_U3404 ( .A(u5_mult_82_n638), .B(u5_mult_82_SUMB_36__35_), 
        .ZN(u5_mult_82_SUMB_37__34_) );
  XNOR2_X2 u5_mult_82_U3403 ( .A(u5_mult_82_SUMB_36__39_), .B(
        u5_mult_82_ab_37__38_), .ZN(u5_mult_82_n637) );
  XNOR2_X2 u5_mult_82_U3402 ( .A(u5_mult_82_CARRYB_36__38_), .B(
        u5_mult_82_n637), .ZN(u5_mult_82_SUMB_37__38_) );
  XNOR2_X2 u5_mult_82_U3401 ( .A(u5_mult_82_ab_32__41_), .B(
        u5_mult_82_CARRYB_31__41_), .ZN(u5_mult_82_n636) );
  XNOR2_X2 u5_mult_82_U3400 ( .A(u5_mult_82_n636), .B(u5_mult_82_SUMB_31__42_), 
        .ZN(u5_mult_82_SUMB_32__41_) );
  NOR2_X1 u5_mult_82_U3399 ( .A1(u5_mult_82_n7006), .A2(u5_mult_82_net66107), 
        .ZN(u5_mult_82_ab_1__48_) );
  INV_X4 u5_mult_82_U3398 ( .A(u5_mult_82_n1716), .ZN(u5_mult_82_n1717) );
  XNOR2_X2 u5_mult_82_U3397 ( .A(u5_mult_82_ab_15__39_), .B(
        u5_mult_82_CARRYB_14__39_), .ZN(u5_mult_82_n635) );
  XNOR2_X2 u5_mult_82_U3396 ( .A(u5_mult_82_n635), .B(u5_mult_82_SUMB_14__40_), 
        .ZN(u5_mult_82_SUMB_15__39_) );
  CLKBUF_X2 u5_mult_82_U3395 ( .A(u5_mult_82_SUMB_13__40_), .Z(u5_mult_82_n634) );
  NAND2_X1 u5_mult_82_U3394 ( .A1(u5_mult_82_ab_40__3_), .A2(
        u5_mult_82_CARRYB_39__3_), .ZN(u5_mult_82_n2668) );
  NAND2_X1 u5_mult_82_U3393 ( .A1(u5_mult_82_CARRYB_39__3_), .A2(
        u5_mult_82_SUMB_39__4_), .ZN(u5_mult_82_n2670) );
  NAND2_X1 u5_mult_82_U3392 ( .A1(u5_mult_82_ab_25__11_), .A2(
        u5_mult_82_SUMB_24__12_), .ZN(u5_mult_82_n2822) );
  NAND2_X1 u5_mult_82_U3391 ( .A1(u5_mult_82_CARRYB_24__11_), .A2(
        u5_mult_82_SUMB_24__12_), .ZN(u5_mult_82_n2823) );
  NOR2_X2 u5_mult_82_U3390 ( .A1(u5_mult_82_n6803), .A2(u5_mult_82_net66107), 
        .ZN(u5_mult_82_ab_1__44_) );
  NOR2_X2 u5_mult_82_U3389 ( .A1(u5_mult_82_n6783), .A2(u5_mult_82_net66107), 
        .ZN(u5_mult_82_ab_1__47_) );
  NAND3_X2 u5_mult_82_U3388 ( .A1(u5_mult_82_n5345), .A2(u5_mult_82_n5346), 
        .A3(u5_mult_82_n5347), .ZN(u5_mult_82_CARRYB_46__18_) );
  CLKBUF_X3 u5_mult_82_U3387 ( .A(u5_mult_82_CARRYB_36__5_), .Z(
        u5_mult_82_n633) );
  XOR2_X1 u5_mult_82_U3386 ( .A(u5_mult_82_SUMB_11__18_), .B(u5_mult_82_n1969), 
        .Z(u5_mult_82_SUMB_12__17_) );
  XNOR2_X2 u5_mult_82_U3385 ( .A(u5_mult_82_ab_45__10_), .B(
        u5_mult_82_CARRYB_44__10_), .ZN(u5_mult_82_n1643) );
  NAND2_X2 u5_mult_82_U3384 ( .A1(u5_mult_82_ab_39__15_), .A2(
        u5_mult_82_CARRYB_38__15_), .ZN(u5_mult_82_n5526) );
  NAND3_X2 u5_mult_82_U3383 ( .A1(u5_mult_82_n5683), .A2(u5_mult_82_n5684), 
        .A3(u5_mult_82_n5685), .ZN(u5_mult_82_CARRYB_15__30_) );
  INV_X2 u5_mult_82_U3382 ( .A(u5_mult_82_CARRYB_30__28_), .ZN(
        u5_mult_82_n1627) );
  NOR2_X2 u5_mult_82_U3381 ( .A1(u5_mult_82_n6803), .A2(u5_mult_82_net65277), 
        .ZN(u5_mult_82_ab_47__44_) );
  NOR2_X2 u5_mult_82_U3380 ( .A1(u5_mult_82_n6803), .A2(u5_mult_82_n6740), 
        .ZN(u5_mult_82_ab_46__44_) );
  NOR2_X2 u5_mult_82_U3379 ( .A1(u5_mult_82_n6803), .A2(u5_mult_82_net65313), 
        .ZN(u5_mult_82_ab_45__44_) );
  NOR2_X2 u5_mult_82_U3378 ( .A1(u5_mult_82_n6803), .A2(u5_mult_82_net65373), 
        .ZN(u5_mult_82_ab_42__44_) );
  NOR2_X2 u5_mult_82_U3377 ( .A1(u5_mult_82_net64217), .A2(u5_mult_82_n6803), 
        .ZN(u5_mult_82_ab_0__44_) );
  NAND3_X2 u5_mult_82_U3376 ( .A1(u5_mult_82_n3130), .A2(u5_mult_82_n3129), 
        .A3(u5_mult_82_n3128), .ZN(u5_mult_82_CARRYB_8__47_) );
  XNOR2_X2 u5_mult_82_U3375 ( .A(u5_mult_82_n1458), .B(
        u5_mult_82_CARRYB_32__7_), .ZN(u5_mult_82_n3788) );
  INV_X2 u5_mult_82_U3374 ( .A(u5_mult_82_n3108), .ZN(u5_mult_82_n1961) );
  INV_X2 u5_mult_82_U3373 ( .A(u5_mult_82_n6478), .ZN(u5_mult_82_CARRYB_1__26_) );
  XNOR2_X2 u5_mult_82_U3372 ( .A(u5_mult_82_n632), .B(
        u5_mult_82_CARRYB_24__12_), .ZN(u5_mult_82_n2280) );
  XNOR2_X2 u5_mult_82_U3371 ( .A(u5_mult_82_ab_2__26_), .B(u5_mult_82_n6478), 
        .ZN(u5_mult_82_n3182) );
  XOR2_X1 u5_mult_82_U3370 ( .A(u5_mult_82_SUMB_38__1_), .B(u5_mult_82_n4844), 
        .Z(u5_N39) );
  NAND2_X1 u5_mult_82_U3369 ( .A1(u5_mult_82_CARRYB_4__25_), .A2(
        u5_mult_82_SUMB_4__26_), .ZN(u5_mult_82_n2479) );
  NAND2_X1 u5_mult_82_U3368 ( .A1(u5_mult_82_CARRYB_3__26_), .A2(
        u5_mult_82_SUMB_3__27_), .ZN(u5_mult_82_n2476) );
  NAND2_X1 u5_mult_82_U3367 ( .A1(u5_mult_82_ab_4__26_), .A2(
        u5_mult_82_SUMB_3__27_), .ZN(u5_mult_82_n2475) );
  NAND2_X2 u5_mult_82_U3366 ( .A1(u5_mult_82_ab_38__2_), .A2(
        u5_mult_82_CARRYB_37__2_), .ZN(u5_mult_82_n4683) );
  XNOR2_X1 u5_mult_82_U3365 ( .A(u5_mult_82_ab_38__2_), .B(
        u5_mult_82_CARRYB_37__2_), .ZN(u5_mult_82_n1908) );
  NAND2_X2 u5_mult_82_U3364 ( .A1(u5_mult_82_n390), .A2(
        u5_mult_82_CARRYB_36__4_), .ZN(u5_mult_82_n2340) );
  XOR2_X2 u5_mult_82_U3363 ( .A(u5_mult_82_SUMB_20__10_), .B(u5_mult_82_n3723), 
        .Z(u5_mult_82_SUMB_21__9_) );
  XOR2_X1 u5_mult_82_U3362 ( .A(u5_mult_82_CARRYB_20__9_), .B(
        u5_mult_82_ab_21__9_), .Z(u5_mult_82_n3723) );
  XNOR2_X2 u5_mult_82_U3361 ( .A(u5_mult_82_SUMB_22__10_), .B(u5_mult_82_n2417), .ZN(u5_mult_82_SUMB_23__9_) );
  XOR2_X2 u5_mult_82_U3360 ( .A(u5_mult_82_n3404), .B(u5_mult_82_SUMB_26__8_), 
        .Z(u5_mult_82_SUMB_27__7_) );
  NAND3_X2 u5_mult_82_U3359 ( .A1(u5_mult_82_n3474), .A2(u5_mult_82_n3475), 
        .A3(u5_mult_82_n3476), .ZN(u5_mult_82_CARRYB_16__19_) );
  NAND2_X2 u5_mult_82_U3358 ( .A1(u5_mult_82_ab_28__13_), .A2(u5_mult_82_n394), 
        .ZN(u5_mult_82_n2596) );
  NAND3_X2 u5_mult_82_U3357 ( .A1(u5_mult_82_n4830), .A2(u5_mult_82_n4831), 
        .A3(u5_mult_82_n4832), .ZN(u5_mult_82_CARRYB_25__14_) );
  NAND3_X4 u5_mult_82_U3356 ( .A1(u5_mult_82_n2561), .A2(u5_mult_82_n2562), 
        .A3(u5_mult_82_n2563), .ZN(u5_mult_82_CARRYB_23__9_) );
  NOR2_X2 u5_mult_82_U3355 ( .A1(u5_mult_82_n6759), .A2(u5_mult_82_net66107), 
        .ZN(u5_mult_82_ab_1__51_) );
  NOR2_X2 u5_mult_82_U3354 ( .A1(u5_mult_82_n6826), .A2(u5_mult_82_net66107), 
        .ZN(u5_mult_82_n3280) );
  CLKBUF_X3 u5_mult_82_U3353 ( .A(u5_mult_82_CARRYB_17__13_), .Z(
        u5_mult_82_n630) );
  BUF_X8 u5_mult_82_U3352 ( .A(u5_mult_82_n1481), .Z(u5_mult_82_n1587) );
  XNOR2_X1 u5_mult_82_U3351 ( .A(u5_mult_82_SUMB_42__2_), .B(
        u5_mult_82_ab_43__1_), .ZN(u5_mult_82_n629) );
  XNOR2_X2 u5_mult_82_U3350 ( .A(u5_mult_82_n1653), .B(u5_mult_82_n629), .ZN(
        u5_mult_82_SUMB_43__1_) );
  XOR2_X1 u5_mult_82_U3349 ( .A(u5_mult_82_CARRYB_52__0_), .B(
        u5_mult_82_SUMB_52__1_), .Z(u5_N53) );
  INV_X4 u5_mult_82_U3348 ( .A(u5_mult_82_n7012), .ZN(u5_mult_82_n6854) );
  XOR2_X2 u5_mult_82_U3347 ( .A(u5_mult_82_n1402), .B(u5_mult_82_n3423), .Z(
        u5_N50) );
  XNOR2_X2 u5_mult_82_U3346 ( .A(u5_mult_82_n4080), .B(u5_mult_82_SUMB_47__2_), 
        .ZN(u5_mult_82_n5813) );
  INV_X4 u5_mult_82_U3345 ( .A(u5_mult_82_n4789), .ZN(u5_mult_82_n4686) );
  XOR2_X1 u5_mult_82_U3344 ( .A(u5_mult_82_CARRYB_38__0_), .B(
        u5_mult_82_ab_39__0_), .Z(u5_mult_82_n4844) );
  NAND2_X2 u5_mult_82_U3343 ( .A1(u5_mult_82_ab_39__0_), .A2(
        u5_mult_82_CARRYB_38__0_), .ZN(u5_mult_82_n4847) );
  NAND2_X1 u5_mult_82_U3342 ( .A1(u5_mult_82_CARRYB_38__0_), .A2(
        u5_mult_82_SUMB_38__1_), .ZN(u5_mult_82_n4845) );
  NAND2_X2 u5_mult_82_U3341 ( .A1(u5_mult_82_SUMB_37__3_), .A2(
        u5_mult_82_CARRYB_37__2_), .ZN(u5_mult_82_n4685) );
  NAND2_X2 u5_mult_82_U3340 ( .A1(u5_mult_82_SUMB_35__3_), .A2(
        u5_mult_82_CARRYB_35__2_), .ZN(u5_mult_82_n876) );
  XNOR2_X1 u5_mult_82_U3339 ( .A(u5_mult_82_ab_39__1_), .B(
        u5_mult_82_SUMB_38__2_), .ZN(u5_mult_82_n627) );
  XNOR2_X2 u5_mult_82_U3338 ( .A(u5_mult_82_n627), .B(u5_mult_82_CARRYB_38__1_), .ZN(u5_mult_82_SUMB_39__1_) );
  INV_X4 u5_mult_82_U3337 ( .A(u5_mult_82_n6973), .ZN(u5_mult_82_n6975) );
  INV_X4 u5_mult_82_U3336 ( .A(u5_mult_82_n7022), .ZN(u5_mult_82_n6978) );
  INV_X16 u5_mult_82_U3335 ( .A(u5_mult_82_n1272), .ZN(u5_mult_82_net65229) );
  INV_X8 u5_mult_82_U3334 ( .A(u5_mult_82_net57179), .ZN(u5_mult_82_n1272) );
  INV_X4 u5_mult_82_U3333 ( .A(u5_mult_82_n1349), .ZN(u5_mult_82_net65197) );
  XOR2_X1 u5_mult_82_U3332 ( .A(u5_mult_82_ab_1__0_), .B(u5_mult_82_ab_0__1_), 
        .Z(u5_N1) );
  INV_X4 u5_mult_82_U3331 ( .A(u5_mult_82_ab_48__15_), .ZN(u5_mult_82_n5521)
         );
  INV_X16 u5_mult_82_U3330 ( .A(u5_mult_82_n1291), .ZN(u5_mult_82_n1290) );
  INV_X8 u5_mult_82_U3329 ( .A(u5_mult_82_n1287), .ZN(u5_mult_82_n1292) );
  INV_X4 u5_mult_82_U3328 ( .A(u5_mult_82_n1292), .ZN(u5_mult_82_n1291) );
  INV_X8 u5_mult_82_U3327 ( .A(u5_mult_82_n7004), .ZN(u5_mult_82_n6745) );
  INV_X16 u5_mult_82_U3326 ( .A(u5_mult_82_net65277), .ZN(u5_mult_82_net65287)
         );
  INV_X8 u5_mult_82_U3325 ( .A(u5_mult_82_net57182), .ZN(u5_mult_82_net65293)
         );
  INV_X4 u5_mult_82_U3324 ( .A(u5_mult_82_ab_44__4_), .ZN(u5_mult_82_n3992) );
  INV_X2 u5_mult_82_U3323 ( .A(u5_mult_82_ab_41__6_), .ZN(u5_mult_82_n4788) );
  INV_X16 u5_mult_82_U3322 ( .A(u5_mult_82_n1327), .ZN(u5_mult_82_n1326) );
  INV_X8 u5_mult_82_U3321 ( .A(u5_mult_82_n1325), .ZN(u5_mult_82_n1328) );
  INV_X4 u5_mult_82_U3320 ( .A(u5_mult_82_n1328), .ZN(u5_mult_82_n1327) );
  INV_X8 u5_mult_82_U3319 ( .A(u5_mult_82_n1277), .ZN(u5_mult_82_n1280) );
  INV_X8 u5_mult_82_U3318 ( .A(u5_mult_82_n1280), .ZN(u5_mult_82_n1279) );
  INV_X16 u5_mult_82_U3317 ( .A(u5_mult_82_n6690), .ZN(u5_mult_82_n6697) );
  INV_X8 u5_mult_82_U3316 ( .A(u5_mult_82_n7001), .ZN(u5_mult_82_n6691) );
  INV_X8 u5_mult_82_U3315 ( .A(u5_mult_82_n6691), .ZN(u5_mult_82_n6690) );
  INV_X16 u5_mult_82_U3314 ( .A(u5_mult_82_n6706), .ZN(u5_mult_82_n6711) );
  INV_X4 u5_mult_82_U3313 ( .A(u5_mult_82_n7002), .ZN(u5_mult_82_n6705) );
  INV_X16 u5_mult_82_U3312 ( .A(u5_mult_82_n6713), .ZN(u5_mult_82_n6718) );
  INV_X4 u5_mult_82_U3311 ( .A(u5_mult_82_n7003), .ZN(u5_mult_82_n6712) );
  INV_X4 u5_mult_82_U3310 ( .A(u5_mult_82_ab_25__33_), .ZN(u5_mult_82_n5548)
         );
  INV_X4 u5_mult_82_U3309 ( .A(u5_mult_82_ab_18__35_), .ZN(u5_mult_82_n3153)
         );
  INV_X16 u5_mult_82_U3308 ( .A(u5_mult_82_n6593), .ZN(u5_mult_82_n6598) );
  INV_X4 u5_mult_82_U3307 ( .A(u5_mult_82_n6996), .ZN(u5_mult_82_n6592) );
  INV_X16 u5_mult_82_U3306 ( .A(u5_mult_82_n6600), .ZN(u5_mult_82_n6605) );
  INV_X4 u5_mult_82_U3305 ( .A(u5_mult_82_n6997), .ZN(u5_mult_82_n6599) );
  AND2_X2 u5_mult_82_U3304 ( .A1(u5_mult_82_ab_52__52_), .A2(
        u5_mult_82_CARRYB_52__51_), .ZN(u5_mult_82_n624) );
  INV_X16 u5_mult_82_U3303 ( .A(u5_mult_82_n6564), .ZN(u5_mult_82_n6569) );
  INV_X4 u5_mult_82_U3302 ( .A(u5_mult_82_n6995), .ZN(u5_mult_82_n6563) );
  AND2_X2 u5_mult_82_U3301 ( .A1(u5_mult_82_ab_0__5_), .A2(u5_mult_82_ab_1__4_), .ZN(u5_mult_82_n623) );
  INV_X16 u5_mult_82_U3300 ( .A(u5_mult_82_n1261), .ZN(u5_mult_82_net64225) );
  AND2_X4 u5_mult_82_U3299 ( .A1(u5_mult_82_SUMB_52__49_), .A2(
        u5_mult_82_CARRYB_52__48_), .ZN(u5_mult_82_n622) );
  AND2_X4 u5_mult_82_U3298 ( .A1(u5_mult_82_SUMB_52__45_), .A2(
        u5_mult_82_CARRYB_52__44_), .ZN(u5_mult_82_n621) );
  AND2_X4 u5_mult_82_U3297 ( .A1(u5_mult_82_SUMB_52__46_), .A2(
        u5_mult_82_CARRYB_52__45_), .ZN(u5_mult_82_n620) );
  AND2_X4 u5_mult_82_U3296 ( .A1(u5_mult_82_SUMB_52__47_), .A2(
        u5_mult_82_CARRYB_52__46_), .ZN(u5_mult_82_n619) );
  AND2_X4 u5_mult_82_U3295 ( .A1(u5_mult_82_SUMB_52__48_), .A2(
        u5_mult_82_CARRYB_52__47_), .ZN(u5_mult_82_n618) );
  AND2_X4 u5_mult_82_U3294 ( .A1(u5_mult_82_SUMB_52__44_), .A2(
        u5_mult_82_CARRYB_52__43_), .ZN(u5_mult_82_n617) );
  XOR2_X2 u5_mult_82_U3293 ( .A(u5_mult_82_CARRYB_52__51_), .B(
        u5_mult_82_ab_52__52_), .Z(u5_mult_82_n616) );
  XOR2_X2 u5_mult_82_U3292 ( .A(u5_mult_82_CARRYB_52__50_), .B(
        u5_mult_82_SUMB_52__51_), .Z(u5_mult_82_n615) );
  XOR2_X2 u5_mult_82_U3291 ( .A(u5_mult_82_ab_1__18_), .B(u5_mult_82_ab_0__19_), .Z(u5_mult_82_n614) );
  INV_X4 u5_mult_82_U3290 ( .A(u5_mult_82_n932), .ZN(u5_mult_82_n1505) );
  XOR2_X2 u5_mult_82_U3289 ( .A(u5_mult_82_SUMB_46__24_), .B(u5_mult_82_n778), 
        .Z(u5_mult_82_SUMB_47__23_) );
  OR2_X4 u5_mult_82_U3288 ( .A1(u5_mult_82_n1264), .A2(u5_mult_82_net66089), 
        .ZN(u5_mult_82_n613) );
  AND2_X2 u5_mult_82_U3287 ( .A1(u5_mult_82_ab_0__39_), .A2(
        u5_mult_82_ab_1__38_), .ZN(u5_mult_82_n612) );
  AND2_X2 u5_mult_82_U3286 ( .A1(u5_mult_82_ab_0__11_), .A2(
        u5_mult_82_ab_1__10_), .ZN(u5_mult_82_n611) );
  AND2_X2 u5_mult_82_U3285 ( .A1(u5_mult_82_ab_0__34_), .A2(
        u5_mult_82_ab_1__33_), .ZN(u5_mult_82_n610) );
  XNOR2_X2 u5_mult_82_U3284 ( .A(u5_mult_82_SUMB_14__38_), .B(u5_mult_82_n961), 
        .ZN(u5_mult_82_n609) );
  AND2_X2 u5_mult_82_U3283 ( .A1(u5_mult_82_SUMB_52__16_), .A2(
        u5_mult_82_CARRYB_52__15_), .ZN(u5_mult_82_n608) );
  AND2_X4 u5_mult_82_U3282 ( .A1(u5_mult_82_SUMB_52__33_), .A2(
        u5_mult_82_CARRYB_52__32_), .ZN(u5_mult_82_n607) );
  AND2_X4 u5_mult_82_U3281 ( .A1(u5_mult_82_SUMB_52__36_), .A2(
        u5_mult_82_CARRYB_52__35_), .ZN(u5_mult_82_n606) );
  AND2_X4 u5_mult_82_U3280 ( .A1(u5_mult_82_SUMB_52__35_), .A2(
        u5_mult_82_CARRYB_52__34_), .ZN(u5_mult_82_n605) );
  AND2_X4 u5_mult_82_U3279 ( .A1(u5_mult_82_SUMB_52__37_), .A2(
        u5_mult_82_CARRYB_52__36_), .ZN(u5_mult_82_n604) );
  AND2_X4 u5_mult_82_U3278 ( .A1(u5_mult_82_SUMB_52__38_), .A2(
        u5_mult_82_CARRYB_52__37_), .ZN(u5_mult_82_n603) );
  AND2_X4 u5_mult_82_U3277 ( .A1(u5_mult_82_SUMB_52__40_), .A2(
        u5_mult_82_CARRYB_52__39_), .ZN(u5_mult_82_n602) );
  AND2_X4 u5_mult_82_U3276 ( .A1(u5_mult_82_SUMB_52__41_), .A2(
        u5_mult_82_CARRYB_52__40_), .ZN(u5_mult_82_n601) );
  AND2_X4 u5_mult_82_U3275 ( .A1(u5_mult_82_SUMB_52__42_), .A2(
        u5_mult_82_CARRYB_52__41_), .ZN(u5_mult_82_n600) );
  AND2_X2 u5_mult_82_U3274 ( .A1(u5_mult_82_ab_0__32_), .A2(
        u5_mult_82_ab_1__31_), .ZN(u5_mult_82_n599) );
  AND2_X4 u5_mult_82_U3273 ( .A1(u5_mult_82_SUMB_52__4_), .A2(
        u5_mult_82_CARRYB_52__3_), .ZN(u5_mult_82_n598) );
  AND2_X2 u5_mult_82_U3272 ( .A1(u5_mult_82_SUMB_52__39_), .A2(
        u5_mult_82_CARRYB_52__38_), .ZN(u5_mult_82_n596) );
  AND2_X2 u5_mult_82_U3271 ( .A1(u5_mult_82_SUMB_52__22_), .A2(
        u5_mult_82_CARRYB_52__21_), .ZN(u5_mult_82_n595) );
  INV_X4 u5_mult_82_U3270 ( .A(u5_mult_82_CARRYB_31__13_), .ZN(
        u5_mult_82_n4724) );
  AND2_X4 u5_mult_82_U3269 ( .A1(u5_mult_82_SUMB_52__8_), .A2(
        u5_mult_82_CARRYB_52__7_), .ZN(u5_mult_82_n594) );
  AND2_X4 u5_mult_82_U3268 ( .A1(u5_mult_82_SUMB_52__31_), .A2(
        u5_mult_82_CARRYB_52__30_), .ZN(u5_mult_82_n593) );
  AND2_X4 u5_mult_82_U3267 ( .A1(u5_mult_82_SUMB_52__10_), .A2(
        u5_mult_82_CARRYB_52__9_), .ZN(u5_mult_82_n592) );
  AND2_X4 u5_mult_82_U3266 ( .A1(u5_mult_82_SUMB_52__23_), .A2(
        u5_mult_82_CARRYB_52__22_), .ZN(u5_mult_82_n591) );
  AND2_X4 u5_mult_82_U3265 ( .A1(u5_mult_82_SUMB_52__34_), .A2(
        u5_mult_82_CARRYB_52__33_), .ZN(u5_mult_82_n590) );
  AND2_X4 u5_mult_82_U3264 ( .A1(u5_mult_82_SUMB_52__12_), .A2(
        u5_mult_82_CARRYB_52__11_), .ZN(u5_mult_82_n589) );
  AND2_X4 u5_mult_82_U3263 ( .A1(u5_mult_82_SUMB_52__9_), .A2(
        u5_mult_82_CARRYB_52__8_), .ZN(u5_mult_82_n588) );
  AND2_X4 u5_mult_82_U3262 ( .A1(u5_mult_82_SUMB_52__26_), .A2(
        u5_mult_82_CARRYB_52__25_), .ZN(u5_mult_82_n587) );
  AND2_X2 u5_mult_82_U3261 ( .A1(u5_mult_82_ab_0__36_), .A2(u5_mult_82_n2748), 
        .ZN(u5_mult_82_n586) );
  AND2_X2 u5_mult_82_U3260 ( .A1(u5_mult_82_SUMB_52__25_), .A2(
        u5_mult_82_CARRYB_52__24_), .ZN(u5_mult_82_n585) );
  AND2_X4 u5_mult_82_U3259 ( .A1(u5_mult_82_SUMB_52__24_), .A2(
        u5_mult_82_CARRYB_52__23_), .ZN(u5_mult_82_n582) );
  AND2_X4 u5_mult_82_U3258 ( .A1(u5_mult_82_SUMB_52__13_), .A2(
        u5_mult_82_CARRYB_52__12_), .ZN(u5_mult_82_n581) );
  INV_X4 u5_mult_82_U3257 ( .A(u5_mult_82_n7022), .ZN(u5_mult_82_n6973) );
  INV_X8 u5_mult_82_U3256 ( .A(u5_mult_82_n6744), .ZN(u5_mult_82_n6743) );
  INV_X16 u5_mult_82_U3255 ( .A(fracta_mul[46]), .ZN(u5_mult_82_n6740) );
  INV_X16 u5_mult_82_U3254 ( .A(u5_mult_82_n6677), .ZN(u5_mult_82_n6682) );
  INV_X4 u5_mult_82_U3253 ( .A(u5_mult_82_n7000), .ZN(u5_mult_82_n6676) );
  INV_X16 u5_mult_82_U3252 ( .A(u5_mult_82_n6724), .ZN(u5_mult_82_n6723) );
  INV_X8 u5_mult_82_U3251 ( .A(u5_mult_82_n6719), .ZN(u5_mult_82_n6725) );
  INV_X8 u5_mult_82_U3250 ( .A(fracta_mul[37]), .ZN(u5_mult_82_n6719) );
  INV_X16 u5_mult_82_U3249 ( .A(u5_mult_82_net65521), .ZN(u5_mult_82_net65519)
         );
  INV_X8 u5_mult_82_U3248 ( .A(u5_mult_82_net65525), .ZN(u5_mult_82_net65523)
         );
  INV_X8 u5_mult_82_U3247 ( .A(fracta_mul[34]), .ZN(u5_mult_82_net65525) );
  INV_X16 u5_mult_82_U3246 ( .A(u5_mult_82_n6670), .ZN(u5_mult_82_n6675) );
  INV_X4 u5_mult_82_U3245 ( .A(u5_mult_82_n6999), .ZN(u5_mult_82_n6669) );
  INV_X16 u5_mult_82_U3244 ( .A(u5_mult_82_n6607), .ZN(u5_mult_82_n6612) );
  INV_X4 u5_mult_82_U3243 ( .A(u5_mult_82_n6998), .ZN(u5_mult_82_n6606) );
  INV_X8 u5_mult_82_U3242 ( .A(u5_mult_82_n6634), .ZN(u5_mult_82_n6640) );
  INV_X8 u5_mult_82_U3241 ( .A(fracta_mul[22]), .ZN(u5_mult_82_n6634) );
  INV_X16 u5_mult_82_U3240 ( .A(u5_mult_82_n6626), .ZN(u5_mult_82_n6621) );
  INV_X4 u5_mult_82_U3239 ( .A(u5_mult_82_n6620), .ZN(u5_mult_82_n6626) );
  INV_X8 u5_mult_82_U3238 ( .A(fracta_mul[20]), .ZN(u5_mult_82_n6620) );
  INV_X16 u5_mult_82_U3237 ( .A(u5_mult_82_n6562), .ZN(u5_mult_82_n6557) );
  INV_X8 u5_mult_82_U3236 ( .A(u5_mult_82_n6556), .ZN(u5_mult_82_n6562) );
  INV_X8 u5_mult_82_U3235 ( .A(fracta_mul[11]), .ZN(u5_mult_82_n6556) );
  INV_X16 u5_mult_82_U3234 ( .A(u5_mult_82_n7020), .ZN(u5_mult_82_n6911) );
  INV_X16 u5_mult_82_U3233 ( .A(u5_mult_82_n7019), .ZN(u5_mult_82_n6890) );
  INV_X16 u5_mult_82_U3232 ( .A(n4787), .ZN(u5_mult_82_n6815) );
  INV_X16 u5_mult_82_U3231 ( .A(u5_mult_82_n6873), .ZN(u5_mult_82_n6872) );
  INV_X16 u5_mult_82_U3230 ( .A(n4742), .ZN(u5_mult_82_n6836) );
  INV_X16 u5_mult_82_U3229 ( .A(n4777), .ZN(u5_mult_82_n6825) );
  INV_X16 u5_mult_82_U3228 ( .A(n4775), .ZN(u5_mult_82_n6809) );
  INV_X16 u5_mult_82_U3227 ( .A(n4811), .ZN(u5_mult_82_n6771) );
  INV_X4 u5_mult_82_U3226 ( .A(u5_mult_82_n1832), .ZN(u5_mult_82_n1833) );
  AND2_X4 u5_mult_82_U3225 ( .A1(u5_mult_82_SUMB_52__43_), .A2(
        u5_mult_82_CARRYB_52__42_), .ZN(u5_mult_82_n580) );
  AND2_X4 u5_mult_82_U3224 ( .A1(u5_mult_82_SUMB_52__3_), .A2(
        u5_mult_82_CARRYB_52__2_), .ZN(u5_mult_82_n579) );
  AND2_X2 u5_mult_82_U3223 ( .A1(u5_mult_82_SUMB_52__15_), .A2(
        u5_mult_82_CARRYB_52__14_), .ZN(u5_mult_82_n578) );
  AND2_X4 u5_mult_82_U3222 ( .A1(u5_mult_82_SUMB_52__17_), .A2(
        u5_mult_82_CARRYB_52__16_), .ZN(u5_mult_82_n577) );
  AND2_X4 u5_mult_82_U3221 ( .A1(u5_mult_82_n725), .A2(
        u5_mult_82_CARRYB_52__6_), .ZN(u5_mult_82_n576) );
  AND2_X4 u5_mult_82_U3220 ( .A1(u5_mult_82_SUMB_52__5_), .A2(
        u5_mult_82_CARRYB_52__4_), .ZN(u5_mult_82_n575) );
  AND2_X4 u5_mult_82_U3219 ( .A1(u5_mult_82_SUMB_52__18_), .A2(
        u5_mult_82_CARRYB_52__17_), .ZN(u5_mult_82_n574) );
  INV_X4 u5_mult_82_U3218 ( .A(u5_mult_82_n6738), .ZN(u5_mult_82_n6737) );
  INV_X16 u5_mult_82_U3217 ( .A(u5_mult_82_n6733), .ZN(u5_mult_82_n6739) );
  INV_X16 u5_mult_82_U3216 ( .A(fracta_mul[44]), .ZN(u5_mult_82_n6733) );
  INV_X4 u5_mult_82_U3215 ( .A(u5_mult_82_n1320), .ZN(u5_mult_82_net65375) );
  INV_X8 u5_mult_82_U3214 ( .A(u5_mult_82_n1321), .ZN(u5_mult_82_net65379) );
  INV_X16 u5_mult_82_U3213 ( .A(fracta_mul[42]), .ZN(u5_mult_82_n1321) );
  INV_X16 u5_mult_82_U3212 ( .A(u5_mult_82_n1351), .ZN(u5_mult_82_net65447) );
  INV_X8 u5_mult_82_U3211 ( .A(u5_mult_82_n1352), .ZN(u5_mult_82_net65451) );
  INV_X8 u5_mult_82_U3210 ( .A(fracta_mul[38]), .ZN(u5_mult_82_n1352) );
  INV_X16 u5_mult_82_U3209 ( .A(u5_mult_82_n6703), .ZN(u5_mult_82_n6702) );
  INV_X16 u5_mult_82_U3208 ( .A(u5_mult_82_n6704), .ZN(u5_mult_82_n6699) );
  INV_X8 u5_mult_82_U3207 ( .A(u5_mult_82_n6698), .ZN(u5_mult_82_n6704) );
  INV_X8 u5_mult_82_U3206 ( .A(fracta_mul[33]), .ZN(u5_mult_82_n6698) );
  INV_X16 u5_mult_82_U3205 ( .A(u5_mult_82_n6688), .ZN(u5_mult_82_n6687) );
  INV_X8 u5_mult_82_U3204 ( .A(u5_mult_82_n6683), .ZN(u5_mult_82_n6689) );
  INV_X8 u5_mult_82_U3203 ( .A(fracta_mul[31]), .ZN(u5_mult_82_n6683) );
  INV_X8 u5_mult_82_U3202 ( .A(u5_mult_82_n6641), .ZN(u5_mult_82_n6647) );
  INV_X8 u5_mult_82_U3201 ( .A(fracta_mul[24]), .ZN(u5_mult_82_n6641) );
  INV_X16 u5_mult_82_U3200 ( .A(u5_mult_82_net65721), .ZN(u5_mult_82_net65711)
         );
  INV_X8 u5_mult_82_U3199 ( .A(u5_mult_82_n1344), .ZN(u5_mult_82_net65721) );
  INV_X8 u5_mult_82_U3198 ( .A(fracta_mul[23]), .ZN(u5_mult_82_n1344) );
  INV_X8 u5_mult_82_U3197 ( .A(u5_mult_82_n6667), .ZN(u5_mult_82_n6666) );
  INV_X16 u5_mult_82_U3196 ( .A(u5_mult_82_n6668), .ZN(u5_mult_82_n6663) );
  INV_X8 u5_mult_82_U3195 ( .A(u5_mult_82_n6662), .ZN(u5_mult_82_n6668) );
  INV_X16 u5_mult_82_U3194 ( .A(fracta_mul[28]), .ZN(u5_mult_82_n6662) );
  INV_X4 u5_mult_82_U3193 ( .A(u5_mult_82_n1380), .ZN(u5_mult_82_net65681) );
  INV_X8 u5_mult_82_U3192 ( .A(u5_mult_82_n1381), .ZN(u5_mult_82_net65685) );
  INV_X16 u5_mult_82_U3191 ( .A(fracta_mul[25]), .ZN(u5_mult_82_n1381) );
  INV_X4 u5_mult_82_U3190 ( .A(u5_mult_82_n6653), .ZN(u5_mult_82_n6652) );
  INV_X16 u5_mult_82_U3189 ( .A(u5_mult_82_n6648), .ZN(u5_mult_82_n6653) );
  INV_X16 u5_mult_82_U3188 ( .A(fracta_mul[26]), .ZN(u5_mult_82_n6648) );
  INV_X16 u5_mult_82_U3187 ( .A(u5_mult_82_n6633), .ZN(u5_mult_82_n6628) );
  INV_X8 u5_mult_82_U3186 ( .A(u5_mult_82_n6627), .ZN(u5_mult_82_n6633) );
  INV_X8 u5_mult_82_U3185 ( .A(fracta_mul[21]), .ZN(u5_mult_82_n6627) );
  INV_X8 u5_mult_82_U3184 ( .A(u5_mult_82_n6577), .ZN(u5_mult_82_n6583) );
  INV_X8 u5_mult_82_U3183 ( .A(fracta_mul[14]), .ZN(u5_mult_82_n6577) );
  INV_X8 u5_mult_82_U3182 ( .A(u6_N11), .ZN(u5_mult_82_n1319) );
  INV_X8 u5_mult_82_U3181 ( .A(u5_mult_82_n1319), .ZN(u5_mult_82_n1318) );
  INV_X8 u5_mult_82_U3180 ( .A(u5_mult_82_n6532), .ZN(u5_mult_82_n6531) );
  INV_X8 u5_mult_82_U3179 ( .A(u5_mult_82_n6527), .ZN(u5_mult_82_n6533) );
  INV_X8 u5_mult_82_U3178 ( .A(fracta_mul[7]), .ZN(u5_mult_82_n6527) );
  INV_X8 u5_mult_82_U3177 ( .A(u5_mult_82_n6539), .ZN(u5_mult_82_n6538) );
  INV_X16 u5_mult_82_U3176 ( .A(u5_mult_82_n6540), .ZN(u5_mult_82_n6535) );
  INV_X8 u5_mult_82_U3175 ( .A(u5_mult_82_n6534), .ZN(u5_mult_82_n6540) );
  INV_X16 u5_mult_82_U3174 ( .A(fracta_mul[8]), .ZN(u5_mult_82_n6534) );
  INV_X16 u5_mult_82_U3173 ( .A(u5_mult_82_net66025), .ZN(u5_mult_82_net66021)
         );
  INV_X8 u5_mult_82_U3172 ( .A(u5_mult_82_n1359), .ZN(u5_mult_82_n1358) );
  INV_X8 u5_mult_82_U3171 ( .A(fracta_mul[6]), .ZN(u5_mult_82_n1359) );
  INV_X16 u5_mult_82_U3170 ( .A(u6_N6), .ZN(u5_mult_82_n1271) );
  INV_X8 u5_mult_82_U3169 ( .A(u5_mult_82_n1271), .ZN(u5_mult_82_n1270) );
  INV_X8 u5_mult_82_U3168 ( .A(u6_N5), .ZN(u5_mult_82_net64373) );
  INV_X8 u5_mult_82_U3167 ( .A(u5_mult_82_net64373), .ZN(u5_mult_82_net64371)
         );
  INV_X8 u5_mult_82_U3166 ( .A(u5_mult_82_n6554), .ZN(u5_mult_82_n6553) );
  INV_X16 u5_mult_82_U3165 ( .A(u5_mult_82_n6555), .ZN(u5_mult_82_n6550) );
  INV_X4 u5_mult_82_U3164 ( .A(u5_mult_82_n6549), .ZN(u5_mult_82_n6555) );
  INV_X8 u5_mult_82_U3163 ( .A(fracta_mul[10]), .ZN(u5_mult_82_n6549) );
  INV_X4 u5_mult_82_U3162 ( .A(u5_mult_82_n6971), .ZN(u5_mult_82_n6970) );
  INV_X8 u5_mult_82_U3161 ( .A(u6_N1), .ZN(u5_mult_82_n6966) );
  INV_X8 u5_mult_82_U3160 ( .A(u5_mult_82_n6966), .ZN(u5_mult_82_n6972) );
  INV_X16 u5_mult_82_U3159 ( .A(u5_mult_82_n6575), .ZN(u5_mult_82_n6572) );
  INV_X16 u5_mult_82_U3158 ( .A(u5_mult_82_n6576), .ZN(u5_mult_82_n6571) );
  INV_X4 u5_mult_82_U3157 ( .A(u5_mult_82_n6570), .ZN(u5_mult_82_n6576) );
  INV_X8 u5_mult_82_U3156 ( .A(fracta_mul[13]), .ZN(u5_mult_82_n6570) );
  INV_X16 u5_mult_82_U3155 ( .A(u5_mult_82_n6992), .ZN(u5_mult_82_n6517) );
  INV_X4 u5_mult_82_U3154 ( .A(fracta_mul[3]), .ZN(u5_mult_82_n6992) );
  INV_X8 u5_mult_82_U3153 ( .A(u6_N15), .ZN(u5_mult_82_n6932) );
  INV_X8 u5_mult_82_U3152 ( .A(u5_mult_82_n6932), .ZN(u5_mult_82_n6938) );
  INV_X8 u5_mult_82_U3151 ( .A(u6_N16), .ZN(u5_mult_82_net64571) );
  INV_X8 u5_mult_82_U3150 ( .A(u5_mult_82_net64571), .ZN(u5_mult_82_net64569)
         );
  INV_X16 u5_mult_82_U3149 ( .A(u6_N13), .ZN(u5_mult_82_net64517) );
  INV_X8 u5_mult_82_U3148 ( .A(u5_mult_82_net64517), .ZN(u5_mult_82_net64515)
         );
  AND2_X4 u5_mult_82_U3147 ( .A1(u5_mult_82_SUMB_52__6_), .A2(
        u5_mult_82_CARRYB_52__5_), .ZN(u5_mult_82_n573) );
  INV_X8 u5_mult_82_U3146 ( .A(u5_mult_82_n6731), .ZN(u5_mult_82_n6730) );
  INV_X16 u5_mult_82_U3145 ( .A(u5_mult_82_n6732), .ZN(u5_mult_82_n6727) );
  INV_X8 u5_mult_82_U3144 ( .A(u5_mult_82_n6726), .ZN(u5_mult_82_n6732) );
  INV_X8 u5_mult_82_U3143 ( .A(fracta_mul[39]), .ZN(u5_mult_82_n6726) );
  INV_X16 u5_mult_82_U3142 ( .A(u5_mult_82_n1343), .ZN(u5_mult_82_net65717) );
  INV_X16 u5_mult_82_U3141 ( .A(u5_mult_82_n6619), .ZN(u5_mult_82_n6614) );
  INV_X4 u5_mult_82_U3140 ( .A(u5_mult_82_n6613), .ZN(u5_mult_82_n6619) );
  INV_X8 u5_mult_82_U3139 ( .A(fracta_mul[19]), .ZN(u5_mult_82_n6613) );
  INV_X8 u5_mult_82_U3138 ( .A(u5_mult_82_n6994), .ZN(u5_mult_82_n6542) );
  INV_X8 u5_mult_82_U3137 ( .A(u5_mult_82_n6542), .ZN(u5_mult_82_n6541) );
  INV_X8 u5_mult_82_U3136 ( .A(u6_N4), .ZN(u5_mult_82_n6945) );
  INV_X8 u5_mult_82_U3135 ( .A(u5_mult_82_n6945), .ZN(u5_mult_82_n6950) );
  INV_X16 u5_mult_82_U3134 ( .A(u6_N8), .ZN(u5_mult_82_net64427) );
  INV_X8 u5_mult_82_U3133 ( .A(u5_mult_82_net64427), .ZN(u5_mult_82_net64425)
         );
  INV_X16 u5_mult_82_U3132 ( .A(u5_mult_82_n1372), .ZN(u5_mult_82_net64451) );
  INV_X8 u5_mult_82_U3131 ( .A(u6_N10), .ZN(u5_mult_82_n1373) );
  INV_X4 u5_mult_82_U3130 ( .A(u5_mult_82_n1373), .ZN(u5_mult_82_n1372) );
  INV_X16 u5_mult_82_U3129 ( .A(u6_N7), .ZN(u5_mult_82_n6939) );
  INV_X8 u5_mult_82_U3128 ( .A(u5_mult_82_n6939), .ZN(u5_mult_82_n6944) );
  INV_X16 u5_mult_82_U3127 ( .A(u6_N9), .ZN(u5_mult_82_n1289) );
  INV_X8 u5_mult_82_U3126 ( .A(u5_mult_82_n1289), .ZN(u5_mult_82_n1288) );
  INV_X16 u5_mult_82_U3125 ( .A(u6_N14), .ZN(u5_mult_82_net64535) );
  INV_X8 u5_mult_82_U3124 ( .A(u5_mult_82_net64535), .ZN(u5_mult_82_net64533)
         );
  INV_X16 u5_mult_82_U3123 ( .A(u6_N12), .ZN(u5_mult_82_net64499) );
  INV_X8 u5_mult_82_U3122 ( .A(u5_mult_82_net64499), .ZN(u5_mult_82_net64497)
         );
  INV_X16 u5_mult_82_U3121 ( .A(n4809), .ZN(u5_mult_82_n6783) );
  INV_X16 u5_mult_82_U3120 ( .A(u5_mult_82_n6783), .ZN(u5_mult_82_n6788) );
  INV_X8 u5_mult_82_U3119 ( .A(u6_N17), .ZN(u5_mult_82_n6926) );
  INV_X8 u5_mult_82_U3118 ( .A(u5_mult_82_n6926), .ZN(u5_mult_82_n6931) );
  INV_X1 u5_mult_82_U3117 ( .A(u2_N157), .ZN(u5_mult_82_n7022) );
  INV_X4 u5_mult_82_U3116 ( .A(u5_mult_82_net65197), .ZN(u5_mult_82_net65191)
         );
  INV_X4 u5_mult_82_U3115 ( .A(u5_mult_82_net65197), .ZN(u5_mult_82_net65189)
         );
  NOR2_X1 u5_mult_82_U3114 ( .A1(u5_mult_82_net64223), .A2(u5_mult_82_n6986), 
        .ZN(u5_N0) );
  NOR2_X2 u5_mult_82_U3113 ( .A1(u5_mult_82_n6989), .A2(u5_mult_82_net66093), 
        .ZN(u5_mult_82_ab_2__0_) );
  NOR2_X1 u5_mult_82_U3112 ( .A1(u5_mult_82_n6989), .A2(u5_mult_82_n6531), 
        .ZN(u5_mult_82_ab_7__0_) );
  NOR2_X2 u5_mult_82_U3111 ( .A1(u5_mult_82_n6989), .A2(u5_mult_82_n6568), 
        .ZN(u5_mult_82_ab_12__0_) );
  NOR2_X2 u5_mult_82_U3110 ( .A1(u5_mult_82_n6988), .A2(u5_mult_82_n6604), 
        .ZN(u5_mult_82_ab_17__0_) );
  NOR2_X2 u5_mult_82_U3109 ( .A1(u5_mult_82_n6988), .A2(u5_mult_82_n6638), 
        .ZN(u5_mult_82_ab_22__0_) );
  NOR2_X2 u5_mult_82_U3108 ( .A1(u5_mult_82_n6988), .A2(u5_mult_82_n6659), 
        .ZN(u5_mult_82_ab_27__0_) );
  NOR2_X2 u5_mult_82_U3107 ( .A1(u5_mult_82_n6987), .A2(u5_mult_82_n6696), 
        .ZN(u5_mult_82_ab_32__0_) );
  NOR2_X2 u5_mult_82_U3106 ( .A1(u5_mult_82_n6987), .A2(u5_mult_82_n6723), 
        .ZN(u5_mult_82_ab_37__0_) );
  NOR2_X1 u5_mult_82_U3105 ( .A1(u5_mult_82_n6986), .A2(u5_mult_82_net65375), 
        .ZN(u5_mult_82_ab_42__0_) );
  NOR2_X1 u5_mult_82_U3104 ( .A1(u5_mult_82_n6986), .A2(u5_mult_82_n6755), 
        .ZN(u5_mult_82_ab_49__0_) );
  NOR2_X1 u5_mult_82_U3103 ( .A1(u5_mult_82_n6970), .A2(u5_mult_82_net66093), 
        .ZN(u5_mult_82_ab_2__1_) );
  NOR2_X1 u5_mult_82_U3102 ( .A1(u5_mult_82_n6969), .A2(u5_mult_82_n6531), 
        .ZN(u5_mult_82_ab_7__1_) );
  NOR2_X2 u5_mult_82_U3101 ( .A1(u5_mult_82_n6969), .A2(u5_mult_82_n6568), 
        .ZN(u5_mult_82_ab_12__1_) );
  NOR2_X2 u5_mult_82_U3100 ( .A1(u5_mult_82_n6968), .A2(u5_mult_82_n6604), 
        .ZN(u5_mult_82_ab_17__1_) );
  NOR2_X2 u5_mult_82_U3099 ( .A1(u5_mult_82_n6968), .A2(u5_mult_82_n6638), 
        .ZN(u5_mult_82_ab_22__1_) );
  NOR2_X2 u5_mult_82_U3098 ( .A1(u5_mult_82_n6968), .A2(u5_mult_82_n6659), 
        .ZN(u5_mult_82_ab_27__1_) );
  NOR2_X2 u5_mult_82_U3097 ( .A1(u5_mult_82_n6967), .A2(u5_mult_82_n6696), 
        .ZN(u5_mult_82_ab_32__1_) );
  NOR2_X1 u5_mult_82_U3096 ( .A1(u5_mult_82_n6967), .A2(u5_mult_82_n6737), 
        .ZN(u5_mult_82_ab_44__1_) );
  NOR2_X1 u5_mult_82_U3095 ( .A1(u5_mult_82_n6967), .A2(u5_mult_82_n6755), 
        .ZN(u5_mult_82_ab_49__1_) );
  NOR2_X1 u5_mult_82_U3094 ( .A1(u5_mult_82_n6967), .A2(u5_mult_82_net65191), 
        .ZN(u5_mult_82_ab_51__1_) );
  INV_X4 u5_mult_82_U3093 ( .A(u5_mult_82_n6973), .ZN(u5_mult_82_n6974) );
  NOR2_X1 u5_mult_82_U3092 ( .A1(u5_mult_82_n6983), .A2(u5_mult_82_n6974), 
        .ZN(u5_mult_82_ab_52__52_) );
  NOR2_X1 u5_mult_82_U3091 ( .A1(u5_mult_82_n6975), .A2(u5_mult_82_n6759), 
        .ZN(u5_mult_82_ab_52__51_) );
  NOR2_X1 u5_mult_82_U3090 ( .A1(u5_mult_82_n6983), .A2(u5_mult_82_net65189), 
        .ZN(u5_mult_82_ab_51__52_) );
  NOR2_X2 u5_mult_82_U3089 ( .A1(u5_mult_82_n6963), .A2(u5_mult_82_net66093), 
        .ZN(u5_mult_82_ab_2__2_) );
  NOR2_X1 u5_mult_82_U3088 ( .A1(u5_mult_82_n6962), .A2(u5_mult_82_n6531), 
        .ZN(u5_mult_82_ab_7__2_) );
  INV_X8 u5_mult_82_U3087 ( .A(u5_mult_82_n6549), .ZN(u5_mult_82_n6554) );
  INV_X8 u5_mult_82_U3086 ( .A(u5_mult_82_n6570), .ZN(u5_mult_82_n6575) );
  NOR2_X2 u5_mult_82_U3085 ( .A1(u5_mult_82_n6962), .A2(u5_mult_82_n6568), 
        .ZN(u5_mult_82_ab_12__2_) );
  INV_X8 u5_mult_82_U3084 ( .A(u5_mult_82_n6577), .ZN(u5_mult_82_n6582) );
  NOR2_X2 u5_mult_82_U3083 ( .A1(u5_mult_82_n6961), .A2(u5_mult_82_n6604), 
        .ZN(u5_mult_82_ab_17__2_) );
  INV_X8 u5_mult_82_U3082 ( .A(u5_mult_82_n6613), .ZN(u5_mult_82_n6618) );
  INV_X8 u5_mult_82_U3081 ( .A(u5_mult_82_n6620), .ZN(u5_mult_82_n6625) );
  INV_X8 u5_mult_82_U3080 ( .A(u5_mult_82_n1344), .ZN(u5_mult_82_n1343) );
  NOR2_X2 u5_mult_82_U3079 ( .A1(u5_mult_82_n6961), .A2(u5_mult_82_n6638), 
        .ZN(u5_mult_82_ab_22__2_) );
  INV_X8 u5_mult_82_U3078 ( .A(u5_mult_82_n6641), .ZN(u5_mult_82_n6646) );
  INV_X8 u5_mult_82_U3077 ( .A(u5_mult_82_n1381), .ZN(u5_mult_82_n1380) );
  INV_X8 u5_mult_82_U3076 ( .A(u5_mult_82_n6662), .ZN(u5_mult_82_n6667) );
  NOR2_X2 u5_mult_82_U3075 ( .A1(u5_mult_82_n6961), .A2(u5_mult_82_n6659), 
        .ZN(u5_mult_82_ab_27__2_) );
  INV_X8 u5_mult_82_U3074 ( .A(u5_mult_82_n6698), .ZN(u5_mult_82_n6703) );
  INV_X8 u5_mult_82_U3073 ( .A(u5_mult_82_net65525), .ZN(u5_mult_82_net65521)
         );
  INV_X8 u5_mult_82_U3072 ( .A(u5_mult_82_n1352), .ZN(u5_mult_82_n1351) );
  NOR2_X2 u5_mult_82_U3071 ( .A1(u5_mult_82_n6960), .A2(u5_mult_82_n6723), 
        .ZN(u5_mult_82_ab_37__2_) );
  NOR2_X1 u5_mult_82_U3070 ( .A1(u5_mult_82_n6960), .A2(u5_mult_82_n6755), 
        .ZN(u5_mult_82_ab_49__2_) );
  NOR2_X1 u5_mult_82_U3069 ( .A1(u5_mult_82_n6960), .A2(u5_mult_82_net65229), 
        .ZN(u5_mult_82_ab_50__2_) );
  NOR2_X1 u5_mult_82_U3068 ( .A1(u5_mult_82_n6952), .A2(u5_mult_82_n6755), 
        .ZN(u5_mult_82_ab_49__3_) );
  INV_X4 u5_mult_82_U3067 ( .A(u5_mult_82_n6423), .ZN(u5_mult_82_CLA_SUM[88])
         );
  NOR2_X2 u5_mult_82_U3066 ( .A1(u5_mult_82_n6960), .A2(u5_mult_82_n6737), 
        .ZN(u5_mult_82_ab_44__2_) );
  NOR2_X2 u5_mult_82_U3065 ( .A1(u5_mult_82_n6952), .A2(u5_mult_82_net65355), 
        .ZN(u5_mult_82_ab_43__3_) );
  INV_X8 u5_mult_82_U3064 ( .A(u5_mult_82_n6740), .ZN(u5_mult_82_n6744) );
  INV_X4 u5_mult_82_U3063 ( .A(u5_mult_82_n6993), .ZN(u5_mult_82_n6519) );
  NOR2_X2 u5_mult_82_U3062 ( .A1(u5_mult_82_n6956), .A2(u5_mult_82_net66093), 
        .ZN(u5_mult_82_ab_2__3_) );
  INV_X4 u5_mult_82_U3061 ( .A(u5_mult_82_n1301), .ZN(u5_mult_82_n1304) );
  NOR2_X1 u5_mult_82_U3060 ( .A1(u5_mult_82_n6955), .A2(u5_mult_82_n6531), 
        .ZN(u5_mult_82_ab_7__3_) );
  NOR2_X2 u5_mult_82_U3059 ( .A1(u5_mult_82_n6955), .A2(u5_mult_82_n6568), 
        .ZN(u5_mult_82_ab_12__3_) );
  INV_X8 u5_mult_82_U3058 ( .A(fracta_mul[15]), .ZN(u5_mult_82_n6584) );
  NOR2_X2 u5_mult_82_U3057 ( .A1(u5_mult_82_n6954), .A2(u5_mult_82_n6604), 
        .ZN(u5_mult_82_ab_17__3_) );
  NOR2_X2 u5_mult_82_U3056 ( .A1(u5_mult_82_n6954), .A2(u5_mult_82_n6638), 
        .ZN(u5_mult_82_ab_22__3_) );
  NOR2_X2 u5_mult_82_U3055 ( .A1(u5_mult_82_n6954), .A2(u5_mult_82_n6659), 
        .ZN(u5_mult_82_ab_27__3_) );
  NOR2_X1 u5_mult_82_U3054 ( .A1(u5_mult_82_n6946), .A2(u5_mult_82_n6680), 
        .ZN(u5_mult_82_ab_30__4_) );
  INV_X8 u5_mult_82_U3053 ( .A(u5_mult_82_n6726), .ZN(u5_mult_82_n6731) );
  INV_X4 u5_mult_82_U3052 ( .A(u5_mult_82_n7005), .ZN(u5_mult_82_n6751) );
  NOR2_X1 u5_mult_82_U3051 ( .A1(u5_mult_82_n6974), .A2(u5_mult_82_n6940), 
        .ZN(u5_mult_82_ab_52__7_) );
  NOR2_X1 u5_mult_82_U3050 ( .A1(u5_mult_82_n6974), .A2(u5_mult_82_net64433), 
        .ZN(u5_mult_82_ab_52__9_) );
  NOR2_X1 u5_mult_82_U3049 ( .A1(u5_mult_82_n6974), .A2(u5_mult_82_net64455), 
        .ZN(u5_mult_82_ab_52__10_) );
  NOR2_X1 u5_mult_82_U3048 ( .A1(u5_mult_82_n6975), .A2(u5_mult_82_net64559), 
        .ZN(u5_mult_82_ab_52__16_) );
  NOR2_X1 u5_mult_82_U3047 ( .A1(u5_mult_82_n6975), .A2(u5_mult_82_n6927), 
        .ZN(u5_mult_82_ab_52__17_) );
  NOR2_X1 u5_mult_82_U3046 ( .A1(u5_mult_82_n6975), .A2(u5_mult_82_n6919), 
        .ZN(u5_mult_82_ab_52__18_) );
  INV_X4 u5_mult_82_U3045 ( .A(u5_mult_82_ab_52__20_), .ZN(u5_mult_82_n2019)
         );
  NAND3_X2 u5_mult_82_U3044 ( .A1(u5_mult_82_n4312), .A2(u5_mult_82_n4313), 
        .A3(u5_mult_82_n4314), .ZN(u5_mult_82_CARRYB_52__21_) );
  NOR2_X1 u5_mult_82_U3043 ( .A1(u5_mult_82_n6976), .A2(u5_mult_82_n6856), 
        .ZN(u5_mult_82_ab_52__30_) );
  NAND2_X2 u5_mult_82_U3042 ( .A1(u5_mult_82_n1053), .A2(u5_mult_82_n1054), 
        .ZN(u5_mult_82_SUMB_51__34_) );
  NOR2_X1 u5_mult_82_U3041 ( .A1(u5_mult_82_n6976), .A2(u5_mult_82_n6837), 
        .ZN(u5_mult_82_ab_52__33_) );
  NOR2_X1 u5_mult_82_U3040 ( .A1(u5_mult_82_n6976), .A2(u5_mult_82_net64881), 
        .ZN(u5_mult_82_ab_52__34_) );
  NOR2_X1 u5_mult_82_U3039 ( .A1(u5_mult_82_n6977), .A2(u5_mult_82_n6777), 
        .ZN(u5_mult_82_ab_52__48_) );
  NOR2_X1 u5_mult_82_U3038 ( .A1(u5_mult_82_n6977), .A2(u5_mult_82_n6772), 
        .ZN(u5_mult_82_ab_52__49_) );
  NOR2_X1 u5_mult_82_U3037 ( .A1(u5_mult_82_n6976), .A2(u5_mult_82_net64935), 
        .ZN(u5_mult_82_ab_52__37_) );
  NOR2_X1 u5_mult_82_U3036 ( .A1(u5_mult_82_n6977), .A2(u5_mult_82_net64957), 
        .ZN(u5_mult_82_ab_52__38_) );
  NOR2_X1 u5_mult_82_U3035 ( .A1(u5_mult_82_n6977), .A2(u5_mult_82_n6831), 
        .ZN(u5_mult_82_ab_52__39_) );
  NOR2_X2 u5_mult_82_U3034 ( .A1(u5_mult_82_n6947), .A2(u5_mult_82_net66093), 
        .ZN(u5_mult_82_ab_2__4_) );
  NOR2_X2 u5_mult_82_U3033 ( .A1(u5_mult_82_n6948), .A2(u5_mult_82_n6530), 
        .ZN(u5_mult_82_ab_7__4_) );
  NOR2_X2 u5_mult_82_U3032 ( .A1(u5_mult_82_n6948), .A2(u5_mult_82_n6567), 
        .ZN(u5_mult_82_ab_12__4_) );
  NOR2_X2 u5_mult_82_U3031 ( .A1(u5_mult_82_n6947), .A2(u5_mult_82_n6603), 
        .ZN(u5_mult_82_ab_17__4_) );
  NOR2_X2 u5_mult_82_U3030 ( .A1(u5_mult_82_net64363), .A2(u5_mult_82_n6610), 
        .ZN(u5_mult_82_ab_18__5_) );
  NOR2_X1 u5_mult_82_U3029 ( .A1(u5_mult_82_n6947), .A2(u5_mult_82_net65717), 
        .ZN(u5_mult_82_ab_23__4_) );
  INV_X4 u5_mult_82_U3028 ( .A(u5_mult_82_net65521), .ZN(u5_mult_82_net65517)
         );
  NOR2_X2 u5_mult_82_U3027 ( .A1(u5_mult_82_net64379), .A2(u5_mult_82_n6695), 
        .ZN(u5_mult_82_ab_32__6_) );
  NOR2_X2 u5_mult_82_U3026 ( .A1(u5_mult_82_net64361), .A2(u5_mult_82_n6716), 
        .ZN(u5_mult_82_ab_36__5_) );
  INV_X4 u5_mult_82_U3025 ( .A(u5_mult_82_n1351), .ZN(u5_mult_82_net65445) );
  NOR2_X2 u5_mult_82_U3024 ( .A1(u5_mult_82_net64379), .A2(u5_mult_82_n6716), 
        .ZN(u5_mult_82_ab_36__6_) );
  NOR2_X1 u5_mult_82_U3023 ( .A1(u5_mult_82_net64361), .A2(u5_mult_82_n6748), 
        .ZN(u5_mult_82_ab_48__5_) );
  NOR2_X1 u5_mult_82_U3022 ( .A1(u5_mult_82_n6946), .A2(u5_mult_82_net65229), 
        .ZN(u5_mult_82_ab_50__4_) );
  NAND3_X2 u5_mult_82_U3021 ( .A1(u5_mult_82_n4169), .A2(u5_mult_82_n4170), 
        .A3(u5_mult_82_n4171), .ZN(u5_mult_82_CARRYB_51__8_) );
  NOR2_X1 u5_mult_82_U3020 ( .A1(u5_mult_82_n6975), .A2(u5_mult_82_net64487), 
        .ZN(u5_mult_82_ab_52__12_) );
  NOR2_X1 u5_mult_82_U3019 ( .A1(u5_mult_82_net64505), .A2(u5_mult_82_net65189), .ZN(u5_mult_82_ab_51__13_) );
  NOR2_X1 u5_mult_82_U3018 ( .A1(u5_mult_82_n6933), .A2(u5_mult_82_net65189), 
        .ZN(u5_mult_82_ab_51__15_) );
  NOR2_X1 u5_mult_82_U3017 ( .A1(u5_mult_82_n6975), .A2(u5_mult_82_n6912), 
        .ZN(u5_mult_82_ab_52__19_) );
  NOR2_X1 u5_mult_82_U3016 ( .A1(u5_mult_82_n6874), .A2(u5_mult_82_net65191), 
        .ZN(u5_mult_82_ab_51__27_) );
  NOR2_X1 u5_mult_82_U3015 ( .A1(u5_mult_82_n6879), .A2(u5_mult_82_net65191), 
        .ZN(u5_mult_82_ab_51__26_) );
  NOR2_X1 u5_mult_82_U3014 ( .A1(u5_mult_82_n6976), .A2(u5_mult_82_n6874), 
        .ZN(u5_mult_82_ab_52__27_) );
  NOR2_X1 u5_mult_82_U3013 ( .A1(u5_mult_82_n6861), .A2(u5_mult_82_net65191), 
        .ZN(u5_mult_82_ab_51__29_) );
  NOR2_X1 u5_mult_82_U3012 ( .A1(u5_mult_82_n6867), .A2(u5_mult_82_net65191), 
        .ZN(u5_mult_82_ab_51__28_) );
  NOR2_X1 u5_mult_82_U3011 ( .A1(u5_mult_82_n6976), .A2(u5_mult_82_n6849), 
        .ZN(u5_mult_82_ab_52__31_) );
  NOR2_X1 u5_mult_82_U3010 ( .A1(u5_mult_82_n6976), .A2(u5_mult_82_n6842), 
        .ZN(u5_mult_82_ab_52__32_) );
  NOR2_X1 u5_mult_82_U3009 ( .A1(u5_mult_82_n6784), .A2(u5_mult_82_net65191), 
        .ZN(u5_mult_82_ab_51__47_) );
  NOR2_X1 u5_mult_82_U3008 ( .A1(u5_mult_82_n6797), .A2(u5_mult_82_net65193), 
        .ZN(u5_mult_82_ab_51__45_) );
  NOR2_X1 u5_mult_82_U3007 ( .A1(u5_mult_82_n6803), .A2(u5_mult_82_net65193), 
        .ZN(u5_mult_82_ab_51__44_) );
  INV_X4 u5_mult_82_U3006 ( .A(u5_mult_82_ab_51__25_), .ZN(u5_mult_82_n3704)
         );
  NOR2_X2 u5_mult_82_U3005 ( .A1(u5_mult_82_n6891), .A2(u5_mult_82_net65191), 
        .ZN(u5_mult_82_ab_51__24_) );
  NOR2_X2 u5_mult_82_U3004 ( .A1(u5_mult_82_n6884), .A2(u5_mult_82_net65229), 
        .ZN(u5_mult_82_ab_50__25_) );
  NOR2_X2 u5_mult_82_U3003 ( .A1(u5_mult_82_net64367), .A2(u5_mult_82_net66093), .ZN(u5_mult_82_ab_2__5_) );
  NOR2_X2 u5_mult_82_U3002 ( .A1(u5_mult_82_net64365), .A2(u5_mult_82_n6530), 
        .ZN(u5_mult_82_ab_7__5_) );
  NOR2_X2 u5_mult_82_U3001 ( .A1(u5_mult_82_net64365), .A2(u5_mult_82_n6567), 
        .ZN(u5_mult_82_ab_12__5_) );
  INV_X4 u5_mult_82_U3000 ( .A(u5_mult_82_n6575), .ZN(u5_mult_82_n6573) );
  INV_X4 u5_mult_82_U2999 ( .A(u5_mult_82_n6582), .ZN(u5_mult_82_n6580) );
  INV_X4 u5_mult_82_U2998 ( .A(u5_mult_82_n6618), .ZN(u5_mult_82_n6616) );
  NOR2_X2 u5_mult_82_U2997 ( .A1(u5_mult_82_net64381), .A2(u5_mult_82_n6637), 
        .ZN(u5_mult_82_ab_22__6_) );
  INV_X4 u5_mult_82_U2996 ( .A(u5_mult_82_n1343), .ZN(u5_mult_82_net65713) );
  INV_X4 u5_mult_82_U2995 ( .A(u5_mult_82_n6646), .ZN(u5_mult_82_n6644) );
  NOR2_X1 u5_mult_82_U2994 ( .A1(u5_mult_82_net64361), .A2(u5_mult_82_n6680), 
        .ZN(u5_mult_82_ab_30__5_) );
  INV_X4 u5_mult_82_U2993 ( .A(u5_mult_82_n6703), .ZN(u5_mult_82_n6701) );
  INV_X4 u5_mult_82_U2992 ( .A(u5_mult_82_n6731), .ZN(u5_mult_82_n6729) );
  INV_X2 u5_mult_82_U2991 ( .A(u5_mult_82_CARRYB_43__4_), .ZN(u5_mult_82_n2978) );
  INV_X4 u5_mult_82_U2990 ( .A(u5_mult_82_ab_43__5_), .ZN(u5_mult_82_n4802) );
  INV_X4 u5_mult_82_U2989 ( .A(u5_mult_82_n6744), .ZN(u5_mult_82_n6742) );
  INV_X4 u5_mult_82_U2988 ( .A(u5_mult_82_ab_44__6_), .ZN(u5_mult_82_n4615) );
  NOR2_X1 u5_mult_82_U2987 ( .A1(u5_mult_82_net64361), .A2(u5_mult_82_n6755), 
        .ZN(u5_mult_82_ab_49__5_) );
  NOR2_X1 u5_mult_82_U2986 ( .A1(u5_mult_82_net64379), .A2(u5_mult_82_net65189), .ZN(u5_mult_82_ab_51__6_) );
  NOR2_X1 u5_mult_82_U2985 ( .A1(u5_mult_82_net64415), .A2(u5_mult_82_net65229), .ZN(u5_mult_82_ab_50__8_) );
  NOR2_X2 u5_mult_82_U2984 ( .A1(u5_mult_82_net64433), .A2(u5_mult_82_net65229), .ZN(u5_mult_82_ab_50__9_) );
  NOR2_X1 u5_mult_82_U2983 ( .A1(u5_mult_82_net64487), .A2(u5_mult_82_net65229), .ZN(u5_mult_82_ab_50__12_) );
  NOR2_X1 u5_mult_82_U2982 ( .A1(u5_mult_82_net64469), .A2(u5_mult_82_net65229), .ZN(u5_mult_82_ab_50__11_) );
  NOR2_X1 u5_mult_82_U2981 ( .A1(u5_mult_82_net64505), .A2(u5_mult_82_net65229), .ZN(u5_mult_82_ab_50__13_) );
  NOR2_X1 u5_mult_82_U2980 ( .A1(u5_mult_82_net64559), .A2(u5_mult_82_net65229), .ZN(u5_mult_82_ab_50__16_) );
  NOR2_X1 u5_mult_82_U2979 ( .A1(u5_mult_82_n6912), .A2(u5_mult_82_net65229), 
        .ZN(u5_mult_82_ab_50__19_) );
  NOR2_X1 u5_mult_82_U2978 ( .A1(u5_mult_82_n6903), .A2(u5_mult_82_net65229), 
        .ZN(u5_mult_82_ab_50__20_) );
  NOR2_X1 u5_mult_82_U2977 ( .A1(u5_mult_82_n6903), .A2(u5_mult_82_net65189), 
        .ZN(u5_mult_82_ab_51__20_) );
  NOR2_X1 u5_mult_82_U2976 ( .A1(u5_mult_82_n6895), .A2(u5_mult_82_net65189), 
        .ZN(u5_mult_82_ab_51__21_) );
  NOR2_X1 u5_mult_82_U2975 ( .A1(u5_mult_82_net64665), .A2(u5_mult_82_net65189), .ZN(u5_mult_82_ab_51__22_) );
  NOR2_X1 u5_mult_82_U2974 ( .A1(u5_mult_82_n6879), .A2(u5_mult_82_net65229), 
        .ZN(u5_mult_82_ab_50__26_) );
  INV_X16 u5_mult_82_U2973 ( .A(u5_mult_82_n1272), .ZN(u5_mult_82_net65225) );
  NOR2_X1 u5_mult_82_U2972 ( .A1(u5_mult_82_n6842), .A2(u5_mult_82_net65191), 
        .ZN(u5_mult_82_ab_51__32_) );
  INV_X4 u5_mult_82_U2971 ( .A(u5_mult_82_n1748), .ZN(u5_mult_82_n1749) );
  NOR2_X1 u5_mult_82_U2970 ( .A1(u5_mult_82_net64935), .A2(u5_mult_82_net65225), .ZN(u5_mult_82_ab_50__37_) );
  INV_X8 u5_mult_82_U2969 ( .A(u5_mult_82_n1269), .ZN(u5_mult_82_n1265) );
  INV_X16 u5_mult_82_U2968 ( .A(u5_mult_82_n6790), .ZN(u5_mult_82_n6789) );
  NOR2_X1 u5_mult_82_U2967 ( .A1(u5_mult_82_n6816), .A2(u5_mult_82_net65223), 
        .ZN(u5_mult_82_ab_50__42_) );
  NOR2_X1 u5_mult_82_U2966 ( .A1(u5_mult_82_n6891), .A2(u5_mult_82_net65229), 
        .ZN(u5_mult_82_ab_50__24_) );
  NOR2_X2 u5_mult_82_U2965 ( .A1(u5_mult_82_n6879), .A2(u5_mult_82_n6749), 
        .ZN(u5_mult_82_ab_48__26_) );
  NOR2_X2 u5_mult_82_U2964 ( .A1(u5_mult_82_net64385), .A2(u5_mult_82_net66093), .ZN(u5_mult_82_ab_2__6_) );
  NOR2_X2 u5_mult_82_U2963 ( .A1(u5_mult_82_net64383), .A2(u5_mult_82_n6530), 
        .ZN(u5_mult_82_ab_7__6_) );
  NOR2_X2 u5_mult_82_U2962 ( .A1(u5_mult_82_net64383), .A2(u5_mult_82_n6567), 
        .ZN(u5_mult_82_ab_12__6_) );
  NOR2_X2 u5_mult_82_U2961 ( .A1(u5_mult_82_n6941), .A2(u5_mult_82_n6637), 
        .ZN(u5_mult_82_ab_22__7_) );
  NOR2_X2 u5_mult_82_U2960 ( .A1(u5_mult_82_n6940), .A2(u5_mult_82_n6716), 
        .ZN(u5_mult_82_ab_36__7_) );
  NAND2_X2 u5_mult_82_U2959 ( .A1(u5_mult_82_net86159), .A2(u5_mult_82_n1298), 
        .ZN(u5_mult_82_n1300) );
  NOR2_X1 u5_mult_82_U2958 ( .A1(u5_mult_82_n6940), .A2(u5_mult_82_net65229), 
        .ZN(u5_mult_82_ab_50__7_) );
  NOR2_X2 u5_mult_82_U2957 ( .A1(u5_mult_82_net64415), .A2(u5_mult_82_n6755), 
        .ZN(u5_mult_82_ab_49__8_) );
  NAND3_X2 u5_mult_82_U2956 ( .A1(u5_mult_82_net81825), .A2(u5_mult_82_n4341), 
        .A3(u5_mult_82_net81827), .ZN(u5_mult_82_CARRYB_48__8_) );
  INV_X4 u5_mult_82_U2955 ( .A(u5_mult_82_ab_48__10_), .ZN(u5_mult_82_n5222)
         );
  NOR2_X2 u5_mult_82_U2954 ( .A1(u5_mult_82_net64487), .A2(u5_mult_82_n6755), 
        .ZN(u5_mult_82_ab_49__12_) );
  NAND3_X2 u5_mult_82_U2953 ( .A1(u5_mult_82_n6108), .A2(u5_mult_82_n6109), 
        .A3(u5_mult_82_n6110), .ZN(u5_mult_82_CARRYB_48__12_) );
  NOR2_X1 u5_mult_82_U2952 ( .A1(u5_mult_82_net64559), .A2(u5_mult_82_n6749), 
        .ZN(u5_mult_82_ab_48__16_) );
  NOR2_X1 u5_mult_82_U2951 ( .A1(u5_mult_82_net64523), .A2(u5_mult_82_net65229), .ZN(u5_mult_82_ab_50__14_) );
  NOR2_X1 u5_mult_82_U2950 ( .A1(u5_mult_82_net64523), .A2(u5_mult_82_n6755), 
        .ZN(u5_mult_82_ab_49__14_) );
  NAND3_X2 u5_mult_82_U2949 ( .A1(u5_mult_82_n3217), .A2(u5_mult_82_n3218), 
        .A3(u5_mult_82_n3219), .ZN(u5_mult_82_CARRYB_48__17_) );
  NOR2_X1 u5_mult_82_U2948 ( .A1(u5_mult_82_n6927), .A2(u5_mult_82_net65229), 
        .ZN(u5_mult_82_ab_50__17_) );
  NOR2_X2 u5_mult_82_U2947 ( .A1(u5_mult_82_n6895), .A2(u5_mult_82_n6754), 
        .ZN(u5_mult_82_ab_49__21_) );
  NOR2_X1 u5_mult_82_U2946 ( .A1(u5_mult_82_net64665), .A2(u5_mult_82_net65229), .ZN(u5_mult_82_ab_50__22_) );
  NOR2_X2 u5_mult_82_U2945 ( .A1(u5_mult_82_n6884), .A2(u5_mult_82_net65285), 
        .ZN(u5_mult_82_ab_47__25_) );
  NOR2_X1 u5_mult_82_U2944 ( .A1(u5_mult_82_net64683), .A2(u5_mult_82_n6754), 
        .ZN(u5_mult_82_ab_49__23_) );
  NOR2_X1 u5_mult_82_U2943 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_net65279), .ZN(u5_mult_82_ab_47__38_) );
  NOR2_X1 u5_mult_82_U2942 ( .A1(u5_mult_82_n6983), .A2(u5_mult_82_n6743), 
        .ZN(u5_mult_82_ab_46__52_) );
  NOR2_X2 u5_mult_82_U2941 ( .A1(u5_mult_82_n6759), .A2(u5_mult_82_net65277), 
        .ZN(u5_mult_82_ab_47__51_) );
  NOR2_X2 u5_mult_82_U2940 ( .A1(u5_mult_82_n6856), .A2(u5_mult_82_net65279), 
        .ZN(u5_mult_82_ab_47__30_) );
  NOR2_X2 u5_mult_82_U2939 ( .A1(u5_mult_82_n6941), .A2(u5_mult_82_net66093), 
        .ZN(u5_mult_82_ab_2__7_) );
  NOR2_X2 u5_mult_82_U2938 ( .A1(u5_mult_82_n6942), .A2(u5_mult_82_n6530), 
        .ZN(u5_mult_82_ab_7__7_) );
  NOR2_X2 u5_mult_82_U2937 ( .A1(u5_mult_82_n6942), .A2(u5_mult_82_n6567), 
        .ZN(u5_mult_82_ab_12__7_) );
  NOR2_X2 u5_mult_82_U2936 ( .A1(u5_mult_82_net64417), .A2(u5_mult_82_n6596), 
        .ZN(u5_mult_82_ab_16__8_) );
  INV_X4 u5_mult_82_U2935 ( .A(u5_mult_82_ab_25__9_), .ZN(u5_mult_82_n2198) );
  NOR2_X1 u5_mult_82_U2934 ( .A1(u5_mult_82_net64451), .A2(u5_mult_82_n6665), 
        .ZN(u5_mult_82_ab_28__10_) );
  NOR2_X1 u5_mult_82_U2933 ( .A1(u5_mult_82_net64433), .A2(u5_mult_82_n6665), 
        .ZN(u5_mult_82_ab_28__9_) );
  NOR2_X1 u5_mult_82_U2932 ( .A1(u5_mult_82_net64433), .A2(u5_mult_82_n6695), 
        .ZN(u5_mult_82_ab_32__9_) );
  NOR2_X1 u5_mult_82_U2931 ( .A1(u5_mult_82_net64415), .A2(u5_mult_82_n6722), 
        .ZN(u5_mult_82_ab_37__8_) );
  INV_X4 u5_mult_82_U2930 ( .A(u5_mult_82_ab_45__8_), .ZN(u5_mult_82_n3500) );
  INV_X4 u5_mult_82_U2929 ( .A(u5_mult_82_ab_47__12_), .ZN(u5_mult_82_n5541)
         );
  NAND3_X2 u5_mult_82_U2928 ( .A1(u5_mult_82_n5679), .A2(u5_mult_82_n5680), 
        .A3(u5_mult_82_n5681), .ZN(u5_mult_82_CARRYB_46__11_) );
  NAND3_X2 u5_mult_82_U2927 ( .A1(u5_mult_82_n5776), .A2(u5_mult_82_n5777), 
        .A3(u5_mult_82_n5778), .ZN(u5_mult_82_CARRYB_46__14_) );
  NOR2_X2 u5_mult_82_U2926 ( .A1(u5_mult_82_net64665), .A2(u5_mult_82_net65285), .ZN(u5_mult_82_ab_47__22_) );
  NOR2_X2 u5_mult_82_U2925 ( .A1(u5_mult_82_n6903), .A2(u5_mult_82_n6741), 
        .ZN(u5_mult_82_ab_46__20_) );
  NOR2_X1 u5_mult_82_U2924 ( .A1(u5_mult_82_n6891), .A2(u5_mult_82_net65285), 
        .ZN(u5_mult_82_ab_47__24_) );
  NOR2_X2 u5_mult_82_U2923 ( .A1(u5_mult_82_n6837), .A2(u5_mult_82_net65279), 
        .ZN(u5_mult_82_ab_47__33_) );
  NOR2_X2 u5_mult_82_U2922 ( .A1(u5_mult_82_net64913), .A2(u5_mult_82_net65279), .ZN(u5_mult_82_ab_47__35_) );
  NOR2_X2 u5_mult_82_U2921 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6747), 
        .ZN(u5_mult_82_ab_48__36_) );
  NAND3_X2 u5_mult_82_U2920 ( .A1(u5_mult_82_n2219), .A2(u5_mult_82_n2220), 
        .A3(u5_mult_82_n2221), .ZN(u5_mult_82_CARRYB_46__39_) );
  NOR2_X2 u5_mult_82_U2919 ( .A1(u5_mult_82_n6826), .A2(u5_mult_82_n6741), 
        .ZN(u5_mult_82_ab_46__40_) );
  NOR2_X2 u5_mult_82_U2918 ( .A1(u5_mult_82_net64417), .A2(u5_mult_82_net66093), .ZN(u5_mult_82_ab_2__8_) );
  NOR2_X2 u5_mult_82_U2917 ( .A1(u5_mult_82_net64419), .A2(u5_mult_82_n6530), 
        .ZN(u5_mult_82_ab_7__8_) );
  NAND3_X2 u5_mult_82_U2916 ( .A1(u5_mult_82_n2778), .A2(u5_mult_82_n2779), 
        .A3(u5_mult_82_n2780), .ZN(u5_mult_82_CARRYB_23__8_) );
  NOR2_X1 u5_mult_82_U2915 ( .A1(u5_mult_82_net64451), .A2(u5_mult_82_n6695), 
        .ZN(u5_mult_82_ab_32__10_) );
  NOR2_X2 u5_mult_82_U2914 ( .A1(u5_mult_82_n6933), .A2(u5_mult_82_n6742), 
        .ZN(u5_mult_82_ab_46__15_) );
  INV_X4 u5_mult_82_U2913 ( .A(u5_mult_82_ab_47__16_), .ZN(u5_mult_82_n3115)
         );
  NOR2_X2 u5_mult_82_U2912 ( .A1(u5_mult_82_n6895), .A2(u5_mult_82_n6741), 
        .ZN(u5_mult_82_ab_46__21_) );
  NOR2_X2 u5_mult_82_U2911 ( .A1(u5_mult_82_n6861), .A2(u5_mult_82_n6734), 
        .ZN(u5_mult_82_ab_44__29_) );
  NOR2_X2 u5_mult_82_U2910 ( .A1(u5_mult_82_n6867), .A2(u5_mult_82_n6734), 
        .ZN(u5_mult_82_ab_44__28_) );
  NOR2_X2 u5_mult_82_U2909 ( .A1(u5_mult_82_net64935), .A2(u5_mult_82_n6741), 
        .ZN(u5_mult_82_ab_46__37_) );
  NOR2_X2 u5_mult_82_U2908 ( .A1(u5_mult_82_n6849), .A2(u5_mult_82_net65351), 
        .ZN(u5_mult_82_ab_43__31_) );
  NOR2_X1 u5_mult_82_U2907 ( .A1(u5_mult_82_net64451), .A2(u5_mult_82_n6716), 
        .ZN(u5_mult_82_ab_36__10_) );
  NOR2_X2 u5_mult_82_U2906 ( .A1(u5_mult_82_net64435), .A2(u5_mult_82_net66093), .ZN(u5_mult_82_ab_2__9_) );
  NOR2_X2 u5_mult_82_U2905 ( .A1(u5_mult_82_net64437), .A2(u5_mult_82_n6530), 
        .ZN(u5_mult_82_ab_7__9_) );
  NOR2_X2 u5_mult_82_U2904 ( .A1(u5_mult_82_net64453), .A2(u5_mult_82_n6596), 
        .ZN(u5_mult_82_ab_16__10_) );
  NOR2_X2 u5_mult_82_U2903 ( .A1(u5_mult_82_net64471), .A2(u5_mult_82_n6596), 
        .ZN(u5_mult_82_ab_16__11_) );
  NAND3_X2 u5_mult_82_U2902 ( .A1(u5_mult_82_n3728), .A2(u5_mult_82_n3729), 
        .A3(u5_mult_82_n3730), .ZN(u5_mult_82_CARRYB_22__9_) );
  NOR2_X2 u5_mult_82_U2901 ( .A1(u5_mult_82_net64489), .A2(u5_mult_82_n6658), 
        .ZN(u5_mult_82_ab_27__12_) );
  NAND3_X2 u5_mult_82_U2900 ( .A1(u5_mult_82_n1980), .A2(u5_mult_82_n1981), 
        .A3(u5_mult_82_n1982), .ZN(u5_mult_82_CARRYB_41__10_) );
  NOR2_X1 u5_mult_82_U2899 ( .A1(u5_mult_82_net64505), .A2(u5_mult_82_n6736), 
        .ZN(u5_mult_82_ab_44__13_) );
  NOR2_X1 u5_mult_82_U2898 ( .A1(u5_mult_82_n6816), .A2(u5_mult_82_net65313), 
        .ZN(u5_mult_82_ab_45__42_) );
  NOR2_X1 u5_mult_82_U2897 ( .A1(u5_mult_82_n6772), .A2(u5_mult_82_n6740), 
        .ZN(u5_mult_82_ab_46__49_) );
  NOR2_X1 u5_mult_82_U2896 ( .A1(u5_mult_82_n6777), .A2(u5_mult_82_n6740), 
        .ZN(u5_mult_82_ab_46__48_) );
  NOR2_X1 u5_mult_82_U2895 ( .A1(u5_mult_82_n6784), .A2(u5_mult_82_n6743), 
        .ZN(u5_mult_82_ab_46__47_) );
  NOR2_X2 u5_mult_82_U2894 ( .A1(u5_mult_82_net64881), .A2(u5_mult_82_net65351), .ZN(u5_mult_82_ab_43__34_) );
  NOR2_X2 u5_mult_82_U2893 ( .A1(u5_mult_82_n6842), .A2(u5_mult_82_net65351), 
        .ZN(u5_mult_82_ab_43__32_) );
  NOR2_X2 u5_mult_82_U2892 ( .A1(u5_mult_82_net64453), .A2(u5_mult_82_net66093), .ZN(u5_mult_82_ab_2__10_) );
  NOR2_X1 u5_mult_82_U2891 ( .A1(u5_mult_82_net64455), .A2(u5_mult_82_n6530), 
        .ZN(u5_mult_82_ab_7__10_) );
  NOR2_X1 u5_mult_82_U2890 ( .A1(u5_mult_82_net64507), .A2(u5_mult_82_net65717), .ZN(u5_mult_82_ab_23__13_) );
  NOR2_X1 u5_mult_82_U2889 ( .A1(u5_mult_82_net64469), .A2(u5_mult_82_net65355), .ZN(u5_mult_82_ab_43__11_) );
  INV_X4 u5_mult_82_U2888 ( .A(u5_mult_82_ab_43__19_), .ZN(u5_mult_82_n2292)
         );
  INV_X4 u5_mult_82_U2887 ( .A(u5_mult_82_ab_42__21_), .ZN(u5_mult_82_n1585)
         );
  NOR2_X2 u5_mult_82_U2886 ( .A1(u5_mult_82_net64665), .A2(u5_mult_82_net65371), .ZN(u5_mult_82_ab_42__22_) );
  INV_X4 u5_mult_82_U2885 ( .A(u5_mult_82_ab_42__27_), .ZN(u5_mult_82_n3701)
         );
  NOR2_X2 u5_mult_82_U2884 ( .A1(u5_mult_82_n6826), .A2(u5_mult_82_net65371), 
        .ZN(u5_mult_82_ab_42__40_) );
  NOR2_X1 u5_mult_82_U2883 ( .A1(u5_mult_82_n6831), .A2(u5_mult_82_net65369), 
        .ZN(u5_mult_82_ab_42__39_) );
  NAND3_X2 u5_mult_82_U2882 ( .A1(u5_mult_82_n2235), .A2(u5_mult_82_n2236), 
        .A3(u5_mult_82_n2237), .ZN(u5_mult_82_CARRYB_44__43_) );
  NOR2_X1 u5_mult_82_U2881 ( .A1(u5_mult_82_n6797), .A2(u5_mult_82_net65313), 
        .ZN(u5_mult_82_ab_45__45_) );
  NAND3_X2 u5_mult_82_U2880 ( .A1(u5_mult_82_n2265), .A2(u5_mult_82_n2266), 
        .A3(u5_mult_82_n2267), .ZN(u5_mult_82_CARRYB_44__44_) );
  NOR2_X2 u5_mult_82_U2879 ( .A1(u5_mult_82_net64475), .A2(u5_mult_82_net66093), .ZN(u5_mult_82_ab_2__11_) );
  NOR2_X2 u5_mult_82_U2878 ( .A1(u5_mult_82_net64473), .A2(u5_mult_82_n6530), 
        .ZN(u5_mult_82_ab_7__11_) );
  NOR2_X1 u5_mult_82_U2877 ( .A1(u5_mult_82_net64491), .A2(u5_mult_82_n6559), 
        .ZN(u5_mult_82_ab_11__12_) );
  NOR2_X1 u5_mult_82_U2876 ( .A1(u5_mult_82_net64509), .A2(u5_mult_82_n6559), 
        .ZN(u5_mult_82_ab_11__13_) );
  NOR2_X2 u5_mult_82_U2875 ( .A1(u5_mult_82_net64489), .A2(u5_mult_82_n6603), 
        .ZN(u5_mult_82_ab_17__12_) );
  NOR2_X2 u5_mult_82_U2874 ( .A1(u5_mult_82_net64507), .A2(u5_mult_82_n6603), 
        .ZN(u5_mult_82_ab_17__13_) );
  NOR2_X1 u5_mult_82_U2873 ( .A1(u5_mult_82_net64489), .A2(u5_mult_82_n6630), 
        .ZN(u5_mult_82_ab_21__12_) );
  NOR2_X2 u5_mult_82_U2872 ( .A1(u5_mult_82_n6934), .A2(u5_mult_82_n6637), 
        .ZN(u5_mult_82_ab_22__15_) );
  NOR2_X2 u5_mult_82_U2871 ( .A1(u5_mult_82_net64507), .A2(u5_mult_82_n6658), 
        .ZN(u5_mult_82_ab_27__13_) );
  NAND3_X2 u5_mult_82_U2870 ( .A1(u5_mult_82_n2602), .A2(u5_mult_82_n2603), 
        .A3(u5_mult_82_n2604), .ZN(u5_mult_82_CARRYB_31__12_) );
  NOR2_X1 u5_mult_82_U2869 ( .A1(u5_mult_82_net64469), .A2(u5_mult_82_n6722), 
        .ZN(u5_mult_82_ab_37__11_) );
  NOR2_X1 u5_mult_82_U2868 ( .A1(u5_mult_82_net64559), .A2(u5_mult_82_net65371), .ZN(u5_mult_82_ab_42__16_) );
  INV_X4 u5_mult_82_U2867 ( .A(u5_mult_82_ab_41__18_), .ZN(u5_mult_82_n4518)
         );
  NOR2_X1 u5_mult_82_U2866 ( .A1(u5_mult_82_n6891), .A2(u5_mult_82_net65389), 
        .ZN(u5_mult_82_ab_41__24_) );
  NOR2_X2 u5_mult_82_U2865 ( .A1(u5_mult_82_n6881), .A2(u5_mult_82_net65407), 
        .ZN(u5_mult_82_ab_40__26_) );
  NOR2_X2 u5_mult_82_U2864 ( .A1(u5_mult_82_n6869), .A2(u5_mult_82_net65405), 
        .ZN(u5_mult_82_ab_40__28_) );
  NOR2_X2 u5_mult_82_U2863 ( .A1(u5_mult_82_n6812), .A2(u5_mult_82_net65403), 
        .ZN(u5_mult_82_ab_40__43_) );
  NOR2_X2 u5_mult_82_U2862 ( .A1(u5_mult_82_n6805), .A2(u5_mult_82_net65403), 
        .ZN(u5_mult_82_ab_40__44_) );
  NOR2_X1 u5_mult_82_U2861 ( .A1(u5_mult_82_n6843), .A2(u5_mult_82_n6727), 
        .ZN(u5_mult_82_ab_39__32_) );
  NOR2_X2 u5_mult_82_U2860 ( .A1(u5_mult_82_net64883), .A2(u5_mult_82_net65441), .ZN(u5_mult_82_ab_38__34_) );
  INV_X4 u5_mult_82_U2859 ( .A(u5_mult_82_ab_22__13_), .ZN(u5_mult_82_n2501)
         );
  NOR2_X2 u5_mult_82_U2858 ( .A1(u5_mult_82_net64525), .A2(u5_mult_82_n6658), 
        .ZN(u5_mult_82_ab_27__14_) );
  NOR2_X1 u5_mult_82_U2857 ( .A1(u5_mult_82_net64523), .A2(u5_mult_82_n6680), 
        .ZN(u5_mult_82_ab_30__14_) );
  NOR2_X1 u5_mult_82_U2856 ( .A1(u5_mult_82_net64487), .A2(u5_mult_82_n6722), 
        .ZN(u5_mult_82_ab_37__12_) );
  NOR2_X2 u5_mult_82_U2855 ( .A1(u5_mult_82_net64523), .A2(u5_mult_82_net65445), .ZN(u5_mult_82_ab_38__14_) );
  NOR2_X2 u5_mult_82_U2854 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_net65405), .ZN(u5_mult_82_ab_40__38_) );
  NOR2_X1 u5_mult_82_U2853 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6727), 
        .ZN(u5_mult_82_ab_39__38_) );
  NOR2_X1 u5_mult_82_U2852 ( .A1(u5_mult_82_n6983), .A2(u5_mult_82_net65411), 
        .ZN(u5_mult_82_ab_40__52_) );
  NOR2_X2 u5_mult_82_U2851 ( .A1(u5_mult_82_n6760), .A2(u5_mult_82_net65385), 
        .ZN(u5_mult_82_ab_41__51_) );
  NOR2_X1 u5_mult_82_U2850 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_net65441), .ZN(u5_mult_82_ab_38__36_) );
  NOR2_X1 u5_mult_82_U2849 ( .A1(u5_mult_82_net64527), .A2(u5_mult_82_n6559), 
        .ZN(u5_mult_82_ab_11__14_) );
  NOR2_X2 u5_mult_82_U2848 ( .A1(u5_mult_82_n6935), .A2(u5_mult_82_n6567), 
        .ZN(u5_mult_82_ab_12__15_) );
  NOR2_X2 u5_mult_82_U2847 ( .A1(u5_mult_82_net64563), .A2(u5_mult_82_n6566), 
        .ZN(u5_mult_82_ab_12__16_) );
  NOR2_X2 u5_mult_82_U2846 ( .A1(u5_mult_82_n6928), .A2(u5_mult_82_n6629), 
        .ZN(u5_mult_82_ab_21__17_) );
  NAND2_X1 u5_mult_82_U2845 ( .A1(u5_mult_82_ab_36__13_), .A2(
        u5_mult_82_SUMB_35__14_), .ZN(u5_mult_82_n1997) );
  NAND3_X2 u5_mult_82_U2844 ( .A1(u5_mult_82_n1996), .A2(u5_mult_82_n1997), 
        .A3(u5_mult_82_n1998), .ZN(u5_mult_82_CARRYB_36__13_) );
  INV_X16 u5_mult_82_U2843 ( .A(u5_mult_82_n6854), .ZN(u5_mult_82_n6851) );
  NOR2_X2 u5_mult_82_U2842 ( .A1(u5_mult_82_n6791), .A2(u5_mult_82_n6729), 
        .ZN(u5_mult_82_ab_39__46_) );
  NOR2_X1 u5_mult_82_U2841 ( .A1(u5_mult_82_n6784), .A2(u5_mult_82_n6728), 
        .ZN(u5_mult_82_ab_39__47_) );
  NAND3_X2 u5_mult_82_U2840 ( .A1(u5_mult_82_n3656), .A2(u5_mult_82_n3657), 
        .A3(u5_mult_82_n3658), .ZN(u5_mult_82_CARRYB_30__15_) );
  NOR2_X2 u5_mult_82_U2839 ( .A1(u5_mult_82_net64223), .A2(u5_mult_82_net64535), .ZN(u5_mult_82_ab_0__14_) );
  INV_X8 u5_mult_82_U2838 ( .A(u5_mult_82_net64513), .ZN(u5_mult_82_net64511)
         );
  NOR2_X1 u5_mult_82_U2837 ( .A1(u5_mult_82_n6935), .A2(u5_mult_82_net66021), 
        .ZN(u5_mult_82_ab_6__15_) );
  INV_X4 u5_mult_82_U2836 ( .A(u5_mult_82_ab_17__15_), .ZN(u5_mult_82_n2066)
         );
  INV_X4 u5_mult_82_U2835 ( .A(u5_mult_82_ab_18__16_), .ZN(u5_mult_82_n2592)
         );
  INV_X4 u5_mult_82_U2834 ( .A(u5_mult_82_ab_17__17_), .ZN(u5_mult_82_n649) );
  NOR2_X2 u5_mult_82_U2833 ( .A1(u5_mult_82_net64667), .A2(u5_mult_82_n6721), 
        .ZN(u5_mult_82_ab_37__22_) );
  NOR2_X1 u5_mult_82_U2832 ( .A1(u5_mult_82_n6891), .A2(u5_mult_82_n6721), 
        .ZN(u5_mult_82_ab_37__24_) );
  NOR2_X2 u5_mult_82_U2831 ( .A1(u5_mult_82_n6885), .A2(u5_mult_82_n6721), 
        .ZN(u5_mult_82_ab_37__25_) );
  NOR2_X2 u5_mult_82_U2830 ( .A1(u5_mult_82_n6857), .A2(u5_mult_82_n6720), 
        .ZN(u5_mult_82_ab_37__30_) );
  INV_X16 u5_mult_82_U2829 ( .A(u5_mult_82_n7014), .ZN(u5_mult_82_n6865) );
  NOR2_X2 u5_mult_82_U2828 ( .A1(u5_mult_82_n6821), .A2(u5_mult_82_n6721), 
        .ZN(u5_mult_82_ab_37__41_) );
  NOR2_X1 u5_mult_82_U2827 ( .A1(u5_mult_82_n6816), .A2(u5_mult_82_n6721), 
        .ZN(u5_mult_82_ab_37__42_) );
  NOR2_X1 u5_mult_82_U2826 ( .A1(u5_mult_82_n6778), .A2(u5_mult_82_n6730), 
        .ZN(u5_mult_82_ab_39__48_) );
  NOR2_X2 u5_mult_82_U2825 ( .A1(u5_mult_82_n6767), .A2(u5_mult_82_net65385), 
        .ZN(u5_mult_82_ab_41__50_) );
  NOR2_X2 u5_mult_82_U2824 ( .A1(u5_mult_82_n6773), .A2(u5_mult_82_net65385), 
        .ZN(u5_mult_82_ab_41__49_) );
  NOR2_X1 u5_mult_82_U2823 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_net65513), .ZN(u5_mult_82_ab_34__36_) );
  NOR2_X2 u5_mult_82_U2822 ( .A1(u5_mult_82_net64223), .A2(u5_mult_82_n6932), 
        .ZN(u5_mult_82_ab_0__15_) );
  INV_X4 u5_mult_82_U2821 ( .A(u5_mult_82_n6582), .ZN(u5_mult_82_n6579) );
  NOR2_X1 u5_mult_82_U2820 ( .A1(u5_mult_82_n6929), .A2(u5_mult_82_n6572), 
        .ZN(u5_mult_82_ab_13__17_) );
  INV_X4 u5_mult_82_U2819 ( .A(u5_mult_82_ab_17__18_), .ZN(u5_mult_82_n2591)
         );
  INV_X4 u5_mult_82_U2818 ( .A(u5_mult_82_n6646), .ZN(u5_mult_82_n6643) );
  NOR2_X1 u5_mult_82_U2817 ( .A1(u5_mult_82_net64559), .A2(u5_mult_82_n6694), 
        .ZN(u5_mult_82_ab_32__16_) );
  NOR2_X2 u5_mult_82_U2816 ( .A1(u5_mult_82_n6913), .A2(u5_mult_82_n6721), 
        .ZN(u5_mult_82_ab_37__19_) );
  INV_X4 u5_mult_82_U2815 ( .A(u5_mult_82_ab_36__24_), .ZN(u5_mult_82_n3744)
         );
  NOR2_X2 u5_mult_82_U2814 ( .A1(u5_mult_82_net64883), .A2(u5_mult_82_net65513), .ZN(u5_mult_82_ab_34__34_) );
  NOR2_X2 u5_mult_82_U2813 ( .A1(u5_mult_82_net64901), .A2(u5_mult_82_net65513), .ZN(u5_mult_82_ab_34__35_) );
  NOR2_X1 u5_mult_82_U2812 ( .A1(u5_mult_82_n6791), .A2(u5_mult_82_n6706), 
        .ZN(u5_mult_82_ab_35__46_) );
  NOR2_X2 u5_mult_82_U2811 ( .A1(u5_mult_82_n6804), .A2(u5_mult_82_n6713), 
        .ZN(u5_mult_82_ab_36__44_) );
  INV_X16 u5_mult_82_U2810 ( .A(u5_mult_82_n6783), .ZN(u5_mult_82_n6787) );
  NAND3_X2 u5_mult_82_U2809 ( .A1(u5_mult_82_n3777), .A2(u5_mult_82_n3778), 
        .A3(u5_mult_82_n3779), .ZN(u5_mult_82_CARRYB_33__40_) );
  NOR2_X2 u5_mult_82_U2808 ( .A1(u5_mult_82_n6920), .A2(u5_mult_82_n6664), 
        .ZN(u5_mult_82_ab_28__18_) );
  NOR2_X2 u5_mult_82_U2807 ( .A1(u5_mult_82_net64223), .A2(u5_mult_82_net64571), .ZN(u5_mult_82_ab_0__16_) );
  INV_X8 u5_mult_82_U2806 ( .A(u5_mult_82_n6937), .ZN(u5_mult_82_n6936) );
  NOR2_X2 u5_mult_82_U2805 ( .A1(u5_mult_82_n6897), .A2(u5_mult_82_n6595), 
        .ZN(u5_mult_82_ab_16__21_) );
  INV_X4 u5_mult_82_U2804 ( .A(u5_mult_82_n1380), .ZN(u5_mult_82_net65677) );
  NOR2_X2 u5_mult_82_U2803 ( .A1(u5_mult_82_n6920), .A2(u5_mult_82_n6694), 
        .ZN(u5_mult_82_ab_32__18_) );
  NOR2_X2 u5_mult_82_U2802 ( .A1(u5_mult_82_n6913), .A2(u5_mult_82_n6694), 
        .ZN(u5_mult_82_ab_32__19_) );
  INV_X4 u5_mult_82_U2801 ( .A(u5_mult_82_n737), .ZN(u5_mult_82_n738) );
  NOR2_X2 u5_mult_82_U2800 ( .A1(u5_mult_82_n6880), .A2(u5_mult_82_net65515), 
        .ZN(u5_mult_82_ab_34__26_) );
  INV_X4 u5_mult_82_U2799 ( .A(u5_mult_82_ab_33__30_), .ZN(u5_mult_82_n5522)
         );
  NOR2_X2 u5_mult_82_U2798 ( .A1(u5_mult_82_n6838), .A2(u5_mult_82_net65513), 
        .ZN(u5_mult_82_ab_34__33_) );
  NOR2_X1 u5_mult_82_U2797 ( .A1(u5_mult_82_n6804), .A2(u5_mult_82_n6701), 
        .ZN(u5_mult_82_ab_33__44_) );
  NOR2_X2 u5_mult_82_U2796 ( .A1(u5_mult_82_n6797), .A2(u5_mult_82_n6706), 
        .ZN(u5_mult_82_ab_35__45_) );
  NOR2_X2 u5_mult_82_U2795 ( .A1(u5_mult_82_n6773), .A2(u5_mult_82_net65513), 
        .ZN(u5_mult_82_ab_34__49_) );
  NOR2_X2 u5_mult_82_U2794 ( .A1(u5_mult_82_n6778), .A2(u5_mult_82_net65519), 
        .ZN(u5_mult_82_ab_34__48_) );
  NOR2_X2 u5_mult_82_U2793 ( .A1(u5_mult_82_n6804), .A2(u5_mult_82_net65515), 
        .ZN(u5_mult_82_ab_34__44_) );
  NOR2_X2 u5_mult_82_U2792 ( .A1(u5_mult_82_n6832), .A2(u5_mult_82_n6699), 
        .ZN(u5_mult_82_ab_33__39_) );
  NAND3_X2 u5_mult_82_U2791 ( .A1(u5_mult_82_n5078), .A2(u5_mult_82_n5079), 
        .A3(u5_mult_82_n5080), .ZN(u5_mult_82_CARRYB_32__39_) );
  NOR2_X1 u5_mult_82_U2790 ( .A1(u5_mult_82_n6816), .A2(u5_mult_82_n6692), 
        .ZN(u5_mult_82_ab_32__42_) );
  NOR2_X2 u5_mult_82_U2789 ( .A1(u5_mult_82_net64219), .A2(u5_mult_82_n6926), 
        .ZN(u5_mult_82_ab_0__17_) );
  INV_X8 u5_mult_82_U2788 ( .A(u5_mult_82_net64567), .ZN(u5_mult_82_net64565)
         );
  NOR2_X2 u5_mult_82_U2787 ( .A1(u5_mult_82_n6915), .A2(u5_mult_82_n6515), 
        .ZN(u5_mult_82_ab_3__19_) );
  NOR2_X2 u5_mult_82_U2786 ( .A1(u5_mult_82_n6898), .A2(u5_mult_82_n6529), 
        .ZN(u5_mult_82_ab_7__21_) );
  NOR2_X2 u5_mult_82_U2785 ( .A1(u5_mult_82_net64669), .A2(u5_mult_82_n6595), 
        .ZN(u5_mult_82_ab_16__22_) );
  NOR2_X2 u5_mult_82_U2784 ( .A1(u5_mult_82_n6906), .A2(u5_mult_82_n6587), 
        .ZN(u5_mult_82_ab_15__20_) );
  NOR2_X2 u5_mult_82_U2783 ( .A1(u5_mult_82_n6905), .A2(u5_mult_82_n6636), 
        .ZN(u5_mult_82_ab_22__20_) );
  NOR2_X1 u5_mult_82_U2782 ( .A1(u5_mult_82_n6914), .A2(u5_mult_82_n6636), 
        .ZN(u5_mult_82_ab_22__19_) );
  NOR2_X2 u5_mult_82_U2781 ( .A1(u5_mult_82_n6896), .A2(u5_mult_82_n6685), 
        .ZN(u5_mult_82_ab_31__21_) );
  INV_X2 u5_mult_82_U2780 ( .A(u5_mult_82_n3605), .ZN(u5_mult_82_n3583) );
  NOR2_X2 u5_mult_82_U2779 ( .A1(u5_mult_82_n6767), .A2(u5_mult_82_net65525), 
        .ZN(u5_mult_82_ab_34__50_) );
  INV_X4 u5_mult_82_U2778 ( .A(u5_mult_82_ab_30__39_), .ZN(u5_mult_82_n2261)
         );
  NOR2_X2 u5_mult_82_U2777 ( .A1(u5_mult_82_n6906), .A2(u5_mult_82_n6515), 
        .ZN(u5_mult_82_ab_3__20_) );
  NOR2_X2 u5_mult_82_U2776 ( .A1(u5_mult_82_n6898), .A2(u5_mult_82_n6515), 
        .ZN(u5_mult_82_ab_3__21_) );
  NOR2_X2 u5_mult_82_U2775 ( .A1(u5_mult_82_net64685), .A2(u5_mult_82_n6694), 
        .ZN(u5_mult_82_ab_32__23_) );
  NOR2_X2 u5_mult_82_U2774 ( .A1(u5_mult_82_n6843), .A2(u5_mult_82_n6684), 
        .ZN(u5_mult_82_ab_31__32_) );
  NOR2_X1 u5_mult_82_U2773 ( .A1(u5_mult_82_n6982), .A2(u5_mult_82_n6702), 
        .ZN(u5_mult_82_ab_33__52_) );
  NOR2_X2 u5_mult_82_U2772 ( .A1(u5_mult_82_n6760), .A2(u5_mult_82_net65525), 
        .ZN(u5_mult_82_ab_34__51_) );
  BUF_X4 u5_mult_82_U2771 ( .A(u5_mult_82_SUMB_27__42_), .Z(u5_mult_82_n1836)
         );
  NAND3_X2 u5_mult_82_U2770 ( .A1(u5_mult_82_n4642), .A2(u5_mult_82_n4643), 
        .A3(u5_mult_82_n4644), .ZN(u5_mult_82_CARRYB_29__37_) );
  NAND3_X2 u5_mult_82_U2769 ( .A1(u5_mult_82_n5667), .A2(u5_mult_82_n5668), 
        .A3(u5_mult_82_n5669), .ZN(u5_mult_82_CARRYB_29__36_) );
  INV_X8 u5_mult_82_U2768 ( .A(u5_mult_82_n6924), .ZN(u5_mult_82_n6923) );
  NOR2_X2 u5_mult_82_U2767 ( .A1(u5_mult_82_n6906), .A2(u5_mult_82_n6566), 
        .ZN(u5_mult_82_ab_12__20_) );
  NOR2_X2 u5_mult_82_U2766 ( .A1(u5_mult_82_net64687), .A2(u5_mult_82_n6595), 
        .ZN(u5_mult_82_ab_16__23_) );
  NOR2_X2 u5_mult_82_U2765 ( .A1(u5_mult_82_n6897), .A2(u5_mult_82_n6636), 
        .ZN(u5_mult_82_ab_22__21_) );
  INV_X4 u5_mult_82_U2764 ( .A(u5_mult_82_ab_22__22_), .ZN(u5_mult_82_n858) );
  NOR2_X2 u5_mult_82_U2763 ( .A1(u5_mult_82_n6904), .A2(u5_mult_82_n6664), 
        .ZN(u5_mult_82_ab_28__20_) );
  NOR2_X2 u5_mult_82_U2762 ( .A1(u5_mult_82_n6896), .A2(u5_mult_82_n6664), 
        .ZN(u5_mult_82_ab_28__21_) );
  NAND3_X2 u5_mult_82_U2761 ( .A1(u5_mult_82_n2352), .A2(u5_mult_82_n2353), 
        .A3(u5_mult_82_n2354), .ZN(u5_mult_82_CARRYB_29__28_) );
  NOR2_X2 u5_mult_82_U2760 ( .A1(u5_mult_82_n6868), .A2(u5_mult_82_n6678), 
        .ZN(u5_mult_82_ab_30__28_) );
  INV_X4 u5_mult_82_U2759 ( .A(u5_mult_82_ab_29__32_), .ZN(u5_mult_82_n1907)
         );
  NOR2_X2 u5_mult_82_U2758 ( .A1(u5_mult_82_net64671), .A2(u5_mult_82_n6515), 
        .ZN(u5_mult_82_ab_3__22_) );
  NOR2_X2 u5_mult_82_U2757 ( .A1(u5_mult_82_net64689), .A2(u5_mult_82_n6515), 
        .ZN(u5_mult_82_ab_3__23_) );
  NOR2_X2 u5_mult_82_U2756 ( .A1(u5_mult_82_net64671), .A2(u5_mult_82_n6529), 
        .ZN(u5_mult_82_ab_7__22_) );
  NOR2_X2 u5_mult_82_U2755 ( .A1(u5_mult_82_net64689), .A2(u5_mult_82_n6529), 
        .ZN(u5_mult_82_ab_7__23_) );
  NOR2_X2 u5_mult_82_U2754 ( .A1(u5_mult_82_n6893), .A2(u5_mult_82_n6551), 
        .ZN(u5_mult_82_ab_10__24_) );
  NOR2_X1 u5_mult_82_U2753 ( .A1(u5_mult_82_n6882), .A2(u5_mult_82_n6558), 
        .ZN(u5_mult_82_ab_11__26_) );
  INV_X4 u5_mult_82_U2752 ( .A(u5_mult_82_ab_10__26_), .ZN(u5_mult_82_n4279)
         );
  INV_X4 u5_mult_82_U2751 ( .A(u5_mult_82_ab_22__23_), .ZN(u5_mult_82_net84453) );
  NOR2_X2 u5_mult_82_U2750 ( .A1(u5_mult_82_n6892), .A2(u5_mult_82_n6650), 
        .ZN(u5_mult_82_ab_26__24_) );
  NOR2_X2 u5_mult_82_U2749 ( .A1(u5_mult_82_net64901), .A2(u5_mult_82_n6671), 
        .ZN(u5_mult_82_ab_29__35_) );
  NOR2_X2 u5_mult_82_U2748 ( .A1(u5_mult_82_n6778), .A2(u5_mult_82_n6670), 
        .ZN(u5_mult_82_ab_29__48_) );
  NOR2_X1 u5_mult_82_U2747 ( .A1(u5_mult_82_n6982), .A2(u5_mult_82_n6666), 
        .ZN(u5_mult_82_ab_28__52_) );
  NOR2_X2 u5_mult_82_U2746 ( .A1(u5_mult_82_n6760), .A2(u5_mult_82_n6670), 
        .ZN(u5_mult_82_ab_29__51_) );
  NOR2_X2 u5_mult_82_U2745 ( .A1(u5_mult_82_n6773), .A2(u5_mult_82_n6670), 
        .ZN(u5_mult_82_ab_29__49_) );
  NOR2_X2 u5_mult_82_U2744 ( .A1(u5_mult_82_n6805), .A2(u5_mult_82_n6655), 
        .ZN(u5_mult_82_ab_27__44_) );
  NOR2_X2 u5_mult_82_U2743 ( .A1(u5_mult_82_n6886), .A2(u5_mult_82_net66091), 
        .ZN(u5_mult_82_ab_2__25_) );
  INV_X4 u5_mult_82_U2742 ( .A(u5_mult_82_ab_16__26_), .ZN(u5_mult_82_n2262)
         );
  NAND3_X2 u5_mult_82_U2741 ( .A1(u5_mult_82_n5972), .A2(u5_mult_82_n5973), 
        .A3(u5_mult_82_n5974), .ZN(u5_mult_82_CARRYB_25__25_) );
  NOR2_X2 u5_mult_82_U2740 ( .A1(u5_mult_82_n6876), .A2(u5_mult_82_n6657), 
        .ZN(u5_mult_82_ab_27__27_) );
  NOR2_X2 u5_mult_82_U2739 ( .A1(u5_mult_82_n6785), .A2(u5_mult_82_n6655), 
        .ZN(u5_mult_82_ab_27__47_) );
  NOR2_X2 u5_mult_82_U2738 ( .A1(u5_mult_82_n6798), .A2(u5_mult_82_n6655), 
        .ZN(u5_mult_82_ab_27__45_) );
  NOR2_X2 u5_mult_82_U2737 ( .A1(u5_mult_82_n6767), .A2(u5_mult_82_n6670), 
        .ZN(u5_mult_82_ab_29__50_) );
  INV_X4 u5_mult_82_U2736 ( .A(u5_mult_82_ab_7__24_), .ZN(u5_mult_82_n3238) );
  NAND3_X2 u5_mult_82_U2735 ( .A1(u5_mult_82_n3446), .A2(u5_mult_82_n3447), 
        .A3(u5_mult_82_n3448), .ZN(u5_mult_82_CARRYB_9__28_) );
  NAND3_X2 u5_mult_82_U2734 ( .A1(u5_mult_82_n3330), .A2(u5_mult_82_n3331), 
        .A3(u5_mult_82_n3332), .ZN(u5_mult_82_CARRYB_16__24_) );
  INV_X4 u5_mult_82_U2733 ( .A(u5_mult_82_ab_24__27_), .ZN(u5_mult_82_n1491)
         );
  NOR2_X2 u5_mult_82_U2732 ( .A1(u5_mult_82_n6844), .A2(u5_mult_82_n6649), 
        .ZN(u5_mult_82_ab_26__32_) );
  NOR2_X2 u5_mult_82_U2731 ( .A1(u5_mult_82_n6858), .A2(u5_mult_82_net65675), 
        .ZN(u5_mult_82_ab_25__30_) );
  NOR2_X2 u5_mult_82_U2730 ( .A1(u5_mult_82_n6851), .A2(u5_mult_82_net65675), 
        .ZN(u5_mult_82_ab_25__31_) );
  NOR2_X2 u5_mult_82_U2729 ( .A1(u5_mult_82_n6839), .A2(u5_mult_82_n6656), 
        .ZN(u5_mult_82_ab_27__33_) );
  NOR2_X1 u5_mult_82_U2728 ( .A1(u5_mult_82_n6817), .A2(u5_mult_82_net65717), 
        .ZN(u5_mult_82_ab_23__42_) );
  INV_X4 u5_mult_82_U2727 ( .A(u5_mult_82_ab_23__43_), .ZN(u5_mult_82_n2498)
         );
  NAND3_X2 u5_mult_82_U2726 ( .A1(u5_mult_82_n3031), .A2(u5_mult_82_n3032), 
        .A3(u5_mult_82_n3033), .ZN(u5_mult_82_CARRYB_24__40_) );
  NOR2_X2 u5_mult_82_U2725 ( .A1(u5_mult_82_n6805), .A2(u5_mult_82_n6644), 
        .ZN(u5_mult_82_ab_24__44_) );
  NOR2_X1 u5_mult_82_U2724 ( .A1(u5_mult_82_n6785), .A2(u5_mult_82_net65717), 
        .ZN(u5_mult_82_ab_23__47_) );
  NOR2_X1 u5_mult_82_U2723 ( .A1(u5_mult_82_n6881), .A2(u5_mult_82_n6615), 
        .ZN(u5_mult_82_ab_19__26_) );
  NOR2_X2 u5_mult_82_U2722 ( .A1(u5_mult_82_n6877), .A2(u5_mult_82_n6515), 
        .ZN(u5_mult_82_ab_3__27_) );
  NAND3_X2 u5_mult_82_U2721 ( .A1(u5_mult_82_n2192), .A2(u5_mult_82_n2193), 
        .A3(u5_mult_82_n2194), .ZN(u5_mult_82_CARRYB_22__25_) );
  NOR2_X2 u5_mult_82_U2720 ( .A1(u5_mult_82_n6832), .A2(u5_mult_82_n6642), 
        .ZN(u5_mult_82_ab_24__39_) );
  INV_X16 u5_mult_82_U2719 ( .A(u5_mult_82_n6854), .ZN(u5_mult_82_n6852) );
  NOR2_X2 u5_mult_82_U2718 ( .A1(u5_mult_82_n6870), .A2(u5_mult_82_n6578), 
        .ZN(u5_mult_82_ab_14__28_) );
  INV_X4 u5_mult_82_U2717 ( .A(u5_mult_82_ab_23__29_), .ZN(u5_mult_82_n1948)
         );
  NOR2_X2 u5_mult_82_U2716 ( .A1(u5_mult_82_n6761), .A2(u5_mult_82_n6641), 
        .ZN(u5_mult_82_ab_24__51_) );
  NOR2_X2 u5_mult_82_U2715 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_net65711), .ZN(u5_mult_82_ab_23__38_) );
  NAND3_X2 u5_mult_82_U2714 ( .A1(u5_mult_82_n2254), .A2(u5_mult_82_n2255), 
        .A3(u5_mult_82_n2256), .ZN(u5_mult_82_CARRYB_22__38_) );
  INV_X1 u5_mult_82_U2713 ( .A(u5_mult_82_ab_21__41_), .ZN(u5_mult_82_n4725)
         );
  NOR2_X2 u5_mult_82_U2712 ( .A1(u5_mult_82_n6863), .A2(u5_mult_82_n6601), 
        .ZN(u5_mult_82_ab_17__29_) );
  NOR2_X2 u5_mult_82_U2711 ( .A1(u5_mult_82_n6859), .A2(u5_mult_82_n6514), 
        .ZN(u5_mult_82_ab_3__30_) );
  NOR2_X2 u5_mult_82_U2710 ( .A1(u5_mult_82_n6852), .A2(u5_mult_82_net66017), 
        .ZN(u5_mult_82_ab_6__31_) );
  NOR2_X2 u5_mult_82_U2709 ( .A1(u5_mult_82_n6840), .A2(u5_mult_82_net66089), 
        .ZN(u5_mult_82_ab_2__33_) );
  NOR2_X2 u5_mult_82_U2708 ( .A1(u5_mult_82_net64887), .A2(u5_mult_82_net66089), .ZN(u5_mult_82_ab_2__34_) );
  NOR2_X1 u5_mult_82_U2707 ( .A1(u5_mult_82_n6844), .A2(u5_mult_82_n6628), 
        .ZN(u5_mult_82_ab_21__32_) );
  NOR2_X2 u5_mult_82_U2706 ( .A1(u5_mult_82_n6851), .A2(u5_mult_82_n6628), 
        .ZN(u5_mult_82_ab_21__31_) );
  NOR2_X1 u5_mult_82_U2705 ( .A1(u5_mult_82_net64903), .A2(u5_mult_82_n6621), 
        .ZN(u5_mult_82_ab_20__35_) );
  NOR2_X2 u5_mult_82_U2704 ( .A1(u5_mult_82_n6768), .A2(u5_mult_82_n6627), 
        .ZN(u5_mult_82_ab_21__50_) );
  NOR2_X2 u5_mult_82_U2703 ( .A1(u5_mult_82_n6779), .A2(u5_mult_82_n6607), 
        .ZN(u5_mult_82_ab_18__48_) );
  INV_X4 u5_mult_82_U2702 ( .A(u5_mult_82_ab_15__29_), .ZN(u5_mult_82_n5219)
         );
  INV_X4 u5_mult_82_U2701 ( .A(u5_mult_82_n6847), .ZN(u5_mult_82_n6846) );
  NOR2_X2 u5_mult_82_U2700 ( .A1(u5_mult_82_n6852), .A2(u5_mult_82_n6550), 
        .ZN(u5_mult_82_ab_10__31_) );
  NOR2_X1 u5_mult_82_U2699 ( .A1(u5_mult_82_n6858), .A2(u5_mult_82_n6614), 
        .ZN(u5_mult_82_ab_19__30_) );
  NAND2_X2 u5_mult_82_U2698 ( .A1(u5_mult_82_ab_19__44_), .A2(
        u5_mult_82_SUMB_18__45_), .ZN(u5_mult_82_n5878) );
  NOR2_X2 u5_mult_82_U2697 ( .A1(u5_mult_82_n6852), .A2(u5_mult_82_n6578), 
        .ZN(u5_mult_82_ab_14__31_) );
  NOR2_X2 u5_mult_82_U2696 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6621), 
        .ZN(u5_mult_82_ab_20__38_) );
  NAND3_X2 u5_mult_82_U2695 ( .A1(u5_mult_82_n4411), .A2(u5_mult_82_n4412), 
        .A3(u5_mult_82_n4413), .ZN(u5_mult_82_CARRYB_19__38_) );
  NOR2_X2 u5_mult_82_U2694 ( .A1(u5_mult_82_n6812), .A2(u5_mult_82_n6600), 
        .ZN(u5_mult_82_ab_17__43_) );
  NOR2_X2 u5_mult_82_U2693 ( .A1(u5_mult_82_n6805), .A2(u5_mult_82_n6607), 
        .ZN(u5_mult_82_ab_18__44_) );
  NOR2_X2 u5_mult_82_U2692 ( .A1(u5_mult_82_n6828), .A2(u5_mult_82_n6607), 
        .ZN(u5_mult_82_ab_18__40_) );
  NOR2_X1 u5_mult_82_U2691 ( .A1(u5_mult_82_n6840), .A2(u5_mult_82_n6571), 
        .ZN(u5_mult_82_ab_13__33_) );
  NOR2_X2 u5_mult_82_U2690 ( .A1(u5_mult_82_n6840), .A2(u5_mult_82_net66017), 
        .ZN(u5_mult_82_ab_6__33_) );
  NOR2_X2 u5_mult_82_U2689 ( .A1(u5_mult_82_n6839), .A2(u5_mult_82_n6601), 
        .ZN(u5_mult_82_ab_17__33_) );
  INV_X4 u5_mult_82_U2688 ( .A(u5_mult_82_ab_17__35_), .ZN(u5_mult_82_n5221)
         );
  NOR2_X2 u5_mult_82_U2687 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6601), 
        .ZN(u5_mult_82_ab_17__38_) );
  NAND3_X2 u5_mult_82_U2686 ( .A1(u5_mult_82_n4609), .A2(u5_mult_82_n4610), 
        .A3(u5_mult_82_n4611), .ZN(u5_mult_82_CARRYB_15__47_) );
  NAND2_X2 u5_mult_82_U2685 ( .A1(u5_mult_82_n3364), .A2(u5_mult_82_n3365), 
        .ZN(u5_mult_82_SUMB_15__48_) );
  NOR2_X2 u5_mult_82_U2684 ( .A1(u5_mult_82_n6785), .A2(u5_mult_82_n6593), 
        .ZN(u5_mult_82_ab_16__47_) );
  INV_X4 u5_mult_82_U2683 ( .A(u5_mult_82_net66089), .ZN(u5_mult_82_net86863)
         );
  INV_X4 u5_mult_82_U2682 ( .A(u5_mult_82_ab_16__35_), .ZN(u5_mult_82_n4906)
         );
  NOR2_X1 u5_mult_82_U2681 ( .A1(u5_mult_82_n6769), .A2(u5_mult_82_n6571), 
        .ZN(u5_mult_82_ab_13__50_) );
  NOR2_X2 u5_mult_82_U2680 ( .A1(u5_mult_82_net64941), .A2(u5_mult_82_n6514), 
        .ZN(u5_mult_82_ab_3__37_) );
  NOR2_X1 u5_mult_82_U2679 ( .A1(u5_mult_82_net64959), .A2(u5_mult_82_n6578), 
        .ZN(u5_mult_82_ab_14__38_) );
  NOR2_X2 u5_mult_82_U2678 ( .A1(u5_mult_82_net64941), .A2(u5_mult_82_n6578), 
        .ZN(u5_mult_82_ab_14__37_) );
  NOR2_X2 u5_mult_82_U2677 ( .A1(u5_mult_82_net64959), .A2(u5_mult_82_n6586), 
        .ZN(u5_mult_82_ab_15__38_) );
  INV_X4 u5_mult_82_U2676 ( .A(u5_mult_82_ab_14__39_), .ZN(u5_mult_82_n960) );
  NAND3_X2 u5_mult_82_U2675 ( .A1(u5_mult_82_n5387), .A2(u5_mult_82_n5386), 
        .A3(u5_mult_82_n5385), .ZN(u5_mult_82_CARRYB_14__40_) );
  NAND3_X2 u5_mult_82_U2674 ( .A1(u5_mult_82_n5352), .A2(u5_mult_82_n5353), 
        .A3(u5_mult_82_n5354), .ZN(u5_mult_82_CARRYB_14__39_) );
  INV_X4 u5_mult_82_U2673 ( .A(u5_mult_82_ab_14__40_), .ZN(u5_mult_82_n3442)
         );
  NOR2_X2 u5_mult_82_U2672 ( .A1(u5_mult_82_n6775), .A2(u5_mult_82_n6564), 
        .ZN(u5_mult_82_ab_12__49_) );
  NOR2_X2 u5_mult_82_U2671 ( .A1(u5_mult_82_net64941), .A2(u5_mult_82_n6544), 
        .ZN(u5_mult_82_ab_9__37_) );
  NAND3_X2 u5_mult_82_U2670 ( .A1(u5_mult_82_n6379), .A2(u5_mult_82_n6380), 
        .A3(u5_mult_82_n6381), .ZN(u5_mult_82_CARRYB_12__45_) );
  NOR2_X2 u5_mult_82_U2669 ( .A1(u5_mult_82_n6780), .A2(u5_mult_82_n6564), 
        .ZN(u5_mult_82_ab_12__48_) );
  NOR2_X2 u5_mult_82_U2668 ( .A1(u5_mult_82_n6786), .A2(u5_mult_82_n6559), 
        .ZN(u5_mult_82_ab_11__47_) );
  INV_X4 u5_mult_82_U2667 ( .A(u5_mult_82_n1762), .ZN(u5_mult_82_n1763) );
  NAND2_X2 u5_mult_82_U2666 ( .A1(u5_mult_82_n1227), .A2(u5_mult_82_n1228), 
        .ZN(u5_mult_82_SUMB_11__38_) );
  NOR2_X2 u5_mult_82_U2665 ( .A1(u5_mult_82_n6833), .A2(u5_mult_82_net66089), 
        .ZN(u5_mult_82_ab_2__39_) );
  NOR2_X1 u5_mult_82_U2664 ( .A1(u5_mult_82_n6823), .A2(u5_mult_82_n6552), 
        .ZN(u5_mult_82_ab_10__41_) );
  NOR2_X1 u5_mult_82_U2663 ( .A1(u5_mult_82_n6806), .A2(u5_mult_82_n6543), 
        .ZN(u5_mult_82_ab_9__44_) );
  NOR2_X2 u5_mult_82_U2662 ( .A1(u5_mult_82_n6829), .A2(u5_mult_82_net66087), 
        .ZN(u5_mult_82_ab_2__40_) );
  INV_X4 u5_mult_82_U2661 ( .A(u5_mult_82_ab_8__40_), .ZN(u5_mult_82_n857) );
  NOR2_X1 u5_mult_82_U2660 ( .A1(u5_mult_82_n6833), .A2(u5_mult_82_n6535), 
        .ZN(u5_mult_82_ab_8__39_) );
  NOR2_X2 u5_mult_82_U2659 ( .A1(u5_mult_82_n6813), .A2(u5_mult_82_n6543), 
        .ZN(u5_mult_82_ab_9__43_) );
  NOR2_X2 u5_mult_82_U2658 ( .A1(u5_mult_82_n6829), .A2(u5_mult_82_n6543), 
        .ZN(u5_mult_82_ab_9__40_) );
  INV_X4 u5_mult_82_U2657 ( .A(u5_mult_82_ab_8__47_), .ZN(u5_mult_82_n1764) );
  NOR2_X2 u5_mult_82_U2656 ( .A1(u5_mult_82_n6762), .A2(u5_mult_82_n6527), 
        .ZN(u5_mult_82_ab_7__51_) );
  NOR2_X2 u5_mult_82_U2655 ( .A1(u5_mult_82_n6769), .A2(u5_mult_82_n6528), 
        .ZN(u5_mult_82_ab_7__50_) );
  NOR2_X2 u5_mult_82_U2654 ( .A1(u5_mult_82_n6818), .A2(u5_mult_82_n6513), 
        .ZN(u5_mult_82_ab_3__42_) );
  NOR2_X1 u5_mult_82_U2653 ( .A1(u5_mult_82_n6806), .A2(u5_mult_82_net66087), 
        .ZN(u5_mult_82_ab_2__44_) );
  NOR2_X2 u5_mult_82_U2652 ( .A1(u5_mult_82_n6775), .A2(u5_mult_82_n6513), 
        .ZN(u5_mult_82_ab_3__49_) );
  NOR2_X2 u5_mult_82_U2651 ( .A1(u5_mult_82_n6799), .A2(u5_mult_82_n6513), 
        .ZN(u5_mult_82_ab_3__45_) );
  NOR2_X2 u5_mult_82_U2650 ( .A1(u5_mult_82_n6780), .A2(u5_mult_82_n6513), 
        .ZN(u5_mult_82_ab_3__48_) );
  NAND3_X2 u5_mult_82_U2649 ( .A1(u5_mult_82_n1929), .A2(u5_mult_82_n1930), 
        .A3(u5_mult_82_n1931), .ZN(u5_mult_82_CARRYB_2__47_) );
  NOR2_X2 u5_mult_82_U2648 ( .A1(u5_mult_82_n6989), .A2(u5_mult_82_n6516), 
        .ZN(u5_mult_82_ab_3__0_) );
  NOR2_X1 u5_mult_82_U2647 ( .A1(u5_mult_82_n6989), .A2(u5_mult_82_n6538), 
        .ZN(u5_mult_82_ab_8__0_) );
  NOR2_X2 u5_mult_82_U2646 ( .A1(u5_mult_82_n6989), .A2(u5_mult_82_n6574), 
        .ZN(u5_mult_82_ab_13__0_) );
  NOR2_X2 u5_mult_82_U2645 ( .A1(u5_mult_82_n6988), .A2(u5_mult_82_n6611), 
        .ZN(u5_mult_82_ab_18__0_) );
  NOR2_X1 u5_mult_82_U2644 ( .A1(u5_mult_82_n6988), .A2(u5_mult_82_net65717), 
        .ZN(u5_mult_82_ab_23__0_) );
  NOR2_X1 u5_mult_82_U2643 ( .A1(u5_mult_82_n6987), .A2(u5_mult_82_n6666), 
        .ZN(u5_mult_82_ab_28__0_) );
  NOR2_X2 u5_mult_82_U2642 ( .A1(u5_mult_82_n6987), .A2(u5_mult_82_n6702), 
        .ZN(u5_mult_82_ab_33__0_) );
  NOR2_X2 u5_mult_82_U2641 ( .A1(u5_mult_82_n6987), .A2(u5_mult_82_net65447), 
        .ZN(u5_mult_82_ab_38__0_) );
  NOR2_X2 u5_mult_82_U2640 ( .A1(u5_mult_82_n6986), .A2(u5_mult_82_net65321), 
        .ZN(u5_mult_82_ab_45__0_) );
  NOR2_X1 u5_mult_82_U2639 ( .A1(u5_mult_82_n6986), .A2(u5_mult_82_net65189), 
        .ZN(u5_mult_82_ab_51__0_) );
  NOR2_X2 u5_mult_82_U2638 ( .A1(u5_mult_82_n6969), .A2(u5_mult_82_n6516), 
        .ZN(u5_mult_82_ab_3__1_) );
  NOR2_X1 u5_mult_82_U2637 ( .A1(u5_mult_82_n6969), .A2(u5_mult_82_n6538), 
        .ZN(u5_mult_82_ab_8__1_) );
  NOR2_X2 u5_mult_82_U2636 ( .A1(u5_mult_82_n6969), .A2(u5_mult_82_n6574), 
        .ZN(u5_mult_82_ab_13__1_) );
  NOR2_X2 u5_mult_82_U2635 ( .A1(u5_mult_82_n6968), .A2(u5_mult_82_n6611), 
        .ZN(u5_mult_82_ab_18__1_) );
  INV_X16 u5_mult_82_U2634 ( .A(u5_mult_82_n6625), .ZN(u5_mult_82_n6624) );
  NOR2_X1 u5_mult_82_U2633 ( .A1(u5_mult_82_n6968), .A2(u5_mult_82_net65717), 
        .ZN(u5_mult_82_ab_23__1_) );
  NOR2_X1 u5_mult_82_U2632 ( .A1(u5_mult_82_n6967), .A2(u5_mult_82_n6666), 
        .ZN(u5_mult_82_ab_28__1_) );
  NOR2_X1 u5_mult_82_U2631 ( .A1(u5_mult_82_n6967), .A2(u5_mult_82_n6702), 
        .ZN(u5_mult_82_ab_33__1_) );
  INV_X1 u5_mult_82_U2630 ( .A(u5_mult_82_ab_38__1_), .ZN(u5_mult_82_n631) );
  NOR2_X2 u5_mult_82_U2629 ( .A1(u5_mult_82_n6961), .A2(u5_mult_82_net65411), 
        .ZN(u5_mult_82_ab_40__2_) );
  NOR2_X1 u5_mult_82_U2628 ( .A1(u5_mult_82_n6974), .A2(u5_mult_82_n6967), 
        .ZN(u5_mult_82_ab_52__1_) );
  NOR2_X1 u5_mult_82_U2627 ( .A1(u5_mult_82_n6967), .A2(u5_mult_82_n6743), 
        .ZN(u5_mult_82_ab_46__1_) );
  NOR2_X2 u5_mult_82_U2626 ( .A1(u5_mult_82_n6962), .A2(u5_mult_82_n6516), 
        .ZN(u5_mult_82_ab_3__2_) );
  INV_X8 u5_mult_82_U2625 ( .A(u5_mult_82_n1359), .ZN(u5_mult_82_net66025) );
  NOR2_X1 u5_mult_82_U2624 ( .A1(u5_mult_82_n6962), .A2(u5_mult_82_n6538), 
        .ZN(u5_mult_82_ab_8__2_) );
  INV_X8 u5_mult_82_U2623 ( .A(u5_mult_82_n6556), .ZN(u5_mult_82_n6561) );
  NOR2_X2 u5_mult_82_U2622 ( .A1(u5_mult_82_n6962), .A2(u5_mult_82_n6574), 
        .ZN(u5_mult_82_ab_13__2_) );
  NOR2_X2 u5_mult_82_U2621 ( .A1(u5_mult_82_n6961), .A2(u5_mult_82_n6611), 
        .ZN(u5_mult_82_ab_18__2_) );
  INV_X8 u5_mult_82_U2620 ( .A(u5_mult_82_n6627), .ZN(u5_mult_82_n6632) );
  NOR2_X1 u5_mult_82_U2619 ( .A1(u5_mult_82_n6961), .A2(u5_mult_82_net65717), 
        .ZN(u5_mult_82_ab_23__2_) );
  NOR2_X1 u5_mult_82_U2618 ( .A1(u5_mult_82_n6960), .A2(u5_mult_82_n6666), 
        .ZN(u5_mult_82_ab_28__2_) );
  INV_X8 u5_mult_82_U2617 ( .A(u5_mult_82_n6683), .ZN(u5_mult_82_n6688) );
  NOR2_X1 u5_mult_82_U2616 ( .A1(u5_mult_82_n6960), .A2(u5_mult_82_n6702), 
        .ZN(u5_mult_82_ab_33__2_) );
  INV_X8 u5_mult_82_U2615 ( .A(u5_mult_82_n6719), .ZN(u5_mult_82_n6724) );
  INV_X16 u5_mult_82_U2614 ( .A(u5_mult_82_n1326), .ZN(u5_mult_82_net65393) );
  NOR2_X1 u5_mult_82_U2613 ( .A1(u5_mult_82_n6974), .A2(u5_mult_82_n6960), 
        .ZN(u5_mult_82_ab_52__2_) );
  INV_X4 u5_mult_82_U2612 ( .A(u5_mult_82_n6398), .ZN(u5_mult_82_CLA_SUM[64])
         );
  NAND2_X2 u5_mult_82_U2611 ( .A1(u5_mult_82_n3608), .A2(u5_mult_82_n3609), 
        .ZN(u5_mult_82_SUMB_51__25_) );
  NOR2_X1 u5_mult_82_U2610 ( .A1(u5_mult_82_n6975), .A2(u5_mult_82_n6891), 
        .ZN(u5_mult_82_ab_52__24_) );
  NOR2_X1 u5_mult_82_U2609 ( .A1(u5_mult_82_n6975), .A2(u5_mult_82_net64683), 
        .ZN(u5_mult_82_ab_52__23_) );
  INV_X16 u5_mult_82_U2608 ( .A(n4802), .ZN(u5_mult_82_n1268) );
  NOR2_X2 u5_mult_82_U2607 ( .A1(u5_mult_82_n6955), .A2(u5_mult_82_n6516), 
        .ZN(u5_mult_82_ab_3__3_) );
  NOR2_X1 u5_mult_82_U2606 ( .A1(u5_mult_82_n6955), .A2(u5_mult_82_n6538), 
        .ZN(u5_mult_82_ab_8__3_) );
  NOR2_X2 u5_mult_82_U2605 ( .A1(u5_mult_82_n6955), .A2(u5_mult_82_n6574), 
        .ZN(u5_mult_82_ab_13__3_) );
  NOR2_X2 u5_mult_82_U2604 ( .A1(u5_mult_82_n6954), .A2(u5_mult_82_n6611), 
        .ZN(u5_mult_82_ab_18__3_) );
  NOR2_X1 u5_mult_82_U2603 ( .A1(u5_mult_82_n6954), .A2(u5_mult_82_net65717), 
        .ZN(u5_mult_82_ab_23__3_) );
  INV_X8 u5_mult_82_U2602 ( .A(fracta_mul[27]), .ZN(u5_mult_82_n6654) );
  NOR2_X2 u5_mult_82_U2601 ( .A1(u5_mult_82_n6954), .A2(u5_mult_82_net65681), 
        .ZN(u5_mult_82_ab_25__3_) );
  NOR2_X1 u5_mult_82_U2600 ( .A1(u5_mult_82_n6953), .A2(u5_mult_82_n6666), 
        .ZN(u5_mult_82_ab_28__3_) );
  NOR2_X2 u5_mult_82_U2599 ( .A1(u5_mult_82_n6953), .A2(u5_mult_82_n6702), 
        .ZN(u5_mult_82_ab_33__3_) );
  INV_X16 u5_mult_82_U2598 ( .A(u5_mult_82_n1375), .ZN(u5_mult_82_n1374) );
  INV_X4 u5_mult_82_U2597 ( .A(u5_mult_82_n1675), .ZN(u5_mult_82_SUMB_41__3_)
         );
  NOR2_X2 u5_mult_82_U2596 ( .A1(u5_mult_82_n6952), .A2(u5_mult_82_net65375), 
        .ZN(u5_mult_82_ab_42__3_) );
  INV_X4 u5_mult_82_U2595 ( .A(u5_mult_82_ab_46__3_), .ZN(u5_mult_82_n3193) );
  NOR2_X1 u5_mult_82_U2594 ( .A1(u5_mult_82_n6974), .A2(u5_mult_82_n6952), 
        .ZN(u5_mult_82_ab_52__3_) );
  NOR2_X1 u5_mult_82_U2593 ( .A1(u5_mult_82_n6974), .A2(u5_mult_82_n6946), 
        .ZN(u5_mult_82_ab_52__4_) );
  INV_X4 u5_mult_82_U2592 ( .A(u5_mult_82_ab_52__5_), .ZN(u5_mult_82_net87687)
         );
  NAND3_X2 u5_mult_82_U2591 ( .A1(u5_mult_82_net80806), .A2(
        u5_mult_82_net80807), .A3(u5_mult_82_net80808), .ZN(
        u5_mult_82_CARRYB_51__6_) );
  NOR2_X1 u5_mult_82_U2590 ( .A1(u5_mult_82_n6974), .A2(u5_mult_82_net64379), 
        .ZN(u5_mult_82_ab_52__6_) );
  NOR2_X1 u5_mult_82_U2589 ( .A1(u5_mult_82_n6975), .A2(u5_mult_82_net64505), 
        .ZN(u5_mult_82_ab_52__13_) );
  NOR2_X1 u5_mult_82_U2588 ( .A1(u5_mult_82_n6975), .A2(u5_mult_82_net64523), 
        .ZN(u5_mult_82_ab_52__14_) );
  NOR2_X1 u5_mult_82_U2587 ( .A1(u5_mult_82_n6975), .A2(u5_mult_82_net64665), 
        .ZN(u5_mult_82_ab_52__22_) );
  NOR2_X1 u5_mult_82_U2586 ( .A1(u5_mult_82_n6976), .A2(u5_mult_82_n6867), 
        .ZN(u5_mult_82_ab_52__28_) );
  NOR2_X1 u5_mult_82_U2585 ( .A1(u5_mult_82_n6976), .A2(u5_mult_82_n6861), 
        .ZN(u5_mult_82_ab_52__29_) );
  NOR2_X2 u5_mult_82_U2584 ( .A1(u5_mult_82_n6976), .A2(u5_mult_82_net64899), 
        .ZN(u5_mult_82_ab_52__35_) );
  NOR2_X1 u5_mult_82_U2583 ( .A1(u5_mult_82_n6976), .A2(u5_mult_82_net64921), 
        .ZN(u5_mult_82_ab_52__36_) );
  NOR2_X1 u5_mult_82_U2582 ( .A1(u5_mult_82_n6977), .A2(u5_mult_82_n6797), 
        .ZN(u5_mult_82_ab_52__45_) );
  NOR2_X1 u5_mult_82_U2581 ( .A1(u5_mult_82_n6977), .A2(u5_mult_82_n6803), 
        .ZN(u5_mult_82_ab_52__44_) );
  NOR2_X1 u5_mult_82_U2580 ( .A1(u5_mult_82_n6983), .A2(u5_mult_82_n6755), 
        .ZN(u5_mult_82_ab_49__52_) );
  NOR2_X1 u5_mult_82_U2579 ( .A1(u5_mult_82_n6759), .A2(u5_mult_82_net65223), 
        .ZN(u5_mult_82_ab_50__51_) );
  NOR2_X1 u5_mult_82_U2578 ( .A1(u5_mult_82_n6977), .A2(u5_mult_82_n6816), 
        .ZN(u5_mult_82_ab_52__42_) );
  NOR2_X1 u5_mult_82_U2577 ( .A1(u5_mult_82_n6977), .A2(u5_mult_82_n6784), 
        .ZN(u5_mult_82_ab_52__47_) );
  NOR2_X1 u5_mult_82_U2576 ( .A1(u5_mult_82_n6977), .A2(u5_mult_82_n6826), 
        .ZN(u5_mult_82_ab_52__40_) );
  NOR2_X2 u5_mult_82_U2575 ( .A1(u5_mult_82_n6948), .A2(u5_mult_82_n6516), 
        .ZN(u5_mult_82_ab_3__4_) );
  NOR2_X2 u5_mult_82_U2574 ( .A1(u5_mult_82_n6948), .A2(u5_mult_82_n6537), 
        .ZN(u5_mult_82_ab_8__4_) );
  NOR2_X1 u5_mult_82_U2573 ( .A1(u5_mult_82_n6948), .A2(u5_mult_82_n6573), 
        .ZN(u5_mult_82_ab_13__4_) );
  NOR2_X2 u5_mult_82_U2572 ( .A1(u5_mult_82_n6947), .A2(u5_mult_82_n6610), 
        .ZN(u5_mult_82_ab_18__4_) );
  NOR2_X1 u5_mult_82_U2571 ( .A1(u5_mult_82_net64363), .A2(u5_mult_82_net65713), .ZN(u5_mult_82_ab_23__5_) );
  NOR2_X1 u5_mult_82_U2570 ( .A1(u5_mult_82_n6946), .A2(u5_mult_82_n6665), 
        .ZN(u5_mult_82_ab_28__4_) );
  INV_X8 u5_mult_82_U2569 ( .A(fracta_mul[43]), .ZN(u5_mult_82_n1375) );
  NAND3_X2 u5_mult_82_U2568 ( .A1(u5_mult_82_n4512), .A2(u5_mult_82_n4513), 
        .A3(u5_mult_82_n4514), .ZN(u5_mult_82_CARRYB_46__3_) );
  NAND3_X2 u5_mult_82_U2567 ( .A1(u5_mult_82_n4661), .A2(u5_mult_82_n4660), 
        .A3(u5_mult_82_n4659), .ZN(u5_mult_82_CARRYB_46__5_) );
  INV_X4 u5_mult_82_U2566 ( .A(u5_mult_82_ab_46__6_), .ZN(u5_mult_82_n4852) );
  INV_X4 u5_mult_82_U2565 ( .A(u5_mult_82_ab_50__9_), .ZN(u5_mult_82_n731) );
  NOR2_X1 u5_mult_82_U2564 ( .A1(u5_mult_82_net64433), .A2(u5_mult_82_net65191), .ZN(u5_mult_82_ab_51__9_) );
  NOR2_X1 u5_mult_82_U2563 ( .A1(u5_mult_82_net64455), .A2(u5_mult_82_net65189), .ZN(u5_mult_82_ab_51__10_) );
  INV_X4 u5_mult_82_U2562 ( .A(u5_mult_82_ab_51__18_), .ZN(u5_mult_82_n3960)
         );
  NAND2_X2 u5_mult_82_U2561 ( .A1(u5_mult_82_ab_50__18_), .A2(
        u5_mult_82_SUMB_49__19_), .ZN(u5_mult_82_n5742) );
  NOR2_X1 u5_mult_82_U2560 ( .A1(u5_mult_82_n6975), .A2(u5_mult_82_n6903), 
        .ZN(u5_mult_82_ab_52__20_) );
  NOR2_X1 u5_mult_82_U2559 ( .A1(u5_mult_82_n6975), .A2(u5_mult_82_n6895), 
        .ZN(u5_mult_82_ab_52__21_) );
  NOR2_X1 u5_mult_82_U2558 ( .A1(u5_mult_82_n6849), .A2(u5_mult_82_net65191), 
        .ZN(u5_mult_82_ab_51__31_) );
  NOR2_X1 u5_mult_82_U2557 ( .A1(u5_mult_82_net64881), .A2(u5_mult_82_net65191), .ZN(u5_mult_82_ab_51__34_) );
  NOR2_X1 u5_mult_82_U2556 ( .A1(u5_mult_82_n6772), .A2(u5_mult_82_net65189), 
        .ZN(u5_mult_82_ab_51__49_) );
  NOR2_X1 u5_mult_82_U2555 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_net65193), .ZN(u5_mult_82_ab_51__38_) );
  NOR2_X1 u5_mult_82_U2554 ( .A1(u5_mult_82_n6831), .A2(u5_mult_82_net65193), 
        .ZN(u5_mult_82_ab_51__39_) );
  INV_X16 u5_mult_82_U2553 ( .A(u5_mult_82_n7018), .ZN(u5_mult_82_n6889) );
  NOR2_X1 u5_mult_82_U2552 ( .A1(u5_mult_82_n6874), .A2(u5_mult_82_net65229), 
        .ZN(u5_mult_82_ab_50__27_) );
  NOR2_X2 u5_mult_82_U2551 ( .A1(u5_mult_82_n6874), .A2(u5_mult_82_n6754), 
        .ZN(u5_mult_82_ab_49__27_) );
  NOR2_X1 u5_mult_82_U2550 ( .A1(u5_mult_82_n6884), .A2(u5_mult_82_net65191), 
        .ZN(u5_mult_82_ab_51__25_) );
  NOR2_X1 u5_mult_82_U2549 ( .A1(u5_mult_82_n6952), .A2(u5_mult_82_n6737), 
        .ZN(u5_mult_82_ab_44__3_) );
  NOR2_X2 u5_mult_82_U2548 ( .A1(u5_mult_82_net64365), .A2(u5_mult_82_n6516), 
        .ZN(u5_mult_82_ab_3__5_) );
  NOR2_X2 u5_mult_82_U2547 ( .A1(u5_mult_82_net64365), .A2(u5_mult_82_n6537), 
        .ZN(u5_mult_82_ab_8__5_) );
  NOR2_X1 u5_mult_82_U2546 ( .A1(u5_mult_82_net64365), .A2(u5_mult_82_n6573), 
        .ZN(u5_mult_82_ab_13__5_) );
  NOR2_X2 u5_mult_82_U2545 ( .A1(u5_mult_82_net64381), .A2(u5_mult_82_n6603), 
        .ZN(u5_mult_82_ab_17__6_) );
  NOR2_X1 u5_mult_82_U2544 ( .A1(u5_mult_82_net64381), .A2(u5_mult_82_net65717), .ZN(u5_mult_82_ab_23__6_) );
  NOR2_X1 u5_mult_82_U2543 ( .A1(u5_mult_82_n6940), .A2(u5_mult_82_n6686), 
        .ZN(u5_mult_82_ab_31__7_) );
  NOR2_X2 u5_mult_82_U2542 ( .A1(u5_mult_82_n6940), .A2(u5_mult_82_n6709), 
        .ZN(u5_mult_82_ab_35__7_) );
  NOR2_X1 u5_mult_82_U2541 ( .A1(u5_mult_82_net64415), .A2(u5_mult_82_net65189), .ZN(u5_mult_82_ab_51__8_) );
  INV_X4 u5_mult_82_U2540 ( .A(u5_mult_82_ab_49__13_), .ZN(u5_mult_82_n2173)
         );
  NOR2_X1 u5_mult_82_U2539 ( .A1(u5_mult_82_n6919), .A2(u5_mult_82_net65189), 
        .ZN(u5_mult_82_ab_51__18_) );
  NOR2_X1 u5_mult_82_U2538 ( .A1(u5_mult_82_n6903), .A2(u5_mult_82_n6754), 
        .ZN(u5_mult_82_ab_49__20_) );
  NOR2_X1 u5_mult_82_U2537 ( .A1(u5_mult_82_n6912), .A2(u5_mult_82_net65189), 
        .ZN(u5_mult_82_ab_51__19_) );
  NOR2_X1 u5_mult_82_U2536 ( .A1(u5_mult_82_n6837), .A2(u5_mult_82_net65191), 
        .ZN(u5_mult_82_ab_51__33_) );
  NOR2_X1 u5_mult_82_U2535 ( .A1(u5_mult_82_n6837), .A2(u5_mult_82_net65225), 
        .ZN(u5_mult_82_ab_50__33_) );
  NOR2_X2 u5_mult_82_U2534 ( .A1(u5_mult_82_net64383), .A2(u5_mult_82_n6516), 
        .ZN(u5_mult_82_ab_3__6_) );
  NOR2_X2 u5_mult_82_U2533 ( .A1(u5_mult_82_net64383), .A2(u5_mult_82_n6537), 
        .ZN(u5_mult_82_ab_8__6_) );
  NOR2_X2 u5_mult_82_U2532 ( .A1(u5_mult_82_net64381), .A2(u5_mult_82_n6644), 
        .ZN(u5_mult_82_ab_24__6_) );
  NOR2_X2 u5_mult_82_U2531 ( .A1(u5_mult_82_n6941), .A2(u5_mult_82_n6651), 
        .ZN(u5_mult_82_ab_26__7_) );
  INV_X8 u5_mult_82_U2530 ( .A(n4729), .ZN(u5_mult_82_n7020) );
  NOR2_X2 u5_mult_82_U2529 ( .A1(u5_mult_82_n6879), .A2(u5_mult_82_net65285), 
        .ZN(u5_mult_82_ab_47__26_) );
  INV_X8 u5_mult_82_U2528 ( .A(n4783), .ZN(u5_mult_82_net64949) );
  NOR2_X2 u5_mult_82_U2527 ( .A1(u5_mult_82_n6942), .A2(u5_mult_82_n6516), 
        .ZN(u5_mult_82_ab_3__7_) );
  NOR2_X2 u5_mult_82_U2526 ( .A1(u5_mult_82_n6942), .A2(u5_mult_82_n6537), 
        .ZN(u5_mult_82_ab_8__7_) );
  NOR2_X2 u5_mult_82_U2525 ( .A1(u5_mult_82_net64417), .A2(u5_mult_82_n6610), 
        .ZN(u5_mult_82_ab_18__8_) );
  NOR2_X1 u5_mult_82_U2524 ( .A1(u5_mult_82_net64433), .A2(u5_mult_82_n6680), 
        .ZN(u5_mult_82_ab_30__9_) );
  NOR2_X2 u5_mult_82_U2523 ( .A1(u5_mult_82_net64415), .A2(u5_mult_82_n6709), 
        .ZN(u5_mult_82_ab_35__8_) );
  NAND2_X2 u5_mult_82_U2522 ( .A1(u5_mult_82_n2982), .A2(u5_mult_82_n2983), 
        .ZN(u5_mult_82_n5820) );
  INV_X4 u5_mult_82_U2521 ( .A(u5_mult_82_n1754), .ZN(u5_mult_82_n1755) );
  INV_X2 u5_mult_82_U2520 ( .A(u5_mult_82_ab_42__8_), .ZN(u5_mult_82_n3589) );
  NOR2_X1 u5_mult_82_U2519 ( .A1(u5_mult_82_net64415), .A2(u5_mult_82_net65283), .ZN(u5_mult_82_ab_47__8_) );
  INV_X4 u5_mult_82_U2518 ( .A(u5_mult_82_ab_46__18_), .ZN(u5_mult_82_n2329)
         );
  INV_X4 u5_mult_82_U2517 ( .A(u5_mult_82_ab_47__17_), .ZN(u5_mult_82_n2595)
         );
  INV_X8 u5_mult_82_U2516 ( .A(n4748), .ZN(u5_mult_82_n6894) );
  INV_X4 u5_mult_82_U2515 ( .A(u5_mult_82_ab_48__31_), .ZN(u5_mult_82_n2127)
         );
  INV_X4 u5_mult_82_U2514 ( .A(u5_mult_82_n2709), .ZN(u5_mult_82_n2710) );
  NOR2_X2 u5_mult_82_U2513 ( .A1(u5_mult_82_n6826), .A2(u5_mult_82_net65313), 
        .ZN(u5_mult_82_ab_45__40_) );
  NOR2_X1 u5_mult_82_U2512 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6742), 
        .ZN(u5_mult_82_ab_46__38_) );
  NOR2_X2 u5_mult_82_U2511 ( .A1(u5_mult_82_n6856), .A2(u5_mult_82_n6734), 
        .ZN(u5_mult_82_ab_44__30_) );
  NOR2_X2 u5_mult_82_U2510 ( .A1(u5_mult_82_net64419), .A2(u5_mult_82_n6516), 
        .ZN(u5_mult_82_ab_3__8_) );
  NOR2_X2 u5_mult_82_U2509 ( .A1(u5_mult_82_net64419), .A2(u5_mult_82_n6537), 
        .ZN(u5_mult_82_ab_8__8_) );
  NOR2_X2 u5_mult_82_U2508 ( .A1(u5_mult_82_net64435), .A2(u5_mult_82_n6610), 
        .ZN(u5_mult_82_ab_18__9_) );
  NOR2_X2 u5_mult_82_U2507 ( .A1(u5_mult_82_net64453), .A2(u5_mult_82_n6610), 
        .ZN(u5_mult_82_ab_18__10_) );
  INV_X2 u5_mult_82_U2506 ( .A(u5_mult_82_ab_24__10_), .ZN(u5_mult_82_n2416)
         );
  NOR2_X2 u5_mult_82_U2505 ( .A1(u5_mult_82_net64471), .A2(u5_mult_82_n6651), 
        .ZN(u5_mult_82_ab_26__11_) );
  NAND2_X2 u5_mult_82_U2504 ( .A1(u5_mult_82_ab_30__10_), .A2(
        u5_mult_82_SUMB_29__11_), .ZN(u5_mult_82_n3214) );
  NAND3_X2 u5_mult_82_U2503 ( .A1(u5_mult_82_n3213), .A2(u5_mult_82_n3214), 
        .A3(u5_mult_82_n3215), .ZN(u5_mult_82_CARRYB_30__10_) );
  NOR2_X1 u5_mult_82_U2502 ( .A1(u5_mult_82_net64433), .A2(u5_mult_82_n6716), 
        .ZN(u5_mult_82_ab_36__9_) );
  NOR2_X2 u5_mult_82_U2501 ( .A1(u5_mult_82_net64469), .A2(u5_mult_82_n6742), 
        .ZN(u5_mult_82_ab_46__11_) );
  NAND3_X2 u5_mult_82_U2500 ( .A1(u5_mult_82_n5676), .A2(u5_mult_82_n5677), 
        .A3(u5_mult_82_n5678), .ZN(u5_mult_82_CARRYB_45__12_) );
  NOR2_X1 u5_mult_82_U2499 ( .A1(u5_mult_82_net64559), .A2(u5_mult_82_n6741), 
        .ZN(u5_mult_82_ab_46__16_) );
  INV_X4 u5_mult_82_U2498 ( .A(u5_mult_82_ab_46__17_), .ZN(u5_mult_82_n4360)
         );
  NOR2_X1 u5_mult_82_U2497 ( .A1(u5_mult_82_n6891), .A2(u5_mult_82_n6741), 
        .ZN(u5_mult_82_ab_46__24_) );
  NOR2_X2 u5_mult_82_U2496 ( .A1(u5_mult_82_net64935), .A2(u5_mult_82_net65315), .ZN(u5_mult_82_ab_45__37_) );
  NOR2_X1 u5_mult_82_U2495 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_net65315), .ZN(u5_mult_82_ab_45__36_) );
  NOR2_X2 u5_mult_82_U2494 ( .A1(u5_mult_82_n6777), .A2(u5_mult_82_net65277), 
        .ZN(u5_mult_82_ab_47__48_) );
  NOR2_X1 u5_mult_82_U2493 ( .A1(u5_mult_82_n6784), .A2(u5_mult_82_net65277), 
        .ZN(u5_mult_82_ab_47__47_) );
  NOR2_X2 u5_mult_82_U2492 ( .A1(u5_mult_82_n6797), .A2(u5_mult_82_net65277), 
        .ZN(u5_mult_82_ab_47__45_) );
  NOR2_X1 u5_mult_82_U2491 ( .A1(u5_mult_82_n6983), .A2(u5_mult_82_n6737), 
        .ZN(u5_mult_82_ab_44__52_) );
  NOR2_X2 u5_mult_82_U2490 ( .A1(u5_mult_82_n6759), .A2(u5_mult_82_net65313), 
        .ZN(u5_mult_82_ab_45__51_) );
  NOR2_X2 u5_mult_82_U2489 ( .A1(u5_mult_82_n6837), .A2(u5_mult_82_n6734), 
        .ZN(u5_mult_82_ab_44__33_) );
  NOR2_X2 u5_mult_82_U2488 ( .A1(u5_mult_82_net64437), .A2(u5_mult_82_n6516), 
        .ZN(u5_mult_82_ab_3__9_) );
  NOR2_X2 u5_mult_82_U2487 ( .A1(u5_mult_82_net64437), .A2(u5_mult_82_n6537), 
        .ZN(u5_mult_82_ab_8__9_) );
  NOR2_X2 u5_mult_82_U2486 ( .A1(u5_mult_82_net64435), .A2(u5_mult_82_n6644), 
        .ZN(u5_mult_82_ab_24__9_) );
  NOR2_X2 u5_mult_82_U2485 ( .A1(u5_mult_82_net64453), .A2(u5_mult_82_net65679), .ZN(u5_mult_82_ab_25__10_) );
  NAND3_X2 u5_mult_82_U2484 ( .A1(u5_mult_82_n2284), .A2(u5_mult_82_n2285), 
        .A3(u5_mult_82_n2286), .ZN(u5_mult_82_CARRYB_25__12_) );
  INV_X4 u5_mult_82_U2483 ( .A(u5_mult_82_ab_30__10_), .ZN(u5_mult_82_n2676)
         );
  INV_X4 u5_mult_82_U2482 ( .A(u5_mult_82_ab_45__11_), .ZN(u5_mult_82_n5281)
         );
  NAND3_X2 u5_mult_82_U2481 ( .A1(u5_mult_82_n5461), .A2(u5_mult_82_n5462), 
        .A3(u5_mult_82_n5463), .ZN(u5_mult_82_CARRYB_45__13_) );
  NOR2_X1 u5_mult_82_U2480 ( .A1(u5_mult_82_n6933), .A2(u5_mult_82_n6736), 
        .ZN(u5_mult_82_ab_44__15_) );
  NOR2_X2 u5_mult_82_U2479 ( .A1(u5_mult_82_net64665), .A2(u5_mult_82_net65321), .ZN(u5_mult_82_ab_45__22_) );
  NOR2_X2 u5_mult_82_U2478 ( .A1(u5_mult_82_net64683), .A2(u5_mult_82_net65321), .ZN(u5_mult_82_ab_45__23_) );
  NOR2_X2 u5_mult_82_U2477 ( .A1(u5_mult_82_n6837), .A2(u5_mult_82_n6742), 
        .ZN(u5_mult_82_ab_46__33_) );
  NOR2_X2 u5_mult_82_U2476 ( .A1(u5_mult_82_net64881), .A2(u5_mult_82_n6734), 
        .ZN(u5_mult_82_ab_44__34_) );
  NOR2_X2 u5_mult_82_U2475 ( .A1(u5_mult_82_net64881), .A2(u5_mult_82_n6742), 
        .ZN(u5_mult_82_ab_46__34_) );
  NAND2_X2 u5_mult_82_U2474 ( .A1(u5_mult_82_ab_45__35_), .A2(
        u5_mult_82_CARRYB_44__35_), .ZN(u5_mult_82_n2653) );
  NOR2_X1 u5_mult_82_U2473 ( .A1(u5_mult_82_n6816), .A2(u5_mult_82_n6743), 
        .ZN(u5_mult_82_ab_46__42_) );
  NOR2_X1 u5_mult_82_U2472 ( .A1(u5_mult_82_net64455), .A2(u5_mult_82_n6516), 
        .ZN(u5_mult_82_ab_3__10_) );
  NOR2_X1 u5_mult_82_U2471 ( .A1(u5_mult_82_net64455), .A2(u5_mult_82_n6537), 
        .ZN(u5_mult_82_ab_8__10_) );
  NOR2_X2 u5_mult_82_U2470 ( .A1(u5_mult_82_net64473), .A2(u5_mult_82_n6567), 
        .ZN(u5_mult_82_ab_12__11_) );
  NOR2_X2 u5_mult_82_U2469 ( .A1(u5_mult_82_net64473), .A2(u5_mult_82_n6573), 
        .ZN(u5_mult_82_ab_13__11_) );
  NOR2_X2 u5_mult_82_U2468 ( .A1(u5_mult_82_net64471), .A2(u5_mult_82_n6610), 
        .ZN(u5_mult_82_ab_18__11_) );
  NOR2_X1 u5_mult_82_U2467 ( .A1(u5_mult_82_net64487), .A2(u5_mult_82_n6680), 
        .ZN(u5_mult_82_ab_30__12_) );
  NOR2_X2 u5_mult_82_U2466 ( .A1(u5_mult_82_net64453), .A2(u5_mult_82_net65409), .ZN(u5_mult_82_ab_40__10_) );
  INV_X2 u5_mult_82_U2465 ( .A(u5_mult_82_ab_43__10_), .ZN(u5_mult_82_net80099) );
  NOR2_X2 u5_mult_82_U2464 ( .A1(u5_mult_82_n6867), .A2(u5_mult_82_net65369), 
        .ZN(u5_mult_82_ab_42__28_) );
  NOR2_X2 u5_mult_82_U2463 ( .A1(u5_mult_82_n6821), .A2(u5_mult_82_net65385), 
        .ZN(u5_mult_82_ab_41__41_) );
  INV_X4 u5_mult_82_U2462 ( .A(u5_mult_82_ab_33__13_), .ZN(u5_mult_82_n3703)
         );
  NOR2_X2 u5_mult_82_U2461 ( .A1(u5_mult_82_net64473), .A2(u5_mult_82_n6516), 
        .ZN(u5_mult_82_ab_3__11_) );
  NOR2_X1 u5_mult_82_U2460 ( .A1(u5_mult_82_net64525), .A2(u5_mult_82_n6644), 
        .ZN(u5_mult_82_ab_24__14_) );
  NOR2_X1 u5_mult_82_U2459 ( .A1(u5_mult_82_n6934), .A2(u5_mult_82_n6644), 
        .ZN(u5_mult_82_ab_24__15_) );
  INV_X4 u5_mult_82_U2458 ( .A(u5_mult_82_ab_32__13_), .ZN(u5_mult_82_n3694)
         );
  NOR2_X1 u5_mult_82_U2457 ( .A1(u5_mult_82_net64487), .A2(u5_mult_82_net65373), .ZN(u5_mult_82_ab_42__12_) );
  NAND2_X2 u5_mult_82_U2456 ( .A1(u5_mult_82_ab_40__31_), .A2(
        u5_mult_82_SUMB_39__32_), .ZN(u5_mult_82_n3086) );
  NOR2_X2 u5_mult_82_U2455 ( .A1(u5_mult_82_n6832), .A2(u5_mult_82_net65387), 
        .ZN(u5_mult_82_ab_41__39_) );
  NOR2_X1 u5_mult_82_U2454 ( .A1(u5_mult_82_n6804), .A2(u5_mult_82_net65385), 
        .ZN(u5_mult_82_ab_41__44_) );
  NOR2_X2 u5_mult_82_U2453 ( .A1(u5_mult_82_net64491), .A2(u5_mult_82_n6516), 
        .ZN(u5_mult_82_ab_3__12_) );
  NOR2_X1 u5_mult_82_U2452 ( .A1(u5_mult_82_net64527), .A2(u5_mult_82_n6552), 
        .ZN(u5_mult_82_ab_10__14_) );
  NOR2_X2 u5_mult_82_U2451 ( .A1(u5_mult_82_net64525), .A2(u5_mult_82_n6596), 
        .ZN(u5_mult_82_ab_16__14_) );
  NOR2_X2 u5_mult_82_U2450 ( .A1(u5_mult_82_n6921), .A2(u5_mult_82_net65407), 
        .ZN(u5_mult_82_ab_40__18_) );
  NOR2_X2 u5_mult_82_U2449 ( .A1(u5_mult_82_net64669), .A2(u5_mult_82_net65407), .ZN(u5_mult_82_ab_40__22_) );
  NOR2_X2 u5_mult_82_U2448 ( .A1(u5_mult_82_n6880), .A2(u5_mult_82_net65443), 
        .ZN(u5_mult_82_ab_38__26_) );
  NOR2_X2 u5_mult_82_U2447 ( .A1(u5_mult_82_n6875), .A2(u5_mult_82_n6728), 
        .ZN(u5_mult_82_ab_39__27_) );
  NOR2_X1 u5_mult_82_U2446 ( .A1(u5_mult_82_n6827), .A2(u5_mult_82_n6729), 
        .ZN(u5_mult_82_ab_39__40_) );
  NAND3_X2 u5_mult_82_U2445 ( .A1(u5_mult_82_n957), .A2(u5_mult_82_n958), .A3(
        u5_mult_82_n959), .ZN(u5_mult_82_CARRYB_39__39_) );
  NOR2_X2 u5_mult_82_U2444 ( .A1(u5_mult_82_n6792), .A2(u5_mult_82_net65403), 
        .ZN(u5_mult_82_ab_40__46_) );
  NAND2_X2 u5_mult_82_U2443 ( .A1(u5_mult_82_n915), .A2(u5_mult_82_n916), .ZN(
        u5_mult_82_SUMB_39__36_) );
  NOR2_X1 u5_mult_82_U2442 ( .A1(u5_mult_82_net64509), .A2(u5_mult_82_net66021), .ZN(u5_mult_82_ab_6__13_) );
  NOR2_X2 u5_mult_82_U2441 ( .A1(u5_mult_82_net64525), .A2(u5_mult_82_n6616), 
        .ZN(u5_mult_82_ab_19__14_) );
  NOR2_X1 u5_mult_82_U2440 ( .A1(u5_mult_82_n6934), .A2(u5_mult_82_n6616), 
        .ZN(u5_mult_82_ab_19__15_) );
  NOR2_X2 u5_mult_82_U2439 ( .A1(u5_mult_82_n6928), .A2(u5_mult_82_n6615), 
        .ZN(u5_mult_82_ab_19__17_) );
  NOR2_X1 u5_mult_82_U2438 ( .A1(u5_mult_82_net64561), .A2(u5_mult_82_n6615), 
        .ZN(u5_mult_82_ab_19__16_) );
  NOR2_X1 u5_mult_82_U2437 ( .A1(u5_mult_82_n6921), .A2(u5_mult_82_n6615), 
        .ZN(u5_mult_82_ab_19__18_) );
  NAND2_X1 u5_mult_82_U2436 ( .A1(u5_mult_82_ab_37__13_), .A2(
        u5_mult_82_CARRYB_36__13_), .ZN(u5_mult_82_n4222) );
  NAND3_X2 u5_mult_82_U2435 ( .A1(u5_mult_82_net82055), .A2(
        u5_mult_82_net82056), .A3(u5_mult_82_n4222), .ZN(
        u5_mult_82_CARRYB_37__13_) );
  NAND2_X2 u5_mult_82_U2434 ( .A1(u5_mult_82_n1356), .A2(u5_mult_82_n6176), 
        .ZN(u5_mult_82_n1353) );
  NOR2_X2 u5_mult_82_U2433 ( .A1(u5_mult_82_n6885), .A2(u5_mult_82_net65443), 
        .ZN(u5_mult_82_ab_38__25_) );
  NOR2_X2 u5_mult_82_U2432 ( .A1(u5_mult_82_n6843), .A2(u5_mult_82_n6720), 
        .ZN(u5_mult_82_ab_37__32_) );
  NOR2_X2 u5_mult_82_U2431 ( .A1(u5_mult_82_n6785), .A2(u5_mult_82_net65403), 
        .ZN(u5_mult_82_ab_40__47_) );
  NOR2_X2 u5_mult_82_U2430 ( .A1(u5_mult_82_n6766), .A2(u5_mult_82_n1321), 
        .ZN(u5_mult_82_ab_42__50_) );
  NOR2_X2 u5_mult_82_U2429 ( .A1(u5_mult_82_n6772), .A2(u5_mult_82_n1321), 
        .ZN(u5_mult_82_ab_42__49_) );
  NOR2_X2 u5_mult_82_U2428 ( .A1(u5_mult_82_n6777), .A2(u5_mult_82_n1321), 
        .ZN(u5_mult_82_ab_42__48_) );
  NAND2_X2 u5_mult_82_U2427 ( .A1(u5_mult_82_ab_36__35_), .A2(
        u5_mult_82_SUMB_35__36_), .ZN(u5_mult_82_n5085) );
  INV_X4 u5_mult_82_U2426 ( .A(u5_mult_82_n6632), .ZN(u5_mult_82_n6629) );
  INV_X4 u5_mult_82_U2425 ( .A(u5_mult_82_ab_25__16_), .ZN(u5_mult_82_n1798)
         );
  INV_X4 u5_mult_82_U2424 ( .A(u5_mult_82_n1497), .ZN(u5_mult_82_n1498) );
  NOR2_X1 u5_mult_82_U2423 ( .A1(u5_mult_82_n6933), .A2(u5_mult_82_n6695), 
        .ZN(u5_mult_82_ab_32__15_) );
  INV_X4 u5_mult_82_U2422 ( .A(u5_mult_82_ab_36__15_), .ZN(u5_mult_82_net83710) );
  NOR2_X2 u5_mult_82_U2421 ( .A1(u5_mult_82_n6927), .A2(u5_mult_82_n6708), 
        .ZN(u5_mult_82_ab_35__17_) );
  INV_X8 u5_mult_82_U2420 ( .A(u5_mult_82_n7018), .ZN(u5_mult_82_n6888) );
  NOR2_X1 u5_mult_82_U2419 ( .A1(u5_mult_82_n6791), .A2(u5_mult_82_n6713), 
        .ZN(u5_mult_82_ab_36__46_) );
  NOR2_X2 u5_mult_82_U2418 ( .A1(u5_mult_82_net64937), .A2(u5_mult_82_n6707), 
        .ZN(u5_mult_82_ab_35__37_) );
  NOR2_X1 u5_mult_82_U2417 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6707), 
        .ZN(u5_mult_82_ab_35__38_) );
  NOR2_X1 u5_mult_82_U2416 ( .A1(u5_mult_82_n6832), .A2(u5_mult_82_n6707), 
        .ZN(u5_mult_82_ab_35__39_) );
  NOR2_X2 u5_mult_82_U2415 ( .A1(u5_mult_82_n6935), .A2(u5_mult_82_net66039), 
        .ZN(u5_mult_82_ab_5__15_) );
  NOR2_X2 u5_mult_82_U2414 ( .A1(u5_mult_82_net64563), .A2(u5_mult_82_net66037), .ZN(u5_mult_82_ab_5__16_) );
  NOR2_X2 u5_mult_82_U2413 ( .A1(u5_mult_82_n6929), .A2(u5_mult_82_net66037), 
        .ZN(u5_mult_82_ab_5__17_) );
  NOR2_X2 u5_mult_82_U2412 ( .A1(u5_mult_82_net64563), .A2(u5_mult_82_n6587), 
        .ZN(u5_mult_82_ab_15__16_) );
  INV_X4 u5_mult_82_U2411 ( .A(u5_mult_82_n1650), .ZN(u5_mult_82_n1651) );
  NOR2_X2 u5_mult_82_U2410 ( .A1(u5_mult_82_n6891), .A2(u5_mult_82_n6708), 
        .ZN(u5_mult_82_ab_35__24_) );
  NOR2_X2 u5_mult_82_U2409 ( .A1(u5_mult_82_n6875), .A2(u5_mult_82_net65515), 
        .ZN(u5_mult_82_ab_34__27_) );
  NOR2_X2 u5_mult_82_U2408 ( .A1(u5_mult_82_n6857), .A2(u5_mult_82_n6714), 
        .ZN(u5_mult_82_ab_36__30_) );
  NAND3_X2 u5_mult_82_U2407 ( .A1(u5_mult_82_n3764), .A2(u5_mult_82_n3765), 
        .A3(u5_mult_82_n3766), .ZN(u5_mult_82_CARRYB_34__40_) );
  NOR2_X2 u5_mult_82_U2406 ( .A1(u5_mult_82_n6827), .A2(u5_mult_82_n6706), 
        .ZN(u5_mult_82_ab_35__40_) );
  NOR2_X1 u5_mult_82_U2405 ( .A1(u5_mult_82_n6797), .A2(u5_mult_82_n6713), 
        .ZN(u5_mult_82_ab_36__45_) );
  NOR2_X2 u5_mult_82_U2404 ( .A1(u5_mult_82_n6778), .A2(u5_mult_82_n6706), 
        .ZN(u5_mult_82_ab_35__48_) );
  NOR2_X1 u5_mult_82_U2403 ( .A1(u5_mult_82_n6804), .A2(u5_mult_82_n6706), 
        .ZN(u5_mult_82_ab_35__44_) );
  NOR2_X2 u5_mult_82_U2402 ( .A1(u5_mult_82_n6922), .A2(u5_mult_82_net66037), 
        .ZN(u5_mult_82_ab_5__18_) );
  INV_X4 u5_mult_82_U2401 ( .A(u5_mult_82_n6561), .ZN(u5_mult_82_n6558) );
  NOR2_X2 u5_mult_82_U2400 ( .A1(u5_mult_82_n6906), .A2(u5_mult_82_n6536), 
        .ZN(u5_mult_82_ab_8__20_) );
  NOR2_X2 u5_mult_82_U2399 ( .A1(u5_mult_82_net64667), .A2(u5_mult_82_n6708), 
        .ZN(u5_mult_82_ab_35__22_) );
  INV_X4 u5_mult_82_U2398 ( .A(u5_mult_82_ab_35__23_), .ZN(u5_mult_82_n2325)
         );
  NOR2_X2 u5_mult_82_U2397 ( .A1(u5_mult_82_n6868), .A2(u5_mult_82_net65513), 
        .ZN(u5_mult_82_ab_34__28_) );
  NOR2_X2 u5_mult_82_U2396 ( .A1(u5_mult_82_n6773), .A2(u5_mult_82_n6706), 
        .ZN(u5_mult_82_ab_35__49_) );
  NOR2_X1 u5_mult_82_U2395 ( .A1(u5_mult_82_n6982), .A2(u5_mult_82_n6717), 
        .ZN(u5_mult_82_ab_36__52_) );
  NOR2_X2 u5_mult_82_U2394 ( .A1(u5_mult_82_n6760), .A2(u5_mult_82_n6719), 
        .ZN(u5_mult_82_ab_37__51_) );
  NOR2_X1 u5_mult_82_U2393 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6684), 
        .ZN(u5_mult_82_ab_31__38_) );
  NOR2_X2 u5_mult_82_U2392 ( .A1(u5_mult_82_net64671), .A2(u5_mult_82_n6587), 
        .ZN(u5_mult_82_ab_15__22_) );
  NOR2_X2 u5_mult_82_U2391 ( .A1(u5_mult_82_n6921), .A2(u5_mult_82_net65677), 
        .ZN(u5_mult_82_ab_25__18_) );
  INV_X4 u5_mult_82_U2390 ( .A(u5_mult_82_ab_25__20_), .ZN(u5_mult_82_n3283)
         );
  NOR2_X2 u5_mult_82_U2389 ( .A1(u5_mult_82_n6904), .A2(u5_mult_82_n6685), 
        .ZN(u5_mult_82_ab_31__20_) );
  NOR2_X2 u5_mult_82_U2388 ( .A1(u5_mult_82_n6920), .A2(u5_mult_82_n6708), 
        .ZN(u5_mult_82_ab_35__18_) );
  INV_X4 u5_mult_82_U2387 ( .A(u5_mult_82_ab_35__20_), .ZN(u5_mult_82_n5512)
         );
  NAND3_X2 u5_mult_82_U2386 ( .A1(u5_mult_82_n5870), .A2(u5_mult_82_n5869), 
        .A3(u5_mult_82_n5868), .ZN(u5_mult_82_CARRYB_32__31_) );
  NOR2_X2 u5_mult_82_U2385 ( .A1(u5_mult_82_n6811), .A2(u5_mult_82_n6685), 
        .ZN(u5_mult_82_ab_31__43_) );
  NOR2_X2 u5_mult_82_U2384 ( .A1(u5_mult_82_n6767), .A2(u5_mult_82_n6706), 
        .ZN(u5_mult_82_ab_35__50_) );
  NOR2_X2 u5_mult_82_U2383 ( .A1(u5_mult_82_n6827), .A2(u5_mult_82_n6686), 
        .ZN(u5_mult_82_ab_31__40_) );
  NOR2_X2 u5_mult_82_U2382 ( .A1(u5_mult_82_n6821), .A2(u5_mult_82_n6685), 
        .ZN(u5_mult_82_ab_31__41_) );
  NOR2_X2 u5_mult_82_U2381 ( .A1(u5_mult_82_n6832), .A2(u5_mult_82_n6684), 
        .ZN(u5_mult_82_ab_31__39_) );
  NOR2_X1 u5_mult_82_U2380 ( .A1(u5_mult_82_n6893), .A2(u5_mult_82_n6579), 
        .ZN(u5_mult_82_ab_14__24_) );
  INV_X4 u5_mult_82_U2379 ( .A(u5_mult_82_ab_30__19_), .ZN(u5_mult_82_net80364) );
  NOR2_X2 u5_mult_82_U2378 ( .A1(u5_mult_82_n6880), .A2(u5_mult_82_n6685), 
        .ZN(u5_mult_82_ab_31__26_) );
  NOR2_X2 u5_mult_82_U2377 ( .A1(u5_mult_82_net64901), .A2(u5_mult_82_n6684), 
        .ZN(u5_mult_82_ab_31__35_) );
  NOR2_X1 u5_mult_82_U2376 ( .A1(u5_mult_82_n6982), .A2(u5_mult_82_n6681), 
        .ZN(u5_mult_82_ab_30__52_) );
  NOR2_X2 u5_mult_82_U2375 ( .A1(u5_mult_82_n6760), .A2(u5_mult_82_n6683), 
        .ZN(u5_mult_82_ab_31__51_) );
  INV_X8 u5_mult_82_U2374 ( .A(u5_mult_82_n6908), .ZN(u5_mult_82_n6907) );
  NAND3_X2 u5_mult_82_U2373 ( .A1(u5_mult_82_n1168), .A2(u5_mult_82_n1169), 
        .A3(u5_mult_82_n1170), .ZN(u5_mult_82_CARRYB_4__22_) );
  NAND3_X2 u5_mult_82_U2372 ( .A1(u5_mult_82_n5231), .A2(u5_mult_82_n5232), 
        .A3(u5_mult_82_n5233), .ZN(u5_mult_82_CARRYB_20__20_) );
  NOR2_X1 u5_mult_82_U2371 ( .A1(u5_mult_82_n6891), .A2(u5_mult_82_n6685), 
        .ZN(u5_mult_82_ab_31__24_) );
  INV_X4 u5_mult_82_U2370 ( .A(u5_mult_82_ab_29__30_), .ZN(u5_mult_82_n1746)
         );
  NOR2_X2 u5_mult_82_U2369 ( .A1(u5_mult_82_net64883), .A2(u5_mult_82_n6678), 
        .ZN(u5_mult_82_ab_30__34_) );
  NOR2_X2 u5_mult_82_U2368 ( .A1(u5_mult_82_n6838), .A2(u5_mult_82_n6678), 
        .ZN(u5_mult_82_ab_30__33_) );
  NOR2_X1 u5_mult_82_U2367 ( .A1(u5_mult_82_n6791), .A2(u5_mult_82_n6670), 
        .ZN(u5_mult_82_ab_29__46_) );
  NOR2_X2 u5_mult_82_U2366 ( .A1(u5_mult_82_n6778), .A2(u5_mult_82_n6677), 
        .ZN(u5_mult_82_ab_30__48_) );
  NOR2_X2 u5_mult_82_U2365 ( .A1(u5_mult_82_n6832), .A2(u5_mult_82_n6663), 
        .ZN(u5_mult_82_ab_28__39_) );
  NOR2_X1 u5_mult_82_U2364 ( .A1(u5_mult_82_n6832), .A2(u5_mult_82_n6656), 
        .ZN(u5_mult_82_ab_27__39_) );
  NOR2_X2 u5_mult_82_U2363 ( .A1(u5_mult_82_n6817), .A2(u5_mult_82_n6655), 
        .ZN(u5_mult_82_ab_27__42_) );
  NOR2_X2 u5_mult_82_U2362 ( .A1(u5_mult_82_n6893), .A2(u5_mult_82_n6522), 
        .ZN(u5_mult_82_ab_4__24_) );
  NOR2_X2 u5_mult_82_U2361 ( .A1(u5_mult_82_net64689), .A2(u5_mult_82_n6551), 
        .ZN(u5_mult_82_ab_10__23_) );
  NOR2_X2 u5_mult_82_U2360 ( .A1(u5_mult_82_net64671), .A2(u5_mult_82_n6551), 
        .ZN(u5_mult_82_ab_10__22_) );
  NOR2_X2 u5_mult_82_U2359 ( .A1(u5_mult_82_n6892), .A2(u5_mult_82_n6609), 
        .ZN(u5_mult_82_ab_18__24_) );
  NOR2_X2 u5_mult_82_U2358 ( .A1(u5_mult_82_net64669), .A2(u5_mult_82_n6650), 
        .ZN(u5_mult_82_ab_26__22_) );
  INV_X4 u5_mult_82_U2357 ( .A(u5_mult_82_ab_28__30_), .ZN(u5_mult_82_n2414)
         );
  NOR2_X2 u5_mult_82_U2356 ( .A1(u5_mult_82_n6773), .A2(u5_mult_82_n6677), 
        .ZN(u5_mult_82_ab_30__49_) );
  NOR2_X2 u5_mult_82_U2355 ( .A1(u5_mult_82_n6767), .A2(u5_mult_82_n6677), 
        .ZN(u5_mult_82_ab_30__50_) );
  NOR2_X2 u5_mult_82_U2354 ( .A1(u5_mult_82_n6822), .A2(u5_mult_82_n6651), 
        .ZN(u5_mult_82_ab_26__41_) );
  NOR2_X1 u5_mult_82_U2353 ( .A1(u5_mult_82_n6805), .A2(u5_mult_82_n6651), 
        .ZN(u5_mult_82_ab_26__44_) );
  NOR2_X2 u5_mult_82_U2352 ( .A1(u5_mult_82_n6887), .A2(u5_mult_82_n6545), 
        .ZN(u5_mult_82_ab_9__25_) );
  NOR2_X2 u5_mult_82_U2351 ( .A1(u5_mult_82_n6877), .A2(u5_mult_82_n6545), 
        .ZN(u5_mult_82_ab_9__27_) );
  NOR2_X2 u5_mult_82_U2350 ( .A1(u5_mult_82_n6887), .A2(u5_mult_82_n6579), 
        .ZN(u5_mult_82_ab_14__25_) );
  NOR2_X2 u5_mult_82_U2349 ( .A1(u5_mult_82_net64687), .A2(u5_mult_82_n6650), 
        .ZN(u5_mult_82_ab_26__23_) );
  INV_X4 u5_mult_82_U2348 ( .A(u5_mult_82_ab_24__26_), .ZN(u5_mult_82_n2175)
         );
  INV_X4 u5_mult_82_U2347 ( .A(u5_mult_82_n1414), .ZN(u5_mult_82_n1415) );
  NOR2_X1 u5_mult_82_U2346 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_net65675), .ZN(u5_mult_82_ab_25__38_) );
  NOR2_X1 u5_mult_82_U2345 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6649), 
        .ZN(u5_mult_82_ab_26__36_) );
  NOR2_X2 u5_mult_82_U2344 ( .A1(u5_mult_82_n6886), .A2(u5_mult_82_net65677), 
        .ZN(u5_mult_82_ab_25__25_) );
  NOR2_X1 u5_mult_82_U2343 ( .A1(u5_mult_82_n6876), .A2(u5_mult_82_net65677), 
        .ZN(u5_mult_82_ab_25__27_) );
  INV_X4 u5_mult_82_U2342 ( .A(u5_mult_82_ab_25__29_), .ZN(u5_mult_82_n3710)
         );
  NAND3_X2 u5_mult_82_U2341 ( .A1(u5_mult_82_n3593), .A2(u5_mult_82_n3594), 
        .A3(u5_mult_82_n3595), .ZN(u5_mult_82_CARRYB_25__46_) );
  NOR2_X1 u5_mult_82_U2340 ( .A1(u5_mult_82_n6877), .A2(u5_mult_82_n6572), 
        .ZN(u5_mult_82_ab_13__27_) );
  NOR2_X1 u5_mult_82_U2339 ( .A1(u5_mult_82_n6839), .A2(u5_mult_82_net65711), 
        .ZN(u5_mult_82_ab_23__33_) );
  NOR2_X2 u5_mult_82_U2338 ( .A1(u5_mult_82_n6768), .A2(u5_mult_82_n1381), 
        .ZN(u5_mult_82_ab_25__50_) );
  NOR2_X2 u5_mult_82_U2337 ( .A1(u5_mult_82_n6774), .A2(u5_mult_82_n6642), 
        .ZN(u5_mult_82_ab_24__49_) );
  NOR2_X2 u5_mult_82_U2336 ( .A1(u5_mult_82_n6785), .A2(u5_mult_82_net65681), 
        .ZN(u5_mult_82_ab_25__47_) );
  NOR2_X2 u5_mult_82_U2335 ( .A1(u5_mult_82_n6761), .A2(u5_mult_82_n1381), 
        .ZN(u5_mult_82_ab_25__51_) );
  NOR2_X1 u5_mult_82_U2334 ( .A1(u5_mult_82_n6822), .A2(u5_mult_82_n6636), 
        .ZN(u5_mult_82_ab_22__41_) );
  NOR2_X2 u5_mult_82_U2333 ( .A1(u5_mult_82_n6817), .A2(u5_mult_82_n6636), 
        .ZN(u5_mult_82_ab_22__42_) );
  NOR2_X1 u5_mult_82_U2332 ( .A1(u5_mult_82_n6798), .A2(u5_mult_82_n6636), 
        .ZN(u5_mult_82_ab_22__45_) );
  NOR2_X1 u5_mult_82_U2331 ( .A1(u5_mult_82_n6812), .A2(u5_mult_82_n6636), 
        .ZN(u5_mult_82_ab_22__43_) );
  INV_X4 u5_mult_82_U2330 ( .A(u5_mult_82_ab_22__44_), .ZN(u5_mult_82_n1102)
         );
  NOR2_X2 u5_mult_82_U2329 ( .A1(u5_mult_82_n6828), .A2(u5_mult_82_n6644), 
        .ZN(u5_mult_82_ab_24__40_) );
  NOR2_X1 u5_mult_82_U2328 ( .A1(u5_mult_82_n6785), .A2(u5_mult_82_n6630), 
        .ZN(u5_mult_82_ab_21__47_) );
  NAND3_X2 u5_mult_82_U2327 ( .A1(u5_mult_82_n2928), .A2(u5_mult_82_n2929), 
        .A3(u5_mult_82_n2930), .ZN(u5_mult_82_CARRYB_21__46_) );
  NOR2_X2 u5_mult_82_U2326 ( .A1(u5_mult_82_n6881), .A2(u5_mult_82_n6609), 
        .ZN(u5_mult_82_ab_18__26_) );
  NOR2_X2 u5_mult_82_U2325 ( .A1(u5_mult_82_n6882), .A2(u5_mult_82_net66037), 
        .ZN(u5_mult_82_ab_5__26_) );
  INV_X4 u5_mult_82_U2324 ( .A(u5_mult_82_ab_5__28_), .ZN(u5_mult_82_n3665) );
  NAND3_X2 u5_mult_82_U2323 ( .A1(u5_mult_82_n3464), .A2(u5_mult_82_n3465), 
        .A3(u5_mult_82_n3466), .ZN(u5_mult_82_CARRYB_6__30_) );
  NOR2_X1 u5_mult_82_U2322 ( .A1(u5_mult_82_n6870), .A2(u5_mult_82_n6571), 
        .ZN(u5_mult_82_ab_13__28_) );
  INV_X4 u5_mult_82_U2321 ( .A(u5_mult_82_n1817), .ZN(u5_mult_82_n1818) );
  NOR2_X1 u5_mult_82_U2320 ( .A1(u5_mult_82_n6864), .A2(u5_mult_82_n6571), 
        .ZN(u5_mult_82_ab_13__29_) );
  NOR2_X1 u5_mult_82_U2319 ( .A1(u5_mult_82_n6869), .A2(u5_mult_82_n6621), 
        .ZN(u5_mult_82_ab_20__28_) );
  NOR2_X1 u5_mult_82_U2318 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6635), 
        .ZN(u5_mult_82_ab_22__36_) );
  NOR2_X2 u5_mult_82_U2317 ( .A1(u5_mult_82_n6831), .A2(u5_mult_82_n6635), 
        .ZN(u5_mult_82_ab_22__39_) );
  NOR2_X2 u5_mult_82_U2316 ( .A1(u5_mult_82_n6768), .A2(u5_mult_82_n6613), 
        .ZN(u5_mult_82_ab_19__50_) );
  NOR2_X2 u5_mult_82_U2315 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6635), 
        .ZN(u5_mult_82_ab_22__38_) );
  INV_X4 u5_mult_82_U2314 ( .A(u5_mult_82_ab_15__30_), .ZN(u5_mult_82_n838) );
  NOR2_X2 u5_mult_82_U2313 ( .A1(u5_mult_82_n6845), .A2(u5_mult_82_net66035), 
        .ZN(u5_mult_82_ab_5__32_) );
  NOR2_X2 u5_mult_82_U2312 ( .A1(u5_mult_82_n6840), .A2(u5_mult_82_net66035), 
        .ZN(u5_mult_82_ab_5__33_) );
  INV_X4 u5_mult_82_U2311 ( .A(u5_mult_82_n6854), .ZN(u5_mult_82_n6853) );
  NOR2_X2 u5_mult_82_U2310 ( .A1(u5_mult_82_net64217), .A2(u5_mult_82_n6842), 
        .ZN(u5_mult_82_ab_0__32_) );
  NOR2_X1 u5_mult_82_U2309 ( .A1(u5_mult_82_n6851), .A2(u5_mult_82_n6614), 
        .ZN(u5_mult_82_ab_19__31_) );
  NOR2_X1 u5_mult_82_U2308 ( .A1(u5_mult_82_net64885), .A2(u5_mult_82_n6614), 
        .ZN(u5_mult_82_ab_19__34_) );
  NOR2_X1 u5_mult_82_U2307 ( .A1(u5_mult_82_n6831), .A2(u5_mult_82_n6621), 
        .ZN(u5_mult_82_ab_20__39_) );
  NOR2_X2 u5_mult_82_U2306 ( .A1(u5_mult_82_n6761), .A2(u5_mult_82_n6613), 
        .ZN(u5_mult_82_ab_19__51_) );
  NOR2_X2 u5_mult_82_U2305 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6628), 
        .ZN(u5_mult_82_ab_21__38_) );
  NOR2_X2 u5_mult_82_U2304 ( .A1(u5_mult_82_n6845), .A2(u5_mult_82_n6578), 
        .ZN(u5_mult_82_ab_14__32_) );
  NAND3_X2 u5_mult_82_U2303 ( .A1(u5_mult_82_n3535), .A2(u5_mult_82_n3534), 
        .A3(u5_mult_82_n3533), .ZN(u5_mult_82_CARRYB_19__33_) );
  NOR2_X2 u5_mult_82_U2302 ( .A1(u5_mult_82_n6817), .A2(u5_mult_82_n6607), 
        .ZN(u5_mult_82_ab_18__42_) );
  NOR2_X2 u5_mult_82_U2301 ( .A1(u5_mult_82_n6792), .A2(u5_mult_82_n6600), 
        .ZN(u5_mult_82_ab_17__46_) );
  NOR2_X2 u5_mult_82_U2300 ( .A1(u5_mult_82_n6798), .A2(u5_mult_82_n6600), 
        .ZN(u5_mult_82_ab_17__45_) );
  NOR2_X2 u5_mult_82_U2299 ( .A1(u5_mult_82_n6779), .A2(u5_mult_82_n6593), 
        .ZN(u5_mult_82_ab_16__48_) );
  NOR2_X2 u5_mult_82_U2298 ( .A1(u5_mult_82_net64887), .A2(u5_mult_82_net66017), .ZN(u5_mult_82_ab_6__34_) );
  NOR2_X2 u5_mult_82_U2297 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6614), 
        .ZN(u5_mult_82_ab_19__38_) );
  NOR2_X1 u5_mult_82_U2296 ( .A1(u5_mult_82_n6831), .A2(u5_mult_82_n6594), 
        .ZN(u5_mult_82_ab_16__39_) );
  NOR2_X2 u5_mult_82_U2295 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6608), 
        .ZN(u5_mult_82_ab_18__38_) );
  NOR2_X2 u5_mult_82_U2294 ( .A1(u5_mult_82_n6840), .A2(u5_mult_82_n6578), 
        .ZN(u5_mult_82_ab_14__33_) );
  NOR2_X2 u5_mult_82_U2293 ( .A1(u5_mult_82_n6823), .A2(u5_mult_82_n6585), 
        .ZN(u5_mult_82_ab_15__41_) );
  NOR2_X2 u5_mult_82_U2292 ( .A1(u5_mult_82_net64905), .A2(u5_mult_82_net66017), .ZN(u5_mult_82_ab_6__35_) );
  NOR2_X2 u5_mult_82_U2291 ( .A1(u5_mult_82_net64905), .A2(u5_mult_82_n6578), 
        .ZN(u5_mult_82_ab_14__35_) );
  INV_X4 u5_mult_82_U2290 ( .A(u5_mult_82_ab_13__46_), .ZN(u5_mult_82_n3152)
         );
  NOR2_X2 u5_mult_82_U2289 ( .A1(u5_mult_82_n6786), .A2(u5_mult_82_n6580), 
        .ZN(u5_mult_82_ab_14__47_) );
  NOR2_X1 u5_mult_82_U2288 ( .A1(u5_mult_82_n6786), .A2(u5_mult_82_n6573), 
        .ZN(u5_mult_82_ab_13__47_) );
  INV_X4 u5_mult_82_U2287 ( .A(u5_mult_82_ab_13__38_), .ZN(u5_mult_82_n2415)
         );
  NOR2_X2 u5_mult_82_U2286 ( .A1(u5_mult_82_net64959), .A2(u5_mult_82_n6535), 
        .ZN(u5_mult_82_ab_8__38_) );
  NOR2_X1 u5_mult_82_U2285 ( .A1(u5_mult_82_net64941), .A2(u5_mult_82_n6535), 
        .ZN(u5_mult_82_ab_8__37_) );
  NOR2_X1 u5_mult_82_U2284 ( .A1(u5_mult_82_n6833), .A2(u5_mult_82_n6557), 
        .ZN(u5_mult_82_ab_11__39_) );
  INV_X4 u5_mult_82_U2283 ( .A(u5_mult_82_ab_11__43_), .ZN(u5_mult_82_n5272)
         );
  NAND3_X2 u5_mult_82_U2282 ( .A1(u5_mult_82_n4741), .A2(u5_mult_82_n4742), 
        .A3(u5_mult_82_n4743), .ZN(u5_mult_82_CARRYB_6__39_) );
  NOR2_X2 u5_mult_82_U2281 ( .A1(u5_mult_82_net64959), .A2(u5_mult_82_n6521), 
        .ZN(u5_mult_82_ab_4__38_) );
  NAND3_X2 u5_mult_82_U2280 ( .A1(u5_mult_82_n3399), .A2(u5_mult_82_n3400), 
        .A3(u5_mult_82_n3401), .ZN(u5_mult_82_CARRYB_11__40_) );
  NOR2_X2 u5_mult_82_U2279 ( .A1(u5_mult_82_n6769), .A2(u5_mult_82_n6543), 
        .ZN(u5_mult_82_ab_9__50_) );
  NOR2_X1 u5_mult_82_U2278 ( .A1(u5_mult_82_n6793), .A2(u5_mult_82_n6559), 
        .ZN(u5_mult_82_ab_11__46_) );
  NOR2_X1 u5_mult_82_U2277 ( .A1(u5_mult_82_n6829), .A2(u5_mult_82_net66019), 
        .ZN(u5_mult_82_ab_6__40_) );
  NOR2_X2 u5_mult_82_U2276 ( .A1(u5_mult_82_net64959), .A2(u5_mult_82_net66035), .ZN(u5_mult_82_ab_5__38_) );
  NOR2_X2 u5_mult_82_U2275 ( .A1(u5_mult_82_n6775), .A2(u5_mult_82_net66017), 
        .ZN(u5_mult_82_ab_6__49_) );
  NOR2_X2 u5_mult_82_U2274 ( .A1(u5_mult_82_n6786), .A2(u5_mult_82_n6530), 
        .ZN(u5_mult_82_ab_7__47_) );
  NOR2_X2 u5_mult_82_U2273 ( .A1(u5_mult_82_n6799), .A2(u5_mult_82_n6530), 
        .ZN(u5_mult_82_ab_7__45_) );
  INV_X4 u5_mult_82_U2272 ( .A(u5_mult_82_ab_7__44_), .ZN(u5_mult_82_n2556) );
  NAND2_X2 u5_mult_82_U2271 ( .A1(u5_mult_82_ab_7__41_), .A2(
        u5_mult_82_SUMB_6__42_), .ZN(u5_mult_82_n6019) );
  INV_X4 u5_mult_82_U2270 ( .A(u5_mult_82_n6510), .ZN(u5_mult_82_CARRYB_1__50_) );
  INV_X4 u5_mult_82_U2269 ( .A(u5_mult_82_n6505), .ZN(u5_mult_82_SUMB_1__47_)
         );
  INV_X4 u5_mult_82_U2268 ( .A(u5_mult_82_n6503), .ZN(u5_mult_82_SUMB_1__46_)
         );
  NAND2_X2 u5_mult_82_U2267 ( .A1(u5_mult_82_ab_1__49_), .A2(
        u5_mult_82_ab_0__50_), .ZN(u5_mult_82_n6508) );
  NOR2_X2 u5_mult_82_U2266 ( .A1(u5_mult_82_n6989), .A2(u5_mult_82_n6524), 
        .ZN(u5_mult_82_ab_4__0_) );
  NOR2_X2 u5_mult_82_U2265 ( .A1(u5_mult_82_n6989), .A2(u5_mult_82_n6547), 
        .ZN(u5_mult_82_ab_9__0_) );
  NOR2_X2 u5_mult_82_U2264 ( .A1(u5_mult_82_n6989), .A2(u5_mult_82_n6581), 
        .ZN(u5_mult_82_ab_14__0_) );
  NOR2_X2 u5_mult_82_U2263 ( .A1(u5_mult_82_n6988), .A2(u5_mult_82_n6617), 
        .ZN(u5_mult_82_ab_19__0_) );
  NOR2_X2 u5_mult_82_U2262 ( .A1(u5_mult_82_n6988), .A2(u5_mult_82_n6645), 
        .ZN(u5_mult_82_ab_24__0_) );
  NOR2_X2 u5_mult_82_U2261 ( .A1(u5_mult_82_n6987), .A2(u5_mult_82_n6674), 
        .ZN(u5_mult_82_ab_29__0_) );
  NOR2_X2 u5_mult_82_U2260 ( .A1(u5_mult_82_n6987), .A2(u5_mult_82_net65519), 
        .ZN(u5_mult_82_ab_34__0_) );
  NOR2_X1 u5_mult_82_U2259 ( .A1(u5_mult_82_n6986), .A2(u5_mult_82_n6974), 
        .ZN(u5_mult_82_ab_52__0_) );
  NOR2_X1 u5_mult_82_U2258 ( .A1(u5_mult_82_n6986), .A2(u5_mult_82_n6743), 
        .ZN(u5_mult_82_ab_46__0_) );
  NAND3_X2 u5_mult_82_U2257 ( .A1(u5_mult_82_net79210), .A2(u5_mult_82_n6036), 
        .A3(u5_mult_82_net79212), .ZN(u5_mult_82_CARRYB_29__20_) );
  NOR2_X2 u5_mult_82_U2256 ( .A1(u5_mult_82_n6913), .A2(u5_mult_82_n6672), 
        .ZN(u5_mult_82_ab_29__19_) );
  NOR2_X1 u5_mult_82_U2255 ( .A1(u5_mult_82_net64223), .A2(u5_mult_82_n6970), 
        .ZN(u5_mult_82_ab_0__1_) );
  NOR2_X2 u5_mult_82_U2254 ( .A1(u5_mult_82_n6969), .A2(u5_mult_82_n6524), 
        .ZN(u5_mult_82_ab_4__1_) );
  INV_X16 u5_mult_82_U2253 ( .A(u5_mult_82_net66025), .ZN(u5_mult_82_net66023)
         );
  NOR2_X2 u5_mult_82_U2252 ( .A1(u5_mult_82_n6969), .A2(u5_mult_82_n6547), 
        .ZN(u5_mult_82_ab_9__1_) );
  INV_X16 u5_mult_82_U2251 ( .A(u5_mult_82_n6561), .ZN(u5_mult_82_n6560) );
  NOR2_X2 u5_mult_82_U2250 ( .A1(u5_mult_82_n6969), .A2(u5_mult_82_n6581), 
        .ZN(u5_mult_82_ab_14__1_) );
  NOR2_X2 u5_mult_82_U2249 ( .A1(u5_mult_82_n6968), .A2(u5_mult_82_n6617), 
        .ZN(u5_mult_82_ab_19__1_) );
  INV_X16 u5_mult_82_U2248 ( .A(u5_mult_82_n6632), .ZN(u5_mult_82_n6631) );
  NOR2_X2 u5_mult_82_U2247 ( .A1(u5_mult_82_n6967), .A2(u5_mult_82_n6674), 
        .ZN(u5_mult_82_ab_29__1_) );
  NOR2_X1 u5_mult_82_U2246 ( .A1(u5_mult_82_n6967), .A2(u5_mult_82_net65519), 
        .ZN(u5_mult_82_ab_34__1_) );
  INV_X4 u5_mult_82_U2245 ( .A(u5_mult_82_ab_48__1_), .ZN(u5_mult_82_n4080) );
  NOR2_X2 u5_mult_82_U2244 ( .A1(u5_mult_82_net64223), .A2(u5_mult_82_n6959), 
        .ZN(u5_mult_82_ab_0__2_) );
  NOR2_X2 u5_mult_82_U2243 ( .A1(u5_mult_82_n6962), .A2(u5_mult_82_n6524), 
        .ZN(u5_mult_82_ab_4__2_) );
  INV_X8 u5_mult_82_U2242 ( .A(u5_mult_82_n6527), .ZN(u5_mult_82_n6532) );
  NOR2_X2 u5_mult_82_U2241 ( .A1(u5_mult_82_n6962), .A2(u5_mult_82_n6547), 
        .ZN(u5_mult_82_ab_9__2_) );
  NOR2_X2 u5_mult_82_U2240 ( .A1(u5_mult_82_n6962), .A2(u5_mult_82_n6581), 
        .ZN(u5_mult_82_ab_14__2_) );
  NOR2_X2 u5_mult_82_U2239 ( .A1(u5_mult_82_n6961), .A2(u5_mult_82_n6617), 
        .ZN(u5_mult_82_ab_19__2_) );
  INV_X8 u5_mult_82_U2238 ( .A(u5_mult_82_n6634), .ZN(u5_mult_82_n6639) );
  NOR2_X2 u5_mult_82_U2237 ( .A1(u5_mult_82_n6961), .A2(u5_mult_82_n6645), 
        .ZN(u5_mult_82_ab_24__2_) );
  NOR2_X2 u5_mult_82_U2236 ( .A1(u5_mult_82_n6960), .A2(u5_mult_82_n6674), 
        .ZN(u5_mult_82_ab_29__2_) );
  NOR2_X1 u5_mult_82_U2235 ( .A1(u5_mult_82_n6960), .A2(u5_mult_82_net65519), 
        .ZN(u5_mult_82_ab_34__2_) );
  NOR2_X2 u5_mult_82_U2234 ( .A1(u5_mult_82_n6953), .A2(u5_mult_82_n6710), 
        .ZN(u5_mult_82_ab_35__3_) );
  NOR2_X1 u5_mult_82_U2233 ( .A1(u5_mult_82_n6960), .A2(u5_mult_82_net65191), 
        .ZN(u5_mult_82_ab_51__2_) );
  NOR2_X1 u5_mult_82_U2232 ( .A1(u5_mult_82_net65189), .A2(u5_mult_82_n6759), 
        .ZN(u5_mult_82_ab_51__51_) );
  NOR2_X1 u5_mult_82_U2231 ( .A1(u5_mult_82_n6983), .A2(u5_mult_82_net65229), 
        .ZN(u5_mult_82_ab_50__52_) );
  NOR2_X1 u5_mult_82_U2230 ( .A1(u5_mult_82_n6976), .A2(u5_mult_82_n6884), 
        .ZN(u5_mult_82_ab_52__25_) );
  INV_X4 u5_mult_82_U2229 ( .A(u5_mult_82_n6926), .ZN(u5_mult_82_n6930) );
  NOR2_X2 u5_mult_82_U2228 ( .A1(u5_mult_82_n6913), .A2(u5_mult_82_net65443), 
        .ZN(u5_mult_82_ab_38__19_) );
  INV_X8 u5_mult_82_U2227 ( .A(u5_mult_82_net64571), .ZN(u5_mult_82_net64567)
         );
  NOR2_X2 u5_mult_82_U2226 ( .A1(u5_mult_82_net64223), .A2(u5_mult_82_n6952), 
        .ZN(u5_mult_82_ab_0__3_) );
  NOR2_X2 u5_mult_82_U2225 ( .A1(u5_mult_82_n6955), .A2(u5_mult_82_n6524), 
        .ZN(u5_mult_82_ab_4__3_) );
  NOR2_X2 u5_mult_82_U2224 ( .A1(u5_mult_82_n6955), .A2(u5_mult_82_n6547), 
        .ZN(u5_mult_82_ab_9__3_) );
  NOR2_X2 u5_mult_82_U2223 ( .A1(u5_mult_82_n6955), .A2(u5_mult_82_n6581), 
        .ZN(u5_mult_82_ab_14__3_) );
  NOR2_X2 u5_mult_82_U2222 ( .A1(u5_mult_82_n6954), .A2(u5_mult_82_n6617), 
        .ZN(u5_mult_82_ab_19__3_) );
  NOR2_X2 u5_mult_82_U2221 ( .A1(u5_mult_82_n6954), .A2(u5_mult_82_n6645), 
        .ZN(u5_mult_82_ab_24__3_) );
  NOR2_X2 u5_mult_82_U2220 ( .A1(u5_mult_82_n6953), .A2(u5_mult_82_n6674), 
        .ZN(u5_mult_82_ab_29__3_) );
  NOR2_X1 u5_mult_82_U2219 ( .A1(u5_mult_82_n6946), .A2(u5_mult_82_net65445), 
        .ZN(u5_mult_82_ab_38__4_) );
  INV_X8 u5_mult_82_U2218 ( .A(u5_mult_82_n6733), .ZN(u5_mult_82_n6738) );
  NAND3_X2 u5_mult_82_U2217 ( .A1(u5_mult_82_n3247), .A2(u5_mult_82_n3248), 
        .A3(u5_mult_82_n3249), .ZN(u5_mult_82_CARRYB_50__3_) );
  NOR2_X1 u5_mult_82_U2216 ( .A1(u5_mult_82_n6976), .A2(u5_mult_82_n6879), 
        .ZN(u5_mult_82_ab_52__26_) );
  INV_X4 u5_mult_82_U2215 ( .A(u5_mult_82_ab_50__25_), .ZN(u5_mult_82_n3274)
         );
  INV_X4 u5_mult_82_U2214 ( .A(u5_mult_82_ab_51__24_), .ZN(u5_mult_82_n3276)
         );
  NOR2_X1 u5_mult_82_U2213 ( .A1(u5_mult_82_n6927), .A2(u5_mult_82_n6715), 
        .ZN(u5_mult_82_ab_36__17_) );
  NOR2_X2 u5_mult_82_U2212 ( .A1(u5_mult_82_net64223), .A2(u5_mult_82_n6945), 
        .ZN(u5_mult_82_ab_0__4_) );
  NOR2_X2 u5_mult_82_U2211 ( .A1(u5_mult_82_n6948), .A2(u5_mult_82_n6523), 
        .ZN(u5_mult_82_ab_4__4_) );
  NOR2_X2 u5_mult_82_U2210 ( .A1(u5_mult_82_n6948), .A2(u5_mult_82_n6546), 
        .ZN(u5_mult_82_ab_9__4_) );
  NOR2_X1 u5_mult_82_U2209 ( .A1(u5_mult_82_n6948), .A2(u5_mult_82_n6580), 
        .ZN(u5_mult_82_ab_14__4_) );
  NOR2_X1 u5_mult_82_U2208 ( .A1(u5_mult_82_net64363), .A2(u5_mult_82_n6644), 
        .ZN(u5_mult_82_ab_24__5_) );
  NOR2_X1 u5_mult_82_U2207 ( .A1(u5_mult_82_n6946), .A2(u5_mult_82_n6673), 
        .ZN(u5_mult_82_ab_29__4_) );
  NOR2_X1 u5_mult_82_U2206 ( .A1(u5_mult_82_net64361), .A2(u5_mult_82_n6673), 
        .ZN(u5_mult_82_ab_29__5_) );
  NOR2_X1 u5_mult_82_U2205 ( .A1(u5_mult_82_net64523), .A2(u5_mult_82_net65189), .ZN(u5_mult_82_ab_51__14_) );
  NOR2_X1 u5_mult_82_U2204 ( .A1(u5_mult_82_net64559), .A2(u5_mult_82_net65189), .ZN(u5_mult_82_ab_51__16_) );
  NOR2_X1 u5_mult_82_U2203 ( .A1(u5_mult_82_n6927), .A2(u5_mult_82_net65189), 
        .ZN(u5_mult_82_ab_51__17_) );
  NOR2_X1 u5_mult_82_U2202 ( .A1(u5_mult_82_net64683), .A2(u5_mult_82_net65229), .ZN(u5_mult_82_ab_50__23_) );
  NOR2_X1 u5_mult_82_U2201 ( .A1(u5_mult_82_n6856), .A2(u5_mult_82_net65191), 
        .ZN(u5_mult_82_ab_51__30_) );
  NOR2_X2 u5_mult_82_U2200 ( .A1(u5_mult_82_net64899), .A2(u5_mult_82_net65193), .ZN(u5_mult_82_ab_51__35_) );
  NOR2_X1 u5_mult_82_U2199 ( .A1(u5_mult_82_net64935), .A2(u5_mult_82_net65193), .ZN(u5_mult_82_ab_51__37_) );
  INV_X4 u5_mult_82_U2198 ( .A(u5_mult_82_n6978), .ZN(u5_mult_82_n6977) );
  NOR2_X1 u5_mult_82_U2197 ( .A1(u5_mult_82_n6777), .A2(u5_mult_82_net65189), 
        .ZN(u5_mult_82_ab_51__48_) );
  NOR2_X1 u5_mult_82_U2196 ( .A1(u5_mult_82_n6816), .A2(u5_mult_82_net65193), 
        .ZN(u5_mult_82_ab_51__42_) );
  NOR2_X1 u5_mult_82_U2195 ( .A1(u5_mult_82_n6826), .A2(u5_mult_82_net65193), 
        .ZN(u5_mult_82_ab_51__40_) );
  NOR2_X1 u5_mult_82_U2194 ( .A1(u5_mult_82_net64559), .A2(u5_mult_82_n6708), 
        .ZN(u5_mult_82_ab_35__16_) );
  INV_X4 u5_mult_82_U2193 ( .A(u5_mult_82_ab_24__21_), .ZN(u5_mult_82_n3281)
         );
  NOR2_X2 u5_mult_82_U2192 ( .A1(u5_mult_82_n6892), .A2(u5_mult_82_net65677), 
        .ZN(u5_mult_82_ab_25__24_) );
  NOR2_X2 u5_mult_82_U2191 ( .A1(u5_mult_82_n6914), .A2(u5_mult_82_net65677), 
        .ZN(u5_mult_82_ab_25__19_) );
  NOR2_X1 u5_mult_82_U2190 ( .A1(u5_mult_82_n6914), .A2(u5_mult_82_n6643), 
        .ZN(u5_mult_82_ab_24__19_) );
  NOR2_X2 u5_mult_82_U2189 ( .A1(u5_mult_82_net64365), .A2(u5_mult_82_n6523), 
        .ZN(u5_mult_82_ab_4__5_) );
  NOR2_X2 u5_mult_82_U2188 ( .A1(u5_mult_82_net64365), .A2(u5_mult_82_n6546), 
        .ZN(u5_mult_82_ab_9__5_) );
  NOR2_X1 u5_mult_82_U2187 ( .A1(u5_mult_82_net64365), .A2(u5_mult_82_n6580), 
        .ZN(u5_mult_82_ab_14__5_) );
  NOR2_X2 u5_mult_82_U2186 ( .A1(u5_mult_82_net64381), .A2(u5_mult_82_n6610), 
        .ZN(u5_mult_82_ab_18__6_) );
  NOR2_X1 u5_mult_82_U2185 ( .A1(u5_mult_82_net64379), .A2(u5_mult_82_n6701), 
        .ZN(u5_mult_82_ab_33__6_) );
  NOR2_X1 u5_mult_82_U2184 ( .A1(u5_mult_82_net64379), .A2(u5_mult_82_net65445), .ZN(u5_mult_82_ab_38__6_) );
  NAND2_X2 u5_mult_82_U2183 ( .A1(u5_mult_82_ab_44__4_), .A2(
        u5_mult_82_CARRYB_43__4_), .ZN(u5_mult_82_n5788) );
  INV_X4 u5_mult_82_U2182 ( .A(u5_mult_82_ab_49__7_), .ZN(u5_mult_82_n1335) );
  NOR2_X1 u5_mult_82_U2181 ( .A1(u5_mult_82_n6940), .A2(u5_mult_82_net65191), 
        .ZN(u5_mult_82_ab_51__7_) );
  NOR2_X1 u5_mult_82_U2180 ( .A1(u5_mult_82_net64433), .A2(u5_mult_82_n6755), 
        .ZN(u5_mult_82_ab_49__9_) );
  NOR2_X1 u5_mult_82_U2179 ( .A1(u5_mult_82_net64455), .A2(u5_mult_82_net65229), .ZN(u5_mult_82_ab_50__10_) );
  NAND2_X2 u5_mult_82_U2178 ( .A1(u5_mult_82_CARRYB_49__19_), .A2(
        u5_mult_82_n1841), .ZN(u5_mult_82_n5568) );
  NOR2_X1 u5_mult_82_U2177 ( .A1(u5_mult_82_n6861), .A2(u5_mult_82_net65225), 
        .ZN(u5_mult_82_ab_50__29_) );
  NOR2_X1 u5_mult_82_U2176 ( .A1(u5_mult_82_n6842), .A2(u5_mult_82_net65225), 
        .ZN(u5_mult_82_ab_50__32_) );
  NOR2_X2 u5_mult_82_U2175 ( .A1(u5_mult_82_net64881), .A2(u5_mult_82_n6753), 
        .ZN(u5_mult_82_ab_49__34_) );
  NOR2_X1 u5_mult_82_U2174 ( .A1(u5_mult_82_n6784), .A2(u5_mult_82_net65223), 
        .ZN(u5_mult_82_ab_50__47_) );
  NOR2_X2 u5_mult_82_U2173 ( .A1(u5_mult_82_n6797), .A2(u5_mult_82_net65223), 
        .ZN(u5_mult_82_ab_50__45_) );
  NOR2_X1 u5_mult_82_U2172 ( .A1(u5_mult_82_n6803), .A2(u5_mult_82_net65223), 
        .ZN(u5_mult_82_ab_50__44_) );
  NOR2_X1 u5_mult_82_U2171 ( .A1(u5_mult_82_n6831), .A2(u5_mult_82_net65225), 
        .ZN(u5_mult_82_ab_50__39_) );
  NOR2_X2 u5_mult_82_U2170 ( .A1(u5_mult_82_n6896), .A2(u5_mult_82_n6700), 
        .ZN(u5_mult_82_ab_33__21_) );
  NOR2_X2 u5_mult_82_U2169 ( .A1(u5_mult_82_n6886), .A2(u5_mult_82_n6643), 
        .ZN(u5_mult_82_ab_24__25_) );
  NOR2_X2 u5_mult_82_U2168 ( .A1(u5_mult_82_n6881), .A2(u5_mult_82_n6643), 
        .ZN(u5_mult_82_ab_24__26_) );
  NOR2_X2 u5_mult_82_U2167 ( .A1(u5_mult_82_net64223), .A2(u5_mult_82_n1271), 
        .ZN(u5_mult_82_ab_0__6_) );
  NOR2_X2 u5_mult_82_U2166 ( .A1(u5_mult_82_net64383), .A2(u5_mult_82_n6523), 
        .ZN(u5_mult_82_ab_4__6_) );
  NOR2_X2 u5_mult_82_U2165 ( .A1(u5_mult_82_net64383), .A2(u5_mult_82_n6546), 
        .ZN(u5_mult_82_ab_9__6_) );
  NOR2_X1 u5_mult_82_U2164 ( .A1(u5_mult_82_n6941), .A2(u5_mult_82_n6616), 
        .ZN(u5_mult_82_ab_19__7_) );
  NOR2_X1 u5_mult_82_U2163 ( .A1(u5_mult_82_n6940), .A2(u5_mult_82_n6736), 
        .ZN(u5_mult_82_ab_44__7_) );
  NOR2_X1 u5_mult_82_U2162 ( .A1(u5_mult_82_net64505), .A2(u5_mult_82_n6748), 
        .ZN(u5_mult_82_ab_48__13_) );
  NOR2_X2 u5_mult_82_U2161 ( .A1(u5_mult_82_n6895), .A2(u5_mult_82_n6749), 
        .ZN(u5_mult_82_ab_48__21_) );
  INV_X4 u5_mult_82_U2160 ( .A(u5_mult_82_ab_21__26_), .ZN(u5_mult_82_n2750)
         );
  NOR2_X1 u5_mult_82_U2159 ( .A1(u5_mult_82_n6876), .A2(u5_mult_82_net65713), 
        .ZN(u5_mult_82_ab_23__27_) );
  NOR2_X1 u5_mult_82_U2158 ( .A1(u5_mult_82_n6892), .A2(u5_mult_82_n6615), 
        .ZN(u5_mult_82_ab_19__24_) );
  NOR2_X2 u5_mult_82_U2157 ( .A1(u5_mult_82_net64223), .A2(u5_mult_82_n6939), 
        .ZN(u5_mult_82_ab_0__7_) );
  NOR2_X2 u5_mult_82_U2156 ( .A1(u5_mult_82_n6942), .A2(u5_mult_82_n6523), 
        .ZN(u5_mult_82_ab_4__7_) );
  NOR2_X2 u5_mult_82_U2155 ( .A1(u5_mult_82_n6942), .A2(u5_mult_82_n6546), 
        .ZN(u5_mult_82_ab_9__7_) );
  NOR2_X1 u5_mult_82_U2154 ( .A1(u5_mult_82_net64417), .A2(u5_mult_82_n6616), 
        .ZN(u5_mult_82_ab_19__8_) );
  NOR2_X1 u5_mult_82_U2153 ( .A1(u5_mult_82_net64435), .A2(u5_mult_82_n6616), 
        .ZN(u5_mult_82_ab_19__9_) );
  NOR2_X1 u5_mult_82_U2152 ( .A1(u5_mult_82_n6941), .A2(u5_mult_82_n6644), 
        .ZN(u5_mult_82_ab_24__7_) );
  INV_X4 u5_mult_82_U2151 ( .A(u5_mult_82_ab_33__7_), .ZN(u5_mult_82_n1458) );
  NAND3_X2 u5_mult_82_U2150 ( .A1(u5_mult_82_n3789), .A2(u5_mult_82_n3790), 
        .A3(u5_mult_82_n3791), .ZN(u5_mult_82_CARRYB_33__7_) );
  INV_X4 u5_mult_82_U2149 ( .A(u5_mult_82_n1687), .ZN(u5_mult_82_n1688) );
  INV_X4 u5_mult_82_U2148 ( .A(u5_mult_82_ab_46__27_), .ZN(u5_mult_82_n1914)
         );
  NOR2_X1 u5_mult_82_U2147 ( .A1(u5_mult_82_n6983), .A2(u5_mult_82_net65321), 
        .ZN(u5_mult_82_ab_45__52_) );
  NOR2_X2 u5_mult_82_U2146 ( .A1(u5_mult_82_n6759), .A2(u5_mult_82_n6741), 
        .ZN(u5_mult_82_ab_46__51_) );
  INV_X4 u5_mult_82_U2145 ( .A(u5_mult_82_ab_46__28_), .ZN(u5_mult_82_n1117)
         );
  NOR2_X2 u5_mult_82_U2144 ( .A1(u5_mult_82_n6849), .A2(u5_mult_82_net65315), 
        .ZN(u5_mult_82_ab_45__31_) );
  NOR2_X2 u5_mult_82_U2143 ( .A1(u5_mult_82_net64223), .A2(u5_mult_82_net64427), .ZN(u5_mult_82_ab_0__8_) );
  NOR2_X2 u5_mult_82_U2142 ( .A1(u5_mult_82_net64419), .A2(u5_mult_82_n6523), 
        .ZN(u5_mult_82_ab_4__8_) );
  NOR2_X2 u5_mult_82_U2141 ( .A1(u5_mult_82_net64419), .A2(u5_mult_82_n6546), 
        .ZN(u5_mult_82_ab_9__8_) );
  NOR2_X2 u5_mult_82_U2140 ( .A1(u5_mult_82_net64435), .A2(u5_mult_82_n6658), 
        .ZN(u5_mult_82_ab_27__9_) );
  INV_X4 u5_mult_82_U2139 ( .A(u5_mult_82_ab_27__11_), .ZN(u5_mult_82_n3590)
         );
  NOR2_X2 u5_mult_82_U2138 ( .A1(u5_mult_82_n6941), .A2(u5_mult_82_net65409), 
        .ZN(u5_mult_82_ab_40__7_) );
  NOR2_X2 u5_mult_82_U2137 ( .A1(u5_mult_82_n6884), .A2(u5_mult_82_net65321), 
        .ZN(u5_mult_82_ab_45__25_) );
  NOR2_X2 u5_mult_82_U2136 ( .A1(u5_mult_82_n6826), .A2(u5_mult_82_n6736), 
        .ZN(u5_mult_82_ab_44__40_) );
  NOR2_X1 u5_mult_82_U2135 ( .A1(u5_mult_82_n6831), .A2(u5_mult_82_n6734), 
        .ZN(u5_mult_82_ab_44__39_) );
  NOR2_X2 u5_mult_82_U2134 ( .A1(u5_mult_82_n6856), .A2(u5_mult_82_net65351), 
        .ZN(u5_mult_82_ab_43__30_) );
  NOR2_X2 u5_mult_82_U2133 ( .A1(u5_mult_82_net64667), .A2(u5_mult_82_n6672), 
        .ZN(u5_mult_82_ab_29__22_) );
  NOR2_X2 u5_mult_82_U2132 ( .A1(u5_mult_82_n6885), .A2(u5_mult_82_n6679), 
        .ZN(u5_mult_82_ab_30__25_) );
  INV_X4 u5_mult_82_U2131 ( .A(u5_mult_82_ab_19__21_), .ZN(u5_mult_82_n700) );
  NOR2_X1 u5_mult_82_U2130 ( .A1(u5_mult_82_n6914), .A2(u5_mult_82_n6615), 
        .ZN(u5_mult_82_ab_19__19_) );
  NOR2_X2 u5_mult_82_U2129 ( .A1(u5_mult_82_net64437), .A2(u5_mult_82_n6523), 
        .ZN(u5_mult_82_ab_4__9_) );
  NOR2_X2 u5_mult_82_U2128 ( .A1(u5_mult_82_net64437), .A2(u5_mult_82_n6546), 
        .ZN(u5_mult_82_ab_9__9_) );
  NOR2_X1 u5_mult_82_U2127 ( .A1(u5_mult_82_net64455), .A2(u5_mult_82_n6573), 
        .ZN(u5_mult_82_ab_13__10_) );
  NOR2_X1 u5_mult_82_U2126 ( .A1(u5_mult_82_net64453), .A2(u5_mult_82_n6616), 
        .ZN(u5_mult_82_ab_19__10_) );
  NOR2_X2 u5_mult_82_U2125 ( .A1(u5_mult_82_net64453), .A2(u5_mult_82_n6644), 
        .ZN(u5_mult_82_ab_24__10_) );
  NAND3_X2 u5_mult_82_U2124 ( .A1(u5_mult_82_n4151), .A2(u5_mult_82_n4152), 
        .A3(u5_mult_82_n4153), .ZN(u5_mult_82_CARRYB_33__10_) );
  NOR2_X2 u5_mult_82_U2123 ( .A1(u5_mult_82_net64417), .A2(u5_mult_82_net65409), .ZN(u5_mult_82_ab_40__8_) );
  INV_X4 u5_mult_82_U2122 ( .A(u5_mult_82_ab_44__12_), .ZN(u5_mult_82_n5246)
         );
  NOR2_X1 u5_mult_82_U2121 ( .A1(u5_mult_82_net64559), .A2(u5_mult_82_net65321), .ZN(u5_mult_82_ab_45__16_) );
  NOR2_X2 u5_mult_82_U2120 ( .A1(u5_mult_82_n6912), .A2(u5_mult_82_net65321), 
        .ZN(u5_mult_82_ab_45__19_) );
  NOR2_X1 u5_mult_82_U2119 ( .A1(u5_mult_82_n6891), .A2(u5_mult_82_n6735), 
        .ZN(u5_mult_82_ab_44__24_) );
  NOR2_X2 u5_mult_82_U2118 ( .A1(u5_mult_82_net64683), .A2(u5_mult_82_net65353), .ZN(u5_mult_82_ab_43__23_) );
  NOR2_X1 u5_mult_82_U2117 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6734), 
        .ZN(u5_mult_82_ab_44__36_) );
  NOR2_X2 u5_mult_82_U2116 ( .A1(u5_mult_82_net64935), .A2(u5_mult_82_n6734), 
        .ZN(u5_mult_82_ab_44__37_) );
  NOR2_X1 u5_mult_82_U2115 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6734), 
        .ZN(u5_mult_82_ab_44__38_) );
  NOR2_X1 u5_mult_82_U2114 ( .A1(u5_mult_82_n6816), .A2(u5_mult_82_net65349), 
        .ZN(u5_mult_82_ab_43__42_) );
  NOR2_X2 u5_mult_82_U2113 ( .A1(u5_mult_82_n6838), .A2(u5_mult_82_net65387), 
        .ZN(u5_mult_82_ab_41__33_) );
  NAND3_X2 u5_mult_82_U2112 ( .A1(u5_mult_82_n5535), .A2(u5_mult_82_n5536), 
        .A3(u5_mult_82_n5537), .ZN(u5_mult_82_CARRYB_27__24_) );
  NOR2_X1 u5_mult_82_U2111 ( .A1(u5_mult_82_n6891), .A2(u5_mult_82_n6664), 
        .ZN(u5_mult_82_ab_28__24_) );
  NOR2_X1 u5_mult_82_U2110 ( .A1(u5_mult_82_n6868), .A2(u5_mult_82_n6663), 
        .ZN(u5_mult_82_ab_28__28_) );
  INV_X4 u5_mult_82_U2109 ( .A(u5_mult_82_ab_30__17_), .ZN(u5_mult_82_n3666)
         );
  NOR2_X2 u5_mult_82_U2108 ( .A1(u5_mult_82_n6858), .A2(u5_mult_82_n6601), 
        .ZN(u5_mult_82_ab_17__30_) );
  NOR2_X2 u5_mult_82_U2107 ( .A1(u5_mult_82_n6869), .A2(u5_mult_82_n6594), 
        .ZN(u5_mult_82_ab_16__28_) );
  NOR2_X2 u5_mult_82_U2106 ( .A1(u5_mult_82_n6882), .A2(u5_mult_82_n6587), 
        .ZN(u5_mult_82_ab_15__26_) );
  NOR2_X2 u5_mult_82_U2105 ( .A1(u5_mult_82_net64223), .A2(u5_mult_82_net64451), .ZN(u5_mult_82_ab_0__10_) );
  NOR2_X1 u5_mult_82_U2104 ( .A1(u5_mult_82_net64455), .A2(u5_mult_82_n6523), 
        .ZN(u5_mult_82_ab_4__10_) );
  NOR2_X1 u5_mult_82_U2103 ( .A1(u5_mult_82_net64473), .A2(u5_mult_82_n6580), 
        .ZN(u5_mult_82_ab_14__11_) );
  NOR2_X2 u5_mult_82_U2102 ( .A1(u5_mult_82_net64491), .A2(u5_mult_82_n6588), 
        .ZN(u5_mult_82_ab_15__12_) );
  NAND3_X2 u5_mult_82_U2101 ( .A1(u5_mult_82_n2045), .A2(u5_mult_82_n2046), 
        .A3(u5_mult_82_n2047), .ZN(u5_mult_82_CARRYB_21__11_) );
  NOR2_X2 u5_mult_82_U2100 ( .A1(u5_mult_82_net64471), .A2(u5_mult_82_n6637), 
        .ZN(u5_mult_82_ab_22__11_) );
  NOR2_X1 u5_mult_82_U2099 ( .A1(u5_mult_82_net64525), .A2(u5_mult_82_net65713), .ZN(u5_mult_82_ab_23__14_) );
  INV_X4 u5_mult_82_U2098 ( .A(u5_mult_82_ab_26__13_), .ZN(u5_mult_82_n2042)
         );
  NOR2_X1 u5_mult_82_U2097 ( .A1(u5_mult_82_net64487), .A2(u5_mult_82_n6701), 
        .ZN(u5_mult_82_ab_33__12_) );
  NAND2_X2 u5_mult_82_U2096 ( .A1(u5_mult_82_n5282), .A2(u5_mult_82_ab_43__16_), .ZN(u5_mult_82_n5285) );
  NAND2_X2 u5_mult_82_U2095 ( .A1(u5_mult_82_n5284), .A2(u5_mult_82_n5285), 
        .ZN(u5_mult_82_n5880) );
  NOR2_X2 u5_mult_82_U2094 ( .A1(u5_mult_82_net64913), .A2(u5_mult_82_net65369), .ZN(u5_mult_82_ab_42__35_) );
  NOR2_X2 u5_mult_82_U2093 ( .A1(u5_mult_82_n6772), .A2(u5_mult_82_net65313), 
        .ZN(u5_mult_82_ab_45__49_) );
  NOR2_X2 u5_mult_82_U2092 ( .A1(u5_mult_82_n6777), .A2(u5_mult_82_net65313), 
        .ZN(u5_mult_82_ab_45__48_) );
  NOR2_X1 u5_mult_82_U2091 ( .A1(u5_mult_82_n6784), .A2(u5_mult_82_net65313), 
        .ZN(u5_mult_82_ab_45__47_) );
  NOR2_X2 u5_mult_82_U2090 ( .A1(u5_mult_82_n6858), .A2(u5_mult_82_n6656), 
        .ZN(u5_mult_82_ab_27__30_) );
  NAND3_X2 u5_mult_82_U2089 ( .A1(u5_mult_82_n5338), .A2(u5_mult_82_n5339), 
        .A3(u5_mult_82_n5340), .ZN(u5_mult_82_CARRYB_15__29_) );
  NOR2_X1 u5_mult_82_U2088 ( .A1(u5_mult_82_n6851), .A2(u5_mult_82_n6608), 
        .ZN(u5_mult_82_ab_18__31_) );
  NOR2_X2 u5_mult_82_U2087 ( .A1(u5_mult_82_n6844), .A2(u5_mult_82_n6608), 
        .ZN(u5_mult_82_ab_18__32_) );
  NOR2_X2 u5_mult_82_U2086 ( .A1(u5_mult_82_net64473), .A2(u5_mult_82_n6523), 
        .ZN(u5_mult_82_ab_4__11_) );
  INV_X4 u5_mult_82_U2085 ( .A(u5_mult_82_ab_28__14_), .ZN(u5_mult_82_n1912)
         );
  NOR2_X1 u5_mult_82_U2084 ( .A1(u5_mult_82_net64469), .A2(u5_mult_82_net65445), .ZN(u5_mult_82_ab_38__11_) );
  NAND3_X2 u5_mult_82_U2083 ( .A1(u5_mult_82_n6162), .A2(u5_mult_82_n6163), 
        .A3(u5_mult_82_n6164), .ZN(u5_mult_82_CARRYB_42__10_) );
  NOR2_X2 u5_mult_82_U2082 ( .A1(u5_mult_82_n6904), .A2(u5_mult_82_net65389), 
        .ZN(u5_mult_82_ab_41__20_) );
  NOR2_X2 u5_mult_82_U2081 ( .A1(u5_mult_82_n6896), .A2(u5_mult_82_net65389), 
        .ZN(u5_mult_82_ab_41__21_) );
  NOR2_X1 u5_mult_82_U2080 ( .A1(u5_mult_82_n6797), .A2(u5_mult_82_net65385), 
        .ZN(u5_mult_82_ab_41__45_) );
  NOR2_X1 u5_mult_82_U2079 ( .A1(u5_mult_82_net64689), .A2(u5_mult_82_n6579), 
        .ZN(u5_mult_82_ab_14__23_) );
  NOR2_X2 u5_mult_82_U2078 ( .A1(u5_mult_82_net64671), .A2(u5_mult_82_n6579), 
        .ZN(u5_mult_82_ab_14__22_) );
  INV_X4 u5_mult_82_U2077 ( .A(u5_mult_82_ab_13__23_), .ZN(u5_mult_82_n2309)
         );
  NOR2_X2 u5_mult_82_U2076 ( .A1(u5_mult_82_net64491), .A2(u5_mult_82_n6523), 
        .ZN(u5_mult_82_ab_4__12_) );
  NAND2_X2 u5_mult_82_U2075 ( .A1(u5_mult_82_ab_28__13_), .A2(u5_mult_82_n1848), .ZN(u5_mult_82_n2597) );
  NOR2_X1 u5_mult_82_U2074 ( .A1(u5_mult_82_net64505), .A2(u5_mult_82_net65391), .ZN(u5_mult_82_ab_41__13_) );
  NOR2_X1 u5_mult_82_U2073 ( .A1(u5_mult_82_n6791), .A2(u5_mult_82_net65385), 
        .ZN(u5_mult_82_ab_41__46_) );
  NOR2_X2 u5_mult_82_U2072 ( .A1(u5_mult_82_n6876), .A2(u5_mult_82_n6643), 
        .ZN(u5_mult_82_ab_24__27_) );
  INV_X2 u5_mult_82_U2071 ( .A(u5_mult_82_ab_23__28_), .ZN(u5_mult_82_n1747)
         );
  NOR2_X2 u5_mult_82_U2070 ( .A1(u5_mult_82_net64887), .A2(u5_mult_82_n6565), 
        .ZN(u5_mult_82_ab_12__34_) );
  NOR2_X2 u5_mult_82_U2069 ( .A1(u5_mult_82_n6915), .A2(u5_mult_82_n6587), 
        .ZN(u5_mult_82_ab_15__19_) );
  INV_X2 u5_mult_82_U2068 ( .A(u5_mult_82_ab_12__23_), .ZN(u5_mult_82_n805) );
  NOR2_X2 u5_mult_82_U2067 ( .A1(u5_mult_82_n6898), .A2(u5_mult_82_n6579), 
        .ZN(u5_mult_82_ab_14__21_) );
  NOR2_X1 u5_mult_82_U2066 ( .A1(u5_mult_82_n6845), .A2(u5_mult_82_n6550), 
        .ZN(u5_mult_82_ab_10__32_) );
  NOR2_X2 u5_mult_82_U2065 ( .A1(u5_mult_82_net64509), .A2(u5_mult_82_n6523), 
        .ZN(u5_mult_82_ab_4__13_) );
  NOR2_X2 u5_mult_82_U2064 ( .A1(u5_mult_82_net64527), .A2(u5_mult_82_n6537), 
        .ZN(u5_mult_82_ab_8__14_) );
  NOR2_X2 u5_mult_82_U2063 ( .A1(u5_mult_82_n6935), .A2(u5_mult_82_n6546), 
        .ZN(u5_mult_82_ab_9__15_) );
  NOR2_X2 u5_mult_82_U2062 ( .A1(u5_mult_82_net64525), .A2(u5_mult_82_n6610), 
        .ZN(u5_mult_82_ab_18__14_) );
  NOR2_X1 u5_mult_82_U2061 ( .A1(u5_mult_82_net64523), .A2(u5_mult_82_n6716), 
        .ZN(u5_mult_82_ab_36__14_) );
  NOR2_X2 u5_mult_82_U2060 ( .A1(u5_mult_82_n6875), .A2(u5_mult_82_net65443), 
        .ZN(u5_mult_82_ab_38__27_) );
  NOR2_X2 u5_mult_82_U2059 ( .A1(u5_mult_82_n6880), .A2(u5_mult_82_n6721), 
        .ZN(u5_mult_82_ab_37__26_) );
  NOR2_X1 u5_mult_82_U2058 ( .A1(u5_mult_82_n6827), .A2(u5_mult_82_net65445), 
        .ZN(u5_mult_82_ab_38__40_) );
  NOR2_X1 u5_mult_82_U2057 ( .A1(u5_mult_82_n6832), .A2(u5_mult_82_n6720), 
        .ZN(u5_mult_82_ab_37__39_) );
  NOR2_X1 u5_mult_82_U2056 ( .A1(u5_mult_82_n6821), .A2(u5_mult_82_net65445), 
        .ZN(u5_mult_82_ab_38__41_) );
  NOR2_X1 u5_mult_82_U2055 ( .A1(u5_mult_82_n6804), .A2(u5_mult_82_net65445), 
        .ZN(u5_mult_82_ab_38__44_) );
  NOR2_X1 u5_mult_82_U2054 ( .A1(u5_mult_82_n6811), .A2(u5_mult_82_net65445), 
        .ZN(u5_mult_82_ab_38__43_) );
  NOR2_X1 u5_mult_82_U2053 ( .A1(u5_mult_82_n6816), .A2(u5_mult_82_net65445), 
        .ZN(u5_mult_82_ab_38__42_) );
  NOR2_X1 u5_mult_82_U2052 ( .A1(u5_mult_82_n6983), .A2(u5_mult_82_n6730), 
        .ZN(u5_mult_82_ab_39__52_) );
  NOR2_X2 u5_mult_82_U2051 ( .A1(u5_mult_82_n6761), .A2(u5_mult_82_net65403), 
        .ZN(u5_mult_82_ab_40__51_) );
  INV_X2 u5_mult_82_U2050 ( .A(u5_mult_82_ab_39__36_), .ZN(u5_mult_82_n3931)
         );
  NOR2_X2 u5_mult_82_U2049 ( .A1(u5_mult_82_n6839), .A2(u5_mult_82_n6635), 
        .ZN(u5_mult_82_ab_22__33_) );
  NOR2_X1 u5_mult_82_U2048 ( .A1(u5_mult_82_n6840), .A2(u5_mult_82_n6557), 
        .ZN(u5_mult_82_ab_11__33_) );
  INV_X4 u5_mult_82_U2047 ( .A(u5_mult_82_ab_11__36_), .ZN(u5_mult_82_n1245)
         );
  NOR2_X2 u5_mult_82_U2046 ( .A1(u5_mult_82_n6852), .A2(u5_mult_82_n6544), 
        .ZN(u5_mult_82_ab_9__31_) );
  NAND3_X2 u5_mult_82_U2045 ( .A1(u5_mult_82_n1015), .A2(u5_mult_82_n1016), 
        .A3(u5_mult_82_n1017), .ZN(u5_mult_82_CARRYB_25__15_) );
  INV_X4 u5_mult_82_U2044 ( .A(u5_mult_82_n1856), .ZN(u5_mult_82_n1857) );
  NAND3_X2 u5_mult_82_U2043 ( .A1(u5_mult_82_n3052), .A2(u5_mult_82_n3053), 
        .A3(u5_mult_82_n3054), .ZN(u5_mult_82_CARRYB_36__38_) );
  NOR2_X1 u5_mult_82_U2042 ( .A1(u5_mult_82_n6784), .A2(u5_mult_82_n6713), 
        .ZN(u5_mult_82_ab_36__47_) );
  NOR2_X2 u5_mult_82_U2041 ( .A1(u5_mult_82_n6779), .A2(u5_mult_82_net65403), 
        .ZN(u5_mult_82_ab_40__48_) );
  NOR2_X2 u5_mult_82_U2040 ( .A1(u5_mult_82_net64937), .A2(u5_mult_82_net65513), .ZN(u5_mult_82_ab_34__37_) );
  INV_X4 u5_mult_82_U2039 ( .A(u5_mult_82_ab_21__33_), .ZN(u5_mult_82_n3745)
         );
  NOR2_X2 u5_mult_82_U2038 ( .A1(u5_mult_82_net64923), .A2(u5_mult_82_n6565), 
        .ZN(u5_mult_82_ab_12__36_) );
  INV_X4 u5_mult_82_U2037 ( .A(u5_mult_82_ab_13__36_), .ZN(u5_mult_82_n1203)
         );
  NOR2_X1 u5_mult_82_U2036 ( .A1(u5_mult_82_n6898), .A2(u5_mult_82_n6558), 
        .ZN(u5_mult_82_ab_11__21_) );
  NOR2_X2 u5_mult_82_U2035 ( .A1(u5_mult_82_net64563), .A2(u5_mult_82_n6551), 
        .ZN(u5_mult_82_ab_10__16_) );
  NOR2_X2 u5_mult_82_U2034 ( .A1(u5_mult_82_n6915), .A2(u5_mult_82_n6545), 
        .ZN(u5_mult_82_ab_9__19_) );
  NOR2_X2 u5_mult_82_U2033 ( .A1(u5_mult_82_n6928), .A2(u5_mult_82_n6595), 
        .ZN(u5_mult_82_ab_16__17_) );
  NOR2_X2 u5_mult_82_U2032 ( .A1(u5_mult_82_n6768), .A2(u5_mult_82_net65403), 
        .ZN(u5_mult_82_ab_40__50_) );
  NOR2_X2 u5_mult_82_U2031 ( .A1(u5_mult_82_n6774), .A2(u5_mult_82_net65403), 
        .ZN(u5_mult_82_ab_40__49_) );
  NOR2_X1 u5_mult_82_U2030 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6699), 
        .ZN(u5_mult_82_ab_33__36_) );
  NOR2_X1 u5_mult_82_U2029 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6614), 
        .ZN(u5_mult_82_ab_19__36_) );
  NAND3_X2 u5_mult_82_U2028 ( .A1(u5_mult_82_n1012), .A2(u5_mult_82_n1013), 
        .A3(u5_mult_82_n1014), .ZN(u5_mult_82_CARRYB_7__26_) );
  NOR2_X2 u5_mult_82_U2027 ( .A1(u5_mult_82_n6882), .A2(u5_mult_82_n6536), 
        .ZN(u5_mult_82_ab_8__26_) );
  NOR2_X2 u5_mult_82_U2026 ( .A1(u5_mult_82_n6864), .A2(u5_mult_82_n6528), 
        .ZN(u5_mult_82_ab_7__29_) );
  NOR2_X2 u5_mult_82_U2025 ( .A1(u5_mult_82_net64565), .A2(u5_mult_82_net66091), .ZN(u5_mult_82_ab_2__16_) );
  NOR2_X1 u5_mult_82_U2024 ( .A1(u5_mult_82_n6891), .A2(u5_mult_82_net65515), 
        .ZN(u5_mult_82_ab_34__24_) );
  NOR2_X1 u5_mult_82_U2023 ( .A1(u5_mult_82_n6868), .A2(u5_mult_82_n6699), 
        .ZN(u5_mult_82_ab_33__28_) );
  INV_X4 u5_mult_82_U2022 ( .A(u5_mult_82_n1574), .ZN(u5_mult_82_n1575) );
  NOR2_X1 u5_mult_82_U2021 ( .A1(u5_mult_82_net64901), .A2(u5_mult_82_n6699), 
        .ZN(u5_mult_82_ab_33__35_) );
  NOR2_X1 u5_mult_82_U2020 ( .A1(u5_mult_82_n6797), .A2(u5_mult_82_net65515), 
        .ZN(u5_mult_82_ab_34__45_) );
  NOR2_X2 u5_mult_82_U2019 ( .A1(u5_mult_82_n6827), .A2(u5_mult_82_n6701), 
        .ZN(u5_mult_82_ab_33__40_) );
  INV_X4 u5_mult_82_U2018 ( .A(u5_mult_82_ab_17__36_), .ZN(u5_mult_82_n3501)
         );
  NOR2_X2 u5_mult_82_U2017 ( .A1(u5_mult_82_net64959), .A2(u5_mult_82_n6528), 
        .ZN(u5_mult_82_ab_7__38_) );
  NOR2_X2 u5_mult_82_U2016 ( .A1(u5_mult_82_net64959), .A2(u5_mult_82_n6565), 
        .ZN(u5_mult_82_ab_12__38_) );
  NOR2_X2 u5_mult_82_U2015 ( .A1(u5_mult_82_n6915), .A2(u5_mult_82_n6558), 
        .ZN(u5_mult_82_ab_11__19_) );
  INV_X4 u5_mult_82_U2014 ( .A(u5_mult_82_ab_4__37_), .ZN(u5_mult_82_n2418) );
  INV_X4 u5_mult_82_U2013 ( .A(u5_mult_82_ab_5__36_), .ZN(u5_mult_82_n1364) );
  NAND2_X2 u5_mult_82_U2012 ( .A1(u5_mult_82_n1364), .A2(u5_mult_82_n1365), 
        .ZN(u5_mult_82_n1367) );
  NOR2_X2 u5_mult_82_U2011 ( .A1(u5_mult_82_n6929), .A2(u5_mult_82_net66091), 
        .ZN(u5_mult_82_ab_2__17_) );
  NOR2_X2 u5_mult_82_U2010 ( .A1(u5_mult_82_n6915), .A2(u5_mult_82_n6522), 
        .ZN(u5_mult_82_ab_4__19_) );
  NOR2_X1 u5_mult_82_U2009 ( .A1(u5_mult_82_n6804), .A2(u5_mult_82_n6686), 
        .ZN(u5_mult_82_ab_31__44_) );
  NOR2_X1 u5_mult_82_U2008 ( .A1(u5_mult_82_n6982), .A2(u5_mult_82_net65519), 
        .ZN(u5_mult_82_ab_34__52_) );
  NOR2_X2 u5_mult_82_U2007 ( .A1(u5_mult_82_n6760), .A2(u5_mult_82_n6706), 
        .ZN(u5_mult_82_ab_35__51_) );
  NOR2_X1 u5_mult_82_U2006 ( .A1(u5_mult_82_n6816), .A2(u5_mult_82_n6686), 
        .ZN(u5_mult_82_ab_31__42_) );
  NOR2_X2 u5_mult_82_U2005 ( .A1(u5_mult_82_n6827), .A2(u5_mult_82_n6677), 
        .ZN(u5_mult_82_ab_30__40_) );
  NOR2_X2 u5_mult_82_U2004 ( .A1(u5_mult_82_net64885), .A2(u5_mult_82_n6601), 
        .ZN(u5_mult_82_ab_17__34_) );
  NOR2_X2 u5_mult_82_U2003 ( .A1(u5_mult_82_n6833), .A2(u5_mult_82_net66035), 
        .ZN(u5_mult_82_ab_5__39_) );
  NOR2_X1 u5_mult_82_U2002 ( .A1(u5_mult_82_n6833), .A2(u5_mult_82_n6550), 
        .ZN(u5_mult_82_ab_10__39_) );
  NOR2_X2 u5_mult_82_U2001 ( .A1(u5_mult_82_net64959), .A2(u5_mult_82_n6557), 
        .ZN(u5_mult_82_ab_11__38_) );
  NOR2_X2 u5_mult_82_U2000 ( .A1(u5_mult_82_n6906), .A2(u5_mult_82_n6545), 
        .ZN(u5_mult_82_ab_9__20_) );
  NOR2_X1 u5_mult_82_U1999 ( .A1(u5_mult_82_n6893), .A2(u5_mult_82_net66019), 
        .ZN(u5_mult_82_ab_6__24_) );
  INV_X4 u5_mult_82_U1998 ( .A(u5_mult_82_ab_4__35_), .ZN(u5_mult_82_net85316)
         );
  NAND3_X2 u5_mult_82_U1997 ( .A1(u5_mult_82_n973), .A2(u5_mult_82_n974), .A3(
        u5_mult_82_n975), .ZN(u5_mult_82_CARRYB_3__33_) );
  NOR2_X2 u5_mult_82_U1996 ( .A1(u5_mult_82_n6923), .A2(u5_mult_82_net66091), 
        .ZN(u5_mult_82_ab_2__18_) );
  NOR2_X2 u5_mult_82_U1995 ( .A1(u5_mult_82_n6906), .A2(u5_mult_82_net66037), 
        .ZN(u5_mult_82_ab_5__20_) );
  NOR2_X2 u5_mult_82_U1994 ( .A1(u5_mult_82_n6850), .A2(u5_mult_82_n6684), 
        .ZN(u5_mult_82_ab_31__31_) );
  NOR2_X2 u5_mult_82_U1993 ( .A1(u5_mult_82_n6821), .A2(u5_mult_82_n6677), 
        .ZN(u5_mult_82_ab_30__41_) );
  NOR2_X2 u5_mult_82_U1992 ( .A1(u5_mult_82_n6832), .A2(u5_mult_82_n6678), 
        .ZN(u5_mult_82_ab_30__39_) );
  NAND3_X2 u5_mult_82_U1991 ( .A1(u5_mult_82_n5024), .A2(u5_mult_82_n5025), 
        .A3(u5_mult_82_n5026), .ZN(u5_mult_82_CARRYB_16__35_) );
  NOR2_X2 u5_mult_82_U1990 ( .A1(u5_mult_82_n6823), .A2(u5_mult_82_net66033), 
        .ZN(u5_mult_82_ab_5__41_) );
  NOR2_X1 u5_mult_82_U1989 ( .A1(u5_mult_82_n6829), .A2(u5_mult_82_n6552), 
        .ZN(u5_mult_82_ab_10__40_) );
  NOR2_X2 u5_mult_82_U1988 ( .A1(u5_mult_82_n6853), .A2(u5_mult_82_net66089), 
        .ZN(u5_mult_82_ab_2__31_) );
  OAI21_X2 u5_mult_82_U1987 ( .B1(u5_mult_82_n1258), .B2(
        u5_mult_82_CARRYB_1__36_), .A(u5_mult_82_n1260), .ZN(u5_mult_82_n1259)
         );
  NOR2_X2 u5_mult_82_U1986 ( .A1(u5_mult_82_n6832), .A2(u5_mult_82_n6671), 
        .ZN(u5_mult_82_ab_29__39_) );
  NOR2_X2 u5_mult_82_U1985 ( .A1(u5_mult_82_n6773), .A2(u5_mult_82_n6684), 
        .ZN(u5_mult_82_ab_31__49_) );
  NOR2_X2 u5_mult_82_U1984 ( .A1(u5_mult_82_n6767), .A2(u5_mult_82_n6683), 
        .ZN(u5_mult_82_ab_31__50_) );
  NOR2_X1 u5_mult_82_U1983 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6663), 
        .ZN(u5_mult_82_ab_28__38_) );
  NOR2_X2 u5_mult_82_U1982 ( .A1(u5_mult_82_n6828), .A2(u5_mult_82_n6600), 
        .ZN(u5_mult_82_ab_17__40_) );
  NOR2_X2 u5_mult_82_U1981 ( .A1(u5_mult_82_n6813), .A2(u5_mult_82_net66033), 
        .ZN(u5_mult_82_ab_5__43_) );
  NOR2_X2 u5_mult_82_U1980 ( .A1(u5_mult_82_n6818), .A2(u5_mult_82_net66033), 
        .ZN(u5_mult_82_ab_5__42_) );
  NOR2_X2 u5_mult_82_U1979 ( .A1(u5_mult_82_n6877), .A2(u5_mult_82_n6522), 
        .ZN(u5_mult_82_ab_4__27_) );
  INV_X8 u5_mult_82_U1978 ( .A(u5_mult_82_n1378), .ZN(u5_mult_82_net64673) );
  NOR2_X2 u5_mult_82_U1977 ( .A1(u5_mult_82_net64939), .A2(u5_mult_82_n6656), 
        .ZN(u5_mult_82_ab_27__37_) );
  NOR2_X1 u5_mult_82_U1976 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_n6656), 
        .ZN(u5_mult_82_ab_27__36_) );
  NOR2_X2 u5_mult_82_U1975 ( .A1(u5_mult_82_n6829), .A2(u5_mult_82_n6580), 
        .ZN(u5_mult_82_ab_14__40_) );
  NOR2_X2 u5_mult_82_U1974 ( .A1(u5_mult_82_n6823), .A2(u5_mult_82_n6573), 
        .ZN(u5_mult_82_ab_13__41_) );
  NOR2_X2 u5_mult_82_U1973 ( .A1(u5_mult_82_n6892), .A2(u5_mult_82_net66091), 
        .ZN(u5_mult_82_ab_2__24_) );
  NOR2_X1 u5_mult_82_U1972 ( .A1(u5_mult_82_n6851), .A2(u5_mult_82_n6656), 
        .ZN(u5_mult_82_ab_27__31_) );
  NOR2_X1 u5_mult_82_U1971 ( .A1(u5_mult_82_net64883), .A2(u5_mult_82_n6663), 
        .ZN(u5_mult_82_ab_28__34_) );
  NAND3_X2 u5_mult_82_U1970 ( .A1(u5_mult_82_n4932), .A2(u5_mult_82_n4933), 
        .A3(u5_mult_82_n4934), .ZN(u5_mult_82_CARRYB_27__35_) );
  NOR2_X2 u5_mult_82_U1969 ( .A1(u5_mult_82_n6779), .A2(u5_mult_82_n6655), 
        .ZN(u5_mult_82_ab_27__48_) );
  NOR2_X1 u5_mult_82_U1968 ( .A1(u5_mult_82_n6817), .A2(u5_mult_82_net65677), 
        .ZN(u5_mult_82_ab_25__42_) );
  INV_X4 u5_mult_82_U1967 ( .A(u5_mult_82_ab_25__43_), .ZN(u5_mult_82_n1430)
         );
  NOR2_X2 u5_mult_82_U1966 ( .A1(u5_mult_82_n6805), .A2(u5_mult_82_net65677), 
        .ZN(u5_mult_82_ab_25__44_) );
  NOR2_X1 u5_mult_82_U1965 ( .A1(u5_mult_82_n6785), .A2(u5_mult_82_n6652), 
        .ZN(u5_mult_82_ab_26__47_) );
  NOR2_X2 u5_mult_82_U1964 ( .A1(u5_mult_82_n6768), .A2(u5_mult_82_n6648), 
        .ZN(u5_mult_82_ab_26__50_) );
  INV_X4 u5_mult_82_U1963 ( .A(u5_mult_82_ab_24__47_), .ZN(u5_mult_82_n1633)
         );
  NOR2_X2 u5_mult_82_U1962 ( .A1(u5_mult_82_n6798), .A2(u5_mult_82_net65677), 
        .ZN(u5_mult_82_ab_25__45_) );
  NOR2_X1 u5_mult_82_U1961 ( .A1(u5_mult_82_n6792), .A2(u5_mult_82_net65717), 
        .ZN(u5_mult_82_ab_23__46_) );
  NOR2_X2 u5_mult_82_U1960 ( .A1(u5_mult_82_n6792), .A2(u5_mult_82_n6643), 
        .ZN(u5_mult_82_ab_24__46_) );
  NOR2_X2 u5_mult_82_U1959 ( .A1(u5_mult_82_n6799), .A2(u5_mult_82_n6520), 
        .ZN(u5_mult_82_ab_4__45_) );
  INV_X4 u5_mult_82_U1958 ( .A(u5_mult_82_ab_25__34_), .ZN(u5_mult_82_n3746)
         );
  NOR2_X2 u5_mult_82_U1957 ( .A1(u5_mult_82_n6761), .A2(u5_mult_82_n6648), 
        .ZN(u5_mult_82_ab_26__51_) );
  NOR2_X2 u5_mult_82_U1956 ( .A1(u5_mult_82_n6828), .A2(u5_mult_82_net65713), 
        .ZN(u5_mult_82_ab_23__40_) );
  INV_X4 u5_mult_82_U1955 ( .A(u5_mult_82_ab_9__42_), .ZN(u5_mult_82_n2361) );
  NOR2_X2 u5_mult_82_U1954 ( .A1(u5_mult_82_n6813), .A2(u5_mult_82_n6537), 
        .ZN(u5_mult_82_ab_8__43_) );
  NOR2_X2 u5_mult_82_U1953 ( .A1(u5_mult_82_n6793), .A2(u5_mult_82_n6537), 
        .ZN(u5_mult_82_ab_8__46_) );
  INV_X4 u5_mult_82_U1952 ( .A(u5_mult_82_ab_21__46_), .ZN(u5_mult_82_n2711)
         );
  NAND2_X1 u5_mult_82_U1951 ( .A1(u5_mult_82_ab_19__46_), .A2(
        u5_mult_82_CARRYB_18__46_), .ZN(u5_mult_82_n2455) );
  INV_X2 u5_mult_82_U1950 ( .A(u5_mult_82_ab_9__47_), .ZN(u5_mult_82_n3508) );
  NOR2_X2 u5_mult_82_U1949 ( .A1(u5_mult_82_n6761), .A2(u5_mult_82_n6620), 
        .ZN(u5_mult_82_ab_20__51_) );
  NOR2_X1 u5_mult_82_U1948 ( .A1(u5_mult_82_n6822), .A2(u5_mult_82_n6615), 
        .ZN(u5_mult_82_ab_19__41_) );
  NOR2_X2 u5_mult_82_U1947 ( .A1(u5_mult_82_n6817), .A2(u5_mult_82_n6615), 
        .ZN(u5_mult_82_ab_19__42_) );
  NOR2_X2 u5_mult_82_U1946 ( .A1(u5_mult_82_n6774), .A2(u5_mult_82_n6600), 
        .ZN(u5_mult_82_ab_17__49_) );
  NOR2_X2 u5_mult_82_U1945 ( .A1(u5_mult_82_n6780), .A2(u5_mult_82_n6520), 
        .ZN(u5_mult_82_ab_4__48_) );
  NOR2_X2 u5_mult_82_U1944 ( .A1(u5_mult_82_n6786), .A2(u5_mult_82_n6552), 
        .ZN(u5_mult_82_ab_10__47_) );
  NOR2_X2 u5_mult_82_U1943 ( .A1(u5_mult_82_n6769), .A2(u5_mult_82_n6520), 
        .ZN(u5_mult_82_ab_4__50_) );
  INV_X4 u5_mult_82_U1942 ( .A(u5_mult_82_ab_18__46_), .ZN(u5_mult_82_n5654)
         );
  INV_X4 u5_mult_82_U1941 ( .A(u5_mult_82_ab_14__49_), .ZN(u5_mult_82_n1766)
         );
  NOR2_X1 u5_mult_82_U1940 ( .A1(u5_mult_82_n6793), .A2(u5_mult_82_n6580), 
        .ZN(u5_mult_82_ab_14__46_) );
  NOR2_X2 u5_mult_82_U1939 ( .A1(u5_mult_82_n6775), .A2(u5_mult_82_n6558), 
        .ZN(u5_mult_82_ab_11__49_) );
  NOR2_X2 u5_mult_82_U1938 ( .A1(u5_mult_82_n6989), .A2(u5_mult_82_net66041), 
        .ZN(u5_mult_82_ab_5__0_) );
  NOR2_X1 u5_mult_82_U1937 ( .A1(u5_mult_82_n6989), .A2(u5_mult_82_n6553), 
        .ZN(u5_mult_82_ab_10__0_) );
  NOR2_X2 u5_mult_82_U1936 ( .A1(u5_mult_82_n6988), .A2(u5_mult_82_n6589), 
        .ZN(u5_mult_82_ab_15__0_) );
  NOR2_X2 u5_mult_82_U1935 ( .A1(u5_mult_82_n6988), .A2(u5_mult_82_n6624), 
        .ZN(u5_mult_82_ab_20__0_) );
  NOR2_X1 u5_mult_82_U1934 ( .A1(u5_mult_82_n6988), .A2(u5_mult_82_net65681), 
        .ZN(u5_mult_82_ab_25__0_) );
  NOR2_X2 u5_mult_82_U1933 ( .A1(u5_mult_82_n6987), .A2(u5_mult_82_n6681), 
        .ZN(u5_mult_82_ab_30__0_) );
  NOR2_X2 u5_mult_82_U1932 ( .A1(u5_mult_82_n6987), .A2(u5_mult_82_n6710), 
        .ZN(u5_mult_82_ab_35__0_) );
  NOR2_X2 u5_mult_82_U1931 ( .A1(u5_mult_82_n6884), .A2(u5_mult_82_net65371), 
        .ZN(u5_mult_82_ab_42__25_) );
  NOR2_X2 u5_mult_82_U1930 ( .A1(u5_mult_82_n6969), .A2(u5_mult_82_net66041), 
        .ZN(u5_mult_82_ab_5__1_) );
  NOR2_X1 u5_mult_82_U1929 ( .A1(u5_mult_82_n6969), .A2(u5_mult_82_n6553), 
        .ZN(u5_mult_82_ab_10__1_) );
  INV_X16 u5_mult_82_U1928 ( .A(u5_mult_82_n6569), .ZN(u5_mult_82_n6568) );
  NOR2_X2 u5_mult_82_U1927 ( .A1(u5_mult_82_n6969), .A2(u5_mult_82_n6589), 
        .ZN(u5_mult_82_ab_15__1_) );
  INV_X16 u5_mult_82_U1926 ( .A(u5_mult_82_n6605), .ZN(u5_mult_82_n6604) );
  NOR2_X2 u5_mult_82_U1925 ( .A1(u5_mult_82_n6968), .A2(u5_mult_82_n6624), 
        .ZN(u5_mult_82_ab_20__1_) );
  INV_X16 u5_mult_82_U1924 ( .A(u5_mult_82_n6639), .ZN(u5_mult_82_n6638) );
  NOR2_X1 u5_mult_82_U1923 ( .A1(u5_mult_82_n6968), .A2(u5_mult_82_net65681), 
        .ZN(u5_mult_82_ab_25__1_) );
  NOR2_X2 u5_mult_82_U1922 ( .A1(u5_mult_82_n6967), .A2(u5_mult_82_n6681), 
        .ZN(u5_mult_82_ab_30__1_) );
  NOR2_X2 u5_mult_82_U1921 ( .A1(u5_mult_82_n6967), .A2(u5_mult_82_n6710), 
        .ZN(u5_mult_82_ab_35__1_) );
  NOR2_X1 u5_mult_82_U1920 ( .A1(u5_mult_82_n6967), .A2(u5_mult_82_net65229), 
        .ZN(u5_mult_82_ab_50__1_) );
  NOR2_X2 u5_mult_82_U1919 ( .A1(u5_mult_82_n6914), .A2(u5_mult_82_n6657), 
        .ZN(u5_mult_82_ab_27__19_) );
  NOR2_X2 u5_mult_82_U1918 ( .A1(u5_mult_82_n6962), .A2(u5_mult_82_net66041), 
        .ZN(u5_mult_82_ab_5__2_) );
  NOR2_X1 u5_mult_82_U1917 ( .A1(u5_mult_82_n6962), .A2(u5_mult_82_n6553), 
        .ZN(u5_mult_82_ab_10__2_) );
  NOR2_X2 u5_mult_82_U1916 ( .A1(u5_mult_82_n6962), .A2(u5_mult_82_n6589), 
        .ZN(u5_mult_82_ab_15__2_) );
  NOR2_X2 u5_mult_82_U1915 ( .A1(u5_mult_82_n6961), .A2(u5_mult_82_n6624), 
        .ZN(u5_mult_82_ab_20__2_) );
  NOR2_X1 u5_mult_82_U1914 ( .A1(u5_mult_82_n6961), .A2(u5_mult_82_net65681), 
        .ZN(u5_mult_82_ab_25__2_) );
  NOR2_X2 u5_mult_82_U1913 ( .A1(u5_mult_82_n6960), .A2(u5_mult_82_n6681), 
        .ZN(u5_mult_82_ab_30__2_) );
  NOR2_X2 u5_mult_82_U1912 ( .A1(u5_mult_82_n6960), .A2(u5_mult_82_n6710), 
        .ZN(u5_mult_82_ab_35__2_) );
  NOR2_X1 u5_mult_82_U1911 ( .A1(u5_mult_82_n6953), .A2(u5_mult_82_n6730), 
        .ZN(u5_mult_82_ab_39__3_) );
  NOR2_X2 u5_mult_82_U1910 ( .A1(u5_mult_82_n6905), .A2(u5_mult_82_n6657), 
        .ZN(u5_mult_82_ab_27__20_) );
  NOR2_X2 u5_mult_82_U1909 ( .A1(u5_mult_82_net64669), .A2(u5_mult_82_n6657), 
        .ZN(u5_mult_82_ab_27__22_) );
  INV_X8 u5_mult_82_U1908 ( .A(u5_mult_82_n6964), .ZN(u5_mult_82_n6963) );
  NOR2_X2 u5_mult_82_U1907 ( .A1(u5_mult_82_n6955), .A2(u5_mult_82_net66041), 
        .ZN(u5_mult_82_ab_5__3_) );
  NOR2_X1 u5_mult_82_U1906 ( .A1(u5_mult_82_n6955), .A2(u5_mult_82_n6553), 
        .ZN(u5_mult_82_ab_10__3_) );
  NOR2_X2 u5_mult_82_U1905 ( .A1(u5_mult_82_n6955), .A2(u5_mult_82_n6589), 
        .ZN(u5_mult_82_ab_15__3_) );
  NOR2_X2 u5_mult_82_U1904 ( .A1(u5_mult_82_n6953), .A2(u5_mult_82_n6681), 
        .ZN(u5_mult_82_ab_30__3_) );
  NOR2_X1 u5_mult_82_U1903 ( .A1(u5_mult_82_n6946), .A2(u5_mult_82_n6755), 
        .ZN(u5_mult_82_ab_49__4_) );
  INV_X4 u5_mult_82_U1902 ( .A(u5_mult_82_n6978), .ZN(u5_mult_82_n6976) );
  NOR2_X2 u5_mult_82_U1901 ( .A1(u5_mult_82_n6913), .A2(u5_mult_82_n6715), 
        .ZN(u5_mult_82_ab_36__19_) );
  INV_X16 u5_mult_82_U1900 ( .A(u5_mult_82_n6894), .ZN(u5_mult_82_n6901) );
  INV_X8 u5_mult_82_U1899 ( .A(u5_mult_82_n6957), .ZN(u5_mult_82_n6956) );
  NOR2_X2 u5_mult_82_U1898 ( .A1(u5_mult_82_n6948), .A2(u5_mult_82_net66039), 
        .ZN(u5_mult_82_ab_5__4_) );
  NOR2_X1 u5_mult_82_U1897 ( .A1(u5_mult_82_n6948), .A2(u5_mult_82_n6552), 
        .ZN(u5_mult_82_ab_10__4_) );
  NOR2_X2 u5_mult_82_U1896 ( .A1(u5_mult_82_n6948), .A2(u5_mult_82_n6588), 
        .ZN(u5_mult_82_ab_15__4_) );
  NOR2_X1 u5_mult_82_U1895 ( .A1(u5_mult_82_n6946), .A2(u5_mult_82_n6729), 
        .ZN(u5_mult_82_ab_39__4_) );
  INV_X4 u5_mult_82_U1894 ( .A(u5_mult_82_ab_45__4_), .ZN(u5_mult_82_n5856) );
  NOR2_X1 u5_mult_82_U1893 ( .A1(u5_mult_82_net64361), .A2(u5_mult_82_net65189), .ZN(u5_mult_82_ab_51__5_) );
  NOR2_X1 u5_mult_82_U1892 ( .A1(u5_mult_82_n6867), .A2(u5_mult_82_net65225), 
        .ZN(u5_mult_82_ab_50__28_) );
  NOR2_X1 u5_mult_82_U1891 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_net65225), .ZN(u5_mult_82_ab_50__36_) );
  NOR2_X1 u5_mult_82_U1890 ( .A1(u5_mult_82_n6983), .A2(u5_mult_82_n6749), 
        .ZN(u5_mult_82_ab_48__52_) );
  NOR2_X2 u5_mult_82_U1889 ( .A1(u5_mult_82_n6759), .A2(u5_mult_82_n6752), 
        .ZN(u5_mult_82_ab_49__51_) );
  NOR2_X2 u5_mult_82_U1888 ( .A1(u5_mult_82_n6875), .A2(u5_mult_82_n6721), 
        .ZN(u5_mult_82_ab_37__27_) );
  NOR2_X2 u5_mult_82_U1887 ( .A1(u5_mult_82_n6868), .A2(u5_mult_82_n6720), 
        .ZN(u5_mult_82_ab_37__28_) );
  NOR2_X2 u5_mult_82_U1886 ( .A1(u5_mult_82_net64223), .A2(u5_mult_82_net64373), .ZN(u5_mult_82_ab_0__5_) );
  NOR2_X2 u5_mult_82_U1885 ( .A1(u5_mult_82_net64365), .A2(u5_mult_82_net66039), .ZN(u5_mult_82_ab_5__5_) );
  NOR2_X1 u5_mult_82_U1884 ( .A1(u5_mult_82_net64365), .A2(u5_mult_82_n6552), 
        .ZN(u5_mult_82_ab_10__5_) );
  NOR2_X2 u5_mult_82_U1883 ( .A1(u5_mult_82_net64365), .A2(u5_mult_82_n6588), 
        .ZN(u5_mult_82_ab_15__5_) );
  NOR2_X2 u5_mult_82_U1882 ( .A1(u5_mult_82_net64381), .A2(u5_mult_82_n6623), 
        .ZN(u5_mult_82_ab_20__6_) );
  INV_X4 u5_mult_82_U1881 ( .A(u5_mult_82_n1373), .ZN(u5_mult_82_net64459) );
  INV_X4 u5_mult_82_U1880 ( .A(u5_mult_82_ab_49__24_), .ZN(u5_mult_82_n4485)
         );
  NOR2_X1 u5_mult_82_U1879 ( .A1(u5_mult_82_n6856), .A2(u5_mult_82_net65225), 
        .ZN(u5_mult_82_ab_50__30_) );
  NOR2_X1 u5_mult_82_U1878 ( .A1(u5_mult_82_n6849), .A2(u5_mult_82_net65225), 
        .ZN(u5_mult_82_ab_50__31_) );
  INV_X4 u5_mult_82_U1877 ( .A(u5_mult_82_net65197), .ZN(u5_mult_82_net65193)
         );
  NOR2_X1 u5_mult_82_U1876 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_net65225), .ZN(u5_mult_82_ab_50__38_) );
  NOR2_X1 u5_mult_82_U1875 ( .A1(u5_mult_82_n6777), .A2(u5_mult_82_net65223), 
        .ZN(u5_mult_82_ab_50__48_) );
  NOR2_X1 u5_mult_82_U1874 ( .A1(u5_mult_82_n6772), .A2(u5_mult_82_net65223), 
        .ZN(u5_mult_82_ab_50__49_) );
  NOR2_X1 u5_mult_82_U1873 ( .A1(u5_mult_82_n6826), .A2(u5_mult_82_net65223), 
        .ZN(u5_mult_82_ab_50__40_) );
  NOR2_X2 u5_mult_82_U1872 ( .A1(u5_mult_82_n6874), .A2(u5_mult_82_n6749), 
        .ZN(u5_mult_82_ab_48__27_) );
  NOR2_X2 u5_mult_82_U1871 ( .A1(u5_mult_82_n6920), .A2(u5_mult_82_net65515), 
        .ZN(u5_mult_82_ab_34__18_) );
  NOR2_X1 u5_mult_82_U1870 ( .A1(u5_mult_82_n6927), .A2(u5_mult_82_net65515), 
        .ZN(u5_mult_82_ab_34__17_) );
  NOR2_X2 u5_mult_82_U1869 ( .A1(u5_mult_82_net64685), .A2(u5_mult_82_net65515), .ZN(u5_mult_82_ab_34__23_) );
  NOR2_X1 u5_mult_82_U1868 ( .A1(u5_mult_82_net64559), .A2(u5_mult_82_net65515), .ZN(u5_mult_82_ab_34__16_) );
  NOR2_X1 u5_mult_82_U1867 ( .A1(u5_mult_82_n6905), .A2(u5_mult_82_net65713), 
        .ZN(u5_mult_82_ab_23__20_) );
  INV_X4 u5_mult_82_U1866 ( .A(u5_mult_82_net64369), .ZN(u5_mult_82_net64367)
         );
  NOR2_X2 u5_mult_82_U1865 ( .A1(u5_mult_82_net64383), .A2(u5_mult_82_net66039), .ZN(u5_mult_82_ab_5__6_) );
  NOR2_X1 u5_mult_82_U1864 ( .A1(u5_mult_82_net64383), .A2(u5_mult_82_n6552), 
        .ZN(u5_mult_82_ab_10__6_) );
  NOR2_X2 u5_mult_82_U1863 ( .A1(u5_mult_82_net64383), .A2(u5_mult_82_n6588), 
        .ZN(u5_mult_82_ab_15__6_) );
  NOR2_X2 u5_mult_82_U1862 ( .A1(u5_mult_82_n6941), .A2(u5_mult_82_n6623), 
        .ZN(u5_mult_82_ab_20__7_) );
  NOR2_X2 u5_mult_82_U1861 ( .A1(u5_mult_82_net64417), .A2(u5_mult_82_n6623), 
        .ZN(u5_mult_82_ab_20__8_) );
  NOR2_X1 u5_mult_82_U1860 ( .A1(u5_mult_82_n6940), .A2(u5_mult_82_n6665), 
        .ZN(u5_mult_82_ab_28__7_) );
  NOR2_X1 u5_mult_82_U1859 ( .A1(u5_mult_82_net64415), .A2(u5_mult_82_n6673), 
        .ZN(u5_mult_82_ab_29__8_) );
  INV_X4 u5_mult_82_U1858 ( .A(u5_mult_82_ab_34__8_), .ZN(u5_mult_82_n2293) );
  INV_X4 u5_mult_82_U1857 ( .A(u5_mult_82_ab_33__9_), .ZN(u5_mult_82_n2324) );
  NOR2_X1 u5_mult_82_U1856 ( .A1(u5_mult_82_net64361), .A2(u5_mult_82_net65373), .ZN(u5_mult_82_ab_42__5_) );
  INV_X4 u5_mult_82_U1855 ( .A(u5_mult_82_ab_48__12_), .ZN(u5_mult_82_n5201)
         );
  INV_X4 u5_mult_82_U1854 ( .A(u5_mult_82_ab_49__11_), .ZN(u5_mult_82_n3061)
         );
  NAND2_X2 u5_mult_82_U1853 ( .A1(u5_mult_82_CARRYB_48__14_), .A2(
        u5_mult_82_n1661), .ZN(u5_mult_82_n5826) );
  NAND3_X2 u5_mult_82_U1852 ( .A1(u5_mult_82_n5826), .A2(u5_mult_82_n5825), 
        .A3(u5_mult_82_n5824), .ZN(u5_mult_82_CARRYB_49__14_) );
  NOR2_X1 u5_mult_82_U1851 ( .A1(u5_mult_82_n6784), .A2(u5_mult_82_n6752), 
        .ZN(u5_mult_82_ab_49__47_) );
  NOR2_X1 u5_mult_82_U1850 ( .A1(u5_mult_82_n6797), .A2(u5_mult_82_n6752), 
        .ZN(u5_mult_82_ab_49__45_) );
  NOR2_X2 u5_mult_82_U1849 ( .A1(u5_mult_82_n6803), .A2(u5_mult_82_n6752), 
        .ZN(u5_mult_82_ab_49__44_) );
  NOR2_X1 u5_mult_82_U1848 ( .A1(u5_mult_82_n6816), .A2(u5_mult_82_n6752), 
        .ZN(u5_mult_82_ab_49__42_) );
  INV_X4 u5_mult_82_U1847 ( .A(u5_mult_82_ab_34__32_), .ZN(u5_mult_82_n1947)
         );
  NAND3_X2 u5_mult_82_U1846 ( .A1(u5_mult_82_n3615), .A2(u5_mult_82_n3616), 
        .A3(u5_mult_82_n3617), .ZN(u5_mult_82_CARRYB_21__23_) );
  INV_X8 u5_mult_82_U1845 ( .A(u5_mult_82_net64387), .ZN(u5_mult_82_net64385)
         );
  NOR2_X2 u5_mult_82_U1844 ( .A1(u5_mult_82_n6942), .A2(u5_mult_82_net66039), 
        .ZN(u5_mult_82_ab_5__7_) );
  NOR2_X1 u5_mult_82_U1843 ( .A1(u5_mult_82_n6942), .A2(u5_mult_82_n6552), 
        .ZN(u5_mult_82_ab_10__7_) );
  NOR2_X2 u5_mult_82_U1842 ( .A1(u5_mult_82_n6942), .A2(u5_mult_82_n6588), 
        .ZN(u5_mult_82_ab_15__7_) );
  NOR2_X2 u5_mult_82_U1841 ( .A1(u5_mult_82_net64419), .A2(u5_mult_82_n6588), 
        .ZN(u5_mult_82_ab_15__8_) );
  NOR2_X2 u5_mult_82_U1840 ( .A1(u5_mult_82_n6875), .A2(u5_mult_82_n6700), 
        .ZN(u5_mult_82_ab_33__27_) );
  NAND3_X2 u5_mult_82_U1839 ( .A1(u5_mult_82_n5412), .A2(u5_mult_82_n5413), 
        .A3(u5_mult_82_n5414), .ZN(u5_mult_82_CARRYB_32__20_) );
  NOR2_X2 u5_mult_82_U1838 ( .A1(u5_mult_82_n6869), .A2(u5_mult_82_n6635), 
        .ZN(u5_mult_82_ab_22__28_) );
  NOR2_X2 u5_mult_82_U1837 ( .A1(u5_mult_82_net64419), .A2(u5_mult_82_net66039), .ZN(u5_mult_82_ab_5__8_) );
  NOR2_X1 u5_mult_82_U1836 ( .A1(u5_mult_82_net64419), .A2(u5_mult_82_n6552), 
        .ZN(u5_mult_82_ab_10__8_) );
  NOR2_X2 u5_mult_82_U1835 ( .A1(u5_mult_82_net64437), .A2(u5_mult_82_n6588), 
        .ZN(u5_mult_82_ab_15__9_) );
  NOR2_X2 u5_mult_82_U1834 ( .A1(u5_mult_82_net64435), .A2(u5_mult_82_n6623), 
        .ZN(u5_mult_82_ab_20__9_) );
  NOR2_X2 u5_mult_82_U1833 ( .A1(u5_mult_82_n6895), .A2(u5_mult_82_net65321), 
        .ZN(u5_mult_82_ab_45__21_) );
  NOR2_X2 u5_mult_82_U1832 ( .A1(u5_mult_82_n6874), .A2(u5_mult_82_n6735), 
        .ZN(u5_mult_82_ab_44__27_) );
  INV_X16 u5_mult_82_U1831 ( .A(u5_mult_82_n1292), .ZN(u5_mult_82_net65313) );
  NOR2_X1 u5_mult_82_U1830 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_net65315), .ZN(u5_mult_82_ab_45__38_) );
  NOR2_X1 u5_mult_82_U1829 ( .A1(u5_mult_82_net64883), .A2(u5_mult_82_n6699), 
        .ZN(u5_mult_82_ab_33__34_) );
  NOR2_X2 u5_mult_82_U1828 ( .A1(u5_mult_82_net64669), .A2(u5_mult_82_n6609), 
        .ZN(u5_mult_82_ab_18__22_) );
  NOR2_X2 u5_mult_82_U1827 ( .A1(u5_mult_82_n6897), .A2(u5_mult_82_n6609), 
        .ZN(u5_mult_82_ab_18__21_) );
  NOR2_X2 u5_mult_82_U1826 ( .A1(u5_mult_82_net64437), .A2(u5_mult_82_net66039), .ZN(u5_mult_82_ab_5__9_) );
  NOR2_X1 u5_mult_82_U1825 ( .A1(u5_mult_82_net64437), .A2(u5_mult_82_n6552), 
        .ZN(u5_mult_82_ab_10__9_) );
  NOR2_X2 u5_mult_82_U1824 ( .A1(u5_mult_82_net64453), .A2(u5_mult_82_n6623), 
        .ZN(u5_mult_82_ab_20__10_) );
  INV_X4 u5_mult_82_U1823 ( .A(u5_mult_82_ab_25__12_), .ZN(u5_mult_82_n632) );
  NAND3_X2 u5_mult_82_U1822 ( .A1(u5_mult_82_n5306), .A2(u5_mult_82_n5307), 
        .A3(u5_mult_82_n5308), .ZN(u5_mult_82_CARRYB_30__11_) );
  NOR2_X1 u5_mult_82_U1821 ( .A1(u5_mult_82_net64469), .A2(u5_mult_82_n6686), 
        .ZN(u5_mult_82_ab_31__11_) );
  NOR2_X1 u5_mult_82_U1820 ( .A1(u5_mult_82_net64451), .A2(u5_mult_82_n6709), 
        .ZN(u5_mult_82_ab_35__10_) );
  INV_X4 u5_mult_82_U1819 ( .A(u5_mult_82_ab_39__8_), .ZN(u5_mult_82_n4702) );
  NOR2_X1 u5_mult_82_U1818 ( .A1(u5_mult_82_n6927), .A2(u5_mult_82_n6735), 
        .ZN(u5_mult_82_ab_44__17_) );
  INV_X1 u5_mult_82_U1817 ( .A(u5_mult_82_ab_46__19_), .ZN(u5_mult_82_n1420)
         );
  NOR2_X2 u5_mult_82_U1816 ( .A1(u5_mult_82_n6879), .A2(u5_mult_82_net65353), 
        .ZN(u5_mult_82_ab_43__26_) );
  NOR2_X2 u5_mult_82_U1815 ( .A1(u5_mult_82_n6861), .A2(u5_mult_82_net65351), 
        .ZN(u5_mult_82_ab_43__29_) );
  NOR2_X1 u5_mult_82_U1814 ( .A1(u5_mult_82_n6816), .A2(u5_mult_82_net65371), 
        .ZN(u5_mult_82_ab_42__42_) );
  NOR2_X1 u5_mult_82_U1813 ( .A1(u5_mult_82_n6983), .A2(u5_mult_82_net65353), 
        .ZN(u5_mult_82_ab_43__52_) );
  NOR2_X2 u5_mult_82_U1812 ( .A1(u5_mult_82_n6759), .A2(u5_mult_82_n6733), 
        .ZN(u5_mult_82_ab_44__51_) );
  INV_X2 u5_mult_82_U1811 ( .A(u5_mult_82_CARRYB_32__31_), .ZN(
        u5_mult_82_n3584) );
  INV_X4 u5_mult_82_U1810 ( .A(u5_mult_82_ab_29__26_), .ZN(u5_mult_82_n4102)
         );
  INV_X4 u5_mult_82_U1809 ( .A(u5_mult_82_n1313), .ZN(u5_mult_82_n1314) );
  NOR2_X2 u5_mult_82_U1808 ( .A1(u5_mult_82_n6914), .A2(u5_mult_82_n6609), 
        .ZN(u5_mult_82_ab_18__19_) );
  NOR2_X2 u5_mult_82_U1807 ( .A1(u5_mult_82_n6877), .A2(u5_mult_82_n6587), 
        .ZN(u5_mult_82_ab_15__27_) );
  NOR2_X1 u5_mult_82_U1806 ( .A1(u5_mult_82_net64455), .A2(u5_mult_82_net66039), .ZN(u5_mult_82_ab_5__10_) );
  NOR2_X1 u5_mult_82_U1805 ( .A1(u5_mult_82_net64455), .A2(u5_mult_82_n6552), 
        .ZN(u5_mult_82_ab_10__10_) );
  NOR2_X1 u5_mult_82_U1804 ( .A1(u5_mult_82_net64471), .A2(u5_mult_82_n6644), 
        .ZN(u5_mult_82_ab_24__11_) );
  INV_X4 u5_mult_82_U1803 ( .A(u5_mult_82_ab_25__14_), .ZN(u5_mult_82_n2131)
         );
  INV_X4 u5_mult_82_U1802 ( .A(u5_mult_82_ab_42__17_), .ZN(u5_mult_82_n4300)
         );
  NOR2_X2 u5_mult_82_U1801 ( .A1(u5_mult_82_n6903), .A2(u5_mult_82_net65371), 
        .ZN(u5_mult_82_ab_42__20_) );
  NOR2_X1 u5_mult_82_U1800 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_net65369), .ZN(u5_mult_82_ab_42__36_) );
  NOR2_X2 u5_mult_82_U1799 ( .A1(u5_mult_82_net64935), .A2(u5_mult_82_net65351), .ZN(u5_mult_82_ab_43__37_) );
  NOR2_X2 u5_mult_82_U1798 ( .A1(u5_mult_82_n6810), .A2(u5_mult_82_net65371), 
        .ZN(u5_mult_82_ab_42__43_) );
  NAND3_X2 u5_mult_82_U1797 ( .A1(u5_mult_82_n1069), .A2(u5_mult_82_n1070), 
        .A3(u5_mult_82_n1071), .ZN(u5_mult_82_CARRYB_41__34_) );
  NOR2_X2 u5_mult_82_U1796 ( .A1(u5_mult_82_net64901), .A2(u5_mult_82_net65387), .ZN(u5_mult_82_ab_41__35_) );
  NOR2_X2 u5_mult_82_U1795 ( .A1(u5_mult_82_n6839), .A2(u5_mult_82_net65405), 
        .ZN(u5_mult_82_ab_40__33_) );
  NOR2_X2 u5_mult_82_U1794 ( .A1(u5_mult_82_n6869), .A2(u5_mult_82_n6656), 
        .ZN(u5_mult_82_ab_27__28_) );
  NOR2_X2 u5_mult_82_U1793 ( .A1(u5_mult_82_n6845), .A2(u5_mult_82_n6586), 
        .ZN(u5_mult_82_ab_15__32_) );
  NOR2_X2 u5_mult_82_U1792 ( .A1(u5_mult_82_n6858), .A2(u5_mult_82_n6594), 
        .ZN(u5_mult_82_ab_16__30_) );
  NOR2_X2 u5_mult_82_U1791 ( .A1(u5_mult_82_net64223), .A2(u5_mult_82_n1319), 
        .ZN(u5_mult_82_ab_0__11_) );
  NOR2_X2 u5_mult_82_U1790 ( .A1(u5_mult_82_net64473), .A2(u5_mult_82_net66039), .ZN(u5_mult_82_ab_5__11_) );
  NOR2_X1 u5_mult_82_U1789 ( .A1(u5_mult_82_net64473), .A2(u5_mult_82_n6552), 
        .ZN(u5_mult_82_ab_10__11_) );
  NOR2_X1 u5_mult_82_U1788 ( .A1(u5_mult_82_net64491), .A2(u5_mult_82_n6573), 
        .ZN(u5_mult_82_ab_13__12_) );
  NOR2_X1 u5_mult_82_U1787 ( .A1(u5_mult_82_net64509), .A2(u5_mult_82_n6580), 
        .ZN(u5_mult_82_ab_14__13_) );
  NOR2_X2 u5_mult_82_U1786 ( .A1(u5_mult_82_net64471), .A2(u5_mult_82_n6623), 
        .ZN(u5_mult_82_ab_20__11_) );
  NOR2_X2 u5_mult_82_U1785 ( .A1(u5_mult_82_n6822), .A2(u5_mult_82_net65403), 
        .ZN(u5_mult_82_ab_40__41_) );
  NOR2_X1 u5_mult_82_U1784 ( .A1(u5_mult_82_n6772), .A2(u5_mult_82_n6737), 
        .ZN(u5_mult_82_ab_44__49_) );
  NOR2_X2 u5_mult_82_U1783 ( .A1(u5_mult_82_n6777), .A2(u5_mult_82_n6733), 
        .ZN(u5_mult_82_ab_44__48_) );
  NOR2_X1 u5_mult_82_U1782 ( .A1(u5_mult_82_n6784), .A2(u5_mult_82_n6733), 
        .ZN(u5_mult_82_ab_44__47_) );
  NOR2_X1 u5_mult_82_U1781 ( .A1(u5_mult_82_n6797), .A2(u5_mult_82_n6734), 
        .ZN(u5_mult_82_ab_44__45_) );
  NOR2_X1 u5_mult_82_U1780 ( .A1(u5_mult_82_n6851), .A2(u5_mult_82_n6649), 
        .ZN(u5_mult_82_ab_26__31_) );
  NAND3_X2 u5_mult_82_U1779 ( .A1(u5_mult_82_n3574), .A2(u5_mult_82_n3575), 
        .A3(u5_mult_82_n3576), .ZN(u5_mult_82_CARRYB_26__17_) );
  NOR2_X2 u5_mult_82_U1778 ( .A1(u5_mult_82_n6928), .A2(u5_mult_82_n6657), 
        .ZN(u5_mult_82_ab_27__17_) );
  INV_X4 u5_mult_82_U1777 ( .A(u5_mult_82_ab_15__33_), .ZN(u5_mult_82_n2011)
         );
  NOR2_X1 u5_mult_82_U1776 ( .A1(u5_mult_82_n6859), .A2(u5_mult_82_n6571), 
        .ZN(u5_mult_82_ab_13__30_) );
  INV_X4 u5_mult_82_U1775 ( .A(u5_mult_82_net64477), .ZN(u5_mult_82_net64475)
         );
  NOR2_X2 u5_mult_82_U1774 ( .A1(u5_mult_82_net64491), .A2(u5_mult_82_net66039), .ZN(u5_mult_82_ab_5__12_) );
  NOR2_X1 u5_mult_82_U1773 ( .A1(u5_mult_82_net64507), .A2(u5_mult_82_n6616), 
        .ZN(u5_mult_82_ab_19__13_) );
  NOR2_X2 u5_mult_82_U1772 ( .A1(u5_mult_82_net64505), .A2(u5_mult_82_n6680), 
        .ZN(u5_mult_82_ab_30__13_) );
  NOR2_X1 u5_mult_82_U1771 ( .A1(u5_mult_82_net64487), .A2(u5_mult_82_n6709), 
        .ZN(u5_mult_82_ab_35__12_) );
  NOR2_X2 u5_mult_82_U1770 ( .A1(u5_mult_82_n6852), .A2(u5_mult_82_n6571), 
        .ZN(u5_mult_82_ab_13__31_) );
  INV_X4 u5_mult_82_U1769 ( .A(u5_mult_82_ab_15__35_), .ZN(u5_mult_82_n1784)
         );
  NOR2_X2 u5_mult_82_U1768 ( .A1(u5_mult_82_net64671), .A2(u5_mult_82_n6566), 
        .ZN(u5_mult_82_ab_12__22_) );
  NOR2_X2 u5_mult_82_U1767 ( .A1(u5_mult_82_n6893), .A2(u5_mult_82_n6566), 
        .ZN(u5_mult_82_ab_12__24_) );
  NOR2_X2 u5_mult_82_U1766 ( .A1(u5_mult_82_net64509), .A2(u5_mult_82_net66039), .ZN(u5_mult_82_ab_5__13_) );
  NOR2_X2 u5_mult_82_U1765 ( .A1(u5_mult_82_n6934), .A2(u5_mult_82_n6623), 
        .ZN(u5_mult_82_ab_20__15_) );
  NOR2_X1 u5_mult_82_U1764 ( .A1(u5_mult_82_n6831), .A2(u5_mult_82_n6649), 
        .ZN(u5_mult_82_ab_26__39_) );
  NAND2_X2 u5_mult_82_U1763 ( .A1(u5_mult_82_ab_26__40_), .A2(u5_mult_82_n2211), .ZN(u5_mult_82_n2213) );
  NOR2_X1 u5_mult_82_U1762 ( .A1(u5_mult_82_n6915), .A2(u5_mult_82_n6579), 
        .ZN(u5_mult_82_ab_14__19_) );
  NOR2_X2 u5_mult_82_U1761 ( .A1(u5_mult_82_net64527), .A2(u5_mult_82_net66039), .ZN(u5_mult_82_ab_5__14_) );
  NOR2_X2 u5_mult_82_U1760 ( .A1(u5_mult_82_n6935), .A2(u5_mult_82_n6537), 
        .ZN(u5_mult_82_ab_8__15_) );
  NOR2_X2 u5_mult_82_U1759 ( .A1(u5_mult_82_net64563), .A2(u5_mult_82_n6536), 
        .ZN(u5_mult_82_ab_8__16_) );
  NOR2_X1 u5_mult_82_U1758 ( .A1(u5_mult_82_net64563), .A2(u5_mult_82_n6579), 
        .ZN(u5_mult_82_ab_14__16_) );
  NOR2_X1 u5_mult_82_U1757 ( .A1(u5_mult_82_n6933), .A2(u5_mult_82_n6701), 
        .ZN(u5_mult_82_ab_33__15_) );
  NOR2_X2 u5_mult_82_U1756 ( .A1(u5_mult_82_n6827), .A2(u5_mult_82_n6713), 
        .ZN(u5_mult_82_ab_36__40_) );
  NOR2_X1 u5_mult_82_U1755 ( .A1(u5_mult_82_n6832), .A2(u5_mult_82_n6714), 
        .ZN(u5_mult_82_ab_36__39_) );
  NOR2_X1 u5_mult_82_U1754 ( .A1(u5_mult_82_n6784), .A2(u5_mult_82_net65443), 
        .ZN(u5_mult_82_ab_38__47_) );
  NOR2_X1 u5_mult_82_U1753 ( .A1(u5_mult_82_n6797), .A2(u5_mult_82_n6721), 
        .ZN(u5_mult_82_ab_37__45_) );
  NOR2_X2 u5_mult_82_U1752 ( .A1(u5_mult_82_n6778), .A2(u5_mult_82_net65447), 
        .ZN(u5_mult_82_ab_38__48_) );
  NOR2_X1 u5_mult_82_U1751 ( .A1(u5_mult_82_n6982), .A2(u5_mult_82_net65447), 
        .ZN(u5_mult_82_ab_38__52_) );
  NOR2_X2 u5_mult_82_U1750 ( .A1(u5_mult_82_n6760), .A2(u5_mult_82_n6726), 
        .ZN(u5_mult_82_ab_39__51_) );
  NAND2_X2 u5_mult_82_U1749 ( .A1(u5_mult_82_ab_25__33_), .A2(u5_mult_82_n3381), .ZN(u5_mult_82_n3383) );
  NAND2_X2 u5_mult_82_U1748 ( .A1(u5_mult_82_n5548), .A2(
        u5_mult_82_CARRYB_24__33_), .ZN(u5_mult_82_n3382) );
  NOR2_X2 u5_mult_82_U1747 ( .A1(u5_mult_82_net64903), .A2(u5_mult_82_net65675), .ZN(u5_mult_82_ab_25__35_) );
  NOR2_X1 u5_mult_82_U1746 ( .A1(u5_mult_82_net64887), .A2(u5_mult_82_n6550), 
        .ZN(u5_mult_82_ab_10__34_) );
  INV_X4 u5_mult_82_U1745 ( .A(u5_mult_82_ab_10__37_), .ZN(u5_mult_82_n2007)
         );
  NAND3_X2 u5_mult_82_U1744 ( .A1(u5_mult_82_n4751), .A2(u5_mult_82_n4750), 
        .A3(u5_mult_82_n4749), .ZN(u5_mult_82_CARRYB_10__36_) );
  NOR2_X1 u5_mult_82_U1743 ( .A1(u5_mult_82_n6840), .A2(u5_mult_82_n6535), 
        .ZN(u5_mult_82_ab_8__33_) );
  NOR2_X1 u5_mult_82_U1742 ( .A1(u5_mult_82_n6845), .A2(u5_mult_82_n6535), 
        .ZN(u5_mult_82_ab_8__32_) );
  NOR2_X1 u5_mult_82_U1741 ( .A1(u5_mult_82_n6852), .A2(u5_mult_82_n6535), 
        .ZN(u5_mult_82_ab_8__31_) );
  NOR2_X2 u5_mult_82_U1740 ( .A1(u5_mult_82_n6929), .A2(u5_mult_82_n6545), 
        .ZN(u5_mult_82_ab_9__17_) );
  NOR2_X2 u5_mult_82_U1739 ( .A1(u5_mult_82_n6773), .A2(u5_mult_82_net65441), 
        .ZN(u5_mult_82_ab_38__49_) );
  NOR2_X1 u5_mult_82_U1738 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_net65513), .ZN(u5_mult_82_ab_34__38_) );
  NOR2_X1 u5_mult_82_U1737 ( .A1(u5_mult_82_net64937), .A2(u5_mult_82_n6699), 
        .ZN(u5_mult_82_ab_33__37_) );
  NOR2_X2 u5_mult_82_U1736 ( .A1(u5_mult_82_n6929), .A2(u5_mult_82_n6587), 
        .ZN(u5_mult_82_ab_15__17_) );
  NOR2_X1 u5_mult_82_U1735 ( .A1(u5_mult_82_n6797), .A2(u5_mult_82_n6701), 
        .ZN(u5_mult_82_ab_33__45_) );
  NOR2_X2 u5_mult_82_U1734 ( .A1(u5_mult_82_n6767), .A2(u5_mult_82_n1352), 
        .ZN(u5_mult_82_ab_38__50_) );
  NOR2_X2 u5_mult_82_U1733 ( .A1(u5_mult_82_n6833), .A2(u5_mult_82_n6544), 
        .ZN(u5_mult_82_ab_9__39_) );
  NOR2_X2 u5_mult_82_U1732 ( .A1(u5_mult_82_n6915), .A2(u5_mult_82_n6551), 
        .ZN(u5_mult_82_ab_10__19_) );
  NOR2_X2 u5_mult_82_U1731 ( .A1(u5_mult_82_n6922), .A2(u5_mult_82_n6515), 
        .ZN(u5_mult_82_ab_3__18_) );
  NOR2_X1 u5_mult_82_U1730 ( .A1(u5_mult_82_n6804), .A2(u5_mult_82_n6692), 
        .ZN(u5_mult_82_ab_32__44_) );
  NOR2_X2 u5_mult_82_U1729 ( .A1(u5_mult_82_n6767), .A2(u5_mult_82_n6698), 
        .ZN(u5_mult_82_ab_33__50_) );
  NOR2_X1 u5_mult_82_U1728 ( .A1(u5_mult_82_n6773), .A2(u5_mult_82_n6699), 
        .ZN(u5_mult_82_ab_33__49_) );
  NOR2_X2 u5_mult_82_U1727 ( .A1(u5_mult_82_n6812), .A2(u5_mult_82_n6630), 
        .ZN(u5_mult_82_ab_21__43_) );
  NOR2_X2 u5_mult_82_U1726 ( .A1(u5_mult_82_n6792), .A2(u5_mult_82_n6622), 
        .ZN(u5_mult_82_ab_20__46_) );
  NOR2_X2 u5_mult_82_U1725 ( .A1(u5_mult_82_n6785), .A2(u5_mult_82_n6623), 
        .ZN(u5_mult_82_ab_20__47_) );
  NOR2_X1 u5_mult_82_U1724 ( .A1(u5_mult_82_n6805), .A2(u5_mult_82_n6630), 
        .ZN(u5_mult_82_ab_21__44_) );
  NOR2_X1 u5_mult_82_U1723 ( .A1(u5_mult_82_n6877), .A2(u5_mult_82_net66019), 
        .ZN(u5_mult_82_ab_6__27_) );
  NOR2_X1 u5_mult_82_U1722 ( .A1(u5_mult_82_net64689), .A2(u5_mult_82_net66019), .ZN(u5_mult_82_ab_6__23_) );
  NOR2_X2 u5_mult_82_U1721 ( .A1(u5_mult_82_n6907), .A2(u5_mult_82_net66091), 
        .ZN(u5_mult_82_ab_2__20_) );
  NOR2_X2 u5_mult_82_U1720 ( .A1(u5_mult_82_n6811), .A2(u5_mult_82_n6677), 
        .ZN(u5_mult_82_ab_30__43_) );
  NOR2_X1 u5_mult_82_U1719 ( .A1(u5_mult_82_n6784), .A2(u5_mult_82_n6692), 
        .ZN(u5_mult_82_ab_32__47_) );
  NOR2_X2 u5_mult_82_U1718 ( .A1(u5_mult_82_n6778), .A2(u5_mult_82_n6692), 
        .ZN(u5_mult_82_ab_32__48_) );
  NOR2_X1 u5_mult_82_U1717 ( .A1(u5_mult_82_n6816), .A2(u5_mult_82_n6677), 
        .ZN(u5_mult_82_ab_30__42_) );
  NOR2_X1 u5_mult_82_U1716 ( .A1(u5_mult_82_n6832), .A2(u5_mult_82_n6614), 
        .ZN(u5_mult_82_ab_19__39_) );
  NOR2_X2 u5_mult_82_U1715 ( .A1(u5_mult_82_n6828), .A2(u5_mult_82_n6615), 
        .ZN(u5_mult_82_ab_19__40_) );
  NOR2_X2 u5_mult_82_U1714 ( .A1(u5_mult_82_n6829), .A2(u5_mult_82_n6520), 
        .ZN(u5_mult_82_ab_4__40_) );
  NOR2_X2 u5_mult_82_U1713 ( .A1(u5_mult_82_n6859), .A2(u5_mult_82_n6521), 
        .ZN(u5_mult_82_ab_4__30_) );
  NOR2_X2 u5_mult_82_U1712 ( .A1(u5_mult_82_net64961), .A2(u5_mult_82_net66089), .ZN(u5_mult_82_ab_2__38_) );
  NOR2_X2 u5_mult_82_U1711 ( .A1(u5_mult_82_net64673), .A2(u5_mult_82_net66091), .ZN(u5_mult_82_ab_2__22_) );
  NAND3_X2 u5_mult_82_U1710 ( .A1(u5_mult_82_n926), .A2(u5_mult_82_n927), .A3(
        u5_mult_82_n928), .ZN(u5_mult_82_CARRYB_27__41_) );
  INV_X4 u5_mult_82_U1709 ( .A(u5_mult_82_ab_3__40_), .ZN(u5_mult_82_n1590) );
  NOR2_X2 u5_mult_82_U1708 ( .A1(u5_mult_82_n6818), .A2(u5_mult_82_n6520), 
        .ZN(u5_mult_82_ab_4__42_) );
  INV_X8 u5_mult_82_U1707 ( .A(u5_mult_82_net64945), .ZN(u5_mult_82_net64943)
         );
  INV_X4 u5_mult_82_U1706 ( .A(u5_mult_82_n1265), .ZN(u5_mult_82_n1264) );
  INV_X8 u5_mult_82_U1705 ( .A(u5_mult_82_n6900), .ZN(u5_mult_82_n6899) );
  NOR2_X1 u5_mult_82_U1704 ( .A1(u5_mult_82_n6829), .A2(u5_mult_82_n6573), 
        .ZN(u5_mult_82_ab_13__40_) );
  NOR2_X2 u5_mult_82_U1703 ( .A1(u5_mult_82_n6806), .A2(u5_mult_82_n6520), 
        .ZN(u5_mult_82_ab_4__44_) );
  INV_X2 u5_mult_82_U1702 ( .A(u5_mult_82_ab_7__43_), .ZN(u5_mult_82_n1785) );
  NOR2_X2 u5_mult_82_U1701 ( .A1(u5_mult_82_net64687), .A2(u5_mult_82_net66091), .ZN(u5_mult_82_ab_2__23_) );
  NOR2_X2 u5_mult_82_U1700 ( .A1(u5_mult_82_n6774), .A2(u5_mult_82_n6655), 
        .ZN(u5_mult_82_ab_27__49_) );
  NOR2_X2 u5_mult_82_U1699 ( .A1(u5_mult_82_n6806), .A2(u5_mult_82_n6585), 
        .ZN(u5_mult_82_ab_15__44_) );
  NOR2_X1 u5_mult_82_U1698 ( .A1(u5_mult_82_n6762), .A2(u5_mult_82_n6585), 
        .ZN(u5_mult_82_ab_15__51_) );
  NOR2_X2 u5_mult_82_U1697 ( .A1(u5_mult_82_n6769), .A2(u5_mult_82_n6578), 
        .ZN(u5_mult_82_ab_14__50_) );
  NOR2_X2 u5_mult_82_U1696 ( .A1(u5_mult_82_n6768), .A2(u5_mult_82_n6655), 
        .ZN(u5_mult_82_ab_27__50_) );
  NOR2_X1 u5_mult_82_U1695 ( .A1(u5_mult_82_n6982), .A2(u5_mult_82_n6652), 
        .ZN(u5_mult_82_ab_26__52_) );
  NOR2_X2 u5_mult_82_U1694 ( .A1(u5_mult_82_n6761), .A2(u5_mult_82_n6655), 
        .ZN(u5_mult_82_ab_27__51_) );
  NOR2_X2 u5_mult_82_U1693 ( .A1(u5_mult_82_n6779), .A2(u5_mult_82_n6637), 
        .ZN(u5_mult_82_ab_22__48_) );
  NAND2_X2 u5_mult_82_U1692 ( .A1(u5_mult_82_ab_2__46_), .A2(
        u5_mult_82_SUMB_1__47_), .ZN(u5_mult_82_n1209) );
  NAND2_X2 u5_mult_82_U1691 ( .A1(u5_mult_82_CARRYB_1__46_), .A2(
        u5_mult_82_SUMB_1__47_), .ZN(u5_mult_82_n1208) );
  NOR2_X2 u5_mult_82_U1690 ( .A1(u5_mult_82_n6774), .A2(u5_mult_82_n6635), 
        .ZN(u5_mult_82_ab_22__49_) );
  NOR2_X2 u5_mult_82_U1689 ( .A1(u5_mult_82_n6761), .A2(u5_mult_82_n6634), 
        .ZN(u5_mult_82_ab_22__51_) );
  NOR2_X2 u5_mult_82_U1688 ( .A1(u5_mult_82_n6768), .A2(u5_mult_82_n6634), 
        .ZN(u5_mult_82_ab_22__50_) );
  INV_X4 u5_mult_82_U1687 ( .A(u5_mult_82_n1821), .ZN(u5_mult_82_n1822) );
  NOR2_X1 u5_mult_82_U1686 ( .A1(u5_mult_82_n6769), .A2(u5_mult_82_n6535), 
        .ZN(u5_mult_82_ab_8__50_) );
  NOR2_X2 u5_mult_82_U1685 ( .A1(u5_mult_82_n6775), .A2(u5_mult_82_n6538), 
        .ZN(u5_mult_82_ab_8__49_) );
  NOR2_X1 u5_mult_82_U1684 ( .A1(u5_mult_82_n6762), .A2(u5_mult_82_n6534), 
        .ZN(u5_mult_82_ab_8__51_) );
  NOR2_X1 u5_mult_82_U1683 ( .A1(u5_mult_82_n6946), .A2(u5_mult_82_n6716), 
        .ZN(u5_mult_82_ab_36__4_) );
  NOR2_X2 u5_mult_82_U1682 ( .A1(u5_mult_82_n6989), .A2(u5_mult_82_net66023), 
        .ZN(u5_mult_82_ab_6__0_) );
  NOR2_X2 u5_mult_82_U1681 ( .A1(u5_mult_82_n6989), .A2(u5_mult_82_n6560), 
        .ZN(u5_mult_82_ab_11__0_) );
  NOR2_X2 u5_mult_82_U1680 ( .A1(u5_mult_82_n6988), .A2(u5_mult_82_n6597), 
        .ZN(u5_mult_82_ab_16__0_) );
  NOR2_X2 u5_mult_82_U1679 ( .A1(u5_mult_82_n6988), .A2(u5_mult_82_n6631), 
        .ZN(u5_mult_82_ab_21__0_) );
  NOR2_X1 u5_mult_82_U1678 ( .A1(u5_mult_82_n6988), .A2(u5_mult_82_n6652), 
        .ZN(u5_mult_82_ab_26__0_) );
  NOR2_X2 u5_mult_82_U1677 ( .A1(u5_mult_82_n6987), .A2(u5_mult_82_n6687), 
        .ZN(u5_mult_82_ab_31__0_) );
  NOR2_X2 u5_mult_82_U1676 ( .A1(u5_mult_82_n6987), .A2(u5_mult_82_n6717), 
        .ZN(u5_mult_82_ab_36__0_) );
  NOR2_X1 u5_mult_82_U1675 ( .A1(u5_mult_82_net64379), .A2(u5_mult_82_n6709), 
        .ZN(u5_mult_82_ab_35__6_) );
  NOR2_X2 u5_mult_82_U1674 ( .A1(u5_mult_82_n6929), .A2(u5_mult_82_n6529), 
        .ZN(u5_mult_82_ab_7__17_) );
  NOR2_X2 u5_mult_82_U1673 ( .A1(u5_mult_82_n6922), .A2(u5_mult_82_n6529), 
        .ZN(u5_mult_82_ab_7__18_) );
  NOR2_X2 u5_mult_82_U1672 ( .A1(u5_mult_82_n6969), .A2(u5_mult_82_net66023), 
        .ZN(u5_mult_82_ab_6__1_) );
  NOR2_X2 u5_mult_82_U1671 ( .A1(u5_mult_82_n6969), .A2(u5_mult_82_n6560), 
        .ZN(u5_mult_82_ab_11__1_) );
  NOR2_X2 u5_mult_82_U1670 ( .A1(u5_mult_82_n6968), .A2(u5_mult_82_n6597), 
        .ZN(u5_mult_82_ab_16__1_) );
  NOR2_X2 u5_mult_82_U1669 ( .A1(u5_mult_82_n6968), .A2(u5_mult_82_n6631), 
        .ZN(u5_mult_82_ab_21__1_) );
  NOR2_X1 u5_mult_82_U1668 ( .A1(u5_mult_82_n6968), .A2(u5_mult_82_n6652), 
        .ZN(u5_mult_82_ab_26__1_) );
  NOR2_X1 u5_mult_82_U1667 ( .A1(u5_mult_82_n6967), .A2(u5_mult_82_n6687), 
        .ZN(u5_mult_82_ab_31__1_) );
  NOR2_X2 u5_mult_82_U1666 ( .A1(u5_mult_82_n6967), .A2(u5_mult_82_n6717), 
        .ZN(u5_mult_82_ab_36__1_) );
  NOR2_X2 u5_mult_82_U1665 ( .A1(u5_mult_82_n6962), .A2(u5_mult_82_net66023), 
        .ZN(u5_mult_82_ab_6__2_) );
  NOR2_X2 u5_mult_82_U1664 ( .A1(u5_mult_82_n6962), .A2(u5_mult_82_n6560), 
        .ZN(u5_mult_82_ab_11__2_) );
  NOR2_X2 u5_mult_82_U1663 ( .A1(u5_mult_82_n6961), .A2(u5_mult_82_n6597), 
        .ZN(u5_mult_82_ab_16__2_) );
  NOR2_X2 u5_mult_82_U1662 ( .A1(u5_mult_82_n6961), .A2(u5_mult_82_n6631), 
        .ZN(u5_mult_82_ab_21__2_) );
  INV_X16 u5_mult_82_U1661 ( .A(u5_mult_82_n6654), .ZN(u5_mult_82_n6660) );
  NOR2_X1 u5_mult_82_U1660 ( .A1(u5_mult_82_n6961), .A2(u5_mult_82_n6652), 
        .ZN(u5_mult_82_ab_26__2_) );
  NOR2_X1 u5_mult_82_U1659 ( .A1(u5_mult_82_n6960), .A2(u5_mult_82_n6687), 
        .ZN(u5_mult_82_ab_31__2_) );
  INV_X4 u5_mult_82_U1658 ( .A(u5_mult_82_ab_47__2_), .ZN(u5_mult_82_n1645) );
  NOR2_X1 u5_mult_82_U1657 ( .A1(u5_mult_82_n6960), .A2(u5_mult_82_n6749), 
        .ZN(u5_mult_82_ab_48__2_) );
  NOR2_X2 u5_mult_82_U1656 ( .A1(u5_mult_82_n6897), .A2(u5_mult_82_n6650), 
        .ZN(u5_mult_82_ab_26__21_) );
  INV_X4 u5_mult_82_U1655 ( .A(u5_mult_82_n6660), .ZN(u5_mult_82_n6657) );
  NOR2_X2 u5_mult_82_U1654 ( .A1(u5_mult_82_n6955), .A2(u5_mult_82_net66023), 
        .ZN(u5_mult_82_ab_6__3_) );
  NOR2_X2 u5_mult_82_U1653 ( .A1(u5_mult_82_n6955), .A2(u5_mult_82_n6560), 
        .ZN(u5_mult_82_ab_11__3_) );
  NOR2_X1 u5_mult_82_U1652 ( .A1(u5_mult_82_n6954), .A2(u5_mult_82_n6652), 
        .ZN(u5_mult_82_ab_26__3_) );
  NOR2_X2 u5_mult_82_U1651 ( .A1(u5_mult_82_n6953), .A2(u5_mult_82_n6717), 
        .ZN(u5_mult_82_ab_36__3_) );
  NOR2_X2 u5_mult_82_U1650 ( .A1(u5_mult_82_n6952), .A2(u5_mult_82_n6749), 
        .ZN(u5_mult_82_ab_48__3_) );
  NOR2_X1 u5_mult_82_U1649 ( .A1(u5_mult_82_n6946), .A2(u5_mult_82_n6695), 
        .ZN(u5_mult_82_ab_32__4_) );
  NOR2_X1 u5_mult_82_U1648 ( .A1(u5_mult_82_n6940), .A2(u5_mult_82_n6680), 
        .ZN(u5_mult_82_ab_30__7_) );
  INV_X8 u5_mult_82_U1647 ( .A(n4740), .ZN(u5_mult_82_n6902) );
  NOR2_X1 u5_mult_82_U1646 ( .A1(u5_mult_82_net64687), .A2(u5_mult_82_net65677), .ZN(u5_mult_82_ab_25__23_) );
  NOR2_X1 u5_mult_82_U1645 ( .A1(u5_mult_82_n6948), .A2(u5_mult_82_net66021), 
        .ZN(u5_mult_82_ab_6__4_) );
  NOR2_X1 u5_mult_82_U1644 ( .A1(u5_mult_82_n6948), .A2(u5_mult_82_n6559), 
        .ZN(u5_mult_82_ab_11__4_) );
  NOR2_X2 u5_mult_82_U1643 ( .A1(u5_mult_82_n6947), .A2(u5_mult_82_net65409), 
        .ZN(u5_mult_82_ab_40__4_) );
  NOR2_X1 u5_mult_82_U1642 ( .A1(u5_mult_82_n6946), .A2(u5_mult_82_net65189), 
        .ZN(u5_mult_82_ab_51__4_) );
  NOR2_X2 u5_mult_82_U1641 ( .A1(u5_mult_82_n6867), .A2(u5_mult_82_n6753), 
        .ZN(u5_mult_82_ab_49__28_) );
  INV_X4 u5_mult_82_U1640 ( .A(u5_mult_82_ab_34__21_), .ZN(u5_mult_82_n1733)
         );
  NOR2_X1 u5_mult_82_U1639 ( .A1(u5_mult_82_net64365), .A2(u5_mult_82_net66021), .ZN(u5_mult_82_ab_6__5_) );
  NOR2_X1 u5_mult_82_U1638 ( .A1(u5_mult_82_net64365), .A2(u5_mult_82_n6559), 
        .ZN(u5_mult_82_ab_11__5_) );
  NOR2_X2 u5_mult_82_U1637 ( .A1(u5_mult_82_net64363), .A2(u5_mult_82_n6623), 
        .ZN(u5_mult_82_ab_20__5_) );
  NOR2_X2 u5_mult_82_U1636 ( .A1(u5_mult_82_net64363), .A2(u5_mult_82_n6651), 
        .ZN(u5_mult_82_ab_26__5_) );
  INV_X4 u5_mult_82_U1635 ( .A(u5_mult_82_ab_48__30_), .ZN(u5_mult_82_n1699)
         );
  NOR2_X1 u5_mult_82_U1634 ( .A1(u5_mult_82_n6983), .A2(u5_mult_82_net65285), 
        .ZN(u5_mult_82_ab_47__52_) );
  NOR2_X2 u5_mult_82_U1633 ( .A1(u5_mult_82_n6759), .A2(u5_mult_82_n6746), 
        .ZN(u5_mult_82_ab_48__51_) );
  INV_X4 u5_mult_82_U1632 ( .A(u5_mult_82_n7010), .ZN(u5_mult_82_n6835) );
  NOR2_X2 u5_mult_82_U1631 ( .A1(u5_mult_82_n6875), .A2(u5_mult_82_n6715), 
        .ZN(u5_mult_82_ab_36__27_) );
  NOR2_X2 u5_mult_82_U1630 ( .A1(u5_mult_82_n6868), .A2(u5_mult_82_n6714), 
        .ZN(u5_mult_82_ab_36__28_) );
  NOR2_X2 u5_mult_82_U1629 ( .A1(u5_mult_82_n6913), .A2(u5_mult_82_net65515), 
        .ZN(u5_mult_82_ab_34__19_) );
  NOR2_X1 u5_mult_82_U1628 ( .A1(u5_mult_82_net64383), .A2(u5_mult_82_net66021), .ZN(u5_mult_82_ab_6__6_) );
  NOR2_X1 u5_mult_82_U1627 ( .A1(u5_mult_82_net64383), .A2(u5_mult_82_n6559), 
        .ZN(u5_mult_82_ab_11__6_) );
  NOR2_X2 u5_mult_82_U1626 ( .A1(u5_mult_82_n6856), .A2(u5_mult_82_n6753), 
        .ZN(u5_mult_82_ab_49__30_) );
  NOR2_X2 u5_mult_82_U1625 ( .A1(u5_mult_82_n6842), .A2(u5_mult_82_n6753), 
        .ZN(u5_mult_82_ab_49__32_) );
  INV_X8 u5_mult_82_U1624 ( .A(u5_mult_82_n7012), .ZN(u5_mult_82_n6855) );
  NOR2_X1 u5_mult_82_U1623 ( .A1(u5_mult_82_n6831), .A2(u5_mult_82_n6747), 
        .ZN(u5_mult_82_ab_48__39_) );
  NOR2_X2 u5_mult_82_U1622 ( .A1(u5_mult_82_n6777), .A2(u5_mult_82_n6752), 
        .ZN(u5_mult_82_ab_49__48_) );
  NOR2_X2 u5_mult_82_U1621 ( .A1(u5_mult_82_n6772), .A2(u5_mult_82_n6752), 
        .ZN(u5_mult_82_ab_49__49_) );
  INV_X8 u5_mult_82_U1620 ( .A(n4790), .ZN(u5_mult_82_n7009) );
  NOR2_X2 u5_mult_82_U1619 ( .A1(u5_mult_82_n6826), .A2(u5_mult_82_n6752), 
        .ZN(u5_mult_82_ab_49__40_) );
  NOR2_X2 u5_mult_82_U1618 ( .A1(u5_mult_82_n6874), .A2(u5_mult_82_net65285), 
        .ZN(u5_mult_82_ab_47__27_) );
  INV_X16 u5_mult_82_U1617 ( .A(u5_mult_82_net64459), .ZN(u5_mult_82_net64453)
         );
  INV_X4 u5_mult_82_U1616 ( .A(u5_mult_82_ab_33__19_), .ZN(u5_mult_82_n5143)
         );
  NOR2_X1 u5_mult_82_U1615 ( .A1(u5_mult_82_net64559), .A2(u5_mult_82_n6700), 
        .ZN(u5_mult_82_ab_33__16_) );
  INV_X4 u5_mult_82_U1614 ( .A(u5_mult_82_ab_20__24_), .ZN(u5_mult_82_n879) );
  NOR2_X1 u5_mult_82_U1613 ( .A1(u5_mult_82_n6942), .A2(u5_mult_82_net66021), 
        .ZN(u5_mult_82_ab_6__7_) );
  NOR2_X1 u5_mult_82_U1612 ( .A1(u5_mult_82_n6942), .A2(u5_mult_82_n6559), 
        .ZN(u5_mult_82_ab_11__7_) );
  NOR2_X1 u5_mult_82_U1611 ( .A1(u5_mult_82_net64417), .A2(u5_mult_82_n6630), 
        .ZN(u5_mult_82_ab_21__8_) );
  NOR2_X1 u5_mult_82_U1610 ( .A1(u5_mult_82_n6784), .A2(u5_mult_82_n6746), 
        .ZN(u5_mult_82_ab_48__47_) );
  NOR2_X1 u5_mult_82_U1609 ( .A1(u5_mult_82_n6797), .A2(u5_mult_82_n6746), 
        .ZN(u5_mult_82_ab_48__45_) );
  NOR2_X1 u5_mult_82_U1608 ( .A1(u5_mult_82_n6816), .A2(u5_mult_82_n6746), 
        .ZN(u5_mult_82_ab_48__42_) );
  INV_X8 u5_mult_82_U1607 ( .A(u5_mult_82_n1319), .ZN(u5_mult_82_net64477) );
  INV_X8 u5_mult_82_U1606 ( .A(u5_mult_82_net64499), .ZN(u5_mult_82_net64495)
         );
  NOR2_X1 u5_mult_82_U1605 ( .A1(u5_mult_82_n6838), .A2(u5_mult_82_n6699), 
        .ZN(u5_mult_82_ab_33__33_) );
  NOR2_X1 u5_mult_82_U1604 ( .A1(u5_mult_82_net64419), .A2(u5_mult_82_net66021), .ZN(u5_mult_82_ab_6__8_) );
  NOR2_X1 u5_mult_82_U1603 ( .A1(u5_mult_82_net64419), .A2(u5_mult_82_n6559), 
        .ZN(u5_mult_82_ab_11__8_) );
  NOR2_X1 u5_mult_82_U1602 ( .A1(u5_mult_82_net64437), .A2(u5_mult_82_n6580), 
        .ZN(u5_mult_82_ab_14__9_) );
  INV_X4 u5_mult_82_U1601 ( .A(u5_mult_82_ab_46__23_), .ZN(u5_mult_82_n3692)
         );
  NOR2_X1 u5_mult_82_U1600 ( .A1(u5_mult_82_net64489), .A2(u5_mult_82_net65717), .ZN(u5_mult_82_ab_23__12_) );
  NOR2_X2 u5_mult_82_U1599 ( .A1(u5_mult_82_net64525), .A2(u5_mult_82_n6637), 
        .ZN(u5_mult_82_ab_22__14_) );
  NOR2_X1 u5_mult_82_U1598 ( .A1(u5_mult_82_net64453), .A2(u5_mult_82_net65713), .ZN(u5_mult_82_ab_23__10_) );
  NOR2_X1 u5_mult_82_U1597 ( .A1(u5_mult_82_n6934), .A2(u5_mult_82_net65713), 
        .ZN(u5_mult_82_ab_23__15_) );
  NOR2_X1 u5_mult_82_U1596 ( .A1(u5_mult_82_net64561), .A2(u5_mult_82_net65713), .ZN(u5_mult_82_ab_23__16_) );
  INV_X8 u5_mult_82_U1595 ( .A(u5_mult_82_net64517), .ZN(u5_mult_82_net64513)
         );
  NOR2_X1 u5_mult_82_U1594 ( .A1(u5_mult_82_net64487), .A2(u5_mult_82_n6716), 
        .ZN(u5_mult_82_ab_36__12_) );
  NOR2_X1 u5_mult_82_U1593 ( .A1(u5_mult_82_net64437), .A2(u5_mult_82_net66021), .ZN(u5_mult_82_ab_6__9_) );
  NOR2_X1 u5_mult_82_U1592 ( .A1(u5_mult_82_net64455), .A2(u5_mult_82_n6580), 
        .ZN(u5_mult_82_ab_14__10_) );
  NAND3_X2 u5_mult_82_U1591 ( .A1(u5_mult_82_n4521), .A2(u5_mult_82_n4522), 
        .A3(u5_mult_82_n4523), .ZN(u5_mult_82_CARRYB_33__9_) );
  NOR2_X2 u5_mult_82_U1590 ( .A1(u5_mult_82_n6884), .A2(u5_mult_82_n6735), 
        .ZN(u5_mult_82_ab_44__25_) );
  NOR2_X2 u5_mult_82_U1589 ( .A1(u5_mult_82_n6874), .A2(u5_mult_82_net65353), 
        .ZN(u5_mult_82_ab_43__27_) );
  NOR2_X2 u5_mult_82_U1588 ( .A1(u5_mult_82_n6867), .A2(u5_mult_82_net65351), 
        .ZN(u5_mult_82_ab_43__28_) );
  NAND2_X2 u5_mult_82_U1587 ( .A1(u5_mult_82_n1628), .A2(
        u5_mult_82_SUMB_30__29_), .ZN(u5_mult_82_n4542) );
  NOR2_X2 u5_mult_82_U1586 ( .A1(u5_mult_82_n6875), .A2(u5_mult_82_n6685), 
        .ZN(u5_mult_82_ab_31__27_) );
  NOR2_X2 u5_mult_82_U1585 ( .A1(u5_mult_82_net64901), .A2(u5_mult_82_n6693), 
        .ZN(u5_mult_82_ab_32__35_) );
  NOR2_X2 u5_mult_82_U1584 ( .A1(u5_mult_82_n6880), .A2(u5_mult_82_n6664), 
        .ZN(u5_mult_82_ab_28__26_) );
  NAND2_X2 u5_mult_82_U1583 ( .A1(u5_mult_82_ab_29__17_), .A2(
        u5_mult_82_CARRYB_28__17_), .ZN(u5_mult_82_n1990) );
  NOR2_X2 u5_mult_82_U1582 ( .A1(u5_mult_82_net64669), .A2(u5_mult_82_n6602), 
        .ZN(u5_mult_82_ab_17__22_) );
  NOR2_X2 u5_mult_82_U1581 ( .A1(u5_mult_82_n6870), .A2(u5_mult_82_n6586), 
        .ZN(u5_mult_82_ab_15__28_) );
  NOR2_X1 u5_mult_82_U1580 ( .A1(u5_mult_82_net64455), .A2(u5_mult_82_net66021), .ZN(u5_mult_82_ab_6__10_) );
  NOR2_X2 u5_mult_82_U1579 ( .A1(u5_mult_82_net64473), .A2(u5_mult_82_n6588), 
        .ZN(u5_mult_82_ab_15__11_) );
  NAND2_X2 u5_mult_82_U1578 ( .A1(u5_mult_82_n3139), .A2(u5_mult_82_n4232), 
        .ZN(u5_mult_82_n4204) );
  NOR2_X1 u5_mult_82_U1577 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_net65351), .ZN(u5_mult_82_ab_43__36_) );
  NOR2_X1 u5_mult_82_U1576 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_net65351), .ZN(u5_mult_82_ab_43__38_) );
  NOR2_X1 u5_mult_82_U1575 ( .A1(u5_mult_82_n6816), .A2(u5_mult_82_net65385), 
        .ZN(u5_mult_82_ab_41__42_) );
  NOR2_X2 u5_mult_82_U1574 ( .A1(u5_mult_82_n6811), .A2(u5_mult_82_net65385), 
        .ZN(u5_mult_82_ab_41__43_) );
  NOR2_X1 u5_mult_82_U1573 ( .A1(u5_mult_82_n6983), .A2(u5_mult_82_net65375), 
        .ZN(u5_mult_82_ab_42__52_) );
  NOR2_X2 u5_mult_82_U1572 ( .A1(u5_mult_82_n6759), .A2(u5_mult_82_net65349), 
        .ZN(u5_mult_82_ab_43__51_) );
  NOR2_X2 u5_mult_82_U1571 ( .A1(u5_mult_82_n6898), .A2(u5_mult_82_n6587), 
        .ZN(u5_mult_82_ab_15__21_) );
  NOR2_X1 u5_mult_82_U1570 ( .A1(u5_mult_82_n6877), .A2(u5_mult_82_n6579), 
        .ZN(u5_mult_82_ab_14__27_) );
  NOR2_X1 u5_mult_82_U1569 ( .A1(u5_mult_82_net64473), .A2(u5_mult_82_net66021), .ZN(u5_mult_82_ab_6__11_) );
  NOR2_X2 u5_mult_82_U1568 ( .A1(u5_mult_82_n6859), .A2(u5_mult_82_n6578), 
        .ZN(u5_mult_82_ab_14__30_) );
  INV_X4 u5_mult_82_U1567 ( .A(u5_mult_82_ab_17__32_), .ZN(u5_mult_82_n4866)
         );
  NOR2_X1 u5_mult_82_U1566 ( .A1(u5_mult_82_net64491), .A2(u5_mult_82_net66021), .ZN(u5_mult_82_ab_6__12_) );
  NOR2_X1 u5_mult_82_U1565 ( .A1(u5_mult_82_net64527), .A2(u5_mult_82_n6573), 
        .ZN(u5_mult_82_ab_13__14_) );
  NOR2_X2 u5_mult_82_U1564 ( .A1(u5_mult_82_n6897), .A2(u5_mult_82_net65407), 
        .ZN(u5_mult_82_ab_40__21_) );
  NOR2_X2 u5_mult_82_U1563 ( .A1(u5_mult_82_n6798), .A2(u5_mult_82_net65403), 
        .ZN(u5_mult_82_ab_40__45_) );
  NOR2_X1 u5_mult_82_U1562 ( .A1(u5_mult_82_n6791), .A2(u5_mult_82_net65369), 
        .ZN(u5_mult_82_ab_42__46_) );
  NOR2_X2 u5_mult_82_U1561 ( .A1(u5_mult_82_n6766), .A2(u5_mult_82_net65349), 
        .ZN(u5_mult_82_ab_43__50_) );
  NOR2_X2 u5_mult_82_U1560 ( .A1(u5_mult_82_n6772), .A2(u5_mult_82_net65349), 
        .ZN(u5_mult_82_ab_43__49_) );
  NOR2_X2 u5_mult_82_U1559 ( .A1(u5_mult_82_n6777), .A2(u5_mult_82_net65349), 
        .ZN(u5_mult_82_ab_43__48_) );
  NOR2_X1 u5_mult_82_U1558 ( .A1(u5_mult_82_n6784), .A2(u5_mult_82_net65349), 
        .ZN(u5_mult_82_ab_43__47_) );
  NOR2_X2 u5_mult_82_U1557 ( .A1(u5_mult_82_n6921), .A2(u5_mult_82_n6595), 
        .ZN(u5_mult_82_ab_16__18_) );
  NOR2_X2 u5_mult_82_U1556 ( .A1(u5_mult_82_n6858), .A2(u5_mult_82_n6642), 
        .ZN(u5_mult_82_ab_24__30_) );
  NOR2_X2 u5_mult_82_U1555 ( .A1(u5_mult_82_net64509), .A2(u5_mult_82_n6530), 
        .ZN(u5_mult_82_ab_7__13_) );
  NOR2_X2 u5_mult_82_U1554 ( .A1(u5_mult_82_n6935), .A2(u5_mult_82_n6588), 
        .ZN(u5_mult_82_ab_15__15_) );
  NOR2_X2 u5_mult_82_U1553 ( .A1(u5_mult_82_net64685), .A2(u5_mult_82_n6728), 
        .ZN(u5_mult_82_ab_39__23_) );
  NOR2_X1 u5_mult_82_U1552 ( .A1(u5_mult_82_net64905), .A2(u5_mult_82_n6571), 
        .ZN(u5_mult_82_ab_13__35_) );
  NOR2_X1 u5_mult_82_U1551 ( .A1(u5_mult_82_net64671), .A2(u5_mult_82_n6558), 
        .ZN(u5_mult_82_ab_11__22_) );
  NOR2_X2 u5_mult_82_U1550 ( .A1(u5_mult_82_net64527), .A2(u5_mult_82_n6530), 
        .ZN(u5_mult_82_ab_7__14_) );
  NOR2_X2 u5_mult_82_U1549 ( .A1(u5_mult_82_n6821), .A2(u5_mult_82_n6713), 
        .ZN(u5_mult_82_ab_36__41_) );
  NOR2_X2 u5_mult_82_U1548 ( .A1(u5_mult_82_net64887), .A2(u5_mult_82_n6528), 
        .ZN(u5_mult_82_ab_7__34_) );
  NOR2_X2 u5_mult_82_U1547 ( .A1(u5_mult_82_net64563), .A2(u5_mult_82_n6529), 
        .ZN(u5_mult_82_ab_7__16_) );
  NOR2_X1 u5_mult_82_U1546 ( .A1(u5_mult_82_n6816), .A2(u5_mult_82_n6713), 
        .ZN(u5_mult_82_ab_36__42_) );
  NOR2_X2 u5_mult_82_U1545 ( .A1(u5_mult_82_n6811), .A2(u5_mult_82_n6713), 
        .ZN(u5_mult_82_ab_36__43_) );
  NOR2_X1 u5_mult_82_U1544 ( .A1(u5_mult_82_n6784), .A2(u5_mult_82_n6706), 
        .ZN(u5_mult_82_ab_35__47_) );
  NOR2_X2 u5_mult_82_U1543 ( .A1(u5_mult_82_n6773), .A2(u5_mult_82_n6720), 
        .ZN(u5_mult_82_ab_37__49_) );
  NOR2_X1 u5_mult_82_U1542 ( .A1(u5_mult_82_n6982), .A2(u5_mult_82_n6723), 
        .ZN(u5_mult_82_ab_37__52_) );
  NOR2_X2 u5_mult_82_U1541 ( .A1(u5_mult_82_n6760), .A2(u5_mult_82_n1352), 
        .ZN(u5_mult_82_ab_38__51_) );
  NOR2_X1 u5_mult_82_U1540 ( .A1(u5_mult_82_n6832), .A2(u5_mult_82_net65513), 
        .ZN(u5_mult_82_ab_34__39_) );
  NOR2_X1 u5_mult_82_U1539 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6699), 
        .ZN(u5_mult_82_ab_33__38_) );
  NOR2_X2 u5_mult_82_U1538 ( .A1(u5_mult_82_net64903), .A2(u5_mult_82_n6642), 
        .ZN(u5_mult_82_ab_24__35_) );
  NAND3_X2 u5_mult_82_U1537 ( .A1(u5_mult_82_n2312), .A2(u5_mult_82_n2313), 
        .A3(u5_mult_82_n2314), .ZN(u5_mult_82_CARRYB_23__40_) );
  NOR2_X2 u5_mult_82_U1536 ( .A1(u5_mult_82_net64905), .A2(u5_mult_82_n6544), 
        .ZN(u5_mult_82_ab_9__35_) );
  NOR2_X2 u5_mult_82_U1535 ( .A1(u5_mult_82_n6898), .A2(u5_mult_82_n6551), 
        .ZN(u5_mult_82_ab_10__21_) );
  NOR2_X2 u5_mult_82_U1534 ( .A1(u5_mult_82_n6845), .A2(u5_mult_82_n6528), 
        .ZN(u5_mult_82_ab_7__32_) );
  NOR2_X1 u5_mult_82_U1533 ( .A1(u5_mult_82_n6791), .A2(u5_mult_82_net65515), 
        .ZN(u5_mult_82_ab_34__46_) );
  NOR2_X2 u5_mult_82_U1532 ( .A1(u5_mult_82_n6767), .A2(u5_mult_82_n6719), 
        .ZN(u5_mult_82_ab_37__50_) );
  NOR2_X2 u5_mult_82_U1531 ( .A1(u5_mult_82_net64937), .A2(u5_mult_82_n6693), 
        .ZN(u5_mult_82_ab_32__37_) );
  NOR2_X1 u5_mult_82_U1530 ( .A1(u5_mult_82_n6844), .A2(u5_mult_82_n6614), 
        .ZN(u5_mult_82_ab_19__32_) );
  NOR2_X2 u5_mult_82_U1529 ( .A1(u5_mult_82_net64885), .A2(u5_mult_82_n6608), 
        .ZN(u5_mult_82_ab_18__34_) );
  NOR2_X1 u5_mult_82_U1528 ( .A1(u5_mult_82_n6852), .A2(u5_mult_82_net66035), 
        .ZN(u5_mult_82_ab_5__31_) );
  NOR2_X1 u5_mult_82_U1527 ( .A1(u5_mult_82_n6798), .A2(u5_mult_82_n6630), 
        .ZN(u5_mult_82_ab_21__45_) );
  NOR2_X1 u5_mult_82_U1526 ( .A1(u5_mult_82_n6797), .A2(u5_mult_82_n6677), 
        .ZN(u5_mult_82_ab_30__45_) );
  NOR2_X1 u5_mult_82_U1525 ( .A1(u5_mult_82_n6779), .A2(u5_mult_82_n6616), 
        .ZN(u5_mult_82_ab_19__48_) );
  INV_X4 u5_mult_82_U1524 ( .A(u5_mult_82_ab_7__40_), .ZN(u5_mult_82_n3999) );
  NOR2_X2 u5_mult_82_U1523 ( .A1(u5_mult_82_n6893), .A2(u5_mult_82_net66037), 
        .ZN(u5_mult_82_ab_5__24_) );
  NOR2_X1 u5_mult_82_U1522 ( .A1(u5_mult_82_n6982), .A2(u5_mult_82_n6674), 
        .ZN(u5_mult_82_ab_29__52_) );
  NOR2_X2 u5_mult_82_U1521 ( .A1(u5_mult_82_n6760), .A2(u5_mult_82_n6677), 
        .ZN(u5_mult_82_ab_30__51_) );
  NOR2_X2 u5_mult_82_U1520 ( .A1(u5_mult_82_n6822), .A2(u5_mult_82_n6607), 
        .ZN(u5_mult_82_ab_18__41_) );
  NOR2_X1 u5_mult_82_U1519 ( .A1(u5_mult_82_n6823), .A2(u5_mult_82_net66019), 
        .ZN(u5_mult_82_ab_6__41_) );
  NOR2_X1 u5_mult_82_U1518 ( .A1(u5_mult_82_n6833), .A2(u5_mult_82_n6571), 
        .ZN(u5_mult_82_ab_13__39_) );
  NOR2_X2 u5_mult_82_U1517 ( .A1(u5_mult_82_n6813), .A2(u5_mult_82_net66087), 
        .ZN(u5_mult_82_ab_2__43_) );
  NOR2_X2 u5_mult_82_U1516 ( .A1(u5_mult_82_n6767), .A2(u5_mult_82_n6662), 
        .ZN(u5_mult_82_ab_28__50_) );
  NOR2_X2 u5_mult_82_U1515 ( .A1(u5_mult_82_n6774), .A2(u5_mult_82_n6649), 
        .ZN(u5_mult_82_ab_26__49_) );
  NOR2_X2 u5_mult_82_U1514 ( .A1(u5_mult_82_n6793), .A2(u5_mult_82_n6573), 
        .ZN(u5_mult_82_ab_13__46_) );
  NAND2_X2 u5_mult_82_U1513 ( .A1(u5_mult_82_ab_12__46_), .A2(u5_mult_82_n4101), .ZN(u5_mult_82_n4891) );
  NOR2_X1 u5_mult_82_U1512 ( .A1(u5_mult_82_n6780), .A2(u5_mult_82_n6559), 
        .ZN(u5_mult_82_ab_11__48_) );
  NOR2_X2 u5_mult_82_U1511 ( .A1(u5_mult_82_n6768), .A2(u5_mult_82_n6620), 
        .ZN(u5_mult_82_ab_20__50_) );
  NOR2_X2 u5_mult_82_U1510 ( .A1(u5_mult_82_n6793), .A2(u5_mult_82_net66033), 
        .ZN(u5_mult_82_ab_5__46_) );
  NOR2_X2 u5_mult_82_U1509 ( .A1(u5_mult_82_n6761), .A2(u5_mult_82_n6627), 
        .ZN(u5_mult_82_ab_21__51_) );
  NOR2_X2 u5_mult_82_U1508 ( .A1(u5_mult_82_n6780), .A2(u5_mult_82_net66033), 
        .ZN(u5_mult_82_ab_5__48_) );
  NOR2_X1 u5_mult_82_U1507 ( .A1(u5_mult_82_net64361), .A2(u5_mult_82_n6709), 
        .ZN(u5_mult_82_ab_35__5_) );
  INV_X16 u5_mult_82_U1506 ( .A(u5_mult_82_n6930), .ZN(u5_mult_82_n6929) );
  NOR2_X2 u5_mult_82_U1505 ( .A1(u5_mult_82_n6929), .A2(u5_mult_82_net66019), 
        .ZN(u5_mult_82_ab_6__17_) );
  NOR2_X1 u5_mult_82_U1504 ( .A1(u5_mult_82_n6915), .A2(u5_mult_82_net66019), 
        .ZN(u5_mult_82_ab_6__19_) );
  INV_X16 u5_mult_82_U1503 ( .A(u5_mult_82_n6985), .ZN(u5_mult_82_n6991) );
  INV_X8 u5_mult_82_U1502 ( .A(u6_N0), .ZN(u5_mult_82_n6985) );
  INV_X4 u5_mult_82_U1501 ( .A(u5_mult_82_n6985), .ZN(u5_mult_82_n6990) );
  NOR2_X2 u5_mult_82_U1500 ( .A1(u5_mult_82_n6960), .A2(u5_mult_82_n6696), 
        .ZN(u5_mult_82_ab_32__2_) );
  NOR2_X1 u5_mult_82_U1499 ( .A1(u5_mult_82_n6897), .A2(u5_mult_82_net65677), 
        .ZN(u5_mult_82_ab_25__21_) );
  INV_X16 u5_mult_82_U1498 ( .A(u5_mult_82_n6966), .ZN(u5_mult_82_n6971) );
  NOR2_X2 u5_mult_82_U1497 ( .A1(u5_mult_82_n6954), .A2(u5_mult_82_n6597), 
        .ZN(u5_mult_82_ab_16__3_) );
  NOR2_X2 u5_mult_82_U1496 ( .A1(u5_mult_82_n6954), .A2(u5_mult_82_n6631), 
        .ZN(u5_mult_82_ab_21__3_) );
  NOR2_X2 u5_mult_82_U1495 ( .A1(u5_mult_82_n6953), .A2(u5_mult_82_n6696), 
        .ZN(u5_mult_82_ab_32__3_) );
  INV_X8 u5_mult_82_U1494 ( .A(u5_mult_82_n6959), .ZN(u5_mult_82_n6964) );
  NOR2_X1 u5_mult_82_U1493 ( .A1(u5_mult_82_net64433), .A2(u5_mult_82_n6686), 
        .ZN(u5_mult_82_ab_31__9_) );
  NOR2_X1 u5_mult_82_U1492 ( .A1(u5_mult_82_net64669), .A2(u5_mult_82_net65677), .ZN(u5_mult_82_ab_25__22_) );
  NOR2_X2 u5_mult_82_U1491 ( .A1(u5_mult_82_n6947), .A2(u5_mult_82_n6596), 
        .ZN(u5_mult_82_ab_16__4_) );
  NOR2_X1 u5_mult_82_U1490 ( .A1(u5_mult_82_n6947), .A2(u5_mult_82_n6630), 
        .ZN(u5_mult_82_ab_21__4_) );
  NOR2_X1 u5_mult_82_U1489 ( .A1(u5_mult_82_net64361), .A2(u5_mult_82_n6686), 
        .ZN(u5_mult_82_ab_31__5_) );
  NOR2_X2 u5_mult_82_U1488 ( .A1(u5_mult_82_net64363), .A2(u5_mult_82_n6596), 
        .ZN(u5_mult_82_ab_16__5_) );
  NOR2_X2 u5_mult_82_U1487 ( .A1(u5_mult_82_net64381), .A2(u5_mult_82_n6630), 
        .ZN(u5_mult_82_ab_21__6_) );
  NOR2_X2 u5_mult_82_U1486 ( .A1(u5_mult_82_net64363), .A2(u5_mult_82_n6658), 
        .ZN(u5_mult_82_ab_27__5_) );
  NOR2_X1 u5_mult_82_U1485 ( .A1(u5_mult_82_net64361), .A2(u5_mult_82_net65229), .ZN(u5_mult_82_ab_50__5_) );
  INV_X16 u5_mult_82_U1484 ( .A(u5_mult_82_n6855), .ZN(u5_mult_82_n6849) );
  NOR2_X2 u5_mult_82_U1483 ( .A1(u5_mult_82_n6867), .A2(u5_mult_82_net65279), 
        .ZN(u5_mult_82_ab_47__28_) );
  INV_X16 u5_mult_82_U1482 ( .A(u5_mult_82_n7016), .ZN(u5_mult_82_n6873) );
  NOR2_X1 u5_mult_82_U1481 ( .A1(u5_mult_82_n6940), .A2(u5_mult_82_n6722), 
        .ZN(u5_mult_82_ab_37__7_) );
  NOR2_X1 u5_mult_82_U1480 ( .A1(u5_mult_82_n6831), .A2(u5_mult_82_n6753), 
        .ZN(u5_mult_82_ab_49__39_) );
  NOR2_X2 u5_mult_82_U1479 ( .A1(u5_mult_82_n6896), .A2(u5_mult_82_n6694), 
        .ZN(u5_mult_82_ab_32__21_) );
  NOR2_X2 u5_mult_82_U1478 ( .A1(u5_mult_82_n6772), .A2(u5_mult_82_n6746), 
        .ZN(u5_mult_82_ab_48__49_) );
  NOR2_X2 u5_mult_82_U1477 ( .A1(u5_mult_82_n6777), .A2(u5_mult_82_n6746), 
        .ZN(u5_mult_82_ab_48__48_) );
  NOR2_X2 u5_mult_82_U1476 ( .A1(u5_mult_82_n6803), .A2(u5_mult_82_n6746), 
        .ZN(u5_mult_82_ab_48__44_) );
  INV_X8 u5_mult_82_U1475 ( .A(u5_mult_82_net64427), .ZN(u5_mult_82_net64423)
         );
  NOR2_X2 u5_mult_82_U1474 ( .A1(u5_mult_82_n6838), .A2(u5_mult_82_n6693), 
        .ZN(u5_mult_82_ab_32__33_) );
  NOR2_X1 u5_mult_82_U1473 ( .A1(u5_mult_82_net64419), .A2(u5_mult_82_n6580), 
        .ZN(u5_mult_82_ab_14__8_) );
  NOR2_X1 u5_mult_82_U1472 ( .A1(u5_mult_82_n6816), .A2(u5_mult_82_net65277), 
        .ZN(u5_mult_82_ab_47__42_) );
  NOR2_X2 u5_mult_82_U1471 ( .A1(u5_mult_82_net64883), .A2(u5_mult_82_n6693), 
        .ZN(u5_mult_82_ab_32__34_) );
  NOR2_X2 u5_mult_82_U1470 ( .A1(u5_mult_82_net64471), .A2(u5_mult_82_n6603), 
        .ZN(u5_mult_82_ab_17__11_) );
  INV_X8 u5_mult_82_U1469 ( .A(u5_mult_82_net64535), .ZN(u5_mult_82_net64531)
         );
  NOR2_X1 u5_mult_82_U1468 ( .A1(u5_mult_82_n6933), .A2(u5_mult_82_n6709), 
        .ZN(u5_mult_82_ab_35__15_) );
  INV_X4 u5_mult_82_U1467 ( .A(u5_mult_82_ab_34__15_), .ZN(u5_mult_82_n3580)
         );
  NOR2_X1 u5_mult_82_U1466 ( .A1(u5_mult_82_net64455), .A2(u5_mult_82_n6546), 
        .ZN(u5_mult_82_ab_9__10_) );
  INV_X4 u5_mult_82_U1465 ( .A(u5_mult_82_ab_43__20_), .ZN(u5_mult_82_n2172)
         );
  NOR2_X2 u5_mult_82_U1464 ( .A1(u5_mult_82_n6884), .A2(u5_mult_82_net65353), 
        .ZN(u5_mult_82_ab_43__25_) );
  NOR2_X2 u5_mult_82_U1463 ( .A1(u5_mult_82_n6862), .A2(u5_mult_82_net65387), 
        .ZN(u5_mult_82_ab_41__29_) );
  INV_X16 u5_mult_82_U1462 ( .A(u5_mult_82_n1375), .ZN(u5_mult_82_net65361) );
  NOR2_X1 u5_mult_82_U1461 ( .A1(u5_mult_82_net64507), .A2(u5_mult_82_n6623), 
        .ZN(u5_mult_82_ab_20__13_) );
  NOR2_X1 u5_mult_82_U1460 ( .A1(u5_mult_82_n6928), .A2(u5_mult_82_n6622), 
        .ZN(u5_mult_82_ab_20__17_) );
  INV_X8 u5_mult_82_U1459 ( .A(u5_mult_82_n6932), .ZN(u5_mult_82_n6937) );
  NOR2_X2 u5_mult_82_U1458 ( .A1(u5_mult_82_net64473), .A2(u5_mult_82_n6546), 
        .ZN(u5_mult_82_ab_9__11_) );
  NOR2_X1 u5_mult_82_U1457 ( .A1(u5_mult_82_net64489), .A2(u5_mult_82_n6623), 
        .ZN(u5_mult_82_ab_20__12_) );
  NOR2_X1 u5_mult_82_U1456 ( .A1(u5_mult_82_net64921), .A2(u5_mult_82_net65405), .ZN(u5_mult_82_ab_40__36_) );
  NOR2_X2 u5_mult_82_U1455 ( .A1(u5_mult_82_net64939), .A2(u5_mult_82_net65405), .ZN(u5_mult_82_ab_40__37_) );
  NOR2_X1 u5_mult_82_U1454 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_net65369), .ZN(u5_mult_82_ab_42__38_) );
  NOR2_X2 u5_mult_82_U1453 ( .A1(u5_mult_82_n6827), .A2(u5_mult_82_net65385), 
        .ZN(u5_mult_82_ab_41__40_) );
  NOR2_X2 u5_mult_82_U1452 ( .A1(u5_mult_82_n6817), .A2(u5_mult_82_net65403), 
        .ZN(u5_mult_82_ab_40__42_) );
  NOR2_X1 u5_mult_82_U1451 ( .A1(u5_mult_82_n6983), .A2(u5_mult_82_net65393), 
        .ZN(u5_mult_82_ab_41__52_) );
  NOR2_X2 u5_mult_82_U1450 ( .A1(u5_mult_82_n6759), .A2(u5_mult_82_net65369), 
        .ZN(u5_mult_82_ab_42__51_) );
  NOR2_X2 u5_mult_82_U1449 ( .A1(u5_mult_82_n6921), .A2(u5_mult_82_n6622), 
        .ZN(u5_mult_82_ab_20__18_) );
  NOR2_X2 u5_mult_82_U1448 ( .A1(u5_mult_82_n6921), .A2(u5_mult_82_n6650), 
        .ZN(u5_mult_82_ab_26__18_) );
  INV_X16 u5_mult_82_U1447 ( .A(u5_mult_82_n6584), .ZN(u5_mult_82_n6591) );
  NOR2_X2 u5_mult_82_U1446 ( .A1(u5_mult_82_net64491), .A2(u5_mult_82_n6546), 
        .ZN(u5_mult_82_ab_9__12_) );
  NOR2_X2 u5_mult_82_U1445 ( .A1(u5_mult_82_net64509), .A2(u5_mult_82_n6546), 
        .ZN(u5_mult_82_ab_9__13_) );
  NOR2_X1 u5_mult_82_U1444 ( .A1(u5_mult_82_n6804), .A2(u5_mult_82_n6729), 
        .ZN(u5_mult_82_ab_39__44_) );
  NOR2_X1 u5_mult_82_U1443 ( .A1(u5_mult_82_n6797), .A2(u5_mult_82_n6729), 
        .ZN(u5_mult_82_ab_39__45_) );
  NOR2_X1 u5_mult_82_U1442 ( .A1(u5_mult_82_n6791), .A2(u5_mult_82_net65349), 
        .ZN(u5_mult_82_ab_43__46_) );
  NOR2_X1 u5_mult_82_U1441 ( .A1(u5_mult_82_n6852), .A2(u5_mult_82_n6565), 
        .ZN(u5_mult_82_ab_12__31_) );
  NOR2_X2 u5_mult_82_U1440 ( .A1(u5_mult_82_n6870), .A2(u5_mult_82_n6565), 
        .ZN(u5_mult_82_ab_12__28_) );
  INV_X4 u5_mult_82_U1439 ( .A(u5_mult_82_n6937), .ZN(u5_mult_82_n6935) );
  NOR2_X1 u5_mult_82_U1438 ( .A1(u5_mult_82_net64523), .A2(u5_mult_82_n6673), 
        .ZN(u5_mult_82_ab_29__14_) );
  NOR2_X2 u5_mult_82_U1437 ( .A1(u5_mult_82_net64527), .A2(u5_mult_82_n6523), 
        .ZN(u5_mult_82_ab_4__14_) );
  NOR2_X2 u5_mult_82_U1436 ( .A1(u5_mult_82_n6922), .A2(u5_mult_82_n6587), 
        .ZN(u5_mult_82_ab_15__18_) );
  NOR2_X2 u5_mult_82_U1435 ( .A1(u5_mult_82_n6821), .A2(u5_mult_82_net65515), 
        .ZN(u5_mult_82_ab_34__41_) );
  NOR2_X2 u5_mult_82_U1434 ( .A1(u5_mult_82_n6778), .A2(u5_mult_82_n6723), 
        .ZN(u5_mult_82_ab_37__48_) );
  INV_X4 u5_mult_82_U1433 ( .A(u5_mult_82_ab_12__18_), .ZN(u5_mult_82_n2593)
         );
  NOR2_X2 u5_mult_82_U1432 ( .A1(u5_mult_82_net64689), .A2(u5_mult_82_n6545), 
        .ZN(u5_mult_82_ab_9__23_) );
  NOR2_X2 u5_mult_82_U1431 ( .A1(u5_mult_82_net64671), .A2(u5_mult_82_n6545), 
        .ZN(u5_mult_82_ab_9__22_) );
  NOR2_X2 u5_mult_82_U1430 ( .A1(u5_mult_82_net64563), .A2(u5_mult_82_n6515), 
        .ZN(u5_mult_82_ab_3__16_) );
  NOR2_X1 u5_mult_82_U1429 ( .A1(u5_mult_82_n6784), .A2(u5_mult_82_net65517), 
        .ZN(u5_mult_82_ab_34__47_) );
  NOR2_X2 u5_mult_82_U1428 ( .A1(u5_mult_82_n6767), .A2(u5_mult_82_n6713), 
        .ZN(u5_mult_82_ab_36__50_) );
  NOR2_X2 u5_mult_82_U1427 ( .A1(u5_mult_82_n6898), .A2(u5_mult_82_n6536), 
        .ZN(u5_mult_82_ab_8__21_) );
  NOR2_X2 u5_mult_82_U1426 ( .A1(u5_mult_82_net64887), .A2(u5_mult_82_net66035), .ZN(u5_mult_82_ab_5__34_) );
  NOR2_X2 u5_mult_82_U1425 ( .A1(u5_mult_82_n6906), .A2(u5_mult_82_n6529), 
        .ZN(u5_mult_82_ab_7__20_) );
  NOR2_X2 u5_mult_82_U1424 ( .A1(u5_mult_82_net64937), .A2(u5_mult_82_n6684), 
        .ZN(u5_mult_82_ab_31__37_) );
  NOR2_X1 u5_mult_82_U1423 ( .A1(u5_mult_82_n6797), .A2(u5_mult_82_n6692), 
        .ZN(u5_mult_82_ab_32__45_) );
  NOR2_X1 u5_mult_82_U1422 ( .A1(u5_mult_82_n6791), .A2(u5_mult_82_n6701), 
        .ZN(u5_mult_82_ab_33__46_) );
  NOR2_X1 u5_mult_82_U1421 ( .A1(u5_mult_82_n6982), .A2(u5_mult_82_n6710), 
        .ZN(u5_mult_82_ab_35__52_) );
  NOR2_X2 u5_mult_82_U1420 ( .A1(u5_mult_82_n6760), .A2(u5_mult_82_n6713), 
        .ZN(u5_mult_82_ab_36__51_) );
  NOR2_X1 u5_mult_82_U1419 ( .A1(u5_mult_82_n6805), .A2(u5_mult_82_n6622), 
        .ZN(u5_mult_82_ab_20__44_) );
  NOR2_X2 u5_mult_82_U1418 ( .A1(u5_mult_82_n6845), .A2(u5_mult_82_n6521), 
        .ZN(u5_mult_82_ab_4__32_) );
  NOR2_X2 u5_mult_82_U1417 ( .A1(u5_mult_82_n6798), .A2(u5_mult_82_n6622), 
        .ZN(u5_mult_82_ab_20__45_) );
  NOR2_X2 u5_mult_82_U1416 ( .A1(u5_mult_82_n6811), .A2(u5_mult_82_n6670), 
        .ZN(u5_mult_82_ab_29__43_) );
  NOR2_X1 u5_mult_82_U1415 ( .A1(u5_mult_82_n6816), .A2(u5_mult_82_n6670), 
        .ZN(u5_mult_82_ab_29__42_) );
  INV_X2 u5_mult_82_U1414 ( .A(u5_mult_82_ab_16__42_), .ZN(u5_mult_82_n5549)
         );
  NOR2_X2 u5_mult_82_U1413 ( .A1(u5_mult_82_n6768), .A2(u5_mult_82_n6593), 
        .ZN(u5_mult_82_ab_16__50_) );
  NOR2_X2 u5_mult_82_U1412 ( .A1(u5_mult_82_n6813), .A2(u5_mult_82_n6520), 
        .ZN(u5_mult_82_ab_4__43_) );
  NOR2_X2 u5_mult_82_U1411 ( .A1(u5_mult_82_n6792), .A2(u5_mult_82_n6655), 
        .ZN(u5_mult_82_ab_27__46_) );
  NOR2_X1 u5_mult_82_U1410 ( .A1(u5_mult_82_n6982), .A2(u5_mult_82_n6659), 
        .ZN(u5_mult_82_ab_27__52_) );
  NOR2_X2 u5_mult_82_U1409 ( .A1(u5_mult_82_n6760), .A2(u5_mult_82_n6662), 
        .ZN(u5_mult_82_ab_28__51_) );
  NOR2_X2 u5_mult_82_U1408 ( .A1(u5_mult_82_n6774), .A2(u5_mult_82_net65675), 
        .ZN(u5_mult_82_ab_25__49_) );
  NOR2_X2 u5_mult_82_U1407 ( .A1(u5_mult_82_n6785), .A2(u5_mult_82_n6636), 
        .ZN(u5_mult_82_ab_22__47_) );
  NOR2_X2 u5_mult_82_U1406 ( .A1(u5_mult_82_n6780), .A2(u5_mult_82_n6551), 
        .ZN(u5_mult_82_ab_10__48_) );
  NOR2_X2 u5_mult_82_U1405 ( .A1(u5_mult_82_n6761), .A2(u5_mult_82_n6607), 
        .ZN(u5_mult_82_ab_18__51_) );
  NOR2_X2 u5_mult_82_U1404 ( .A1(u5_mult_82_n6775), .A2(u5_mult_82_net66087), 
        .ZN(u5_mult_82_ab_2__49_) );
  NOR2_X1 u5_mult_82_U1403 ( .A1(u5_mult_82_n6922), .A2(u5_mult_82_n6558), 
        .ZN(u5_mult_82_ab_11__18_) );
  NOR2_X2 u5_mult_82_U1402 ( .A1(u5_mult_82_n6922), .A2(u5_mult_82_n6522), 
        .ZN(u5_mult_82_ab_4__18_) );
  INV_X8 u5_mult_82_U1401 ( .A(u6_N2), .ZN(u5_mult_82_n6959) );
  INV_X4 u5_mult_82_U1400 ( .A(u5_mult_82_n6959), .ZN(u5_mult_82_n6965) );
  INV_X4 u5_mult_82_U1399 ( .A(u5_mult_82_n6965), .ZN(u5_mult_82_n6960) );
  NOR2_X2 u5_mult_82_U1398 ( .A1(u5_mult_82_n6953), .A2(u5_mult_82_net65519), 
        .ZN(u5_mult_82_ab_34__3_) );
  NOR2_X1 u5_mult_82_U1397 ( .A1(u5_mult_82_n6929), .A2(u5_mult_82_n6522), 
        .ZN(u5_mult_82_ab_4__17_) );
  NOR2_X2 u5_mult_82_U1396 ( .A1(u5_mult_82_n6898), .A2(u5_mult_82_n6522), 
        .ZN(u5_mult_82_ab_4__21_) );
  NOR2_X2 u5_mult_82_U1395 ( .A1(u5_mult_82_n6947), .A2(u5_mult_82_n6637), 
        .ZN(u5_mult_82_ab_22__4_) );
  NOR2_X2 u5_mult_82_U1394 ( .A1(u5_mult_82_n6947), .A2(u5_mult_82_n6658), 
        .ZN(u5_mult_82_ab_27__4_) );
  NOR2_X2 u5_mult_82_U1393 ( .A1(u5_mult_82_net64363), .A2(u5_mult_82_n6603), 
        .ZN(u5_mult_82_ab_17__5_) );
  NOR2_X1 u5_mult_82_U1392 ( .A1(u5_mult_82_n6940), .A2(u5_mult_82_n6673), 
        .ZN(u5_mult_82_ab_29__7_) );
  NOR2_X1 u5_mult_82_U1391 ( .A1(u5_mult_82_net64671), .A2(u5_mult_82_net66019), .ZN(u5_mult_82_ab_6__22_) );
  NOR2_X2 u5_mult_82_U1390 ( .A1(u5_mult_82_n6941), .A2(u5_mult_82_n6596), 
        .ZN(u5_mult_82_ab_16__7_) );
  NOR2_X2 u5_mult_82_U1389 ( .A1(u5_mult_82_net64563), .A2(u5_mult_82_n6522), 
        .ZN(u5_mult_82_ab_4__16_) );
  NOR2_X2 u5_mult_82_U1388 ( .A1(u5_mult_82_n6826), .A2(u5_mult_82_net65277), 
        .ZN(u5_mult_82_ab_47__40_) );
  INV_X16 u5_mult_82_U1387 ( .A(u5_mult_82_n1268), .ZN(u5_mult_82_n1267) );
  NOR2_X2 u5_mult_82_U1386 ( .A1(u5_mult_82_net64435), .A2(u5_mult_82_n6603), 
        .ZN(u5_mult_82_ab_17__9_) );
  NOR2_X2 u5_mult_82_U1385 ( .A1(u5_mult_82_n6772), .A2(u5_mult_82_net65277), 
        .ZN(u5_mult_82_ab_47__49_) );
  NOR2_X2 u5_mult_82_U1384 ( .A1(u5_mult_82_n6838), .A2(u5_mult_82_n6684), 
        .ZN(u5_mult_82_ab_31__33_) );
  NOR2_X2 u5_mult_82_U1383 ( .A1(u5_mult_82_net64883), .A2(u5_mult_82_n6684), 
        .ZN(u5_mult_82_ab_31__34_) );
  NOR2_X2 u5_mult_82_U1382 ( .A1(u5_mult_82_n6896), .A2(u5_mult_82_n6679), 
        .ZN(u5_mult_82_ab_30__21_) );
  NOR2_X1 u5_mult_82_U1381 ( .A1(u5_mult_82_net64437), .A2(u5_mult_82_n6559), 
        .ZN(u5_mult_82_ab_11__9_) );
  NOR2_X1 u5_mult_82_U1380 ( .A1(u5_mult_82_n6797), .A2(u5_mult_82_n6740), 
        .ZN(u5_mult_82_ab_46__45_) );
  NOR2_X1 u5_mult_82_U1379 ( .A1(u5_mult_82_net64455), .A2(u5_mult_82_n6559), 
        .ZN(u5_mult_82_ab_11__10_) );
  NOR2_X1 u5_mult_82_U1378 ( .A1(u5_mult_82_n6928), .A2(u5_mult_82_n6636), 
        .ZN(u5_mult_82_ab_22__17_) );
  NOR2_X2 u5_mult_82_U1377 ( .A1(u5_mult_82_net64935), .A2(u5_mult_82_net65369), .ZN(u5_mult_82_ab_42__37_) );
  NOR2_X1 u5_mult_82_U1376 ( .A1(u5_mult_82_net64509), .A2(u5_mult_82_n6552), 
        .ZN(u5_mult_82_ab_10__13_) );
  NOR2_X1 u5_mult_82_U1375 ( .A1(u5_mult_82_n6811), .A2(u5_mult_82_n6729), 
        .ZN(u5_mult_82_ab_39__43_) );
  NOR2_X1 u5_mult_82_U1374 ( .A1(u5_mult_82_n6816), .A2(u5_mult_82_n6729), 
        .ZN(u5_mult_82_ab_39__42_) );
  NOR2_X1 u5_mult_82_U1373 ( .A1(u5_mult_82_n6821), .A2(u5_mult_82_n6729), 
        .ZN(u5_mult_82_ab_39__41_) );
  NOR2_X2 u5_mult_82_U1372 ( .A1(u5_mult_82_n6877), .A2(u5_mult_82_n6566), 
        .ZN(u5_mult_82_ab_12__27_) );
  NOR2_X2 u5_mult_82_U1371 ( .A1(u5_mult_82_n6896), .A2(u5_mult_82_n6728), 
        .ZN(u5_mult_82_ab_39__21_) );
  NOR2_X2 u5_mult_82_U1370 ( .A1(u5_mult_82_net64667), .A2(u5_mult_82_n6728), 
        .ZN(u5_mult_82_ab_39__22_) );
  NOR2_X1 u5_mult_82_U1369 ( .A1(u5_mult_82_n6797), .A2(u5_mult_82_net65445), 
        .ZN(u5_mult_82_ab_38__45_) );
  NOR2_X1 u5_mult_82_U1368 ( .A1(u5_mult_82_n6791), .A2(u5_mult_82_net65445), 
        .ZN(u5_mult_82_ab_38__46_) );
  NOR2_X1 u5_mult_82_U1367 ( .A1(u5_mult_82_n6784), .A2(u5_mult_82_net65385), 
        .ZN(u5_mult_82_ab_41__47_) );
  NOR2_X1 u5_mult_82_U1366 ( .A1(u5_mult_82_n6845), .A2(u5_mult_82_n6557), 
        .ZN(u5_mult_82_ab_11__32_) );
  NOR2_X2 u5_mult_82_U1365 ( .A1(u5_mult_82_n6778), .A2(u5_mult_82_net65385), 
        .ZN(u5_mult_82_ab_41__48_) );
  NOR2_X1 u5_mult_82_U1364 ( .A1(u5_mult_82_n6915), .A2(u5_mult_82_n6572), 
        .ZN(u5_mult_82_ab_13__19_) );
  NOR2_X2 u5_mult_82_U1363 ( .A1(u5_mult_82_n6773), .A2(u5_mult_82_n6713), 
        .ZN(u5_mult_82_ab_36__49_) );
  NOR2_X2 u5_mult_82_U1362 ( .A1(u5_mult_82_net64689), .A2(u5_mult_82_n6536), 
        .ZN(u5_mult_82_ab_8__23_) );
  NOR2_X1 u5_mult_82_U1361 ( .A1(u5_mult_82_n6791), .A2(u5_mult_82_n6692), 
        .ZN(u5_mult_82_ab_32__46_) );
  NOR2_X1 u5_mult_82_U1360 ( .A1(u5_mult_82_n6804), .A2(u5_mult_82_n6677), 
        .ZN(u5_mult_82_ab_30__44_) );
  NOR2_X1 u5_mult_82_U1359 ( .A1(u5_mult_82_n6797), .A2(u5_mult_82_n6686), 
        .ZN(u5_mult_82_ab_31__45_) );
  NOR2_X2 u5_mult_82_U1358 ( .A1(u5_mult_82_n6845), .A2(u5_mult_82_n6514), 
        .ZN(u5_mult_82_ab_3__32_) );
  NOR2_X2 u5_mult_82_U1357 ( .A1(u5_mult_82_n6778), .A2(u5_mult_82_n6687), 
        .ZN(u5_mult_82_ab_31__48_) );
  NOR2_X1 u5_mult_82_U1356 ( .A1(u5_mult_82_n6806), .A2(u5_mult_82_n6513), 
        .ZN(u5_mult_82_ab_3__44_) );
  NOR2_X1 u5_mult_82_U1355 ( .A1(u5_mult_82_n6798), .A2(u5_mult_82_net65713), 
        .ZN(u5_mult_82_ab_23__45_) );
  NOR2_X2 u5_mult_82_U1354 ( .A1(u5_mult_82_n6768), .A2(u5_mult_82_n6641), 
        .ZN(u5_mult_82_ab_24__50_) );
  NOR2_X1 u5_mult_82_U1353 ( .A1(u5_mult_82_n6774), .A2(u5_mult_82_net65711), 
        .ZN(u5_mult_82_ab_23__49_) );
  NOR2_X2 u5_mult_82_U1352 ( .A1(u5_mult_82_n6780), .A2(u5_mult_82_n6543), 
        .ZN(u5_mult_82_ab_9__48_) );
  NOR2_X2 u5_mult_82_U1351 ( .A1(u5_mult_82_n6761), .A2(u5_mult_82_n6600), 
        .ZN(u5_mult_82_ab_17__51_) );
  XNOR2_X2 u5_mult_82_U1350 ( .A(u5_mult_82_ab_7__46_), .B(
        u5_mult_82_CARRYB_6__46_), .ZN(u5_mult_82_n572) );
  XNOR2_X2 u5_mult_82_U1349 ( .A(u5_mult_82_n572), .B(u5_mult_82_SUMB_6__47_), 
        .ZN(u5_mult_82_SUMB_7__46_) );
  NAND2_X2 u5_mult_82_U1348 ( .A1(u5_mult_82_CARRYB_46__15_), .A2(
        u5_mult_82_SUMB_46__16_), .ZN(u5_mult_82_n5851) );
  NAND2_X1 u5_mult_82_U1347 ( .A1(u5_mult_82_CARRYB_49__14_), .A2(
        u5_mult_82_SUMB_49__15_), .ZN(u5_mult_82_n5941) );
  INV_X1 u5_mult_82_U1346 ( .A(u5_mult_82_SUMB_49__15_), .ZN(u5_mult_82_n784)
         );
  NAND2_X1 u5_mult_82_U1345 ( .A1(u5_mult_82_n4362), .A2(
        u5_mult_82_SUMB_49__15_), .ZN(u5_mult_82_n785) );
  NAND2_X2 u5_mult_82_U1344 ( .A1(u5_mult_82_CARRYB_14__46_), .A2(
        u5_mult_82_SUMB_14__47_), .ZN(u5_mult_82_n4879) );
  NAND2_X2 u5_mult_82_U1343 ( .A1(u5_mult_82_CARRYB_33__32_), .A2(
        u5_mult_82_n74), .ZN(u5_mult_82_n2719) );
  NAND3_X4 u5_mult_82_U1342 ( .A1(u5_mult_82_n4400), .A2(u5_mult_82_n4399), 
        .A3(u5_mult_82_n4398), .ZN(u5_mult_82_CARRYB_50__17_) );
  NAND3_X2 u5_mult_82_U1341 ( .A1(u5_mult_82_n3636), .A2(u5_mult_82_n3637), 
        .A3(u5_mult_82_n3638), .ZN(u5_mult_82_CARRYB_49__17_) );
  NAND2_X2 u5_mult_82_U1340 ( .A1(u5_mult_82_ab_45__17_), .A2(
        u5_mult_82_SUMB_44__18_), .ZN(u5_mult_82_n4015) );
  NAND2_X1 u5_mult_82_U1339 ( .A1(u5_mult_82_ab_46__17_), .A2(
        u5_mult_82_CARRYB_45__17_), .ZN(u5_mult_82_n5861) );
  NAND2_X2 u5_mult_82_U1338 ( .A1(u5_mult_82_ab_21__34_), .A2(u5_mult_82_n1725), .ZN(u5_mult_82_n5543) );
  NAND2_X1 u5_mult_82_U1337 ( .A1(u5_mult_82_CARRYB_20__35_), .A2(
        u5_mult_82_SUMB_20__36_), .ZN(u5_mult_82_n4988) );
  NAND2_X1 u5_mult_82_U1336 ( .A1(u5_mult_82_ab_28__30_), .A2(
        u5_mult_82_SUMB_27__31_), .ZN(u5_mult_82_n3226) );
  NAND2_X1 u5_mult_82_U1335 ( .A1(u5_mult_82_SUMB_28__31_), .A2(
        u5_mult_82_CARRYB_28__30_), .ZN(u5_mult_82_n4536) );
  NAND2_X1 u5_mult_82_U1334 ( .A1(u5_mult_82_ab_48__18_), .A2(
        u5_mult_82_CARRYB_47__18_), .ZN(u5_mult_82_n5712) );
  NAND2_X1 u5_mult_82_U1333 ( .A1(u5_mult_82_ab_22__25_), .A2(
        u5_mult_82_CARRYB_21__25_), .ZN(u5_mult_82_n2192) );
  XNOR2_X2 u5_mult_82_U1332 ( .A(u5_mult_82_ab_19__33_), .B(
        u5_mult_82_CARRYB_18__33_), .ZN(u5_mult_82_n1463) );
  NAND3_X4 u5_mult_82_U1331 ( .A1(u5_mult_82_n6250), .A2(u5_mult_82_n6251), 
        .A3(u5_mult_82_n6252), .ZN(u5_mult_82_CARRYB_28__27_) );
  NAND2_X2 u5_mult_82_U1330 ( .A1(u5_mult_82_ab_33__26_), .A2(
        u5_mult_82_CARRYB_32__26_), .ZN(u5_mult_82_n3385) );
  NAND2_X4 u5_mult_82_U1329 ( .A1(u5_mult_82_ab_32__26_), .A2(u5_mult_82_n1500), .ZN(u5_mult_82_n3955) );
  NOR2_X1 u5_mult_82_U1328 ( .A1(u5_mult_82_net64685), .A2(u5_mult_82_net65443), .ZN(u5_mult_82_ab_38__23_) );
  NAND3_X4 u5_mult_82_U1327 ( .A1(u5_mult_82_n569), .A2(u5_mult_82_n570), .A3(
        u5_mult_82_n571), .ZN(u5_mult_82_CARRYB_40__21_) );
  NAND2_X2 u5_mult_82_U1326 ( .A1(u5_mult_82_CARRYB_39__21_), .A2(
        u5_mult_82_SUMB_39__22_), .ZN(u5_mult_82_n571) );
  NAND2_X2 u5_mult_82_U1325 ( .A1(u5_mult_82_ab_40__21_), .A2(
        u5_mult_82_SUMB_39__22_), .ZN(u5_mult_82_n570) );
  NAND2_X1 u5_mult_82_U1324 ( .A1(u5_mult_82_ab_40__21_), .A2(
        u5_mult_82_CARRYB_39__21_), .ZN(u5_mult_82_n569) );
  NAND3_X4 u5_mult_82_U1323 ( .A1(u5_mult_82_n566), .A2(u5_mult_82_n567), .A3(
        u5_mult_82_n568), .ZN(u5_mult_82_CARRYB_39__22_) );
  NAND2_X2 u5_mult_82_U1322 ( .A1(u5_mult_82_CARRYB_38__22_), .A2(
        u5_mult_82_SUMB_38__23_), .ZN(u5_mult_82_n568) );
  NAND2_X2 u5_mult_82_U1321 ( .A1(u5_mult_82_ab_39__22_), .A2(
        u5_mult_82_SUMB_38__23_), .ZN(u5_mult_82_n567) );
  NAND2_X2 u5_mult_82_U1320 ( .A1(u5_mult_82_ab_39__22_), .A2(
        u5_mult_82_CARRYB_38__22_), .ZN(u5_mult_82_n566) );
  XOR2_X2 u5_mult_82_U1319 ( .A(u5_mult_82_n565), .B(u5_mult_82_SUMB_38__23_), 
        .Z(u5_mult_82_SUMB_39__22_) );
  XOR2_X2 u5_mult_82_U1318 ( .A(u5_mult_82_ab_39__22_), .B(
        u5_mult_82_CARRYB_38__22_), .Z(u5_mult_82_n565) );
  NAND3_X2 u5_mult_82_U1317 ( .A1(u5_mult_82_n562), .A2(u5_mult_82_n563), .A3(
        u5_mult_82_n564), .ZN(u5_mult_82_CARRYB_38__23_) );
  NAND2_X2 u5_mult_82_U1316 ( .A1(u5_mult_82_ab_38__23_), .A2(
        u5_mult_82_CARRYB_37__23_), .ZN(u5_mult_82_n564) );
  NAND2_X1 u5_mult_82_U1315 ( .A1(u5_mult_82_CARRYB_37__23_), .A2(
        u5_mult_82_SUMB_37__24_), .ZN(u5_mult_82_n562) );
  XOR2_X2 u5_mult_82_U1314 ( .A(u5_mult_82_SUMB_37__24_), .B(u5_mult_82_n561), 
        .Z(u5_mult_82_SUMB_38__23_) );
  XOR2_X2 u5_mult_82_U1313 ( .A(u5_mult_82_CARRYB_37__23_), .B(
        u5_mult_82_ab_38__23_), .Z(u5_mult_82_n561) );
  NAND2_X2 u5_mult_82_U1312 ( .A1(u5_mult_82_ab_10__44_), .A2(
        u5_mult_82_SUMB_9__45_), .ZN(u5_mult_82_n6356) );
  NAND2_X2 u5_mult_82_U1311 ( .A1(u5_mult_82_CARRYB_45__6_), .A2(
        u5_mult_82_SUMB_45__7_), .ZN(u5_mult_82_n6168) );
  NAND2_X2 u5_mult_82_U1310 ( .A1(u5_mult_82_ab_47__10_), .A2(
        u5_mult_82_SUMB_46__11_), .ZN(u5_mult_82_n4181) );
  NAND2_X4 u5_mult_82_U1309 ( .A1(u5_mult_82_n1559), .A2(
        u5_mult_82_CARRYB_18__43_), .ZN(u5_mult_82_n5842) );
  NAND2_X2 u5_mult_82_U1308 ( .A1(u5_mult_82_ab_1__52_), .A2(u5_mult_82_n965), 
        .ZN(u5_mult_82_n901) );
  NAND2_X4 u5_mult_82_U1307 ( .A1(u5_mult_82_n1205), .A2(u5_mult_82_n1206), 
        .ZN(u5_mult_82_n2565) );
  XNOR2_X2 u5_mult_82_U1306 ( .A(u5_mult_82_CARRYB_43__11_), .B(
        u5_mult_82_ab_44__11_), .ZN(u5_mult_82_net79780) );
  NOR2_X2 u5_mult_82_U1305 ( .A1(u5_mult_82_net64505), .A2(u5_mult_82_n6729), 
        .ZN(u5_mult_82_ab_39__13_) );
  NOR2_X1 u5_mult_82_U1304 ( .A1(u5_mult_82_net64669), .A2(u5_mult_82_n6643), 
        .ZN(u5_mult_82_ab_24__22_) );
  NOR2_X2 u5_mult_82_U1303 ( .A1(u5_mult_82_n6892), .A2(u5_mult_82_n6636), 
        .ZN(u5_mult_82_ab_22__24_) );
  NAND3_X2 u5_mult_82_U1302 ( .A1(u5_mult_82_n558), .A2(u5_mult_82_n559), .A3(
        u5_mult_82_n560), .ZN(u5_mult_82_CARRYB_52__4_) );
  NAND2_X1 u5_mult_82_U1301 ( .A1(u5_mult_82_ab_52__4_), .A2(
        u5_mult_82_CARRYB_51__4_), .ZN(u5_mult_82_n560) );
  NAND2_X2 u5_mult_82_U1300 ( .A1(u5_mult_82_ab_52__4_), .A2(
        u5_mult_82_SUMB_51__5_), .ZN(u5_mult_82_n559) );
  NAND2_X1 u5_mult_82_U1299 ( .A1(u5_mult_82_CARRYB_51__4_), .A2(
        u5_mult_82_SUMB_51__5_), .ZN(u5_mult_82_n558) );
  XOR2_X2 u5_mult_82_U1298 ( .A(u5_mult_82_SUMB_51__5_), .B(u5_mult_82_n557), 
        .Z(u5_mult_82_SUMB_52__4_) );
  XOR2_X2 u5_mult_82_U1297 ( .A(u5_mult_82_CARRYB_51__4_), .B(
        u5_mult_82_ab_52__4_), .Z(u5_mult_82_n557) );
  INV_X1 u5_mult_82_U1296 ( .A(u5_mult_82_CARRYB_38__13_), .ZN(u5_mult_82_n554) );
  INV_X1 u5_mult_82_U1295 ( .A(u5_mult_82_ab_39__13_), .ZN(u5_mult_82_n553) );
  NAND2_X2 u5_mult_82_U1294 ( .A1(u5_mult_82_n555), .A2(u5_mult_82_n556), .ZN(
        u5_mult_82_n1284) );
  NAND2_X2 u5_mult_82_U1293 ( .A1(u5_mult_82_n553), .A2(
        u5_mult_82_CARRYB_38__13_), .ZN(u5_mult_82_n556) );
  NAND2_X2 u5_mult_82_U1292 ( .A1(u5_mult_82_ab_39__13_), .A2(u5_mult_82_n554), 
        .ZN(u5_mult_82_n555) );
  NAND3_X4 u5_mult_82_U1291 ( .A1(u5_mult_82_n550), .A2(u5_mult_82_n551), .A3(
        u5_mult_82_n552), .ZN(u5_mult_82_CARRYB_36__14_) );
  NAND2_X2 u5_mult_82_U1290 ( .A1(u5_mult_82_ab_36__14_), .A2(
        u5_mult_82_SUMB_35__15_), .ZN(u5_mult_82_n552) );
  NAND2_X2 u5_mult_82_U1289 ( .A1(u5_mult_82_CARRYB_35__14_), .A2(
        u5_mult_82_SUMB_35__15_), .ZN(u5_mult_82_n551) );
  NAND2_X1 u5_mult_82_U1288 ( .A1(u5_mult_82_CARRYB_35__14_), .A2(
        u5_mult_82_ab_36__14_), .ZN(u5_mult_82_n550) );
  NAND3_X4 u5_mult_82_U1287 ( .A1(u5_mult_82_n547), .A2(u5_mult_82_n548), .A3(
        u5_mult_82_n549), .ZN(u5_mult_82_CARRYB_35__15_) );
  NAND2_X2 u5_mult_82_U1286 ( .A1(u5_mult_82_CARRYB_34__15_), .A2(
        u5_mult_82_SUMB_34__16_), .ZN(u5_mult_82_n549) );
  NAND2_X2 u5_mult_82_U1285 ( .A1(u5_mult_82_ab_35__15_), .A2(
        u5_mult_82_SUMB_34__16_), .ZN(u5_mult_82_n548) );
  NAND2_X1 u5_mult_82_U1284 ( .A1(u5_mult_82_ab_35__15_), .A2(
        u5_mult_82_CARRYB_34__15_), .ZN(u5_mult_82_n547) );
  XOR2_X2 u5_mult_82_U1283 ( .A(u5_mult_82_n546), .B(u5_mult_82_SUMB_35__15_), 
        .Z(u5_mult_82_SUMB_36__14_) );
  XOR2_X2 u5_mult_82_U1282 ( .A(u5_mult_82_CARRYB_35__14_), .B(
        u5_mult_82_ab_36__14_), .Z(u5_mult_82_n546) );
  XOR2_X2 u5_mult_82_U1281 ( .A(u5_mult_82_n545), .B(u5_mult_82_SUMB_34__16_), 
        .Z(u5_mult_82_SUMB_35__15_) );
  XOR2_X2 u5_mult_82_U1280 ( .A(u5_mult_82_ab_35__15_), .B(
        u5_mult_82_CARRYB_34__15_), .Z(u5_mult_82_n545) );
  NAND3_X2 u5_mult_82_U1279 ( .A1(u5_mult_82_n542), .A2(u5_mult_82_n543), .A3(
        u5_mult_82_n544), .ZN(u5_mult_82_CARRYB_24__22_) );
  NAND2_X1 u5_mult_82_U1278 ( .A1(u5_mult_82_ab_24__22_), .A2(
        u5_mult_82_CARRYB_23__22_), .ZN(u5_mult_82_n544) );
  NAND2_X2 u5_mult_82_U1277 ( .A1(u5_mult_82_ab_24__22_), .A2(
        u5_mult_82_SUMB_23__23_), .ZN(u5_mult_82_n543) );
  NAND2_X1 u5_mult_82_U1276 ( .A1(u5_mult_82_CARRYB_23__22_), .A2(
        u5_mult_82_SUMB_23__23_), .ZN(u5_mult_82_n542) );
  XOR2_X2 u5_mult_82_U1275 ( .A(u5_mult_82_SUMB_23__23_), .B(u5_mult_82_n541), 
        .Z(u5_mult_82_SUMB_24__22_) );
  XOR2_X2 u5_mult_82_U1274 ( .A(u5_mult_82_CARRYB_23__22_), .B(
        u5_mult_82_ab_24__22_), .Z(u5_mult_82_n541) );
  INV_X1 u5_mult_82_U1273 ( .A(u5_mult_82_ab_22__24_), .ZN(u5_mult_82_n538) );
  INV_X4 u5_mult_82_U1272 ( .A(u5_mult_82_CARRYB_21__24_), .ZN(u5_mult_82_n537) );
  NAND2_X2 u5_mult_82_U1271 ( .A1(u5_mult_82_n539), .A2(u5_mult_82_n540), .ZN(
        u5_mult_82_n1348) );
  NAND2_X4 u5_mult_82_U1270 ( .A1(u5_mult_82_n537), .A2(u5_mult_82_n538), .ZN(
        u5_mult_82_n540) );
  NAND2_X1 u5_mult_82_U1269 ( .A1(u5_mult_82_CARRYB_21__24_), .A2(
        u5_mult_82_ab_22__24_), .ZN(u5_mult_82_n539) );
  NAND2_X2 u5_mult_82_U1268 ( .A1(u5_mult_82_n58), .A2(u5_mult_82_SUMB_31__28_), .ZN(u5_mult_82_n4545) );
  NAND2_X2 u5_mult_82_U1267 ( .A1(u5_mult_82_ab_6__37_), .A2(
        u5_mult_82_SUMB_5__38_), .ZN(u5_mult_82_n3291) );
  NAND2_X2 u5_mult_82_U1266 ( .A1(u5_mult_82_ab_8__36_), .A2(
        u5_mult_82_SUMB_7__37_), .ZN(u5_mult_82_n5622) );
  NAND2_X1 u5_mult_82_U1265 ( .A1(u5_mult_82_n3277), .A2(
        u5_mult_82_SUMB_7__37_), .ZN(u5_mult_82_n2737) );
  NAND2_X1 u5_mult_82_U1264 ( .A1(u5_mult_82_CARRYB_10__35_), .A2(
        u5_mult_82_SUMB_10__36_), .ZN(u5_mult_82_n4754) );
  CLKBUF_X3 u5_mult_82_U1263 ( .A(u5_mult_82_CARRYB_26__25_), .Z(
        u5_mult_82_n733) );
  NAND2_X1 u5_mult_82_U1262 ( .A1(u5_mult_82_CARRYB_44__13_), .A2(
        u5_mult_82_SUMB_44__14_), .ZN(u5_mult_82_n5463) );
  CLKBUF_X3 u5_mult_82_U1261 ( .A(u5_mult_82_SUMB_47__12_), .Z(
        u5_mult_82_n1541) );
  NAND2_X2 u5_mult_82_U1260 ( .A1(u5_mult_82_CARRYB_45__11_), .A2(
        u5_mult_82_SUMB_45__12_), .ZN(u5_mult_82_n5681) );
  NAND2_X1 u5_mult_82_U1259 ( .A1(u5_mult_82_CARRYB_47__35_), .A2(
        u5_mult_82_n1503), .ZN(u5_mult_82_n3091) );
  AND2_X2 u5_mult_82_U1258 ( .A1(u5_mult_82_SUMB_52__32_), .A2(
        u5_mult_82_CARRYB_52__31_), .ZN(u5_mult_82_n597) );
  XNOR2_X2 u5_mult_82_U1257 ( .A(u5_mult_82_SUMB_46__11_), .B(
        u5_mult_82_ab_47__10_), .ZN(u5_mult_82_n1696) );
  INV_X8 u5_mult_82_U1256 ( .A(u5_mult_82_net64217), .ZN(u5_mult_82_net86084)
         );
  XNOR2_X2 u5_mult_82_U1255 ( .A(u5_mult_82_ab_21__30_), .B(
        u5_mult_82_CARRYB_20__30_), .ZN(u5_mult_82_n1773) );
  XOR2_X2 u5_mult_82_U1254 ( .A(u5_mult_82_ab_10__50_), .B(
        u5_mult_82_CARRYB_9__50_), .Z(u5_mult_82_n1039) );
  NAND3_X4 u5_mult_82_U1253 ( .A1(u5_mult_82_n4911), .A2(u5_mult_82_n4912), 
        .A3(u5_mult_82_n4913), .ZN(u5_mult_82_CARRYB_51__19_) );
  XNOR2_X2 u5_mult_82_U1252 ( .A(u5_mult_82_ab_13__25_), .B(
        u5_mult_82_CARRYB_12__25_), .ZN(u5_mult_82_n536) );
  XNOR2_X2 u5_mult_82_U1251 ( .A(u5_mult_82_n536), .B(u5_mult_82_SUMB_12__26_), 
        .ZN(u5_mult_82_SUMB_13__25_) );
  NAND3_X4 u5_mult_82_U1250 ( .A1(u5_mult_82_n3388), .A2(u5_mult_82_n3389), 
        .A3(u5_mult_82_n3390), .ZN(u5_mult_82_CARRYB_34__25_) );
  NAND3_X2 u5_mult_82_U1249 ( .A1(u5_mult_82_n3956), .A2(u5_mult_82_n3955), 
        .A3(u5_mult_82_n3954), .ZN(u5_mult_82_CARRYB_32__26_) );
  NAND2_X1 u5_mult_82_U1248 ( .A1(u5_mult_82_CARRYB_3__34_), .A2(
        u5_mult_82_SUMB_3__35_), .ZN(u5_mult_82_net83295) );
  INV_X4 u5_mult_82_U1247 ( .A(u5_mult_82_n6408), .ZN(u5_mult_82_CLA_SUM[74])
         );
  NAND2_X1 u5_mult_82_U1246 ( .A1(u5_mult_82_CARRYB_20__22_), .A2(
        u5_mult_82_SUMB_20__23_), .ZN(u5_mult_82_n5498) );
  NAND2_X1 u5_mult_82_U1245 ( .A1(u5_mult_82_SUMB_25__20_), .A2(
        u5_mult_82_CARRYB_25__19_), .ZN(u5_mult_82_n3158) );
  INV_X4 u5_mult_82_U1244 ( .A(u5_mult_82_CARRYB_42__13_), .ZN(u5_mult_82_n533) );
  INV_X2 u5_mult_82_U1243 ( .A(u5_mult_82_ab_43__13_), .ZN(u5_mult_82_n532) );
  NAND2_X2 u5_mult_82_U1242 ( .A1(u5_mult_82_n534), .A2(u5_mult_82_n535), .ZN(
        u5_mult_82_n5520) );
  NAND2_X4 u5_mult_82_U1241 ( .A1(u5_mult_82_n532), .A2(u5_mult_82_n533), .ZN(
        u5_mult_82_n535) );
  NAND2_X2 u5_mult_82_U1240 ( .A1(u5_mult_82_ab_43__13_), .A2(
        u5_mult_82_CARRYB_42__13_), .ZN(u5_mult_82_n534) );
  NAND2_X4 u5_mult_82_U1239 ( .A1(u5_mult_82_SUMB_34__30_), .A2(
        u5_mult_82_ab_35__29_), .ZN(u5_mult_82_n1205) );
  CLKBUF_X3 u5_mult_82_U1238 ( .A(u5_mult_82_SUMB_15__46_), .Z(u5_mult_82_n531) );
  NAND3_X2 u5_mult_82_U1237 ( .A1(u5_mult_82_n528), .A2(u5_mult_82_n529), .A3(
        u5_mult_82_n530), .ZN(u5_mult_82_CARRYB_32__44_) );
  NAND2_X1 u5_mult_82_U1236 ( .A1(u5_mult_82_ab_32__44_), .A2(
        u5_mult_82_SUMB_31__45_), .ZN(u5_mult_82_n530) );
  NAND2_X1 u5_mult_82_U1235 ( .A1(u5_mult_82_ab_32__44_), .A2(
        u5_mult_82_CARRYB_31__44_), .ZN(u5_mult_82_n529) );
  NAND2_X1 u5_mult_82_U1234 ( .A1(u5_mult_82_SUMB_31__45_), .A2(
        u5_mult_82_CARRYB_31__44_), .ZN(u5_mult_82_n528) );
  XOR2_X2 u5_mult_82_U1233 ( .A(u5_mult_82_CARRYB_31__44_), .B(u5_mult_82_n527), .Z(u5_mult_82_SUMB_32__44_) );
  XOR2_X2 u5_mult_82_U1232 ( .A(u5_mult_82_SUMB_31__45_), .B(
        u5_mult_82_ab_32__44_), .Z(u5_mult_82_n527) );
  NAND3_X2 u5_mult_82_U1231 ( .A1(u5_mult_82_n524), .A2(u5_mult_82_n525), .A3(
        u5_mult_82_n526), .ZN(u5_mult_82_CARRYB_22__45_) );
  NAND2_X1 u5_mult_82_U1230 ( .A1(u5_mult_82_ab_22__45_), .A2(
        u5_mult_82_SUMB_21__46_), .ZN(u5_mult_82_n526) );
  NAND2_X2 u5_mult_82_U1229 ( .A1(u5_mult_82_ab_22__45_), .A2(
        u5_mult_82_CARRYB_21__45_), .ZN(u5_mult_82_n525) );
  NAND2_X2 u5_mult_82_U1228 ( .A1(u5_mult_82_SUMB_21__46_), .A2(
        u5_mult_82_CARRYB_21__45_), .ZN(u5_mult_82_n524) );
  XOR2_X2 u5_mult_82_U1227 ( .A(u5_mult_82_CARRYB_21__45_), .B(u5_mult_82_n523), .Z(u5_mult_82_SUMB_22__45_) );
  XOR2_X2 u5_mult_82_U1226 ( .A(u5_mult_82_SUMB_21__46_), .B(
        u5_mult_82_ab_22__45_), .Z(u5_mult_82_n523) );
  NAND3_X2 u5_mult_82_U1225 ( .A1(u5_mult_82_n520), .A2(u5_mult_82_n521), .A3(
        u5_mult_82_n522), .ZN(u5_mult_82_CARRYB_44__41_) );
  NAND2_X1 u5_mult_82_U1224 ( .A1(u5_mult_82_ab_44__41_), .A2(
        u5_mult_82_CARRYB_43__41_), .ZN(u5_mult_82_n522) );
  NAND2_X2 u5_mult_82_U1223 ( .A1(u5_mult_82_ab_44__41_), .A2(
        u5_mult_82_SUMB_43__42_), .ZN(u5_mult_82_n521) );
  NAND2_X1 u5_mult_82_U1222 ( .A1(u5_mult_82_CARRYB_43__41_), .A2(
        u5_mult_82_SUMB_43__42_), .ZN(u5_mult_82_n520) );
  XOR2_X2 u5_mult_82_U1221 ( .A(u5_mult_82_SUMB_43__42_), .B(u5_mult_82_n519), 
        .Z(u5_mult_82_SUMB_44__41_) );
  XOR2_X2 u5_mult_82_U1220 ( .A(u5_mult_82_CARRYB_43__41_), .B(
        u5_mult_82_ab_44__41_), .Z(u5_mult_82_n519) );
  NAND3_X2 u5_mult_82_U1219 ( .A1(u5_mult_82_n516), .A2(u5_mult_82_n517), .A3(
        u5_mult_82_n518), .ZN(u5_mult_82_CARRYB_50__38_) );
  NAND2_X1 u5_mult_82_U1218 ( .A1(u5_mult_82_CARRYB_49__38_), .A2(
        u5_mult_82_SUMB_49__39_), .ZN(u5_mult_82_n518) );
  NAND2_X1 u5_mult_82_U1217 ( .A1(u5_mult_82_ab_50__38_), .A2(
        u5_mult_82_SUMB_49__39_), .ZN(u5_mult_82_n517) );
  NAND2_X1 u5_mult_82_U1216 ( .A1(u5_mult_82_ab_50__38_), .A2(
        u5_mult_82_CARRYB_49__38_), .ZN(u5_mult_82_n516) );
  NAND3_X4 u5_mult_82_U1215 ( .A1(u5_mult_82_n513), .A2(u5_mult_82_n514), .A3(
        u5_mult_82_n515), .ZN(u5_mult_82_CARRYB_49__39_) );
  NAND2_X2 u5_mult_82_U1214 ( .A1(u5_mult_82_ab_49__39_), .A2(
        u5_mult_82_SUMB_48__40_), .ZN(u5_mult_82_n515) );
  NAND2_X2 u5_mult_82_U1213 ( .A1(u5_mult_82_CARRYB_48__39_), .A2(
        u5_mult_82_SUMB_48__40_), .ZN(u5_mult_82_n514) );
  NAND2_X1 u5_mult_82_U1212 ( .A1(u5_mult_82_CARRYB_48__39_), .A2(
        u5_mult_82_ab_49__39_), .ZN(u5_mult_82_n513) );
  XOR2_X2 u5_mult_82_U1211 ( .A(u5_mult_82_n512), .B(u5_mult_82_SUMB_49__39_), 
        .Z(u5_mult_82_SUMB_50__38_) );
  XOR2_X2 u5_mult_82_U1210 ( .A(u5_mult_82_ab_50__38_), .B(
        u5_mult_82_CARRYB_49__38_), .Z(u5_mult_82_n512) );
  XOR2_X2 u5_mult_82_U1209 ( .A(u5_mult_82_n511), .B(u5_mult_82_SUMB_48__40_), 
        .Z(u5_mult_82_SUMB_49__39_) );
  XOR2_X2 u5_mult_82_U1208 ( .A(u5_mult_82_CARRYB_48__39_), .B(
        u5_mult_82_ab_49__39_), .Z(u5_mult_82_n511) );
  INV_X1 u5_mult_82_U1207 ( .A(u5_mult_82_SUMB_24__46_), .ZN(u5_mult_82_n508)
         );
  INV_X4 u5_mult_82_U1206 ( .A(u5_mult_82_n1240), .ZN(u5_mult_82_n507) );
  NAND2_X2 u5_mult_82_U1205 ( .A1(u5_mult_82_n509), .A2(u5_mult_82_n510), .ZN(
        u5_mult_82_SUMB_25__45_) );
  NAND2_X2 u5_mult_82_U1204 ( .A1(u5_mult_82_n507), .A2(u5_mult_82_n508), .ZN(
        u5_mult_82_n510) );
  NAND2_X2 u5_mult_82_U1203 ( .A1(u5_mult_82_n1240), .A2(
        u5_mult_82_SUMB_24__46_), .ZN(u5_mult_82_n509) );
  NAND2_X1 u5_mult_82_U1202 ( .A1(u5_mult_82_CARRYB_39__31_), .A2(
        u5_mult_82_SUMB_39__32_), .ZN(u5_mult_82_n3085) );
  XNOR2_X2 u5_mult_82_U1201 ( .A(u5_mult_82_CARRYB_50__23_), .B(
        u5_mult_82_n1247), .ZN(u5_mult_82_SUMB_51__23_) );
  XNOR2_X2 u5_mult_82_U1200 ( .A(u5_mult_82_CARRYB_38__20_), .B(
        u5_mult_82_ab_39__20_), .ZN(u5_mult_82_n1391) );
  INV_X8 u5_mult_82_U1199 ( .A(u5_mult_82_n6405), .ZN(u5_mult_82_CLA_SUM[71])
         );
  NAND2_X1 u5_mult_82_U1198 ( .A1(u5_mult_82_CARRYB_27__42_), .A2(
        u5_mult_82_SUMB_27__43_), .ZN(u5_mult_82_n2179) );
  NAND2_X1 u5_mult_82_U1197 ( .A1(u5_mult_82_CARRYB_40__37_), .A2(
        u5_mult_82_SUMB_40__38_), .ZN(u5_mult_82_n955) );
  NAND2_X2 u5_mult_82_U1196 ( .A1(u5_mult_82_CARRYB_45__10_), .A2(
        u5_mult_82_SUMB_45__11_), .ZN(u5_mult_82_n6264) );
  NAND2_X4 u5_mult_82_U1195 ( .A1(u5_mult_82_CARRYB_37__18_), .A2(
        u5_mult_82_n741), .ZN(u5_mult_82_n4759) );
  XNOR2_X2 u5_mult_82_U1194 ( .A(u5_mult_82_n2330), .B(u5_mult_82_SUMB_45__27_), .ZN(u5_mult_82_SUMB_46__26_) );
  NAND2_X2 u5_mult_82_U1193 ( .A1(u5_mult_82_ab_41__28_), .A2(
        u5_mult_82_SUMB_40__29_), .ZN(u5_mult_82_n5583) );
  XOR2_X2 u5_mult_82_U1192 ( .A(u5_mult_82_n455), .B(u5_mult_82_n4281), .Z(
        u5_mult_82_SUMB_43__17_) );
  NAND3_X4 u5_mult_82_U1191 ( .A1(u5_mult_82_n5732), .A2(u5_mult_82_n5733), 
        .A3(u5_mult_82_n5734), .ZN(u5_mult_82_CARRYB_28__36_) );
  NAND2_X1 u5_mult_82_U1190 ( .A1(u5_mult_82_CARRYB_11__26_), .A2(
        u5_mult_82_SUMB_11__27_), .ZN(u5_mult_82_n2200) );
  NAND2_X1 u5_mult_82_U1189 ( .A1(u5_mult_82_SUMB_30__16_), .A2(
        u5_mult_82_CARRYB_30__15_), .ZN(u5_mult_82_n2000) );
  NAND2_X1 u5_mult_82_U1188 ( .A1(u5_mult_82_CARRYB_42__16_), .A2(
        u5_mult_82_n5283), .ZN(u5_mult_82_n5284) );
  NAND2_X1 u5_mult_82_U1187 ( .A1(u5_mult_82_CARRYB_48__12_), .A2(
        u5_mult_82_n1843), .ZN(u5_mult_82_n5990) );
  XNOR2_X2 u5_mult_82_U1186 ( .A(u5_mult_82_CARRYB_42__12_), .B(
        u5_mult_82_ab_43__12_), .ZN(u5_mult_82_n712) );
  NAND2_X2 u5_mult_82_U1185 ( .A1(u5_mult_82_CARRYB_42__12_), .A2(
        u5_mult_82_ab_43__12_), .ZN(u5_mult_82_n5004) );
  NAND3_X4 u5_mult_82_U1184 ( .A1(u5_mult_82_n504), .A2(u5_mult_82_n505), .A3(
        u5_mult_82_n506), .ZN(u5_mult_82_CARRYB_35__16_) );
  NAND2_X2 u5_mult_82_U1183 ( .A1(u5_mult_82_CARRYB_34__16_), .A2(
        u5_mult_82_SUMB_34__17_), .ZN(u5_mult_82_n506) );
  NAND2_X2 u5_mult_82_U1182 ( .A1(u5_mult_82_ab_35__16_), .A2(
        u5_mult_82_SUMB_34__17_), .ZN(u5_mult_82_n505) );
  NAND2_X1 u5_mult_82_U1181 ( .A1(u5_mult_82_ab_35__16_), .A2(
        u5_mult_82_CARRYB_34__16_), .ZN(u5_mult_82_n504) );
  NAND3_X2 u5_mult_82_U1180 ( .A1(u5_mult_82_n501), .A2(u5_mult_82_n502), .A3(
        u5_mult_82_n503), .ZN(u5_mult_82_CARRYB_34__17_) );
  NAND2_X2 u5_mult_82_U1179 ( .A1(u5_mult_82_CARRYB_33__17_), .A2(
        u5_mult_82_SUMB_33__18_), .ZN(u5_mult_82_n503) );
  NAND2_X2 u5_mult_82_U1178 ( .A1(u5_mult_82_ab_34__17_), .A2(
        u5_mult_82_SUMB_33__18_), .ZN(u5_mult_82_n502) );
  NAND2_X1 u5_mult_82_U1177 ( .A1(u5_mult_82_ab_34__17_), .A2(
        u5_mult_82_CARRYB_33__17_), .ZN(u5_mult_82_n501) );
  XOR2_X2 u5_mult_82_U1176 ( .A(u5_mult_82_ab_35__16_), .B(
        u5_mult_82_CARRYB_34__16_), .Z(u5_mult_82_n500) );
  XOR2_X2 u5_mult_82_U1175 ( .A(u5_mult_82_n499), .B(u5_mult_82_SUMB_33__18_), 
        .Z(u5_mult_82_SUMB_34__17_) );
  XOR2_X2 u5_mult_82_U1174 ( .A(u5_mult_82_ab_34__17_), .B(
        u5_mult_82_CARRYB_33__17_), .Z(u5_mult_82_n499) );
  NAND3_X2 u5_mult_82_U1173 ( .A1(u5_mult_82_n496), .A2(u5_mult_82_n497), .A3(
        u5_mult_82_n498), .ZN(u5_mult_82_CARRYB_42__12_) );
  NAND2_X1 u5_mult_82_U1172 ( .A1(u5_mult_82_ab_42__12_), .A2(
        u5_mult_82_CARRYB_41__12_), .ZN(u5_mult_82_n498) );
  NAND2_X2 u5_mult_82_U1171 ( .A1(u5_mult_82_ab_42__12_), .A2(
        u5_mult_82_SUMB_41__13_), .ZN(u5_mult_82_n497) );
  NAND2_X1 u5_mult_82_U1170 ( .A1(u5_mult_82_CARRYB_41__12_), .A2(
        u5_mult_82_SUMB_41__13_), .ZN(u5_mult_82_n496) );
  XOR2_X2 u5_mult_82_U1169 ( .A(u5_mult_82_SUMB_41__13_), .B(u5_mult_82_n495), 
        .Z(u5_mult_82_SUMB_42__12_) );
  XOR2_X2 u5_mult_82_U1168 ( .A(u5_mult_82_CARRYB_41__12_), .B(
        u5_mult_82_ab_42__12_), .Z(u5_mult_82_n495) );
  NAND2_X2 u5_mult_82_U1167 ( .A1(u5_mult_82_ab_29__19_), .A2(
        u5_mult_82_SUMB_28__20_), .ZN(u5_mult_82_n493) );
  NAND2_X1 u5_mult_82_U1166 ( .A1(u5_mult_82_ab_29__19_), .A2(
        u5_mult_82_CARRYB_28__19_), .ZN(u5_mult_82_n492) );
  NAND3_X4 u5_mult_82_U1165 ( .A1(u5_mult_82_n489), .A2(u5_mult_82_n490), .A3(
        u5_mult_82_n491), .ZN(u5_mult_82_CARRYB_28__20_) );
  NAND2_X2 u5_mult_82_U1164 ( .A1(u5_mult_82_SUMB_27__21_), .A2(
        u5_mult_82_CARRYB_27__20_), .ZN(u5_mult_82_n491) );
  NAND2_X2 u5_mult_82_U1163 ( .A1(u5_mult_82_ab_28__20_), .A2(
        u5_mult_82_CARRYB_27__20_), .ZN(u5_mult_82_n490) );
  NAND2_X2 u5_mult_82_U1162 ( .A1(u5_mult_82_ab_28__20_), .A2(
        u5_mult_82_SUMB_27__21_), .ZN(u5_mult_82_n489) );
  XOR2_X2 u5_mult_82_U1161 ( .A(u5_mult_82_n488), .B(u5_mult_82_SUMB_28__20_), 
        .Z(u5_mult_82_SUMB_29__19_) );
  XOR2_X2 u5_mult_82_U1160 ( .A(u5_mult_82_ab_29__19_), .B(
        u5_mult_82_CARRYB_28__19_), .Z(u5_mult_82_n488) );
  XOR2_X2 u5_mult_82_U1159 ( .A(u5_mult_82_n487), .B(u5_mult_82_CARRYB_27__20_), .Z(u5_mult_82_SUMB_28__20_) );
  XOR2_X2 u5_mult_82_U1158 ( .A(u5_mult_82_ab_28__20_), .B(
        u5_mult_82_SUMB_27__21_), .Z(u5_mult_82_n487) );
  NAND2_X2 u5_mult_82_U1157 ( .A1(u5_mult_82_ab_32__27_), .A2(
        u5_mult_82_SUMB_31__28_), .ZN(u5_mult_82_n4544) );
  NAND2_X4 u5_mult_82_U1156 ( .A1(u5_mult_82_ab_5__36_), .A2(
        u5_mult_82_CARRYB_4__36_), .ZN(u5_mult_82_n1366) );
  AND2_X2 u5_mult_82_U1155 ( .A1(u5_mult_82_SUMB_52__28_), .A2(
        u5_mult_82_CARRYB_52__27_), .ZN(u5_mult_82_n486) );
  AND2_X2 u5_mult_82_U1154 ( .A1(u5_mult_82_SUMB_52__27_), .A2(
        u5_mult_82_CARRYB_52__26_), .ZN(u5_mult_82_n485) );
  AND2_X2 u5_mult_82_U1153 ( .A1(u5_mult_82_SUMB_52__20_), .A2(
        u5_mult_82_CARRYB_52__19_), .ZN(u5_mult_82_n484) );
  NAND3_X4 u5_mult_82_U1152 ( .A1(u5_mult_82_n5756), .A2(u5_mult_82_n5757), 
        .A3(u5_mult_82_n5758), .ZN(u5_mult_82_n2112) );
  NAND3_X4 u5_mult_82_U1151 ( .A1(u5_mult_82_n6227), .A2(u5_mult_82_n6228), 
        .A3(u5_mult_82_n6229), .ZN(u5_mult_82_n4553) );
  XOR2_X2 u5_mult_82_U1150 ( .A(u5_mult_82_n500), .B(u5_mult_82_SUMB_34__17_), 
        .Z(u5_mult_82_n483) );
  NAND2_X4 u5_mult_82_U1149 ( .A1(u5_mult_82_ab_37__15_), .A2(
        u5_mult_82_CARRYB_36__15_), .ZN(u5_mult_82_n6176) );
  NAND3_X2 u5_mult_82_U1148 ( .A1(u5_mult_82_n4625), .A2(u5_mult_82_net81427), 
        .A3(u5_mult_82_net81428), .ZN(u5_mult_82_CARRYB_38__13_) );
  NAND3_X4 u5_mult_82_U1147 ( .A1(u5_mult_82_n6315), .A2(u5_mult_82_n6314), 
        .A3(u5_mult_82_n6313), .ZN(u5_mult_82_CARRYB_18__35_) );
  NAND2_X4 u5_mult_82_U1146 ( .A1(u5_mult_82_ab_31__19_), .A2(
        u5_mult_82_CARRYB_30__19_), .ZN(u5_mult_82_n2756) );
  NAND2_X4 u5_mult_82_U1145 ( .A1(u5_mult_82_ab_21__22_), .A2(
        u5_mult_82_CARRYB_20__22_), .ZN(u5_mult_82_n970) );
  XNOR2_X1 u5_mult_82_U1144 ( .A(u5_mult_82_SUMB_27__41_), .B(u5_mult_82_n1106), .ZN(u5_mult_82_n482) );
  XOR2_X2 u5_mult_82_U1143 ( .A(u5_mult_82_ab_1__43_), .B(u5_mult_82_ab_0__44_), .Z(u5_mult_82_n481) );
  AND2_X2 u5_mult_82_U1142 ( .A1(u5_mult_82_ab_0__2_), .A2(u5_mult_82_ab_1__1_), .ZN(u5_mult_82_n480) );
  XOR2_X1 u5_mult_82_U1141 ( .A(u5_mult_82_ab_1__1_), .B(u5_mult_82_ab_0__2_), 
        .Z(u5_mult_82_n479) );
  XOR2_X2 u5_mult_82_U1140 ( .A(u5_mult_82_ab_1__4_), .B(u5_mult_82_ab_0__5_), 
        .Z(u5_mult_82_n478) );
  AND2_X2 u5_mult_82_U1139 ( .A1(u5_mult_82_ab_0__9_), .A2(u5_mult_82_ab_1__8_), .ZN(u5_mult_82_n477) );
  XOR2_X1 u5_mult_82_U1138 ( .A(u5_mult_82_ab_1__10_), .B(u5_mult_82_ab_0__11_), .Z(u5_mult_82_n476) );
  AND2_X2 u5_mult_82_U1137 ( .A1(u5_mult_82_ab_0__16_), .A2(
        u5_mult_82_ab_1__15_), .ZN(u5_mult_82_n475) );
  AND2_X2 u5_mult_82_U1136 ( .A1(u5_mult_82_ab_0__23_), .A2(
        u5_mult_82_ab_1__22_), .ZN(u5_mult_82_n474) );
  XOR2_X2 u5_mult_82_U1135 ( .A(u5_mult_82_ab_1__21_), .B(u5_mult_82_ab_0__22_), .Z(u5_mult_82_n473) );
  AND2_X2 u5_mult_82_U1134 ( .A1(u5_mult_82_ab_0__21_), .A2(
        u5_mult_82_ab_1__20_), .ZN(u5_mult_82_n472) );
  AND2_X2 u5_mult_82_U1133 ( .A1(u5_mult_82_ab_0__18_), .A2(
        u5_mult_82_ab_1__17_), .ZN(u5_mult_82_n471) );
  INV_X32 u5_mult_82_U1132 ( .A(u5_mult_82_net66107), .ZN(u5_mult_82_net66121)
         );
  NOR2_X4 u5_mult_82_U1131 ( .A1(u5_mult_82_net64913), .A2(u5_mult_82_n1262), 
        .ZN(u5_mult_82_n2748) );
  AND2_X2 u5_mult_82_U1130 ( .A1(u5_mult_82_ab_0__29_), .A2(
        u5_mult_82_ab_1__28_), .ZN(u5_mult_82_n470) );
  XOR2_X2 u5_mult_82_U1129 ( .A(u5_mult_82_ab_1__28_), .B(u5_mult_82_ab_0__29_), .Z(u5_mult_82_n469) );
  AND2_X2 u5_mult_82_U1128 ( .A1(u5_mult_82_ab_0__41_), .A2(u5_mult_82_n3280), 
        .ZN(u5_mult_82_n467) );
  XOR2_X2 u5_mult_82_U1127 ( .A(u5_mult_82_ab_1__41_), .B(u5_mult_82_ab_0__42_), .Z(u5_mult_82_n466) );
  CLKBUF_X2 u5_mult_82_U1126 ( .A(u5_mult_82_CARRYB_44__27_), .Z(
        u5_mult_82_n465) );
  XNOR2_X2 u5_mult_82_U1125 ( .A(u5_mult_82_n464), .B(u5_mult_82_n2260), .ZN(
        u5_mult_82_SUMB_22__38_) );
  XNOR2_X2 u5_mult_82_U1124 ( .A(u5_mult_82_ab_39__18_), .B(
        u5_mult_82_CARRYB_38__18_), .ZN(u5_mult_82_n463) );
  XNOR2_X2 u5_mult_82_U1123 ( .A(u5_mult_82_n463), .B(u5_mult_82_n735), .ZN(
        u5_mult_82_SUMB_39__18_) );
  XNOR2_X2 u5_mult_82_U1122 ( .A(u5_mult_82_CARRYB_4__37_), .B(
        u5_mult_82_ab_5__37_), .ZN(u5_mult_82_n462) );
  XNOR2_X2 u5_mult_82_U1121 ( .A(u5_mult_82_n462), .B(u5_mult_82_SUMB_4__38_), 
        .ZN(u5_mult_82_SUMB_5__37_) );
  XNOR2_X2 u5_mult_82_U1120 ( .A(u5_mult_82_ab_9__29_), .B(
        u5_mult_82_CARRYB_8__29_), .ZN(u5_mult_82_n461) );
  XNOR2_X2 u5_mult_82_U1119 ( .A(u5_mult_82_ab_7__30_), .B(
        u5_mult_82_CARRYB_6__30_), .ZN(u5_mult_82_n460) );
  XNOR2_X2 u5_mult_82_U1118 ( .A(u5_mult_82_n460), .B(u5_mult_82_n1534), .ZN(
        u5_mult_82_SUMB_7__30_) );
  XNOR2_X2 u5_mult_82_U1117 ( .A(u5_mult_82_SUMB_23__30_), .B(
        u5_mult_82_CARRYB_23__29_), .ZN(u5_mult_82_n459) );
  XNOR2_X2 u5_mult_82_U1116 ( .A(u5_mult_82_n459), .B(u5_mult_82_ab_24__29_), 
        .ZN(u5_mult_82_SUMB_24__29_) );
  XNOR2_X2 u5_mult_82_U1115 ( .A(u5_mult_82_ab_51__19_), .B(
        u5_mult_82_CARRYB_50__19_), .ZN(u5_mult_82_n685) );
  XNOR2_X1 u5_mult_82_U1114 ( .A(u5_mult_82_SUMB_27__18_), .B(
        u5_mult_82_ab_28__17_), .ZN(u5_mult_82_n458) );
  XNOR2_X2 u5_mult_82_U1113 ( .A(u5_mult_82_CARRYB_27__17_), .B(
        u5_mult_82_n458), .ZN(u5_mult_82_SUMB_28__17_) );
  XNOR2_X1 u5_mult_82_U1112 ( .A(u5_mult_82_n879), .B(
        u5_mult_82_CARRYB_19__24_), .ZN(u5_mult_82_n5607) );
  CLKBUF_X2 u5_mult_82_U1111 ( .A(u5_mult_82_CARRYB_23__20_), .Z(
        u5_mult_82_n457) );
  XNOR2_X2 u5_mult_82_U1110 ( .A(u5_mult_82_ab_35__21_), .B(
        u5_mult_82_CARRYB_34__21_), .ZN(u5_mult_82_n456) );
  XNOR2_X2 u5_mult_82_U1109 ( .A(u5_mult_82_n456), .B(u5_mult_82_SUMB_34__22_), 
        .ZN(u5_mult_82_SUMB_35__21_) );
  INV_X4 u5_mult_82_U1108 ( .A(u5_mult_82_n138), .ZN(u5_mult_82_n455) );
  NAND2_X1 u5_mult_82_U1107 ( .A1(u5_mult_82_ab_16__24_), .A2(
        u5_mult_82_SUMB_15__25_), .ZN(u5_mult_82_n3331) );
  NAND2_X1 u5_mult_82_U1106 ( .A1(u5_mult_82_CARRYB_15__24_), .A2(
        u5_mult_82_SUMB_15__25_), .ZN(u5_mult_82_n3330) );
  XNOR2_X2 u5_mult_82_U1105 ( .A(u5_mult_82_ab_49__18_), .B(
        u5_mult_82_CARRYB_48__18_), .ZN(u5_mult_82_n454) );
  XNOR2_X2 u5_mult_82_U1104 ( .A(u5_mult_82_n454), .B(u5_mult_82_SUMB_48__19_), 
        .ZN(u5_mult_82_SUMB_49__18_) );
  XNOR2_X2 u5_mult_82_U1103 ( .A(u5_mult_82_ab_45__20_), .B(
        u5_mult_82_CARRYB_44__20_), .ZN(u5_mult_82_n453) );
  XNOR2_X2 u5_mult_82_U1102 ( .A(u5_mult_82_n453), .B(u5_mult_82_SUMB_44__21_), 
        .ZN(u5_mult_82_SUMB_45__20_) );
  XOR2_X2 u5_mult_82_U1101 ( .A(u5_mult_82_n3281), .B(
        u5_mult_82_CARRYB_23__21_), .Z(u5_mult_82_n452) );
  XNOR2_X2 u5_mult_82_U1100 ( .A(u5_mult_82_n452), .B(u5_mult_82_SUMB_23__22_), 
        .ZN(u5_mult_82_SUMB_24__21_) );
  XNOR2_X2 u5_mult_82_U1099 ( .A(u5_mult_82_CARRYB_48__19_), .B(
        u5_mult_82_ab_49__19_), .ZN(u5_mult_82_n451) );
  XNOR2_X2 u5_mult_82_U1098 ( .A(u5_mult_82_SUMB_48__20_), .B(u5_mult_82_n451), 
        .ZN(u5_mult_82_SUMB_49__19_) );
  XNOR2_X2 u5_mult_82_U1097 ( .A(u5_mult_82_ab_22__35_), .B(
        u5_mult_82_CARRYB_21__35_), .ZN(u5_mult_82_n450) );
  XNOR2_X2 u5_mult_82_U1096 ( .A(u5_mult_82_n450), .B(u5_mult_82_SUMB_21__36_), 
        .ZN(u5_mult_82_SUMB_22__35_) );
  XOR2_X2 u5_mult_82_U1095 ( .A(u5_mult_82_n4394), .B(u5_mult_82_SUMB_49__18_), 
        .Z(u5_mult_82_SUMB_50__17_) );
  NAND2_X2 u5_mult_82_U1094 ( .A1(u5_mult_82_ab_48__11_), .A2(
        u5_mult_82_SUMB_47__12_), .ZN(u5_mult_82_n6235) );
  XNOR2_X2 u5_mult_82_U1093 ( .A(u5_mult_82_ab_40__19_), .B(
        u5_mult_82_CARRYB_39__19_), .ZN(u5_mult_82_n449) );
  XNOR2_X2 u5_mult_82_U1092 ( .A(u5_mult_82_n449), .B(u5_mult_82_n427), .ZN(
        u5_mult_82_SUMB_40__19_) );
  INV_X4 u5_mult_82_U1091 ( .A(u5_mult_82_n447), .ZN(u5_mult_82_n448) );
  INV_X2 u5_mult_82_U1090 ( .A(u5_mult_82_SUMB_10__31_), .ZN(u5_mult_82_n447)
         );
  INV_X4 u5_mult_82_U1089 ( .A(u5_mult_82_n445), .ZN(u5_mult_82_n446) );
  INV_X2 u5_mult_82_U1088 ( .A(u5_mult_82_CARRYB_20__39_), .ZN(u5_mult_82_n445) );
  XNOR2_X1 u5_mult_82_U1087 ( .A(u5_mult_82_CARRYB_10__44_), .B(
        u5_mult_82_ab_11__44_), .ZN(u5_mult_82_n444) );
  XNOR2_X2 u5_mult_82_U1086 ( .A(u5_mult_82_SUMB_10__45_), .B(u5_mult_82_n444), 
        .ZN(u5_mult_82_SUMB_11__44_) );
  NAND2_X2 u5_mult_82_U1085 ( .A1(u5_mult_82_ab_45__34_), .A2(u5_mult_82_n42), 
        .ZN(u5_mult_82_n2608) );
  CLKBUF_X2 u5_mult_82_U1084 ( .A(u5_mult_82_SUMB_36__34_), .Z(u5_mult_82_n443) );
  INV_X4 u5_mult_82_U1083 ( .A(u5_mult_82_n441), .ZN(u5_mult_82_n442) );
  INV_X2 u5_mult_82_U1082 ( .A(u5_mult_82_SUMB_34__35_), .ZN(u5_mult_82_n441)
         );
  INV_X2 u5_mult_82_U1081 ( .A(u5_mult_82_n439), .ZN(u5_mult_82_n440) );
  INV_X2 u5_mult_82_U1080 ( .A(u5_mult_82_SUMB_15__44_), .ZN(u5_mult_82_n439)
         );
  NAND2_X2 u5_mult_82_U1079 ( .A1(u5_mult_82_ab_7__49_), .A2(
        u5_mult_82_SUMB_6__50_), .ZN(u5_mult_82_n5096) );
  INV_X4 u5_mult_82_U1078 ( .A(u5_mult_82_n437), .ZN(u5_mult_82_n438) );
  INV_X2 u5_mult_82_U1077 ( .A(u5_mult_82_SUMB_45__18_), .ZN(u5_mult_82_n437)
         );
  XNOR2_X1 u5_mult_82_U1076 ( .A(u5_mult_82_SUMB_6__50_), .B(
        u5_mult_82_ab_7__49_), .ZN(u5_mult_82_n436) );
  XNOR2_X2 u5_mult_82_U1075 ( .A(u5_mult_82_n1765), .B(u5_mult_82_n436), .ZN(
        u5_mult_82_SUMB_7__49_) );
  XNOR2_X2 u5_mult_82_U1074 ( .A(u5_mult_82_SUMB_5__51_), .B(
        u5_mult_82_ab_6__50_), .ZN(u5_mult_82_n435) );
  XOR2_X2 u5_mult_82_U1073 ( .A(u5_mult_82_CARRYB_42__20_), .B(
        u5_mult_82_n2172), .Z(u5_mult_82_n434) );
  XNOR2_X2 u5_mult_82_U1072 ( .A(u5_mult_82_SUMB_42__21_), .B(u5_mult_82_n434), 
        .ZN(u5_mult_82_SUMB_43__20_) );
  INV_X4 u5_mult_82_U1071 ( .A(u5_mult_82_n432), .ZN(u5_mult_82_n433) );
  INV_X2 u5_mult_82_U1070 ( .A(u5_mult_82_SUMB_23__33_), .ZN(u5_mult_82_n432)
         );
  NAND2_X1 u5_mult_82_U1069 ( .A1(u5_mult_82_CARRYB_19__16_), .A2(
        u5_mult_82_SUMB_19__17_), .ZN(u5_mult_82_n2842) );
  INV_X4 u5_mult_82_U1068 ( .A(u5_mult_82_n430), .ZN(u5_mult_82_n431) );
  INV_X2 u5_mult_82_U1067 ( .A(u5_mult_82_SUMB_28__18_), .ZN(u5_mult_82_n430)
         );
  XOR2_X2 u5_mult_82_U1066 ( .A(u5_mult_82_n2262), .B(
        u5_mult_82_CARRYB_15__26_), .Z(u5_mult_82_n429) );
  XNOR2_X2 u5_mult_82_U1065 ( .A(u5_mult_82_n429), .B(u5_mult_82_net86785), 
        .ZN(u5_mult_82_SUMB_16__26_) );
  NAND2_X1 u5_mult_82_U1064 ( .A1(u5_mult_82_SUMB_12__50_), .A2(
        u5_mult_82_CARRYB_12__49_), .ZN(u5_mult_82_n1200) );
  NAND2_X1 u5_mult_82_U1063 ( .A1(u5_mult_82_ab_13__49_), .A2(
        u5_mult_82_CARRYB_12__49_), .ZN(u5_mult_82_n1201) );
  NAND2_X1 u5_mult_82_U1062 ( .A1(u5_mult_82_ab_10__50_), .A2(
        u5_mult_82_CARRYB_9__50_), .ZN(u5_mult_82_n1041) );
  NAND2_X1 u5_mult_82_U1061 ( .A1(u5_mult_82_CARRYB_9__50_), .A2(
        u5_mult_82_SUMB_9__51_), .ZN(u5_mult_82_n1043) );
  NAND2_X1 u5_mult_82_U1060 ( .A1(u5_mult_82_ab_26__20_), .A2(
        u5_mult_82_SUMB_25__21_), .ZN(u5_mult_82_n4585) );
  XOR2_X2 u5_mult_82_U1059 ( .A(u5_mult_82_n397), .B(u5_mult_82_n2816), .Z(
        u5_mult_82_SUMB_24__12_) );
  NAND2_X2 u5_mult_82_U1058 ( .A1(u5_mult_82_ab_50__27_), .A2(
        u5_mult_82_CARRYB_49__27_), .ZN(u5_mult_82_n3751) );
  NAND2_X1 u5_mult_82_U1057 ( .A1(u5_mult_82_CARRYB_49__27_), .A2(
        u5_mult_82_SUMB_49__28_), .ZN(u5_mult_82_n3753) );
  NAND2_X1 u5_mult_82_U1056 ( .A1(u5_mult_82_ab_27__41_), .A2(
        u5_mult_82_CARRYB_26__41_), .ZN(u5_mult_82_n928) );
  NAND2_X1 u5_mult_82_U1055 ( .A1(u5_mult_82_CARRYB_26__41_), .A2(
        u5_mult_82_SUMB_26__42_), .ZN(u5_mult_82_n926) );
  XNOR2_X2 u5_mult_82_U1054 ( .A(u5_mult_82_SUMB_33__11_), .B(u5_mult_82_n428), 
        .ZN(u5_mult_82_SUMB_34__10_) );
  XOR2_X2 u5_mult_82_U1053 ( .A(u5_mult_82_ab_26__30_), .B(
        u5_mult_82_CARRYB_25__30_), .Z(u5_mult_82_n6278) );
  NOR2_X2 u5_mult_82_U1052 ( .A1(u5_mult_82_n6762), .A2(u5_mult_82_n1359), 
        .ZN(u5_mult_82_ab_6__51_) );
  NOR2_X4 u5_mult_82_U1051 ( .A1(u5_mult_82_n6762), .A2(u5_mult_82_net66033), 
        .ZN(u5_mult_82_ab_5__51_) );
  NOR2_X4 u5_mult_82_U1050 ( .A1(u5_mult_82_n6762), .A2(u5_mult_82_n6520), 
        .ZN(u5_mult_82_ab_4__51_) );
  NOR2_X4 u5_mult_82_U1049 ( .A1(u5_mult_82_n6762), .A2(u5_mult_82_n6513), 
        .ZN(u5_mult_82_ab_3__51_) );
  INV_X16 u5_mult_82_U1048 ( .A(u5_mult_82_n6763), .ZN(u5_mult_82_n6762) );
  XOR2_X1 u5_mult_82_U1047 ( .A(u5_mult_82_ab_29__28_), .B(
        u5_mult_82_CARRYB_28__28_), .Z(u5_mult_82_n2351) );
  NAND2_X1 u5_mult_82_U1046 ( .A1(u5_mult_82_CARRYB_28__28_), .A2(
        u5_mult_82_SUMB_28__29_), .ZN(u5_mult_82_n2354) );
  NAND2_X1 u5_mult_82_U1045 ( .A1(u5_mult_82_n5552), .A2(
        u5_mult_82_SUMB_15__45_), .ZN(u5_mult_82_n6130) );
  NAND2_X1 u5_mult_82_U1044 ( .A1(u5_mult_82_ab_5__50_), .A2(
        u5_mult_82_SUMB_4__51_), .ZN(u5_mult_82_n6292) );
  INV_X4 u5_mult_82_U1043 ( .A(u5_mult_82_n426), .ZN(u5_mult_82_n427) );
  XNOR2_X2 u5_mult_82_U1042 ( .A(u5_mult_82_SUMB_36__22_), .B(
        u5_mult_82_ab_37__21_), .ZN(u5_mult_82_n425) );
  XNOR2_X2 u5_mult_82_U1041 ( .A(u5_mult_82_CARRYB_36__21_), .B(
        u5_mult_82_n425), .ZN(u5_mult_82_SUMB_37__21_) );
  INV_X4 u5_mult_82_U1040 ( .A(u5_mult_82_n423), .ZN(u5_mult_82_n424) );
  INV_X2 u5_mult_82_U1039 ( .A(u5_mult_82_CARRYB_13__47_), .ZN(u5_mult_82_n423) );
  XOR2_X2 u5_mult_82_U1038 ( .A(u5_mult_82_CARRYB_30__13_), .B(
        u5_mult_82_ab_31__13_), .Z(u5_mult_82_n651) );
  INV_X8 u5_mult_82_U1037 ( .A(u5_mult_82_n420), .ZN(u5_mult_82_n421) );
  INV_X2 u5_mult_82_U1036 ( .A(u5_mult_82_CARRYB_14__38_), .ZN(u5_mult_82_n420) );
  NAND2_X2 u5_mult_82_U1035 ( .A1(u5_mult_82_ab_35__21_), .A2(
        u5_mult_82_SUMB_34__22_), .ZN(u5_mult_82_n4246) );
  NAND2_X2 u5_mult_82_U1034 ( .A1(u5_mult_82_ab_50__20_), .A2(
        u5_mult_82_CARRYB_49__20_), .ZN(u5_mult_82_n4908) );
  XOR2_X2 u5_mult_82_U1033 ( .A(u5_mult_82_ab_32__31_), .B(
        u5_mult_82_CARRYB_31__31_), .Z(u5_mult_82_n419) );
  XNOR2_X2 u5_mult_82_U1032 ( .A(u5_mult_82_n419), .B(u5_mult_82_n1799), .ZN(
        u5_mult_82_SUMB_32__31_) );
  XNOR2_X2 u5_mult_82_U1031 ( .A(u5_mult_82_ab_32__27_), .B(u5_mult_82_n58), 
        .ZN(u5_mult_82_n2413) );
  NAND2_X2 u5_mult_82_U1030 ( .A1(u5_mult_82_ab_32__27_), .A2(u5_mult_82_n58), 
        .ZN(u5_mult_82_n4543) );
  INV_X32 u5_mult_82_U1029 ( .A(u5_mult_82_ab_12__47_), .ZN(u5_mult_82_n418)
         );
  XNOR2_X2 u5_mult_82_U1028 ( .A(u5_mult_82_CARRYB_11__47_), .B(
        u5_mult_82_n418), .ZN(u5_mult_82_n4587) );
  CLKBUF_X2 u5_mult_82_U1027 ( .A(u5_mult_82_SUMB_43__5_), .Z(u5_mult_82_n417)
         );
  INV_X4 u5_mult_82_U1026 ( .A(u5_mult_82_n415), .ZN(u5_mult_82_n416) );
  INV_X2 u5_mult_82_U1025 ( .A(u5_mult_82_CARRYB_14__50_), .ZN(u5_mult_82_n415) );
  XNOR2_X2 u5_mult_82_U1024 ( .A(u5_mult_82_ab_42__14_), .B(
        u5_mult_82_CARRYB_41__14_), .ZN(u5_mult_82_n414) );
  XNOR2_X2 u5_mult_82_U1023 ( .A(u5_mult_82_n414), .B(u5_mult_82_SUMB_41__15_), 
        .ZN(u5_mult_82_SUMB_42__14_) );
  NAND2_X1 u5_mult_82_U1022 ( .A1(u5_mult_82_SUMB_50__24_), .A2(
        u5_mult_82_CARRYB_50__23_), .ZN(u5_mult_82_n4456) );
  NAND2_X1 u5_mult_82_U1021 ( .A1(u5_mult_82_CARRYB_19__42_), .A2(
        u5_mult_82_SUMB_19__43_), .ZN(u5_mult_82_n5845) );
  XNOR2_X2 u5_mult_82_U1020 ( .A(u5_mult_82_ab_49__25_), .B(
        u5_mult_82_CARRYB_48__25_), .ZN(u5_mult_82_n413) );
  XNOR2_X2 u5_mult_82_U1019 ( .A(u5_mult_82_n413), .B(u5_mult_82_n1663), .ZN(
        u5_mult_82_SUMB_49__25_) );
  CLKBUF_X3 u5_mult_82_U1018 ( .A(u5_mult_82_SUMB_50__23_), .Z(
        u5_mult_82_n1434) );
  NAND2_X1 u5_mult_82_U1017 ( .A1(u5_mult_82_ab_34__11_), .A2(
        u5_mult_82_SUMB_33__12_), .ZN(u5_mult_82_n3578) );
  XNOR2_X1 u5_mult_82_U1016 ( .A(u5_mult_82_SUMB_33__12_), .B(u5_mult_82_n2118), .ZN(u5_mult_82_SUMB_34__11_) );
  XNOR2_X2 u5_mult_82_U1015 ( .A(u5_mult_82_CARRYB_24__15_), .B(
        u5_mult_82_ab_25__15_), .ZN(u5_mult_82_n782) );
  NAND2_X2 u5_mult_82_U1014 ( .A1(u5_mult_82_SUMB_28__31_), .A2(
        u5_mult_82_ab_29__30_), .ZN(u5_mult_82_n4535) );
  NAND2_X2 u5_mult_82_U1013 ( .A1(u5_mult_82_ab_2__51_), .A2(
        u5_mult_82_ab_1__52_), .ZN(u5_mult_82_n900) );
  NAND3_X1 u5_mult_82_U1012 ( .A1(u5_mult_82_n899), .A2(u5_mult_82_n900), .A3(
        u5_mult_82_n901), .ZN(u5_mult_82_n411) );
  XNOR2_X2 u5_mult_82_U1011 ( .A(u5_mult_82_n639), .B(u5_mult_82_SUMB_39__33_), 
        .ZN(u5_mult_82_SUMB_40__32_) );
  NAND2_X1 u5_mult_82_U1010 ( .A1(u5_mult_82_ab_41__31_), .A2(
        u5_mult_82_SUMB_40__32_), .ZN(u5_mult_82_n3089) );
  NAND2_X2 u5_mult_82_U1009 ( .A1(u5_mult_82_CARRYB_43__12_), .A2(
        u5_mult_82_SUMB_43__13_), .ZN(u5_mult_82_n5406) );
  NAND2_X1 u5_mult_82_U1008 ( .A1(u5_mult_82_ab_44__26_), .A2(
        u5_mult_82_SUMB_43__27_), .ZN(u5_mult_82_n4922) );
  XNOR2_X2 u5_mult_82_U1007 ( .A(u5_mult_82_ab_52__19_), .B(
        u5_mult_82_CARRYB_51__19_), .ZN(u5_mult_82_n409) );
  XNOR2_X2 u5_mult_82_U1006 ( .A(u5_mult_82_n409), .B(u5_mult_82_SUMB_51__20_), 
        .ZN(u5_mult_82_SUMB_52__19_) );
  XNOR2_X2 u5_mult_82_U1005 ( .A(u5_mult_82_net83142), .B(
        u5_mult_82_SUMB_44__10_), .ZN(u5_mult_82_SUMB_45__9_) );
  XNOR2_X2 u5_mult_82_U1004 ( .A(u5_mult_82_ab_45__26_), .B(
        u5_mult_82_CARRYB_44__26_), .ZN(u5_mult_82_n408) );
  XNOR2_X2 u5_mult_82_U1003 ( .A(u5_mult_82_n408), .B(u5_mult_82_SUMB_44__27_), 
        .ZN(u5_mult_82_SUMB_45__26_) );
  CLKBUF_X2 u5_mult_82_U1002 ( .A(u5_mult_82_CARRYB_49__18_), .Z(
        u5_mult_82_n407) );
  NAND3_X2 u5_mult_82_U1001 ( .A1(u5_mult_82_n4695), .A2(u5_mult_82_n4696), 
        .A3(u5_mult_82_n4697), .ZN(u5_mult_82_n406) );
  INV_X32 u5_mult_82_U1000 ( .A(u5_mult_82_ab_52__11_), .ZN(u5_mult_82_n405)
         );
  XNOR2_X2 u5_mult_82_U999 ( .A(u5_mult_82_CARRYB_51__11_), .B(u5_mult_82_n405), .ZN(u5_mult_82_n4698) );
  XNOR2_X2 u5_mult_82_U998 ( .A(u5_mult_82_n1514), .B(u5_mult_82_ab_33__10_), 
        .ZN(u5_mult_82_n1506) );
  XOR2_X2 u5_mult_82_U997 ( .A(u5_mult_82_n2418), .B(u5_mult_82_CARRYB_3__37_), 
        .Z(u5_mult_82_n404) );
  XNOR2_X2 u5_mult_82_U996 ( .A(u5_mult_82_n404), .B(u5_mult_82_SUMB_3__38_), 
        .ZN(u5_mult_82_SUMB_4__37_) );
  NAND2_X2 u5_mult_82_U995 ( .A1(u5_mult_82_SUMB_37__16_), .A2(
        u5_mult_82_ab_38__15_), .ZN(u5_mult_82_n3881) );
  NAND2_X2 u5_mult_82_U994 ( .A1(u5_mult_82_SUMB_37__16_), .A2(
        u5_mult_82_CARRYB_37__15_), .ZN(u5_mult_82_n3882) );
  NAND3_X4 u5_mult_82_U993 ( .A1(u5_mult_82_n3880), .A2(u5_mult_82_n3881), 
        .A3(u5_mult_82_n3882), .ZN(u5_mult_82_CARRYB_38__15_) );
  INV_X8 u5_mult_82_U992 ( .A(u5_mult_82_n6415), .ZN(u5_mult_82_CLA_CARRY[81])
         );
  XNOR2_X2 u5_mult_82_U991 ( .A(u5_mult_82_CARRYB_49__15_), .B(
        u5_mult_82_ab_50__15_), .ZN(u5_mult_82_n403) );
  XNOR2_X2 u5_mult_82_U990 ( .A(u5_mult_82_SUMB_49__16_), .B(u5_mult_82_n403), 
        .ZN(u5_mult_82_SUMB_50__15_) );
  NAND3_X2 u5_mult_82_U989 ( .A1(u5_mult_82_n5946), .A2(u5_mult_82_n5947), 
        .A3(u5_mult_82_n5948), .ZN(u5_mult_82_CARRYB_33__31_) );
  XNOR2_X2 u5_mult_82_U988 ( .A(u5_mult_82_n3074), .B(u5_mult_82_ab_29__21_), 
        .ZN(u5_mult_82_n2753) );
  XNOR2_X2 u5_mult_82_U987 ( .A(u5_mult_82_n1708), .B(u5_mult_82_ab_23__40_), 
        .ZN(u5_mult_82_n401) );
  XNOR2_X2 u5_mult_82_U986 ( .A(u5_mult_82_n401), .B(u5_mult_82_CARRYB_22__40_), .ZN(u5_mult_82_SUMB_23__40_) );
  XNOR2_X2 u5_mult_82_U985 ( .A(u5_mult_82_ab_16__43_), .B(
        u5_mult_82_CARRYB_15__43_), .ZN(u5_mult_82_n400) );
  XNOR2_X2 u5_mult_82_U984 ( .A(u5_mult_82_n400), .B(u5_mult_82_n440), .ZN(
        u5_mult_82_SUMB_16__43_) );
  INV_X4 u5_mult_82_U983 ( .A(u5_mult_82_n398), .ZN(u5_mult_82_n399) );
  INV_X2 u5_mult_82_U982 ( .A(u5_mult_82_SUMB_28__10_), .ZN(u5_mult_82_n398)
         );
  INV_X4 u5_mult_82_U981 ( .A(u5_mult_82_n396), .ZN(u5_mult_82_n397) );
  INV_X2 u5_mult_82_U980 ( .A(u5_mult_82_SUMB_23__13_), .ZN(u5_mult_82_n396)
         );
  XNOR2_X2 u5_mult_82_U979 ( .A(u5_mult_82_ab_33__11_), .B(
        u5_mult_82_CARRYB_32__11_), .ZN(u5_mult_82_n395) );
  XNOR2_X2 u5_mult_82_U978 ( .A(u5_mult_82_n395), .B(u5_mult_82_SUMB_32__12_), 
        .ZN(u5_mult_82_SUMB_33__11_) );
  INV_X8 u5_mult_82_U977 ( .A(u5_mult_82_n393), .ZN(u5_mult_82_n394) );
  INV_X4 u5_mult_82_U976 ( .A(u5_mult_82_CARRYB_27__13_), .ZN(u5_mult_82_n393)
         );
  NAND2_X1 u5_mult_82_U975 ( .A1(u5_mult_82_CARRYB_36__10_), .A2(
        u5_mult_82_SUMB_36__11_), .ZN(u5_mult_82_n988) );
  XNOR2_X2 u5_mult_82_U974 ( .A(u5_mult_82_ab_16__20_), .B(
        u5_mult_82_CARRYB_15__20_), .ZN(u5_mult_82_n2129) );
  NAND2_X2 u5_mult_82_U973 ( .A1(u5_mult_82_ab_41__12_), .A2(
        u5_mult_82_CARRYB_40__12_), .ZN(u5_mult_82_net86288) );
  NAND2_X1 u5_mult_82_U972 ( .A1(u5_mult_82_ab_39__13_), .A2(
        u5_mult_82_SUMB_38__14_), .ZN(u5_mult_82_net82468) );
  NAND2_X1 u5_mult_82_U971 ( .A1(u5_mult_82_CARRYB_38__13_), .A2(
        u5_mult_82_SUMB_38__14_), .ZN(u5_mult_82_net82469) );
  CLKBUF_X3 u5_mult_82_U970 ( .A(u5_mult_82_SUMB_38__14_), .Z(u5_mult_82_n1286) );
  XNOR2_X2 u5_mult_82_U969 ( .A(u5_mult_82_CARRYB_45__2_), .B(
        u5_mult_82_ab_46__2_), .ZN(u5_mult_82_n746) );
  NAND3_X4 u5_mult_82_U968 ( .A1(u5_mult_82_n5628), .A2(u5_mult_82_n5629), 
        .A3(u5_mult_82_n5630), .ZN(u5_mult_82_CARRYB_45__2_) );
  INV_X4 u5_mult_82_U967 ( .A(u5_mult_82_n391), .ZN(u5_mult_82_n392) );
  INV_X4 u5_mult_82_U966 ( .A(u5_mult_82_SUMB_13__22_), .ZN(u5_mult_82_n391)
         );
  NAND2_X1 u5_mult_82_U965 ( .A1(u5_mult_82_ab_34__14_), .A2(
        u5_mult_82_SUMB_33__15_), .ZN(u5_mult_82_n4952) );
  INV_X4 u5_mult_82_U964 ( .A(u5_mult_82_n389), .ZN(u5_mult_82_n390) );
  INV_X2 u5_mult_82_U963 ( .A(u5_mult_82_SUMB_36__5_), .ZN(u5_mult_82_n389) );
  CLKBUF_X2 u5_mult_82_U962 ( .A(u5_mult_82_CARRYB_32__9_), .Z(u5_mult_82_n388) );
  XNOR2_X2 u5_mult_82_U961 ( .A(u5_mult_82_ab_21__14_), .B(
        u5_mult_82_CARRYB_20__14_), .ZN(u5_mult_82_n387) );
  XNOR2_X2 u5_mult_82_U960 ( .A(u5_mult_82_n387), .B(u5_mult_82_n1717), .ZN(
        u5_mult_82_SUMB_21__14_) );
  XNOR2_X2 u5_mult_82_U959 ( .A(u5_mult_82_ab_4__26_), .B(
        u5_mult_82_CARRYB_3__26_), .ZN(u5_mult_82_n386) );
  XNOR2_X2 u5_mult_82_U958 ( .A(u5_mult_82_n386), .B(u5_mult_82_SUMB_3__27_), 
        .ZN(u5_mult_82_SUMB_4__26_) );
  XNOR2_X2 u5_mult_82_U957 ( .A(u5_mult_82_ab_6__28_), .B(
        u5_mult_82_CARRYB_5__28_), .ZN(u5_mult_82_n385) );
  XNOR2_X2 u5_mult_82_U956 ( .A(u5_mult_82_n385), .B(u5_mult_82_SUMB_5__29_), 
        .ZN(u5_mult_82_SUMB_6__28_) );
  XNOR2_X2 u5_mult_82_U955 ( .A(u5_mult_82_CARRYB_4__29_), .B(
        u5_mult_82_ab_5__29_), .ZN(u5_mult_82_n384) );
  XNOR2_X2 u5_mult_82_U954 ( .A(u5_mult_82_n380), .B(u5_mult_82_n384), .ZN(
        u5_mult_82_SUMB_5__29_) );
  NAND2_X2 u5_mult_82_U953 ( .A1(u5_mult_82_ab_46__6_), .A2(
        u5_mult_82_SUMB_45__7_), .ZN(u5_mult_82_n6167) );
  NAND2_X2 u5_mult_82_U952 ( .A1(u5_mult_82_CARRYB_38__7_), .A2(
        u5_mult_82_SUMB_38__8_), .ZN(u5_mult_82_n2989) );
  INV_X2 u5_mult_82_U951 ( .A(u5_mult_82_SUMB_40__5_), .ZN(u5_mult_82_n1028)
         );
  CLKBUF_X2 u5_mult_82_U950 ( .A(u5_mult_82_SUMB_38__6_), .Z(u5_mult_82_n383)
         );
  INV_X4 u5_mult_82_U949 ( .A(u5_mult_82_n381), .ZN(u5_mult_82_n382) );
  INV_X2 u5_mult_82_U948 ( .A(u5_mult_82_SUMB_9__27_), .ZN(u5_mult_82_n381) );
  INV_X8 u5_mult_82_U947 ( .A(u5_mult_82_n379), .ZN(u5_mult_82_n380) );
  INV_X4 u5_mult_82_U946 ( .A(u5_mult_82_SUMB_4__30_), .ZN(u5_mult_82_n379) );
  XOR2_X2 u5_mult_82_U945 ( .A(u5_mult_82_n5813), .B(u5_mult_82_n376), .Z(
        u5_mult_82_SUMB_48__1_) );
  XNOR2_X2 u5_mult_82_U944 ( .A(u5_mult_82_ab_35__9_), .B(
        u5_mult_82_CARRYB_34__9_), .ZN(u5_mult_82_n378) );
  XNOR2_X2 u5_mult_82_U943 ( .A(u5_mult_82_n378), .B(u5_mult_82_SUMB_34__10_), 
        .ZN(u5_mult_82_SUMB_35__9_) );
  XNOR2_X2 u5_mult_82_U942 ( .A(u5_mult_82_ab_30__11_), .B(
        u5_mult_82_CARRYB_29__11_), .ZN(u5_mult_82_n377) );
  XNOR2_X2 u5_mult_82_U941 ( .A(u5_mult_82_n377), .B(u5_mult_82_SUMB_29__12_), 
        .ZN(u5_mult_82_SUMB_30__11_) );
  NAND2_X1 u5_mult_82_U940 ( .A1(u5_mult_82_CARRYB_34__11_), .A2(
        u5_mult_82_SUMB_34__12_), .ZN(u5_mult_82_n1939) );
  NAND2_X1 u5_mult_82_U939 ( .A1(u5_mult_82_CARRYB_40__8_), .A2(
        u5_mult_82_SUMB_40__9_), .ZN(u5_mult_82_n2878) );
  CLKBUF_X2 u5_mult_82_U938 ( .A(u5_mult_82_CARRYB_47__1_), .Z(u5_mult_82_n376) );
  INV_X4 u5_mult_82_U937 ( .A(u5_mult_82_n2981), .ZN(u5_mult_82_n375) );
  NAND2_X2 u5_mult_82_U936 ( .A1(u5_mult_82_ab_8__24_), .A2(
        u5_mult_82_CARRYB_7__24_), .ZN(u5_mult_82_n3988) );
  NAND2_X1 u5_mult_82_U935 ( .A1(u5_mult_82_CARRYB_7__24_), .A2(
        u5_mult_82_SUMB_7__25_), .ZN(u5_mult_82_n3990) );
  NAND3_X4 u5_mult_82_U934 ( .A1(u5_mult_82_n3820), .A2(u5_mult_82_n3821), 
        .A3(u5_mult_82_n3822), .ZN(u5_mult_82_CARRYB_7__24_) );
  NAND2_X1 u5_mult_82_U933 ( .A1(u5_mult_82_CARRYB_45__5_), .A2(
        u5_mult_82_SUMB_45__6_), .ZN(u5_mult_82_n4661) );
  NAND2_X1 u5_mult_82_U932 ( .A1(u5_mult_82_ab_46__5_), .A2(
        u5_mult_82_SUMB_45__6_), .ZN(u5_mult_82_n4660) );
  XNOR2_X1 u5_mult_82_U931 ( .A(u5_mult_82_CARRYB_50__1_), .B(
        u5_mult_82_ab_51__1_), .ZN(u5_mult_82_n373) );
  XNOR2_X2 u5_mult_82_U930 ( .A(u5_mult_82_n373), .B(u5_mult_82_SUMB_50__2_), 
        .ZN(u5_mult_82_SUMB_51__1_) );
  XOR2_X2 u5_mult_82_U929 ( .A(u5_mult_82_ab_1__34_), .B(u5_mult_82_ab_0__35_), 
        .Z(u5_mult_82_n804) );
  CLKBUF_X3 u5_mult_82_U928 ( .A(u5_mult_82_SUMB_15__16_), .Z(u5_mult_82_n1454) );
  XNOR2_X1 u5_mult_82_U927 ( .A(u5_mult_82_SUMB_44__2_), .B(
        u5_mult_82_ab_45__1_), .ZN(u5_mult_82_n372) );
  XNOR2_X2 u5_mult_82_U926 ( .A(u5_mult_82_CARRYB_44__1_), .B(u5_mult_82_n372), 
        .ZN(u5_mult_82_SUMB_45__1_) );
  XOR2_X2 u5_mult_82_U925 ( .A(u5_mult_82_CARRYB_47__0_), .B(u5_mult_82_n2028), 
        .Z(u5_N48) );
  XNOR2_X2 u5_mult_82_U924 ( .A(u5_mult_82_SUMB_46__1_), .B(u5_mult_82_n626), 
        .ZN(u5_N47) );
  NAND2_X2 u5_mult_82_U923 ( .A1(u5_mult_82_CARRYB_24__29_), .A2(
        u5_mult_82_n54), .ZN(u5_mult_82_n5442) );
  NAND2_X1 u5_mult_82_U922 ( .A1(u5_mult_82_CARRYB_38__20_), .A2(
        u5_mult_82_SUMB_38__21_), .ZN(u5_mult_82_n4977) );
  XNOR2_X2 u5_mult_82_U921 ( .A(u5_mult_82_n4363), .B(u5_mult_82_SUMB_45__15_), 
        .ZN(u5_mult_82_n1537) );
  NAND2_X2 u5_mult_82_U920 ( .A1(u5_mult_82_CARRYB_7__36_), .A2(
        u5_mult_82_SUMB_7__37_), .ZN(u5_mult_82_n5623) );
  NAND2_X1 u5_mult_82_U919 ( .A1(u5_mult_82_ab_46__19_), .A2(
        u5_mult_82_CARRYB_45__19_), .ZN(u5_mult_82_n3848) );
  NAND2_X1 u5_mult_82_U918 ( .A1(u5_mult_82_CARRYB_45__19_), .A2(
        u5_mult_82_SUMB_45__20_), .ZN(u5_mult_82_n3850) );
  NAND3_X4 u5_mult_82_U917 ( .A1(u5_mult_82_n3957), .A2(u5_mult_82_n3958), 
        .A3(u5_mult_82_n3959), .ZN(u5_mult_82_CARRYB_33__25_) );
  NAND2_X1 u5_mult_82_U916 ( .A1(u5_mult_82_ab_35__19_), .A2(
        u5_mult_82_CARRYB_34__19_), .ZN(u5_mult_82_n6336) );
  CLKBUF_X1 u5_mult_82_U915 ( .A(u5_mult_82_CARRYB_22__26_), .Z(
        u5_mult_82_n402) );
  NAND2_X2 u5_mult_82_U914 ( .A1(u5_mult_82_ab_25__29_), .A2(u5_mult_82_n54), 
        .ZN(u5_mult_82_n5441) );
  NAND2_X1 u5_mult_82_U913 ( .A1(u5_mult_82_CARRYB_14__35_), .A2(
        u5_mult_82_SUMB_14__36_), .ZN(u5_mult_82_n5053) );
  NAND2_X1 u5_mult_82_U912 ( .A1(u5_mult_82_ab_41__19_), .A2(
        u5_mult_82_SUMB_40__20_), .ZN(u5_mult_82_n1133) );
  XNOR2_X2 u5_mult_82_U911 ( .A(u5_mult_82_ab_28__31_), .B(
        u5_mult_82_CARRYB_27__31_), .ZN(u5_mult_82_n1745) );
  XNOR2_X2 u5_mult_82_U910 ( .A(u5_mult_82_n411), .B(u5_mult_82_n1528), .ZN(
        u5_mult_82_SUMB_3__51_) );
  XNOR2_X2 u5_mult_82_U909 ( .A(u5_mult_82_n5248), .B(u5_mult_82_ab_19__44_), 
        .ZN(u5_mult_82_n1403) );
  XOR2_X2 u5_mult_82_U908 ( .A(u5_mult_82_ab_40__23_), .B(
        u5_mult_82_CARRYB_39__23_), .Z(u5_mult_82_n2239) );
  NAND3_X4 u5_mult_82_U907 ( .A1(u5_mult_82_n5709), .A2(u5_mult_82_n5710), 
        .A3(u5_mult_82_n5711), .ZN(u5_mult_82_CARRYB_47__19_) );
  NAND2_X2 u5_mult_82_U906 ( .A1(u5_mult_82_CARRYB_47__36_), .A2(
        u5_mult_82_SUMB_47__37_), .ZN(u5_mult_82_n3004) );
  XNOR2_X1 u5_mult_82_U905 ( .A(u5_mult_82_n2714), .B(u5_mult_82_SUMB_47__37_), 
        .ZN(u5_mult_82_SUMB_48__36_) );
  INV_X8 u5_mult_82_U904 ( .A(u5_mult_82_n1474), .ZN(u5_mult_82_n1475) );
  NAND2_X2 u5_mult_82_U903 ( .A1(u5_mult_82_ab_40__29_), .A2(
        u5_mult_82_CARRYB_39__29_), .ZN(u5_mult_82_n4331) );
  NAND3_X4 u5_mult_82_U902 ( .A1(u5_mult_82_n4329), .A2(u5_mult_82_n4330), 
        .A3(u5_mult_82_n4331), .ZN(u5_mult_82_CARRYB_40__29_) );
  NAND2_X1 u5_mult_82_U901 ( .A1(u5_mult_82_ab_45__13_), .A2(
        u5_mult_82_SUMB_44__14_), .ZN(u5_mult_82_n5462) );
  BUF_X2 u5_mult_82_U900 ( .A(u5_mult_82_CARRYB_45__19_), .Z(u5_mult_82_n730)
         );
  INV_X4 u5_mult_82_U899 ( .A(u5_mult_82_n5674), .ZN(u5_mult_82_n4157) );
  NAND2_X2 u5_mult_82_U898 ( .A1(u5_mult_82_ab_47__17_), .A2(
        u5_mult_82_SUMB_46__18_), .ZN(u5_mult_82_n5349) );
  NAND2_X2 u5_mult_82_U897 ( .A1(u5_mult_82_CARRYB_46__17_), .A2(
        u5_mult_82_SUMB_46__18_), .ZN(u5_mult_82_n5350) );
  NAND3_X4 u5_mult_82_U896 ( .A1(u5_mult_82_n5348), .A2(u5_mult_82_n5349), 
        .A3(u5_mult_82_n5350), .ZN(u5_mult_82_CARRYB_47__17_) );
  NAND2_X2 u5_mult_82_U895 ( .A1(u5_mult_82_CARRYB_45__34_), .A2(
        u5_mult_82_SUMB_45__35_), .ZN(u5_mult_82_n2658) );
  NAND2_X4 u5_mult_82_U894 ( .A1(u5_mult_82_ab_46__35_), .A2(u5_mult_82_n1570), 
        .ZN(u5_mult_82_n2918) );
  NAND3_X1 u5_mult_82_U893 ( .A1(u5_mult_82_n5642), .A2(u5_mult_82_n5643), 
        .A3(u5_mult_82_n5644), .ZN(u5_mult_82_n762) );
  BUF_X8 u5_mult_82_U892 ( .A(u5_mult_82_CARRYB_45__23_), .Z(u5_mult_82_n1595)
         );
  NAND2_X2 u5_mult_82_U891 ( .A1(u5_mult_82_ab_15__48_), .A2(
        u5_mult_82_SUMB_14__49_), .ZN(u5_mult_82_n4327) );
  NAND3_X4 u5_mult_82_U890 ( .A1(u5_mult_82_n2881), .A2(u5_mult_82_n2882), 
        .A3(u5_mult_82_n2883), .ZN(u5_mult_82_CARRYB_38__17_) );
  NAND2_X1 u5_mult_82_U889 ( .A1(u5_mult_82_CARRYB_15__37_), .A2(
        u5_mult_82_SUMB_15__38_), .ZN(u5_mult_82_n6305) );
  NAND3_X2 u5_mult_82_U888 ( .A1(u5_mult_82_n5039), .A2(u5_mult_82_n5038), 
        .A3(u5_mult_82_n5040), .ZN(u5_mult_82_CARRYB_18__36_) );
  BUF_X8 u5_mult_82_U887 ( .A(u5_mult_82_SUMB_29__30_), .Z(u5_mult_82_n410) );
  NAND2_X2 u5_mult_82_U886 ( .A1(u5_mult_82_ab_32__28_), .A2(
        u5_mult_82_SUMB_31__29_), .ZN(u5_mult_82_n5250) );
  NAND2_X2 u5_mult_82_U885 ( .A1(u5_mult_82_CARRYB_48__10_), .A2(
        u5_mult_82_SUMB_48__11_), .ZN(u5_mult_82_n6239) );
  NAND3_X4 u5_mult_82_U884 ( .A1(u5_mult_82_n6231), .A2(u5_mult_82_n6233), 
        .A3(u5_mult_82_n6232), .ZN(u5_mult_82_CARRYB_47__12_) );
  NAND2_X2 u5_mult_82_U883 ( .A1(u5_mult_82_ab_47__12_), .A2(u5_mult_82_n369), 
        .ZN(u5_mult_82_n6233) );
  INV_X32 u5_mult_82_U882 ( .A(u5_mult_82_ab_22__31_), .ZN(u5_mult_82_n371) );
  XNOR2_X2 u5_mult_82_U881 ( .A(u5_mult_82_CARRYB_21__31_), .B(u5_mult_82_n371), .ZN(u5_mult_82_n5265) );
  XNOR2_X2 u5_mult_82_U880 ( .A(u5_mult_82_ab_50__27_), .B(
        u5_mult_82_CARRYB_49__27_), .ZN(u5_mult_82_n370) );
  XNOR2_X2 u5_mult_82_U879 ( .A(u5_mult_82_n370), .B(u5_mult_82_SUMB_49__28_), 
        .ZN(u5_mult_82_SUMB_50__27_) );
  NAND2_X1 u5_mult_82_U878 ( .A1(u5_mult_82_ab_24__36_), .A2(
        u5_mult_82_CARRYB_23__36_), .ZN(u5_mult_82_n5737) );
  BUF_X8 u5_mult_82_U877 ( .A(u5_mult_82_CARRYB_50__19_), .Z(u5_mult_82_n2715)
         );
  NAND2_X1 u5_mult_82_U876 ( .A1(u5_mult_82_SUMB_52__14_), .A2(
        u5_mult_82_CARRYB_52__13_), .ZN(u5_mult_82_n6399) );
  NAND2_X2 u5_mult_82_U875 ( .A1(u5_mult_82_ab_46__12_), .A2(
        u5_mult_82_CARRYB_45__12_), .ZN(u5_mult_82_n5464) );
  INV_X1 u5_mult_82_U874 ( .A(u5_mult_82_ab_45__13_), .ZN(u5_mult_82_n3588) );
  NAND3_X1 u5_mult_82_U873 ( .A1(u5_mult_82_n5466), .A2(u5_mult_82_n5465), 
        .A3(u5_mult_82_n5464), .ZN(u5_mult_82_n369) );
  INV_X4 u5_mult_82_U872 ( .A(u5_mult_82_n3588), .ZN(u5_mult_82_n366) );
  INV_X2 u5_mult_82_U871 ( .A(u5_mult_82_CARRYB_44__13_), .ZN(u5_mult_82_n365)
         );
  NAND2_X2 u5_mult_82_U870 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n368), .ZN(
        u5_mult_82_n5460) );
  NAND2_X2 u5_mult_82_U869 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n366), .ZN(
        u5_mult_82_n368) );
  NAND2_X1 u5_mult_82_U868 ( .A1(u5_mult_82_CARRYB_44__13_), .A2(
        u5_mult_82_n3588), .ZN(u5_mult_82_n367) );
  NAND2_X2 u5_mult_82_U867 ( .A1(u5_mult_82_CARRYB_40__22_), .A2(
        u5_mult_82_ab_41__22_), .ZN(u5_mult_82_n2248) );
  NAND3_X4 u5_mult_82_U866 ( .A1(u5_mult_82_n362), .A2(u5_mult_82_n363), .A3(
        u5_mult_82_n364), .ZN(u5_mult_82_CARRYB_42__20_) );
  NAND2_X2 u5_mult_82_U865 ( .A1(u5_mult_82_CARRYB_41__20_), .A2(
        u5_mult_82_SUMB_41__21_), .ZN(u5_mult_82_n364) );
  NAND2_X2 u5_mult_82_U864 ( .A1(u5_mult_82_ab_42__20_), .A2(
        u5_mult_82_SUMB_41__21_), .ZN(u5_mult_82_n363) );
  NAND2_X1 u5_mult_82_U863 ( .A1(u5_mult_82_ab_42__20_), .A2(
        u5_mult_82_CARRYB_41__20_), .ZN(u5_mult_82_n362) );
  NAND3_X4 u5_mult_82_U862 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n360), .A3(
        u5_mult_82_n361), .ZN(u5_mult_82_CARRYB_41__21_) );
  NAND2_X2 u5_mult_82_U861 ( .A1(u5_mult_82_ab_41__21_), .A2(
        u5_mult_82_SUMB_40__22_), .ZN(u5_mult_82_n361) );
  NAND2_X2 u5_mult_82_U860 ( .A1(u5_mult_82_CARRYB_40__21_), .A2(
        u5_mult_82_SUMB_40__22_), .ZN(u5_mult_82_n360) );
  NAND2_X1 u5_mult_82_U859 ( .A1(u5_mult_82_CARRYB_40__21_), .A2(
        u5_mult_82_ab_41__21_), .ZN(u5_mult_82_n359) );
  XOR2_X2 u5_mult_82_U858 ( .A(u5_mult_82_n358), .B(u5_mult_82_SUMB_41__21_), 
        .Z(u5_mult_82_SUMB_42__20_) );
  XOR2_X2 u5_mult_82_U857 ( .A(u5_mult_82_ab_42__20_), .B(
        u5_mult_82_CARRYB_41__20_), .Z(u5_mult_82_n358) );
  XOR2_X2 u5_mult_82_U856 ( .A(u5_mult_82_n357), .B(u5_mult_82_SUMB_40__22_), 
        .Z(u5_mult_82_SUMB_41__21_) );
  XOR2_X2 u5_mult_82_U855 ( .A(u5_mult_82_CARRYB_40__21_), .B(
        u5_mult_82_ab_41__21_), .Z(u5_mult_82_n357) );
  NAND3_X4 u5_mult_82_U854 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n355), .A3(
        u5_mult_82_n356), .ZN(u5_mult_82_CARRYB_40__22_) );
  NAND2_X1 u5_mult_82_U853 ( .A1(u5_mult_82_ab_40__22_), .A2(
        u5_mult_82_CARRYB_39__22_), .ZN(u5_mult_82_n356) );
  NAND2_X2 u5_mult_82_U852 ( .A1(u5_mult_82_ab_40__22_), .A2(
        u5_mult_82_SUMB_39__23_), .ZN(u5_mult_82_n355) );
  NAND2_X2 u5_mult_82_U851 ( .A1(u5_mult_82_CARRYB_39__22_), .A2(
        u5_mult_82_SUMB_39__23_), .ZN(u5_mult_82_n354) );
  XOR2_X2 u5_mult_82_U850 ( .A(u5_mult_82_SUMB_39__23_), .B(u5_mult_82_n353), 
        .Z(u5_mult_82_SUMB_40__22_) );
  XOR2_X2 u5_mult_82_U849 ( .A(u5_mult_82_CARRYB_39__22_), .B(
        u5_mult_82_ab_40__22_), .Z(u5_mult_82_n353) );
  CLKBUF_X3 u5_mult_82_U848 ( .A(u5_mult_82_SUMB_26__27_), .Z(u5_mult_82_n1769) );
  CLKBUF_X3 u5_mult_82_U847 ( .A(u5_mult_82_CARRYB_28__26_), .Z(
        u5_mult_82_n1515) );
  NAND2_X2 u5_mult_82_U846 ( .A1(u5_mult_82_ab_30__26_), .A2(
        u5_mult_82_CARRYB_29__26_), .ZN(u5_mult_82_n6271) );
  NAND3_X4 u5_mult_82_U845 ( .A1(u5_mult_82_n3117), .A2(u5_mult_82_n3118), 
        .A3(u5_mult_82_n3119), .ZN(u5_mult_82_CARRYB_28__35_) );
  NAND2_X2 u5_mult_82_U844 ( .A1(u5_mult_82_ab_12__33_), .A2(
        u5_mult_82_CARRYB_11__33_), .ZN(u5_mult_82_n5702) );
  NAND2_X1 u5_mult_82_U843 ( .A1(u5_mult_82_CARRYB_11__33_), .A2(
        u5_mult_82_SUMB_11__34_), .ZN(u5_mult_82_n5704) );
  NAND2_X1 u5_mult_82_U842 ( .A1(u5_mult_82_ab_46__14_), .A2(
        u5_mult_82_SUMB_45__15_), .ZN(u5_mult_82_n5777) );
  NAND2_X1 u5_mult_82_U841 ( .A1(u5_mult_82_ab_47__14_), .A2(
        u5_mult_82_CARRYB_46__14_), .ZN(u5_mult_82_n5770) );
  BUF_X4 u5_mult_82_U840 ( .A(u5_mult_82_SUMB_49__27_), .Z(u5_mult_82_n694) );
  NAND3_X4 u5_mult_82_U839 ( .A1(u5_mult_82_n3935), .A2(u5_mult_82_n3936), 
        .A3(u5_mult_82_n3937), .ZN(u5_mult_82_CARRYB_39__34_) );
  NAND2_X2 u5_mult_82_U838 ( .A1(u5_mult_82_CARRYB_26__38_), .A2(
        u5_mult_82_SUMB_26__39_), .ZN(u5_mult_82_n1060) );
  NAND2_X2 u5_mult_82_U837 ( .A1(u5_mult_82_CARRYB_34__21_), .A2(
        u5_mult_82_SUMB_34__22_), .ZN(u5_mult_82_n4247) );
  XNOR2_X2 u5_mult_82_U836 ( .A(u5_mult_82_ab_33__40_), .B(
        u5_mult_82_CARRYB_32__40_), .ZN(u5_mult_82_n352) );
  XNOR2_X2 u5_mult_82_U835 ( .A(u5_mult_82_n352), .B(u5_mult_82_SUMB_32__41_), 
        .ZN(u5_mult_82_SUMB_33__40_) );
  XOR2_X2 u5_mult_82_U834 ( .A(u5_mult_82_n4418), .B(u5_mult_82_SUMB_40__31_), 
        .Z(u5_mult_82_SUMB_41__30_) );
  NAND2_X2 u5_mult_82_U833 ( .A1(u5_mult_82_ab_45__28_), .A2(
        u5_mult_82_CARRYB_44__28_), .ZN(u5_mult_82_n4570) );
  XNOR2_X2 u5_mult_82_U832 ( .A(u5_mult_82_ab_19__38_), .B(
        u5_mult_82_CARRYB_18__38_), .ZN(u5_mult_82_n351) );
  XNOR2_X2 u5_mult_82_U831 ( .A(u5_mult_82_n351), .B(u5_mult_82_SUMB_18__39_), 
        .ZN(u5_mult_82_SUMB_19__38_) );
  NAND2_X2 u5_mult_82_U830 ( .A1(u5_mult_82_ab_22__38_), .A2(
        u5_mult_82_SUMB_21__39_), .ZN(u5_mult_82_n2255) );
  BUF_X8 u5_mult_82_U829 ( .A(u5_mult_82_CARRYB_32__23_), .Z(u5_mult_82_n1727)
         );
  CLKBUF_X3 u5_mult_82_U828 ( .A(u5_mult_82_SUMB_35__23_), .Z(u5_mult_82_n1387) );
  NAND2_X2 u5_mult_82_U827 ( .A1(u5_mult_82_ab_36__18_), .A2(
        u5_mult_82_CARRYB_35__18_), .ZN(u5_mult_82_n5962) );
  NAND2_X2 u5_mult_82_U826 ( .A1(u5_mult_82_ab_44__14_), .A2(
        u5_mult_82_SUMB_43__15_), .ZN(u5_mult_82_n5458) );
  NAND2_X4 u5_mult_82_U825 ( .A1(u5_mult_82_n455), .A2(u5_mult_82_ab_43__17_), 
        .ZN(u5_mult_82_n4283) );
  NAND2_X2 u5_mult_82_U824 ( .A1(u5_mult_82_ab_30__31_), .A2(
        u5_mult_82_SUMB_29__32_), .ZN(u5_mult_82_n5163) );
  NAND2_X2 u5_mult_82_U823 ( .A1(u5_mult_82_CARRYB_8__51_), .A2(
        u5_mult_82_ab_8__52_), .ZN(u5_mult_82_n2086) );
  NAND2_X2 u5_mult_82_U822 ( .A1(u5_mult_82_CARRYB_8__51_), .A2(
        u5_mult_82_ab_9__51_), .ZN(u5_mult_82_n2084) );
  NAND2_X2 u5_mult_82_U821 ( .A1(u5_mult_82_ab_12__50_), .A2(
        u5_mult_82_SUMB_11__51_), .ZN(u5_mult_82_n3602) );
  XOR2_X1 u5_mult_82_U820 ( .A(u5_mult_82_CARRYB_16__50_), .B(u5_mult_82_n2581), .Z(u5_mult_82_SUMB_17__50_) );
  INV_X1 u5_mult_82_U819 ( .A(u5_mult_82_ab_18__37_), .ZN(u5_mult_82_n2006) );
  INV_X2 u5_mult_82_U818 ( .A(u5_mult_82_ab_29__31_), .ZN(u5_mult_82_n2051) );
  NAND3_X2 u5_mult_82_U817 ( .A1(u5_mult_82_n5035), .A2(u5_mult_82_n5036), 
        .A3(u5_mult_82_n5037), .ZN(u5_mult_82_n350) );
  NAND3_X2 u5_mult_82_U816 ( .A1(u5_mult_82_n2813), .A2(u5_mult_82_n2814), 
        .A3(u5_mult_82_n2815), .ZN(u5_mult_82_n349) );
  NAND3_X4 u5_mult_82_U815 ( .A1(u5_mult_82_n346), .A2(u5_mult_82_n347), .A3(
        u5_mult_82_n348), .ZN(u5_mult_82_CARRYB_27__31_) );
  NAND2_X2 u5_mult_82_U814 ( .A1(u5_mult_82_ab_27__31_), .A2(
        u5_mult_82_SUMB_26__32_), .ZN(u5_mult_82_n348) );
  NAND2_X2 u5_mult_82_U813 ( .A1(u5_mult_82_CARRYB_26__31_), .A2(
        u5_mult_82_SUMB_26__32_), .ZN(u5_mult_82_n347) );
  NAND2_X1 u5_mult_82_U812 ( .A1(u5_mult_82_CARRYB_26__31_), .A2(
        u5_mult_82_ab_27__31_), .ZN(u5_mult_82_n346) );
  NAND3_X4 u5_mult_82_U811 ( .A1(u5_mult_82_n343), .A2(u5_mult_82_n344), .A3(
        u5_mult_82_n345), .ZN(u5_mult_82_CARRYB_26__32_) );
  NAND2_X2 u5_mult_82_U810 ( .A1(u5_mult_82_CARRYB_25__32_), .A2(
        u5_mult_82_SUMB_25__33_), .ZN(u5_mult_82_n345) );
  NAND2_X2 u5_mult_82_U809 ( .A1(u5_mult_82_ab_26__32_), .A2(
        u5_mult_82_SUMB_25__33_), .ZN(u5_mult_82_n344) );
  NAND2_X1 u5_mult_82_U808 ( .A1(u5_mult_82_ab_26__32_), .A2(
        u5_mult_82_CARRYB_25__32_), .ZN(u5_mult_82_n343) );
  XOR2_X2 u5_mult_82_U807 ( .A(u5_mult_82_n342), .B(u5_mult_82_SUMB_26__32_), 
        .Z(u5_mult_82_SUMB_27__31_) );
  XOR2_X1 u5_mult_82_U806 ( .A(u5_mult_82_CARRYB_26__31_), .B(
        u5_mult_82_ab_27__31_), .Z(u5_mult_82_n342) );
  XOR2_X2 u5_mult_82_U805 ( .A(u5_mult_82_n341), .B(u5_mult_82_SUMB_25__33_), 
        .Z(u5_mult_82_SUMB_26__32_) );
  XOR2_X2 u5_mult_82_U804 ( .A(u5_mult_82_ab_26__32_), .B(
        u5_mult_82_CARRYB_25__32_), .Z(u5_mult_82_n341) );
  INV_X4 u5_mult_82_U803 ( .A(u5_mult_82_n350), .ZN(u5_mult_82_n338) );
  INV_X4 u5_mult_82_U802 ( .A(u5_mult_82_n2006), .ZN(u5_mult_82_n337) );
  NAND2_X2 u5_mult_82_U801 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n340), .ZN(
        u5_mult_82_n3392) );
  NAND2_X2 u5_mult_82_U800 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n338), .ZN(
        u5_mult_82_n340) );
  NAND2_X1 u5_mult_82_U799 ( .A1(u5_mult_82_n2006), .A2(
        u5_mult_82_CARRYB_17__37_), .ZN(u5_mult_82_n339) );
  INV_X4 u5_mult_82_U798 ( .A(u5_mult_82_CARRYB_28__31_), .ZN(u5_mult_82_n334)
         );
  INV_X8 u5_mult_82_U797 ( .A(u5_mult_82_n2051), .ZN(u5_mult_82_n333) );
  NAND2_X4 u5_mult_82_U796 ( .A1(u5_mult_82_n335), .A2(u5_mult_82_n336), .ZN(
        u5_mult_82_n6117) );
  NAND2_X4 u5_mult_82_U795 ( .A1(u5_mult_82_n333), .A2(u5_mult_82_n334), .ZN(
        u5_mult_82_n336) );
  NAND2_X2 u5_mult_82_U794 ( .A1(u5_mult_82_n2051), .A2(u5_mult_82_n349), .ZN(
        u5_mult_82_n335) );
  INV_X4 u5_mult_82_U793 ( .A(u5_mult_82_SUMB_41__20_), .ZN(u5_mult_82_n1750)
         );
  AND2_X2 u5_mult_82_U792 ( .A1(u5_mult_82_SUMB_52__21_), .A2(
        u5_mult_82_CARRYB_52__20_), .ZN(u5_mult_82_n584) );
  INV_X32 u5_mult_82_U791 ( .A(u5_mult_82_ab_52__21_), .ZN(u5_mult_82_n332) );
  XNOR2_X2 u5_mult_82_U790 ( .A(u5_mult_82_n332), .B(u5_mult_82_CARRYB_51__21_), .ZN(u5_mult_82_n4308) );
  NAND2_X2 u5_mult_82_U789 ( .A1(u5_mult_82_ab_46__10_), .A2(
        u5_mult_82_SUMB_45__11_), .ZN(u5_mult_82_n6263) );
  NAND3_X4 u5_mult_82_U788 ( .A1(u5_mult_82_n6262), .A2(u5_mult_82_n6263), 
        .A3(u5_mult_82_n6264), .ZN(u5_mult_82_CARRYB_46__10_) );
  NAND3_X4 u5_mult_82_U787 ( .A1(u5_mult_82_net82676), .A2(u5_mult_82_n3883), 
        .A3(u5_mult_82_net82678), .ZN(u5_mult_82_CARRYB_39__14_) );
  INV_X32 u5_mult_82_U786 ( .A(u5_mult_82_ab_17__41_), .ZN(u5_mult_82_n331) );
  XNOR2_X2 u5_mult_82_U785 ( .A(u5_mult_82_CARRYB_16__41_), .B(u5_mult_82_n331), .ZN(u5_mult_82_n940) );
  NAND2_X2 u5_mult_82_U784 ( .A1(u5_mult_82_ab_23__28_), .A2(
        u5_mult_82_CARRYB_22__28_), .ZN(u5_mult_82_n4297) );
  XNOR2_X1 u5_mult_82_U783 ( .A(u5_mult_82_n1747), .B(
        u5_mult_82_CARRYB_22__28_), .ZN(u5_mult_82_n4293) );
  NAND2_X2 u5_mult_82_U782 ( .A1(u5_mult_82_ab_33__23_), .A2(
        u5_mult_82_SUMB_32__24_), .ZN(u5_mult_82_n4009) );
  XNOR2_X1 u5_mult_82_U781 ( .A(u5_mult_82_ab_29__34_), .B(
        u5_mult_82_CARRYB_28__34_), .ZN(u5_mult_82_n330) );
  XNOR2_X2 u5_mult_82_U780 ( .A(u5_mult_82_n330), .B(u5_mult_82_SUMB_28__35_), 
        .ZN(u5_mult_82_SUMB_29__34_) );
  NAND2_X2 u5_mult_82_U779 ( .A1(u5_mult_82_ab_44__21_), .A2(
        u5_mult_82_SUMB_43__22_), .ZN(u5_mult_82_n5180) );
  CLKBUF_X3 u5_mult_82_U778 ( .A(u5_mult_82_SUMB_18__34_), .Z(u5_mult_82_n1626) );
  BUF_X8 u5_mult_82_U777 ( .A(u5_mult_82_CARRYB_32__25_), .Z(u5_mult_82_n1432)
         );
  INV_X32 u5_mult_82_U776 ( .A(u5_mult_82_ab_31__22_), .ZN(u5_mult_82_n329) );
  XNOR2_X2 u5_mult_82_U775 ( .A(u5_mult_82_n329), .B(u5_mult_82_CARRYB_30__22_), .ZN(u5_mult_82_n6298) );
  XNOR2_X2 u5_mult_82_U774 ( .A(u5_mult_82_ab_40__21_), .B(
        u5_mult_82_CARRYB_39__21_), .ZN(u5_mult_82_n328) );
  XNOR2_X2 u5_mult_82_U773 ( .A(u5_mult_82_n328), .B(u5_mult_82_SUMB_39__22_), 
        .ZN(u5_mult_82_SUMB_40__21_) );
  INV_X8 u5_mult_82_U772 ( .A(u5_mult_82_n6500), .ZN(u5_mult_82_CARRYB_1__45_)
         );
  NAND2_X4 u5_mult_82_U771 ( .A1(u5_mult_82_ab_0__46_), .A2(
        u5_mult_82_ab_1__45_), .ZN(u5_mult_82_n6500) );
  NAND2_X2 u5_mult_82_U770 ( .A1(u5_mult_82_ab_46__11_), .A2(
        u5_mult_82_SUMB_45__12_), .ZN(u5_mult_82_n5680) );
  BUF_X8 u5_mult_82_U769 ( .A(u5_mult_82_CARRYB_6__40_), .Z(u5_mult_82_n1726)
         );
  NAND3_X4 u5_mult_82_U768 ( .A1(u5_mult_82_n3527), .A2(u5_mult_82_n3528), 
        .A3(u5_mult_82_n3529), .ZN(u5_mult_82_CARRYB_2__42_) );
  NAND3_X2 u5_mult_82_U767 ( .A1(u5_mult_82_n325), .A2(u5_mult_82_n326), .A3(
        u5_mult_82_n327), .ZN(u5_mult_82_CARRYB_3__42_) );
  NAND2_X1 u5_mult_82_U766 ( .A1(u5_mult_82_ab_3__42_), .A2(
        u5_mult_82_CARRYB_2__42_), .ZN(u5_mult_82_n327) );
  NAND2_X2 u5_mult_82_U765 ( .A1(u5_mult_82_ab_3__42_), .A2(
        u5_mult_82_SUMB_2__43_), .ZN(u5_mult_82_n326) );
  NAND2_X1 u5_mult_82_U764 ( .A1(u5_mult_82_CARRYB_2__42_), .A2(
        u5_mult_82_SUMB_2__43_), .ZN(u5_mult_82_n325) );
  XOR2_X2 u5_mult_82_U763 ( .A(u5_mult_82_SUMB_2__43_), .B(u5_mult_82_n324), 
        .Z(u5_mult_82_SUMB_3__42_) );
  XOR2_X2 u5_mult_82_U762 ( .A(u5_mult_82_CARRYB_2__42_), .B(
        u5_mult_82_ab_3__42_), .Z(u5_mult_82_n324) );
  NAND2_X1 u5_mult_82_U761 ( .A1(u5_mult_82_SUMB_28__26_), .A2(
        u5_mult_82_CARRYB_28__25_), .ZN(u5_mult_82_n5450) );
  NAND2_X1 u5_mult_82_U760 ( .A1(u5_mult_82_ab_29__25_), .A2(
        u5_mult_82_SUMB_28__26_), .ZN(u5_mult_82_n5449) );
  XNOR2_X2 u5_mult_82_U759 ( .A(u5_mult_82_ab_45__28_), .B(
        u5_mult_82_CARRYB_44__28_), .ZN(u5_mult_82_n1741) );
  NAND2_X2 u5_mult_82_U758 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_ab_21__39_), 
        .ZN(u5_mult_82_n4944) );
  NAND3_X4 u5_mult_82_U757 ( .A1(u5_mult_82_n6302), .A2(u5_mult_82_n6303), 
        .A3(u5_mult_82_n6304), .ZN(u5_mult_82_CARRYB_31__22_) );
  NAND2_X2 u5_mult_82_U756 ( .A1(u5_mult_82_CARRYB_10__50_), .A2(
        u5_mult_82_SUMB_10__51_), .ZN(u5_mult_82_n3601) );
  NAND2_X2 u5_mult_82_U755 ( .A1(u5_mult_82_CARRYB_48__36_), .A2(
        u5_mult_82_SUMB_48__37_), .ZN(u5_mult_82_n2704) );
  INV_X4 u5_mult_82_U754 ( .A(u5_mult_82_CARRYB_35__22_), .ZN(u5_mult_82_n717)
         );
  NAND2_X1 u5_mult_82_U753 ( .A1(u5_mult_82_CARRYB_7__45_), .A2(
        u5_mult_82_n3278), .ZN(u5_mult_82_n2524) );
  NAND2_X1 u5_mult_82_U752 ( .A1(u5_mult_82_CARRYB_11__43_), .A2(
        u5_mult_82_SUMB_11__44_), .ZN(u5_mult_82_n5780) );
  NAND3_X4 u5_mult_82_U751 ( .A1(u5_mult_82_n5567), .A2(u5_mult_82_n5566), 
        .A3(u5_mult_82_n5568), .ZN(u5_mult_82_CARRYB_50__19_) );
  NAND3_X4 u5_mult_82_U750 ( .A1(u5_mult_82_n4208), .A2(u5_mult_82_n4209), 
        .A3(u5_mult_82_n4210), .ZN(u5_mult_82_CARRYB_46__13_) );
  NAND3_X4 u5_mult_82_U749 ( .A1(u5_mult_82_n2888), .A2(u5_mult_82_n2889), 
        .A3(u5_mult_82_n2890), .ZN(u5_mult_82_CARRYB_40__16_) );
  NAND3_X4 u5_mult_82_U748 ( .A1(u5_mult_82_n321), .A2(u5_mult_82_n322), .A3(
        u5_mult_82_n323), .ZN(u5_mult_82_CARRYB_17__45_) );
  NAND2_X1 u5_mult_82_U747 ( .A1(u5_mult_82_ab_17__45_), .A2(
        u5_mult_82_CARRYB_16__45_), .ZN(u5_mult_82_n323) );
  NAND2_X2 u5_mult_82_U746 ( .A1(u5_mult_82_ab_17__45_), .A2(
        u5_mult_82_SUMB_16__46_), .ZN(u5_mult_82_n322) );
  NAND2_X2 u5_mult_82_U745 ( .A1(u5_mult_82_CARRYB_16__45_), .A2(
        u5_mult_82_SUMB_16__46_), .ZN(u5_mult_82_n321) );
  XOR2_X2 u5_mult_82_U744 ( .A(u5_mult_82_SUMB_16__46_), .B(u5_mult_82_n320), 
        .Z(u5_mult_82_SUMB_17__45_) );
  XOR2_X2 u5_mult_82_U743 ( .A(u5_mult_82_CARRYB_16__45_), .B(
        u5_mult_82_ab_17__45_), .Z(u5_mult_82_n320) );
  XNOR2_X2 u5_mult_82_U742 ( .A(u5_mult_82_ab_31__23_), .B(
        u5_mult_82_CARRYB_30__23_), .ZN(u5_mult_82_n319) );
  XNOR2_X2 u5_mult_82_U741 ( .A(u5_mult_82_n319), .B(u5_mult_82_SUMB_30__24_), 
        .ZN(u5_mult_82_SUMB_31__23_) );
  NAND2_X2 u5_mult_82_U740 ( .A1(u5_mult_82_CARRYB_22__24_), .A2(
        u5_mult_82_SUMB_22__25_), .ZN(u5_mult_82_n2196) );
  BUF_X8 u5_mult_82_U739 ( .A(u5_mult_82_SUMB_22__23_), .Z(u5_mult_82_n1101)
         );
  INV_X2 u5_mult_82_U738 ( .A(u5_mult_82_CARRYB_36__15_), .ZN(u5_mult_82_n1355) );
  NAND2_X1 u5_mult_82_U737 ( .A1(u5_mult_82_ab_45__11_), .A2(
        u5_mult_82_CARRYB_44__11_), .ZN(u5_mult_82_n5407) );
  NAND2_X1 u5_mult_82_U736 ( .A1(u5_mult_82_CARRYB_46__11_), .A2(
        u5_mult_82_SUMB_46__12_), .ZN(u5_mult_82_n6208) );
  NAND2_X2 u5_mult_82_U735 ( .A1(u5_mult_82_ab_11__50_), .A2(
        u5_mult_82_CARRYB_10__50_), .ZN(u5_mult_82_n3599) );
  XNOR2_X1 u5_mult_82_U734 ( .A(u5_mult_82_CARRYB_10__50_), .B(
        u5_mult_82_ab_11__50_), .ZN(u5_mult_82_n2752) );
  NAND2_X2 u5_mult_82_U733 ( .A1(u5_mult_82_CARRYB_38__15_), .A2(
        u5_mult_82_SUMB_38__16_), .ZN(u5_mult_82_n5528) );
  NAND2_X2 u5_mult_82_U732 ( .A1(u5_mult_82_ab_39__15_), .A2(
        u5_mult_82_SUMB_38__16_), .ZN(u5_mult_82_n5527) );
  XNOR2_X1 u5_mult_82_U731 ( .A(u5_mult_82_CARRYB_22__24_), .B(
        u5_mult_82_ab_23__24_), .ZN(u5_mult_82_n318) );
  XNOR2_X2 u5_mult_82_U730 ( .A(u5_mult_82_n318), .B(u5_mult_82_SUMB_22__25_), 
        .ZN(u5_mult_82_SUMB_23__24_) );
  NAND2_X2 u5_mult_82_U729 ( .A1(u5_mult_82_ab_51__18_), .A2(
        u5_mult_82_SUMB_50__19_), .ZN(u5_mult_82_n5570) );
  INV_X4 u5_mult_82_U728 ( .A(u5_mult_82_n1840), .ZN(u5_mult_82_n1841) );
  XNOR2_X1 u5_mult_82_U727 ( .A(u5_mult_82_ab_50__19_), .B(
        u5_mult_82_CARRYB_49__19_), .ZN(u5_mult_82_n4147) );
  INV_X2 u5_mult_82_U726 ( .A(u5_mult_82_n1841), .ZN(u5_mult_82_n315) );
  INV_X1 u5_mult_82_U725 ( .A(u5_mult_82_n4147), .ZN(u5_mult_82_n314) );
  NAND2_X4 u5_mult_82_U724 ( .A1(u5_mult_82_n316), .A2(u5_mult_82_n317), .ZN(
        u5_mult_82_SUMB_50__19_) );
  NAND2_X4 u5_mult_82_U723 ( .A1(u5_mult_82_n314), .A2(u5_mult_82_n315), .ZN(
        u5_mult_82_n317) );
  NAND2_X1 u5_mult_82_U722 ( .A1(u5_mult_82_n4147), .A2(u5_mult_82_n1841), 
        .ZN(u5_mult_82_n316) );
  NAND3_X2 u5_mult_82_U721 ( .A1(u5_mult_82_n311), .A2(u5_mult_82_n312), .A3(
        u5_mult_82_n313), .ZN(u5_mult_82_CARRYB_20__39_) );
  NAND2_X1 u5_mult_82_U720 ( .A1(u5_mult_82_CARRYB_19__39_), .A2(
        u5_mult_82_SUMB_19__40_), .ZN(u5_mult_82_n313) );
  NAND2_X1 u5_mult_82_U719 ( .A1(u5_mult_82_ab_20__39_), .A2(
        u5_mult_82_SUMB_19__40_), .ZN(u5_mult_82_n312) );
  NAND2_X1 u5_mult_82_U718 ( .A1(u5_mult_82_ab_20__39_), .A2(
        u5_mult_82_CARRYB_19__39_), .ZN(u5_mult_82_n311) );
  NAND3_X2 u5_mult_82_U717 ( .A1(u5_mult_82_n308), .A2(u5_mult_82_n309), .A3(
        u5_mult_82_n310), .ZN(u5_mult_82_CARRYB_19__40_) );
  NAND2_X2 u5_mult_82_U716 ( .A1(u5_mult_82_CARRYB_18__40_), .A2(
        u5_mult_82_SUMB_18__41_), .ZN(u5_mult_82_n310) );
  NAND2_X2 u5_mult_82_U715 ( .A1(u5_mult_82_ab_19__40_), .A2(
        u5_mult_82_SUMB_18__41_), .ZN(u5_mult_82_n309) );
  NAND2_X1 u5_mult_82_U714 ( .A1(u5_mult_82_ab_19__40_), .A2(
        u5_mult_82_CARRYB_18__40_), .ZN(u5_mult_82_n308) );
  XOR2_X2 u5_mult_82_U713 ( .A(u5_mult_82_n307), .B(u5_mult_82_SUMB_19__40_), 
        .Z(u5_mult_82_SUMB_20__39_) );
  XOR2_X2 u5_mult_82_U712 ( .A(u5_mult_82_ab_20__39_), .B(
        u5_mult_82_CARRYB_19__39_), .Z(u5_mult_82_n307) );
  XOR2_X2 u5_mult_82_U711 ( .A(u5_mult_82_n306), .B(u5_mult_82_SUMB_18__41_), 
        .Z(u5_mult_82_SUMB_19__40_) );
  XOR2_X2 u5_mult_82_U710 ( .A(u5_mult_82_ab_19__40_), .B(
        u5_mult_82_CARRYB_18__40_), .Z(u5_mult_82_n306) );
  NAND3_X4 u5_mult_82_U709 ( .A1(u5_mult_82_n4626), .A2(u5_mult_82_n4627), 
        .A3(u5_mult_82_n4628), .ZN(u5_mult_82_CARRYB_16__26_) );
  NAND2_X2 u5_mult_82_U708 ( .A1(u5_mult_82_ab_33__19_), .A2(
        u5_mult_82_SUMB_32__20_), .ZN(u5_mult_82_n5416) );
  NAND2_X2 u5_mult_82_U707 ( .A1(u5_mult_82_n5641), .A2(
        u5_mult_82_SUMB_42__23_), .ZN(u5_mult_82_n5655) );
  INV_X32 u5_mult_82_U706 ( .A(u5_mult_82_ab_31__25_), .ZN(u5_mult_82_n305) );
  XNOR2_X2 u5_mult_82_U705 ( .A(u5_mult_82_n305), .B(u5_mult_82_CARRYB_30__25_), .ZN(u5_mult_82_n4235) );
  NAND2_X1 u5_mult_82_U704 ( .A1(u5_mult_82_CARRYB_50__8_), .A2(
        u5_mult_82_SUMB_50__9_), .ZN(u5_mult_82_n4171) );
  NAND2_X2 u5_mult_82_U703 ( .A1(u5_mult_82_SUMB_43__22_), .A2(
        u5_mult_82_CARRYB_43__21_), .ZN(u5_mult_82_n5182) );
  CLKBUF_X3 u5_mult_82_U702 ( .A(u5_mult_82_SUMB_36__18_), .Z(u5_mult_82_n304)
         );
  NAND2_X2 u5_mult_82_U701 ( .A1(u5_mult_82_net64225), .A2(n4791), .ZN(
        u5_mult_82_n1256) );
  NAND2_X2 u5_mult_82_U700 ( .A1(u5_mult_82_CARRYB_10__29_), .A2(
        u5_mult_82_SUMB_10__30_), .ZN(u5_mult_82_n2307) );
  INV_X4 u5_mult_82_U699 ( .A(u5_mult_82_n302), .ZN(u5_mult_82_n303) );
  INV_X2 u5_mult_82_U698 ( .A(u5_mult_82_CARRYB_17__29_), .ZN(u5_mult_82_n302)
         );
  NAND2_X1 u5_mult_82_U697 ( .A1(u5_mult_82_ab_14__34_), .A2(
        u5_mult_82_SUMB_13__35_), .ZN(u5_mult_82_n4856) );
  XNOR2_X2 u5_mult_82_U696 ( .A(u5_mult_82_n4907), .B(u5_mult_82_SUMB_22__31_), 
        .ZN(u5_mult_82_SUMB_23__30_) );
  NAND2_X2 u5_mult_82_U695 ( .A1(u5_mult_82_SUMB_19__33_), .A2(
        u5_mult_82_CARRYB_19__32_), .ZN(u5_mult_82_n3538) );
  NAND2_X4 u5_mult_82_U694 ( .A1(u5_mult_82_n3536), .A2(u5_mult_82_n1127), 
        .ZN(u5_mult_82_n3151) );
  NAND2_X4 u5_mult_82_U693 ( .A1(u5_mult_82_ab_25__28_), .A2(
        u5_mult_82_CARRYB_24__28_), .ZN(u5_mult_82_n1139) );
  NOR2_X1 u5_mult_82_U692 ( .A1(u5_mult_82_n6869), .A2(u5_mult_82_n6642), .ZN(
        u5_mult_82_ab_24__28_) );
  NAND3_X4 u5_mult_82_U691 ( .A1(u5_mult_82_n299), .A2(u5_mult_82_n300), .A3(
        u5_mult_82_n301), .ZN(u5_mult_82_CARRYB_24__28_) );
  NAND2_X1 u5_mult_82_U690 ( .A1(u5_mult_82_ab_24__28_), .A2(
        u5_mult_82_CARRYB_23__28_), .ZN(u5_mult_82_n301) );
  NAND2_X2 u5_mult_82_U689 ( .A1(u5_mult_82_ab_24__28_), .A2(
        u5_mult_82_SUMB_23__29_), .ZN(u5_mult_82_n300) );
  NAND2_X2 u5_mult_82_U688 ( .A1(u5_mult_82_CARRYB_23__28_), .A2(
        u5_mult_82_SUMB_23__29_), .ZN(u5_mult_82_n299) );
  XOR2_X2 u5_mult_82_U687 ( .A(u5_mult_82_SUMB_23__29_), .B(u5_mult_82_n298), 
        .Z(u5_mult_82_SUMB_24__28_) );
  XOR2_X2 u5_mult_82_U686 ( .A(u5_mult_82_CARRYB_23__28_), .B(
        u5_mult_82_ab_24__28_), .Z(u5_mult_82_n298) );
  XNOR2_X2 u5_mult_82_U685 ( .A(u5_mult_82_ab_48__24_), .B(
        u5_mult_82_CARRYB_47__24_), .ZN(u5_mult_82_n1409) );
  NAND2_X2 u5_mult_82_U684 ( .A1(u5_mult_82_ab_48__24_), .A2(
        u5_mult_82_CARRYB_47__24_), .ZN(u5_mult_82_n4301) );
  NOR2_X2 u5_mult_82_U683 ( .A1(u5_mult_82_n6815), .A2(u5_mult_82_net66107), 
        .ZN(u5_mult_82_ab_1__42_) );
  INV_X32 u5_mult_82_U682 ( .A(u5_mult_82_ab_24__24_), .ZN(u5_mult_82_n297) );
  XNOR2_X2 u5_mult_82_U681 ( .A(u5_mult_82_CARRYB_23__24_), .B(u5_mult_82_n297), .ZN(u5_mult_82_n1215) );
  NAND2_X2 u5_mult_82_U680 ( .A1(u5_mult_82_CARRYB_5__45_), .A2(
        u5_mult_82_SUMB_5__46_), .ZN(u5_mult_82_n6151) );
  NAND2_X1 u5_mult_82_U679 ( .A1(u5_mult_82_SUMB_50__22_), .A2(
        u5_mult_82_CARRYB_50__21_), .ZN(u5_mult_82_n5103) );
  NAND2_X1 u5_mult_82_U678 ( .A1(u5_mult_82_ab_51__21_), .A2(
        u5_mult_82_CARRYB_50__21_), .ZN(u5_mult_82_n5101) );
  NAND2_X4 u5_mult_82_U677 ( .A1(u5_mult_82_n3142), .A2(u5_mult_82_n3141), 
        .ZN(u5_mult_82_n5050) );
  NAND3_X4 u5_mult_82_U676 ( .A1(u5_mult_82_n5846), .A2(u5_mult_82_n5847), 
        .A3(u5_mult_82_n5848), .ZN(u5_mult_82_CARRYB_24__38_) );
  NAND2_X2 u5_mult_82_U675 ( .A1(u5_mult_82_ab_8__47_), .A2(
        u5_mult_82_SUMB_7__48_), .ZN(u5_mult_82_n3129) );
  INV_X4 u5_mult_82_U674 ( .A(u5_mult_82_SUMB_49__20_), .ZN(u5_mult_82_n1840)
         );
  NAND2_X2 u5_mult_82_U673 ( .A1(u5_mult_82_SUMB_3__50_), .A2(
        u5_mult_82_ab_4__49_), .ZN(u5_mult_82_n6317) );
  NAND3_X4 u5_mult_82_U672 ( .A1(u5_mult_82_net82047), .A2(u5_mult_82_net82048), .A3(u5_mult_82_n4217), .ZN(u5_mult_82_CARRYB_28__19_) );
  NAND3_X4 u5_mult_82_U671 ( .A1(u5_mult_82_n4951), .A2(u5_mult_82_n4952), 
        .A3(u5_mult_82_n4953), .ZN(u5_mult_82_CARRYB_34__14_) );
  NAND2_X2 u5_mult_82_U670 ( .A1(u5_mult_82_n4079), .A2(
        u5_mult_82_SUMB_34__15_), .ZN(u5_mult_82_n3785) );
  INV_X8 u5_mult_82_U669 ( .A(u5_mult_82_n1609), .ZN(u5_mult_82_n1610) );
  NAND2_X1 u5_mult_82_U668 ( .A1(u5_mult_82_SUMB_6__41_), .A2(
        u5_mult_82_ab_7__40_), .ZN(u5_mult_82_n4021) );
  INV_X8 u5_mult_82_U667 ( .A(u5_mult_82_n6504), .ZN(u5_mult_82_CARRYB_1__47_)
         );
  INV_X8 u5_mult_82_U666 ( .A(u5_mult_82_n701), .ZN(u5_mult_82_n702) );
  NAND2_X2 u5_mult_82_U665 ( .A1(u5_mult_82_CARRYB_25__16_), .A2(
        u5_mult_82_SUMB_25__17_), .ZN(u5_mult_82_n2783) );
  NAND3_X4 u5_mult_82_U664 ( .A1(u5_mult_82_n2781), .A2(u5_mult_82_n2782), 
        .A3(u5_mult_82_n2783), .ZN(u5_mult_82_CARRYB_26__16_) );
  NAND2_X4 u5_mult_82_U663 ( .A1(u5_mult_82_SUMB_21__19_), .A2(
        u5_mult_82_CARRYB_21__18_), .ZN(u5_mult_82_n4740) );
  NAND2_X1 u5_mult_82_U662 ( .A1(u5_mult_82_ab_2__45_), .A2(
        u5_mult_82_CARRYB_1__45_), .ZN(u5_mult_82_n2689) );
  NAND2_X1 u5_mult_82_U661 ( .A1(u5_mult_82_ab_8__40_), .A2(
        u5_mult_82_CARRYB_7__40_), .ZN(u5_mult_82_n6021) );
  XNOR2_X1 u5_mult_82_U660 ( .A(u5_mult_82_CARRYB_2__43_), .B(
        u5_mult_82_ab_3__43_), .ZN(u5_mult_82_n1712) );
  NAND3_X4 u5_mult_82_U659 ( .A1(u5_mult_82_n294), .A2(u5_mult_82_n295), .A3(
        u5_mult_82_n296), .ZN(u5_mult_82_CARRYB_6__40_) );
  NAND2_X2 u5_mult_82_U658 ( .A1(u5_mult_82_CARRYB_5__40_), .A2(
        u5_mult_82_SUMB_5__41_), .ZN(u5_mult_82_n296) );
  NAND2_X2 u5_mult_82_U657 ( .A1(u5_mult_82_ab_6__40_), .A2(
        u5_mult_82_SUMB_5__41_), .ZN(u5_mult_82_n295) );
  NAND2_X1 u5_mult_82_U656 ( .A1(u5_mult_82_ab_6__40_), .A2(
        u5_mult_82_CARRYB_5__40_), .ZN(u5_mult_82_n294) );
  NAND3_X2 u5_mult_82_U655 ( .A1(u5_mult_82_n291), .A2(u5_mult_82_n292), .A3(
        u5_mult_82_n293), .ZN(u5_mult_82_CARRYB_5__41_) );
  NAND2_X1 u5_mult_82_U654 ( .A1(u5_mult_82_CARRYB_4__41_), .A2(
        u5_mult_82_SUMB_4__42_), .ZN(u5_mult_82_n293) );
  NAND2_X1 u5_mult_82_U653 ( .A1(u5_mult_82_ab_5__41_), .A2(
        u5_mult_82_SUMB_4__42_), .ZN(u5_mult_82_n292) );
  NAND2_X1 u5_mult_82_U652 ( .A1(u5_mult_82_ab_5__41_), .A2(
        u5_mult_82_CARRYB_4__41_), .ZN(u5_mult_82_n291) );
  XOR2_X2 u5_mult_82_U651 ( .A(u5_mult_82_n290), .B(u5_mult_82_SUMB_5__41_), 
        .Z(u5_mult_82_SUMB_6__40_) );
  XOR2_X2 u5_mult_82_U650 ( .A(u5_mult_82_ab_6__40_), .B(
        u5_mult_82_CARRYB_5__40_), .Z(u5_mult_82_n290) );
  XOR2_X2 u5_mult_82_U649 ( .A(u5_mult_82_n289), .B(u5_mult_82_SUMB_4__42_), 
        .Z(u5_mult_82_SUMB_5__41_) );
  XOR2_X2 u5_mult_82_U648 ( .A(u5_mult_82_ab_5__41_), .B(
        u5_mult_82_CARRYB_4__41_), .Z(u5_mult_82_n289) );
  XOR2_X2 u5_mult_82_U647 ( .A(u5_mult_82_ab_37__10_), .B(
        u5_mult_82_CARRYB_36__10_), .Z(u5_mult_82_n982) );
  NAND2_X2 u5_mult_82_U646 ( .A1(u5_mult_82_CARRYB_12__25_), .A2(
        u5_mult_82_SUMB_12__26_), .ZN(u5_mult_82_n2204) );
  NAND2_X2 u5_mult_82_U645 ( .A1(u5_mult_82_ab_42__7_), .A2(
        u5_mult_82_CARRYB_41__7_), .ZN(u5_mult_82_n6027) );
  NAND3_X4 u5_mult_82_U644 ( .A1(u5_mult_82_n652), .A2(u5_mult_82_n653), .A3(
        u5_mult_82_n654), .ZN(u5_mult_82_CARRYB_31__13_) );
  NAND3_X4 u5_mult_82_U643 ( .A1(u5_mult_82_n986), .A2(u5_mult_82_n987), .A3(
        u5_mult_82_n988), .ZN(u5_mult_82_CARRYB_37__10_) );
  NAND2_X2 u5_mult_82_U642 ( .A1(u5_mult_82_CARRYB_6__28_), .A2(
        u5_mult_82_SUMB_6__29_), .ZN(u5_mult_82_n2623) );
  INV_X4 u5_mult_82_U641 ( .A(u5_mult_82_n287), .ZN(u5_mult_82_n288) );
  INV_X4 u5_mult_82_U640 ( .A(u5_mult_82_SUMB_4__36_), .ZN(u5_mult_82_n287) );
  XOR2_X1 u5_mult_82_U639 ( .A(u5_mult_82_n2087), .B(u5_mult_82_CARRYB_9__51_), 
        .Z(u5_mult_82_SUMB_10__51_) );
  XOR2_X1 u5_mult_82_U638 ( .A(u5_mult_82_n2095), .B(u5_mult_82_CARRYB_13__51_), .Z(u5_mult_82_SUMB_14__51_) );
  NAND2_X1 u5_mult_82_U637 ( .A1(u5_mult_82_ab_18__49_), .A2(
        u5_mult_82_SUMB_17__50_), .ZN(u5_mult_82_n1198) );
  NAND2_X1 u5_mult_82_U636 ( .A1(u5_mult_82_SUMB_17__50_), .A2(
        u5_mult_82_CARRYB_17__49_), .ZN(u5_mult_82_n1196) );
  NAND2_X2 u5_mult_82_U635 ( .A1(u5_mult_82_CARRYB_16__48_), .A2(
        u5_mult_82_SUMB_16__49_), .ZN(u5_mult_82_n4428) );
  INV_X16 u5_mult_82_U634 ( .A(n4791), .ZN(u5_mult_82_net64961) );
  NAND2_X2 u5_mult_82_U633 ( .A1(u5_mult_82_SUMB_18__48_), .A2(
        u5_mult_82_CARRYB_18__47_), .ZN(u5_mult_82_n3105) );
  XNOR2_X2 u5_mult_82_U632 ( .A(u5_mult_82_ab_32__40_), .B(
        u5_mult_82_CARRYB_31__40_), .ZN(u5_mult_82_n2691) );
  NAND2_X2 u5_mult_82_U631 ( .A1(u5_mult_82_SUMB_15__47_), .A2(
        u5_mult_82_CARRYB_15__46_), .ZN(u5_mult_82_n4614) );
  NAND2_X2 u5_mult_82_U630 ( .A1(u5_mult_82_ab_25__36_), .A2(
        u5_mult_82_CARRYB_24__36_), .ZN(u5_mult_82_n5557) );
  XNOR2_X2 u5_mult_82_U629 ( .A(u5_mult_82_CARRYB_17__33_), .B(
        u5_mult_82_ab_18__33_), .ZN(u5_mult_82_n286) );
  XNOR2_X2 u5_mult_82_U628 ( .A(u5_mult_82_SUMB_17__34_), .B(u5_mult_82_n286), 
        .ZN(u5_mult_82_SUMB_18__33_) );
  NAND2_X2 u5_mult_82_U627 ( .A1(u5_mult_82_ab_17__37_), .A2(
        u5_mult_82_CARRYB_16__37_), .ZN(u5_mult_82_n5035) );
  NAND2_X4 u5_mult_82_U626 ( .A1(u5_mult_82_ab_43__22_), .A2(u5_mult_82_n5641), 
        .ZN(u5_mult_82_n5657) );
  XNOR2_X2 u5_mult_82_U625 ( .A(u5_mult_82_ab_15__46_), .B(
        u5_mult_82_CARRYB_14__46_), .ZN(u5_mult_82_n1913) );
  NAND2_X4 u5_mult_82_U624 ( .A1(u5_mult_82_n1559), .A2(u5_mult_82_ab_19__43_), 
        .ZN(u5_mult_82_n5841) );
  XNOR2_X2 u5_mult_82_U623 ( .A(u5_mult_82_ab_40__13_), .B(
        u5_mult_82_CARRYB_39__13_), .ZN(u5_mult_82_n1377) );
  NAND2_X2 u5_mult_82_U622 ( .A1(u5_mult_82_CARRYB_28__19_), .A2(
        u5_mult_82_SUMB_28__20_), .ZN(u5_mult_82_n494) );
  NAND3_X4 u5_mult_82_U621 ( .A1(u5_mult_82_n492), .A2(u5_mult_82_n493), .A3(
        u5_mult_82_n494), .ZN(u5_mult_82_CARRYB_29__19_) );
  NAND2_X4 u5_mult_82_U620 ( .A1(u5_mult_82_ab_16__34_), .A2(u5_mult_82_n3140), 
        .ZN(u5_mult_82_n3142) );
  NAND3_X4 u5_mult_82_U619 ( .A1(u5_mult_82_n5131), .A2(u5_mult_82_n5132), 
        .A3(u5_mult_82_n5133), .ZN(u5_mult_82_CARRYB_39__11_) );
  NAND2_X4 u5_mult_82_U618 ( .A1(u5_mult_82_n6835), .A2(u5_mult_82_net66121), 
        .ZN(u5_mult_82_n2311) );
  XNOR2_X2 u5_mult_82_U617 ( .A(u5_mult_82_SUMB_23__24_), .B(u5_mult_82_n643), 
        .ZN(u5_mult_82_SUMB_24__23_) );
  NAND2_X1 u5_mult_82_U616 ( .A1(u5_mult_82_SUMB_12__39_), .A2(
        u5_mult_82_CARRYB_12__38_), .ZN(u5_mult_82_n6161) );
  INV_X32 u5_mult_82_U615 ( .A(u5_mult_82_ab_32__22_), .ZN(u5_mult_82_n285) );
  XNOR2_X2 u5_mult_82_U614 ( .A(u5_mult_82_n285), .B(u5_mult_82_CARRYB_31__22_), .ZN(u5_mult_82_n3519) );
  XNOR2_X2 u5_mult_82_U613 ( .A(u5_mult_82_ab_11__38_), .B(
        u5_mult_82_CARRYB_10__38_), .ZN(u5_mult_82_n1603) );
  NAND3_X4 u5_mult_82_U612 ( .A1(u5_mult_82_n5794), .A2(u5_mult_82_n5795), 
        .A3(u5_mult_82_n5796), .ZN(u5_mult_82_CARRYB_15__31_) );
  XNOR2_X2 u5_mult_82_U611 ( .A(u5_mult_82_ab_22__38_), .B(
        u5_mult_82_CARRYB_21__38_), .ZN(u5_mult_82_n464) );
  NAND2_X2 u5_mult_82_U610 ( .A1(u5_mult_82_ab_22__38_), .A2(
        u5_mult_82_CARRYB_21__38_), .ZN(u5_mult_82_n2254) );
  NAND2_X1 u5_mult_82_U609 ( .A1(u5_mult_82_ab_16__33_), .A2(
        u5_mult_82_SUMB_15__34_), .ZN(u5_mult_82_n6046) );
  INV_X16 u5_mult_82_U608 ( .A(u5_mult_82_n6763), .ZN(u5_mult_82_n6761) );
  INV_X1 u5_mult_82_U607 ( .A(u5_mult_82_n6764), .ZN(u5_mult_82_n6760) );
  INV_X4 u5_mult_82_U606 ( .A(u5_mult_82_n6758), .ZN(u5_mult_82_n6763) );
  INV_X4 u5_mult_82_U605 ( .A(u5_mult_82_SUMB_20__35_), .ZN(u5_mult_82_n1724)
         );
  NAND2_X2 u5_mult_82_U604 ( .A1(u5_mult_82_ab_21__35_), .A2(
        u5_mult_82_CARRYB_20__35_), .ZN(u5_mult_82_n4986) );
  NAND3_X2 u5_mult_82_U603 ( .A1(u5_mult_82_n282), .A2(u5_mult_82_n283), .A3(
        u5_mult_82_n284), .ZN(u5_mult_82_CARRYB_20__35_) );
  NAND2_X1 u5_mult_82_U602 ( .A1(u5_mult_82_ab_20__35_), .A2(
        u5_mult_82_CARRYB_19__35_), .ZN(u5_mult_82_n284) );
  NAND2_X1 u5_mult_82_U601 ( .A1(u5_mult_82_ab_20__35_), .A2(
        u5_mult_82_SUMB_19__36_), .ZN(u5_mult_82_n283) );
  NAND2_X1 u5_mult_82_U600 ( .A1(u5_mult_82_CARRYB_19__35_), .A2(
        u5_mult_82_SUMB_19__36_), .ZN(u5_mult_82_n282) );
  XOR2_X2 u5_mult_82_U599 ( .A(u5_mult_82_SUMB_19__36_), .B(u5_mult_82_n281), 
        .Z(u5_mult_82_SUMB_20__35_) );
  XOR2_X2 u5_mult_82_U598 ( .A(u5_mult_82_CARRYB_19__35_), .B(
        u5_mult_82_ab_20__35_), .Z(u5_mult_82_n281) );
  NAND2_X2 u5_mult_82_U597 ( .A1(u5_mult_82_CARRYB_34__19_), .A2(
        u5_mult_82_SUMB_34__20_), .ZN(u5_mult_82_n6338) );
  NAND2_X2 u5_mult_82_U596 ( .A1(u5_mult_82_CARRYB_18__22_), .A2(
        u5_mult_82_SUMB_18__23_), .ZN(u5_mult_82_n3246) );
  NAND2_X2 u5_mult_82_U595 ( .A1(u5_mult_82_ab_13__25_), .A2(
        u5_mult_82_SUMB_12__26_), .ZN(u5_mult_82_n2203) );
  XNOR2_X2 u5_mult_82_U594 ( .A(u5_mult_82_CARRYB_36__20_), .B(
        u5_mult_82_ab_37__20_), .ZN(u5_mult_82_n280) );
  XNOR2_X2 u5_mult_82_U593 ( .A(u5_mult_82_SUMB_36__21_), .B(u5_mult_82_n280), 
        .ZN(u5_mult_82_SUMB_37__20_) );
  NAND2_X2 u5_mult_82_U592 ( .A1(u5_mult_82_ab_1__50_), .A2(
        u5_mult_82_ab_0__51_), .ZN(u5_mult_82_n6510) );
  NAND3_X2 u5_mult_82_U591 ( .A1(u5_mult_82_n277), .A2(u5_mult_82_n278), .A3(
        u5_mult_82_n279), .ZN(u5_mult_82_CARRYB_23__47_) );
  NAND2_X1 u5_mult_82_U590 ( .A1(u5_mult_82_CARRYB_22__47_), .A2(
        u5_mult_82_SUMB_22__48_), .ZN(u5_mult_82_n279) );
  NAND2_X1 u5_mult_82_U589 ( .A1(u5_mult_82_ab_23__47_), .A2(
        u5_mult_82_SUMB_22__48_), .ZN(u5_mult_82_n278) );
  NAND2_X1 u5_mult_82_U588 ( .A1(u5_mult_82_ab_23__47_), .A2(
        u5_mult_82_CARRYB_22__47_), .ZN(u5_mult_82_n277) );
  NAND3_X2 u5_mult_82_U587 ( .A1(u5_mult_82_n274), .A2(u5_mult_82_n275), .A3(
        u5_mult_82_n276), .ZN(u5_mult_82_CARRYB_22__48_) );
  NAND2_X2 u5_mult_82_U586 ( .A1(u5_mult_82_CARRYB_21__48_), .A2(
        u5_mult_82_SUMB_21__49_), .ZN(u5_mult_82_n276) );
  NAND2_X2 u5_mult_82_U585 ( .A1(u5_mult_82_ab_22__48_), .A2(
        u5_mult_82_SUMB_21__49_), .ZN(u5_mult_82_n275) );
  NAND2_X2 u5_mult_82_U584 ( .A1(u5_mult_82_ab_22__48_), .A2(
        u5_mult_82_CARRYB_21__48_), .ZN(u5_mult_82_n274) );
  XOR2_X2 u5_mult_82_U583 ( .A(u5_mult_82_n273), .B(u5_mult_82_SUMB_22__48_), 
        .Z(u5_mult_82_SUMB_23__47_) );
  XOR2_X1 u5_mult_82_U582 ( .A(u5_mult_82_ab_23__47_), .B(
        u5_mult_82_CARRYB_22__47_), .Z(u5_mult_82_n273) );
  XOR2_X2 u5_mult_82_U581 ( .A(u5_mult_82_n272), .B(u5_mult_82_SUMB_21__49_), 
        .Z(u5_mult_82_SUMB_22__48_) );
  XOR2_X2 u5_mult_82_U580 ( .A(u5_mult_82_ab_22__48_), .B(
        u5_mult_82_CARRYB_21__48_), .Z(u5_mult_82_n272) );
  INV_X4 u5_mult_82_U579 ( .A(u5_mult_82_SUMB_34__26_), .ZN(u5_mult_82_n1814)
         );
  AND2_X2 u5_mult_82_U578 ( .A1(u5_mult_82_SUMB_52__11_), .A2(
        u5_mult_82_CARRYB_52__10_), .ZN(u5_mult_82_n583) );
  INV_X32 u5_mult_82_U577 ( .A(u5_mult_82_net86084), .ZN(u5_mult_82_net64223)
         );
  NAND2_X1 u5_mult_82_U576 ( .A1(u5_mult_82_ab_49__12_), .A2(u5_mult_82_n1843), 
        .ZN(u5_mult_82_n5989) );
  INV_X32 u5_mult_82_U575 ( .A(u5_mult_82_ab_32__20_), .ZN(u5_mult_82_n271) );
  XNOR2_X2 u5_mult_82_U574 ( .A(u5_mult_82_n271), .B(u5_mult_82_CARRYB_31__20_), .ZN(u5_mult_82_n5410) );
  XNOR2_X2 u5_mult_82_U573 ( .A(u5_mult_82_ab_42__15_), .B(
        u5_mult_82_CARRYB_41__15_), .ZN(u5_mult_82_n1494) );
  NOR2_X4 u5_mult_82_U572 ( .A1(u5_mult_82_n6863), .A2(u5_mult_82_n6649), .ZN(
        u5_mult_82_ab_26__29_) );
  NAND2_X4 u5_mult_82_U571 ( .A1(u5_mult_82_ab_43__18_), .A2(
        u5_mult_82_CARRYB_42__18_), .ZN(u5_mult_82_n4232) );
  NOR2_X1 u5_mult_82_U570 ( .A1(u5_mult_82_n6919), .A2(u5_mult_82_net65371), 
        .ZN(u5_mult_82_ab_42__18_) );
  INV_X4 u5_mult_82_U569 ( .A(u5_mult_82_ab_26__29_), .ZN(u5_mult_82_n268) );
  INV_X4 u5_mult_82_U568 ( .A(u5_mult_82_CARRYB_25__29_), .ZN(u5_mult_82_n267)
         );
  NAND2_X2 u5_mult_82_U567 ( .A1(u5_mult_82_n269), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_n2749) );
  NAND2_X4 u5_mult_82_U566 ( .A1(u5_mult_82_n267), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_n270) );
  NAND2_X1 u5_mult_82_U565 ( .A1(u5_mult_82_CARRYB_25__29_), .A2(
        u5_mult_82_ab_26__29_), .ZN(u5_mult_82_n269) );
  NAND3_X4 u5_mult_82_U564 ( .A1(u5_mult_82_n264), .A2(u5_mult_82_n265), .A3(
        u5_mult_82_n266), .ZN(u5_mult_82_CARRYB_42__18_) );
  NAND2_X1 u5_mult_82_U563 ( .A1(u5_mult_82_ab_42__18_), .A2(
        u5_mult_82_CARRYB_41__18_), .ZN(u5_mult_82_n266) );
  NAND2_X2 u5_mult_82_U562 ( .A1(u5_mult_82_ab_42__18_), .A2(
        u5_mult_82_SUMB_41__19_), .ZN(u5_mult_82_n265) );
  NAND2_X1 u5_mult_82_U561 ( .A1(u5_mult_82_CARRYB_41__18_), .A2(
        u5_mult_82_SUMB_41__19_), .ZN(u5_mult_82_n264) );
  XNOR2_X2 u5_mult_82_U560 ( .A(u5_mult_82_ab_12__44_), .B(
        u5_mult_82_CARRYB_11__44_), .ZN(u5_mult_82_n263) );
  XNOR2_X2 u5_mult_82_U559 ( .A(u5_mult_82_n263), .B(u5_mult_82_SUMB_11__45_), 
        .ZN(u5_mult_82_SUMB_12__44_) );
  INV_X8 u5_mult_82_U558 ( .A(u5_mult_82_n6509), .ZN(u5_mult_82_SUMB_1__49_)
         );
  CLKBUF_X3 u5_mult_82_U557 ( .A(u5_mult_82_CARRYB_5__46_), .Z(u5_mult_82_n736) );
  XNOR2_X2 u5_mult_82_U556 ( .A(u5_mult_82_ab_1__36_), .B(u5_mult_82_n4414), 
        .ZN(u5_mult_82_n6491) );
  NAND2_X1 u5_mult_82_U555 ( .A1(u5_mult_82_ab_45__10_), .A2(
        u5_mult_82_CARRYB_44__10_), .ZN(u5_mult_82_n2567) );
  NAND3_X2 u5_mult_82_U554 ( .A1(u5_mult_82_n5699), .A2(u5_mult_82_n5700), 
        .A3(u5_mult_82_n5701), .ZN(u5_mult_82_CARRYB_10__35_) );
  NAND2_X2 u5_mult_82_U553 ( .A1(u5_mult_82_ab_50__11_), .A2(u5_mult_82_n1419), 
        .ZN(u5_mult_82_n5992) );
  XOR2_X2 u5_mult_82_U552 ( .A(u5_mult_82_CARRYB_27__42_), .B(
        u5_mult_82_ab_28__42_), .Z(u5_mult_82_n2176) );
  XNOR2_X2 u5_mult_82_U551 ( .A(u5_mult_82_ab_35__41_), .B(
        u5_mult_82_CARRYB_34__41_), .ZN(u5_mult_82_n262) );
  XNOR2_X2 u5_mult_82_U550 ( .A(u5_mult_82_n262), .B(u5_mult_82_SUMB_34__42_), 
        .ZN(u5_mult_82_SUMB_35__41_) );
  NAND2_X2 u5_mult_82_U549 ( .A1(u5_mult_82_n762), .A2(u5_mult_82_SUMB_11__45_), .ZN(u5_mult_82_n939) );
  NOR2_X2 u5_mult_82_U548 ( .A1(u5_mult_82_net64505), .A2(u5_mult_82_net65283), 
        .ZN(u5_mult_82_ab_47__13_) );
  INV_X1 u5_mult_82_U547 ( .A(u5_mult_82_SUMB_38__20_), .ZN(u5_mult_82_n259)
         );
  INV_X4 u5_mult_82_U546 ( .A(u5_mult_82_n767), .ZN(u5_mult_82_n258) );
  NAND2_X2 u5_mult_82_U545 ( .A1(u5_mult_82_n767), .A2(u5_mult_82_SUMB_38__20_), .ZN(u5_mult_82_n260) );
  NAND3_X2 u5_mult_82_U544 ( .A1(u5_mult_82_n255), .A2(u5_mult_82_n256), .A3(
        u5_mult_82_n257), .ZN(u5_mult_82_CARRYB_47__13_) );
  NAND2_X1 u5_mult_82_U543 ( .A1(u5_mult_82_ab_47__13_), .A2(
        u5_mult_82_CARRYB_46__13_), .ZN(u5_mult_82_n257) );
  NAND2_X2 u5_mult_82_U542 ( .A1(u5_mult_82_ab_47__13_), .A2(
        u5_mult_82_SUMB_46__14_), .ZN(u5_mult_82_n256) );
  NAND2_X2 u5_mult_82_U541 ( .A1(u5_mult_82_CARRYB_46__13_), .A2(
        u5_mult_82_SUMB_46__14_), .ZN(u5_mult_82_n255) );
  XOR2_X2 u5_mult_82_U540 ( .A(u5_mult_82_SUMB_46__14_), .B(u5_mult_82_n254), 
        .Z(u5_mult_82_SUMB_47__13_) );
  XOR2_X2 u5_mult_82_U539 ( .A(u5_mult_82_CARRYB_46__13_), .B(
        u5_mult_82_ab_47__13_), .Z(u5_mult_82_n254) );
  BUF_X8 u5_mult_82_U538 ( .A(u5_mult_82_CARRYB_16__20_), .Z(u5_mult_82_n1625)
         );
  NAND2_X4 u5_mult_82_U537 ( .A1(u5_mult_82_SUMB_25__15_), .A2(
        u5_mult_82_ab_26__14_), .ZN(u5_mult_82_n4066) );
  NAND3_X2 u5_mult_82_U536 ( .A1(u5_mult_82_n4763), .A2(u5_mult_82_n4764), 
        .A3(u5_mult_82_n4765), .ZN(u5_mult_82_CARRYB_32__13_) );
  XNOR2_X2 u5_mult_82_U535 ( .A(u5_mult_82_ab_16__41_), .B(
        u5_mult_82_CARRYB_15__41_), .ZN(u5_mult_82_n253) );
  XNOR2_X2 u5_mult_82_U534 ( .A(u5_mult_82_n253), .B(u5_mult_82_SUMB_15__42_), 
        .ZN(u5_mult_82_SUMB_16__41_) );
  NAND2_X2 u5_mult_82_U533 ( .A1(u5_mult_82_CARRYB_19__24_), .A2(
        u5_mult_82_SUMB_19__25_), .ZN(u5_mult_82_n5613) );
  INV_X2 u5_mult_82_U532 ( .A(u5_mult_82_SUMB_20__25_), .ZN(
        u5_mult_82_net87429) );
  INV_X4 u5_mult_82_U531 ( .A(u5_mult_82_n1315), .ZN(u5_mult_82_n250) );
  INV_X4 u5_mult_82_U530 ( .A(u5_mult_82_n1317), .ZN(u5_mult_82_n249) );
  NAND2_X4 u5_mult_82_U529 ( .A1(u5_mult_82_n251), .A2(u5_mult_82_n252), .ZN(
        u5_mult_82_SUMB_20__25_) );
  NAND2_X4 u5_mult_82_U528 ( .A1(u5_mult_82_n249), .A2(u5_mult_82_n250), .ZN(
        u5_mult_82_n252) );
  NAND2_X2 u5_mult_82_U527 ( .A1(u5_mult_82_n1317), .A2(u5_mult_82_n1315), 
        .ZN(u5_mult_82_n251) );
  INV_X4 u5_mult_82_U526 ( .A(u5_mult_82_net84453), .ZN(u5_mult_82_n246) );
  INV_X4 u5_mult_82_U525 ( .A(u5_mult_82_SUMB_21__24_), .ZN(u5_mult_82_n245)
         );
  NAND2_X2 u5_mult_82_U524 ( .A1(u5_mult_82_n247), .A2(u5_mult_82_n248), .ZN(
        u5_mult_82_n3614) );
  NAND2_X4 u5_mult_82_U523 ( .A1(u5_mult_82_n245), .A2(u5_mult_82_n246), .ZN(
        u5_mult_82_n248) );
  NAND2_X1 u5_mult_82_U522 ( .A1(u5_mult_82_SUMB_21__24_), .A2(
        u5_mult_82_net84453), .ZN(u5_mult_82_n247) );
  INV_X4 u5_mult_82_U521 ( .A(u5_mult_82_n1842), .ZN(u5_mult_82_n1843) );
  NAND3_X4 u5_mult_82_U520 ( .A1(u5_mult_82_n5188), .A2(u5_mult_82_n5189), 
        .A3(u5_mult_82_n5190), .ZN(u5_mult_82_CARRYB_39__18_) );
  NAND2_X4 u5_mult_82_U519 ( .A1(u5_mult_82_CARRYB_38__18_), .A2(
        u5_mult_82_n735), .ZN(u5_mult_82_n5190) );
  NAND2_X2 u5_mult_82_U518 ( .A1(u5_mult_82_ab_18__28_), .A2(u5_mult_82_n31), 
        .ZN(u5_mult_82_n5798) );
  NAND3_X2 u5_mult_82_U517 ( .A1(u5_mult_82_n242), .A2(u5_mult_82_n243), .A3(
        u5_mult_82_n244), .ZN(u5_mult_82_CARRYB_35__17_) );
  NAND2_X2 u5_mult_82_U516 ( .A1(u5_mult_82_CARRYB_34__17_), .A2(
        u5_mult_82_SUMB_34__18_), .ZN(u5_mult_82_n244) );
  NAND2_X2 u5_mult_82_U515 ( .A1(u5_mult_82_ab_35__17_), .A2(
        u5_mult_82_SUMB_34__18_), .ZN(u5_mult_82_n243) );
  NAND2_X1 u5_mult_82_U514 ( .A1(u5_mult_82_ab_35__17_), .A2(
        u5_mult_82_CARRYB_34__17_), .ZN(u5_mult_82_n242) );
  NAND3_X2 u5_mult_82_U513 ( .A1(u5_mult_82_n239), .A2(u5_mult_82_n240), .A3(
        u5_mult_82_n241), .ZN(u5_mult_82_CARRYB_34__18_) );
  NAND2_X2 u5_mult_82_U512 ( .A1(u5_mult_82_CARRYB_33__18_), .A2(
        u5_mult_82_SUMB_33__19_), .ZN(u5_mult_82_n241) );
  NAND2_X2 u5_mult_82_U511 ( .A1(u5_mult_82_ab_34__18_), .A2(
        u5_mult_82_SUMB_33__19_), .ZN(u5_mult_82_n240) );
  NAND2_X1 u5_mult_82_U510 ( .A1(u5_mult_82_ab_34__18_), .A2(
        u5_mult_82_CARRYB_33__18_), .ZN(u5_mult_82_n239) );
  XOR2_X2 u5_mult_82_U509 ( .A(u5_mult_82_n238), .B(u5_mult_82_SUMB_34__18_), 
        .Z(u5_mult_82_SUMB_35__17_) );
  XOR2_X1 u5_mult_82_U508 ( .A(u5_mult_82_ab_35__17_), .B(
        u5_mult_82_CARRYB_34__17_), .Z(u5_mult_82_n238) );
  XOR2_X2 u5_mult_82_U507 ( .A(u5_mult_82_n237), .B(u5_mult_82_SUMB_33__19_), 
        .Z(u5_mult_82_SUMB_34__18_) );
  XOR2_X2 u5_mult_82_U506 ( .A(u5_mult_82_ab_34__18_), .B(
        u5_mult_82_CARRYB_33__18_), .Z(u5_mult_82_n237) );
  NAND2_X1 u5_mult_82_U505 ( .A1(u5_mult_82_CARRYB_34__26_), .A2(
        u5_mult_82_n1647), .ZN(u5_mult_82_n5994) );
  NAND2_X2 u5_mult_82_U504 ( .A1(u5_mult_82_ab_48__20_), .A2(
        u5_mult_82_SUMB_47__21_), .ZN(u5_mult_82_n5749) );
  NAND2_X2 u5_mult_82_U503 ( .A1(u5_mult_82_CARRYB_47__20_), .A2(
        u5_mult_82_SUMB_47__21_), .ZN(u5_mult_82_n5750) );
  XOR2_X2 u5_mult_82_U502 ( .A(u5_mult_82_CARRYB_37__24_), .B(
        u5_mult_82_ab_38__24_), .Z(u5_mult_82_n3632) );
  NAND2_X2 u5_mult_82_U501 ( .A1(u5_mult_82_ab_28__40_), .A2(
        u5_mult_82_SUMB_27__41_), .ZN(u5_mult_82_n1108) );
  NAND2_X1 u5_mult_82_U500 ( .A1(u5_mult_82_CARRYB_34__36_), .A2(
        u5_mult_82_SUMB_34__37_), .ZN(u5_mult_82_n5083) );
  XNOR2_X2 u5_mult_82_U499 ( .A(u5_mult_82_n931), .B(u5_mult_82_SUMB_36__36_), 
        .ZN(u5_mult_82_SUMB_37__35_) );
  INV_X8 u5_mult_82_U498 ( .A(u5_mult_82_n6413), .ZN(u5_mult_82_CLA_SUM[79])
         );
  NAND3_X2 u5_mult_82_U497 ( .A1(u5_mult_82_n5029), .A2(u5_mult_82_n5030), 
        .A3(u5_mult_82_n5031), .ZN(u5_mult_82_CARRYB_35__25_) );
  NAND3_X2 u5_mult_82_U496 ( .A1(u5_mult_82_n5517), .A2(u5_mult_82_n5518), 
        .A3(u5_mult_82_n5519), .ZN(u5_mult_82_CARRYB_21__37_) );
  NAND2_X2 u5_mult_82_U495 ( .A1(u5_mult_82_CARRYB_28__32_), .A2(
        u5_mult_82_SUMB_28__33_), .ZN(u5_mult_82_n2429) );
  NAND2_X1 u5_mult_82_U494 ( .A1(u5_mult_82_ab_29__32_), .A2(
        u5_mult_82_SUMB_28__33_), .ZN(u5_mult_82_n2428) );
  NAND2_X2 u5_mult_82_U493 ( .A1(u5_mult_82_ab_19__27_), .A2(
        u5_mult_82_SUMB_18__28_), .ZN(u5_mult_82_n5801) );
  NAND2_X2 u5_mult_82_U492 ( .A1(u5_mult_82_ab_34__10_), .A2(
        u5_mult_82_CARRYB_33__10_), .ZN(u5_mult_82_n4072) );
  NAND2_X1 u5_mult_82_U491 ( .A1(u5_mult_82_CARRYB_33__10_), .A2(
        u5_mult_82_SUMB_33__11_), .ZN(u5_mult_82_n4070) );
  XNOR2_X1 u5_mult_82_U490 ( .A(u5_mult_82_CARRYB_33__10_), .B(
        u5_mult_82_ab_34__10_), .ZN(u5_mult_82_n428) );
  INV_X4 u5_mult_82_U489 ( .A(u5_mult_82_SUMB_39__20_), .ZN(u5_mult_82_n426)
         );
  INV_X2 u5_mult_82_U488 ( .A(u5_mult_82_SUMB_48__13_), .ZN(u5_mult_82_n1842)
         );
  NAND3_X4 u5_mult_82_U487 ( .A1(u5_mult_82_n234), .A2(u5_mult_82_n235), .A3(
        u5_mult_82_n236), .ZN(u5_mult_82_CARRYB_45__23_) );
  NAND2_X2 u5_mult_82_U486 ( .A1(u5_mult_82_CARRYB_44__23_), .A2(
        u5_mult_82_SUMB_44__24_), .ZN(u5_mult_82_n236) );
  NAND2_X2 u5_mult_82_U485 ( .A1(u5_mult_82_ab_45__23_), .A2(
        u5_mult_82_SUMB_44__24_), .ZN(u5_mult_82_n235) );
  NAND2_X1 u5_mult_82_U484 ( .A1(u5_mult_82_ab_45__23_), .A2(
        u5_mult_82_CARRYB_44__23_), .ZN(u5_mult_82_n234) );
  NAND3_X4 u5_mult_82_U483 ( .A1(u5_mult_82_n231), .A2(u5_mult_82_n232), .A3(
        u5_mult_82_n233), .ZN(u5_mult_82_CARRYB_44__24_) );
  NAND2_X2 u5_mult_82_U482 ( .A1(u5_mult_82_CARRYB_43__24_), .A2(
        u5_mult_82_SUMB_43__25_), .ZN(u5_mult_82_n233) );
  NAND2_X2 u5_mult_82_U481 ( .A1(u5_mult_82_ab_44__24_), .A2(
        u5_mult_82_SUMB_43__25_), .ZN(u5_mult_82_n232) );
  NAND2_X1 u5_mult_82_U480 ( .A1(u5_mult_82_ab_44__24_), .A2(
        u5_mult_82_CARRYB_43__24_), .ZN(u5_mult_82_n231) );
  XOR2_X2 u5_mult_82_U479 ( .A(u5_mult_82_n230), .B(u5_mult_82_SUMB_44__24_), 
        .Z(u5_mult_82_SUMB_45__23_) );
  XOR2_X2 u5_mult_82_U478 ( .A(u5_mult_82_ab_45__23_), .B(
        u5_mult_82_CARRYB_44__23_), .Z(u5_mult_82_n230) );
  XOR2_X2 u5_mult_82_U477 ( .A(u5_mult_82_n229), .B(u5_mult_82_SUMB_43__25_), 
        .Z(u5_mult_82_SUMB_44__24_) );
  XOR2_X2 u5_mult_82_U476 ( .A(u5_mult_82_CARRYB_43__24_), .B(
        u5_mult_82_ab_44__24_), .Z(u5_mult_82_n229) );
  NAND2_X4 u5_mult_82_U475 ( .A1(u5_mult_82_n261), .A2(u5_mult_82_n260), .ZN(
        u5_mult_82_SUMB_39__19_) );
  NAND2_X2 u5_mult_82_U474 ( .A1(u5_mult_82_CARRYB_23__38_), .A2(
        u5_mult_82_SUMB_23__39_), .ZN(u5_mult_82_n5846) );
  XNOR2_X2 u5_mult_82_U473 ( .A(u5_mult_82_ab_41__7_), .B(
        u5_mult_82_CARRYB_40__7_), .ZN(u5_mult_82_n1768) );
  NAND3_X2 u5_mult_82_U472 ( .A1(u5_mult_82_n4289), .A2(u5_mult_82_n4290), 
        .A3(u5_mult_82_n4291), .ZN(u5_mult_82_CARRYB_45__15_) );
  NAND2_X2 u5_mult_82_U471 ( .A1(u5_mult_82_CARRYB_36__18_), .A2(
        u5_mult_82_SUMB_36__19_), .ZN(u5_mult_82_n5011) );
  NAND2_X1 u5_mult_82_U470 ( .A1(u5_mult_82_ab_38__23_), .A2(
        u5_mult_82_SUMB_37__24_), .ZN(u5_mult_82_n563) );
  NAND2_X1 u5_mult_82_U469 ( .A1(u5_mult_82_ab_51__25_), .A2(
        u5_mult_82_SUMB_50__26_), .ZN(u5_mult_82_n4188) );
  NAND2_X1 u5_mult_82_U468 ( .A1(u5_mult_82_n3606), .A2(
        u5_mult_82_SUMB_50__26_), .ZN(u5_mult_82_n3609) );
  INV_X4 u5_mult_82_U467 ( .A(u5_mult_82_n6410), .ZN(u5_mult_82_CLA_SUM[76])
         );
  INV_X4 u5_mult_82_U466 ( .A(u5_mult_82_SUMB_38__19_), .ZN(u5_mult_82_n734)
         );
  NAND2_X1 u5_mult_82_U465 ( .A1(u5_mult_82_ab_43__5_), .A2(
        u5_mult_82_CARRYB_42__5_), .ZN(u5_mult_82_n5244) );
  CLKBUF_X3 u5_mult_82_U464 ( .A(u5_mult_82_CARRYB_42__5_), .Z(
        u5_mult_82_n1835) );
  NAND2_X2 u5_mult_82_U463 ( .A1(u5_mult_82_CARRYB_21__12_), .A2(
        u5_mult_82_ab_22__12_), .ZN(u5_mult_82_n2470) );
  NAND2_X1 u5_mult_82_U462 ( .A1(u5_mult_82_CARRYB_35__25_), .A2(
        u5_mult_82_SUMB_35__26_), .ZN(u5_mult_82_n4554) );
  XNOR2_X2 u5_mult_82_U461 ( .A(u5_mult_82_ab_39__16_), .B(
        u5_mult_82_CARRYB_38__16_), .ZN(u5_mult_82_n1470) );
  INV_X32 u5_mult_82_U460 ( .A(u5_mult_82_ab_47__34_), .ZN(u5_mult_82_n228) );
  XNOR2_X2 u5_mult_82_U459 ( .A(u5_mult_82_n228), .B(u5_mult_82_CARRYB_46__34_), .ZN(u5_mult_82_n2920) );
  NAND2_X1 u5_mult_82_U458 ( .A1(u5_mult_82_ab_28__41_), .A2(
        u5_mult_82_CARRYB_27__41_), .ZN(u5_mult_82_n2447) );
  NOR2_X1 u5_mult_82_U457 ( .A1(u5_mult_82_n6768), .A2(u5_mult_82_n1344), .ZN(
        u5_mult_82_ab_23__50_) );
  NAND3_X2 u5_mult_82_U456 ( .A1(u5_mult_82_n225), .A2(u5_mult_82_n226), .A3(
        u5_mult_82_n227), .ZN(u5_mult_82_CARRYB_23__50_) );
  NAND2_X1 u5_mult_82_U455 ( .A1(u5_mult_82_ab_23__50_), .A2(
        u5_mult_82_SUMB_22__51_), .ZN(u5_mult_82_n227) );
  NAND2_X2 u5_mult_82_U454 ( .A1(u5_mult_82_ab_23__50_), .A2(
        u5_mult_82_CARRYB_22__50_), .ZN(u5_mult_82_n226) );
  NAND2_X1 u5_mult_82_U453 ( .A1(u5_mult_82_SUMB_22__51_), .A2(
        u5_mult_82_CARRYB_22__50_), .ZN(u5_mult_82_n225) );
  XOR2_X2 u5_mult_82_U452 ( .A(u5_mult_82_CARRYB_22__50_), .B(u5_mult_82_n224), 
        .Z(u5_mult_82_SUMB_23__50_) );
  XOR2_X2 u5_mult_82_U451 ( .A(u5_mult_82_SUMB_22__51_), .B(
        u5_mult_82_ab_23__50_), .Z(u5_mult_82_n224) );
  NAND3_X2 u5_mult_82_U450 ( .A1(u5_mult_82_n221), .A2(u5_mult_82_n222), .A3(
        u5_mult_82_n223), .ZN(u5_mult_82_CARRYB_30__49_) );
  NAND2_X1 u5_mult_82_U449 ( .A1(u5_mult_82_CARRYB_29__49_), .A2(
        u5_mult_82_SUMB_29__50_), .ZN(u5_mult_82_n223) );
  NAND2_X1 u5_mult_82_U448 ( .A1(u5_mult_82_ab_30__49_), .A2(
        u5_mult_82_SUMB_29__50_), .ZN(u5_mult_82_n222) );
  NAND2_X1 u5_mult_82_U447 ( .A1(u5_mult_82_ab_30__49_), .A2(
        u5_mult_82_CARRYB_29__49_), .ZN(u5_mult_82_n221) );
  NAND3_X4 u5_mult_82_U446 ( .A1(u5_mult_82_n218), .A2(u5_mult_82_n219), .A3(
        u5_mult_82_n220), .ZN(u5_mult_82_CARRYB_29__50_) );
  NAND2_X2 u5_mult_82_U445 ( .A1(u5_mult_82_CARRYB_28__50_), .A2(
        u5_mult_82_SUMB_28__51_), .ZN(u5_mult_82_n220) );
  NAND2_X2 u5_mult_82_U444 ( .A1(u5_mult_82_ab_29__50_), .A2(
        u5_mult_82_SUMB_28__51_), .ZN(u5_mult_82_n219) );
  NAND2_X2 u5_mult_82_U443 ( .A1(u5_mult_82_ab_29__50_), .A2(
        u5_mult_82_CARRYB_28__50_), .ZN(u5_mult_82_n218) );
  XOR2_X2 u5_mult_82_U442 ( .A(u5_mult_82_n217), .B(u5_mult_82_SUMB_29__50_), 
        .Z(u5_mult_82_SUMB_30__49_) );
  XOR2_X2 u5_mult_82_U441 ( .A(u5_mult_82_ab_30__49_), .B(
        u5_mult_82_CARRYB_29__49_), .Z(u5_mult_82_n217) );
  XOR2_X2 u5_mult_82_U440 ( .A(u5_mult_82_n216), .B(u5_mult_82_SUMB_28__51_), 
        .Z(u5_mult_82_SUMB_29__50_) );
  XOR2_X2 u5_mult_82_U439 ( .A(u5_mult_82_ab_29__50_), .B(
        u5_mult_82_CARRYB_28__50_), .Z(u5_mult_82_n216) );
  INV_X4 u5_mult_82_U438 ( .A(u5_mult_82_n214), .ZN(u5_mult_82_n215) );
  INV_X2 u5_mult_82_U437 ( .A(u5_mult_82_ab_1__52_), .ZN(u5_mult_82_n214) );
  NAND3_X4 u5_mult_82_U436 ( .A1(u5_mult_82_n5997), .A2(u5_mult_82_n5998), 
        .A3(u5_mult_82_n5999), .ZN(u5_mult_82_CARRYB_22__39_) );
  CLKBUF_X3 u5_mult_82_U435 ( .A(u5_mult_82_SUMB_46__3_), .Z(u5_mult_82_n412)
         );
  NAND2_X2 u5_mult_82_U434 ( .A1(u5_mult_82_CARRYB_30__14_), .A2(
        u5_mult_82_SUMB_30__15_), .ZN(u5_mult_82_n3660) );
  NAND2_X2 u5_mult_82_U433 ( .A1(u5_mult_82_ab_8__28_), .A2(
        u5_mult_82_SUMB_7__29_), .ZN(u5_mult_82_n2508) );
  NAND3_X2 u5_mult_82_U432 ( .A1(u5_mult_82_n4768), .A2(u5_mult_82_n4769), 
        .A3(u5_mult_82_n4770), .ZN(u5_mult_82_CARRYB_38__10_) );
  XNOR2_X2 u5_mult_82_U431 ( .A(u5_mult_82_net84580), .B(
        u5_mult_82_SUMB_31__18_), .ZN(u5_mult_82_SUMB_32__17_) );
  NAND3_X4 u5_mult_82_U430 ( .A1(u5_mult_82_n4560), .A2(u5_mult_82_n4561), 
        .A3(u5_mult_82_n4562), .ZN(u5_mult_82_CARRYB_29__18_) );
  NAND2_X4 u5_mult_82_U429 ( .A1(u5_mult_82_n3540), .A2(u5_mult_82_n3539), 
        .ZN(u5_mult_82_n3542) );
  INV_X4 u5_mult_82_U428 ( .A(u5_mult_82_CARRYB_18__44_), .ZN(u5_mult_82_n5247) );
  NAND2_X1 u5_mult_82_U427 ( .A1(u5_mult_82_ab_41__36_), .A2(
        u5_mult_82_SUMB_40__37_), .ZN(u5_mult_82_n2975) );
  NAND2_X2 u5_mult_82_U426 ( .A1(u5_mult_82_n697), .A2(
        u5_mult_82_CARRYB_44__14_), .ZN(u5_mult_82_n4207) );
  AND2_X4 u5_mult_82_U425 ( .A1(u5_mult_82_n2212), .A2(u5_mult_82_n2213), .ZN(
        u5_mult_82_n213) );
  XNOR2_X2 u5_mult_82_U424 ( .A(u5_mult_82_n213), .B(u5_mult_82_SUMB_25__41_), 
        .ZN(u5_mult_82_SUMB_26__40_) );
  NAND2_X1 u5_mult_82_U423 ( .A1(u5_mult_82_CARRYB_37__1_), .A2(
        u5_mult_82_SUMB_37__2_), .ZN(u5_mult_82_n2550) );
  XNOR2_X2 u5_mult_82_U422 ( .A(u5_mult_82_CARRYB_37__1_), .B(u5_mult_82_n631), 
        .ZN(u5_mult_82_n2547) );
  NOR2_X1 u5_mult_82_U421 ( .A1(u5_mult_82_n6967), .A2(u5_mult_82_n6723), .ZN(
        u5_mult_82_ab_37__1_) );
  NOR2_X1 u5_mult_82_U420 ( .A1(u5_mult_82_n6968), .A2(u5_mult_82_n6645), .ZN(
        u5_mult_82_ab_24__1_) );
  NOR2_X1 u5_mult_82_U419 ( .A1(u5_mult_82_n6941), .A2(u5_mult_82_n6603), .ZN(
        u5_mult_82_ab_17__7_) );
  INV_X2 u5_mult_82_U418 ( .A(u5_mult_82_CARRYB_46__1_), .ZN(u5_mult_82_n1807)
         );
  NAND3_X2 u5_mult_82_U417 ( .A1(u5_mult_82_n210), .A2(u5_mult_82_n211), .A3(
        u5_mult_82_n212), .ZN(u5_mult_82_CARRYB_37__1_) );
  NAND2_X1 u5_mult_82_U416 ( .A1(u5_mult_82_ab_37__1_), .A2(
        u5_mult_82_SUMB_36__2_), .ZN(u5_mult_82_n212) );
  NAND2_X2 u5_mult_82_U415 ( .A1(u5_mult_82_ab_37__1_), .A2(
        u5_mult_82_CARRYB_36__1_), .ZN(u5_mult_82_n211) );
  NAND2_X2 u5_mult_82_U414 ( .A1(u5_mult_82_SUMB_36__2_), .A2(
        u5_mult_82_CARRYB_36__1_), .ZN(u5_mult_82_n210) );
  XOR2_X2 u5_mult_82_U413 ( .A(u5_mult_82_CARRYB_36__1_), .B(u5_mult_82_n209), 
        .Z(u5_mult_82_SUMB_37__1_) );
  XOR2_X2 u5_mult_82_U412 ( .A(u5_mult_82_SUMB_36__2_), .B(
        u5_mult_82_ab_37__1_), .Z(u5_mult_82_n209) );
  NAND3_X2 u5_mult_82_U411 ( .A1(u5_mult_82_n2551), .A2(u5_mult_82_n2552), 
        .A3(u5_mult_82_n2553), .ZN(u5_mult_82_n208) );
  NAND3_X2 u5_mult_82_U410 ( .A1(u5_mult_82_n205), .A2(u5_mult_82_n206), .A3(
        u5_mult_82_n207), .ZN(u5_mult_82_CARRYB_26__1_) );
  NAND2_X1 u5_mult_82_U409 ( .A1(u5_mult_82_ab_26__1_), .A2(
        u5_mult_82_CARRYB_25__1_), .ZN(u5_mult_82_n207) );
  NAND2_X2 u5_mult_82_U408 ( .A1(u5_mult_82_ab_26__1_), .A2(
        u5_mult_82_SUMB_25__2_), .ZN(u5_mult_82_n206) );
  NAND2_X1 u5_mult_82_U407 ( .A1(u5_mult_82_CARRYB_25__1_), .A2(
        u5_mult_82_SUMB_25__2_), .ZN(u5_mult_82_n205) );
  XOR2_X2 u5_mult_82_U406 ( .A(u5_mult_82_SUMB_25__2_), .B(u5_mult_82_n204), 
        .Z(u5_mult_82_SUMB_26__1_) );
  XOR2_X2 u5_mult_82_U405 ( .A(u5_mult_82_CARRYB_25__1_), .B(
        u5_mult_82_ab_26__1_), .Z(u5_mult_82_n204) );
  NAND3_X2 u5_mult_82_U404 ( .A1(u5_mult_82_n201), .A2(u5_mult_82_n202), .A3(
        u5_mult_82_n203), .ZN(u5_mult_82_CARRYB_25__1_) );
  NAND2_X1 u5_mult_82_U403 ( .A1(u5_mult_82_ab_25__1_), .A2(
        u5_mult_82_CARRYB_24__1_), .ZN(u5_mult_82_n203) );
  NAND2_X2 u5_mult_82_U402 ( .A1(u5_mult_82_ab_25__1_), .A2(
        u5_mult_82_SUMB_24__2_), .ZN(u5_mult_82_n202) );
  NAND2_X1 u5_mult_82_U401 ( .A1(u5_mult_82_CARRYB_24__1_), .A2(
        u5_mult_82_SUMB_24__2_), .ZN(u5_mult_82_n201) );
  XOR2_X2 u5_mult_82_U400 ( .A(u5_mult_82_SUMB_24__2_), .B(u5_mult_82_n200), 
        .Z(u5_mult_82_SUMB_25__1_) );
  XOR2_X2 u5_mult_82_U399 ( .A(u5_mult_82_CARRYB_24__1_), .B(
        u5_mult_82_ab_25__1_), .Z(u5_mult_82_n200) );
  NAND3_X2 u5_mult_82_U398 ( .A1(u5_mult_82_n197), .A2(u5_mult_82_n198), .A3(
        u5_mult_82_n199), .ZN(u5_mult_82_CARRYB_24__1_) );
  NAND2_X1 u5_mult_82_U397 ( .A1(u5_mult_82_ab_24__1_), .A2(
        u5_mult_82_CARRYB_23__1_), .ZN(u5_mult_82_n199) );
  NAND2_X2 u5_mult_82_U396 ( .A1(u5_mult_82_ab_24__1_), .A2(
        u5_mult_82_SUMB_23__2_), .ZN(u5_mult_82_n198) );
  NAND2_X1 u5_mult_82_U395 ( .A1(u5_mult_82_CARRYB_23__1_), .A2(
        u5_mult_82_SUMB_23__2_), .ZN(u5_mult_82_n197) );
  XOR2_X2 u5_mult_82_U394 ( .A(u5_mult_82_SUMB_23__2_), .B(u5_mult_82_n196), 
        .Z(u5_mult_82_SUMB_24__1_) );
  XOR2_X2 u5_mult_82_U393 ( .A(u5_mult_82_CARRYB_23__1_), .B(
        u5_mult_82_ab_24__1_), .Z(u5_mult_82_n196) );
  NAND3_X2 u5_mult_82_U392 ( .A1(u5_mult_82_n193), .A2(u5_mult_82_n194), .A3(
        u5_mult_82_n195), .ZN(u5_mult_82_CARRYB_17__7_) );
  NAND2_X1 u5_mult_82_U391 ( .A1(u5_mult_82_ab_17__7_), .A2(
        u5_mult_82_CARRYB_16__7_), .ZN(u5_mult_82_n195) );
  NAND2_X2 u5_mult_82_U390 ( .A1(u5_mult_82_ab_17__7_), .A2(
        u5_mult_82_SUMB_16__8_), .ZN(u5_mult_82_n194) );
  NAND2_X1 u5_mult_82_U389 ( .A1(u5_mult_82_CARRYB_16__7_), .A2(
        u5_mult_82_SUMB_16__8_), .ZN(u5_mult_82_n193) );
  XOR2_X2 u5_mult_82_U388 ( .A(u5_mult_82_SUMB_16__8_), .B(u5_mult_82_n192), 
        .Z(u5_mult_82_SUMB_17__7_) );
  XOR2_X2 u5_mult_82_U387 ( .A(u5_mult_82_CARRYB_16__7_), .B(
        u5_mult_82_ab_17__7_), .Z(u5_mult_82_n192) );
  NAND3_X2 u5_mult_82_U386 ( .A1(u5_mult_82_n189), .A2(u5_mult_82_n190), .A3(
        u5_mult_82_n191), .ZN(u5_mult_82_CARRYB_46__1_) );
  NAND2_X2 u5_mult_82_U385 ( .A1(u5_mult_82_ab_46__1_), .A2(
        u5_mult_82_SUMB_45__2_), .ZN(u5_mult_82_n191) );
  NAND2_X1 u5_mult_82_U384 ( .A1(u5_mult_82_ab_46__1_), .A2(
        u5_mult_82_CARRYB_45__1_), .ZN(u5_mult_82_n190) );
  NAND2_X1 u5_mult_82_U383 ( .A1(u5_mult_82_SUMB_45__2_), .A2(
        u5_mult_82_CARRYB_45__1_), .ZN(u5_mult_82_n189) );
  XOR2_X2 u5_mult_82_U382 ( .A(u5_mult_82_CARRYB_45__1_), .B(u5_mult_82_n188), 
        .Z(u5_mult_82_SUMB_46__1_) );
  XOR2_X2 u5_mult_82_U381 ( .A(u5_mult_82_SUMB_45__2_), .B(
        u5_mult_82_ab_46__1_), .Z(u5_mult_82_n188) );
  NAND3_X2 u5_mult_82_U380 ( .A1(u5_mult_82_n185), .A2(u5_mult_82_n186), .A3(
        u5_mult_82_n187), .ZN(u5_mult_82_CARRYB_13__10_) );
  NAND2_X2 u5_mult_82_U379 ( .A1(u5_mult_82_ab_13__10_), .A2(
        u5_mult_82_CARRYB_12__10_), .ZN(u5_mult_82_n187) );
  NAND2_X2 u5_mult_82_U378 ( .A1(u5_mult_82_ab_13__10_), .A2(
        u5_mult_82_SUMB_12__11_), .ZN(u5_mult_82_n186) );
  NAND2_X2 u5_mult_82_U377 ( .A1(u5_mult_82_CARRYB_12__10_), .A2(
        u5_mult_82_SUMB_12__11_), .ZN(u5_mult_82_n185) );
  XOR2_X2 u5_mult_82_U376 ( .A(u5_mult_82_SUMB_12__11_), .B(u5_mult_82_n184), 
        .Z(u5_mult_82_SUMB_13__10_) );
  XOR2_X2 u5_mult_82_U375 ( .A(u5_mult_82_CARRYB_12__10_), .B(
        u5_mult_82_ab_13__10_), .Z(u5_mult_82_n184) );
  XNOR2_X2 u5_mult_82_U374 ( .A(u5_mult_82_ab_37__34_), .B(
        u5_mult_82_CARRYB_36__34_), .ZN(u5_mult_82_n638) );
  NAND2_X1 u5_mult_82_U373 ( .A1(u5_mult_82_CARRYB_47__19_), .A2(
        u5_mult_82_SUMB_47__20_), .ZN(u5_mult_82_n4393) );
  NAND2_X2 u5_mult_82_U372 ( .A1(u5_mult_82_ab_30__38_), .A2(
        u5_mult_82_CARRYB_29__38_), .ZN(u5_mult_82_n2402) );
  NOR2_X2 u5_mult_82_U371 ( .A1(u5_mult_82_net64957), .A2(u5_mult_82_n6671), 
        .ZN(u5_mult_82_ab_29__38_) );
  NAND3_X2 u5_mult_82_U370 ( .A1(u5_mult_82_n181), .A2(u5_mult_82_n182), .A3(
        u5_mult_82_n183), .ZN(u5_mult_82_CARRYB_29__38_) );
  NAND2_X1 u5_mult_82_U369 ( .A1(u5_mult_82_ab_29__38_), .A2(
        u5_mult_82_SUMB_28__39_), .ZN(u5_mult_82_n183) );
  NAND2_X1 u5_mult_82_U368 ( .A1(u5_mult_82_ab_29__38_), .A2(
        u5_mult_82_CARRYB_28__38_), .ZN(u5_mult_82_n182) );
  NAND2_X1 u5_mult_82_U367 ( .A1(u5_mult_82_SUMB_28__39_), .A2(
        u5_mult_82_CARRYB_28__38_), .ZN(u5_mult_82_n181) );
  XOR2_X2 u5_mult_82_U366 ( .A(u5_mult_82_CARRYB_28__38_), .B(u5_mult_82_n180), 
        .Z(u5_mult_82_SUMB_29__38_) );
  XOR2_X2 u5_mult_82_U365 ( .A(u5_mult_82_SUMB_28__39_), .B(
        u5_mult_82_ab_29__38_), .Z(u5_mult_82_n180) );
  NAND3_X2 u5_mult_82_U364 ( .A1(u5_mult_82_n177), .A2(u5_mult_82_n178), .A3(
        u5_mult_82_n179), .ZN(u5_mult_82_CARRYB_26__39_) );
  NAND2_X1 u5_mult_82_U363 ( .A1(u5_mult_82_ab_26__39_), .A2(
        u5_mult_82_CARRYB_25__39_), .ZN(u5_mult_82_n179) );
  NAND2_X2 u5_mult_82_U362 ( .A1(u5_mult_82_ab_26__39_), .A2(
        u5_mult_82_SUMB_25__40_), .ZN(u5_mult_82_n178) );
  NAND2_X1 u5_mult_82_U361 ( .A1(u5_mult_82_CARRYB_25__39_), .A2(
        u5_mult_82_SUMB_25__40_), .ZN(u5_mult_82_n177) );
  XOR2_X2 u5_mult_82_U360 ( .A(u5_mult_82_SUMB_25__40_), .B(u5_mult_82_n176), 
        .Z(u5_mult_82_SUMB_26__39_) );
  XOR2_X2 u5_mult_82_U359 ( .A(u5_mult_82_CARRYB_25__39_), .B(
        u5_mult_82_ab_26__39_), .Z(u5_mult_82_n176) );
  NAND3_X2 u5_mult_82_U358 ( .A1(u5_mult_82_n173), .A2(u5_mult_82_n174), .A3(
        u5_mult_82_n175), .ZN(u5_mult_82_CARRYB_34__34_) );
  NAND2_X1 u5_mult_82_U357 ( .A1(u5_mult_82_CARRYB_33__34_), .A2(
        u5_mult_82_SUMB_33__35_), .ZN(u5_mult_82_n175) );
  NAND2_X2 u5_mult_82_U356 ( .A1(u5_mult_82_ab_34__34_), .A2(
        u5_mult_82_SUMB_33__35_), .ZN(u5_mult_82_n174) );
  NAND2_X1 u5_mult_82_U355 ( .A1(u5_mult_82_ab_34__34_), .A2(
        u5_mult_82_CARRYB_33__34_), .ZN(u5_mult_82_n173) );
  NAND3_X4 u5_mult_82_U354 ( .A1(u5_mult_82_n170), .A2(u5_mult_82_n171), .A3(
        u5_mult_82_n172), .ZN(u5_mult_82_CARRYB_33__35_) );
  NAND2_X2 u5_mult_82_U353 ( .A1(u5_mult_82_ab_33__35_), .A2(
        u5_mult_82_SUMB_32__36_), .ZN(u5_mult_82_n172) );
  NAND2_X2 u5_mult_82_U352 ( .A1(u5_mult_82_CARRYB_32__35_), .A2(
        u5_mult_82_SUMB_32__36_), .ZN(u5_mult_82_n171) );
  NAND2_X2 u5_mult_82_U351 ( .A1(u5_mult_82_CARRYB_32__35_), .A2(
        u5_mult_82_ab_33__35_), .ZN(u5_mult_82_n170) );
  XOR2_X2 u5_mult_82_U350 ( .A(u5_mult_82_n169), .B(u5_mult_82_SUMB_32__36_), 
        .Z(u5_mult_82_SUMB_33__35_) );
  XOR2_X2 u5_mult_82_U349 ( .A(u5_mult_82_CARRYB_32__35_), .B(
        u5_mult_82_ab_33__35_), .Z(u5_mult_82_n169) );
  INV_X32 u5_mult_82_U348 ( .A(u5_mult_82_ab_38__37_), .ZN(u5_mult_82_n168) );
  XNOR2_X2 u5_mult_82_U347 ( .A(u5_mult_82_n168), .B(u5_mult_82_CARRYB_37__37_), .ZN(u5_mult_82_n4470) );
  NAND2_X2 u5_mult_82_U346 ( .A1(u5_mult_82_ab_26__16_), .A2(
        u5_mult_82_SUMB_25__17_), .ZN(u5_mult_82_n2782) );
  NAND3_X4 u5_mult_82_U345 ( .A1(u5_mult_82_n165), .A2(u5_mult_82_n166), .A3(
        u5_mult_82_n167), .ZN(u5_mult_82_CARRYB_40__37_) );
  NAND2_X2 u5_mult_82_U344 ( .A1(u5_mult_82_CARRYB_39__37_), .A2(
        u5_mult_82_SUMB_39__38_), .ZN(u5_mult_82_n167) );
  NAND2_X2 u5_mult_82_U343 ( .A1(u5_mult_82_ab_40__37_), .A2(
        u5_mult_82_SUMB_39__38_), .ZN(u5_mult_82_n166) );
  NAND2_X1 u5_mult_82_U342 ( .A1(u5_mult_82_ab_40__37_), .A2(
        u5_mult_82_CARRYB_39__37_), .ZN(u5_mult_82_n165) );
  NAND3_X2 u5_mult_82_U341 ( .A1(u5_mult_82_n162), .A2(u5_mult_82_n163), .A3(
        u5_mult_82_n164), .ZN(u5_mult_82_CARRYB_39__38_) );
  NAND2_X2 u5_mult_82_U340 ( .A1(u5_mult_82_CARRYB_38__38_), .A2(
        u5_mult_82_SUMB_38__39_), .ZN(u5_mult_82_n164) );
  NAND2_X2 u5_mult_82_U339 ( .A1(u5_mult_82_ab_39__38_), .A2(
        u5_mult_82_SUMB_38__39_), .ZN(u5_mult_82_n163) );
  NAND2_X1 u5_mult_82_U338 ( .A1(u5_mult_82_ab_39__38_), .A2(
        u5_mult_82_CARRYB_38__38_), .ZN(u5_mult_82_n162) );
  XOR2_X2 u5_mult_82_U337 ( .A(u5_mult_82_n161), .B(u5_mult_82_SUMB_39__38_), 
        .Z(u5_mult_82_SUMB_40__37_) );
  XOR2_X2 u5_mult_82_U336 ( .A(u5_mult_82_ab_40__37_), .B(
        u5_mult_82_CARRYB_39__37_), .Z(u5_mult_82_n161) );
  XOR2_X2 u5_mult_82_U335 ( .A(u5_mult_82_n160), .B(u5_mult_82_SUMB_38__39_), 
        .Z(u5_mult_82_SUMB_39__38_) );
  XOR2_X2 u5_mult_82_U334 ( .A(u5_mult_82_ab_39__38_), .B(
        u5_mult_82_CARRYB_38__38_), .Z(u5_mult_82_n160) );
  NAND3_X2 u5_mult_82_U333 ( .A1(u5_mult_82_n157), .A2(u5_mult_82_n158), .A3(
        u5_mult_82_n159), .ZN(u5_mult_82_CARRYB_35__40_) );
  NAND2_X1 u5_mult_82_U332 ( .A1(u5_mult_82_CARRYB_34__40_), .A2(
        u5_mult_82_SUMB_34__41_), .ZN(u5_mult_82_n159) );
  NAND2_X2 u5_mult_82_U331 ( .A1(u5_mult_82_ab_35__40_), .A2(
        u5_mult_82_SUMB_34__41_), .ZN(u5_mult_82_n158) );
  NAND2_X1 u5_mult_82_U330 ( .A1(u5_mult_82_ab_35__40_), .A2(
        u5_mult_82_CARRYB_34__40_), .ZN(u5_mult_82_n157) );
  NAND3_X2 u5_mult_82_U329 ( .A1(u5_mult_82_n154), .A2(u5_mult_82_n155), .A3(
        u5_mult_82_n156), .ZN(u5_mult_82_CARRYB_34__41_) );
  NAND2_X2 u5_mult_82_U328 ( .A1(u5_mult_82_CARRYB_33__41_), .A2(
        u5_mult_82_SUMB_33__42_), .ZN(u5_mult_82_n156) );
  NAND2_X2 u5_mult_82_U327 ( .A1(u5_mult_82_ab_34__41_), .A2(
        u5_mult_82_SUMB_33__42_), .ZN(u5_mult_82_n155) );
  NAND2_X1 u5_mult_82_U326 ( .A1(u5_mult_82_ab_34__41_), .A2(
        u5_mult_82_CARRYB_33__41_), .ZN(u5_mult_82_n154) );
  XOR2_X2 u5_mult_82_U325 ( .A(u5_mult_82_n153), .B(u5_mult_82_SUMB_34__41_), 
        .Z(u5_mult_82_SUMB_35__40_) );
  XOR2_X2 u5_mult_82_U324 ( .A(u5_mult_82_ab_35__40_), .B(
        u5_mult_82_CARRYB_34__40_), .Z(u5_mult_82_n153) );
  XOR2_X2 u5_mult_82_U323 ( .A(u5_mult_82_n152), .B(u5_mult_82_SUMB_33__42_), 
        .Z(u5_mult_82_SUMB_34__41_) );
  XOR2_X2 u5_mult_82_U322 ( .A(u5_mult_82_ab_34__41_), .B(
        u5_mult_82_CARRYB_33__41_), .Z(u5_mult_82_n152) );
  NAND2_X2 u5_mult_82_U321 ( .A1(u5_mult_82_CARRYB_39__6_), .A2(
        u5_mult_82_ab_40__6_), .ZN(u5_mult_82_n5819) );
  NOR2_X4 u5_mult_82_U320 ( .A1(u5_mult_82_n6880), .A2(u5_mult_82_n6708), .ZN(
        u5_mult_82_ab_35__26_) );
  INV_X1 u5_mult_82_U319 ( .A(u5_mult_82_ab_35__26_), .ZN(u5_mult_82_n149) );
  INV_X1 u5_mult_82_U318 ( .A(u5_mult_82_CARRYB_34__26_), .ZN(u5_mult_82_n148)
         );
  NAND2_X2 u5_mult_82_U317 ( .A1(u5_mult_82_n150), .A2(u5_mult_82_n151), .ZN(
        u5_mult_82_n1482) );
  NAND2_X2 u5_mult_82_U316 ( .A1(u5_mult_82_n148), .A2(u5_mult_82_n149), .ZN(
        u5_mult_82_n151) );
  NAND2_X1 u5_mult_82_U315 ( .A1(u5_mult_82_CARRYB_34__26_), .A2(
        u5_mult_82_ab_35__26_), .ZN(u5_mult_82_n150) );
  NAND2_X2 u5_mult_82_U314 ( .A1(u5_mult_82_CARRYB_15__20_), .A2(
        u5_mult_82_SUMB_15__21_), .ZN(u5_mult_82_n3894) );
  NAND2_X2 u5_mult_82_U313 ( .A1(u5_mult_82_CARRYB_50__1_), .A2(
        u5_mult_82_SUMB_50__2_), .ZN(u5_mult_82_n994) );
  NAND2_X2 u5_mult_82_U312 ( .A1(u5_mult_82_CARRYB_22__22_), .A2(
        u5_mult_82_SUMB_22__23_), .ZN(u5_mult_82_n5334) );
  BUF_X8 u5_mult_82_U311 ( .A(u5_mult_82_SUMB_39__7_), .Z(u5_mult_82_n374) );
  NAND2_X4 u5_mult_82_U310 ( .A1(u5_mult_82_n697), .A2(u5_mult_82_ab_45__14_), 
        .ZN(u5_mult_82_n4206) );
  INV_X4 u5_mult_82_U309 ( .A(u5_mult_82_SUMB_9__37_), .ZN(u5_mult_82_n1868)
         );
  NAND2_X1 u5_mult_82_U308 ( .A1(u5_mult_82_ab_15__33_), .A2(
        u5_mult_82_SUMB_14__34_), .ZN(u5_mult_82_n4860) );
  NAND2_X1 u5_mult_82_U307 ( .A1(u5_mult_82_CARRYB_20__30_), .A2(
        u5_mult_82_SUMB_20__31_), .ZN(u5_mult_82_n2531) );
  NAND3_X4 u5_mult_82_U306 ( .A1(u5_mult_82_n145), .A2(u5_mult_82_n146), .A3(
        u5_mult_82_n147), .ZN(u5_mult_82_CARRYB_12__19_) );
  NAND2_X2 u5_mult_82_U305 ( .A1(u5_mult_82_CARRYB_11__19_), .A2(
        u5_mult_82_SUMB_11__20_), .ZN(u5_mult_82_n147) );
  NAND2_X2 u5_mult_82_U304 ( .A1(u5_mult_82_ab_12__19_), .A2(
        u5_mult_82_SUMB_11__20_), .ZN(u5_mult_82_n146) );
  NAND2_X1 u5_mult_82_U303 ( .A1(u5_mult_82_ab_12__19_), .A2(
        u5_mult_82_CARRYB_11__19_), .ZN(u5_mult_82_n145) );
  NAND3_X2 u5_mult_82_U302 ( .A1(u5_mult_82_n142), .A2(u5_mult_82_n143), .A3(
        u5_mult_82_n144), .ZN(u5_mult_82_CARRYB_11__20_) );
  NAND2_X2 u5_mult_82_U301 ( .A1(u5_mult_82_CARRYB_10__20_), .A2(
        u5_mult_82_SUMB_10__21_), .ZN(u5_mult_82_n144) );
  NAND2_X2 u5_mult_82_U300 ( .A1(u5_mult_82_ab_11__20_), .A2(
        u5_mult_82_SUMB_10__21_), .ZN(u5_mult_82_n143) );
  NAND2_X1 u5_mult_82_U299 ( .A1(u5_mult_82_ab_11__20_), .A2(
        u5_mult_82_CARRYB_10__20_), .ZN(u5_mult_82_n142) );
  XOR2_X2 u5_mult_82_U298 ( .A(u5_mult_82_n141), .B(u5_mult_82_SUMB_11__20_), 
        .Z(u5_mult_82_SUMB_12__19_) );
  XOR2_X2 u5_mult_82_U297 ( .A(u5_mult_82_ab_12__19_), .B(
        u5_mult_82_CARRYB_11__19_), .Z(u5_mult_82_n141) );
  XOR2_X2 u5_mult_82_U296 ( .A(u5_mult_82_n140), .B(u5_mult_82_SUMB_10__21_), 
        .Z(u5_mult_82_SUMB_11__20_) );
  XOR2_X2 u5_mult_82_U295 ( .A(u5_mult_82_ab_11__20_), .B(
        u5_mult_82_CARRYB_10__20_), .Z(u5_mult_82_n140) );
  INV_X2 u5_mult_82_U294 ( .A(u5_mult_82_CARRYB_28__34_), .ZN(u5_mult_82_n1664) );
  BUF_X8 u5_mult_82_U293 ( .A(u5_mult_82_SUMB_45__23_), .Z(u5_mult_82_n3772)
         );
  NAND2_X1 u5_mult_82_U292 ( .A1(u5_mult_82_ab_3__33_), .A2(
        u5_mult_82_SUMB_2__34_), .ZN(u5_mult_82_n974) );
  NAND2_X1 u5_mult_82_U291 ( .A1(u5_mult_82_ab_4__33_), .A2(
        u5_mult_82_CARRYB_3__33_), .ZN(u5_mult_82_n4503) );
  XNOR2_X1 u5_mult_82_U290 ( .A(u5_mult_82_n461), .B(u5_mult_82_SUMB_8__30_), 
        .ZN(u5_mult_82_SUMB_9__29_) );
  BUF_X4 u5_mult_82_U289 ( .A(u5_mult_82_CARRYB_16__25_), .Z(u5_mult_82_n2631)
         );
  NAND2_X2 u5_mult_82_U288 ( .A1(u5_mult_82_CARRYB_29__17_), .A2(
        u5_mult_82_SUMB_29__18_), .ZN(u5_mult_82_n4565) );
  NAND3_X4 u5_mult_82_U287 ( .A1(u5_mult_82_n3912), .A2(u5_mult_82_n3913), 
        .A3(u5_mult_82_n3914), .ZN(u5_mult_82_CARRYB_42__24_) );
  NAND2_X2 u5_mult_82_U286 ( .A1(u5_mult_82_ab_50__18_), .A2(
        u5_mult_82_CARRYB_49__18_), .ZN(u5_mult_82_n5743) );
  NAND2_X1 u5_mult_82_U285 ( .A1(u5_mult_82_ab_29__40_), .A2(
        u5_mult_82_CARRYB_28__40_), .ZN(u5_mult_82_n2450) );
  XNOR2_X2 u5_mult_82_U284 ( .A(u5_mult_82_CARRYB_41__18_), .B(
        u5_mult_82_ab_42__18_), .ZN(u5_mult_82_n139) );
  XOR2_X2 u5_mult_82_U283 ( .A(u5_mult_82_SUMB_41__19_), .B(u5_mult_82_n139), 
        .Z(u5_mult_82_n138) );
  NAND2_X2 u5_mult_82_U282 ( .A1(u5_mult_82_ab_31__13_), .A2(
        u5_mult_82_CARRYB_30__13_), .ZN(u5_mult_82_n654) );
  NAND2_X1 u5_mult_82_U281 ( .A1(u5_mult_82_CARRYB_30__13_), .A2(
        u5_mult_82_SUMB_30__14_), .ZN(u5_mult_82_n652) );
  BUF_X8 u5_mult_82_U280 ( .A(u5_mult_82_SUMB_2__51_), .Z(u5_mult_82_n422) );
  NAND2_X1 u5_mult_82_U279 ( .A1(u5_mult_82_SUMB_23__46_), .A2(
        u5_mult_82_CARRYB_23__45_), .ZN(u5_mult_82_n3374) );
  NAND2_X2 u5_mult_82_U278 ( .A1(u5_mult_82_ab_24__45_), .A2(
        u5_mult_82_SUMB_23__46_), .ZN(u5_mult_82_n3376) );
  NAND3_X2 u5_mult_82_U277 ( .A1(u5_mult_82_n4472), .A2(u5_mult_82_n4473), 
        .A3(u5_mult_82_n4474), .ZN(u5_mult_82_CARRYB_38__37_) );
  NAND3_X4 u5_mult_82_U276 ( .A1(u5_mult_82_n3774), .A2(u5_mult_82_n3775), 
        .A3(u5_mult_82_n3776), .ZN(u5_mult_82_CARRYB_32__41_) );
  NAND2_X2 u5_mult_82_U275 ( .A1(u5_mult_82_n3891), .A2(u5_mult_82_n1008), 
        .ZN(u5_mult_82_n1009) );
  NAND3_X2 u5_mult_82_U274 ( .A1(u5_mult_82_n135), .A2(u5_mult_82_n136), .A3(
        u5_mult_82_n137), .ZN(u5_mult_82_CARRYB_44__39_) );
  NAND2_X1 u5_mult_82_U273 ( .A1(u5_mult_82_ab_44__39_), .A2(
        u5_mult_82_CARRYB_43__39_), .ZN(u5_mult_82_n137) );
  NAND2_X1 u5_mult_82_U272 ( .A1(u5_mult_82_ab_44__39_), .A2(
        u5_mult_82_SUMB_43__40_), .ZN(u5_mult_82_n136) );
  NAND2_X1 u5_mult_82_U271 ( .A1(u5_mult_82_CARRYB_43__39_), .A2(
        u5_mult_82_SUMB_43__40_), .ZN(u5_mult_82_n135) );
  XOR2_X2 u5_mult_82_U270 ( .A(u5_mult_82_SUMB_43__40_), .B(u5_mult_82_n134), 
        .Z(u5_mult_82_SUMB_44__39_) );
  XOR2_X2 u5_mult_82_U269 ( .A(u5_mult_82_CARRYB_43__39_), .B(
        u5_mult_82_ab_44__39_), .Z(u5_mult_82_n134) );
  NAND3_X2 u5_mult_82_U268 ( .A1(u5_mult_82_n131), .A2(u5_mult_82_n132), .A3(
        u5_mult_82_n133), .ZN(u5_mult_82_CARRYB_31__45_) );
  NAND2_X1 u5_mult_82_U267 ( .A1(u5_mult_82_ab_31__45_), .A2(
        u5_mult_82_SUMB_30__46_), .ZN(u5_mult_82_n133) );
  NAND2_X2 u5_mult_82_U266 ( .A1(u5_mult_82_ab_31__45_), .A2(
        u5_mult_82_CARRYB_30__45_), .ZN(u5_mult_82_n132) );
  NAND2_X1 u5_mult_82_U265 ( .A1(u5_mult_82_SUMB_30__46_), .A2(
        u5_mult_82_CARRYB_30__45_), .ZN(u5_mult_82_n131) );
  XOR2_X2 u5_mult_82_U264 ( .A(u5_mult_82_CARRYB_30__45_), .B(u5_mult_82_n130), 
        .Z(u5_mult_82_SUMB_31__45_) );
  XOR2_X2 u5_mult_82_U263 ( .A(u5_mult_82_SUMB_30__46_), .B(
        u5_mult_82_ab_31__45_), .Z(u5_mult_82_n130) );
  NAND3_X2 u5_mult_82_U262 ( .A1(u5_mult_82_n127), .A2(u5_mult_82_n128), .A3(
        u5_mult_82_n129), .ZN(u5_mult_82_CARRYB_52__35_) );
  NAND2_X1 u5_mult_82_U261 ( .A1(u5_mult_82_ab_52__35_), .A2(
        u5_mult_82_SUMB_51__36_), .ZN(u5_mult_82_n129) );
  NAND2_X2 u5_mult_82_U260 ( .A1(u5_mult_82_ab_52__35_), .A2(
        u5_mult_82_CARRYB_51__35_), .ZN(u5_mult_82_n128) );
  NAND2_X1 u5_mult_82_U259 ( .A1(u5_mult_82_SUMB_51__36_), .A2(
        u5_mult_82_CARRYB_51__35_), .ZN(u5_mult_82_n127) );
  XOR2_X2 u5_mult_82_U258 ( .A(u5_mult_82_CARRYB_51__35_), .B(u5_mult_82_n126), 
        .Z(u5_mult_82_SUMB_52__35_) );
  XOR2_X2 u5_mult_82_U257 ( .A(u5_mult_82_SUMB_51__36_), .B(
        u5_mult_82_ab_52__35_), .Z(u5_mult_82_n126) );
  NAND3_X4 u5_mult_82_U256 ( .A1(u5_mult_82_n123), .A2(u5_mult_82_n124), .A3(
        u5_mult_82_n125), .ZN(u5_mult_82_CARRYB_23__46_) );
  NAND2_X2 u5_mult_82_U255 ( .A1(u5_mult_82_ab_23__46_), .A2(
        u5_mult_82_SUMB_22__47_), .ZN(u5_mult_82_n125) );
  NAND2_X2 u5_mult_82_U254 ( .A1(u5_mult_82_CARRYB_22__46_), .A2(
        u5_mult_82_SUMB_22__47_), .ZN(u5_mult_82_n124) );
  NAND2_X1 u5_mult_82_U253 ( .A1(u5_mult_82_CARRYB_22__46_), .A2(
        u5_mult_82_ab_23__46_), .ZN(u5_mult_82_n123) );
  NAND3_X4 u5_mult_82_U252 ( .A1(u5_mult_82_n120), .A2(u5_mult_82_n121), .A3(
        u5_mult_82_n122), .ZN(u5_mult_82_CARRYB_22__47_) );
  NAND2_X1 u5_mult_82_U251 ( .A1(u5_mult_82_CARRYB_21__47_), .A2(
        u5_mult_82_SUMB_21__48_), .ZN(u5_mult_82_n122) );
  NAND2_X1 u5_mult_82_U250 ( .A1(u5_mult_82_ab_22__47_), .A2(
        u5_mult_82_SUMB_21__48_), .ZN(u5_mult_82_n121) );
  NAND2_X1 u5_mult_82_U249 ( .A1(u5_mult_82_ab_22__47_), .A2(
        u5_mult_82_CARRYB_21__47_), .ZN(u5_mult_82_n120) );
  XOR2_X2 u5_mult_82_U248 ( .A(u5_mult_82_n119), .B(u5_mult_82_SUMB_22__47_), 
        .Z(u5_mult_82_SUMB_23__46_) );
  XOR2_X2 u5_mult_82_U247 ( .A(u5_mult_82_CARRYB_22__46_), .B(
        u5_mult_82_ab_23__46_), .Z(u5_mult_82_n119) );
  XOR2_X2 u5_mult_82_U246 ( .A(u5_mult_82_n118), .B(u5_mult_82_SUMB_21__48_), 
        .Z(u5_mult_82_SUMB_22__47_) );
  XOR2_X2 u5_mult_82_U245 ( .A(u5_mult_82_ab_22__47_), .B(
        u5_mult_82_CARRYB_21__47_), .Z(u5_mult_82_n118) );
  XOR2_X2 u5_mult_82_U244 ( .A(u5_mult_82_ab_19__20_), .B(
        u5_mult_82_CARRYB_18__20_), .Z(u5_mult_82_n2794) );
  NAND2_X2 u5_mult_82_U243 ( .A1(u5_mult_82_CARRYB_23__17_), .A2(
        u5_mult_82_SUMB_23__18_), .ZN(u5_mult_82_n5304) );
  NAND3_X4 u5_mult_82_U242 ( .A1(u5_mult_82_n5302), .A2(u5_mult_82_n5303), 
        .A3(u5_mult_82_n5304), .ZN(u5_mult_82_CARRYB_24__17_) );
  NAND2_X2 u5_mult_82_U241 ( .A1(u5_mult_82_ab_28__15_), .A2(
        u5_mult_82_SUMB_27__16_), .ZN(u5_mult_82_n4900) );
  NAND2_X4 u5_mult_82_U240 ( .A1(u5_mult_82_SUMB_27__34_), .A2(
        u5_mult_82_n1614), .ZN(u5_mult_82_n2426) );
  NAND2_X4 u5_mult_82_U239 ( .A1(u5_mult_82_n3541), .A2(u5_mult_82_n3542), 
        .ZN(u5_mult_82_SUMB_50__11_) );
  NAND2_X2 u5_mult_82_U238 ( .A1(u5_mult_82_CARRYB_39__24_), .A2(
        u5_mult_82_SUMB_39__25_), .ZN(u5_mult_82_n3859) );
  INV_X16 u5_mult_82_U237 ( .A(u5_mult_82_n6814), .ZN(u5_mult_82_n6811) );
  INV_X16 u5_mult_82_U236 ( .A(u5_mult_82_n6814), .ZN(u5_mult_82_n6810) );
  INV_X16 u5_mult_82_U235 ( .A(u5_mult_82_n6814), .ZN(u5_mult_82_n6813) );
  NAND2_X4 u5_mult_82_U234 ( .A1(u5_mult_82_ab_29__21_), .A2(u5_mult_82_n3074), 
        .ZN(u5_mult_82_n5437) );
  NAND2_X2 u5_mult_82_U233 ( .A1(u5_mult_82_CARRYB_20__24_), .A2(
        u5_mult_82_SUMB_20__25_), .ZN(u5_mult_82_net80542) );
  NAND2_X2 u5_mult_82_U232 ( .A1(u5_mult_82_ab_15__37_), .A2(
        u5_mult_82_SUMB_14__38_), .ZN(u5_mult_82_n963) );
  NAND2_X2 u5_mult_82_U231 ( .A1(u5_mult_82_ab_5__45_), .A2(
        u5_mult_82_SUMB_4__46_), .ZN(u5_mult_82_n4994) );
  NOR2_X2 u5_mult_82_U230 ( .A1(u5_mult_82_n6849), .A2(u5_mult_82_net66107), 
        .ZN(u5_mult_82_ab_1__31_) );
  XNOR2_X2 u5_mult_82_U229 ( .A(u5_mult_82_SUMB_35__38_), .B(
        u5_mult_82_ab_36__37_), .ZN(u5_mult_82_n117) );
  XNOR2_X2 u5_mult_82_U228 ( .A(u5_mult_82_CARRYB_35__37_), .B(u5_mult_82_n117), .ZN(u5_mult_82_SUMB_36__37_) );
  XNOR2_X2 u5_mult_82_U227 ( .A(u5_mult_82_CARRYB_47__28_), .B(
        u5_mult_82_ab_48__28_), .ZN(u5_mult_82_n116) );
  XNOR2_X2 u5_mult_82_U226 ( .A(u5_mult_82_SUMB_47__29_), .B(u5_mult_82_n116), 
        .ZN(u5_mult_82_SUMB_48__28_) );
  NAND2_X4 u5_mult_82_U225 ( .A1(u5_mult_82_n258), .A2(u5_mult_82_n259), .ZN(
        u5_mult_82_n261) );
  INV_X32 u5_mult_82_U224 ( .A(u5_mult_82_net66121), .ZN(u5_mult_82_n1262) );
  NAND2_X2 u5_mult_82_U223 ( .A1(u5_mult_82_CARRYB_21__25_), .A2(
        u5_mult_82_SUMB_21__26_), .ZN(u5_mult_82_n2194) );
  BUF_X8 u5_mult_82_U222 ( .A(u5_mult_82_CARRYB_9__27_), .Z(u5_mult_82_n1390)
         );
  NAND2_X2 u5_mult_82_U221 ( .A1(u5_mult_82_ab_24__17_), .A2(
        u5_mult_82_SUMB_23__18_), .ZN(u5_mult_82_n5303) );
  NAND2_X2 u5_mult_82_U220 ( .A1(u5_mult_82_ab_46__31_), .A2(u5_mult_82_n1566), 
        .ZN(u5_mult_82_n3833) );
  NAND2_X2 u5_mult_82_U219 ( .A1(u5_mult_82_n1566), .A2(
        u5_mult_82_SUMB_45__32_), .ZN(u5_mult_82_n3835) );
  XNOR2_X2 u5_mult_82_U218 ( .A(u5_mult_82_CARRYB_52__35_), .B(
        u5_mult_82_SUMB_52__36_), .ZN(u5_mult_82_n6423) );
  NAND2_X2 u5_mult_82_U217 ( .A1(u5_mult_82_ab_11__29_), .A2(
        u5_mult_82_SUMB_10__30_), .ZN(u5_mult_82_n2306) );
  NAND3_X4 u5_mult_82_U216 ( .A1(u5_mult_82_n2305), .A2(u5_mult_82_n2306), 
        .A3(u5_mult_82_n2307), .ZN(u5_mult_82_CARRYB_11__29_) );
  NOR2_X1 u5_mult_82_U215 ( .A1(u5_mult_82_n6861), .A2(u5_mult_82_n6753), .ZN(
        u5_mult_82_ab_49__29_) );
  INV_X8 u5_mult_82_U214 ( .A(u5_mult_82_CARRYB_48__29_), .ZN(u5_mult_82_n113)
         );
  INV_X4 u5_mult_82_U213 ( .A(u5_mult_82_ab_49__29_), .ZN(u5_mult_82_n112) );
  NAND2_X4 u5_mult_82_U212 ( .A1(u5_mult_82_n114), .A2(u5_mult_82_n115), .ZN(
        u5_mult_82_n2326) );
  NAND2_X4 u5_mult_82_U211 ( .A1(u5_mult_82_n112), .A2(u5_mult_82_n113), .ZN(
        u5_mult_82_n115) );
  NAND2_X2 u5_mult_82_U210 ( .A1(u5_mult_82_ab_49__29_), .A2(
        u5_mult_82_CARRYB_48__29_), .ZN(u5_mult_82_n114) );
  NAND2_X4 u5_mult_82_U209 ( .A1(u5_mult_82_n5561), .A2(u5_mult_82_n5562), 
        .ZN(u5_mult_82_n5564) );
  XNOR2_X2 u5_mult_82_U208 ( .A(u5_mult_82_ab_14__17_), .B(
        u5_mult_82_CARRYB_13__17_), .ZN(u5_mult_82_n111) );
  XNOR2_X2 u5_mult_82_U207 ( .A(u5_mult_82_n111), .B(u5_mult_82_SUMB_13__18_), 
        .ZN(u5_mult_82_SUMB_14__17_) );
  NOR2_X2 u5_mult_82_U206 ( .A1(u5_mult_82_n6842), .A2(u5_mult_82_n1262), .ZN(
        u5_mult_82_ab_1__32_) );
  INV_X1 u5_mult_82_U205 ( .A(u5_mult_82_ab_0__33_), .ZN(u5_mult_82_n108) );
  INV_X2 u5_mult_82_U204 ( .A(u5_mult_82_ab_1__32_), .ZN(u5_mult_82_n107) );
  NAND2_X2 u5_mult_82_U203 ( .A1(u5_mult_82_n109), .A2(u5_mult_82_n110), .ZN(
        u5_mult_82_n468) );
  NAND2_X2 u5_mult_82_U202 ( .A1(u5_mult_82_n107), .A2(u5_mult_82_ab_0__33_), 
        .ZN(u5_mult_82_n110) );
  NAND2_X2 u5_mult_82_U201 ( .A1(u5_mult_82_ab_1__32_), .A2(u5_mult_82_n108), 
        .ZN(u5_mult_82_n109) );
  INV_X32 u5_mult_82_U200 ( .A(u5_mult_82_ab_29__18_), .ZN(u5_mult_82_n106) );
  XNOR2_X2 u5_mult_82_U199 ( .A(u5_mult_82_CARRYB_28__18_), .B(u5_mult_82_n106), .ZN(u5_mult_82_n4558) );
  NAND2_X2 u5_mult_82_U198 ( .A1(u5_mult_82_CARRYB_40__19_), .A2(
        u5_mult_82_SUMB_40__20_), .ZN(u5_mult_82_n1134) );
  XNOR2_X2 u5_mult_82_U197 ( .A(u5_mult_82_ab_36__32_), .B(
        u5_mult_82_CARRYB_35__32_), .ZN(u5_mult_82_n105) );
  XNOR2_X2 u5_mult_82_U196 ( .A(u5_mult_82_n105), .B(u5_mult_82_SUMB_35__33_), 
        .ZN(u5_mult_82_SUMB_36__32_) );
  NAND2_X2 u5_mult_82_U195 ( .A1(u5_mult_82_ab_46__3_), .A2(
        u5_mult_82_CARRYB_45__3_), .ZN(u5_mult_82_n4512) );
  INV_X4 u5_mult_82_U194 ( .A(u5_mult_82_n103), .ZN(u5_mult_82_n104) );
  INV_X2 u5_mult_82_U193 ( .A(u5_mult_82_CARRYB_6__24_), .ZN(u5_mult_82_n103)
         );
  INV_X1 u5_mult_82_U192 ( .A(u5_mult_82_SUMB_24__20_), .ZN(u5_mult_82_n100)
         );
  INV_X4 u5_mult_82_U191 ( .A(u5_mult_82_n930), .ZN(u5_mult_82_n99) );
  NAND2_X2 u5_mult_82_U190 ( .A1(u5_mult_82_n101), .A2(u5_mult_82_n102), .ZN(
        u5_mult_82_SUMB_25__19_) );
  NAND2_X2 u5_mult_82_U189 ( .A1(u5_mult_82_n99), .A2(u5_mult_82_n100), .ZN(
        u5_mult_82_n102) );
  NAND2_X1 u5_mult_82_U188 ( .A1(u5_mult_82_n930), .A2(u5_mult_82_SUMB_24__20_), .ZN(u5_mult_82_n101) );
  NOR2_X2 u5_mult_82_U187 ( .A1(u5_mult_82_net64379), .A2(u5_mult_82_net65283), 
        .ZN(u5_mult_82_ab_47__6_) );
  INV_X4 u5_mult_82_U186 ( .A(u5_mult_82_ab_0__40_), .ZN(u5_mult_82_n96) );
  INV_X4 u5_mult_82_U185 ( .A(u5_mult_82_n2311), .ZN(u5_mult_82_n95) );
  NAND2_X2 u5_mult_82_U184 ( .A1(u5_mult_82_n97), .A2(u5_mult_82_n98), .ZN(
        u5_mult_82_n2310) );
  NAND2_X2 u5_mult_82_U183 ( .A1(u5_mult_82_n95), .A2(u5_mult_82_n96), .ZN(
        u5_mult_82_n98) );
  NAND2_X2 u5_mult_82_U182 ( .A1(u5_mult_82_n2311), .A2(u5_mult_82_ab_0__40_), 
        .ZN(u5_mult_82_n97) );
  INV_X1 u5_mult_82_U181 ( .A(u5_mult_82_ab_47__6_), .ZN(u5_mult_82_n92) );
  INV_X4 u5_mult_82_U180 ( .A(u5_mult_82_CARRYB_46__6_), .ZN(u5_mult_82_n91)
         );
  NAND2_X2 u5_mult_82_U179 ( .A1(u5_mult_82_n93), .A2(u5_mult_82_n94), .ZN(
        u5_mult_82_n4146) );
  NAND2_X2 u5_mult_82_U178 ( .A1(u5_mult_82_n91), .A2(u5_mult_82_n92), .ZN(
        u5_mult_82_n94) );
  NAND2_X1 u5_mult_82_U177 ( .A1(u5_mult_82_CARRYB_46__6_), .A2(
        u5_mult_82_ab_47__6_), .ZN(u5_mult_82_n93) );
  NAND2_X4 u5_mult_82_U176 ( .A1(u5_mult_82_ab_15__36_), .A2(u5_mult_82_n1859), 
        .ZN(u5_mult_82_n5022) );
  NAND2_X4 u5_mult_82_U175 ( .A1(u5_mult_82_ab_29__39_), .A2(u5_mult_82_n1810), 
        .ZN(u5_mult_82_n2400) );
  NAND2_X2 u5_mult_82_U174 ( .A1(u5_mult_82_ab_36__24_), .A2(
        u5_mult_82_CARRYB_35__24_), .ZN(u5_mult_82_n5032) );
  INV_X4 u5_mult_82_U173 ( .A(u5_mult_82_n1615), .ZN(u5_mult_82_n1616) );
  INV_X1 u5_mult_82_U172 ( .A(u5_mult_82_ab_36__34_), .ZN(u5_mult_82_n1906) );
  INV_X4 u5_mult_82_U171 ( .A(u5_mult_82_CARRYB_35__34_), .ZN(u5_mult_82_n88)
         );
  INV_X4 u5_mult_82_U170 ( .A(u5_mult_82_n1906), .ZN(u5_mult_82_n87) );
  NAND2_X4 u5_mult_82_U169 ( .A1(u5_mult_82_n89), .A2(u5_mult_82_n90), .ZN(
        u5_mult_82_n3924) );
  NAND2_X4 u5_mult_82_U168 ( .A1(u5_mult_82_n87), .A2(u5_mult_82_n88), .ZN(
        u5_mult_82_n90) );
  NAND2_X2 u5_mult_82_U167 ( .A1(u5_mult_82_n1906), .A2(
        u5_mult_82_CARRYB_35__34_), .ZN(u5_mult_82_n89) );
  BUF_X4 u5_mult_82_U166 ( .A(u5_mult_82_CARRYB_23__13_), .Z(u5_mult_82_n1596)
         );
  NOR2_X2 u5_mult_82_U165 ( .A1(u5_mult_82_n6820), .A2(u5_mult_82_net66107), 
        .ZN(u5_mult_82_ab_1__41_) );
  NAND2_X2 u5_mult_82_U164 ( .A1(u5_mult_82_ab_44__16_), .A2(
        u5_mult_82_CARRYB_43__16_), .ZN(u5_mult_82_n4286) );
  INV_X2 u5_mult_82_U163 ( .A(u5_mult_82_SUMB_16__36_), .ZN(u5_mult_82_n2358)
         );
  OR2_X2 u5_mult_82_U162 ( .A1(u5_mult_82_n6186), .A2(u5_mult_82_n2358), .ZN(
        u5_mult_82_n2360) );
  CLKBUF_X2 u5_mult_82_U161 ( .A(u5_mult_82_SUMB_31__21_), .Z(u5_mult_82_n86)
         );
  XOR2_X1 u5_mult_82_U160 ( .A(u5_mult_82_CARRYB_8__51_), .B(
        u5_mult_82_ab_9__51_), .Z(u5_mult_82_n2083) );
  INV_X8 u5_mult_82_U159 ( .A(u5_mult_82_n84), .ZN(u5_mult_82_n85) );
  INV_X4 u5_mult_82_U158 ( .A(u5_mult_82_SUMB_24__19_), .ZN(u5_mult_82_n84) );
  XNOR2_X2 u5_mult_82_U157 ( .A(u5_mult_82_ab_45__15_), .B(
        u5_mult_82_CARRYB_44__15_), .ZN(u5_mult_82_n83) );
  XNOR2_X2 u5_mult_82_U156 ( .A(u5_mult_82_n83), .B(u5_mult_82_SUMB_44__16_), 
        .ZN(u5_mult_82_SUMB_45__15_) );
  INV_X4 u5_mult_82_U155 ( .A(u5_mult_82_n81), .ZN(u5_mult_82_n82) );
  INV_X2 u5_mult_82_U154 ( .A(u5_mult_82_SUMB_34__24_), .ZN(u5_mult_82_n81) );
  XNOR2_X2 u5_mult_82_U153 ( .A(u5_mult_82_ab_29__33_), .B(
        u5_mult_82_CARRYB_28__33_), .ZN(u5_mult_82_n80) );
  INV_X4 u5_mult_82_U152 ( .A(u5_mult_82_n79), .ZN(u5_mult_82_SUMB_29__33_) );
  XNOR2_X2 u5_mult_82_U151 ( .A(u5_mult_82_n80), .B(u5_mult_82_n1549), .ZN(
        u5_mult_82_n79) );
  NAND2_X2 u5_mult_82_U150 ( .A1(u5_mult_82_ab_1__30_), .A2(
        u5_mult_82_ab_0__31_), .ZN(u5_mult_82_n6484) );
  NAND2_X2 u5_mult_82_U149 ( .A1(u5_mult_82_ab_0__44_), .A2(
        u5_mult_82_ab_1__43_), .ZN(u5_mult_82_n6497) );
  NAND2_X2 u5_mult_82_U148 ( .A1(u5_mult_82_ab_1__46_), .A2(
        u5_mult_82_ab_0__47_), .ZN(u5_mult_82_n6502) );
  NAND2_X1 u5_mult_82_U147 ( .A1(u5_mult_82_ab_0__40_), .A2(
        u5_mult_82_net66121), .ZN(u5_mult_82_n2133) );
  NOR2_X2 u5_mult_82_U146 ( .A1(u5_mult_82_net64217), .A2(u5_mult_82_n6849), 
        .ZN(u5_mult_82_ab_0__31_) );
  NOR2_X2 u5_mult_82_U145 ( .A1(u5_mult_82_net64217), .A2(u5_mult_82_n6815), 
        .ZN(u5_mult_82_ab_0__42_) );
  NOR2_X2 u5_mult_82_U144 ( .A1(u5_mult_82_net64217), .A2(u5_mult_82_n7008), 
        .ZN(u5_mult_82_ab_0__45_) );
  NOR2_X2 u5_mult_82_U143 ( .A1(u5_mult_82_net64217), .A2(u5_mult_82_n1263), 
        .ZN(u5_mult_82_ab_0__36_) );
  NOR2_X2 u5_mult_82_U142 ( .A1(u5_mult_82_net64217), .A2(u5_mult_82_n6783), 
        .ZN(u5_mult_82_ab_0__47_) );
  BUF_X8 u5_mult_82_U141 ( .A(u5_mult_82_SUMB_24__15_), .Z(u5_mult_82_n1795)
         );
  XOR2_X2 u5_mult_82_U140 ( .A(u5_mult_82_n4828), .B(u5_mult_82_n1795), .Z(
        u5_mult_82_n78) );
  XNOR2_X2 u5_mult_82_U139 ( .A(u5_mult_82_ab_18__28_), .B(
        u5_mult_82_CARRYB_17__28_), .ZN(u5_mult_82_n77) );
  XNOR2_X2 u5_mult_82_U138 ( .A(u5_mult_82_n77), .B(u5_mult_82_n31), .ZN(
        u5_mult_82_SUMB_18__28_) );
  INV_X4 u5_mult_82_U137 ( .A(u5_mult_82_n75), .ZN(u5_mult_82_n76) );
  INV_X2 u5_mult_82_U136 ( .A(u5_mult_82_SUMB_16__39_), .ZN(u5_mult_82_n75) );
  XNOR2_X2 u5_mult_82_U135 ( .A(u5_mult_82_CARRYB_15__37_), .B(
        u5_mult_82_ab_16__37_), .ZN(u5_mult_82_n1756) );
  XNOR2_X2 u5_mult_82_U134 ( .A(u5_mult_82_SUMB_16__24_), .B(u5_mult_82_n2847), 
        .ZN(u5_mult_82_SUMB_17__23_) );
  XNOR2_X1 u5_mult_82_U133 ( .A(u5_mult_82_CARRYB_22__11_), .B(
        u5_mult_82_ab_23__11_), .ZN(u5_mult_82_n2074) );
  NAND3_X2 u5_mult_82_U132 ( .A1(u5_mult_82_n4983), .A2(u5_mult_82_n4984), 
        .A3(u5_mult_82_n4985), .ZN(u5_mult_82_CARRYB_41__18_) );
  INV_X4 u5_mult_82_U131 ( .A(u5_mult_82_n73), .ZN(u5_mult_82_n74) );
  INV_X4 u5_mult_82_U130 ( .A(u5_mult_82_n71), .ZN(u5_mult_82_n72) );
  INV_X2 u5_mult_82_U129 ( .A(u5_mult_82_SUMB_32__33_), .ZN(u5_mult_82_n71) );
  XNOR2_X2 u5_mult_82_U128 ( .A(u5_mult_82_n1578), .B(u5_mult_82_SUMB_22__27_), 
        .ZN(u5_mult_82_n70) );
  XNOR2_X2 u5_mult_82_U127 ( .A(u5_mult_82_ab_18__39_), .B(
        u5_mult_82_CARRYB_17__39_), .ZN(u5_mult_82_n69) );
  XNOR2_X2 u5_mult_82_U126 ( .A(u5_mult_82_n69), .B(u5_mult_82_SUMB_17__40_), 
        .ZN(u5_mult_82_SUMB_18__39_) );
  NOR2_X2 u5_mult_82_U125 ( .A1(u5_mult_82_n6772), .A2(u5_mult_82_net66107), 
        .ZN(u5_mult_82_ab_1__49_) );
  NOR2_X1 u5_mult_82_U124 ( .A1(u5_mult_82_n6810), .A2(u5_mult_82_net66107), 
        .ZN(u5_mult_82_ab_1__43_) );
  NAND2_X1 u5_mult_82_U123 ( .A1(u5_mult_82_CARRYB_12__48_), .A2(
        u5_mult_82_SUMB_12__49_), .ZN(u5_mult_82_n909) );
  NAND2_X1 u5_mult_82_U122 ( .A1(u5_mult_82_ab_13__48_), .A2(
        u5_mult_82_CARRYB_12__48_), .ZN(u5_mult_82_n907) );
  XNOR2_X2 u5_mult_82_U121 ( .A(u5_mult_82_SUMB_2__44_), .B(u5_mult_82_n1712), 
        .ZN(u5_mult_82_SUMB_3__43_) );
  NOR2_X4 u5_mult_82_U120 ( .A1(u5_mult_82_net66107), .A2(u5_mult_82_n7008), 
        .ZN(u5_mult_82_n68) );
  XNOR2_X2 u5_mult_82_U119 ( .A(u5_mult_82_ab_29__23_), .B(
        u5_mult_82_CARRYB_28__23_), .ZN(u5_mult_82_n67) );
  XNOR2_X2 u5_mult_82_U118 ( .A(u5_mult_82_n67), .B(u5_mult_82_n1522), .ZN(
        u5_mult_82_SUMB_29__23_) );
  XOR2_X2 u5_mult_82_U117 ( .A(u5_mult_82_CARRYB_31__38_), .B(
        u5_mult_82_ab_32__38_), .Z(u5_mult_82_n4924) );
  INV_X4 u5_mult_82_U116 ( .A(u5_mult_82_n65), .ZN(u5_mult_82_n66) );
  INV_X2 u5_mult_82_U115 ( .A(u5_mult_82_SUMB_19__41_), .ZN(u5_mult_82_n65) );
  CLKBUF_X2 u5_mult_82_U114 ( .A(u5_mult_82_CARRYB_3__49_), .Z(
        u5_mult_82_n1468) );
  NOR2_X4 u5_mult_82_U113 ( .A1(u5_mult_82_net64217), .A2(u5_mult_82_n7007), 
        .ZN(u5_mult_82_n64) );
  XNOR2_X1 u5_mult_82_U112 ( .A(u5_mult_82_CARRYB_22__22_), .B(
        u5_mult_82_ab_23__22_), .ZN(u5_mult_82_n63) );
  XNOR2_X2 u5_mult_82_U111 ( .A(u5_mult_82_n1101), .B(u5_mult_82_n63), .ZN(
        u5_mult_82_SUMB_23__22_) );
  XNOR2_X2 u5_mult_82_U110 ( .A(u5_mult_82_ab_21__35_), .B(
        u5_mult_82_CARRYB_20__35_), .ZN(u5_mult_82_n62) );
  XNOR2_X2 u5_mult_82_U109 ( .A(u5_mult_82_n62), .B(u5_mult_82_SUMB_20__36_), 
        .ZN(u5_mult_82_SUMB_21__35_) );
  XNOR2_X2 u5_mult_82_U108 ( .A(u5_mult_82_ab_22__27_), .B(
        u5_mult_82_CARRYB_21__27_), .ZN(u5_mult_82_n61) );
  XNOR2_X2 u5_mult_82_U107 ( .A(u5_mult_82_n61), .B(u5_mult_82_SUMB_21__28_), 
        .ZN(u5_mult_82_SUMB_22__27_) );
  NAND3_X2 u5_mult_82_U106 ( .A1(u5_mult_82_n4385), .A2(u5_mult_82_n4386), 
        .A3(u5_mult_82_n4387), .ZN(u5_mult_82_CARRYB_42__8_) );
  XOR2_X2 u5_mult_82_U105 ( .A(u5_mult_82_ab_23__21_), .B(
        u5_mult_82_CARRYB_22__21_), .Z(u5_mult_82_n3162) );
  CLKBUF_X3 u5_mult_82_U104 ( .A(u5_mult_82_SUMB_25__27_), .Z(u5_mult_82_n60)
         );
  XNOR2_X2 u5_mult_82_U103 ( .A(u5_mult_82_ab_9__36_), .B(
        u5_mult_82_CARRYB_8__36_), .ZN(u5_mult_82_n59) );
  XNOR2_X2 u5_mult_82_U102 ( .A(u5_mult_82_n59), .B(u5_mult_82_n1763), .ZN(
        u5_mult_82_SUMB_9__36_) );
  INV_X8 u5_mult_82_U101 ( .A(u5_mult_82_n57), .ZN(u5_mult_82_n58) );
  INV_X4 u5_mult_82_U100 ( .A(u5_mult_82_CARRYB_31__27_), .ZN(u5_mult_82_n57)
         );
  NAND2_X1 u5_mult_82_U99 ( .A1(u5_mult_82_CARRYB_13__25_), .A2(
        u5_mult_82_SUMB_13__26_), .ZN(u5_mult_82_n5151) );
  XNOR2_X2 u5_mult_82_U98 ( .A(u5_mult_82_ab_18__38_), .B(
        u5_mult_82_CARRYB_17__38_), .ZN(u5_mult_82_n56) );
  XNOR2_X2 u5_mult_82_U97 ( .A(u5_mult_82_n56), .B(u5_mult_82_n1512), .ZN(
        u5_mult_82_SUMB_18__38_) );
  CLKBUF_X3 u5_mult_82_U96 ( .A(u5_mult_82_SUMB_37__8_), .Z(u5_mult_82_n55) );
  INV_X8 u5_mult_82_U95 ( .A(u5_mult_82_n53), .ZN(u5_mult_82_n54) );
  INV_X4 u5_mult_82_U94 ( .A(u5_mult_82_SUMB_24__30_), .ZN(u5_mult_82_n53) );
  XNOR2_X2 u5_mult_82_U93 ( .A(u5_mult_82_ab_38__35_), .B(
        u5_mult_82_CARRYB_37__35_), .ZN(u5_mult_82_n52) );
  XNOR2_X2 u5_mult_82_U92 ( .A(u5_mult_82_n52), .B(u5_mult_82_SUMB_37__36_), 
        .ZN(u5_mult_82_SUMB_38__35_) );
  CLKBUF_X2 u5_mult_82_U91 ( .A(u5_mult_82_SUMB_23__5_), .Z(u5_mult_82_n51) );
  XNOR2_X2 u5_mult_82_U90 ( .A(u5_mult_82_SUMB_31__29_), .B(u5_mult_82_n1443), 
        .ZN(u5_mult_82_SUMB_32__28_) );
  XNOR2_X2 u5_mult_82_U89 ( .A(u5_mult_82_CARRYB_48__26_), .B(
        u5_mult_82_ab_49__26_), .ZN(u5_mult_82_n50) );
  XNOR2_X2 u5_mult_82_U88 ( .A(u5_mult_82_n50), .B(u5_mult_82_SUMB_48__27_), 
        .ZN(u5_mult_82_SUMB_49__26_) );
  NAND2_X1 u5_mult_82_U87 ( .A1(u5_mult_82_CARRYB_19__26_), .A2(
        u5_mult_82_SUMB_19__27_), .ZN(u5_mult_82_net85541) );
  INV_X8 u5_mult_82_U86 ( .A(u5_mult_82_n48), .ZN(u5_mult_82_n49) );
  INV_X4 u5_mult_82_U85 ( .A(u5_mult_82_SUMB_41__2_), .ZN(u5_mult_82_n48) );
  XNOR2_X2 u5_mult_82_U84 ( .A(u5_mult_82_n2733), .B(u5_mult_82_SUMB_5__38_), 
        .ZN(u5_mult_82_SUMB_6__37_) );
  NAND2_X1 u5_mult_82_U83 ( .A1(u5_mult_82_CARRYB_6__36_), .A2(
        u5_mult_82_SUMB_6__37_), .ZN(u5_mult_82_n891) );
  NAND2_X1 u5_mult_82_U82 ( .A1(u5_mult_82_ab_7__36_), .A2(
        u5_mult_82_SUMB_6__37_), .ZN(u5_mult_82_n890) );
  CLKBUF_X2 u5_mult_82_U81 ( .A(u5_mult_82_SUMB_41__8_), .Z(u5_mult_82_n47) );
  XNOR2_X2 u5_mult_82_U80 ( .A(u5_mult_82_CARRYB_11__26_), .B(
        u5_mult_82_ab_12__26_), .ZN(u5_mult_82_n46) );
  XNOR2_X2 u5_mult_82_U79 ( .A(u5_mult_82_n46), .B(u5_mult_82_SUMB_11__27_), 
        .ZN(u5_mult_82_SUMB_12__26_) );
  CLKBUF_X3 u5_mult_82_U78 ( .A(u5_mult_82_SUMB_47__26_), .Z(u5_mult_82_n727)
         );
  XNOR2_X1 u5_mult_82_U77 ( .A(u5_mult_82_n1520), .B(u5_mult_82_n727), .ZN(
        u5_mult_82_n45) );
  INV_X32 u5_mult_82_U76 ( .A(u5_mult_82_ab_46__25_), .ZN(u5_mult_82_n44) );
  XNOR2_X2 u5_mult_82_U75 ( .A(u5_mult_82_n44), .B(u5_mult_82_CARRYB_45__25_), 
        .ZN(u5_mult_82_n1144) );
  NAND3_X2 u5_mult_82_U74 ( .A1(u5_mult_82_n3929), .A2(u5_mult_82_n3928), .A3(
        u5_mult_82_n3930), .ZN(u5_mult_82_CARRYB_36__34_) );
  NAND2_X1 u5_mult_82_U73 ( .A1(u5_mult_82_CARRYB_37__7_), .A2(
        u5_mult_82_SUMB_37__8_), .ZN(u5_mult_82_n3963) );
  XNOR2_X2 u5_mult_82_U72 ( .A(u5_mult_82_ab_28__11_), .B(
        u5_mult_82_CARRYB_27__11_), .ZN(u5_mult_82_n43) );
  XNOR2_X2 u5_mult_82_U71 ( .A(u5_mult_82_n43), .B(u5_mult_82_SUMB_27__12_), 
        .ZN(u5_mult_82_SUMB_28__11_) );
  INV_X4 u5_mult_82_U70 ( .A(u5_mult_82_SUMB_33__33_), .ZN(u5_mult_82_n73) );
  XNOR2_X2 u5_mult_82_U69 ( .A(u5_mult_82_n2716), .B(u5_mult_82_n73), .ZN(
        u5_mult_82_SUMB_34__32_) );
  INV_X4 u5_mult_82_U68 ( .A(u5_mult_82_n41), .ZN(u5_mult_82_n42) );
  INV_X2 u5_mult_82_U67 ( .A(u5_mult_82_CARRYB_44__34_), .ZN(u5_mult_82_n41)
         );
  XNOR2_X1 u5_mult_82_U66 ( .A(u5_mult_82_CARRYB_2__50_), .B(
        u5_mult_82_ab_3__50_), .ZN(u5_mult_82_n40) );
  XNOR2_X2 u5_mult_82_U65 ( .A(u5_mult_82_n40), .B(u5_mult_82_n422), .ZN(
        u5_mult_82_SUMB_3__50_) );
  BUF_X8 u5_mult_82_U64 ( .A(u5_mult_82_SUMB_27__30_), .Z(u5_mult_82_n1809) );
  CLKBUF_X2 u5_mult_82_U63 ( .A(u5_mult_82_SUMB_38__8_), .Z(u5_mult_82_n39) );
  XNOR2_X2 u5_mult_82_U62 ( .A(u5_mult_82_ab_19__23_), .B(
        u5_mult_82_CARRYB_18__23_), .ZN(u5_mult_82_n38) );
  XNOR2_X2 u5_mult_82_U61 ( .A(u5_mult_82_n38), .B(u5_mult_82_SUMB_18__24_), 
        .ZN(u5_mult_82_SUMB_19__23_) );
  INV_X8 u5_mult_82_U60 ( .A(u5_mult_82_n36), .ZN(u5_mult_82_n37) );
  INV_X2 u5_mult_82_U59 ( .A(u5_mult_82_SUMB_18__26_), .ZN(u5_mult_82_n36) );
  CLKBUF_X2 u5_mult_82_U58 ( .A(u5_mult_82_SUMB_46__6_), .Z(u5_mult_82_n35) );
  CLKBUF_X2 u5_mult_82_U57 ( .A(u5_mult_82_CARRYB_6__35_), .Z(u5_mult_82_n34)
         );
  CLKBUF_X2 u5_mult_82_U56 ( .A(u5_mult_82_SUMB_7__45_), .Z(u5_mult_82_n33) );
  BUF_X2 u5_mult_82_U55 ( .A(u5_mult_82_SUMB_18__29_), .Z(u5_mult_82_n32) );
  INV_X4 u5_mult_82_U54 ( .A(u5_mult_82_n30), .ZN(u5_mult_82_n31) );
  INV_X2 u5_mult_82_U53 ( .A(u5_mult_82_SUMB_17__29_), .ZN(u5_mult_82_n30) );
  INV_X1 u5_mult_82_U52 ( .A(u5_mult_82_SUMB_5__39_), .ZN(u5_mult_82_n1477) );
  XNOR2_X2 u5_mult_82_U51 ( .A(u5_mult_82_n1477), .B(u5_mult_82_n5614), .ZN(
        u5_mult_82_SUMB_6__38_) );
  NAND2_X1 u5_mult_82_U50 ( .A1(u5_mult_82_ab_4__31_), .A2(
        u5_mult_82_SUMB_3__32_), .ZN(u5_mult_82_n4266) );
  XNOR2_X2 u5_mult_82_U49 ( .A(u5_mult_82_CARRYB_15__24_), .B(
        u5_mult_82_ab_16__24_), .ZN(u5_mult_82_n29) );
  XNOR2_X2 u5_mult_82_U48 ( .A(u5_mult_82_SUMB_15__25_), .B(u5_mult_82_n29), 
        .ZN(u5_mult_82_SUMB_16__24_) );
  XNOR2_X2 u5_mult_82_U47 ( .A(u5_mult_82_ab_34__34_), .B(
        u5_mult_82_CARRYB_33__34_), .ZN(u5_mult_82_n28) );
  XNOR2_X2 u5_mult_82_U46 ( .A(u5_mult_82_n28), .B(u5_mult_82_SUMB_33__35_), 
        .ZN(u5_mult_82_SUMB_34__34_) );
  CLKBUF_X2 u5_mult_82_U45 ( .A(u5_mult_82_SUMB_41__7_), .Z(u5_mult_82_n27) );
  NAND2_X1 u5_mult_82_U44 ( .A1(u5_mult_82_CARRYB_46__0_), .A2(
        u5_mult_82_SUMB_46__1_), .ZN(u5_mult_82_n4276) );
  XNOR2_X1 u5_mult_82_U43 ( .A(u5_mult_82_CARRYB_46__0_), .B(
        u5_mult_82_ab_47__0_), .ZN(u5_mult_82_n626) );
  XNOR2_X2 u5_mult_82_U42 ( .A(u5_mult_82_ab_7__31_), .B(
        u5_mult_82_CARRYB_6__31_), .ZN(u5_mult_82_n26) );
  XNOR2_X2 u5_mult_82_U41 ( .A(u5_mult_82_n26), .B(u5_mult_82_SUMB_6__32_), 
        .ZN(u5_mult_82_SUMB_7__31_) );
  FA_X1 u5_mult_82_U40 ( .A(u5_mult_82_ab_41__20_), .B(
        u5_mult_82_CARRYB_40__20_), .CI(u5_mult_82_SUMB_40__21_), .S(
        u5_mult_82_n25) );
  INV_X32 u5_mult_82_U39 ( .A(u5_mult_82_ab_26__27_), .ZN(u5_mult_82_n24) );
  XNOR2_X2 u5_mult_82_U38 ( .A(u5_mult_82_CARRYB_25__27_), .B(u5_mult_82_n24), 
        .ZN(u5_mult_82_n1236) );
  XNOR2_X1 u5_mult_82_U37 ( .A(u5_mult_82_CARRYB_5__50_), .B(u5_mult_82_n435), 
        .ZN(u5_mult_82_SUMB_6__50_) );
  XNOR2_X2 u5_mult_82_U36 ( .A(u5_mult_82_ab_39__30_), .B(
        u5_mult_82_CARRYB_38__30_), .ZN(u5_mult_82_n23) );
  XNOR2_X2 u5_mult_82_U35 ( .A(u5_mult_82_n23), .B(u5_mult_82_SUMB_38__31_), 
        .ZN(u5_mult_82_SUMB_39__30_) );
  XNOR2_X2 u5_mult_82_U34 ( .A(u5_mult_82_CARRYB_25__25_), .B(
        u5_mult_82_ab_26__25_), .ZN(u5_mult_82_n22) );
  XNOR2_X2 u5_mult_82_U33 ( .A(u5_mult_82_SUMB_25__26_), .B(u5_mult_82_n22), 
        .ZN(u5_mult_82_SUMB_26__25_) );
  XOR2_X2 u5_mult_82_U32 ( .A(u5_mult_82_n858), .B(u5_mult_82_CARRYB_21__22_), 
        .Z(u5_mult_82_n21) );
  XNOR2_X2 u5_mult_82_U31 ( .A(u5_mult_82_n21), .B(u5_mult_82_SUMB_21__23_), 
        .ZN(u5_mult_82_SUMB_22__22_) );
  INV_X8 u5_mult_82_U30 ( .A(u5_mult_82_n19), .ZN(u5_mult_82_n20) );
  INV_X4 u5_mult_82_U29 ( .A(u5_mult_82_SUMB_28__28_), .ZN(u5_mult_82_n19) );
  XNOR2_X2 u5_mult_82_U28 ( .A(u5_mult_82_ab_33__41_), .B(
        u5_mult_82_CARRYB_32__41_), .ZN(u5_mult_82_n18) );
  XNOR2_X2 u5_mult_82_U27 ( .A(u5_mult_82_n18), .B(u5_mult_82_n1846), .ZN(
        u5_mult_82_SUMB_33__41_) );
  XOR2_X2 u5_mult_82_U26 ( .A(u5_mult_82_n4817), .B(u5_mult_82_CARRYB_20__33_), 
        .Z(u5_mult_82_n17) );
  XNOR2_X1 u5_mult_82_U25 ( .A(u5_mult_82_ab_16__45_), .B(
        u5_mult_82_CARRYB_15__45_), .ZN(u5_mult_82_n16) );
  XNOR2_X2 u5_mult_82_U24 ( .A(u5_mult_82_n16), .B(u5_mult_82_n531), .ZN(
        u5_mult_82_SUMB_16__45_) );
  XNOR2_X2 u5_mult_82_U23 ( .A(u5_mult_82_ab_46__32_), .B(
        u5_mult_82_CARRYB_45__32_), .ZN(u5_mult_82_n15) );
  XNOR2_X2 u5_mult_82_U22 ( .A(u5_mult_82_n15), .B(u5_mult_82_SUMB_45__33_), 
        .ZN(u5_mult_82_SUMB_46__32_) );
  NAND2_X1 u5_mult_82_U21 ( .A1(u5_mult_82_ab_25__25_), .A2(
        u5_mult_82_SUMB_24__26_), .ZN(u5_mult_82_n5973) );
  FA_X1 u5_mult_82_U20 ( .A(u5_mult_82_ab_42__0_), .B(u5_mult_82_CARRYB_41__0_), .CI(u5_mult_82_SUMB_41__1_), .CO(u5_mult_82_n14) );
  INV_X2 u5_mult_82_U19 ( .A(u5_mult_82_n12), .ZN(u5_mult_82_n13) );
  INV_X1 u5_mult_82_U18 ( .A(u5_mult_82_CARRYB_35__2_), .ZN(u5_mult_82_n12) );
  INV_X2 u5_mult_82_U17 ( .A(u5_mult_82_n10), .ZN(u5_mult_82_n11) );
  INV_X1 u5_mult_82_U16 ( .A(u5_mult_82_CARRYB_30__3_), .ZN(u5_mult_82_n10) );
  XNOR2_X1 u5_mult_82_U15 ( .A(u5_mult_82_SUMB_36__7_), .B(
        u5_mult_82_ab_37__6_), .ZN(u5_mult_82_n2123) );
  CLKBUF_X2 u5_mult_82_U14 ( .A(u5_mult_82_SUMB_15__28_), .Z(u5_mult_82_n9) );
  NAND2_X2 u5_mult_82_U13 ( .A1(u5_mult_82_ab_16__43_), .A2(
        u5_mult_82_CARRYB_15__43_), .ZN(u5_mult_82_n2727) );
  XNOR2_X1 u5_mult_82_U12 ( .A(u5_mult_82_ab_36__36_), .B(
        u5_mult_82_CARRYB_35__36_), .ZN(u5_mult_82_n8) );
  XNOR2_X2 u5_mult_82_U11 ( .A(u5_mult_82_n8), .B(u5_mult_82_n710), .ZN(
        u5_mult_82_SUMB_36__36_) );
  CLKBUF_X3 u5_mult_82_U10 ( .A(u5_mult_82_SUMB_48__36_), .Z(u5_mult_82_n7) );
  XNOR2_X2 u5_mult_82_U9 ( .A(u5_mult_82_CARRYB_35__13_), .B(
        u5_mult_82_ab_36__13_), .ZN(u5_mult_82_n6) );
  XNOR2_X2 u5_mult_82_U8 ( .A(u5_mult_82_SUMB_35__14_), .B(u5_mult_82_n6), 
        .ZN(u5_mult_82_SUMB_36__13_) );
  INV_X4 u5_mult_82_U7 ( .A(u5_mult_82_n4), .ZN(u5_mult_82_n5) );
  INV_X2 u5_mult_82_U6 ( .A(u5_mult_82_SUMB_46__37_), .ZN(u5_mult_82_n4) );
  CLKBUF_X2 u5_mult_82_U5 ( .A(u5_mult_82_SUMB_34__36_), .Z(u5_mult_82_n3) );
  NAND2_X1 u5_mult_82_U4 ( .A1(u5_mult_82_SUMB_10__41_), .A2(
        u5_mult_82_CARRYB_10__40_), .ZN(u5_mult_82_n3399) );
  XNOR2_X1 u5_mult_82_U3 ( .A(u5_mult_82_SUMB_10__41_), .B(
        u5_mult_82_ab_11__40_), .ZN(u5_mult_82_n1695) );
  NAND2_X1 u5_mult_82_U2 ( .A1(u5_mult_82_n1726), .A2(u5_mult_82_SUMB_6__41_), 
        .ZN(u5_mult_82_n4020) );
  FA_X1 u5_mult_82_S2_3_35 ( .A(u5_mult_82_ab_3__35_), .B(
        u5_mult_82_CARRYB_2__35_), .CI(u5_mult_82_SUMB_2__36_), .CO(
        u5_mult_82_CARRYB_3__35_), .S(u5_mult_82_SUMB_3__35_) );
  FA_X1 u5_mult_82_S2_51_5 ( .A(u5_mult_82_ab_51__5_), .B(
        u5_mult_82_CARRYB_50__5_), .CI(u5_mult_82_SUMB_50__6_), .CO(
        u5_mult_82_CARRYB_51__5_), .S(u5_mult_82_SUMB_51__5_) );
  FA_X1 u5_mult_82_S2_50_5 ( .A(u5_mult_82_CARRYB_49__5_), .B(
        u5_mult_82_ab_50__5_), .CI(u5_mult_82_SUMB_49__6_), .CO(
        u5_mult_82_CARRYB_50__5_), .S(u5_mult_82_SUMB_50__5_) );
  FA_X1 u5_mult_82_S2_51_4 ( .A(u5_mult_82_ab_51__4_), .B(
        u5_mult_82_CARRYB_50__4_), .CI(u5_mult_82_SUMB_50__5_), .CO(
        u5_mult_82_CARRYB_51__4_), .S(u5_mult_82_SUMB_51__4_) );
  FA_X1 u5_mult_82_S2_5_34 ( .A(u5_mult_82_ab_5__34_), .B(
        u5_mult_82_CARRYB_4__34_), .CI(u5_mult_82_SUMB_4__35_), .CO(
        u5_mult_82_CARRYB_5__34_), .S(u5_mult_82_SUMB_5__34_) );
  FA_X1 u5_mult_82_S2_6_34 ( .A(u5_mult_82_ab_6__34_), .B(
        u5_mult_82_CARRYB_5__34_), .CI(u5_mult_82_SUMB_5__35_), .CO(
        u5_mult_82_CARRYB_6__34_), .S(u5_mult_82_SUMB_6__34_) );
  FA_X1 u5_mult_82_S2_6_33 ( .A(u5_mult_82_ab_6__33_), .B(
        u5_mult_82_CARRYB_5__33_), .CI(u5_mult_82_SUMB_5__34_), .CO(
        u5_mult_82_CARRYB_6__33_), .S(u5_mult_82_SUMB_6__33_) );
  FA_X1 u5_mult_82_S2_7_34 ( .A(u5_mult_82_ab_7__34_), .B(
        u5_mult_82_CARRYB_6__34_), .CI(u5_mult_82_SUMB_6__35_), .CO(
        u5_mult_82_CARRYB_7__34_), .S(u5_mult_82_SUMB_7__34_) );
  FA_X1 u5_mult_82_S2_27_20 ( .A(u5_mult_82_ab_27__20_), .B(
        u5_mult_82_CARRYB_26__20_), .CI(u5_mult_82_SUMB_26__21_), .CO(
        u5_mult_82_CARRYB_27__20_), .S(u5_mult_82_SUMB_27__20_) );
  FA_X1 u5_mult_82_S2_26_21 ( .A(u5_mult_82_CARRYB_25__21_), .B(
        u5_mult_82_ab_26__21_), .CI(u5_mult_82_SUMB_25__22_), .CO(
        u5_mult_82_CARRYB_26__21_), .S(u5_mult_82_SUMB_26__21_) );
  FA_X1 u5_mult_82_S2_25_22 ( .A(u5_mult_82_CARRYB_24__22_), .B(
        u5_mult_82_ab_25__22_), .CI(u5_mult_82_SUMB_24__23_), .CO(
        u5_mult_82_CARRYB_25__22_), .S(u5_mult_82_SUMB_25__22_) );
  FA_X1 u5_mult_82_S2_26_22 ( .A(u5_mult_82_ab_26__22_), .B(
        u5_mult_82_CARRYB_25__22_), .CI(u5_mult_82_SUMB_25__23_), .CO(
        u5_mult_82_CARRYB_26__22_), .S(u5_mult_82_SUMB_26__22_) );
  FA_X1 u5_mult_82_S2_19_26 ( .A(u5_mult_82_ab_19__26_), .B(
        u5_mult_82_CARRYB_18__26_), .CI(u5_mult_82_SUMB_18__27_), .CO(
        u5_mult_82_CARRYB_19__26_), .S(u5_mult_82_SUMB_19__26_) );
  FA_X1 u5_mult_82_S2_18_26 ( .A(u5_mult_82_CARRYB_17__26_), .B(
        u5_mult_82_ab_18__26_), .CI(u5_mult_82_SUMB_17__27_), .CO(
        u5_mult_82_CARRYB_18__26_), .S(u5_mult_82_SUMB_18__26_) );
  FA_X1 u5_mult_82_S2_16_28 ( .A(u5_mult_82_ab_16__28_), .B(
        u5_mult_82_CARRYB_15__28_), .CI(u5_mult_82_SUMB_15__29_), .CO(
        u5_mult_82_CARRYB_16__28_), .S(u5_mult_82_SUMB_16__28_) );
  FA_X1 u5_mult_82_S2_43_11 ( .A(u5_mult_82_CARRYB_42__11_), .B(
        u5_mult_82_ab_43__11_), .CI(u5_mult_82_SUMB_42__12_), .CO(
        u5_mult_82_CARRYB_43__11_), .S(u5_mult_82_SUMB_43__11_) );
  FA_X1 u5_mult_82_S2_41_13 ( .A(u5_mult_82_CARRYB_40__13_), .B(
        u5_mult_82_ab_41__13_), .CI(u5_mult_82_SUMB_40__14_), .CO(
        u5_mult_82_CARRYB_41__13_), .S(u5_mult_82_SUMB_41__13_) );
  FA_X1 u5_mult_82_S2_15_27 ( .A(u5_mult_82_ab_15__27_), .B(
        u5_mult_82_CARRYB_14__27_), .CI(u5_mult_82_SUMB_14__28_), .CO(
        u5_mult_82_CARRYB_15__27_), .S(u5_mult_82_SUMB_15__27_) );
  FA_X1 u5_mult_82_S2_14_28 ( .A(u5_mult_82_ab_14__28_), .B(
        u5_mult_82_CARRYB_13__28_), .CI(u5_mult_82_SUMB_13__29_), .CO(
        u5_mult_82_CARRYB_14__28_), .S(u5_mult_82_SUMB_14__28_) );
  FA_X1 u5_mult_82_S2_15_28 ( .A(u5_mult_82_ab_15__28_), .B(
        u5_mult_82_CARRYB_14__28_), .CI(u5_mult_82_SUMB_14__29_), .CO(
        u5_mult_82_CARRYB_15__28_), .S(u5_mult_82_SUMB_15__28_) );
  FA_X1 u5_mult_82_S2_13_29 ( .A(u5_mult_82_ab_13__29_), .B(
        u5_mult_82_CARRYB_12__29_), .CI(u5_mult_82_SUMB_12__30_), .CO(
        u5_mult_82_CARRYB_13__29_), .S(u5_mult_82_SUMB_13__29_) );
  FA_X1 u5_mult_82_S2_13_30 ( .A(u5_mult_82_ab_13__30_), .B(
        u5_mult_82_CARRYB_12__30_), .CI(u5_mult_82_SUMB_12__31_), .CO(
        u5_mult_82_CARRYB_13__30_), .S(u5_mult_82_SUMB_13__30_) );
  FA_X1 u5_mult_82_S2_12_31 ( .A(u5_mult_82_ab_12__31_), .B(
        u5_mult_82_CARRYB_11__31_), .CI(u5_mult_82_SUMB_11__32_), .CO(
        u5_mult_82_CARRYB_12__31_), .S(u5_mult_82_SUMB_12__31_) );
  FA_X1 u5_mult_82_S2_10_32 ( .A(u5_mult_82_SUMB_9__33_), .B(
        u5_mult_82_ab_10__32_), .CI(u5_mult_82_CARRYB_9__32_), .CO(
        u5_mult_82_CARRYB_10__32_), .S(u5_mult_82_SUMB_10__32_) );
  FA_X1 u5_mult_82_S2_11_32 ( .A(u5_mult_82_CARRYB_10__32_), .B(
        u5_mult_82_ab_11__32_), .CI(u5_mult_82_SUMB_10__33_), .CO(
        u5_mult_82_CARRYB_11__32_), .S(u5_mult_82_SUMB_11__32_) );
  FA_X1 u5_mult_82_S2_9_33 ( .A(u5_mult_82_ab_9__33_), .B(
        u5_mult_82_SUMB_8__34_), .CI(u5_mult_82_CARRYB_8__33_), .CO(
        u5_mult_82_CARRYB_9__33_), .S(u5_mult_82_SUMB_9__33_) );
  FA_X1 u5_mult_82_S2_10_33 ( .A(u5_mult_82_ab_10__33_), .B(
        u5_mult_82_CARRYB_9__33_), .CI(u5_mult_82_SUMB_9__34_), .CO(
        u5_mult_82_CARRYB_10__33_), .S(u5_mult_82_SUMB_10__33_) );
  FA_X1 u5_mult_82_S2_8_33 ( .A(u5_mult_82_ab_8__33_), .B(
        u5_mult_82_CARRYB_7__33_), .CI(u5_mult_82_SUMB_7__34_), .CO(
        u5_mult_82_CARRYB_8__33_), .S(u5_mult_82_SUMB_8__33_) );
  FA_X1 u5_mult_82_S2_9_32 ( .A(u5_mult_82_ab_9__32_), .B(
        u5_mult_82_CARRYB_8__32_), .CI(u5_mult_82_SUMB_8__33_), .CO(
        u5_mult_82_CARRYB_9__32_), .S(u5_mult_82_SUMB_9__32_) );
  FA_X1 u5_mult_82_S2_6_35 ( .A(u5_mult_82_ab_6__35_), .B(
        u5_mult_82_CARRYB_5__35_), .CI(u5_mult_82_SUMB_5__36_), .CO(
        u5_mult_82_CARRYB_6__35_), .S(u5_mult_82_SUMB_6__35_) );
  FA_X1 u5_mult_82_S2_34_16 ( .A(u5_mult_82_CARRYB_33__16_), .B(
        u5_mult_82_ab_34__16_), .CI(u5_mult_82_SUMB_33__17_), .CO(
        u5_mult_82_CARRYB_34__16_), .S(u5_mult_82_SUMB_34__16_) );
  FA_X1 u5_mult_82_S2_47_8 ( .A(u5_mult_82_ab_47__8_), .B(
        u5_mult_82_CARRYB_46__8_), .CI(u5_mult_82_SUMB_46__9_), .CO(
        u5_mult_82_CARRYB_47__8_), .S(u5_mult_82_SUMB_47__8_) );
  FA_X1 u5_mult_82_S2_23_23 ( .A(u5_mult_82_ab_23__23_), .B(
        u5_mult_82_CARRYB_22__23_), .CI(u5_mult_82_SUMB_22__24_), .CO(
        u5_mult_82_CARRYB_23__23_), .S(u5_mult_82_SUMB_23__23_) );
  FA_X1 u5_mult_82_S2_38_14 ( .A(u5_mult_82_ab_38__14_), .B(
        u5_mult_82_CARRYB_37__14_), .CI(u5_mult_82_SUMB_37__15_), .CO(
        u5_mult_82_CARRYB_38__14_), .S(u5_mult_82_SUMB_38__14_) );
  FA_X1 u5_mult_82_S2_2_49 ( .A(u5_mult_82_ab_2__49_), .B(
        u5_mult_82_CARRYB_1__49_), .CI(u5_mult_82_SUMB_1__50_), .CO(
        u5_mult_82_CARRYB_2__49_), .S(u5_mult_82_SUMB_2__49_) );
  FA_X1 u5_mult_82_S2_2_48 ( .A(u5_mult_82_ab_2__48_), .B(
        u5_mult_82_CARRYB_1__48_), .CI(u5_mult_82_SUMB_1__49_), .CO(
        u5_mult_82_CARRYB_2__48_), .S(u5_mult_82_SUMB_2__48_) );
  FA_X1 u5_mult_82_S2_2_44 ( .A(u5_mult_82_ab_2__44_), .B(
        u5_mult_82_CARRYB_1__44_), .CI(u5_mult_82_SUMB_1__45_), .CO(
        u5_mult_82_CARRYB_2__44_), .S(u5_mult_82_SUMB_2__44_) );
  FA_X1 u5_mult_82_S2_2_43 ( .A(u5_mult_82_ab_2__43_), .B(
        u5_mult_82_CARRYB_1__43_), .CI(u5_mult_82_SUMB_1__44_), .CO(
        u5_mult_82_CARRYB_2__43_), .S(u5_mult_82_SUMB_2__43_) );
  FA_X1 u5_mult_82_S2_2_41 ( .A(u5_mult_82_ab_2__41_), .B(
        u5_mult_82_CARRYB_1__41_), .CI(u5_mult_82_SUMB_1__42_), .CO(
        u5_mult_82_CARRYB_2__41_), .S(u5_mult_82_SUMB_2__41_) );
  FA_X1 u5_mult_82_S2_2_40 ( .A(u5_mult_82_ab_2__40_), .B(u5_mult_82_n467), 
        .CI(u5_mult_82_n466), .CO(u5_mult_82_CARRYB_2__40_), .S(
        u5_mult_82_SUMB_2__40_) );
  FA_X1 u5_mult_82_S2_2_39 ( .A(u5_mult_82_SUMB_1__40_), .B(u5_mult_82_n2132), 
        .CI(u5_mult_82_ab_2__39_), .CO(u5_mult_82_CARRYB_2__39_), .S(
        u5_mult_82_SUMB_2__39_) );
  FA_X1 u5_mult_82_S2_2_38 ( .A(u5_mult_82_ab_2__38_), .B(u5_mult_82_n612), 
        .CI(u5_mult_82_n2310), .CO(u5_mult_82_CARRYB_2__38_), .S(
        u5_mult_82_SUMB_2__38_) );
  FA_X1 u5_mult_82_S2_2_37 ( .A(u5_mult_82_ab_2__37_), .B(
        u5_mult_82_CARRYB_1__37_), .CI(u5_mult_82_SUMB_1__38_), .CO(
        u5_mult_82_CARRYB_2__37_), .S(u5_mult_82_SUMB_2__37_) );
  FA_X1 u5_mult_82_S2_2_34 ( .A(u5_mult_82_ab_2__34_), .B(
        u5_mult_82_CARRYB_1__34_), .CI(u5_mult_82_SUMB_1__35_), .CO(
        u5_mult_82_CARRYB_2__34_), .S(u5_mult_82_SUMB_2__34_) );
  FA_X1 u5_mult_82_S2_2_33 ( .A(u5_mult_82_ab_2__33_), .B(u5_mult_82_n610), 
        .CI(u5_mult_82_n804), .CO(u5_mult_82_CARRYB_2__33_), .S(
        u5_mult_82_SUMB_2__33_) );
  FA_X1 u5_mult_82_S2_2_31 ( .A(u5_mult_82_ab_2__31_), .B(u5_mult_82_n599), 
        .CI(u5_mult_82_n468), .CO(u5_mult_82_CARRYB_2__31_), .S(
        u5_mult_82_SUMB_2__31_) );
  FA_X1 u5_mult_82_S2_2_25 ( .A(u5_mult_82_ab_2__25_), .B(
        u5_mult_82_CARRYB_1__25_), .CI(u5_mult_82_SUMB_1__26_), .CO(
        u5_mult_82_CARRYB_2__25_), .S(u5_mult_82_SUMB_2__25_) );
  FA_X1 u5_mult_82_S2_2_24 ( .A(u5_mult_82_ab_2__24_), .B(
        u5_mult_82_CARRYB_1__24_), .CI(u5_mult_82_SUMB_1__25_), .CO(
        u5_mult_82_CARRYB_2__24_), .S(u5_mult_82_SUMB_2__24_) );
  FA_X1 u5_mult_82_S2_2_23 ( .A(u5_mult_82_ab_2__23_), .B(
        u5_mult_82_CARRYB_1__23_), .CI(u5_mult_82_SUMB_1__24_), .CO(
        u5_mult_82_CARRYB_2__23_), .S(u5_mult_82_SUMB_2__23_) );
  FA_X1 u5_mult_82_S2_2_22 ( .A(u5_mult_82_ab_2__22_), .B(u5_mult_82_n474), 
        .CI(u5_mult_82_SUMB_1__23_), .CO(u5_mult_82_CARRYB_2__22_), .S(
        u5_mult_82_SUMB_2__22_) );
  FA_X1 u5_mult_82_S2_2_21 ( .A(u5_mult_82_ab_2__21_), .B(
        u5_mult_82_CARRYB_1__21_), .CI(u5_mult_82_SUMB_1__22_), .CO(
        u5_mult_82_CARRYB_2__21_), .S(u5_mult_82_SUMB_2__21_) );
  FA_X1 u5_mult_82_S2_2_20 ( .A(u5_mult_82_ab_2__20_), .B(u5_mult_82_n472), 
        .CI(u5_mult_82_n473), .CO(u5_mult_82_CARRYB_2__20_), .S(
        u5_mult_82_SUMB_2__20_) );
  FA_X1 u5_mult_82_S2_2_19 ( .A(u5_mult_82_ab_2__19_), .B(
        u5_mult_82_CARRYB_1__19_), .CI(u5_mult_82_SUMB_1__20_), .CO(
        u5_mult_82_CARRYB_2__19_), .S(u5_mult_82_SUMB_2__19_) );
  FA_X1 u5_mult_82_S2_2_18 ( .A(u5_mult_82_ab_2__18_), .B(
        u5_mult_82_CARRYB_1__18_), .CI(u5_mult_82_SUMB_1__19_), .CO(
        u5_mult_82_CARRYB_2__18_), .S(u5_mult_82_SUMB_2__18_) );
  FA_X1 u5_mult_82_S2_2_17 ( .A(u5_mult_82_ab_2__17_), .B(u5_mult_82_n471), 
        .CI(u5_mult_82_n614), .CO(u5_mult_82_CARRYB_2__17_), .S(
        u5_mult_82_SUMB_2__17_) );
  FA_X1 u5_mult_82_S2_2_16 ( .A(u5_mult_82_ab_2__16_), .B(
        u5_mult_82_CARRYB_1__16_), .CI(u5_mult_82_SUMB_1__17_), .CO(
        u5_mult_82_CARRYB_2__16_), .S(u5_mult_82_SUMB_2__16_) );
  FA_X1 u5_mult_82_S2_2_15 ( .A(u5_mult_82_ab_2__15_), .B(u5_mult_82_n475), 
        .CI(u5_mult_82_SUMB_1__16_), .CO(u5_mult_82_CARRYB_2__15_), .S(
        u5_mult_82_SUMB_2__15_) );
  FA_X1 u5_mult_82_S2_2_14 ( .A(u5_mult_82_ab_2__14_), .B(
        u5_mult_82_CARRYB_1__14_), .CI(u5_mult_82_SUMB_1__15_), .CO(
        u5_mult_82_CARRYB_2__14_), .S(u5_mult_82_SUMB_2__14_) );
  FA_X1 u5_mult_82_S2_2_13 ( .A(u5_mult_82_ab_2__13_), .B(
        u5_mult_82_CARRYB_1__13_), .CI(u5_mult_82_SUMB_1__14_), .CO(
        u5_mult_82_CARRYB_2__13_), .S(u5_mult_82_SUMB_2__13_) );
  FA_X1 u5_mult_82_S2_2_12 ( .A(u5_mult_82_ab_2__12_), .B(
        u5_mult_82_CARRYB_1__12_), .CI(u5_mult_82_SUMB_1__13_), .CO(
        u5_mult_82_CARRYB_2__12_), .S(u5_mult_82_SUMB_2__12_) );
  FA_X1 u5_mult_82_S2_2_11 ( .A(u5_mult_82_ab_2__11_), .B(
        u5_mult_82_CARRYB_1__11_), .CI(u5_mult_82_SUMB_1__12_), .CO(
        u5_mult_82_CARRYB_2__11_), .S(u5_mult_82_SUMB_2__11_) );
  FA_X1 u5_mult_82_S2_2_10 ( .A(u5_mult_82_ab_2__10_), .B(u5_mult_82_n611), 
        .CI(u5_mult_82_SUMB_1__11_), .CO(u5_mult_82_CARRYB_2__10_), .S(
        u5_mult_82_SUMB_2__10_) );
  FA_X1 u5_mult_82_S2_2_9 ( .A(u5_mult_82_ab_2__9_), .B(
        u5_mult_82_CARRYB_1__9_), .CI(u5_mult_82_n476), .CO(
        u5_mult_82_CARRYB_2__9_), .S(u5_mult_82_SUMB_2__9_) );
  FA_X1 u5_mult_82_S2_2_8 ( .A(u5_mult_82_ab_2__8_), .B(u5_mult_82_n477), .CI(
        u5_mult_82_SUMB_1__9_), .CO(u5_mult_82_CARRYB_2__8_), .S(
        u5_mult_82_SUMB_2__8_) );
  FA_X1 u5_mult_82_S2_2_7 ( .A(u5_mult_82_ab_2__7_), .B(
        u5_mult_82_CARRYB_1__7_), .CI(u5_mult_82_SUMB_1__8_), .CO(
        u5_mult_82_CARRYB_2__7_), .S(u5_mult_82_SUMB_2__7_) );
  FA_X1 u5_mult_82_S2_2_6 ( .A(u5_mult_82_ab_2__6_), .B(
        u5_mult_82_CARRYB_1__6_), .CI(u5_mult_82_SUMB_1__7_), .CO(
        u5_mult_82_CARRYB_2__6_), .S(u5_mult_82_SUMB_2__6_) );
  FA_X1 u5_mult_82_S2_2_5 ( .A(u5_mult_82_ab_2__5_), .B(
        u5_mult_82_CARRYB_1__5_), .CI(u5_mult_82_SUMB_1__6_), .CO(
        u5_mult_82_CARRYB_2__5_), .S(u5_mult_82_SUMB_2__5_) );
  FA_X1 u5_mult_82_S2_2_4 ( .A(u5_mult_82_ab_2__4_), .B(u5_mult_82_n623), .CI(
        u5_mult_82_SUMB_1__5_), .CO(u5_mult_82_CARRYB_2__4_), .S(
        u5_mult_82_SUMB_2__4_) );
  FA_X1 u5_mult_82_S2_2_3 ( .A(u5_mult_82_ab_2__3_), .B(
        u5_mult_82_CARRYB_1__3_), .CI(u5_mult_82_n478), .CO(
        u5_mult_82_CARRYB_2__3_), .S(u5_mult_82_SUMB_2__3_) );
  FA_X1 u5_mult_82_S2_2_2 ( .A(u5_mult_82_ab_2__2_), .B(
        u5_mult_82_CARRYB_1__2_), .CI(u5_mult_82_SUMB_1__3_), .CO(
        u5_mult_82_CARRYB_2__2_), .S(u5_mult_82_SUMB_2__2_) );
  FA_X1 u5_mult_82_S2_2_1 ( .A(u5_mult_82_ab_2__1_), .B(u5_mult_82_n480), .CI(
        u5_mult_82_SUMB_1__2_), .CO(u5_mult_82_CARRYB_2__1_), .S(
        u5_mult_82_SUMB_2__1_) );
  FA_X1 u5_mult_82_S1_2_0 ( .A(u5_mult_82_ab_2__0_), .B(
        u5_mult_82_CARRYB_1__0_), .CI(u5_mult_82_n479), .CO(
        u5_mult_82_CARRYB_2__0_), .S(u5_N2) );
  FA_X1 u5_mult_82_S2_3_49 ( .A(u5_mult_82_ab_3__49_), .B(
        u5_mult_82_CARRYB_2__49_), .CI(u5_mult_82_SUMB_2__50_), .CO(
        u5_mult_82_CARRYB_3__49_), .S(u5_mult_82_SUMB_3__49_) );
  FA_X1 u5_mult_82_S2_3_48 ( .A(u5_mult_82_ab_3__48_), .B(
        u5_mult_82_CARRYB_2__48_), .CI(u5_mult_82_SUMB_2__49_), .CO(
        u5_mult_82_CARRYB_3__48_), .S(u5_mult_82_SUMB_3__48_) );
  FA_X1 u5_mult_82_S2_3_45 ( .A(u5_mult_82_ab_3__45_), .B(
        u5_mult_82_CARRYB_2__45_), .CI(u5_mult_82_SUMB_2__46_), .CO(
        u5_mult_82_CARRYB_3__45_), .S(u5_mult_82_SUMB_3__45_) );
  FA_X1 u5_mult_82_S2_3_44 ( .A(u5_mult_82_CARRYB_2__44_), .B(
        u5_mult_82_ab_3__44_), .CI(u5_mult_82_SUMB_2__45_), .CO(
        u5_mult_82_CARRYB_3__44_), .S(u5_mult_82_SUMB_3__44_) );
  FA_X1 u5_mult_82_S2_3_38 ( .A(u5_mult_82_CARRYB_2__38_), .B(
        u5_mult_82_ab_3__38_), .CI(u5_mult_82_SUMB_2__39_), .CO(
        u5_mult_82_CARRYB_3__38_), .S(u5_mult_82_SUMB_3__38_) );
  FA_X1 u5_mult_82_S2_3_37 ( .A(u5_mult_82_ab_3__37_), .B(
        u5_mult_82_CARRYB_2__37_), .CI(u5_mult_82_SUMB_2__38_), .CO(
        u5_mult_82_CARRYB_3__37_), .S(u5_mult_82_SUMB_3__37_) );
  FA_X1 u5_mult_82_S2_3_32 ( .A(u5_mult_82_ab_3__32_), .B(
        u5_mult_82_CARRYB_2__32_), .CI(u5_mult_82_SUMB_2__33_), .CO(
        u5_mult_82_CARRYB_3__32_), .S(u5_mult_82_SUMB_3__32_) );
  FA_X1 u5_mult_82_S2_3_30 ( .A(u5_mult_82_ab_3__30_), .B(
        u5_mult_82_CARRYB_2__30_), .CI(u5_mult_82_SUMB_2__31_), .CO(
        u5_mult_82_CARRYB_3__30_), .S(u5_mult_82_SUMB_3__30_) );
  FA_X1 u5_mult_82_S2_3_27 ( .A(u5_mult_82_ab_3__27_), .B(
        u5_mult_82_CARRYB_2__27_), .CI(u5_mult_82_SUMB_2__28_), .CO(
        u5_mult_82_CARRYB_3__27_), .S(u5_mult_82_SUMB_3__27_) );
  FA_X1 u5_mult_82_S2_3_23 ( .A(u5_mult_82_ab_3__23_), .B(
        u5_mult_82_CARRYB_2__23_), .CI(u5_mult_82_SUMB_2__24_), .CO(
        u5_mult_82_CARRYB_3__23_), .S(u5_mult_82_SUMB_3__23_) );
  FA_X1 u5_mult_82_S2_3_22 ( .A(u5_mult_82_ab_3__22_), .B(
        u5_mult_82_CARRYB_2__22_), .CI(u5_mult_82_SUMB_2__23_), .CO(
        u5_mult_82_CARRYB_3__22_), .S(u5_mult_82_SUMB_3__22_) );
  FA_X1 u5_mult_82_S2_3_21 ( .A(u5_mult_82_ab_3__21_), .B(
        u5_mult_82_CARRYB_2__21_), .CI(u5_mult_82_SUMB_2__22_), .CO(
        u5_mult_82_CARRYB_3__21_), .S(u5_mult_82_SUMB_3__21_) );
  FA_X1 u5_mult_82_S2_3_20 ( .A(u5_mult_82_ab_3__20_), .B(
        u5_mult_82_CARRYB_2__20_), .CI(u5_mult_82_SUMB_2__21_), .CO(
        u5_mult_82_CARRYB_3__20_), .S(u5_mult_82_SUMB_3__20_) );
  FA_X1 u5_mult_82_S2_3_19 ( .A(u5_mult_82_ab_3__19_), .B(
        u5_mult_82_CARRYB_2__19_), .CI(u5_mult_82_SUMB_2__20_), .CO(
        u5_mult_82_CARRYB_3__19_), .S(u5_mult_82_SUMB_3__19_) );
  FA_X1 u5_mult_82_S2_3_18 ( .A(u5_mult_82_ab_3__18_), .B(
        u5_mult_82_CARRYB_2__18_), .CI(u5_mult_82_SUMB_2__19_), .CO(
        u5_mult_82_CARRYB_3__18_), .S(u5_mult_82_SUMB_3__18_) );
  FA_X1 u5_mult_82_S2_3_17 ( .A(u5_mult_82_ab_3__17_), .B(
        u5_mult_82_CARRYB_2__17_), .CI(u5_mult_82_SUMB_2__18_), .CO(
        u5_mult_82_CARRYB_3__17_), .S(u5_mult_82_SUMB_3__17_) );
  FA_X1 u5_mult_82_S2_3_16 ( .A(u5_mult_82_ab_3__16_), .B(
        u5_mult_82_CARRYB_2__16_), .CI(u5_mult_82_SUMB_2__17_), .CO(
        u5_mult_82_CARRYB_3__16_), .S(u5_mult_82_SUMB_3__16_) );
  FA_X1 u5_mult_82_S2_3_15 ( .A(u5_mult_82_ab_3__15_), .B(
        u5_mult_82_CARRYB_2__15_), .CI(u5_mult_82_SUMB_2__16_), .CO(
        u5_mult_82_CARRYB_3__15_), .S(u5_mult_82_SUMB_3__15_) );
  FA_X1 u5_mult_82_S2_3_14 ( .A(u5_mult_82_ab_3__14_), .B(
        u5_mult_82_CARRYB_2__14_), .CI(u5_mult_82_SUMB_2__15_), .CO(
        u5_mult_82_CARRYB_3__14_), .S(u5_mult_82_SUMB_3__14_) );
  FA_X1 u5_mult_82_S2_3_13 ( .A(u5_mult_82_ab_3__13_), .B(
        u5_mult_82_CARRYB_2__13_), .CI(u5_mult_82_SUMB_2__14_), .CO(
        u5_mult_82_CARRYB_3__13_), .S(u5_mult_82_SUMB_3__13_) );
  FA_X1 u5_mult_82_S2_3_12 ( .A(u5_mult_82_ab_3__12_), .B(
        u5_mult_82_CARRYB_2__12_), .CI(u5_mult_82_SUMB_2__13_), .CO(
        u5_mult_82_CARRYB_3__12_), .S(u5_mult_82_SUMB_3__12_) );
  FA_X1 u5_mult_82_S2_3_11 ( .A(u5_mult_82_ab_3__11_), .B(
        u5_mult_82_CARRYB_2__11_), .CI(u5_mult_82_SUMB_2__12_), .CO(
        u5_mult_82_CARRYB_3__11_), .S(u5_mult_82_SUMB_3__11_) );
  FA_X1 u5_mult_82_S2_3_10 ( .A(u5_mult_82_ab_3__10_), .B(
        u5_mult_82_CARRYB_2__10_), .CI(u5_mult_82_SUMB_2__11_), .CO(
        u5_mult_82_CARRYB_3__10_), .S(u5_mult_82_SUMB_3__10_) );
  FA_X1 u5_mult_82_S2_3_9 ( .A(u5_mult_82_ab_3__9_), .B(
        u5_mult_82_CARRYB_2__9_), .CI(u5_mult_82_SUMB_2__10_), .CO(
        u5_mult_82_CARRYB_3__9_), .S(u5_mult_82_SUMB_3__9_) );
  FA_X1 u5_mult_82_S2_3_8 ( .A(u5_mult_82_ab_3__8_), .B(
        u5_mult_82_CARRYB_2__8_), .CI(u5_mult_82_SUMB_2__9_), .CO(
        u5_mult_82_CARRYB_3__8_), .S(u5_mult_82_SUMB_3__8_) );
  FA_X1 u5_mult_82_S2_3_7 ( .A(u5_mult_82_ab_3__7_), .B(
        u5_mult_82_CARRYB_2__7_), .CI(u5_mult_82_SUMB_2__8_), .CO(
        u5_mult_82_CARRYB_3__7_), .S(u5_mult_82_SUMB_3__7_) );
  FA_X1 u5_mult_82_S2_3_6 ( .A(u5_mult_82_ab_3__6_), .B(
        u5_mult_82_CARRYB_2__6_), .CI(u5_mult_82_SUMB_2__7_), .CO(
        u5_mult_82_CARRYB_3__6_), .S(u5_mult_82_SUMB_3__6_) );
  FA_X1 u5_mult_82_S2_3_5 ( .A(u5_mult_82_ab_3__5_), .B(
        u5_mult_82_CARRYB_2__5_), .CI(u5_mult_82_SUMB_2__6_), .CO(
        u5_mult_82_CARRYB_3__5_), .S(u5_mult_82_SUMB_3__5_) );
  FA_X1 u5_mult_82_S2_3_4 ( .A(u5_mult_82_ab_3__4_), .B(
        u5_mult_82_CARRYB_2__4_), .CI(u5_mult_82_SUMB_2__5_), .CO(
        u5_mult_82_CARRYB_3__4_), .S(u5_mult_82_SUMB_3__4_) );
  FA_X1 u5_mult_82_S2_3_3 ( .A(u5_mult_82_ab_3__3_), .B(
        u5_mult_82_CARRYB_2__3_), .CI(u5_mult_82_SUMB_2__4_), .CO(
        u5_mult_82_CARRYB_3__3_), .S(u5_mult_82_SUMB_3__3_) );
  FA_X1 u5_mult_82_S2_3_2 ( .A(u5_mult_82_ab_3__2_), .B(
        u5_mult_82_CARRYB_2__2_), .CI(u5_mult_82_SUMB_2__3_), .CO(
        u5_mult_82_CARRYB_3__2_), .S(u5_mult_82_SUMB_3__2_) );
  FA_X1 u5_mult_82_S2_3_1 ( .A(u5_mult_82_ab_3__1_), .B(
        u5_mult_82_CARRYB_2__1_), .CI(u5_mult_82_SUMB_2__2_), .CO(
        u5_mult_82_CARRYB_3__1_), .S(u5_mult_82_SUMB_3__1_) );
  FA_X1 u5_mult_82_S1_3_0 ( .A(u5_mult_82_ab_3__0_), .B(
        u5_mult_82_CARRYB_2__0_), .CI(u5_mult_82_SUMB_2__1_), .CO(
        u5_mult_82_CARRYB_3__0_), .S(u5_N3) );
  FA_X1 u5_mult_82_S3_4_51 ( .A(u5_mult_82_ab_4__51_), .B(u5_mult_82_ab_3__52_), .CI(u5_mult_82_CARRYB_3__51_), .CO(u5_mult_82_CARRYB_4__51_), .S(
        u5_mult_82_SUMB_4__51_) );
  FA_X1 u5_mult_82_S2_4_50 ( .A(u5_mult_82_SUMB_3__51_), .B(
        u5_mult_82_ab_4__50_), .CI(u5_mult_82_CARRYB_3__50_), .CO(
        u5_mult_82_CARRYB_4__50_), .S(u5_mult_82_SUMB_4__50_) );
  FA_X1 u5_mult_82_S2_4_48 ( .A(u5_mult_82_CARRYB_3__48_), .B(
        u5_mult_82_ab_4__48_), .CI(u5_mult_82_SUMB_3__49_), .CO(
        u5_mult_82_CARRYB_4__48_), .S(u5_mult_82_SUMB_4__48_) );
  FA_X1 u5_mult_82_S2_4_45 ( .A(u5_mult_82_ab_4__45_), .B(
        u5_mult_82_CARRYB_3__45_), .CI(u5_mult_82_SUMB_3__46_), .CO(
        u5_mult_82_CARRYB_4__45_), .S(u5_mult_82_SUMB_4__45_) );
  FA_X1 u5_mult_82_S2_4_44 ( .A(u5_mult_82_ab_4__44_), .B(
        u5_mult_82_CARRYB_3__44_), .CI(u5_mult_82_SUMB_3__45_), .CO(
        u5_mult_82_CARRYB_4__44_), .S(u5_mult_82_SUMB_4__44_) );
  FA_X1 u5_mult_82_S2_4_43 ( .A(u5_mult_82_ab_4__43_), .B(
        u5_mult_82_CARRYB_3__43_), .CI(u5_mult_82_SUMB_3__44_), .CO(
        u5_mult_82_CARRYB_4__43_), .S(u5_mult_82_SUMB_4__43_) );
  FA_X1 u5_mult_82_S2_4_42 ( .A(u5_mult_82_CARRYB_3__42_), .B(
        u5_mult_82_ab_4__42_), .CI(u5_mult_82_SUMB_3__43_), .CO(
        u5_mult_82_CARRYB_4__42_), .S(u5_mult_82_SUMB_4__42_) );
  FA_X1 u5_mult_82_S2_4_40 ( .A(u5_mult_82_ab_4__40_), .B(
        u5_mult_82_CARRYB_3__40_), .CI(u5_mult_82_SUMB_3__41_), .CO(
        u5_mult_82_CARRYB_4__40_), .S(u5_mult_82_SUMB_4__40_) );
  FA_X1 u5_mult_82_S2_4_32 ( .A(u5_mult_82_ab_4__32_), .B(
        u5_mult_82_CARRYB_3__32_), .CI(u5_mult_82_SUMB_3__33_), .CO(
        u5_mult_82_CARRYB_4__32_), .S(u5_mult_82_SUMB_4__32_) );
  FA_X1 u5_mult_82_S2_4_30 ( .A(u5_mult_82_ab_4__30_), .B(
        u5_mult_82_CARRYB_3__30_), .CI(u5_mult_82_SUMB_3__31_), .CO(
        u5_mult_82_CARRYB_4__30_), .S(u5_mult_82_SUMB_4__30_) );
  FA_X1 u5_mult_82_S2_4_27 ( .A(u5_mult_82_ab_4__27_), .B(
        u5_mult_82_CARRYB_3__27_), .CI(u5_mult_82_SUMB_3__28_), .CO(
        u5_mult_82_CARRYB_4__27_), .S(u5_mult_82_SUMB_4__27_) );
  FA_X1 u5_mult_82_S2_4_25 ( .A(u5_mult_82_ab_4__25_), .B(
        u5_mult_82_CARRYB_3__25_), .CI(u5_mult_82_SUMB_3__26_), .CO(
        u5_mult_82_CARRYB_4__25_), .S(u5_mult_82_SUMB_4__25_) );
  FA_X1 u5_mult_82_S2_4_24 ( .A(u5_mult_82_CARRYB_3__24_), .B(
        u5_mult_82_ab_4__24_), .CI(u5_mult_82_SUMB_3__25_), .CO(
        u5_mult_82_CARRYB_4__24_), .S(u5_mult_82_SUMB_4__24_) );
  FA_X1 u5_mult_82_S2_4_21 ( .A(u5_mult_82_ab_4__21_), .B(
        u5_mult_82_CARRYB_3__21_), .CI(u5_mult_82_SUMB_3__22_), .CO(
        u5_mult_82_CARRYB_4__21_), .S(u5_mult_82_SUMB_4__21_) );
  FA_X1 u5_mult_82_S2_4_19 ( .A(u5_mult_82_ab_4__19_), .B(
        u5_mult_82_CARRYB_3__19_), .CI(u5_mult_82_SUMB_3__20_), .CO(
        u5_mult_82_CARRYB_4__19_), .S(u5_mult_82_SUMB_4__19_) );
  FA_X1 u5_mult_82_S2_4_18 ( .A(u5_mult_82_ab_4__18_), .B(
        u5_mult_82_CARRYB_3__18_), .CI(u5_mult_82_SUMB_3__19_), .CO(
        u5_mult_82_CARRYB_4__18_), .S(u5_mult_82_SUMB_4__18_) );
  FA_X1 u5_mult_82_S2_4_17 ( .A(u5_mult_82_ab_4__17_), .B(
        u5_mult_82_CARRYB_3__17_), .CI(u5_mult_82_SUMB_3__18_), .CO(
        u5_mult_82_CARRYB_4__17_), .S(u5_mult_82_SUMB_4__17_) );
  FA_X1 u5_mult_82_S2_4_16 ( .A(u5_mult_82_ab_4__16_), .B(
        u5_mult_82_CARRYB_3__16_), .CI(u5_mult_82_SUMB_3__17_), .CO(
        u5_mult_82_CARRYB_4__16_), .S(u5_mult_82_SUMB_4__16_) );
  FA_X1 u5_mult_82_S2_4_15 ( .A(u5_mult_82_ab_4__15_), .B(
        u5_mult_82_CARRYB_3__15_), .CI(u5_mult_82_SUMB_3__16_), .CO(
        u5_mult_82_CARRYB_4__15_), .S(u5_mult_82_SUMB_4__15_) );
  FA_X1 u5_mult_82_S2_4_14 ( .A(u5_mult_82_ab_4__14_), .B(
        u5_mult_82_CARRYB_3__14_), .CI(u5_mult_82_SUMB_3__15_), .CO(
        u5_mult_82_CARRYB_4__14_), .S(u5_mult_82_SUMB_4__14_) );
  FA_X1 u5_mult_82_S2_4_13 ( .A(u5_mult_82_ab_4__13_), .B(
        u5_mult_82_CARRYB_3__13_), .CI(u5_mult_82_SUMB_3__14_), .CO(
        u5_mult_82_CARRYB_4__13_), .S(u5_mult_82_SUMB_4__13_) );
  FA_X1 u5_mult_82_S2_4_12 ( .A(u5_mult_82_ab_4__12_), .B(
        u5_mult_82_CARRYB_3__12_), .CI(u5_mult_82_SUMB_3__13_), .CO(
        u5_mult_82_CARRYB_4__12_), .S(u5_mult_82_SUMB_4__12_) );
  FA_X1 u5_mult_82_S2_4_11 ( .A(u5_mult_82_ab_4__11_), .B(
        u5_mult_82_CARRYB_3__11_), .CI(u5_mult_82_SUMB_3__12_), .CO(
        u5_mult_82_CARRYB_4__11_), .S(u5_mult_82_SUMB_4__11_) );
  FA_X1 u5_mult_82_S2_4_10 ( .A(u5_mult_82_ab_4__10_), .B(
        u5_mult_82_CARRYB_3__10_), .CI(u5_mult_82_SUMB_3__11_), .CO(
        u5_mult_82_CARRYB_4__10_), .S(u5_mult_82_SUMB_4__10_) );
  FA_X1 u5_mult_82_S2_4_9 ( .A(u5_mult_82_ab_4__9_), .B(
        u5_mult_82_CARRYB_3__9_), .CI(u5_mult_82_SUMB_3__10_), .CO(
        u5_mult_82_CARRYB_4__9_), .S(u5_mult_82_SUMB_4__9_) );
  FA_X1 u5_mult_82_S2_4_8 ( .A(u5_mult_82_ab_4__8_), .B(
        u5_mult_82_CARRYB_3__8_), .CI(u5_mult_82_SUMB_3__9_), .CO(
        u5_mult_82_CARRYB_4__8_), .S(u5_mult_82_SUMB_4__8_) );
  FA_X1 u5_mult_82_S2_4_7 ( .A(u5_mult_82_ab_4__7_), .B(
        u5_mult_82_CARRYB_3__7_), .CI(u5_mult_82_SUMB_3__8_), .CO(
        u5_mult_82_CARRYB_4__7_), .S(u5_mult_82_SUMB_4__7_) );
  FA_X1 u5_mult_82_S2_4_6 ( .A(u5_mult_82_ab_4__6_), .B(
        u5_mult_82_CARRYB_3__6_), .CI(u5_mult_82_SUMB_3__7_), .CO(
        u5_mult_82_CARRYB_4__6_), .S(u5_mult_82_SUMB_4__6_) );
  FA_X1 u5_mult_82_S2_4_5 ( .A(u5_mult_82_ab_4__5_), .B(
        u5_mult_82_CARRYB_3__5_), .CI(u5_mult_82_SUMB_3__6_), .CO(
        u5_mult_82_CARRYB_4__5_), .S(u5_mult_82_SUMB_4__5_) );
  FA_X1 u5_mult_82_S2_4_4 ( .A(u5_mult_82_ab_4__4_), .B(
        u5_mult_82_CARRYB_3__4_), .CI(u5_mult_82_SUMB_3__5_), .CO(
        u5_mult_82_CARRYB_4__4_), .S(u5_mult_82_SUMB_4__4_) );
  FA_X1 u5_mult_82_S2_4_3 ( .A(u5_mult_82_ab_4__3_), .B(
        u5_mult_82_CARRYB_3__3_), .CI(u5_mult_82_SUMB_3__4_), .CO(
        u5_mult_82_CARRYB_4__3_), .S(u5_mult_82_SUMB_4__3_) );
  FA_X1 u5_mult_82_S2_4_2 ( .A(u5_mult_82_ab_4__2_), .B(
        u5_mult_82_CARRYB_3__2_), .CI(u5_mult_82_SUMB_3__3_), .CO(
        u5_mult_82_CARRYB_4__2_), .S(u5_mult_82_SUMB_4__2_) );
  FA_X1 u5_mult_82_S2_4_1 ( .A(u5_mult_82_ab_4__1_), .B(
        u5_mult_82_CARRYB_3__1_), .CI(u5_mult_82_SUMB_3__2_), .CO(
        u5_mult_82_CARRYB_4__1_), .S(u5_mult_82_SUMB_4__1_) );
  FA_X1 u5_mult_82_S1_4_0 ( .A(u5_mult_82_ab_4__0_), .B(
        u5_mult_82_CARRYB_3__0_), .CI(u5_mult_82_SUMB_3__1_), .CO(
        u5_mult_82_CARRYB_4__0_), .S(u5_N4) );
  FA_X1 u5_mult_82_S2_5_48 ( .A(u5_mult_82_SUMB_4__49_), .B(
        u5_mult_82_ab_5__48_), .CI(u5_mult_82_CARRYB_4__48_), .CO(
        u5_mult_82_CARRYB_5__48_), .S(u5_mult_82_SUMB_5__48_) );
  FA_X1 u5_mult_82_S2_5_46 ( .A(u5_mult_82_ab_5__46_), .B(
        u5_mult_82_CARRYB_4__46_), .CI(u5_mult_82_SUMB_4__47_), .CO(
        u5_mult_82_CARRYB_5__46_), .S(u5_mult_82_SUMB_5__46_) );
  FA_X1 u5_mult_82_S2_5_43 ( .A(u5_mult_82_ab_5__43_), .B(
        u5_mult_82_CARRYB_4__43_), .CI(u5_mult_82_SUMB_4__44_), .CO(
        u5_mult_82_CARRYB_5__43_), .S(u5_mult_82_SUMB_5__43_) );
  FA_X1 u5_mult_82_S2_5_42 ( .A(u5_mult_82_ab_5__42_), .B(
        u5_mult_82_CARRYB_4__42_), .CI(u5_mult_82_SUMB_4__43_), .CO(
        u5_mult_82_CARRYB_5__42_), .S(u5_mult_82_SUMB_5__42_) );
  FA_X1 u5_mult_82_S2_5_39 ( .A(u5_mult_82_ab_5__39_), .B(
        u5_mult_82_CARRYB_4__39_), .CI(u5_mult_82_SUMB_4__40_), .CO(
        u5_mult_82_CARRYB_5__39_), .S(u5_mult_82_SUMB_5__39_) );
  FA_X1 u5_mult_82_S2_5_33 ( .A(u5_mult_82_ab_5__33_), .B(
        u5_mult_82_CARRYB_4__33_), .CI(u5_mult_82_SUMB_4__34_), .CO(
        u5_mult_82_CARRYB_5__33_), .S(u5_mult_82_SUMB_5__33_) );
  FA_X1 u5_mult_82_S2_5_32 ( .A(u5_mult_82_ab_5__32_), .B(
        u5_mult_82_CARRYB_4__32_), .CI(u5_mult_82_SUMB_4__33_), .CO(
        u5_mult_82_CARRYB_5__32_), .S(u5_mult_82_SUMB_5__32_) );
  FA_X1 u5_mult_82_S2_5_31 ( .A(u5_mult_82_ab_5__31_), .B(
        u5_mult_82_CARRYB_4__31_), .CI(u5_mult_82_SUMB_4__32_), .CO(
        u5_mult_82_CARRYB_5__31_), .S(u5_mult_82_SUMB_5__31_) );
  FA_X1 u5_mult_82_S2_5_26 ( .A(u5_mult_82_ab_5__26_), .B(
        u5_mult_82_CARRYB_4__26_), .CI(u5_mult_82_SUMB_4__27_), .CO(
        u5_mult_82_CARRYB_5__26_), .S(u5_mult_82_SUMB_5__26_) );
  FA_X1 u5_mult_82_S2_5_24 ( .A(u5_mult_82_CARRYB_4__24_), .B(
        u5_mult_82_ab_5__24_), .CI(u5_mult_82_SUMB_4__25_), .CO(
        u5_mult_82_CARRYB_5__24_), .S(u5_mult_82_SUMB_5__24_) );
  FA_X1 u5_mult_82_S2_5_23 ( .A(u5_mult_82_ab_5__23_), .B(
        u5_mult_82_CARRYB_4__23_), .CI(u5_mult_82_SUMB_4__24_), .CO(
        u5_mult_82_CARRYB_5__23_), .S(u5_mult_82_SUMB_5__23_) );
  FA_X1 u5_mult_82_S2_5_20 ( .A(u5_mult_82_ab_5__20_), .B(
        u5_mult_82_CARRYB_4__20_), .CI(u5_mult_82_SUMB_4__21_), .CO(
        u5_mult_82_CARRYB_5__20_), .S(u5_mult_82_SUMB_5__20_) );
  FA_X1 u5_mult_82_S2_5_18 ( .A(u5_mult_82_ab_5__18_), .B(
        u5_mult_82_CARRYB_4__18_), .CI(u5_mult_82_SUMB_4__19_), .CO(
        u5_mult_82_CARRYB_5__18_), .S(u5_mult_82_SUMB_5__18_) );
  FA_X1 u5_mult_82_S2_5_17 ( .A(u5_mult_82_ab_5__17_), .B(
        u5_mult_82_CARRYB_4__17_), .CI(u5_mult_82_SUMB_4__18_), .CO(
        u5_mult_82_CARRYB_5__17_), .S(u5_mult_82_SUMB_5__17_) );
  FA_X1 u5_mult_82_S2_5_16 ( .A(u5_mult_82_ab_5__16_), .B(
        u5_mult_82_CARRYB_4__16_), .CI(u5_mult_82_SUMB_4__17_), .CO(
        u5_mult_82_CARRYB_5__16_), .S(u5_mult_82_SUMB_5__16_) );
  FA_X1 u5_mult_82_S2_5_15 ( .A(u5_mult_82_ab_5__15_), .B(
        u5_mult_82_CARRYB_4__15_), .CI(u5_mult_82_SUMB_4__16_), .CO(
        u5_mult_82_CARRYB_5__15_), .S(u5_mult_82_SUMB_5__15_) );
  FA_X1 u5_mult_82_S2_5_14 ( .A(u5_mult_82_ab_5__14_), .B(
        u5_mult_82_CARRYB_4__14_), .CI(u5_mult_82_SUMB_4__15_), .CO(
        u5_mult_82_CARRYB_5__14_), .S(u5_mult_82_SUMB_5__14_) );
  FA_X1 u5_mult_82_S2_5_13 ( .A(u5_mult_82_ab_5__13_), .B(
        u5_mult_82_CARRYB_4__13_), .CI(u5_mult_82_SUMB_4__14_), .CO(
        u5_mult_82_CARRYB_5__13_), .S(u5_mult_82_SUMB_5__13_) );
  FA_X1 u5_mult_82_S2_5_12 ( .A(u5_mult_82_ab_5__12_), .B(
        u5_mult_82_CARRYB_4__12_), .CI(u5_mult_82_SUMB_4__13_), .CO(
        u5_mult_82_CARRYB_5__12_), .S(u5_mult_82_SUMB_5__12_) );
  FA_X1 u5_mult_82_S2_5_11 ( .A(u5_mult_82_ab_5__11_), .B(
        u5_mult_82_CARRYB_4__11_), .CI(u5_mult_82_SUMB_4__12_), .CO(
        u5_mult_82_CARRYB_5__11_), .S(u5_mult_82_SUMB_5__11_) );
  FA_X1 u5_mult_82_S2_5_10 ( .A(u5_mult_82_ab_5__10_), .B(
        u5_mult_82_CARRYB_4__10_), .CI(u5_mult_82_SUMB_4__11_), .CO(
        u5_mult_82_CARRYB_5__10_), .S(u5_mult_82_SUMB_5__10_) );
  FA_X1 u5_mult_82_S2_5_9 ( .A(u5_mult_82_ab_5__9_), .B(
        u5_mult_82_CARRYB_4__9_), .CI(u5_mult_82_SUMB_4__10_), .CO(
        u5_mult_82_CARRYB_5__9_), .S(u5_mult_82_SUMB_5__9_) );
  FA_X1 u5_mult_82_S2_5_8 ( .A(u5_mult_82_ab_5__8_), .B(
        u5_mult_82_CARRYB_4__8_), .CI(u5_mult_82_SUMB_4__9_), .CO(
        u5_mult_82_CARRYB_5__8_), .S(u5_mult_82_SUMB_5__8_) );
  FA_X1 u5_mult_82_S2_5_7 ( .A(u5_mult_82_ab_5__7_), .B(
        u5_mult_82_CARRYB_4__7_), .CI(u5_mult_82_SUMB_4__8_), .CO(
        u5_mult_82_CARRYB_5__7_), .S(u5_mult_82_SUMB_5__7_) );
  FA_X1 u5_mult_82_S2_5_6 ( .A(u5_mult_82_ab_5__6_), .B(
        u5_mult_82_CARRYB_4__6_), .CI(u5_mult_82_SUMB_4__7_), .CO(
        u5_mult_82_CARRYB_5__6_), .S(u5_mult_82_SUMB_5__6_) );
  FA_X1 u5_mult_82_S2_5_5 ( .A(u5_mult_82_ab_5__5_), .B(
        u5_mult_82_CARRYB_4__5_), .CI(u5_mult_82_SUMB_4__6_), .CO(
        u5_mult_82_CARRYB_5__5_), .S(u5_mult_82_SUMB_5__5_) );
  FA_X1 u5_mult_82_S2_5_4 ( .A(u5_mult_82_ab_5__4_), .B(
        u5_mult_82_CARRYB_4__4_), .CI(u5_mult_82_SUMB_4__5_), .CO(
        u5_mult_82_CARRYB_5__4_), .S(u5_mult_82_SUMB_5__4_) );
  FA_X1 u5_mult_82_S2_5_3 ( .A(u5_mult_82_ab_5__3_), .B(
        u5_mult_82_CARRYB_4__3_), .CI(u5_mult_82_SUMB_4__4_), .CO(
        u5_mult_82_CARRYB_5__3_), .S(u5_mult_82_SUMB_5__3_) );
  FA_X1 u5_mult_82_S2_5_2 ( .A(u5_mult_82_ab_5__2_), .B(
        u5_mult_82_CARRYB_4__2_), .CI(u5_mult_82_SUMB_4__3_), .CO(
        u5_mult_82_CARRYB_5__2_), .S(u5_mult_82_SUMB_5__2_) );
  FA_X1 u5_mult_82_S2_5_1 ( .A(u5_mult_82_ab_5__1_), .B(
        u5_mult_82_CARRYB_4__1_), .CI(u5_mult_82_SUMB_4__2_), .CO(
        u5_mult_82_CARRYB_5__1_), .S(u5_mult_82_SUMB_5__1_) );
  FA_X1 u5_mult_82_S1_5_0 ( .A(u5_mult_82_ab_5__0_), .B(
        u5_mult_82_CARRYB_4__0_), .CI(u5_mult_82_SUMB_4__1_), .CO(
        u5_mult_82_CARRYB_5__0_), .S(u5_N5) );
  FA_X1 u5_mult_82_S3_6_51 ( .A(u5_mult_82_ab_6__51_), .B(u5_mult_82_ab_5__52_), .CI(u5_mult_82_CARRYB_5__51_), .CO(u5_mult_82_CARRYB_6__51_), .S(
        u5_mult_82_SUMB_6__51_) );
  FA_X1 u5_mult_82_S2_6_49 ( .A(u5_mult_82_ab_6__49_), .B(
        u5_mult_82_CARRYB_5__49_), .CI(u5_mult_82_SUMB_5__50_), .CO(
        u5_mult_82_CARRYB_6__49_), .S(u5_mult_82_SUMB_6__49_) );
  FA_X1 u5_mult_82_S2_6_41 ( .A(u5_mult_82_ab_6__41_), .B(
        u5_mult_82_CARRYB_5__41_), .CI(u5_mult_82_SUMB_5__42_), .CO(
        u5_mult_82_CARRYB_6__41_), .S(u5_mult_82_SUMB_6__41_) );
  FA_X1 u5_mult_82_S2_6_31 ( .A(u5_mult_82_ab_6__31_), .B(
        u5_mult_82_CARRYB_5__31_), .CI(u5_mult_82_SUMB_5__32_), .CO(
        u5_mult_82_CARRYB_6__31_), .S(u5_mult_82_SUMB_6__31_) );
  FA_X1 u5_mult_82_S2_6_27 ( .A(u5_mult_82_CARRYB_5__27_), .B(
        u5_mult_82_ab_6__27_), .CI(u5_mult_82_SUMB_5__28_), .CO(
        u5_mult_82_CARRYB_6__27_), .S(u5_mult_82_SUMB_6__27_) );
  FA_X1 u5_mult_82_S2_6_24 ( .A(u5_mult_82_ab_6__24_), .B(
        u5_mult_82_CARRYB_5__24_), .CI(u5_mult_82_SUMB_5__25_), .CO(
        u5_mult_82_CARRYB_6__24_), .S(u5_mult_82_SUMB_6__24_) );
  FA_X1 u5_mult_82_S2_6_23 ( .A(u5_mult_82_ab_6__23_), .B(
        u5_mult_82_CARRYB_5__23_), .CI(u5_mult_82_SUMB_5__24_), .CO(
        u5_mult_82_CARRYB_6__23_), .S(u5_mult_82_SUMB_6__23_) );
  FA_X1 u5_mult_82_S2_6_22 ( .A(u5_mult_82_ab_6__22_), .B(
        u5_mult_82_CARRYB_5__22_), .CI(u5_mult_82_SUMB_5__23_), .CO(
        u5_mult_82_CARRYB_6__22_), .S(u5_mult_82_SUMB_6__22_) );
  FA_X1 u5_mult_82_S2_6_21 ( .A(u5_mult_82_ab_6__21_), .B(
        u5_mult_82_CARRYB_5__21_), .CI(u5_mult_82_SUMB_5__22_), .CO(
        u5_mult_82_CARRYB_6__21_), .S(u5_mult_82_SUMB_6__21_) );
  FA_X1 u5_mult_82_S2_6_19 ( .A(u5_mult_82_ab_6__19_), .B(
        u5_mult_82_CARRYB_5__19_), .CI(u5_mult_82_SUMB_5__20_), .CO(
        u5_mult_82_CARRYB_6__19_), .S(u5_mult_82_SUMB_6__19_) );
  FA_X1 u5_mult_82_S2_6_17 ( .A(u5_mult_82_ab_6__17_), .B(
        u5_mult_82_CARRYB_5__17_), .CI(u5_mult_82_SUMB_5__18_), .CO(
        u5_mult_82_CARRYB_6__17_), .S(u5_mult_82_SUMB_6__17_) );
  FA_X1 u5_mult_82_S2_6_15 ( .A(u5_mult_82_ab_6__15_), .B(
        u5_mult_82_CARRYB_5__15_), .CI(u5_mult_82_SUMB_5__16_), .CO(
        u5_mult_82_CARRYB_6__15_), .S(u5_mult_82_SUMB_6__15_) );
  FA_X1 u5_mult_82_S2_6_14 ( .A(u5_mult_82_ab_6__14_), .B(
        u5_mult_82_CARRYB_5__14_), .CI(u5_mult_82_SUMB_5__15_), .CO(
        u5_mult_82_CARRYB_6__14_), .S(u5_mult_82_SUMB_6__14_) );
  FA_X1 u5_mult_82_S2_6_13 ( .A(u5_mult_82_ab_6__13_), .B(
        u5_mult_82_CARRYB_5__13_), .CI(u5_mult_82_SUMB_5__14_), .CO(
        u5_mult_82_CARRYB_6__13_), .S(u5_mult_82_SUMB_6__13_) );
  FA_X1 u5_mult_82_S2_6_12 ( .A(u5_mult_82_ab_6__12_), .B(
        u5_mult_82_CARRYB_5__12_), .CI(u5_mult_82_SUMB_5__13_), .CO(
        u5_mult_82_CARRYB_6__12_), .S(u5_mult_82_SUMB_6__12_) );
  FA_X1 u5_mult_82_S2_6_11 ( .A(u5_mult_82_ab_6__11_), .B(
        u5_mult_82_CARRYB_5__11_), .CI(u5_mult_82_SUMB_5__12_), .CO(
        u5_mult_82_CARRYB_6__11_), .S(u5_mult_82_SUMB_6__11_) );
  FA_X1 u5_mult_82_S2_6_10 ( .A(u5_mult_82_ab_6__10_), .B(
        u5_mult_82_CARRYB_5__10_), .CI(u5_mult_82_SUMB_5__11_), .CO(
        u5_mult_82_CARRYB_6__10_), .S(u5_mult_82_SUMB_6__10_) );
  FA_X1 u5_mult_82_S2_6_9 ( .A(u5_mult_82_ab_6__9_), .B(
        u5_mult_82_CARRYB_5__9_), .CI(u5_mult_82_SUMB_5__10_), .CO(
        u5_mult_82_CARRYB_6__9_), .S(u5_mult_82_SUMB_6__9_) );
  FA_X1 u5_mult_82_S2_6_8 ( .A(u5_mult_82_ab_6__8_), .B(
        u5_mult_82_CARRYB_5__8_), .CI(u5_mult_82_SUMB_5__9_), .CO(
        u5_mult_82_CARRYB_6__8_), .S(u5_mult_82_SUMB_6__8_) );
  FA_X1 u5_mult_82_S2_6_7 ( .A(u5_mult_82_ab_6__7_), .B(
        u5_mult_82_CARRYB_5__7_), .CI(u5_mult_82_SUMB_5__8_), .CO(
        u5_mult_82_CARRYB_6__7_), .S(u5_mult_82_SUMB_6__7_) );
  FA_X1 u5_mult_82_S2_6_6 ( .A(u5_mult_82_ab_6__6_), .B(
        u5_mult_82_CARRYB_5__6_), .CI(u5_mult_82_SUMB_5__7_), .CO(
        u5_mult_82_CARRYB_6__6_), .S(u5_mult_82_SUMB_6__6_) );
  FA_X1 u5_mult_82_S2_6_5 ( .A(u5_mult_82_ab_6__5_), .B(
        u5_mult_82_CARRYB_5__5_), .CI(u5_mult_82_SUMB_5__6_), .CO(
        u5_mult_82_CARRYB_6__5_), .S(u5_mult_82_SUMB_6__5_) );
  FA_X1 u5_mult_82_S2_6_4 ( .A(u5_mult_82_ab_6__4_), .B(
        u5_mult_82_CARRYB_5__4_), .CI(u5_mult_82_SUMB_5__5_), .CO(
        u5_mult_82_CARRYB_6__4_), .S(u5_mult_82_SUMB_6__4_) );
  FA_X1 u5_mult_82_S2_6_3 ( .A(u5_mult_82_ab_6__3_), .B(
        u5_mult_82_CARRYB_5__3_), .CI(u5_mult_82_SUMB_5__4_), .CO(
        u5_mult_82_CARRYB_6__3_), .S(u5_mult_82_SUMB_6__3_) );
  FA_X1 u5_mult_82_S2_6_2 ( .A(u5_mult_82_ab_6__2_), .B(
        u5_mult_82_CARRYB_5__2_), .CI(u5_mult_82_SUMB_5__3_), .CO(
        u5_mult_82_CARRYB_6__2_), .S(u5_mult_82_SUMB_6__2_) );
  FA_X1 u5_mult_82_S2_6_1 ( .A(u5_mult_82_ab_6__1_), .B(
        u5_mult_82_CARRYB_5__1_), .CI(u5_mult_82_SUMB_5__2_), .CO(
        u5_mult_82_CARRYB_6__1_), .S(u5_mult_82_SUMB_6__1_) );
  FA_X1 u5_mult_82_S1_6_0 ( .A(u5_mult_82_ab_6__0_), .B(
        u5_mult_82_CARRYB_5__0_), .CI(u5_mult_82_SUMB_5__1_), .CO(
        u5_mult_82_CARRYB_6__0_), .S(u5_N6) );
  FA_X1 u5_mult_82_S3_7_51 ( .A(u5_mult_82_ab_7__51_), .B(u5_mult_82_ab_6__52_), .CI(u5_mult_82_CARRYB_6__51_), .CO(u5_mult_82_CARRYB_7__51_), .S(
        u5_mult_82_SUMB_7__51_) );
  FA_X1 u5_mult_82_S2_7_50 ( .A(u5_mult_82_ab_7__50_), .B(
        u5_mult_82_CARRYB_6__50_), .CI(u5_mult_82_SUMB_6__51_), .CO(
        u5_mult_82_CARRYB_7__50_), .S(u5_mult_82_SUMB_7__50_) );
  FA_X1 u5_mult_82_S2_7_47 ( .A(u5_mult_82_CARRYB_6__47_), .B(
        u5_mult_82_ab_7__47_), .CI(u5_mult_82_SUMB_6__48_), .CO(
        u5_mult_82_CARRYB_7__47_), .S(u5_mult_82_SUMB_7__47_) );
  FA_X1 u5_mult_82_S2_7_45 ( .A(u5_mult_82_ab_7__45_), .B(
        u5_mult_82_CARRYB_6__45_), .CI(u5_mult_82_SUMB_6__46_), .CO(
        u5_mult_82_CARRYB_7__45_), .S(u5_mult_82_SUMB_7__45_) );
  FA_X1 u5_mult_82_S2_7_32 ( .A(u5_mult_82_ab_7__32_), .B(
        u5_mult_82_CARRYB_6__32_), .CI(u5_mult_82_SUMB_6__33_), .CO(
        u5_mult_82_CARRYB_7__32_), .S(u5_mult_82_SUMB_7__32_) );
  FA_X1 u5_mult_82_S2_7_29 ( .A(u5_mult_82_ab_7__29_), .B(
        u5_mult_82_CARRYB_6__29_), .CI(u5_mult_82_SUMB_6__30_), .CO(
        u5_mult_82_CARRYB_7__29_), .S(u5_mult_82_SUMB_7__29_) );
  FA_X1 u5_mult_82_S2_7_23 ( .A(u5_mult_82_CARRYB_6__23_), .B(
        u5_mult_82_ab_7__23_), .CI(u5_mult_82_SUMB_6__24_), .CO(
        u5_mult_82_CARRYB_7__23_), .S(u5_mult_82_SUMB_7__23_) );
  FA_X1 u5_mult_82_S2_7_22 ( .A(u5_mult_82_CARRYB_6__22_), .B(
        u5_mult_82_ab_7__22_), .CI(u5_mult_82_SUMB_6__23_), .CO(
        u5_mult_82_CARRYB_7__22_), .S(u5_mult_82_SUMB_7__22_) );
  FA_X1 u5_mult_82_S2_7_21 ( .A(u5_mult_82_ab_7__21_), .B(
        u5_mult_82_CARRYB_6__21_), .CI(u5_mult_82_SUMB_6__22_), .CO(
        u5_mult_82_CARRYB_7__21_), .S(u5_mult_82_SUMB_7__21_) );
  FA_X1 u5_mult_82_S2_7_20 ( .A(u5_mult_82_ab_7__20_), .B(
        u5_mult_82_CARRYB_6__20_), .CI(u5_mult_82_SUMB_6__21_), .CO(
        u5_mult_82_CARRYB_7__20_), .S(u5_mult_82_SUMB_7__20_) );
  FA_X1 u5_mult_82_S2_7_18 ( .A(u5_mult_82_ab_7__18_), .B(
        u5_mult_82_CARRYB_6__18_), .CI(u5_mult_82_SUMB_6__19_), .CO(
        u5_mult_82_CARRYB_7__18_), .S(u5_mult_82_SUMB_7__18_) );
  FA_X1 u5_mult_82_S2_7_17 ( .A(u5_mult_82_ab_7__17_), .B(
        u5_mult_82_CARRYB_6__17_), .CI(u5_mult_82_SUMB_6__18_), .CO(
        u5_mult_82_CARRYB_7__17_), .S(u5_mult_82_SUMB_7__17_) );
  FA_X1 u5_mult_82_S2_7_16 ( .A(u5_mult_82_ab_7__16_), .B(
        u5_mult_82_CARRYB_6__16_), .CI(u5_mult_82_SUMB_6__17_), .CO(
        u5_mult_82_CARRYB_7__16_), .S(u5_mult_82_SUMB_7__16_) );
  FA_X1 u5_mult_82_S2_7_14 ( .A(u5_mult_82_ab_7__14_), .B(
        u5_mult_82_CARRYB_6__14_), .CI(u5_mult_82_SUMB_6__15_), .CO(
        u5_mult_82_CARRYB_7__14_), .S(u5_mult_82_SUMB_7__14_) );
  FA_X1 u5_mult_82_S2_7_13 ( .A(u5_mult_82_ab_7__13_), .B(
        u5_mult_82_CARRYB_6__13_), .CI(u5_mult_82_SUMB_6__14_), .CO(
        u5_mult_82_CARRYB_7__13_), .S(u5_mult_82_SUMB_7__13_) );
  FA_X1 u5_mult_82_S2_7_12 ( .A(u5_mult_82_ab_7__12_), .B(
        u5_mult_82_CARRYB_6__12_), .CI(u5_mult_82_SUMB_6__13_), .CO(
        u5_mult_82_CARRYB_7__12_), .S(u5_mult_82_SUMB_7__12_) );
  FA_X1 u5_mult_82_S2_7_11 ( .A(u5_mult_82_ab_7__11_), .B(
        u5_mult_82_CARRYB_6__11_), .CI(u5_mult_82_SUMB_6__12_), .CO(
        u5_mult_82_CARRYB_7__11_), .S(u5_mult_82_SUMB_7__11_) );
  FA_X1 u5_mult_82_S2_7_10 ( .A(u5_mult_82_ab_7__10_), .B(
        u5_mult_82_CARRYB_6__10_), .CI(u5_mult_82_SUMB_6__11_), .CO(
        u5_mult_82_CARRYB_7__10_), .S(u5_mult_82_SUMB_7__10_) );
  FA_X1 u5_mult_82_S2_7_9 ( .A(u5_mult_82_ab_7__9_), .B(
        u5_mult_82_CARRYB_6__9_), .CI(u5_mult_82_SUMB_6__10_), .CO(
        u5_mult_82_CARRYB_7__9_), .S(u5_mult_82_SUMB_7__9_) );
  FA_X1 u5_mult_82_S2_7_8 ( .A(u5_mult_82_ab_7__8_), .B(
        u5_mult_82_CARRYB_6__8_), .CI(u5_mult_82_SUMB_6__9_), .CO(
        u5_mult_82_CARRYB_7__8_), .S(u5_mult_82_SUMB_7__8_) );
  FA_X1 u5_mult_82_S2_7_7 ( .A(u5_mult_82_ab_7__7_), .B(
        u5_mult_82_CARRYB_6__7_), .CI(u5_mult_82_SUMB_6__8_), .CO(
        u5_mult_82_CARRYB_7__7_), .S(u5_mult_82_SUMB_7__7_) );
  FA_X1 u5_mult_82_S2_7_6 ( .A(u5_mult_82_ab_7__6_), .B(
        u5_mult_82_CARRYB_6__6_), .CI(u5_mult_82_SUMB_6__7_), .CO(
        u5_mult_82_CARRYB_7__6_), .S(u5_mult_82_SUMB_7__6_) );
  FA_X1 u5_mult_82_S2_7_5 ( .A(u5_mult_82_ab_7__5_), .B(
        u5_mult_82_CARRYB_6__5_), .CI(u5_mult_82_SUMB_6__6_), .CO(
        u5_mult_82_CARRYB_7__5_), .S(u5_mult_82_SUMB_7__5_) );
  FA_X1 u5_mult_82_S2_7_4 ( .A(u5_mult_82_ab_7__4_), .B(
        u5_mult_82_CARRYB_6__4_), .CI(u5_mult_82_SUMB_6__5_), .CO(
        u5_mult_82_CARRYB_7__4_), .S(u5_mult_82_SUMB_7__4_) );
  FA_X1 u5_mult_82_S2_7_3 ( .A(u5_mult_82_ab_7__3_), .B(
        u5_mult_82_CARRYB_6__3_), .CI(u5_mult_82_SUMB_6__4_), .CO(
        u5_mult_82_CARRYB_7__3_), .S(u5_mult_82_SUMB_7__3_) );
  FA_X1 u5_mult_82_S2_7_2 ( .A(u5_mult_82_ab_7__2_), .B(
        u5_mult_82_CARRYB_6__2_), .CI(u5_mult_82_SUMB_6__3_), .CO(
        u5_mult_82_CARRYB_7__2_), .S(u5_mult_82_SUMB_7__2_) );
  FA_X1 u5_mult_82_S2_7_1 ( .A(u5_mult_82_ab_7__1_), .B(
        u5_mult_82_CARRYB_6__1_), .CI(u5_mult_82_SUMB_6__2_), .CO(
        u5_mult_82_CARRYB_7__1_), .S(u5_mult_82_SUMB_7__1_) );
  FA_X1 u5_mult_82_S1_7_0 ( .A(u5_mult_82_ab_7__0_), .B(
        u5_mult_82_CARRYB_6__0_), .CI(u5_mult_82_SUMB_6__1_), .CO(
        u5_mult_82_CARRYB_7__0_), .S(u5_N7) );
  FA_X1 u5_mult_82_S3_8_51 ( .A(u5_mult_82_ab_8__51_), .B(
        u5_mult_82_CARRYB_7__51_), .CI(u5_mult_82_ab_7__52_), .CO(
        u5_mult_82_CARRYB_8__51_), .S(u5_mult_82_SUMB_8__51_) );
  FA_X1 u5_mult_82_S2_8_50 ( .A(u5_mult_82_ab_8__50_), .B(
        u5_mult_82_CARRYB_7__50_), .CI(u5_mult_82_SUMB_7__51_), .CO(
        u5_mult_82_CARRYB_8__50_), .S(u5_mult_82_SUMB_8__50_) );
  FA_X1 u5_mult_82_S2_8_49 ( .A(u5_mult_82_ab_8__49_), .B(
        u5_mult_82_CARRYB_7__49_), .CI(u5_mult_82_SUMB_7__50_), .CO(
        u5_mult_82_CARRYB_8__49_), .S(u5_mult_82_SUMB_8__49_) );
  FA_X1 u5_mult_82_S2_8_46 ( .A(u5_mult_82_ab_8__46_), .B(
        u5_mult_82_CARRYB_7__46_), .CI(u5_mult_82_SUMB_7__47_), .CO(
        u5_mult_82_CARRYB_8__46_), .S(u5_mult_82_SUMB_8__46_) );
  FA_X1 u5_mult_82_S2_8_43 ( .A(u5_mult_82_ab_8__43_), .B(
        u5_mult_82_CARRYB_7__43_), .CI(u5_mult_82_SUMB_7__44_), .CO(
        u5_mult_82_CARRYB_8__43_), .S(u5_mult_82_SUMB_8__43_) );
  FA_X1 u5_mult_82_S2_8_39 ( .A(u5_mult_82_ab_8__39_), .B(
        u5_mult_82_CARRYB_7__39_), .CI(u5_mult_82_SUMB_7__40_), .CO(
        u5_mult_82_CARRYB_8__39_), .S(u5_mult_82_SUMB_8__39_) );
  FA_X1 u5_mult_82_S2_8_37 ( .A(u5_mult_82_ab_8__37_), .B(
        u5_mult_82_CARRYB_7__37_), .CI(u5_mult_82_SUMB_7__38_), .CO(
        u5_mult_82_CARRYB_8__37_), .S(u5_mult_82_SUMB_8__37_) );
  FA_X1 u5_mult_82_S2_8_32 ( .A(u5_mult_82_CARRYB_7__32_), .B(
        u5_mult_82_ab_8__32_), .CI(u5_mult_82_SUMB_7__33_), .CO(
        u5_mult_82_CARRYB_8__32_), .S(u5_mult_82_SUMB_8__32_) );
  FA_X1 u5_mult_82_S2_8_31 ( .A(u5_mult_82_ab_8__31_), .B(
        u5_mult_82_CARRYB_7__31_), .CI(u5_mult_82_SUMB_7__32_), .CO(
        u5_mult_82_CARRYB_8__31_), .S(u5_mult_82_SUMB_8__31_) );
  FA_X1 u5_mult_82_S2_8_26 ( .A(u5_mult_82_CARRYB_7__26_), .B(
        u5_mult_82_ab_8__26_), .CI(u5_mult_82_SUMB_7__27_), .CO(
        u5_mult_82_CARRYB_8__26_), .S(u5_mult_82_SUMB_8__26_) );
  FA_X1 u5_mult_82_S2_8_23 ( .A(u5_mult_82_ab_8__23_), .B(
        u5_mult_82_CARRYB_7__23_), .CI(u5_mult_82_SUMB_7__24_), .CO(
        u5_mult_82_CARRYB_8__23_), .S(u5_mult_82_SUMB_8__23_) );
  FA_X1 u5_mult_82_S2_8_21 ( .A(u5_mult_82_ab_8__21_), .B(
        u5_mult_82_CARRYB_7__21_), .CI(u5_mult_82_SUMB_7__22_), .CO(
        u5_mult_82_CARRYB_8__21_), .S(u5_mult_82_SUMB_8__21_) );
  FA_X1 u5_mult_82_S2_8_20 ( .A(u5_mult_82_ab_8__20_), .B(
        u5_mult_82_CARRYB_7__20_), .CI(u5_mult_82_SUMB_7__21_), .CO(
        u5_mult_82_CARRYB_8__20_), .S(u5_mult_82_SUMB_8__20_) );
  FA_X1 u5_mult_82_S2_8_18 ( .A(u5_mult_82_ab_8__18_), .B(
        u5_mult_82_CARRYB_7__18_), .CI(u5_mult_82_SUMB_7__19_), .CO(
        u5_mult_82_CARRYB_8__18_), .S(u5_mult_82_SUMB_8__18_) );
  FA_X1 u5_mult_82_S2_8_16 ( .A(u5_mult_82_ab_8__16_), .B(
        u5_mult_82_CARRYB_7__16_), .CI(u5_mult_82_SUMB_7__17_), .CO(
        u5_mult_82_CARRYB_8__16_), .S(u5_mult_82_SUMB_8__16_) );
  FA_X1 u5_mult_82_S2_8_15 ( .A(u5_mult_82_ab_8__15_), .B(
        u5_mult_82_CARRYB_7__15_), .CI(u5_mult_82_SUMB_7__16_), .CO(
        u5_mult_82_CARRYB_8__15_), .S(u5_mult_82_SUMB_8__15_) );
  FA_X1 u5_mult_82_S2_8_14 ( .A(u5_mult_82_ab_8__14_), .B(
        u5_mult_82_CARRYB_7__14_), .CI(u5_mult_82_SUMB_7__15_), .CO(
        u5_mult_82_CARRYB_8__14_), .S(u5_mult_82_SUMB_8__14_) );
  FA_X1 u5_mult_82_S2_8_13 ( .A(u5_mult_82_ab_8__13_), .B(
        u5_mult_82_CARRYB_7__13_), .CI(u5_mult_82_SUMB_7__14_), .CO(
        u5_mult_82_CARRYB_8__13_), .S(u5_mult_82_SUMB_8__13_) );
  FA_X1 u5_mult_82_S2_8_12 ( .A(u5_mult_82_ab_8__12_), .B(
        u5_mult_82_CARRYB_7__12_), .CI(u5_mult_82_SUMB_7__13_), .CO(
        u5_mult_82_CARRYB_8__12_), .S(u5_mult_82_SUMB_8__12_) );
  FA_X1 u5_mult_82_S2_8_11 ( .A(u5_mult_82_ab_8__11_), .B(
        u5_mult_82_CARRYB_7__11_), .CI(u5_mult_82_SUMB_7__12_), .CO(
        u5_mult_82_CARRYB_8__11_), .S(u5_mult_82_SUMB_8__11_) );
  FA_X1 u5_mult_82_S2_8_10 ( .A(u5_mult_82_ab_8__10_), .B(
        u5_mult_82_CARRYB_7__10_), .CI(u5_mult_82_SUMB_7__11_), .CO(
        u5_mult_82_CARRYB_8__10_), .S(u5_mult_82_SUMB_8__10_) );
  FA_X1 u5_mult_82_S2_8_9 ( .A(u5_mult_82_ab_8__9_), .B(
        u5_mult_82_CARRYB_7__9_), .CI(u5_mult_82_SUMB_7__10_), .CO(
        u5_mult_82_CARRYB_8__9_), .S(u5_mult_82_SUMB_8__9_) );
  FA_X1 u5_mult_82_S2_8_8 ( .A(u5_mult_82_ab_8__8_), .B(
        u5_mult_82_CARRYB_7__8_), .CI(u5_mult_82_SUMB_7__9_), .CO(
        u5_mult_82_CARRYB_8__8_), .S(u5_mult_82_SUMB_8__8_) );
  FA_X1 u5_mult_82_S2_8_7 ( .A(u5_mult_82_ab_8__7_), .B(
        u5_mult_82_CARRYB_7__7_), .CI(u5_mult_82_SUMB_7__8_), .CO(
        u5_mult_82_CARRYB_8__7_), .S(u5_mult_82_SUMB_8__7_) );
  FA_X1 u5_mult_82_S2_8_6 ( .A(u5_mult_82_ab_8__6_), .B(
        u5_mult_82_CARRYB_7__6_), .CI(u5_mult_82_SUMB_7__7_), .CO(
        u5_mult_82_CARRYB_8__6_), .S(u5_mult_82_SUMB_8__6_) );
  FA_X1 u5_mult_82_S2_8_5 ( .A(u5_mult_82_ab_8__5_), .B(
        u5_mult_82_CARRYB_7__5_), .CI(u5_mult_82_SUMB_7__6_), .CO(
        u5_mult_82_CARRYB_8__5_), .S(u5_mult_82_SUMB_8__5_) );
  FA_X1 u5_mult_82_S2_8_4 ( .A(u5_mult_82_ab_8__4_), .B(
        u5_mult_82_CARRYB_7__4_), .CI(u5_mult_82_SUMB_7__5_), .CO(
        u5_mult_82_CARRYB_8__4_), .S(u5_mult_82_SUMB_8__4_) );
  FA_X1 u5_mult_82_S2_8_3 ( .A(u5_mult_82_ab_8__3_), .B(
        u5_mult_82_CARRYB_7__3_), .CI(u5_mult_82_SUMB_7__4_), .CO(
        u5_mult_82_CARRYB_8__3_), .S(u5_mult_82_SUMB_8__3_) );
  FA_X1 u5_mult_82_S2_8_2 ( .A(u5_mult_82_ab_8__2_), .B(
        u5_mult_82_CARRYB_7__2_), .CI(u5_mult_82_SUMB_7__3_), .CO(
        u5_mult_82_CARRYB_8__2_), .S(u5_mult_82_SUMB_8__2_) );
  FA_X1 u5_mult_82_S2_8_1 ( .A(u5_mult_82_ab_8__1_), .B(
        u5_mult_82_CARRYB_7__1_), .CI(u5_mult_82_SUMB_7__2_), .CO(
        u5_mult_82_CARRYB_8__1_), .S(u5_mult_82_SUMB_8__1_) );
  FA_X1 u5_mult_82_S1_8_0 ( .A(u5_mult_82_ab_8__0_), .B(
        u5_mult_82_CARRYB_7__0_), .CI(u5_mult_82_SUMB_7__1_), .CO(
        u5_mult_82_CARRYB_8__0_), .S(u5_N8) );
  FA_X1 u5_mult_82_S2_9_50 ( .A(u5_mult_82_ab_9__50_), .B(
        u5_mult_82_CARRYB_8__50_), .CI(u5_mult_82_SUMB_8__51_), .CO(
        u5_mult_82_CARRYB_9__50_), .S(u5_mult_82_SUMB_9__50_) );
  FA_X1 u5_mult_82_S2_9_48 ( .A(u5_mult_82_ab_9__48_), .B(
        u5_mult_82_CARRYB_8__48_), .CI(u5_mult_82_SUMB_8__49_), .CO(
        u5_mult_82_CARRYB_9__48_), .S(u5_mult_82_SUMB_9__48_) );
  FA_X1 u5_mult_82_S2_9_44 ( .A(u5_mult_82_ab_9__44_), .B(
        u5_mult_82_CARRYB_8__44_), .CI(u5_mult_82_SUMB_8__45_), .CO(
        u5_mult_82_CARRYB_9__44_), .S(u5_mult_82_SUMB_9__44_) );
  FA_X1 u5_mult_82_S2_9_43 ( .A(u5_mult_82_ab_9__43_), .B(
        u5_mult_82_CARRYB_8__43_), .CI(u5_mult_82_SUMB_8__44_), .CO(
        u5_mult_82_CARRYB_9__43_), .S(u5_mult_82_SUMB_9__43_) );
  FA_X1 u5_mult_82_S2_9_40 ( .A(u5_mult_82_ab_9__40_), .B(
        u5_mult_82_CARRYB_8__40_), .CI(u5_mult_82_SUMB_8__41_), .CO(
        u5_mult_82_CARRYB_9__40_), .S(u5_mult_82_SUMB_9__40_) );
  FA_X1 u5_mult_82_S2_9_39 ( .A(u5_mult_82_ab_9__39_), .B(
        u5_mult_82_CARRYB_8__39_), .CI(u5_mult_82_SUMB_8__40_), .CO(
        u5_mult_82_CARRYB_9__39_), .S(u5_mult_82_SUMB_9__39_) );
  FA_X1 u5_mult_82_S2_9_37 ( .A(u5_mult_82_CARRYB_8__37_), .B(
        u5_mult_82_ab_9__37_), .CI(u5_mult_82_SUMB_8__38_), .CO(
        u5_mult_82_CARRYB_9__37_), .S(u5_mult_82_SUMB_9__37_) );
  FA_X1 u5_mult_82_S2_9_35 ( .A(u5_mult_82_ab_9__35_), .B(
        u5_mult_82_CARRYB_8__35_), .CI(u5_mult_82_SUMB_8__36_), .CO(
        u5_mult_82_CARRYB_9__35_), .S(u5_mult_82_SUMB_9__35_) );
  FA_X1 u5_mult_82_S2_9_31 ( .A(u5_mult_82_ab_9__31_), .B(
        u5_mult_82_CARRYB_8__31_), .CI(u5_mult_82_SUMB_8__32_), .CO(
        u5_mult_82_CARRYB_9__31_), .S(u5_mult_82_SUMB_9__31_) );
  FA_X1 u5_mult_82_S2_9_27 ( .A(u5_mult_82_ab_9__27_), .B(
        u5_mult_82_CARRYB_8__27_), .CI(u5_mult_82_SUMB_8__28_), .CO(
        u5_mult_82_CARRYB_9__27_), .S(u5_mult_82_SUMB_9__27_) );
  FA_X1 u5_mult_82_S2_9_25 ( .A(u5_mult_82_ab_9__25_), .B(
        u5_mult_82_CARRYB_8__25_), .CI(u5_mult_82_SUMB_8__26_), .CO(
        u5_mult_82_CARRYB_9__25_), .S(u5_mult_82_SUMB_9__25_) );
  FA_X1 u5_mult_82_S2_9_23 ( .A(u5_mult_82_CARRYB_8__23_), .B(
        u5_mult_82_ab_9__23_), .CI(u5_mult_82_SUMB_8__24_), .CO(
        u5_mult_82_CARRYB_9__23_), .S(u5_mult_82_SUMB_9__23_) );
  FA_X1 u5_mult_82_S2_9_22 ( .A(u5_mult_82_ab_9__22_), .B(
        u5_mult_82_CARRYB_8__22_), .CI(u5_mult_82_SUMB_8__23_), .CO(
        u5_mult_82_CARRYB_9__22_), .S(u5_mult_82_SUMB_9__22_) );
  FA_X1 u5_mult_82_S2_9_20 ( .A(u5_mult_82_CARRYB_8__20_), .B(
        u5_mult_82_ab_9__20_), .CI(u5_mult_82_SUMB_8__21_), .CO(
        u5_mult_82_CARRYB_9__20_), .S(u5_mult_82_SUMB_9__20_) );
  FA_X1 u5_mult_82_S2_9_19 ( .A(u5_mult_82_ab_9__19_), .B(
        u5_mult_82_CARRYB_8__19_), .CI(u5_mult_82_SUMB_8__20_), .CO(
        u5_mult_82_CARRYB_9__19_), .S(u5_mult_82_SUMB_9__19_) );
  FA_X1 u5_mult_82_S2_9_17 ( .A(u5_mult_82_ab_9__17_), .B(
        u5_mult_82_CARRYB_8__17_), .CI(u5_mult_82_SUMB_8__18_), .CO(
        u5_mult_82_CARRYB_9__17_), .S(u5_mult_82_SUMB_9__17_) );
  FA_X1 u5_mult_82_S2_9_15 ( .A(u5_mult_82_ab_9__15_), .B(
        u5_mult_82_CARRYB_8__15_), .CI(u5_mult_82_SUMB_8__16_), .CO(
        u5_mult_82_CARRYB_9__15_), .S(u5_mult_82_SUMB_9__15_) );
  FA_X1 u5_mult_82_S2_9_14 ( .A(u5_mult_82_ab_9__14_), .B(
        u5_mult_82_CARRYB_8__14_), .CI(u5_mult_82_SUMB_8__15_), .CO(
        u5_mult_82_CARRYB_9__14_), .S(u5_mult_82_SUMB_9__14_) );
  FA_X1 u5_mult_82_S2_9_13 ( .A(u5_mult_82_ab_9__13_), .B(
        u5_mult_82_CARRYB_8__13_), .CI(u5_mult_82_SUMB_8__14_), .CO(
        u5_mult_82_CARRYB_9__13_), .S(u5_mult_82_SUMB_9__13_) );
  FA_X1 u5_mult_82_S2_9_12 ( .A(u5_mult_82_ab_9__12_), .B(
        u5_mult_82_CARRYB_8__12_), .CI(u5_mult_82_SUMB_8__13_), .CO(
        u5_mult_82_CARRYB_9__12_), .S(u5_mult_82_SUMB_9__12_) );
  FA_X1 u5_mult_82_S2_9_11 ( .A(u5_mult_82_ab_9__11_), .B(
        u5_mult_82_CARRYB_8__11_), .CI(u5_mult_82_SUMB_8__12_), .CO(
        u5_mult_82_CARRYB_9__11_), .S(u5_mult_82_SUMB_9__11_) );
  FA_X1 u5_mult_82_S2_9_10 ( .A(u5_mult_82_ab_9__10_), .B(
        u5_mult_82_CARRYB_8__10_), .CI(u5_mult_82_SUMB_8__11_), .CO(
        u5_mult_82_CARRYB_9__10_), .S(u5_mult_82_SUMB_9__10_) );
  FA_X1 u5_mult_82_S2_9_9 ( .A(u5_mult_82_ab_9__9_), .B(
        u5_mult_82_CARRYB_8__9_), .CI(u5_mult_82_SUMB_8__10_), .CO(
        u5_mult_82_CARRYB_9__9_), .S(u5_mult_82_SUMB_9__9_) );
  FA_X1 u5_mult_82_S2_9_8 ( .A(u5_mult_82_ab_9__8_), .B(
        u5_mult_82_CARRYB_8__8_), .CI(u5_mult_82_SUMB_8__9_), .CO(
        u5_mult_82_CARRYB_9__8_), .S(u5_mult_82_SUMB_9__8_) );
  FA_X1 u5_mult_82_S2_9_7 ( .A(u5_mult_82_ab_9__7_), .B(
        u5_mult_82_CARRYB_8__7_), .CI(u5_mult_82_SUMB_8__8_), .CO(
        u5_mult_82_CARRYB_9__7_), .S(u5_mult_82_SUMB_9__7_) );
  FA_X1 u5_mult_82_S2_9_6 ( .A(u5_mult_82_ab_9__6_), .B(
        u5_mult_82_CARRYB_8__6_), .CI(u5_mult_82_SUMB_8__7_), .CO(
        u5_mult_82_CARRYB_9__6_), .S(u5_mult_82_SUMB_9__6_) );
  FA_X1 u5_mult_82_S2_9_5 ( .A(u5_mult_82_ab_9__5_), .B(
        u5_mult_82_CARRYB_8__5_), .CI(u5_mult_82_SUMB_8__6_), .CO(
        u5_mult_82_CARRYB_9__5_), .S(u5_mult_82_SUMB_9__5_) );
  FA_X1 u5_mult_82_S2_9_4 ( .A(u5_mult_82_ab_9__4_), .B(
        u5_mult_82_CARRYB_8__4_), .CI(u5_mult_82_SUMB_8__5_), .CO(
        u5_mult_82_CARRYB_9__4_), .S(u5_mult_82_SUMB_9__4_) );
  FA_X1 u5_mult_82_S2_9_3 ( .A(u5_mult_82_ab_9__3_), .B(
        u5_mult_82_CARRYB_8__3_), .CI(u5_mult_82_SUMB_8__4_), .CO(
        u5_mult_82_CARRYB_9__3_), .S(u5_mult_82_SUMB_9__3_) );
  FA_X1 u5_mult_82_S2_9_2 ( .A(u5_mult_82_ab_9__2_), .B(
        u5_mult_82_CARRYB_8__2_), .CI(u5_mult_82_SUMB_8__3_), .CO(
        u5_mult_82_CARRYB_9__2_), .S(u5_mult_82_SUMB_9__2_) );
  FA_X1 u5_mult_82_S2_9_1 ( .A(u5_mult_82_ab_9__1_), .B(
        u5_mult_82_CARRYB_8__1_), .CI(u5_mult_82_SUMB_8__2_), .CO(
        u5_mult_82_CARRYB_9__1_), .S(u5_mult_82_SUMB_9__1_) );
  FA_X1 u5_mult_82_S1_9_0 ( .A(u5_mult_82_ab_9__0_), .B(
        u5_mult_82_CARRYB_8__0_), .CI(u5_mult_82_SUMB_8__1_), .CO(
        u5_mult_82_CARRYB_9__0_), .S(u5_N9) );
  FA_X1 u5_mult_82_S2_10_48 ( .A(u5_mult_82_ab_10__48_), .B(
        u5_mult_82_CARRYB_9__48_), .CI(u5_mult_82_SUMB_9__49_), .CO(
        u5_mult_82_CARRYB_10__48_), .S(u5_mult_82_SUMB_10__48_) );
  FA_X1 u5_mult_82_S2_10_47 ( .A(u5_mult_82_ab_10__47_), .B(
        u5_mult_82_CARRYB_9__47_), .CI(u5_mult_82_SUMB_9__48_), .CO(
        u5_mult_82_CARRYB_10__47_), .S(u5_mult_82_SUMB_10__47_) );
  FA_X1 u5_mult_82_S2_10_41 ( .A(u5_mult_82_ab_10__41_), .B(
        u5_mult_82_CARRYB_9__41_), .CI(u5_mult_82_SUMB_9__42_), .CO(
        u5_mult_82_CARRYB_10__41_), .S(u5_mult_82_SUMB_10__41_) );
  FA_X1 u5_mult_82_S2_10_40 ( .A(u5_mult_82_ab_10__40_), .B(
        u5_mult_82_CARRYB_9__40_), .CI(u5_mult_82_SUMB_9__41_), .CO(
        u5_mult_82_CARRYB_10__40_), .S(u5_mult_82_SUMB_10__40_) );
  FA_X1 u5_mult_82_S2_10_39 ( .A(u5_mult_82_ab_10__39_), .B(
        u5_mult_82_CARRYB_9__39_), .CI(u5_mult_82_SUMB_9__40_), .CO(
        u5_mult_82_CARRYB_10__39_), .S(u5_mult_82_SUMB_10__39_) );
  FA_X1 u5_mult_82_S2_10_34 ( .A(u5_mult_82_ab_10__34_), .B(
        u5_mult_82_CARRYB_9__34_), .CI(u5_mult_82_SUMB_9__35_), .CO(
        u5_mult_82_CARRYB_10__34_), .S(u5_mult_82_SUMB_10__34_) );
  FA_X1 u5_mult_82_S2_10_31 ( .A(u5_mult_82_ab_10__31_), .B(
        u5_mult_82_CARRYB_9__31_), .CI(u5_mult_82_SUMB_9__32_), .CO(
        u5_mult_82_CARRYB_10__31_), .S(u5_mult_82_SUMB_10__31_) );
  FA_X1 u5_mult_82_S2_10_24 ( .A(u5_mult_82_ab_10__24_), .B(
        u5_mult_82_CARRYB_9__24_), .CI(u5_mult_82_SUMB_9__25_), .CO(
        u5_mult_82_CARRYB_10__24_), .S(u5_mult_82_SUMB_10__24_) );
  FA_X1 u5_mult_82_S2_10_23 ( .A(u5_mult_82_ab_10__23_), .B(
        u5_mult_82_CARRYB_9__23_), .CI(u5_mult_82_SUMB_9__24_), .CO(
        u5_mult_82_CARRYB_10__23_), .S(u5_mult_82_SUMB_10__23_) );
  FA_X1 u5_mult_82_S2_10_22 ( .A(u5_mult_82_ab_10__22_), .B(
        u5_mult_82_CARRYB_9__22_), .CI(u5_mult_82_SUMB_9__23_), .CO(
        u5_mult_82_CARRYB_10__22_), .S(u5_mult_82_SUMB_10__22_) );
  FA_X1 u5_mult_82_S2_10_21 ( .A(u5_mult_82_ab_10__21_), .B(
        u5_mult_82_CARRYB_9__21_), .CI(u5_mult_82_SUMB_9__22_), .CO(
        u5_mult_82_CARRYB_10__21_), .S(u5_mult_82_SUMB_10__21_) );
  FA_X1 u5_mult_82_S2_10_19 ( .A(u5_mult_82_ab_10__19_), .B(
        u5_mult_82_CARRYB_9__19_), .CI(u5_mult_82_SUMB_9__20_), .CO(
        u5_mult_82_CARRYB_10__19_), .S(u5_mult_82_SUMB_10__19_) );
  FA_X1 u5_mult_82_S2_10_16 ( .A(u5_mult_82_ab_10__16_), .B(
        u5_mult_82_CARRYB_9__16_), .CI(u5_mult_82_SUMB_9__17_), .CO(
        u5_mult_82_CARRYB_10__16_), .S(u5_mult_82_SUMB_10__16_) );
  FA_X1 u5_mult_82_S2_10_14 ( .A(u5_mult_82_ab_10__14_), .B(
        u5_mult_82_CARRYB_9__14_), .CI(u5_mult_82_SUMB_9__15_), .CO(
        u5_mult_82_CARRYB_10__14_), .S(u5_mult_82_SUMB_10__14_) );
  FA_X1 u5_mult_82_S2_10_13 ( .A(u5_mult_82_ab_10__13_), .B(
        u5_mult_82_CARRYB_9__13_), .CI(u5_mult_82_SUMB_9__14_), .CO(
        u5_mult_82_CARRYB_10__13_), .S(u5_mult_82_SUMB_10__13_) );
  FA_X1 u5_mult_82_S2_10_11 ( .A(u5_mult_82_ab_10__11_), .B(
        u5_mult_82_CARRYB_9__11_), .CI(u5_mult_82_SUMB_9__12_), .CO(
        u5_mult_82_CARRYB_10__11_), .S(u5_mult_82_SUMB_10__11_) );
  FA_X1 u5_mult_82_S2_10_10 ( .A(u5_mult_82_ab_10__10_), .B(
        u5_mult_82_CARRYB_9__10_), .CI(u5_mult_82_SUMB_9__11_), .CO(
        u5_mult_82_CARRYB_10__10_), .S(u5_mult_82_SUMB_10__10_) );
  FA_X1 u5_mult_82_S2_10_9 ( .A(u5_mult_82_ab_10__9_), .B(
        u5_mult_82_CARRYB_9__9_), .CI(u5_mult_82_SUMB_9__10_), .CO(
        u5_mult_82_CARRYB_10__9_), .S(u5_mult_82_SUMB_10__9_) );
  FA_X1 u5_mult_82_S2_10_8 ( .A(u5_mult_82_ab_10__8_), .B(
        u5_mult_82_CARRYB_9__8_), .CI(u5_mult_82_SUMB_9__9_), .CO(
        u5_mult_82_CARRYB_10__8_), .S(u5_mult_82_SUMB_10__8_) );
  FA_X1 u5_mult_82_S2_10_7 ( .A(u5_mult_82_ab_10__7_), .B(
        u5_mult_82_CARRYB_9__7_), .CI(u5_mult_82_SUMB_9__8_), .CO(
        u5_mult_82_CARRYB_10__7_), .S(u5_mult_82_SUMB_10__7_) );
  FA_X1 u5_mult_82_S2_10_6 ( .A(u5_mult_82_ab_10__6_), .B(
        u5_mult_82_CARRYB_9__6_), .CI(u5_mult_82_SUMB_9__7_), .CO(
        u5_mult_82_CARRYB_10__6_), .S(u5_mult_82_SUMB_10__6_) );
  FA_X1 u5_mult_82_S2_10_5 ( .A(u5_mult_82_ab_10__5_), .B(
        u5_mult_82_CARRYB_9__5_), .CI(u5_mult_82_SUMB_9__6_), .CO(
        u5_mult_82_CARRYB_10__5_), .S(u5_mult_82_SUMB_10__5_) );
  FA_X1 u5_mult_82_S2_10_4 ( .A(u5_mult_82_ab_10__4_), .B(
        u5_mult_82_CARRYB_9__4_), .CI(u5_mult_82_SUMB_9__5_), .CO(
        u5_mult_82_CARRYB_10__4_), .S(u5_mult_82_SUMB_10__4_) );
  FA_X1 u5_mult_82_S2_10_3 ( .A(u5_mult_82_ab_10__3_), .B(
        u5_mult_82_CARRYB_9__3_), .CI(u5_mult_82_SUMB_9__4_), .CO(
        u5_mult_82_CARRYB_10__3_), .S(u5_mult_82_SUMB_10__3_) );
  FA_X1 u5_mult_82_S2_10_2 ( .A(u5_mult_82_ab_10__2_), .B(
        u5_mult_82_CARRYB_9__2_), .CI(u5_mult_82_SUMB_9__3_), .CO(
        u5_mult_82_CARRYB_10__2_), .S(u5_mult_82_SUMB_10__2_) );
  FA_X1 u5_mult_82_S2_10_1 ( .A(u5_mult_82_ab_10__1_), .B(
        u5_mult_82_CARRYB_9__1_), .CI(u5_mult_82_SUMB_9__2_), .CO(
        u5_mult_82_CARRYB_10__1_), .S(u5_mult_82_SUMB_10__1_) );
  FA_X1 u5_mult_82_S1_10_0 ( .A(u5_mult_82_ab_10__0_), .B(
        u5_mult_82_CARRYB_9__0_), .CI(u5_mult_82_SUMB_9__1_), .CO(
        u5_mult_82_CARRYB_10__0_), .S(u5_N10) );
  FA_X1 u5_mult_82_S2_11_48 ( .A(u5_mult_82_ab_11__48_), .B(
        u5_mult_82_CARRYB_10__48_), .CI(u5_mult_82_SUMB_10__49_), .CO(
        u5_mult_82_CARRYB_11__48_), .S(u5_mult_82_SUMB_11__48_) );
  FA_X1 u5_mult_82_S2_11_47 ( .A(u5_mult_82_ab_11__47_), .B(
        u5_mult_82_CARRYB_10__47_), .CI(u5_mult_82_SUMB_10__48_), .CO(
        u5_mult_82_CARRYB_11__47_), .S(u5_mult_82_SUMB_11__47_) );
  FA_X1 u5_mult_82_S2_11_46 ( .A(u5_mult_82_ab_11__46_), .B(
        u5_mult_82_CARRYB_10__46_), .CI(u5_mult_82_SUMB_10__47_), .CO(
        u5_mult_82_CARRYB_11__46_), .S(u5_mult_82_SUMB_11__46_) );
  FA_X1 u5_mult_82_S2_11_39 ( .A(u5_mult_82_CARRYB_10__39_), .B(
        u5_mult_82_ab_11__39_), .CI(u5_mult_82_SUMB_10__40_), .CO(
        u5_mult_82_CARRYB_11__39_), .S(u5_mult_82_SUMB_11__39_) );
  FA_X1 u5_mult_82_S2_11_33 ( .A(u5_mult_82_ab_11__33_), .B(
        u5_mult_82_CARRYB_10__33_), .CI(u5_mult_82_SUMB_10__34_), .CO(
        u5_mult_82_CARRYB_11__33_), .S(u5_mult_82_SUMB_11__33_) );
  FA_X1 u5_mult_82_S2_11_28 ( .A(u5_mult_82_ab_11__28_), .B(
        u5_mult_82_CARRYB_10__28_), .CI(u5_mult_82_SUMB_10__29_), .CO(
        u5_mult_82_CARRYB_11__28_), .S(u5_mult_82_SUMB_11__28_) );
  FA_X1 u5_mult_82_S2_11_26 ( .A(u5_mult_82_ab_11__26_), .B(
        u5_mult_82_CARRYB_10__26_), .CI(u5_mult_82_SUMB_10__27_), .CO(
        u5_mult_82_CARRYB_11__26_), .S(u5_mult_82_SUMB_11__26_) );
  FA_X1 u5_mult_82_S2_11_23 ( .A(u5_mult_82_ab_11__23_), .B(
        u5_mult_82_CARRYB_10__23_), .CI(u5_mult_82_SUMB_10__24_), .CO(
        u5_mult_82_CARRYB_11__23_), .S(u5_mult_82_SUMB_11__23_) );
  FA_X1 u5_mult_82_S2_11_22 ( .A(u5_mult_82_ab_11__22_), .B(
        u5_mult_82_CARRYB_10__22_), .CI(u5_mult_82_SUMB_10__23_), .CO(
        u5_mult_82_CARRYB_11__22_), .S(u5_mult_82_SUMB_11__22_) );
  FA_X1 u5_mult_82_S2_11_21 ( .A(u5_mult_82_ab_11__21_), .B(
        u5_mult_82_CARRYB_10__21_), .CI(u5_mult_82_SUMB_10__22_), .CO(
        u5_mult_82_CARRYB_11__21_), .S(u5_mult_82_SUMB_11__21_) );
  FA_X1 u5_mult_82_S2_11_18 ( .A(u5_mult_82_ab_11__18_), .B(
        u5_mult_82_CARRYB_10__18_), .CI(u5_mult_82_SUMB_10__19_), .CO(
        u5_mult_82_CARRYB_11__18_), .S(u5_mult_82_SUMB_11__18_) );
  FA_X1 u5_mult_82_S2_11_14 ( .A(u5_mult_82_ab_11__14_), .B(
        u5_mult_82_CARRYB_10__14_), .CI(u5_mult_82_SUMB_10__15_), .CO(
        u5_mult_82_CARRYB_11__14_), .S(u5_mult_82_SUMB_11__14_) );
  FA_X1 u5_mult_82_S2_11_13 ( .A(u5_mult_82_ab_11__13_), .B(
        u5_mult_82_CARRYB_10__13_), .CI(u5_mult_82_SUMB_10__14_), .CO(
        u5_mult_82_CARRYB_11__13_), .S(u5_mult_82_SUMB_11__13_) );
  FA_X1 u5_mult_82_S2_11_12 ( .A(u5_mult_82_ab_11__12_), .B(
        u5_mult_82_CARRYB_10__12_), .CI(u5_mult_82_SUMB_10__13_), .CO(
        u5_mult_82_CARRYB_11__12_), .S(u5_mult_82_SUMB_11__12_) );
  FA_X1 u5_mult_82_S2_11_10 ( .A(u5_mult_82_ab_11__10_), .B(
        u5_mult_82_CARRYB_10__10_), .CI(u5_mult_82_SUMB_10__11_), .CO(
        u5_mult_82_CARRYB_11__10_), .S(u5_mult_82_SUMB_11__10_) );
  FA_X1 u5_mult_82_S2_11_9 ( .A(u5_mult_82_ab_11__9_), .B(
        u5_mult_82_CARRYB_10__9_), .CI(u5_mult_82_SUMB_10__10_), .CO(
        u5_mult_82_CARRYB_11__9_), .S(u5_mult_82_SUMB_11__9_) );
  FA_X1 u5_mult_82_S2_11_8 ( .A(u5_mult_82_ab_11__8_), .B(
        u5_mult_82_CARRYB_10__8_), .CI(u5_mult_82_SUMB_10__9_), .CO(
        u5_mult_82_CARRYB_11__8_), .S(u5_mult_82_SUMB_11__8_) );
  FA_X1 u5_mult_82_S2_11_7 ( .A(u5_mult_82_ab_11__7_), .B(
        u5_mult_82_CARRYB_10__7_), .CI(u5_mult_82_SUMB_10__8_), .CO(
        u5_mult_82_CARRYB_11__7_), .S(u5_mult_82_SUMB_11__7_) );
  FA_X1 u5_mult_82_S2_11_6 ( .A(u5_mult_82_ab_11__6_), .B(
        u5_mult_82_CARRYB_10__6_), .CI(u5_mult_82_SUMB_10__7_), .CO(
        u5_mult_82_CARRYB_11__6_), .S(u5_mult_82_SUMB_11__6_) );
  FA_X1 u5_mult_82_S2_11_5 ( .A(u5_mult_82_ab_11__5_), .B(
        u5_mult_82_CARRYB_10__5_), .CI(u5_mult_82_SUMB_10__6_), .CO(
        u5_mult_82_CARRYB_11__5_), .S(u5_mult_82_SUMB_11__5_) );
  FA_X1 u5_mult_82_S2_11_4 ( .A(u5_mult_82_ab_11__4_), .B(
        u5_mult_82_CARRYB_10__4_), .CI(u5_mult_82_SUMB_10__5_), .CO(
        u5_mult_82_CARRYB_11__4_), .S(u5_mult_82_SUMB_11__4_) );
  FA_X1 u5_mult_82_S2_11_3 ( .A(u5_mult_82_ab_11__3_), .B(
        u5_mult_82_CARRYB_10__3_), .CI(u5_mult_82_SUMB_10__4_), .CO(
        u5_mult_82_CARRYB_11__3_), .S(u5_mult_82_SUMB_11__3_) );
  FA_X1 u5_mult_82_S2_11_2 ( .A(u5_mult_82_ab_11__2_), .B(
        u5_mult_82_CARRYB_10__2_), .CI(u5_mult_82_SUMB_10__3_), .CO(
        u5_mult_82_CARRYB_11__2_), .S(u5_mult_82_SUMB_11__2_) );
  FA_X1 u5_mult_82_S2_11_1 ( .A(u5_mult_82_ab_11__1_), .B(
        u5_mult_82_CARRYB_10__1_), .CI(u5_mult_82_SUMB_10__2_), .CO(
        u5_mult_82_CARRYB_11__1_), .S(u5_mult_82_SUMB_11__1_) );
  FA_X1 u5_mult_82_S1_11_0 ( .A(u5_mult_82_ab_11__0_), .B(
        u5_mult_82_CARRYB_10__0_), .CI(u5_mult_82_SUMB_10__1_), .CO(
        u5_mult_82_CARRYB_11__0_), .S(u5_N11) );
  FA_X1 u5_mult_82_S2_12_49 ( .A(u5_mult_82_ab_12__49_), .B(
        u5_mult_82_CARRYB_11__49_), .CI(u5_mult_82_SUMB_11__50_), .CO(
        u5_mult_82_CARRYB_12__49_), .S(u5_mult_82_SUMB_12__49_) );
  FA_X1 u5_mult_82_S2_12_48 ( .A(u5_mult_82_CARRYB_11__48_), .B(
        u5_mult_82_ab_12__48_), .CI(u5_mult_82_SUMB_11__49_), .CO(
        u5_mult_82_CARRYB_12__48_), .S(u5_mult_82_SUMB_12__48_) );
  FA_X1 u5_mult_82_S2_12_36 ( .A(u5_mult_82_ab_12__36_), .B(
        u5_mult_82_CARRYB_11__36_), .CI(u5_mult_82_SUMB_11__37_), .CO(
        u5_mult_82_CARRYB_12__36_), .S(u5_mult_82_SUMB_12__36_) );
  FA_X1 u5_mult_82_S2_12_34 ( .A(u5_mult_82_ab_12__34_), .B(
        u5_mult_82_CARRYB_11__34_), .CI(u5_mult_82_SUMB_11__35_), .CO(
        u5_mult_82_CARRYB_12__34_), .S(u5_mult_82_SUMB_12__34_) );
  FA_X1 u5_mult_82_S2_12_28 ( .A(u5_mult_82_ab_12__28_), .B(
        u5_mult_82_CARRYB_11__28_), .CI(u5_mult_82_SUMB_11__29_), .CO(
        u5_mult_82_CARRYB_12__28_), .S(u5_mult_82_SUMB_12__28_) );
  FA_X1 u5_mult_82_S2_12_27 ( .A(u5_mult_82_ab_12__27_), .B(
        u5_mult_82_CARRYB_11__27_), .CI(u5_mult_82_SUMB_11__28_), .CO(
        u5_mult_82_CARRYB_12__27_), .S(u5_mult_82_SUMB_12__27_) );
  FA_X1 u5_mult_82_S2_12_24 ( .A(u5_mult_82_ab_12__24_), .B(
        u5_mult_82_CARRYB_11__24_), .CI(u5_mult_82_SUMB_11__25_), .CO(
        u5_mult_82_CARRYB_12__24_), .S(u5_mult_82_SUMB_12__24_) );
  FA_X1 u5_mult_82_S2_12_22 ( .A(u5_mult_82_ab_12__22_), .B(
        u5_mult_82_CARRYB_11__22_), .CI(u5_mult_82_SUMB_11__23_), .CO(
        u5_mult_82_CARRYB_12__22_), .S(u5_mult_82_SUMB_12__22_) );
  FA_X1 u5_mult_82_S2_12_20 ( .A(u5_mult_82_ab_12__20_), .B(
        u5_mult_82_CARRYB_11__20_), .CI(u5_mult_82_SUMB_11__21_), .CO(
        u5_mult_82_CARRYB_12__20_), .S(u5_mult_82_SUMB_12__20_) );
  FA_X1 u5_mult_82_S2_12_16 ( .A(u5_mult_82_ab_12__16_), .B(
        u5_mult_82_CARRYB_11__16_), .CI(u5_mult_82_SUMB_11__17_), .CO(
        u5_mult_82_CARRYB_12__16_), .S(u5_mult_82_SUMB_12__16_) );
  FA_X1 u5_mult_82_S2_12_15 ( .A(u5_mult_82_ab_12__15_), .B(
        u5_mult_82_CARRYB_11__15_), .CI(u5_mult_82_SUMB_11__16_), .CO(
        u5_mult_82_CARRYB_12__15_), .S(u5_mult_82_SUMB_12__15_) );
  FA_X1 u5_mult_82_S2_12_13 ( .A(u5_mult_82_ab_12__13_), .B(
        u5_mult_82_CARRYB_11__13_), .CI(u5_mult_82_SUMB_11__14_), .CO(
        u5_mult_82_CARRYB_12__13_), .S(u5_mult_82_SUMB_12__13_) );
  FA_X1 u5_mult_82_S2_12_11 ( .A(u5_mult_82_ab_12__11_), .B(
        u5_mult_82_CARRYB_11__11_), .CI(u5_mult_82_SUMB_11__12_), .CO(
        u5_mult_82_CARRYB_12__11_), .S(u5_mult_82_SUMB_12__11_) );
  FA_X1 u5_mult_82_S2_12_9 ( .A(u5_mult_82_ab_12__9_), .B(
        u5_mult_82_CARRYB_11__9_), .CI(u5_mult_82_SUMB_11__10_), .CO(
        u5_mult_82_CARRYB_12__9_), .S(u5_mult_82_SUMB_12__9_) );
  FA_X1 u5_mult_82_S2_12_8 ( .A(u5_mult_82_ab_12__8_), .B(
        u5_mult_82_CARRYB_11__8_), .CI(u5_mult_82_SUMB_11__9_), .CO(
        u5_mult_82_CARRYB_12__8_), .S(u5_mult_82_SUMB_12__8_) );
  FA_X1 u5_mult_82_S2_12_7 ( .A(u5_mult_82_ab_12__7_), .B(
        u5_mult_82_CARRYB_11__7_), .CI(u5_mult_82_SUMB_11__8_), .CO(
        u5_mult_82_CARRYB_12__7_), .S(u5_mult_82_SUMB_12__7_) );
  FA_X1 u5_mult_82_S2_12_6 ( .A(u5_mult_82_ab_12__6_), .B(
        u5_mult_82_CARRYB_11__6_), .CI(u5_mult_82_SUMB_11__7_), .CO(
        u5_mult_82_CARRYB_12__6_), .S(u5_mult_82_SUMB_12__6_) );
  FA_X1 u5_mult_82_S2_12_5 ( .A(u5_mult_82_ab_12__5_), .B(
        u5_mult_82_CARRYB_11__5_), .CI(u5_mult_82_SUMB_11__6_), .CO(
        u5_mult_82_CARRYB_12__5_), .S(u5_mult_82_SUMB_12__5_) );
  FA_X1 u5_mult_82_S2_12_4 ( .A(u5_mult_82_ab_12__4_), .B(
        u5_mult_82_CARRYB_11__4_), .CI(u5_mult_82_SUMB_11__5_), .CO(
        u5_mult_82_CARRYB_12__4_), .S(u5_mult_82_SUMB_12__4_) );
  FA_X1 u5_mult_82_S2_12_3 ( .A(u5_mult_82_ab_12__3_), .B(
        u5_mult_82_CARRYB_11__3_), .CI(u5_mult_82_SUMB_11__4_), .CO(
        u5_mult_82_CARRYB_12__3_), .S(u5_mult_82_SUMB_12__3_) );
  FA_X1 u5_mult_82_S2_12_2 ( .A(u5_mult_82_ab_12__2_), .B(
        u5_mult_82_CARRYB_11__2_), .CI(u5_mult_82_SUMB_11__3_), .CO(
        u5_mult_82_CARRYB_12__2_), .S(u5_mult_82_SUMB_12__2_) );
  FA_X1 u5_mult_82_S2_12_1 ( .A(u5_mult_82_ab_12__1_), .B(
        u5_mult_82_CARRYB_11__1_), .CI(u5_mult_82_SUMB_11__2_), .CO(
        u5_mult_82_CARRYB_12__1_), .S(u5_mult_82_SUMB_12__1_) );
  FA_X1 u5_mult_82_S1_12_0 ( .A(u5_mult_82_ab_12__0_), .B(
        u5_mult_82_CARRYB_11__0_), .CI(u5_mult_82_SUMB_11__1_), .CO(
        u5_mult_82_CARRYB_12__0_), .S(u5_N12) );
  FA_X1 u5_mult_82_S2_13_50 ( .A(u5_mult_82_ab_13__50_), .B(
        u5_mult_82_SUMB_12__51_), .CI(u5_mult_82_CARRYB_12__50_), .CO(
        u5_mult_82_CARRYB_13__50_), .S(u5_mult_82_SUMB_13__50_) );
  FA_X1 u5_mult_82_S2_13_47 ( .A(u5_mult_82_ab_13__47_), .B(
        u5_mult_82_CARRYB_12__47_), .CI(u5_mult_82_SUMB_12__48_), .CO(
        u5_mult_82_CARRYB_13__47_), .S(u5_mult_82_SUMB_13__47_) );
  FA_X1 u5_mult_82_S2_13_43 ( .A(u5_mult_82_ab_13__43_), .B(
        u5_mult_82_CARRYB_12__43_), .CI(u5_mult_82_SUMB_12__44_), .CO(
        u5_mult_82_CARRYB_13__43_), .S(u5_mult_82_SUMB_13__43_) );
  FA_X1 u5_mult_82_S2_13_42 ( .A(u5_mult_82_ab_13__42_), .B(
        u5_mult_82_CARRYB_12__42_), .CI(u5_mult_82_SUMB_12__43_), .CO(
        u5_mult_82_CARRYB_13__42_), .S(u5_mult_82_SUMB_13__42_) );
  FA_X1 u5_mult_82_S2_13_40 ( .A(u5_mult_82_ab_13__40_), .B(
        u5_mult_82_CARRYB_12__40_), .CI(u5_mult_82_SUMB_12__41_), .CO(
        u5_mult_82_CARRYB_13__40_), .S(u5_mult_82_SUMB_13__40_) );
  FA_X1 u5_mult_82_S2_13_39 ( .A(u5_mult_82_ab_13__39_), .B(
        u5_mult_82_CARRYB_12__39_), .CI(u5_mult_82_SUMB_12__40_), .CO(
        u5_mult_82_CARRYB_13__39_), .S(u5_mult_82_SUMB_13__39_) );
  FA_X1 u5_mult_82_S2_13_35 ( .A(u5_mult_82_ab_13__35_), .B(
        u5_mult_82_CARRYB_12__35_), .CI(u5_mult_82_SUMB_12__36_), .CO(
        u5_mult_82_CARRYB_13__35_), .S(u5_mult_82_SUMB_13__35_) );
  FA_X1 u5_mult_82_S2_13_33 ( .A(u5_mult_82_ab_13__33_), .B(
        u5_mult_82_CARRYB_12__33_), .CI(u5_mult_82_SUMB_12__34_), .CO(
        u5_mult_82_CARRYB_13__33_), .S(u5_mult_82_SUMB_13__33_) );
  FA_X1 u5_mult_82_S2_13_28 ( .A(u5_mult_82_ab_13__28_), .B(
        u5_mult_82_CARRYB_12__28_), .CI(u5_mult_82_SUMB_12__29_), .CO(
        u5_mult_82_CARRYB_13__28_), .S(u5_mult_82_SUMB_13__28_) );
  FA_X1 u5_mult_82_S2_13_27 ( .A(u5_mult_82_ab_13__27_), .B(
        u5_mult_82_CARRYB_12__27_), .CI(u5_mult_82_SUMB_12__28_), .CO(
        u5_mult_82_CARRYB_13__27_), .S(u5_mult_82_SUMB_13__27_) );
  FA_X1 u5_mult_82_S2_13_19 ( .A(u5_mult_82_ab_13__19_), .B(
        u5_mult_82_CARRYB_12__19_), .CI(u5_mult_82_SUMB_12__20_), .CO(
        u5_mult_82_CARRYB_13__19_), .S(u5_mult_82_SUMB_13__19_) );
  FA_X1 u5_mult_82_S2_13_17 ( .A(u5_mult_82_ab_13__17_), .B(
        u5_mult_82_CARRYB_12__17_), .CI(u5_mult_82_SUMB_12__18_), .CO(
        u5_mult_82_CARRYB_13__17_), .S(u5_mult_82_SUMB_13__17_) );
  FA_X1 u5_mult_82_S2_13_15 ( .A(u5_mult_82_ab_13__15_), .B(
        u5_mult_82_CARRYB_12__15_), .CI(u5_mult_82_SUMB_12__16_), .CO(
        u5_mult_82_CARRYB_13__15_), .S(u5_mult_82_SUMB_13__15_) );
  FA_X1 u5_mult_82_S2_13_14 ( .A(u5_mult_82_ab_13__14_), .B(
        u5_mult_82_CARRYB_12__14_), .CI(u5_mult_82_SUMB_12__15_), .CO(
        u5_mult_82_CARRYB_13__14_), .S(u5_mult_82_SUMB_13__14_) );
  FA_X1 u5_mult_82_S2_13_13 ( .A(u5_mult_82_CARRYB_12__13_), .B(
        u5_mult_82_ab_13__13_), .CI(u5_mult_82_SUMB_12__14_), .CO(
        u5_mult_82_CARRYB_13__13_), .S(u5_mult_82_SUMB_13__13_) );
  FA_X1 u5_mult_82_S2_13_12 ( .A(u5_mult_82_ab_13__12_), .B(
        u5_mult_82_CARRYB_12__12_), .CI(u5_mult_82_SUMB_12__13_), .CO(
        u5_mult_82_CARRYB_13__12_), .S(u5_mult_82_SUMB_13__12_) );
  FA_X1 u5_mult_82_S2_13_9 ( .A(u5_mult_82_ab_13__9_), .B(
        u5_mult_82_CARRYB_12__9_), .CI(u5_mult_82_SUMB_12__10_), .CO(
        u5_mult_82_CARRYB_13__9_), .S(u5_mult_82_SUMB_13__9_) );
  FA_X1 u5_mult_82_S2_13_8 ( .A(u5_mult_82_ab_13__8_), .B(
        u5_mult_82_CARRYB_12__8_), .CI(u5_mult_82_SUMB_12__9_), .CO(
        u5_mult_82_CARRYB_13__8_), .S(u5_mult_82_SUMB_13__8_) );
  FA_X1 u5_mult_82_S2_13_7 ( .A(u5_mult_82_ab_13__7_), .B(
        u5_mult_82_CARRYB_12__7_), .CI(u5_mult_82_SUMB_12__8_), .CO(
        u5_mult_82_CARRYB_13__7_), .S(u5_mult_82_SUMB_13__7_) );
  FA_X1 u5_mult_82_S2_13_6 ( .A(u5_mult_82_ab_13__6_), .B(
        u5_mult_82_CARRYB_12__6_), .CI(u5_mult_82_SUMB_12__7_), .CO(
        u5_mult_82_CARRYB_13__6_), .S(u5_mult_82_SUMB_13__6_) );
  FA_X1 u5_mult_82_S2_13_5 ( .A(u5_mult_82_ab_13__5_), .B(
        u5_mult_82_CARRYB_12__5_), .CI(u5_mult_82_SUMB_12__6_), .CO(
        u5_mult_82_CARRYB_13__5_), .S(u5_mult_82_SUMB_13__5_) );
  FA_X1 u5_mult_82_S2_13_4 ( .A(u5_mult_82_ab_13__4_), .B(
        u5_mult_82_CARRYB_12__4_), .CI(u5_mult_82_SUMB_12__5_), .CO(
        u5_mult_82_CARRYB_13__4_), .S(u5_mult_82_SUMB_13__4_) );
  FA_X1 u5_mult_82_S2_13_3 ( .A(u5_mult_82_ab_13__3_), .B(
        u5_mult_82_CARRYB_12__3_), .CI(u5_mult_82_SUMB_12__4_), .CO(
        u5_mult_82_CARRYB_13__3_), .S(u5_mult_82_SUMB_13__3_) );
  FA_X1 u5_mult_82_S2_13_2 ( .A(u5_mult_82_ab_13__2_), .B(
        u5_mult_82_CARRYB_12__2_), .CI(u5_mult_82_SUMB_12__3_), .CO(
        u5_mult_82_CARRYB_13__2_), .S(u5_mult_82_SUMB_13__2_) );
  FA_X1 u5_mult_82_S2_13_1 ( .A(u5_mult_82_ab_13__1_), .B(
        u5_mult_82_CARRYB_12__1_), .CI(u5_mult_82_SUMB_12__2_), .CO(
        u5_mult_82_CARRYB_13__1_), .S(u5_mult_82_SUMB_13__1_) );
  FA_X1 u5_mult_82_S1_13_0 ( .A(u5_mult_82_ab_13__0_), .B(
        u5_mult_82_CARRYB_12__0_), .CI(u5_mult_82_SUMB_12__1_), .CO(
        u5_mult_82_CARRYB_13__0_), .S(u5_N13) );
  FA_X1 u5_mult_82_S2_14_50 ( .A(u5_mult_82_ab_14__50_), .B(
        u5_mult_82_CARRYB_13__50_), .CI(u5_mult_82_SUMB_13__51_), .CO(
        u5_mult_82_CARRYB_14__50_), .S(u5_mult_82_SUMB_14__50_) );
  FA_X1 u5_mult_82_S2_14_46 ( .A(u5_mult_82_ab_14__46_), .B(
        u5_mult_82_CARRYB_13__46_), .CI(u5_mult_82_SUMB_13__47_), .CO(
        u5_mult_82_CARRYB_14__46_), .S(u5_mult_82_SUMB_14__46_) );
  FA_X1 u5_mult_82_S2_14_38 ( .A(u5_mult_82_CARRYB_13__38_), .B(
        u5_mult_82_ab_14__38_), .CI(u5_mult_82_SUMB_13__39_), .CO(
        u5_mult_82_CARRYB_14__38_), .S(u5_mult_82_SUMB_14__38_) );
  FA_X1 u5_mult_82_S2_14_37 ( .A(u5_mult_82_ab_14__37_), .B(
        u5_mult_82_CARRYB_13__37_), .CI(u5_mult_82_SUMB_13__38_), .CO(
        u5_mult_82_CARRYB_14__37_), .S(u5_mult_82_SUMB_14__37_) );
  FA_X1 u5_mult_82_S2_14_35 ( .A(u5_mult_82_ab_14__35_), .B(
        u5_mult_82_CARRYB_13__35_), .CI(u5_mult_82_SUMB_13__36_), .CO(
        u5_mult_82_CARRYB_14__35_), .S(u5_mult_82_SUMB_14__35_) );
  FA_X1 u5_mult_82_S2_14_33 ( .A(u5_mult_82_ab_14__33_), .B(
        u5_mult_82_CARRYB_13__33_), .CI(u5_mult_82_SUMB_13__34_), .CO(
        u5_mult_82_CARRYB_14__33_), .S(u5_mult_82_SUMB_14__33_) );
  FA_X1 u5_mult_82_S2_14_32 ( .A(u5_mult_82_ab_14__32_), .B(
        u5_mult_82_CARRYB_13__32_), .CI(u5_mult_82_SUMB_13__33_), .CO(
        u5_mult_82_CARRYB_14__32_), .S(u5_mult_82_SUMB_14__32_) );
  FA_X1 u5_mult_82_S2_14_31 ( .A(u5_mult_82_ab_14__31_), .B(
        u5_mult_82_CARRYB_13__31_), .CI(u5_mult_82_SUMB_13__32_), .CO(
        u5_mult_82_CARRYB_14__31_), .S(u5_mult_82_SUMB_14__31_) );
  FA_X1 u5_mult_82_S2_14_30 ( .A(u5_mult_82_ab_14__30_), .B(
        u5_mult_82_CARRYB_13__30_), .CI(u5_mult_82_SUMB_13__31_), .CO(
        u5_mult_82_CARRYB_14__30_), .S(u5_mult_82_SUMB_14__30_) );
  FA_X1 u5_mult_82_S2_14_27 ( .A(u5_mult_82_ab_14__27_), .B(
        u5_mult_82_CARRYB_13__27_), .CI(u5_mult_82_SUMB_13__28_), .CO(
        u5_mult_82_CARRYB_14__27_), .S(u5_mult_82_SUMB_14__27_) );
  FA_X1 u5_mult_82_S2_14_24 ( .A(u5_mult_82_ab_14__24_), .B(
        u5_mult_82_CARRYB_13__24_), .CI(u5_mult_82_SUMB_13__25_), .CO(
        u5_mult_82_CARRYB_14__24_), .S(u5_mult_82_SUMB_14__24_) );
  FA_X1 u5_mult_82_S2_14_23 ( .A(u5_mult_82_ab_14__23_), .B(
        u5_mult_82_CARRYB_13__23_), .CI(u5_mult_82_SUMB_13__24_), .CO(
        u5_mult_82_CARRYB_14__23_), .S(u5_mult_82_SUMB_14__23_) );
  FA_X1 u5_mult_82_S2_14_19 ( .A(u5_mult_82_CARRYB_13__19_), .B(
        u5_mult_82_ab_14__19_), .CI(u5_mult_82_SUMB_13__20_), .CO(
        u5_mult_82_CARRYB_14__19_), .S(u5_mult_82_SUMB_14__19_) );
  FA_X1 u5_mult_82_S2_14_18 ( .A(u5_mult_82_ab_14__18_), .B(
        u5_mult_82_CARRYB_13__18_), .CI(u5_mult_82_SUMB_13__19_), .CO(
        u5_mult_82_CARRYB_14__18_), .S(u5_mult_82_SUMB_14__18_) );
  FA_X1 u5_mult_82_S2_14_16 ( .A(u5_mult_82_ab_14__16_), .B(
        u5_mult_82_CARRYB_13__16_), .CI(u5_mult_82_SUMB_13__17_), .CO(
        u5_mult_82_CARRYB_14__16_), .S(u5_mult_82_SUMB_14__16_) );
  FA_X1 u5_mult_82_S2_14_13 ( .A(u5_mult_82_ab_14__13_), .B(
        u5_mult_82_CARRYB_13__13_), .CI(u5_mult_82_SUMB_13__14_), .CO(
        u5_mult_82_CARRYB_14__13_), .S(u5_mult_82_SUMB_14__13_) );
  FA_X1 u5_mult_82_S2_14_12 ( .A(u5_mult_82_ab_14__12_), .B(
        u5_mult_82_CARRYB_13__12_), .CI(u5_mult_82_SUMB_13__13_), .CO(
        u5_mult_82_CARRYB_14__12_), .S(u5_mult_82_SUMB_14__12_) );
  FA_X1 u5_mult_82_S2_14_11 ( .A(u5_mult_82_ab_14__11_), .B(
        u5_mult_82_CARRYB_13__11_), .CI(u5_mult_82_SUMB_13__12_), .CO(
        u5_mult_82_CARRYB_14__11_), .S(u5_mult_82_SUMB_14__11_) );
  FA_X1 u5_mult_82_S2_14_10 ( .A(u5_mult_82_ab_14__10_), .B(
        u5_mult_82_CARRYB_13__10_), .CI(u5_mult_82_SUMB_13__11_), .CO(
        u5_mult_82_CARRYB_14__10_), .S(u5_mult_82_SUMB_14__10_) );
  FA_X1 u5_mult_82_S2_14_9 ( .A(u5_mult_82_ab_14__9_), .B(
        u5_mult_82_CARRYB_13__9_), .CI(u5_mult_82_SUMB_13__10_), .CO(
        u5_mult_82_CARRYB_14__9_), .S(u5_mult_82_SUMB_14__9_) );
  FA_X1 u5_mult_82_S2_14_8 ( .A(u5_mult_82_ab_14__8_), .B(
        u5_mult_82_CARRYB_13__8_), .CI(u5_mult_82_SUMB_13__9_), .CO(
        u5_mult_82_CARRYB_14__8_), .S(u5_mult_82_SUMB_14__8_) );
  FA_X1 u5_mult_82_S2_14_7 ( .A(u5_mult_82_ab_14__7_), .B(
        u5_mult_82_CARRYB_13__7_), .CI(u5_mult_82_SUMB_13__8_), .CO(
        u5_mult_82_CARRYB_14__7_), .S(u5_mult_82_SUMB_14__7_) );
  FA_X1 u5_mult_82_S2_14_6 ( .A(u5_mult_82_ab_14__6_), .B(
        u5_mult_82_CARRYB_13__6_), .CI(u5_mult_82_SUMB_13__7_), .CO(
        u5_mult_82_CARRYB_14__6_), .S(u5_mult_82_SUMB_14__6_) );
  FA_X1 u5_mult_82_S2_14_5 ( .A(u5_mult_82_ab_14__5_), .B(
        u5_mult_82_CARRYB_13__5_), .CI(u5_mult_82_SUMB_13__6_), .CO(
        u5_mult_82_CARRYB_14__5_), .S(u5_mult_82_SUMB_14__5_) );
  FA_X1 u5_mult_82_S2_14_4 ( .A(u5_mult_82_ab_14__4_), .B(
        u5_mult_82_CARRYB_13__4_), .CI(u5_mult_82_SUMB_13__5_), .CO(
        u5_mult_82_CARRYB_14__4_), .S(u5_mult_82_SUMB_14__4_) );
  FA_X1 u5_mult_82_S2_14_3 ( .A(u5_mult_82_ab_14__3_), .B(
        u5_mult_82_CARRYB_13__3_), .CI(u5_mult_82_SUMB_13__4_), .CO(
        u5_mult_82_CARRYB_14__3_), .S(u5_mult_82_SUMB_14__3_) );
  FA_X1 u5_mult_82_S2_14_2 ( .A(u5_mult_82_ab_14__2_), .B(
        u5_mult_82_CARRYB_13__2_), .CI(u5_mult_82_SUMB_13__3_), .CO(
        u5_mult_82_CARRYB_14__2_), .S(u5_mult_82_SUMB_14__2_) );
  FA_X1 u5_mult_82_S2_14_1 ( .A(u5_mult_82_ab_14__1_), .B(
        u5_mult_82_CARRYB_13__1_), .CI(u5_mult_82_SUMB_13__2_), .CO(
        u5_mult_82_CARRYB_14__1_), .S(u5_mult_82_SUMB_14__1_) );
  FA_X1 u5_mult_82_S1_14_0 ( .A(u5_mult_82_ab_14__0_), .B(
        u5_mult_82_CARRYB_13__0_), .CI(u5_mult_82_SUMB_13__1_), .CO(
        u5_mult_82_CARRYB_14__0_), .S(u5_N14) );
  FA_X1 u5_mult_82_S3_15_51 ( .A(u5_mult_82_ab_15__51_), .B(
        u5_mult_82_CARRYB_14__51_), .CI(u5_mult_82_ab_14__52_), .CO(
        u5_mult_82_CARRYB_15__51_), .S(u5_mult_82_SUMB_15__51_) );
  FA_X1 u5_mult_82_S2_15_44 ( .A(u5_mult_82_ab_15__44_), .B(
        u5_mult_82_CARRYB_14__44_), .CI(u5_mult_82_SUMB_14__45_), .CO(
        u5_mult_82_CARRYB_15__44_), .S(u5_mult_82_SUMB_15__44_) );
  FA_X1 u5_mult_82_S2_15_41 ( .A(u5_mult_82_ab_15__41_), .B(
        u5_mult_82_CARRYB_14__41_), .CI(u5_mult_82_SUMB_14__42_), .CO(
        u5_mult_82_CARRYB_15__41_), .S(u5_mult_82_SUMB_15__41_) );
  FA_X1 u5_mult_82_S2_15_32 ( .A(u5_mult_82_ab_15__32_), .B(
        u5_mult_82_CARRYB_14__32_), .CI(u5_mult_82_SUMB_14__33_), .CO(
        u5_mult_82_CARRYB_15__32_), .S(u5_mult_82_SUMB_15__32_) );
  FA_X1 u5_mult_82_S2_15_26 ( .A(u5_mult_82_ab_15__26_), .B(
        u5_mult_82_CARRYB_14__26_), .CI(u5_mult_82_SUMB_14__27_), .CO(
        u5_mult_82_CARRYB_15__26_), .S(u5_mult_82_SUMB_15__26_) );
  FA_X1 u5_mult_82_S2_15_25 ( .A(u5_mult_82_ab_15__25_), .B(
        u5_mult_82_CARRYB_14__25_), .CI(u5_mult_82_SUMB_14__26_), .CO(
        u5_mult_82_CARRYB_15__25_), .S(u5_mult_82_SUMB_15__25_) );
  FA_X1 u5_mult_82_S2_15_22 ( .A(u5_mult_82_ab_15__22_), .B(
        u5_mult_82_CARRYB_14__22_), .CI(u5_mult_82_SUMB_14__23_), .CO(
        u5_mult_82_CARRYB_15__22_), .S(u5_mult_82_SUMB_15__22_) );
  FA_X1 u5_mult_82_S2_15_21 ( .A(u5_mult_82_ab_15__21_), .B(
        u5_mult_82_CARRYB_14__21_), .CI(u5_mult_82_SUMB_14__22_), .CO(
        u5_mult_82_CARRYB_15__21_), .S(u5_mult_82_SUMB_15__21_) );
  FA_X1 u5_mult_82_S2_15_20 ( .A(u5_mult_82_ab_15__20_), .B(
        u5_mult_82_CARRYB_14__20_), .CI(u5_mult_82_SUMB_14__21_), .CO(
        u5_mult_82_CARRYB_15__20_), .S(u5_mult_82_SUMB_15__20_) );
  FA_X1 u5_mult_82_S2_15_19 ( .A(u5_mult_82_ab_15__19_), .B(
        u5_mult_82_CARRYB_14__19_), .CI(u5_mult_82_SUMB_14__20_), .CO(
        u5_mult_82_CARRYB_15__19_), .S(u5_mult_82_SUMB_15__19_) );
  FA_X1 u5_mult_82_S2_15_18 ( .A(u5_mult_82_ab_15__18_), .B(
        u5_mult_82_CARRYB_14__18_), .CI(u5_mult_82_SUMB_14__19_), .CO(
        u5_mult_82_CARRYB_15__18_), .S(u5_mult_82_SUMB_15__18_) );
  FA_X1 u5_mult_82_S2_15_17 ( .A(u5_mult_82_ab_15__17_), .B(
        u5_mult_82_CARRYB_14__17_), .CI(u5_mult_82_SUMB_14__18_), .CO(
        u5_mult_82_CARRYB_15__17_), .S(u5_mult_82_SUMB_15__17_) );
  FA_X1 u5_mult_82_S2_15_16 ( .A(u5_mult_82_ab_15__16_), .B(
        u5_mult_82_CARRYB_14__16_), .CI(u5_mult_82_SUMB_14__17_), .CO(
        u5_mult_82_CARRYB_15__16_), .S(u5_mult_82_SUMB_15__16_) );
  FA_X1 u5_mult_82_S2_15_15 ( .A(u5_mult_82_ab_15__15_), .B(
        u5_mult_82_CARRYB_14__15_), .CI(u5_mult_82_SUMB_14__16_), .CO(
        u5_mult_82_CARRYB_15__15_), .S(u5_mult_82_SUMB_15__15_) );
  FA_X1 u5_mult_82_S2_15_12 ( .A(u5_mult_82_ab_15__12_), .B(
        u5_mult_82_CARRYB_14__12_), .CI(u5_mult_82_SUMB_14__13_), .CO(
        u5_mult_82_CARRYB_15__12_), .S(u5_mult_82_SUMB_15__12_) );
  FA_X1 u5_mult_82_S2_15_11 ( .A(u5_mult_82_ab_15__11_), .B(
        u5_mult_82_CARRYB_14__11_), .CI(u5_mult_82_SUMB_14__12_), .CO(
        u5_mult_82_CARRYB_15__11_), .S(u5_mult_82_SUMB_15__11_) );
  FA_X1 u5_mult_82_S2_15_9 ( .A(u5_mult_82_ab_15__9_), .B(
        u5_mult_82_CARRYB_14__9_), .CI(u5_mult_82_SUMB_14__10_), .CO(
        u5_mult_82_CARRYB_15__9_), .S(u5_mult_82_SUMB_15__9_) );
  FA_X1 u5_mult_82_S2_15_8 ( .A(u5_mult_82_ab_15__8_), .B(
        u5_mult_82_CARRYB_14__8_), .CI(u5_mult_82_SUMB_14__9_), .CO(
        u5_mult_82_CARRYB_15__8_), .S(u5_mult_82_SUMB_15__8_) );
  FA_X1 u5_mult_82_S2_15_7 ( .A(u5_mult_82_ab_15__7_), .B(
        u5_mult_82_CARRYB_14__7_), .CI(u5_mult_82_SUMB_14__8_), .CO(
        u5_mult_82_CARRYB_15__7_), .S(u5_mult_82_SUMB_15__7_) );
  FA_X1 u5_mult_82_S2_15_6 ( .A(u5_mult_82_ab_15__6_), .B(
        u5_mult_82_CARRYB_14__6_), .CI(u5_mult_82_SUMB_14__7_), .CO(
        u5_mult_82_CARRYB_15__6_), .S(u5_mult_82_SUMB_15__6_) );
  FA_X1 u5_mult_82_S2_15_5 ( .A(u5_mult_82_ab_15__5_), .B(
        u5_mult_82_CARRYB_14__5_), .CI(u5_mult_82_SUMB_14__6_), .CO(
        u5_mult_82_CARRYB_15__5_), .S(u5_mult_82_SUMB_15__5_) );
  FA_X1 u5_mult_82_S2_15_4 ( .A(u5_mult_82_ab_15__4_), .B(
        u5_mult_82_CARRYB_14__4_), .CI(u5_mult_82_SUMB_14__5_), .CO(
        u5_mult_82_CARRYB_15__4_), .S(u5_mult_82_SUMB_15__4_) );
  FA_X1 u5_mult_82_S2_15_3 ( .A(u5_mult_82_ab_15__3_), .B(
        u5_mult_82_CARRYB_14__3_), .CI(u5_mult_82_SUMB_14__4_), .CO(
        u5_mult_82_CARRYB_15__3_), .S(u5_mult_82_SUMB_15__3_) );
  FA_X1 u5_mult_82_S2_15_2 ( .A(u5_mult_82_ab_15__2_), .B(
        u5_mult_82_CARRYB_14__2_), .CI(u5_mult_82_SUMB_14__3_), .CO(
        u5_mult_82_CARRYB_15__2_), .S(u5_mult_82_SUMB_15__2_) );
  FA_X1 u5_mult_82_S2_15_1 ( .A(u5_mult_82_ab_15__1_), .B(
        u5_mult_82_CARRYB_14__1_), .CI(u5_mult_82_SUMB_14__2_), .CO(
        u5_mult_82_CARRYB_15__1_), .S(u5_mult_82_SUMB_15__1_) );
  FA_X1 u5_mult_82_S1_15_0 ( .A(u5_mult_82_ab_15__0_), .B(
        u5_mult_82_CARRYB_14__0_), .CI(u5_mult_82_SUMB_14__1_), .CO(
        u5_mult_82_CARRYB_15__0_), .S(u5_N15) );
  FA_X1 u5_mult_82_S3_16_51 ( .A(u5_mult_82_ab_16__51_), .B(
        u5_mult_82_CARRYB_15__51_), .CI(u5_mult_82_ab_15__52_), .CO(
        u5_mult_82_CARRYB_16__51_), .S(u5_mult_82_SUMB_16__51_) );
  FA_X1 u5_mult_82_S2_16_50 ( .A(u5_mult_82_ab_16__50_), .B(
        u5_mult_82_CARRYB_15__50_), .CI(u5_mult_82_SUMB_15__51_), .CO(
        u5_mult_82_CARRYB_16__50_), .S(u5_mult_82_SUMB_16__50_) );
  FA_X1 u5_mult_82_S2_16_48 ( .A(u5_mult_82_ab_16__48_), .B(
        u5_mult_82_CARRYB_15__48_), .CI(u5_mult_82_SUMB_15__49_), .CO(
        u5_mult_82_CARRYB_16__48_), .S(u5_mult_82_SUMB_16__48_) );
  FA_X1 u5_mult_82_S2_16_47 ( .A(u5_mult_82_ab_16__47_), .B(
        u5_mult_82_CARRYB_15__47_), .CI(u5_mult_82_SUMB_15__48_), .CO(
        u5_mult_82_CARRYB_16__47_), .S(u5_mult_82_SUMB_16__47_) );
  FA_X1 u5_mult_82_S2_16_39 ( .A(u5_mult_82_CARRYB_15__39_), .B(
        u5_mult_82_ab_16__39_), .CI(u5_mult_82_SUMB_15__40_), .CO(
        u5_mult_82_CARRYB_16__39_), .S(u5_mult_82_SUMB_16__39_) );
  FA_X1 u5_mult_82_S2_16_30 ( .A(u5_mult_82_ab_16__30_), .B(
        u5_mult_82_CARRYB_15__30_), .CI(u5_mult_82_SUMB_15__31_), .CO(
        u5_mult_82_CARRYB_16__30_), .S(u5_mult_82_SUMB_16__30_) );
  FA_X1 u5_mult_82_S2_16_23 ( .A(u5_mult_82_ab_16__23_), .B(
        u5_mult_82_SUMB_15__24_), .CI(u5_mult_82_CARRYB_15__23_), .CO(
        u5_mult_82_CARRYB_16__23_), .S(u5_mult_82_SUMB_16__23_) );
  FA_X1 u5_mult_82_S2_16_22 ( .A(u5_mult_82_ab_16__22_), .B(
        u5_mult_82_CARRYB_15__22_), .CI(u5_mult_82_SUMB_15__23_), .CO(
        u5_mult_82_CARRYB_16__22_), .S(u5_mult_82_SUMB_16__22_) );
  FA_X1 u5_mult_82_S2_16_21 ( .A(u5_mult_82_ab_16__21_), .B(
        u5_mult_82_CARRYB_15__21_), .CI(u5_mult_82_SUMB_15__22_), .CO(
        u5_mult_82_CARRYB_16__21_), .S(u5_mult_82_SUMB_16__21_) );
  FA_X1 u5_mult_82_S2_16_18 ( .A(u5_mult_82_ab_16__18_), .B(
        u5_mult_82_CARRYB_15__18_), .CI(u5_mult_82_SUMB_15__19_), .CO(
        u5_mult_82_CARRYB_16__18_), .S(u5_mult_82_SUMB_16__18_) );
  FA_X1 u5_mult_82_S2_16_17 ( .A(u5_mult_82_ab_16__17_), .B(
        u5_mult_82_CARRYB_15__17_), .CI(u5_mult_82_SUMB_15__18_), .CO(
        u5_mult_82_CARRYB_16__17_), .S(u5_mult_82_SUMB_16__17_) );
  FA_X1 u5_mult_82_S2_16_14 ( .A(u5_mult_82_ab_16__14_), .B(
        u5_mult_82_CARRYB_15__14_), .CI(u5_mult_82_SUMB_15__15_), .CO(
        u5_mult_82_CARRYB_16__14_), .S(u5_mult_82_SUMB_16__14_) );
  FA_X1 u5_mult_82_S2_16_13 ( .A(u5_mult_82_ab_16__13_), .B(
        u5_mult_82_CARRYB_15__13_), .CI(u5_mult_82_SUMB_15__14_), .CO(
        u5_mult_82_CARRYB_16__13_), .S(u5_mult_82_SUMB_16__13_) );
  FA_X1 u5_mult_82_S2_16_11 ( .A(u5_mult_82_ab_16__11_), .B(
        u5_mult_82_CARRYB_15__11_), .CI(u5_mult_82_SUMB_15__12_), .CO(
        u5_mult_82_CARRYB_16__11_), .S(u5_mult_82_SUMB_16__11_) );
  FA_X1 u5_mult_82_S2_16_10 ( .A(u5_mult_82_ab_16__10_), .B(
        u5_mult_82_CARRYB_15__10_), .CI(u5_mult_82_SUMB_15__11_), .CO(
        u5_mult_82_CARRYB_16__10_), .S(u5_mult_82_SUMB_16__10_) );
  FA_X1 u5_mult_82_S2_16_8 ( .A(u5_mult_82_ab_16__8_), .B(
        u5_mult_82_CARRYB_15__8_), .CI(u5_mult_82_SUMB_15__9_), .CO(
        u5_mult_82_CARRYB_16__8_), .S(u5_mult_82_SUMB_16__8_) );
  FA_X1 u5_mult_82_S2_16_7 ( .A(u5_mult_82_ab_16__7_), .B(
        u5_mult_82_CARRYB_15__7_), .CI(u5_mult_82_SUMB_15__8_), .CO(
        u5_mult_82_CARRYB_16__7_), .S(u5_mult_82_SUMB_16__7_) );
  FA_X1 u5_mult_82_S2_16_6 ( .A(u5_mult_82_ab_16__6_), .B(
        u5_mult_82_CARRYB_15__6_), .CI(u5_mult_82_SUMB_15__7_), .CO(
        u5_mult_82_CARRYB_16__6_), .S(u5_mult_82_SUMB_16__6_) );
  FA_X1 u5_mult_82_S2_16_5 ( .A(u5_mult_82_ab_16__5_), .B(
        u5_mult_82_CARRYB_15__5_), .CI(u5_mult_82_SUMB_15__6_), .CO(
        u5_mult_82_CARRYB_16__5_), .S(u5_mult_82_SUMB_16__5_) );
  FA_X1 u5_mult_82_S2_16_4 ( .A(u5_mult_82_ab_16__4_), .B(
        u5_mult_82_CARRYB_15__4_), .CI(u5_mult_82_SUMB_15__5_), .CO(
        u5_mult_82_CARRYB_16__4_), .S(u5_mult_82_SUMB_16__4_) );
  FA_X1 u5_mult_82_S2_16_3 ( .A(u5_mult_82_ab_16__3_), .B(
        u5_mult_82_CARRYB_15__3_), .CI(u5_mult_82_SUMB_15__4_), .CO(
        u5_mult_82_CARRYB_16__3_), .S(u5_mult_82_SUMB_16__3_) );
  FA_X1 u5_mult_82_S2_16_2 ( .A(u5_mult_82_ab_16__2_), .B(
        u5_mult_82_CARRYB_15__2_), .CI(u5_mult_82_SUMB_15__3_), .CO(
        u5_mult_82_CARRYB_16__2_), .S(u5_mult_82_SUMB_16__2_) );
  FA_X1 u5_mult_82_S2_16_1 ( .A(u5_mult_82_ab_16__1_), .B(
        u5_mult_82_CARRYB_15__1_), .CI(u5_mult_82_SUMB_15__2_), .CO(
        u5_mult_82_CARRYB_16__1_), .S(u5_mult_82_SUMB_16__1_) );
  FA_X1 u5_mult_82_S1_16_0 ( .A(u5_mult_82_ab_16__0_), .B(
        u5_mult_82_CARRYB_15__0_), .CI(u5_mult_82_SUMB_15__1_), .CO(
        u5_mult_82_CARRYB_16__0_), .S(u5_N16) );
  FA_X1 u5_mult_82_S3_17_51 ( .A(u5_mult_82_ab_17__51_), .B(
        u5_mult_82_ab_16__52_), .CI(u5_mult_82_CARRYB_16__51_), .CO(
        u5_mult_82_CARRYB_17__51_), .S(u5_mult_82_SUMB_17__51_) );
  FA_X1 u5_mult_82_S2_17_49 ( .A(u5_mult_82_CARRYB_16__49_), .B(
        u5_mult_82_ab_17__49_), .CI(u5_mult_82_SUMB_16__50_), .CO(
        u5_mult_82_CARRYB_17__49_), .S(u5_mult_82_SUMB_17__49_) );
  FA_X1 u5_mult_82_S2_17_46 ( .A(u5_mult_82_ab_17__46_), .B(
        u5_mult_82_CARRYB_16__46_), .CI(u5_mult_82_SUMB_16__47_), .CO(
        u5_mult_82_CARRYB_17__46_), .S(u5_mult_82_SUMB_17__46_) );
  FA_X1 u5_mult_82_S2_17_43 ( .A(u5_mult_82_CARRYB_16__43_), .B(
        u5_mult_82_ab_17__43_), .CI(u5_mult_82_SUMB_16__44_), .CO(
        u5_mult_82_CARRYB_17__43_), .S(u5_mult_82_SUMB_17__43_) );
  FA_X1 u5_mult_82_S2_17_40 ( .A(u5_mult_82_ab_17__40_), .B(
        u5_mult_82_CARRYB_16__40_), .CI(u5_mult_82_SUMB_16__41_), .CO(
        u5_mult_82_CARRYB_17__40_), .S(u5_mult_82_SUMB_17__40_) );
  FA_X1 u5_mult_82_S2_17_39 ( .A(u5_mult_82_ab_17__39_), .B(
        u5_mult_82_CARRYB_16__39_), .CI(u5_mult_82_SUMB_16__40_), .CO(
        u5_mult_82_CARRYB_17__39_), .S(u5_mult_82_SUMB_17__39_) );
  FA_X1 u5_mult_82_S2_17_34 ( .A(u5_mult_82_ab_17__34_), .B(
        u5_mult_82_CARRYB_16__34_), .CI(u5_mult_82_SUMB_16__35_), .CO(
        u5_mult_82_CARRYB_17__34_), .S(u5_mult_82_SUMB_17__34_) );
  FA_X1 u5_mult_82_S2_17_33 ( .A(u5_mult_82_ab_17__33_), .B(
        u5_mult_82_CARRYB_16__33_), .CI(u5_mult_82_SUMB_16__34_), .CO(
        u5_mult_82_CARRYB_17__33_), .S(u5_mult_82_SUMB_17__33_) );
  FA_X1 u5_mult_82_S2_17_30 ( .A(u5_mult_82_CARRYB_16__30_), .B(
        u5_mult_82_ab_17__30_), .CI(u5_mult_82_SUMB_16__31_), .CO(
        u5_mult_82_CARRYB_17__30_), .S(u5_mult_82_SUMB_17__30_) );
  FA_X1 u5_mult_82_S2_17_29 ( .A(u5_mult_82_ab_17__29_), .B(
        u5_mult_82_CARRYB_16__29_), .CI(u5_mult_82_SUMB_16__30_), .CO(
        u5_mult_82_CARRYB_17__29_), .S(u5_mult_82_SUMB_17__29_) );
  FA_X1 u5_mult_82_S2_17_22 ( .A(u5_mult_82_ab_17__22_), .B(
        u5_mult_82_CARRYB_16__22_), .CI(u5_mult_82_SUMB_16__23_), .CO(
        u5_mult_82_CARRYB_17__22_), .S(u5_mult_82_SUMB_17__22_) );
  FA_X1 u5_mult_82_S2_17_13 ( .A(u5_mult_82_ab_17__13_), .B(
        u5_mult_82_CARRYB_16__13_), .CI(u5_mult_82_SUMB_16__14_), .CO(
        u5_mult_82_CARRYB_17__13_), .S(u5_mult_82_SUMB_17__13_) );
  FA_X1 u5_mult_82_S2_17_12 ( .A(u5_mult_82_ab_17__12_), .B(
        u5_mult_82_CARRYB_16__12_), .CI(u5_mult_82_SUMB_16__13_), .CO(
        u5_mult_82_CARRYB_17__12_), .S(u5_mult_82_SUMB_17__12_) );
  FA_X1 u5_mult_82_S2_17_11 ( .A(u5_mult_82_CARRYB_16__11_), .B(
        u5_mult_82_ab_17__11_), .CI(u5_mult_82_SUMB_16__12_), .CO(
        u5_mult_82_CARRYB_17__11_), .S(u5_mult_82_SUMB_17__11_) );
  FA_X1 u5_mult_82_S2_17_9 ( .A(u5_mult_82_ab_17__9_), .B(
        u5_mult_82_CARRYB_16__9_), .CI(u5_mult_82_SUMB_16__10_), .CO(
        u5_mult_82_CARRYB_17__9_), .S(u5_mult_82_SUMB_17__9_) );
  FA_X1 u5_mult_82_S2_17_8 ( .A(u5_mult_82_ab_17__8_), .B(
        u5_mult_82_CARRYB_16__8_), .CI(u5_mult_82_SUMB_16__9_), .CO(
        u5_mult_82_CARRYB_17__8_), .S(u5_mult_82_SUMB_17__8_) );
  FA_X1 u5_mult_82_S2_17_6 ( .A(u5_mult_82_ab_17__6_), .B(
        u5_mult_82_CARRYB_16__6_), .CI(u5_mult_82_SUMB_16__7_), .CO(
        u5_mult_82_CARRYB_17__6_), .S(u5_mult_82_SUMB_17__6_) );
  FA_X1 u5_mult_82_S2_17_5 ( .A(u5_mult_82_ab_17__5_), .B(
        u5_mult_82_CARRYB_16__5_), .CI(u5_mult_82_SUMB_16__6_), .CO(
        u5_mult_82_CARRYB_17__5_), .S(u5_mult_82_SUMB_17__5_) );
  FA_X1 u5_mult_82_S2_17_4 ( .A(u5_mult_82_ab_17__4_), .B(
        u5_mult_82_CARRYB_16__4_), .CI(u5_mult_82_SUMB_16__5_), .CO(
        u5_mult_82_CARRYB_17__4_), .S(u5_mult_82_SUMB_17__4_) );
  FA_X1 u5_mult_82_S2_17_3 ( .A(u5_mult_82_ab_17__3_), .B(
        u5_mult_82_CARRYB_16__3_), .CI(u5_mult_82_SUMB_16__4_), .CO(
        u5_mult_82_CARRYB_17__3_), .S(u5_mult_82_SUMB_17__3_) );
  FA_X1 u5_mult_82_S2_17_2 ( .A(u5_mult_82_ab_17__2_), .B(
        u5_mult_82_CARRYB_16__2_), .CI(u5_mult_82_SUMB_16__3_), .CO(
        u5_mult_82_CARRYB_17__2_), .S(u5_mult_82_SUMB_17__2_) );
  FA_X1 u5_mult_82_S2_17_1 ( .A(u5_mult_82_ab_17__1_), .B(
        u5_mult_82_CARRYB_16__1_), .CI(u5_mult_82_SUMB_16__2_), .CO(
        u5_mult_82_CARRYB_17__1_), .S(u5_mult_82_SUMB_17__1_) );
  FA_X1 u5_mult_82_S1_17_0 ( .A(u5_mult_82_ab_17__0_), .B(
        u5_mult_82_CARRYB_16__0_), .CI(u5_mult_82_SUMB_16__1_), .CO(
        u5_mult_82_CARRYB_17__0_), .S(u5_N17) );
  FA_X1 u5_mult_82_S3_18_51 ( .A(u5_mult_82_ab_18__51_), .B(
        u5_mult_82_CARRYB_17__51_), .CI(u5_mult_82_ab_17__52_), .CO(
        u5_mult_82_CARRYB_18__51_), .S(u5_mult_82_SUMB_18__51_) );
  FA_X1 u5_mult_82_S2_18_48 ( .A(u5_mult_82_CARRYB_17__48_), .B(
        u5_mult_82_ab_18__48_), .CI(u5_mult_82_SUMB_17__49_), .CO(
        u5_mult_82_CARRYB_18__48_), .S(u5_mult_82_SUMB_18__48_) );
  FA_X1 u5_mult_82_S2_18_44 ( .A(u5_mult_82_ab_18__44_), .B(
        u5_mult_82_CARRYB_17__44_), .CI(u5_mult_82_SUMB_17__45_), .CO(
        u5_mult_82_CARRYB_18__44_), .S(u5_mult_82_SUMB_18__44_) );
  FA_X1 u5_mult_82_S2_18_42 ( .A(u5_mult_82_ab_18__42_), .B(
        u5_mult_82_CARRYB_17__42_), .CI(u5_mult_82_SUMB_17__43_), .CO(
        u5_mult_82_CARRYB_18__42_), .S(u5_mult_82_SUMB_18__42_) );
  FA_X1 u5_mult_82_S2_18_41 ( .A(u5_mult_82_ab_18__41_), .B(
        u5_mult_82_CARRYB_17__41_), .CI(u5_mult_82_SUMB_17__42_), .CO(
        u5_mult_82_CARRYB_18__41_), .S(u5_mult_82_SUMB_18__41_) );
  FA_X1 u5_mult_82_S2_18_40 ( .A(u5_mult_82_CARRYB_17__40_), .B(
        u5_mult_82_ab_18__40_), .CI(u5_mult_82_SUMB_17__41_), .CO(
        u5_mult_82_CARRYB_18__40_), .S(u5_mult_82_SUMB_18__40_) );
  FA_X1 u5_mult_82_S2_18_34 ( .A(u5_mult_82_ab_18__34_), .B(
        u5_mult_82_CARRYB_17__34_), .CI(u5_mult_82_SUMB_17__35_), .CO(
        u5_mult_82_CARRYB_18__34_), .S(u5_mult_82_SUMB_18__34_) );
  FA_X1 u5_mult_82_S2_18_32 ( .A(u5_mult_82_ab_18__32_), .B(
        u5_mult_82_CARRYB_17__32_), .CI(u5_mult_82_SUMB_17__33_), .CO(
        u5_mult_82_CARRYB_18__32_), .S(u5_mult_82_SUMB_18__32_) );
  FA_X1 u5_mult_82_S2_18_31 ( .A(u5_mult_82_ab_18__31_), .B(
        u5_mult_82_CARRYB_17__31_), .CI(u5_mult_82_SUMB_17__32_), .CO(
        u5_mult_82_CARRYB_18__31_), .S(u5_mult_82_SUMB_18__31_) );
  FA_X1 u5_mult_82_S2_18_24 ( .A(u5_mult_82_ab_18__24_), .B(
        u5_mult_82_CARRYB_17__24_), .CI(u5_mult_82_SUMB_17__25_), .CO(
        u5_mult_82_CARRYB_18__24_), .S(u5_mult_82_SUMB_18__24_) );
  FA_X1 u5_mult_82_S2_18_22 ( .A(u5_mult_82_ab_18__22_), .B(
        u5_mult_82_CARRYB_17__22_), .CI(u5_mult_82_SUMB_17__23_), .CO(
        u5_mult_82_CARRYB_18__22_), .S(u5_mult_82_SUMB_18__22_) );
  FA_X1 u5_mult_82_S2_18_21 ( .A(u5_mult_82_ab_18__21_), .B(
        u5_mult_82_CARRYB_17__21_), .CI(u5_mult_82_SUMB_17__22_), .CO(
        u5_mult_82_CARRYB_18__21_), .S(u5_mult_82_SUMB_18__21_) );
  FA_X1 u5_mult_82_S2_18_19 ( .A(u5_mult_82_ab_18__19_), .B(
        u5_mult_82_CARRYB_17__19_), .CI(u5_mult_82_SUMB_17__20_), .CO(
        u5_mult_82_CARRYB_18__19_), .S(u5_mult_82_SUMB_18__19_) );
  FA_X1 u5_mult_82_S2_18_18 ( .A(u5_mult_82_CARRYB_17__18_), .B(
        u5_mult_82_ab_18__18_), .CI(u5_mult_82_SUMB_17__19_), .CO(
        u5_mult_82_CARRYB_18__18_), .S(u5_mult_82_SUMB_18__18_) );
  FA_X1 u5_mult_82_S2_18_17 ( .A(u5_mult_82_ab_18__17_), .B(
        u5_mult_82_CARRYB_17__17_), .CI(u5_mult_82_SUMB_17__18_), .CO(
        u5_mult_82_CARRYB_18__17_), .S(u5_mult_82_SUMB_18__17_) );
  FA_X1 u5_mult_82_S2_18_14 ( .A(u5_mult_82_CARRYB_17__14_), .B(
        u5_mult_82_ab_18__14_), .CI(u5_mult_82_SUMB_17__15_), .CO(
        u5_mult_82_CARRYB_18__14_), .S(u5_mult_82_SUMB_18__14_) );
  FA_X1 u5_mult_82_S2_18_11 ( .A(u5_mult_82_ab_18__11_), .B(
        u5_mult_82_CARRYB_17__11_), .CI(u5_mult_82_SUMB_17__12_), .CO(
        u5_mult_82_CARRYB_18__11_), .S(u5_mult_82_SUMB_18__11_) );
  FA_X1 u5_mult_82_S2_18_10 ( .A(u5_mult_82_ab_18__10_), .B(
        u5_mult_82_CARRYB_17__10_), .CI(u5_mult_82_SUMB_17__11_), .CO(
        u5_mult_82_CARRYB_18__10_), .S(u5_mult_82_SUMB_18__10_) );
  FA_X1 u5_mult_82_S2_18_9 ( .A(u5_mult_82_ab_18__9_), .B(
        u5_mult_82_CARRYB_17__9_), .CI(u5_mult_82_SUMB_17__10_), .CO(
        u5_mult_82_CARRYB_18__9_), .S(u5_mult_82_SUMB_18__9_) );
  FA_X1 u5_mult_82_S2_18_8 ( .A(u5_mult_82_ab_18__8_), .B(
        u5_mult_82_CARRYB_17__8_), .CI(u5_mult_82_SUMB_17__9_), .CO(
        u5_mult_82_CARRYB_18__8_), .S(u5_mult_82_SUMB_18__8_) );
  FA_X1 u5_mult_82_S2_18_7 ( .A(u5_mult_82_ab_18__7_), .B(
        u5_mult_82_CARRYB_17__7_), .CI(u5_mult_82_SUMB_17__8_), .CO(
        u5_mult_82_CARRYB_18__7_), .S(u5_mult_82_SUMB_18__7_) );
  FA_X1 u5_mult_82_S2_18_6 ( .A(u5_mult_82_ab_18__6_), .B(
        u5_mult_82_CARRYB_17__6_), .CI(u5_mult_82_SUMB_17__7_), .CO(
        u5_mult_82_CARRYB_18__6_), .S(u5_mult_82_SUMB_18__6_) );
  FA_X1 u5_mult_82_S2_18_5 ( .A(u5_mult_82_ab_18__5_), .B(
        u5_mult_82_CARRYB_17__5_), .CI(u5_mult_82_SUMB_17__6_), .CO(
        u5_mult_82_CARRYB_18__5_), .S(u5_mult_82_SUMB_18__5_) );
  FA_X1 u5_mult_82_S2_18_4 ( .A(u5_mult_82_ab_18__4_), .B(
        u5_mult_82_CARRYB_17__4_), .CI(u5_mult_82_SUMB_17__5_), .CO(
        u5_mult_82_CARRYB_18__4_), .S(u5_mult_82_SUMB_18__4_) );
  FA_X1 u5_mult_82_S2_18_3 ( .A(u5_mult_82_ab_18__3_), .B(
        u5_mult_82_CARRYB_17__3_), .CI(u5_mult_82_SUMB_17__4_), .CO(
        u5_mult_82_CARRYB_18__3_), .S(u5_mult_82_SUMB_18__3_) );
  FA_X1 u5_mult_82_S2_18_2 ( .A(u5_mult_82_ab_18__2_), .B(
        u5_mult_82_CARRYB_17__2_), .CI(u5_mult_82_SUMB_17__3_), .CO(
        u5_mult_82_CARRYB_18__2_), .S(u5_mult_82_SUMB_18__2_) );
  FA_X1 u5_mult_82_S2_18_1 ( .A(u5_mult_82_ab_18__1_), .B(
        u5_mult_82_CARRYB_17__1_), .CI(u5_mult_82_SUMB_17__2_), .CO(
        u5_mult_82_CARRYB_18__1_), .S(u5_mult_82_SUMB_18__1_) );
  FA_X1 u5_mult_82_S1_18_0 ( .A(u5_mult_82_ab_18__0_), .B(
        u5_mult_82_CARRYB_17__0_), .CI(u5_mult_82_SUMB_17__1_), .CO(
        u5_mult_82_CARRYB_18__0_), .S(u5_N18) );
  FA_X1 u5_mult_82_S3_19_51 ( .A(u5_mult_82_ab_19__51_), .B(
        u5_mult_82_CARRYB_18__51_), .CI(u5_mult_82_ab_18__52_), .CO(
        u5_mult_82_CARRYB_19__51_), .S(u5_mult_82_SUMB_19__51_) );
  FA_X1 u5_mult_82_S2_19_50 ( .A(u5_mult_82_ab_19__50_), .B(
        u5_mult_82_CARRYB_18__50_), .CI(u5_mult_82_SUMB_18__51_), .CO(
        u5_mult_82_CARRYB_19__50_), .S(u5_mult_82_SUMB_19__50_) );
  FA_X1 u5_mult_82_S2_19_48 ( .A(u5_mult_82_ab_19__48_), .B(
        u5_mult_82_CARRYB_18__48_), .CI(u5_mult_82_SUMB_18__49_), .CO(
        u5_mult_82_CARRYB_19__48_), .S(u5_mult_82_SUMB_19__48_) );
  FA_X1 u5_mult_82_S2_19_42 ( .A(u5_mult_82_ab_19__42_), .B(
        u5_mult_82_CARRYB_18__42_), .CI(u5_mult_82_SUMB_18__43_), .CO(
        u5_mult_82_CARRYB_19__42_), .S(u5_mult_82_SUMB_19__42_) );
  FA_X1 u5_mult_82_S2_19_41 ( .A(u5_mult_82_ab_19__41_), .B(
        u5_mult_82_CARRYB_18__41_), .CI(u5_mult_82_SUMB_18__42_), .CO(
        u5_mult_82_CARRYB_19__41_), .S(u5_mult_82_SUMB_19__41_) );
  FA_X1 u5_mult_82_S2_19_39 ( .A(u5_mult_82_ab_19__39_), .B(
        u5_mult_82_CARRYB_18__39_), .CI(u5_mult_82_SUMB_18__40_), .CO(
        u5_mult_82_CARRYB_19__39_), .S(u5_mult_82_SUMB_19__39_) );
  FA_X1 u5_mult_82_S2_19_36 ( .A(u5_mult_82_CARRYB_18__36_), .B(
        u5_mult_82_ab_19__36_), .CI(u5_mult_82_SUMB_18__37_), .CO(
        u5_mult_82_CARRYB_19__36_), .S(u5_mult_82_SUMB_19__36_) );
  FA_X1 u5_mult_82_S2_19_34 ( .A(u5_mult_82_CARRYB_18__34_), .B(
        u5_mult_82_ab_19__34_), .CI(u5_mult_82_SUMB_18__35_), .CO(
        u5_mult_82_CARRYB_19__34_), .S(u5_mult_82_SUMB_19__34_) );
  FA_X1 u5_mult_82_S2_19_32 ( .A(u5_mult_82_CARRYB_18__32_), .B(
        u5_mult_82_ab_19__32_), .CI(u5_mult_82_SUMB_18__33_), .CO(
        u5_mult_82_CARRYB_19__32_), .S(u5_mult_82_SUMB_19__32_) );
  FA_X1 u5_mult_82_S2_19_31 ( .A(u5_mult_82_ab_19__31_), .B(
        u5_mult_82_CARRYB_18__31_), .CI(u5_mult_82_SUMB_18__32_), .CO(
        u5_mult_82_CARRYB_19__31_), .S(u5_mult_82_SUMB_19__31_) );
  FA_X1 u5_mult_82_S2_19_30 ( .A(u5_mult_82_CARRYB_18__30_), .B(
        u5_mult_82_ab_19__30_), .CI(u5_mult_82_SUMB_18__31_), .CO(
        u5_mult_82_CARRYB_19__30_), .S(u5_mult_82_SUMB_19__30_) );
  FA_X1 u5_mult_82_S2_19_24 ( .A(u5_mult_82_ab_19__24_), .B(
        u5_mult_82_CARRYB_18__24_), .CI(u5_mult_82_SUMB_18__25_), .CO(
        u5_mult_82_CARRYB_19__24_), .S(u5_mult_82_SUMB_19__24_) );
  FA_X1 u5_mult_82_S2_19_19 ( .A(u5_mult_82_ab_19__19_), .B(
        u5_mult_82_CARRYB_18__19_), .CI(u5_mult_82_SUMB_18__20_), .CO(
        u5_mult_82_CARRYB_19__19_), .S(u5_mult_82_SUMB_19__19_) );
  FA_X1 u5_mult_82_S2_19_18 ( .A(u5_mult_82_ab_19__18_), .B(
        u5_mult_82_CARRYB_18__18_), .CI(u5_mult_82_SUMB_18__19_), .CO(
        u5_mult_82_CARRYB_19__18_), .S(u5_mult_82_SUMB_19__18_) );
  FA_X1 u5_mult_82_S2_19_17 ( .A(u5_mult_82_CARRYB_18__17_), .B(
        u5_mult_82_ab_19__17_), .CI(u5_mult_82_SUMB_18__18_), .CO(
        u5_mult_82_CARRYB_19__17_), .S(u5_mult_82_SUMB_19__17_) );
  FA_X1 u5_mult_82_S2_19_16 ( .A(u5_mult_82_ab_19__16_), .B(
        u5_mult_82_CARRYB_18__16_), .CI(u5_mult_82_SUMB_18__17_), .CO(
        u5_mult_82_CARRYB_19__16_), .S(u5_mult_82_SUMB_19__16_) );
  FA_X1 u5_mult_82_S2_19_15 ( .A(u5_mult_82_ab_19__15_), .B(
        u5_mult_82_CARRYB_18__15_), .CI(u5_mult_82_SUMB_18__16_), .CO(
        u5_mult_82_CARRYB_19__15_), .S(u5_mult_82_SUMB_19__15_) );
  FA_X1 u5_mult_82_S2_19_13 ( .A(u5_mult_82_ab_19__13_), .B(
        u5_mult_82_CARRYB_18__13_), .CI(u5_mult_82_SUMB_18__14_), .CO(
        u5_mult_82_CARRYB_19__13_), .S(u5_mult_82_SUMB_19__13_) );
  FA_X1 u5_mult_82_S2_19_10 ( .A(u5_mult_82_CARRYB_18__10_), .B(
        u5_mult_82_ab_19__10_), .CI(u5_mult_82_SUMB_18__11_), .CO(
        u5_mult_82_CARRYB_19__10_), .S(u5_mult_82_SUMB_19__10_) );
  FA_X1 u5_mult_82_S2_19_9 ( .A(u5_mult_82_ab_19__9_), .B(
        u5_mult_82_CARRYB_18__9_), .CI(u5_mult_82_SUMB_18__10_), .CO(
        u5_mult_82_CARRYB_19__9_), .S(u5_mult_82_SUMB_19__9_) );
  FA_X1 u5_mult_82_S2_19_8 ( .A(u5_mult_82_ab_19__8_), .B(
        u5_mult_82_CARRYB_18__8_), .CI(u5_mult_82_SUMB_18__9_), .CO(
        u5_mult_82_CARRYB_19__8_), .S(u5_mult_82_SUMB_19__8_) );
  FA_X1 u5_mult_82_S2_19_7 ( .A(u5_mult_82_ab_19__7_), .B(
        u5_mult_82_CARRYB_18__7_), .CI(u5_mult_82_SUMB_18__8_), .CO(
        u5_mult_82_CARRYB_19__7_), .S(u5_mult_82_SUMB_19__7_) );
  FA_X1 u5_mult_82_S2_19_6 ( .A(u5_mult_82_ab_19__6_), .B(
        u5_mult_82_CARRYB_18__6_), .CI(u5_mult_82_SUMB_18__7_), .CO(
        u5_mult_82_CARRYB_19__6_), .S(u5_mult_82_SUMB_19__6_) );
  FA_X1 u5_mult_82_S2_19_3 ( .A(u5_mult_82_ab_19__3_), .B(
        u5_mult_82_CARRYB_18__3_), .CI(u5_mult_82_SUMB_18__4_), .CO(
        u5_mult_82_CARRYB_19__3_), .S(u5_mult_82_SUMB_19__3_) );
  FA_X1 u5_mult_82_S2_19_2 ( .A(u5_mult_82_ab_19__2_), .B(
        u5_mult_82_CARRYB_18__2_), .CI(u5_mult_82_SUMB_18__3_), .CO(
        u5_mult_82_CARRYB_19__2_), .S(u5_mult_82_SUMB_19__2_) );
  FA_X1 u5_mult_82_S2_19_1 ( .A(u5_mult_82_ab_19__1_), .B(
        u5_mult_82_CARRYB_18__1_), .CI(u5_mult_82_SUMB_18__2_), .CO(
        u5_mult_82_CARRYB_19__1_), .S(u5_mult_82_SUMB_19__1_) );
  FA_X1 u5_mult_82_S1_19_0 ( .A(u5_mult_82_ab_19__0_), .B(
        u5_mult_82_CARRYB_18__0_), .CI(u5_mult_82_SUMB_18__1_), .CO(
        u5_mult_82_CARRYB_19__0_), .S(u5_N19) );
  FA_X1 u5_mult_82_S3_20_51 ( .A(u5_mult_82_ab_20__51_), .B(
        u5_mult_82_CARRYB_19__51_), .CI(u5_mult_82_ab_19__52_), .CO(
        u5_mult_82_CARRYB_20__51_), .S(u5_mult_82_SUMB_20__51_) );
  FA_X1 u5_mult_82_S2_20_50 ( .A(u5_mult_82_ab_20__50_), .B(
        u5_mult_82_CARRYB_19__50_), .CI(u5_mult_82_SUMB_19__51_), .CO(
        u5_mult_82_CARRYB_20__50_), .S(u5_mult_82_SUMB_20__50_) );
  FA_X1 u5_mult_82_S2_20_48 ( .A(u5_mult_82_ab_20__48_), .B(
        u5_mult_82_CARRYB_19__48_), .CI(u5_mult_82_SUMB_19__49_), .CO(
        u5_mult_82_CARRYB_20__48_), .S(u5_mult_82_SUMB_20__48_) );
  FA_X1 u5_mult_82_S2_20_47 ( .A(u5_mult_82_ab_20__47_), .B(
        u5_mult_82_CARRYB_19__47_), .CI(u5_mult_82_SUMB_19__48_), .CO(
        u5_mult_82_CARRYB_20__47_), .S(u5_mult_82_SUMB_20__47_) );
  FA_X1 u5_mult_82_S2_20_46 ( .A(u5_mult_82_ab_20__46_), .B(
        u5_mult_82_CARRYB_19__46_), .CI(u5_mult_82_SUMB_19__47_), .CO(
        u5_mult_82_CARRYB_20__46_), .S(u5_mult_82_SUMB_20__46_) );
  FA_X1 u5_mult_82_S2_20_45 ( .A(u5_mult_82_CARRYB_19__45_), .B(
        u5_mult_82_ab_20__45_), .CI(u5_mult_82_SUMB_19__46_), .CO(
        u5_mult_82_CARRYB_20__45_), .S(u5_mult_82_SUMB_20__45_) );
  FA_X1 u5_mult_82_S2_20_44 ( .A(u5_mult_82_ab_20__44_), .B(
        u5_mult_82_CARRYB_19__44_), .CI(u5_mult_82_SUMB_19__45_), .CO(
        u5_mult_82_CARRYB_20__44_), .S(u5_mult_82_SUMB_20__44_) );
  FA_X1 u5_mult_82_S2_20_28 ( .A(u5_mult_82_ab_20__28_), .B(
        u5_mult_82_CARRYB_19__28_), .CI(u5_mult_82_SUMB_19__29_), .CO(
        u5_mult_82_CARRYB_20__28_), .S(u5_mult_82_SUMB_20__28_) );
  FA_X1 u5_mult_82_S2_20_18 ( .A(u5_mult_82_CARRYB_19__18_), .B(
        u5_mult_82_ab_20__18_), .CI(u5_mult_82_SUMB_19__19_), .CO(
        u5_mult_82_CARRYB_20__18_), .S(u5_mult_82_SUMB_20__18_) );
  FA_X1 u5_mult_82_S2_20_17 ( .A(u5_mult_82_CARRYB_19__17_), .B(
        u5_mult_82_ab_20__17_), .CI(u5_mult_82_SUMB_19__18_), .CO(
        u5_mult_82_CARRYB_20__17_), .S(u5_mult_82_SUMB_20__17_) );
  FA_X1 u5_mult_82_S2_20_15 ( .A(u5_mult_82_ab_20__15_), .B(
        u5_mult_82_CARRYB_19__15_), .CI(u5_mult_82_SUMB_19__16_), .CO(
        u5_mult_82_CARRYB_20__15_), .S(u5_mult_82_SUMB_20__15_) );
  FA_X1 u5_mult_82_S2_20_13 ( .A(u5_mult_82_ab_20__13_), .B(
        u5_mult_82_CARRYB_19__13_), .CI(u5_mult_82_SUMB_19__14_), .CO(
        u5_mult_82_CARRYB_20__13_), .S(u5_mult_82_SUMB_20__13_) );
  FA_X1 u5_mult_82_S2_20_12 ( .A(u5_mult_82_ab_20__12_), .B(
        u5_mult_82_CARRYB_19__12_), .CI(u5_mult_82_SUMB_19__13_), .CO(
        u5_mult_82_CARRYB_20__12_), .S(u5_mult_82_SUMB_20__12_) );
  FA_X1 u5_mult_82_S2_20_11 ( .A(u5_mult_82_ab_20__11_), .B(
        u5_mult_82_CARRYB_19__11_), .CI(u5_mult_82_SUMB_19__12_), .CO(
        u5_mult_82_CARRYB_20__11_), .S(u5_mult_82_SUMB_20__11_) );
  FA_X1 u5_mult_82_S2_20_10 ( .A(u5_mult_82_ab_20__10_), .B(
        u5_mult_82_CARRYB_19__10_), .CI(u5_mult_82_SUMB_19__11_), .CO(
        u5_mult_82_CARRYB_20__10_), .S(u5_mult_82_SUMB_20__10_) );
  FA_X1 u5_mult_82_S2_20_9 ( .A(u5_mult_82_CARRYB_19__9_), .B(
        u5_mult_82_ab_20__9_), .CI(u5_mult_82_SUMB_19__10_), .CO(
        u5_mult_82_CARRYB_20__9_), .S(u5_mult_82_SUMB_20__9_) );
  FA_X1 u5_mult_82_S2_20_8 ( .A(u5_mult_82_ab_20__8_), .B(
        u5_mult_82_CARRYB_19__8_), .CI(u5_mult_82_SUMB_19__9_), .CO(
        u5_mult_82_CARRYB_20__8_), .S(u5_mult_82_SUMB_20__8_) );
  FA_X1 u5_mult_82_S2_20_7 ( .A(u5_mult_82_CARRYB_19__7_), .B(
        u5_mult_82_ab_20__7_), .CI(u5_mult_82_SUMB_19__8_), .CO(
        u5_mult_82_CARRYB_20__7_), .S(u5_mult_82_SUMB_20__7_) );
  FA_X1 u5_mult_82_S2_20_6 ( .A(u5_mult_82_ab_20__6_), .B(
        u5_mult_82_CARRYB_19__6_), .CI(u5_mult_82_SUMB_19__7_), .CO(
        u5_mult_82_CARRYB_20__6_), .S(u5_mult_82_SUMB_20__6_) );
  FA_X1 u5_mult_82_S2_20_5 ( .A(u5_mult_82_ab_20__5_), .B(
        u5_mult_82_CARRYB_19__5_), .CI(u5_mult_82_SUMB_19__6_), .CO(
        u5_mult_82_CARRYB_20__5_), .S(u5_mult_82_SUMB_20__5_) );
  FA_X1 u5_mult_82_S2_20_2 ( .A(u5_mult_82_ab_20__2_), .B(
        u5_mult_82_CARRYB_19__2_), .CI(u5_mult_82_SUMB_19__3_), .CO(
        u5_mult_82_CARRYB_20__2_), .S(u5_mult_82_SUMB_20__2_) );
  FA_X1 u5_mult_82_S2_20_1 ( .A(u5_mult_82_ab_20__1_), .B(
        u5_mult_82_CARRYB_19__1_), .CI(u5_mult_82_SUMB_19__2_), .CO(
        u5_mult_82_CARRYB_20__1_), .S(u5_mult_82_SUMB_20__1_) );
  FA_X1 u5_mult_82_S1_20_0 ( .A(u5_mult_82_ab_20__0_), .B(
        u5_mult_82_CARRYB_19__0_), .CI(u5_mult_82_SUMB_19__1_), .CO(
        u5_mult_82_CARRYB_20__0_), .S(u5_N20) );
  FA_X1 u5_mult_82_S3_21_51 ( .A(u5_mult_82_ab_21__51_), .B(
        u5_mult_82_CARRYB_20__51_), .CI(u5_mult_82_ab_20__52_), .CO(
        u5_mult_82_CARRYB_21__51_), .S(u5_mult_82_SUMB_21__51_) );
  FA_X1 u5_mult_82_S2_21_50 ( .A(u5_mult_82_ab_21__50_), .B(
        u5_mult_82_CARRYB_20__50_), .CI(u5_mult_82_SUMB_20__51_), .CO(
        u5_mult_82_CARRYB_21__50_), .S(u5_mult_82_SUMB_21__50_) );
  FA_X1 u5_mult_82_S2_21_48 ( .A(u5_mult_82_ab_21__48_), .B(
        u5_mult_82_SUMB_20__49_), .CI(u5_mult_82_CARRYB_20__48_), .CO(
        u5_mult_82_CARRYB_21__48_), .S(u5_mult_82_SUMB_21__48_) );
  FA_X1 u5_mult_82_S2_21_47 ( .A(u5_mult_82_ab_21__47_), .B(
        u5_mult_82_CARRYB_20__47_), .CI(u5_mult_82_SUMB_20__48_), .CO(
        u5_mult_82_CARRYB_21__47_), .S(u5_mult_82_SUMB_21__47_) );
  FA_X1 u5_mult_82_S2_21_45 ( .A(u5_mult_82_ab_21__45_), .B(
        u5_mult_82_CARRYB_20__45_), .CI(u5_mult_82_SUMB_20__46_), .CO(
        u5_mult_82_CARRYB_21__45_), .S(u5_mult_82_SUMB_21__45_) );
  FA_X1 u5_mult_82_S2_21_44 ( .A(u5_mult_82_CARRYB_20__44_), .B(
        u5_mult_82_ab_21__44_), .CI(u5_mult_82_SUMB_20__45_), .CO(
        u5_mult_82_CARRYB_21__44_), .S(u5_mult_82_SUMB_21__44_) );
  FA_X1 u5_mult_82_S2_21_43 ( .A(u5_mult_82_ab_21__43_), .B(
        u5_mult_82_CARRYB_20__43_), .CI(u5_mult_82_SUMB_20__44_), .CO(
        u5_mult_82_CARRYB_21__43_), .S(u5_mult_82_SUMB_21__43_) );
  FA_X1 u5_mult_82_S2_21_32 ( .A(u5_mult_82_ab_21__32_), .B(
        u5_mult_82_CARRYB_20__32_), .CI(u5_mult_82_SUMB_20__33_), .CO(
        u5_mult_82_CARRYB_21__32_), .S(u5_mult_82_SUMB_21__32_) );
  FA_X1 u5_mult_82_S2_21_31 ( .A(u5_mult_82_ab_21__31_), .B(
        u5_mult_82_CARRYB_20__31_), .CI(u5_mult_82_SUMB_20__32_), .CO(
        u5_mult_82_CARRYB_21__31_), .S(u5_mult_82_SUMB_21__31_) );
  FA_X1 u5_mult_82_S2_21_27 ( .A(u5_mult_82_ab_21__27_), .B(
        u5_mult_82_CARRYB_20__27_), .CI(u5_mult_82_SUMB_20__28_), .CO(
        u5_mult_82_CARRYB_21__27_), .S(u5_mult_82_SUMB_21__27_) );
  FA_X1 u5_mult_82_S2_21_17 ( .A(u5_mult_82_ab_21__17_), .B(
        u5_mult_82_CARRYB_20__17_), .CI(u5_mult_82_SUMB_20__18_), .CO(
        u5_mult_82_CARRYB_21__17_), .S(u5_mult_82_SUMB_21__17_) );
  FA_X1 u5_mult_82_S2_21_12 ( .A(u5_mult_82_ab_21__12_), .B(
        u5_mult_82_CARRYB_20__12_), .CI(u5_mult_82_SUMB_20__13_), .CO(
        u5_mult_82_CARRYB_21__12_), .S(u5_mult_82_SUMB_21__12_) );
  FA_X1 u5_mult_82_S2_21_8 ( .A(u5_mult_82_CARRYB_20__8_), .B(
        u5_mult_82_ab_21__8_), .CI(u5_mult_82_SUMB_20__9_), .CO(
        u5_mult_82_CARRYB_21__8_), .S(u5_mult_82_SUMB_21__8_) );
  FA_X1 u5_mult_82_S2_21_6 ( .A(u5_mult_82_ab_21__6_), .B(
        u5_mult_82_CARRYB_20__6_), .CI(u5_mult_82_SUMB_20__7_), .CO(
        u5_mult_82_CARRYB_21__6_), .S(u5_mult_82_SUMB_21__6_) );
  FA_X1 u5_mult_82_S2_21_4 ( .A(u5_mult_82_ab_21__4_), .B(
        u5_mult_82_CARRYB_20__4_), .CI(u5_mult_82_SUMB_20__5_), .CO(
        u5_mult_82_CARRYB_21__4_), .S(u5_mult_82_SUMB_21__4_) );
  FA_X1 u5_mult_82_S2_21_3 ( .A(u5_mult_82_ab_21__3_), .B(
        u5_mult_82_CARRYB_20__3_), .CI(u5_mult_82_SUMB_20__4_), .CO(
        u5_mult_82_CARRYB_21__3_), .S(u5_mult_82_SUMB_21__3_) );
  FA_X1 u5_mult_82_S2_21_2 ( .A(u5_mult_82_ab_21__2_), .B(
        u5_mult_82_CARRYB_20__2_), .CI(u5_mult_82_SUMB_20__3_), .CO(
        u5_mult_82_CARRYB_21__2_), .S(u5_mult_82_SUMB_21__2_) );
  FA_X1 u5_mult_82_S2_21_1 ( .A(u5_mult_82_ab_21__1_), .B(
        u5_mult_82_CARRYB_20__1_), .CI(u5_mult_82_SUMB_20__2_), .CO(
        u5_mult_82_CARRYB_21__1_), .S(u5_mult_82_SUMB_21__1_) );
  FA_X1 u5_mult_82_S1_21_0 ( .A(u5_mult_82_ab_21__0_), .B(
        u5_mult_82_CARRYB_20__0_), .CI(u5_mult_82_SUMB_20__1_), .CO(
        u5_mult_82_CARRYB_21__0_), .S(u5_N21) );
  FA_X1 u5_mult_82_S3_22_51 ( .A(u5_mult_82_ab_22__51_), .B(
        u5_mult_82_CARRYB_21__51_), .CI(u5_mult_82_ab_21__52_), .CO(
        u5_mult_82_CARRYB_22__51_), .S(u5_mult_82_SUMB_22__51_) );
  FA_X1 u5_mult_82_S2_22_50 ( .A(u5_mult_82_ab_22__50_), .B(
        u5_mult_82_CARRYB_21__50_), .CI(u5_mult_82_SUMB_21__51_), .CO(
        u5_mult_82_CARRYB_22__50_), .S(u5_mult_82_SUMB_22__50_) );
  FA_X1 u5_mult_82_S2_22_49 ( .A(u5_mult_82_ab_22__49_), .B(
        u5_mult_82_CARRYB_21__49_), .CI(u5_mult_82_SUMB_21__50_), .CO(
        u5_mult_82_CARRYB_22__49_), .S(u5_mult_82_SUMB_22__49_) );
  FA_X1 u5_mult_82_S2_22_43 ( .A(u5_mult_82_ab_22__43_), .B(
        u5_mult_82_CARRYB_21__43_), .CI(u5_mult_82_SUMB_21__44_), .CO(
        u5_mult_82_CARRYB_22__43_), .S(u5_mult_82_SUMB_22__43_) );
  FA_X1 u5_mult_82_S2_22_42 ( .A(u5_mult_82_ab_22__42_), .B(
        u5_mult_82_CARRYB_21__42_), .CI(u5_mult_82_SUMB_21__43_), .CO(
        u5_mult_82_CARRYB_22__42_), .S(u5_mult_82_SUMB_22__42_) );
  FA_X1 u5_mult_82_S2_22_41 ( .A(u5_mult_82_ab_22__41_), .B(
        u5_mult_82_CARRYB_21__41_), .CI(u5_mult_82_SUMB_21__42_), .CO(
        u5_mult_82_CARRYB_22__41_), .S(u5_mult_82_SUMB_22__41_) );
  FA_X1 u5_mult_82_S2_22_36 ( .A(u5_mult_82_ab_22__36_), .B(
        u5_mult_82_CARRYB_21__36_), .CI(u5_mult_82_SUMB_21__37_), .CO(
        u5_mult_82_CARRYB_22__36_), .S(u5_mult_82_SUMB_22__36_) );
  FA_X1 u5_mult_82_S2_22_33 ( .A(u5_mult_82_CARRYB_21__33_), .B(
        u5_mult_82_ab_22__33_), .CI(u5_mult_82_SUMB_21__34_), .CO(
        u5_mult_82_CARRYB_22__33_), .S(u5_mult_82_SUMB_22__33_) );
  FA_X1 u5_mult_82_S2_22_28 ( .A(u5_mult_82_ab_22__28_), .B(
        u5_mult_82_CARRYB_21__28_), .CI(u5_mult_82_SUMB_21__29_), .CO(
        u5_mult_82_CARRYB_22__28_), .S(u5_mult_82_SUMB_22__28_) );
  FA_X1 u5_mult_82_S2_22_21 ( .A(u5_mult_82_ab_22__21_), .B(
        u5_mult_82_CARRYB_21__21_), .CI(u5_mult_82_SUMB_21__22_), .CO(
        u5_mult_82_CARRYB_22__21_), .S(u5_mult_82_SUMB_22__21_) );
  FA_X1 u5_mult_82_S2_22_20 ( .A(u5_mult_82_ab_22__20_), .B(
        u5_mult_82_CARRYB_21__20_), .CI(u5_mult_82_SUMB_21__21_), .CO(
        u5_mult_82_CARRYB_22__20_), .S(u5_mult_82_SUMB_22__20_) );
  FA_X1 u5_mult_82_S2_22_19 ( .A(u5_mult_82_ab_22__19_), .B(
        u5_mult_82_CARRYB_21__19_), .CI(u5_mult_82_SUMB_21__20_), .CO(
        u5_mult_82_CARRYB_22__19_), .S(u5_mult_82_SUMB_22__19_) );
  FA_X1 u5_mult_82_S2_22_17 ( .A(u5_mult_82_ab_22__17_), .B(
        u5_mult_82_SUMB_21__18_), .CI(u5_mult_82_CARRYB_21__17_), .CO(
        u5_mult_82_CARRYB_22__17_), .S(u5_mult_82_SUMB_22__17_) );
  FA_X1 u5_mult_82_S2_22_15 ( .A(u5_mult_82_CARRYB_21__15_), .B(
        u5_mult_82_ab_22__15_), .CI(u5_mult_82_SUMB_21__16_), .CO(
        u5_mult_82_CARRYB_22__15_), .S(u5_mult_82_SUMB_22__15_) );
  FA_X1 u5_mult_82_S2_22_14 ( .A(u5_mult_82_ab_22__14_), .B(
        u5_mult_82_CARRYB_21__14_), .CI(u5_mult_82_SUMB_21__15_), .CO(
        u5_mult_82_CARRYB_22__14_), .S(u5_mult_82_SUMB_22__14_) );
  FA_X1 u5_mult_82_S2_22_11 ( .A(u5_mult_82_ab_22__11_), .B(
        u5_mult_82_CARRYB_21__11_), .CI(u5_mult_82_SUMB_21__12_), .CO(
        u5_mult_82_CARRYB_22__11_), .S(u5_mult_82_SUMB_22__11_) );
  FA_X1 u5_mult_82_S2_22_7 ( .A(u5_mult_82_ab_22__7_), .B(
        u5_mult_82_CARRYB_21__7_), .CI(u5_mult_82_SUMB_21__8_), .CO(
        u5_mult_82_CARRYB_22__7_), .S(u5_mult_82_SUMB_22__7_) );
  FA_X1 u5_mult_82_S2_22_6 ( .A(u5_mult_82_ab_22__6_), .B(
        u5_mult_82_CARRYB_21__6_), .CI(u5_mult_82_SUMB_21__7_), .CO(
        u5_mult_82_CARRYB_22__6_), .S(u5_mult_82_SUMB_22__6_) );
  FA_X1 u5_mult_82_S2_22_4 ( .A(u5_mult_82_ab_22__4_), .B(
        u5_mult_82_CARRYB_21__4_), .CI(u5_mult_82_SUMB_21__5_), .CO(
        u5_mult_82_CARRYB_22__4_), .S(u5_mult_82_SUMB_22__4_) );
  FA_X1 u5_mult_82_S2_22_3 ( .A(u5_mult_82_ab_22__3_), .B(
        u5_mult_82_CARRYB_21__3_), .CI(u5_mult_82_SUMB_21__4_), .CO(
        u5_mult_82_CARRYB_22__3_), .S(u5_mult_82_SUMB_22__3_) );
  FA_X1 u5_mult_82_S2_22_2 ( .A(u5_mult_82_ab_22__2_), .B(
        u5_mult_82_CARRYB_21__2_), .CI(u5_mult_82_SUMB_21__3_), .CO(
        u5_mult_82_CARRYB_22__2_), .S(u5_mult_82_SUMB_22__2_) );
  FA_X1 u5_mult_82_S2_22_1 ( .A(u5_mult_82_ab_22__1_), .B(
        u5_mult_82_CARRYB_21__1_), .CI(u5_mult_82_SUMB_21__2_), .CO(
        u5_mult_82_CARRYB_22__1_), .S(u5_mult_82_SUMB_22__1_) );
  FA_X1 u5_mult_82_S1_22_0 ( .A(u5_mult_82_ab_22__0_), .B(
        u5_mult_82_CARRYB_21__0_), .CI(u5_mult_82_SUMB_21__1_), .CO(
        u5_mult_82_CARRYB_22__0_), .S(u5_N22) );
  FA_X1 u5_mult_82_S3_23_51 ( .A(u5_mult_82_ab_23__51_), .B(
        u5_mult_82_CARRYB_22__51_), .CI(u5_mult_82_ab_22__52_), .CO(
        u5_mult_82_CARRYB_23__51_), .S(u5_mult_82_SUMB_23__51_) );
  FA_X1 u5_mult_82_S2_23_49 ( .A(u5_mult_82_ab_23__49_), .B(
        u5_mult_82_CARRYB_22__49_), .CI(u5_mult_82_SUMB_22__50_), .CO(
        u5_mult_82_CARRYB_23__49_), .S(u5_mult_82_SUMB_23__49_) );
  FA_X1 u5_mult_82_S2_23_45 ( .A(u5_mult_82_ab_23__45_), .B(
        u5_mult_82_CARRYB_22__45_), .CI(u5_mult_82_SUMB_22__46_), .CO(
        u5_mult_82_CARRYB_23__45_), .S(u5_mult_82_SUMB_23__45_) );
  FA_X1 u5_mult_82_S2_23_42 ( .A(u5_mult_82_ab_23__42_), .B(
        u5_mult_82_CARRYB_22__42_), .CI(u5_mult_82_SUMB_22__43_), .CO(
        u5_mult_82_CARRYB_23__42_), .S(u5_mult_82_SUMB_23__42_) );
  FA_X1 u5_mult_82_S2_23_33 ( .A(u5_mult_82_ab_23__33_), .B(
        u5_mult_82_CARRYB_22__33_), .CI(u5_mult_82_SUMB_22__34_), .CO(
        u5_mult_82_CARRYB_23__33_), .S(u5_mult_82_SUMB_23__33_) );
  FA_X1 u5_mult_82_S2_23_27 ( .A(u5_mult_82_ab_23__27_), .B(
        u5_mult_82_CARRYB_22__27_), .CI(u5_mult_82_SUMB_22__28_), .CO(
        u5_mult_82_CARRYB_23__27_), .S(u5_mult_82_SUMB_23__27_) );
  FA_X1 u5_mult_82_S2_23_20 ( .A(u5_mult_82_ab_23__20_), .B(
        u5_mult_82_CARRYB_22__20_), .CI(u5_mult_82_SUMB_22__21_), .CO(
        u5_mult_82_CARRYB_23__20_), .S(u5_mult_82_SUMB_23__20_) );
  FA_X1 u5_mult_82_S2_23_16 ( .A(u5_mult_82_CARRYB_22__16_), .B(
        u5_mult_82_ab_23__16_), .CI(u5_mult_82_SUMB_22__17_), .CO(
        u5_mult_82_CARRYB_23__16_), .S(u5_mult_82_SUMB_23__16_) );
  FA_X1 u5_mult_82_S2_23_15 ( .A(u5_mult_82_ab_23__15_), .B(
        u5_mult_82_CARRYB_22__15_), .CI(u5_mult_82_SUMB_22__16_), .CO(
        u5_mult_82_CARRYB_23__15_), .S(u5_mult_82_SUMB_23__15_) );
  FA_X1 u5_mult_82_S2_23_14 ( .A(u5_mult_82_ab_23__14_), .B(
        u5_mult_82_CARRYB_22__14_), .CI(u5_mult_82_SUMB_22__15_), .CO(
        u5_mult_82_CARRYB_23__14_), .S(u5_mult_82_SUMB_23__14_) );
  FA_X1 u5_mult_82_S2_23_13 ( .A(u5_mult_82_ab_23__13_), .B(
        u5_mult_82_CARRYB_22__13_), .CI(u5_mult_82_SUMB_22__14_), .CO(
        u5_mult_82_CARRYB_23__13_), .S(u5_mult_82_SUMB_23__13_) );
  FA_X1 u5_mult_82_S2_23_12 ( .A(u5_mult_82_ab_23__12_), .B(
        u5_mult_82_CARRYB_22__12_), .CI(u5_mult_82_SUMB_22__13_), .CO(
        u5_mult_82_CARRYB_23__12_), .S(u5_mult_82_SUMB_23__12_) );
  FA_X1 u5_mult_82_S2_23_10 ( .A(u5_mult_82_ab_23__10_), .B(
        u5_mult_82_CARRYB_22__10_), .CI(u5_mult_82_SUMB_22__11_), .CO(
        u5_mult_82_CARRYB_23__10_), .S(u5_mult_82_SUMB_23__10_) );
  FA_X1 u5_mult_82_S2_23_6 ( .A(u5_mult_82_CARRYB_22__6_), .B(
        u5_mult_82_ab_23__6_), .CI(u5_mult_82_SUMB_22__7_), .CO(
        u5_mult_82_CARRYB_23__6_), .S(u5_mult_82_SUMB_23__6_) );
  FA_X1 u5_mult_82_S2_23_5 ( .A(u5_mult_82_ab_23__5_), .B(
        u5_mult_82_CARRYB_22__5_), .CI(u5_mult_82_SUMB_22__6_), .CO(
        u5_mult_82_CARRYB_23__5_), .S(u5_mult_82_SUMB_23__5_) );
  FA_X1 u5_mult_82_S2_23_4 ( .A(u5_mult_82_ab_23__4_), .B(
        u5_mult_82_CARRYB_22__4_), .CI(u5_mult_82_SUMB_22__5_), .CO(
        u5_mult_82_CARRYB_23__4_), .S(u5_mult_82_SUMB_23__4_) );
  FA_X1 u5_mult_82_S2_23_3 ( .A(u5_mult_82_ab_23__3_), .B(
        u5_mult_82_CARRYB_22__3_), .CI(u5_mult_82_SUMB_22__4_), .CO(
        u5_mult_82_CARRYB_23__3_), .S(u5_mult_82_SUMB_23__3_) );
  FA_X1 u5_mult_82_S2_23_2 ( .A(u5_mult_82_ab_23__2_), .B(
        u5_mult_82_CARRYB_22__2_), .CI(u5_mult_82_SUMB_22__3_), .CO(
        u5_mult_82_CARRYB_23__2_), .S(u5_mult_82_SUMB_23__2_) );
  FA_X1 u5_mult_82_S2_23_1 ( .A(u5_mult_82_ab_23__1_), .B(
        u5_mult_82_CARRYB_22__1_), .CI(u5_mult_82_SUMB_22__2_), .CO(
        u5_mult_82_CARRYB_23__1_), .S(u5_mult_82_SUMB_23__1_) );
  FA_X1 u5_mult_82_S1_23_0 ( .A(u5_mult_82_ab_23__0_), .B(
        u5_mult_82_CARRYB_22__0_), .CI(u5_mult_82_SUMB_22__1_), .CO(
        u5_mult_82_CARRYB_23__0_), .S(u5_N23) );
  FA_X1 u5_mult_82_S3_24_51 ( .A(u5_mult_82_ab_24__51_), .B(
        u5_mult_82_CARRYB_23__51_), .CI(u5_mult_82_ab_23__52_), .CO(
        u5_mult_82_CARRYB_24__51_), .S(u5_mult_82_SUMB_24__51_) );
  FA_X1 u5_mult_82_S2_24_50 ( .A(u5_mult_82_CARRYB_23__50_), .B(
        u5_mult_82_ab_24__50_), .CI(u5_mult_82_SUMB_23__51_), .CO(
        u5_mult_82_CARRYB_24__50_), .S(u5_mult_82_SUMB_24__50_) );
  FA_X1 u5_mult_82_S2_24_49 ( .A(u5_mult_82_ab_24__49_), .B(
        u5_mult_82_CARRYB_23__49_), .CI(u5_mult_82_SUMB_23__50_), .CO(
        u5_mult_82_CARRYB_24__49_), .S(u5_mult_82_SUMB_24__49_) );
  FA_X1 u5_mult_82_S2_24_44 ( .A(u5_mult_82_ab_24__44_), .B(
        u5_mult_82_CARRYB_23__44_), .CI(u5_mult_82_SUMB_23__45_), .CO(
        u5_mult_82_CARRYB_24__44_), .S(u5_mult_82_SUMB_24__44_) );
  FA_X1 u5_mult_82_S2_24_43 ( .A(u5_mult_82_CARRYB_23__43_), .B(
        u5_mult_82_ab_24__43_), .CI(u5_mult_82_SUMB_23__44_), .CO(
        u5_mult_82_CARRYB_24__43_), .S(u5_mult_82_SUMB_24__43_) );
  FA_X1 u5_mult_82_S2_24_35 ( .A(u5_mult_82_SUMB_23__36_), .B(
        u5_mult_82_ab_24__35_), .CI(u5_mult_82_CARRYB_23__35_), .CO(
        u5_mult_82_CARRYB_24__35_), .S(u5_mult_82_SUMB_24__35_) );
  FA_X1 u5_mult_82_S2_24_30 ( .A(u5_mult_82_ab_24__30_), .B(
        u5_mult_82_CARRYB_23__30_), .CI(u5_mult_82_SUMB_23__31_), .CO(
        u5_mult_82_CARRYB_24__30_), .S(u5_mult_82_SUMB_24__30_) );
  FA_X1 u5_mult_82_S2_24_19 ( .A(u5_mult_82_ab_24__19_), .B(
        u5_mult_82_CARRYB_23__19_), .CI(u5_mult_82_SUMB_23__20_), .CO(
        u5_mult_82_CARRYB_24__19_), .S(u5_mult_82_SUMB_24__19_) );
  FA_X1 u5_mult_82_S2_24_15 ( .A(u5_mult_82_CARRYB_23__15_), .B(
        u5_mult_82_ab_24__15_), .CI(u5_mult_82_SUMB_23__16_), .CO(
        u5_mult_82_CARRYB_24__15_), .S(u5_mult_82_SUMB_24__15_) );
  FA_X1 u5_mult_82_S2_24_14 ( .A(u5_mult_82_CARRYB_23__14_), .B(
        u5_mult_82_ab_24__14_), .CI(u5_mult_82_SUMB_23__15_), .CO(
        u5_mult_82_CARRYB_24__14_), .S(u5_mult_82_SUMB_24__14_) );
  FA_X1 u5_mult_82_S2_24_11 ( .A(u5_mult_82_ab_24__11_), .B(
        u5_mult_82_CARRYB_23__11_), .CI(u5_mult_82_SUMB_23__12_), .CO(
        u5_mult_82_CARRYB_24__11_), .S(u5_mult_82_SUMB_24__11_) );
  FA_X1 u5_mult_82_S2_24_7 ( .A(u5_mult_82_CARRYB_23__7_), .B(
        u5_mult_82_ab_24__7_), .CI(u5_mult_82_SUMB_23__8_), .CO(
        u5_mult_82_CARRYB_24__7_), .S(u5_mult_82_SUMB_24__7_) );
  FA_X1 u5_mult_82_S2_24_5 ( .A(u5_mult_82_ab_24__5_), .B(
        u5_mult_82_CARRYB_23__5_), .CI(u5_mult_82_SUMB_23__6_), .CO(
        u5_mult_82_CARRYB_24__5_), .S(u5_mult_82_SUMB_24__5_) );
  FA_X1 u5_mult_82_S2_24_3 ( .A(u5_mult_82_ab_24__3_), .B(
        u5_mult_82_CARRYB_23__3_), .CI(u5_mult_82_SUMB_23__4_), .CO(
        u5_mult_82_CARRYB_24__3_), .S(u5_mult_82_SUMB_24__3_) );
  FA_X1 u5_mult_82_S2_24_2 ( .A(u5_mult_82_ab_24__2_), .B(
        u5_mult_82_CARRYB_23__2_), .CI(u5_mult_82_SUMB_23__3_), .CO(
        u5_mult_82_CARRYB_24__2_), .S(u5_mult_82_SUMB_24__2_) );
  FA_X1 u5_mult_82_S1_24_0 ( .A(u5_mult_82_ab_24__0_), .B(
        u5_mult_82_CARRYB_23__0_), .CI(u5_mult_82_SUMB_23__1_), .CO(
        u5_mult_82_CARRYB_24__0_), .S(u5_N24) );
  FA_X1 u5_mult_82_S3_25_51 ( .A(u5_mult_82_ab_25__51_), .B(
        u5_mult_82_CARRYB_24__51_), .CI(u5_mult_82_ab_24__52_), .CO(
        u5_mult_82_CARRYB_25__51_), .S(u5_mult_82_SUMB_25__51_) );
  FA_X1 u5_mult_82_S2_25_50 ( .A(u5_mult_82_ab_25__50_), .B(
        u5_mult_82_CARRYB_24__50_), .CI(u5_mult_82_SUMB_24__51_), .CO(
        u5_mult_82_CARRYB_25__50_), .S(u5_mult_82_SUMB_25__50_) );
  FA_X1 u5_mult_82_S2_25_49 ( .A(u5_mult_82_ab_25__49_), .B(
        u5_mult_82_CARRYB_24__49_), .CI(u5_mult_82_SUMB_24__50_), .CO(
        u5_mult_82_CARRYB_25__49_), .S(u5_mult_82_SUMB_25__49_) );
  FA_X1 u5_mult_82_S2_25_42 ( .A(u5_mult_82_ab_25__42_), .B(
        u5_mult_82_CARRYB_24__42_), .CI(u5_mult_82_SUMB_24__43_), .CO(
        u5_mult_82_CARRYB_25__42_), .S(u5_mult_82_SUMB_25__42_) );
  FA_X1 u5_mult_82_S2_25_38 ( .A(u5_mult_82_ab_25__38_), .B(
        u5_mult_82_CARRYB_24__38_), .CI(u5_mult_82_SUMB_24__39_), .CO(
        u5_mult_82_CARRYB_25__38_), .S(u5_mult_82_SUMB_25__38_) );
  FA_X1 u5_mult_82_S2_25_35 ( .A(u5_mult_82_CARRYB_24__35_), .B(
        u5_mult_82_ab_25__35_), .CI(u5_mult_82_SUMB_24__36_), .CO(
        u5_mult_82_CARRYB_25__35_), .S(u5_mult_82_SUMB_25__35_) );
  FA_X1 u5_mult_82_S2_25_31 ( .A(u5_mult_82_ab_25__31_), .B(
        u5_mult_82_CARRYB_24__31_), .CI(u5_mult_82_SUMB_24__32_), .CO(
        u5_mult_82_CARRYB_25__31_), .S(u5_mult_82_SUMB_25__31_) );
  FA_X1 u5_mult_82_S2_25_30 ( .A(u5_mult_82_ab_25__30_), .B(
        u5_mult_82_CARRYB_24__30_), .CI(u5_mult_82_SUMB_24__31_), .CO(
        u5_mult_82_CARRYB_25__30_), .S(u5_mult_82_SUMB_25__30_) );
  FA_X1 u5_mult_82_S2_25_27 ( .A(u5_mult_82_ab_25__27_), .B(
        u5_mult_82_CARRYB_24__27_), .CI(u5_mult_82_SUMB_24__28_), .CO(
        u5_mult_82_CARRYB_25__27_), .S(u5_mult_82_SUMB_25__27_) );
  FA_X1 u5_mult_82_S2_25_23 ( .A(u5_mult_82_ab_25__23_), .B(
        u5_mult_82_CARRYB_24__23_), .CI(u5_mult_82_SUMB_24__24_), .CO(
        u5_mult_82_CARRYB_25__23_), .S(u5_mult_82_SUMB_25__23_) );
  FA_X1 u5_mult_82_S2_25_21 ( .A(u5_mult_82_ab_25__21_), .B(
        u5_mult_82_CARRYB_24__21_), .CI(u5_mult_82_SUMB_24__22_), .CO(
        u5_mult_82_CARRYB_25__21_), .S(u5_mult_82_SUMB_25__21_) );
  FA_X1 u5_mult_82_S2_25_10 ( .A(u5_mult_82_ab_25__10_), .B(
        u5_mult_82_CARRYB_24__10_), .CI(u5_mult_82_SUMB_24__11_), .CO(
        u5_mult_82_CARRYB_25__10_), .S(u5_mult_82_SUMB_25__10_) );
  FA_X1 u5_mult_82_S2_25_8 ( .A(u5_mult_82_ab_25__8_), .B(
        u5_mult_82_CARRYB_24__8_), .CI(u5_mult_82_SUMB_24__9_), .CO(
        u5_mult_82_CARRYB_25__8_), .S(u5_mult_82_SUMB_25__8_) );
  FA_X1 u5_mult_82_S2_25_6 ( .A(u5_mult_82_ab_25__6_), .B(
        u5_mult_82_CARRYB_24__6_), .CI(u5_mult_82_SUMB_24__7_), .CO(
        u5_mult_82_CARRYB_25__6_), .S(u5_mult_82_SUMB_25__6_) );
  FA_X1 u5_mult_82_S2_25_2 ( .A(u5_mult_82_ab_25__2_), .B(
        u5_mult_82_CARRYB_24__2_), .CI(u5_mult_82_SUMB_24__3_), .CO(
        u5_mult_82_CARRYB_25__2_), .S(u5_mult_82_SUMB_25__2_) );
  FA_X1 u5_mult_82_S1_25_0 ( .A(u5_mult_82_ab_25__0_), .B(
        u5_mult_82_CARRYB_24__0_), .CI(u5_mult_82_SUMB_24__1_), .CO(
        u5_mult_82_CARRYB_25__0_), .S(u5_N25) );
  FA_X1 u5_mult_82_S3_26_51 ( .A(u5_mult_82_ab_26__51_), .B(
        u5_mult_82_CARRYB_25__51_), .CI(u5_mult_82_ab_25__52_), .CO(
        u5_mult_82_CARRYB_26__51_), .S(u5_mult_82_SUMB_26__51_) );
  FA_X1 u5_mult_82_S2_26_50 ( .A(u5_mult_82_ab_26__50_), .B(
        u5_mult_82_CARRYB_25__50_), .CI(u5_mult_82_SUMB_25__51_), .CO(
        u5_mult_82_CARRYB_26__50_), .S(u5_mult_82_SUMB_26__50_) );
  FA_X1 u5_mult_82_S2_26_49 ( .A(u5_mult_82_ab_26__49_), .B(
        u5_mult_82_CARRYB_25__49_), .CI(u5_mult_82_SUMB_25__50_), .CO(
        u5_mult_82_CARRYB_26__49_), .S(u5_mult_82_SUMB_26__49_) );
  FA_X1 u5_mult_82_S2_26_47 ( .A(u5_mult_82_ab_26__47_), .B(
        u5_mult_82_CARRYB_25__47_), .CI(u5_mult_82_SUMB_25__48_), .CO(
        u5_mult_82_CARRYB_26__47_), .S(u5_mult_82_SUMB_26__47_) );
  FA_X1 u5_mult_82_S2_26_44 ( .A(u5_mult_82_CARRYB_25__44_), .B(
        u5_mult_82_ab_26__44_), .CI(u5_mult_82_SUMB_25__45_), .CO(
        u5_mult_82_CARRYB_26__44_), .S(u5_mult_82_SUMB_26__44_) );
  FA_X1 u5_mult_82_S2_26_41 ( .A(u5_mult_82_ab_26__41_), .B(
        u5_mult_82_CARRYB_25__41_), .CI(u5_mult_82_SUMB_25__42_), .CO(
        u5_mult_82_CARRYB_26__41_), .S(u5_mult_82_SUMB_26__41_) );
  FA_X1 u5_mult_82_S2_26_36 ( .A(u5_mult_82_ab_26__36_), .B(
        u5_mult_82_CARRYB_25__36_), .CI(u5_mult_82_SUMB_25__37_), .CO(
        u5_mult_82_CARRYB_26__36_), .S(u5_mult_82_SUMB_26__36_) );
  FA_X1 u5_mult_82_S2_26_31 ( .A(u5_mult_82_ab_26__31_), .B(
        u5_mult_82_CARRYB_25__31_), .CI(u5_mult_82_SUMB_25__32_), .CO(
        u5_mult_82_CARRYB_26__31_), .S(u5_mult_82_SUMB_26__31_) );
  FA_X1 u5_mult_82_S2_26_24 ( .A(u5_mult_82_ab_26__24_), .B(
        u5_mult_82_CARRYB_25__24_), .CI(u5_mult_82_SUMB_25__25_), .CO(
        u5_mult_82_CARRYB_26__24_), .S(u5_mult_82_SUMB_26__24_) );
  FA_X1 u5_mult_82_S2_26_23 ( .A(u5_mult_82_CARRYB_25__23_), .B(
        u5_mult_82_ab_26__23_), .CI(u5_mult_82_SUMB_25__24_), .CO(
        u5_mult_82_CARRYB_26__23_), .S(u5_mult_82_SUMB_26__23_) );
  FA_X1 u5_mult_82_S2_26_18 ( .A(u5_mult_82_ab_26__18_), .B(
        u5_mult_82_CARRYB_25__18_), .CI(u5_mult_82_SUMB_25__19_), .CO(
        u5_mult_82_CARRYB_26__18_), .S(u5_mult_82_SUMB_26__18_) );
  FA_X1 u5_mult_82_S2_26_11 ( .A(u5_mult_82_ab_26__11_), .B(
        u5_mult_82_CARRYB_25__11_), .CI(u5_mult_82_SUMB_25__12_), .CO(
        u5_mult_82_CARRYB_26__11_), .S(u5_mult_82_SUMB_26__11_) );
  FA_X1 u5_mult_82_S2_26_7 ( .A(u5_mult_82_ab_26__7_), .B(
        u5_mult_82_CARRYB_25__7_), .CI(u5_mult_82_SUMB_25__8_), .CO(
        u5_mult_82_CARRYB_26__7_), .S(u5_mult_82_SUMB_26__7_) );
  FA_X1 u5_mult_82_S2_26_5 ( .A(u5_mult_82_ab_26__5_), .B(
        u5_mult_82_CARRYB_25__5_), .CI(u5_mult_82_SUMB_25__6_), .CO(
        u5_mult_82_CARRYB_26__5_), .S(u5_mult_82_SUMB_26__5_) );
  FA_X1 u5_mult_82_S2_26_3 ( .A(u5_mult_82_ab_26__3_), .B(
        u5_mult_82_CARRYB_25__3_), .CI(u5_mult_82_SUMB_25__4_), .CO(
        u5_mult_82_CARRYB_26__3_), .S(u5_mult_82_SUMB_26__3_) );
  FA_X1 u5_mult_82_S2_26_2 ( .A(u5_mult_82_ab_26__2_), .B(
        u5_mult_82_CARRYB_25__2_), .CI(u5_mult_82_SUMB_25__3_), .CO(
        u5_mult_82_CARRYB_26__2_), .S(u5_mult_82_SUMB_26__2_) );
  FA_X1 u5_mult_82_S1_26_0 ( .A(u5_mult_82_ab_26__0_), .B(
        u5_mult_82_CARRYB_25__0_), .CI(u5_mult_82_SUMB_25__1_), .CO(
        u5_mult_82_CARRYB_26__0_), .S(u5_N26) );
  FA_X1 u5_mult_82_S3_27_51 ( .A(u5_mult_82_ab_27__51_), .B(
        u5_mult_82_CARRYB_26__51_), .CI(u5_mult_82_ab_26__52_), .CO(
        u5_mult_82_CARRYB_27__51_), .S(u5_mult_82_SUMB_27__51_) );
  FA_X1 u5_mult_82_S2_27_50 ( .A(u5_mult_82_ab_27__50_), .B(
        u5_mult_82_CARRYB_26__50_), .CI(u5_mult_82_SUMB_26__51_), .CO(
        u5_mult_82_CARRYB_27__50_), .S(u5_mult_82_SUMB_27__50_) );
  FA_X1 u5_mult_82_S2_27_49 ( .A(u5_mult_82_ab_27__49_), .B(
        u5_mult_82_CARRYB_26__49_), .CI(u5_mult_82_SUMB_26__50_), .CO(
        u5_mult_82_CARRYB_27__49_), .S(u5_mult_82_SUMB_27__49_) );
  FA_X1 u5_mult_82_S2_27_48 ( .A(u5_mult_82_ab_27__48_), .B(
        u5_mult_82_CARRYB_26__48_), .CI(u5_mult_82_SUMB_26__49_), .CO(
        u5_mult_82_CARRYB_27__48_), .S(u5_mult_82_SUMB_27__48_) );
  FA_X1 u5_mult_82_S2_27_47 ( .A(u5_mult_82_ab_27__47_), .B(
        u5_mult_82_CARRYB_26__47_), .CI(u5_mult_82_SUMB_26__48_), .CO(
        u5_mult_82_CARRYB_27__47_), .S(u5_mult_82_SUMB_27__47_) );
  FA_X1 u5_mult_82_S2_27_46 ( .A(u5_mult_82_ab_27__46_), .B(
        u5_mult_82_CARRYB_26__46_), .CI(u5_mult_82_SUMB_26__47_), .CO(
        u5_mult_82_CARRYB_27__46_), .S(u5_mult_82_SUMB_27__46_) );
  FA_X1 u5_mult_82_S2_27_45 ( .A(u5_mult_82_ab_27__45_), .B(
        u5_mult_82_CARRYB_26__45_), .CI(u5_mult_82_SUMB_26__46_), .CO(
        u5_mult_82_CARRYB_27__45_), .S(u5_mult_82_SUMB_27__45_) );
  FA_X1 u5_mult_82_S2_27_44 ( .A(u5_mult_82_ab_27__44_), .B(
        u5_mult_82_CARRYB_26__44_), .CI(u5_mult_82_SUMB_26__45_), .CO(
        u5_mult_82_CARRYB_27__44_), .S(u5_mult_82_SUMB_27__44_) );
  FA_X1 u5_mult_82_S2_27_42 ( .A(u5_mult_82_ab_27__42_), .B(
        u5_mult_82_CARRYB_26__42_), .CI(u5_mult_82_SUMB_26__43_), .CO(
        u5_mult_82_CARRYB_27__42_), .S(u5_mult_82_SUMB_27__42_) );
  FA_X1 u5_mult_82_S2_27_39 ( .A(u5_mult_82_ab_27__39_), .B(
        u5_mult_82_CARRYB_26__39_), .CI(u5_mult_82_SUMB_26__40_), .CO(
        u5_mult_82_CARRYB_27__39_), .S(u5_mult_82_SUMB_27__39_) );
  FA_X1 u5_mult_82_S2_27_37 ( .A(u5_mult_82_ab_27__37_), .B(
        u5_mult_82_CARRYB_26__37_), .CI(u5_mult_82_SUMB_26__38_), .CO(
        u5_mult_82_CARRYB_27__37_), .S(u5_mult_82_SUMB_27__37_) );
  FA_X1 u5_mult_82_S2_27_36 ( .A(u5_mult_82_ab_27__36_), .B(
        u5_mult_82_CARRYB_26__36_), .CI(u5_mult_82_SUMB_26__37_), .CO(
        u5_mult_82_CARRYB_27__36_), .S(u5_mult_82_SUMB_27__36_) );
  FA_X1 u5_mult_82_S2_27_33 ( .A(u5_mult_82_ab_27__33_), .B(
        u5_mult_82_CARRYB_26__33_), .CI(u5_mult_82_SUMB_26__34_), .CO(
        u5_mult_82_CARRYB_27__33_), .S(u5_mult_82_SUMB_27__33_) );
  FA_X1 u5_mult_82_S2_27_30 ( .A(u5_mult_82_ab_27__30_), .B(
        u5_mult_82_CARRYB_26__30_), .CI(u5_mult_82_SUMB_26__31_), .CO(
        u5_mult_82_CARRYB_27__30_), .S(u5_mult_82_SUMB_27__30_) );
  FA_X1 u5_mult_82_S2_27_28 ( .A(u5_mult_82_ab_27__28_), .B(
        u5_mult_82_CARRYB_26__28_), .CI(u5_mult_82_SUMB_26__29_), .CO(
        u5_mult_82_CARRYB_27__28_), .S(u5_mult_82_SUMB_27__28_) );
  FA_X1 u5_mult_82_S2_27_27 ( .A(u5_mult_82_CARRYB_26__27_), .B(
        u5_mult_82_ab_27__27_), .CI(u5_mult_82_SUMB_26__28_), .CO(
        u5_mult_82_CARRYB_27__27_), .S(u5_mult_82_SUMB_27__27_) );
  FA_X1 u5_mult_82_S2_27_22 ( .A(u5_mult_82_ab_27__22_), .B(
        u5_mult_82_CARRYB_26__22_), .CI(u5_mult_82_SUMB_26__23_), .CO(
        u5_mult_82_CARRYB_27__22_), .S(u5_mult_82_SUMB_27__22_) );
  FA_X1 u5_mult_82_S2_27_19 ( .A(u5_mult_82_ab_27__19_), .B(
        u5_mult_82_CARRYB_26__19_), .CI(u5_mult_82_SUMB_26__20_), .CO(
        u5_mult_82_CARRYB_27__19_), .S(u5_mult_82_SUMB_27__19_) );
  FA_X1 u5_mult_82_S2_27_17 ( .A(u5_mult_82_ab_27__17_), .B(
        u5_mult_82_CARRYB_26__17_), .CI(u5_mult_82_SUMB_26__18_), .CO(
        u5_mult_82_CARRYB_27__17_), .S(u5_mult_82_SUMB_27__17_) );
  FA_X1 u5_mult_82_S2_27_14 ( .A(u5_mult_82_ab_27__14_), .B(
        u5_mult_82_CARRYB_26__14_), .CI(u5_mult_82_SUMB_26__15_), .CO(
        u5_mult_82_CARRYB_27__14_), .S(u5_mult_82_SUMB_27__14_) );
  FA_X1 u5_mult_82_S2_27_13 ( .A(u5_mult_82_ab_27__13_), .B(
        u5_mult_82_CARRYB_26__13_), .CI(u5_mult_82_SUMB_26__14_), .CO(
        u5_mult_82_CARRYB_27__13_), .S(u5_mult_82_SUMB_27__13_) );
  FA_X1 u5_mult_82_S2_27_12 ( .A(u5_mult_82_ab_27__12_), .B(
        u5_mult_82_CARRYB_26__12_), .CI(u5_mult_82_SUMB_26__13_), .CO(
        u5_mult_82_CARRYB_27__12_), .S(u5_mult_82_SUMB_27__12_) );
  FA_X1 u5_mult_82_S2_27_9 ( .A(u5_mult_82_ab_27__9_), .B(
        u5_mult_82_CARRYB_26__9_), .CI(u5_mult_82_SUMB_26__10_), .CO(
        u5_mult_82_CARRYB_27__9_), .S(u5_mult_82_SUMB_27__9_) );
  FA_X1 u5_mult_82_S2_27_5 ( .A(u5_mult_82_CARRYB_26__5_), .B(
        u5_mult_82_ab_27__5_), .CI(u5_mult_82_SUMB_26__6_), .CO(
        u5_mult_82_CARRYB_27__5_), .S(u5_mult_82_SUMB_27__5_) );
  FA_X1 u5_mult_82_S2_27_4 ( .A(u5_mult_82_ab_27__4_), .B(
        u5_mult_82_CARRYB_26__4_), .CI(u5_mult_82_SUMB_26__5_), .CO(
        u5_mult_82_CARRYB_27__4_), .S(u5_mult_82_SUMB_27__4_) );
  FA_X1 u5_mult_82_S2_27_3 ( .A(u5_mult_82_ab_27__3_), .B(
        u5_mult_82_CARRYB_26__3_), .CI(u5_mult_82_SUMB_26__4_), .CO(
        u5_mult_82_CARRYB_27__3_), .S(u5_mult_82_SUMB_27__3_) );
  FA_X1 u5_mult_82_S2_27_2 ( .A(u5_mult_82_ab_27__2_), .B(
        u5_mult_82_CARRYB_26__2_), .CI(u5_mult_82_SUMB_26__3_), .CO(
        u5_mult_82_CARRYB_27__2_), .S(u5_mult_82_SUMB_27__2_) );
  FA_X1 u5_mult_82_S2_27_1 ( .A(u5_mult_82_ab_27__1_), .B(
        u5_mult_82_CARRYB_26__1_), .CI(u5_mult_82_SUMB_26__2_), .CO(
        u5_mult_82_CARRYB_27__1_), .S(u5_mult_82_SUMB_27__1_) );
  FA_X1 u5_mult_82_S1_27_0 ( .A(u5_mult_82_ab_27__0_), .B(
        u5_mult_82_CARRYB_26__0_), .CI(u5_mult_82_SUMB_26__1_), .CO(
        u5_mult_82_CARRYB_27__0_), .S(u5_N27) );
  FA_X1 u5_mult_82_S3_28_51 ( .A(u5_mult_82_ab_28__51_), .B(
        u5_mult_82_CARRYB_27__51_), .CI(u5_mult_82_ab_27__52_), .CO(
        u5_mult_82_CARRYB_28__51_), .S(u5_mult_82_SUMB_28__51_) );
  FA_X1 u5_mult_82_S2_28_50 ( .A(u5_mult_82_ab_28__50_), .B(
        u5_mult_82_CARRYB_27__50_), .CI(u5_mult_82_SUMB_27__51_), .CO(
        u5_mult_82_CARRYB_28__50_), .S(u5_mult_82_SUMB_28__50_) );
  FA_X1 u5_mult_82_S2_28_49 ( .A(u5_mult_82_CARRYB_27__49_), .B(
        u5_mult_82_ab_28__49_), .CI(u5_mult_82_SUMB_27__50_), .CO(
        u5_mult_82_CARRYB_28__49_), .S(u5_mult_82_SUMB_28__49_) );
  FA_X1 u5_mult_82_S2_28_48 ( .A(u5_mult_82_ab_28__48_), .B(
        u5_mult_82_CARRYB_27__48_), .CI(u5_mult_82_SUMB_27__49_), .CO(
        u5_mult_82_CARRYB_28__48_), .S(u5_mult_82_SUMB_28__48_) );
  FA_X1 u5_mult_82_S2_28_47 ( .A(u5_mult_82_ab_28__47_), .B(
        u5_mult_82_CARRYB_27__47_), .CI(u5_mult_82_SUMB_27__48_), .CO(
        u5_mult_82_CARRYB_28__47_), .S(u5_mult_82_SUMB_28__47_) );
  FA_X1 u5_mult_82_S2_28_46 ( .A(u5_mult_82_ab_28__46_), .B(
        u5_mult_82_CARRYB_27__46_), .CI(u5_mult_82_SUMB_27__47_), .CO(
        u5_mult_82_CARRYB_28__46_), .S(u5_mult_82_SUMB_28__46_) );
  FA_X1 u5_mult_82_S2_28_45 ( .A(u5_mult_82_ab_28__45_), .B(
        u5_mult_82_CARRYB_27__45_), .CI(u5_mult_82_SUMB_27__46_), .CO(
        u5_mult_82_CARRYB_28__45_), .S(u5_mult_82_SUMB_28__45_) );
  FA_X1 u5_mult_82_S2_28_44 ( .A(u5_mult_82_CARRYB_27__44_), .B(
        u5_mult_82_ab_28__44_), .CI(u5_mult_82_SUMB_27__45_), .CO(
        u5_mult_82_CARRYB_28__44_), .S(u5_mult_82_SUMB_28__44_) );
  FA_X1 u5_mult_82_S2_28_38 ( .A(u5_mult_82_ab_28__38_), .B(
        u5_mult_82_CARRYB_27__38_), .CI(u5_mult_82_SUMB_27__39_), .CO(
        u5_mult_82_CARRYB_28__38_), .S(u5_mult_82_SUMB_28__38_) );
  FA_X1 u5_mult_82_S2_28_34 ( .A(u5_mult_82_ab_28__34_), .B(
        u5_mult_82_SUMB_27__35_), .CI(u5_mult_82_CARRYB_27__34_), .CO(
        u5_mult_82_CARRYB_28__34_), .S(u5_mult_82_SUMB_28__34_) );
  FA_X1 u5_mult_82_S2_28_28 ( .A(u5_mult_82_ab_28__28_), .B(
        u5_mult_82_CARRYB_27__28_), .CI(u5_mult_82_SUMB_27__29_), .CO(
        u5_mult_82_CARRYB_28__28_), .S(u5_mult_82_SUMB_28__28_) );
  FA_X1 u5_mult_82_S2_28_26 ( .A(u5_mult_82_ab_28__26_), .B(
        u5_mult_82_CARRYB_27__26_), .CI(u5_mult_82_SUMB_27__27_), .CO(
        u5_mult_82_CARRYB_28__26_), .S(u5_mult_82_SUMB_28__26_) );
  FA_X1 u5_mult_82_S2_28_24 ( .A(u5_mult_82_ab_28__24_), .B(
        u5_mult_82_CARRYB_27__24_), .CI(u5_mult_82_SUMB_27__25_), .CO(
        u5_mult_82_CARRYB_28__24_), .S(u5_mult_82_SUMB_28__24_) );
  FA_X1 u5_mult_82_S2_28_21 ( .A(u5_mult_82_ab_28__21_), .B(
        u5_mult_82_CARRYB_27__21_), .CI(u5_mult_82_SUMB_27__22_), .CO(
        u5_mult_82_CARRYB_28__21_), .S(u5_mult_82_SUMB_28__21_) );
  FA_X1 u5_mult_82_S2_28_18 ( .A(u5_mult_82_ab_28__18_), .B(
        u5_mult_82_CARRYB_27__18_), .CI(u5_mult_82_SUMB_27__19_), .CO(
        u5_mult_82_CARRYB_28__18_), .S(u5_mult_82_SUMB_28__18_) );
  FA_X1 u5_mult_82_S2_28_10 ( .A(u5_mult_82_ab_28__10_), .B(
        u5_mult_82_CARRYB_27__10_), .CI(u5_mult_82_SUMB_27__11_), .CO(
        u5_mult_82_CARRYB_28__10_), .S(u5_mult_82_SUMB_28__10_) );
  FA_X1 u5_mult_82_S2_28_9 ( .A(u5_mult_82_CARRYB_27__9_), .B(
        u5_mult_82_ab_28__9_), .CI(u5_mult_82_SUMB_27__10_), .CO(
        u5_mult_82_CARRYB_28__9_), .S(u5_mult_82_SUMB_28__9_) );
  FA_X1 u5_mult_82_S2_28_8 ( .A(u5_mult_82_ab_28__8_), .B(
        u5_mult_82_CARRYB_27__8_), .CI(u5_mult_82_SUMB_27__9_), .CO(
        u5_mult_82_CARRYB_28__8_), .S(u5_mult_82_SUMB_28__8_) );
  FA_X1 u5_mult_82_S2_28_7 ( .A(u5_mult_82_ab_28__7_), .B(
        u5_mult_82_CARRYB_27__7_), .CI(u5_mult_82_SUMB_27__8_), .CO(
        u5_mult_82_CARRYB_28__7_), .S(u5_mult_82_SUMB_28__7_) );
  FA_X1 u5_mult_82_S2_28_4 ( .A(u5_mult_82_ab_28__4_), .B(
        u5_mult_82_CARRYB_27__4_), .CI(u5_mult_82_SUMB_27__5_), .CO(
        u5_mult_82_CARRYB_28__4_), .S(u5_mult_82_SUMB_28__4_) );
  FA_X1 u5_mult_82_S2_28_3 ( .A(u5_mult_82_ab_28__3_), .B(
        u5_mult_82_CARRYB_27__3_), .CI(u5_mult_82_SUMB_27__4_), .CO(
        u5_mult_82_CARRYB_28__3_), .S(u5_mult_82_SUMB_28__3_) );
  FA_X1 u5_mult_82_S2_28_2 ( .A(u5_mult_82_CARRYB_27__2_), .B(
        u5_mult_82_ab_28__2_), .CI(u5_mult_82_SUMB_27__3_), .CO(
        u5_mult_82_CARRYB_28__2_), .S(u5_mult_82_SUMB_28__2_) );
  FA_X1 u5_mult_82_S2_28_1 ( .A(u5_mult_82_ab_28__1_), .B(
        u5_mult_82_CARRYB_27__1_), .CI(u5_mult_82_SUMB_27__2_), .CO(
        u5_mult_82_CARRYB_28__1_), .S(u5_mult_82_SUMB_28__1_) );
  FA_X1 u5_mult_82_S1_28_0 ( .A(u5_mult_82_ab_28__0_), .B(
        u5_mult_82_CARRYB_27__0_), .CI(u5_mult_82_SUMB_27__1_), .CO(
        u5_mult_82_CARRYB_28__0_), .S(u5_N28) );
  FA_X1 u5_mult_82_S3_29_51 ( .A(u5_mult_82_ab_29__51_), .B(
        u5_mult_82_CARRYB_28__51_), .CI(u5_mult_82_ab_28__52_), .CO(
        u5_mult_82_CARRYB_29__51_), .S(u5_mult_82_SUMB_29__51_) );
  FA_X1 u5_mult_82_S2_29_49 ( .A(u5_mult_82_ab_29__49_), .B(
        u5_mult_82_CARRYB_28__49_), .CI(u5_mult_82_SUMB_28__50_), .CO(
        u5_mult_82_CARRYB_29__49_), .S(u5_mult_82_SUMB_29__49_) );
  FA_X1 u5_mult_82_S2_29_48 ( .A(u5_mult_82_ab_29__48_), .B(
        u5_mult_82_CARRYB_28__48_), .CI(u5_mult_82_SUMB_28__49_), .CO(
        u5_mult_82_CARRYB_29__48_), .S(u5_mult_82_SUMB_29__48_) );
  FA_X1 u5_mult_82_S2_29_46 ( .A(u5_mult_82_ab_29__46_), .B(
        u5_mult_82_CARRYB_28__46_), .CI(u5_mult_82_SUMB_28__47_), .CO(
        u5_mult_82_CARRYB_29__46_), .S(u5_mult_82_SUMB_29__46_) );
  FA_X1 u5_mult_82_S2_29_45 ( .A(u5_mult_82_ab_29__45_), .B(
        u5_mult_82_CARRYB_28__45_), .CI(u5_mult_82_SUMB_28__46_), .CO(
        u5_mult_82_CARRYB_29__45_), .S(u5_mult_82_SUMB_29__45_) );
  FA_X1 u5_mult_82_S2_29_44 ( .A(u5_mult_82_ab_29__44_), .B(
        u5_mult_82_CARRYB_28__44_), .CI(u5_mult_82_SUMB_28__45_), .CO(
        u5_mult_82_CARRYB_29__44_), .S(u5_mult_82_SUMB_29__44_) );
  FA_X1 u5_mult_82_S2_29_43 ( .A(u5_mult_82_ab_29__43_), .B(
        u5_mult_82_CARRYB_28__43_), .CI(u5_mult_82_SUMB_28__44_), .CO(
        u5_mult_82_CARRYB_29__43_), .S(u5_mult_82_SUMB_29__43_) );
  FA_X1 u5_mult_82_S2_29_42 ( .A(u5_mult_82_ab_29__42_), .B(
        u5_mult_82_CARRYB_28__42_), .CI(u5_mult_82_SUMB_28__43_), .CO(
        u5_mult_82_CARRYB_29__42_), .S(u5_mult_82_SUMB_29__42_) );
  FA_X1 u5_mult_82_S2_29_35 ( .A(u5_mult_82_CARRYB_28__35_), .B(
        u5_mult_82_ab_29__35_), .CI(u5_mult_82_SUMB_28__36_), .CO(
        u5_mult_82_CARRYB_29__35_), .S(u5_mult_82_SUMB_29__35_) );
  FA_X1 u5_mult_82_S2_29_22 ( .A(u5_mult_82_CARRYB_28__22_), .B(
        u5_mult_82_ab_29__22_), .CI(u5_mult_82_SUMB_28__23_), .CO(
        u5_mult_82_CARRYB_29__22_), .S(u5_mult_82_SUMB_29__22_) );
  FA_X1 u5_mult_82_S2_29_14 ( .A(u5_mult_82_CARRYB_28__14_), .B(
        u5_mult_82_ab_29__14_), .CI(u5_mult_82_SUMB_28__15_), .CO(
        u5_mult_82_CARRYB_29__14_), .S(u5_mult_82_SUMB_29__14_) );
  FA_X1 u5_mult_82_S2_29_8 ( .A(u5_mult_82_ab_29__8_), .B(
        u5_mult_82_CARRYB_28__8_), .CI(u5_mult_82_SUMB_28__9_), .CO(
        u5_mult_82_CARRYB_29__8_), .S(u5_mult_82_SUMB_29__8_) );
  FA_X1 u5_mult_82_S2_29_7 ( .A(u5_mult_82_ab_29__7_), .B(
        u5_mult_82_CARRYB_28__7_), .CI(u5_mult_82_SUMB_28__8_), .CO(
        u5_mult_82_CARRYB_29__7_), .S(u5_mult_82_SUMB_29__7_) );
  FA_X1 u5_mult_82_S2_29_5 ( .A(u5_mult_82_ab_29__5_), .B(
        u5_mult_82_CARRYB_28__5_), .CI(u5_mult_82_SUMB_28__6_), .CO(
        u5_mult_82_CARRYB_29__5_), .S(u5_mult_82_SUMB_29__5_) );
  FA_X1 u5_mult_82_S2_29_4 ( .A(u5_mult_82_ab_29__4_), .B(
        u5_mult_82_CARRYB_28__4_), .CI(u5_mult_82_SUMB_28__5_), .CO(
        u5_mult_82_CARRYB_29__4_), .S(u5_mult_82_SUMB_29__4_) );
  FA_X1 u5_mult_82_S2_29_3 ( .A(u5_mult_82_ab_29__3_), .B(
        u5_mult_82_CARRYB_28__3_), .CI(u5_mult_82_SUMB_28__4_), .CO(
        u5_mult_82_CARRYB_29__3_), .S(u5_mult_82_SUMB_29__3_) );
  FA_X1 u5_mult_82_S2_29_2 ( .A(u5_mult_82_ab_29__2_), .B(
        u5_mult_82_CARRYB_28__2_), .CI(u5_mult_82_SUMB_28__3_), .CO(
        u5_mult_82_CARRYB_29__2_), .S(u5_mult_82_SUMB_29__2_) );
  FA_X1 u5_mult_82_S2_29_1 ( .A(u5_mult_82_ab_29__1_), .B(
        u5_mult_82_CARRYB_28__1_), .CI(u5_mult_82_SUMB_28__2_), .CO(
        u5_mult_82_CARRYB_29__1_), .S(u5_mult_82_SUMB_29__1_) );
  FA_X1 u5_mult_82_S1_29_0 ( .A(u5_mult_82_ab_29__0_), .B(
        u5_mult_82_CARRYB_28__0_), .CI(u5_mult_82_SUMB_28__1_), .CO(
        u5_mult_82_CARRYB_29__0_), .S(u5_N29) );
  FA_X1 u5_mult_82_S3_30_51 ( .A(u5_mult_82_ab_30__51_), .B(
        u5_mult_82_CARRYB_29__51_), .CI(u5_mult_82_ab_29__52_), .CO(
        u5_mult_82_CARRYB_30__51_), .S(u5_mult_82_SUMB_30__51_) );
  FA_X1 u5_mult_82_S2_30_50 ( .A(u5_mult_82_ab_30__50_), .B(
        u5_mult_82_CARRYB_29__50_), .CI(u5_mult_82_SUMB_29__51_), .CO(
        u5_mult_82_CARRYB_30__50_), .S(u5_mult_82_SUMB_30__50_) );
  FA_X1 u5_mult_82_S2_30_48 ( .A(u5_mult_82_ab_30__48_), .B(
        u5_mult_82_CARRYB_29__48_), .CI(u5_mult_82_SUMB_29__49_), .CO(
        u5_mult_82_CARRYB_30__48_), .S(u5_mult_82_SUMB_30__48_) );
  FA_X1 u5_mult_82_S2_30_47 ( .A(u5_mult_82_ab_30__47_), .B(
        u5_mult_82_CARRYB_29__47_), .CI(u5_mult_82_SUMB_29__48_), .CO(
        u5_mult_82_CARRYB_30__47_), .S(u5_mult_82_SUMB_30__47_) );
  FA_X1 u5_mult_82_S2_30_46 ( .A(u5_mult_82_CARRYB_29__46_), .B(
        u5_mult_82_ab_30__46_), .CI(u5_mult_82_SUMB_29__47_), .CO(
        u5_mult_82_CARRYB_30__46_), .S(u5_mult_82_SUMB_30__46_) );
  FA_X1 u5_mult_82_S2_30_45 ( .A(u5_mult_82_ab_30__45_), .B(
        u5_mult_82_CARRYB_29__45_), .CI(u5_mult_82_SUMB_29__46_), .CO(
        u5_mult_82_CARRYB_30__45_), .S(u5_mult_82_SUMB_30__45_) );
  FA_X1 u5_mult_82_S2_30_44 ( .A(u5_mult_82_ab_30__44_), .B(
        u5_mult_82_CARRYB_29__44_), .CI(u5_mult_82_SUMB_29__45_), .CO(
        u5_mult_82_CARRYB_30__44_), .S(u5_mult_82_SUMB_30__44_) );
  FA_X1 u5_mult_82_S2_30_43 ( .A(u5_mult_82_CARRYB_29__43_), .B(
        u5_mult_82_ab_30__43_), .CI(u5_mult_82_SUMB_29__44_), .CO(
        u5_mult_82_CARRYB_30__43_), .S(u5_mult_82_SUMB_30__43_) );
  FA_X1 u5_mult_82_S2_30_42 ( .A(u5_mult_82_CARRYB_29__42_), .B(
        u5_mult_82_ab_30__42_), .CI(u5_mult_82_SUMB_29__43_), .CO(
        u5_mult_82_CARRYB_30__42_), .S(u5_mult_82_SUMB_30__42_) );
  FA_X1 u5_mult_82_S2_30_41 ( .A(u5_mult_82_ab_30__41_), .B(
        u5_mult_82_CARRYB_29__41_), .CI(u5_mult_82_SUMB_29__42_), .CO(
        u5_mult_82_CARRYB_30__41_), .S(u5_mult_82_SUMB_30__41_) );
  FA_X1 u5_mult_82_S2_30_40 ( .A(u5_mult_82_ab_30__40_), .B(
        u5_mult_82_CARRYB_29__40_), .CI(u5_mult_82_SUMB_29__41_), .CO(
        u5_mult_82_CARRYB_30__40_), .S(u5_mult_82_SUMB_30__40_) );
  FA_X1 u5_mult_82_S2_30_35 ( .A(u5_mult_82_CARRYB_29__35_), .B(
        u5_mult_82_ab_30__35_), .CI(u5_mult_82_SUMB_29__36_), .CO(
        u5_mult_82_CARRYB_30__35_), .S(u5_mult_82_SUMB_30__35_) );
  FA_X1 u5_mult_82_S2_30_34 ( .A(u5_mult_82_ab_30__34_), .B(
        u5_mult_82_CARRYB_29__34_), .CI(u5_mult_82_SUMB_29__35_), .CO(
        u5_mult_82_CARRYB_30__34_), .S(u5_mult_82_SUMB_30__34_) );
  FA_X1 u5_mult_82_S2_30_33 ( .A(u5_mult_82_ab_30__33_), .B(
        u5_mult_82_CARRYB_29__33_), .CI(u5_mult_82_SUMB_29__34_), .CO(
        u5_mult_82_CARRYB_30__33_), .S(u5_mult_82_SUMB_30__33_) );
  FA_X1 u5_mult_82_S2_30_28 ( .A(u5_mult_82_ab_30__28_), .B(
        u5_mult_82_CARRYB_29__28_), .CI(u5_mult_82_SUMB_29__29_), .CO(
        u5_mult_82_CARRYB_30__28_), .S(u5_mult_82_SUMB_30__28_) );
  FA_X1 u5_mult_82_S2_30_25 ( .A(u5_mult_82_CARRYB_29__25_), .B(
        u5_mult_82_ab_30__25_), .CI(u5_mult_82_SUMB_29__26_), .CO(
        u5_mult_82_CARRYB_30__25_), .S(u5_mult_82_SUMB_30__25_) );
  FA_X1 u5_mult_82_S2_30_21 ( .A(u5_mult_82_ab_30__21_), .B(
        u5_mult_82_CARRYB_29__21_), .CI(u5_mult_82_SUMB_29__22_), .CO(
        u5_mult_82_CARRYB_30__21_), .S(u5_mult_82_SUMB_30__21_) );
  FA_X1 u5_mult_82_S2_30_14 ( .A(u5_mult_82_ab_30__14_), .B(
        u5_mult_82_CARRYB_29__14_), .CI(u5_mult_82_SUMB_29__15_), .CO(
        u5_mult_82_CARRYB_30__14_), .S(u5_mult_82_SUMB_30__14_) );
  FA_X1 u5_mult_82_S2_30_13 ( .A(u5_mult_82_ab_30__13_), .B(
        u5_mult_82_CARRYB_29__13_), .CI(u5_mult_82_SUMB_29__14_), .CO(
        u5_mult_82_CARRYB_30__13_), .S(u5_mult_82_SUMB_30__13_) );
  FA_X1 u5_mult_82_S2_30_12 ( .A(u5_mult_82_ab_30__12_), .B(
        u5_mult_82_CARRYB_29__12_), .CI(u5_mult_82_SUMB_29__13_), .CO(
        u5_mult_82_CARRYB_30__12_), .S(u5_mult_82_SUMB_30__12_) );
  FA_X1 u5_mult_82_S2_30_9 ( .A(u5_mult_82_ab_30__9_), .B(
        u5_mult_82_CARRYB_29__9_), .CI(u5_mult_82_SUMB_29__10_), .CO(
        u5_mult_82_CARRYB_30__9_), .S(u5_mult_82_SUMB_30__9_) );
  FA_X1 u5_mult_82_S2_30_7 ( .A(u5_mult_82_CARRYB_29__7_), .B(
        u5_mult_82_ab_30__7_), .CI(u5_mult_82_SUMB_29__8_), .CO(
        u5_mult_82_CARRYB_30__7_), .S(u5_mult_82_SUMB_30__7_) );
  FA_X1 u5_mult_82_S2_30_5 ( .A(u5_mult_82_ab_30__5_), .B(
        u5_mult_82_CARRYB_29__5_), .CI(u5_mult_82_SUMB_29__6_), .CO(
        u5_mult_82_CARRYB_30__5_), .S(u5_mult_82_SUMB_30__5_) );
  FA_X1 u5_mult_82_S2_30_4 ( .A(u5_mult_82_SUMB_29__5_), .B(
        u5_mult_82_ab_30__4_), .CI(u5_mult_82_CARRYB_29__4_), .CO(
        u5_mult_82_CARRYB_30__4_), .S(u5_mult_82_SUMB_30__4_) );
  FA_X1 u5_mult_82_S2_30_3 ( .A(u5_mult_82_ab_30__3_), .B(
        u5_mult_82_CARRYB_29__3_), .CI(u5_mult_82_SUMB_29__4_), .CO(
        u5_mult_82_CARRYB_30__3_), .S(u5_mult_82_SUMB_30__3_) );
  FA_X1 u5_mult_82_S2_30_2 ( .A(u5_mult_82_CARRYB_29__2_), .B(
        u5_mult_82_ab_30__2_), .CI(u5_mult_82_SUMB_29__3_), .CO(
        u5_mult_82_CARRYB_30__2_), .S(u5_mult_82_SUMB_30__2_) );
  FA_X1 u5_mult_82_S2_30_1 ( .A(u5_mult_82_ab_30__1_), .B(
        u5_mult_82_CARRYB_29__1_), .CI(u5_mult_82_SUMB_29__2_), .CO(
        u5_mult_82_CARRYB_30__1_), .S(u5_mult_82_SUMB_30__1_) );
  FA_X1 u5_mult_82_S1_30_0 ( .A(u5_mult_82_ab_30__0_), .B(
        u5_mult_82_CARRYB_29__0_), .CI(u5_mult_82_SUMB_29__1_), .CO(
        u5_mult_82_CARRYB_30__0_), .S(u5_N30) );
  FA_X1 u5_mult_82_S3_31_51 ( .A(u5_mult_82_ab_31__51_), .B(
        u5_mult_82_CARRYB_30__51_), .CI(u5_mult_82_ab_30__52_), .CO(
        u5_mult_82_CARRYB_31__51_), .S(u5_mult_82_SUMB_31__51_) );
  FA_X1 u5_mult_82_S2_31_50 ( .A(u5_mult_82_ab_31__50_), .B(
        u5_mult_82_CARRYB_30__50_), .CI(u5_mult_82_SUMB_30__51_), .CO(
        u5_mult_82_CARRYB_31__50_), .S(u5_mult_82_SUMB_31__50_) );
  FA_X1 u5_mult_82_S2_31_49 ( .A(u5_mult_82_ab_31__49_), .B(
        u5_mult_82_CARRYB_30__49_), .CI(u5_mult_82_SUMB_30__50_), .CO(
        u5_mult_82_CARRYB_31__49_), .S(u5_mult_82_SUMB_31__49_) );
  FA_X1 u5_mult_82_S2_31_48 ( .A(u5_mult_82_ab_31__48_), .B(
        u5_mult_82_CARRYB_30__48_), .CI(u5_mult_82_SUMB_30__49_), .CO(
        u5_mult_82_CARRYB_31__48_), .S(u5_mult_82_SUMB_31__48_) );
  FA_X1 u5_mult_82_S2_31_47 ( .A(u5_mult_82_ab_31__47_), .B(
        u5_mult_82_CARRYB_30__47_), .CI(u5_mult_82_SUMB_30__48_), .CO(
        u5_mult_82_CARRYB_31__47_), .S(u5_mult_82_SUMB_31__47_) );
  FA_X1 u5_mult_82_S2_31_46 ( .A(u5_mult_82_ab_31__46_), .B(
        u5_mult_82_CARRYB_30__46_), .CI(u5_mult_82_SUMB_30__47_), .CO(
        u5_mult_82_CARRYB_31__46_), .S(u5_mult_82_SUMB_31__46_) );
  FA_X1 u5_mult_82_S2_31_44 ( .A(u5_mult_82_ab_31__44_), .B(
        u5_mult_82_CARRYB_30__44_), .CI(u5_mult_82_SUMB_30__45_), .CO(
        u5_mult_82_CARRYB_31__44_), .S(u5_mult_82_SUMB_31__44_) );
  FA_X1 u5_mult_82_S2_31_43 ( .A(u5_mult_82_ab_31__43_), .B(
        u5_mult_82_CARRYB_30__43_), .CI(u5_mult_82_SUMB_30__44_), .CO(
        u5_mult_82_CARRYB_31__43_), .S(u5_mult_82_SUMB_31__43_) );
  FA_X1 u5_mult_82_S2_31_42 ( .A(u5_mult_82_CARRYB_30__42_), .B(
        u5_mult_82_ab_31__42_), .CI(u5_mult_82_SUMB_30__43_), .CO(
        u5_mult_82_CARRYB_31__42_), .S(u5_mult_82_SUMB_31__42_) );
  FA_X1 u5_mult_82_S2_31_41 ( .A(u5_mult_82_CARRYB_30__41_), .B(
        u5_mult_82_ab_31__41_), .CI(u5_mult_82_SUMB_30__42_), .CO(
        u5_mult_82_CARRYB_31__41_), .S(u5_mult_82_SUMB_31__41_) );
  FA_X1 u5_mult_82_S2_31_40 ( .A(u5_mult_82_ab_31__40_), .B(
        u5_mult_82_CARRYB_30__40_), .CI(u5_mult_82_SUMB_30__41_), .CO(
        u5_mult_82_CARRYB_31__40_), .S(u5_mult_82_SUMB_31__40_) );
  FA_X1 u5_mult_82_S2_31_38 ( .A(u5_mult_82_ab_31__38_), .B(
        u5_mult_82_CARRYB_30__38_), .CI(u5_mult_82_SUMB_30__39_), .CO(
        u5_mult_82_CARRYB_31__38_), .S(u5_mult_82_SUMB_31__38_) );
  FA_X1 u5_mult_82_S2_31_37 ( .A(u5_mult_82_ab_31__37_), .B(
        u5_mult_82_CARRYB_30__37_), .CI(u5_mult_82_SUMB_30__38_), .CO(
        u5_mult_82_CARRYB_31__37_), .S(u5_mult_82_SUMB_31__37_) );
  FA_X1 u5_mult_82_S2_31_35 ( .A(u5_mult_82_ab_31__35_), .B(
        u5_mult_82_CARRYB_30__35_), .CI(u5_mult_82_SUMB_30__36_), .CO(
        u5_mult_82_CARRYB_31__35_), .S(u5_mult_82_SUMB_31__35_) );
  FA_X1 u5_mult_82_S2_31_34 ( .A(u5_mult_82_ab_31__34_), .B(
        u5_mult_82_CARRYB_30__34_), .CI(u5_mult_82_SUMB_30__35_), .CO(
        u5_mult_82_CARRYB_31__34_), .S(u5_mult_82_SUMB_31__34_) );
  FA_X1 u5_mult_82_S2_31_33 ( .A(u5_mult_82_ab_31__33_), .B(
        u5_mult_82_CARRYB_30__33_), .CI(u5_mult_82_SUMB_30__34_), .CO(
        u5_mult_82_CARRYB_31__33_), .S(u5_mult_82_SUMB_31__33_) );
  FA_X1 u5_mult_82_S2_31_32 ( .A(u5_mult_82_ab_31__32_), .B(
        u5_mult_82_CARRYB_30__32_), .CI(u5_mult_82_SUMB_30__33_), .CO(
        u5_mult_82_CARRYB_31__32_), .S(u5_mult_82_SUMB_31__32_) );
  FA_X1 u5_mult_82_S2_31_31 ( .A(u5_mult_82_CARRYB_30__31_), .B(
        u5_mult_82_ab_31__31_), .CI(u5_mult_82_SUMB_30__32_), .CO(
        u5_mult_82_CARRYB_31__31_), .S(u5_mult_82_SUMB_31__31_) );
  FA_X1 u5_mult_82_S2_31_27 ( .A(u5_mult_82_ab_31__27_), .B(
        u5_mult_82_CARRYB_30__27_), .CI(u5_mult_82_SUMB_30__28_), .CO(
        u5_mult_82_CARRYB_31__27_), .S(u5_mult_82_SUMB_31__27_) );
  FA_X1 u5_mult_82_S2_31_26 ( .A(u5_mult_82_ab_31__26_), .B(
        u5_mult_82_CARRYB_30__26_), .CI(u5_mult_82_SUMB_30__27_), .CO(
        u5_mult_82_CARRYB_31__26_), .S(u5_mult_82_SUMB_31__26_) );
  FA_X1 u5_mult_82_S2_31_24 ( .A(u5_mult_82_ab_31__24_), .B(
        u5_mult_82_CARRYB_30__24_), .CI(u5_mult_82_SUMB_30__25_), .CO(
        u5_mult_82_CARRYB_31__24_), .S(u5_mult_82_SUMB_31__24_) );
  FA_X1 u5_mult_82_S2_31_21 ( .A(u5_mult_82_ab_31__21_), .B(
        u5_mult_82_CARRYB_30__21_), .CI(u5_mult_82_SUMB_30__22_), .CO(
        u5_mult_82_CARRYB_31__21_), .S(u5_mult_82_SUMB_31__21_) );
  FA_X1 u5_mult_82_S2_31_20 ( .A(u5_mult_82_ab_31__20_), .B(
        u5_mult_82_CARRYB_30__20_), .CI(u5_mult_82_SUMB_30__21_), .CO(
        u5_mult_82_CARRYB_31__20_), .S(u5_mult_82_SUMB_31__20_) );
  FA_X1 u5_mult_82_S2_31_11 ( .A(u5_mult_82_ab_31__11_), .B(
        u5_mult_82_CARRYB_30__11_), .CI(u5_mult_82_SUMB_30__12_), .CO(
        u5_mult_82_CARRYB_31__11_), .S(u5_mult_82_SUMB_31__11_) );
  FA_X1 u5_mult_82_S2_31_9 ( .A(u5_mult_82_CARRYB_30__9_), .B(
        u5_mult_82_ab_31__9_), .CI(u5_mult_82_SUMB_30__10_), .CO(
        u5_mult_82_CARRYB_31__9_), .S(u5_mult_82_SUMB_31__9_) );
  FA_X1 u5_mult_82_S2_31_7 ( .A(u5_mult_82_ab_31__7_), .B(
        u5_mult_82_SUMB_30__8_), .CI(u5_mult_82_CARRYB_30__7_), .CO(
        u5_mult_82_CARRYB_31__7_), .S(u5_mult_82_SUMB_31__7_) );
  FA_X1 u5_mult_82_S2_31_5 ( .A(u5_mult_82_CARRYB_30__5_), .B(
        u5_mult_82_ab_31__5_), .CI(u5_mult_82_SUMB_30__6_), .CO(
        u5_mult_82_CARRYB_31__5_), .S(u5_mult_82_SUMB_31__5_) );
  FA_X1 u5_mult_82_S2_31_4 ( .A(u5_mult_82_ab_31__4_), .B(
        u5_mult_82_CARRYB_30__4_), .CI(u5_mult_82_SUMB_30__5_), .CO(
        u5_mult_82_CARRYB_31__4_), .S(u5_mult_82_SUMB_31__4_) );
  FA_X1 u5_mult_82_S2_31_2 ( .A(u5_mult_82_ab_31__2_), .B(
        u5_mult_82_CARRYB_30__2_), .CI(u5_mult_82_SUMB_30__3_), .CO(
        u5_mult_82_CARRYB_31__2_), .S(u5_mult_82_SUMB_31__2_) );
  FA_X1 u5_mult_82_S2_31_1 ( .A(u5_mult_82_ab_31__1_), .B(
        u5_mult_82_CARRYB_30__1_), .CI(u5_mult_82_SUMB_30__2_), .CO(
        u5_mult_82_CARRYB_31__1_), .S(u5_mult_82_SUMB_31__1_) );
  FA_X1 u5_mult_82_S1_31_0 ( .A(u5_mult_82_ab_31__0_), .B(
        u5_mult_82_CARRYB_30__0_), .CI(u5_mult_82_SUMB_30__1_), .CO(
        u5_mult_82_CARRYB_31__0_), .S(u5_N31) );
  FA_X1 u5_mult_82_S2_32_50 ( .A(u5_mult_82_ab_32__50_), .B(
        u5_mult_82_CARRYB_31__50_), .CI(u5_mult_82_SUMB_31__51_), .CO(
        u5_mult_82_CARRYB_32__50_), .S(u5_mult_82_SUMB_32__50_) );
  FA_X1 u5_mult_82_S2_32_49 ( .A(u5_mult_82_ab_32__49_), .B(
        u5_mult_82_CARRYB_31__49_), .CI(u5_mult_82_SUMB_31__50_), .CO(
        u5_mult_82_CARRYB_32__49_), .S(u5_mult_82_SUMB_32__49_) );
  FA_X1 u5_mult_82_S2_32_48 ( .A(u5_mult_82_ab_32__48_), .B(
        u5_mult_82_CARRYB_31__48_), .CI(u5_mult_82_SUMB_31__49_), .CO(
        u5_mult_82_CARRYB_32__48_), .S(u5_mult_82_SUMB_32__48_) );
  FA_X1 u5_mult_82_S2_32_47 ( .A(u5_mult_82_ab_32__47_), .B(
        u5_mult_82_CARRYB_31__47_), .CI(u5_mult_82_SUMB_31__48_), .CO(
        u5_mult_82_CARRYB_32__47_), .S(u5_mult_82_SUMB_32__47_) );
  FA_X1 u5_mult_82_S2_32_46 ( .A(u5_mult_82_ab_32__46_), .B(
        u5_mult_82_CARRYB_31__46_), .CI(u5_mult_82_SUMB_31__47_), .CO(
        u5_mult_82_CARRYB_32__46_), .S(u5_mult_82_SUMB_32__46_) );
  FA_X1 u5_mult_82_S2_32_45 ( .A(u5_mult_82_ab_32__45_), .B(
        u5_mult_82_CARRYB_31__45_), .CI(u5_mult_82_SUMB_31__46_), .CO(
        u5_mult_82_CARRYB_32__45_), .S(u5_mult_82_SUMB_32__45_) );
  FA_X1 u5_mult_82_S2_32_42 ( .A(u5_mult_82_ab_32__42_), .B(
        u5_mult_82_CARRYB_31__42_), .CI(u5_mult_82_SUMB_31__43_), .CO(
        u5_mult_82_CARRYB_32__42_), .S(u5_mult_82_SUMB_32__42_) );
  FA_X1 u5_mult_82_S2_32_37 ( .A(u5_mult_82_ab_32__37_), .B(
        u5_mult_82_CARRYB_31__37_), .CI(u5_mult_82_SUMB_31__38_), .CO(
        u5_mult_82_CARRYB_32__37_), .S(u5_mult_82_SUMB_32__37_) );
  FA_X1 u5_mult_82_S2_32_35 ( .A(u5_mult_82_ab_32__35_), .B(
        u5_mult_82_CARRYB_31__35_), .CI(u5_mult_82_SUMB_31__36_), .CO(
        u5_mult_82_CARRYB_32__35_), .S(u5_mult_82_SUMB_32__35_) );
  FA_X1 u5_mult_82_S2_32_34 ( .A(u5_mult_82_CARRYB_31__34_), .B(
        u5_mult_82_ab_32__34_), .CI(u5_mult_82_SUMB_31__35_), .CO(
        u5_mult_82_CARRYB_32__34_), .S(u5_mult_82_SUMB_32__34_) );
  FA_X1 u5_mult_82_S2_32_33 ( .A(u5_mult_82_ab_32__33_), .B(
        u5_mult_82_CARRYB_31__33_), .CI(u5_mult_82_SUMB_31__34_), .CO(
        u5_mult_82_CARRYB_32__33_), .S(u5_mult_82_SUMB_32__33_) );
  FA_X1 u5_mult_82_S2_32_23 ( .A(u5_mult_82_ab_32__23_), .B(
        u5_mult_82_CARRYB_31__23_), .CI(u5_mult_82_SUMB_31__24_), .CO(
        u5_mult_82_CARRYB_32__23_), .S(u5_mult_82_SUMB_32__23_) );
  FA_X1 u5_mult_82_S2_32_21 ( .A(u5_mult_82_ab_32__21_), .B(
        u5_mult_82_CARRYB_31__21_), .CI(u5_mult_82_SUMB_31__22_), .CO(
        u5_mult_82_CARRYB_32__21_), .S(u5_mult_82_SUMB_32__21_) );
  FA_X1 u5_mult_82_S2_32_19 ( .A(u5_mult_82_ab_32__19_), .B(
        u5_mult_82_CARRYB_31__19_), .CI(u5_mult_82_SUMB_31__20_), .CO(
        u5_mult_82_CARRYB_32__19_), .S(u5_mult_82_SUMB_32__19_) );
  FA_X1 u5_mult_82_S2_32_18 ( .A(u5_mult_82_ab_32__18_), .B(
        u5_mult_82_CARRYB_31__18_), .CI(u5_mult_82_SUMB_31__19_), .CO(
        u5_mult_82_CARRYB_32__18_), .S(u5_mult_82_SUMB_32__18_) );
  FA_X1 u5_mult_82_S2_32_16 ( .A(u5_mult_82_ab_32__16_), .B(
        u5_mult_82_CARRYB_31__16_), .CI(u5_mult_82_SUMB_31__17_), .CO(
        u5_mult_82_CARRYB_32__16_), .S(u5_mult_82_SUMB_32__16_) );
  FA_X1 u5_mult_82_S2_32_15 ( .A(u5_mult_82_CARRYB_31__15_), .B(
        u5_mult_82_ab_32__15_), .CI(u5_mult_82_SUMB_31__16_), .CO(
        u5_mult_82_CARRYB_32__15_), .S(u5_mult_82_SUMB_32__15_) );
  FA_X1 u5_mult_82_S2_32_10 ( .A(u5_mult_82_ab_32__10_), .B(
        u5_mult_82_CARRYB_31__10_), .CI(u5_mult_82_SUMB_31__11_), .CO(
        u5_mult_82_CARRYB_32__10_), .S(u5_mult_82_SUMB_32__10_) );
  FA_X1 u5_mult_82_S2_32_9 ( .A(u5_mult_82_CARRYB_31__9_), .B(
        u5_mult_82_ab_32__9_), .CI(u5_mult_82_SUMB_31__10_), .CO(
        u5_mult_82_CARRYB_32__9_), .S(u5_mult_82_SUMB_32__9_) );
  FA_X1 u5_mult_82_S2_32_6 ( .A(u5_mult_82_ab_32__6_), .B(
        u5_mult_82_CARRYB_31__6_), .CI(u5_mult_82_SUMB_31__7_), .CO(
        u5_mult_82_CARRYB_32__6_), .S(u5_mult_82_SUMB_32__6_) );
  FA_X1 u5_mult_82_S2_32_4 ( .A(u5_mult_82_ab_32__4_), .B(
        u5_mult_82_CARRYB_31__4_), .CI(u5_mult_82_SUMB_31__5_), .CO(
        u5_mult_82_CARRYB_32__4_), .S(u5_mult_82_SUMB_32__4_) );
  FA_X1 u5_mult_82_S2_32_3 ( .A(u5_mult_82_ab_32__3_), .B(
        u5_mult_82_CARRYB_31__3_), .CI(u5_mult_82_SUMB_31__4_), .CO(
        u5_mult_82_CARRYB_32__3_), .S(u5_mult_82_SUMB_32__3_) );
  FA_X1 u5_mult_82_S2_32_2 ( .A(u5_mult_82_ab_32__2_), .B(
        u5_mult_82_CARRYB_31__2_), .CI(u5_mult_82_SUMB_31__3_), .CO(
        u5_mult_82_CARRYB_32__2_), .S(u5_mult_82_SUMB_32__2_) );
  FA_X1 u5_mult_82_S2_32_1 ( .A(u5_mult_82_ab_32__1_), .B(
        u5_mult_82_CARRYB_31__1_), .CI(u5_mult_82_SUMB_31__2_), .CO(
        u5_mult_82_CARRYB_32__1_), .S(u5_mult_82_SUMB_32__1_) );
  FA_X1 u5_mult_82_S1_32_0 ( .A(u5_mult_82_ab_32__0_), .B(
        u5_mult_82_CARRYB_31__0_), .CI(u5_mult_82_SUMB_31__1_), .CO(
        u5_mult_82_CARRYB_32__0_), .S(u5_N32) );
  FA_X1 u5_mult_82_S2_33_50 ( .A(u5_mult_82_ab_33__50_), .B(
        u5_mult_82_CARRYB_32__50_), .CI(u5_mult_82_SUMB_32__51_), .CO(
        u5_mult_82_CARRYB_33__50_), .S(u5_mult_82_SUMB_33__50_) );
  FA_X1 u5_mult_82_S2_33_49 ( .A(u5_mult_82_ab_33__49_), .B(
        u5_mult_82_CARRYB_32__49_), .CI(u5_mult_82_SUMB_32__50_), .CO(
        u5_mult_82_CARRYB_33__49_), .S(u5_mult_82_SUMB_33__49_) );
  FA_X1 u5_mult_82_S2_33_48 ( .A(u5_mult_82_ab_33__48_), .B(
        u5_mult_82_CARRYB_32__48_), .CI(u5_mult_82_SUMB_32__49_), .CO(
        u5_mult_82_CARRYB_33__48_), .S(u5_mult_82_SUMB_33__48_) );
  FA_X1 u5_mult_82_S2_33_47 ( .A(u5_mult_82_CARRYB_32__47_), .B(
        u5_mult_82_ab_33__47_), .CI(u5_mult_82_SUMB_32__48_), .CO(
        u5_mult_82_CARRYB_33__47_), .S(u5_mult_82_SUMB_33__47_) );
  FA_X1 u5_mult_82_S2_33_46 ( .A(u5_mult_82_ab_33__46_), .B(
        u5_mult_82_CARRYB_32__46_), .CI(u5_mult_82_SUMB_32__47_), .CO(
        u5_mult_82_CARRYB_33__46_), .S(u5_mult_82_SUMB_33__46_) );
  FA_X1 u5_mult_82_S2_33_45 ( .A(u5_mult_82_CARRYB_32__45_), .B(
        u5_mult_82_ab_33__45_), .CI(u5_mult_82_SUMB_32__46_), .CO(
        u5_mult_82_CARRYB_33__45_), .S(u5_mult_82_SUMB_33__45_) );
  FA_X1 u5_mult_82_S2_33_44 ( .A(u5_mult_82_ab_33__44_), .B(
        u5_mult_82_CARRYB_32__44_), .CI(u5_mult_82_SUMB_32__45_), .CO(
        u5_mult_82_CARRYB_33__44_), .S(u5_mult_82_SUMB_33__44_) );
  FA_X1 u5_mult_82_S2_33_43 ( .A(u5_mult_82_ab_33__43_), .B(
        u5_mult_82_CARRYB_32__43_), .CI(u5_mult_82_SUMB_32__44_), .CO(
        u5_mult_82_CARRYB_33__43_), .S(u5_mult_82_SUMB_33__43_) );
  FA_X1 u5_mult_82_S2_33_38 ( .A(u5_mult_82_ab_33__38_), .B(
        u5_mult_82_CARRYB_32__38_), .CI(u5_mult_82_SUMB_32__39_), .CO(
        u5_mult_82_CARRYB_33__38_), .S(u5_mult_82_SUMB_33__38_) );
  FA_X1 u5_mult_82_S2_33_37 ( .A(u5_mult_82_ab_33__37_), .B(
        u5_mult_82_CARRYB_32__37_), .CI(u5_mult_82_SUMB_32__38_), .CO(
        u5_mult_82_CARRYB_33__37_), .S(u5_mult_82_SUMB_33__37_) );
  FA_X1 u5_mult_82_S2_33_36 ( .A(u5_mult_82_ab_33__36_), .B(
        u5_mult_82_CARRYB_32__36_), .CI(u5_mult_82_SUMB_32__37_), .CO(
        u5_mult_82_CARRYB_33__36_), .S(u5_mult_82_SUMB_33__36_) );
  FA_X1 u5_mult_82_S2_33_34 ( .A(u5_mult_82_ab_33__34_), .B(
        u5_mult_82_CARRYB_32__34_), .CI(u5_mult_82_SUMB_32__35_), .CO(
        u5_mult_82_CARRYB_33__34_), .S(u5_mult_82_SUMB_33__34_) );
  FA_X1 u5_mult_82_S2_33_33 ( .A(u5_mult_82_ab_33__33_), .B(
        u5_mult_82_CARRYB_32__33_), .CI(u5_mult_82_SUMB_32__34_), .CO(
        u5_mult_82_CARRYB_33__33_), .S(u5_mult_82_SUMB_33__33_) );
  FA_X1 u5_mult_82_S2_33_28 ( .A(u5_mult_82_ab_33__28_), .B(
        u5_mult_82_CARRYB_32__28_), .CI(u5_mult_82_SUMB_32__29_), .CO(
        u5_mult_82_CARRYB_33__28_), .S(u5_mult_82_SUMB_33__28_) );
  FA_X1 u5_mult_82_S2_33_27 ( .A(u5_mult_82_ab_33__27_), .B(
        u5_mult_82_CARRYB_32__27_), .CI(u5_mult_82_SUMB_32__28_), .CO(
        u5_mult_82_CARRYB_33__27_), .S(u5_mult_82_SUMB_33__27_) );
  FA_X1 u5_mult_82_S2_33_21 ( .A(u5_mult_82_ab_33__21_), .B(
        u5_mult_82_CARRYB_32__21_), .CI(u5_mult_82_SUMB_32__22_), .CO(
        u5_mult_82_CARRYB_33__21_), .S(u5_mult_82_SUMB_33__21_) );
  FA_X1 u5_mult_82_S2_33_16 ( .A(u5_mult_82_ab_33__16_), .B(
        u5_mult_82_CARRYB_32__16_), .CI(u5_mult_82_SUMB_32__17_), .CO(
        u5_mult_82_CARRYB_33__16_), .S(u5_mult_82_SUMB_33__16_) );
  FA_X1 u5_mult_82_S2_33_15 ( .A(u5_mult_82_ab_33__15_), .B(
        u5_mult_82_CARRYB_32__15_), .CI(u5_mult_82_SUMB_32__16_), .CO(
        u5_mult_82_CARRYB_33__15_), .S(u5_mult_82_SUMB_33__15_) );
  FA_X1 u5_mult_82_S2_33_12 ( .A(u5_mult_82_SUMB_32__13_), .B(
        u5_mult_82_ab_33__12_), .CI(u5_mult_82_CARRYB_32__12_), .CO(
        u5_mult_82_CARRYB_33__12_), .S(u5_mult_82_SUMB_33__12_) );
  FA_X1 u5_mult_82_S2_33_6 ( .A(u5_mult_82_ab_33__6_), .B(
        u5_mult_82_CARRYB_32__6_), .CI(u5_mult_82_SUMB_32__7_), .CO(
        u5_mult_82_CARRYB_33__6_), .S(u5_mult_82_SUMB_33__6_) );
  FA_X1 u5_mult_82_S2_33_3 ( .A(u5_mult_82_ab_33__3_), .B(
        u5_mult_82_CARRYB_32__3_), .CI(u5_mult_82_SUMB_32__4_), .CO(
        u5_mult_82_CARRYB_33__3_), .S(u5_mult_82_SUMB_33__3_) );
  FA_X1 u5_mult_82_S2_33_2 ( .A(u5_mult_82_ab_33__2_), .B(
        u5_mult_82_CARRYB_32__2_), .CI(u5_mult_82_SUMB_32__3_), .CO(
        u5_mult_82_CARRYB_33__2_), .S(u5_mult_82_SUMB_33__2_) );
  FA_X1 u5_mult_82_S2_33_1 ( .A(u5_mult_82_ab_33__1_), .B(
        u5_mult_82_CARRYB_32__1_), .CI(u5_mult_82_SUMB_32__2_), .CO(
        u5_mult_82_CARRYB_33__1_), .S(u5_mult_82_SUMB_33__1_) );
  FA_X1 u5_mult_82_S1_33_0 ( .A(u5_mult_82_ab_33__0_), .B(
        u5_mult_82_CARRYB_32__0_), .CI(u5_mult_82_SUMB_32__1_), .CO(
        u5_mult_82_CARRYB_33__0_), .S(u5_N33) );
  FA_X1 u5_mult_82_S3_34_51 ( .A(u5_mult_82_ab_34__51_), .B(
        u5_mult_82_CARRYB_33__51_), .CI(u5_mult_82_ab_33__52_), .CO(
        u5_mult_82_CARRYB_34__51_), .S(u5_mult_82_SUMB_34__51_) );
  FA_X1 u5_mult_82_S2_34_50 ( .A(u5_mult_82_ab_34__50_), .B(
        u5_mult_82_CARRYB_33__50_), .CI(u5_mult_82_SUMB_33__51_), .CO(
        u5_mult_82_CARRYB_34__50_), .S(u5_mult_82_SUMB_34__50_) );
  FA_X1 u5_mult_82_S2_34_49 ( .A(u5_mult_82_ab_34__49_), .B(
        u5_mult_82_CARRYB_33__49_), .CI(u5_mult_82_SUMB_33__50_), .CO(
        u5_mult_82_CARRYB_34__49_), .S(u5_mult_82_SUMB_34__49_) );
  FA_X1 u5_mult_82_S2_34_48 ( .A(u5_mult_82_ab_34__48_), .B(
        u5_mult_82_CARRYB_33__48_), .CI(u5_mult_82_SUMB_33__49_), .CO(
        u5_mult_82_CARRYB_34__48_), .S(u5_mult_82_SUMB_34__48_) );
  FA_X1 u5_mult_82_S2_34_47 ( .A(u5_mult_82_CARRYB_33__47_), .B(
        u5_mult_82_ab_34__47_), .CI(u5_mult_82_SUMB_33__48_), .CO(
        u5_mult_82_CARRYB_34__47_), .S(u5_mult_82_SUMB_34__47_) );
  FA_X1 u5_mult_82_S2_34_46 ( .A(u5_mult_82_ab_34__46_), .B(
        u5_mult_82_CARRYB_33__46_), .CI(u5_mult_82_SUMB_33__47_), .CO(
        u5_mult_82_CARRYB_34__46_), .S(u5_mult_82_SUMB_34__46_) );
  FA_X1 u5_mult_82_S2_34_45 ( .A(u5_mult_82_CARRYB_33__45_), .B(
        u5_mult_82_ab_34__45_), .CI(u5_mult_82_SUMB_33__46_), .CO(
        u5_mult_82_CARRYB_34__45_), .S(u5_mult_82_SUMB_34__45_) );
  FA_X1 u5_mult_82_S2_34_39 ( .A(u5_mult_82_ab_34__39_), .B(
        u5_mult_82_CARRYB_33__39_), .CI(u5_mult_82_SUMB_33__40_), .CO(
        u5_mult_82_CARRYB_34__39_), .S(u5_mult_82_SUMB_34__39_) );
  FA_X1 u5_mult_82_S2_34_38 ( .A(u5_mult_82_ab_34__38_), .B(
        u5_mult_82_CARRYB_33__38_), .CI(u5_mult_82_SUMB_33__39_), .CO(
        u5_mult_82_CARRYB_34__38_), .S(u5_mult_82_SUMB_34__38_) );
  FA_X1 u5_mult_82_S2_34_37 ( .A(u5_mult_82_CARRYB_33__37_), .B(
        u5_mult_82_ab_34__37_), .CI(u5_mult_82_SUMB_33__38_), .CO(
        u5_mult_82_CARRYB_34__37_), .S(u5_mult_82_SUMB_34__37_) );
  FA_X1 u5_mult_82_S2_34_36 ( .A(u5_mult_82_ab_34__36_), .B(
        u5_mult_82_CARRYB_33__36_), .CI(u5_mult_82_SUMB_33__37_), .CO(
        u5_mult_82_CARRYB_34__36_), .S(u5_mult_82_SUMB_34__36_) );
  FA_X1 u5_mult_82_S2_34_35 ( .A(u5_mult_82_ab_34__35_), .B(
        u5_mult_82_CARRYB_33__35_), .CI(u5_mult_82_SUMB_33__36_), .CO(
        u5_mult_82_CARRYB_34__35_), .S(u5_mult_82_SUMB_34__35_) );
  FA_X1 u5_mult_82_S2_34_33 ( .A(u5_mult_82_CARRYB_33__33_), .B(
        u5_mult_82_ab_34__33_), .CI(u5_mult_82_SUMB_33__34_), .CO(
        u5_mult_82_CARRYB_34__33_), .S(u5_mult_82_SUMB_34__33_) );
  FA_X1 u5_mult_82_S2_34_28 ( .A(u5_mult_82_ab_34__28_), .B(
        u5_mult_82_CARRYB_33__28_), .CI(u5_mult_82_SUMB_33__29_), .CO(
        u5_mult_82_CARRYB_34__28_), .S(u5_mult_82_SUMB_34__28_) );
  FA_X1 u5_mult_82_S2_34_27 ( .A(u5_mult_82_CARRYB_33__27_), .B(
        u5_mult_82_ab_34__27_), .CI(u5_mult_82_SUMB_33__28_), .CO(
        u5_mult_82_CARRYB_34__27_), .S(u5_mult_82_SUMB_34__27_) );
  FA_X1 u5_mult_82_S2_34_26 ( .A(u5_mult_82_ab_34__26_), .B(
        u5_mult_82_CARRYB_33__26_), .CI(u5_mult_82_SUMB_33__27_), .CO(
        u5_mult_82_CARRYB_34__26_), .S(u5_mult_82_SUMB_34__26_) );
  FA_X1 u5_mult_82_S2_34_24 ( .A(u5_mult_82_ab_34__24_), .B(
        u5_mult_82_CARRYB_33__24_), .CI(u5_mult_82_SUMB_33__25_), .CO(
        u5_mult_82_CARRYB_34__24_), .S(u5_mult_82_SUMB_34__24_) );
  FA_X1 u5_mult_82_S2_34_23 ( .A(u5_mult_82_ab_34__23_), .B(
        u5_mult_82_CARRYB_33__23_), .CI(u5_mult_82_SUMB_33__24_), .CO(
        u5_mult_82_CARRYB_34__23_), .S(u5_mult_82_SUMB_34__23_) );
  FA_X1 u5_mult_82_S2_34_19 ( .A(u5_mult_82_ab_34__19_), .B(
        u5_mult_82_CARRYB_33__19_), .CI(u5_mult_82_SUMB_33__20_), .CO(
        u5_mult_82_CARRYB_34__19_), .S(u5_mult_82_SUMB_34__19_) );
  FA_X1 u5_mult_82_S2_34_3 ( .A(u5_mult_82_ab_34__3_), .B(
        u5_mult_82_CARRYB_33__3_), .CI(u5_mult_82_SUMB_33__4_), .CO(
        u5_mult_82_CARRYB_34__3_), .S(u5_mult_82_SUMB_34__3_) );
  FA_X1 u5_mult_82_S2_34_2 ( .A(u5_mult_82_ab_34__2_), .B(
        u5_mult_82_CARRYB_33__2_), .CI(u5_mult_82_SUMB_33__3_), .CO(
        u5_mult_82_CARRYB_34__2_), .S(u5_mult_82_SUMB_34__2_) );
  FA_X1 u5_mult_82_S2_34_1 ( .A(u5_mult_82_ab_34__1_), .B(
        u5_mult_82_CARRYB_33__1_), .CI(u5_mult_82_SUMB_33__2_), .CO(
        u5_mult_82_CARRYB_34__1_), .S(u5_mult_82_SUMB_34__1_) );
  FA_X1 u5_mult_82_S1_34_0 ( .A(u5_mult_82_ab_34__0_), .B(
        u5_mult_82_CARRYB_33__0_), .CI(u5_mult_82_SUMB_33__1_), .CO(
        u5_mult_82_CARRYB_34__0_), .S(u5_N34) );
  FA_X1 u5_mult_82_S3_35_51 ( .A(u5_mult_82_ab_35__51_), .B(
        u5_mult_82_CARRYB_34__51_), .CI(u5_mult_82_ab_34__52_), .CO(
        u5_mult_82_CARRYB_35__51_), .S(u5_mult_82_SUMB_35__51_) );
  FA_X1 u5_mult_82_S2_35_50 ( .A(u5_mult_82_ab_35__50_), .B(
        u5_mult_82_CARRYB_34__50_), .CI(u5_mult_82_SUMB_34__51_), .CO(
        u5_mult_82_CARRYB_35__50_), .S(u5_mult_82_SUMB_35__50_) );
  FA_X1 u5_mult_82_S2_35_49 ( .A(u5_mult_82_CARRYB_34__49_), .B(
        u5_mult_82_ab_35__49_), .CI(u5_mult_82_SUMB_34__50_), .CO(
        u5_mult_82_CARRYB_35__49_), .S(u5_mult_82_SUMB_35__49_) );
  FA_X1 u5_mult_82_S2_35_48 ( .A(u5_mult_82_ab_35__48_), .B(
        u5_mult_82_CARRYB_34__48_), .CI(u5_mult_82_SUMB_34__49_), .CO(
        u5_mult_82_CARRYB_35__48_), .S(u5_mult_82_SUMB_35__48_) );
  FA_X1 u5_mult_82_S2_35_47 ( .A(u5_mult_82_ab_35__47_), .B(
        u5_mult_82_CARRYB_34__47_), .CI(u5_mult_82_SUMB_34__48_), .CO(
        u5_mult_82_CARRYB_35__47_), .S(u5_mult_82_SUMB_35__47_) );
  FA_X1 u5_mult_82_S2_35_46 ( .A(u5_mult_82_ab_35__46_), .B(
        u5_mult_82_CARRYB_34__46_), .CI(u5_mult_82_SUMB_34__47_), .CO(
        u5_mult_82_CARRYB_35__46_), .S(u5_mult_82_SUMB_35__46_) );
  FA_X1 u5_mult_82_S2_35_44 ( .A(u5_mult_82_ab_35__44_), .B(
        u5_mult_82_CARRYB_34__44_), .CI(u5_mult_82_SUMB_34__45_), .CO(
        u5_mult_82_CARRYB_35__44_), .S(u5_mult_82_SUMB_35__44_) );
  FA_X1 u5_mult_82_S2_35_39 ( .A(u5_mult_82_ab_35__39_), .B(
        u5_mult_82_CARRYB_34__39_), .CI(u5_mult_82_SUMB_34__40_), .CO(
        u5_mult_82_CARRYB_35__39_), .S(u5_mult_82_SUMB_35__39_) );
  FA_X1 u5_mult_82_S2_35_38 ( .A(u5_mult_82_ab_35__38_), .B(
        u5_mult_82_CARRYB_34__38_), .CI(u5_mult_82_SUMB_34__39_), .CO(
        u5_mult_82_CARRYB_35__38_), .S(u5_mult_82_SUMB_35__38_) );
  FA_X1 u5_mult_82_S2_35_37 ( .A(u5_mult_82_ab_35__37_), .B(
        u5_mult_82_CARRYB_34__37_), .CI(u5_mult_82_SUMB_34__38_), .CO(
        u5_mult_82_CARRYB_35__37_), .S(u5_mult_82_SUMB_35__37_) );
  FA_X1 u5_mult_82_S2_35_24 ( .A(u5_mult_82_ab_35__24_), .B(
        u5_mult_82_CARRYB_34__24_), .CI(u5_mult_82_SUMB_34__25_), .CO(
        u5_mult_82_CARRYB_35__24_), .S(u5_mult_82_SUMB_35__24_) );
  FA_X1 u5_mult_82_S2_35_22 ( .A(u5_mult_82_ab_35__22_), .B(
        u5_mult_82_CARRYB_34__22_), .CI(u5_mult_82_SUMB_34__23_), .CO(
        u5_mult_82_CARRYB_35__22_), .S(u5_mult_82_SUMB_35__22_) );
  FA_X1 u5_mult_82_S2_35_18 ( .A(u5_mult_82_ab_35__18_), .B(
        u5_mult_82_CARRYB_34__18_), .CI(u5_mult_82_SUMB_34__19_), .CO(
        u5_mult_82_CARRYB_35__18_), .S(u5_mult_82_SUMB_35__18_) );
  FA_X1 u5_mult_82_S2_35_12 ( .A(u5_mult_82_CARRYB_34__12_), .B(
        u5_mult_82_ab_35__12_), .CI(u5_mult_82_SUMB_34__13_), .CO(
        u5_mult_82_CARRYB_35__12_), .S(u5_mult_82_SUMB_35__12_) );
  FA_X1 u5_mult_82_S2_35_10 ( .A(u5_mult_82_ab_35__10_), .B(
        u5_mult_82_CARRYB_34__10_), .CI(u5_mult_82_SUMB_34__11_), .CO(
        u5_mult_82_CARRYB_35__10_), .S(u5_mult_82_SUMB_35__10_) );
  FA_X1 u5_mult_82_S2_35_8 ( .A(u5_mult_82_CARRYB_34__8_), .B(
        u5_mult_82_ab_35__8_), .CI(u5_mult_82_SUMB_34__9_), .CO(
        u5_mult_82_CARRYB_35__8_), .S(u5_mult_82_SUMB_35__8_) );
  FA_X1 u5_mult_82_S2_35_7 ( .A(u5_mult_82_ab_35__7_), .B(
        u5_mult_82_CARRYB_34__7_), .CI(u5_mult_82_SUMB_34__8_), .CO(
        u5_mult_82_CARRYB_35__7_), .S(u5_mult_82_SUMB_35__7_) );
  FA_X1 u5_mult_82_S2_35_6 ( .A(u5_mult_82_SUMB_34__7_), .B(
        u5_mult_82_CARRYB_34__6_), .CI(u5_mult_82_ab_35__6_), .CO(
        u5_mult_82_CARRYB_35__6_), .S(u5_mult_82_SUMB_35__6_) );
  FA_X1 u5_mult_82_S2_35_5 ( .A(u5_mult_82_CARRYB_34__5_), .B(
        u5_mult_82_ab_35__5_), .CI(u5_mult_82_SUMB_34__6_), .CO(
        u5_mult_82_CARRYB_35__5_), .S(u5_mult_82_SUMB_35__5_) );
  FA_X1 u5_mult_82_S2_35_3 ( .A(u5_mult_82_ab_35__3_), .B(
        u5_mult_82_CARRYB_34__3_), .CI(u5_mult_82_SUMB_34__4_), .CO(
        u5_mult_82_CARRYB_35__3_), .S(u5_mult_82_SUMB_35__3_) );
  FA_X1 u5_mult_82_S2_35_2 ( .A(u5_mult_82_ab_35__2_), .B(
        u5_mult_82_SUMB_34__3_), .CI(u5_mult_82_CARRYB_34__2_), .CO(
        u5_mult_82_CARRYB_35__2_), .S(u5_mult_82_SUMB_35__2_) );
  FA_X1 u5_mult_82_S2_35_1 ( .A(u5_mult_82_ab_35__1_), .B(
        u5_mult_82_CARRYB_34__1_), .CI(u5_mult_82_SUMB_34__2_), .CO(
        u5_mult_82_CARRYB_35__1_), .S(u5_mult_82_SUMB_35__1_) );
  FA_X1 u5_mult_82_S1_35_0 ( .A(u5_mult_82_ab_35__0_), .B(
        u5_mult_82_CARRYB_34__0_), .CI(u5_mult_82_SUMB_34__1_), .CO(
        u5_mult_82_CARRYB_35__0_), .S(u5_N35) );
  FA_X1 u5_mult_82_S3_36_51 ( .A(u5_mult_82_ab_36__51_), .B(
        u5_mult_82_CARRYB_35__51_), .CI(u5_mult_82_ab_35__52_), .CO(
        u5_mult_82_CARRYB_36__51_), .S(u5_mult_82_SUMB_36__51_) );
  FA_X1 u5_mult_82_S2_36_50 ( .A(u5_mult_82_ab_36__50_), .B(
        u5_mult_82_CARRYB_35__50_), .CI(u5_mult_82_SUMB_35__51_), .CO(
        u5_mult_82_CARRYB_36__50_), .S(u5_mult_82_SUMB_36__50_) );
  FA_X1 u5_mult_82_S2_36_49 ( .A(u5_mult_82_ab_36__49_), .B(
        u5_mult_82_CARRYB_35__49_), .CI(u5_mult_82_SUMB_35__50_), .CO(
        u5_mult_82_CARRYB_36__49_), .S(u5_mult_82_SUMB_36__49_) );
  FA_X1 u5_mult_82_S2_36_48 ( .A(u5_mult_82_ab_36__48_), .B(
        u5_mult_82_CARRYB_35__48_), .CI(u5_mult_82_SUMB_35__49_), .CO(
        u5_mult_82_CARRYB_36__48_), .S(u5_mult_82_SUMB_36__48_) );
  FA_X1 u5_mult_82_S2_36_47 ( .A(u5_mult_82_ab_36__47_), .B(
        u5_mult_82_CARRYB_35__47_), .CI(u5_mult_82_SUMB_35__48_), .CO(
        u5_mult_82_CARRYB_36__47_), .S(u5_mult_82_SUMB_36__47_) );
  FA_X1 u5_mult_82_S2_36_46 ( .A(u5_mult_82_ab_36__46_), .B(
        u5_mult_82_CARRYB_35__46_), .CI(u5_mult_82_SUMB_35__47_), .CO(
        u5_mult_82_CARRYB_36__46_), .S(u5_mult_82_SUMB_36__46_) );
  FA_X1 u5_mult_82_S2_36_45 ( .A(u5_mult_82_ab_36__45_), .B(
        u5_mult_82_CARRYB_35__45_), .CI(u5_mult_82_SUMB_35__46_), .CO(
        u5_mult_82_CARRYB_36__45_), .S(u5_mult_82_SUMB_36__45_) );
  FA_X1 u5_mult_82_S2_36_43 ( .A(u5_mult_82_ab_36__43_), .B(
        u5_mult_82_CARRYB_35__43_), .CI(u5_mult_82_SUMB_35__44_), .CO(
        u5_mult_82_CARRYB_36__43_), .S(u5_mult_82_SUMB_36__43_) );
  FA_X1 u5_mult_82_S2_36_42 ( .A(u5_mult_82_ab_36__42_), .B(
        u5_mult_82_CARRYB_35__42_), .CI(u5_mult_82_SUMB_35__43_), .CO(
        u5_mult_82_CARRYB_36__42_), .S(u5_mult_82_SUMB_36__42_) );
  FA_X1 u5_mult_82_S2_36_41 ( .A(u5_mult_82_ab_36__41_), .B(
        u5_mult_82_CARRYB_35__41_), .CI(u5_mult_82_SUMB_35__42_), .CO(
        u5_mult_82_CARRYB_36__41_), .S(u5_mult_82_SUMB_36__41_) );
  FA_X1 u5_mult_82_S2_36_40 ( .A(u5_mult_82_ab_36__40_), .B(
        u5_mult_82_CARRYB_35__40_), .CI(u5_mult_82_SUMB_35__41_), .CO(
        u5_mult_82_CARRYB_36__40_), .S(u5_mult_82_SUMB_36__40_) );
  FA_X1 u5_mult_82_S2_36_39 ( .A(u5_mult_82_CARRYB_35__39_), .B(
        u5_mult_82_ab_36__39_), .CI(u5_mult_82_SUMB_35__40_), .CO(
        u5_mult_82_CARRYB_36__39_), .S(u5_mult_82_SUMB_36__39_) );
  FA_X1 u5_mult_82_S2_36_30 ( .A(u5_mult_82_ab_36__30_), .B(
        u5_mult_82_CARRYB_35__30_), .CI(u5_mult_82_SUMB_35__31_), .CO(
        u5_mult_82_CARRYB_36__30_), .S(u5_mult_82_SUMB_36__30_) );
  FA_X1 u5_mult_82_S2_36_28 ( .A(u5_mult_82_ab_36__28_), .B(
        u5_mult_82_CARRYB_35__28_), .CI(u5_mult_82_SUMB_35__29_), .CO(
        u5_mult_82_CARRYB_36__28_), .S(u5_mult_82_SUMB_36__28_) );
  FA_X1 u5_mult_82_S2_36_27 ( .A(u5_mult_82_CARRYB_35__27_), .B(
        u5_mult_82_ab_36__27_), .CI(u5_mult_82_SUMB_35__28_), .CO(
        u5_mult_82_CARRYB_36__27_), .S(u5_mult_82_SUMB_36__27_) );
  FA_X1 u5_mult_82_S2_36_19 ( .A(u5_mult_82_ab_36__19_), .B(
        u5_mult_82_CARRYB_35__19_), .CI(u5_mult_82_SUMB_35__20_), .CO(
        u5_mult_82_CARRYB_36__19_), .S(u5_mult_82_SUMB_36__19_) );
  FA_X1 u5_mult_82_S2_36_17 ( .A(u5_mult_82_ab_36__17_), .B(
        u5_mult_82_CARRYB_35__17_), .CI(u5_mult_82_SUMB_35__18_), .CO(
        u5_mult_82_CARRYB_36__17_), .S(u5_mult_82_SUMB_36__17_) );
  FA_X1 u5_mult_82_S2_36_12 ( .A(u5_mult_82_ab_36__12_), .B(
        u5_mult_82_CARRYB_35__12_), .CI(u5_mult_82_SUMB_35__13_), .CO(
        u5_mult_82_CARRYB_36__12_), .S(u5_mult_82_SUMB_36__12_) );
  FA_X1 u5_mult_82_S2_36_10 ( .A(u5_mult_82_ab_36__10_), .B(
        u5_mult_82_CARRYB_35__10_), .CI(u5_mult_82_SUMB_35__11_), .CO(
        u5_mult_82_CARRYB_36__10_), .S(u5_mult_82_SUMB_36__10_) );
  FA_X1 u5_mult_82_S2_36_9 ( .A(u5_mult_82_ab_36__9_), .B(
        u5_mult_82_CARRYB_35__9_), .CI(u5_mult_82_SUMB_35__10_), .CO(
        u5_mult_82_CARRYB_36__9_), .S(u5_mult_82_SUMB_36__9_) );
  FA_X1 u5_mult_82_S2_36_7 ( .A(u5_mult_82_ab_36__7_), .B(
        u5_mult_82_CARRYB_35__7_), .CI(u5_mult_82_SUMB_35__8_), .CO(
        u5_mult_82_CARRYB_36__7_), .S(u5_mult_82_SUMB_36__7_) );
  FA_X1 u5_mult_82_S2_36_6 ( .A(u5_mult_82_ab_36__6_), .B(
        u5_mult_82_CARRYB_35__6_), .CI(u5_mult_82_SUMB_35__7_), .CO(
        u5_mult_82_CARRYB_36__6_), .S(u5_mult_82_SUMB_36__6_) );
  FA_X1 u5_mult_82_S2_36_5 ( .A(u5_mult_82_SUMB_35__6_), .B(
        u5_mult_82_ab_36__5_), .CI(u5_mult_82_CARRYB_35__5_), .CO(
        u5_mult_82_CARRYB_36__5_), .S(u5_mult_82_SUMB_36__5_) );
  FA_X1 u5_mult_82_S2_36_4 ( .A(u5_mult_82_CARRYB_35__4_), .B(
        u5_mult_82_ab_36__4_), .CI(u5_mult_82_SUMB_35__5_), .CO(
        u5_mult_82_CARRYB_36__4_), .S(u5_mult_82_SUMB_36__4_) );
  FA_X1 u5_mult_82_S2_36_3 ( .A(u5_mult_82_ab_36__3_), .B(
        u5_mult_82_SUMB_35__4_), .CI(u5_mult_82_CARRYB_35__3_), .CO(
        u5_mult_82_CARRYB_36__3_), .S(u5_mult_82_SUMB_36__3_) );
  FA_X1 u5_mult_82_S2_36_1 ( .A(u5_mult_82_ab_36__1_), .B(
        u5_mult_82_CARRYB_35__1_), .CI(u5_mult_82_SUMB_35__2_), .CO(
        u5_mult_82_CARRYB_36__1_), .S(u5_mult_82_SUMB_36__1_) );
  FA_X1 u5_mult_82_S1_36_0 ( .A(u5_mult_82_CARRYB_35__0_), .B(
        u5_mult_82_ab_36__0_), .CI(u5_mult_82_SUMB_35__1_), .CO(
        u5_mult_82_CARRYB_36__0_), .S(u5_N36) );
  FA_X1 u5_mult_82_S3_37_51 ( .A(u5_mult_82_ab_37__51_), .B(
        u5_mult_82_CARRYB_36__51_), .CI(u5_mult_82_ab_36__52_), .CO(
        u5_mult_82_CARRYB_37__51_), .S(u5_mult_82_SUMB_37__51_) );
  FA_X1 u5_mult_82_S2_37_50 ( .A(u5_mult_82_ab_37__50_), .B(
        u5_mult_82_CARRYB_36__50_), .CI(u5_mult_82_SUMB_36__51_), .CO(
        u5_mult_82_CARRYB_37__50_), .S(u5_mult_82_SUMB_37__50_) );
  FA_X1 u5_mult_82_S2_37_49 ( .A(u5_mult_82_ab_37__49_), .B(
        u5_mult_82_CARRYB_36__49_), .CI(u5_mult_82_SUMB_36__50_), .CO(
        u5_mult_82_CARRYB_37__49_), .S(u5_mult_82_SUMB_37__49_) );
  FA_X1 u5_mult_82_S2_37_48 ( .A(u5_mult_82_ab_37__48_), .B(
        u5_mult_82_CARRYB_36__48_), .CI(u5_mult_82_SUMB_36__49_), .CO(
        u5_mult_82_CARRYB_37__48_), .S(u5_mult_82_SUMB_37__48_) );
  FA_X1 u5_mult_82_S2_37_47 ( .A(u5_mult_82_ab_37__47_), .B(
        u5_mult_82_CARRYB_36__47_), .CI(u5_mult_82_SUMB_36__48_), .CO(
        u5_mult_82_CARRYB_37__47_), .S(u5_mult_82_SUMB_37__47_) );
  FA_X1 u5_mult_82_S2_37_45 ( .A(u5_mult_82_ab_37__45_), .B(
        u5_mult_82_CARRYB_36__45_), .CI(u5_mult_82_SUMB_36__46_), .CO(
        u5_mult_82_CARRYB_37__45_), .S(u5_mult_82_SUMB_37__45_) );
  FA_X1 u5_mult_82_S2_37_44 ( .A(u5_mult_82_ab_37__44_), .B(
        u5_mult_82_CARRYB_36__44_), .CI(u5_mult_82_SUMB_36__45_), .CO(
        u5_mult_82_CARRYB_37__44_), .S(u5_mult_82_SUMB_37__44_) );
  FA_X1 u5_mult_82_S2_37_43 ( .A(u5_mult_82_ab_37__43_), .B(
        u5_mult_82_CARRYB_36__43_), .CI(u5_mult_82_SUMB_36__44_), .CO(
        u5_mult_82_CARRYB_37__43_), .S(u5_mult_82_SUMB_37__43_) );
  FA_X1 u5_mult_82_S2_37_42 ( .A(u5_mult_82_ab_37__42_), .B(
        u5_mult_82_CARRYB_36__42_), .CI(u5_mult_82_SUMB_36__43_), .CO(
        u5_mult_82_CARRYB_37__42_), .S(u5_mult_82_SUMB_37__42_) );
  FA_X1 u5_mult_82_S2_37_41 ( .A(u5_mult_82_ab_37__41_), .B(
        u5_mult_82_CARRYB_36__41_), .CI(u5_mult_82_SUMB_36__42_), .CO(
        u5_mult_82_CARRYB_37__41_), .S(u5_mult_82_SUMB_37__41_) );
  FA_X1 u5_mult_82_S2_37_39 ( .A(u5_mult_82_ab_37__39_), .B(
        u5_mult_82_CARRYB_36__39_), .CI(u5_mult_82_SUMB_36__40_), .CO(
        u5_mult_82_CARRYB_37__39_), .S(u5_mult_82_SUMB_37__39_) );
  FA_X1 u5_mult_82_S2_37_32 ( .A(u5_mult_82_ab_37__32_), .B(
        u5_mult_82_CARRYB_36__32_), .CI(u5_mult_82_SUMB_36__33_), .CO(
        u5_mult_82_CARRYB_37__32_), .S(u5_mult_82_SUMB_37__32_) );
  FA_X1 u5_mult_82_S2_37_30 ( .A(u5_mult_82_ab_37__30_), .B(
        u5_mult_82_CARRYB_36__30_), .CI(u5_mult_82_SUMB_36__31_), .CO(
        u5_mult_82_CARRYB_37__30_), .S(u5_mult_82_SUMB_37__30_) );
  FA_X1 u5_mult_82_S2_37_28 ( .A(u5_mult_82_ab_37__28_), .B(
        u5_mult_82_CARRYB_36__28_), .CI(u5_mult_82_SUMB_36__29_), .CO(
        u5_mult_82_CARRYB_37__28_), .S(u5_mult_82_SUMB_37__28_) );
  FA_X1 u5_mult_82_S2_37_27 ( .A(u5_mult_82_ab_37__27_), .B(
        u5_mult_82_CARRYB_36__27_), .CI(u5_mult_82_SUMB_36__28_), .CO(
        u5_mult_82_CARRYB_37__27_), .S(u5_mult_82_SUMB_37__27_) );
  FA_X1 u5_mult_82_S2_37_26 ( .A(u5_mult_82_ab_37__26_), .B(
        u5_mult_82_CARRYB_36__26_), .CI(u5_mult_82_SUMB_36__27_), .CO(
        u5_mult_82_CARRYB_37__26_), .S(u5_mult_82_SUMB_37__26_) );
  FA_X1 u5_mult_82_S2_37_25 ( .A(u5_mult_82_ab_37__25_), .B(
        u5_mult_82_CARRYB_36__25_), .CI(u5_mult_82_SUMB_36__26_), .CO(
        u5_mult_82_CARRYB_37__25_), .S(u5_mult_82_SUMB_37__25_) );
  FA_X1 u5_mult_82_S2_37_24 ( .A(u5_mult_82_ab_37__24_), .B(
        u5_mult_82_CARRYB_36__24_), .CI(u5_mult_82_SUMB_36__25_), .CO(
        u5_mult_82_CARRYB_37__24_), .S(u5_mult_82_SUMB_37__24_) );
  FA_X1 u5_mult_82_S2_37_22 ( .A(u5_mult_82_ab_37__22_), .B(
        u5_mult_82_CARRYB_36__22_), .CI(u5_mult_82_SUMB_36__23_), .CO(
        u5_mult_82_CARRYB_37__22_), .S(u5_mult_82_SUMB_37__22_) );
  FA_X1 u5_mult_82_S2_37_19 ( .A(u5_mult_82_ab_37__19_), .B(
        u5_mult_82_CARRYB_36__19_), .CI(u5_mult_82_SUMB_36__20_), .CO(
        u5_mult_82_CARRYB_37__19_), .S(u5_mult_82_SUMB_37__19_) );
  FA_X1 u5_mult_82_S2_37_12 ( .A(u5_mult_82_SUMB_36__13_), .B(
        u5_mult_82_ab_37__12_), .CI(u5_mult_82_CARRYB_36__12_), .CO(
        u5_mult_82_CARRYB_37__12_), .S(u5_mult_82_SUMB_37__12_) );
  FA_X1 u5_mult_82_S2_37_11 ( .A(u5_mult_82_ab_37__11_), .B(
        u5_mult_82_CARRYB_36__11_), .CI(u5_mult_82_SUMB_36__12_), .CO(
        u5_mult_82_CARRYB_37__11_), .S(u5_mult_82_SUMB_37__11_) );
  FA_X1 u5_mult_82_S2_37_8 ( .A(u5_mult_82_ab_37__8_), .B(
        u5_mult_82_CARRYB_36__8_), .CI(u5_mult_82_SUMB_36__9_), .CO(
        u5_mult_82_CARRYB_37__8_), .S(u5_mult_82_SUMB_37__8_) );
  FA_X1 u5_mult_82_S2_37_7 ( .A(u5_mult_82_SUMB_36__8_), .B(
        u5_mult_82_ab_37__7_), .CI(u5_mult_82_CARRYB_36__7_), .CO(
        u5_mult_82_CARRYB_37__7_), .S(u5_mult_82_SUMB_37__7_) );
  FA_X1 u5_mult_82_S2_37_2 ( .A(u5_mult_82_ab_37__2_), .B(
        u5_mult_82_CARRYB_36__2_), .CI(u5_mult_82_SUMB_36__3_), .CO(
        u5_mult_82_CARRYB_37__2_), .S(u5_mult_82_SUMB_37__2_) );
  FA_X1 u5_mult_82_S1_37_0 ( .A(u5_mult_82_ab_37__0_), .B(
        u5_mult_82_CARRYB_36__0_), .CI(u5_mult_82_SUMB_36__1_), .CO(
        u5_mult_82_CARRYB_37__0_), .S(u5_N37) );
  FA_X1 u5_mult_82_S3_38_51 ( .A(u5_mult_82_ab_38__51_), .B(
        u5_mult_82_CARRYB_37__51_), .CI(u5_mult_82_ab_37__52_), .CO(
        u5_mult_82_CARRYB_38__51_), .S(u5_mult_82_SUMB_38__51_) );
  FA_X1 u5_mult_82_S2_38_50 ( .A(u5_mult_82_ab_38__50_), .B(
        u5_mult_82_CARRYB_37__50_), .CI(u5_mult_82_SUMB_37__51_), .CO(
        u5_mult_82_CARRYB_38__50_), .S(u5_mult_82_SUMB_38__50_) );
  FA_X1 u5_mult_82_S2_38_49 ( .A(u5_mult_82_ab_38__49_), .B(
        u5_mult_82_CARRYB_37__49_), .CI(u5_mult_82_SUMB_37__50_), .CO(
        u5_mult_82_CARRYB_38__49_), .S(u5_mult_82_SUMB_38__49_) );
  FA_X1 u5_mult_82_S2_38_48 ( .A(u5_mult_82_ab_38__48_), .B(
        u5_mult_82_CARRYB_37__48_), .CI(u5_mult_82_SUMB_37__49_), .CO(
        u5_mult_82_CARRYB_38__48_), .S(u5_mult_82_SUMB_38__48_) );
  FA_X1 u5_mult_82_S2_38_47 ( .A(u5_mult_82_CARRYB_37__47_), .B(
        u5_mult_82_ab_38__47_), .CI(u5_mult_82_SUMB_37__48_), .CO(
        u5_mult_82_CARRYB_38__47_), .S(u5_mult_82_SUMB_38__47_) );
  FA_X1 u5_mult_82_S2_38_46 ( .A(u5_mult_82_ab_38__46_), .B(
        u5_mult_82_CARRYB_37__46_), .CI(u5_mult_82_SUMB_37__47_), .CO(
        u5_mult_82_CARRYB_38__46_), .S(u5_mult_82_SUMB_38__46_) );
  FA_X1 u5_mult_82_S2_38_45 ( .A(u5_mult_82_CARRYB_37__45_), .B(
        u5_mult_82_ab_38__45_), .CI(u5_mult_82_SUMB_37__46_), .CO(
        u5_mult_82_CARRYB_38__45_), .S(u5_mult_82_SUMB_38__45_) );
  FA_X1 u5_mult_82_S2_38_44 ( .A(u5_mult_82_CARRYB_37__44_), .B(
        u5_mult_82_ab_38__44_), .CI(u5_mult_82_SUMB_37__45_), .CO(
        u5_mult_82_CARRYB_38__44_), .S(u5_mult_82_SUMB_38__44_) );
  FA_X1 u5_mult_82_S2_38_43 ( .A(u5_mult_82_ab_38__43_), .B(
        u5_mult_82_CARRYB_37__43_), .CI(u5_mult_82_SUMB_37__44_), .CO(
        u5_mult_82_CARRYB_38__43_), .S(u5_mult_82_SUMB_38__43_) );
  FA_X1 u5_mult_82_S2_38_42 ( .A(u5_mult_82_ab_38__42_), .B(
        u5_mult_82_CARRYB_37__42_), .CI(u5_mult_82_SUMB_37__43_), .CO(
        u5_mult_82_CARRYB_38__42_), .S(u5_mult_82_SUMB_38__42_) );
  FA_X1 u5_mult_82_S2_38_41 ( .A(u5_mult_82_ab_38__41_), .B(
        u5_mult_82_CARRYB_37__41_), .CI(u5_mult_82_SUMB_37__42_), .CO(
        u5_mult_82_CARRYB_38__41_), .S(u5_mult_82_SUMB_38__41_) );
  FA_X1 u5_mult_82_S2_38_40 ( .A(u5_mult_82_ab_38__40_), .B(
        u5_mult_82_CARRYB_37__40_), .CI(u5_mult_82_SUMB_37__41_), .CO(
        u5_mult_82_CARRYB_38__40_), .S(u5_mult_82_SUMB_38__40_) );
  FA_X1 u5_mult_82_S2_38_36 ( .A(u5_mult_82_CARRYB_37__36_), .B(
        u5_mult_82_ab_38__36_), .CI(u5_mult_82_SUMB_37__37_), .CO(
        u5_mult_82_CARRYB_38__36_), .S(u5_mult_82_SUMB_38__36_) );
  FA_X1 u5_mult_82_S2_38_34 ( .A(u5_mult_82_ab_38__34_), .B(
        u5_mult_82_CARRYB_37__34_), .CI(u5_mult_82_SUMB_37__35_), .CO(
        u5_mult_82_CARRYB_38__34_), .S(u5_mult_82_SUMB_38__34_) );
  FA_X1 u5_mult_82_S2_38_27 ( .A(u5_mult_82_ab_38__27_), .B(
        u5_mult_82_CARRYB_37__27_), .CI(u5_mult_82_SUMB_37__28_), .CO(
        u5_mult_82_CARRYB_38__27_), .S(u5_mult_82_SUMB_38__27_) );
  FA_X1 u5_mult_82_S2_38_26 ( .A(u5_mult_82_CARRYB_37__26_), .B(
        u5_mult_82_ab_38__26_), .CI(u5_mult_82_SUMB_37__27_), .CO(
        u5_mult_82_CARRYB_38__26_), .S(u5_mult_82_SUMB_38__26_) );
  FA_X1 u5_mult_82_S2_38_25 ( .A(u5_mult_82_ab_38__25_), .B(
        u5_mult_82_CARRYB_37__25_), .CI(u5_mult_82_SUMB_37__26_), .CO(
        u5_mult_82_CARRYB_38__25_), .S(u5_mult_82_SUMB_38__25_) );
  FA_X1 u5_mult_82_S2_38_19 ( .A(u5_mult_82_ab_38__19_), .B(
        u5_mult_82_CARRYB_37__19_), .CI(u5_mult_82_SUMB_37__20_), .CO(
        u5_mult_82_CARRYB_38__19_), .S(u5_mult_82_SUMB_38__19_) );
  FA_X1 u5_mult_82_S2_38_11 ( .A(u5_mult_82_CARRYB_37__11_), .B(
        u5_mult_82_ab_38__11_), .CI(u5_mult_82_SUMB_37__12_), .CO(
        u5_mult_82_CARRYB_38__11_), .S(u5_mult_82_SUMB_38__11_) );
  FA_X1 u5_mult_82_S2_38_6 ( .A(u5_mult_82_ab_38__6_), .B(
        u5_mult_82_CARRYB_37__6_), .CI(u5_mult_82_SUMB_37__7_), .CO(
        u5_mult_82_CARRYB_38__6_), .S(u5_mult_82_SUMB_38__6_) );
  FA_X1 u5_mult_82_S2_38_4 ( .A(u5_mult_82_CARRYB_37__4_), .B(
        u5_mult_82_ab_38__4_), .CI(u5_mult_82_SUMB_37__5_), .CO(
        u5_mult_82_CARRYB_38__4_), .S(u5_mult_82_SUMB_38__4_) );
  FA_X1 u5_mult_82_S1_38_0 ( .A(u5_mult_82_CARRYB_37__0_), .B(
        u5_mult_82_ab_38__0_), .CI(u5_mult_82_SUMB_37__1_), .CO(
        u5_mult_82_CARRYB_38__0_), .S(u5_N38) );
  FA_X1 u5_mult_82_S3_39_51 ( .A(u5_mult_82_ab_39__51_), .B(
        u5_mult_82_CARRYB_38__51_), .CI(u5_mult_82_ab_38__52_), .CO(
        u5_mult_82_CARRYB_39__51_), .S(u5_mult_82_SUMB_39__51_) );
  FA_X1 u5_mult_82_S2_39_50 ( .A(u5_mult_82_ab_39__50_), .B(
        u5_mult_82_CARRYB_38__50_), .CI(u5_mult_82_SUMB_38__51_), .CO(
        u5_mult_82_CARRYB_39__50_), .S(u5_mult_82_SUMB_39__50_) );
  FA_X1 u5_mult_82_S2_39_49 ( .A(u5_mult_82_ab_39__49_), .B(
        u5_mult_82_CARRYB_38__49_), .CI(u5_mult_82_SUMB_38__50_), .CO(
        u5_mult_82_CARRYB_39__49_), .S(u5_mult_82_SUMB_39__49_) );
  FA_X1 u5_mult_82_S2_39_48 ( .A(u5_mult_82_ab_39__48_), .B(
        u5_mult_82_CARRYB_38__48_), .CI(u5_mult_82_SUMB_38__49_), .CO(
        u5_mult_82_CARRYB_39__48_), .S(u5_mult_82_SUMB_39__48_) );
  FA_X1 u5_mult_82_S2_39_47 ( .A(u5_mult_82_ab_39__47_), .B(
        u5_mult_82_CARRYB_38__47_), .CI(u5_mult_82_SUMB_38__48_), .CO(
        u5_mult_82_CARRYB_39__47_), .S(u5_mult_82_SUMB_39__47_) );
  FA_X1 u5_mult_82_S2_39_46 ( .A(u5_mult_82_ab_39__46_), .B(
        u5_mult_82_CARRYB_38__46_), .CI(u5_mult_82_SUMB_38__47_), .CO(
        u5_mult_82_CARRYB_39__46_), .S(u5_mult_82_SUMB_39__46_) );
  FA_X1 u5_mult_82_S2_39_45 ( .A(u5_mult_82_ab_39__45_), .B(
        u5_mult_82_CARRYB_38__45_), .CI(u5_mult_82_SUMB_38__46_), .CO(
        u5_mult_82_CARRYB_39__45_), .S(u5_mult_82_SUMB_39__45_) );
  FA_X1 u5_mult_82_S2_39_44 ( .A(u5_mult_82_ab_39__44_), .B(
        u5_mult_82_CARRYB_38__44_), .CI(u5_mult_82_SUMB_38__45_), .CO(
        u5_mult_82_CARRYB_39__44_), .S(u5_mult_82_SUMB_39__44_) );
  FA_X1 u5_mult_82_S2_39_43 ( .A(u5_mult_82_ab_39__43_), .B(
        u5_mult_82_CARRYB_38__43_), .CI(u5_mult_82_SUMB_38__44_), .CO(
        u5_mult_82_CARRYB_39__43_), .S(u5_mult_82_SUMB_39__43_) );
  FA_X1 u5_mult_82_S2_39_42 ( .A(u5_mult_82_ab_39__42_), .B(
        u5_mult_82_CARRYB_38__42_), .CI(u5_mult_82_SUMB_38__43_), .CO(
        u5_mult_82_CARRYB_39__42_), .S(u5_mult_82_SUMB_39__42_) );
  FA_X1 u5_mult_82_S2_39_41 ( .A(u5_mult_82_ab_39__41_), .B(
        u5_mult_82_CARRYB_38__41_), .CI(u5_mult_82_SUMB_38__42_), .CO(
        u5_mult_82_CARRYB_39__41_), .S(u5_mult_82_SUMB_39__41_) );
  FA_X1 u5_mult_82_S2_39_40 ( .A(u5_mult_82_ab_39__40_), .B(
        u5_mult_82_CARRYB_38__40_), .CI(u5_mult_82_SUMB_38__41_), .CO(
        u5_mult_82_CARRYB_39__40_), .S(u5_mult_82_SUMB_39__40_) );
  FA_X1 u5_mult_82_S2_39_32 ( .A(u5_mult_82_CARRYB_38__32_), .B(
        u5_mult_82_ab_39__32_), .CI(u5_mult_82_SUMB_38__33_), .CO(
        u5_mult_82_CARRYB_39__32_), .S(u5_mult_82_SUMB_39__32_) );
  FA_X1 u5_mult_82_S2_39_27 ( .A(u5_mult_82_CARRYB_38__27_), .B(
        u5_mult_82_ab_39__27_), .CI(u5_mult_82_SUMB_38__28_), .CO(
        u5_mult_82_CARRYB_39__27_), .S(u5_mult_82_SUMB_39__27_) );
  FA_X1 u5_mult_82_S2_39_23 ( .A(u5_mult_82_ab_39__23_), .B(
        u5_mult_82_CARRYB_38__23_), .CI(u5_mult_82_SUMB_38__24_), .CO(
        u5_mult_82_CARRYB_39__23_), .S(u5_mult_82_SUMB_39__23_) );
  FA_X1 u5_mult_82_S2_39_21 ( .A(u5_mult_82_ab_39__21_), .B(
        u5_mult_82_CARRYB_38__21_), .CI(u5_mult_82_SUMB_38__22_), .CO(
        u5_mult_82_CARRYB_39__21_), .S(u5_mult_82_SUMB_39__21_) );
  FA_X1 u5_mult_82_S2_39_4 ( .A(u5_mult_82_ab_39__4_), .B(
        u5_mult_82_CARRYB_38__4_), .CI(u5_mult_82_SUMB_38__5_), .CO(
        u5_mult_82_CARRYB_39__4_), .S(u5_mult_82_SUMB_39__4_) );
  FA_X1 u5_mult_82_S2_39_3 ( .A(u5_mult_82_ab_39__3_), .B(
        u5_mult_82_CARRYB_38__3_), .CI(u5_mult_82_SUMB_38__4_), .CO(
        u5_mult_82_CARRYB_39__3_), .S(u5_mult_82_SUMB_39__3_) );
  FA_X1 u5_mult_82_S3_40_51 ( .A(u5_mult_82_ab_40__51_), .B(
        u5_mult_82_CARRYB_39__51_), .CI(u5_mult_82_ab_39__52_), .CO(
        u5_mult_82_CARRYB_40__51_), .S(u5_mult_82_SUMB_40__51_) );
  FA_X1 u5_mult_82_S2_40_50 ( .A(u5_mult_82_ab_40__50_), .B(
        u5_mult_82_CARRYB_39__50_), .CI(u5_mult_82_SUMB_39__51_), .CO(
        u5_mult_82_CARRYB_40__50_), .S(u5_mult_82_SUMB_40__50_) );
  FA_X1 u5_mult_82_S2_40_49 ( .A(u5_mult_82_ab_40__49_), .B(
        u5_mult_82_CARRYB_39__49_), .CI(u5_mult_82_SUMB_39__50_), .CO(
        u5_mult_82_CARRYB_40__49_), .S(u5_mult_82_SUMB_40__49_) );
  FA_X1 u5_mult_82_S2_40_48 ( .A(u5_mult_82_ab_40__48_), .B(
        u5_mult_82_CARRYB_39__48_), .CI(u5_mult_82_SUMB_39__49_), .CO(
        u5_mult_82_CARRYB_40__48_), .S(u5_mult_82_SUMB_40__48_) );
  FA_X1 u5_mult_82_S2_40_47 ( .A(u5_mult_82_ab_40__47_), .B(
        u5_mult_82_CARRYB_39__47_), .CI(u5_mult_82_SUMB_39__48_), .CO(
        u5_mult_82_CARRYB_40__47_), .S(u5_mult_82_SUMB_40__47_) );
  FA_X1 u5_mult_82_S2_40_46 ( .A(u5_mult_82_ab_40__46_), .B(
        u5_mult_82_CARRYB_39__46_), .CI(u5_mult_82_SUMB_39__47_), .CO(
        u5_mult_82_CARRYB_40__46_), .S(u5_mult_82_SUMB_40__46_) );
  FA_X1 u5_mult_82_S2_40_45 ( .A(u5_mult_82_ab_40__45_), .B(
        u5_mult_82_CARRYB_39__45_), .CI(u5_mult_82_SUMB_39__46_), .CO(
        u5_mult_82_CARRYB_40__45_), .S(u5_mult_82_SUMB_40__45_) );
  FA_X1 u5_mult_82_S2_40_44 ( .A(u5_mult_82_ab_40__44_), .B(
        u5_mult_82_CARRYB_39__44_), .CI(u5_mult_82_SUMB_39__45_), .CO(
        u5_mult_82_CARRYB_40__44_), .S(u5_mult_82_SUMB_40__44_) );
  FA_X1 u5_mult_82_S2_40_43 ( .A(u5_mult_82_ab_40__43_), .B(
        u5_mult_82_CARRYB_39__43_), .CI(u5_mult_82_SUMB_39__44_), .CO(
        u5_mult_82_CARRYB_40__43_), .S(u5_mult_82_SUMB_40__43_) );
  FA_X1 u5_mult_82_S2_40_42 ( .A(u5_mult_82_ab_40__42_), .B(
        u5_mult_82_CARRYB_39__42_), .CI(u5_mult_82_SUMB_39__43_), .CO(
        u5_mult_82_CARRYB_40__42_), .S(u5_mult_82_SUMB_40__42_) );
  FA_X1 u5_mult_82_S2_40_41 ( .A(u5_mult_82_ab_40__41_), .B(
        u5_mult_82_CARRYB_39__41_), .CI(u5_mult_82_SUMB_39__42_), .CO(
        u5_mult_82_CARRYB_40__41_), .S(u5_mult_82_SUMB_40__41_) );
  FA_X1 u5_mult_82_S2_40_36 ( .A(u5_mult_82_ab_40__36_), .B(
        u5_mult_82_CARRYB_39__36_), .CI(u5_mult_82_SUMB_39__37_), .CO(
        u5_mult_82_CARRYB_40__36_), .S(u5_mult_82_SUMB_40__36_) );
  FA_X1 u5_mult_82_S2_40_33 ( .A(u5_mult_82_ab_40__33_), .B(
        u5_mult_82_CARRYB_39__33_), .CI(u5_mult_82_SUMB_39__34_), .CO(
        u5_mult_82_CARRYB_40__33_), .S(u5_mult_82_SUMB_40__33_) );
  FA_X1 u5_mult_82_S2_40_28 ( .A(u5_mult_82_ab_40__28_), .B(
        u5_mult_82_CARRYB_39__28_), .CI(u5_mult_82_SUMB_39__29_), .CO(
        u5_mult_82_CARRYB_40__28_), .S(u5_mult_82_SUMB_40__28_) );
  FA_X1 u5_mult_82_S2_40_26 ( .A(u5_mult_82_CARRYB_39__26_), .B(
        u5_mult_82_ab_40__26_), .CI(u5_mult_82_SUMB_39__27_), .CO(
        u5_mult_82_CARRYB_40__26_), .S(u5_mult_82_SUMB_40__26_) );
  FA_X1 u5_mult_82_S2_40_18 ( .A(u5_mult_82_ab_40__18_), .B(
        u5_mult_82_CARRYB_39__18_), .CI(u5_mult_82_SUMB_39__19_), .CO(
        u5_mult_82_CARRYB_40__18_), .S(u5_mult_82_SUMB_40__18_) );
  FA_X1 u5_mult_82_S2_40_10 ( .A(u5_mult_82_ab_40__10_), .B(
        u5_mult_82_CARRYB_39__10_), .CI(u5_mult_82_SUMB_39__11_), .CO(
        u5_mult_82_CARRYB_40__10_), .S(u5_mult_82_SUMB_40__10_) );
  FA_X1 u5_mult_82_S2_40_8 ( .A(u5_mult_82_ab_40__8_), .B(
        u5_mult_82_CARRYB_39__8_), .CI(u5_mult_82_SUMB_39__9_), .CO(
        u5_mult_82_CARRYB_40__8_), .S(u5_mult_82_SUMB_40__8_) );
  FA_X1 u5_mult_82_S2_40_7 ( .A(u5_mult_82_ab_40__7_), .B(
        u5_mult_82_CARRYB_39__7_), .CI(u5_mult_82_SUMB_39__8_), .CO(
        u5_mult_82_CARRYB_40__7_), .S(u5_mult_82_SUMB_40__7_) );
  FA_X1 u5_mult_82_S2_40_4 ( .A(u5_mult_82_CARRYB_39__4_), .B(
        u5_mult_82_ab_40__4_), .CI(u5_mult_82_SUMB_39__5_), .CO(
        u5_mult_82_CARRYB_40__4_), .S(u5_mult_82_SUMB_40__4_) );
  FA_X1 u5_mult_82_S2_40_2 ( .A(u5_mult_82_CARRYB_39__2_), .B(
        u5_mult_82_ab_40__2_), .CI(u5_mult_82_SUMB_39__3_), .CO(
        u5_mult_82_CARRYB_40__2_), .S(u5_mult_82_SUMB_40__2_) );
  FA_X1 u5_mult_82_S2_40_1 ( .A(u5_mult_82_SUMB_39__2_), .B(
        u5_mult_82_ab_40__1_), .CI(u5_mult_82_CARRYB_39__1_), .CO(
        u5_mult_82_CARRYB_40__1_), .S(u5_mult_82_SUMB_40__1_) );
  FA_X1 u5_mult_82_S3_41_51 ( .A(u5_mult_82_ab_41__51_), .B(
        u5_mult_82_CARRYB_40__51_), .CI(u5_mult_82_ab_40__52_), .CO(
        u5_mult_82_CARRYB_41__51_), .S(u5_mult_82_SUMB_41__51_) );
  FA_X1 u5_mult_82_S2_41_50 ( .A(u5_mult_82_ab_41__50_), .B(
        u5_mult_82_CARRYB_40__50_), .CI(u5_mult_82_SUMB_40__51_), .CO(
        u5_mult_82_CARRYB_41__50_), .S(u5_mult_82_SUMB_41__50_) );
  FA_X1 u5_mult_82_S2_41_49 ( .A(u5_mult_82_ab_41__49_), .B(
        u5_mult_82_CARRYB_40__49_), .CI(u5_mult_82_SUMB_40__50_), .CO(
        u5_mult_82_CARRYB_41__49_), .S(u5_mult_82_SUMB_41__49_) );
  FA_X1 u5_mult_82_S2_41_48 ( .A(u5_mult_82_ab_41__48_), .B(
        u5_mult_82_CARRYB_40__48_), .CI(u5_mult_82_SUMB_40__49_), .CO(
        u5_mult_82_CARRYB_41__48_), .S(u5_mult_82_SUMB_41__48_) );
  FA_X1 u5_mult_82_S2_41_47 ( .A(u5_mult_82_ab_41__47_), .B(
        u5_mult_82_CARRYB_40__47_), .CI(u5_mult_82_SUMB_40__48_), .CO(
        u5_mult_82_CARRYB_41__47_), .S(u5_mult_82_SUMB_41__47_) );
  FA_X1 u5_mult_82_S2_41_46 ( .A(u5_mult_82_ab_41__46_), .B(
        u5_mult_82_CARRYB_40__46_), .CI(u5_mult_82_SUMB_40__47_), .CO(
        u5_mult_82_CARRYB_41__46_), .S(u5_mult_82_SUMB_41__46_) );
  FA_X1 u5_mult_82_S2_41_45 ( .A(u5_mult_82_CARRYB_40__45_), .B(
        u5_mult_82_ab_41__45_), .CI(u5_mult_82_SUMB_40__46_), .CO(
        u5_mult_82_CARRYB_41__45_), .S(u5_mult_82_SUMB_41__45_) );
  FA_X1 u5_mult_82_S2_41_44 ( .A(u5_mult_82_ab_41__44_), .B(
        u5_mult_82_CARRYB_40__44_), .CI(u5_mult_82_SUMB_40__45_), .CO(
        u5_mult_82_CARRYB_41__44_), .S(u5_mult_82_SUMB_41__44_) );
  FA_X1 u5_mult_82_S2_41_43 ( .A(u5_mult_82_CARRYB_40__43_), .B(
        u5_mult_82_ab_41__43_), .CI(u5_mult_82_SUMB_40__44_), .CO(
        u5_mult_82_CARRYB_41__43_), .S(u5_mult_82_SUMB_41__43_) );
  FA_X1 u5_mult_82_S2_41_42 ( .A(u5_mult_82_CARRYB_40__42_), .B(
        u5_mult_82_ab_41__42_), .CI(u5_mult_82_SUMB_40__43_), .CO(
        u5_mult_82_CARRYB_41__42_), .S(u5_mult_82_SUMB_41__42_) );
  FA_X1 u5_mult_82_S2_41_41 ( .A(u5_mult_82_ab_41__41_), .B(
        u5_mult_82_CARRYB_40__41_), .CI(u5_mult_82_SUMB_40__42_), .CO(
        u5_mult_82_CARRYB_41__41_), .S(u5_mult_82_SUMB_41__41_) );
  FA_X1 u5_mult_82_S2_41_40 ( .A(u5_mult_82_ab_41__40_), .B(
        u5_mult_82_CARRYB_40__40_), .CI(u5_mult_82_SUMB_40__41_), .CO(
        u5_mult_82_CARRYB_41__40_), .S(u5_mult_82_SUMB_41__40_) );
  FA_X1 u5_mult_82_S2_41_38 ( .A(u5_mult_82_ab_41__38_), .B(
        u5_mult_82_CARRYB_40__38_), .CI(u5_mult_82_SUMB_40__39_), .CO(
        u5_mult_82_CARRYB_41__38_), .S(u5_mult_82_SUMB_41__38_) );
  FA_X1 u5_mult_82_S2_41_35 ( .A(u5_mult_82_ab_41__35_), .B(
        u5_mult_82_CARRYB_40__35_), .CI(u5_mult_82_SUMB_40__36_), .CO(
        u5_mult_82_CARRYB_41__35_), .S(u5_mult_82_SUMB_41__35_) );
  FA_X1 u5_mult_82_S2_41_33 ( .A(u5_mult_82_ab_41__33_), .B(
        u5_mult_82_CARRYB_40__33_), .CI(u5_mult_82_SUMB_40__34_), .CO(
        u5_mult_82_CARRYB_41__33_), .S(u5_mult_82_SUMB_41__33_) );
  FA_X1 u5_mult_82_S2_41_29 ( .A(u5_mult_82_ab_41__29_), .B(
        u5_mult_82_CARRYB_40__29_), .CI(u5_mult_82_SUMB_40__30_), .CO(
        u5_mult_82_CARRYB_41__29_), .S(u5_mult_82_SUMB_41__29_) );
  FA_X1 u5_mult_82_S2_41_24 ( .A(u5_mult_82_ab_41__24_), .B(
        u5_mult_82_CARRYB_40__24_), .CI(u5_mult_82_SUMB_40__25_), .CO(
        u5_mult_82_CARRYB_41__24_), .S(u5_mult_82_SUMB_41__24_) );
  FA_X1 u5_mult_82_S2_41_20 ( .A(u5_mult_82_ab_41__20_), .B(
        u5_mult_82_CARRYB_40__20_), .CI(u5_mult_82_SUMB_40__21_), .CO(
        u5_mult_82_CARRYB_41__20_), .S(u5_mult_82_SUMB_41__20_) );
  FA_X1 u5_mult_82_S3_42_51 ( .A(u5_mult_82_ab_42__51_), .B(
        u5_mult_82_CARRYB_41__51_), .CI(u5_mult_82_ab_41__52_), .CO(
        u5_mult_82_CARRYB_42__51_), .S(u5_mult_82_SUMB_42__51_) );
  FA_X1 u5_mult_82_S2_42_50 ( .A(u5_mult_82_ab_42__50_), .B(
        u5_mult_82_CARRYB_41__50_), .CI(u5_mult_82_SUMB_41__51_), .CO(
        u5_mult_82_CARRYB_42__50_), .S(u5_mult_82_SUMB_42__50_) );
  FA_X1 u5_mult_82_S2_42_49 ( .A(u5_mult_82_ab_42__49_), .B(
        u5_mult_82_CARRYB_41__49_), .CI(u5_mult_82_SUMB_41__50_), .CO(
        u5_mult_82_CARRYB_42__49_), .S(u5_mult_82_SUMB_42__49_) );
  FA_X1 u5_mult_82_S2_42_48 ( .A(u5_mult_82_ab_42__48_), .B(
        u5_mult_82_CARRYB_41__48_), .CI(u5_mult_82_SUMB_41__49_), .CO(
        u5_mult_82_CARRYB_42__48_), .S(u5_mult_82_SUMB_42__48_) );
  FA_X1 u5_mult_82_S2_42_47 ( .A(u5_mult_82_ab_42__47_), .B(
        u5_mult_82_CARRYB_41__47_), .CI(u5_mult_82_SUMB_41__48_), .CO(
        u5_mult_82_CARRYB_42__47_), .S(u5_mult_82_SUMB_42__47_) );
  FA_X1 u5_mult_82_S2_42_46 ( .A(u5_mult_82_ab_42__46_), .B(
        u5_mult_82_CARRYB_41__46_), .CI(u5_mult_82_SUMB_41__47_), .CO(
        u5_mult_82_CARRYB_42__46_), .S(u5_mult_82_SUMB_42__46_) );
  FA_X1 u5_mult_82_S2_42_45 ( .A(u5_mult_82_ab_42__45_), .B(
        u5_mult_82_CARRYB_41__45_), .CI(u5_mult_82_SUMB_41__46_), .CO(
        u5_mult_82_CARRYB_42__45_), .S(u5_mult_82_SUMB_42__45_) );
  FA_X1 u5_mult_82_S2_42_44 ( .A(u5_mult_82_ab_42__44_), .B(
        u5_mult_82_CARRYB_41__44_), .CI(u5_mult_82_SUMB_41__45_), .CO(
        u5_mult_82_CARRYB_42__44_), .S(u5_mult_82_SUMB_42__44_) );
  FA_X1 u5_mult_82_S2_42_43 ( .A(u5_mult_82_CARRYB_41__43_), .B(
        u5_mult_82_ab_42__43_), .CI(u5_mult_82_SUMB_41__44_), .CO(
        u5_mult_82_CARRYB_42__43_), .S(u5_mult_82_SUMB_42__43_) );
  FA_X1 u5_mult_82_S2_42_42 ( .A(u5_mult_82_CARRYB_41__42_), .B(
        u5_mult_82_ab_42__42_), .CI(u5_mult_82_SUMB_41__43_), .CO(
        u5_mult_82_CARRYB_42__42_), .S(u5_mult_82_SUMB_42__42_) );
  FA_X1 u5_mult_82_S2_42_40 ( .A(u5_mult_82_ab_42__40_), .B(
        u5_mult_82_CARRYB_41__40_), .CI(u5_mult_82_SUMB_41__41_), .CO(
        u5_mult_82_CARRYB_42__40_), .S(u5_mult_82_SUMB_42__40_) );
  FA_X1 u5_mult_82_S2_42_39 ( .A(u5_mult_82_ab_42__39_), .B(
        u5_mult_82_CARRYB_41__39_), .CI(u5_mult_82_SUMB_41__40_), .CO(
        u5_mult_82_CARRYB_42__39_), .S(u5_mult_82_SUMB_42__39_) );
  FA_X1 u5_mult_82_S2_42_38 ( .A(u5_mult_82_ab_42__38_), .B(
        u5_mult_82_CARRYB_41__38_), .CI(u5_mult_82_SUMB_41__39_), .CO(
        u5_mult_82_CARRYB_42__38_), .S(u5_mult_82_SUMB_42__38_) );
  FA_X1 u5_mult_82_S2_42_37 ( .A(u5_mult_82_ab_42__37_), .B(
        u5_mult_82_CARRYB_41__37_), .CI(u5_mult_82_SUMB_41__38_), .CO(
        u5_mult_82_CARRYB_42__37_), .S(u5_mult_82_SUMB_42__37_) );
  FA_X1 u5_mult_82_S2_42_36 ( .A(u5_mult_82_ab_42__36_), .B(
        u5_mult_82_CARRYB_41__36_), .CI(u5_mult_82_SUMB_41__37_), .CO(
        u5_mult_82_CARRYB_42__36_), .S(u5_mult_82_SUMB_42__36_) );
  FA_X1 u5_mult_82_S2_42_35 ( .A(u5_mult_82_CARRYB_41__35_), .B(
        u5_mult_82_ab_42__35_), .CI(u5_mult_82_SUMB_41__36_), .CO(
        u5_mult_82_CARRYB_42__35_), .S(u5_mult_82_SUMB_42__35_) );
  FA_X1 u5_mult_82_S2_42_28 ( .A(u5_mult_82_ab_42__28_), .B(
        u5_mult_82_CARRYB_41__28_), .CI(u5_mult_82_SUMB_41__29_), .CO(
        u5_mult_82_CARRYB_42__28_), .S(u5_mult_82_SUMB_42__28_) );
  FA_X1 u5_mult_82_S2_42_25 ( .A(u5_mult_82_ab_42__25_), .B(
        u5_mult_82_CARRYB_41__25_), .CI(u5_mult_82_SUMB_41__26_), .CO(
        u5_mult_82_CARRYB_42__25_), .S(u5_mult_82_SUMB_42__25_) );
  FA_X1 u5_mult_82_S2_42_22 ( .A(u5_mult_82_ab_42__22_), .B(
        u5_mult_82_CARRYB_41__22_), .CI(u5_mult_82_SUMB_41__23_), .CO(
        u5_mult_82_CARRYB_42__22_), .S(u5_mult_82_SUMB_42__22_) );
  FA_X1 u5_mult_82_S2_42_16 ( .A(u5_mult_82_ab_42__16_), .B(
        u5_mult_82_CARRYB_41__16_), .CI(u5_mult_82_SUMB_41__17_), .CO(
        u5_mult_82_CARRYB_42__16_), .S(u5_mult_82_SUMB_42__16_) );
  FA_X1 u5_mult_82_S2_42_5 ( .A(u5_mult_82_CARRYB_41__5_), .B(
        u5_mult_82_ab_42__5_), .CI(u5_mult_82_SUMB_41__6_), .CO(
        u5_mult_82_CARRYB_42__5_), .S(u5_mult_82_SUMB_42__5_) );
  FA_X1 u5_mult_82_S2_42_1 ( .A(u5_mult_82_ab_42__1_), .B(
        u5_mult_82_CARRYB_41__1_), .CI(u5_mult_82_n49), .CO(
        u5_mult_82_CARRYB_42__1_), .S(u5_mult_82_SUMB_42__1_) );
  FA_X1 u5_mult_82_S1_42_0 ( .A(u5_mult_82_ab_42__0_), .B(
        u5_mult_82_CARRYB_41__0_), .CI(u5_mult_82_SUMB_41__1_), .CO(
        u5_mult_82_CARRYB_42__0_), .S(u5_N42) );
  FA_X1 u5_mult_82_S3_43_51 ( .A(u5_mult_82_ab_43__51_), .B(
        u5_mult_82_CARRYB_42__51_), .CI(u5_mult_82_ab_42__52_), .CO(
        u5_mult_82_CARRYB_43__51_), .S(u5_mult_82_SUMB_43__51_) );
  FA_X1 u5_mult_82_S2_43_50 ( .A(u5_mult_82_ab_43__50_), .B(
        u5_mult_82_CARRYB_42__50_), .CI(u5_mult_82_SUMB_42__51_), .CO(
        u5_mult_82_CARRYB_43__50_), .S(u5_mult_82_SUMB_43__50_) );
  FA_X1 u5_mult_82_S2_43_49 ( .A(u5_mult_82_ab_43__49_), .B(
        u5_mult_82_CARRYB_42__49_), .CI(u5_mult_82_SUMB_42__50_), .CO(
        u5_mult_82_CARRYB_43__49_), .S(u5_mult_82_SUMB_43__49_) );
  FA_X1 u5_mult_82_S2_43_48 ( .A(u5_mult_82_ab_43__48_), .B(
        u5_mult_82_CARRYB_42__48_), .CI(u5_mult_82_SUMB_42__49_), .CO(
        u5_mult_82_CARRYB_43__48_), .S(u5_mult_82_SUMB_43__48_) );
  FA_X1 u5_mult_82_S2_43_47 ( .A(u5_mult_82_ab_43__47_), .B(
        u5_mult_82_CARRYB_42__47_), .CI(u5_mult_82_SUMB_42__48_), .CO(
        u5_mult_82_CARRYB_43__47_), .S(u5_mult_82_SUMB_43__47_) );
  FA_X1 u5_mult_82_S2_43_46 ( .A(u5_mult_82_ab_43__46_), .B(
        u5_mult_82_CARRYB_42__46_), .CI(u5_mult_82_SUMB_42__47_), .CO(
        u5_mult_82_CARRYB_43__46_), .S(u5_mult_82_SUMB_43__46_) );
  FA_X1 u5_mult_82_S2_43_45 ( .A(u5_mult_82_ab_43__45_), .B(
        u5_mult_82_CARRYB_42__45_), .CI(u5_mult_82_SUMB_42__46_), .CO(
        u5_mult_82_CARRYB_43__45_), .S(u5_mult_82_SUMB_43__45_) );
  FA_X1 u5_mult_82_S2_43_42 ( .A(u5_mult_82_ab_43__42_), .B(
        u5_mult_82_CARRYB_42__42_), .CI(u5_mult_82_SUMB_42__43_), .CO(
        u5_mult_82_CARRYB_43__42_), .S(u5_mult_82_SUMB_43__42_) );
  FA_X1 u5_mult_82_S2_43_38 ( .A(u5_mult_82_ab_43__38_), .B(
        u5_mult_82_CARRYB_42__38_), .CI(u5_mult_82_SUMB_42__39_), .CO(
        u5_mult_82_CARRYB_43__38_), .S(u5_mult_82_SUMB_43__38_) );
  FA_X1 u5_mult_82_S2_43_37 ( .A(u5_mult_82_ab_43__37_), .B(
        u5_mult_82_CARRYB_42__37_), .CI(u5_mult_82_SUMB_42__38_), .CO(
        u5_mult_82_CARRYB_43__37_), .S(u5_mult_82_SUMB_43__37_) );
  FA_X1 u5_mult_82_S2_43_36 ( .A(u5_mult_82_ab_43__36_), .B(
        u5_mult_82_CARRYB_42__36_), .CI(u5_mult_82_SUMB_42__37_), .CO(
        u5_mult_82_CARRYB_43__36_), .S(u5_mult_82_SUMB_43__36_) );
  FA_X1 u5_mult_82_S2_43_34 ( .A(u5_mult_82_ab_43__34_), .B(
        u5_mult_82_CARRYB_42__34_), .CI(u5_mult_82_SUMB_42__35_), .CO(
        u5_mult_82_CARRYB_43__34_), .S(u5_mult_82_SUMB_43__34_) );
  FA_X1 u5_mult_82_S2_43_32 ( .A(u5_mult_82_ab_43__32_), .B(
        u5_mult_82_CARRYB_42__32_), .CI(u5_mult_82_SUMB_42__33_), .CO(
        u5_mult_82_CARRYB_43__32_), .S(u5_mult_82_SUMB_43__32_) );
  FA_X1 u5_mult_82_S2_43_31 ( .A(u5_mult_82_ab_43__31_), .B(
        u5_mult_82_CARRYB_42__31_), .CI(u5_mult_82_SUMB_42__32_), .CO(
        u5_mult_82_CARRYB_43__31_), .S(u5_mult_82_SUMB_43__31_) );
  FA_X1 u5_mult_82_S2_43_30 ( .A(u5_mult_82_SUMB_42__31_), .B(
        u5_mult_82_CARRYB_42__30_), .CI(u5_mult_82_ab_43__30_), .CO(
        u5_mult_82_CARRYB_43__30_), .S(u5_mult_82_SUMB_43__30_) );
  FA_X1 u5_mult_82_S2_43_29 ( .A(u5_mult_82_ab_43__29_), .B(
        u5_mult_82_CARRYB_42__29_), .CI(u5_mult_82_SUMB_42__30_), .CO(
        u5_mult_82_CARRYB_43__29_), .S(u5_mult_82_SUMB_43__29_) );
  FA_X1 u5_mult_82_S2_43_28 ( .A(u5_mult_82_ab_43__28_), .B(
        u5_mult_82_CARRYB_42__28_), .CI(u5_mult_82_SUMB_42__29_), .CO(
        u5_mult_82_CARRYB_43__28_), .S(u5_mult_82_SUMB_43__28_) );
  FA_X1 u5_mult_82_S2_43_27 ( .A(u5_mult_82_ab_43__27_), .B(
        u5_mult_82_CARRYB_42__27_), .CI(u5_mult_82_SUMB_42__28_), .CO(
        u5_mult_82_CARRYB_43__27_), .S(u5_mult_82_SUMB_43__27_) );
  FA_X1 u5_mult_82_S2_43_26 ( .A(u5_mult_82_ab_43__26_), .B(
        u5_mult_82_CARRYB_42__26_), .CI(u5_mult_82_SUMB_42__27_), .CO(
        u5_mult_82_CARRYB_43__26_), .S(u5_mult_82_SUMB_43__26_) );
  FA_X1 u5_mult_82_S2_43_25 ( .A(u5_mult_82_CARRYB_42__25_), .B(
        u5_mult_82_ab_43__25_), .CI(u5_mult_82_SUMB_42__26_), .CO(
        u5_mult_82_CARRYB_43__25_), .S(u5_mult_82_SUMB_43__25_) );
  FA_X1 u5_mult_82_S2_43_23 ( .A(u5_mult_82_ab_43__23_), .B(
        u5_mult_82_CARRYB_42__23_), .CI(u5_mult_82_SUMB_42__24_), .CO(
        u5_mult_82_CARRYB_43__23_), .S(u5_mult_82_SUMB_43__23_) );
  FA_X1 u5_mult_82_S2_43_3 ( .A(u5_mult_82_CARRYB_42__3_), .B(
        u5_mult_82_ab_43__3_), .CI(u5_mult_82_SUMB_42__4_), .CO(
        u5_mult_82_CARRYB_43__3_), .S(u5_mult_82_SUMB_43__3_) );
  FA_X1 u5_mult_82_S3_44_51 ( .A(u5_mult_82_ab_44__51_), .B(
        u5_mult_82_CARRYB_43__51_), .CI(u5_mult_82_ab_43__52_), .CO(
        u5_mult_82_CARRYB_44__51_), .S(u5_mult_82_SUMB_44__51_) );
  FA_X1 u5_mult_82_S2_44_50 ( .A(u5_mult_82_ab_44__50_), .B(
        u5_mult_82_CARRYB_43__50_), .CI(u5_mult_82_SUMB_43__51_), .CO(
        u5_mult_82_CARRYB_44__50_), .S(u5_mult_82_SUMB_44__50_) );
  FA_X1 u5_mult_82_S2_44_49 ( .A(u5_mult_82_ab_44__49_), .B(
        u5_mult_82_CARRYB_43__49_), .CI(u5_mult_82_SUMB_43__50_), .CO(
        u5_mult_82_CARRYB_44__49_), .S(u5_mult_82_SUMB_44__49_) );
  FA_X1 u5_mult_82_S2_44_48 ( .A(u5_mult_82_ab_44__48_), .B(
        u5_mult_82_CARRYB_43__48_), .CI(u5_mult_82_SUMB_43__49_), .CO(
        u5_mult_82_CARRYB_44__48_), .S(u5_mult_82_SUMB_44__48_) );
  FA_X1 u5_mult_82_S2_44_47 ( .A(u5_mult_82_ab_44__47_), .B(
        u5_mult_82_CARRYB_43__47_), .CI(u5_mult_82_SUMB_43__48_), .CO(
        u5_mult_82_CARRYB_44__47_), .S(u5_mult_82_SUMB_44__47_) );
  FA_X1 u5_mult_82_S2_44_46 ( .A(u5_mult_82_ab_44__46_), .B(
        u5_mult_82_CARRYB_43__46_), .CI(u5_mult_82_SUMB_43__47_), .CO(
        u5_mult_82_CARRYB_44__46_), .S(u5_mult_82_SUMB_44__46_) );
  FA_X1 u5_mult_82_S2_44_45 ( .A(u5_mult_82_CARRYB_43__45_), .B(
        u5_mult_82_ab_44__45_), .CI(u5_mult_82_SUMB_43__46_), .CO(
        u5_mult_82_CARRYB_44__45_), .S(u5_mult_82_SUMB_44__45_) );
  FA_X1 u5_mult_82_S2_44_40 ( .A(u5_mult_82_ab_44__40_), .B(
        u5_mult_82_CARRYB_43__40_), .CI(u5_mult_82_SUMB_43__41_), .CO(
        u5_mult_82_CARRYB_44__40_), .S(u5_mult_82_SUMB_44__40_) );
  FA_X1 u5_mult_82_S2_44_38 ( .A(u5_mult_82_ab_44__38_), .B(
        u5_mult_82_CARRYB_43__38_), .CI(u5_mult_82_SUMB_43__39_), .CO(
        u5_mult_82_CARRYB_44__38_), .S(u5_mult_82_SUMB_44__38_) );
  FA_X1 u5_mult_82_S2_44_37 ( .A(u5_mult_82_ab_44__37_), .B(
        u5_mult_82_CARRYB_43__37_), .CI(u5_mult_82_SUMB_43__38_), .CO(
        u5_mult_82_CARRYB_44__37_), .S(u5_mult_82_SUMB_44__37_) );
  FA_X1 u5_mult_82_S2_44_36 ( .A(u5_mult_82_ab_44__36_), .B(
        u5_mult_82_CARRYB_43__36_), .CI(u5_mult_82_SUMB_43__37_), .CO(
        u5_mult_82_CARRYB_44__36_), .S(u5_mult_82_SUMB_44__36_) );
  FA_X1 u5_mult_82_S2_44_34 ( .A(u5_mult_82_ab_44__34_), .B(
        u5_mult_82_CARRYB_43__34_), .CI(u5_mult_82_SUMB_43__35_), .CO(
        u5_mult_82_CARRYB_44__34_), .S(u5_mult_82_SUMB_44__34_) );
  FA_X1 u5_mult_82_S2_44_33 ( .A(u5_mult_82_ab_44__33_), .B(
        u5_mult_82_CARRYB_43__33_), .CI(u5_mult_82_SUMB_43__34_), .CO(
        u5_mult_82_CARRYB_44__33_), .S(u5_mult_82_SUMB_44__33_) );
  FA_X1 u5_mult_82_S2_44_30 ( .A(u5_mult_82_ab_44__30_), .B(
        u5_mult_82_CARRYB_43__30_), .CI(u5_mult_82_SUMB_43__31_), .CO(
        u5_mult_82_CARRYB_44__30_), .S(u5_mult_82_SUMB_44__30_) );
  FA_X1 u5_mult_82_S2_44_29 ( .A(u5_mult_82_ab_44__29_), .B(
        u5_mult_82_CARRYB_43__29_), .CI(u5_mult_82_SUMB_43__30_), .CO(
        u5_mult_82_CARRYB_44__29_), .S(u5_mult_82_SUMB_44__29_) );
  FA_X1 u5_mult_82_S2_44_28 ( .A(u5_mult_82_ab_44__28_), .B(
        u5_mult_82_CARRYB_43__28_), .CI(u5_mult_82_SUMB_43__29_), .CO(
        u5_mult_82_CARRYB_44__28_), .S(u5_mult_82_SUMB_44__28_) );
  FA_X1 u5_mult_82_S2_44_27 ( .A(u5_mult_82_ab_44__27_), .B(
        u5_mult_82_CARRYB_43__27_), .CI(u5_mult_82_SUMB_43__28_), .CO(
        u5_mult_82_CARRYB_44__27_), .S(u5_mult_82_SUMB_44__27_) );
  FA_X1 u5_mult_82_S2_44_25 ( .A(u5_mult_82_ab_44__25_), .B(
        u5_mult_82_CARRYB_43__25_), .CI(u5_mult_82_SUMB_43__26_), .CO(
        u5_mult_82_CARRYB_44__25_), .S(u5_mult_82_SUMB_44__25_) );
  FA_X1 u5_mult_82_S2_44_17 ( .A(u5_mult_82_SUMB_43__18_), .B(
        u5_mult_82_CARRYB_43__17_), .CI(u5_mult_82_ab_44__17_), .CO(
        u5_mult_82_CARRYB_44__17_), .S(u5_mult_82_SUMB_44__17_) );
  FA_X1 u5_mult_82_S2_44_15 ( .A(u5_mult_82_ab_44__15_), .B(
        u5_mult_82_CARRYB_43__15_), .CI(u5_mult_82_SUMB_43__16_), .CO(
        u5_mult_82_CARRYB_44__15_), .S(u5_mult_82_SUMB_44__15_) );
  FA_X1 u5_mult_82_S2_44_13 ( .A(u5_mult_82_ab_44__13_), .B(
        u5_mult_82_CARRYB_43__13_), .CI(u5_mult_82_SUMB_43__14_), .CO(
        u5_mult_82_CARRYB_44__13_), .S(u5_mult_82_SUMB_44__13_) );
  FA_X1 u5_mult_82_S2_44_7 ( .A(u5_mult_82_CARRYB_43__7_), .B(
        u5_mult_82_ab_44__7_), .CI(u5_mult_82_SUMB_43__8_), .CO(
        u5_mult_82_CARRYB_44__7_), .S(u5_mult_82_SUMB_44__7_) );
  FA_X1 u5_mult_82_S2_44_3 ( .A(u5_mult_82_SUMB_43__4_), .B(
        u5_mult_82_ab_44__3_), .CI(u5_mult_82_CARRYB_43__3_), .CO(
        u5_mult_82_CARRYB_44__3_), .S(u5_mult_82_SUMB_44__3_) );
  FA_X1 u5_mult_82_S2_44_1 ( .A(u5_mult_82_ab_44__1_), .B(
        u5_mult_82_CARRYB_43__1_), .CI(u5_mult_82_SUMB_43__2_), .CO(
        u5_mult_82_CARRYB_44__1_), .S(u5_mult_82_SUMB_44__1_) );
  FA_X1 u5_mult_82_S3_45_51 ( .A(u5_mult_82_ab_45__51_), .B(
        u5_mult_82_CARRYB_44__51_), .CI(u5_mult_82_ab_44__52_), .CO(
        u5_mult_82_CARRYB_45__51_), .S(u5_mult_82_SUMB_45__51_) );
  FA_X1 u5_mult_82_S2_45_50 ( .A(u5_mult_82_ab_45__50_), .B(
        u5_mult_82_CARRYB_44__50_), .CI(u5_mult_82_SUMB_44__51_), .CO(
        u5_mult_82_CARRYB_45__50_), .S(u5_mult_82_SUMB_45__50_) );
  FA_X1 u5_mult_82_S2_45_49 ( .A(u5_mult_82_ab_45__49_), .B(
        u5_mult_82_CARRYB_44__49_), .CI(u5_mult_82_SUMB_44__50_), .CO(
        u5_mult_82_CARRYB_45__49_), .S(u5_mult_82_SUMB_45__49_) );
  FA_X1 u5_mult_82_S2_45_48 ( .A(u5_mult_82_ab_45__48_), .B(
        u5_mult_82_CARRYB_44__48_), .CI(u5_mult_82_SUMB_44__49_), .CO(
        u5_mult_82_CARRYB_45__48_), .S(u5_mult_82_SUMB_45__48_) );
  FA_X1 u5_mult_82_S2_45_47 ( .A(u5_mult_82_ab_45__47_), .B(
        u5_mult_82_CARRYB_44__47_), .CI(u5_mult_82_SUMB_44__48_), .CO(
        u5_mult_82_CARRYB_45__47_), .S(u5_mult_82_SUMB_45__47_) );
  FA_X1 u5_mult_82_S2_45_46 ( .A(u5_mult_82_ab_45__46_), .B(
        u5_mult_82_CARRYB_44__46_), .CI(u5_mult_82_SUMB_44__47_), .CO(
        u5_mult_82_CARRYB_45__46_), .S(u5_mult_82_SUMB_45__46_) );
  FA_X1 u5_mult_82_S2_45_45 ( .A(u5_mult_82_ab_45__45_), .B(
        u5_mult_82_CARRYB_44__45_), .CI(u5_mult_82_SUMB_44__46_), .CO(
        u5_mult_82_CARRYB_45__45_), .S(u5_mult_82_SUMB_45__45_) );
  FA_X1 u5_mult_82_S2_45_44 ( .A(u5_mult_82_ab_45__44_), .B(
        u5_mult_82_CARRYB_44__44_), .CI(u5_mult_82_SUMB_44__45_), .CO(
        u5_mult_82_CARRYB_45__44_), .S(u5_mult_82_SUMB_45__44_) );
  FA_X1 u5_mult_82_S2_45_42 ( .A(u5_mult_82_ab_45__42_), .B(
        u5_mult_82_CARRYB_44__42_), .CI(u5_mult_82_SUMB_44__43_), .CO(
        u5_mult_82_CARRYB_45__42_), .S(u5_mult_82_SUMB_45__42_) );
  FA_X1 u5_mult_82_S2_45_41 ( .A(u5_mult_82_CARRYB_44__41_), .B(
        u5_mult_82_ab_45__41_), .CI(u5_mult_82_SUMB_44__42_), .CO(
        u5_mult_82_CARRYB_45__41_), .S(u5_mult_82_SUMB_45__41_) );
  FA_X1 u5_mult_82_S2_45_40 ( .A(u5_mult_82_CARRYB_44__40_), .B(
        u5_mult_82_ab_45__40_), .CI(u5_mult_82_SUMB_44__41_), .CO(
        u5_mult_82_CARRYB_45__40_), .S(u5_mult_82_SUMB_45__40_) );
  FA_X1 u5_mult_82_S2_45_38 ( .A(u5_mult_82_ab_45__38_), .B(
        u5_mult_82_CARRYB_44__38_), .CI(u5_mult_82_SUMB_44__39_), .CO(
        u5_mult_82_CARRYB_45__38_), .S(u5_mult_82_SUMB_45__38_) );
  FA_X1 u5_mult_82_S2_45_37 ( .A(u5_mult_82_ab_45__37_), .B(
        u5_mult_82_CARRYB_44__37_), .CI(u5_mult_82_SUMB_44__38_), .CO(
        u5_mult_82_CARRYB_45__37_), .S(u5_mult_82_SUMB_45__37_) );
  FA_X1 u5_mult_82_S2_45_36 ( .A(u5_mult_82_ab_45__36_), .B(
        u5_mult_82_CARRYB_44__36_), .CI(u5_mult_82_SUMB_44__37_), .CO(
        u5_mult_82_CARRYB_45__36_), .S(u5_mult_82_SUMB_45__36_) );
  FA_X1 u5_mult_82_S2_45_31 ( .A(u5_mult_82_CARRYB_44__31_), .B(
        u5_mult_82_ab_45__31_), .CI(u5_mult_82_SUMB_44__32_), .CO(
        u5_mult_82_CARRYB_45__31_), .S(u5_mult_82_SUMB_45__31_) );
  FA_X1 u5_mult_82_S2_45_25 ( .A(u5_mult_82_ab_45__25_), .B(
        u5_mult_82_CARRYB_44__25_), .CI(u5_mult_82_SUMB_44__26_), .CO(
        u5_mult_82_CARRYB_45__25_), .S(u5_mult_82_SUMB_45__25_) );
  FA_X1 u5_mult_82_S2_45_22 ( .A(u5_mult_82_ab_45__22_), .B(
        u5_mult_82_CARRYB_44__22_), .CI(u5_mult_82_SUMB_44__23_), .CO(
        u5_mult_82_CARRYB_45__22_), .S(u5_mult_82_SUMB_45__22_) );
  FA_X1 u5_mult_82_S2_45_21 ( .A(u5_mult_82_ab_45__21_), .B(
        u5_mult_82_CARRYB_44__21_), .CI(u5_mult_82_SUMB_44__22_), .CO(
        u5_mult_82_CARRYB_45__21_), .S(u5_mult_82_SUMB_45__21_) );
  FA_X1 u5_mult_82_S2_45_19 ( .A(u5_mult_82_CARRYB_44__19_), .B(
        u5_mult_82_ab_45__19_), .CI(u5_mult_82_SUMB_44__20_), .CO(
        u5_mult_82_CARRYB_45__19_), .S(u5_mult_82_SUMB_45__19_) );
  FA_X1 u5_mult_82_S2_45_16 ( .A(u5_mult_82_ab_45__16_), .B(
        u5_mult_82_CARRYB_44__16_), .CI(u5_mult_82_SUMB_44__17_), .CO(
        u5_mult_82_CARRYB_45__16_), .S(u5_mult_82_SUMB_45__16_) );
  FA_X1 u5_mult_82_S1_45_0 ( .A(u5_mult_82_CARRYB_44__0_), .B(
        u5_mult_82_ab_45__0_), .CI(u5_mult_82_SUMB_44__1_), .CO(
        u5_mult_82_CARRYB_45__0_), .S(u5_N45) );
  FA_X1 u5_mult_82_S3_46_51 ( .A(u5_mult_82_ab_46__51_), .B(
        u5_mult_82_CARRYB_45__51_), .CI(u5_mult_82_ab_45__52_), .CO(
        u5_mult_82_CARRYB_46__51_), .S(u5_mult_82_SUMB_46__51_) );
  FA_X1 u5_mult_82_S2_46_50 ( .A(u5_mult_82_ab_46__50_), .B(
        u5_mult_82_CARRYB_45__50_), .CI(u5_mult_82_SUMB_45__51_), .CO(
        u5_mult_82_CARRYB_46__50_), .S(u5_mult_82_SUMB_46__50_) );
  FA_X1 u5_mult_82_S2_46_49 ( .A(u5_mult_82_ab_46__49_), .B(
        u5_mult_82_CARRYB_45__49_), .CI(u5_mult_82_SUMB_45__50_), .CO(
        u5_mult_82_CARRYB_46__49_), .S(u5_mult_82_SUMB_46__49_) );
  FA_X1 u5_mult_82_S2_46_48 ( .A(u5_mult_82_ab_46__48_), .B(
        u5_mult_82_CARRYB_45__48_), .CI(u5_mult_82_SUMB_45__49_), .CO(
        u5_mult_82_CARRYB_46__48_), .S(u5_mult_82_SUMB_46__48_) );
  FA_X1 u5_mult_82_S2_46_47 ( .A(u5_mult_82_ab_46__47_), .B(
        u5_mult_82_CARRYB_45__47_), .CI(u5_mult_82_SUMB_45__48_), .CO(
        u5_mult_82_CARRYB_46__47_), .S(u5_mult_82_SUMB_46__47_) );
  FA_X1 u5_mult_82_S2_46_46 ( .A(u5_mult_82_ab_46__46_), .B(
        u5_mult_82_CARRYB_45__46_), .CI(u5_mult_82_SUMB_45__47_), .CO(
        u5_mult_82_CARRYB_46__46_), .S(u5_mult_82_SUMB_46__46_) );
  FA_X1 u5_mult_82_S2_46_45 ( .A(u5_mult_82_ab_46__45_), .B(
        u5_mult_82_CARRYB_45__45_), .CI(u5_mult_82_SUMB_45__46_), .CO(
        u5_mult_82_CARRYB_46__45_), .S(u5_mult_82_SUMB_46__45_) );
  FA_X1 u5_mult_82_S2_46_44 ( .A(u5_mult_82_ab_46__44_), .B(
        u5_mult_82_CARRYB_45__44_), .CI(u5_mult_82_SUMB_45__45_), .CO(
        u5_mult_82_CARRYB_46__44_), .S(u5_mult_82_SUMB_46__44_) );
  FA_X1 u5_mult_82_S2_46_43 ( .A(u5_mult_82_ab_46__43_), .B(
        u5_mult_82_CARRYB_45__43_), .CI(u5_mult_82_SUMB_45__44_), .CO(
        u5_mult_82_CARRYB_46__43_), .S(u5_mult_82_SUMB_46__43_) );
  FA_X1 u5_mult_82_S2_46_42 ( .A(u5_mult_82_ab_46__42_), .B(
        u5_mult_82_CARRYB_45__42_), .CI(u5_mult_82_SUMB_45__43_), .CO(
        u5_mult_82_CARRYB_46__42_), .S(u5_mult_82_SUMB_46__42_) );
  FA_X1 u5_mult_82_S2_46_41 ( .A(u5_mult_82_ab_46__41_), .B(
        u5_mult_82_CARRYB_45__41_), .CI(u5_mult_82_SUMB_45__42_), .CO(
        u5_mult_82_CARRYB_46__41_), .S(u5_mult_82_SUMB_46__41_) );
  FA_X1 u5_mult_82_S2_46_40 ( .A(u5_mult_82_ab_46__40_), .B(
        u5_mult_82_CARRYB_45__40_), .CI(u5_mult_82_SUMB_45__41_), .CO(
        u5_mult_82_CARRYB_46__40_), .S(u5_mult_82_SUMB_46__40_) );
  FA_X1 u5_mult_82_S2_46_38 ( .A(u5_mult_82_CARRYB_45__38_), .B(
        u5_mult_82_ab_46__38_), .CI(u5_mult_82_SUMB_45__39_), .CO(
        u5_mult_82_CARRYB_46__38_), .S(u5_mult_82_SUMB_46__38_) );
  FA_X1 u5_mult_82_S2_46_37 ( .A(u5_mult_82_ab_46__37_), .B(
        u5_mult_82_CARRYB_45__37_), .CI(u5_mult_82_SUMB_45__38_), .CO(
        u5_mult_82_CARRYB_46__37_), .S(u5_mult_82_SUMB_46__37_) );
  FA_X1 u5_mult_82_S2_46_24 ( .A(u5_mult_82_ab_46__24_), .B(
        u5_mult_82_CARRYB_45__24_), .CI(u5_mult_82_SUMB_45__25_), .CO(
        u5_mult_82_CARRYB_46__24_), .S(u5_mult_82_SUMB_46__24_) );
  FA_X1 u5_mult_82_S2_46_21 ( .A(u5_mult_82_ab_46__21_), .B(
        u5_mult_82_CARRYB_45__21_), .CI(u5_mult_82_SUMB_45__22_), .CO(
        u5_mult_82_CARRYB_46__21_), .S(u5_mult_82_SUMB_46__21_) );
  FA_X1 u5_mult_82_S2_46_20 ( .A(u5_mult_82_ab_46__20_), .B(
        u5_mult_82_CARRYB_45__20_), .CI(u5_mult_82_SUMB_45__21_), .CO(
        u5_mult_82_CARRYB_46__20_), .S(u5_mult_82_SUMB_46__20_) );
  FA_X1 u5_mult_82_S2_46_16 ( .A(u5_mult_82_CARRYB_45__16_), .B(
        u5_mult_82_ab_46__16_), .CI(u5_mult_82_SUMB_45__17_), .CO(
        u5_mult_82_CARRYB_46__16_), .S(u5_mult_82_SUMB_46__16_) );
  FA_X1 u5_mult_82_S2_46_15 ( .A(u5_mult_82_ab_46__15_), .B(
        u5_mult_82_CARRYB_45__15_), .CI(u5_mult_82_SUMB_45__16_), .CO(
        u5_mult_82_CARRYB_46__15_), .S(u5_mult_82_SUMB_46__15_) );
  FA_X1 u5_mult_82_S1_46_0 ( .A(u5_mult_82_SUMB_45__1_), .B(
        u5_mult_82_ab_46__0_), .CI(u5_mult_82_CARRYB_45__0_), .CO(
        u5_mult_82_CARRYB_46__0_), .S(u5_N46) );
  FA_X1 u5_mult_82_S3_47_51 ( .A(u5_mult_82_ab_47__51_), .B(
        u5_mult_82_CARRYB_46__51_), .CI(u5_mult_82_ab_46__52_), .CO(
        u5_mult_82_CARRYB_47__51_), .S(u5_mult_82_SUMB_47__51_) );
  FA_X1 u5_mult_82_S2_47_50 ( .A(u5_mult_82_ab_47__50_), .B(
        u5_mult_82_CARRYB_46__50_), .CI(u5_mult_82_SUMB_46__51_), .CO(
        u5_mult_82_CARRYB_47__50_), .S(u5_mult_82_SUMB_47__50_) );
  FA_X1 u5_mult_82_S2_47_49 ( .A(u5_mult_82_ab_47__49_), .B(
        u5_mult_82_CARRYB_46__49_), .CI(u5_mult_82_SUMB_46__50_), .CO(
        u5_mult_82_CARRYB_47__49_), .S(u5_mult_82_SUMB_47__49_) );
  FA_X1 u5_mult_82_S2_47_48 ( .A(u5_mult_82_ab_47__48_), .B(
        u5_mult_82_CARRYB_46__48_), .CI(u5_mult_82_SUMB_46__49_), .CO(
        u5_mult_82_CARRYB_47__48_), .S(u5_mult_82_SUMB_47__48_) );
  FA_X1 u5_mult_82_S2_47_47 ( .A(u5_mult_82_ab_47__47_), .B(
        u5_mult_82_CARRYB_46__47_), .CI(u5_mult_82_SUMB_46__48_), .CO(
        u5_mult_82_CARRYB_47__47_), .S(u5_mult_82_SUMB_47__47_) );
  FA_X1 u5_mult_82_S2_47_46 ( .A(u5_mult_82_ab_47__46_), .B(
        u5_mult_82_CARRYB_46__46_), .CI(u5_mult_82_SUMB_46__47_), .CO(
        u5_mult_82_CARRYB_47__46_), .S(u5_mult_82_SUMB_47__46_) );
  FA_X1 u5_mult_82_S2_47_45 ( .A(u5_mult_82_ab_47__45_), .B(
        u5_mult_82_CARRYB_46__45_), .CI(u5_mult_82_SUMB_46__46_), .CO(
        u5_mult_82_CARRYB_47__45_), .S(u5_mult_82_SUMB_47__45_) );
  FA_X1 u5_mult_82_S2_47_44 ( .A(u5_mult_82_ab_47__44_), .B(
        u5_mult_82_CARRYB_46__44_), .CI(u5_mult_82_SUMB_46__45_), .CO(
        u5_mult_82_CARRYB_47__44_), .S(u5_mult_82_SUMB_47__44_) );
  FA_X1 u5_mult_82_S2_47_43 ( .A(u5_mult_82_ab_47__43_), .B(
        u5_mult_82_CARRYB_46__43_), .CI(u5_mult_82_SUMB_46__44_), .CO(
        u5_mult_82_CARRYB_47__43_), .S(u5_mult_82_SUMB_47__43_) );
  FA_X1 u5_mult_82_S2_47_42 ( .A(u5_mult_82_ab_47__42_), .B(
        u5_mult_82_CARRYB_46__42_), .CI(u5_mult_82_SUMB_46__43_), .CO(
        u5_mult_82_CARRYB_47__42_), .S(u5_mult_82_SUMB_47__42_) );
  FA_X1 u5_mult_82_S2_47_41 ( .A(u5_mult_82_CARRYB_46__41_), .B(
        u5_mult_82_ab_47__41_), .CI(u5_mult_82_SUMB_46__42_), .CO(
        u5_mult_82_CARRYB_47__41_), .S(u5_mult_82_SUMB_47__41_) );
  FA_X1 u5_mult_82_S2_47_40 ( .A(u5_mult_82_ab_47__40_), .B(
        u5_mult_82_CARRYB_46__40_), .CI(u5_mult_82_SUMB_46__41_), .CO(
        u5_mult_82_CARRYB_47__40_), .S(u5_mult_82_SUMB_47__40_) );
  FA_X1 u5_mult_82_S2_47_38 ( .A(u5_mult_82_ab_47__38_), .B(
        u5_mult_82_CARRYB_46__38_), .CI(u5_mult_82_SUMB_46__39_), .CO(
        u5_mult_82_CARRYB_47__38_), .S(u5_mult_82_SUMB_47__38_) );
  FA_X1 u5_mult_82_S2_47_35 ( .A(u5_mult_82_ab_47__35_), .B(
        u5_mult_82_CARRYB_46__35_), .CI(u5_mult_82_SUMB_46__36_), .CO(
        u5_mult_82_CARRYB_47__35_), .S(u5_mult_82_SUMB_47__35_) );
  FA_X1 u5_mult_82_S2_47_33 ( .A(u5_mult_82_ab_47__33_), .B(
        u5_mult_82_CARRYB_46__33_), .CI(u5_mult_82_SUMB_46__34_), .CO(
        u5_mult_82_CARRYB_47__33_), .S(u5_mult_82_SUMB_47__33_) );
  FA_X1 u5_mult_82_S2_47_30 ( .A(u5_mult_82_ab_47__30_), .B(
        u5_mult_82_CARRYB_46__30_), .CI(u5_mult_82_SUMB_46__31_), .CO(
        u5_mult_82_CARRYB_47__30_), .S(u5_mult_82_SUMB_47__30_) );
  FA_X1 u5_mult_82_S2_47_28 ( .A(u5_mult_82_ab_47__28_), .B(
        u5_mult_82_CARRYB_46__28_), .CI(u5_mult_82_SUMB_46__29_), .CO(
        u5_mult_82_CARRYB_47__28_), .S(u5_mult_82_SUMB_47__28_) );
  FA_X1 u5_mult_82_S2_47_27 ( .A(u5_mult_82_ab_47__27_), .B(
        u5_mult_82_CARRYB_46__27_), .CI(u5_mult_82_SUMB_46__28_), .CO(
        u5_mult_82_CARRYB_47__27_), .S(u5_mult_82_SUMB_47__27_) );
  FA_X1 u5_mult_82_S2_47_26 ( .A(u5_mult_82_ab_47__26_), .B(
        u5_mult_82_CARRYB_46__26_), .CI(u5_mult_82_SUMB_46__27_), .CO(
        u5_mult_82_CARRYB_47__26_), .S(u5_mult_82_SUMB_47__26_) );
  FA_X1 u5_mult_82_S2_47_25 ( .A(u5_mult_82_ab_47__25_), .B(
        u5_mult_82_CARRYB_46__25_), .CI(u5_mult_82_SUMB_46__26_), .CO(
        u5_mult_82_CARRYB_47__25_), .S(u5_mult_82_SUMB_47__25_) );
  FA_X1 u5_mult_82_S2_47_24 ( .A(u5_mult_82_ab_47__24_), .B(
        u5_mult_82_CARRYB_46__24_), .CI(u5_mult_82_SUMB_46__25_), .CO(
        u5_mult_82_CARRYB_47__24_), .S(u5_mult_82_SUMB_47__24_) );
  FA_X1 u5_mult_82_S2_47_22 ( .A(u5_mult_82_ab_47__22_), .B(
        u5_mult_82_CARRYB_46__22_), .CI(u5_mult_82_SUMB_46__23_), .CO(
        u5_mult_82_CARRYB_47__22_), .S(u5_mult_82_SUMB_47__22_) );
  FA_X1 u5_mult_82_S3_48_51 ( .A(u5_mult_82_ab_48__51_), .B(
        u5_mult_82_CARRYB_47__51_), .CI(u5_mult_82_ab_47__52_), .CO(
        u5_mult_82_CARRYB_48__51_), .S(u5_mult_82_SUMB_48__51_) );
  FA_X1 u5_mult_82_S2_48_50 ( .A(u5_mult_82_ab_48__50_), .B(
        u5_mult_82_CARRYB_47__50_), .CI(u5_mult_82_SUMB_47__51_), .CO(
        u5_mult_82_CARRYB_48__50_), .S(u5_mult_82_SUMB_48__50_) );
  FA_X1 u5_mult_82_S2_48_49 ( .A(u5_mult_82_ab_48__49_), .B(
        u5_mult_82_CARRYB_47__49_), .CI(u5_mult_82_SUMB_47__50_), .CO(
        u5_mult_82_CARRYB_48__49_), .S(u5_mult_82_SUMB_48__49_) );
  FA_X1 u5_mult_82_S2_48_48 ( .A(u5_mult_82_ab_48__48_), .B(
        u5_mult_82_CARRYB_47__48_), .CI(u5_mult_82_SUMB_47__49_), .CO(
        u5_mult_82_CARRYB_48__48_), .S(u5_mult_82_SUMB_48__48_) );
  FA_X1 u5_mult_82_S2_48_47 ( .A(u5_mult_82_ab_48__47_), .B(
        u5_mult_82_CARRYB_47__47_), .CI(u5_mult_82_SUMB_47__48_), .CO(
        u5_mult_82_CARRYB_48__47_), .S(u5_mult_82_SUMB_48__47_) );
  FA_X1 u5_mult_82_S2_48_46 ( .A(u5_mult_82_ab_48__46_), .B(
        u5_mult_82_CARRYB_47__46_), .CI(u5_mult_82_SUMB_47__47_), .CO(
        u5_mult_82_CARRYB_48__46_), .S(u5_mult_82_SUMB_48__46_) );
  FA_X1 u5_mult_82_S2_48_45 ( .A(u5_mult_82_ab_48__45_), .B(
        u5_mult_82_CARRYB_47__45_), .CI(u5_mult_82_SUMB_47__46_), .CO(
        u5_mult_82_CARRYB_48__45_), .S(u5_mult_82_SUMB_48__45_) );
  FA_X1 u5_mult_82_S2_48_44 ( .A(u5_mult_82_ab_48__44_), .B(
        u5_mult_82_CARRYB_47__44_), .CI(u5_mult_82_SUMB_47__45_), .CO(
        u5_mult_82_CARRYB_48__44_), .S(u5_mult_82_SUMB_48__44_) );
  FA_X1 u5_mult_82_S2_48_43 ( .A(u5_mult_82_ab_48__43_), .B(
        u5_mult_82_CARRYB_47__43_), .CI(u5_mult_82_SUMB_47__44_), .CO(
        u5_mult_82_CARRYB_48__43_), .S(u5_mult_82_SUMB_48__43_) );
  FA_X1 u5_mult_82_S2_48_42 ( .A(u5_mult_82_ab_48__42_), .B(
        u5_mult_82_CARRYB_47__42_), .CI(u5_mult_82_SUMB_47__43_), .CO(
        u5_mult_82_CARRYB_48__42_), .S(u5_mult_82_SUMB_48__42_) );
  FA_X1 u5_mult_82_S2_48_41 ( .A(u5_mult_82_ab_48__41_), .B(
        u5_mult_82_CARRYB_47__41_), .CI(u5_mult_82_SUMB_47__42_), .CO(
        u5_mult_82_CARRYB_48__41_), .S(u5_mult_82_SUMB_48__41_) );
  FA_X1 u5_mult_82_S2_48_40 ( .A(u5_mult_82_ab_48__40_), .B(
        u5_mult_82_CARRYB_47__40_), .CI(u5_mult_82_SUMB_47__41_), .CO(
        u5_mult_82_CARRYB_48__40_), .S(u5_mult_82_SUMB_48__40_) );
  FA_X1 u5_mult_82_S2_48_39 ( .A(u5_mult_82_ab_48__39_), .B(
        u5_mult_82_CARRYB_47__39_), .CI(u5_mult_82_SUMB_47__40_), .CO(
        u5_mult_82_CARRYB_48__39_), .S(u5_mult_82_SUMB_48__39_) );
  FA_X1 u5_mult_82_S2_48_27 ( .A(u5_mult_82_CARRYB_47__27_), .B(
        u5_mult_82_ab_48__27_), .CI(u5_mult_82_SUMB_47__28_), .CO(
        u5_mult_82_CARRYB_48__27_), .S(u5_mult_82_SUMB_48__27_) );
  FA_X1 u5_mult_82_S2_48_26 ( .A(u5_mult_82_ab_48__26_), .B(
        u5_mult_82_CARRYB_47__26_), .CI(u5_mult_82_SUMB_47__27_), .CO(
        u5_mult_82_CARRYB_48__26_), .S(u5_mult_82_SUMB_48__26_) );
  FA_X1 u5_mult_82_S2_48_21 ( .A(u5_mult_82_ab_48__21_), .B(
        u5_mult_82_CARRYB_47__21_), .CI(u5_mult_82_SUMB_47__22_), .CO(
        u5_mult_82_CARRYB_48__21_), .S(u5_mult_82_SUMB_48__21_) );
  FA_X1 u5_mult_82_S2_48_16 ( .A(u5_mult_82_ab_48__16_), .B(
        u5_mult_82_CARRYB_47__16_), .CI(u5_mult_82_SUMB_47__17_), .CO(
        u5_mult_82_CARRYB_48__16_), .S(u5_mult_82_SUMB_48__16_) );
  FA_X1 u5_mult_82_S2_48_13 ( .A(u5_mult_82_ab_48__13_), .B(
        u5_mult_82_CARRYB_47__13_), .CI(u5_mult_82_SUMB_47__14_), .CO(
        u5_mult_82_CARRYB_48__13_), .S(u5_mult_82_SUMB_48__13_) );
  FA_X1 u5_mult_82_S2_48_5 ( .A(u5_mult_82_CARRYB_47__5_), .B(
        u5_mult_82_ab_48__5_), .CI(u5_mult_82_SUMB_47__6_), .CO(
        u5_mult_82_CARRYB_48__5_), .S(u5_mult_82_SUMB_48__5_) );
  FA_X1 u5_mult_82_S2_48_3 ( .A(u5_mult_82_ab_48__3_), .B(
        u5_mult_82_CARRYB_47__3_), .CI(u5_mult_82_SUMB_47__4_), .CO(
        u5_mult_82_CARRYB_48__3_), .S(u5_mult_82_SUMB_48__3_) );
  FA_X1 u5_mult_82_S2_48_2 ( .A(u5_mult_82_ab_48__2_), .B(
        u5_mult_82_CARRYB_47__2_), .CI(u5_mult_82_SUMB_47__3_), .CO(
        u5_mult_82_CARRYB_48__2_), .S(u5_mult_82_SUMB_48__2_) );
  FA_X1 u5_mult_82_S3_49_51 ( .A(u5_mult_82_ab_49__51_), .B(
        u5_mult_82_CARRYB_48__51_), .CI(u5_mult_82_ab_48__52_), .CO(
        u5_mult_82_CARRYB_49__51_), .S(u5_mult_82_SUMB_49__51_) );
  FA_X1 u5_mult_82_S2_49_50 ( .A(u5_mult_82_ab_49__50_), .B(
        u5_mult_82_CARRYB_48__50_), .CI(u5_mult_82_SUMB_48__51_), .CO(
        u5_mult_82_CARRYB_49__50_), .S(u5_mult_82_SUMB_49__50_) );
  FA_X1 u5_mult_82_S2_49_49 ( .A(u5_mult_82_ab_49__49_), .B(
        u5_mult_82_CARRYB_48__49_), .CI(u5_mult_82_SUMB_48__50_), .CO(
        u5_mult_82_CARRYB_49__49_), .S(u5_mult_82_SUMB_49__49_) );
  FA_X1 u5_mult_82_S2_49_48 ( .A(u5_mult_82_ab_49__48_), .B(
        u5_mult_82_CARRYB_48__48_), .CI(u5_mult_82_SUMB_48__49_), .CO(
        u5_mult_82_CARRYB_49__48_), .S(u5_mult_82_SUMB_49__48_) );
  FA_X1 u5_mult_82_S2_49_47 ( .A(u5_mult_82_ab_49__47_), .B(
        u5_mult_82_CARRYB_48__47_), .CI(u5_mult_82_SUMB_48__48_), .CO(
        u5_mult_82_CARRYB_49__47_), .S(u5_mult_82_SUMB_49__47_) );
  FA_X1 u5_mult_82_S2_49_46 ( .A(u5_mult_82_ab_49__46_), .B(
        u5_mult_82_CARRYB_48__46_), .CI(u5_mult_82_SUMB_48__47_), .CO(
        u5_mult_82_CARRYB_49__46_), .S(u5_mult_82_SUMB_49__46_) );
  FA_X1 u5_mult_82_S2_49_45 ( .A(u5_mult_82_ab_49__45_), .B(
        u5_mult_82_CARRYB_48__45_), .CI(u5_mult_82_SUMB_48__46_), .CO(
        u5_mult_82_CARRYB_49__45_), .S(u5_mult_82_SUMB_49__45_) );
  FA_X1 u5_mult_82_S2_49_44 ( .A(u5_mult_82_ab_49__44_), .B(
        u5_mult_82_CARRYB_48__44_), .CI(u5_mult_82_SUMB_48__45_), .CO(
        u5_mult_82_CARRYB_49__44_), .S(u5_mult_82_SUMB_49__44_) );
  FA_X1 u5_mult_82_S2_49_43 ( .A(u5_mult_82_ab_49__43_), .B(
        u5_mult_82_CARRYB_48__43_), .CI(u5_mult_82_SUMB_48__44_), .CO(
        u5_mult_82_CARRYB_49__43_), .S(u5_mult_82_SUMB_49__43_) );
  FA_X1 u5_mult_82_S2_49_42 ( .A(u5_mult_82_ab_49__42_), .B(
        u5_mult_82_CARRYB_48__42_), .CI(u5_mult_82_SUMB_48__43_), .CO(
        u5_mult_82_CARRYB_49__42_), .S(u5_mult_82_SUMB_49__42_) );
  FA_X1 u5_mult_82_S2_49_41 ( .A(u5_mult_82_ab_49__41_), .B(
        u5_mult_82_CARRYB_48__41_), .CI(u5_mult_82_SUMB_48__42_), .CO(
        u5_mult_82_CARRYB_49__41_), .S(u5_mult_82_SUMB_49__41_) );
  FA_X1 u5_mult_82_S2_49_40 ( .A(u5_mult_82_ab_49__40_), .B(
        u5_mult_82_CARRYB_48__40_), .CI(u5_mult_82_SUMB_48__41_), .CO(
        u5_mult_82_CARRYB_49__40_), .S(u5_mult_82_SUMB_49__40_) );
  FA_X1 u5_mult_82_S2_49_34 ( .A(u5_mult_82_ab_49__34_), .B(
        u5_mult_82_CARRYB_48__34_), .CI(u5_mult_82_SUMB_48__35_), .CO(
        u5_mult_82_CARRYB_49__34_), .S(u5_mult_82_SUMB_49__34_) );
  FA_X1 u5_mult_82_S2_49_32 ( .A(u5_mult_82_ab_49__32_), .B(
        u5_mult_82_CARRYB_48__32_), .CI(u5_mult_82_SUMB_48__33_), .CO(
        u5_mult_82_CARRYB_49__32_), .S(u5_mult_82_SUMB_49__32_) );
  FA_X1 u5_mult_82_S2_49_30 ( .A(u5_mult_82_ab_49__30_), .B(
        u5_mult_82_CARRYB_48__30_), .CI(u5_mult_82_SUMB_48__31_), .CO(
        u5_mult_82_CARRYB_49__30_), .S(u5_mult_82_SUMB_49__30_) );
  FA_X1 u5_mult_82_S2_49_28 ( .A(u5_mult_82_ab_49__28_), .B(
        u5_mult_82_CARRYB_48__28_), .CI(u5_mult_82_SUMB_48__29_), .CO(
        u5_mult_82_CARRYB_49__28_), .S(u5_mult_82_SUMB_49__28_) );
  FA_X1 u5_mult_82_S2_49_27 ( .A(u5_mult_82_ab_49__27_), .B(
        u5_mult_82_CARRYB_48__27_), .CI(u5_mult_82_SUMB_48__28_), .CO(
        u5_mult_82_CARRYB_49__27_), .S(u5_mult_82_SUMB_49__27_) );
  FA_X1 u5_mult_82_S2_49_22 ( .A(u5_mult_82_ab_49__22_), .B(
        u5_mult_82_CARRYB_48__22_), .CI(u5_mult_82_SUMB_48__23_), .CO(
        u5_mult_82_CARRYB_49__22_), .S(u5_mult_82_SUMB_49__22_) );
  FA_X1 u5_mult_82_S2_49_20 ( .A(u5_mult_82_ab_49__20_), .B(
        u5_mult_82_CARRYB_48__20_), .CI(u5_mult_82_SUMB_48__21_), .CO(
        u5_mult_82_CARRYB_49__20_), .S(u5_mult_82_SUMB_49__20_) );
  FA_X1 u5_mult_82_S2_49_9 ( .A(u5_mult_82_ab_49__9_), .B(
        u5_mult_82_CARRYB_48__9_), .CI(u5_mult_82_SUMB_48__10_), .CO(
        u5_mult_82_CARRYB_49__9_), .S(u5_mult_82_SUMB_49__9_) );
  FA_X1 u5_mult_82_S2_49_4 ( .A(u5_mult_82_ab_49__4_), .B(
        u5_mult_82_CARRYB_48__4_), .CI(u5_mult_82_SUMB_48__5_), .CO(
        u5_mult_82_CARRYB_49__4_), .S(u5_mult_82_SUMB_49__4_) );
  FA_X1 u5_mult_82_S2_49_3 ( .A(u5_mult_82_ab_49__3_), .B(
        u5_mult_82_CARRYB_48__3_), .CI(u5_mult_82_SUMB_48__4_), .CO(
        u5_mult_82_CARRYB_49__3_), .S(u5_mult_82_SUMB_49__3_) );
  FA_X1 u5_mult_82_S2_49_2 ( .A(u5_mult_82_CARRYB_48__2_), .B(
        u5_mult_82_ab_49__2_), .CI(u5_mult_82_SUMB_48__3_), .CO(
        u5_mult_82_CARRYB_49__2_), .S(u5_mult_82_SUMB_49__2_) );
  FA_X1 u5_mult_82_S2_49_1 ( .A(u5_mult_82_CARRYB_48__1_), .B(
        u5_mult_82_ab_49__1_), .CI(u5_mult_82_SUMB_48__2_), .CO(
        u5_mult_82_CARRYB_49__1_), .S(u5_mult_82_SUMB_49__1_) );
  FA_X1 u5_mult_82_S1_49_0 ( .A(u5_mult_82_CARRYB_48__0_), .B(
        u5_mult_82_ab_49__0_), .CI(u5_mult_82_SUMB_48__1_), .CO(
        u5_mult_82_CARRYB_49__0_), .S(u5_N49) );
  FA_X1 u5_mult_82_S3_50_51 ( .A(u5_mult_82_ab_50__51_), .B(
        u5_mult_82_CARRYB_49__51_), .CI(u5_mult_82_ab_49__52_), .CO(
        u5_mult_82_CARRYB_50__51_), .S(u5_mult_82_SUMB_50__51_) );
  FA_X1 u5_mult_82_S2_50_50 ( .A(u5_mult_82_ab_50__50_), .B(
        u5_mult_82_CARRYB_49__50_), .CI(u5_mult_82_SUMB_49__51_), .CO(
        u5_mult_82_CARRYB_50__50_), .S(u5_mult_82_SUMB_50__50_) );
  FA_X1 u5_mult_82_S2_50_49 ( .A(u5_mult_82_ab_50__49_), .B(
        u5_mult_82_CARRYB_49__49_), .CI(u5_mult_82_SUMB_49__50_), .CO(
        u5_mult_82_CARRYB_50__49_), .S(u5_mult_82_SUMB_50__49_) );
  FA_X1 u5_mult_82_S2_50_48 ( .A(u5_mult_82_ab_50__48_), .B(
        u5_mult_82_CARRYB_49__48_), .CI(u5_mult_82_SUMB_49__49_), .CO(
        u5_mult_82_CARRYB_50__48_), .S(u5_mult_82_SUMB_50__48_) );
  FA_X1 u5_mult_82_S2_50_47 ( .A(u5_mult_82_ab_50__47_), .B(
        u5_mult_82_CARRYB_49__47_), .CI(u5_mult_82_SUMB_49__48_), .CO(
        u5_mult_82_CARRYB_50__47_), .S(u5_mult_82_SUMB_50__47_) );
  FA_X1 u5_mult_82_S2_50_46 ( .A(u5_mult_82_ab_50__46_), .B(
        u5_mult_82_CARRYB_49__46_), .CI(u5_mult_82_SUMB_49__47_), .CO(
        u5_mult_82_CARRYB_50__46_), .S(u5_mult_82_SUMB_50__46_) );
  FA_X1 u5_mult_82_S2_50_45 ( .A(u5_mult_82_ab_50__45_), .B(
        u5_mult_82_CARRYB_49__45_), .CI(u5_mult_82_SUMB_49__46_), .CO(
        u5_mult_82_CARRYB_50__45_), .S(u5_mult_82_SUMB_50__45_) );
  FA_X1 u5_mult_82_S2_50_44 ( .A(u5_mult_82_ab_50__44_), .B(
        u5_mult_82_CARRYB_49__44_), .CI(u5_mult_82_SUMB_49__45_), .CO(
        u5_mult_82_CARRYB_50__44_), .S(u5_mult_82_SUMB_50__44_) );
  FA_X1 u5_mult_82_S2_50_43 ( .A(u5_mult_82_ab_50__43_), .B(
        u5_mult_82_CARRYB_49__43_), .CI(u5_mult_82_SUMB_49__44_), .CO(
        u5_mult_82_CARRYB_50__43_), .S(u5_mult_82_SUMB_50__43_) );
  FA_X1 u5_mult_82_S2_50_42 ( .A(u5_mult_82_ab_50__42_), .B(
        u5_mult_82_CARRYB_49__42_), .CI(u5_mult_82_SUMB_49__43_), .CO(
        u5_mult_82_CARRYB_50__42_), .S(u5_mult_82_SUMB_50__42_) );
  FA_X1 u5_mult_82_S2_50_41 ( .A(u5_mult_82_ab_50__41_), .B(
        u5_mult_82_CARRYB_49__41_), .CI(u5_mult_82_SUMB_49__42_), .CO(
        u5_mult_82_CARRYB_50__41_), .S(u5_mult_82_SUMB_50__41_) );
  FA_X1 u5_mult_82_S2_50_40 ( .A(u5_mult_82_ab_50__40_), .B(
        u5_mult_82_CARRYB_49__40_), .CI(u5_mult_82_SUMB_49__41_), .CO(
        u5_mult_82_CARRYB_50__40_), .S(u5_mult_82_SUMB_50__40_) );
  FA_X1 u5_mult_82_S2_50_39 ( .A(u5_mult_82_ab_50__39_), .B(
        u5_mult_82_CARRYB_49__39_), .CI(u5_mult_82_SUMB_49__40_), .CO(
        u5_mult_82_CARRYB_50__39_), .S(u5_mult_82_SUMB_50__39_) );
  FA_X1 u5_mult_82_S2_50_36 ( .A(u5_mult_82_ab_50__36_), .B(
        u5_mult_82_CARRYB_49__36_), .CI(u5_mult_82_SUMB_49__37_), .CO(
        u5_mult_82_CARRYB_50__36_), .S(u5_mult_82_SUMB_50__36_) );
  FA_X1 u5_mult_82_S2_50_33 ( .A(u5_mult_82_ab_50__33_), .B(
        u5_mult_82_CARRYB_49__33_), .CI(u5_mult_82_SUMB_49__34_), .CO(
        u5_mult_82_CARRYB_50__33_), .S(u5_mult_82_SUMB_50__33_) );
  FA_X1 u5_mult_82_S2_50_32 ( .A(u5_mult_82_ab_50__32_), .B(
        u5_mult_82_CARRYB_49__32_), .CI(u5_mult_82_SUMB_49__33_), .CO(
        u5_mult_82_CARRYB_50__32_), .S(u5_mult_82_SUMB_50__32_) );
  FA_X1 u5_mult_82_S2_50_31 ( .A(u5_mult_82_ab_50__31_), .B(
        u5_mult_82_CARRYB_49__31_), .CI(u5_mult_82_SUMB_49__32_), .CO(
        u5_mult_82_CARRYB_50__31_), .S(u5_mult_82_SUMB_50__31_) );
  FA_X1 u5_mult_82_S2_50_30 ( .A(u5_mult_82_ab_50__30_), .B(
        u5_mult_82_CARRYB_49__30_), .CI(u5_mult_82_SUMB_49__31_), .CO(
        u5_mult_82_CARRYB_50__30_), .S(u5_mult_82_SUMB_50__30_) );
  FA_X1 u5_mult_82_S2_50_29 ( .A(u5_mult_82_ab_50__29_), .B(
        u5_mult_82_CARRYB_49__29_), .CI(u5_mult_82_SUMB_49__30_), .CO(
        u5_mult_82_CARRYB_50__29_), .S(u5_mult_82_SUMB_50__29_) );
  FA_X1 u5_mult_82_S2_50_28 ( .A(u5_mult_82_CARRYB_49__28_), .B(
        u5_mult_82_ab_50__28_), .CI(u5_mult_82_SUMB_49__29_), .CO(
        u5_mult_82_CARRYB_50__28_), .S(u5_mult_82_SUMB_50__28_) );
  FA_X1 u5_mult_82_S2_50_23 ( .A(u5_mult_82_ab_50__23_), .B(
        u5_mult_82_CARRYB_49__23_), .CI(u5_mult_82_SUMB_49__24_), .CO(
        u5_mult_82_CARRYB_50__23_), .S(u5_mult_82_SUMB_50__23_) );
  FA_X1 u5_mult_82_S2_50_10 ( .A(u5_mult_82_CARRYB_49__10_), .B(
        u5_mult_82_ab_50__10_), .CI(u5_mult_82_SUMB_49__11_), .CO(
        u5_mult_82_CARRYB_50__10_), .S(u5_mult_82_SUMB_50__10_) );
  FA_X1 u5_mult_82_S2_50_1 ( .A(u5_mult_82_CARRYB_49__1_), .B(
        u5_mult_82_ab_50__1_), .CI(u5_mult_82_SUMB_49__2_), .CO(
        u5_mult_82_CARRYB_50__1_), .S(u5_mult_82_SUMB_50__1_) );
  FA_X1 u5_mult_82_S3_51_51 ( .A(u5_mult_82_ab_51__51_), .B(
        u5_mult_82_CARRYB_50__51_), .CI(u5_mult_82_ab_50__52_), .CO(
        u5_mult_82_CARRYB_51__51_), .S(u5_mult_82_SUMB_51__51_) );
  FA_X1 u5_mult_82_S2_51_50 ( .A(u5_mult_82_ab_51__50_), .B(
        u5_mult_82_CARRYB_50__50_), .CI(u5_mult_82_SUMB_50__51_), .CO(
        u5_mult_82_CARRYB_51__50_), .S(u5_mult_82_SUMB_51__50_) );
  FA_X1 u5_mult_82_S2_51_49 ( .A(u5_mult_82_ab_51__49_), .B(
        u5_mult_82_CARRYB_50__49_), .CI(u5_mult_82_SUMB_50__50_), .CO(
        u5_mult_82_CARRYB_51__49_), .S(u5_mult_82_SUMB_51__49_) );
  FA_X1 u5_mult_82_S2_51_48 ( .A(u5_mult_82_ab_51__48_), .B(
        u5_mult_82_CARRYB_50__48_), .CI(u5_mult_82_SUMB_50__49_), .CO(
        u5_mult_82_CARRYB_51__48_), .S(u5_mult_82_SUMB_51__48_) );
  FA_X1 u5_mult_82_S2_51_47 ( .A(u5_mult_82_ab_51__47_), .B(
        u5_mult_82_CARRYB_50__47_), .CI(u5_mult_82_SUMB_50__48_), .CO(
        u5_mult_82_CARRYB_51__47_), .S(u5_mult_82_SUMB_51__47_) );
  FA_X1 u5_mult_82_S2_51_46 ( .A(u5_mult_82_ab_51__46_), .B(
        u5_mult_82_CARRYB_50__46_), .CI(u5_mult_82_SUMB_50__47_), .CO(
        u5_mult_82_CARRYB_51__46_), .S(u5_mult_82_SUMB_51__46_) );
  FA_X1 u5_mult_82_S2_51_45 ( .A(u5_mult_82_ab_51__45_), .B(
        u5_mult_82_CARRYB_50__45_), .CI(u5_mult_82_SUMB_50__46_), .CO(
        u5_mult_82_CARRYB_51__45_), .S(u5_mult_82_SUMB_51__45_) );
  FA_X1 u5_mult_82_S2_51_44 ( .A(u5_mult_82_ab_51__44_), .B(
        u5_mult_82_CARRYB_50__44_), .CI(u5_mult_82_SUMB_50__45_), .CO(
        u5_mult_82_CARRYB_51__44_), .S(u5_mult_82_SUMB_51__44_) );
  FA_X1 u5_mult_82_S2_51_43 ( .A(u5_mult_82_ab_51__43_), .B(
        u5_mult_82_CARRYB_50__43_), .CI(u5_mult_82_SUMB_50__44_), .CO(
        u5_mult_82_CARRYB_51__43_), .S(u5_mult_82_SUMB_51__43_) );
  FA_X1 u5_mult_82_S2_51_42 ( .A(u5_mult_82_ab_51__42_), .B(
        u5_mult_82_CARRYB_50__42_), .CI(u5_mult_82_SUMB_50__43_), .CO(
        u5_mult_82_CARRYB_51__42_), .S(u5_mult_82_SUMB_51__42_) );
  FA_X1 u5_mult_82_S2_51_41 ( .A(u5_mult_82_ab_51__41_), .B(
        u5_mult_82_CARRYB_50__41_), .CI(u5_mult_82_SUMB_50__42_), .CO(
        u5_mult_82_CARRYB_51__41_), .S(u5_mult_82_SUMB_51__41_) );
  FA_X1 u5_mult_82_S2_51_40 ( .A(u5_mult_82_ab_51__40_), .B(
        u5_mult_82_CARRYB_50__40_), .CI(u5_mult_82_SUMB_50__41_), .CO(
        u5_mult_82_CARRYB_51__40_), .S(u5_mult_82_SUMB_51__40_) );
  FA_X1 u5_mult_82_S2_51_39 ( .A(u5_mult_82_ab_51__39_), .B(
        u5_mult_82_CARRYB_50__39_), .CI(u5_mult_82_SUMB_50__40_), .CO(
        u5_mult_82_CARRYB_51__39_), .S(u5_mult_82_SUMB_51__39_) );
  FA_X1 u5_mult_82_S2_51_38 ( .A(u5_mult_82_ab_51__38_), .B(
        u5_mult_82_CARRYB_50__38_), .CI(u5_mult_82_SUMB_50__39_), .CO(
        u5_mult_82_CARRYB_51__38_), .S(u5_mult_82_SUMB_51__38_) );
  FA_X1 u5_mult_82_S2_51_37 ( .A(u5_mult_82_ab_51__37_), .B(
        u5_mult_82_CARRYB_50__37_), .CI(u5_mult_82_SUMB_50__38_), .CO(
        u5_mult_82_CARRYB_51__37_), .S(u5_mult_82_SUMB_51__37_) );
  FA_X1 u5_mult_82_S2_51_35 ( .A(u5_mult_82_ab_51__35_), .B(
        u5_mult_82_CARRYB_50__35_), .CI(u5_mult_82_SUMB_50__36_), .CO(
        u5_mult_82_CARRYB_51__35_), .S(u5_mult_82_SUMB_51__35_) );
  FA_X1 u5_mult_82_S2_51_31 ( .A(u5_mult_82_ab_51__31_), .B(
        u5_mult_82_CARRYB_50__31_), .CI(u5_mult_82_SUMB_50__32_), .CO(
        u5_mult_82_CARRYB_51__31_), .S(u5_mult_82_SUMB_51__31_) );
  FA_X1 u5_mult_82_S2_51_30 ( .A(u5_mult_82_ab_51__30_), .B(
        u5_mult_82_CARRYB_50__30_), .CI(u5_mult_82_SUMB_50__31_), .CO(
        u5_mult_82_CARRYB_51__30_), .S(u5_mult_82_SUMB_51__30_) );
  FA_X1 u5_mult_82_S2_51_29 ( .A(u5_mult_82_ab_51__29_), .B(
        u5_mult_82_CARRYB_50__29_), .CI(u5_mult_82_SUMB_50__30_), .CO(
        u5_mult_82_CARRYB_51__29_), .S(u5_mult_82_SUMB_51__29_) );
  FA_X1 u5_mult_82_S2_51_27 ( .A(u5_mult_82_ab_51__27_), .B(
        u5_mult_82_CARRYB_50__27_), .CI(u5_mult_82_SUMB_50__28_), .CO(
        u5_mult_82_CARRYB_51__27_), .S(u5_mult_82_SUMB_51__27_) );
  FA_X1 u5_mult_82_S2_51_17 ( .A(u5_mult_82_ab_51__17_), .B(
        u5_mult_82_CARRYB_50__17_), .CI(u5_mult_82_SUMB_50__18_), .CO(
        u5_mult_82_CARRYB_51__17_), .S(u5_mult_82_SUMB_51__17_) );
  FA_X1 u5_mult_82_S2_51_16 ( .A(u5_mult_82_CARRYB_50__16_), .B(
        u5_mult_82_ab_51__16_), .CI(u5_mult_82_SUMB_50__17_), .CO(
        u5_mult_82_CARRYB_51__16_), .S(u5_mult_82_SUMB_51__16_) );
  FA_X1 u5_mult_82_S2_51_14 ( .A(u5_mult_82_ab_51__14_), .B(
        u5_mult_82_CARRYB_50__14_), .CI(u5_mult_82_SUMB_50__15_), .CO(
        u5_mult_82_CARRYB_51__14_), .S(u5_mult_82_SUMB_51__14_) );
  FA_X1 u5_mult_82_S2_51_10 ( .A(u5_mult_82_CARRYB_50__10_), .B(
        u5_mult_82_ab_51__10_), .CI(u5_mult_82_SUMB_50__11_), .CO(
        u5_mult_82_CARRYB_51__10_), .S(u5_mult_82_SUMB_51__10_) );
  FA_X1 u5_mult_82_S2_51_9 ( .A(u5_mult_82_ab_51__9_), .B(
        u5_mult_82_CARRYB_50__9_), .CI(u5_mult_82_SUMB_50__10_), .CO(
        u5_mult_82_CARRYB_51__9_), .S(u5_mult_82_SUMB_51__9_) );
  FA_X1 u5_mult_82_S2_51_2 ( .A(u5_mult_82_CARRYB_50__2_), .B(
        u5_mult_82_ab_51__2_), .CI(u5_mult_82_SUMB_50__3_), .CO(
        u5_mult_82_CARRYB_51__2_), .S(u5_mult_82_SUMB_51__2_) );
  FA_X1 u5_mult_82_S1_51_0 ( .A(u5_mult_82_CARRYB_50__0_), .B(
        u5_mult_82_ab_51__0_), .CI(u5_mult_82_SUMB_50__1_), .CO(
        u5_mult_82_CARRYB_51__0_), .S(u5_N51) );
  FA_X1 u5_mult_82_S5_51 ( .A(u5_mult_82_ab_52__51_), .B(
        u5_mult_82_CARRYB_51__51_), .CI(u5_mult_82_ab_51__52_), .CO(
        u5_mult_82_CARRYB_52__51_), .S(u5_mult_82_SUMB_52__51_) );
  FA_X1 u5_mult_82_S4_50 ( .A(u5_mult_82_ab_52__50_), .B(
        u5_mult_82_CARRYB_51__50_), .CI(u5_mult_82_SUMB_51__51_), .CO(
        u5_mult_82_CARRYB_52__50_), .S(u5_mult_82_SUMB_52__50_) );
  FA_X1 u5_mult_82_S4_49 ( .A(u5_mult_82_ab_52__49_), .B(
        u5_mult_82_CARRYB_51__49_), .CI(u5_mult_82_SUMB_51__50_), .CO(
        u5_mult_82_CARRYB_52__49_), .S(u5_mult_82_SUMB_52__49_) );
  FA_X1 u5_mult_82_S4_48 ( .A(u5_mult_82_ab_52__48_), .B(
        u5_mult_82_CARRYB_51__48_), .CI(u5_mult_82_SUMB_51__49_), .CO(
        u5_mult_82_CARRYB_52__48_), .S(u5_mult_82_SUMB_52__48_) );
  FA_X1 u5_mult_82_S4_47 ( .A(u5_mult_82_ab_52__47_), .B(
        u5_mult_82_CARRYB_51__47_), .CI(u5_mult_82_SUMB_51__48_), .CO(
        u5_mult_82_CARRYB_52__47_), .S(u5_mult_82_SUMB_52__47_) );
  FA_X1 u5_mult_82_S4_46 ( .A(u5_mult_82_ab_52__46_), .B(
        u5_mult_82_CARRYB_51__46_), .CI(u5_mult_82_SUMB_51__47_), .CO(
        u5_mult_82_CARRYB_52__46_), .S(u5_mult_82_SUMB_52__46_) );
  FA_X1 u5_mult_82_S4_45 ( .A(u5_mult_82_ab_52__45_), .B(
        u5_mult_82_CARRYB_51__45_), .CI(u5_mult_82_SUMB_51__46_), .CO(
        u5_mult_82_CARRYB_52__45_), .S(u5_mult_82_SUMB_52__45_) );
  FA_X1 u5_mult_82_S4_44 ( .A(u5_mult_82_ab_52__44_), .B(
        u5_mult_82_CARRYB_51__44_), .CI(u5_mult_82_SUMB_51__45_), .CO(
        u5_mult_82_CARRYB_52__44_), .S(u5_mult_82_SUMB_52__44_) );
  FA_X1 u5_mult_82_S4_43 ( .A(u5_mult_82_ab_52__43_), .B(
        u5_mult_82_CARRYB_51__43_), .CI(u5_mult_82_SUMB_51__44_), .CO(
        u5_mult_82_CARRYB_52__43_), .S(u5_mult_82_SUMB_52__43_) );
  FA_X1 u5_mult_82_S4_42 ( .A(u5_mult_82_ab_52__42_), .B(
        u5_mult_82_CARRYB_51__42_), .CI(u5_mult_82_SUMB_51__43_), .CO(
        u5_mult_82_CARRYB_52__42_), .S(u5_mult_82_SUMB_52__42_) );
  FA_X1 u5_mult_82_S4_41 ( .A(u5_mult_82_ab_52__41_), .B(
        u5_mult_82_CARRYB_51__41_), .CI(u5_mult_82_SUMB_51__42_), .CO(
        u5_mult_82_CARRYB_52__41_), .S(u5_mult_82_SUMB_52__41_) );
  FA_X1 u5_mult_82_S4_40 ( .A(u5_mult_82_ab_52__40_), .B(
        u5_mult_82_CARRYB_51__40_), .CI(u5_mult_82_SUMB_51__41_), .CO(
        u5_mult_82_CARRYB_52__40_), .S(u5_mult_82_SUMB_52__40_) );
  FA_X1 u5_mult_82_S4_39 ( .A(u5_mult_82_ab_52__39_), .B(
        u5_mult_82_CARRYB_51__39_), .CI(u5_mult_82_SUMB_51__40_), .CO(
        u5_mult_82_CARRYB_52__39_), .S(u5_mult_82_SUMB_52__39_) );
  FA_X1 u5_mult_82_S4_38 ( .A(u5_mult_82_ab_52__38_), .B(
        u5_mult_82_CARRYB_51__38_), .CI(u5_mult_82_SUMB_51__39_), .CO(
        u5_mult_82_CARRYB_52__38_), .S(u5_mult_82_SUMB_52__38_) );
  FA_X1 u5_mult_82_S4_37 ( .A(u5_mult_82_ab_52__37_), .B(
        u5_mult_82_CARRYB_51__37_), .CI(u5_mult_82_SUMB_51__38_), .CO(
        u5_mult_82_CARRYB_52__37_), .S(u5_mult_82_SUMB_52__37_) );
  FA_X1 u5_mult_82_S4_36 ( .A(u5_mult_82_ab_52__36_), .B(
        u5_mult_82_CARRYB_51__36_), .CI(u5_mult_82_SUMB_51__37_), .CO(
        u5_mult_82_CARRYB_52__36_), .S(u5_mult_82_SUMB_52__36_) );
  FA_X1 u5_mult_82_S4_34 ( .A(u5_mult_82_ab_52__34_), .B(
        u5_mult_82_CARRYB_51__34_), .CI(u5_mult_82_SUMB_51__35_), .CO(
        u5_mult_82_CARRYB_52__34_), .S(u5_mult_82_SUMB_52__34_) );
  FA_X1 u5_mult_82_S4_33 ( .A(u5_mult_82_ab_52__33_), .B(
        u5_mult_82_CARRYB_51__33_), .CI(u5_mult_82_SUMB_51__34_), .CO(
        u5_mult_82_CARRYB_52__33_), .S(u5_mult_82_SUMB_52__33_) );
  FA_X1 u5_mult_82_S4_30 ( .A(u5_mult_82_ab_52__30_), .B(
        u5_mult_82_CARRYB_51__30_), .CI(u5_mult_82_SUMB_51__31_), .CO(
        u5_mult_82_CARRYB_52__30_), .S(u5_mult_82_SUMB_52__30_) );
  FA_X1 u5_mult_82_S4_29 ( .A(u5_mult_82_ab_52__29_), .B(
        u5_mult_82_CARRYB_51__29_), .CI(u5_mult_82_SUMB_51__30_), .CO(
        u5_mult_82_CARRYB_52__29_), .S(u5_mult_82_SUMB_52__29_) );
  FA_X1 u5_mult_82_S4_28 ( .A(u5_mult_82_ab_52__28_), .B(
        u5_mult_82_CARRYB_51__28_), .CI(u5_mult_82_SUMB_51__29_), .CO(
        u5_mult_82_CARRYB_52__28_), .S(u5_mult_82_SUMB_52__28_) );
  FA_X1 u5_mult_82_S4_26 ( .A(u5_mult_82_ab_52__26_), .B(
        u5_mult_82_CARRYB_51__26_), .CI(u5_mult_82_SUMB_51__27_), .CO(
        u5_mult_82_CARRYB_52__26_), .S(u5_mult_82_SUMB_52__26_) );
  FA_X1 u5_mult_82_S4_25 ( .A(u5_mult_82_ab_52__25_), .B(
        u5_mult_82_CARRYB_51__25_), .CI(u5_mult_82_SUMB_51__26_), .CO(
        u5_mult_82_CARRYB_52__25_), .S(u5_mult_82_SUMB_52__25_) );
  FA_X1 u5_mult_82_S4_24 ( .A(u5_mult_82_ab_52__24_), .B(
        u5_mult_82_CARRYB_51__24_), .CI(u5_mult_82_SUMB_51__25_), .CO(
        u5_mult_82_CARRYB_52__24_), .S(u5_mult_82_SUMB_52__24_) );
  FA_X1 u5_mult_82_S4_23 ( .A(u5_mult_82_ab_52__23_), .B(
        u5_mult_82_CARRYB_51__23_), .CI(u5_mult_82_SUMB_51__24_), .CO(
        u5_mult_82_CARRYB_52__23_), .S(u5_mult_82_SUMB_52__23_) );
  FA_X1 u5_mult_82_S4_22 ( .A(u5_mult_82_ab_52__22_), .B(
        u5_mult_82_CARRYB_51__22_), .CI(u5_mult_82_SUMB_51__23_), .CO(
        u5_mult_82_CARRYB_52__22_), .S(u5_mult_82_SUMB_52__22_) );
  FA_X1 u5_mult_82_S4_18 ( .A(u5_mult_82_ab_52__18_), .B(
        u5_mult_82_CARRYB_51__18_), .CI(u5_mult_82_SUMB_51__19_), .CO(
        u5_mult_82_CARRYB_52__18_), .S(u5_mult_82_SUMB_52__18_) );
  FA_X1 u5_mult_82_S4_17 ( .A(u5_mult_82_SUMB_51__18_), .B(
        u5_mult_82_CARRYB_51__17_), .CI(u5_mult_82_ab_52__17_), .CO(
        u5_mult_82_CARRYB_52__17_), .S(u5_mult_82_SUMB_52__17_) );
  FA_X1 u5_mult_82_S4_16 ( .A(u5_mult_82_ab_52__16_), .B(
        u5_mult_82_CARRYB_51__16_), .CI(u5_mult_82_SUMB_51__17_), .CO(
        u5_mult_82_CARRYB_52__16_), .S(u5_mult_82_SUMB_52__16_) );
  FA_X1 u5_mult_82_S4_14 ( .A(u5_mult_82_ab_52__14_), .B(
        u5_mult_82_CARRYB_51__14_), .CI(u5_mult_82_SUMB_51__15_), .CO(
        u5_mult_82_CARRYB_52__14_), .S(u5_mult_82_SUMB_52__14_) );
  FA_X1 u5_mult_82_S4_13 ( .A(u5_mult_82_ab_52__13_), .B(
        u5_mult_82_CARRYB_51__13_), .CI(u5_mult_82_SUMB_51__14_), .CO(
        u5_mult_82_CARRYB_52__13_), .S(u5_mult_82_SUMB_52__13_) );
  FA_X1 u5_mult_82_S4_10 ( .A(u5_mult_82_ab_52__10_), .B(
        u5_mult_82_CARRYB_51__10_), .CI(u5_mult_82_SUMB_51__11_), .CO(
        u5_mult_82_CARRYB_52__10_), .S(u5_mult_82_SUMB_52__10_) );
  FA_X1 u5_mult_82_S4_9 ( .A(u5_mult_82_ab_52__9_), .B(
        u5_mult_82_CARRYB_51__9_), .CI(u5_mult_82_SUMB_51__10_), .CO(
        u5_mult_82_CARRYB_52__9_), .S(u5_mult_82_SUMB_52__9_) );
  FA_X1 u5_mult_82_S4_7 ( .A(u5_mult_82_ab_52__7_), .B(
        u5_mult_82_CARRYB_51__7_), .CI(u5_mult_82_SUMB_51__8_), .CO(
        u5_mult_82_CARRYB_52__7_), .S(u5_mult_82_SUMB_52__7_) );
  FA_X1 u5_mult_82_S4_6 ( .A(u5_mult_82_ab_52__6_), .B(
        u5_mult_82_CARRYB_51__6_), .CI(u5_mult_82_SUMB_51__7_), .CO(
        u5_mult_82_CARRYB_52__6_), .S(u5_mult_82_SUMB_52__6_) );
  FA_X1 u5_mult_82_S4_3 ( .A(u5_mult_82_ab_52__3_), .B(
        u5_mult_82_CARRYB_51__3_), .CI(u5_mult_82_SUMB_51__4_), .CO(
        u5_mult_82_CARRYB_52__3_), .S(u5_mult_82_SUMB_52__3_) );
  FA_X1 u5_mult_82_S4_2 ( .A(u5_mult_82_SUMB_51__3_), .B(u5_mult_82_ab_52__2_), 
        .CI(u5_mult_82_CARRYB_51__2_), .CO(u5_mult_82_CARRYB_52__2_), .S(
        u5_mult_82_SUMB_52__2_) );
  FA_X1 u5_mult_82_S4_1 ( .A(u5_mult_82_CARRYB_51__1_), .B(
        u5_mult_82_ab_52__1_), .CI(u5_mult_82_SUMB_51__2_), .CO(
        u5_mult_82_CARRYB_52__1_), .S(u5_mult_82_SUMB_52__1_) );
  FA_X1 u5_mult_82_S4_0 ( .A(u5_mult_82_CARRYB_51__0_), .B(
        u5_mult_82_ab_52__0_), .CI(u5_mult_82_SUMB_51__1_), .CO(
        u5_mult_82_CARRYB_52__0_), .S(u5_N52) );
  NAND2_X2 u5_mult_82_FS_1_U796 ( .A1(u5_mult_82_n622), .A2(
        u5_mult_82_CLA_SUM[102]), .ZN(u5_mult_82_FS_1_n543) );
  INV_X4 u5_mult_82_FS_1_U795 ( .A(u5_mult_82_n622), .ZN(u5_mult_82_FS_1_n742)
         );
  INV_X4 u5_mult_82_FS_1_U794 ( .A(u5_mult_82_CLA_SUM[102]), .ZN(
        u5_mult_82_FS_1_n743) );
  NAND2_X2 u5_mult_82_FS_1_U793 ( .A1(u5_mult_82_FS_1_n742), .A2(
        u5_mult_82_FS_1_n743), .ZN(u5_mult_82_FS_1_n542) );
  NAND2_X2 u5_mult_82_FS_1_U792 ( .A1(u5_mult_82_FS_1_n543), .A2(
        u5_mult_82_FS_1_n542), .ZN(u5_mult_82_FS_1_n551) );
  INV_X4 u5_mult_82_FS_1_U791 ( .A(u5_mult_82_n621), .ZN(u5_mult_82_FS_1_n740)
         );
  INV_X4 u5_mult_82_FS_1_U790 ( .A(u5_mult_82_CLA_SUM[98]), .ZN(
        u5_mult_82_FS_1_n741) );
  NAND2_X2 u5_mult_82_FS_1_U789 ( .A1(u5_mult_82_FS_1_n740), .A2(
        u5_mult_82_FS_1_n741), .ZN(u5_mult_82_FS_1_n101) );
  INV_X4 u5_mult_82_FS_1_U788 ( .A(u5_mult_82_FS_1_n101), .ZN(
        u5_mult_82_FS_1_n97) );
  INV_X4 u5_mult_82_FS_1_U787 ( .A(u5_mult_82_n619), .ZN(u5_mult_82_FS_1_n738)
         );
  INV_X4 u5_mult_82_FS_1_U786 ( .A(u5_mult_82_CLA_SUM[100]), .ZN(
        u5_mult_82_FS_1_n739) );
  NAND2_X2 u5_mult_82_FS_1_U785 ( .A1(u5_mult_82_FS_1_n738), .A2(
        u5_mult_82_FS_1_n739), .ZN(u5_mult_82_FS_1_n74) );
  INV_X4 u5_mult_82_FS_1_U784 ( .A(u5_mult_82_FS_1_n74), .ZN(
        u5_mult_82_FS_1_n625) );
  INV_X4 u5_mult_82_FS_1_U783 ( .A(u5_mult_82_n620), .ZN(u5_mult_82_FS_1_n736)
         );
  INV_X4 u5_mult_82_FS_1_U782 ( .A(u5_mult_82_CLA_SUM[99]), .ZN(
        u5_mult_82_FS_1_n737) );
  NAND2_X2 u5_mult_82_FS_1_U781 ( .A1(u5_mult_82_FS_1_n736), .A2(
        u5_mult_82_FS_1_n737), .ZN(u5_mult_82_FS_1_n91) );
  INV_X4 u5_mult_82_FS_1_U780 ( .A(u5_mult_82_FS_1_n91), .ZN(
        u5_mult_82_FS_1_n626) );
  NOR3_X4 u5_mult_82_FS_1_U779 ( .A1(u5_mult_82_FS_1_n97), .A2(
        u5_mult_82_FS_1_n625), .A3(u5_mult_82_FS_1_n626), .ZN(
        u5_mult_82_FS_1_n592) );
  INV_X4 u5_mult_82_FS_1_U778 ( .A(u5_mult_82_CLA_SUM[101]), .ZN(
        u5_mult_82_FS_1_n734) );
  INV_X4 u5_mult_82_FS_1_U777 ( .A(u5_mult_82_n618), .ZN(u5_mult_82_FS_1_n735)
         );
  NAND2_X2 u5_mult_82_FS_1_U776 ( .A1(u5_mult_82_FS_1_n734), .A2(
        u5_mult_82_FS_1_n735), .ZN(u5_mult_82_FS_1_n85) );
  INV_X4 u5_mult_82_FS_1_U775 ( .A(u5_mult_82_n607), .ZN(u5_mult_82_FS_1_n732)
         );
  INV_X4 u5_mult_82_FS_1_U774 ( .A(u5_mult_82_n606), .ZN(u5_mult_82_FS_1_n730)
         );
  INV_X4 u5_mult_82_FS_1_U773 ( .A(u5_mult_82_CLA_SUM[89]), .ZN(
        u5_mult_82_FS_1_n731) );
  INV_X4 u5_mult_82_FS_1_U772 ( .A(u5_mult_82_n590), .ZN(u5_mult_82_FS_1_n728)
         );
  INV_X4 u5_mult_82_FS_1_U771 ( .A(u5_mult_82_CLA_SUM[87]), .ZN(
        u5_mult_82_FS_1_n729) );
  INV_X4 u5_mult_82_FS_1_U770 ( .A(u5_mult_82_FS_1_n232), .ZN(
        u5_mult_82_FS_1_n724) );
  INV_X4 u5_mult_82_FS_1_U769 ( .A(u5_mult_82_n605), .ZN(u5_mult_82_FS_1_n726)
         );
  INV_X4 u5_mult_82_FS_1_U768 ( .A(u5_mult_82_CLA_SUM[88]), .ZN(
        u5_mult_82_FS_1_n727) );
  INV_X4 u5_mult_82_FS_1_U767 ( .A(u5_mult_82_FS_1_n216), .ZN(
        u5_mult_82_FS_1_n725) );
  NOR2_X4 u5_mult_82_FS_1_U766 ( .A1(u5_mult_82_FS_1_n724), .A2(
        u5_mult_82_FS_1_n725), .ZN(u5_mult_82_FS_1_n723) );
  NAND3_X4 u5_mult_82_FS_1_U765 ( .A1(u5_mult_82_FS_1_n723), .A2(
        u5_mult_82_FS_1_n202), .A3(u5_mult_82_FS_1_n240), .ZN(
        u5_mult_82_FS_1_n205) );
  INV_X4 u5_mult_82_FS_1_U764 ( .A(u5_mult_82_n593), .ZN(u5_mult_82_FS_1_n721)
         );
  INV_X4 u5_mult_82_FS_1_U763 ( .A(u5_mult_82_CLA_SUM[84]), .ZN(
        u5_mult_82_FS_1_n722) );
  INV_X4 u5_mult_82_FS_1_U762 ( .A(u5_mult_82_FS_1_n270), .ZN(
        u5_mult_82_FS_1_n717) );
  INV_X4 u5_mult_82_FS_1_U761 ( .A(u5_mult_82_n597), .ZN(u5_mult_82_FS_1_n719)
         );
  INV_X4 u5_mult_82_FS_1_U760 ( .A(u5_mult_82_CLA_SUM[85]), .ZN(
        u5_mult_82_FS_1_n720) );
  NOR2_X4 u5_mult_82_FS_1_U759 ( .A1(u5_mult_82_FS_1_n606), .A2(
        u5_mult_82_FS_1_n271), .ZN(u5_mult_82_FS_1_n718) );
  NAND3_X4 u5_mult_82_FS_1_U758 ( .A1(u5_mult_82_FS_1_n250), .A2(
        u5_mult_82_FS_1_n717), .A3(u5_mult_82_FS_1_n718), .ZN(
        u5_mult_82_FS_1_n241) );
  INV_X4 u5_mult_82_FS_1_U757 ( .A(u5_mult_82_n601), .ZN(u5_mult_82_FS_1_n715)
         );
  INV_X4 u5_mult_82_FS_1_U756 ( .A(u5_mult_82_CLA_SUM[94]), .ZN(
        u5_mult_82_FS_1_n716) );
  INV_X4 u5_mult_82_FS_1_U755 ( .A(u5_mult_82_n600), .ZN(u5_mult_82_FS_1_n713)
         );
  INV_X4 u5_mult_82_FS_1_U754 ( .A(u5_mult_82_CLA_SUM[95]), .ZN(
        u5_mult_82_FS_1_n714) );
  NAND2_X2 u5_mult_82_FS_1_U753 ( .A1(u5_mult_82_FS_1_n713), .A2(
        u5_mult_82_FS_1_n714), .ZN(u5_mult_82_FS_1_n144) );
  INV_X4 u5_mult_82_FS_1_U752 ( .A(u5_mult_82_n617), .ZN(u5_mult_82_FS_1_n711)
         );
  INV_X4 u5_mult_82_FS_1_U751 ( .A(u5_mult_82_CLA_SUM[97]), .ZN(
        u5_mult_82_FS_1_n712) );
  NAND2_X2 u5_mult_82_FS_1_U750 ( .A1(u5_mult_82_FS_1_n711), .A2(
        u5_mult_82_FS_1_n712), .ZN(u5_mult_82_FS_1_n710) );
  INV_X4 u5_mult_82_FS_1_U749 ( .A(u5_mult_82_FS_1_n710), .ZN(
        u5_mult_82_FS_1_n109) );
  INV_X4 u5_mult_82_FS_1_U748 ( .A(u5_mult_82_n580), .ZN(u5_mult_82_FS_1_n708)
         );
  INV_X4 u5_mult_82_FS_1_U747 ( .A(u5_mult_82_CLA_SUM[96]), .ZN(
        u5_mult_82_FS_1_n709) );
  NAND2_X2 u5_mult_82_FS_1_U746 ( .A1(u5_mult_82_FS_1_n708), .A2(
        u5_mult_82_FS_1_n709), .ZN(u5_mult_82_FS_1_n153) );
  INV_X4 u5_mult_82_FS_1_U745 ( .A(u5_mult_82_FS_1_n153), .ZN(
        u5_mult_82_FS_1_n131) );
  NOR2_X4 u5_mult_82_FS_1_U744 ( .A1(u5_mult_82_FS_1_n109), .A2(
        u5_mult_82_FS_1_n131), .ZN(u5_mult_82_FS_1_n707) );
  NAND3_X4 u5_mult_82_FS_1_U743 ( .A1(u5_mult_82_FS_1_n143), .A2(
        u5_mult_82_FS_1_n144), .A3(u5_mult_82_FS_1_n707), .ZN(
        u5_mult_82_FS_1_n607) );
  INV_X4 u5_mult_82_FS_1_U742 ( .A(u5_mult_82_n604), .ZN(u5_mult_82_FS_1_n705)
         );
  INV_X4 u5_mult_82_FS_1_U741 ( .A(u5_mult_82_CLA_SUM[90]), .ZN(
        u5_mult_82_FS_1_n706) );
  NAND2_X2 u5_mult_82_FS_1_U740 ( .A1(u5_mult_82_FS_1_n705), .A2(
        u5_mult_82_FS_1_n706), .ZN(u5_mult_82_FS_1_n198) );
  INV_X4 u5_mult_82_FS_1_U739 ( .A(u5_mult_82_n602), .ZN(u5_mult_82_FS_1_n703)
         );
  INV_X4 u5_mult_82_FS_1_U738 ( .A(u5_mult_82_CLA_SUM[93]), .ZN(
        u5_mult_82_FS_1_n704) );
  NAND2_X2 u5_mult_82_FS_1_U737 ( .A1(u5_mult_82_FS_1_n703), .A2(
        u5_mult_82_FS_1_n704), .ZN(u5_mult_82_FS_1_n170) );
  INV_X4 u5_mult_82_FS_1_U736 ( .A(u5_mult_82_n603), .ZN(u5_mult_82_FS_1_n701)
         );
  INV_X4 u5_mult_82_FS_1_U735 ( .A(u5_mult_82_CLA_SUM[91]), .ZN(
        u5_mult_82_FS_1_n702) );
  INV_X4 u5_mult_82_FS_1_U734 ( .A(u5_mult_82_FS_1_n191), .ZN(
        u5_mult_82_FS_1_n188) );
  NAND3_X4 u5_mult_82_FS_1_U733 ( .A1(u5_mult_82_FS_1_n198), .A2(
        u5_mult_82_FS_1_n170), .A3(u5_mult_82_FS_1_n613), .ZN(
        u5_mult_82_FS_1_n165) );
  NOR2_X4 u5_mult_82_FS_1_U732 ( .A1(u5_mult_82_FS_1_n607), .A2(
        u5_mult_82_FS_1_n165), .ZN(u5_mult_82_FS_1_n700) );
  INV_X4 u5_mult_82_FS_1_U731 ( .A(u5_mult_82_n485), .ZN(u5_mult_82_FS_1_n697)
         );
  INV_X4 u5_mult_82_FS_1_U730 ( .A(u5_mult_82_CLA_SUM[80]), .ZN(
        u5_mult_82_FS_1_n698) );
  INV_X4 u5_mult_82_FS_1_U729 ( .A(u5_mult_82_n486), .ZN(u5_mult_82_FS_1_n695)
         );
  INV_X4 u5_mult_82_FS_1_U728 ( .A(u5_mult_82_CLA_SUM[81]), .ZN(
        u5_mult_82_FS_1_n696) );
  NAND2_X2 u5_mult_82_FS_1_U727 ( .A1(u5_mult_82_FS_1_n695), .A2(
        u5_mult_82_FS_1_n696), .ZN(u5_mult_82_FS_1_n305) );
  INV_X4 u5_mult_82_FS_1_U726 ( .A(u5_mult_82_n587), .ZN(u5_mult_82_FS_1_n693)
         );
  INV_X4 u5_mult_82_FS_1_U725 ( .A(u5_mult_82_CLA_SUM[79]), .ZN(
        u5_mult_82_FS_1_n694) );
  NOR2_X4 u5_mult_82_FS_1_U724 ( .A1(u5_mult_82_FS_1_n14), .A2(
        u5_mult_82_FS_1_n316), .ZN(u5_mult_82_FS_1_n311) );
  NOR2_X4 u5_mult_82_FS_1_U723 ( .A1(u5_mult_82_CLA_SUM[68]), .A2(
        u5_mult_82_n578), .ZN(u5_mult_82_FS_1_n426) );
  NOR2_X4 u5_mult_82_FS_1_U722 ( .A1(u5_mult_82_CLA_SUM[67]), .A2(
        u5_mult_82_CLA_CARRY[66]), .ZN(u5_mult_82_FS_1_n429) );
  INV_X4 u5_mult_82_FS_1_U721 ( .A(u5_mult_82_FS_1_n429), .ZN(
        u5_mult_82_FS_1_n689) );
  INV_X4 u5_mult_82_FS_1_U720 ( .A(u5_mult_82_n608), .ZN(u5_mult_82_FS_1_n691)
         );
  INV_X4 u5_mult_82_FS_1_U719 ( .A(u5_mult_82_n5565), .ZN(u5_mult_82_FS_1_n692) );
  NOR2_X4 u5_mult_82_FS_1_U718 ( .A1(u5_mult_82_CLA_SUM[66]), .A2(
        u5_mult_82_n581), .ZN(u5_mult_82_FS_1_n430) );
  NOR2_X4 u5_mult_82_FS_1_U717 ( .A1(u5_mult_82_FS_1_n409), .A2(
        u5_mult_82_FS_1_n430), .ZN(u5_mult_82_FS_1_n690) );
  NOR2_X4 u5_mult_82_FS_1_U716 ( .A1(u5_mult_82_FS_1_n389), .A2(
        u5_mult_82_FS_1_n563), .ZN(u5_mult_82_FS_1_n671) );
  INV_X4 u5_mult_82_FS_1_U715 ( .A(u5_mult_82_n584), .ZN(u5_mult_82_FS_1_n687)
         );
  INV_X4 u5_mult_82_FS_1_U714 ( .A(u5_mult_82_CLA_SUM[74]), .ZN(
        u5_mult_82_FS_1_n688) );
  INV_X4 u5_mult_82_FS_1_U713 ( .A(u5_mult_82_n582), .ZN(u5_mult_82_FS_1_n685)
         );
  INV_X4 u5_mult_82_FS_1_U712 ( .A(u5_mult_82_CLA_SUM[77]), .ZN(
        u5_mult_82_FS_1_n686) );
  INV_X4 u5_mult_82_FS_1_U711 ( .A(u5_mult_82_n595), .ZN(u5_mult_82_FS_1_n683)
         );
  INV_X4 u5_mult_82_FS_1_U710 ( .A(u5_mult_82_n591), .ZN(u5_mult_82_FS_1_n681)
         );
  NOR2_X4 u5_mult_82_FS_1_U709 ( .A1(u5_mult_82_FS_1_n343), .A2(
        u5_mult_82_FS_1_n342), .ZN(u5_mult_82_FS_1_n679) );
  NAND3_X4 u5_mult_82_FS_1_U708 ( .A1(u5_mult_82_FS_1_n363), .A2(
        u5_mult_82_FS_1_n349), .A3(u5_mult_82_FS_1_n679), .ZN(
        u5_mult_82_FS_1_n572) );
  INV_X4 u5_mult_82_FS_1_U707 ( .A(u5_mult_82_CLA_CARRY[71]), .ZN(
        u5_mult_82_FS_1_n677) );
  NOR2_X4 u5_mult_82_FS_1_U706 ( .A1(u5_mult_82_CLA_SUM[71]), .A2(
        u5_mult_82_n574), .ZN(u5_mult_82_FS_1_n384) );
  INV_X4 u5_mult_82_FS_1_U705 ( .A(u5_mult_82_n484), .ZN(u5_mult_82_FS_1_n675)
         );
  INV_X4 u5_mult_82_FS_1_U704 ( .A(u5_mult_82_FS_1_n369), .ZN(
        u5_mult_82_FS_1_n674) );
  NOR2_X4 u5_mult_82_FS_1_U703 ( .A1(u5_mult_82_CLA_SUM[70]), .A2(
        u5_mult_82_n577), .ZN(u5_mult_82_FS_1_n390) );
  NOR2_X4 u5_mult_82_FS_1_U702 ( .A1(u5_mult_82_FS_1_n674), .A2(
        u5_mult_82_FS_1_n390), .ZN(u5_mult_82_FS_1_n673) );
  INV_X4 u5_mult_82_FS_1_U701 ( .A(u5_mult_82_n588), .ZN(u5_mult_82_FS_1_n669)
         );
  INV_X4 u5_mult_82_FS_1_U700 ( .A(u5_mult_82_n592), .ZN(u5_mult_82_FS_1_n667)
         );
  NOR2_X4 u5_mult_82_FS_1_U699 ( .A1(u5_mult_82_FS_1_n19), .A2(
        u5_mult_82_FS_1_n34), .ZN(u5_mult_82_FS_1_n666) );
  NOR2_X4 u5_mult_82_FS_1_U698 ( .A1(u5_mult_82_CLA_SUM[58]), .A2(
        u5_mult_82_n575), .ZN(u5_mult_82_FS_1_n487) );
  NOR2_X4 u5_mult_82_FS_1_U697 ( .A1(u5_mult_82_CLA_SUM[55]), .A2(
        u5_mult_82_n1604), .ZN(u5_mult_82_FS_1_n499) );
  NOR2_X4 u5_mult_82_FS_1_U696 ( .A1(u5_mult_82_FS_1_n50), .A2(u5_mult_82_n573), .ZN(u5_mult_82_FS_1_n483) );
  NOR2_X4 u5_mult_82_FS_1_U695 ( .A1(u5_mult_82_CLA_SUM[60]), .A2(
        u5_mult_82_n576), .ZN(u5_mult_82_FS_1_n474) );
  INV_X4 u5_mult_82_FS_1_U694 ( .A(u5_mult_82_n594), .ZN(u5_mult_82_FS_1_n662)
         );
  INV_X4 u5_mult_82_FS_1_U693 ( .A(u5_mult_82_CLA_SUM[61]), .ZN(
        u5_mult_82_FS_1_n663) );
  NOR2_X4 u5_mult_82_FS_1_U692 ( .A1(u5_mult_82_FS_1_n474), .A2(
        u5_mult_82_FS_1_n470), .ZN(u5_mult_82_FS_1_n661) );
  NOR2_X4 u5_mult_82_FS_1_U691 ( .A1(u5_mult_82_FS_1_n658), .A2(
        u5_mult_82_FS_1_n659), .ZN(u5_mult_82_FS_1_n655) );
  INV_X4 u5_mult_82_FS_1_U690 ( .A(u5_mult_82_n598), .ZN(u5_mult_82_FS_1_n656)
         );
  INV_X4 u5_mult_82_FS_1_U689 ( .A(u5_mult_82_CLA_SUM[57]), .ZN(
        u5_mult_82_FS_1_n657) );
  NOR2_X4 u5_mult_82_FS_1_U688 ( .A1(u5_mult_82_FS_1_n506), .A2(
        u5_mult_82_FS_1_n644), .ZN(u5_mult_82_FS_1_n494) );
  NAND3_X4 u5_mult_82_FS_1_U687 ( .A1(u5_mult_82_FS_1_n655), .A2(
        u5_mult_82_FS_1_n281), .A3(u5_mult_82_FS_1_n494), .ZN(
        u5_mult_82_FS_1_n222) );
  INV_X4 u5_mult_82_FS_1_U686 ( .A(u5_mult_82_FS_1_n651), .ZN(
        u5_mult_82_FS_1_n645) );
  NOR2_X4 u5_mult_82_FS_1_U685 ( .A1(u5_mult_82_CLA_SUM[58]), .A2(
        u5_mult_82_n575), .ZN(u5_mult_82_FS_1_n648) );
  INV_X4 u5_mult_82_FS_1_U684 ( .A(u5_mult_82_FS_1_n654), .ZN(
        u5_mult_82_FS_1_n653) );
  NAND3_X4 u5_mult_82_FS_1_U683 ( .A1(u5_mult_82_FS_1_n281), .A2(
        u5_mult_82_FS_1_n652), .A3(u5_mult_82_FS_1_n645), .ZN(
        u5_mult_82_FS_1_n221) );
  NAND2_X2 u5_mult_82_FS_1_U682 ( .A1(u5_mult_82_n598), .A2(
        u5_mult_82_CLA_SUM[57]), .ZN(u5_mult_82_FS_1_n501) );
  NAND3_X4 u5_mult_82_FS_1_U681 ( .A1(u5_mult_82_FS_1_n281), .A2(
        u5_mult_82_FS_1_n650), .A3(u5_mult_82_FS_1_n649), .ZN(
        u5_mult_82_FS_1_n223) );
  OAI21_X4 u5_mult_82_FS_1_U680 ( .B1(u5_mult_82_FS_1_n640), .B2(
        u5_mult_82_FS_1_n641), .A(u5_mult_82_FS_1_n642), .ZN(
        u5_mult_82_FS_1_n122) );
  NAND2_X2 u5_mult_82_FS_1_U679 ( .A1(u5_mult_82_n576), .A2(
        u5_mult_82_CLA_SUM[60]), .ZN(u5_mult_82_FS_1_n475) );
  INV_X4 u5_mult_82_FS_1_U678 ( .A(u5_mult_82_CLA_SUM[58]), .ZN(
        u5_mult_82_FS_1_n638) );
  INV_X4 u5_mult_82_FS_1_U677 ( .A(u5_mult_82_n575), .ZN(u5_mult_82_FS_1_n639)
         );
  NOR2_X4 u5_mult_82_FS_1_U676 ( .A1(u5_mult_82_FS_1_n638), .A2(
        u5_mult_82_FS_1_n639), .ZN(u5_mult_82_FS_1_n634) );
  NOR2_X4 u5_mult_82_FS_1_U675 ( .A1(u5_mult_82_FS_1_n636), .A2(
        u5_mult_82_FS_1_n637), .ZN(u5_mult_82_FS_1_n635) );
  NAND3_X4 u5_mult_82_FS_1_U674 ( .A1(u5_mult_82_FS_1_n281), .A2(
        u5_mult_82_FS_1_n477), .A3(u5_mult_82_FS_1_n15), .ZN(
        u5_mult_82_FS_1_n218) );
  NAND2_X2 u5_mult_82_FS_1_U673 ( .A1(u5_mult_82_n621), .A2(
        u5_mult_82_CLA_SUM[98]), .ZN(u5_mult_82_FS_1_n99) );
  NAND2_X2 u5_mult_82_FS_1_U672 ( .A1(u5_mult_82_n620), .A2(
        u5_mult_82_CLA_SUM[99]), .ZN(u5_mult_82_FS_1_n76) );
  NAND2_X2 u5_mult_82_FS_1_U671 ( .A1(u5_mult_82_FS_1_n99), .A2(
        u5_mult_82_FS_1_n76), .ZN(u5_mult_82_FS_1_n623) );
  NAND2_X2 u5_mult_82_FS_1_U670 ( .A1(u5_mult_82_n619), .A2(
        u5_mult_82_CLA_SUM[100]), .ZN(u5_mult_82_FS_1_n72) );
  NAND2_X2 u5_mult_82_FS_1_U669 ( .A1(u5_mult_82_n618), .A2(
        u5_mult_82_CLA_SUM[101]), .ZN(u5_mult_82_FS_1_n86) );
  NAND2_X2 u5_mult_82_FS_1_U668 ( .A1(u5_mult_82_FS_1_n72), .A2(
        u5_mult_82_FS_1_n86), .ZN(u5_mult_82_FS_1_n624) );
  INV_X4 u5_mult_82_FS_1_U667 ( .A(u5_mult_82_FS_1_n202), .ZN(
        u5_mult_82_FS_1_n621) );
  NOR3_X4 u5_mult_82_FS_1_U666 ( .A1(u5_mult_82_FS_1_n621), .A2(
        u5_mult_82_FS_1_n607), .A3(u5_mult_82_FS_1_n165), .ZN(
        u5_mult_82_FS_1_n608) );
  NAND2_X2 u5_mult_82_FS_1_U665 ( .A1(u5_mult_82_n607), .A2(u5_mult_82_n1075), 
        .ZN(u5_mult_82_FS_1_n239) );
  NAND2_X2 u5_mult_82_FS_1_U664 ( .A1(u5_mult_82_FS_1_n239), .A2(
        u5_mult_82_FS_1_n225), .ZN(u5_mult_82_FS_1_n620) );
  INV_X4 u5_mult_82_FS_1_U663 ( .A(u5_mult_82_FS_1_n620), .ZN(
        u5_mult_82_FS_1_n615) );
  NAND2_X2 u5_mult_82_FS_1_U662 ( .A1(u5_mult_82_n605), .A2(
        u5_mult_82_CLA_SUM[88]), .ZN(u5_mult_82_FS_1_n213) );
  INV_X4 u5_mult_82_FS_1_U661 ( .A(u5_mult_82_FS_1_n213), .ZN(
        u5_mult_82_FS_1_n618) );
  NAND2_X2 u5_mult_82_FS_1_U660 ( .A1(u5_mult_82_n606), .A2(
        u5_mult_82_CLA_SUM[89]), .ZN(u5_mult_82_FS_1_n210) );
  INV_X4 u5_mult_82_FS_1_U659 ( .A(u5_mult_82_FS_1_n210), .ZN(
        u5_mult_82_FS_1_n619) );
  NOR2_X4 u5_mult_82_FS_1_U658 ( .A1(u5_mult_82_FS_1_n618), .A2(
        u5_mult_82_FS_1_n619), .ZN(u5_mult_82_FS_1_n617) );
  NAND2_X2 u5_mult_82_FS_1_U657 ( .A1(u5_mult_82_n603), .A2(
        u5_mult_82_CLA_SUM[91]), .ZN(u5_mult_82_FS_1_n182) );
  NAND2_X2 u5_mult_82_FS_1_U656 ( .A1(u5_mult_82_FS_1_n197), .A2(
        u5_mult_82_FS_1_n182), .ZN(u5_mult_82_FS_1_n614) );
  NAND2_X2 u5_mult_82_FS_1_U655 ( .A1(u5_mult_82_FS_1_n614), .A2(
        u5_mult_82_FS_1_n613), .ZN(u5_mult_82_FS_1_n612) );
  INV_X4 u5_mult_82_FS_1_U654 ( .A(u5_mult_82_FS_1_n612), .ZN(
        u5_mult_82_FS_1_n610) );
  NAND2_X2 u5_mult_82_FS_1_U653 ( .A1(u5_mult_82_n602), .A2(
        u5_mult_82_CLA_SUM[93]), .ZN(u5_mult_82_FS_1_n171) );
  NAND2_X2 u5_mult_82_FS_1_U652 ( .A1(u5_mult_82_n596), .A2(
        u5_mult_82_CLA_SUM[92]), .ZN(u5_mult_82_FS_1_n174) );
  NAND2_X2 u5_mult_82_FS_1_U651 ( .A1(u5_mult_82_FS_1_n171), .A2(
        u5_mult_82_FS_1_n174), .ZN(u5_mult_82_FS_1_n611) );
  OAI21_X4 u5_mult_82_FS_1_U650 ( .B1(u5_mult_82_FS_1_n610), .B2(
        u5_mult_82_FS_1_n611), .A(u5_mult_82_FS_1_n170), .ZN(
        u5_mult_82_FS_1_n166) );
  AOI21_X4 u5_mult_82_FS_1_U649 ( .B1(u5_mult_82_FS_1_n608), .B2(
        u5_mult_82_FS_1_n203), .A(u5_mult_82_FS_1_n609), .ZN(
        u5_mult_82_FS_1_n593) );
  INV_X4 u5_mult_82_FS_1_U648 ( .A(u5_mult_82_FS_1_n607), .ZN(
        u5_mult_82_FS_1_n598) );
  INV_X4 u5_mult_82_FS_1_U647 ( .A(u5_mult_82_FS_1_n165), .ZN(
        u5_mult_82_FS_1_n599) );
  NAND2_X2 u5_mult_82_FS_1_U646 ( .A1(u5_mult_82_n593), .A2(
        u5_mult_82_CLA_SUM[84]), .ZN(u5_mult_82_FS_1_n254) );
  NAND2_X2 u5_mult_82_FS_1_U645 ( .A1(u5_mult_82_n597), .A2(
        u5_mult_82_CLA_SUM[85]), .ZN(u5_mult_82_FS_1_n261) );
  INV_X4 u5_mult_82_FS_1_U644 ( .A(u5_mult_82_FS_1_n261), .ZN(
        u5_mult_82_FS_1_n603) );
  AOI21_X4 u5_mult_82_FS_1_U643 ( .B1(u5_mult_82_FS_1_n601), .B2(
        u5_mult_82_FS_1_n602), .A(u5_mult_82_FS_1_n603), .ZN(
        u5_mult_82_FS_1_n600) );
  NAND2_X2 u5_mult_82_FS_1_U642 ( .A1(u5_mult_82_n580), .A2(
        u5_mult_82_CLA_SUM[96]), .ZN(u5_mult_82_FS_1_n113) );
  INV_X4 u5_mult_82_FS_1_U641 ( .A(u5_mult_82_FS_1_n113), .ZN(
        u5_mult_82_FS_1_n596) );
  INV_X4 u5_mult_82_FS_1_U640 ( .A(u5_mult_82_FS_1_n144), .ZN(
        u5_mult_82_FS_1_n141) );
  NAND2_X2 u5_mult_82_FS_1_U639 ( .A1(u5_mult_82_n601), .A2(
        u5_mult_82_CLA_SUM[94]), .ZN(u5_mult_82_FS_1_n142) );
  NAND2_X2 u5_mult_82_FS_1_U638 ( .A1(u5_mult_82_n600), .A2(
        u5_mult_82_CLA_SUM[95]), .ZN(u5_mult_82_FS_1_n128) );
  OAI21_X4 u5_mult_82_FS_1_U637 ( .B1(u5_mult_82_FS_1_n141), .B2(
        u5_mult_82_FS_1_n142), .A(u5_mult_82_FS_1_n128), .ZN(
        u5_mult_82_FS_1_n597) );
  OAI21_X4 u5_mult_82_FS_1_U636 ( .B1(u5_mult_82_FS_1_n596), .B2(
        u5_mult_82_FS_1_n597), .A(u5_mult_82_FS_1_n707), .ZN(
        u5_mult_82_FS_1_n595) );
  NAND2_X2 u5_mult_82_FS_1_U635 ( .A1(u5_mult_82_n617), .A2(
        u5_mult_82_CLA_SUM[97]), .ZN(u5_mult_82_FS_1_n110) );
  INV_X4 u5_mult_82_FS_1_U634 ( .A(u5_mult_82_FS_1_n85), .ZN(
        u5_mult_82_FS_1_n591) );
  AOI21_X4 u5_mult_82_FS_1_U633 ( .B1(u5_mult_82_FS_1_n589), .B2(
        u5_mult_82_FS_1_n590), .A(u5_mult_82_FS_1_n591), .ZN(
        u5_mult_82_FS_1_n588) );
  NOR2_X4 u5_mult_82_FS_1_U632 ( .A1(u5_mult_82_FS_1_n579), .A2(
        u5_mult_82_FS_1_n580), .ZN(u5_mult_82_FS_1_n366) );
  NAND2_X2 u5_mult_82_FS_1_U631 ( .A1(u5_mult_82_CLA_CARRY[71]), .A2(
        u5_mult_82_CLA_SUM[72]), .ZN(u5_mult_82_FS_1_n381) );
  AOI21_X4 u5_mult_82_FS_1_U630 ( .B1(u5_mult_82_FS_1_n569), .B2(
        u5_mult_82_FS_1_n570), .A(u5_mult_82_FS_1_n571), .ZN(
        u5_mult_82_FS_1_n567) );
  INV_X4 u5_mult_82_FS_1_U629 ( .A(u5_mult_82_FS_1_n349), .ZN(
        u5_mult_82_FS_1_n568) );
  OAI21_X4 u5_mult_82_FS_1_U628 ( .B1(u5_mult_82_FS_1_n560), .B2(
        u5_mult_82_FS_1_n561), .A(u5_mult_82_FS_1_n562), .ZN(
        u5_mult_82_FS_1_n84) );
  NOR2_X4 u5_mult_82_FS_1_U627 ( .A1(u5_mult_82_FS_1_n301), .A2(
        u5_mult_82_FS_1_n316), .ZN(u5_mult_82_FS_1_n557) );
  NAND2_X2 u5_mult_82_FS_1_U626 ( .A1(u5_mult_82_n486), .A2(
        u5_mult_82_CLA_SUM[81]), .ZN(u5_mult_82_FS_1_n304) );
  NAND2_X2 u5_mult_82_FS_1_U625 ( .A1(u5_mult_82_n485), .A2(
        u5_mult_82_CLA_SUM[80]), .ZN(u5_mult_82_FS_1_n300) );
  NAND2_X2 u5_mult_82_FS_1_U624 ( .A1(u5_mult_82_FS_1_n304), .A2(
        u5_mult_82_FS_1_n300), .ZN(u5_mult_82_FS_1_n559) );
  INV_X4 u5_mult_82_FS_1_U623 ( .A(u5_mult_82_FS_1_n305), .ZN(
        u5_mult_82_FS_1_n556) );
  NOR2_X4 u5_mult_82_FS_1_U622 ( .A1(u5_mult_82_FS_1_n555), .A2(
        u5_mult_82_FS_1_n556), .ZN(u5_mult_82_FS_1_n554) );
  NAND2_X2 u5_mult_82_FS_1_U621 ( .A1(u5_mult_82_CLA_CARRY[102]), .A2(
        u5_mult_82_n615), .ZN(u5_mult_82_FS_1_n544) );
  INV_X4 u5_mult_82_FS_1_U620 ( .A(u5_mult_82_CLA_CARRY[102]), .ZN(
        u5_mult_82_FS_1_n549) );
  INV_X4 u5_mult_82_FS_1_U619 ( .A(u5_mult_82_n615), .ZN(u5_mult_82_FS_1_n550)
         );
  NAND2_X2 u5_mult_82_FS_1_U618 ( .A1(u5_mult_82_FS_1_n549), .A2(
        u5_mult_82_FS_1_n550), .ZN(u5_mult_82_FS_1_n545) );
  NAND2_X2 u5_mult_82_FS_1_U617 ( .A1(u5_mult_82_FS_1_n544), .A2(
        u5_mult_82_FS_1_n545), .ZN(u5_mult_82_FS_1_n546) );
  XNOR2_X2 u5_mult_82_FS_1_U616 ( .A(u5_mult_82_FS_1_n547), .B(
        u5_mult_82_FS_1_n546), .ZN(u5_N103) );
  INV_X4 u5_mult_82_FS_1_U615 ( .A(u5_mult_82_FS_1_n545), .ZN(
        u5_mult_82_FS_1_n541) );
  OAI21_X4 u5_mult_82_FS_1_U614 ( .B1(u5_mult_82_FS_1_n541), .B2(
        u5_mult_82_FS_1_n543), .A(u5_mult_82_FS_1_n544), .ZN(
        u5_mult_82_FS_1_n530) );
  INV_X4 u5_mult_82_FS_1_U613 ( .A(u5_mult_82_FS_1_n530), .ZN(
        u5_mult_82_FS_1_n537) );
  INV_X4 u5_mult_82_FS_1_U612 ( .A(u5_mult_82_FS_1_n542), .ZN(
        u5_mult_82_FS_1_n540) );
  NOR2_X4 u5_mult_82_FS_1_U611 ( .A1(u5_mult_82_FS_1_n540), .A2(
        u5_mult_82_FS_1_n541), .ZN(u5_mult_82_FS_1_n524) );
  NAND2_X2 u5_mult_82_FS_1_U610 ( .A1(u5_mult_82_FS_1_n539), .A2(
        u5_mult_82_FS_1_n524), .ZN(u5_mult_82_FS_1_n538) );
  INV_X4 u5_mult_82_FS_1_U609 ( .A(u5_mult_82_CLA_CARRY[103]), .ZN(
        u5_mult_82_FS_1_n535) );
  INV_X4 u5_mult_82_FS_1_U608 ( .A(u5_mult_82_n616), .ZN(u5_mult_82_FS_1_n536)
         );
  NAND2_X2 u5_mult_82_FS_1_U607 ( .A1(u5_mult_82_FS_1_n535), .A2(
        u5_mult_82_FS_1_n536), .ZN(u5_mult_82_FS_1_n523) );
  NAND2_X2 u5_mult_82_FS_1_U606 ( .A1(u5_mult_82_CLA_CARRY[103]), .A2(
        u5_mult_82_n616), .ZN(u5_mult_82_FS_1_n529) );
  NAND2_X2 u5_mult_82_FS_1_U605 ( .A1(u5_mult_82_FS_1_n523), .A2(
        u5_mult_82_FS_1_n529), .ZN(u5_mult_82_FS_1_n534) );
  XNOR2_X2 u5_mult_82_FS_1_U604 ( .A(u5_mult_82_FS_1_n533), .B(
        u5_mult_82_FS_1_n534), .ZN(u5_N104) );
  NAND2_X2 u5_mult_82_FS_1_U603 ( .A1(u5_mult_82_FS_1_n524), .A2(
        u5_mult_82_FS_1_n523), .ZN(u5_mult_82_FS_1_n532) );
  NOR2_X4 u5_mult_82_FS_1_U602 ( .A1(u5_mult_82_FS_1_n531), .A2(
        u5_mult_82_FS_1_n532), .ZN(u5_mult_82_FS_1_n526) );
  NAND2_X2 u5_mult_82_FS_1_U601 ( .A1(u5_mult_82_FS_1_n523), .A2(
        u5_mult_82_FS_1_n530), .ZN(u5_mult_82_FS_1_n528) );
  NAND2_X2 u5_mult_82_FS_1_U600 ( .A1(u5_mult_82_FS_1_n528), .A2(
        u5_mult_82_FS_1_n529), .ZN(u5_mult_82_FS_1_n527) );
  NOR3_X4 u5_mult_82_FS_1_U599 ( .A1(u5_mult_82_FS_1_n284), .A2(
        u5_mult_82_FS_1_n121), .A3(u5_mult_82_FS_1_n283), .ZN(
        u5_mult_82_FS_1_n521) );
  NAND3_X2 u5_mult_82_FS_1_U598 ( .A1(u5_mult_82_FS_1_n516), .A2(
        u5_mult_82_FS_1_n518), .A3(u5_mult_82_FS_1_n517), .ZN(
        u5_mult_82_FS_1_n515) );
  XNOR2_X2 u5_mult_82_FS_1_U597 ( .A(u5_mult_82_FS_1_n515), .B(
        u5_mult_82_FS_1_n514), .ZN(u5_N105) );
  XNOR2_X2 u5_mult_82_FS_1_U596 ( .A(u5_mult_82_FS_1_n4), .B(
        u5_mult_82_FS_1_n510), .ZN(u5_N55) );
  XNOR2_X2 u5_mult_82_FS_1_U595 ( .A(u5_mult_82_FS_1_n504), .B(
        u5_mult_82_FS_1_n503), .ZN(u5_N57) );
  NAND2_X2 u5_mult_82_FS_1_U594 ( .A1(u5_mult_82_n575), .A2(
        u5_mult_82_CLA_SUM[58]), .ZN(u5_mult_82_FS_1_n484) );
  INV_X4 u5_mult_82_FS_1_U593 ( .A(u5_mult_82_FS_1_n484), .ZN(
        u5_mult_82_FS_1_n502) );
  INV_X4 u5_mult_82_FS_1_U592 ( .A(u5_mult_82_FS_1_n462), .ZN(
        u5_mult_82_FS_1_n493) );
  XNOR2_X2 u5_mult_82_FS_1_U591 ( .A(u5_mult_82_FS_1_n492), .B(
        u5_mult_82_FS_1_n5), .ZN(u5_N58) );
  NAND2_X2 u5_mult_82_FS_1_U590 ( .A1(u5_mult_82_FS_1_n491), .A2(
        u5_mult_82_FS_1_n485), .ZN(u5_mult_82_FS_1_n490) );
  XNOR2_X2 u5_mult_82_FS_1_U589 ( .A(u5_mult_82_FS_1_n489), .B(
        u5_mult_82_FS_1_n490), .ZN(u5_N59) );
  INV_X4 u5_mult_82_FS_1_U588 ( .A(u5_mult_82_FS_1_n486), .ZN(
        u5_mult_82_FS_1_n479) );
  INV_X4 u5_mult_82_FS_1_U587 ( .A(u5_mult_82_FS_1_n485), .ZN(
        u5_mult_82_FS_1_n481) );
  OAI21_X4 u5_mult_82_FS_1_U586 ( .B1(u5_mult_82_FS_1_n466), .B2(
        u5_mult_82_FS_1_n479), .A(u5_mult_82_FS_1_n480), .ZN(
        u5_mult_82_FS_1_n476) );
  XNOR2_X2 u5_mult_82_FS_1_U585 ( .A(u5_mult_82_FS_1_n476), .B(
        u5_mult_82_FS_1_n6), .ZN(u5_N60) );
  INV_X4 u5_mult_82_FS_1_U584 ( .A(u5_mult_82_FS_1_n476), .ZN(
        u5_mult_82_FS_1_n473) );
  XNOR2_X2 u5_mult_82_FS_1_U583 ( .A(u5_mult_82_FS_1_n471), .B(
        u5_mult_82_FS_1_n472), .ZN(u5_N61) );
  XNOR2_X2 u5_mult_82_FS_1_U582 ( .A(u5_mult_82_FS_1_n464), .B(
        u5_mult_82_FS_1_n465), .ZN(u5_N62) );
  INV_X4 u5_mult_82_FS_1_U581 ( .A(u5_mult_82_FS_1_n458), .ZN(
        u5_mult_82_FS_1_n457) );
  XNOR2_X2 u5_mult_82_FS_1_U580 ( .A(u5_mult_82_FS_1_n453), .B(
        u5_mult_82_FS_1_n454), .ZN(u5_N63) );
  NAND2_X2 u5_mult_82_FS_1_U579 ( .A1(u5_mult_82_FS_1_n447), .A2(
        u5_mult_82_FS_1_n450), .ZN(u5_mult_82_FS_1_n448) );
  XNOR2_X2 u5_mult_82_FS_1_U578 ( .A(u5_mult_82_FS_1_n448), .B(
        u5_mult_82_FS_1_n449), .ZN(u5_N64) );
  INV_X4 u5_mult_82_FS_1_U577 ( .A(u5_mult_82_FS_1_n447), .ZN(
        u5_mult_82_FS_1_n446) );
  XNOR2_X2 u5_mult_82_FS_1_U576 ( .A(u5_mult_82_FS_1_n438), .B(
        u5_mult_82_FS_1_n439), .ZN(u5_N65) );
  NAND2_X2 u5_mult_82_FS_1_U575 ( .A1(u5_mult_82_n581), .A2(
        u5_mult_82_CLA_SUM[66]), .ZN(u5_mult_82_FS_1_n431) );
  INV_X4 u5_mult_82_FS_1_U574 ( .A(u5_mult_82_FS_1_n431), .ZN(
        u5_mult_82_FS_1_n437) );
  NOR3_X4 u5_mult_82_FS_1_U573 ( .A1(u5_mult_82_FS_1_n121), .A2(
        u5_mult_82_FS_1_n283), .A3(u5_mult_82_FS_1_n284), .ZN(
        u5_mult_82_FS_1_n435) );
  NAND2_X2 u5_mult_82_FS_1_U572 ( .A1(u5_mult_82_FS_1_n689), .A2(
        u5_mult_82_FS_1_n432), .ZN(u5_mult_82_FS_1_n434) );
  XNOR2_X2 u5_mult_82_FS_1_U571 ( .A(u5_mult_82_FS_1_n433), .B(
        u5_mult_82_FS_1_n434), .ZN(u5_N67) );
  INV_X4 u5_mult_82_FS_1_U570 ( .A(u5_mult_82_FS_1_n432), .ZN(
        u5_mult_82_FS_1_n416) );
  NAND2_X2 u5_mult_82_FS_1_U569 ( .A1(u5_mult_82_FS_1_n427), .A2(
        u5_mult_82_FS_1_n428), .ZN(u5_mult_82_FS_1_n424) );
  NAND2_X2 u5_mult_82_FS_1_U568 ( .A1(u5_mult_82_FS_1_n583), .A2(
        u5_mult_82_FS_1_n423), .ZN(u5_mult_82_FS_1_n425) );
  XNOR2_X2 u5_mult_82_FS_1_U567 ( .A(u5_mult_82_FS_1_n424), .B(
        u5_mult_82_FS_1_n425), .ZN(u5_N68) );
  INV_X4 u5_mult_82_FS_1_U566 ( .A(u5_mult_82_FS_1_n423), .ZN(
        u5_mult_82_FS_1_n411) );
  NOR2_X4 u5_mult_82_FS_1_U565 ( .A1(u5_mult_82_FS_1_n411), .A2(
        u5_mult_82_FS_1_n412), .ZN(u5_mult_82_FS_1_n406) );
  INV_X4 u5_mult_82_FS_1_U564 ( .A(u5_mult_82_FS_1_n410), .ZN(
        u5_mult_82_FS_1_n408) );
  XNOR2_X2 u5_mult_82_FS_1_U563 ( .A(u5_mult_82_FS_1_n406), .B(
        u5_mult_82_FS_1_n407), .ZN(u5_N69) );
  NAND2_X2 u5_mult_82_FS_1_U562 ( .A1(u5_mult_82_FS_1_n402), .A2(
        u5_mult_82_FS_1_n403), .ZN(u5_mult_82_FS_1_n405) );
  XNOR2_X2 u5_mult_82_FS_1_U561 ( .A(u5_mult_82_FS_1_n404), .B(
        u5_mult_82_FS_1_n405), .ZN(u5_N70) );
  NAND2_X2 u5_mult_82_FS_1_U560 ( .A1(u5_mult_82_FS_1_n371), .A2(
        u5_mult_82_FS_1_n403), .ZN(u5_mult_82_FS_1_n399) );
  NAND2_X2 u5_mult_82_FS_1_U559 ( .A1(u5_mult_82_n574), .A2(
        u5_mult_82_CLA_SUM[71]), .ZN(u5_mult_82_FS_1_n380) );
  NAND2_X2 u5_mult_82_FS_1_U558 ( .A1(u5_mult_82_FS_1_n396), .A2(
        u5_mult_82_FS_1_n380), .ZN(u5_mult_82_FS_1_n401) );
  XNOR2_X2 u5_mult_82_FS_1_U557 ( .A(u5_mult_82_FS_1_n400), .B(
        u5_mult_82_FS_1_n401), .ZN(u5_N71) );
  INV_X4 u5_mult_82_FS_1_U556 ( .A(u5_mult_82_FS_1_n399), .ZN(
        u5_mult_82_FS_1_n398) );
  NAND2_X2 u5_mult_82_FS_1_U555 ( .A1(u5_mult_82_FS_1_n396), .A2(
        u5_mult_82_FS_1_n398), .ZN(u5_mult_82_FS_1_n393) );
  INV_X4 u5_mult_82_FS_1_U554 ( .A(u5_mult_82_FS_1_n380), .ZN(
        u5_mult_82_FS_1_n397) );
  XNOR2_X2 u5_mult_82_FS_1_U553 ( .A(u5_mult_82_FS_1_n391), .B(
        u5_mult_82_FS_1_n392), .ZN(u5_N72) );
  NAND2_X2 u5_mult_82_FS_1_U552 ( .A1(u5_mult_82_FS_1_n387), .A2(
        u5_mult_82_FS_1_n388), .ZN(u5_mult_82_FS_1_n386) );
  INV_X4 u5_mult_82_FS_1_U551 ( .A(u5_mult_82_FS_1_n375), .ZN(
        u5_mult_82_FS_1_n374) );
  XNOR2_X2 u5_mult_82_FS_1_U550 ( .A(u5_mult_82_FS_1_n373), .B(
        u5_mult_82_FS_1_n374), .ZN(u5_N73) );
  XNOR2_X2 u5_mult_82_FS_1_U549 ( .A(u5_mult_82_FS_1_n364), .B(
        u5_mult_82_FS_1_n365), .ZN(u5_N74) );
  OAI21_X4 u5_mult_82_FS_1_U548 ( .B1(u5_mult_82_FS_1_n339), .B2(
        u5_mult_82_FS_1_n361), .A(u5_mult_82_FS_1_n2), .ZN(
        u5_mult_82_FS_1_n360) );
  XNOR2_X2 u5_mult_82_FS_1_U547 ( .A(u5_mult_82_FS_1_n358), .B(
        u5_mult_82_FS_1_n359), .ZN(u5_N75) );
  NOR2_X4 u5_mult_82_FS_1_U546 ( .A1(u5_mult_82_FS_1_n353), .A2(
        u5_mult_82_FS_1_n354), .ZN(u5_mult_82_FS_1_n350) );
  INV_X4 u5_mult_82_FS_1_U545 ( .A(u5_mult_82_FS_1_n352), .ZN(
        u5_mult_82_FS_1_n345) );
  XNOR2_X2 u5_mult_82_FS_1_U544 ( .A(u5_mult_82_FS_1_n350), .B(
        u5_mult_82_FS_1_n351), .ZN(u5_N76) );
  NOR2_X4 u5_mult_82_FS_1_U543 ( .A1(u5_mult_82_FS_1_n348), .A2(
        u5_mult_82_FS_1_n9), .ZN(u5_mult_82_FS_1_n344) );
  INV_X4 u5_mult_82_FS_1_U542 ( .A(u5_mult_82_FS_1_n341), .ZN(
        u5_mult_82_FS_1_n340) );
  XNOR2_X2 u5_mult_82_FS_1_U541 ( .A(u5_mult_82_FS_1_n333), .B(
        u5_mult_82_FS_1_n334), .ZN(u5_N77) );
  XNOR2_X2 u5_mult_82_FS_1_U540 ( .A(u5_mult_82_FS_1_n328), .B(
        u5_mult_82_FS_1_n329), .ZN(u5_N78) );
  NAND2_X2 u5_mult_82_FS_1_U539 ( .A1(u5_mult_82_FS_1_n327), .A2(
        u5_mult_82_FS_1_n302), .ZN(u5_mult_82_FS_1_n318) );
  INV_X4 u5_mult_82_FS_1_U538 ( .A(u5_mult_82_FS_1_n326), .ZN(
        u5_mult_82_FS_1_n313) );
  XNOR2_X2 u5_mult_82_FS_1_U537 ( .A(u5_mult_82_FS_1_n318), .B(
        u5_mult_82_FS_1_n319), .ZN(u5_N79) );
  NOR2_X4 u5_mult_82_FS_1_U536 ( .A1(u5_mult_82_FS_1_n316), .A2(
        u5_mult_82_FS_1_n317), .ZN(u5_mult_82_FS_1_n303) );
  INV_X4 u5_mult_82_FS_1_U535 ( .A(u5_mult_82_FS_1_n302), .ZN(
        u5_mult_82_FS_1_n315) );
  NAND4_X2 u5_mult_82_FS_1_U534 ( .A1(u5_mult_82_FS_1_n308), .A2(
        u5_mult_82_FS_1_n295), .A3(u5_mult_82_FS_1_n309), .A4(
        u5_mult_82_FS_1_n293), .ZN(u5_mult_82_FS_1_n306) );
  XNOR2_X2 u5_mult_82_FS_1_U533 ( .A(u5_mult_82_FS_1_n306), .B(
        u5_mult_82_FS_1_n307), .ZN(u5_N80) );
  INV_X4 u5_mult_82_FS_1_U532 ( .A(u5_mult_82_FS_1_n300), .ZN(
        u5_mult_82_FS_1_n299) );
  INV_X4 u5_mult_82_FS_1_U531 ( .A(u5_mult_82_FS_1_n295), .ZN(
        u5_mult_82_FS_1_n294) );
  NOR2_X4 u5_mult_82_FS_1_U530 ( .A1(u5_mult_82_FS_1_n284), .A2(
        u5_mult_82_FS_1_n283), .ZN(u5_mult_82_FS_1_n282) );
  OAI21_X4 u5_mult_82_FS_1_U529 ( .B1(u5_mult_82_FS_1_n278), .B2(
        u5_mult_82_FS_1_n279), .A(u5_mult_82_FS_1_n149), .ZN(
        u5_mult_82_FS_1_n277) );
  NAND3_X4 u5_mult_82_FS_1_U528 ( .A1(u5_mult_82_FS_1_n277), .A2(
        u5_mult_82_FS_1_n23), .A3(u5_mult_82_FS_1_n83), .ZN(
        u5_mult_82_FS_1_n276) );
  NAND2_X2 u5_mult_82_FS_1_U527 ( .A1(u5_mult_82_CLA_SUM[82]), .A2(
        u5_mult_82_CLA_CARRY[81]), .ZN(u5_mult_82_FS_1_n274) );
  INV_X4 u5_mult_82_FS_1_U526 ( .A(u5_mult_82_FS_1_n274), .ZN(
        u5_mult_82_FS_1_n269) );
  XNOR2_X2 u5_mult_82_FS_1_U525 ( .A(u5_mult_82_FS_1_n272), .B(
        u5_mult_82_FS_1_n273), .ZN(u5_N83) );
  NOR2_X4 u5_mult_82_FS_1_U524 ( .A1(u5_mult_82_FS_1_n270), .A2(
        u5_mult_82_FS_1_n3), .ZN(u5_mult_82_FS_1_n268) );
  OAI21_X4 u5_mult_82_FS_1_U523 ( .B1(u5_mult_82_FS_1_n269), .B2(
        u5_mult_82_FS_1_n150), .A(u5_mult_82_FS_1_n268), .ZN(
        u5_mult_82_FS_1_n258) );
  INV_X4 u5_mult_82_FS_1_U522 ( .A(u5_mult_82_FS_1_n268), .ZN(
        u5_mult_82_FS_1_n267) );
  XNOR2_X2 u5_mult_82_FS_1_U521 ( .A(u5_mult_82_FS_1_n262), .B(
        u5_mult_82_FS_1_n263), .ZN(u5_N84) );
  INV_X4 u5_mult_82_FS_1_U520 ( .A(u5_mult_82_FS_1_n259), .ZN(
        u5_mult_82_FS_1_n256) );
  INV_X4 u5_mult_82_FS_1_U519 ( .A(u5_mult_82_FS_1_n255), .ZN(
        u5_mult_82_FS_1_n249) );
  XNOR2_X2 u5_mult_82_FS_1_U518 ( .A(u5_mult_82_FS_1_n245), .B(
        u5_mult_82_FS_1_n246), .ZN(u5_N85) );
  NAND2_X2 u5_mult_82_FS_1_U517 ( .A1(u5_mult_82_FS_1_n240), .A2(
        u5_mult_82_FS_1_n239), .ZN(u5_mult_82_FS_1_n242) );
  XNOR2_X2 u5_mult_82_FS_1_U516 ( .A(u5_mult_82_FS_1_n243), .B(
        u5_mult_82_FS_1_n242), .ZN(u5_N86) );
  INV_X4 u5_mult_82_FS_1_U515 ( .A(u5_mult_82_FS_1_n241), .ZN(
        u5_mult_82_FS_1_n206) );
  NAND2_X2 u5_mult_82_FS_1_U514 ( .A1(u5_mult_82_FS_1_n206), .A2(
        u5_mult_82_FS_1_n240), .ZN(u5_mult_82_FS_1_n234) );
  INV_X4 u5_mult_82_FS_1_U513 ( .A(u5_mult_82_FS_1_n240), .ZN(
        u5_mult_82_FS_1_n238) );
  XNOR2_X2 u5_mult_82_FS_1_U512 ( .A(u5_mult_82_FS_1_n236), .B(
        u5_mult_82_FS_1_n235), .ZN(u5_N87) );
  INV_X4 u5_mult_82_FS_1_U511 ( .A(u5_mult_82_FS_1_n234), .ZN(
        u5_mult_82_FS_1_n233) );
  NAND2_X2 u5_mult_82_FS_1_U510 ( .A1(u5_mult_82_FS_1_n233), .A2(
        u5_mult_82_FS_1_n232), .ZN(u5_mult_82_FS_1_n224) );
  NAND2_X2 u5_mult_82_FS_1_U509 ( .A1(u5_mult_82_FS_1_n231), .A2(
        u5_mult_82_FS_1_n232), .ZN(u5_mult_82_FS_1_n226) );
  XNOR2_X2 u5_mult_82_FS_1_U508 ( .A(u5_mult_82_FS_1_n229), .B(
        u5_mult_82_FS_1_n230), .ZN(u5_N88) );
  NAND3_X4 u5_mult_82_FS_1_U507 ( .A1(u5_mult_82_FS_1_n224), .A2(
        u5_mult_82_FS_1_n225), .A3(u5_mult_82_FS_1_n226), .ZN(
        u5_mult_82_FS_1_n215) );
  AOI21_X4 u5_mult_82_FS_1_U506 ( .B1(u5_mult_82_FS_1_n217), .B2(
        u5_mult_82_FS_1_n152), .A(u5_mult_82_FS_1_n81), .ZN(
        u5_mult_82_FS_1_n159) );
  NOR2_X4 u5_mult_82_FS_1_U505 ( .A1(u5_mult_82_FS_1_n600), .A2(
        u5_mult_82_FS_1_n205), .ZN(u5_mult_82_FS_1_n204) );
  AOI21_X4 u5_mult_82_FS_1_U504 ( .B1(u5_mult_82_FS_1_n202), .B2(
        u5_mult_82_FS_1_n203), .A(u5_mult_82_FS_1_n204), .ZN(
        u5_mult_82_FS_1_n164) );
  XNOR2_X2 u5_mult_82_FS_1_U503 ( .A(u5_mult_82_FS_1_n201), .B(
        u5_mult_82_FS_1_n200), .ZN(u5_N90) );
  INV_X4 u5_mult_82_FS_1_U502 ( .A(u5_mult_82_FS_1_n199), .ZN(
        u5_mult_82_FS_1_n167) );
  INV_X4 u5_mult_82_FS_1_U501 ( .A(u5_mult_82_FS_1_n198), .ZN(
        u5_mult_82_FS_1_n196) );
  NAND2_X2 u5_mult_82_FS_1_U500 ( .A1(u5_mult_82_FS_1_n176), .A2(
        u5_mult_82_FS_1_n174), .ZN(u5_mult_82_FS_1_n184) );
  INV_X4 u5_mult_82_FS_1_U499 ( .A(u5_mult_82_FS_1_n192), .ZN(
        u5_mult_82_FS_1_n190) );
  INV_X4 u5_mult_82_FS_1_U498 ( .A(u5_mult_82_FS_1_n182), .ZN(
        u5_mult_82_FS_1_n187) );
  NOR2_X4 u5_mult_82_FS_1_U497 ( .A1(u5_mult_82_FS_1_n189), .A2(
        u5_mult_82_FS_1_n188), .ZN(u5_mult_82_FS_1_n179) );
  XNOR2_X2 u5_mult_82_FS_1_U496 ( .A(u5_mult_82_FS_1_n185), .B(
        u5_mult_82_FS_1_n184), .ZN(u5_N92) );
  NOR2_X4 u5_mult_82_FS_1_U495 ( .A1(u5_mult_82_FS_1_n179), .A2(
        u5_mult_82_FS_1_n180), .ZN(u5_mult_82_FS_1_n177) );
  NAND2_X2 u5_mult_82_FS_1_U494 ( .A1(u5_mult_82_FS_1_n178), .A2(
        u5_mult_82_FS_1_n176), .ZN(u5_mult_82_FS_1_n173) );
  NAND2_X2 u5_mult_82_FS_1_U493 ( .A1(u5_mult_82_FS_1_n170), .A2(
        u5_mult_82_FS_1_n171), .ZN(u5_mult_82_FS_1_n169) );
  XNOR2_X2 u5_mult_82_FS_1_U492 ( .A(u5_mult_82_FS_1_n168), .B(
        u5_mult_82_FS_1_n169), .ZN(u5_N93) );
  NAND2_X2 u5_mult_82_FS_1_U491 ( .A1(u5_mult_82_FS_1_n142), .A2(
        u5_mult_82_FS_1_n143), .ZN(u5_mult_82_FS_1_n162) );
  NAND2_X2 u5_mult_82_FS_1_U490 ( .A1(u5_mult_82_FS_1_n167), .A2(
        u5_mult_82_FS_1_n599), .ZN(u5_mult_82_FS_1_n147) );
  OAI21_X4 u5_mult_82_FS_1_U489 ( .B1(u5_mult_82_FS_1_n164), .B2(
        u5_mult_82_FS_1_n165), .A(u5_mult_82_FS_1_n166), .ZN(
        u5_mult_82_FS_1_n145) );
  XNOR2_X2 u5_mult_82_FS_1_U488 ( .A(u5_mult_82_FS_1_n163), .B(
        u5_mult_82_FS_1_n162), .ZN(u5_N94) );
  NAND2_X2 u5_mult_82_FS_1_U487 ( .A1(u5_mult_82_FS_1_n144), .A2(
        u5_mult_82_FS_1_n128), .ZN(u5_mult_82_FS_1_n154) );
  XNOR2_X2 u5_mult_82_FS_1_U486 ( .A(u5_mult_82_FS_1_n155), .B(
        u5_mult_82_FS_1_n154), .ZN(u5_N95) );
  NAND2_X2 u5_mult_82_FS_1_U485 ( .A1(u5_mult_82_FS_1_n153), .A2(
        u5_mult_82_FS_1_n113), .ZN(u5_mult_82_FS_1_n138) );
  INV_X4 u5_mult_82_FS_1_U484 ( .A(u5_mult_82_FS_1_n147), .ZN(
        u5_mult_82_FS_1_n146) );
  NAND3_X4 u5_mult_82_FS_1_U483 ( .A1(u5_mult_82_FS_1_n143), .A2(
        u5_mult_82_FS_1_n144), .A3(u5_mult_82_FS_1_n146), .ZN(
        u5_mult_82_FS_1_n134) );
  NAND3_X4 u5_mult_82_FS_1_U482 ( .A1(u5_mult_82_FS_1_n145), .A2(
        u5_mult_82_FS_1_n144), .A3(u5_mult_82_FS_1_n143), .ZN(
        u5_mult_82_FS_1_n137) );
  INV_X4 u5_mult_82_FS_1_U481 ( .A(u5_mult_82_FS_1_n128), .ZN(
        u5_mult_82_FS_1_n136) );
  NOR2_X4 u5_mult_82_FS_1_U480 ( .A1(u5_mult_82_FS_1_n141), .A2(
        u5_mult_82_FS_1_n142), .ZN(u5_mult_82_FS_1_n129) );
  XNOR2_X2 u5_mult_82_FS_1_U479 ( .A(u5_mult_82_FS_1_n139), .B(
        u5_mult_82_FS_1_n138), .ZN(u5_N96) );
  INV_X4 u5_mult_82_FS_1_U478 ( .A(u5_mult_82_FS_1_n137), .ZN(
        u5_mult_82_FS_1_n130) );
  NAND2_X2 u5_mult_82_FS_1_U477 ( .A1(u5_mult_82_FS_1_n134), .A2(
        u5_mult_82_FS_1_n135), .ZN(u5_mult_82_FS_1_n133) );
  NOR2_X4 u5_mult_82_FS_1_U476 ( .A1(u5_mult_82_FS_1_n130), .A2(
        u5_mult_82_FS_1_n133), .ZN(u5_mult_82_FS_1_n132) );
  NOR2_X4 u5_mult_82_FS_1_U475 ( .A1(u5_mult_82_FS_1_n131), .A2(
        u5_mult_82_FS_1_n132), .ZN(u5_mult_82_FS_1_n111) );
  NOR2_X4 u5_mult_82_FS_1_U474 ( .A1(u5_mult_82_FS_1_n129), .A2(
        u5_mult_82_FS_1_n130), .ZN(u5_mult_82_FS_1_n114) );
  NAND2_X2 u5_mult_82_FS_1_U473 ( .A1(u5_mult_82_FS_1_n83), .A2(
        u5_mult_82_FS_1_n128), .ZN(u5_mult_82_FS_1_n127) );
  NAND3_X2 u5_mult_82_FS_1_U472 ( .A1(u5_mult_82_FS_1_n114), .A2(
        u5_mult_82_FS_1_n115), .A3(u5_mult_82_FS_1_n116), .ZN(
        u5_mult_82_FS_1_n112) );
  INV_X4 u5_mult_82_FS_1_U471 ( .A(u5_mult_82_FS_1_n110), .ZN(
        u5_mult_82_FS_1_n108) );
  NOR2_X4 u5_mult_82_FS_1_U470 ( .A1(u5_mult_82_FS_1_n108), .A2(
        u5_mult_82_FS_1_n109), .ZN(u5_mult_82_FS_1_n107) );
  NAND2_X2 u5_mult_82_FS_1_U469 ( .A1(u5_mult_82_FS_1_n101), .A2(
        u5_mult_82_FS_1_n99), .ZN(u5_mult_82_FS_1_n102) );
  XNOR2_X2 u5_mult_82_FS_1_U468 ( .A(u5_mult_82_FS_1_n103), .B(
        u5_mult_82_FS_1_n102), .ZN(u5_N98) );
  NAND2_X2 u5_mult_82_FS_1_U467 ( .A1(u5_mult_82_FS_1_n91), .A2(
        u5_mult_82_FS_1_n76), .ZN(u5_mult_82_FS_1_n94) );
  NAND2_X2 u5_mult_82_FS_1_U466 ( .A1(u5_mult_82_FS_1_n100), .A2(
        u5_mult_82_FS_1_n101), .ZN(u5_mult_82_FS_1_n93) );
  OAI21_X4 u5_mult_82_FS_1_U465 ( .B1(u5_mult_82_FS_1_n97), .B2(
        u5_mult_82_FS_1_n98), .A(u5_mult_82_FS_1_n99), .ZN(u5_mult_82_FS_1_n90) );
  XNOR2_X2 u5_mult_82_FS_1_U464 ( .A(u5_mult_82_FS_1_n95), .B(
        u5_mult_82_FS_1_n94), .ZN(u5_N99) );
  NAND2_X2 u5_mult_82_FS_1_U463 ( .A1(u5_mult_82_FS_1_n74), .A2(
        u5_mult_82_FS_1_n72), .ZN(u5_mult_82_FS_1_n87) );
  INV_X4 u5_mult_82_FS_1_U462 ( .A(u5_mult_82_FS_1_n93), .ZN(
        u5_mult_82_FS_1_n92) );
  NAND2_X2 u5_mult_82_FS_1_U461 ( .A1(u5_mult_82_FS_1_n92), .A2(
        u5_mult_82_FS_1_n91), .ZN(u5_mult_82_FS_1_n75) );
  XNOR2_X2 u5_mult_82_FS_1_U460 ( .A(u5_mult_82_FS_1_n88), .B(
        u5_mult_82_FS_1_n87), .ZN(u5_N100) );
  NAND2_X2 u5_mult_82_FS_1_U459 ( .A1(u5_mult_82_FS_1_n85), .A2(
        u5_mult_82_FS_1_n86), .ZN(u5_mult_82_FS_1_n68) );
  OAI21_X4 u5_mult_82_FS_1_U458 ( .B1(u5_mult_82_FS_1_n80), .B2(
        u5_mult_82_FS_1_n81), .A(u5_mult_82_FS_1_n77), .ZN(u5_mult_82_FS_1_n79) );
  INV_X16 u5_mult_82_FS_1_U457 ( .A(u5_mult_82_FS_1_n276), .ZN(
        u5_mult_82_FS_1_n89) );
  NOR2_X1 u5_mult_82_FS_1_U456 ( .A1(u5_mult_82_CLA_SUM[54]), .A2(
        u5_mult_82_CLA_CARRY[53]), .ZN(u5_mult_82_FS_1_n512) );
  NAND3_X2 u5_mult_82_FS_1_U455 ( .A1(u5_mult_82_FS_1_n215), .A2(
        u5_mult_82_FS_1_n216), .A3(u5_mult_82_FS_1_n159), .ZN(
        u5_mult_82_FS_1_n214) );
  NAND2_X1 u5_mult_82_FS_1_U454 ( .A1(u5_mult_82_FS_1_n501), .A2(
        u5_mult_82_FS_1_n500), .ZN(u5_mult_82_FS_1_n462) );
  NOR3_X1 u5_mult_82_FS_1_U453 ( .A1(u5_mult_82_FS_1_n421), .A2(
        u5_mult_82_FS_1_n125), .A3(u5_mult_82_FS_1_n422), .ZN(
        u5_mult_82_FS_1_n413) );
  NAND2_X1 u5_mult_82_FS_1_U452 ( .A1(u5_mult_82_FS_1_n417), .A2(
        u5_mult_82_FS_1_n40), .ZN(u5_mult_82_FS_1_n428) );
  NAND3_X2 u5_mult_82_FS_1_U451 ( .A1(u5_mult_82_FS_1_n222), .A2(
        u5_mult_82_FS_1_n282), .A3(u5_mult_82_FS_1_n218), .ZN(
        u5_mult_82_FS_1_n278) );
  NAND2_X1 u5_mult_82_FS_1_U450 ( .A1(u5_mult_82_FS_1_n223), .A2(
        u5_mult_82_FS_1_n222), .ZN(u5_mult_82_FS_1_n421) );
  NAND2_X4 u5_mult_82_FS_1_U449 ( .A1(u5_mult_82_FS_1_n715), .A2(
        u5_mult_82_FS_1_n716), .ZN(u5_mult_82_FS_1_n143) );
  NAND2_X1 u5_mult_82_FS_1_U448 ( .A1(u5_mult_82_FS_1_n12), .A2(
        u5_mult_82_FS_1_n159), .ZN(u5_mult_82_FS_1_n157) );
  NOR2_X2 u5_mult_82_FS_1_U447 ( .A1(u5_mult_82_CLA_SUM[56]), .A2(
        u5_mult_82_n579), .ZN(u5_mult_82_FS_1_n506) );
  NAND2_X1 u5_mult_82_FS_1_U446 ( .A1(u5_mult_82_n579), .A2(
        u5_mult_82_CLA_SUM[56]), .ZN(u5_mult_82_FS_1_n507) );
  AOI21_X4 u5_mult_82_FS_1_U445 ( .B1(u5_mult_82_FS_1_n497), .B2(
        u5_mult_82_FS_1_n498), .A(u5_mult_82_FS_1_n487), .ZN(
        u5_mult_82_FS_1_n664) );
  NOR3_X4 u5_mult_82_FS_1_U444 ( .A1(u5_mult_82_FS_1_n124), .A2(
        u5_mult_82_FS_1_n125), .A3(u5_mult_82_FS_1_n219), .ZN(
        u5_mult_82_FS_1_n436) );
  OAI211_X4 u5_mult_82_FS_1_U443 ( .C1(u5_mult_82_FS_1_n89), .C2(
        u5_mult_82_FS_1_n75), .A(u5_mult_82_FS_1_n77), .B(u5_mult_82_FS_1_n76), 
        .ZN(u5_mult_82_FS_1_n88) );
  OAI211_X4 u5_mult_82_FS_1_U442 ( .C1(u5_mult_82_FS_1_n172), .C2(
        u5_mult_82_FS_1_n173), .A(u5_mult_82_FS_1_n175), .B(
        u5_mult_82_FS_1_n174), .ZN(u5_mult_82_FS_1_n168) );
  OAI211_X4 u5_mult_82_FS_1_U441 ( .C1(u5_mult_82_FS_1_n89), .C2(
        u5_mult_82_FS_1_n224), .A(u5_mult_82_FS_1_n225), .B(
        u5_mult_82_FS_1_n226), .ZN(u5_mult_82_FS_1_n229) );
  OAI21_X2 u5_mult_82_FS_1_U440 ( .B1(u5_mult_82_FS_1_n89), .B2(
        u5_mult_82_FS_1_n199), .A(u5_mult_82_FS_1_n18), .ZN(
        u5_mult_82_FS_1_n201) );
  OAI21_X2 u5_mult_82_FS_1_U439 ( .B1(u5_mult_82_FS_1_n89), .B2(
        u5_mult_82_FS_1_n234), .A(u5_mult_82_FS_1_n237), .ZN(
        u5_mult_82_FS_1_n236) );
  OAI21_X2 u5_mult_82_FS_1_U438 ( .B1(u5_mult_82_FS_1_n89), .B2(
        u5_mult_82_FS_1_n93), .A(u5_mult_82_FS_1_n96), .ZN(u5_mult_82_FS_1_n95) );
  OAI21_X2 u5_mult_82_FS_1_U437 ( .B1(u5_mult_82_FS_1_n89), .B2(
        u5_mult_82_FS_1_n241), .A(u5_mult_82_FS_1_n600), .ZN(
        u5_mult_82_FS_1_n243) );
  OAI21_X2 u5_mult_82_FS_1_U436 ( .B1(u5_mult_82_FS_1_n89), .B2(
        u5_mult_82_FS_1_n147), .A(u5_mult_82_FS_1_n161), .ZN(
        u5_mult_82_FS_1_n163) );
  OAI21_X2 u5_mult_82_FS_1_U435 ( .B1(u5_mult_82_FS_1_n89), .B2(
        u5_mult_82_FS_1_n181), .A(u5_mult_82_FS_1_n186), .ZN(
        u5_mult_82_FS_1_n185) );
  OAI21_X2 u5_mult_82_FS_1_U434 ( .B1(u5_mult_82_FS_1_n89), .B2(
        u5_mult_82_FS_1_n3), .A(u5_mult_82_FS_1_n274), .ZN(
        u5_mult_82_FS_1_n272) );
  XNOR2_X1 u5_mult_82_FS_1_U433 ( .A(u5_mult_82_FS_1_n89), .B(
        u5_mult_82_FS_1_n275), .ZN(u5_N82) );
  INV_X8 u5_mult_82_FS_1_U432 ( .A(u5_mult_82_FS_1_n467), .ZN(
        u5_mult_82_FS_1_n280) );
  INV_X4 u5_mult_82_FS_1_U431 ( .A(u5_mult_82_FS_1_n64), .ZN(
        u5_mult_82_FS_1_n65) );
  NAND2_X1 u5_mult_82_FS_1_U430 ( .A1(u5_mult_82_FS_1_n294), .A2(
        u5_mult_82_FS_1_n292), .ZN(u5_mult_82_FS_1_n289) );
  NOR3_X2 u5_mult_82_FS_1_U429 ( .A1(u5_mult_82_FS_1_n7), .A2(
        u5_mult_82_FS_1_n298), .A3(u5_mult_82_FS_1_n299), .ZN(
        u5_mult_82_FS_1_n287) );
  INV_X4 u5_mult_82_FS_1_U428 ( .A(u5_mult_82_FS_1_n62), .ZN(
        u5_mult_82_FS_1_n63) );
  INV_X4 u5_mult_82_FS_1_U427 ( .A(u5_mult_82_FS_1_n209), .ZN(
        u5_mult_82_FS_1_n59) );
  NOR2_X4 u5_mult_82_FS_1_U426 ( .A1(u5_mult_82_FS_1_n78), .A2(
        u5_mult_82_FS_1_n79), .ZN(u5_mult_82_FS_1_n70) );
  NOR3_X4 u5_mult_82_FS_1_U425 ( .A1(u5_mult_82_FS_1_n124), .A2(
        u5_mult_82_FS_1_n125), .A3(u5_mult_82_FS_1_n219), .ZN(
        u5_mult_82_FS_1_n118) );
  INV_X1 u5_mult_82_FS_1_U424 ( .A(u5_mult_82_FS_1_n68), .ZN(
        u5_mult_82_FS_1_n55) );
  NAND2_X2 u5_mult_82_FS_1_U423 ( .A1(u5_mult_82_FS_1_n56), .A2(
        u5_mult_82_FS_1_n57), .ZN(u5_N101) );
  NAND2_X1 u5_mult_82_FS_1_U422 ( .A1(u5_mult_82_FS_1_n191), .A2(
        u5_mult_82_FS_1_n182), .ZN(u5_mult_82_FS_1_n193) );
  INV_X4 u5_mult_82_FS_1_U421 ( .A(u5_mult_82_FS_1_n193), .ZN(
        u5_mult_82_FS_1_n51) );
  NAND2_X2 u5_mult_82_FS_1_U420 ( .A1(u5_mult_82_FS_1_n53), .A2(
        u5_mult_82_FS_1_n54), .ZN(u5_N91) );
  NAND2_X2 u5_mult_82_FS_1_U419 ( .A1(u5_mult_82_FS_1_n51), .A2(
        u5_mult_82_FS_1_n52), .ZN(u5_mult_82_FS_1_n54) );
  NAND2_X1 u5_mult_82_FS_1_U418 ( .A1(u5_mult_82_FS_1_n193), .A2(
        u5_mult_82_FS_1_n194), .ZN(u5_mult_82_FS_1_n53) );
  NAND2_X4 u5_mult_82_FS_1_U417 ( .A1(u5_mult_82_FS_1_n628), .A2(
        u5_mult_82_FS_1_n627), .ZN(u5_mult_82_FS_1_n552) );
  BUF_X4 u5_mult_82_FS_1_U416 ( .A(u5_mult_82_n5330), .Z(u5_mult_82_FS_1_n50)
         );
  NAND2_X4 u5_mult_82_FS_1_U415 ( .A1(u5_mult_82_FS_1_n656), .A2(
        u5_mult_82_FS_1_n657), .ZN(u5_mult_82_FS_1_n509) );
  NAND2_X4 u5_mult_82_FS_1_U414 ( .A1(u5_mult_82_CLA_CARRY[53]), .A2(
        u5_mult_82_CLA_SUM[54]), .ZN(u5_mult_82_FS_1_n497) );
  INV_X4 u5_mult_82_FS_1_U413 ( .A(u5_mult_82_n624), .ZN(u5_mult_82_FS_1_n514)
         );
  NAND2_X2 u5_mult_82_FS_1_U412 ( .A1(u5_mult_82_FS_1_n223), .A2(
        u5_mult_82_FS_1_n221), .ZN(u5_mult_82_FS_1_n279) );
  NAND2_X4 u5_mult_82_FS_1_U411 ( .A1(u5_mult_82_FS_1_n436), .A2(
        u5_mult_82_FS_1_n435), .ZN(u5_mult_82_FS_1_n296) );
  NAND2_X2 u5_mult_82_FS_1_U410 ( .A1(u5_mult_82_FS_1_n118), .A2(
        u5_mult_82_FS_1_n119), .ZN(u5_mult_82_FS_1_n117) );
  OAI21_X2 u5_mult_82_FS_1_U409 ( .B1(u5_mult_82_FS_1_n320), .B2(
        u5_mult_82_FS_1_n393), .A(u5_mult_82_FS_1_n394), .ZN(
        u5_mult_82_FS_1_n392) );
  OAI21_X2 u5_mult_82_FS_1_U408 ( .B1(u5_mult_82_FS_1_n320), .B2(
        u5_mult_82_FS_1_n338), .A(u5_mult_82_FS_1_n361), .ZN(
        u5_mult_82_FS_1_n365) );
  OAI21_X2 u5_mult_82_FS_1_U407 ( .B1(u5_mult_82_FS_1_n320), .B2(
        u5_mult_82_FS_1_n357), .A(u5_mult_82_FS_1_n348), .ZN(
        u5_mult_82_FS_1_n359) );
  OAI21_X2 u5_mult_82_FS_1_U406 ( .B1(u5_mult_82_FS_1_n320), .B2(
        u5_mult_82_FS_1_n321), .A(u5_mult_82_FS_1_n322), .ZN(
        u5_mult_82_FS_1_n319) );
  OAI21_X2 u5_mult_82_FS_1_U405 ( .B1(u5_mult_82_FS_1_n320), .B2(
        u5_mult_82_FS_1_n430), .A(u5_mult_82_FS_1_n431), .ZN(
        u5_mult_82_FS_1_n433) );
  OAI21_X2 u5_mult_82_FS_1_U404 ( .B1(u5_mult_82_FS_1_n320), .B2(
        u5_mult_82_FS_1_n399), .A(u5_mult_82_FS_1_n383), .ZN(
        u5_mult_82_FS_1_n400) );
  OAI21_X2 u5_mult_82_FS_1_U403 ( .B1(u5_mult_82_FS_1_n320), .B2(
        u5_mult_82_FS_1_n389), .A(u5_mult_82_FS_1_n28), .ZN(
        u5_mult_82_FS_1_n404) );
  INV_X8 u5_mult_82_FS_1_U402 ( .A(u5_mult_82_FS_1_n477), .ZN(
        u5_mult_82_FS_1_n470) );
  NOR2_X4 u5_mult_82_FS_1_U401 ( .A1(u5_mult_82_FS_1_n653), .A2(
        u5_mult_82_FS_1_n49), .ZN(u5_mult_82_FS_1_n652) );
  NAND2_X4 u5_mult_82_FS_1_U400 ( .A1(u5_mult_82_CLA_SUM[55]), .A2(
        u5_mult_82_n1604), .ZN(u5_mult_82_FS_1_n498) );
  NAND3_X4 u5_mult_82_FS_1_U399 ( .A1(u5_mult_82_FS_1_n222), .A2(
        u5_mult_82_FS_1_n221), .A3(u5_mult_82_FS_1_n223), .ZN(
        u5_mult_82_FS_1_n265) );
  NOR2_X4 u5_mult_82_FS_1_U398 ( .A1(u5_mult_82_FS_1_n499), .A2(
        u5_mult_82_FS_1_n483), .ZN(u5_mult_82_FS_1_n660) );
  NAND3_X1 u5_mult_82_FS_1_U397 ( .A1(u5_mult_82_FS_1_n123), .A2(
        u5_mult_82_FS_1_n218), .A3(u5_mult_82_FS_1_n122), .ZN(
        u5_mult_82_FS_1_n264) );
  NAND2_X4 u5_mult_82_FS_1_U396 ( .A1(u5_mult_82_FS_1_n118), .A2(
        u5_mult_82_FS_1_n629), .ZN(u5_mult_82_FS_1_n628) );
  NOR2_X4 u5_mult_82_FS_1_U395 ( .A1(u5_mult_82_FS_1_n219), .A2(
        u5_mult_82_FS_1_n125), .ZN(u5_mult_82_FS_1_n64) );
  INV_X2 u5_mult_82_FS_1_U394 ( .A(u5_mult_82_FS_1_n506), .ZN(
        u5_mult_82_FS_1_n511) );
  NAND2_X1 u5_mult_82_FS_1_U393 ( .A1(u5_mult_82_n573), .A2(
        u5_mult_82_FS_1_n50), .ZN(u5_mult_82_FS_1_n485) );
  NAND2_X4 u5_mult_82_FS_1_U392 ( .A1(u5_mult_82_FS_1_n31), .A2(
        u5_mult_82_FS_1_n542), .ZN(u5_mult_82_FS_1_n548) );
  AOI21_X4 u5_mult_82_FS_1_U391 ( .B1(u5_mult_82_FS_1_n111), .B2(
        u5_mult_82_FS_1_n112), .A(u5_mult_82_FS_1_n596), .ZN(
        u5_mult_82_FS_1_n106) );
  NAND2_X4 u5_mult_82_FS_1_U390 ( .A1(u5_mult_82_FS_1_n663), .A2(
        u5_mult_82_FS_1_n662), .ZN(u5_mult_82_FS_1_n477) );
  NAND2_X4 u5_mult_82_FS_1_U389 ( .A1(u5_mult_82_FS_1_n667), .A2(
        u5_mult_82_FS_1_n668), .ZN(u5_mult_82_FS_1_n444) );
  NAND2_X1 u5_mult_82_FS_1_U388 ( .A1(u5_mult_82_FS_1_n477), .A2(
        u5_mult_82_FS_1_n478), .ZN(u5_mult_82_FS_1_n471) );
  AOI22_X4 u5_mult_82_FS_1_U387 ( .A1(u5_mult_82_FS_1_n126), .A2(
        u5_mult_82_FS_1_n525), .B1(u5_mult_82_FS_1_n150), .B2(
        u5_mult_82_FS_1_n525), .ZN(u5_mult_82_FS_1_n553) );
  OAI21_X1 u5_mult_82_FS_1_U386 ( .B1(u5_mult_82_FS_1_n366), .B2(
        u5_mult_82_FS_1_n8), .A(u5_mult_82_FS_1_n402), .ZN(
        u5_mult_82_FS_1_n395) );
  NOR2_X4 u5_mult_82_FS_1_U385 ( .A1(u5_mult_82_FS_1_n220), .A2(
        u5_mult_82_FS_1_n219), .ZN(u5_mult_82_FS_1_n217) );
  NAND2_X4 u5_mult_82_FS_1_U384 ( .A1(u5_mult_82_FS_1_n670), .A2(
        u5_mult_82_FS_1_n669), .ZN(u5_mult_82_FS_1_n455) );
  NAND2_X4 u5_mult_82_FS_1_U383 ( .A1(u5_mult_82_CLA_SUM[62]), .A2(
        u5_mult_82_n588), .ZN(u5_mult_82_FS_1_n452) );
  NAND2_X4 u5_mult_82_FS_1_U382 ( .A1(u5_mult_82_FS_1_n520), .A2(
        u5_mult_82_FS_1_n521), .ZN(u5_mult_82_FS_1_n82) );
  NAND2_X4 u5_mult_82_FS_1_U381 ( .A1(u5_mult_82_n592), .A2(
        u5_mult_82_CLA_SUM[63]), .ZN(u5_mult_82_FS_1_n447) );
  NAND2_X1 u5_mult_82_FS_1_U380 ( .A1(u5_mult_82_FS_1_n454), .A2(
        u5_mult_82_FS_1_n444), .ZN(u5_mult_82_FS_1_n450) );
  NAND2_X1 u5_mult_82_FS_1_U379 ( .A1(u5_mult_82_FS_1_n444), .A2(
        u5_mult_82_FS_1_n447), .ZN(u5_mult_82_FS_1_n453) );
  NAND3_X1 u5_mult_82_FS_1_U378 ( .A1(u5_mult_82_FS_1_n584), .A2(
        u5_mult_82_n578), .A3(u5_mult_82_CLA_SUM[68]), .ZN(
        u5_mult_82_FS_1_n581) );
  INV_X2 u5_mult_82_FS_1_U377 ( .A(u5_mult_82_FS_1_n584), .ZN(
        u5_mult_82_FS_1_n409) );
  OAI211_X2 u5_mult_82_FS_1_U376 ( .C1(u5_mult_82_FS_1_n320), .C2(
        u5_mult_82_FS_1_n326), .A(u5_mult_82_FS_1_n314), .B(
        u5_mult_82_FS_1_n325), .ZN(u5_mult_82_FS_1_n328) );
  NOR2_X4 u5_mult_82_FS_1_U375 ( .A1(u5_mult_82_FS_1_n500), .A2(
        u5_mult_82_FS_1_n648), .ZN(u5_mult_82_FS_1_n654) );
  NAND3_X4 u5_mult_82_FS_1_U374 ( .A1(u5_mult_82_FS_1_n673), .A2(
        u5_mult_82_FS_1_n396), .A3(u5_mult_82_FS_1_n382), .ZN(
        u5_mult_82_FS_1_n367) );
  NAND2_X4 u5_mult_82_FS_1_U373 ( .A1(u5_mult_82_FS_1_n677), .A2(
        u5_mult_82_FS_1_n678), .ZN(u5_mult_82_FS_1_n382) );
  NOR2_X1 u5_mult_82_FS_1_U372 ( .A1(u5_mult_82_FS_1_n429), .A2(
        u5_mult_82_FS_1_n430), .ZN(u5_mult_82_FS_1_n417) );
  NAND2_X4 u5_mult_82_FS_1_U371 ( .A1(u5_mult_82_FS_1_n691), .A2(
        u5_mult_82_FS_1_n692), .ZN(u5_mult_82_FS_1_n584) );
  NOR2_X1 u5_mult_82_FS_1_U370 ( .A1(u5_mult_82_FS_1_n483), .A2(
        u5_mult_82_FS_1_n484), .ZN(u5_mult_82_FS_1_n482) );
  NAND2_X1 u5_mult_82_FS_1_U369 ( .A1(u5_mult_82_n578), .A2(
        u5_mult_82_CLA_SUM[68]), .ZN(u5_mult_82_FS_1_n423) );
  NOR2_X4 u5_mult_82_FS_1_U368 ( .A1(u5_mult_82_FS_1_n643), .A2(
        u5_mult_82_FS_1_n452), .ZN(u5_mult_82_FS_1_n640) );
  NAND3_X1 u5_mult_82_FS_1_U367 ( .A1(u5_mult_82_FS_1_n20), .A2(
        u5_mult_82_FS_1_n182), .A3(u5_mult_82_FS_1_n83), .ZN(
        u5_mult_82_FS_1_n183) );
  NAND3_X1 u5_mult_82_FS_1_U366 ( .A1(u5_mult_82_FS_1_n83), .A2(
        u5_mult_82_FS_1_n76), .A3(u5_mult_82_FS_1_n20), .ZN(
        u5_mult_82_FS_1_n78) );
  NAND2_X1 u5_mult_82_FS_1_U365 ( .A1(u5_mult_82_n608), .A2(u5_mult_82_n5565), 
        .ZN(u5_mult_82_FS_1_n410) );
  INV_X4 u5_mult_82_FS_1_U364 ( .A(u5_mult_82_FS_1_n107), .ZN(
        u5_mult_82_FS_1_n42) );
  INV_X4 u5_mult_82_FS_1_U363 ( .A(u5_mult_82_FS_1_n106), .ZN(
        u5_mult_82_FS_1_n41) );
  NAND2_X2 u5_mult_82_FS_1_U362 ( .A1(u5_mult_82_FS_1_n43), .A2(
        u5_mult_82_FS_1_n44), .ZN(u5_N97) );
  NAND2_X4 u5_mult_82_FS_1_U361 ( .A1(u5_mult_82_FS_1_n41), .A2(
        u5_mult_82_FS_1_n42), .ZN(u5_mult_82_FS_1_n44) );
  NAND2_X2 u5_mult_82_FS_1_U360 ( .A1(u5_mult_82_FS_1_n106), .A2(
        u5_mult_82_FS_1_n107), .ZN(u5_mult_82_FS_1_n43) );
  NOR2_X4 u5_mult_82_FS_1_U359 ( .A1(u5_mult_82_FS_1_n366), .A2(
        u5_mult_82_FS_1_n46), .ZN(u5_mult_82_FS_1_n560) );
  INV_X1 u5_mult_82_FS_1_U358 ( .A(u5_mult_82_FS_1_n483), .ZN(
        u5_mult_82_FS_1_n491) );
  NAND2_X1 u5_mult_82_FS_1_U357 ( .A1(u5_mult_82_FS_1_n304), .A2(
        u5_mult_82_FS_1_n305), .ZN(u5_mult_82_FS_1_n285) );
  NAND2_X4 u5_mult_82_FS_1_U356 ( .A1(u5_mult_82_FS_1_n436), .A2(
        u5_mult_82_FS_1_n435), .ZN(u5_mult_82_FS_1_n40) );
  INV_X4 u5_mult_82_FS_1_U355 ( .A(u5_mult_82_FS_1_n285), .ZN(
        u5_mult_82_FS_1_n36) );
  NAND2_X2 u5_mult_82_FS_1_U354 ( .A1(u5_mult_82_FS_1_n38), .A2(
        u5_mult_82_FS_1_n39), .ZN(u5_N81) );
  NAND2_X2 u5_mult_82_FS_1_U353 ( .A1(u5_mult_82_FS_1_n36), .A2(
        u5_mult_82_FS_1_n37), .ZN(u5_mult_82_FS_1_n39) );
  NAND2_X1 u5_mult_82_FS_1_U352 ( .A1(u5_mult_82_FS_1_n285), .A2(
        u5_mult_82_FS_1_n286), .ZN(u5_mult_82_FS_1_n38) );
  OAI21_X4 u5_mult_82_FS_1_U351 ( .B1(u5_mult_82_FS_1_n89), .B2(
        u5_mult_82_FS_1_n192), .A(u5_mult_82_FS_1_n189), .ZN(
        u5_mult_82_FS_1_n194) );
  NAND2_X1 u5_mult_82_FS_1_U350 ( .A1(u5_mult_82_FS_1_n446), .A2(
        u5_mult_82_FS_1_n445), .ZN(u5_mult_82_FS_1_n442) );
  NAND2_X1 u5_mult_82_FS_1_U349 ( .A1(u5_mult_82_FS_1_n445), .A2(
        u5_mult_82_FS_1_n441), .ZN(u5_mult_82_FS_1_n449) );
  NAND2_X1 u5_mult_82_FS_1_U348 ( .A1(u5_mult_82_FS_1_n122), .A2(
        u5_mult_82_FS_1_n123), .ZN(u5_mult_82_FS_1_n120) );
  NAND2_X1 u5_mult_82_FS_1_U347 ( .A1(u5_mult_82_FS_1_n420), .A2(
        u5_mult_82_FS_1_n1), .ZN(u5_mult_82_FS_1_n419) );
  NOR2_X1 u5_mult_82_FS_1_U346 ( .A1(u5_mult_82_FS_1_n389), .A2(
        u5_mult_82_FS_1_n8), .ZN(u5_mult_82_FS_1_n387) );
  NAND3_X2 u5_mult_82_FS_1_U345 ( .A1(u5_mult_82_FS_1_n441), .A2(
        u5_mult_82_FS_1_n442), .A3(u5_mult_82_FS_1_n443), .ZN(
        u5_mult_82_FS_1_n438) );
  INV_X4 u5_mult_82_FS_1_U344 ( .A(u5_mult_82_FS_1_n208), .ZN(
        u5_mult_82_FS_1_n58) );
  NAND2_X4 u5_mult_82_FS_1_U343 ( .A1(u5_mult_82_FS_1_n548), .A2(
        u5_mult_82_FS_1_n543), .ZN(u5_mult_82_FS_1_n547) );
  INV_X16 u5_mult_82_FS_1_U342 ( .A(u5_mult_82_FS_1_n221), .ZN(
        u5_mult_82_FS_1_n125) );
  NAND2_X4 u5_mult_82_FS_1_U341 ( .A1(u5_mult_82_FS_1_n671), .A2(
        u5_mult_82_FS_1_n672), .ZN(u5_mult_82_FS_1_n81) );
  NAND3_X2 u5_mult_82_FS_1_U340 ( .A1(u5_mult_82_FS_1_n160), .A2(
        u5_mult_82_FS_1_n143), .A3(u5_mult_82_FS_1_n158), .ZN(
        u5_mult_82_FS_1_n156) );
  AOI21_X2 u5_mult_82_FS_1_U339 ( .B1(u5_mult_82_FS_1_n413), .B2(
        u5_mult_82_FS_1_n414), .A(u5_mult_82_FS_1_n415), .ZN(
        u5_mult_82_FS_1_n412) );
  OAI21_X1 u5_mult_82_FS_1_U338 ( .B1(u5_mult_82_FS_1_n385), .B2(
        u5_mult_82_FS_1_n380), .A(u5_mult_82_FS_1_n381), .ZN(
        u5_mult_82_FS_1_n379) );
  NOR2_X4 u5_mult_82_FS_1_U337 ( .A1(u5_mult_82_FS_1_n377), .A2(
        u5_mult_82_FS_1_n10), .ZN(u5_mult_82_FS_1_n373) );
  INV_X8 u5_mult_82_FS_1_U336 ( .A(u5_mult_82_FS_1_n222), .ZN(
        u5_mult_82_FS_1_n124) );
  NOR2_X2 u5_mult_82_FS_1_U335 ( .A1(u5_mult_82_FS_1_n81), .A2(
        u5_mult_82_FS_1_n267), .ZN(u5_mult_82_FS_1_n266) );
  NAND2_X4 u5_mult_82_FS_1_U334 ( .A1(u5_mult_82_FS_1_n335), .A2(
        u5_mult_82_FS_1_n336), .ZN(u5_mult_82_FS_1_n334) );
  NAND2_X1 u5_mult_82_FS_1_U333 ( .A1(u5_mult_82_FS_1_n376), .A2(
        u5_mult_82_FS_1_n369), .ZN(u5_mult_82_FS_1_n375) );
  NAND2_X4 u5_mult_82_FS_1_U332 ( .A1(u5_mult_82_FS_1_n683), .A2(
        u5_mult_82_FS_1_n684), .ZN(u5_mult_82_FS_1_n356) );
  NAND3_X4 u5_mult_82_FS_1_U331 ( .A1(u5_mult_82_FS_1_n666), .A2(
        u5_mult_82_FS_1_n455), .A3(u5_mult_82_FS_1_n444), .ZN(
        u5_mult_82_FS_1_n665) );
  NAND2_X1 u5_mult_82_FS_1_U330 ( .A1(u5_mult_82_FS_1_n455), .A2(
        u5_mult_82_FS_1_n452), .ZN(u5_mult_82_FS_1_n464) );
  NOR2_X4 u5_mult_82_FS_1_U329 ( .A1(u5_mult_82_FS_1_n121), .A2(
        u5_mult_82_FS_1_n630), .ZN(u5_mult_82_FS_1_n152) );
  NAND2_X2 u5_mult_82_FS_1_U328 ( .A1(u5_mult_82_FS_1_n208), .A2(
        u5_mult_82_FS_1_n209), .ZN(u5_mult_82_FS_1_n60) );
  NOR2_X2 u5_mult_82_FS_1_U327 ( .A1(u5_mult_82_FS_1_n469), .A2(
        u5_mult_82_FS_1_n470), .ZN(u5_mult_82_FS_1_n459) );
  NAND3_X4 u5_mult_82_FS_1_U326 ( .A1(u5_mult_82_FS_1_n645), .A2(
        u5_mult_82_FS_1_n646), .A3(u5_mult_82_FS_1_n647), .ZN(
        u5_mult_82_FS_1_n467) );
  NOR2_X2 u5_mult_82_FS_1_U325 ( .A1(u5_mult_82_FS_1_n474), .A2(
        u5_mult_82_FS_1_n470), .ZN(u5_mult_82_FS_1_n647) );
  INV_X16 u5_mult_82_FS_1_U324 ( .A(u5_mult_82_FS_1_n665), .ZN(
        u5_mult_82_FS_1_n281) );
  NAND2_X1 u5_mult_82_FS_1_U323 ( .A1(u5_mult_82_CLA_CARRY[66]), .A2(
        u5_mult_82_CLA_SUM[67]), .ZN(u5_mult_82_FS_1_n432) );
  NOR2_X4 u5_mult_82_FS_1_U322 ( .A1(u5_mult_82_FS_1_n474), .A2(
        u5_mult_82_FS_1_n470), .ZN(u5_mult_82_FS_1_n48) );
  OAI21_X4 u5_mult_82_FS_1_U321 ( .B1(u5_mult_82_FS_1_n70), .B2(
        u5_mult_82_FS_1_n71), .A(u5_mult_82_FS_1_n72), .ZN(u5_mult_82_FS_1_n69) );
  INV_X4 u5_mult_82_FS_1_U320 ( .A(u5_mult_82_FS_1_n69), .ZN(
        u5_mult_82_FS_1_n35) );
  NAND2_X4 u5_mult_82_FS_1_U319 ( .A1(u5_mult_82_CLA_SUM[74]), .A2(
        u5_mult_82_n584), .ZN(u5_mult_82_FS_1_n362) );
  INV_X4 u5_mult_82_FS_1_U318 ( .A(u5_mult_82_FS_1_n66), .ZN(
        u5_mult_82_FS_1_n67) );
  NAND2_X4 u5_mult_82_FS_1_U317 ( .A1(u5_mult_82_n484), .A2(
        u5_mult_82_CLA_SUM[73]), .ZN(u5_mult_82_FS_1_n376) );
  NAND2_X4 u5_mult_82_FS_1_U316 ( .A1(u5_mult_82_FS_1_n310), .A2(
        u5_mult_82_FS_1_n22), .ZN(u5_mult_82_FS_1_n293) );
  NAND2_X4 u5_mult_82_FS_1_U315 ( .A1(u5_mult_82_FS_1_n681), .A2(
        u5_mult_82_FS_1_n682), .ZN(u5_mult_82_FS_1_n680) );
  OAI211_X4 u5_mult_82_FS_1_U314 ( .C1(u5_mult_82_FS_1_n140), .C2(
        u5_mult_82_FS_1_n134), .A(u5_mult_82_FS_1_n137), .B(
        u5_mult_82_FS_1_n135), .ZN(u5_mult_82_FS_1_n139) );
  NAND2_X4 u5_mult_82_FS_1_U313 ( .A1(u5_mult_82_FS_1_n675), .A2(
        u5_mult_82_FS_1_n676), .ZN(u5_mult_82_FS_1_n369) );
  NAND2_X4 u5_mult_82_FS_1_U312 ( .A1(u5_mult_82_FS_1_n441), .A2(
        u5_mult_82_FS_1_n447), .ZN(u5_mult_82_FS_1_n641) );
  INV_X8 u5_mult_82_FS_1_U311 ( .A(u5_mult_82_FS_1_n572), .ZN(
        u5_mult_82_FS_1_n330) );
  NOR2_X4 u5_mult_82_FS_1_U310 ( .A1(u5_mult_82_n583), .A2(
        u5_mult_82_CLA_SUM[64]), .ZN(u5_mult_82_FS_1_n34) );
  NAND2_X4 u5_mult_82_FS_1_U309 ( .A1(u5_mult_82_n583), .A2(
        u5_mult_82_CLA_SUM[64]), .ZN(u5_mult_82_FS_1_n441) );
  NOR2_X4 u5_mult_82_FS_1_U308 ( .A1(u5_mult_82_FS_1_n567), .A2(
        u5_mult_82_FS_1_n568), .ZN(u5_mult_82_FS_1_n566) );
  NOR2_X2 u5_mult_82_FS_1_U307 ( .A1(u5_mult_82_FS_1_n343), .A2(
        u5_mult_82_FS_1_n342), .ZN(u5_mult_82_FS_1_n569) );
  NOR2_X1 u5_mult_82_FS_1_U306 ( .A1(u5_mult_82_FS_1_n342), .A2(
        u5_mult_82_FS_1_n343), .ZN(u5_mult_82_FS_1_n341) );
  NOR2_X1 u5_mult_82_FS_1_U305 ( .A1(u5_mult_82_FS_1_n342), .A2(
        u5_mult_82_FS_1_n347), .ZN(u5_mult_82_FS_1_n346) );
  NOR2_X1 u5_mult_82_FS_1_U304 ( .A1(u5_mult_82_FS_1_n345), .A2(
        u5_mult_82_FS_1_n342), .ZN(u5_mult_82_FS_1_n351) );
  INV_X1 u5_mult_82_FS_1_U303 ( .A(u5_mult_82_FS_1_n390), .ZN(
        u5_mult_82_FS_1_n403) );
  NAND3_X2 u5_mult_82_FS_1_U302 ( .A1(u5_mult_82_FS_1_n496), .A2(
        u5_mult_82_FS_1_n495), .A3(u5_mult_82_FS_1_n494), .ZN(
        u5_mult_82_FS_1_n460) );
  NOR2_X2 u5_mult_82_FS_1_U301 ( .A1(u5_mult_82_FS_1_n512), .A2(
        u5_mult_82_FS_1_n510), .ZN(u5_N54) );
  AOI21_X2 u5_mult_82_FS_1_U300 ( .B1(u5_mult_82_FS_1_n249), .B2(
        u5_mult_82_FS_1_n250), .A(u5_mult_82_FS_1_n251), .ZN(
        u5_mult_82_FS_1_n248) );
  OAI21_X4 u5_mult_82_FS_1_U299 ( .B1(u5_mult_82_FS_1_n565), .B2(
        u5_mult_82_FS_1_n564), .A(u5_mult_82_FS_1_n314), .ZN(
        u5_mult_82_FS_1_n561) );
  NAND2_X1 u5_mult_82_FS_1_U298 ( .A1(u5_mult_82_FS_1_n382), .A2(
        u5_mult_82_FS_1_n381), .ZN(u5_mult_82_FS_1_n391) );
  NOR2_X1 u5_mult_82_FS_1_U297 ( .A1(u5_mult_82_FS_1_n487), .A2(
        u5_mult_82_FS_1_n483), .ZN(u5_mult_82_FS_1_n486) );
  NAND2_X4 u5_mult_82_FS_1_U296 ( .A1(u5_mult_82_CLA_CARRY[82]), .A2(
        u5_mult_82_CLA_SUM[83]), .ZN(u5_mult_82_FS_1_n253) );
  NAND2_X4 u5_mult_82_FS_1_U295 ( .A1(u5_mult_82_FS_1_n371), .A2(
        u5_mult_82_FS_1_n372), .ZN(u5_mult_82_FS_1_n338) );
  NAND2_X1 u5_mult_82_FS_1_U294 ( .A1(u5_mult_82_FS_1_n349), .A2(
        u5_mult_82_FS_1_n33), .ZN(u5_mult_82_FS_1_n333) );
  NAND2_X4 u5_mult_82_FS_1_U293 ( .A1(u5_mult_82_n591), .A2(
        u5_mult_82_CLA_SUM[76]), .ZN(u5_mult_82_FS_1_n352) );
  INV_X8 u5_mult_82_FS_1_U292 ( .A(u5_mult_82_FS_1_n356), .ZN(
        u5_mult_82_FS_1_n343) );
  NAND2_X2 u5_mult_82_FS_1_U291 ( .A1(u5_mult_82_FS_1_n369), .A2(
        u5_mult_82_FS_1_n370), .ZN(u5_mult_82_FS_1_n368) );
  NAND2_X1 u5_mult_82_FS_1_U290 ( .A1(u5_mult_82_n577), .A2(
        u5_mult_82_FS_1_n26), .ZN(u5_mult_82_FS_1_n402) );
  NAND2_X4 u5_mult_82_FS_1_U289 ( .A1(u5_mult_82_FS_1_n33), .A2(
        u5_mult_82_FS_1_n352), .ZN(u5_mult_82_FS_1_n571) );
  AOI21_X1 u5_mult_82_FS_1_U288 ( .B1(u5_mult_82_FS_1_n17), .B2(
        u5_mult_82_FS_1_n396), .A(u5_mult_82_FS_1_n397), .ZN(
        u5_mult_82_FS_1_n394) );
  NAND2_X4 u5_mult_82_FS_1_U287 ( .A1(u5_mult_82_FS_1_n58), .A2(
        u5_mult_82_FS_1_n59), .ZN(u5_mult_82_FS_1_n61) );
  INV_X8 u5_mult_82_FS_1_U286 ( .A(u5_mult_82_FS_1_n293), .ZN(
        u5_mult_82_FS_1_n291) );
  NAND3_X2 u5_mult_82_FS_1_U285 ( .A1(u5_mult_82_FS_1_n552), .A2(
        u5_mult_82_FS_1_n553), .A3(u5_mult_82_FS_1_n531), .ZN(
        u5_mult_82_FS_1_n539) );
  NAND3_X2 u5_mult_82_FS_1_U284 ( .A1(u5_mult_82_FS_1_n552), .A2(
        u5_mult_82_FS_1_n553), .A3(u5_mult_82_FS_1_n531), .ZN(
        u5_mult_82_FS_1_n31) );
  INV_X8 u5_mult_82_FS_1_U283 ( .A(u5_mult_82_FS_1_n680), .ZN(
        u5_mult_82_FS_1_n342) );
  NOR2_X2 u5_mult_82_FS_1_U282 ( .A1(u5_mult_82_FS_1_n367), .A2(
        u5_mult_82_FS_1_n572), .ZN(u5_mult_82_FS_1_n672) );
  INV_X8 u5_mult_82_FS_1_U281 ( .A(u5_mult_82_FS_1_n384), .ZN(
        u5_mult_82_FS_1_n396) );
  NOR3_X1 u5_mult_82_FS_1_U280 ( .A1(u5_mult_82_FS_1_n383), .A2(
        u5_mult_82_FS_1_n384), .A3(u5_mult_82_FS_1_n385), .ZN(
        u5_mult_82_FS_1_n378) );
  NOR2_X1 u5_mult_82_FS_1_U279 ( .A1(u5_mult_82_FS_1_n385), .A2(
        u5_mult_82_FS_1_n384), .ZN(u5_mult_82_FS_1_n388) );
  AOI22_X2 u5_mult_82_FS_1_U278 ( .A1(u5_mult_82_FS_1_n150), .A2(
        u5_mult_82_FS_1_n519), .B1(u5_mult_82_FS_1_n519), .B2(
        u5_mult_82_FS_1_n228), .ZN(u5_mult_82_FS_1_n518) );
  NOR2_X4 u5_mult_82_FS_1_U277 ( .A1(u5_mult_82_FS_1_n367), .A2(
        u5_mult_82_FS_1_n572), .ZN(u5_mult_82_FS_1_n45) );
  NAND2_X1 u5_mult_82_FS_1_U276 ( .A1(u5_mult_82_FS_1_n363), .A2(
        u5_mult_82_FS_1_n2), .ZN(u5_mult_82_FS_1_n364) );
  NAND2_X4 u5_mult_82_FS_1_U275 ( .A1(u5_mult_82_FS_1_n721), .A2(
        u5_mult_82_FS_1_n722), .ZN(u5_mult_82_FS_1_n250) );
  NAND3_X2 u5_mult_82_FS_1_U274 ( .A1(u5_mult_82_FS_1_n576), .A2(
        u5_mult_82_FS_1_n381), .A3(u5_mult_82_FS_1_n376), .ZN(
        u5_mult_82_FS_1_n575) );
  OAI211_X4 u5_mult_82_FS_1_U273 ( .C1(u5_mult_82_FS_1_n604), .C2(
        u5_mult_82_FS_1_n605), .A(u5_mult_82_FS_1_n253), .B(
        u5_mult_82_FS_1_n254), .ZN(u5_mult_82_FS_1_n602) );
  INV_X1 u5_mult_82_FS_1_U272 ( .A(u5_mult_82_FS_1_n382), .ZN(
        u5_mult_82_FS_1_n385) );
  NAND3_X1 u5_mult_82_FS_1_U271 ( .A1(u5_mult_82_FS_1_n552), .A2(
        u5_mult_82_FS_1_n531), .A3(u5_mult_82_FS_1_n553), .ZN(
        u5_mult_82_FS_1_n32) );
  NAND2_X4 u5_mult_82_FS_1_U270 ( .A1(u5_mult_82_n585), .A2(
        u5_mult_82_CLA_SUM[78]), .ZN(u5_mult_82_FS_1_n317) );
  OAI21_X1 u5_mult_82_FS_1_U269 ( .B1(u5_mult_82_FS_1_n252), .B2(
        u5_mult_82_FS_1_n253), .A(u5_mult_82_FS_1_n254), .ZN(
        u5_mult_82_FS_1_n251) );
  INV_X2 u5_mult_82_FS_1_U268 ( .A(u5_mult_82_FS_1_n177), .ZN(
        u5_mult_82_FS_1_n178) );
  NAND2_X1 u5_mult_82_FS_1_U267 ( .A1(u5_mult_82_FS_1_n253), .A2(
        u5_mult_82_FS_1_n717), .ZN(u5_mult_82_FS_1_n273) );
  INV_X2 u5_mult_82_FS_1_U266 ( .A(u5_mult_82_FS_1_n563), .ZN(
        u5_mult_82_FS_1_n562) );
  INV_X8 u5_mult_82_FS_1_U265 ( .A(u5_mult_82_FS_1_n145), .ZN(
        u5_mult_82_FS_1_n161) );
  INV_X4 u5_mult_82_FS_1_U264 ( .A(u5_mult_82_FS_1_n29), .ZN(
        u5_mult_82_FS_1_n30) );
  NAND2_X4 u5_mult_82_FS_1_U263 ( .A1(u5_mult_82_FS_1_n685), .A2(
        u5_mult_82_FS_1_n686), .ZN(u5_mult_82_FS_1_n349) );
  INV_X2 u5_mult_82_FS_1_U262 ( .A(u5_mult_82_FS_1_n27), .ZN(
        u5_mult_82_FS_1_n28) );
  INV_X1 u5_mult_82_FS_1_U261 ( .A(u5_mult_82_FS_1_n366), .ZN(
        u5_mult_82_FS_1_n27) );
  NAND2_X4 u5_mult_82_FS_1_U260 ( .A1(u5_mult_82_FS_1_n687), .A2(
        u5_mult_82_FS_1_n688), .ZN(u5_mult_82_FS_1_n363) );
  BUF_X8 u5_mult_82_FS_1_U259 ( .A(u5_mult_82_CLA_SUM[70]), .Z(
        u5_mult_82_FS_1_n26) );
  NAND2_X1 u5_mult_82_FS_1_U258 ( .A1(u5_mult_82_FS_1_n356), .A2(
        u5_mult_82_FS_1_n347), .ZN(u5_mult_82_FS_1_n358) );
  NOR2_X2 u5_mult_82_FS_1_U257 ( .A1(u5_mult_82_FS_1_n587), .A2(
        u5_mult_82_FS_1_n81), .ZN(u5_mult_82_FS_1_n627) );
  NAND2_X1 u5_mult_82_FS_1_U256 ( .A1(u5_mult_82_FS_1_n566), .A2(
        u5_mult_82_FS_1_n22), .ZN(u5_mult_82_FS_1_n295) );
  OAI21_X4 u5_mult_82_FS_1_U255 ( .B1(u5_mult_82_CLA_SUM[71]), .B2(
        u5_mult_82_n574), .A(u5_mult_82_FS_1_n382), .ZN(u5_mult_82_FS_1_n578)
         );
  INV_X4 u5_mult_82_FS_1_U254 ( .A(u5_mult_82_FS_1_n664), .ZN(
        u5_mult_82_FS_1_n658) );
  NOR3_X1 u5_mult_82_FS_1_U253 ( .A1(u5_mult_82_FS_1_n338), .A2(
        u5_mult_82_FS_1_n339), .A3(u5_mult_82_FS_1_n340), .ZN(
        u5_mult_82_FS_1_n337) );
  NAND2_X1 u5_mult_82_FS_1_U252 ( .A1(u5_mult_82_FS_1_n250), .A2(
        u5_mult_82_FS_1_n254), .ZN(u5_mult_82_FS_1_n262) );
  NAND2_X4 u5_mult_82_FS_1_U251 ( .A1(u5_mult_82_FS_1_n697), .A2(
        u5_mult_82_FS_1_n698), .ZN(u5_mult_82_FS_1_n292) );
  NOR2_X1 u5_mult_82_FS_1_U250 ( .A1(u5_mult_82_FS_1_n187), .A2(
        u5_mult_82_FS_1_n179), .ZN(u5_mult_82_FS_1_n186) );
  NAND2_X4 u5_mult_82_FS_1_U249 ( .A1(u5_mult_82_FS_1_n693), .A2(
        u5_mult_82_FS_1_n694), .ZN(u5_mult_82_FS_1_n327) );
  NOR2_X1 u5_mult_82_FS_1_U248 ( .A1(u5_mult_82_FS_1_n408), .A2(
        u5_mult_82_FS_1_n409), .ZN(u5_mult_82_FS_1_n407) );
  NAND2_X4 u5_mult_82_FS_1_U247 ( .A1(u5_mult_82_CLA_SUM[79]), .A2(
        u5_mult_82_n587), .ZN(u5_mult_82_FS_1_n302) );
  NAND2_X4 u5_mult_82_FS_1_U246 ( .A1(u5_mult_82_FS_1_n719), .A2(
        u5_mult_82_FS_1_n720), .ZN(u5_mult_82_FS_1_n260) );
  NAND2_X4 u5_mult_82_FS_1_U245 ( .A1(u5_mult_82_FS_1_n661), .A2(
        u5_mult_82_FS_1_n660), .ZN(u5_mult_82_FS_1_n659) );
  NAND2_X1 u5_mult_82_FS_1_U244 ( .A1(u5_mult_82_FS_1_n260), .A2(
        u5_mult_82_FS_1_n261), .ZN(u5_mult_82_FS_1_n245) );
  AOI21_X4 u5_mult_82_FS_1_U243 ( .B1(u5_mult_82_FS_1_n557), .B2(
        u5_mult_82_FS_1_n558), .A(u5_mult_82_FS_1_n559), .ZN(
        u5_mult_82_FS_1_n555) );
  OAI21_X4 u5_mult_82_FS_1_U242 ( .B1(u5_mult_82_FS_1_n196), .B2(
        u5_mult_82_FS_1_n164), .A(u5_mult_82_FS_1_n197), .ZN(
        u5_mult_82_FS_1_n195) );
  NAND2_X2 u5_mult_82_FS_1_U241 ( .A1(u5_mult_82_FS_1_n161), .A2(
        u5_mult_82_FS_1_n147), .ZN(u5_mult_82_FS_1_n158) );
  NAND2_X1 u5_mult_82_FS_1_U240 ( .A1(u5_mult_82_FS_1_n216), .A2(
        u5_mult_82_FS_1_n232), .ZN(u5_mult_82_FS_1_n616) );
  NAND2_X1 u5_mult_82_FS_1_U239 ( .A1(u5_mult_82_FS_1_n215), .A2(
        u5_mult_82_FS_1_n216), .ZN(u5_mult_82_FS_1_n212) );
  NAND2_X1 u5_mult_82_FS_1_U238 ( .A1(u5_mult_82_FS_1_n216), .A2(
        u5_mult_82_FS_1_n213), .ZN(u5_mult_82_FS_1_n230) );
  NAND2_X4 u5_mult_82_FS_1_U237 ( .A1(u5_mult_82_FS_1_n728), .A2(
        u5_mult_82_FS_1_n729), .ZN(u5_mult_82_FS_1_n232) );
  NAND3_X4 u5_mult_82_FS_1_U236 ( .A1(u5_mult_82_CLA_SUM[71]), .A2(
        u5_mult_82_n574), .A3(u5_mult_82_FS_1_n382), .ZN(u5_mult_82_FS_1_n576)
         );
  NAND2_X4 u5_mult_82_FS_1_U235 ( .A1(u5_mult_82_FS_1_n161), .A2(
        u5_mult_82_FS_1_n83), .ZN(u5_mult_82_FS_1_n29) );
  INV_X4 u5_mult_82_FS_1_U234 ( .A(u5_mult_82_FS_1_n195), .ZN(
        u5_mult_82_FS_1_n189) );
  INV_X2 u5_mult_82_FS_1_U233 ( .A(u5_mult_82_FS_1_n426), .ZN(
        u5_mult_82_FS_1_n583) );
  INV_X8 u5_mult_82_FS_1_U232 ( .A(u5_mult_82_FS_1_n566), .ZN(
        u5_mult_82_FS_1_n314) );
  INV_X1 u5_mult_82_FS_1_U231 ( .A(u5_mult_82_FS_1_n34), .ZN(
        u5_mult_82_FS_1_n445) );
  INV_X4 u5_mult_82_FS_1_U230 ( .A(u5_mult_82_FS_1_n84), .ZN(
        u5_mult_82_FS_1_n126) );
  INV_X4 u5_mult_82_FS_1_U229 ( .A(u5_mult_82_FS_1_n45), .ZN(
        u5_mult_82_FS_1_n46) );
  NAND3_X2 u5_mult_82_FS_1_U228 ( .A1(u5_mult_82_FS_1_n311), .A2(
        u5_mult_82_FS_1_n305), .A3(u5_mult_82_FS_1_n292), .ZN(
        u5_mult_82_FS_1_n563) );
  NAND2_X1 u5_mult_82_FS_1_U227 ( .A1(u5_mult_82_FS_1_n323), .A2(
        u5_mult_82_FS_1_n313), .ZN(u5_mult_82_FS_1_n321) );
  AOI21_X1 u5_mult_82_FS_1_U226 ( .B1(u5_mult_82_FS_1_n310), .B2(
        u5_mult_82_FS_1_n323), .A(u5_mult_82_FS_1_n324), .ZN(
        u5_mult_82_FS_1_n322) );
  NAND2_X1 u5_mult_82_FS_1_U225 ( .A1(u5_mult_82_FS_1_n323), .A2(
        u5_mult_82_FS_1_n317), .ZN(u5_mult_82_FS_1_n329) );
  NAND4_X4 u5_mult_82_FS_1_U224 ( .A1(u5_mult_82_FS_1_n593), .A2(
        u5_mult_82_FS_1_n594), .A3(u5_mult_82_FS_1_n595), .A4(
        u5_mult_82_FS_1_n110), .ZN(u5_mult_82_FS_1_n105) );
  NAND2_X4 u5_mult_82_FS_1_U223 ( .A1(u5_mult_82_FS_1_n90), .A2(
        u5_mult_82_FS_1_n91), .ZN(u5_mult_82_FS_1_n77) );
  NAND3_X2 u5_mult_82_FS_1_U222 ( .A1(u5_mult_82_FS_1_n444), .A2(
        u5_mult_82_FS_1_n445), .A3(u5_mult_82_FS_1_n454), .ZN(
        u5_mult_82_FS_1_n443) );
  INV_X8 u5_mult_82_FS_1_U221 ( .A(u5_mult_82_CLA_SUM[63]), .ZN(
        u5_mult_82_FS_1_n668) );
  INV_X8 u5_mult_82_FS_1_U220 ( .A(u5_mult_82_FS_1_n522), .ZN(
        u5_mult_82_FS_1_n519) );
  INV_X4 u5_mult_82_FS_1_U219 ( .A(u5_mult_82_FS_1_n389), .ZN(
        u5_mult_82_FS_1_n371) );
  INV_X4 u5_mult_82_FS_1_U218 ( .A(u5_mult_82_FS_1_n325), .ZN(
        u5_mult_82_FS_1_n310) );
  NAND2_X4 u5_mult_82_FS_1_U217 ( .A1(u5_mult_82_FS_1_n167), .A2(
        u5_mult_82_FS_1_n198), .ZN(u5_mult_82_FS_1_n192) );
  NAND3_X2 u5_mult_82_FS_1_U216 ( .A1(u5_mult_82_FS_1_n457), .A2(
        u5_mult_82_FS_1_n456), .A3(u5_mult_82_FS_1_n455), .ZN(
        u5_mult_82_FS_1_n451) );
  NAND2_X4 u5_mult_82_FS_1_U215 ( .A1(u5_mult_82_FS_1_n732), .A2(
        u5_mult_82_FS_1_n733), .ZN(u5_mult_82_FS_1_n240) );
  INV_X8 u5_mult_82_FS_1_U214 ( .A(u5_mult_82_FS_1_n292), .ZN(
        u5_mult_82_FS_1_n301) );
  NAND2_X1 u5_mult_82_FS_1_U213 ( .A1(u5_mult_82_FS_1_n292), .A2(
        u5_mult_82_FS_1_n300), .ZN(u5_mult_82_FS_1_n307) );
  INV_X16 u5_mult_82_FS_1_U212 ( .A(u5_mult_82_FS_1_n223), .ZN(
        u5_mult_82_FS_1_n219) );
  INV_X4 u5_mult_82_FS_1_U211 ( .A(u5_mult_82_FS_1_n260), .ZN(
        u5_mult_82_FS_1_n606) );
  NOR2_X2 u5_mult_82_FS_1_U210 ( .A1(u5_mult_82_FS_1_n252), .A2(
        u5_mult_82_FS_1_n606), .ZN(u5_mult_82_FS_1_n601) );
  INV_X8 u5_mult_82_FS_1_U209 ( .A(u5_mult_82_FS_1_n122), .ZN(
        u5_mult_82_FS_1_n284) );
  NAND2_X2 u5_mult_82_FS_1_U208 ( .A1(u5_mult_82_FS_1_n247), .A2(
        u5_mult_82_FS_1_n248), .ZN(u5_mult_82_FS_1_n246) );
  NOR2_X2 u5_mult_82_FS_1_U207 ( .A1(u5_mult_82_FS_1_n179), .A2(
        u5_mult_82_FS_1_n183), .ZN(u5_mult_82_FS_1_n172) );
  NAND2_X4 u5_mult_82_FS_1_U206 ( .A1(u5_mult_82_FS_1_n726), .A2(
        u5_mult_82_FS_1_n727), .ZN(u5_mult_82_FS_1_n216) );
  OAI21_X1 u5_mult_82_FS_1_U205 ( .B1(u5_mult_82_FS_1_n238), .B2(
        u5_mult_82_FS_1_n600), .A(u5_mult_82_FS_1_n239), .ZN(
        u5_mult_82_FS_1_n231) );
  NAND2_X2 u5_mult_82_FS_1_U204 ( .A1(u5_mult_82_FS_1_n592), .A2(
        u5_mult_82_FS_1_n105), .ZN(u5_mult_82_FS_1_n590) );
  NAND2_X4 u5_mult_82_FS_1_U203 ( .A1(u5_mult_82_FS_1_n291), .A2(
        u5_mult_82_FS_1_n292), .ZN(u5_mult_82_FS_1_n290) );
  NAND3_X2 u5_mult_82_FS_1_U202 ( .A1(u5_mult_82_FS_1_n77), .A2(
        u5_mult_82_FS_1_n76), .A3(u5_mult_82_FS_1_n75), .ZN(
        u5_mult_82_FS_1_n73) );
  INV_X8 u5_mult_82_FS_1_U201 ( .A(u5_mult_82_FS_1_n554), .ZN(
        u5_mult_82_FS_1_n83) );
  INV_X8 u5_mult_82_FS_1_U200 ( .A(u5_mult_82_FS_1_n83), .ZN(
        u5_mult_82_FS_1_n150) );
  INV_X8 u5_mult_82_FS_1_U199 ( .A(u5_mult_82_FS_1_n104), .ZN(
        u5_mult_82_FS_1_n100) );
  INV_X1 u5_mult_82_FS_1_U198 ( .A(u5_mult_82_FS_1_n100), .ZN(
        u5_mult_82_FS_1_n24) );
  INV_X2 u5_mult_82_FS_1_U197 ( .A(u5_mult_82_FS_1_n463), .ZN(
        u5_mult_82_FS_1_n469) );
  NOR2_X1 u5_mult_82_FS_1_U196 ( .A1(u5_mult_82_FS_1_n462), .A2(
        u5_mult_82_FS_1_n463), .ZN(u5_mult_82_FS_1_n461) );
  AOI21_X4 u5_mult_82_FS_1_U195 ( .B1(u5_mult_82_FS_1_n256), .B2(
        u5_mult_82_FS_1_n250), .A(u5_mult_82_FS_1_n257), .ZN(
        u5_mult_82_FS_1_n247) );
  INV_X1 u5_mult_82_FS_1_U194 ( .A(u5_mult_82_FS_1_n459), .ZN(
        u5_mult_82_FS_1_n468) );
  INV_X4 u5_mult_82_FS_1_U193 ( .A(u5_mult_82_FS_1_n370), .ZN(
        u5_mult_82_FS_1_n564) );
  NAND3_X2 u5_mult_82_FS_1_U192 ( .A1(u5_mult_82_FS_1_n633), .A2(
        u5_mult_82_FS_1_n632), .A3(u5_mult_82_FS_1_n631), .ZN(
        u5_mult_82_FS_1_n463) );
  NAND2_X2 u5_mult_82_FS_1_U191 ( .A1(u5_mult_82_FS_1_n63), .A2(
        u5_mult_82_FS_1_n288), .ZN(u5_mult_82_FS_1_n286) );
  INV_X8 u5_mult_82_FS_1_U190 ( .A(u5_mult_82_FS_1_n84), .ZN(
        u5_mult_82_FS_1_n228) );
  INV_X8 u5_mult_82_FS_1_U189 ( .A(u5_mult_82_FS_1_n228), .ZN(
        u5_mult_82_FS_1_n23) );
  OR2_X2 u5_mult_82_FS_1_U188 ( .A1(u5_mult_82_FS_1_n343), .A2(
        u5_mult_82_FS_1_n357), .ZN(u5_mult_82_FS_1_n355) );
  NOR2_X2 u5_mult_82_FS_1_U187 ( .A1(u5_mult_82_FS_1_n419), .A2(
        u5_mult_82_FS_1_n121), .ZN(u5_mult_82_FS_1_n414) );
  NOR2_X2 u5_mult_82_FS_1_U186 ( .A1(u5_mult_82_FS_1_n120), .A2(
        u5_mult_82_FS_1_n121), .ZN(u5_mult_82_FS_1_n119) );
  NOR2_X2 u5_mult_82_FS_1_U185 ( .A1(u5_mult_82_FS_1_n630), .A2(
        u5_mult_82_FS_1_n121), .ZN(u5_mult_82_FS_1_n629) );
  NOR2_X2 u5_mult_82_FS_1_U184 ( .A1(u5_mult_82_FS_1_n651), .A2(
        u5_mult_82_FS_1_n501), .ZN(u5_mult_82_FS_1_n649) );
  OAI211_X2 u5_mult_82_FS_1_U183 ( .C1(u5_mult_82_CLA_SUM[60]), .C2(
        u5_mult_82_n576), .A(u5_mult_82_n573), .B(u5_mult_82_FS_1_n50), .ZN(
        u5_mult_82_FS_1_n631) );
  OAI21_X2 u5_mult_82_FS_1_U182 ( .B1(u5_mult_82_FS_1_n560), .B2(
        u5_mult_82_FS_1_n561), .A(u5_mult_82_FS_1_n562), .ZN(
        u5_mult_82_FS_1_n20) );
  NOR2_X4 u5_mult_82_FS_1_U181 ( .A1(u5_mult_82_n589), .A2(u5_mult_82_n5651), 
        .ZN(u5_mult_82_FS_1_n19) );
  NAND2_X2 u5_mult_82_FS_1_U180 ( .A1(u5_mult_82_FS_1_n440), .A2(
        u5_mult_82_FS_1_n123), .ZN(u5_mult_82_FS_1_n439) );
  INV_X8 u5_mult_82_FS_1_U179 ( .A(u5_mult_82_FS_1_n123), .ZN(
        u5_mult_82_FS_1_n283) );
  NAND3_X2 u5_mult_82_FS_1_U178 ( .A1(u5_mult_82_FS_1_n225), .A2(
        u5_mult_82_FS_1_n83), .A3(u5_mult_82_FS_1_n226), .ZN(
        u5_mult_82_FS_1_n227) );
  NAND2_X1 u5_mult_82_FS_1_U177 ( .A1(u5_mult_82_FS_1_n232), .A2(
        u5_mult_82_FS_1_n225), .ZN(u5_mult_82_FS_1_n235) );
  OAI21_X4 u5_mult_82_FS_1_U176 ( .B1(u5_mult_82_FS_1_n366), .B2(
        u5_mult_82_FS_1_n367), .A(u5_mult_82_FS_1_n368), .ZN(
        u5_mult_82_FS_1_n331) );
  NAND2_X4 u5_mult_82_FS_1_U175 ( .A1(u5_mult_82_FS_1_n330), .A2(
        u5_mult_82_FS_1_n331), .ZN(u5_mult_82_FS_1_n325) );
  INV_X1 u5_mult_82_FS_1_U174 ( .A(u5_mult_82_FS_1_n383), .ZN(
        u5_mult_82_FS_1_n17) );
  INV_X8 u5_mult_82_FS_1_U173 ( .A(u5_mult_82_FS_1_n297), .ZN(
        u5_mult_82_FS_1_n312) );
  NAND2_X4 u5_mult_82_FS_1_U172 ( .A1(u5_mult_82_FS_1_n313), .A2(
        u5_mult_82_FS_1_n22), .ZN(u5_mult_82_FS_1_n297) );
  INV_X4 u5_mult_82_FS_1_U171 ( .A(u5_mult_82_FS_1_n16), .ZN(
        u5_mult_82_FS_1_n176) );
  NOR2_X4 u5_mult_82_FS_1_U170 ( .A1(u5_mult_82_n596), .A2(
        u5_mult_82_CLA_SUM[92]), .ZN(u5_mult_82_FS_1_n16) );
  NAND2_X2 u5_mult_82_FS_1_U169 ( .A1(u5_mult_82_FS_1_n228), .A2(
        u5_mult_82_FS_1_n268), .ZN(u5_mult_82_FS_1_n259) );
  NAND3_X2 u5_mult_82_FS_1_U168 ( .A1(u5_mult_82_FS_1_n633), .A2(
        u5_mult_82_FS_1_n632), .A3(u5_mult_82_FS_1_n631), .ZN(
        u5_mult_82_FS_1_n15) );
  INV_X8 u5_mult_82_FS_1_U167 ( .A(u5_mult_82_FS_1_n587), .ZN(
        u5_mult_82_FS_1_n525) );
  INV_X8 u5_mult_82_FS_1_U166 ( .A(u5_mult_82_FS_1_n338), .ZN(
        u5_mult_82_FS_1_n332) );
  NOR3_X2 u5_mult_82_FS_1_U165 ( .A1(u5_mult_82_FS_1_n344), .A2(
        u5_mult_82_FS_1_n345), .A3(u5_mult_82_FS_1_n346), .ZN(
        u5_mult_82_FS_1_n335) );
  NAND2_X2 u5_mult_82_FS_1_U164 ( .A1(u5_mult_82_FS_1_n40), .A2(
        u5_mult_82_FS_1_n337), .ZN(u5_mult_82_FS_1_n336) );
  NAND3_X4 u5_mult_82_FS_1_U163 ( .A1(u5_mult_82_FS_1_n592), .A2(
        u5_mult_82_FS_1_n85), .A3(u5_mult_82_FS_1_n100), .ZN(
        u5_mult_82_FS_1_n587) );
  NAND2_X4 u5_mult_82_FS_1_U162 ( .A1(u5_mult_82_FS_1_n35), .A2(
        u5_mult_82_FS_1_n55), .ZN(u5_mult_82_FS_1_n57) );
  INV_X8 u5_mult_82_FS_1_U161 ( .A(u5_mult_82_CLA_SUM[76]), .ZN(
        u5_mult_82_FS_1_n682) );
  INV_X2 u5_mult_82_FS_1_U160 ( .A(u5_mult_82_FS_1_n648), .ZN(
        u5_mult_82_FS_1_n646) );
  NAND2_X4 u5_mult_82_FS_1_U159 ( .A1(u5_mult_82_n590), .A2(
        u5_mult_82_CLA_SUM[87]), .ZN(u5_mult_82_FS_1_n225) );
  NAND2_X4 u5_mult_82_FS_1_U158 ( .A1(u5_mult_82_FS_1_n206), .A2(
        u5_mult_82_FS_1_n207), .ZN(u5_mult_82_FS_1_n199) );
  NAND2_X4 u5_mult_82_FS_1_U157 ( .A1(u5_mult_82_FS_1_n701), .A2(
        u5_mult_82_FS_1_n702), .ZN(u5_mult_82_FS_1_n191) );
  NOR2_X4 u5_mult_82_FS_1_U156 ( .A1(u5_mult_82_FS_1_n205), .A2(
        u5_mult_82_FS_1_n241), .ZN(u5_mult_82_FS_1_n699) );
  NAND2_X4 u5_mult_82_FS_1_U155 ( .A1(u5_mult_82_FS_1_n699), .A2(
        u5_mult_82_FS_1_n700), .ZN(u5_mult_82_FS_1_n104) );
  INV_X8 u5_mult_82_FS_1_U154 ( .A(u5_mult_82_CLA_SUM[82]), .ZN(
        u5_mult_82_FS_1_n605) );
  INV_X1 u5_mult_82_FS_1_U153 ( .A(u5_mult_82_FS_1_n90), .ZN(
        u5_mult_82_FS_1_n96) );
  NOR2_X2 u5_mult_82_FS_1_U152 ( .A1(u5_mult_82_CLA_SUM[83]), .A2(
        u5_mult_82_CLA_CARRY[82]), .ZN(u5_mult_82_FS_1_n270) );
  OAI21_X2 u5_mult_82_FS_1_U151 ( .B1(u5_mult_82_FS_1_n615), .B2(
        u5_mult_82_FS_1_n616), .A(u5_mult_82_FS_1_n617), .ZN(
        u5_mult_82_FS_1_n203) );
  NAND2_X2 u5_mult_82_FS_1_U150 ( .A1(u5_mult_82_FS_1_n68), .A2(
        u5_mult_82_FS_1_n69), .ZN(u5_mult_82_FS_1_n56) );
  INV_X2 u5_mult_82_FS_1_U149 ( .A(u5_mult_82_FS_1_n311), .ZN(
        u5_mult_82_FS_1_n21) );
  INV_X4 u5_mult_82_FS_1_U148 ( .A(u5_mult_82_CLA_SUM[75]), .ZN(
        u5_mult_82_FS_1_n684) );
  NAND2_X2 u5_mult_82_FS_1_U147 ( .A1(u5_mult_82_n595), .A2(
        u5_mult_82_CLA_SUM[75]), .ZN(u5_mult_82_FS_1_n347) );
  INV_X16 u5_mult_82_FS_1_U146 ( .A(u5_mult_82_FS_1_n218), .ZN(
        u5_mult_82_FS_1_n121) );
  INV_X4 u5_mult_82_FS_1_U145 ( .A(u5_mult_82_FS_1_n265), .ZN(
        u5_mult_82_FS_1_n520) );
  NAND2_X4 u5_mult_82_FS_1_U144 ( .A1(u5_mult_82_FS_1_n538), .A2(
        u5_mult_82_FS_1_n537), .ZN(u5_mult_82_FS_1_n533) );
  NAND2_X2 u5_mult_82_FS_1_U143 ( .A1(u5_mult_82_n589), .A2(u5_mult_82_n5651), 
        .ZN(u5_mult_82_FS_1_n123) );
  INV_X1 u5_mult_82_FS_1_U142 ( .A(u5_mult_82_FS_1_n19), .ZN(
        u5_mult_82_FS_1_n440) );
  INV_X4 u5_mult_82_FS_1_U141 ( .A(u5_mult_82_FS_1_n331), .ZN(
        u5_mult_82_FS_1_n361) );
  INV_X1 u5_mult_82_FS_1_U140 ( .A(u5_mult_82_FS_1_n363), .ZN(
        u5_mult_82_FS_1_n339) );
  INV_X8 u5_mult_82_FS_1_U139 ( .A(u5_mult_82_FS_1_n588), .ZN(
        u5_mult_82_FS_1_n531) );
  INV_X4 u5_mult_82_FS_1_U138 ( .A(u5_mult_82_FS_1_n14), .ZN(
        u5_mult_82_FS_1_n323) );
  NOR2_X4 u5_mult_82_FS_1_U137 ( .A1(u5_mult_82_CLA_SUM[78]), .A2(
        u5_mult_82_n585), .ZN(u5_mult_82_FS_1_n14) );
  XNOR2_X2 u5_mult_82_FS_1_U136 ( .A(u5_mult_82_FS_1_n32), .B(
        u5_mult_82_FS_1_n551), .ZN(u5_N102) );
  NAND2_X2 u5_mult_82_FS_1_U135 ( .A1(u5_mult_82_FS_1_n60), .A2(
        u5_mult_82_FS_1_n61), .ZN(u5_N89) );
  XNOR2_X2 u5_mult_82_FS_1_U134 ( .A(u5_mult_82_FS_1_n11), .B(
        u5_mult_82_FS_1_n40), .ZN(u5_N66) );
  NAND2_X2 u5_mult_82_FS_1_U133 ( .A1(u5_mult_82_FS_1_n312), .A2(
        u5_mult_82_FS_1_n40), .ZN(u5_mult_82_FS_1_n309) );
  OAI21_X2 u5_mult_82_FS_1_U132 ( .B1(u5_mult_82_FS_1_n14), .B2(
        u5_mult_82_FS_1_n314), .A(u5_mult_82_FS_1_n317), .ZN(
        u5_mult_82_FS_1_n324) );
  OAI21_X2 u5_mult_82_FS_1_U131 ( .B1(u5_mult_82_FS_1_n343), .B2(
        u5_mult_82_FS_1_n348), .A(u5_mult_82_FS_1_n347), .ZN(
        u5_mult_82_FS_1_n354) );
  NAND2_X2 u5_mult_82_FS_1_U130 ( .A1(u5_mult_82_FS_1_n117), .A2(
        u5_mult_82_FS_1_n149), .ZN(u5_mult_82_FS_1_n116) );
  OAI21_X2 u5_mult_82_FS_1_U129 ( .B1(u5_mult_82_FS_1_n473), .B2(
        u5_mult_82_FS_1_n474), .A(u5_mult_82_FS_1_n475), .ZN(
        u5_mult_82_FS_1_n472) );
  OAI21_X2 u5_mult_82_FS_1_U128 ( .B1(u5_mult_82_FS_1_n505), .B2(
        u5_mult_82_FS_1_n506), .A(u5_mult_82_FS_1_n507), .ZN(
        u5_mult_82_FS_1_n504) );
  AND2_X2 u5_mult_82_FS_1_U127 ( .A1(u5_mult_82_FS_1_n507), .A2(
        u5_mult_82_FS_1_n511), .ZN(u5_mult_82_FS_1_n13) );
  XNOR2_X2 u5_mult_82_FS_1_U126 ( .A(u5_mult_82_FS_1_n505), .B(
        u5_mult_82_FS_1_n13), .ZN(u5_N56) );
  AND2_X2 u5_mult_82_FS_1_U125 ( .A1(u5_mult_82_FS_1_n143), .A2(
        u5_mult_82_FS_1_n158), .ZN(u5_mult_82_FS_1_n12) );
  INV_X4 u5_mult_82_FS_1_U124 ( .A(u5_mult_82_FS_1_n21), .ZN(
        u5_mult_82_FS_1_n22) );
  INV_X4 u5_mult_82_FS_1_U123 ( .A(u5_mult_82_FS_1_n426), .ZN(
        u5_mult_82_FS_1_n418) );
  OR2_X4 u5_mult_82_FS_1_U122 ( .A1(u5_mult_82_FS_1_n430), .A2(
        u5_mult_82_FS_1_n437), .ZN(u5_mult_82_FS_1_n11) );
  OR2_X4 u5_mult_82_FS_1_U121 ( .A1(u5_mult_82_FS_1_n378), .A2(
        u5_mult_82_FS_1_n379), .ZN(u5_mult_82_FS_1_n10) );
  OR2_X4 u5_mult_82_FS_1_U120 ( .A1(u5_mult_82_FS_1_n343), .A2(
        u5_mult_82_FS_1_n342), .ZN(u5_mult_82_FS_1_n9) );
  NOR2_X2 u5_mult_82_FS_1_U119 ( .A1(u5_mult_82_FS_1_n416), .A2(
        u5_mult_82_FS_1_n422), .ZN(u5_mult_82_FS_1_n427) );
  NOR2_X2 u5_mult_82_FS_1_U118 ( .A1(u5_mult_82_FS_1_n303), .A2(
        u5_mult_82_FS_1_n315), .ZN(u5_mult_82_FS_1_n308) );
  NOR2_X2 u5_mult_82_FS_1_U117 ( .A1(u5_mult_82_FS_1_n269), .A2(
        u5_mult_82_FS_1_n3), .ZN(u5_mult_82_FS_1_n275) );
  NOR2_X2 u5_mult_82_FS_1_U116 ( .A1(u5_mult_82_FS_1_n481), .A2(
        u5_mult_82_FS_1_n482), .ZN(u5_mult_82_FS_1_n480) );
  INV_X8 u5_mult_82_FS_1_U115 ( .A(u5_mult_82_FS_1_n296), .ZN(
        u5_mult_82_FS_1_n320) );
  OAI21_X2 u5_mult_82_FS_1_U114 ( .B1(u5_mult_82_FS_1_n264), .B2(
        u5_mult_82_FS_1_n265), .A(u5_mult_82_FS_1_n266), .ZN(
        u5_mult_82_FS_1_n255) );
  AOI21_X2 u5_mult_82_FS_1_U113 ( .B1(u5_mult_82_FS_1_n622), .B2(
        u5_mult_82_FS_1_n623), .A(u5_mult_82_FS_1_n624), .ZN(
        u5_mult_82_FS_1_n589) );
  NAND2_X2 u5_mult_82_FS_1_U112 ( .A1(u5_mult_82_FS_1_n142), .A2(
        u5_mult_82_FS_1_n156), .ZN(u5_mult_82_FS_1_n66) );
  NOR2_X1 u5_mult_82_FS_1_U111 ( .A1(u5_mult_82_FS_1_n283), .A2(
        u5_mult_82_FS_1_n416), .ZN(u5_mult_82_FS_1_n420) );
  NAND3_X2 u5_mult_82_FS_1_U110 ( .A1(u5_mult_82_n581), .A2(
        u5_mult_82_CLA_SUM[66]), .A3(u5_mult_82_FS_1_n418), .ZN(
        u5_mult_82_FS_1_n585) );
  NOR2_X1 u5_mult_82_FS_1_U109 ( .A1(u5_mult_82_FS_1_n429), .A2(
        u5_mult_82_FS_1_n431), .ZN(u5_mult_82_FS_1_n422) );
  NOR2_X2 u5_mult_82_FS_1_U108 ( .A1(u5_mult_82_FS_1_n526), .A2(
        u5_mult_82_FS_1_n527), .ZN(u5_mult_82_FS_1_n516) );
  NOR2_X2 u5_mult_82_FS_1_U107 ( .A1(u5_mult_82_FS_1_n124), .A2(
        u5_mult_82_FS_1_n65), .ZN(u5_mult_82_FS_1_n151) );
  AOI211_X2 u5_mult_82_FS_1_U106 ( .C1(u5_mult_82_FS_1_n148), .C2(
        u5_mult_82_FS_1_n149), .A(u5_mult_82_FS_1_n150), .B(
        u5_mult_82_FS_1_n228), .ZN(u5_mult_82_FS_1_n140) );
  NOR2_X2 u5_mult_82_FS_1_U105 ( .A1(u5_mult_82_FS_1_n301), .A2(
        u5_mult_82_FS_1_n302), .ZN(u5_mult_82_FS_1_n298) );
  NAND3_X2 u5_mult_82_FS_1_U104 ( .A1(u5_mult_82_FS_1_n523), .A2(
        u5_mult_82_FS_1_n524), .A3(u5_mult_82_FS_1_n525), .ZN(
        u5_mult_82_FS_1_n522) );
  INV_X2 u5_mult_82_FS_1_U103 ( .A(u5_mult_82_FS_1_n444), .ZN(
        u5_mult_82_FS_1_n643) );
  NOR2_X2 u5_mult_82_FS_1_U102 ( .A1(u5_mult_82_FS_1_n625), .A2(
        u5_mult_82_FS_1_n626), .ZN(u5_mult_82_FS_1_n622) );
  NOR3_X2 u5_mult_82_FS_1_U101 ( .A1(u5_mult_82_FS_1_n648), .A2(
        u5_mult_82_FS_1_n474), .A3(u5_mult_82_FS_1_n470), .ZN(
        u5_mult_82_FS_1_n650) );
  NAND4_X2 u5_mult_82_FS_1_U100 ( .A1(u5_mult_82_FS_1_n418), .A2(
        u5_mult_82_CLA_SUM[67]), .A3(u5_mult_82_CLA_CARRY[66]), .A4(
        u5_mult_82_FS_1_n584), .ZN(u5_mult_82_FS_1_n582) );
  NOR2_X2 u5_mult_82_FS_1_U99 ( .A1(u5_mult_82_CLA_SUM[60]), .A2(
        u5_mult_82_n576), .ZN(u5_mult_82_FS_1_n637) );
  NOR2_X2 u5_mult_82_FS_1_U98 ( .A1(u5_mult_82_FS_1_n50), .A2(u5_mult_82_n573), 
        .ZN(u5_mult_82_FS_1_n636) );
  NOR2_X1 u5_mult_82_FS_1_U97 ( .A1(u5_mult_82_FS_1_n19), .A2(
        u5_mult_82_FS_1_n34), .ZN(u5_mult_82_FS_1_n642) );
  INV_X4 u5_mult_82_FS_1_U96 ( .A(u5_mult_82_FS_1_n573), .ZN(
        u5_mult_82_FS_1_n370) );
  NOR2_X2 u5_mult_82_FS_1_U95 ( .A1(u5_mult_82_FS_1_n459), .A2(
        u5_mult_82_FS_1_n280), .ZN(u5_mult_82_FS_1_n458) );
  NAND2_X4 u5_mult_82_FS_1_U94 ( .A1(u5_mult_82_FS_1_n634), .A2(
        u5_mult_82_FS_1_n635), .ZN(u5_mult_82_FS_1_n633) );
  NAND2_X2 u5_mult_82_FS_1_U93 ( .A1(u5_mult_82_FS_1_n332), .A2(
        u5_mult_82_FS_1_n363), .ZN(u5_mult_82_FS_1_n357) );
  NOR2_X2 u5_mult_82_FS_1_U92 ( .A1(u5_mult_82_FS_1_n50), .A2(u5_mult_82_n573), 
        .ZN(u5_mult_82_FS_1_n651) );
  INV_X4 u5_mult_82_FS_1_U91 ( .A(u5_mult_82_FS_1_n600), .ZN(
        u5_mult_82_FS_1_n244) );
  NAND2_X4 u5_mult_82_FS_1_U90 ( .A1(u5_mult_82_CLA_SUM[70]), .A2(
        u5_mult_82_n577), .ZN(u5_mult_82_FS_1_n577) );
  INV_X2 u5_mult_82_FS_1_U89 ( .A(u5_mult_82_FS_1_n403), .ZN(
        u5_mult_82_FS_1_n8) );
  NAND2_X2 u5_mult_82_FS_1_U88 ( .A1(u5_mult_82_FS_1_n67), .A2(
        u5_mult_82_FS_1_n157), .ZN(u5_mult_82_FS_1_n155) );
  NAND2_X2 u5_mult_82_FS_1_U87 ( .A1(u5_mult_82_FS_1_n581), .A2(
        u5_mult_82_FS_1_n582), .ZN(u5_mult_82_FS_1_n580) );
  INV_X8 u5_mult_82_FS_1_U86 ( .A(u5_mult_82_FS_1_n81), .ZN(
        u5_mult_82_FS_1_n149) );
  AND2_X2 u5_mult_82_FS_1_U85 ( .A1(u5_mult_82_FS_1_n303), .A2(
        u5_mult_82_FS_1_n292), .ZN(u5_mult_82_FS_1_n7) );
  NAND2_X4 u5_mult_82_FS_1_U84 ( .A1(u5_mult_82_n582), .A2(
        u5_mult_82_CLA_SUM[77]), .ZN(u5_mult_82_FS_1_n33) );
  NAND2_X2 u5_mult_82_FS_1_U83 ( .A1(u5_mult_82_FS_1_n122), .A2(
        u5_mult_82_FS_1_n123), .ZN(u5_mult_82_FS_1_n630) );
  OR2_X1 u5_mult_82_FS_1_U82 ( .A1(u5_mult_82_FS_1_n488), .A2(
        u5_mult_82_FS_1_n474), .ZN(u5_mult_82_FS_1_n6) );
  INV_X4 u5_mult_82_FS_1_U81 ( .A(u5_mult_82_FS_1_n205), .ZN(
        u5_mult_82_FS_1_n207) );
  OR2_X1 u5_mult_82_FS_1_U80 ( .A1(u5_mult_82_FS_1_n502), .A2(
        u5_mult_82_FS_1_n487), .ZN(u5_mult_82_FS_1_n5) );
  NOR2_X4 u5_mult_82_FS_1_U79 ( .A1(u5_mult_82_FS_1_n188), .A2(
        u5_mult_82_FS_1_n16), .ZN(u5_mult_82_FS_1_n613) );
  NOR2_X4 u5_mult_82_FS_1_U78 ( .A1(u5_mult_82_FS_1_n136), .A2(
        u5_mult_82_FS_1_n129), .ZN(u5_mult_82_FS_1_n135) );
  CLKBUF_X3 u5_mult_82_FS_1_U77 ( .A(u5_mult_82_FS_1_n164), .Z(
        u5_mult_82_FS_1_n18) );
  NAND2_X4 u5_mult_82_FS_1_U76 ( .A1(u5_mult_82_FS_1_n730), .A2(
        u5_mult_82_FS_1_n731), .ZN(u5_mult_82_FS_1_n202) );
  NAND2_X4 u5_mult_82_FS_1_U75 ( .A1(u5_mult_82_FS_1_n202), .A2(
        u5_mult_82_FS_1_n210), .ZN(u5_mult_82_FS_1_n209) );
  OAI211_X4 u5_mult_82_FS_1_U74 ( .C1(u5_mult_82_FS_1_n211), .C2(
        u5_mult_82_FS_1_n212), .A(u5_mult_82_FS_1_n214), .B(
        u5_mult_82_FS_1_n213), .ZN(u5_mult_82_FS_1_n208) );
  INV_X4 u5_mult_82_FS_1_U73 ( .A(u5_mult_82_FS_1_n395), .ZN(
        u5_mult_82_FS_1_n383) );
  NOR2_X2 u5_mult_82_FS_1_U72 ( .A1(u5_mult_82_CLA_SUM[82]), .A2(
        u5_mult_82_CLA_CARRY[81]), .ZN(u5_mult_82_FS_1_n271) );
  NOR2_X4 u5_mult_82_FS_1_U71 ( .A1(u5_mult_82_CLA_SUM[82]), .A2(
        u5_mult_82_CLA_CARRY[81]), .ZN(u5_mult_82_FS_1_n3) );
  INV_X2 u5_mult_82_FS_1_U70 ( .A(u5_mult_82_FS_1_n475), .ZN(
        u5_mult_82_FS_1_n488) );
  AND2_X4 u5_mult_82_FS_1_U69 ( .A1(u5_mult_82_FS_1_n475), .A2(
        u5_mult_82_FS_1_n478), .ZN(u5_mult_82_FS_1_n632) );
  NAND2_X2 u5_mult_82_FS_1_U68 ( .A1(u5_mult_82_FS_1_n47), .A2(
        u5_mult_82_FS_1_n498), .ZN(u5_mult_82_FS_1_n496) );
  NAND2_X1 u5_mult_82_FS_1_U67 ( .A1(u5_mult_82_FS_1_n460), .A2(
        u5_mult_82_FS_1_n461), .ZN(u5_mult_82_FS_1_n456) );
  NAND2_X4 u5_mult_82_FS_1_U66 ( .A1(u5_mult_82_FS_1_n493), .A2(
        u5_mult_82_FS_1_n460), .ZN(u5_mult_82_FS_1_n492) );
  INV_X8 u5_mult_82_FS_1_U65 ( .A(u5_mult_82_FS_1_n492), .ZN(
        u5_mult_82_FS_1_n466) );
  OAI21_X2 u5_mult_82_FS_1_U64 ( .B1(u5_mult_82_FS_1_n466), .B2(
        u5_mult_82_FS_1_n487), .A(u5_mult_82_FS_1_n484), .ZN(
        u5_mult_82_FS_1_n489) );
  OAI21_X2 u5_mult_82_FS_1_U63 ( .B1(u5_mult_82_FS_1_n466), .B2(
        u5_mult_82_FS_1_n467), .A(u5_mult_82_FS_1_n468), .ZN(
        u5_mult_82_FS_1_n465) );
  INV_X2 u5_mult_82_FS_1_U62 ( .A(u5_mult_82_FS_1_n509), .ZN(
        u5_mult_82_FS_1_n644) );
  NAND2_X2 u5_mult_82_FS_1_U61 ( .A1(u5_mult_82_FS_1_n509), .A2(
        u5_mult_82_FS_1_n501), .ZN(u5_mult_82_FS_1_n503) );
  NAND3_X2 u5_mult_82_FS_1_U60 ( .A1(u5_mult_82_FS_1_n509), .A2(
        u5_mult_82_n579), .A3(u5_mult_82_CLA_SUM[56]), .ZN(
        u5_mult_82_FS_1_n500) );
  INV_X2 u5_mult_82_FS_1_U59 ( .A(u5_mult_82_FS_1_n499), .ZN(
        u5_mult_82_FS_1_n495) );
  INV_X4 u5_mult_82_FS_1_U58 ( .A(u5_mult_82_FS_1_n508), .ZN(
        u5_mult_82_FS_1_n505) );
  OR2_X2 u5_mult_82_FS_1_U57 ( .A1(u5_mult_82_FS_1_n513), .A2(
        u5_mult_82_FS_1_n499), .ZN(u5_mult_82_FS_1_n4) );
  INV_X2 u5_mult_82_FS_1_U56 ( .A(u5_mult_82_FS_1_n498), .ZN(
        u5_mult_82_FS_1_n513) );
  NAND2_X4 u5_mult_82_FS_1_U55 ( .A1(u5_mult_82_FS_1_n151), .A2(
        u5_mult_82_FS_1_n152), .ZN(u5_mult_82_FS_1_n148) );
  INV_X2 u5_mult_82_FS_1_U54 ( .A(u5_mult_82_n1075), .ZN(u5_mult_82_FS_1_n733)
         );
  INV_X8 u5_mult_82_FS_1_U53 ( .A(u5_mult_82_CLA_SUM[72]), .ZN(
        u5_mult_82_FS_1_n678) );
  NAND2_X4 u5_mult_82_FS_1_U52 ( .A1(u5_mult_82_FS_1_n362), .A2(
        u5_mult_82_FS_1_n347), .ZN(u5_mult_82_FS_1_n570) );
  OAI21_X4 u5_mult_82_FS_1_U51 ( .B1(u5_mult_82_CLA_SUM[83]), .B2(
        u5_mult_82_CLA_CARRY[82]), .A(u5_mult_82_CLA_CARRY[81]), .ZN(
        u5_mult_82_FS_1_n604) );
  INV_X8 u5_mult_82_FS_1_U50 ( .A(u5_mult_82_FS_1_n250), .ZN(
        u5_mult_82_FS_1_n252) );
  NAND4_X1 u5_mult_82_FS_1_U49 ( .A1(u5_mult_82_FS_1_n259), .A2(
        u5_mult_82_FS_1_n255), .A3(u5_mult_82_FS_1_n258), .A4(
        u5_mult_82_FS_1_n253), .ZN(u5_mult_82_FS_1_n263) );
  NOR2_X4 u5_mult_82_FS_1_U48 ( .A1(u5_mult_82_FS_1_n574), .A2(
        u5_mult_82_FS_1_n575), .ZN(u5_mult_82_FS_1_n573) );
  NAND2_X4 u5_mult_82_FS_1_U47 ( .A1(u5_mult_82_FS_1_n369), .A2(
        u5_mult_82_FS_1_n330), .ZN(u5_mult_82_FS_1_n565) );
  INV_X8 u5_mult_82_FS_1_U46 ( .A(u5_mult_82_CLA_SUM[73]), .ZN(
        u5_mult_82_FS_1_n676) );
  NOR2_X4 u5_mult_82_FS_1_U45 ( .A1(u5_mult_82_FS_1_n607), .A2(
        u5_mult_82_FS_1_n166), .ZN(u5_mult_82_FS_1_n609) );
  OAI21_X2 u5_mult_82_FS_1_U44 ( .B1(u5_mult_82_FS_1_n89), .B2(
        u5_mult_82_FS_1_n24), .A(u5_mult_82_FS_1_n98), .ZN(
        u5_mult_82_FS_1_n103) );
  INV_X2 u5_mult_82_FS_1_U43 ( .A(u5_mult_82_FS_1_n286), .ZN(
        u5_mult_82_FS_1_n37) );
  NAND2_X2 u5_mult_82_FS_1_U42 ( .A1(u5_mult_82_FS_1_n190), .A2(
        u5_mult_82_FS_1_n191), .ZN(u5_mult_82_FS_1_n181) );
  NAND2_X4 u5_mult_82_FS_1_U41 ( .A1(u5_mult_82_FS_1_n181), .A2(
        u5_mult_82_FS_1_n182), .ZN(u5_mult_82_FS_1_n180) );
  NAND2_X1 u5_mult_82_FS_1_U40 ( .A1(u5_mult_82_FS_1_n198), .A2(
        u5_mult_82_FS_1_n197), .ZN(u5_mult_82_FS_1_n200) );
  INV_X8 u5_mult_82_FS_1_U39 ( .A(u5_mult_82_FS_1_n82), .ZN(
        u5_mult_82_FS_1_n80) );
  NAND3_X1 u5_mult_82_FS_1_U38 ( .A1(u5_mult_82_FS_1_n149), .A2(
        u5_mult_82_FS_1_n519), .A3(u5_mult_82_FS_1_n82), .ZN(
        u5_mult_82_FS_1_n517) );
  NAND2_X4 u5_mult_82_FS_1_U37 ( .A1(u5_mult_82_FS_1_n332), .A2(
        u5_mult_82_FS_1_n330), .ZN(u5_mult_82_FS_1_n326) );
  NAND2_X1 u5_mult_82_FS_1_U36 ( .A1(u5_mult_82_n594), .A2(
        u5_mult_82_CLA_SUM[61]), .ZN(u5_mult_82_FS_1_n478) );
  NOR2_X4 u5_mult_82_FS_1_U35 ( .A1(u5_mult_82_FS_1_n577), .A2(
        u5_mult_82_FS_1_n578), .ZN(u5_mult_82_FS_1_n574) );
  NAND2_X2 u5_mult_82_FS_1_U34 ( .A1(u5_mult_82_FS_1_n451), .A2(
        u5_mult_82_FS_1_n452), .ZN(u5_mult_82_FS_1_n454) );
  NAND3_X4 u5_mult_82_FS_1_U33 ( .A1(u5_mult_82_FS_1_n290), .A2(
        u5_mult_82_FS_1_n289), .A3(u5_mult_82_FS_1_n287), .ZN(
        u5_mult_82_FS_1_n62) );
  NAND3_X2 u5_mult_82_FS_1_U32 ( .A1(u5_mult_82_FS_1_n292), .A2(
        u5_mult_82_FS_1_n312), .A3(u5_mult_82_FS_1_n296), .ZN(
        u5_mult_82_FS_1_n288) );
  NOR2_X4 u5_mult_82_FS_1_U31 ( .A1(u5_mult_82_FS_1_n386), .A2(
        u5_mult_82_FS_1_n320), .ZN(u5_mult_82_FS_1_n377) );
  NOR2_X2 u5_mult_82_FS_1_U30 ( .A1(u5_mult_82_FS_1_n320), .A2(
        u5_mult_82_FS_1_n355), .ZN(u5_mult_82_FS_1_n353) );
  INV_X4 u5_mult_82_FS_1_U29 ( .A(u5_mult_82_FS_1_n48), .ZN(
        u5_mult_82_FS_1_n49) );
  NAND4_X4 u5_mult_82_FS_1_U28 ( .A1(u5_mult_82_FS_1_n207), .A2(
        u5_mult_82_FS_1_n599), .A3(u5_mult_82_FS_1_n244), .A4(
        u5_mult_82_FS_1_n598), .ZN(u5_mult_82_FS_1_n594) );
  NAND2_X4 u5_mult_82_FS_1_U27 ( .A1(u5_mult_82_n604), .A2(
        u5_mult_82_CLA_SUM[90]), .ZN(u5_mult_82_FS_1_n197) );
  INV_X4 u5_mult_82_FS_1_U26 ( .A(u5_mult_82_FS_1_n105), .ZN(
        u5_mult_82_FS_1_n98) );
  INV_X8 u5_mult_82_FS_1_U25 ( .A(u5_mult_82_FS_1_n360), .ZN(
        u5_mult_82_FS_1_n348) );
  INV_X1 u5_mult_82_FS_1_U24 ( .A(u5_mult_82_FS_1_n367), .ZN(
        u5_mult_82_FS_1_n372) );
  INV_X4 u5_mult_82_FS_1_U23 ( .A(u5_mult_82_CLA_SUM[62]), .ZN(
        u5_mult_82_FS_1_n670) );
  OAI21_X4 u5_mult_82_FS_1_U22 ( .B1(u5_mult_82_FS_1_n585), .B2(
        u5_mult_82_FS_1_n586), .A(u5_mult_82_FS_1_n410), .ZN(
        u5_mult_82_FS_1_n579) );
  NAND2_X1 u5_mult_82_FS_1_U21 ( .A1(u5_mult_82_CLA_SUM[74]), .A2(
        u5_mult_82_n584), .ZN(u5_mult_82_FS_1_n2) );
  INV_X4 u5_mult_82_FS_1_U20 ( .A(u5_mult_82_FS_1_n194), .ZN(
        u5_mult_82_FS_1_n52) );
  NOR2_X4 u5_mult_82_FS_1_U19 ( .A1(u5_mult_82_FS_1_n252), .A2(
        u5_mult_82_FS_1_n258), .ZN(u5_mult_82_FS_1_n257) );
  NAND2_X4 u5_mult_82_FS_1_U18 ( .A1(u5_mult_82_FS_1_n73), .A2(
        u5_mult_82_FS_1_n74), .ZN(u5_mult_82_FS_1_n71) );
  NAND2_X4 u5_mult_82_FS_1_U17 ( .A1(u5_mult_82_FS_1_n317), .A2(
        u5_mult_82_FS_1_n302), .ZN(u5_mult_82_FS_1_n558) );
  INV_X8 u5_mult_82_FS_1_U16 ( .A(u5_mult_82_FS_1_n327), .ZN(
        u5_mult_82_FS_1_n316) );
  NAND3_X2 u5_mult_82_FS_1_U15 ( .A1(u5_mult_82_FS_1_n690), .A2(
        u5_mult_82_FS_1_n689), .A3(u5_mult_82_FS_1_n583), .ZN(
        u5_mult_82_FS_1_n389) );
  OAI21_X1 u5_mult_82_FS_1_U14 ( .B1(u5_mult_82_FS_1_n416), .B2(
        u5_mult_82_FS_1_n417), .A(u5_mult_82_FS_1_n583), .ZN(
        u5_mult_82_FS_1_n415) );
  OAI21_X2 u5_mult_82_FS_1_U13 ( .B1(u5_mult_82_CLA_SUM[67]), .B2(
        u5_mult_82_CLA_CARRY[66]), .A(u5_mult_82_FS_1_n584), .ZN(
        u5_mult_82_FS_1_n586) );
  NAND2_X4 u5_mult_82_FS_1_U12 ( .A1(u5_mult_82_FS_1_n221), .A2(
        u5_mult_82_FS_1_n222), .ZN(u5_mult_82_FS_1_n220) );
  INV_X1 u5_mult_82_FS_1_U11 ( .A(u5_mult_82_FS_1_n284), .ZN(
        u5_mult_82_FS_1_n1) );
  NOR2_X1 u5_mult_82_FS_1_U10 ( .A1(u5_mult_82_FS_1_n228), .A2(
        u5_mult_82_FS_1_n127), .ZN(u5_mult_82_FS_1_n115) );
  NAND2_X2 u5_mult_82_FS_1_U9 ( .A1(u5_mult_82_FS_1_n30), .A2(
        u5_mult_82_FS_1_n20), .ZN(u5_mult_82_FS_1_n160) );
  NOR2_X1 u5_mult_82_FS_1_U8 ( .A1(u5_mult_82_FS_1_n227), .A2(
        u5_mult_82_FS_1_n228), .ZN(u5_mult_82_FS_1_n211) );
  INV_X1 u5_mult_82_FS_1_U7 ( .A(u5_mult_82_FS_1_n231), .ZN(
        u5_mult_82_FS_1_n237) );
  OAI21_X1 u5_mult_82_FS_1_U6 ( .B1(u5_mult_82_FS_1_n47), .B2(
        u5_mult_82_FS_1_n499), .A(u5_mult_82_FS_1_n498), .ZN(
        u5_mult_82_FS_1_n508) );
  NAND2_X2 u5_mult_82_FS_1_U5 ( .A1(u5_mult_82_CLA_SUM[54]), .A2(
        u5_mult_82_CLA_CARRY[53]), .ZN(u5_mult_82_FS_1_n47) );
  INV_X2 u5_mult_82_FS_1_U4 ( .A(u5_mult_82_FS_1_n47), .ZN(
        u5_mult_82_FS_1_n510) );
  NAND2_X4 u5_mult_82_FS_1_U3 ( .A1(u5_mult_82_FS_1_n25), .A2(
        u5_mult_82_FS_1_n159), .ZN(u5_mult_82_FS_1_n175) );
  NOR2_X4 u5_mult_82_FS_1_U2 ( .A1(u5_mult_82_FS_1_n177), .A2(
        u5_mult_82_FS_1_n16), .ZN(u5_mult_82_FS_1_n25) );
  INV_X4 u4_sub_470_U114 ( .A(net44696), .ZN(u4_sub_470_n100) );
  NAND2_X2 u4_sub_470_U113 ( .A1(u4_exp_in_pl1_0_), .A2(u4_sub_470_n100), .ZN(
        u4_sub_470_n43) );
  INV_X4 u4_sub_470_U112 ( .A(u4_exp_in_pl1_0_), .ZN(u4_sub_470_n99) );
  NAND2_X2 u4_sub_470_U111 ( .A1(net44696), .A2(u4_sub_470_n99), .ZN(
        u4_sub_470_n92) );
  NAND2_X2 u4_sub_470_U110 ( .A1(u4_sub_470_n43), .A2(u4_sub_470_n92), .ZN(
        u4_exp_next_mi_0_) );
  INV_X4 u4_sub_470_U109 ( .A(u4_fi_ldz_mi1_5_), .ZN(u4_sub_470_n96) );
  NAND2_X2 u4_sub_470_U108 ( .A1(u4_exp_in_pl1_5_), .A2(u4_sub_470_n96), .ZN(
        u4_sub_470_n16) );
  INV_X4 u4_sub_470_U107 ( .A(u4_fi_ldz_mi1_4_), .ZN(u4_sub_470_n98) );
  NAND2_X2 u4_sub_470_U106 ( .A1(u4_exp_in_pl1_4_), .A2(u4_sub_470_n98), .ZN(
        u4_sub_470_n22) );
  NAND2_X2 u4_sub_470_U105 ( .A1(u4_sub_470_n16), .A2(u4_sub_470_n22), .ZN(
        u4_sub_470_n68) );
  INV_X4 u4_sub_470_U104 ( .A(u4_exp_in_pl1_6_), .ZN(u4_sub_470_n97) );
  NAND2_X2 u4_sub_470_U103 ( .A1(u4_fi_ldz_mi1_6_), .A2(u4_sub_470_n97), .ZN(
        u4_sub_470_n12) );
  INV_X4 u4_sub_470_U102 ( .A(u4_sub_470_n12), .ZN(u4_sub_470_n64) );
  OAI211_X2 u4_sub_470_U101 ( .C1(u4_exp_in_pl1_5_), .C2(u4_sub_470_n96), .A(
        u4_sub_470_n68), .B(u4_sub_470_n69), .ZN(u4_sub_470_n76) );
  INV_X4 u4_sub_470_U100 ( .A(u4_exp_in_pl1_5_), .ZN(u4_sub_470_n70) );
  NAND2_X2 u4_sub_470_U99 ( .A1(u4_fi_ldz_mi1_5_), .A2(u4_sub_470_n70), .ZN(
        u4_sub_470_n25) );
  INV_X4 u4_sub_470_U98 ( .A(u4_fi_ldz_2a_2_), .ZN(u4_sub_470_n95) );
  NAND2_X2 u4_sub_470_U97 ( .A1(u4_exp_in_pl1_2_), .A2(u4_sub_470_n95), .ZN(
        u4_sub_470_n30) );
  INV_X4 u4_sub_470_U96 ( .A(u4_sub_470_n30), .ZN(u4_sub_470_n93) );
  INV_X4 u4_sub_470_U95 ( .A(u4_exp_in_pl1_3_), .ZN(u4_sub_470_n94) );
  NAND2_X2 u4_sub_470_U94 ( .A1(u4_fi_ldz_mi1_3_), .A2(u4_sub_470_n94), .ZN(
        u4_sub_470_n33) );
  NAND2_X2 u4_sub_470_U93 ( .A1(u4_sub_470_n93), .A2(u4_sub_470_n33), .ZN(
        u4_sub_470_n79) );
  INV_X4 u4_sub_470_U92 ( .A(u4_sub_470_n42), .ZN(u4_sub_470_n61) );
  INV_X4 u4_sub_470_U91 ( .A(u4_exp_in_pl1_1_), .ZN(u4_sub_470_n87) );
  NAND2_X2 u4_sub_470_U90 ( .A1(u4_fi_ldz_mi1_1_), .A2(u4_sub_470_n87), .ZN(
        u4_sub_470_n39) );
  INV_X4 u4_sub_470_U89 ( .A(u4_sub_470_n33), .ZN(u4_sub_470_n56) );
  INV_X4 u4_sub_470_U88 ( .A(u4_exp_in_pl1_2_), .ZN(u4_sub_470_n91) );
  NAND2_X2 u4_sub_470_U87 ( .A1(u4_fi_ldz_2a_2_), .A2(u4_sub_470_n91), .ZN(
        u4_sub_470_n31) );
  INV_X4 u4_sub_470_U86 ( .A(u4_sub_470_n31), .ZN(u4_sub_470_n86) );
  INV_X4 u4_sub_470_U85 ( .A(u4_fi_ldz_mi1_1_), .ZN(u4_sub_470_n89) );
  NAND2_X2 u4_sub_470_U84 ( .A1(u4_exp_in_pl1_1_), .A2(u4_sub_470_n89), .ZN(
        u4_sub_470_n38) );
  NAND2_X2 u4_sub_470_U83 ( .A1(u4_sub_470_n38), .A2(u4_sub_470_n43), .ZN(
        u4_sub_470_n88) );
  INV_X4 u4_sub_470_U82 ( .A(u4_sub_470_n88), .ZN(u4_sub_470_n58) );
  NOR2_X4 u4_sub_470_U81 ( .A1(u4_sub_470_n58), .A2(u4_sub_470_n37), .ZN(
        u4_sub_470_n82) );
  INV_X4 u4_sub_470_U80 ( .A(u4_fi_ldz_mi1_3_), .ZN(u4_sub_470_n85) );
  NAND2_X2 u4_sub_470_U79 ( .A1(u4_exp_in_pl1_3_), .A2(u4_sub_470_n85), .ZN(
        u4_sub_470_n34) );
  INV_X4 u4_sub_470_U78 ( .A(u4_sub_470_n34), .ZN(u4_sub_470_n84) );
  AOI21_X4 u4_sub_470_U77 ( .B1(u4_sub_470_n82), .B2(u4_sub_470_n83), .A(
        u4_sub_470_n84), .ZN(u4_sub_470_n81) );
  NAND3_X4 u4_sub_470_U76 ( .A1(u4_sub_470_n79), .A2(u4_sub_470_n80), .A3(
        u4_sub_470_n81), .ZN(u4_sub_470_n23) );
  INV_X4 u4_sub_470_U75 ( .A(u4_exp_in_pl1_4_), .ZN(u4_sub_470_n78) );
  NAND2_X2 u4_sub_470_U74 ( .A1(u4_fi_ldz_mi1_4_), .A2(u4_sub_470_n78), .ZN(
        u4_sub_470_n24) );
  INV_X4 u4_sub_470_U73 ( .A(u4_sub_470_n20), .ZN(u4_sub_470_n62) );
  NAND4_X2 u4_sub_470_U72 ( .A1(u4_sub_470_n25), .A2(u4_sub_470_n12), .A3(
        u4_sub_470_n23), .A4(u4_sub_470_n62), .ZN(u4_sub_470_n77) );
  INV_X4 u4_sub_470_U71 ( .A(u4_fi_ldz_mi1_6_), .ZN(u4_sub_470_n18) );
  NAND4_X2 u4_sub_470_U70 ( .A1(u4_sub_470_n76), .A2(u4_sub_470_n8), .A3(
        u4_sub_470_n77), .A4(u4_sub_470_n49), .ZN(u4_sub_470_n5) );
  INV_X4 u4_sub_470_U69 ( .A(u4_sub_470_n5), .ZN(u4_sub_470_n2) );
  INV_X4 u4_sub_470_U68 ( .A(u4_sub_470_n3), .ZN(u4_sub_470_n74) );
  INV_X4 u4_sub_470_U67 ( .A(u4_sub_470_n4), .ZN(u4_sub_470_n75) );
  NOR2_X4 u4_sub_470_U66 ( .A1(u4_sub_470_n74), .A2(u4_sub_470_n75), .ZN(
        u4_sub_470_n50) );
  XNOR2_X2 u4_sub_470_U65 ( .A(u4_sub_470_n71), .B(u4_sub_470_n73), .ZN(
        u4_exp_next_mi_10_) );
  INV_X4 u4_sub_470_U64 ( .A(u4_sub_470_n72), .ZN(u4_sub_470_n71) );
  NOR2_X4 u4_sub_470_U63 ( .A1(u4_sub_470_n71), .A2(u4_sub_470_n7), .ZN(
        u4_sub_470_n65) );
  NAND2_X2 u4_sub_470_U62 ( .A1(u4_fi_ldz_mi1_5_), .A2(u4_sub_470_n70), .ZN(
        u4_sub_470_n67) );
  NAND2_X2 u4_sub_470_U61 ( .A1(u4_sub_470_n65), .A2(u4_sub_470_n66), .ZN(
        u4_sub_470_n46) );
  INV_X4 u4_sub_470_U60 ( .A(u4_sub_470_n25), .ZN(u4_sub_470_n15) );
  NAND2_X2 u4_sub_470_U59 ( .A1(u4_sub_470_n31), .A2(u4_sub_470_n33), .ZN(
        u4_sub_470_n59) );
  NAND2_X2 u4_sub_470_U58 ( .A1(u4_sub_470_n61), .A2(u4_sub_470_n39), .ZN(
        u4_sub_470_n60) );
  NAND2_X2 u4_sub_470_U57 ( .A1(u4_sub_470_n31), .A2(u4_sub_470_n33), .ZN(
        u4_sub_470_n57) );
  NOR3_X4 u4_sub_470_U56 ( .A1(u4_sub_470_n53), .A2(u4_sub_470_n54), .A3(
        u4_sub_470_n55), .ZN(u4_sub_470_n52) );
  NOR3_X4 u4_sub_470_U55 ( .A1(u4_sub_470_n46), .A2(u4_sub_470_n47), .A3(
        u4_sub_470_n48), .ZN(u4_sub_470_n44) );
  XNOR2_X2 u4_sub_470_U54 ( .A(u4_sub_470_n44), .B(u4_sub_470_n45), .ZN(
        u4_exp_next_mi_11_) );
  NAND2_X2 u4_sub_470_U53 ( .A1(u4_sub_470_n38), .A2(u4_sub_470_n39), .ZN(
        u4_sub_470_n41) );
  NAND2_X2 u4_sub_470_U52 ( .A1(u4_sub_470_n42), .A2(u4_sub_470_n43), .ZN(
        u4_sub_470_n40) );
  XNOR2_X2 u4_sub_470_U51 ( .A(u4_sub_470_n41), .B(u4_sub_470_n40), .ZN(
        u4_exp_next_mi_1_) );
  NAND2_X2 u4_sub_470_U50 ( .A1(u4_sub_470_n31), .A2(u4_sub_470_n30), .ZN(
        u4_sub_470_n35) );
  INV_X4 u4_sub_470_U49 ( .A(u4_sub_470_n40), .ZN(u4_sub_470_n36) );
  INV_X4 u4_sub_470_U48 ( .A(u4_sub_470_n39), .ZN(u4_sub_470_n37) );
  OAI21_X4 u4_sub_470_U47 ( .B1(u4_sub_470_n36), .B2(u4_sub_470_n37), .A(
        u4_sub_470_n38), .ZN(u4_sub_470_n32) );
  XNOR2_X2 u4_sub_470_U46 ( .A(u4_sub_470_n35), .B(u4_sub_470_n32), .ZN(
        u4_exp_next_mi_2_) );
  NAND2_X2 u4_sub_470_U45 ( .A1(u4_sub_470_n33), .A2(u4_sub_470_n34), .ZN(
        u4_sub_470_n27) );
  NAND2_X2 u4_sub_470_U44 ( .A1(u4_sub_470_n31), .A2(u4_sub_470_n32), .ZN(
        u4_sub_470_n29) );
  NAND2_X2 u4_sub_470_U43 ( .A1(u4_sub_470_n29), .A2(u4_sub_470_n30), .ZN(
        u4_sub_470_n28) );
  XNOR2_X2 u4_sub_470_U42 ( .A(u4_sub_470_n27), .B(u4_sub_470_n28), .ZN(
        u4_exp_next_mi_3_) );
  NAND2_X2 u4_sub_470_U41 ( .A1(u4_sub_470_n22), .A2(u4_sub_470_n24), .ZN(
        u4_sub_470_n26) );
  XNOR2_X2 u4_sub_470_U40 ( .A(u4_sub_470_n23), .B(u4_sub_470_n26), .ZN(
        u4_exp_next_mi_4_) );
  NAND2_X2 u4_sub_470_U39 ( .A1(u4_sub_470_n25), .A2(u4_sub_470_n16), .ZN(
        u4_sub_470_n19) );
  INV_X4 u4_sub_470_U38 ( .A(u4_sub_470_n24), .ZN(u4_sub_470_n20) );
  INV_X4 u4_sub_470_U37 ( .A(u4_sub_470_n23), .ZN(u4_sub_470_n21) );
  OAI21_X4 u4_sub_470_U36 ( .B1(u4_sub_470_n20), .B2(u4_sub_470_n21), .A(
        u4_sub_470_n22), .ZN(u4_sub_470_n17) );
  XNOR2_X2 u4_sub_470_U35 ( .A(u4_sub_470_n19), .B(u4_sub_470_n17), .ZN(
        u4_exp_next_mi_5_) );
  NAND2_X2 u4_sub_470_U34 ( .A1(u4_exp_in_pl1_6_), .A2(u4_sub_470_n18), .ZN(
        u4_sub_470_n9) );
  NAND2_X2 u4_sub_470_U33 ( .A1(u4_sub_470_n12), .A2(u4_sub_470_n9), .ZN(
        u4_sub_470_n13) );
  INV_X4 u4_sub_470_U32 ( .A(u4_sub_470_n17), .ZN(u4_sub_470_n14) );
  OAI21_X4 u4_sub_470_U31 ( .B1(u4_sub_470_n14), .B2(u4_sub_470_n15), .A(
        u4_sub_470_n16), .ZN(u4_sub_470_n11) );
  XNOR2_X2 u4_sub_470_U30 ( .A(u4_sub_470_n13), .B(u4_sub_470_n11), .ZN(
        u4_exp_next_mi_6_) );
  NAND2_X2 u4_sub_470_U29 ( .A1(u4_sub_470_n11), .A2(u4_sub_470_n12), .ZN(
        u4_sub_470_n10) );
  NAND2_X2 u4_sub_470_U28 ( .A1(u4_sub_470_n9), .A2(u4_sub_470_n10), .ZN(
        u4_sub_470_n6) );
  XNOR2_X2 u4_sub_470_U27 ( .A(u4_sub_470_n6), .B(u4_sub_470_n7), .ZN(
        u4_exp_next_mi_7_) );
  XNOR2_X2 u4_sub_470_U26 ( .A(u4_sub_470_n74), .B(u4_sub_470_n5), .ZN(
        u4_exp_next_mi_8_) );
  XNOR2_X2 u4_sub_470_U25 ( .A(u4_sub_470_n75), .B(u4_sub_470_n1), .ZN(
        u4_exp_next_mi_9_) );
  INV_X4 u4_sub_470_U24 ( .A(u4_exp_in_pl1_11_), .ZN(u4_sub_470_n45) );
  INV_X4 u4_sub_470_U23 ( .A(u4_sub_470_n64), .ZN(u4_sub_470_n69) );
  NAND2_X2 u4_sub_470_U22 ( .A1(u4_sub_470_n2), .A2(u4_sub_470_n3), .ZN(
        u4_sub_470_n1) );
  NAND2_X2 u4_sub_470_U21 ( .A1(u4_sub_470_n2), .A2(u4_sub_470_n50), .ZN(
        u4_sub_470_n73) );
  NAND2_X2 u4_sub_470_U20 ( .A1(u4_sub_470_n49), .A2(u4_sub_470_n50), .ZN(
        u4_sub_470_n48) );
  INV_X4 u4_sub_470_U19 ( .A(u4_sub_470_n92), .ZN(u4_sub_470_n42) );
  NAND2_X2 u4_sub_470_U18 ( .A1(u4_exp_in_pl1_6_), .A2(u4_sub_470_n18), .ZN(
        u4_sub_470_n49) );
  INV_X4 u4_sub_470_U17 ( .A(u4_sub_470_n8), .ZN(u4_sub_470_n7) );
  NAND3_X4 u4_sub_470_U16 ( .A1(u4_sub_470_n68), .A2(u4_sub_470_n69), .A3(
        u4_sub_470_n67), .ZN(u4_sub_470_n66) );
  NAND2_X2 u4_sub_470_U15 ( .A1(u4_sub_470_n62), .A2(u4_sub_470_n63), .ZN(
        u4_sub_470_n51) );
  INV_X2 u4_sub_470_U14 ( .A(u4_exp_in_pl1_10_), .ZN(u4_sub_470_n72) );
  INV_X2 u4_sub_470_U13 ( .A(u4_exp_in_pl1_9_), .ZN(u4_sub_470_n4) );
  INV_X2 u4_sub_470_U12 ( .A(u4_exp_in_pl1_8_), .ZN(u4_sub_470_n3) );
  INV_X2 u4_sub_470_U11 ( .A(u4_exp_in_pl1_7_), .ZN(u4_sub_470_n8) );
  NAND3_X2 u4_sub_470_U10 ( .A1(u4_sub_470_n61), .A2(u4_sub_470_n39), .A3(
        u4_sub_470_n90), .ZN(u4_sub_470_n80) );
  OAI21_X1 u4_sub_470_U9 ( .B1(u4_sub_470_n59), .B2(u4_sub_470_n60), .A(
        u4_sub_470_n34), .ZN(u4_sub_470_n53) );
  NOR2_X2 u4_sub_470_U8 ( .A1(u4_sub_470_n51), .A2(u4_sub_470_n52), .ZN(
        u4_sub_470_n47) );
  NOR2_X2 u4_sub_470_U7 ( .A1(u4_sub_470_n56), .A2(u4_sub_470_n86), .ZN(
        u4_sub_470_n83) );
  NOR2_X2 u4_sub_470_U6 ( .A1(u4_sub_470_n56), .A2(u4_sub_470_n86), .ZN(
        u4_sub_470_n90) );
  NOR2_X1 u4_sub_470_U5 ( .A1(u4_sub_470_n56), .A2(u4_sub_470_n30), .ZN(
        u4_sub_470_n55) );
  NOR2_X1 u4_sub_470_U4 ( .A1(u4_sub_470_n64), .A2(u4_sub_470_n15), .ZN(
        u4_sub_470_n63) );
  NOR3_X1 u4_sub_470_U3 ( .A1(u4_sub_470_n57), .A2(u4_sub_470_n58), .A3(
        u4_sub_470_n37), .ZN(u4_sub_470_n54) );
  INV_X4 u4_add_464_U35 ( .A(u4_exp_out_0_), .ZN(u4_exp_out_pl1_0_) );
  NAND2_X2 u4_add_464_U34 ( .A1(net96080), .A2(net87237), .ZN(u4_add_464_n23)
         );
  NOR2_X4 u4_add_464_U33 ( .A1(u4_add_464_n13), .A2(u4_add_464_n23), .ZN(
        u4_add_464_n10) );
  NAND2_X2 u4_add_464_U32 ( .A1(u4_exp_out_6_), .A2(u4_add_464_n10), .ZN(
        u4_add_464_n8) );
  INV_X4 u4_add_464_U31 ( .A(u4_add_464_n8), .ZN(u4_add_464_n2) );
  NAND2_X2 u4_add_464_U30 ( .A1(u4_add_464_n2), .A2(u4_exp_out_7_), .ZN(
        u4_add_464_n22) );
  XNOR2_X2 u4_add_464_U29 ( .A(u4_add_464_n19), .B(u4_add_464_n20), .ZN(
        u4_exp_out_pl1_10_) );
  XNOR2_X2 u4_add_464_U28 ( .A(u4_exp_out_1_), .B(u4_exp_out_0_), .ZN(
        u4_add_464_n18) );
  INV_X4 u4_add_464_U27 ( .A(u4_add_464_n18), .ZN(u4_exp_out_pl1_1_) );
  NAND2_X2 u4_add_464_U26 ( .A1(u4_exp_out_1_), .A2(u4_exp_out_0_), .ZN(
        u4_add_464_n17) );
  XNOR2_X2 u4_add_464_U25 ( .A(u4_exp_out_2_), .B(u4_add_464_n17), .ZN(
        u4_exp_out_pl1_2_) );
  XNOR2_X2 u4_add_464_U24 ( .A(u4_exp_out_3_), .B(u4_add_464_n16), .ZN(
        u4_exp_out_pl1_3_) );
  INV_X4 u4_add_464_U23 ( .A(net96080), .ZN(u4_add_464_n15) );
  XNOR2_X2 u4_add_464_U22 ( .A(u4_add_464_n14), .B(u4_add_464_n15), .ZN(
        u4_exp_out_pl1_4_) );
  INV_X4 u4_add_464_U21 ( .A(u4_add_464_n13), .ZN(u4_add_464_n12) );
  NAND3_X2 u4_add_464_U20 ( .A1(u4_add_464_n12), .A2(net96080), .A3(
        u4_exp_out_0_), .ZN(u4_add_464_n11) );
  XNOR2_X2 u4_add_464_U19 ( .A(net87237), .B(u4_add_464_n11), .ZN(
        u4_exp_out_pl1_5_) );
  NAND2_X2 u4_add_464_U18 ( .A1(u4_add_464_n10), .A2(u4_exp_out_0_), .ZN(
        u4_add_464_n9) );
  XNOR2_X2 u4_add_464_U17 ( .A(u4_exp_out_6_), .B(u4_add_464_n9), .ZN(
        u4_exp_out_pl1_6_) );
  NOR2_X4 u4_add_464_U16 ( .A1(u4_exp_out_pl1_0_), .A2(u4_add_464_n8), .ZN(
        u4_add_464_n7) );
  INV_X4 u4_add_464_U15 ( .A(u4_exp_out_7_), .ZN(u4_add_464_n4) );
  XNOR2_X2 u4_add_464_U14 ( .A(u4_add_464_n7), .B(u4_add_464_n4), .ZN(
        u4_exp_out_pl1_7_) );
  NAND3_X2 u4_add_464_U13 ( .A1(u4_add_464_n2), .A2(u4_exp_out_7_), .A3(
        u4_exp_out_0_), .ZN(u4_add_464_n6) );
  XNOR2_X2 u4_add_464_U12 ( .A(u4_exp_out_8_), .B(u4_add_464_n6), .ZN(
        u4_exp_out_pl1_8_) );
  INV_X4 u4_add_464_U11 ( .A(u4_exp_out_8_), .ZN(u4_add_464_n5) );
  NAND3_X2 u4_add_464_U10 ( .A1(u4_add_464_n2), .A2(u4_add_464_n3), .A3(
        u4_exp_out_0_), .ZN(u4_add_464_n1) );
  INV_X2 u4_add_464_U9 ( .A(u4_exp_out_10_), .ZN(u4_add_464_n20) );
  NAND3_X1 u4_add_464_U8 ( .A1(u4_exp_out_9_), .A2(u4_exp_out_8_), .A3(
        u4_exp_out_0_), .ZN(u4_add_464_n21) );
  XNOR2_X1 u4_add_464_U7 ( .A(u4_exp_out_9_), .B(u4_add_464_n1), .ZN(
        u4_exp_out_pl1_9_) );
  NOR2_X1 u4_add_464_U6 ( .A1(u4_exp_out_pl1_0_), .A2(u4_add_464_n13), .ZN(
        u4_add_464_n14) );
  NAND3_X1 u4_add_464_U5 ( .A1(u4_exp_out_2_), .A2(u4_exp_out_0_), .A3(
        u4_exp_out_1_), .ZN(u4_add_464_n16) );
  NAND3_X1 u4_add_464_U4 ( .A1(u4_exp_out_2_), .A2(u4_exp_out_3_), .A3(
        u4_exp_out_1_), .ZN(u4_add_464_n13) );
  NOR2_X2 u4_add_464_U3 ( .A1(u4_add_464_n4), .A2(u4_add_464_n5), .ZN(
        u4_add_464_n3) );
  NOR2_X2 u4_add_464_U2 ( .A1(u4_add_464_n21), .A2(u4_add_464_n22), .ZN(
        u4_add_464_n19) );
  INV_X4 u4_add_396_U226 ( .A(u4_fract_out_0_), .ZN(u4_fract_out_pl1_0_) );
  NAND4_X2 u4_add_396_U225 ( .A1(u4_fract_out_4_), .A2(u4_fract_out_3_), .A3(
        u4_fract_out_2_), .A4(u4_fract_out_1_), .ZN(u4_add_396_n172) );
  NAND3_X4 u4_add_396_U224 ( .A1(u4_fract_out_6_), .A2(u4_fract_out_7_), .A3(
        u4_fract_out_5_), .ZN(u4_add_396_n173) );
  NOR2_X4 u4_add_396_U223 ( .A1(u4_add_396_n172), .A2(u4_add_396_n173), .ZN(
        u4_add_396_n26) );
  NAND2_X2 u4_add_396_U222 ( .A1(u4_add_396_n26), .A2(u4_fract_out_0_), .ZN(
        u4_add_396_n5) );
  INV_X4 u4_add_396_U221 ( .A(u4_add_396_n5), .ZN(u4_add_396_n153) );
  NAND3_X4 u4_add_396_U220 ( .A1(u4_fract_out_8_), .A2(u4_fract_out_9_), .A3(
        u4_add_396_n153), .ZN(u4_add_396_n171) );
  INV_X4 u4_add_396_U219 ( .A(u4_add_396_n171), .ZN(u4_add_396_n170) );
  INV_X4 u4_add_396_U218 ( .A(u4_fract_out_10_), .ZN(u4_add_396_n31) );
  XNOR2_X2 u4_add_396_U217 ( .A(u4_add_396_n170), .B(u4_add_396_n31), .ZN(
        u4_fract_out_pl1_10_) );
  NAND2_X2 u4_add_396_U216 ( .A1(u4_add_396_n170), .A2(u4_fract_out_10_), .ZN(
        u4_add_396_n169) );
  XNOR2_X2 u4_add_396_U215 ( .A(u4_fract_out_11_), .B(u4_add_396_n169), .ZN(
        u4_fract_out_pl1_11_) );
  NAND4_X2 u4_add_396_U214 ( .A1(u4_fract_out_9_), .A2(u4_fract_out_8_), .A3(
        u4_fract_out_11_), .A4(u4_fract_out_10_), .ZN(u4_add_396_n155) );
  INV_X4 u4_add_396_U213 ( .A(u4_add_396_n155), .ZN(u4_add_396_n168) );
  NAND2_X2 u4_add_396_U212 ( .A1(u4_add_396_n168), .A2(u4_add_396_n153), .ZN(
        u4_add_396_n167) );
  INV_X4 u4_add_396_U211 ( .A(u4_add_396_n167), .ZN(u4_add_396_n163) );
  INV_X4 u4_add_396_U210 ( .A(u4_fract_out_12_), .ZN(u4_add_396_n164) );
  XNOR2_X2 u4_add_396_U209 ( .A(u4_add_396_n163), .B(u4_add_396_n164), .ZN(
        u4_fract_out_pl1_12_) );
  NAND2_X2 u4_add_396_U208 ( .A1(u4_add_396_n163), .A2(u4_fract_out_12_), .ZN(
        u4_add_396_n166) );
  XNOR2_X2 u4_add_396_U207 ( .A(u4_fract_out_13_), .B(u4_add_396_n166), .ZN(
        u4_fract_out_pl1_13_) );
  INV_X4 u4_add_396_U206 ( .A(u4_fract_out_13_), .ZN(u4_add_396_n165) );
  NAND2_X2 u4_add_396_U205 ( .A1(u4_add_396_n162), .A2(u4_add_396_n163), .ZN(
        u4_add_396_n161) );
  XNOR2_X2 u4_add_396_U204 ( .A(u4_fract_out_14_), .B(u4_add_396_n161), .ZN(
        u4_fract_out_pl1_14_) );
  INV_X4 u4_add_396_U203 ( .A(u4_fract_out_14_), .ZN(u4_add_396_n160) );
  INV_X4 u4_add_396_U202 ( .A(u4_fract_out_15_), .ZN(u4_add_396_n159) );
  XNOR2_X2 u4_add_396_U201 ( .A(u4_add_396_n158), .B(u4_add_396_n159), .ZN(
        u4_fract_out_pl1_15_) );
  NAND2_X2 u4_add_396_U200 ( .A1(u4_fract_out_12_), .A2(u4_fract_out_13_), 
        .ZN(u4_add_396_n156) );
  NAND2_X2 u4_add_396_U199 ( .A1(u4_fract_out_15_), .A2(u4_fract_out_14_), 
        .ZN(u4_add_396_n157) );
  NAND2_X2 u4_add_396_U198 ( .A1(u4_add_396_n153), .A2(u4_add_396_n154), .ZN(
        u4_add_396_n152) );
  INV_X4 u4_add_396_U197 ( .A(u4_add_396_n152), .ZN(u4_add_396_n102) );
  INV_X4 u4_add_396_U196 ( .A(u4_fract_out_16_), .ZN(u4_add_396_n149) );
  XNOR2_X2 u4_add_396_U195 ( .A(u4_add_396_n102), .B(u4_add_396_n149), .ZN(
        u4_fract_out_pl1_16_) );
  NAND2_X2 u4_add_396_U194 ( .A1(u4_add_396_n102), .A2(u4_fract_out_16_), .ZN(
        u4_add_396_n151) );
  XNOR2_X2 u4_add_396_U193 ( .A(u4_fract_out_17_), .B(u4_add_396_n151), .ZN(
        u4_fract_out_pl1_17_) );
  INV_X4 u4_add_396_U192 ( .A(u4_fract_out_17_), .ZN(u4_add_396_n150) );
  NOR2_X4 u4_add_396_U191 ( .A1(u4_add_396_n149), .A2(u4_add_396_n150), .ZN(
        u4_add_396_n148) );
  NAND2_X2 u4_add_396_U190 ( .A1(u4_add_396_n148), .A2(u4_add_396_n102), .ZN(
        u4_add_396_n147) );
  INV_X4 u4_add_396_U189 ( .A(u4_add_396_n147), .ZN(u4_add_396_n128) );
  INV_X4 u4_add_396_U188 ( .A(u4_fract_out_18_), .ZN(u4_add_396_n144) );
  XNOR2_X2 u4_add_396_U187 ( .A(u4_add_396_n128), .B(u4_add_396_n144), .ZN(
        u4_fract_out_pl1_18_) );
  NAND2_X2 u4_add_396_U186 ( .A1(u4_add_396_n128), .A2(u4_fract_out_18_), .ZN(
        u4_add_396_n146) );
  XNOR2_X2 u4_add_396_U185 ( .A(u4_fract_out_19_), .B(u4_add_396_n146), .ZN(
        u4_fract_out_pl1_19_) );
  INV_X4 u4_add_396_U184 ( .A(u4_fract_out_19_), .ZN(u4_add_396_n145) );
  NAND2_X2 u4_add_396_U183 ( .A1(u4_add_396_n143), .A2(u4_add_396_n128), .ZN(
        u4_add_396_n142) );
  INV_X4 u4_add_396_U182 ( .A(u4_add_396_n142), .ZN(u4_add_396_n139) );
  INV_X4 u4_add_396_U181 ( .A(u4_fract_out_20_), .ZN(u4_add_396_n131) );
  XNOR2_X2 u4_add_396_U180 ( .A(u4_add_396_n139), .B(u4_add_396_n131), .ZN(
        u4_fract_out_pl1_20_) );
  NAND2_X2 u4_add_396_U179 ( .A1(u4_add_396_n139), .A2(u4_fract_out_20_), .ZN(
        u4_add_396_n141) );
  XNOR2_X2 u4_add_396_U178 ( .A(u4_fract_out_21_), .B(u4_add_396_n141), .ZN(
        u4_fract_out_pl1_21_) );
  INV_X4 u4_add_396_U177 ( .A(u4_fract_out_21_), .ZN(u4_add_396_n140) );
  NAND2_X2 u4_add_396_U176 ( .A1(u4_add_396_n138), .A2(u4_add_396_n139), .ZN(
        u4_add_396_n137) );
  XNOR2_X2 u4_add_396_U175 ( .A(u4_fract_out_22_), .B(u4_add_396_n137), .ZN(
        u4_fract_out_pl1_22_) );
  INV_X4 u4_add_396_U174 ( .A(u4_add_396_n137), .ZN(u4_add_396_n136) );
  NAND2_X2 u4_add_396_U173 ( .A1(u4_add_396_n136), .A2(u4_fract_out_22_), .ZN(
        u4_add_396_n135) );
  XNOR2_X2 u4_add_396_U172 ( .A(u4_fract_out_23_), .B(u4_add_396_n135), .ZN(
        u4_fract_out_pl1_23_) );
  INV_X4 u4_add_396_U171 ( .A(u4_fract_out_23_), .ZN(u4_add_396_n133) );
  NAND2_X2 u4_add_396_U170 ( .A1(u4_fract_out_22_), .A2(u4_fract_out_21_), 
        .ZN(u4_add_396_n134) );
  NAND2_X2 u4_add_396_U169 ( .A1(u4_fract_out_19_), .A2(u4_fract_out_18_), 
        .ZN(u4_add_396_n132) );
  NAND2_X2 u4_add_396_U168 ( .A1(u4_add_396_n128), .A2(u4_add_396_n1), .ZN(
        u4_add_396_n127) );
  XNOR2_X2 u4_add_396_U167 ( .A(u4_fract_out_24_), .B(u4_add_396_n127), .ZN(
        u4_fract_out_pl1_24_) );
  INV_X4 u4_add_396_U166 ( .A(u4_add_396_n127), .ZN(u4_add_396_n117) );
  NAND2_X2 u4_add_396_U165 ( .A1(u4_add_396_n117), .A2(u4_fract_out_24_), .ZN(
        u4_add_396_n126) );
  XNOR2_X2 u4_add_396_U164 ( .A(u4_fract_out_25_), .B(u4_add_396_n126), .ZN(
        u4_fract_out_pl1_25_) );
  INV_X4 u4_add_396_U163 ( .A(u4_fract_out_24_), .ZN(u4_add_396_n124) );
  INV_X4 u4_add_396_U162 ( .A(u4_fract_out_25_), .ZN(u4_add_396_n125) );
  NAND2_X2 u4_add_396_U161 ( .A1(u4_add_396_n123), .A2(u4_add_396_n117), .ZN(
        u4_add_396_n122) );
  INV_X4 u4_add_396_U160 ( .A(u4_add_396_n122), .ZN(u4_add_396_n120) );
  INV_X4 u4_add_396_U159 ( .A(u4_fract_out_26_), .ZN(u4_add_396_n121) );
  XNOR2_X2 u4_add_396_U158 ( .A(u4_add_396_n120), .B(u4_add_396_n121), .ZN(
        u4_fract_out_pl1_26_) );
  NAND2_X2 u4_add_396_U157 ( .A1(u4_add_396_n120), .A2(u4_fract_out_26_), .ZN(
        u4_add_396_n119) );
  XNOR2_X2 u4_add_396_U156 ( .A(u4_fract_out_27_), .B(u4_add_396_n119), .ZN(
        u4_fract_out_pl1_27_) );
  NAND4_X2 u4_add_396_U155 ( .A1(u4_fract_out_27_), .A2(u4_fract_out_26_), 
        .A3(u4_fract_out_25_), .A4(u4_fract_out_24_), .ZN(u4_add_396_n103) );
  INV_X4 u4_add_396_U154 ( .A(u4_add_396_n103), .ZN(u4_add_396_n118) );
  NAND2_X2 u4_add_396_U153 ( .A1(u4_add_396_n117), .A2(u4_add_396_n118), .ZN(
        u4_add_396_n116) );
  XNOR2_X2 u4_add_396_U152 ( .A(u4_fract_out_28_), .B(u4_add_396_n116), .ZN(
        u4_fract_out_pl1_28_) );
  INV_X4 u4_add_396_U151 ( .A(u4_add_396_n116), .ZN(u4_add_396_n112) );
  NAND2_X2 u4_add_396_U150 ( .A1(u4_add_396_n112), .A2(u4_fract_out_28_), .ZN(
        u4_add_396_n115) );
  XNOR2_X2 u4_add_396_U149 ( .A(u4_fract_out_29_), .B(u4_add_396_n115), .ZN(
        u4_fract_out_pl1_29_) );
  NAND2_X2 u4_add_396_U148 ( .A1(u4_fract_out_1_), .A2(u4_fract_out_0_), .ZN(
        u4_add_396_n81) );
  XNOR2_X2 u4_add_396_U147 ( .A(u4_fract_out_2_), .B(u4_add_396_n81), .ZN(
        u4_fract_out_pl1_2_) );
  INV_X4 u4_add_396_U146 ( .A(u4_fract_out_28_), .ZN(u4_add_396_n113) );
  INV_X4 u4_add_396_U145 ( .A(u4_fract_out_29_), .ZN(u4_add_396_n114) );
  NAND2_X2 u4_add_396_U144 ( .A1(u4_add_396_n111), .A2(u4_add_396_n112), .ZN(
        u4_add_396_n110) );
  INV_X4 u4_add_396_U143 ( .A(u4_add_396_n110), .ZN(u4_add_396_n108) );
  INV_X4 u4_add_396_U142 ( .A(u4_fract_out_30_), .ZN(u4_add_396_n109) );
  XNOR2_X2 u4_add_396_U141 ( .A(u4_add_396_n108), .B(u4_add_396_n109), .ZN(
        u4_fract_out_pl1_30_) );
  NAND2_X2 u4_add_396_U140 ( .A1(u4_add_396_n108), .A2(u4_fract_out_30_), .ZN(
        u4_add_396_n107) );
  XNOR2_X2 u4_add_396_U139 ( .A(u4_fract_out_31_), .B(u4_add_396_n107), .ZN(
        u4_fract_out_pl1_31_) );
  NAND2_X2 u4_add_396_U138 ( .A1(u4_fract_out_17_), .A2(u4_fract_out_16_), 
        .ZN(u4_add_396_n106) );
  INV_X4 u4_add_396_U137 ( .A(u4_fract_out_31_), .ZN(u4_add_396_n104) );
  NOR2_X4 u4_add_396_U136 ( .A1(u4_add_396_n103), .A2(u4_add_396_n104), .ZN(
        u4_add_396_n101) );
  NAND4_X2 u4_add_396_U135 ( .A1(u4_add_396_n1), .A2(u4_add_396_n100), .A3(
        u4_add_396_n101), .A4(u4_add_396_n102), .ZN(u4_add_396_n89) );
  INV_X4 u4_add_396_U134 ( .A(u4_add_396_n89), .ZN(u4_add_396_n96) );
  INV_X4 u4_add_396_U133 ( .A(u4_fract_out_32_), .ZN(u4_add_396_n97) );
  XNOR2_X2 u4_add_396_U132 ( .A(u4_add_396_n96), .B(u4_add_396_n97), .ZN(
        u4_fract_out_pl1_32_) );
  NAND2_X2 u4_add_396_U131 ( .A1(u4_add_396_n96), .A2(u4_fract_out_32_), .ZN(
        u4_add_396_n99) );
  XNOR2_X2 u4_add_396_U130 ( .A(u4_fract_out_33_), .B(u4_add_396_n99), .ZN(
        u4_fract_out_pl1_33_) );
  INV_X4 u4_add_396_U129 ( .A(u4_fract_out_33_), .ZN(u4_add_396_n98) );
  NOR2_X4 u4_add_396_U128 ( .A1(u4_add_396_n97), .A2(u4_add_396_n98), .ZN(
        u4_add_396_n95) );
  NAND2_X2 u4_add_396_U127 ( .A1(u4_add_396_n95), .A2(u4_add_396_n96), .ZN(
        u4_add_396_n94) );
  INV_X4 u4_add_396_U126 ( .A(u4_add_396_n94), .ZN(u4_add_396_n92) );
  INV_X4 u4_add_396_U125 ( .A(u4_fract_out_34_), .ZN(u4_add_396_n93) );
  XNOR2_X2 u4_add_396_U124 ( .A(u4_add_396_n92), .B(u4_add_396_n93), .ZN(
        u4_fract_out_pl1_34_) );
  NAND2_X2 u4_add_396_U123 ( .A1(u4_add_396_n92), .A2(u4_fract_out_34_), .ZN(
        u4_add_396_n91) );
  XNOR2_X2 u4_add_396_U122 ( .A(u4_fract_out_35_), .B(u4_add_396_n91), .ZN(
        u4_fract_out_pl1_35_) );
  NAND4_X2 u4_add_396_U121 ( .A1(u4_fract_out_35_), .A2(u4_fract_out_32_), 
        .A3(u4_fract_out_33_), .A4(u4_fract_out_34_), .ZN(u4_add_396_n90) );
  NOR2_X4 u4_add_396_U120 ( .A1(u4_add_396_n89), .A2(u4_add_396_n90), .ZN(
        u4_add_396_n75) );
  INV_X4 u4_add_396_U119 ( .A(u4_fract_out_36_), .ZN(u4_add_396_n86) );
  XNOR2_X2 u4_add_396_U118 ( .A(u4_add_396_n75), .B(u4_add_396_n86), .ZN(
        u4_fract_out_pl1_36_) );
  NAND2_X2 u4_add_396_U117 ( .A1(u4_add_396_n75), .A2(u4_fract_out_36_), .ZN(
        u4_add_396_n88) );
  XNOR2_X2 u4_add_396_U116 ( .A(u4_fract_out_37_), .B(u4_add_396_n88), .ZN(
        u4_fract_out_pl1_37_) );
  INV_X4 u4_add_396_U115 ( .A(u4_fract_out_37_), .ZN(u4_add_396_n87) );
  NOR2_X4 u4_add_396_U114 ( .A1(u4_add_396_n86), .A2(u4_add_396_n87), .ZN(
        u4_add_396_n85) );
  NAND2_X2 u4_add_396_U113 ( .A1(u4_add_396_n85), .A2(u4_add_396_n75), .ZN(
        u4_add_396_n84) );
  XNOR2_X2 u4_add_396_U112 ( .A(u4_fract_out_38_), .B(u4_add_396_n84), .ZN(
        u4_fract_out_pl1_38_) );
  INV_X4 u4_add_396_U111 ( .A(u4_add_396_n84), .ZN(u4_add_396_n83) );
  NAND2_X2 u4_add_396_U110 ( .A1(u4_add_396_n83), .A2(u4_fract_out_38_), .ZN(
        u4_add_396_n82) );
  XNOR2_X2 u4_add_396_U109 ( .A(u4_fract_out_39_), .B(u4_add_396_n82), .ZN(
        u4_fract_out_pl1_39_) );
  INV_X4 u4_add_396_U108 ( .A(u4_fract_out_2_), .ZN(u4_add_396_n80) );
  INV_X4 u4_add_396_U107 ( .A(u4_fract_out_3_), .ZN(u4_add_396_n79) );
  XNOR2_X2 u4_add_396_U106 ( .A(u4_add_396_n78), .B(u4_add_396_n79), .ZN(
        u4_fract_out_pl1_3_) );
  NAND2_X2 u4_add_396_U105 ( .A1(u4_fract_out_37_), .A2(u4_fract_out_38_), 
        .ZN(u4_add_396_n76) );
  NAND2_X2 u4_add_396_U104 ( .A1(u4_fract_out_39_), .A2(u4_fract_out_36_), 
        .ZN(u4_add_396_n77) );
  NAND2_X2 u4_add_396_U103 ( .A1(u4_add_396_n74), .A2(u4_add_396_n75), .ZN(
        u4_add_396_n51) );
  XNOR2_X2 u4_add_396_U102 ( .A(u4_fract_out_40_), .B(u4_add_396_n51), .ZN(
        u4_fract_out_pl1_40_) );
  INV_X4 u4_add_396_U101 ( .A(u4_add_396_n51), .ZN(u4_add_396_n64) );
  NAND2_X2 u4_add_396_U100 ( .A1(u4_add_396_n64), .A2(u4_fract_out_40_), .ZN(
        u4_add_396_n73) );
  XNOR2_X2 u4_add_396_U99 ( .A(u4_fract_out_41_), .B(u4_add_396_n73), .ZN(
        u4_fract_out_pl1_41_) );
  INV_X4 u4_add_396_U98 ( .A(u4_fract_out_40_), .ZN(u4_add_396_n71) );
  INV_X4 u4_add_396_U97 ( .A(u4_fract_out_41_), .ZN(u4_add_396_n72) );
  NAND2_X2 u4_add_396_U96 ( .A1(u4_add_396_n70), .A2(u4_add_396_n64), .ZN(
        u4_add_396_n69) );
  INV_X4 u4_add_396_U95 ( .A(u4_add_396_n69), .ZN(u4_add_396_n67) );
  INV_X4 u4_add_396_U94 ( .A(u4_fract_out_42_), .ZN(u4_add_396_n68) );
  XNOR2_X2 u4_add_396_U93 ( .A(u4_add_396_n67), .B(u4_add_396_n68), .ZN(
        u4_fract_out_pl1_42_) );
  NAND2_X2 u4_add_396_U92 ( .A1(u4_add_396_n67), .A2(u4_fract_out_42_), .ZN(
        u4_add_396_n66) );
  XNOR2_X2 u4_add_396_U91 ( .A(u4_fract_out_43_), .B(u4_add_396_n66), .ZN(
        u4_fract_out_pl1_43_) );
  NAND4_X2 u4_add_396_U90 ( .A1(u4_fract_out_43_), .A2(u4_fract_out_42_), .A3(
        u4_fract_out_41_), .A4(u4_fract_out_40_), .ZN(u4_add_396_n52) );
  INV_X4 u4_add_396_U89 ( .A(u4_add_396_n52), .ZN(u4_add_396_n65) );
  NAND2_X2 u4_add_396_U88 ( .A1(u4_add_396_n64), .A2(u4_add_396_n65), .ZN(
        u4_add_396_n63) );
  XNOR2_X2 u4_add_396_U87 ( .A(u4_fract_out_44_), .B(u4_add_396_n63), .ZN(
        u4_fract_out_pl1_44_) );
  INV_X4 u4_add_396_U86 ( .A(u4_add_396_n63), .ZN(u4_add_396_n59) );
  NAND2_X2 u4_add_396_U85 ( .A1(u4_add_396_n59), .A2(u4_fract_out_44_), .ZN(
        u4_add_396_n62) );
  XNOR2_X2 u4_add_396_U84 ( .A(u4_fract_out_45_), .B(u4_add_396_n62), .ZN(
        u4_fract_out_pl1_45_) );
  INV_X4 u4_add_396_U83 ( .A(u4_fract_out_44_), .ZN(u4_add_396_n60) );
  INV_X4 u4_add_396_U82 ( .A(u4_fract_out_45_), .ZN(u4_add_396_n61) );
  NAND2_X2 u4_add_396_U81 ( .A1(u4_add_396_n58), .A2(u4_add_396_n59), .ZN(
        u4_add_396_n57) );
  INV_X4 u4_add_396_U80 ( .A(u4_add_396_n57), .ZN(u4_add_396_n55) );
  INV_X4 u4_add_396_U79 ( .A(u4_fract_out_46_), .ZN(u4_add_396_n56) );
  XNOR2_X2 u4_add_396_U78 ( .A(u4_add_396_n55), .B(u4_add_396_n56), .ZN(
        u4_fract_out_pl1_46_) );
  NAND2_X2 u4_add_396_U77 ( .A1(u4_add_396_n55), .A2(u4_fract_out_46_), .ZN(
        u4_add_396_n54) );
  XNOR2_X2 u4_add_396_U76 ( .A(u4_fract_out_47_), .B(u4_add_396_n54), .ZN(
        u4_fract_out_pl1_47_) );
  NAND4_X2 u4_add_396_U75 ( .A1(u4_fract_out_47_), .A2(u4_fract_out_44_), .A3(
        u4_fract_out_45_), .A4(u4_fract_out_46_), .ZN(u4_add_396_n53) );
  NOR3_X4 u4_add_396_U74 ( .A1(u4_add_396_n51), .A2(u4_add_396_n52), .A3(
        u4_add_396_n53), .ZN(u4_add_396_n48) );
  INV_X4 u4_add_396_U73 ( .A(u4_fract_out_48_), .ZN(u4_add_396_n50) );
  XNOR2_X2 u4_add_396_U72 ( .A(u4_add_396_n48), .B(u4_add_396_n50), .ZN(
        u4_fract_out_pl1_48_) );
  NAND2_X2 u4_add_396_U71 ( .A1(u4_add_396_n48), .A2(u4_fract_out_48_), .ZN(
        u4_add_396_n49) );
  XNOR2_X2 u4_add_396_U70 ( .A(u4_fract_out_49_), .B(u4_add_396_n49), .ZN(
        u4_fract_out_pl1_49_) );
  NAND4_X2 u4_add_396_U69 ( .A1(u4_fract_out_3_), .A2(u4_fract_out_2_), .A3(
        u4_fract_out_1_), .A4(u4_fract_out_0_), .ZN(u4_add_396_n15) );
  INV_X4 u4_add_396_U68 ( .A(u4_add_396_n15), .ZN(u4_add_396_n11) );
  INV_X4 u4_add_396_U67 ( .A(u4_fract_out_4_), .ZN(u4_add_396_n14) );
  XNOR2_X2 u4_add_396_U66 ( .A(u4_add_396_n11), .B(u4_add_396_n14), .ZN(
        u4_fract_out_pl1_4_) );
  NAND3_X4 u4_add_396_U65 ( .A1(u4_fract_out_49_), .A2(u4_fract_out_48_), .A3(
        u4_add_396_n48), .ZN(u4_add_396_n47) );
  XNOR2_X2 u4_add_396_U64 ( .A(u4_fract_out_50_), .B(u4_add_396_n47), .ZN(
        u4_fract_out_pl1_50_) );
  INV_X4 u4_add_396_U63 ( .A(u4_add_396_n47), .ZN(u4_add_396_n46) );
  NAND2_X2 u4_add_396_U62 ( .A1(u4_add_396_n46), .A2(u4_fract_out_50_), .ZN(
        u4_add_396_n45) );
  XNOR2_X2 u4_add_396_U61 ( .A(u4_fract_out_51_), .B(u4_add_396_n45), .ZN(
        u4_fract_out_pl1_51_) );
  NAND3_X4 u4_add_396_U60 ( .A1(u4_fract_out_49_), .A2(u4_fract_out_47_), .A3(
        u4_fract_out_48_), .ZN(u4_add_396_n43) );
  NAND2_X2 u4_add_396_U59 ( .A1(u4_fract_out_51_), .A2(u4_fract_out_50_), .ZN(
        u4_add_396_n44) );
  NAND3_X4 u4_add_396_U58 ( .A1(u4_fract_out_43_), .A2(u4_fract_out_41_), .A3(
        u4_fract_out_42_), .ZN(u4_add_396_n41) );
  NAND3_X4 u4_add_396_U57 ( .A1(u4_fract_out_45_), .A2(u4_fract_out_46_), .A3(
        u4_fract_out_44_), .ZN(u4_add_396_n42) );
  NOR2_X4 u4_add_396_U56 ( .A1(u4_add_396_n41), .A2(u4_add_396_n42), .ZN(
        u4_add_396_n34) );
  NAND3_X4 u4_add_396_U55 ( .A1(u4_fract_out_37_), .A2(u4_fract_out_35_), .A3(
        u4_fract_out_36_), .ZN(u4_add_396_n39) );
  NAND3_X4 u4_add_396_U54 ( .A1(u4_fract_out_39_), .A2(u4_fract_out_38_), .A3(
        u4_fract_out_40_), .ZN(u4_add_396_n40) );
  NOR2_X4 u4_add_396_U53 ( .A1(u4_add_396_n39), .A2(u4_add_396_n40), .ZN(
        u4_add_396_n35) );
  NAND3_X4 u4_add_396_U52 ( .A1(u4_fract_out_33_), .A2(u4_fract_out_34_), .A3(
        u4_fract_out_32_), .ZN(u4_add_396_n38) );
  NOR2_X4 u4_add_396_U51 ( .A1(u4_add_396_n37), .A2(u4_add_396_n38), .ZN(
        u4_add_396_n36) );
  NAND4_X2 u4_add_396_U50 ( .A1(u4_add_396_n33), .A2(u4_add_396_n34), .A3(
        u4_add_396_n35), .A4(u4_add_396_n36), .ZN(u4_add_396_n16) );
  INV_X4 u4_add_396_U49 ( .A(u4_fract_out_8_), .ZN(u4_add_396_n6) );
  NAND2_X2 u4_add_396_U48 ( .A1(u4_fract_out_11_), .A2(u4_fract_out_9_), .ZN(
        u4_add_396_n32) );
  NAND3_X4 u4_add_396_U47 ( .A1(u4_fract_out_17_), .A2(u4_fract_out_15_), .A3(
        u4_fract_out_16_), .ZN(u4_add_396_n30) );
  NOR2_X4 u4_add_396_U46 ( .A1(u4_add_396_n29), .A2(u4_add_396_n30), .ZN(
        u4_add_396_n28) );
  NAND4_X2 u4_add_396_U45 ( .A1(u4_add_396_n25), .A2(u4_add_396_n26), .A3(
        u4_add_396_n27), .A4(u4_add_396_n28), .ZN(u4_add_396_n17) );
  NAND3_X4 u4_add_396_U44 ( .A1(u4_fract_out_25_), .A2(u4_fract_out_26_), .A3(
        u4_fract_out_24_), .ZN(u4_add_396_n23) );
  NAND2_X2 u4_add_396_U43 ( .A1(u4_fract_out_28_), .A2(u4_fract_out_27_), .ZN(
        u4_add_396_n24) );
  NOR2_X4 u4_add_396_U42 ( .A1(u4_add_396_n23), .A2(u4_add_396_n24), .ZN(
        u4_add_396_n19) );
  NAND3_X4 u4_add_396_U41 ( .A1(u4_fract_out_19_), .A2(u4_fract_out_18_), .A3(
        u4_fract_out_20_), .ZN(u4_add_396_n21) );
  NAND3_X4 u4_add_396_U40 ( .A1(u4_fract_out_22_), .A2(u4_fract_out_21_), .A3(
        u4_fract_out_23_), .ZN(u4_add_396_n22) );
  NOR2_X4 u4_add_396_U39 ( .A1(u4_add_396_n21), .A2(u4_add_396_n22), .ZN(
        u4_add_396_n20) );
  NAND2_X2 u4_add_396_U38 ( .A1(u4_add_396_n19), .A2(u4_add_396_n20), .ZN(
        u4_add_396_n18) );
  NOR3_X4 u4_add_396_U37 ( .A1(u4_add_396_n16), .A2(u4_add_396_n17), .A3(
        u4_add_396_n18), .ZN(u4_fract_out_pl1_52_) );
  INV_X4 u4_add_396_U36 ( .A(u4_fract_out_5_), .ZN(u4_add_396_n13) );
  XNOR2_X2 u4_add_396_U35 ( .A(u4_add_396_n12), .B(u4_add_396_n13), .ZN(
        u4_fract_out_pl1_5_) );
  NAND3_X4 u4_add_396_U34 ( .A1(u4_fract_out_5_), .A2(u4_fract_out_4_), .A3(
        u4_add_396_n11), .ZN(u4_add_396_n10) );
  INV_X4 u4_add_396_U33 ( .A(u4_add_396_n10), .ZN(u4_add_396_n8) );
  INV_X4 u4_add_396_U32 ( .A(u4_fract_out_6_), .ZN(u4_add_396_n9) );
  XNOR2_X2 u4_add_396_U31 ( .A(u4_add_396_n8), .B(u4_add_396_n9), .ZN(
        u4_fract_out_pl1_6_) );
  NAND2_X2 u4_add_396_U30 ( .A1(u4_add_396_n8), .A2(u4_fract_out_6_), .ZN(
        u4_add_396_n7) );
  XNOR2_X2 u4_add_396_U29 ( .A(u4_fract_out_7_), .B(u4_add_396_n7), .ZN(
        u4_fract_out_pl1_7_) );
  XNOR2_X2 u4_add_396_U28 ( .A(u4_fract_out_8_), .B(u4_add_396_n5), .ZN(
        u4_fract_out_pl1_8_) );
  INV_X4 u4_add_396_U27 ( .A(u4_fract_out_9_), .ZN(u4_add_396_n4) );
  XNOR2_X2 u4_add_396_U26 ( .A(u4_add_396_n3), .B(u4_add_396_n4), .ZN(
        u4_fract_out_pl1_9_) );
  XOR2_X1 u4_add_396_U25 ( .A(u4_fract_out_1_), .B(u4_fract_out_0_), .Z(
        u4_fract_out_pl1_1_) );
  AND2_X2 u4_add_396_U24 ( .A1(u4_add_396_n129), .A2(u4_add_396_n130), .ZN(
        u4_add_396_n1) );
  NOR2_X1 u4_add_396_U23 ( .A1(u4_add_396_n5), .A2(u4_add_396_n6), .ZN(
        u4_add_396_n3) );
  NOR2_X1 u4_add_396_U22 ( .A1(u4_add_396_n14), .A2(u4_add_396_n15), .ZN(
        u4_add_396_n12) );
  NOR2_X2 u4_add_396_U21 ( .A1(u4_add_396_n60), .A2(u4_add_396_n61), .ZN(
        u4_add_396_n58) );
  NOR2_X2 u4_add_396_U20 ( .A1(u4_add_396_n71), .A2(u4_add_396_n72), .ZN(
        u4_add_396_n70) );
  NOR2_X2 u4_add_396_U19 ( .A1(u4_add_396_n113), .A2(u4_add_396_n114), .ZN(
        u4_add_396_n111) );
  NOR2_X1 u4_add_396_U18 ( .A1(u4_add_396_n131), .A2(u4_add_396_n140), .ZN(
        u4_add_396_n138) );
  NOR3_X2 u4_add_396_U17 ( .A1(u4_add_396_n155), .A2(u4_add_396_n156), .A3(
        u4_add_396_n157), .ZN(u4_add_396_n154) );
  NOR2_X2 u4_add_396_U16 ( .A1(u4_add_396_n160), .A2(u4_add_396_n161), .ZN(
        u4_add_396_n158) );
  NOR2_X2 u4_add_396_U15 ( .A1(u4_add_396_n80), .A2(u4_add_396_n81), .ZN(
        u4_add_396_n78) );
  NOR2_X2 u4_add_396_U14 ( .A1(u4_add_396_n133), .A2(u4_add_396_n134), .ZN(
        u4_add_396_n129) );
  NOR2_X2 u4_add_396_U13 ( .A1(u4_add_396_n131), .A2(u4_add_396_n132), .ZN(
        u4_add_396_n130) );
  NAND3_X1 u4_add_396_U12 ( .A1(u4_fract_out_30_), .A2(u4_fract_out_29_), .A3(
        u4_fract_out_31_), .ZN(u4_add_396_n37) );
  NOR2_X2 u4_add_396_U11 ( .A1(u4_fract_out_pl1_0_), .A2(u4_add_396_n6), .ZN(
        u4_add_396_n25) );
  NOR2_X2 u4_add_396_U10 ( .A1(u4_add_396_n31), .A2(u4_add_396_n32), .ZN(
        u4_add_396_n27) );
  NAND3_X1 u4_add_396_U9 ( .A1(u4_fract_out_13_), .A2(u4_fract_out_14_), .A3(
        u4_fract_out_12_), .ZN(u4_add_396_n29) );
  NOR2_X2 u4_add_396_U8 ( .A1(u4_add_396_n76), .A2(u4_add_396_n77), .ZN(
        u4_add_396_n74) );
  NOR2_X2 u4_add_396_U7 ( .A1(u4_add_396_n124), .A2(u4_add_396_n125), .ZN(
        u4_add_396_n123) );
  NOR2_X2 u4_add_396_U6 ( .A1(u4_add_396_n164), .A2(u4_add_396_n165), .ZN(
        u4_add_396_n162) );
  NOR2_X2 u4_add_396_U5 ( .A1(u4_add_396_n43), .A2(u4_add_396_n44), .ZN(
        u4_add_396_n33) );
  NOR2_X2 u4_add_396_U4 ( .A1(u4_add_396_n144), .A2(u4_add_396_n145), .ZN(
        u4_add_396_n143) );
  NAND3_X1 u4_add_396_U3 ( .A1(u4_fract_out_29_), .A2(u4_fract_out_28_), .A3(
        u4_fract_out_30_), .ZN(u4_add_396_n105) );
  NOR2_X2 u4_add_396_U2 ( .A1(u4_add_396_n105), .A2(u4_add_396_n106), .ZN(
        u4_add_396_n100) );
  INV_X4 u1_gt_239_U860 ( .A(n8401), .ZN(u1_gt_239_n859) );
  NAND2_X2 u1_gt_239_U859 ( .A1(n8456), .A2(u1_gt_239_n859), .ZN(
        u1_gt_239_n235) );
  INV_X4 u1_gt_239_U858 ( .A(n8402), .ZN(u1_gt_239_n858) );
  NAND2_X2 u1_gt_239_U857 ( .A1(n8457), .A2(u1_gt_239_n858), .ZN(
        u1_gt_239_n766) );
  INV_X4 u1_gt_239_U856 ( .A(n8459), .ZN(u1_gt_239_n857) );
  NOR2_X4 u1_gt_239_U855 ( .A1(n8404), .A2(u1_gt_239_n857), .ZN(u1_gt_239_n854) );
  INV_X4 u1_gt_239_U854 ( .A(n8458), .ZN(u1_gt_239_n856) );
  NOR2_X4 u1_gt_239_U853 ( .A1(n8403), .A2(u1_gt_239_n856), .ZN(u1_gt_239_n855) );
  NOR2_X4 u1_gt_239_U852 ( .A1(u1_gt_239_n854), .A2(u1_gt_239_n855), .ZN(
        u1_gt_239_n853) );
  NAND3_X4 u1_gt_239_U851 ( .A1(u1_gt_239_n235), .A2(u1_gt_239_n766), .A3(
        u1_gt_239_n853), .ZN(u1_gt_239_n113) );
  INV_X4 u1_gt_239_U850 ( .A(n8372), .ZN(u1_gt_239_n504) );
  INV_X4 u1_gt_239_U849 ( .A(n8370), .ZN(u1_gt_239_n852) );
  NAND2_X2 u1_gt_239_U848 ( .A1(n8423), .A2(u1_gt_239_n852), .ZN(
        u1_gt_239_n245) );
  INV_X4 u1_gt_239_U847 ( .A(u1_gt_239_n245), .ZN(u1_gt_239_n89) );
  NOR2_X4 u1_gt_239_U846 ( .A1(u1_gt_239_n86), .A2(u1_gt_239_n31), .ZN(
        u1_gt_239_n849) );
  INV_X4 u1_gt_239_U845 ( .A(n8371), .ZN(u1_gt_239_n851) );
  INV_X4 u1_gt_239_U844 ( .A(n8378), .ZN(u1_gt_239_n727) );
  NAND2_X2 u1_gt_239_U843 ( .A1(n8431), .A2(u1_gt_239_n727), .ZN(
        u1_gt_239_n850) );
  NAND3_X2 u1_gt_239_U842 ( .A1(u1_gt_239_n849), .A2(u1_gt_239_n144), .A3(
        u1_gt_239_n850), .ZN(u1_gt_239_n848) );
  NOR2_X4 u1_gt_239_U841 ( .A1(u1_gt_239_n113), .A2(u1_gt_239_n848), .ZN(
        u1_gt_239_n829) );
  INV_X4 u1_gt_239_U840 ( .A(n8426), .ZN(u1_gt_239_n847) );
  NAND2_X2 u1_gt_239_U839 ( .A1(n8373), .A2(u1_gt_239_n847), .ZN(
        u1_gt_239_n309) );
  INV_X4 u1_gt_239_U838 ( .A(n8374), .ZN(u1_gt_239_n846) );
  INV_X4 u1_gt_239_U837 ( .A(n8373), .ZN(u1_gt_239_n845) );
  NAND2_X2 u1_gt_239_U836 ( .A1(u1_gt_239_n222), .A2(u1_gt_239_n201), .ZN(
        u1_gt_239_n840) );
  INV_X4 u1_gt_239_U835 ( .A(n8428), .ZN(u1_gt_239_n312) );
  NOR2_X4 u1_gt_239_U834 ( .A1(n8375), .A2(u1_gt_239_n312), .ZN(u1_gt_239_n843) );
  INV_X4 u1_gt_239_U833 ( .A(n8427), .ZN(u1_gt_239_n844) );
  NAND2_X2 u1_gt_239_U832 ( .A1(n8374), .A2(u1_gt_239_n844), .ZN(
        u1_gt_239_n311) );
  INV_X4 u1_gt_239_U831 ( .A(n8377), .ZN(u1_gt_239_n91) );
  INV_X4 u1_gt_239_U830 ( .A(n8376), .ZN(u1_gt_239_n533) );
  INV_X4 u1_gt_239_U829 ( .A(n8379), .ZN(u1_gt_239_n842) );
  NAND3_X2 u1_gt_239_U828 ( .A1(u1_gt_239_n78), .A2(u1_gt_239_n77), .A3(
        u1_gt_239_n79), .ZN(u1_gt_239_n841) );
  INV_X4 u1_gt_239_U827 ( .A(n8385), .ZN(u1_gt_239_n397) );
  INV_X4 u1_gt_239_U826 ( .A(n8387), .ZN(u1_gt_239_n146) );
  NAND2_X2 u1_gt_239_U825 ( .A1(n8440), .A2(u1_gt_239_n146), .ZN(
        u1_gt_239_n120) );
  INV_X4 u1_gt_239_U824 ( .A(n8386), .ZN(u1_gt_239_n517) );
  NAND2_X2 u1_gt_239_U823 ( .A1(n8439), .A2(u1_gt_239_n517), .ZN(
        u1_gt_239_n165) );
  INV_X4 u1_gt_239_U822 ( .A(n8388), .ZN(u1_gt_239_n377) );
  NAND2_X2 u1_gt_239_U821 ( .A1(n8441), .A2(u1_gt_239_n377), .ZN(
        u1_gt_239_n121) );
  INV_X4 u1_gt_239_U820 ( .A(n8390), .ZN(u1_gt_239_n362) );
  NAND2_X2 u1_gt_239_U819 ( .A1(n8444), .A2(u1_gt_239_n362), .ZN(
        u1_gt_239_n194) );
  INV_X4 u1_gt_239_U818 ( .A(u1_gt_239_n194), .ZN(u1_gt_239_n162) );
  INV_X4 u1_gt_239_U817 ( .A(n8389), .ZN(u1_gt_239_n438) );
  NAND2_X2 u1_gt_239_U816 ( .A1(n8443), .A2(u1_gt_239_n438), .ZN(
        u1_gt_239_n192) );
  NAND2_X2 u1_gt_239_U815 ( .A1(u1_gt_239_n838), .A2(u1_gt_239_n839), .ZN(
        u1_gt_239_n832) );
  INV_X4 u1_gt_239_U814 ( .A(n8382), .ZN(u1_gt_239_n837) );
  INV_X4 u1_gt_239_U813 ( .A(n8384), .ZN(u1_gt_239_n836) );
  NAND2_X2 u1_gt_239_U812 ( .A1(n8437), .A2(u1_gt_239_n836), .ZN(
        u1_gt_239_n197) );
  INV_X4 u1_gt_239_U811 ( .A(n8383), .ZN(u1_gt_239_n499) );
  NAND3_X2 u1_gt_239_U810 ( .A1(u1_gt_239_n18), .A2(u1_gt_239_n197), .A3(
        u1_gt_239_n17), .ZN(u1_gt_239_n833) );
  INV_X4 u1_gt_239_U809 ( .A(n8380), .ZN(u1_gt_239_n290) );
  INV_X4 u1_gt_239_U808 ( .A(n8381), .ZN(u1_gt_239_n835) );
  NAND2_X2 u1_gt_239_U807 ( .A1(u1_gt_239_n15), .A2(u1_gt_239_n13), .ZN(
        u1_gt_239_n834) );
  NOR3_X4 u1_gt_239_U806 ( .A1(u1_gt_239_n832), .A2(u1_gt_239_n833), .A3(
        u1_gt_239_n834), .ZN(u1_gt_239_n831) );
  NAND3_X2 u1_gt_239_U805 ( .A1(u1_gt_239_n829), .A2(u1_gt_239_n830), .A3(
        u1_gt_239_n831), .ZN(u1_gt_239_n794) );
  INV_X4 u1_gt_239_U804 ( .A(n8394), .ZN(u1_gt_239_n350) );
  INV_X4 u1_gt_239_U803 ( .A(n8395), .ZN(u1_gt_239_n637) );
  NAND2_X2 u1_gt_239_U802 ( .A1(n8449), .A2(u1_gt_239_n637), .ZN(
        u1_gt_239_n566) );
  INV_X4 u1_gt_239_U801 ( .A(n8393), .ZN(u1_gt_239_n155) );
  NAND3_X2 u1_gt_239_U800 ( .A1(u1_gt_239_n213), .A2(u1_gt_239_n566), .A3(
        u1_gt_239_n212), .ZN(u1_gt_239_n828) );
  INV_X4 u1_gt_239_U799 ( .A(n8392), .ZN(u1_gt_239_n411) );
  NAND2_X2 u1_gt_239_U798 ( .A1(n8446), .A2(u1_gt_239_n411), .ZN(
        u1_gt_239_n342) );
  INV_X4 u1_gt_239_U797 ( .A(u1_gt_239_n342), .ZN(u1_gt_239_n160) );
  INV_X4 u1_gt_239_U796 ( .A(n8391), .ZN(u1_gt_239_n203) );
  INV_X4 u1_gt_239_U795 ( .A(n8400), .ZN(u1_gt_239_n827) );
  INV_X4 u1_gt_239_U794 ( .A(n8405), .ZN(u1_gt_239_n543) );
  NAND2_X2 u1_gt_239_U793 ( .A1(n8460), .A2(u1_gt_239_n543), .ZN(
        u1_gt_239_n276) );
  INV_X4 u1_gt_239_U792 ( .A(n8399), .ZN(u1_gt_239_n218) );
  NAND3_X2 u1_gt_239_U791 ( .A1(u1_gt_239_n232), .A2(u1_gt_239_n276), .A3(
        u1_gt_239_n9), .ZN(u1_gt_239_n823) );
  INV_X4 u1_gt_239_U790 ( .A(n8397), .ZN(u1_gt_239_n826) );
  NAND2_X2 u1_gt_239_U789 ( .A1(n8451), .A2(u1_gt_239_n826), .ZN(
        u1_gt_239_n567) );
  INV_X4 u1_gt_239_U788 ( .A(n8398), .ZN(u1_gt_239_n825) );
  NAND2_X2 u1_gt_239_U787 ( .A1(n8452), .A2(u1_gt_239_n825), .ZN(
        u1_gt_239_n568) );
  INV_X4 u1_gt_239_U786 ( .A(n8396), .ZN(u1_gt_239_n461) );
  NAND2_X2 u1_gt_239_U785 ( .A1(n8450), .A2(u1_gt_239_n461), .ZN(
        u1_gt_239_n569) );
  NAND3_X2 u1_gt_239_U784 ( .A1(u1_gt_239_n567), .A2(u1_gt_239_n568), .A3(
        u1_gt_239_n569), .ZN(u1_gt_239_n824) );
  NOR2_X4 u1_gt_239_U783 ( .A1(u1_gt_239_n823), .A2(u1_gt_239_n824), .ZN(
        u1_gt_239_n818) );
  INV_X4 u1_gt_239_U782 ( .A(n8356), .ZN(u1_gt_239_n699) );
  NAND2_X2 u1_gt_239_U781 ( .A1(n8409), .A2(u1_gt_239_n699), .ZN(
        u1_gt_239_n707) );
  INV_X4 u1_gt_239_U780 ( .A(n8357), .ZN(u1_gt_239_n177) );
  NAND2_X2 u1_gt_239_U779 ( .A1(n8410), .A2(u1_gt_239_n177), .ZN(
        u1_gt_239_n560) );
  INV_X4 u1_gt_239_U778 ( .A(n8408), .ZN(u1_gt_239_n822) );
  NAND2_X2 u1_gt_239_U777 ( .A1(n8463), .A2(u1_gt_239_n822), .ZN(
        u1_gt_239_n659) );
  NAND3_X2 u1_gt_239_U776 ( .A1(u1_gt_239_n707), .A2(u1_gt_239_n560), .A3(
        u1_gt_239_n659), .ZN(u1_gt_239_n820) );
  INV_X4 u1_gt_239_U775 ( .A(n8406), .ZN(u1_gt_239_n277) );
  NAND2_X2 u1_gt_239_U774 ( .A1(n8461), .A2(u1_gt_239_n277), .ZN(
        u1_gt_239_n421) );
  INV_X4 u1_gt_239_U773 ( .A(n8407), .ZN(u1_gt_239_n423) );
  NAND2_X2 u1_gt_239_U772 ( .A1(n8462), .A2(u1_gt_239_n423), .ZN(
        u1_gt_239_n473) );
  NAND2_X2 u1_gt_239_U771 ( .A1(u1_gt_239_n421), .A2(u1_gt_239_n473), .ZN(
        u1_gt_239_n821) );
  NOR2_X4 u1_gt_239_U770 ( .A1(u1_gt_239_n820), .A2(u1_gt_239_n821), .ZN(
        u1_gt_239_n819) );
  NAND3_X2 u1_gt_239_U769 ( .A1(u1_gt_239_n817), .A2(u1_gt_239_n818), .A3(
        u1_gt_239_n819), .ZN(u1_gt_239_n795) );
  INV_X4 u1_gt_239_U768 ( .A(n4285), .ZN(u1_gt_239_n816) );
  NAND2_X2 u1_gt_239_U767 ( .A1(n8453), .A2(u1_gt_239_n816), .ZN(
        u1_gt_239_n815) );
  NAND2_X2 u1_gt_239_U766 ( .A1(n4333), .A2(u1_gt_239_n815), .ZN(
        u1_gt_239_n811) );
  INV_X4 u1_gt_239_U765 ( .A(n8464), .ZN(u1_gt_239_n814) );
  NOR2_X4 u1_gt_239_U764 ( .A1(n4333), .A2(u1_gt_239_n814), .ZN(u1_gt_239_n813) );
  NOR3_X4 u1_gt_239_U763 ( .A1(u1_gt_239_n811), .A2(u1_gt_239_n812), .A3(
        u1_gt_239_n813), .ZN(u1_gt_239_n797) );
  INV_X4 u1_gt_239_U762 ( .A(n8442), .ZN(u1_gt_239_n802) );
  NAND2_X2 u1_gt_239_U761 ( .A1(n4397), .A2(u1_gt_239_n802), .ZN(
        u1_gt_239_n808) );
  INV_X4 u1_gt_239_U760 ( .A(n8453), .ZN(u1_gt_239_n810) );
  NAND2_X2 u1_gt_239_U759 ( .A1(n4285), .A2(u1_gt_239_n810), .ZN(
        u1_gt_239_n809) );
  NAND2_X2 u1_gt_239_U758 ( .A1(u1_gt_239_n808), .A2(u1_gt_239_n809), .ZN(
        u1_gt_239_n798) );
  INV_X4 u1_gt_239_U757 ( .A(n8360), .ZN(u1_gt_239_n807) );
  NAND2_X2 u1_gt_239_U756 ( .A1(n8413), .A2(u1_gt_239_n807), .ZN(
        u1_gt_239_n806) );
  INV_X4 u1_gt_239_U755 ( .A(u1_gt_239_n806), .ZN(u1_gt_239_n663) );
  INV_X4 u1_gt_239_U754 ( .A(n8359), .ZN(u1_gt_239_n805) );
  NAND2_X2 u1_gt_239_U753 ( .A1(n8412), .A2(u1_gt_239_n805), .ZN(
        u1_gt_239_n804) );
  INV_X4 u1_gt_239_U752 ( .A(u1_gt_239_n804), .ZN(u1_gt_239_n662) );
  INV_X4 u1_gt_239_U751 ( .A(n8358), .ZN(u1_gt_239_n114) );
  NAND2_X2 u1_gt_239_U750 ( .A1(n8411), .A2(u1_gt_239_n114), .ZN(
        u1_gt_239_n803) );
  INV_X4 u1_gt_239_U749 ( .A(u1_gt_239_n803), .ZN(u1_gt_239_n562) );
  INV_X4 u1_gt_239_U748 ( .A(n8367), .ZN(u1_gt_239_n653) );
  OAI211_X2 u1_gt_239_U747 ( .C1(u1_gt_239_n797), .C2(u1_gt_239_n798), .A(
        u1_gt_239_n799), .B(u1_gt_239_n800), .ZN(u1_gt_239_n796) );
  NOR3_X4 u1_gt_239_U746 ( .A1(u1_gt_239_n794), .A2(u1_gt_239_n795), .A3(
        u1_gt_239_n796), .ZN(u1_gt_239_n741) );
  NAND2_X2 u1_gt_239_U745 ( .A1(n8360), .A2(u1_gt_239_n26), .ZN(u1_gt_239_n793) );
  INV_X4 u1_gt_239_U744 ( .A(u1_gt_239_n113), .ZN(u1_gt_239_n582) );
  NAND2_X2 u1_gt_239_U743 ( .A1(u1_gt_239_n792), .A2(u1_gt_239_n582), .ZN(
        u1_gt_239_n788) );
  NOR2_X4 u1_gt_239_U742 ( .A1(u1_gt_239_n241), .A2(u1_gt_239_n204), .ZN(
        u1_gt_239_n791) );
  NAND2_X2 u1_gt_239_U741 ( .A1(u1_gt_239_n791), .A2(u1_gt_239_n223), .ZN(
        u1_gt_239_n789) );
  NAND2_X2 u1_gt_239_U740 ( .A1(u1_gt_239_n201), .A2(u1_gt_239_n222), .ZN(
        u1_gt_239_n790) );
  NOR3_X4 u1_gt_239_U739 ( .A1(u1_gt_239_n788), .A2(u1_gt_239_n789), .A3(
        u1_gt_239_n790), .ZN(u1_gt_239_n769) );
  INV_X4 u1_gt_239_U738 ( .A(u1_gt_239_n79), .ZN(u1_gt_239_n112) );
  NOR2_X4 u1_gt_239_U737 ( .A1(u1_gt_239_n137), .A2(u1_gt_239_n34), .ZN(
        u1_gt_239_n787) );
  NAND3_X2 u1_gt_239_U736 ( .A1(u1_gt_239_n785), .A2(u1_gt_239_n786), .A3(
        u1_gt_239_n787), .ZN(u1_gt_239_n783) );
  NAND2_X2 u1_gt_239_U735 ( .A1(u1_gt_239_n119), .A2(u1_gt_239_n13), .ZN(
        u1_gt_239_n784) );
  NOR3_X4 u1_gt_239_U734 ( .A1(u1_gt_239_n783), .A2(u1_gt_239_n16), .A3(
        u1_gt_239_n784), .ZN(u1_gt_239_n770) );
  NAND3_X2 u1_gt_239_U733 ( .A1(u1_gt_239_n567), .A2(u1_gt_239_n568), .A3(
        u1_gt_239_n569), .ZN(u1_gt_239_n779) );
  NAND2_X2 u1_gt_239_U732 ( .A1(u1_gt_239_n213), .A2(u1_gt_239_n566), .ZN(
        u1_gt_239_n780) );
  NOR3_X4 u1_gt_239_U731 ( .A1(u1_gt_239_n778), .A2(u1_gt_239_n779), .A3(
        u1_gt_239_n780), .ZN(u1_gt_239_n771) );
  INV_X4 u1_gt_239_U730 ( .A(u1_gt_239_n659), .ZN(u1_gt_239_n110) );
  INV_X4 u1_gt_239_U729 ( .A(u1_gt_239_n560), .ZN(u1_gt_239_n108) );
  INV_X4 u1_gt_239_U728 ( .A(u1_gt_239_n707), .ZN(u1_gt_239_n107) );
  NAND2_X2 u1_gt_239_U727 ( .A1(u1_gt_239_n776), .A2(u1_gt_239_n777), .ZN(
        u1_gt_239_n773) );
  NAND3_X2 u1_gt_239_U726 ( .A1(u1_gt_239_n421), .A2(u1_gt_239_n276), .A3(
        u1_gt_239_n473), .ZN(u1_gt_239_n774) );
  NAND2_X2 u1_gt_239_U725 ( .A1(u1_gt_239_n9), .A2(u1_gt_239_n232), .ZN(
        u1_gt_239_n775) );
  NOR3_X4 u1_gt_239_U724 ( .A1(u1_gt_239_n773), .A2(u1_gt_239_n774), .A3(
        u1_gt_239_n775), .ZN(u1_gt_239_n772) );
  NAND4_X2 u1_gt_239_U723 ( .A1(u1_gt_239_n769), .A2(u1_gt_239_n770), .A3(
        u1_gt_239_n771), .A4(u1_gt_239_n772), .ZN(u1_gt_239_n743) );
  INV_X4 u1_gt_239_U722 ( .A(u1_gt_239_n766), .ZN(u1_gt_239_n765) );
  NOR2_X4 u1_gt_239_U721 ( .A1(n8458), .A2(u1_gt_239_n765), .ZN(u1_gt_239_n764) );
  NAND2_X2 u1_gt_239_U720 ( .A1(u1_gt_239_n764), .A2(u1_gt_239_n235), .ZN(
        u1_gt_239_n762) );
  NAND2_X2 u1_gt_239_U719 ( .A1(u1_gt_239_n9), .A2(u1_gt_239_n232), .ZN(
        u1_gt_239_n763) );
  NOR3_X4 u1_gt_239_U718 ( .A1(u1_gt_239_n761), .A2(u1_gt_239_n762), .A3(
        u1_gt_239_n763), .ZN(u1_gt_239_n745) );
  NOR2_X4 u1_gt_239_U717 ( .A1(u1_gt_239_n87), .A2(u1_gt_239_n760), .ZN(
        u1_gt_239_n751) );
  INV_X4 u1_gt_239_U716 ( .A(u1_gt_239_n569), .ZN(u1_gt_239_n476) );
  INV_X4 u1_gt_239_U715 ( .A(u1_gt_239_n566), .ZN(u1_gt_239_n452) );
  NOR2_X4 u1_gt_239_U714 ( .A1(u1_gt_239_n476), .A2(u1_gt_239_n452), .ZN(
        u1_gt_239_n758) );
  INV_X4 u1_gt_239_U713 ( .A(u1_gt_239_n568), .ZN(u1_gt_239_n474) );
  INV_X4 u1_gt_239_U712 ( .A(u1_gt_239_n567), .ZN(u1_gt_239_n475) );
  NOR2_X4 u1_gt_239_U711 ( .A1(u1_gt_239_n474), .A2(u1_gt_239_n475), .ZN(
        u1_gt_239_n759) );
  NAND2_X2 u1_gt_239_U710 ( .A1(u1_gt_239_n758), .A2(u1_gt_239_n759), .ZN(
        u1_gt_239_n755) );
  NAND2_X2 u1_gt_239_U709 ( .A1(u1_gt_239_n192), .A2(u1_gt_239_n194), .ZN(
        u1_gt_239_n756) );
  NAND2_X2 u1_gt_239_U708 ( .A1(u1_gt_239_n24), .A2(u1_gt_239_n165), .ZN(
        u1_gt_239_n757) );
  NOR3_X4 u1_gt_239_U707 ( .A1(u1_gt_239_n755), .A2(u1_gt_239_n756), .A3(
        u1_gt_239_n757), .ZN(u1_gt_239_n752) );
  NAND2_X2 u1_gt_239_U706 ( .A1(n8446), .A2(u1_gt_239_n411), .ZN(
        u1_gt_239_n754) );
  AND4_X2 u1_gt_239_U705 ( .A1(u1_gt_239_n754), .A2(u1_gt_239_n245), .A3(
        u1_gt_239_n145), .A4(u1_gt_239_n25), .ZN(u1_gt_239_n753) );
  NAND3_X4 u1_gt_239_U704 ( .A1(u1_gt_239_n751), .A2(u1_gt_239_n752), .A3(
        u1_gt_239_n753), .ZN(u1_gt_239_n183) );
  NAND2_X2 u1_gt_239_U703 ( .A1(u1_gt_239_n222), .A2(n8403), .ZN(
        u1_gt_239_n748) );
  NOR3_X4 u1_gt_239_U702 ( .A1(u1_gt_239_n747), .A2(u1_gt_239_n748), .A3(
        u1_gt_239_n27), .ZN(u1_gt_239_n746) );
  NAND3_X2 u1_gt_239_U701 ( .A1(u1_gt_239_n745), .A2(u1_gt_239_n116), .A3(
        u1_gt_239_n746), .ZN(u1_gt_239_n744) );
  NAND2_X2 u1_gt_239_U700 ( .A1(u1_gt_239_n743), .A2(u1_gt_239_n744), .ZN(
        u1_gt_239_n742) );
  NAND2_X2 u1_gt_239_U699 ( .A1(u1_gt_239_n739), .A2(u1_gt_239_n740), .ZN(
        u1_gt_239_n737) );
  NAND2_X2 u1_gt_239_U698 ( .A1(u1_gt_239_n222), .A2(n8401), .ZN(
        u1_gt_239_n738) );
  NOR3_X4 u1_gt_239_U697 ( .A1(u1_gt_239_n737), .A2(u1_gt_239_n738), .A3(
        u1_gt_239_n27), .ZN(u1_gt_239_n729) );
  INV_X4 u1_gt_239_U696 ( .A(u1_gt_239_n232), .ZN(u1_gt_239_n102) );
  NAND2_X2 u1_gt_239_U695 ( .A1(u1_gt_239_n733), .A2(u1_gt_239_n734), .ZN(
        u1_gt_239_n732) );
  NOR2_X4 u1_gt_239_U694 ( .A1(u1_gt_239_n731), .A2(u1_gt_239_n732), .ZN(
        u1_gt_239_n730) );
  NAND3_X2 u1_gt_239_U693 ( .A1(u1_gt_239_n729), .A2(u1_gt_239_n116), .A3(
        u1_gt_239_n730), .ZN(u1_gt_239_n728) );
  INV_X4 u1_gt_239_U692 ( .A(u1_gt_239_n728), .ZN(u1_gt_239_n670) );
  NAND3_X2 u1_gt_239_U691 ( .A1(u1_gt_239_n245), .A2(u1_gt_239_n145), .A3(
        u1_gt_239_n144), .ZN(u1_gt_239_n726) );
  NOR2_X4 u1_gt_239_U690 ( .A1(u1_gt_239_n726), .A2(u1_gt_239_n727), .ZN(
        u1_gt_239_n725) );
  NAND2_X2 u1_gt_239_U689 ( .A1(u1_gt_239_n725), .A2(u1_gt_239_n582), .ZN(
        u1_gt_239_n721) );
  NOR2_X4 u1_gt_239_U688 ( .A1(u1_gt_239_n241), .A2(u1_gt_239_n204), .ZN(
        u1_gt_239_n724) );
  NAND2_X2 u1_gt_239_U687 ( .A1(u1_gt_239_n724), .A2(u1_gt_239_n223), .ZN(
        u1_gt_239_n722) );
  NAND2_X2 u1_gt_239_U686 ( .A1(u1_gt_239_n201), .A2(u1_gt_239_n222), .ZN(
        u1_gt_239_n723) );
  NOR3_X4 u1_gt_239_U685 ( .A1(u1_gt_239_n721), .A2(u1_gt_239_n722), .A3(
        u1_gt_239_n723), .ZN(u1_gt_239_n700) );
  NAND3_X2 u1_gt_239_U684 ( .A1(u1_gt_239_n718), .A2(u1_gt_239_n719), .A3(
        u1_gt_239_n720), .ZN(u1_gt_239_n716) );
  NAND2_X2 u1_gt_239_U683 ( .A1(u1_gt_239_n18), .A2(u1_gt_239_n13), .ZN(
        u1_gt_239_n717) );
  NOR3_X4 u1_gt_239_U682 ( .A1(u1_gt_239_n716), .A2(u1_gt_239_n16), .A3(
        u1_gt_239_n717), .ZN(u1_gt_239_n701) );
  NAND2_X2 u1_gt_239_U681 ( .A1(u1_gt_239_n714), .A2(u1_gt_239_n715), .ZN(
        u1_gt_239_n710) );
  NOR2_X4 u1_gt_239_U680 ( .A1(u1_gt_239_n103), .A2(u1_gt_239_n104), .ZN(
        u1_gt_239_n713) );
  NAND2_X2 u1_gt_239_U679 ( .A1(u1_gt_239_n713), .A2(u1_gt_239_n342), .ZN(
        u1_gt_239_n711) );
  NAND2_X2 u1_gt_239_U678 ( .A1(u1_gt_239_n194), .A2(u1_gt_239_n11), .ZN(
        u1_gt_239_n712) );
  NOR3_X4 u1_gt_239_U677 ( .A1(u1_gt_239_n710), .A2(u1_gt_239_n711), .A3(
        u1_gt_239_n712), .ZN(u1_gt_239_n702) );
  NOR3_X4 u1_gt_239_U676 ( .A1(n8431), .A2(u1_gt_239_n663), .A3(u1_gt_239_n1), 
        .ZN(u1_gt_239_n709) );
  NAND2_X2 u1_gt_239_U675 ( .A1(u1_gt_239_n708), .A2(u1_gt_239_n709), .ZN(
        u1_gt_239_n704) );
  NAND3_X2 u1_gt_239_U674 ( .A1(u1_gt_239_n276), .A2(u1_gt_239_n421), .A3(
        u1_gt_239_n473), .ZN(u1_gt_239_n705) );
  NAND2_X2 u1_gt_239_U673 ( .A1(u1_gt_239_n659), .A2(u1_gt_239_n707), .ZN(
        u1_gt_239_n706) );
  NOR3_X4 u1_gt_239_U672 ( .A1(u1_gt_239_n704), .A2(u1_gt_239_n705), .A3(
        u1_gt_239_n706), .ZN(u1_gt_239_n703) );
  NAND4_X2 u1_gt_239_U671 ( .A1(u1_gt_239_n700), .A2(u1_gt_239_n701), .A3(
        u1_gt_239_n702), .A4(u1_gt_239_n703), .ZN(u1_gt_239_n672) );
  NAND2_X2 u1_gt_239_U670 ( .A1(u1_gt_239_n698), .A2(u1_gt_239_n582), .ZN(
        u1_gt_239_n694) );
  NOR2_X4 u1_gt_239_U669 ( .A1(u1_gt_239_n87), .A2(u1_gt_239_n86), .ZN(
        u1_gt_239_n697) );
  NAND2_X2 u1_gt_239_U668 ( .A1(u1_gt_239_n697), .A2(u1_gt_239_n223), .ZN(
        u1_gt_239_n695) );
  NAND2_X2 u1_gt_239_U667 ( .A1(u1_gt_239_n222), .A2(u1_gt_239_n77), .ZN(
        u1_gt_239_n696) );
  NOR3_X4 u1_gt_239_U666 ( .A1(u1_gt_239_n694), .A2(u1_gt_239_n695), .A3(
        u1_gt_239_n696), .ZN(u1_gt_239_n674) );
  NOR2_X4 u1_gt_239_U665 ( .A1(u1_gt_239_n142), .A2(u1_gt_239_n141), .ZN(
        u1_gt_239_n692) );
  NAND2_X2 u1_gt_239_U664 ( .A1(u1_gt_239_n690), .A2(u1_gt_239_n691), .ZN(
        u1_gt_239_n689) );
  NOR2_X4 u1_gt_239_U663 ( .A1(u1_gt_239_n688), .A2(u1_gt_239_n689), .ZN(
        u1_gt_239_n675) );
  NAND3_X2 u1_gt_239_U662 ( .A1(u1_gt_239_n213), .A2(u1_gt_239_n566), .A3(
        u1_gt_239_n212), .ZN(u1_gt_239_n684) );
  NOR2_X4 u1_gt_239_U661 ( .A1(u1_gt_239_n683), .A2(u1_gt_239_n684), .ZN(
        u1_gt_239_n676) );
  INV_X4 u1_gt_239_U660 ( .A(u1_gt_239_n421), .ZN(u1_gt_239_n111) );
  INV_X4 u1_gt_239_U659 ( .A(u1_gt_239_n276), .ZN(u1_gt_239_n101) );
  NOR2_X4 u1_gt_239_U658 ( .A1(u1_gt_239_n111), .A2(u1_gt_239_n101), .ZN(
        u1_gt_239_n681) );
  NAND3_X2 u1_gt_239_U657 ( .A1(u1_gt_239_n569), .A2(u1_gt_239_n567), .A3(
        u1_gt_239_n9), .ZN(u1_gt_239_n679) );
  NAND2_X2 u1_gt_239_U656 ( .A1(u1_gt_239_n568), .A2(u1_gt_239_n232), .ZN(
        u1_gt_239_n680) );
  NOR3_X4 u1_gt_239_U655 ( .A1(u1_gt_239_n678), .A2(u1_gt_239_n679), .A3(
        u1_gt_239_n680), .ZN(u1_gt_239_n677) );
  NAND4_X2 u1_gt_239_U654 ( .A1(u1_gt_239_n674), .A2(u1_gt_239_n675), .A3(
        u1_gt_239_n676), .A4(u1_gt_239_n677), .ZN(u1_gt_239_n673) );
  NAND2_X2 u1_gt_239_U653 ( .A1(u1_gt_239_n672), .A2(u1_gt_239_n673), .ZN(
        u1_gt_239_n671) );
  NOR2_X4 u1_gt_239_U652 ( .A1(u1_gt_239_n103), .A2(u1_gt_239_n104), .ZN(
        u1_gt_239_n667) );
  NAND2_X2 u1_gt_239_U651 ( .A1(u1_gt_239_n667), .A2(u1_gt_239_n342), .ZN(
        u1_gt_239_n665) );
  NAND2_X2 u1_gt_239_U650 ( .A1(u1_gt_239_n194), .A2(u1_gt_239_n11), .ZN(
        u1_gt_239_n666) );
  NOR3_X4 u1_gt_239_U649 ( .A1(u1_gt_239_n664), .A2(u1_gt_239_n665), .A3(
        u1_gt_239_n666), .ZN(u1_gt_239_n654) );
  NOR3_X4 u1_gt_239_U648 ( .A1(u1_gt_239_n662), .A2(n8420), .A3(u1_gt_239_n663), .ZN(u1_gt_239_n661) );
  NAND2_X2 u1_gt_239_U647 ( .A1(u1_gt_239_n660), .A2(u1_gt_239_n661), .ZN(
        u1_gt_239_n656) );
  NAND3_X2 u1_gt_239_U646 ( .A1(u1_gt_239_n232), .A2(u1_gt_239_n276), .A3(
        u1_gt_239_n473), .ZN(u1_gt_239_n657) );
  NAND2_X2 u1_gt_239_U645 ( .A1(u1_gt_239_n421), .A2(u1_gt_239_n659), .ZN(
        u1_gt_239_n658) );
  NOR3_X4 u1_gt_239_U644 ( .A1(u1_gt_239_n656), .A2(u1_gt_239_n657), .A3(
        u1_gt_239_n658), .ZN(u1_gt_239_n655) );
  NAND2_X2 u1_gt_239_U643 ( .A1(u1_gt_239_n654), .A2(u1_gt_239_n655), .ZN(
        u1_gt_239_n601) );
  NAND2_X2 u1_gt_239_U642 ( .A1(u1_gt_239_n651), .A2(u1_gt_239_n652), .ZN(
        u1_gt_239_n650) );
  NAND2_X2 u1_gt_239_U641 ( .A1(u1_gt_239_n201), .A2(u1_gt_239_n222), .ZN(
        u1_gt_239_n648) );
  NAND2_X2 u1_gt_239_U640 ( .A1(u1_gt_239_n77), .A2(u1_gt_239_n78), .ZN(
        u1_gt_239_n649) );
  NOR3_X4 u1_gt_239_U639 ( .A1(u1_gt_239_n648), .A2(u1_gt_239_n27), .A3(
        u1_gt_239_n649), .ZN(u1_gt_239_n641) );
  NOR3_X4 u1_gt_239_U638 ( .A1(u1_gt_239_n345), .A2(u1_gt_239_n142), .A3(
        u1_gt_239_n141), .ZN(u1_gt_239_n645) );
  NOR3_X4 u1_gt_239_U637 ( .A1(u1_gt_239_n20), .A2(u1_gt_239_n163), .A3(
        u1_gt_239_n22), .ZN(u1_gt_239_n646) );
  NOR2_X4 u1_gt_239_U636 ( .A1(u1_gt_239_n137), .A2(u1_gt_239_n34), .ZN(
        u1_gt_239_n647) );
  NAND3_X2 u1_gt_239_U635 ( .A1(u1_gt_239_n645), .A2(u1_gt_239_n646), .A3(
        u1_gt_239_n647), .ZN(u1_gt_239_n643) );
  NAND2_X2 u1_gt_239_U634 ( .A1(u1_gt_239_n119), .A2(u1_gt_239_n13), .ZN(
        u1_gt_239_n644) );
  NOR3_X4 u1_gt_239_U633 ( .A1(u1_gt_239_n643), .A2(u1_gt_239_n16), .A3(
        u1_gt_239_n644), .ZN(u1_gt_239_n642) );
  NAND3_X2 u1_gt_239_U632 ( .A1(u1_gt_239_n640), .A2(u1_gt_239_n641), .A3(
        u1_gt_239_n642), .ZN(u1_gt_239_n602) );
  NAND2_X2 u1_gt_239_U631 ( .A1(u1_gt_239_n13), .A2(u1_gt_239_n18), .ZN(
        u1_gt_239_n639) );
  NAND2_X2 u1_gt_239_U630 ( .A1(u1_gt_239_n638), .A2(u1_gt_239_n223), .ZN(
        u1_gt_239_n633) );
  NOR2_X4 u1_gt_239_U629 ( .A1(u1_gt_239_n637), .A2(u1_gt_239_n31), .ZN(
        u1_gt_239_n635) );
  NOR3_X4 u1_gt_239_U628 ( .A1(u1_gt_239_n633), .A2(u1_gt_239_n634), .A3(
        u1_gt_239_n29), .ZN(u1_gt_239_n624) );
  NOR3_X4 u1_gt_239_U627 ( .A1(u1_gt_239_n10), .A2(u1_gt_239_n163), .A3(
        u1_gt_239_n162), .ZN(u1_gt_239_n632) );
  NAND3_X2 u1_gt_239_U626 ( .A1(u1_gt_239_n630), .A2(u1_gt_239_n631), .A3(
        u1_gt_239_n632), .ZN(u1_gt_239_n626) );
  NAND2_X2 u1_gt_239_U625 ( .A1(u1_gt_239_n628), .A2(u1_gt_239_n629), .ZN(
        u1_gt_239_n627) );
  NOR2_X4 u1_gt_239_U624 ( .A1(u1_gt_239_n626), .A2(u1_gt_239_n627), .ZN(
        u1_gt_239_n625) );
  NAND3_X2 u1_gt_239_U623 ( .A1(u1_gt_239_n623), .A2(u1_gt_239_n624), .A3(
        u1_gt_239_n625), .ZN(u1_gt_239_n603) );
  NOR2_X4 u1_gt_239_U622 ( .A1(u1_gt_239_n87), .A2(u1_gt_239_n86), .ZN(
        u1_gt_239_n622) );
  NAND2_X2 u1_gt_239_U621 ( .A1(u1_gt_239_n222), .A2(u1_gt_239_n622), .ZN(
        u1_gt_239_n620) );
  NAND3_X2 u1_gt_239_U620 ( .A1(u1_gt_239_n245), .A2(n8397), .A3(u1_gt_239_n25), .ZN(u1_gt_239_n621) );
  NOR3_X4 u1_gt_239_U619 ( .A1(u1_gt_239_n620), .A2(u1_gt_239_n621), .A3(
        u1_gt_239_n27), .ZN(u1_gt_239_n605) );
  NOR2_X4 u1_gt_239_U618 ( .A1(u1_gt_239_n204), .A2(u1_gt_239_n241), .ZN(
        u1_gt_239_n618) );
  NOR2_X4 u1_gt_239_U617 ( .A1(u1_gt_239_n136), .A2(u1_gt_239_n137), .ZN(
        u1_gt_239_n619) );
  NAND2_X2 u1_gt_239_U616 ( .A1(u1_gt_239_n18), .A2(u1_gt_239_n17), .ZN(
        u1_gt_239_n617) );
  NOR2_X4 u1_gt_239_U615 ( .A1(u1_gt_239_n616), .A2(u1_gt_239_n617), .ZN(
        u1_gt_239_n606) );
  NAND2_X2 u1_gt_239_U614 ( .A1(u1_gt_239_n614), .A2(u1_gt_239_n615), .ZN(
        u1_gt_239_n612) );
  NAND3_X2 u1_gt_239_U613 ( .A1(u1_gt_239_n197), .A2(u1_gt_239_n165), .A3(
        u1_gt_239_n24), .ZN(u1_gt_239_n613) );
  NOR2_X4 u1_gt_239_U612 ( .A1(u1_gt_239_n612), .A2(u1_gt_239_n613), .ZN(
        u1_gt_239_n607) );
  INV_X4 u1_gt_239_U611 ( .A(n8451), .ZN(u1_gt_239_n611) );
  NAND4_X2 u1_gt_239_U610 ( .A1(u1_gt_239_n213), .A2(u1_gt_239_n566), .A3(
        u1_gt_239_n569), .A4(u1_gt_239_n611), .ZN(u1_gt_239_n609) );
  NAND3_X2 u1_gt_239_U609 ( .A1(u1_gt_239_n342), .A2(u1_gt_239_n212), .A3(
        u1_gt_239_n11), .ZN(u1_gt_239_n610) );
  NOR2_X4 u1_gt_239_U608 ( .A1(u1_gt_239_n609), .A2(u1_gt_239_n610), .ZN(
        u1_gt_239_n608) );
  NAND4_X2 u1_gt_239_U607 ( .A1(u1_gt_239_n605), .A2(u1_gt_239_n606), .A3(
        u1_gt_239_n607), .A4(u1_gt_239_n608), .ZN(u1_gt_239_n604) );
  OAI211_X2 u1_gt_239_U606 ( .C1(u1_gt_239_n601), .C2(u1_gt_239_n602), .A(
        u1_gt_239_n603), .B(u1_gt_239_n604), .ZN(u1_gt_239_n549) );
  INV_X4 u1_gt_239_U605 ( .A(n8366), .ZN(u1_gt_239_n585) );
  INV_X4 u1_gt_239_U604 ( .A(n8421), .ZN(u1_gt_239_n59) );
  NAND2_X2 u1_gt_239_U603 ( .A1(n8368), .A2(u1_gt_239_n59), .ZN(u1_gt_239_n586) );
  INV_X4 u1_gt_239_U602 ( .A(n8416), .ZN(u1_gt_239_n599) );
  NAND2_X2 u1_gt_239_U601 ( .A1(n8363), .A2(u1_gt_239_n599), .ZN(
        u1_gt_239_n596) );
  INV_X4 u1_gt_239_U600 ( .A(n8415), .ZN(u1_gt_239_n598) );
  NAND2_X2 u1_gt_239_U599 ( .A1(n8362), .A2(u1_gt_239_n598), .ZN(
        u1_gt_239_n597) );
  NAND2_X2 u1_gt_239_U598 ( .A1(u1_gt_239_n596), .A2(u1_gt_239_n597), .ZN(
        u1_gt_239_n595) );
  NOR2_X4 u1_gt_239_U597 ( .A1(u1_gt_239_n2), .A2(u1_gt_239_n595), .ZN(
        u1_gt_239_n588) );
  INV_X4 u1_gt_239_U596 ( .A(n8363), .ZN(u1_gt_239_n594) );
  NAND2_X2 u1_gt_239_U595 ( .A1(n8416), .A2(u1_gt_239_n594), .ZN(u1_gt_239_n52) );
  INV_X4 u1_gt_239_U594 ( .A(n8417), .ZN(u1_gt_239_n593) );
  NAND3_X2 u1_gt_239_U593 ( .A1(u1_gt_239_n52), .A2(u1_gt_239_n593), .A3(n8364), .ZN(u1_gt_239_n589) );
  INV_X4 u1_gt_239_U592 ( .A(n8364), .ZN(u1_gt_239_n592) );
  NAND2_X2 u1_gt_239_U591 ( .A1(n8417), .A2(u1_gt_239_n592), .ZN(u1_gt_239_n53) );
  INV_X4 u1_gt_239_U590 ( .A(n8418), .ZN(u1_gt_239_n591) );
  NAND4_X2 u1_gt_239_U589 ( .A1(n8365), .A2(u1_gt_239_n52), .A3(u1_gt_239_n53), 
        .A4(u1_gt_239_n591), .ZN(u1_gt_239_n590) );
  NAND3_X4 u1_gt_239_U588 ( .A1(u1_gt_239_n588), .A2(u1_gt_239_n589), .A3(
        u1_gt_239_n590), .ZN(u1_gt_239_n45) );
  INV_X4 u1_gt_239_U587 ( .A(u1_gt_239_n45), .ZN(u1_gt_239_n587) );
  OAI211_X2 u1_gt_239_U586 ( .C1(n8419), .C2(u1_gt_239_n585), .A(
        u1_gt_239_n586), .B(u1_gt_239_n587), .ZN(u1_gt_239_n584) );
  INV_X4 u1_gt_239_U585 ( .A(u1_gt_239_n584), .ZN(u1_gt_239_n58) );
  NAND2_X2 u1_gt_239_U584 ( .A1(n8359), .A2(u1_gt_239_n144), .ZN(
        u1_gt_239_n583) );
  NAND2_X2 u1_gt_239_U583 ( .A1(u1_gt_239_n581), .A2(u1_gt_239_n582), .ZN(
        u1_gt_239_n577) );
  NAND2_X2 u1_gt_239_U582 ( .A1(u1_gt_239_n580), .A2(u1_gt_239_n223), .ZN(
        u1_gt_239_n578) );
  NAND2_X2 u1_gt_239_U581 ( .A1(u1_gt_239_n201), .A2(u1_gt_239_n222), .ZN(
        u1_gt_239_n579) );
  NOR3_X4 u1_gt_239_U580 ( .A1(u1_gt_239_n577), .A2(u1_gt_239_n578), .A3(
        u1_gt_239_n579), .ZN(u1_gt_239_n552) );
  NAND3_X2 u1_gt_239_U579 ( .A1(u1_gt_239_n574), .A2(u1_gt_239_n575), .A3(
        u1_gt_239_n576), .ZN(u1_gt_239_n572) );
  NAND2_X2 u1_gt_239_U578 ( .A1(u1_gt_239_n119), .A2(u1_gt_239_n13), .ZN(
        u1_gt_239_n573) );
  NOR3_X4 u1_gt_239_U577 ( .A1(u1_gt_239_n572), .A2(u1_gt_239_n16), .A3(
        u1_gt_239_n573), .ZN(u1_gt_239_n553) );
  NAND3_X2 u1_gt_239_U576 ( .A1(u1_gt_239_n567), .A2(u1_gt_239_n568), .A3(
        u1_gt_239_n569), .ZN(u1_gt_239_n564) );
  NAND2_X2 u1_gt_239_U575 ( .A1(u1_gt_239_n213), .A2(u1_gt_239_n566), .ZN(
        u1_gt_239_n565) );
  NOR3_X4 u1_gt_239_U574 ( .A1(u1_gt_239_n563), .A2(u1_gt_239_n564), .A3(
        u1_gt_239_n565), .ZN(u1_gt_239_n554) );
  NAND3_X2 u1_gt_239_U573 ( .A1(u1_gt_239_n421), .A2(u1_gt_239_n276), .A3(
        u1_gt_239_n473), .ZN(u1_gt_239_n557) );
  NAND2_X2 u1_gt_239_U572 ( .A1(u1_gt_239_n9), .A2(u1_gt_239_n232), .ZN(
        u1_gt_239_n558) );
  NOR3_X4 u1_gt_239_U571 ( .A1(u1_gt_239_n556), .A2(u1_gt_239_n557), .A3(
        u1_gt_239_n558), .ZN(u1_gt_239_n555) );
  NAND4_X2 u1_gt_239_U570 ( .A1(u1_gt_239_n552), .A2(u1_gt_239_n553), .A3(
        u1_gt_239_n554), .A4(u1_gt_239_n555), .ZN(u1_gt_239_n551) );
  NAND2_X2 u1_gt_239_U569 ( .A1(u1_gt_239_n58), .A2(u1_gt_239_n551), .ZN(
        u1_gt_239_n550) );
  NAND3_X2 u1_gt_239_U568 ( .A1(u1_gt_239_n546), .A2(u1_gt_239_n547), .A3(
        u1_gt_239_n548), .ZN(u1_gt_239_n379) );
  NAND3_X2 u1_gt_239_U567 ( .A1(u1_gt_239_n13), .A2(u1_gt_239_n18), .A3(
        u1_gt_239_n15), .ZN(u1_gt_239_n545) );
  NOR3_X4 u1_gt_239_U566 ( .A1(u1_gt_239_n545), .A2(u1_gt_239_n33), .A3(
        u1_gt_239_n27), .ZN(u1_gt_239_n544) );
  NAND2_X2 u1_gt_239_U565 ( .A1(u1_gt_239_n544), .A2(u1_gt_239_n116), .ZN(
        u1_gt_239_n534) );
  INV_X4 u1_gt_239_U564 ( .A(n8460), .ZN(u1_gt_239_n542) );
  NAND3_X2 u1_gt_239_U563 ( .A1(u1_gt_239_n232), .A2(u1_gt_239_n542), .A3(
        u1_gt_239_n9), .ZN(u1_gt_239_n540) );
  NAND2_X2 u1_gt_239_U562 ( .A1(u1_gt_239_n212), .A2(u1_gt_239_n213), .ZN(
        u1_gt_239_n541) );
  NAND2_X2 u1_gt_239_U561 ( .A1(u1_gt_239_n121), .A2(u1_gt_239_n11), .ZN(
        u1_gt_239_n539) );
  NAND3_X2 u1_gt_239_U560 ( .A1(u1_gt_239_n536), .A2(u1_gt_239_n537), .A3(
        u1_gt_239_n538), .ZN(u1_gt_239_n535) );
  NOR2_X4 u1_gt_239_U559 ( .A1(u1_gt_239_n534), .A2(u1_gt_239_n535), .ZN(
        u1_gt_239_n518) );
  NAND2_X2 u1_gt_239_U558 ( .A1(u1_gt_239_n144), .A2(u1_gt_239_n145), .ZN(
        u1_gt_239_n532) );
  NAND2_X2 u1_gt_239_U557 ( .A1(u1_gt_239_n530), .A2(u1_gt_239_n531), .ZN(
        u1_gt_239_n520) );
  INV_X4 u1_gt_239_U556 ( .A(n8434), .ZN(u1_gt_239_n526) );
  NAND3_X2 u1_gt_239_U555 ( .A1(u1_gt_239_n15), .A2(u1_gt_239_n526), .A3(
        u1_gt_239_n79), .ZN(u1_gt_239_n524) );
  NAND2_X2 u1_gt_239_U554 ( .A1(u1_gt_239_n77), .A2(u1_gt_239_n78), .ZN(
        u1_gt_239_n525) );
  NAND2_X2 u1_gt_239_U553 ( .A1(u1_gt_239_n522), .A2(u1_gt_239_n523), .ZN(
        u1_gt_239_n521) );
  NAND2_X2 u1_gt_239_U552 ( .A1(u1_gt_239_n520), .A2(u1_gt_239_n521), .ZN(
        u1_gt_239_n519) );
  NAND2_X2 u1_gt_239_U551 ( .A1(u1_gt_239_n25), .A2(u1_gt_239_n145), .ZN(
        u1_gt_239_n516) );
  NAND2_X2 u1_gt_239_U550 ( .A1(u1_gt_239_n512), .A2(u1_gt_239_n513), .ZN(
        u1_gt_239_n511) );
  NOR2_X4 u1_gt_239_U549 ( .A1(u1_gt_239_n510), .A2(u1_gt_239_n511), .ZN(
        u1_gt_239_n509) );
  NAND3_X2 u1_gt_239_U548 ( .A1(u1_gt_239_n507), .A2(u1_gt_239_n508), .A3(
        u1_gt_239_n509), .ZN(u1_gt_239_n506) );
  INV_X4 u1_gt_239_U547 ( .A(u1_gt_239_n506), .ZN(u1_gt_239_n491) );
  INV_X4 u1_gt_239_U546 ( .A(n8425), .ZN(u1_gt_239_n505) );
  NAND2_X2 u1_gt_239_U545 ( .A1(u1_gt_239_n26), .A2(u1_gt_239_n505), .ZN(
        u1_gt_239_n503) );
  NAND3_X2 u1_gt_239_U544 ( .A1(u1_gt_239_n500), .A2(u1_gt_239_n501), .A3(
        u1_gt_239_n502), .ZN(u1_gt_239_n494) );
  NAND2_X2 u1_gt_239_U543 ( .A1(u1_gt_239_n223), .A2(u1_gt_239_n498), .ZN(
        u1_gt_239_n495) );
  NAND2_X2 u1_gt_239_U542 ( .A1(u1_gt_239_n222), .A2(u1_gt_239_n497), .ZN(
        u1_gt_239_n496) );
  NOR3_X4 u1_gt_239_U541 ( .A1(u1_gt_239_n494), .A2(u1_gt_239_n495), .A3(
        u1_gt_239_n496), .ZN(u1_gt_239_n493) );
  NAND2_X2 u1_gt_239_U540 ( .A1(u1_gt_239_n489), .A2(u1_gt_239_n490), .ZN(
        u1_gt_239_n380) );
  NAND2_X2 u1_gt_239_U539 ( .A1(u1_gt_239_n145), .A2(u1_gt_239_n201), .ZN(
        u1_gt_239_n488) );
  NOR2_X4 u1_gt_239_U538 ( .A1(u1_gt_239_n28), .A2(u1_gt_239_n488), .ZN(
        u1_gt_239_n478) );
  NAND3_X2 u1_gt_239_U537 ( .A1(u1_gt_239_n245), .A2(u1_gt_239_n25), .A3(n8408), .ZN(u1_gt_239_n487) );
  NAND2_X2 u1_gt_239_U536 ( .A1(u1_gt_239_n483), .A2(u1_gt_239_n484), .ZN(
        u1_gt_239_n482) );
  NOR2_X4 u1_gt_239_U535 ( .A1(u1_gt_239_n481), .A2(u1_gt_239_n482), .ZN(
        u1_gt_239_n480) );
  NAND4_X2 u1_gt_239_U534 ( .A1(u1_gt_239_n477), .A2(u1_gt_239_n478), .A3(
        u1_gt_239_n479), .A4(u1_gt_239_n480), .ZN(u1_gt_239_n462) );
  INV_X4 u1_gt_239_U533 ( .A(u1_gt_239_n473), .ZN(u1_gt_239_n109) );
  NAND4_X2 u1_gt_239_U532 ( .A1(u1_gt_239_n469), .A2(u1_gt_239_n470), .A3(
        u1_gt_239_n471), .A4(u1_gt_239_n472), .ZN(u1_gt_239_n463) );
  NOR2_X4 u1_gt_239_U531 ( .A1(u1_gt_239_n160), .A2(u1_gt_239_n10), .ZN(
        u1_gt_239_n465) );
  NAND2_X2 u1_gt_239_U530 ( .A1(u1_gt_239_n192), .A2(u1_gt_239_n194), .ZN(
        u1_gt_239_n468) );
  NAND3_X2 u1_gt_239_U529 ( .A1(u1_gt_239_n465), .A2(u1_gt_239_n466), .A3(
        u1_gt_239_n467), .ZN(u1_gt_239_n464) );
  NOR3_X4 u1_gt_239_U528 ( .A1(u1_gt_239_n462), .A2(u1_gt_239_n463), .A3(
        u1_gt_239_n464), .ZN(u1_gt_239_n427) );
  NOR2_X4 u1_gt_239_U527 ( .A1(u1_gt_239_n461), .A2(u1_gt_239_n31), .ZN(
        u1_gt_239_n459) );
  NAND2_X2 u1_gt_239_U526 ( .A1(u1_gt_239_n77), .A2(u1_gt_239_n78), .ZN(
        u1_gt_239_n457) );
  NAND2_X2 u1_gt_239_U525 ( .A1(u1_gt_239_n13), .A2(u1_gt_239_n119), .ZN(
        u1_gt_239_n456) );
  NOR3_X4 u1_gt_239_U524 ( .A1(u1_gt_239_n456), .A2(u1_gt_239_n137), .A3(
        u1_gt_239_n33), .ZN(u1_gt_239_n455) );
  NAND3_X4 u1_gt_239_U523 ( .A1(u1_gt_239_n453), .A2(u1_gt_239_n454), .A3(
        u1_gt_239_n455), .ZN(u1_gt_239_n443) );
  NAND3_X2 u1_gt_239_U522 ( .A1(u1_gt_239_n449), .A2(u1_gt_239_n450), .A3(
        u1_gt_239_n451), .ZN(u1_gt_239_n444) );
  NAND3_X2 u1_gt_239_U521 ( .A1(u1_gt_239_n446), .A2(u1_gt_239_n447), .A3(
        u1_gt_239_n448), .ZN(u1_gt_239_n445) );
  NOR3_X4 u1_gt_239_U520 ( .A1(u1_gt_239_n443), .A2(u1_gt_239_n444), .A3(
        u1_gt_239_n445), .ZN(u1_gt_239_n428) );
  NOR2_X4 u1_gt_239_U519 ( .A1(u1_gt_239_n136), .A2(u1_gt_239_n137), .ZN(
        u1_gt_239_n441) );
  NAND4_X2 u1_gt_239_U518 ( .A1(u1_gt_239_n439), .A2(u1_gt_239_n440), .A3(
        u1_gt_239_n441), .A4(u1_gt_239_n442), .ZN(u1_gt_239_n430) );
  INV_X4 u1_gt_239_U517 ( .A(u1_gt_239_n437), .ZN(u1_gt_239_n435) );
  NAND2_X2 u1_gt_239_U516 ( .A1(u1_gt_239_n145), .A2(u1_gt_239_n25), .ZN(
        u1_gt_239_n436) );
  NOR2_X4 u1_gt_239_U515 ( .A1(u1_gt_239_n435), .A2(u1_gt_239_n436), .ZN(
        u1_gt_239_n434) );
  NAND2_X2 u1_gt_239_U514 ( .A1(u1_gt_239_n434), .A2(u1_gt_239_n223), .ZN(
        u1_gt_239_n431) );
  NAND2_X2 u1_gt_239_U513 ( .A1(u1_gt_239_n222), .A2(u1_gt_239_n433), .ZN(
        u1_gt_239_n432) );
  NOR3_X4 u1_gt_239_U512 ( .A1(u1_gt_239_n430), .A2(u1_gt_239_n431), .A3(
        u1_gt_239_n432), .ZN(u1_gt_239_n429) );
  NAND3_X2 u1_gt_239_U511 ( .A1(u1_gt_239_n119), .A2(u1_gt_239_n13), .A3(
        u1_gt_239_n17), .ZN(u1_gt_239_n425) );
  NAND2_X2 u1_gt_239_U510 ( .A1(u1_gt_239_n79), .A2(u1_gt_239_n15), .ZN(
        u1_gt_239_n426) );
  NAND2_X2 u1_gt_239_U509 ( .A1(u1_gt_239_n424), .A2(u1_gt_239_n116), .ZN(
        u1_gt_239_n412) );
  NOR2_X4 u1_gt_239_U508 ( .A1(u1_gt_239_n113), .A2(u1_gt_239_n423), .ZN(
        u1_gt_239_n415) );
  NAND3_X2 u1_gt_239_U507 ( .A1(u1_gt_239_n120), .A2(u1_gt_239_n121), .A3(
        u1_gt_239_n11), .ZN(u1_gt_239_n418) );
  NAND2_X2 u1_gt_239_U506 ( .A1(u1_gt_239_n212), .A2(u1_gt_239_n213), .ZN(
        u1_gt_239_n419) );
  NOR3_X4 u1_gt_239_U505 ( .A1(u1_gt_239_n417), .A2(u1_gt_239_n418), .A3(
        u1_gt_239_n419), .ZN(u1_gt_239_n416) );
  NAND3_X2 u1_gt_239_U504 ( .A1(u1_gt_239_n414), .A2(u1_gt_239_n415), .A3(
        u1_gt_239_n416), .ZN(u1_gt_239_n413) );
  NOR2_X4 u1_gt_239_U503 ( .A1(u1_gt_239_n412), .A2(u1_gt_239_n413), .ZN(
        u1_gt_239_n384) );
  NOR3_X4 u1_gt_239_U502 ( .A1(u1_gt_239_n28), .A2(u1_gt_239_n204), .A3(
        u1_gt_239_n29), .ZN(u1_gt_239_n398) );
  NOR3_X4 u1_gt_239_U501 ( .A1(u1_gt_239_n87), .A2(u1_gt_239_n30), .A3(
        u1_gt_239_n411), .ZN(u1_gt_239_n410) );
  NAND3_X2 u1_gt_239_U500 ( .A1(u1_gt_239_n409), .A2(u1_gt_239_n410), .A3(
        u1_gt_239_n79), .ZN(u1_gt_239_n407) );
  NAND2_X2 u1_gt_239_U499 ( .A1(u1_gt_239_n78), .A2(u1_gt_239_n15), .ZN(
        u1_gt_239_n408) );
  NOR2_X4 u1_gt_239_U498 ( .A1(u1_gt_239_n407), .A2(u1_gt_239_n408), .ZN(
        u1_gt_239_n399) );
  NOR2_X4 u1_gt_239_U497 ( .A1(u1_gt_239_n142), .A2(u1_gt_239_n141), .ZN(
        u1_gt_239_n406) );
  NAND3_X2 u1_gt_239_U496 ( .A1(u1_gt_239_n406), .A2(u1_gt_239_n24), .A3(
        u1_gt_239_n17), .ZN(u1_gt_239_n405) );
  NOR3_X4 u1_gt_239_U495 ( .A1(u1_gt_239_n405), .A2(u1_gt_239_n136), .A3(
        u1_gt_239_n135), .ZN(u1_gt_239_n400) );
  INV_X4 u1_gt_239_U494 ( .A(n8446), .ZN(u1_gt_239_n404) );
  NAND3_X2 u1_gt_239_U493 ( .A1(u1_gt_239_n194), .A2(u1_gt_239_n404), .A3(
        u1_gt_239_n11), .ZN(u1_gt_239_n402) );
  NAND3_X2 u1_gt_239_U492 ( .A1(u1_gt_239_n120), .A2(u1_gt_239_n192), .A3(
        u1_gt_239_n121), .ZN(u1_gt_239_n403) );
  NAND4_X2 u1_gt_239_U491 ( .A1(u1_gt_239_n398), .A2(u1_gt_239_n399), .A3(
        u1_gt_239_n400), .A4(u1_gt_239_n401), .ZN(u1_gt_239_n386) );
  NOR2_X4 u1_gt_239_U490 ( .A1(u1_gt_239_n204), .A2(u1_gt_239_n28), .ZN(
        u1_gt_239_n388) );
  NAND2_X2 u1_gt_239_U489 ( .A1(u1_gt_239_n144), .A2(u1_gt_239_n145), .ZN(
        u1_gt_239_n396) );
  NOR3_X4 u1_gt_239_U488 ( .A1(u1_gt_239_n29), .A2(u1_gt_239_n3), .A3(
        u1_gt_239_n396), .ZN(u1_gt_239_n389) );
  NAND2_X2 u1_gt_239_U487 ( .A1(u1_gt_239_n393), .A2(u1_gt_239_n394), .ZN(
        u1_gt_239_n392) );
  NOR2_X4 u1_gt_239_U486 ( .A1(u1_gt_239_n391), .A2(u1_gt_239_n392), .ZN(
        u1_gt_239_n390) );
  NAND3_X2 u1_gt_239_U485 ( .A1(u1_gt_239_n388), .A2(u1_gt_239_n389), .A3(
        u1_gt_239_n390), .ZN(u1_gt_239_n387) );
  NAND2_X2 u1_gt_239_U484 ( .A1(u1_gt_239_n386), .A2(u1_gt_239_n387), .ZN(
        u1_gt_239_n385) );
  NAND2_X2 u1_gt_239_U483 ( .A1(u1_gt_239_n382), .A2(u1_gt_239_n383), .ZN(
        u1_gt_239_n381) );
  NAND2_X2 u1_gt_239_U482 ( .A1(u1_gt_239_n77), .A2(u1_gt_239_n78), .ZN(
        u1_gt_239_n378) );
  NAND2_X2 u1_gt_239_U481 ( .A1(u1_gt_239_n25), .A2(u1_gt_239_n145), .ZN(
        u1_gt_239_n376) );
  NAND2_X2 u1_gt_239_U480 ( .A1(u1_gt_239_n79), .A2(u1_gt_239_n15), .ZN(
        u1_gt_239_n373) );
  NOR2_X4 u1_gt_239_U479 ( .A1(u1_gt_239_n372), .A2(u1_gt_239_n373), .ZN(
        u1_gt_239_n370) );
  NAND4_X2 u1_gt_239_U478 ( .A1(u1_gt_239_n368), .A2(u1_gt_239_n369), .A3(
        u1_gt_239_n370), .A4(u1_gt_239_n371), .ZN(u1_gt_239_n367) );
  INV_X4 u1_gt_239_U477 ( .A(u1_gt_239_n367), .ZN(u1_gt_239_n352) );
  NAND4_X2 u1_gt_239_U476 ( .A1(u1_gt_239_n363), .A2(u1_gt_239_n364), .A3(
        u1_gt_239_n365), .A4(u1_gt_239_n366), .ZN(u1_gt_239_n354) );
  INV_X4 u1_gt_239_U475 ( .A(u1_gt_239_n361), .ZN(u1_gt_239_n359) );
  NAND2_X2 u1_gt_239_U474 ( .A1(u1_gt_239_n145), .A2(u1_gt_239_n26), .ZN(
        u1_gt_239_n360) );
  NOR2_X4 u1_gt_239_U473 ( .A1(u1_gt_239_n359), .A2(u1_gt_239_n360), .ZN(
        u1_gt_239_n358) );
  NAND2_X2 u1_gt_239_U472 ( .A1(u1_gt_239_n358), .A2(u1_gt_239_n223), .ZN(
        u1_gt_239_n355) );
  NOR3_X4 u1_gt_239_U471 ( .A1(u1_gt_239_n33), .A2(u1_gt_239_n204), .A3(
        u1_gt_239_n241), .ZN(u1_gt_239_n357) );
  NAND2_X2 u1_gt_239_U470 ( .A1(u1_gt_239_n222), .A2(u1_gt_239_n357), .ZN(
        u1_gt_239_n356) );
  NOR3_X4 u1_gt_239_U469 ( .A1(u1_gt_239_n354), .A2(u1_gt_239_n355), .A3(
        u1_gt_239_n356), .ZN(u1_gt_239_n353) );
  NAND2_X2 u1_gt_239_U468 ( .A1(u1_gt_239_n351), .A2(u1_gt_239_n223), .ZN(
        u1_gt_239_n346) );
  NOR2_X4 u1_gt_239_U467 ( .A1(u1_gt_239_n350), .A2(u1_gt_239_n31), .ZN(
        u1_gt_239_n348) );
  NOR3_X4 u1_gt_239_U466 ( .A1(u1_gt_239_n346), .A2(u1_gt_239_n347), .A3(
        u1_gt_239_n29), .ZN(u1_gt_239_n337) );
  NAND4_X2 u1_gt_239_U465 ( .A1(u1_gt_239_n344), .A2(u1_gt_239_n17), .A3(
        u1_gt_239_n18), .A4(u1_gt_239_n197), .ZN(u1_gt_239_n339) );
  INV_X4 u1_gt_239_U464 ( .A(n8448), .ZN(u1_gt_239_n343) );
  NAND4_X2 u1_gt_239_U463 ( .A1(u1_gt_239_n11), .A2(u1_gt_239_n342), .A3(
        u1_gt_239_n212), .A4(u1_gt_239_n343), .ZN(u1_gt_239_n340) );
  NAND3_X2 u1_gt_239_U462 ( .A1(u1_gt_239_n192), .A2(u1_gt_239_n194), .A3(
        u1_gt_239_n121), .ZN(u1_gt_239_n341) );
  NOR3_X4 u1_gt_239_U461 ( .A1(u1_gt_239_n339), .A2(u1_gt_239_n340), .A3(
        u1_gt_239_n341), .ZN(u1_gt_239_n338) );
  NAND3_X2 u1_gt_239_U460 ( .A1(u1_gt_239_n336), .A2(u1_gt_239_n337), .A3(
        u1_gt_239_n338), .ZN(u1_gt_239_n335) );
  NAND2_X2 u1_gt_239_U459 ( .A1(u1_gt_239_n334), .A2(u1_gt_239_n335), .ZN(
        u1_gt_239_n302) );
  NAND2_X2 u1_gt_239_U458 ( .A1(u1_gt_239_n332), .A2(u1_gt_239_n333), .ZN(
        u1_gt_239_n330) );
  NAND2_X2 u1_gt_239_U457 ( .A1(u1_gt_239_n222), .A2(n8400), .ZN(
        u1_gt_239_n331) );
  NOR3_X4 u1_gt_239_U456 ( .A1(u1_gt_239_n330), .A2(u1_gt_239_n331), .A3(
        u1_gt_239_n27), .ZN(u1_gt_239_n324) );
  NAND3_X2 u1_gt_239_U455 ( .A1(u1_gt_239_n324), .A2(u1_gt_239_n116), .A3(
        u1_gt_239_n325), .ZN(u1_gt_239_n323) );
  INV_X4 u1_gt_239_U454 ( .A(u1_gt_239_n323), .ZN(u1_gt_239_n303) );
  NAND3_X2 u1_gt_239_U453 ( .A1(u1_gt_239_n245), .A2(n8384), .A3(u1_gt_239_n26), .ZN(u1_gt_239_n322) );
  INV_X4 u1_gt_239_U452 ( .A(n8437), .ZN(u1_gt_239_n321) );
  NAND4_X2 u1_gt_239_U451 ( .A1(u1_gt_239_n13), .A2(u1_gt_239_n119), .A3(
        u1_gt_239_n17), .A4(u1_gt_239_n321), .ZN(u1_gt_239_n318) );
  NAND3_X2 u1_gt_239_U450 ( .A1(u1_gt_239_n320), .A2(u1_gt_239_n15), .A3(
        u1_gt_239_n79), .ZN(u1_gt_239_n319) );
  NOR2_X4 u1_gt_239_U449 ( .A1(u1_gt_239_n318), .A2(u1_gt_239_n319), .ZN(
        u1_gt_239_n317) );
  INV_X4 u1_gt_239_U448 ( .A(u1_gt_239_n70), .ZN(u1_gt_239_n307) );
  NAND2_X2 u1_gt_239_U447 ( .A1(n8375), .A2(u1_gt_239_n312), .ZN(
        u1_gt_239_n310) );
  NAND3_X2 u1_gt_239_U446 ( .A1(u1_gt_239_n309), .A2(u1_gt_239_n310), .A3(
        u1_gt_239_n311), .ZN(u1_gt_239_n308) );
  NAND2_X2 u1_gt_239_U445 ( .A1(u1_gt_239_n307), .A2(u1_gt_239_n308), .ZN(
        u1_gt_239_n306) );
  NAND2_X2 u1_gt_239_U444 ( .A1(u1_gt_239_n305), .A2(u1_gt_239_n306), .ZN(
        u1_gt_239_n304) );
  INV_X4 u1_gt_239_U443 ( .A(n8404), .ZN(u1_gt_239_n301) );
  NAND3_X2 u1_gt_239_U442 ( .A1(u1_gt_239_n13), .A2(u1_gt_239_n119), .A3(
        u1_gt_239_n15), .ZN(u1_gt_239_n300) );
  NAND2_X2 u1_gt_239_U441 ( .A1(u1_gt_239_n298), .A2(u1_gt_239_n299), .ZN(
        u1_gt_239_n280) );
  NOR2_X4 u1_gt_239_U440 ( .A1(u1_gt_239_n103), .A2(u1_gt_239_n104), .ZN(
        u1_gt_239_n297) );
  NAND2_X2 u1_gt_239_U439 ( .A1(u1_gt_239_n294), .A2(u1_gt_239_n295), .ZN(
        u1_gt_239_n293) );
  NOR2_X4 u1_gt_239_U438 ( .A1(u1_gt_239_n292), .A2(u1_gt_239_n293), .ZN(
        u1_gt_239_n291) );
  NAND2_X2 u1_gt_239_U437 ( .A1(u1_gt_239_n291), .A2(u1_gt_239_n116), .ZN(
        u1_gt_239_n281) );
  NOR2_X4 u1_gt_239_U436 ( .A1(u1_gt_239_n31), .A2(u1_gt_239_n290), .ZN(
        u1_gt_239_n289) );
  INV_X4 u1_gt_239_U435 ( .A(n8433), .ZN(u1_gt_239_n287) );
  NAND2_X2 u1_gt_239_U434 ( .A1(u1_gt_239_n78), .A2(u1_gt_239_n287), .ZN(
        u1_gt_239_n286) );
  NOR3_X4 u1_gt_239_U433 ( .A1(u1_gt_239_n285), .A2(u1_gt_239_n33), .A3(
        u1_gt_239_n286), .ZN(u1_gt_239_n284) );
  NAND2_X2 u1_gt_239_U432 ( .A1(u1_gt_239_n283), .A2(u1_gt_239_n284), .ZN(
        u1_gt_239_n282) );
  OAI21_X4 u1_gt_239_U431 ( .B1(u1_gt_239_n280), .B2(u1_gt_239_n281), .A(
        u1_gt_239_n282), .ZN(u1_gt_239_n255) );
  NAND3_X2 u1_gt_239_U430 ( .A1(u1_gt_239_n13), .A2(u1_gt_239_n18), .A3(
        u1_gt_239_n15), .ZN(u1_gt_239_n279) );
  NAND2_X2 u1_gt_239_U429 ( .A1(u1_gt_239_n278), .A2(u1_gt_239_n116), .ZN(
        u1_gt_239_n257) );
  INV_X4 u1_gt_239_U428 ( .A(n8461), .ZN(u1_gt_239_n275) );
  NAND3_X2 u1_gt_239_U427 ( .A1(u1_gt_239_n232), .A2(u1_gt_239_n275), .A3(
        u1_gt_239_n276), .ZN(u1_gt_239_n272) );
  NAND2_X2 u1_gt_239_U426 ( .A1(u1_gt_239_n213), .A2(u1_gt_239_n9), .ZN(
        u1_gt_239_n273) );
  NOR2_X4 u1_gt_239_U425 ( .A1(u1_gt_239_n272), .A2(u1_gt_239_n273), .ZN(
        u1_gt_239_n268) );
  NAND3_X2 u1_gt_239_U424 ( .A1(u1_gt_239_n121), .A2(u1_gt_239_n212), .A3(
        u1_gt_239_n11), .ZN(u1_gt_239_n270) );
  NAND2_X2 u1_gt_239_U423 ( .A1(u1_gt_239_n17), .A2(u1_gt_239_n120), .ZN(
        u1_gt_239_n271) );
  NOR2_X4 u1_gt_239_U422 ( .A1(u1_gt_239_n270), .A2(u1_gt_239_n271), .ZN(
        u1_gt_239_n269) );
  NAND3_X2 u1_gt_239_U421 ( .A1(u1_gt_239_n267), .A2(u1_gt_239_n268), .A3(
        u1_gt_239_n269), .ZN(u1_gt_239_n258) );
  INV_X4 u1_gt_239_U420 ( .A(n8424), .ZN(u1_gt_239_n266) );
  NAND2_X2 u1_gt_239_U419 ( .A1(n8371), .A2(u1_gt_239_n266), .ZN(
        u1_gt_239_n265) );
  NOR2_X4 u1_gt_239_U418 ( .A1(u1_gt_239_n31), .A2(u1_gt_239_n265), .ZN(
        u1_gt_239_n260) );
  INV_X4 u1_gt_239_U417 ( .A(n8423), .ZN(u1_gt_239_n264) );
  NAND2_X2 u1_gt_239_U416 ( .A1(n8370), .A2(u1_gt_239_n264), .ZN(
        u1_gt_239_n262) );
  INV_X4 u1_gt_239_U415 ( .A(n8422), .ZN(u1_gt_239_n61) );
  NAND2_X2 u1_gt_239_U414 ( .A1(n8369), .A2(u1_gt_239_n61), .ZN(u1_gt_239_n263) );
  NAND2_X2 u1_gt_239_U413 ( .A1(u1_gt_239_n262), .A2(u1_gt_239_n263), .ZN(
        u1_gt_239_n261) );
  OAI21_X4 u1_gt_239_U412 ( .B1(u1_gt_239_n257), .B2(u1_gt_239_n258), .A(
        u1_gt_239_n259), .ZN(u1_gt_239_n256) );
  NAND2_X2 u1_gt_239_U411 ( .A1(u1_gt_239_n253), .A2(u1_gt_239_n254), .ZN(
        u1_gt_239_n62) );
  NAND4_X2 u1_gt_239_U410 ( .A1(u1_gt_239_n250), .A2(u1_gt_239_n17), .A3(
        u1_gt_239_n251), .A4(u1_gt_239_n252), .ZN(u1_gt_239_n246) );
  NAND3_X2 u1_gt_239_U409 ( .A1(n8398), .A2(u1_gt_239_n222), .A3(
        u1_gt_239_n249), .ZN(u1_gt_239_n247) );
  NAND2_X2 u1_gt_239_U408 ( .A1(u1_gt_239_n223), .A2(u1_gt_239_n79), .ZN(
        u1_gt_239_n248) );
  NOR3_X4 u1_gt_239_U407 ( .A1(u1_gt_239_n246), .A2(u1_gt_239_n247), .A3(
        u1_gt_239_n248), .ZN(u1_gt_239_n236) );
  NAND3_X2 u1_gt_239_U406 ( .A1(u1_gt_239_n145), .A2(u1_gt_239_n26), .A3(
        u1_gt_239_n201), .ZN(u1_gt_239_n243) );
  NAND2_X2 u1_gt_239_U405 ( .A1(n8379), .A2(u1_gt_239_n245), .ZN(
        u1_gt_239_n244) );
  NOR2_X4 u1_gt_239_U404 ( .A1(u1_gt_239_n243), .A2(u1_gt_239_n244), .ZN(
        u1_gt_239_n242) );
  NAND2_X2 u1_gt_239_U403 ( .A1(u1_gt_239_n242), .A2(u1_gt_239_n223), .ZN(
        u1_gt_239_n238) );
  NAND2_X2 u1_gt_239_U402 ( .A1(u1_gt_239_n222), .A2(u1_gt_239_n240), .ZN(
        u1_gt_239_n239) );
  INV_X4 u1_gt_239_U401 ( .A(u1_gt_239_n235), .ZN(u1_gt_239_n234) );
  NAND2_X2 u1_gt_239_U400 ( .A1(u1_gt_239_n229), .A2(u1_gt_239_n230), .ZN(
        u1_gt_239_n228) );
  NOR2_X4 u1_gt_239_U399 ( .A1(u1_gt_239_n227), .A2(u1_gt_239_n228), .ZN(
        u1_gt_239_n226) );
  NAND2_X2 u1_gt_239_U398 ( .A1(u1_gt_239_n226), .A2(u1_gt_239_n116), .ZN(
        u1_gt_239_n219) );
  NAND3_X2 u1_gt_239_U397 ( .A1(u1_gt_239_n222), .A2(n8402), .A3(
        u1_gt_239_n223), .ZN(u1_gt_239_n221) );
  NOR3_X4 u1_gt_239_U396 ( .A1(u1_gt_239_n219), .A2(u1_gt_239_n220), .A3(
        u1_gt_239_n221), .ZN(u1_gt_239_n181) );
  NAND2_X2 u1_gt_239_U395 ( .A1(u1_gt_239_n15), .A2(u1_gt_239_n13), .ZN(
        u1_gt_239_n217) );
  INV_X4 u1_gt_239_U394 ( .A(n8454), .ZN(u1_gt_239_n214) );
  NAND2_X2 u1_gt_239_U393 ( .A1(u1_gt_239_n213), .A2(u1_gt_239_n214), .ZN(
        u1_gt_239_n209) );
  NAND2_X2 u1_gt_239_U392 ( .A1(u1_gt_239_n11), .A2(u1_gt_239_n212), .ZN(
        u1_gt_239_n210) );
  NOR3_X4 u1_gt_239_U391 ( .A1(u1_gt_239_n208), .A2(u1_gt_239_n209), .A3(
        u1_gt_239_n210), .ZN(u1_gt_239_n207) );
  NAND3_X2 u1_gt_239_U390 ( .A1(u1_gt_239_n205), .A2(u1_gt_239_n206), .A3(
        u1_gt_239_n207), .ZN(u1_gt_239_n184) );
  NOR2_X4 u1_gt_239_U389 ( .A1(u1_gt_239_n88), .A2(u1_gt_239_n86), .ZN(
        u1_gt_239_n200) );
  NAND2_X2 u1_gt_239_U388 ( .A1(u1_gt_239_n78), .A2(u1_gt_239_n15), .ZN(
        u1_gt_239_n199) );
  NOR3_X4 u1_gt_239_U387 ( .A1(u1_gt_239_n198), .A2(u1_gt_239_n33), .A3(
        u1_gt_239_n199), .ZN(u1_gt_239_n187) );
  NAND3_X2 u1_gt_239_U386 ( .A1(u1_gt_239_n197), .A2(u1_gt_239_n24), .A3(
        u1_gt_239_n17), .ZN(u1_gt_239_n195) );
  NAND2_X2 u1_gt_239_U385 ( .A1(u1_gt_239_n13), .A2(u1_gt_239_n18), .ZN(
        u1_gt_239_n196) );
  NOR2_X4 u1_gt_239_U384 ( .A1(u1_gt_239_n195), .A2(u1_gt_239_n196), .ZN(
        u1_gt_239_n188) );
  INV_X4 u1_gt_239_U383 ( .A(n8445), .ZN(u1_gt_239_n193) );
  NAND3_X2 u1_gt_239_U382 ( .A1(u1_gt_239_n192), .A2(u1_gt_239_n193), .A3(
        u1_gt_239_n194), .ZN(u1_gt_239_n190) );
  NAND3_X2 u1_gt_239_U381 ( .A1(u1_gt_239_n120), .A2(u1_gt_239_n165), .A3(
        u1_gt_239_n121), .ZN(u1_gt_239_n191) );
  NAND4_X2 u1_gt_239_U380 ( .A1(u1_gt_239_n186), .A2(u1_gt_239_n187), .A3(
        u1_gt_239_n188), .A4(u1_gt_239_n189), .ZN(u1_gt_239_n185) );
  OAI21_X4 u1_gt_239_U379 ( .B1(u1_gt_239_n183), .B2(u1_gt_239_n184), .A(
        u1_gt_239_n185), .ZN(u1_gt_239_n182) );
  NAND3_X2 u1_gt_239_U378 ( .A1(u1_gt_239_n18), .A2(u1_gt_239_n120), .A3(
        u1_gt_239_n17), .ZN(u1_gt_239_n179) );
  NAND3_X2 u1_gt_239_U377 ( .A1(u1_gt_239_n15), .A2(u1_gt_239_n13), .A3(
        u1_gt_239_n79), .ZN(u1_gt_239_n180) );
  NOR2_X4 u1_gt_239_U376 ( .A1(u1_gt_239_n179), .A2(u1_gt_239_n180), .ZN(
        u1_gt_239_n178) );
  NAND2_X2 u1_gt_239_U375 ( .A1(u1_gt_239_n178), .A2(u1_gt_239_n116), .ZN(
        u1_gt_239_n166) );
  NAND2_X2 u1_gt_239_U374 ( .A1(u1_gt_239_n175), .A2(u1_gt_239_n176), .ZN(
        u1_gt_239_n171) );
  NOR3_X4 u1_gt_239_U373 ( .A1(u1_gt_239_n10), .A2(u1_gt_239_n104), .A3(
        u1_gt_239_n20), .ZN(u1_gt_239_n173) );
  NOR3_X4 u1_gt_239_U372 ( .A1(u1_gt_239_n8), .A2(u1_gt_239_n102), .A3(
        u1_gt_239_n103), .ZN(u1_gt_239_n174) );
  NAND2_X2 u1_gt_239_U371 ( .A1(u1_gt_239_n173), .A2(u1_gt_239_n174), .ZN(
        u1_gt_239_n172) );
  NOR2_X4 u1_gt_239_U370 ( .A1(u1_gt_239_n171), .A2(u1_gt_239_n172), .ZN(
        u1_gt_239_n170) );
  NAND3_X2 u1_gt_239_U369 ( .A1(u1_gt_239_n168), .A2(u1_gt_239_n169), .A3(
        u1_gt_239_n170), .ZN(u1_gt_239_n167) );
  NOR2_X4 u1_gt_239_U368 ( .A1(u1_gt_239_n166), .A2(u1_gt_239_n167), .ZN(
        u1_gt_239_n123) );
  NAND3_X2 u1_gt_239_U367 ( .A1(u1_gt_239_n165), .A2(u1_gt_239_n120), .A3(
        u1_gt_239_n24), .ZN(u1_gt_239_n164) );
  NAND4_X2 u1_gt_239_U366 ( .A1(u1_gt_239_n156), .A2(u1_gt_239_n157), .A3(
        u1_gt_239_n158), .A4(u1_gt_239_n159), .ZN(u1_gt_239_n125) );
  NOR2_X4 u1_gt_239_U365 ( .A1(u1_gt_239_n155), .A2(u1_gt_239_n31), .ZN(
        u1_gt_239_n153) );
  NOR2_X4 u1_gt_239_U364 ( .A1(u1_gt_239_n152), .A2(u1_gt_239_n29), .ZN(
        u1_gt_239_n148) );
  NAND2_X2 u1_gt_239_U363 ( .A1(u1_gt_239_n77), .A2(u1_gt_239_n78), .ZN(
        u1_gt_239_n151) );
  NAND2_X2 u1_gt_239_U362 ( .A1(u1_gt_239_n77), .A2(u1_gt_239_n78), .ZN(
        u1_gt_239_n147) );
  NAND2_X2 u1_gt_239_U361 ( .A1(u1_gt_239_n26), .A2(u1_gt_239_n145), .ZN(
        u1_gt_239_n143) );
  NOR3_X4 u1_gt_239_U360 ( .A1(u1_gt_239_n29), .A2(u1_gt_239_n5), .A3(
        u1_gt_239_n143), .ZN(u1_gt_239_n129) );
  NOR2_X4 u1_gt_239_U359 ( .A1(u1_gt_239_n137), .A2(u1_gt_239_n34), .ZN(
        u1_gt_239_n133) );
  NAND2_X2 u1_gt_239_U358 ( .A1(u1_gt_239_n133), .A2(u1_gt_239_n134), .ZN(
        u1_gt_239_n132) );
  NOR2_X4 u1_gt_239_U357 ( .A1(u1_gt_239_n131), .A2(u1_gt_239_n132), .ZN(
        u1_gt_239_n130) );
  NAND3_X2 u1_gt_239_U356 ( .A1(u1_gt_239_n128), .A2(u1_gt_239_n129), .A3(
        u1_gt_239_n130), .ZN(u1_gt_239_n127) );
  OAI21_X4 u1_gt_239_U355 ( .B1(u1_gt_239_n125), .B2(u1_gt_239_n126), .A(
        u1_gt_239_n127), .ZN(u1_gt_239_n124) );
  NAND3_X2 u1_gt_239_U354 ( .A1(u1_gt_239_n120), .A2(u1_gt_239_n121), .A3(
        u1_gt_239_n17), .ZN(u1_gt_239_n117) );
  NAND3_X2 u1_gt_239_U353 ( .A1(u1_gt_239_n13), .A2(u1_gt_239_n119), .A3(
        u1_gt_239_n15), .ZN(u1_gt_239_n118) );
  NOR2_X4 u1_gt_239_U352 ( .A1(u1_gt_239_n117), .A2(u1_gt_239_n118), .ZN(
        u1_gt_239_n115) );
  NAND2_X2 u1_gt_239_U351 ( .A1(u1_gt_239_n115), .A2(u1_gt_239_n116), .ZN(
        u1_gt_239_n92) );
  NOR3_X4 u1_gt_239_U350 ( .A1(u1_gt_239_n109), .A2(u1_gt_239_n110), .A3(
        u1_gt_239_n111), .ZN(u1_gt_239_n105) );
  NOR3_X4 u1_gt_239_U349 ( .A1(u1_gt_239_n107), .A2(n8411), .A3(u1_gt_239_n108), .ZN(u1_gt_239_n106) );
  NAND2_X2 u1_gt_239_U348 ( .A1(u1_gt_239_n105), .A2(u1_gt_239_n106), .ZN(
        u1_gt_239_n97) );
  NOR3_X4 u1_gt_239_U347 ( .A1(u1_gt_239_n10), .A2(u1_gt_239_n103), .A3(
        u1_gt_239_n104), .ZN(u1_gt_239_n99) );
  NOR3_X4 u1_gt_239_U346 ( .A1(u1_gt_239_n8), .A2(u1_gt_239_n101), .A3(
        u1_gt_239_n102), .ZN(u1_gt_239_n100) );
  NAND2_X2 u1_gt_239_U345 ( .A1(u1_gt_239_n99), .A2(u1_gt_239_n100), .ZN(
        u1_gt_239_n98) );
  NOR2_X4 u1_gt_239_U344 ( .A1(u1_gt_239_n97), .A2(u1_gt_239_n98), .ZN(
        u1_gt_239_n96) );
  NAND3_X2 u1_gt_239_U343 ( .A1(u1_gt_239_n94), .A2(u1_gt_239_n95), .A3(
        u1_gt_239_n96), .ZN(u1_gt_239_n93) );
  NOR2_X4 u1_gt_239_U342 ( .A1(u1_gt_239_n92), .A2(u1_gt_239_n93), .ZN(
        u1_gt_239_n68) );
  NAND2_X2 u1_gt_239_U341 ( .A1(u1_gt_239_n77), .A2(u1_gt_239_n90), .ZN(
        u1_gt_239_n71) );
  NOR2_X4 u1_gt_239_U340 ( .A1(u1_gt_239_n88), .A2(u1_gt_239_n31), .ZN(
        u1_gt_239_n84) );
  NOR2_X4 u1_gt_239_U339 ( .A1(u1_gt_239_n86), .A2(u1_gt_239_n87), .ZN(
        u1_gt_239_n85) );
  NAND3_X4 u1_gt_239_U338 ( .A1(u1_gt_239_n84), .A2(n8382), .A3(u1_gt_239_n85), 
        .ZN(u1_gt_239_n83) );
  NOR2_X4 u1_gt_239_U337 ( .A1(u1_gt_239_n83), .A2(u1_gt_239_n29), .ZN(
        u1_gt_239_n73) );
  INV_X4 u1_gt_239_U336 ( .A(n8435), .ZN(u1_gt_239_n82) );
  NAND4_X2 u1_gt_239_U335 ( .A1(u1_gt_239_n79), .A2(u1_gt_239_n15), .A3(
        u1_gt_239_n13), .A4(u1_gt_239_n82), .ZN(u1_gt_239_n75) );
  NAND2_X2 u1_gt_239_U334 ( .A1(u1_gt_239_n77), .A2(u1_gt_239_n78), .ZN(
        u1_gt_239_n76) );
  NOR3_X4 u1_gt_239_U333 ( .A1(u1_gt_239_n75), .A2(u1_gt_239_n27), .A3(
        u1_gt_239_n76), .ZN(u1_gt_239_n74) );
  NAND2_X2 u1_gt_239_U332 ( .A1(u1_gt_239_n73), .A2(u1_gt_239_n74), .ZN(
        u1_gt_239_n72) );
  NAND4_X2 u1_gt_239_U331 ( .A1(u1_gt_239_n64), .A2(u1_gt_239_n65), .A3(
        u1_gt_239_n66), .A4(u1_gt_239_n67), .ZN(u1_gt_239_n63) );
  NAND2_X2 u1_gt_239_U330 ( .A1(u1_gt_239_n60), .A2(u1_gt_239_n58), .ZN(
        u1_gt_239_n39) );
  NAND2_X2 u1_gt_239_U329 ( .A1(u1_gt_239_n57), .A2(u1_gt_239_n58), .ZN(
        u1_gt_239_n40) );
  XNOR2_X2 u1_gt_239_U328 ( .A(n8361), .B(n8414), .ZN(u1_gt_239_n54) );
  INV_X4 u1_gt_239_U327 ( .A(n8362), .ZN(u1_gt_239_n56) );
  NAND2_X2 u1_gt_239_U326 ( .A1(n8415), .A2(u1_gt_239_n56), .ZN(u1_gt_239_n55)
         );
  OAI22_X2 u1_gt_239_U325 ( .A1(u1_gt_239_n2), .A2(u1_gt_239_n54), .B1(
        u1_gt_239_n2), .B2(u1_gt_239_n55), .ZN(u1_gt_239_n49) );
  NAND2_X2 u1_gt_239_U324 ( .A1(n8419), .A2(u1_gt_239_n585), .ZN(u1_gt_239_n48) );
  INV_X4 u1_gt_239_U323 ( .A(n8365), .ZN(u1_gt_239_n47) );
  NAND2_X2 u1_gt_239_U322 ( .A1(n8418), .A2(u1_gt_239_n47), .ZN(u1_gt_239_n46)
         );
  NAND4_X2 u1_gt_239_U321 ( .A1(u1_gt_239_n39), .A2(u1_gt_239_n40), .A3(
        u1_gt_239_n41), .A4(u1_gt_239_n42), .ZN(u1_gt_239_n38) );
  AOI21_X4 u1_gt_239_U320 ( .B1(u1_gt_239_n36), .B2(u1_gt_239_n37), .A(
        u1_gt_239_n38), .ZN(u1_fractb_lt_fracta) );
  INV_X32 u1_gt_239_U319 ( .A(u1_gt_239_n32), .ZN(u1_gt_239_n31) );
  INV_X32 u1_gt_239_U318 ( .A(u1_gt_239_n222), .ZN(u1_gt_239_n29) );
  NAND2_X4 u1_gt_239_U317 ( .A1(n8425), .A2(u1_gt_239_n504), .ZN(
        u1_gt_239_n145) );
  INV_X16 u1_gt_239_U316 ( .A(u1_gt_239_n145), .ZN(u1_gt_239_n86) );
  NAND2_X4 u1_gt_239_U315 ( .A1(n8424), .A2(u1_gt_239_n851), .ZN(
        u1_gt_239_n144) );
  NAND2_X4 u1_gt_239_U314 ( .A1(n8424), .A2(u1_gt_239_n851), .ZN(u1_gt_239_n26) );
  NAND2_X4 u1_gt_239_U313 ( .A1(n8424), .A2(u1_gt_239_n851), .ZN(u1_gt_239_n25) );
  NAND3_X4 u1_gt_239_U312 ( .A1(u1_gt_239_n309), .A2(u1_gt_239_n846), .A3(
        n8427), .ZN(u1_gt_239_n222) );
  NAND2_X4 u1_gt_239_U311 ( .A1(n8426), .A2(u1_gt_239_n845), .ZN(
        u1_gt_239_n201) );
  NAND3_X4 u1_gt_239_U310 ( .A1(u1_gt_239_n843), .A2(u1_gt_239_n309), .A3(
        u1_gt_239_n311), .ZN(u1_gt_239_n223) );
  NAND2_X4 u1_gt_239_U309 ( .A1(n8430), .A2(u1_gt_239_n91), .ZN(u1_gt_239_n78)
         );
  NAND2_X4 u1_gt_239_U308 ( .A1(n8429), .A2(u1_gt_239_n533), .ZN(u1_gt_239_n77) );
  NAND2_X4 u1_gt_239_U307 ( .A1(n8432), .A2(u1_gt_239_n842), .ZN(u1_gt_239_n79) );
  NAND2_X4 u1_gt_239_U306 ( .A1(n8438), .A2(u1_gt_239_n397), .ZN(
        u1_gt_239_n139) );
  INV_X32 u1_gt_239_U305 ( .A(u1_gt_239_n23), .ZN(u1_gt_239_n24) );
  INV_X8 u1_gt_239_U304 ( .A(u1_gt_239_n120), .ZN(u1_gt_239_n216) );
  INV_X32 u1_gt_239_U303 ( .A(u1_gt_239_n21), .ZN(u1_gt_239_n22) );
  INV_X8 u1_gt_239_U302 ( .A(u1_gt_239_n121), .ZN(u1_gt_239_n161) );
  INV_X32 u1_gt_239_U301 ( .A(u1_gt_239_n19), .ZN(u1_gt_239_n20) );
  NAND2_X4 u1_gt_239_U300 ( .A1(n8435), .A2(u1_gt_239_n837), .ZN(
        u1_gt_239_n119) );
  NAND2_X4 u1_gt_239_U299 ( .A1(n8435), .A2(u1_gt_239_n837), .ZN(u1_gt_239_n18) );
  NAND2_X4 u1_gt_239_U298 ( .A1(n8436), .A2(u1_gt_239_n499), .ZN(
        u1_gt_239_n122) );
  INV_X32 u1_gt_239_U297 ( .A(u1_gt_239_n14), .ZN(u1_gt_239_n15) );
  NAND2_X4 u1_gt_239_U296 ( .A1(n8434), .A2(u1_gt_239_n835), .ZN(u1_gt_239_n81) );
  INV_X32 u1_gt_239_U295 ( .A(u1_gt_239_n12), .ZN(u1_gt_239_n13) );
  NAND2_X4 u1_gt_239_U294 ( .A1(n8448), .A2(u1_gt_239_n350), .ZN(
        u1_gt_239_n213) );
  NAND2_X4 u1_gt_239_U293 ( .A1(n8447), .A2(u1_gt_239_n155), .ZN(
        u1_gt_239_n212) );
  NAND2_X4 u1_gt_239_U292 ( .A1(n8445), .A2(u1_gt_239_n203), .ZN(
        u1_gt_239_n211) );
  NAND2_X4 u1_gt_239_U291 ( .A1(n8455), .A2(u1_gt_239_n827), .ZN(
        u1_gt_239_n232) );
  NAND2_X4 u1_gt_239_U290 ( .A1(n8454), .A2(u1_gt_239_n218), .ZN(
        u1_gt_239_n274) );
  INV_X16 u1_gt_239_U289 ( .A(u1_gt_239_n78), .ZN(u1_gt_239_n241) );
  INV_X16 u1_gt_239_U288 ( .A(u1_gt_239_n77), .ZN(u1_gt_239_n204) );
  INV_X16 u1_gt_239_U287 ( .A(u1_gt_239_n197), .ZN(u1_gt_239_n141) );
  INV_X32 u1_gt_239_U286 ( .A(u1_gt_239_n15), .ZN(u1_gt_239_n137) );
  INV_X16 u1_gt_239_U285 ( .A(u1_gt_239_n212), .ZN(u1_gt_239_n104) );
  INV_X16 u1_gt_239_U284 ( .A(u1_gt_239_n213), .ZN(u1_gt_239_n103) );
  INV_X16 u1_gt_239_U283 ( .A(u1_gt_239_n183), .ZN(u1_gt_239_n116) );
  INV_X32 u1_gt_239_U282 ( .A(u1_gt_239_n13), .ZN(u1_gt_239_n136) );
  INV_X16 u1_gt_239_U281 ( .A(u1_gt_239_n119), .ZN(u1_gt_239_n135) );
  INV_X16 u1_gt_239_U280 ( .A(u1_gt_239_n144), .ZN(u1_gt_239_n88) );
  INV_X4 u1_gt_239_U279 ( .A(n8414), .ZN(u1_gt_239_n600) );
  INV_X4 u1_gt_239_U278 ( .A(u1_gt_239_n814), .ZN(u1_gt_239_n812) );
  INV_X16 u1_gt_239_U277 ( .A(u1_gt_239_n223), .ZN(u1_gt_239_n28) );
  INV_X16 u1_gt_239_U276 ( .A(u1_gt_239_n35), .ZN(u1_gt_239_n33) );
  OR3_X2 u1_gt_239_U275 ( .A1(u1_gt_239_n87), .A2(u1_gt_239_n31), .A3(
        u1_gt_239_n517), .ZN(u1_gt_239_n7) );
  OR3_X2 u1_gt_239_U274 ( .A1(u1_gt_239_n87), .A2(u1_gt_239_n30), .A3(
        u1_gt_239_n377), .ZN(u1_gt_239_n6) );
  OR3_X4 u1_gt_239_U273 ( .A1(u1_gt_239_n87), .A2(u1_gt_239_n30), .A3(
        u1_gt_239_n146), .ZN(u1_gt_239_n5) );
  OR3_X2 u1_gt_239_U272 ( .A1(u1_gt_239_n87), .A2(u1_gt_239_n30), .A3(
        u1_gt_239_n533), .ZN(u1_gt_239_n4) );
  OR3_X2 u1_gt_239_U271 ( .A1(u1_gt_239_n87), .A2(u1_gt_239_n30), .A3(
        u1_gt_239_n397), .ZN(u1_gt_239_n3) );
  INV_X16 u1_gt_239_U270 ( .A(u1_gt_239_n211), .ZN(u1_gt_239_n10) );
  INV_X16 u1_gt_239_U269 ( .A(u1_gt_239_n10), .ZN(u1_gt_239_n11) );
  AND2_X4 u1_gt_239_U268 ( .A1(u1_gt_239_n600), .A2(n8361), .ZN(u1_gt_239_n2)
         );
  INV_X16 u1_gt_239_U267 ( .A(u1_gt_239_n122), .ZN(u1_gt_239_n16) );
  INV_X16 u1_gt_239_U266 ( .A(u1_gt_239_n16), .ZN(u1_gt_239_n17) );
  INV_X8 u1_gt_239_U265 ( .A(u1_gt_239_n274), .ZN(u1_gt_239_n8) );
  INV_X16 u1_gt_239_U264 ( .A(u1_gt_239_n8), .ZN(u1_gt_239_n9) );
  NOR3_X2 u1_gt_239_U263 ( .A1(u1_gt_239_n379), .A2(u1_gt_239_n380), .A3(
        u1_gt_239_n381), .ZN(u1_gt_239_n36) );
  NOR3_X2 u1_gt_239_U262 ( .A1(u1_gt_239_n326), .A2(u1_gt_239_n22), .A3(
        u1_gt_239_n16), .ZN(u1_gt_239_n325) );
  NOR2_X2 u1_gt_239_U261 ( .A1(u1_gt_239_n322), .A2(u1_gt_239_n28), .ZN(
        u1_gt_239_n316) );
  NOR3_X1 u1_gt_239_U260 ( .A1(u1_gt_239_n29), .A2(u1_gt_239_n87), .A3(
        u1_gt_239_n86), .ZN(u1_gt_239_n315) );
  NAND3_X2 u1_gt_239_U259 ( .A1(u1_gt_239_n315), .A2(u1_gt_239_n316), .A3(
        u1_gt_239_n317), .ZN(u1_gt_239_n305) );
  NOR3_X2 u1_gt_239_U258 ( .A1(u1_gt_239_n33), .A2(u1_gt_239_n136), .A3(
        u1_gt_239_n137), .ZN(u1_gt_239_n336) );
  NOR2_X2 u1_gt_239_U257 ( .A1(u1_gt_239_n352), .A2(u1_gt_239_n353), .ZN(
        u1_gt_239_n334) );
  NOR2_X2 u1_gt_239_U256 ( .A1(u1_gt_239_n136), .A2(u1_gt_239_n137), .ZN(
        u1_gt_239_n249) );
  NOR2_X2 u1_gt_239_U255 ( .A1(n8452), .A2(u1_gt_239_n103), .ZN(u1_gt_239_n252) );
  NOR3_X2 u1_gt_239_U254 ( .A1(u1_gt_239_n135), .A2(u1_gt_239_n20), .A3(
        u1_gt_239_n22), .ZN(u1_gt_239_n250) );
  NOR2_X2 u1_gt_239_U253 ( .A1(u1_gt_239_n104), .A2(u1_gt_239_n10), .ZN(
        u1_gt_239_n251) );
  NOR3_X1 u1_gt_239_U252 ( .A1(u1_gt_239_n204), .A2(n8432), .A3(u1_gt_239_n241), .ZN(u1_gt_239_n240) );
  NOR3_X2 u1_gt_239_U251 ( .A1(u1_gt_239_n217), .A2(u1_gt_239_n29), .A3(
        u1_gt_239_n218), .ZN(u1_gt_239_n206) );
  NOR2_X2 u1_gt_239_U250 ( .A1(u1_gt_239_n34), .A2(u1_gt_239_n28), .ZN(
        u1_gt_239_n205) );
  NOR2_X2 u1_gt_239_U249 ( .A1(u1_gt_239_n137), .A2(u1_gt_239_n34), .ZN(
        u1_gt_239_n225) );
  NOR2_X2 u1_gt_239_U248 ( .A1(u1_gt_239_n136), .A2(u1_gt_239_n135), .ZN(
        u1_gt_239_n224) );
  NAND3_X1 u1_gt_239_U247 ( .A1(u1_gt_239_n224), .A2(u1_gt_239_n17), .A3(
        u1_gt_239_n225), .ZN(u1_gt_239_n220) );
  NAND3_X1 u1_gt_239_U246 ( .A1(u1_gt_239_n231), .A2(u1_gt_239_n232), .A3(
        u1_gt_239_n233), .ZN(u1_gt_239_n227) );
  NOR2_X2 u1_gt_239_U245 ( .A1(u1_gt_239_n190), .A2(u1_gt_239_n191), .ZN(
        u1_gt_239_n189) );
  NOR3_X2 u1_gt_239_U244 ( .A1(u1_gt_239_n27), .A2(u1_gt_239_n204), .A3(
        u1_gt_239_n29), .ZN(u1_gt_239_n186) );
  NOR2_X2 u1_gt_239_U243 ( .A1(u1_gt_239_n31), .A2(u1_gt_239_n203), .ZN(
        u1_gt_239_n202) );
  NAND3_X1 u1_gt_239_U242 ( .A1(u1_gt_239_n200), .A2(u1_gt_239_n201), .A3(
        u1_gt_239_n202), .ZN(u1_gt_239_n198) );
  NOR3_X2 u1_gt_239_U241 ( .A1(u1_gt_239_n34), .A2(u1_gt_239_n136), .A3(
        u1_gt_239_n137), .ZN(u1_gt_239_n150) );
  NOR2_X2 u1_gt_239_U240 ( .A1(u1_gt_239_n28), .A2(u1_gt_239_n151), .ZN(
        u1_gt_239_n149) );
  NAND3_X2 u1_gt_239_U239 ( .A1(u1_gt_239_n148), .A2(u1_gt_239_n149), .A3(
        u1_gt_239_n150), .ZN(u1_gt_239_n126) );
  NOR2_X2 u1_gt_239_U238 ( .A1(u1_gt_239_n28), .A2(u1_gt_239_n147), .ZN(
        u1_gt_239_n128) );
  NOR2_X1 u1_gt_239_U237 ( .A1(u1_gt_239_n113), .A2(u1_gt_239_n177), .ZN(
        u1_gt_239_n169) );
  NOR2_X2 u1_gt_239_U236 ( .A1(u1_gt_239_n28), .A2(u1_gt_239_n29), .ZN(
        u1_gt_239_n168) );
  NOR2_X2 u1_gt_239_U235 ( .A1(u1_gt_239_n16), .A2(u1_gt_239_n164), .ZN(
        u1_gt_239_n156) );
  NOR2_X1 u1_gt_239_U234 ( .A1(u1_gt_239_n141), .A2(u1_gt_239_n135), .ZN(
        u1_gt_239_n157) );
  NOR3_X1 u1_gt_239_U233 ( .A1(u1_gt_239_n10), .A2(n8447), .A3(u1_gt_239_n160), 
        .ZN(u1_gt_239_n159) );
  NOR3_X1 u1_gt_239_U232 ( .A1(u1_gt_239_n20), .A2(u1_gt_239_n162), .A3(
        u1_gt_239_n163), .ZN(u1_gt_239_n158) );
  NOR2_X2 u1_gt_239_U231 ( .A1(u1_gt_239_n87), .A2(u1_gt_239_n29), .ZN(
        u1_gt_239_n314) );
  NOR3_X1 u1_gt_239_U230 ( .A1(u1_gt_239_n88), .A2(u1_gt_239_n86), .A3(
        u1_gt_239_n30), .ZN(u1_gt_239_n313) );
  NAND3_X2 u1_gt_239_U229 ( .A1(u1_gt_239_n313), .A2(u1_gt_239_n223), .A3(
        u1_gt_239_n314), .ZN(u1_gt_239_n70) );
  NOR3_X2 u1_gt_239_U228 ( .A1(u1_gt_239_n28), .A2(u1_gt_239_n33), .A3(
        u1_gt_239_n29), .ZN(u1_gt_239_n95) );
  NOR2_X1 u1_gt_239_U227 ( .A1(u1_gt_239_n113), .A2(u1_gt_239_n114), .ZN(
        u1_gt_239_n94) );
  NOR2_X2 u1_gt_239_U226 ( .A1(n8430), .A2(u1_gt_239_n91), .ZN(u1_gt_239_n90)
         );
  NOR3_X1 u1_gt_239_U225 ( .A1(u1_gt_239_n113), .A2(u1_gt_239_n29), .A3(
        u1_gt_239_n277), .ZN(u1_gt_239_n267) );
  NOR3_X2 u1_gt_239_U224 ( .A1(u1_gt_239_n279), .A2(u1_gt_239_n33), .A3(
        u1_gt_239_n27), .ZN(u1_gt_239_n278) );
  NOR3_X1 u1_gt_239_U223 ( .A1(u1_gt_239_n28), .A2(u1_gt_239_n204), .A3(
        u1_gt_239_n29), .ZN(u1_gt_239_n283) );
  NAND3_X1 u1_gt_239_U222 ( .A1(u1_gt_239_n288), .A2(u1_gt_239_n201), .A3(
        u1_gt_239_n289), .ZN(u1_gt_239_n285) );
  NOR3_X2 u1_gt_239_U221 ( .A1(u1_gt_239_n300), .A2(u1_gt_239_n33), .A3(
        u1_gt_239_n27), .ZN(u1_gt_239_n299) );
  NOR3_X1 u1_gt_239_U220 ( .A1(u1_gt_239_n113), .A2(u1_gt_239_n29), .A3(
        u1_gt_239_n301), .ZN(u1_gt_239_n298) );
  NOR2_X2 u1_gt_239_U219 ( .A1(u1_gt_239_n22), .A2(u1_gt_239_n16), .ZN(
        u1_gt_239_n294) );
  NAND3_X2 u1_gt_239_U218 ( .A1(u1_gt_239_n296), .A2(u1_gt_239_n9), .A3(
        u1_gt_239_n297), .ZN(u1_gt_239_n292) );
  NOR3_X2 u1_gt_239_U217 ( .A1(u1_gt_239_n499), .A2(u1_gt_239_n88), .A3(
        u1_gt_239_n30), .ZN(u1_gt_239_n498) );
  NOR2_X1 u1_gt_239_U216 ( .A1(u1_gt_239_n87), .A2(u1_gt_239_n86), .ZN(
        u1_gt_239_n497) );
  NOR2_X2 u1_gt_239_U215 ( .A1(u1_gt_239_n136), .A2(u1_gt_239_n137), .ZN(
        u1_gt_239_n500) );
  NOR2_X2 u1_gt_239_U214 ( .A1(n8436), .A2(u1_gt_239_n135), .ZN(u1_gt_239_n501) );
  NOR3_X1 u1_gt_239_U213 ( .A1(u1_gt_239_n33), .A2(u1_gt_239_n204), .A3(
        u1_gt_239_n241), .ZN(u1_gt_239_n502) );
  NOR2_X1 u1_gt_239_U212 ( .A1(u1_gt_239_n16), .A2(u1_gt_239_n135), .ZN(
        u1_gt_239_n515) );
  NAND3_X1 u1_gt_239_U211 ( .A1(u1_gt_239_n514), .A2(u1_gt_239_n24), .A3(
        u1_gt_239_n515), .ZN(u1_gt_239_n510) );
  NOR3_X2 u1_gt_239_U210 ( .A1(u1_gt_239_n524), .A2(u1_gt_239_n27), .A3(
        u1_gt_239_n525), .ZN(u1_gt_239_n523) );
  NOR2_X2 u1_gt_239_U209 ( .A1(n8429), .A2(u1_gt_239_n28), .ZN(u1_gt_239_n530)
         );
  NOR3_X2 u1_gt_239_U208 ( .A1(u1_gt_239_n29), .A2(u1_gt_239_n4), .A3(
        u1_gt_239_n532), .ZN(u1_gt_239_n531) );
  NOR2_X1 u1_gt_239_U207 ( .A1(u1_gt_239_n86), .A2(u1_gt_239_n87), .ZN(
        u1_gt_239_n529) );
  NOR2_X2 u1_gt_239_U206 ( .A1(u1_gt_239_n88), .A2(u1_gt_239_n31), .ZN(
        u1_gt_239_n528) );
  NAND3_X2 u1_gt_239_U205 ( .A1(u1_gt_239_n528), .A2(n8381), .A3(
        u1_gt_239_n529), .ZN(u1_gt_239_n527) );
  NOR3_X2 u1_gt_239_U204 ( .A1(u1_gt_239_n539), .A2(u1_gt_239_n22), .A3(
        u1_gt_239_n16), .ZN(u1_gt_239_n538) );
  NOR3_X1 u1_gt_239_U203 ( .A1(u1_gt_239_n113), .A2(u1_gt_239_n29), .A3(
        u1_gt_239_n543), .ZN(u1_gt_239_n536) );
  NOR3_X2 u1_gt_239_U202 ( .A1(u1_gt_239_n87), .A2(u1_gt_239_n30), .A3(
        u1_gt_239_n438), .ZN(u1_gt_239_n437) );
  NOR2_X2 u1_gt_239_U201 ( .A1(u1_gt_239_n142), .A2(u1_gt_239_n345), .ZN(
        u1_gt_239_n439) );
  NOR3_X2 u1_gt_239_U200 ( .A1(u1_gt_239_n20), .A2(n8443), .A3(u1_gt_239_n22), 
        .ZN(u1_gt_239_n440) );
  NOR3_X1 u1_gt_239_U199 ( .A1(u1_gt_239_n16), .A2(u1_gt_239_n141), .A3(
        u1_gt_239_n135), .ZN(u1_gt_239_n442) );
  NOR3_X1 u1_gt_239_U198 ( .A1(u1_gt_239_n33), .A2(u1_gt_239_n204), .A3(
        u1_gt_239_n241), .ZN(u1_gt_239_n433) );
  NOR3_X2 u1_gt_239_U197 ( .A1(u1_gt_239_n468), .A2(u1_gt_239_n20), .A3(
        u1_gt_239_n22), .ZN(u1_gt_239_n466) );
  NOR3_X1 u1_gt_239_U196 ( .A1(u1_gt_239_n104), .A2(u1_gt_239_n452), .A3(
        u1_gt_239_n103), .ZN(u1_gt_239_n467) );
  NOR2_X2 u1_gt_239_U195 ( .A1(u1_gt_239_n204), .A2(u1_gt_239_n29), .ZN(
        u1_gt_239_n477) );
  NOR2_X2 u1_gt_239_U194 ( .A1(u1_gt_239_n113), .A2(u1_gt_239_n487), .ZN(
        u1_gt_239_n479) );
  NOR2_X2 u1_gt_239_U193 ( .A1(u1_gt_239_n16), .A2(u1_gt_239_n135), .ZN(
        u1_gt_239_n486) );
  NAND3_X1 u1_gt_239_U192 ( .A1(u1_gt_239_n485), .A2(u1_gt_239_n24), .A3(
        u1_gt_239_n486), .ZN(u1_gt_239_n481) );
  NOR2_X2 u1_gt_239_U191 ( .A1(u1_gt_239_n8), .A2(u1_gt_239_n474), .ZN(
        u1_gt_239_n470) );
  NOR2_X2 u1_gt_239_U190 ( .A1(u1_gt_239_n475), .A2(u1_gt_239_n476), .ZN(
        u1_gt_239_n469) );
  NOR3_X1 u1_gt_239_U189 ( .A1(u1_gt_239_n109), .A2(u1_gt_239_n101), .A3(
        u1_gt_239_n102), .ZN(u1_gt_239_n472) );
  NOR2_X2 u1_gt_239_U188 ( .A1(n8463), .A2(u1_gt_239_n111), .ZN(u1_gt_239_n471) );
  NOR2_X2 u1_gt_239_U187 ( .A1(u1_gt_239_n88), .A2(u1_gt_239_n86), .ZN(
        u1_gt_239_n409) );
  NOR2_X2 u1_gt_239_U186 ( .A1(u1_gt_239_n136), .A2(u1_gt_239_n137), .ZN(
        u1_gt_239_n394) );
  NAND3_X2 u1_gt_239_U185 ( .A1(u1_gt_239_n18), .A2(u1_gt_239_n395), .A3(
        u1_gt_239_n17), .ZN(u1_gt_239_n391) );
  NOR2_X2 u1_gt_239_U184 ( .A1(u1_gt_239_n28), .A2(u1_gt_239_n29), .ZN(
        u1_gt_239_n414) );
  NAND3_X1 u1_gt_239_U183 ( .A1(u1_gt_239_n420), .A2(u1_gt_239_n421), .A3(
        u1_gt_239_n422), .ZN(u1_gt_239_n417) );
  NOR2_X1 u1_gt_239_U182 ( .A1(u1_gt_239_n86), .A2(u1_gt_239_n87), .ZN(
        u1_gt_239_n460) );
  NAND3_X2 u1_gt_239_U181 ( .A1(u1_gt_239_n459), .A2(u1_gt_239_n26), .A3(
        u1_gt_239_n460), .ZN(u1_gt_239_n458) );
  NOR2_X2 u1_gt_239_U180 ( .A1(u1_gt_239_n137), .A2(u1_gt_239_n34), .ZN(
        u1_gt_239_n739) );
  NOR2_X2 u1_gt_239_U179 ( .A1(u1_gt_239_n135), .A2(u1_gt_239_n136), .ZN(
        u1_gt_239_n740) );
  NOR2_X2 u1_gt_239_U178 ( .A1(u1_gt_239_n10), .A2(u1_gt_239_n20), .ZN(
        u1_gt_239_n734) );
  NOR2_X2 u1_gt_239_U177 ( .A1(u1_gt_239_n22), .A2(u1_gt_239_n16), .ZN(
        u1_gt_239_n733) );
  NOR2_X1 u1_gt_239_U176 ( .A1(u1_gt_239_n103), .A2(u1_gt_239_n104), .ZN(
        u1_gt_239_n736) );
  NOR2_X2 u1_gt_239_U175 ( .A1(n8456), .A2(u1_gt_239_n102), .ZN(u1_gt_239_n735) );
  NAND3_X2 u1_gt_239_U174 ( .A1(u1_gt_239_n735), .A2(u1_gt_239_n9), .A3(
        u1_gt_239_n736), .ZN(u1_gt_239_n731) );
  NOR3_X2 u1_gt_239_U173 ( .A1(u1_gt_239_n20), .A2(u1_gt_239_n163), .A3(
        u1_gt_239_n22), .ZN(u1_gt_239_n719) );
  NOR2_X2 u1_gt_239_U172 ( .A1(u1_gt_239_n16), .A2(u1_gt_239_n135), .ZN(
        u1_gt_239_n693) );
  NAND3_X1 u1_gt_239_U171 ( .A1(u1_gt_239_n692), .A2(u1_gt_239_n24), .A3(
        u1_gt_239_n693), .ZN(u1_gt_239_n688) );
  NOR2_X1 u1_gt_239_U170 ( .A1(u1_gt_239_n160), .A2(u1_gt_239_n10), .ZN(
        u1_gt_239_n687) );
  NAND3_X2 u1_gt_239_U169 ( .A1(u1_gt_239_n685), .A2(u1_gt_239_n686), .A3(
        u1_gt_239_n687), .ZN(u1_gt_239_n683) );
  NAND3_X2 u1_gt_239_U168 ( .A1(u1_gt_239_n681), .A2(u1_gt_239_n473), .A3(
        u1_gt_239_n682), .ZN(u1_gt_239_n678) );
  NOR3_X1 u1_gt_239_U167 ( .A1(u1_gt_239_n8), .A2(u1_gt_239_n102), .A3(
        u1_gt_239_n474), .ZN(u1_gt_239_n715) );
  NOR3_X1 u1_gt_239_U166 ( .A1(u1_gt_239_n476), .A2(u1_gt_239_n475), .A3(
        u1_gt_239_n452), .ZN(u1_gt_239_n714) );
  NOR2_X2 u1_gt_239_U165 ( .A1(u1_gt_239_n663), .A2(u1_gt_239_n662), .ZN(
        u1_gt_239_n799) );
  NOR3_X1 u1_gt_239_U164 ( .A1(u1_gt_239_n828), .A2(u1_gt_239_n160), .A3(
        u1_gt_239_n10), .ZN(u1_gt_239_n817) );
  NOR3_X2 u1_gt_239_U163 ( .A1(u1_gt_239_n840), .A2(u1_gt_239_n27), .A3(
        u1_gt_239_n841), .ZN(u1_gt_239_n830) );
  NOR2_X2 u1_gt_239_U162 ( .A1(u1_gt_239_n136), .A2(u1_gt_239_n135), .ZN(
        u1_gt_239_n749) );
  NAND3_X2 u1_gt_239_U161 ( .A1(u1_gt_239_n749), .A2(u1_gt_239_n17), .A3(
        u1_gt_239_n750), .ZN(u1_gt_239_n747) );
  NOR2_X2 u1_gt_239_U160 ( .A1(u1_gt_239_n345), .A2(u1_gt_239_n141), .ZN(
        u1_gt_239_n785) );
  NAND3_X2 u1_gt_239_U159 ( .A1(u1_gt_239_n781), .A2(u1_gt_239_n11), .A3(
        u1_gt_239_n782), .ZN(u1_gt_239_n778) );
  NOR2_X1 u1_gt_239_U158 ( .A1(u1_gt_239_n103), .A2(u1_gt_239_n104), .ZN(
        u1_gt_239_n768) );
  NOR2_X2 u1_gt_239_U157 ( .A1(u1_gt_239_n20), .A2(u1_gt_239_n22), .ZN(
        u1_gt_239_n767) );
  NAND3_X2 u1_gt_239_U156 ( .A1(u1_gt_239_n767), .A2(u1_gt_239_n11), .A3(
        u1_gt_239_n768), .ZN(u1_gt_239_n761) );
  NAND3_X1 u1_gt_239_U155 ( .A1(u1_gt_239_n559), .A2(u1_gt_239_n560), .A3(
        u1_gt_239_n561), .ZN(u1_gt_239_n556) );
  NOR3_X2 u1_gt_239_U154 ( .A1(u1_gt_239_n20), .A2(u1_gt_239_n142), .A3(
        u1_gt_239_n22), .ZN(u1_gt_239_n575) );
  NOR2_X2 u1_gt_239_U153 ( .A1(u1_gt_239_n137), .A2(u1_gt_239_n34), .ZN(
        u1_gt_239_n576) );
  NOR2_X2 u1_gt_239_U152 ( .A1(u1_gt_239_n345), .A2(u1_gt_239_n141), .ZN(
        u1_gt_239_n574) );
  NOR2_X1 u1_gt_239_U151 ( .A1(u1_gt_239_n162), .A2(u1_gt_239_n163), .ZN(
        u1_gt_239_n570) );
  NOR2_X1 u1_gt_239_U150 ( .A1(u1_gt_239_n104), .A2(u1_gt_239_n160), .ZN(
        u1_gt_239_n571) );
  NAND3_X2 u1_gt_239_U149 ( .A1(u1_gt_239_n570), .A2(u1_gt_239_n11), .A3(
        u1_gt_239_n571), .ZN(u1_gt_239_n563) );
  NOR3_X2 u1_gt_239_U148 ( .A1(u1_gt_239_n639), .A2(u1_gt_239_n137), .A3(
        u1_gt_239_n33), .ZN(u1_gt_239_n623) );
  NAND3_X2 u1_gt_239_U147 ( .A1(u1_gt_239_n635), .A2(u1_gt_239_n25), .A3(
        u1_gt_239_n636), .ZN(u1_gt_239_n634) );
  NOR3_X2 u1_gt_239_U146 ( .A1(u1_gt_239_n20), .A2(u1_gt_239_n142), .A3(
        u1_gt_239_n22), .ZN(u1_gt_239_n629) );
  NOR2_X2 u1_gt_239_U145 ( .A1(u1_gt_239_n20), .A2(u1_gt_239_n22), .ZN(
        u1_gt_239_n614) );
  NAND3_X2 u1_gt_239_U144 ( .A1(u1_gt_239_n618), .A2(u1_gt_239_n79), .A3(
        u1_gt_239_n619), .ZN(u1_gt_239_n616) );
  NOR2_X2 u1_gt_239_U143 ( .A1(u1_gt_239_n86), .A2(u1_gt_239_n31), .ZN(
        u1_gt_239_n651) );
  NOR2_X2 u1_gt_239_U142 ( .A1(u1_gt_239_n88), .A2(u1_gt_239_n653), .ZN(
        u1_gt_239_n652) );
  NOR2_X2 u1_gt_239_U141 ( .A1(u1_gt_239_n113), .A2(u1_gt_239_n650), .ZN(
        u1_gt_239_n640) );
  NOR3_X1 u1_gt_239_U140 ( .A1(u1_gt_239_n108), .A2(u1_gt_239_n662), .A3(
        u1_gt_239_n562), .ZN(u1_gt_239_n708) );
  NOR3_X2 u1_gt_239_U139 ( .A1(u1_gt_239_n699), .A2(u1_gt_239_n88), .A3(
        u1_gt_239_n30), .ZN(u1_gt_239_n698) );
  NOR3_X2 u1_gt_239_U138 ( .A1(u1_gt_239_n345), .A2(u1_gt_239_n22), .A3(
        u1_gt_239_n142), .ZN(u1_gt_239_n838) );
  NOR3_X1 u1_gt_239_U137 ( .A1(u1_gt_239_n20), .A2(u1_gt_239_n162), .A3(
        u1_gt_239_n163), .ZN(u1_gt_239_n839) );
  NOR3_X2 u1_gt_239_U136 ( .A1(u1_gt_239_n793), .A2(u1_gt_239_n86), .A3(
        u1_gt_239_n30), .ZN(u1_gt_239_n792) );
  NOR3_X2 u1_gt_239_U135 ( .A1(u1_gt_239_n562), .A2(n8413), .A3(u1_gt_239_n662), .ZN(u1_gt_239_n777) );
  NOR3_X1 u1_gt_239_U134 ( .A1(u1_gt_239_n110), .A2(u1_gt_239_n108), .A3(
        u1_gt_239_n107), .ZN(u1_gt_239_n776) );
  NOR2_X2 u1_gt_239_U133 ( .A1(u1_gt_239_n241), .A2(u1_gt_239_n204), .ZN(
        u1_gt_239_n580) );
  NOR3_X2 u1_gt_239_U132 ( .A1(u1_gt_239_n583), .A2(u1_gt_239_n86), .A3(
        u1_gt_239_n30), .ZN(u1_gt_239_n581) );
  NOR2_X1 u1_gt_239_U131 ( .A1(u1_gt_239_n476), .A2(u1_gt_239_n452), .ZN(
        u1_gt_239_n669) );
  NOR2_X1 u1_gt_239_U130 ( .A1(u1_gt_239_n475), .A2(u1_gt_239_n474), .ZN(
        u1_gt_239_n668) );
  NAND3_X2 u1_gt_239_U129 ( .A1(u1_gt_239_n668), .A2(u1_gt_239_n9), .A3(
        u1_gt_239_n669), .ZN(u1_gt_239_n664) );
  NOR3_X2 u1_gt_239_U128 ( .A1(u1_gt_239_n107), .A2(u1_gt_239_n562), .A3(
        u1_gt_239_n108), .ZN(u1_gt_239_n660) );
  NOR2_X2 u1_gt_239_U127 ( .A1(u1_gt_239_n255), .A2(u1_gt_239_n256), .ZN(
        u1_gt_239_n254) );
  NOR2_X2 u1_gt_239_U126 ( .A1(u1_gt_239_n62), .A2(u1_gt_239_n63), .ZN(
        u1_gt_239_n37) );
  NOR2_X2 u1_gt_239_U125 ( .A1(u1_gt_239_n45), .A2(u1_gt_239_n46), .ZN(
        u1_gt_239_n44) );
  NOR2_X2 u1_gt_239_U124 ( .A1(u1_gt_239_n45), .A2(u1_gt_239_n48), .ZN(
        u1_gt_239_n43) );
  NOR2_X2 u1_gt_239_U123 ( .A1(u1_gt_239_n43), .A2(u1_gt_239_n44), .ZN(
        u1_gt_239_n42) );
  NOR2_X1 u1_gt_239_U122 ( .A1(u1_gt_239_n45), .A2(u1_gt_239_n52), .ZN(
        u1_gt_239_n51) );
  NOR2_X2 u1_gt_239_U121 ( .A1(u1_gt_239_n45), .A2(u1_gt_239_n53), .ZN(
        u1_gt_239_n50) );
  NOR3_X2 u1_gt_239_U120 ( .A1(u1_gt_239_n49), .A2(u1_gt_239_n50), .A3(
        u1_gt_239_n51), .ZN(u1_gt_239_n41) );
  NOR2_X1 u1_gt_239_U119 ( .A1(n8369), .A2(u1_gt_239_n61), .ZN(u1_gt_239_n60)
         );
  NOR2_X1 u1_gt_239_U118 ( .A1(n8368), .A2(u1_gt_239_n59), .ZN(u1_gt_239_n57)
         );
  NOR3_X2 u1_gt_239_U117 ( .A1(u1_gt_239_n503), .A2(u1_gt_239_n31), .A3(
        u1_gt_239_n504), .ZN(u1_gt_239_n492) );
  NOR2_X2 u1_gt_239_U116 ( .A1(u1_gt_239_n518), .A2(u1_gt_239_n519), .ZN(
        u1_gt_239_n489) );
  NOR3_X2 u1_gt_239_U115 ( .A1(u1_gt_239_n491), .A2(u1_gt_239_n492), .A3(
        u1_gt_239_n493), .ZN(u1_gt_239_n490) );
  NOR2_X2 u1_gt_239_U114 ( .A1(u1_gt_239_n384), .A2(u1_gt_239_n385), .ZN(
        u1_gt_239_n383) );
  NOR3_X2 u1_gt_239_U113 ( .A1(u1_gt_239_n427), .A2(u1_gt_239_n428), .A3(
        u1_gt_239_n429), .ZN(u1_gt_239_n382) );
  NOR2_X2 u1_gt_239_U112 ( .A1(u1_gt_239_n549), .A2(u1_gt_239_n550), .ZN(
        u1_gt_239_n548) );
  NOR2_X2 u1_gt_239_U111 ( .A1(u1_gt_239_n741), .A2(u1_gt_239_n742), .ZN(
        u1_gt_239_n546) );
  NOR2_X2 u1_gt_239_U110 ( .A1(u1_gt_239_n670), .A2(u1_gt_239_n671), .ZN(
        u1_gt_239_n547) );
  NOR2_X2 u1_gt_239_U109 ( .A1(u1_gt_239_n137), .A2(u1_gt_239_n34), .ZN(
        u1_gt_239_n332) );
  NOR2_X2 u1_gt_239_U108 ( .A1(u1_gt_239_n135), .A2(u1_gt_239_n136), .ZN(
        u1_gt_239_n333) );
  NOR2_X2 u1_gt_239_U107 ( .A1(u1_gt_239_n103), .A2(u1_gt_239_n104), .ZN(
        u1_gt_239_n327) );
  NOR2_X2 u1_gt_239_U106 ( .A1(u1_gt_239_n10), .A2(u1_gt_239_n20), .ZN(
        u1_gt_239_n329) );
  NOR2_X2 u1_gt_239_U105 ( .A1(n8455), .A2(u1_gt_239_n8), .ZN(u1_gt_239_n328)
         );
  NAND3_X2 u1_gt_239_U104 ( .A1(u1_gt_239_n327), .A2(u1_gt_239_n328), .A3(
        u1_gt_239_n329), .ZN(u1_gt_239_n326) );
  NOR2_X1 u1_gt_239_U103 ( .A1(u1_gt_239_n241), .A2(u1_gt_239_n204), .ZN(
        u1_gt_239_n320) );
  NOR2_X1 u1_gt_239_U102 ( .A1(u1_gt_239_n86), .A2(u1_gt_239_n87), .ZN(
        u1_gt_239_n349) );
  NAND3_X2 u1_gt_239_U101 ( .A1(u1_gt_239_n348), .A2(u1_gt_239_n144), .A3(
        u1_gt_239_n349), .ZN(u1_gt_239_n347) );
  NOR2_X1 u1_gt_239_U100 ( .A1(u1_gt_239_n241), .A2(u1_gt_239_n204), .ZN(
        u1_gt_239_n351) );
  NOR3_X2 u1_gt_239_U99 ( .A1(u1_gt_239_n345), .A2(u1_gt_239_n22), .A3(
        u1_gt_239_n142), .ZN(u1_gt_239_n344) );
  NOR3_X2 u1_gt_239_U98 ( .A1(u1_gt_239_n345), .A2(u1_gt_239_n22), .A3(
        u1_gt_239_n142), .ZN(u1_gt_239_n363) );
  NOR3_X1 u1_gt_239_U97 ( .A1(u1_gt_239_n20), .A2(n8444), .A3(u1_gt_239_n163), 
        .ZN(u1_gt_239_n364) );
  NOR2_X2 u1_gt_239_U96 ( .A1(u1_gt_239_n136), .A2(u1_gt_239_n137), .ZN(
        u1_gt_239_n365) );
  NOR2_X1 u1_gt_239_U95 ( .A1(u1_gt_239_n28), .A2(u1_gt_239_n378), .ZN(
        u1_gt_239_n368) );
  NOR3_X1 u1_gt_239_U94 ( .A1(u1_gt_239_n16), .A2(u1_gt_239_n136), .A3(
        u1_gt_239_n135), .ZN(u1_gt_239_n371) );
  NOR3_X2 u1_gt_239_U93 ( .A1(u1_gt_239_n29), .A2(u1_gt_239_n6), .A3(
        u1_gt_239_n376), .ZN(u1_gt_239_n369) );
  NOR2_X2 u1_gt_239_U92 ( .A1(n8441), .A2(u1_gt_239_n22), .ZN(u1_gt_239_n374)
         );
  NAND3_X1 u1_gt_239_U91 ( .A1(u1_gt_239_n374), .A2(u1_gt_239_n165), .A3(
        u1_gt_239_n375), .ZN(u1_gt_239_n372) );
  NOR2_X2 u1_gt_239_U90 ( .A1(u1_gt_239_n20), .A2(u1_gt_239_n22), .ZN(
        u1_gt_239_n215) );
  NAND3_X2 u1_gt_239_U89 ( .A1(u1_gt_239_n119), .A2(u1_gt_239_n215), .A3(
        u1_gt_239_n17), .ZN(u1_gt_239_n208) );
  NAND3_X2 u1_gt_239_U88 ( .A1(u1_gt_239_n78), .A2(u1_gt_239_n197), .A3(
        u1_gt_239_n77), .ZN(u1_gt_239_n760) );
  NOR2_X2 u1_gt_239_U87 ( .A1(u1_gt_239_n104), .A2(u1_gt_239_n10), .ZN(
        u1_gt_239_n230) );
  NOR2_X2 u1_gt_239_U86 ( .A1(u1_gt_239_n20), .A2(u1_gt_239_n22), .ZN(
        u1_gt_239_n229) );
  NOR2_X2 u1_gt_239_U85 ( .A1(n8457), .A2(u1_gt_239_n234), .ZN(u1_gt_239_n231)
         );
  NOR2_X1 u1_gt_239_U84 ( .A1(u1_gt_239_n8), .A2(u1_gt_239_n103), .ZN(
        u1_gt_239_n233) );
  NOR2_X1 u1_gt_239_U83 ( .A1(u1_gt_239_n86), .A2(u1_gt_239_n87), .ZN(
        u1_gt_239_n154) );
  NAND3_X2 u1_gt_239_U82 ( .A1(u1_gt_239_n153), .A2(u1_gt_239_n25), .A3(
        u1_gt_239_n154), .ZN(u1_gt_239_n152) );
  NOR2_X1 u1_gt_239_U81 ( .A1(u1_gt_239_n141), .A2(u1_gt_239_n16), .ZN(
        u1_gt_239_n140) );
  NOR2_X2 u1_gt_239_U80 ( .A1(n8440), .A2(u1_gt_239_n142), .ZN(u1_gt_239_n138)
         );
  NAND3_X2 u1_gt_239_U79 ( .A1(u1_gt_239_n138), .A2(u1_gt_239_n24), .A3(
        u1_gt_239_n140), .ZN(u1_gt_239_n131) );
  NOR2_X2 u1_gt_239_U78 ( .A1(u1_gt_239_n135), .A2(u1_gt_239_n136), .ZN(
        u1_gt_239_n134) );
  NOR3_X2 u1_gt_239_U77 ( .A1(u1_gt_239_n109), .A2(u1_gt_239_n101), .A3(
        u1_gt_239_n111), .ZN(u1_gt_239_n175) );
  NOR3_X1 u1_gt_239_U76 ( .A1(u1_gt_239_n110), .A2(n8410), .A3(u1_gt_239_n107), 
        .ZN(u1_gt_239_n176) );
  NOR2_X1 u1_gt_239_U75 ( .A1(u1_gt_239_n88), .A2(u1_gt_239_n86), .ZN(
        u1_gt_239_n288) );
  NOR2_X2 u1_gt_239_U74 ( .A1(u1_gt_239_n10), .A2(u1_gt_239_n20), .ZN(
        u1_gt_239_n295) );
  NOR2_X2 u1_gt_239_U73 ( .A1(n8459), .A2(u1_gt_239_n102), .ZN(u1_gt_239_n296)
         );
  NOR2_X1 u1_gt_239_U72 ( .A1(n8439), .A2(u1_gt_239_n141), .ZN(u1_gt_239_n514)
         );
  NOR2_X2 u1_gt_239_U71 ( .A1(u1_gt_239_n136), .A2(u1_gt_239_n137), .ZN(
        u1_gt_239_n513) );
  NOR2_X2 u1_gt_239_U70 ( .A1(u1_gt_239_n33), .A2(u1_gt_239_n241), .ZN(
        u1_gt_239_n512) );
  NOR2_X1 u1_gt_239_U69 ( .A1(u1_gt_239_n142), .A2(u1_gt_239_n141), .ZN(
        u1_gt_239_n485) );
  NOR2_X2 u1_gt_239_U68 ( .A1(u1_gt_239_n136), .A2(u1_gt_239_n137), .ZN(
        u1_gt_239_n484) );
  NOR2_X2 u1_gt_239_U67 ( .A1(u1_gt_239_n34), .A2(u1_gt_239_n241), .ZN(
        u1_gt_239_n483) );
  NOR2_X2 u1_gt_239_U66 ( .A1(u1_gt_239_n33), .A2(u1_gt_239_n241), .ZN(
        u1_gt_239_n393) );
  NOR2_X2 u1_gt_239_U65 ( .A1(n8438), .A2(u1_gt_239_n141), .ZN(u1_gt_239_n395)
         );
  NOR2_X1 u1_gt_239_U64 ( .A1(u1_gt_239_n102), .A2(u1_gt_239_n8), .ZN(
        u1_gt_239_n422) );
  NOR2_X1 u1_gt_239_U63 ( .A1(n8462), .A2(u1_gt_239_n101), .ZN(u1_gt_239_n420)
         );
  NOR2_X2 u1_gt_239_U62 ( .A1(u1_gt_239_n137), .A2(u1_gt_239_n34), .ZN(
        u1_gt_239_n720) );
  NOR3_X2 u1_gt_239_U61 ( .A1(u1_gt_239_n345), .A2(u1_gt_239_n142), .A3(
        u1_gt_239_n141), .ZN(u1_gt_239_n718) );
  NOR2_X2 u1_gt_239_U60 ( .A1(u1_gt_239_n136), .A2(u1_gt_239_n137), .ZN(
        u1_gt_239_n691) );
  NOR2_X2 u1_gt_239_U59 ( .A1(u1_gt_239_n34), .A2(u1_gt_239_n241), .ZN(
        u1_gt_239_n690) );
  NOR2_X2 u1_gt_239_U58 ( .A1(u1_gt_239_n20), .A2(u1_gt_239_n22), .ZN(
        u1_gt_239_n685) );
  NOR2_X1 u1_gt_239_U57 ( .A1(u1_gt_239_n162), .A2(u1_gt_239_n163), .ZN(
        u1_gt_239_n686) );
  NOR2_X2 u1_gt_239_U56 ( .A1(n8409), .A2(u1_gt_239_n110), .ZN(u1_gt_239_n682)
         );
  NOR2_X2 u1_gt_239_U55 ( .A1(u1_gt_239_n137), .A2(u1_gt_239_n34), .ZN(
        u1_gt_239_n750) );
  NOR3_X2 u1_gt_239_U54 ( .A1(u1_gt_239_n20), .A2(u1_gt_239_n142), .A3(
        u1_gt_239_n22), .ZN(u1_gt_239_n786) );
  NOR2_X1 u1_gt_239_U53 ( .A1(u1_gt_239_n104), .A2(u1_gt_239_n160), .ZN(
        u1_gt_239_n782) );
  NOR2_X1 u1_gt_239_U52 ( .A1(u1_gt_239_n162), .A2(u1_gt_239_n163), .ZN(
        u1_gt_239_n781) );
  NOR2_X2 u1_gt_239_U51 ( .A1(n8412), .A2(u1_gt_239_n562), .ZN(u1_gt_239_n559)
         );
  NOR2_X2 u1_gt_239_U50 ( .A1(u1_gt_239_n107), .A2(u1_gt_239_n110), .ZN(
        u1_gt_239_n561) );
  NOR2_X2 u1_gt_239_U49 ( .A1(u1_gt_239_n86), .A2(u1_gt_239_n87), .ZN(
        u1_gt_239_n636) );
  NOR2_X2 u1_gt_239_U48 ( .A1(u1_gt_239_n241), .A2(u1_gt_239_n204), .ZN(
        u1_gt_239_n638) );
  NOR3_X2 u1_gt_239_U47 ( .A1(u1_gt_239_n16), .A2(u1_gt_239_n345), .A3(
        u1_gt_239_n141), .ZN(u1_gt_239_n628) );
  NOR2_X1 u1_gt_239_U46 ( .A1(u1_gt_239_n104), .A2(u1_gt_239_n160), .ZN(
        u1_gt_239_n630) );
  NOR2_X2 u1_gt_239_U45 ( .A1(n8449), .A2(u1_gt_239_n103), .ZN(u1_gt_239_n631)
         );
  NOR2_X1 u1_gt_239_U44 ( .A1(u1_gt_239_n162), .A2(u1_gt_239_n163), .ZN(
        u1_gt_239_n615) );
  NOR3_X2 u1_gt_239_U43 ( .A1(u1_gt_239_n87), .A2(u1_gt_239_n30), .A3(
        u1_gt_239_n362), .ZN(u1_gt_239_n361) );
  NOR3_X2 u1_gt_239_U42 ( .A1(u1_gt_239_n302), .A2(u1_gt_239_n303), .A3(
        u1_gt_239_n304), .ZN(u1_gt_239_n253) );
  NOR2_X2 u1_gt_239_U41 ( .A1(u1_gt_239_n238), .A2(u1_gt_239_n239), .ZN(
        u1_gt_239_n237) );
  AOI21_X1 u1_gt_239_U40 ( .B1(u1_gt_239_n236), .B2(u1_gt_239_n116), .A(
        u1_gt_239_n237), .ZN(u1_gt_239_n64) );
  NOR2_X2 u1_gt_239_U39 ( .A1(u1_gt_239_n181), .A2(u1_gt_239_n182), .ZN(
        u1_gt_239_n65) );
  NOR2_X2 u1_gt_239_U38 ( .A1(u1_gt_239_n123), .A2(u1_gt_239_n124), .ZN(
        u1_gt_239_n66) );
  OAI21_X2 u1_gt_239_U37 ( .B1(u1_gt_239_n70), .B2(u1_gt_239_n71), .A(
        u1_gt_239_n72), .ZN(u1_gt_239_n69) );
  NOR2_X2 u1_gt_239_U36 ( .A1(u1_gt_239_n68), .A2(u1_gt_239_n69), .ZN(
        u1_gt_239_n67) );
  NOR2_X2 u1_gt_239_U35 ( .A1(u1_gt_239_n260), .A2(u1_gt_239_n261), .ZN(
        u1_gt_239_n259) );
  NOR3_X1 u1_gt_239_U34 ( .A1(u1_gt_239_n29), .A2(u1_gt_239_n7), .A3(
        u1_gt_239_n516), .ZN(u1_gt_239_n508) );
  NOR2_X1 u1_gt_239_U33 ( .A1(u1_gt_239_n204), .A2(u1_gt_239_n28), .ZN(
        u1_gt_239_n507) );
  NOR2_X1 u1_gt_239_U32 ( .A1(u1_gt_239_n527), .A2(u1_gt_239_n29), .ZN(
        u1_gt_239_n522) );
  NOR2_X2 u1_gt_239_U31 ( .A1(u1_gt_239_n540), .A2(u1_gt_239_n541), .ZN(
        u1_gt_239_n537) );
  NOR2_X2 u1_gt_239_U30 ( .A1(u1_gt_239_n402), .A2(u1_gt_239_n403), .ZN(
        u1_gt_239_n401) );
  NOR2_X2 u1_gt_239_U29 ( .A1(u1_gt_239_n425), .A2(u1_gt_239_n426), .ZN(
        u1_gt_239_n424) );
  NOR3_X1 u1_gt_239_U28 ( .A1(u1_gt_239_n16), .A2(u1_gt_239_n345), .A3(
        u1_gt_239_n141), .ZN(u1_gt_239_n448) );
  NOR2_X2 u1_gt_239_U27 ( .A1(u1_gt_239_n22), .A2(u1_gt_239_n142), .ZN(
        u1_gt_239_n446) );
  NOR2_X2 u1_gt_239_U26 ( .A1(u1_gt_239_n163), .A2(u1_gt_239_n20), .ZN(
        u1_gt_239_n447) );
  NOR3_X1 u1_gt_239_U25 ( .A1(u1_gt_239_n10), .A2(u1_gt_239_n160), .A3(
        u1_gt_239_n162), .ZN(u1_gt_239_n451) );
  NOR2_X1 u1_gt_239_U24 ( .A1(u1_gt_239_n103), .A2(u1_gt_239_n104), .ZN(
        u1_gt_239_n449) );
  NOR2_X1 u1_gt_239_U23 ( .A1(n8450), .A2(u1_gt_239_n452), .ZN(u1_gt_239_n450)
         );
  NOR2_X2 u1_gt_239_U22 ( .A1(u1_gt_239_n458), .A2(u1_gt_239_n29), .ZN(
        u1_gt_239_n453) );
  NOR2_X2 u1_gt_239_U21 ( .A1(u1_gt_239_n28), .A2(u1_gt_239_n457), .ZN(
        u1_gt_239_n454) );
  NOR2_X2 u1_gt_239_U20 ( .A1(n4397), .A2(u1_gt_239_n802), .ZN(u1_gt_239_n801)
         );
  NOR3_X2 u1_gt_239_U19 ( .A1(u1_gt_239_n562), .A2(u1_gt_239_n1), .A3(
        u1_gt_239_n801), .ZN(u1_gt_239_n800) );
  NOR2_X2 u1_gt_239_U18 ( .A1(u1_gt_239_n345), .A2(u1_gt_239_n141), .ZN(
        u1_gt_239_n375) );
  INV_X8 u1_gt_239_U17 ( .A(u1_gt_239_n89), .ZN(u1_gt_239_n32) );
  INV_X4 u1_gt_239_U16 ( .A(u1_gt_239_n192), .ZN(u1_gt_239_n163) );
  INV_X8 u1_gt_239_U15 ( .A(u1_gt_239_n161), .ZN(u1_gt_239_n19) );
  INV_X8 u1_gt_239_U14 ( .A(u1_gt_239_n165), .ZN(u1_gt_239_n142) );
  INV_X8 u1_gt_239_U13 ( .A(u1_gt_239_n216), .ZN(u1_gt_239_n21) );
  INV_X16 u1_gt_239_U12 ( .A(u1_gt_239_n24), .ZN(u1_gt_239_n345) );
  INV_X8 u1_gt_239_U11 ( .A(u1_gt_239_n223), .ZN(u1_gt_239_n27) );
  INV_X16 u1_gt_239_U10 ( .A(u1_gt_239_n201), .ZN(u1_gt_239_n87) );
  INV_X16 u1_gt_239_U9 ( .A(u1_gt_239_n35), .ZN(u1_gt_239_n34) );
  NAND2_X2 u1_gt_239_U8 ( .A1(n8433), .A2(u1_gt_239_n290), .ZN(u1_gt_239_n80)
         );
  INV_X4 u1_gt_239_U7 ( .A(u1_gt_239_n80), .ZN(u1_gt_239_n14) );
  INV_X4 u1_gt_239_U6 ( .A(u1_gt_239_n139), .ZN(u1_gt_239_n23) );
  INV_X4 u1_gt_239_U5 ( .A(u1_gt_239_n81), .ZN(u1_gt_239_n12) );
  INV_X8 u1_gt_239_U4 ( .A(u1_gt_239_n112), .ZN(u1_gt_239_n35) );
  NOR3_X1 u1_gt_239_U3 ( .A1(u1_gt_239_n16), .A2(u1_gt_239_n141), .A3(
        u1_gt_239_n135), .ZN(u1_gt_239_n366) );
  INV_X16 u1_gt_239_U2 ( .A(u1_gt_239_n32), .ZN(u1_gt_239_n30) );
  AND2_X2 u1_gt_239_U1 ( .A1(n8420), .A2(u1_gt_239_n653), .ZN(u1_gt_239_n1) );
  INV_X4 u4_sub_496_U95 ( .A(u4_ldz_all_0_), .ZN(u4_sub_496_n52) );
  NAND2_X2 u4_sub_496_U94 ( .A1(u4_exp_in_pl1_0_), .A2(u4_sub_496_n52), .ZN(
        u4_sub_496_n32) );
  INV_X4 u4_sub_496_U93 ( .A(u4_exp_in_pl1_0_), .ZN(u4_sub_496_n51) );
  NAND2_X2 u4_sub_496_U92 ( .A1(u4_ldz_all_0_), .A2(u4_sub_496_n51), .ZN(
        u4_sub_496_n42) );
  NAND2_X2 u4_sub_496_U91 ( .A1(u4_sub_496_n32), .A2(u4_sub_496_n42), .ZN(
        u4_div_exp2_0_) );
  INV_X4 u4_sub_496_U90 ( .A(u4_sub_496_net61360), .ZN(u4_sub_496_net61437) );
  NOR2_X4 u4_sub_496_U89 ( .A1(u4_sub_496_net61437), .A2(u4_sub_496_net61438), 
        .ZN(u4_sub_496_n35) );
  NAND2_X2 u4_sub_496_U88 ( .A1(u4_sub_496_net61430), .A2(u4_sub_496_net61352), 
        .ZN(u4_sub_496_net61429) );
  INV_X4 u4_sub_496_U87 ( .A(u4_exp_in_pl1_2_), .ZN(u4_sub_496_n49) );
  NAND2_X2 u4_sub_496_U86 ( .A1(u4_ldz_all_2_), .A2(u4_sub_496_n49), .ZN(
        u4_sub_496_n21) );
  INV_X4 u4_sub_496_U85 ( .A(u4_exp_in_pl1_1_), .ZN(u4_sub_496_n48) );
  NAND2_X2 u4_sub_496_U84 ( .A1(u4_ldz_all_1_), .A2(u4_sub_496_n48), .ZN(
        u4_sub_496_n33) );
  INV_X4 u4_sub_496_U83 ( .A(u4_sub_496_n33), .ZN(u4_sub_496_n27) );
  INV_X4 u4_sub_496_U82 ( .A(u4_ldz_all_1_), .ZN(u4_sub_496_n47) );
  NAND2_X2 u4_sub_496_U81 ( .A1(u4_exp_in_pl1_1_), .A2(u4_sub_496_n47), .ZN(
        u4_sub_496_n28) );
  INV_X4 u4_sub_496_U80 ( .A(u4_ldz_all_2_), .ZN(u4_sub_496_n46) );
  NAND2_X2 u4_sub_496_U79 ( .A1(u4_exp_in_pl1_2_), .A2(u4_sub_496_n46), .ZN(
        u4_sub_496_n19) );
  OAI211_X2 u4_sub_496_U78 ( .C1(u4_sub_496_n27), .C2(u4_sub_496_n32), .A(
        u4_sub_496_n28), .B(u4_sub_496_n19), .ZN(u4_sub_496_n44) );
  INV_X4 u4_sub_496_U77 ( .A(u4_exp_in_pl1_3_), .ZN(u4_sub_496_n45) );
  NAND3_X2 u4_sub_496_U76 ( .A1(u4_sub_496_n21), .A2(u4_sub_496_n44), .A3(
        u4_sub_496_n24), .ZN(u4_sub_496_n39) );
  NAND2_X2 u4_sub_496_U75 ( .A1(u4_exp_in_pl1_3_), .A2(u4_sub_496_n43), .ZN(
        u4_sub_496_n23) );
  INV_X4 u4_sub_496_U74 ( .A(u4_sub_496_n31), .ZN(u4_sub_496_n41) );
  INV_X4 u4_sub_496_U73 ( .A(u4_exp_in_pl1_4_), .ZN(u4_sub_496_n38) );
  NAND2_X2 u4_sub_496_U72 ( .A1(u4_ldz_all_4_), .A2(u4_sub_496_n38), .ZN(
        u4_sub_496_net61389) );
  NAND2_X2 u4_sub_496_U71 ( .A1(u4_sub_496_net61355), .A2(u4_sub_496_net61354), 
        .ZN(u4_sub_496_n37) );
  XNOR2_X2 u4_sub_496_U70 ( .A(u4_exp_in_pl1_10_), .B(u4_sub_496_n34), .ZN(
        u4_div_exp2_10_) );
  NAND2_X2 u4_sub_496_U69 ( .A1(u4_sub_496_n28), .A2(u4_sub_496_n33), .ZN(
        u4_sub_496_n30) );
  NAND2_X2 u4_sub_496_U68 ( .A1(u4_sub_496_n31), .A2(u4_sub_496_n32), .ZN(
        u4_sub_496_n29) );
  XNOR2_X2 u4_sub_496_U67 ( .A(u4_sub_496_n30), .B(u4_sub_496_n29), .ZN(
        u4_div_exp2_1_) );
  NAND2_X2 u4_sub_496_U66 ( .A1(u4_sub_496_n21), .A2(u4_sub_496_n19), .ZN(
        u4_sub_496_n25) );
  INV_X4 u4_sub_496_U65 ( .A(u4_sub_496_n29), .ZN(u4_sub_496_n26) );
  OAI21_X4 u4_sub_496_U64 ( .B1(u4_sub_496_n26), .B2(u4_sub_496_n27), .A(
        u4_sub_496_n28), .ZN(u4_sub_496_n22) );
  XNOR2_X2 u4_sub_496_U63 ( .A(u4_sub_496_n25), .B(u4_sub_496_n22), .ZN(
        u4_div_exp2_2_) );
  NAND2_X2 u4_sub_496_U62 ( .A1(u4_sub_496_n23), .A2(u4_sub_496_n24), .ZN(
        u4_sub_496_n17) );
  NAND2_X2 u4_sub_496_U61 ( .A1(u4_sub_496_n21), .A2(u4_sub_496_n22), .ZN(
        u4_sub_496_n20) );
  NAND2_X2 u4_sub_496_U60 ( .A1(u4_sub_496_n19), .A2(u4_sub_496_n20), .ZN(
        u4_sub_496_n18) );
  XNOR2_X2 u4_sub_496_U59 ( .A(u4_sub_496_n17), .B(u4_sub_496_n18), .ZN(
        u4_div_exp2_3_) );
  XNOR2_X2 u4_sub_496_U58 ( .A(u4_sub_496_net61387), .B(u4_sub_496_n16), .ZN(
        u4_div_exp2_4_) );
  INV_X4 u4_sub_496_U57 ( .A(u4_sub_496_net61370), .ZN(u4_sub_496_net61369) );
  XNOR2_X2 u4_sub_496_U56 ( .A(u4_sub_496_net61365), .B(u4_sub_496_net61437), 
        .ZN(u4_div_exp2_8_) );
  INV_X4 u4_sub_496_U55 ( .A(u4_sub_496_n15), .ZN(u4_sub_496_n14) );
  NOR2_X4 u4_sub_496_U54 ( .A1(u4_sub_496_n14), .A2(u4_sub_496_net61358), .ZN(
        u4_sub_496_n12) );
  NAND2_X2 u4_sub_496_U53 ( .A1(u4_sub_496_n12), .A2(u4_sub_496_n13), .ZN(
        u4_sub_496_n11) );
  XNOR2_X2 u4_sub_496_U52 ( .A(u4_sub_496_n11), .B(u4_sub_496_net61347), .ZN(
        u4_div_exp2_9_) );
  INV_X4 u4_sub_496_U51 ( .A(u4_exp_in_pl1_8_), .ZN(u4_sub_496_net61360) );
  INV_X4 u4_sub_496_U50 ( .A(u4_exp_in_pl1_9_), .ZN(u4_sub_496_net61349) );
  INV_X4 u4_sub_496_U49 ( .A(u4_sub_496_n42), .ZN(u4_sub_496_n31) );
  NAND2_X2 u4_sub_496_U48 ( .A1(u4_sub_496_net61363), .A2(u4_sub_496_net61364), 
        .ZN(u4_sub_496_net61368) );
  INV_X4 u4_sub_496_U47 ( .A(u4_sub_496_net61370), .ZN(u4_sub_496_net61411) );
  NAND2_X2 u4_sub_496_U46 ( .A1(u4_sub_496_net61364), .A2(u4_sub_496_net61363), 
        .ZN(u4_sub_496_n36) );
  NAND2_X2 u4_sub_496_U45 ( .A1(u4_sub_496_net61363), .A2(u4_sub_496_net61364), 
        .ZN(u4_sub_496_n15) );
  INV_X4 u4_sub_496_U44 ( .A(u4_sub_496_net61349), .ZN(u4_sub_496_net61347) );
  NAND3_X4 u4_sub_496_U43 ( .A1(u4_sub_496_n39), .A2(u4_sub_496_n23), .A3(
        u4_sub_496_n40), .ZN(u4_sub_496_n16) );
  NAND2_X2 u4_sub_496_U42 ( .A1(u4_sub_496_net61359), .A2(u4_sub_496_net61360), 
        .ZN(u4_sub_496_net61358) );
  NAND2_X2 u4_sub_496_U41 ( .A1(u4_sub_496_net61359), .A2(u4_sub_496_net61349), 
        .ZN(u4_sub_496_net61438) );
  INV_X4 u4_sub_496_U40 ( .A(u4_exp_in_pl1_7_), .ZN(u4_sub_496_net61359) );
  INV_X4 u4_sub_496_U39 ( .A(u4_sub_496_net61359), .ZN(u4_sub_496_net61372) );
  NAND2_X2 u4_sub_496_U38 ( .A1(u4_ldz_all_6_), .A2(u4_sub_496_n10), .ZN(
        u4_sub_496_net61354) );
  NAND2_X2 u4_sub_496_U37 ( .A1(u4_ldz_all_6_), .A2(u4_sub_496_n10), .ZN(
        u4_sub_496_net61364) );
  INV_X4 u4_sub_496_U36 ( .A(u4_exp_in_pl1_6_), .ZN(u4_sub_496_n10) );
  NAND2_X2 u4_sub_496_U35 ( .A1(u4_sub_496_net61354), .A2(u4_sub_496_net61376), 
        .ZN(u4_sub_496_net61379) );
  XNOR2_X2 u4_sub_496_U34 ( .A(u4_sub_496_n7), .B(u4_sub_496_net61372), .ZN(
        u4_div_exp2_7_) );
  NAND2_X1 u4_sub_496_U33 ( .A1(u4_sub_496_net61386), .A2(u4_sub_496_net61389), 
        .ZN(u4_sub_496_net61387) );
  INV_X2 u4_sub_496_U32 ( .A(u4_sub_496_net61386), .ZN(u4_sub_496_net61430) );
  INV_X4 u4_sub_496_U31 ( .A(u4_sub_496_net61385), .ZN(u4_sub_496_net61355) );
  NAND2_X4 u4_sub_496_U30 ( .A1(u4_sub_496_net61385), .A2(u4_sub_496_net61386), 
        .ZN(u4_sub_496_net61383) );
  INV_X4 u4_sub_496_U29 ( .A(u4_exp_in_pl1_5_), .ZN(u4_sub_496_n5) );
  INV_X4 u4_sub_496_U28 ( .A(u4_ldz_all_5_), .ZN(u4_sub_496_n6) );
  NAND2_X2 u4_sub_496_U27 ( .A1(u4_sub_496_net61352), .A2(u4_sub_496_net61382), 
        .ZN(u4_sub_496_n4) );
  INV_X4 u4_sub_496_U26 ( .A(u4_sub_496_net61352), .ZN(u4_sub_496_net61381) );
  INV_X4 u4_sub_496_U25 ( .A(u4_sub_496_n2), .ZN(u4_sub_496_net61374) );
  OAI21_X4 u4_sub_496_U24 ( .B1(u4_sub_496_n3), .B2(u4_sub_496_net61381), .A(
        u4_sub_496_net61382), .ZN(u4_sub_496_n2) );
  NAND2_X4 u4_sub_496_U23 ( .A1(u4_ldz_all_5_), .A2(u4_sub_496_n5), .ZN(
        u4_sub_496_net61352) );
  NAND3_X1 u4_sub_496_U22 ( .A1(u4_sub_496_net61354), .A2(u4_sub_496_net61355), 
        .A3(u4_sub_496_net61352), .ZN(u4_sub_496_n13) );
  NAND2_X4 u4_sub_496_U21 ( .A1(u4_exp_in_pl1_4_), .A2(u4_sub_496_n50), .ZN(
        u4_sub_496_net61386) );
  INV_X4 u4_sub_496_U20 ( .A(u4_ldz_all_4_), .ZN(u4_sub_496_n50) );
  NAND2_X4 u4_sub_496_U19 ( .A1(u4_exp_in_pl1_6_), .A2(u4_sub_496_n9), .ZN(
        u4_sub_496_net61376) );
  OAI21_X4 u4_sub_496_U18 ( .B1(u4_sub_496_net61374), .B2(u4_sub_496_n8), .A(
        u4_sub_496_net61376), .ZN(u4_sub_496_n7) );
  NAND4_X4 u4_sub_496_U17 ( .A1(u4_sub_496_n41), .A2(u4_sub_496_n33), .A3(
        u4_sub_496_n21), .A4(u4_sub_496_n24), .ZN(u4_sub_496_n40) );
  NAND3_X2 u4_sub_496_U16 ( .A1(u4_sub_496_net61382), .A2(u4_sub_496_net61376), 
        .A3(u4_sub_496_net61429), .ZN(u4_sub_496_net61363) );
  INV_X8 u4_sub_496_U15 ( .A(u4_sub_496_net61383), .ZN(u4_sub_496_n3) );
  INV_X1 u4_sub_496_U14 ( .A(u4_sub_496_n3), .ZN(u4_sub_496_n1) );
  INV_X4 u4_sub_496_U13 ( .A(u4_ldz_all_6_), .ZN(u4_sub_496_n9) );
  XNOR2_X2 u4_sub_496_U12 ( .A(u4_sub_496_net61379), .B(u4_sub_496_n2), .ZN(
        u4_div_exp2_6_) );
  XNOR2_X2 u4_sub_496_U11 ( .A(u4_sub_496_n4), .B(u4_sub_496_n1), .ZN(
        u4_div_exp2_5_) );
  NAND2_X4 u4_sub_496_U10 ( .A1(u4_exp_in_pl1_5_), .A2(u4_sub_496_n6), .ZN(
        u4_sub_496_net61382) );
  NOR2_X2 u4_sub_496_U9 ( .A1(u4_exp_in_pl1_6_), .A2(u4_sub_496_n9), .ZN(
        u4_sub_496_n8) );
  NOR2_X2 u4_sub_496_U8 ( .A1(u4_sub_496_net61381), .A2(u4_sub_496_n37), .ZN(
        u4_sub_496_net61370) );
  NAND3_X2 u4_sub_496_U7 ( .A1(u4_sub_496_n35), .A2(u4_sub_496_n36), .A3(
        u4_sub_496_net61411), .ZN(u4_sub_496_n34) );
  NAND3_X2 u4_sub_496_U6 ( .A1(u4_sub_496_net61359), .A2(u4_sub_496_net61368), 
        .A3(u4_sub_496_net61369), .ZN(u4_sub_496_net61365) );
  NAND2_X2 u4_sub_496_U5 ( .A1(u4_sub_496_n16), .A2(u4_sub_496_net61389), .ZN(
        u4_sub_496_net61385) );
  INV_X1 u4_sub_496_U4 ( .A(u4_ldz_all_3_), .ZN(u4_sub_496_n43) );
  NAND2_X2 u4_sub_496_U3 ( .A1(u4_ldz_all_3_), .A2(u4_sub_496_n45), .ZN(
        u4_sub_496_n24) );
  INV_X32 u4_sll_454_U577 ( .A(u4_sll_454_net63277), .ZN(u4_sll_454_net63259)
         );
  INV_X32 u4_sll_454_U576 ( .A(u4_sll_454_net66455), .ZN(u4_sll_454_net66445)
         );
  INV_X32 u4_sll_454_U575 ( .A(u4_sll_454_net66455), .ZN(u4_sll_454_net66443)
         );
  INV_X32 u4_sll_454_U574 ( .A(u4_sll_454_net66451), .ZN(u4_sll_454_net66441)
         );
  INV_X32 u4_sll_454_U573 ( .A(u4_sll_454_net66451), .ZN(u4_sll_454_net66439)
         );
  INV_X32 u4_sll_454_U572 ( .A(u4_sll_454_net66455), .ZN(u4_sll_454_net66429)
         );
  INV_X32 u4_sll_454_U571 ( .A(u4_sll_454_net66509), .ZN(u4_sll_454_net66501)
         );
  INV_X32 u4_sll_454_U570 ( .A(u4_sll_454_net66509), .ZN(u4_sll_454_net66499)
         );
  INV_X32 u4_sll_454_U569 ( .A(u4_sll_454_net66509), .ZN(u4_sll_454_net66497)
         );
  INV_X32 u4_sll_454_U568 ( .A(u4_sll_454_net66509), .ZN(u4_sll_454_net66495)
         );
  INV_X32 u4_sll_454_U567 ( .A(u4_sll_454_net66509), .ZN(u4_sll_454_net66493)
         );
  INV_X32 u4_sll_454_U566 ( .A(u4_sll_454_net66509), .ZN(u4_sll_454_net66485)
         );
  INV_X32 u4_sll_454_U565 ( .A(u4_sll_454_net66591), .ZN(u4_sll_454_net66557)
         );
  INV_X32 u4_sll_454_U564 ( .A(u4_sll_454_net66563), .ZN(u4_sll_454_net66551)
         );
  INV_X32 u4_sll_454_U563 ( .A(u4_sll_454_net66563), .ZN(u4_sll_454_net66549)
         );
  INV_X32 u4_sll_454_U562 ( .A(u4_sll_454_net66619), .ZN(u4_sll_454_net66609)
         );
  INV_X32 u4_sll_454_U561 ( .A(u4_sll_454_net66619), .ZN(u4_sll_454_net66607)
         );
  INV_X32 u4_sll_454_U560 ( .A(u4_sll_454_net66699), .ZN(u4_sll_454_net66673)
         );
  INV_X32 u4_sll_454_U559 ( .A(u4_sll_454_net66673), .ZN(u4_sll_454_net66667)
         );
  INV_X32 u4_sll_454_U558 ( .A(u4_sll_454_net66675), .ZN(u4_sll_454_net66663)
         );
  INV_X32 u4_sll_454_U557 ( .A(u4_sll_454_net66757), .ZN(u4_sll_454_net66723)
         );
  INV_X4 u4_sll_454_U556 ( .A(net33546), .ZN(u4_sll_454_n233) );
  NOR2_X4 u4_sll_454_U555 ( .A1(u4_sll_454_net66373), .A2(u4_sll_454_n233), 
        .ZN(u4_sll_454_ML_int_1__0_) );
  INV_X4 u4_sll_454_U554 ( .A(u4_sll_454_ML_int_1__0_), .ZN(u4_sll_454_n232)
         );
  INV_X4 u4_sll_454_U553 ( .A(u4_sll_454_ML_int_1__1_), .ZN(u4_sll_454_n231)
         );
  INV_X4 u4_sll_454_U552 ( .A(u4_sll_454_ML_int_2__0_), .ZN(u4_sll_454_n230)
         );
  INV_X4 u4_sll_454_U551 ( .A(u4_sll_454_ML_int_2__1_), .ZN(u4_sll_454_n229)
         );
  NOR2_X4 u4_sll_454_U550 ( .A1(u4_sll_454_net66667), .A2(u4_sll_454_n229), 
        .ZN(u4_sll_454_ML_int_3__1_) );
  INV_X4 u4_sll_454_U549 ( .A(u4_sll_454_ML_int_2__2_), .ZN(u4_sll_454_n228)
         );
  NOR2_X4 u4_sll_454_U548 ( .A1(u4_sll_454_net66667), .A2(u4_sll_454_n228), 
        .ZN(u4_sll_454_ML_int_3__2_) );
  INV_X4 u4_sll_454_U547 ( .A(u4_sll_454_ML_int_2__3_), .ZN(u4_sll_454_n227)
         );
  NOR2_X4 u4_sll_454_U546 ( .A1(u4_sll_454_net66667), .A2(u4_sll_454_n227), 
        .ZN(u4_sll_454_ML_int_3__3_) );
  INV_X4 u4_sll_454_U545 ( .A(u4_sll_454_ML_int_3__0_), .ZN(u4_sll_454_n226)
         );
  INV_X4 u4_sll_454_U544 ( .A(u4_sll_454_ML_int_3__1_), .ZN(u4_sll_454_n225)
         );
  INV_X4 u4_sll_454_U543 ( .A(u4_sll_454_ML_int_3__2_), .ZN(u4_sll_454_n224)
         );
  NOR2_X4 u4_sll_454_U542 ( .A1(u4_sll_454_net66611), .A2(u4_sll_454_n224), 
        .ZN(u4_sll_454_ML_int_4__2_) );
  INV_X4 u4_sll_454_U541 ( .A(u4_sll_454_ML_int_3__3_), .ZN(u4_sll_454_n223)
         );
  NOR2_X4 u4_sll_454_U540 ( .A1(u4_sll_454_net66611), .A2(u4_sll_454_n223), 
        .ZN(u4_sll_454_ML_int_4__3_) );
  INV_X4 u4_sll_454_U539 ( .A(u4_sll_454_ML_int_3__4_), .ZN(u4_sll_454_n222)
         );
  NOR2_X4 u4_sll_454_U538 ( .A1(u4_sll_454_net66611), .A2(u4_sll_454_n222), 
        .ZN(u4_sll_454_ML_int_4__4_) );
  INV_X4 u4_sll_454_U537 ( .A(u4_sll_454_ML_int_3__5_), .ZN(u4_sll_454_n221)
         );
  NOR2_X4 u4_sll_454_U536 ( .A1(u4_sll_454_net66611), .A2(u4_sll_454_n221), 
        .ZN(u4_sll_454_ML_int_4__5_) );
  INV_X4 u4_sll_454_U535 ( .A(u4_sll_454_ML_int_3__6_), .ZN(u4_sll_454_n220)
         );
  NOR2_X4 u4_sll_454_U534 ( .A1(u4_sll_454_net66611), .A2(u4_sll_454_n220), 
        .ZN(u4_sll_454_ML_int_4__6_) );
  INV_X4 u4_sll_454_U533 ( .A(u4_sll_454_ML_int_3__7_), .ZN(u4_sll_454_n219)
         );
  NOR2_X4 u4_sll_454_U532 ( .A1(u4_sll_454_net66613), .A2(u4_sll_454_n219), 
        .ZN(u4_sll_454_ML_int_4__7_) );
  INV_X4 u4_sll_454_U531 ( .A(u4_sll_454_ML_int_4__0_), .ZN(u4_sll_454_n218)
         );
  NOR2_X4 u4_sll_454_U530 ( .A1(u4_sll_454_net66557), .A2(u4_sll_454_n218), 
        .ZN(u4_sll_454_ML_int_5__0_) );
  INV_X4 u4_sll_454_U529 ( .A(u4_sll_454_ML_int_4__1_), .ZN(u4_sll_454_n217)
         );
  NOR2_X4 u4_sll_454_U528 ( .A1(u4_sll_454_net66557), .A2(u4_sll_454_n217), 
        .ZN(u4_sll_454_ML_int_5__1_) );
  INV_X4 u4_sll_454_U527 ( .A(u4_sll_454_ML_int_4__2_), .ZN(u4_sll_454_n216)
         );
  NOR2_X4 u4_sll_454_U526 ( .A1(u4_sll_454_net66557), .A2(u4_sll_454_n216), 
        .ZN(u4_sll_454_ML_int_5__2_) );
  INV_X4 u4_sll_454_U525 ( .A(u4_sll_454_ML_int_4__3_), .ZN(u4_sll_454_n215)
         );
  NOR2_X4 u4_sll_454_U524 ( .A1(u4_sll_454_net66557), .A2(u4_sll_454_n215), 
        .ZN(u4_sll_454_ML_int_5__3_) );
  INV_X4 u4_sll_454_U523 ( .A(u4_sll_454_ML_int_4__4_), .ZN(u4_sll_454_n214)
         );
  NOR2_X4 u4_sll_454_U522 ( .A1(u4_sll_454_net66557), .A2(u4_sll_454_n214), 
        .ZN(u4_sll_454_ML_int_5__4_) );
  INV_X4 u4_sll_454_U521 ( .A(u4_sll_454_ML_int_4__5_), .ZN(u4_sll_454_n213)
         );
  NOR2_X4 u4_sll_454_U520 ( .A1(u4_sll_454_net66557), .A2(u4_sll_454_n213), 
        .ZN(u4_sll_454_ML_int_5__5_) );
  INV_X4 u4_sll_454_U519 ( .A(u4_sll_454_ML_int_4__6_), .ZN(u4_sll_454_n212)
         );
  NOR2_X4 u4_sll_454_U518 ( .A1(u4_sll_454_net66557), .A2(u4_sll_454_n212), 
        .ZN(u4_sll_454_ML_int_5__6_) );
  INV_X4 u4_sll_454_U517 ( .A(u4_sll_454_ML_int_4__7_), .ZN(u4_sll_454_n211)
         );
  NOR2_X4 u4_sll_454_U516 ( .A1(u4_sll_454_net66557), .A2(u4_sll_454_n211), 
        .ZN(u4_sll_454_ML_int_5__7_) );
  INV_X4 u4_sll_454_U515 ( .A(u4_sll_454_ML_int_4__8_), .ZN(u4_sll_454_n210)
         );
  NOR2_X4 u4_sll_454_U514 ( .A1(u4_sll_454_net66557), .A2(u4_sll_454_n210), 
        .ZN(u4_sll_454_ML_int_5__8_) );
  INV_X4 u4_sll_454_U513 ( .A(u4_sll_454_ML_int_4__9_), .ZN(u4_sll_454_n209)
         );
  NOR2_X4 u4_sll_454_U512 ( .A1(u4_sll_454_net66557), .A2(u4_sll_454_n209), 
        .ZN(u4_sll_454_ML_int_5__9_) );
  INV_X4 u4_sll_454_U511 ( .A(u4_sll_454_ML_int_4__10_), .ZN(u4_sll_454_n208)
         );
  NOR2_X4 u4_sll_454_U510 ( .A1(u4_sll_454_net66557), .A2(u4_sll_454_n208), 
        .ZN(u4_sll_454_ML_int_5__10_) );
  INV_X4 u4_sll_454_U509 ( .A(u4_sll_454_ML_int_4__11_), .ZN(u4_sll_454_n207)
         );
  NOR2_X4 u4_sll_454_U508 ( .A1(u4_sll_454_net66551), .A2(u4_sll_454_n207), 
        .ZN(u4_sll_454_ML_int_5__11_) );
  INV_X4 u4_sll_454_U507 ( .A(u4_sll_454_ML_int_4__12_), .ZN(
        u4_sll_454__UDW__89915_net72603) );
  NOR2_X4 u4_sll_454_U506 ( .A1(u4_sll_454_net66551), .A2(
        u4_sll_454__UDW__89915_net72603), .ZN(u4_sll_454_ML_int_5__12_) );
  INV_X4 u4_sll_454_U505 ( .A(u4_sll_454_ML_int_4__13_), .ZN(u4_sll_454_n206)
         );
  NOR2_X4 u4_sll_454_U504 ( .A1(u4_sll_454_net66551), .A2(u4_sll_454_n206), 
        .ZN(u4_sll_454_ML_int_5__13_) );
  INV_X4 u4_sll_454_U503 ( .A(u4_sll_454_ML_int_4__14_), .ZN(u4_sll_454_n205)
         );
  NOR2_X4 u4_sll_454_U502 ( .A1(u4_sll_454_net66551), .A2(u4_sll_454_n205), 
        .ZN(u4_sll_454_ML_int_5__14_) );
  INV_X4 u4_sll_454_U501 ( .A(u4_sll_454_ML_int_4__15_), .ZN(u4_sll_454_n204)
         );
  NOR2_X4 u4_sll_454_U500 ( .A1(u4_sll_454_net66551), .A2(u4_sll_454_n204), 
        .ZN(u4_sll_454_ML_int_5__15_) );
  INV_X4 u4_sll_454_U499 ( .A(u4_sll_454_ML_int_5__0_), .ZN(u4_sll_454_n203)
         );
  NOR2_X4 u4_sll_454_U498 ( .A1(u4_sll_454_net66485), .A2(u4_sll_454_n203), 
        .ZN(u4_sll_454_ML_int_6__0_) );
  INV_X4 u4_sll_454_U497 ( .A(u4_sll_454_ML_int_5__1_), .ZN(u4_sll_454_n202)
         );
  NOR2_X4 u4_sll_454_U496 ( .A1(u4_sll_454_net66485), .A2(u4_sll_454_n202), 
        .ZN(u4_sll_454_ML_int_6__1_) );
  INV_X4 u4_sll_454_U495 ( .A(u4_sll_454_ML_int_5__2_), .ZN(u4_sll_454_n201)
         );
  NOR2_X4 u4_sll_454_U494 ( .A1(u4_sll_454_net66485), .A2(u4_sll_454_n201), 
        .ZN(u4_sll_454_ML_int_6__2_) );
  INV_X4 u4_sll_454_U493 ( .A(u4_sll_454_ML_int_5__3_), .ZN(u4_sll_454_n200)
         );
  NOR2_X4 u4_sll_454_U492 ( .A1(u4_sll_454_net66485), .A2(u4_sll_454_n200), 
        .ZN(u4_sll_454_ML_int_6__3_) );
  INV_X4 u4_sll_454_U491 ( .A(u4_sll_454_ML_int_5__4_), .ZN(u4_sll_454_n199)
         );
  NOR2_X4 u4_sll_454_U490 ( .A1(u4_sll_454_net66485), .A2(u4_sll_454_n199), 
        .ZN(u4_sll_454_ML_int_6__4_) );
  INV_X4 u4_sll_454_U489 ( .A(u4_sll_454_ML_int_5__5_), .ZN(u4_sll_454_n198)
         );
  NOR2_X4 u4_sll_454_U488 ( .A1(u4_sll_454_net66485), .A2(u4_sll_454_n198), 
        .ZN(u4_sll_454_ML_int_6__5_) );
  INV_X4 u4_sll_454_U487 ( .A(u4_sll_454_ML_int_5__6_), .ZN(u4_sll_454_n197)
         );
  NOR2_X4 u4_sll_454_U486 ( .A1(u4_sll_454_net66485), .A2(u4_sll_454_n197), 
        .ZN(u4_sll_454_ML_int_6__6_) );
  INV_X4 u4_sll_454_U485 ( .A(u4_sll_454_ML_int_5__7_), .ZN(u4_sll_454_n196)
         );
  NOR2_X4 u4_sll_454_U484 ( .A1(u4_sll_454_net66501), .A2(u4_sll_454_n196), 
        .ZN(u4_sll_454_ML_int_6__7_) );
  INV_X4 u4_sll_454_U483 ( .A(u4_sll_454_ML_int_5__8_), .ZN(u4_sll_454_n195)
         );
  NOR2_X4 u4_sll_454_U482 ( .A1(u4_sll_454_net66501), .A2(u4_sll_454_n195), 
        .ZN(u4_sll_454_ML_int_6__8_) );
  INV_X4 u4_sll_454_U481 ( .A(u4_sll_454_ML_int_5__9_), .ZN(u4_sll_454_n194)
         );
  NOR2_X4 u4_sll_454_U480 ( .A1(u4_sll_454_net66501), .A2(u4_sll_454_n194), 
        .ZN(u4_sll_454_ML_int_6__9_) );
  INV_X4 u4_sll_454_U479 ( .A(u4_sll_454_ML_int_5__10_), .ZN(u4_sll_454_n193)
         );
  NOR2_X4 u4_sll_454_U478 ( .A1(u4_sll_454_net66501), .A2(u4_sll_454_n193), 
        .ZN(u4_sll_454_ML_int_6__10_) );
  INV_X4 u4_sll_454_U477 ( .A(u4_sll_454_ML_int_5__11_), .ZN(u4_sll_454_n192)
         );
  NOR2_X4 u4_sll_454_U476 ( .A1(u4_sll_454_net66485), .A2(u4_sll_454_n192), 
        .ZN(u4_sll_454_ML_int_6__11_) );
  INV_X4 u4_sll_454_U475 ( .A(u4_sll_454_ML_int_5__12_), .ZN(
        u4_sll_454__UDW__89963_net72763) );
  NOR2_X4 u4_sll_454_U474 ( .A1(u4_sll_454_net66485), .A2(
        u4_sll_454__UDW__89963_net72763), .ZN(u4_sll_454_ML_int_6__12_) );
  INV_X4 u4_sll_454_U473 ( .A(u4_sll_454_ML_int_5__13_), .ZN(u4_sll_454_n191)
         );
  NOR2_X4 u4_sll_454_U472 ( .A1(u4_sll_454_net66485), .A2(u4_sll_454_n191), 
        .ZN(u4_sll_454_ML_int_6__13_) );
  INV_X4 u4_sll_454_U471 ( .A(u4_sll_454_ML_int_5__14_), .ZN(u4_sll_454_n190)
         );
  NOR2_X4 u4_sll_454_U470 ( .A1(u4_sll_454_net66485), .A2(u4_sll_454_n190), 
        .ZN(u4_sll_454_ML_int_6__14_) );
  INV_X4 u4_sll_454_U469 ( .A(u4_sll_454_ML_int_5__15_), .ZN(u4_sll_454_n189)
         );
  NOR2_X4 u4_sll_454_U468 ( .A1(u4_sll_454_net66485), .A2(u4_sll_454_n189), 
        .ZN(u4_sll_454_ML_int_6__15_) );
  INV_X4 u4_sll_454_U467 ( .A(u4_sll_454_ML_int_5__16_), .ZN(u4_sll_454_n188)
         );
  NOR2_X4 u4_sll_454_U466 ( .A1(u4_sll_454_net66485), .A2(u4_sll_454_n188), 
        .ZN(u4_sll_454_ML_int_6__16_) );
  INV_X4 u4_sll_454_U465 ( .A(u4_sll_454_ML_int_5__17_), .ZN(u4_sll_454_n187)
         );
  NOR2_X4 u4_sll_454_U464 ( .A1(u4_sll_454_net66485), .A2(u4_sll_454_n187), 
        .ZN(u4_sll_454_ML_int_6__17_) );
  INV_X4 u4_sll_454_U463 ( .A(u4_sll_454_ML_int_5__18_), .ZN(u4_sll_454_n186)
         );
  NOR2_X4 u4_sll_454_U462 ( .A1(u4_sll_454_net66485), .A2(u4_sll_454_n186), 
        .ZN(u4_sll_454_ML_int_6__18_) );
  INV_X4 u4_sll_454_U461 ( .A(u4_sll_454_ML_int_5__19_), .ZN(u4_sll_454_n185)
         );
  NOR2_X4 u4_sll_454_U460 ( .A1(u4_sll_454_net66485), .A2(u4_sll_454_n185), 
        .ZN(u4_sll_454_ML_int_6__19_) );
  INV_X4 u4_sll_454_U459 ( .A(u4_sll_454_ML_int_5__20_), .ZN(u4_sll_454_n184)
         );
  NOR2_X4 u4_sll_454_U458 ( .A1(u4_sll_454_net66485), .A2(u4_sll_454_n184), 
        .ZN(u4_sll_454_ML_int_6__20_) );
  INV_X4 u4_sll_454_U457 ( .A(u4_sll_454_ML_int_5__21_), .ZN(u4_sll_454_n183)
         );
  NOR2_X4 u4_sll_454_U456 ( .A1(u4_sll_454_net66485), .A2(u4_sll_454_n183), 
        .ZN(u4_sll_454_ML_int_6__21_) );
  INV_X4 u4_sll_454_U455 ( .A(u4_sll_454_ML_int_5__22_), .ZN(u4_sll_454_n182)
         );
  NOR2_X4 u4_sll_454_U454 ( .A1(u4_sll_454_net66487), .A2(u4_sll_454_n182), 
        .ZN(u4_sll_454_ML_int_6__22_) );
  INV_X4 u4_sll_454_U453 ( .A(u4_sll_454_ML_int_5__23_), .ZN(u4_sll_454_n181)
         );
  NOR2_X4 u4_sll_454_U452 ( .A1(u4_sll_454_net66487), .A2(u4_sll_454_n181), 
        .ZN(u4_sll_454_ML_int_6__23_) );
  INV_X4 u4_sll_454_U451 ( .A(u4_sll_454_ML_int_5__24_), .ZN(u4_sll_454_n180)
         );
  NOR2_X4 u4_sll_454_U450 ( .A1(u4_sll_454_net66487), .A2(u4_sll_454_n180), 
        .ZN(u4_sll_454_ML_int_6__24_) );
  INV_X4 u4_sll_454_U449 ( .A(u4_sll_454_ML_int_5__25_), .ZN(u4_sll_454_n179)
         );
  NOR2_X4 u4_sll_454_U448 ( .A1(u4_sll_454_net66487), .A2(u4_sll_454_n179), 
        .ZN(u4_sll_454_ML_int_6__25_) );
  INV_X4 u4_sll_454_U447 ( .A(u4_sll_454_ML_int_5__26_), .ZN(u4_sll_454_n178)
         );
  NOR2_X4 u4_sll_454_U446 ( .A1(u4_sll_454_net66487), .A2(u4_sll_454_n178), 
        .ZN(u4_sll_454_ML_int_6__26_) );
  INV_X4 u4_sll_454_U445 ( .A(u4_sll_454_ML_int_5__27_), .ZN(u4_sll_454_n177)
         );
  NOR2_X4 u4_sll_454_U444 ( .A1(u4_sll_454_net66487), .A2(u4_sll_454_n177), 
        .ZN(u4_sll_454_ML_int_6__27_) );
  INV_X4 u4_sll_454_U443 ( .A(u4_sll_454_ML_int_5__28_), .ZN(
        u4_sll_454__UDW__90011_net72923) );
  NOR2_X4 u4_sll_454_U442 ( .A1(u4_sll_454_net66487), .A2(
        u4_sll_454__UDW__90011_net72923), .ZN(u4_sll_454_ML_int_6__28_) );
  INV_X4 u4_sll_454_U441 ( .A(u4_sll_454_ML_int_5__29_), .ZN(u4_sll_454_n176)
         );
  NOR2_X4 u4_sll_454_U440 ( .A1(u4_sll_454_net66487), .A2(u4_sll_454_n176), 
        .ZN(u4_sll_454_ML_int_6__29_) );
  INV_X4 u4_sll_454_U439 ( .A(u4_sll_454_ML_int_5__30_), .ZN(u4_sll_454_n175)
         );
  NOR2_X4 u4_sll_454_U438 ( .A1(u4_sll_454_net66487), .A2(u4_sll_454_n175), 
        .ZN(u4_sll_454_ML_int_6__30_) );
  INV_X4 u4_sll_454_U437 ( .A(u4_sll_454_ML_int_5__31_), .ZN(u4_sll_454_n174)
         );
  NOR2_X4 u4_sll_454_U436 ( .A1(u4_sll_454_net66487), .A2(u4_sll_454_n174), 
        .ZN(u4_sll_454_ML_int_6__31_) );
  INV_X4 u4_sll_454_U435 ( .A(u4_sll_454_ML_int_6__0_), .ZN(u4_sll_454_n173)
         );
  NOR2_X4 u4_sll_454_U434 ( .A1(u4_sll_454_net66429), .A2(u4_sll_454_n173), 
        .ZN(u4_sll_454_ML_int_7__0_) );
  INV_X4 u4_sll_454_U433 ( .A(u4_sll_454_ML_int_6__1_), .ZN(u4_sll_454_n172)
         );
  NOR2_X4 u4_sll_454_U432 ( .A1(u4_sll_454_net66429), .A2(u4_sll_454_n172), 
        .ZN(u4_sll_454_ML_int_7__1_) );
  INV_X4 u4_sll_454_U431 ( .A(u4_sll_454_ML_int_6__2_), .ZN(u4_sll_454_n171)
         );
  INV_X4 u4_sll_454_U430 ( .A(u4_sll_454_ML_int_6__3_), .ZN(u4_sll_454_n170)
         );
  INV_X4 u4_sll_454_U429 ( .A(u4_sll_454_ML_int_6__4_), .ZN(u4_sll_454_n169)
         );
  INV_X4 u4_sll_454_U428 ( .A(u4_sll_454_ML_int_6__5_), .ZN(u4_sll_454_n168)
         );
  INV_X4 u4_sll_454_U427 ( .A(u4_sll_454_ML_int_6__6_), .ZN(u4_sll_454_n167)
         );
  INV_X4 u4_sll_454_U426 ( .A(u4_sll_454_ML_int_6__7_), .ZN(u4_sll_454_n166)
         );
  INV_X4 u4_sll_454_U425 ( .A(u4_sll_454_ML_int_6__8_), .ZN(u4_sll_454_n165)
         );
  INV_X4 u4_sll_454_U424 ( .A(u4_sll_454_ML_int_6__9_), .ZN(u4_sll_454_n164)
         );
  INV_X4 u4_sll_454_U423 ( .A(u4_sll_454_ML_int_6__10_), .ZN(u4_sll_454_n163)
         );
  INV_X4 u4_sll_454_U422 ( .A(u4_sll_454_ML_int_6__11_), .ZN(u4_sll_454_n162)
         );
  NOR2_X4 u4_sll_454_U421 ( .A1(u4_sll_454_net66429), .A2(u4_sll_454_n162), 
        .ZN(u4_sll_454_ML_int_7__11_) );
  INV_X4 u4_sll_454_U420 ( .A(u4_sll_454_ML_int_6__12_), .ZN(u4_sll_454_n161)
         );
  INV_X4 u4_sll_454_U419 ( .A(u4_sll_454_ML_int_6__13_), .ZN(u4_sll_454_n160)
         );
  INV_X4 u4_sll_454_U418 ( .A(u4_sll_454_ML_int_6__14_), .ZN(u4_sll_454_n159)
         );
  INV_X4 u4_sll_454_U417 ( .A(u4_sll_454_ML_int_6__15_), .ZN(u4_sll_454_n158)
         );
  INV_X4 u4_sll_454_U416 ( .A(u4_sll_454_ML_int_6__16_), .ZN(u4_sll_454_n157)
         );
  INV_X4 u4_sll_454_U415 ( .A(u4_sll_454_ML_int_6__17_), .ZN(u4_sll_454_n156)
         );
  INV_X4 u4_sll_454_U414 ( .A(u4_sll_454_ML_int_6__18_), .ZN(u4_sll_454_n155)
         );
  NOR2_X4 u4_sll_454_U413 ( .A1(u4_sll_454_net66429), .A2(u4_sll_454_n155), 
        .ZN(u4_sll_454_ML_int_7__18_) );
  INV_X4 u4_sll_454_U412 ( .A(u4_sll_454_ML_int_6__19_), .ZN(u4_sll_454_n154)
         );
  INV_X4 u4_sll_454_U411 ( .A(u4_sll_454_ML_int_6__20_), .ZN(u4_sll_454_n153)
         );
  NOR2_X4 u4_sll_454_U410 ( .A1(u4_sll_454_net66429), .A2(u4_sll_454_n153), 
        .ZN(u4_sll_454_ML_int_7__20_) );
  INV_X4 u4_sll_454_U409 ( .A(u4_sll_454_ML_int_6__21_), .ZN(u4_sll_454_n152)
         );
  NOR2_X4 u4_sll_454_U408 ( .A1(u4_sll_454_net66429), .A2(u4_sll_454_n152), 
        .ZN(u4_sll_454_ML_int_7__21_) );
  INV_X4 u4_sll_454_U407 ( .A(u4_sll_454_ML_int_6__22_), .ZN(u4_sll_454_n151)
         );
  INV_X4 u4_sll_454_U406 ( .A(u4_sll_454_ML_int_6__23_), .ZN(u4_sll_454_n150)
         );
  INV_X4 u4_sll_454_U405 ( .A(u4_sll_454_ML_int_6__24_), .ZN(u4_sll_454_n149)
         );
  INV_X4 u4_sll_454_U404 ( .A(u4_sll_454_ML_int_6__25_), .ZN(u4_sll_454_n148)
         );
  INV_X4 u4_sll_454_U403 ( .A(u4_sll_454_ML_int_6__26_), .ZN(u4_sll_454_n147)
         );
  INV_X4 u4_sll_454_U402 ( .A(u4_sll_454_ML_int_6__27_), .ZN(u4_sll_454_n146)
         );
  INV_X4 u4_sll_454_U401 ( .A(u4_sll_454_ML_int_6__28_), .ZN(u4_sll_454_n145)
         );
  INV_X4 u4_sll_454_U400 ( .A(u4_sll_454_ML_int_6__29_), .ZN(u4_sll_454_n144)
         );
  INV_X4 u4_sll_454_U399 ( .A(u4_sll_454_ML_int_6__30_), .ZN(u4_sll_454_n143)
         );
  INV_X4 u4_sll_454_U398 ( .A(u4_sll_454_ML_int_6__31_), .ZN(u4_sll_454_n142)
         );
  INV_X4 u4_sll_454_U397 ( .A(u4_sll_454_ML_int_6__32_), .ZN(u4_sll_454_n141)
         );
  INV_X4 u4_sll_454_U396 ( .A(u4_sll_454_ML_int_6__34_), .ZN(u4_sll_454_n139)
         );
  INV_X4 u4_sll_454_U395 ( .A(u4_sll_454_ML_int_6__35_), .ZN(u4_sll_454_n138)
         );
  INV_X4 u4_sll_454_U394 ( .A(u4_sll_454_ML_int_6__36_), .ZN(u4_sll_454_n137)
         );
  INV_X4 u4_sll_454_U393 ( .A(u4_sll_454_ML_int_6__37_), .ZN(u4_sll_454_n136)
         );
  INV_X4 u4_sll_454_U392 ( .A(u4_sll_454_ML_int_6__38_), .ZN(u4_sll_454_n135)
         );
  INV_X4 u4_sll_454_U391 ( .A(u4_sll_454_ML_int_6__39_), .ZN(u4_sll_454_n134)
         );
  INV_X4 u4_sll_454_U390 ( .A(u4_sll_454_ML_int_6__40_), .ZN(u4_sll_454_n133)
         );
  INV_X4 u4_sll_454_U389 ( .A(u4_sll_454_ML_int_6__41_), .ZN(u4_sll_454_n132)
         );
  INV_X4 u4_sll_454_U388 ( .A(u4_sll_454_ML_int_6__42_), .ZN(u4_sll_454_n131)
         );
  NOR2_X4 u4_sll_454_U387 ( .A1(u4_sll_454_net66433), .A2(u4_sll_454_n131), 
        .ZN(u4_sll_454_ML_int_7__42_) );
  INV_X4 u4_sll_454_U386 ( .A(u4_sll_454_ML_int_6__43_), .ZN(u4_sll_454_n130)
         );
  INV_X4 u4_sll_454_U385 ( .A(u4_sll_454_ML_int_6__45_), .ZN(u4_sll_454_n129)
         );
  NOR2_X4 u4_sll_454_U384 ( .A1(u4_sll_454_net66435), .A2(u4_sll_454_n129), 
        .ZN(u4_sll_454_ML_int_7__45_) );
  INV_X4 u4_sll_454_U383 ( .A(u4_sll_454_ML_int_6__46_), .ZN(u4_sll_454_n128)
         );
  NOR2_X4 u4_sll_454_U382 ( .A1(u4_sll_454_net66435), .A2(u4_sll_454_n128), 
        .ZN(u4_sll_454_ML_int_7__46_) );
  INV_X4 u4_sll_454_U381 ( .A(u4_sll_454_ML_int_6__47_), .ZN(u4_sll_454_n127)
         );
  INV_X4 u4_sll_454_U380 ( .A(u4_sll_454_ML_int_6__48_), .ZN(u4_sll_454_n126)
         );
  INV_X4 u4_sll_454_U379 ( .A(u4_sll_454_ML_int_6__49_), .ZN(u4_sll_454_n125)
         );
  INV_X4 u4_sll_454_U378 ( .A(u4_sll_454_ML_int_6__50_), .ZN(u4_sll_454_n124)
         );
  INV_X4 u4_sll_454_U377 ( .A(u4_sll_454_ML_int_6__51_), .ZN(u4_sll_454_n123)
         );
  INV_X4 u4_sll_454_U376 ( .A(u4_sll_454_ML_int_6__52_), .ZN(u4_sll_454_n122)
         );
  INV_X4 u4_sll_454_U375 ( .A(u4_sll_454_ML_int_6__53_), .ZN(u4_sll_454_n121)
         );
  INV_X4 u4_sll_454_U374 ( .A(u4_sll_454_ML_int_6__54_), .ZN(u4_sll_454_n120)
         );
  INV_X4 u4_sll_454_U373 ( .A(u4_sll_454_ML_int_6__55_), .ZN(u4_sll_454_n119)
         );
  INV_X4 u4_sll_454_U372 ( .A(u4_sll_454_ML_int_6__56_), .ZN(u4_sll_454_n118)
         );
  INV_X4 u4_sll_454_U371 ( .A(u4_sll_454_ML_int_6__57_), .ZN(u4_sll_454_n117)
         );
  INV_X4 u4_sll_454_U370 ( .A(u4_sll_454_ML_int_6__58_), .ZN(u4_sll_454_n116)
         );
  INV_X4 u4_sll_454_U369 ( .A(u4_sll_454_ML_int_6__59_), .ZN(u4_sll_454_n115)
         );
  INV_X4 u4_sll_454_U368 ( .A(u4_sll_454_ML_int_6__60_), .ZN(u4_sll_454_n114)
         );
  INV_X4 u4_sll_454_U367 ( .A(u4_sll_454_ML_int_6__61_), .ZN(u4_sll_454_n113)
         );
  INV_X4 u4_sll_454_U366 ( .A(u4_sll_454_ML_int_6__62_), .ZN(u4_sll_454_n112)
         );
  INV_X4 u4_sll_454_U365 ( .A(u4_sll_454_ML_int_6__63_), .ZN(u4_sll_454_n111)
         );
  INV_X4 u4_sll_454_U364 ( .A(u4_sll_454_ML_int_7__0_), .ZN(u4_sll_454_n110)
         );
  NOR2_X4 u4_sll_454_U363 ( .A1(u4_sll_454_net63273), .A2(u4_sll_454_n110), 
        .ZN(u4_N6014) );
  INV_X4 u4_sll_454_U362 ( .A(u4_sll_454_ML_int_7__1_), .ZN(u4_sll_454_n109)
         );
  NOR2_X4 u4_sll_454_U361 ( .A1(u4_sll_454_net63273), .A2(u4_sll_454_n109), 
        .ZN(u4_N6015) );
  INV_X4 u4_sll_454_U360 ( .A(u4_sll_454_ML_int_7__2_), .ZN(u4_sll_454_n108)
         );
  INV_X4 u4_sll_454_U359 ( .A(u4_sll_454_ML_int_7__3_), .ZN(u4_sll_454_n107)
         );
  INV_X4 u4_sll_454_U358 ( .A(u4_sll_454_ML_int_7__4_), .ZN(u4_sll_454_n106)
         );
  INV_X4 u4_sll_454_U357 ( .A(u4_sll_454_ML_int_7__5_), .ZN(u4_sll_454_n105)
         );
  INV_X4 u4_sll_454_U356 ( .A(u4_sll_454_ML_int_7__6_), .ZN(u4_sll_454_n104)
         );
  INV_X4 u4_sll_454_U355 ( .A(u4_sll_454_ML_int_7__7_), .ZN(u4_sll_454_n103)
         );
  INV_X4 u4_sll_454_U354 ( .A(u4_sll_454_ML_int_7__8_), .ZN(u4_sll_454_n102)
         );
  INV_X4 u4_sll_454_U353 ( .A(u4_sll_454_ML_int_7__9_), .ZN(u4_sll_454_n101)
         );
  NOR2_X4 u4_sll_454_U352 ( .A1(u4_sll_454_net63271), .A2(u4_sll_454_n101), 
        .ZN(u4_N6023) );
  INV_X4 u4_sll_454_U351 ( .A(u4_sll_454_ML_int_7__10_), .ZN(u4_sll_454_n100)
         );
  INV_X4 u4_sll_454_U350 ( .A(u4_sll_454_ML_int_7__11_), .ZN(u4_sll_454_n99)
         );
  NOR2_X4 u4_sll_454_U349 ( .A1(u4_sll_454_net63271), .A2(u4_sll_454_n99), 
        .ZN(u4_N6025) );
  INV_X4 u4_sll_454_U348 ( .A(u4_sll_454_ML_int_7__12_), .ZN(u4_sll_454_n98)
         );
  INV_X4 u4_sll_454_U347 ( .A(u4_sll_454_ML_int_7__13_), .ZN(u4_sll_454_n97)
         );
  INV_X4 u4_sll_454_U346 ( .A(u4_sll_454_ML_int_7__14_), .ZN(u4_sll_454_n96)
         );
  INV_X4 u4_sll_454_U345 ( .A(u4_sll_454_ML_int_7__15_), .ZN(u4_sll_454_n95)
         );
  INV_X4 u4_sll_454_U344 ( .A(u4_sll_454_ML_int_7__16_), .ZN(u4_sll_454_n94)
         );
  INV_X4 u4_sll_454_U343 ( .A(u4_sll_454_ML_int_7__17_), .ZN(u4_sll_454_n93)
         );
  INV_X4 u4_sll_454_U342 ( .A(u4_sll_454_ML_int_7__18_), .ZN(u4_sll_454_n92)
         );
  NOR2_X4 u4_sll_454_U341 ( .A1(u4_sll_454_net63271), .A2(u4_sll_454_n92), 
        .ZN(u4_N6032) );
  INV_X4 u4_sll_454_U340 ( .A(u4_sll_454_ML_int_7__19_), .ZN(u4_sll_454_n91)
         );
  NOR2_X4 u4_sll_454_U339 ( .A1(u4_sll_454_net63271), .A2(u4_sll_454_n91), 
        .ZN(u4_N6033) );
  INV_X4 u4_sll_454_U338 ( .A(u4_sll_454_ML_int_7__20_), .ZN(u4_sll_454_n90)
         );
  NOR2_X4 u4_sll_454_U337 ( .A1(u4_sll_454_net63271), .A2(u4_sll_454_n90), 
        .ZN(u4_N6034) );
  INV_X4 u4_sll_454_U336 ( .A(u4_sll_454_ML_int_7__21_), .ZN(u4_sll_454_n89)
         );
  NOR2_X4 u4_sll_454_U335 ( .A1(u4_sll_454_net63271), .A2(u4_sll_454_n89), 
        .ZN(u4_N6035) );
  INV_X4 u4_sll_454_U334 ( .A(u4_sll_454_ML_int_7__22_), .ZN(u4_sll_454_n88)
         );
  NOR2_X4 u4_sll_454_U333 ( .A1(u4_sll_454_net63271), .A2(u4_sll_454_n88), 
        .ZN(u4_N6036) );
  INV_X4 u4_sll_454_U332 ( .A(u4_sll_454_ML_int_7__23_), .ZN(u4_sll_454_n87)
         );
  NOR2_X4 u4_sll_454_U331 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n87), 
        .ZN(u4_N6037) );
  INV_X4 u4_sll_454_U330 ( .A(u4_sll_454_ML_int_7__24_), .ZN(u4_sll_454_n86)
         );
  NOR2_X4 u4_sll_454_U329 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n86), 
        .ZN(u4_N6038) );
  INV_X4 u4_sll_454_U328 ( .A(u4_sll_454_ML_int_7__25_), .ZN(u4_sll_454_n85)
         );
  NOR2_X4 u4_sll_454_U327 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n85), 
        .ZN(u4_N6039) );
  INV_X4 u4_sll_454_U326 ( .A(u4_sll_454_ML_int_7__26_), .ZN(u4_sll_454_n84)
         );
  NOR2_X4 u4_sll_454_U325 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n84), 
        .ZN(u4_N6040) );
  INV_X4 u4_sll_454_U324 ( .A(u4_sll_454_ML_int_7__27_), .ZN(u4_sll_454_n83)
         );
  NOR2_X4 u4_sll_454_U323 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n83), 
        .ZN(u4_N6041) );
  INV_X4 u4_sll_454_U322 ( .A(u4_sll_454_ML_int_7__28_), .ZN(u4_sll_454_n82)
         );
  INV_X4 u4_sll_454_U321 ( .A(u4_sll_454_ML_int_7__29_), .ZN(u4_sll_454_n81)
         );
  NOR2_X4 u4_sll_454_U320 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n81), 
        .ZN(u4_N6043) );
  INV_X4 u4_sll_454_U319 ( .A(u4_sll_454_ML_int_7__30_), .ZN(u4_sll_454_n80)
         );
  INV_X4 u4_sll_454_U318 ( .A(u4_sll_454_ML_int_7__31_), .ZN(u4_sll_454_n79)
         );
  NOR2_X4 u4_sll_454_U317 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n79), 
        .ZN(u4_N6045) );
  INV_X4 u4_sll_454_U316 ( .A(u4_sll_454_ML_int_7__32_), .ZN(u4_sll_454_n78)
         );
  NOR2_X4 u4_sll_454_U315 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n78), 
        .ZN(u4_N6046) );
  INV_X4 u4_sll_454_U314 ( .A(u4_sll_454_ML_int_7__33_), .ZN(u4_sll_454_n77)
         );
  NOR2_X4 u4_sll_454_U313 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n77), 
        .ZN(u4_N6047) );
  INV_X4 u4_sll_454_U312 ( .A(u4_sll_454_ML_int_7__34_), .ZN(u4_sll_454_n76)
         );
  INV_X4 u4_sll_454_U311 ( .A(u4_sll_454_ML_int_7__35_), .ZN(u4_sll_454_n75)
         );
  INV_X4 u4_sll_454_U310 ( .A(u4_sll_454_ML_int_7__36_), .ZN(u4_sll_454_n74)
         );
  INV_X4 u4_sll_454_U309 ( .A(u4_sll_454_ML_int_7__37_), .ZN(u4_sll_454_n73)
         );
  INV_X4 u4_sll_454_U308 ( .A(u4_sll_454_ML_int_7__38_), .ZN(u4_sll_454_n72)
         );
  INV_X4 u4_sll_454_U307 ( .A(u4_sll_454_ML_int_7__39_), .ZN(u4_sll_454_n71)
         );
  INV_X4 u4_sll_454_U306 ( .A(u4_sll_454_ML_int_7__40_), .ZN(u4_sll_454_n70)
         );
  NOR2_X4 u4_sll_454_U305 ( .A1(u4_sll_454_net63267), .A2(u4_sll_454_n70), 
        .ZN(u4_N6054) );
  INV_X4 u4_sll_454_U304 ( .A(u4_sll_454_ML_int_7__41_), .ZN(u4_sll_454_n69)
         );
  INV_X4 u4_sll_454_U303 ( .A(u4_sll_454_ML_int_7__42_), .ZN(u4_sll_454_n68)
         );
  NOR2_X4 u4_sll_454_U302 ( .A1(u4_sll_454_net63267), .A2(u4_sll_454_n68), 
        .ZN(u4_N6056) );
  INV_X4 u4_sll_454_U301 ( .A(u4_sll_454_ML_int_7__43_), .ZN(u4_sll_454_n67)
         );
  INV_X4 u4_sll_454_U300 ( .A(u4_sll_454_ML_int_7__45_), .ZN(u4_sll_454_n66)
         );
  NOR2_X4 u4_sll_454_U299 ( .A1(u4_sll_454_net63267), .A2(u4_sll_454_n66), 
        .ZN(u4_N6059) );
  INV_X4 u4_sll_454_U298 ( .A(u4_sll_454_ML_int_7__46_), .ZN(u4_sll_454_n65)
         );
  NOR2_X4 u4_sll_454_U297 ( .A1(u4_sll_454_net63267), .A2(u4_sll_454_n65), 
        .ZN(u4_N6060) );
  INV_X4 u4_sll_454_U296 ( .A(u4_sll_454_ML_int_7__47_), .ZN(u4_sll_454_n64)
         );
  INV_X4 u4_sll_454_U295 ( .A(u4_sll_454_ML_int_7__48_), .ZN(u4_sll_454_n63)
         );
  INV_X4 u4_sll_454_U294 ( .A(u4_sll_454_ML_int_7__49_), .ZN(u4_sll_454_n62)
         );
  INV_X4 u4_sll_454_U293 ( .A(u4_sll_454_ML_int_7__50_), .ZN(u4_sll_454_n61)
         );
  INV_X4 u4_sll_454_U292 ( .A(u4_sll_454_ML_int_7__51_), .ZN(u4_sll_454_n60)
         );
  INV_X4 u4_sll_454_U291 ( .A(u4_sll_454_ML_int_7__52_), .ZN(u4_sll_454_n59)
         );
  INV_X4 u4_sll_454_U290 ( .A(u4_sll_454_ML_int_7__53_), .ZN(u4_sll_454_n58)
         );
  INV_X4 u4_sll_454_U289 ( .A(u4_sll_454_ML_int_7__54_), .ZN(u4_sll_454_n57)
         );
  INV_X4 u4_sll_454_U288 ( .A(u4_sll_454_ML_int_7__55_), .ZN(u4_sll_454_n56)
         );
  INV_X4 u4_sll_454_U287 ( .A(u4_sll_454_ML_int_7__56_), .ZN(u4_sll_454_n55)
         );
  INV_X4 u4_sll_454_U286 ( .A(u4_sll_454_ML_int_7__57_), .ZN(u4_sll_454_n54)
         );
  INV_X4 u4_sll_454_U285 ( .A(u4_sll_454_ML_int_7__58_), .ZN(u4_sll_454_n53)
         );
  INV_X4 u4_sll_454_U284 ( .A(u4_sll_454_ML_int_7__59_), .ZN(u4_sll_454_n52)
         );
  INV_X4 u4_sll_454_U283 ( .A(u4_sll_454_ML_int_7__60_), .ZN(u4_sll_454_n51)
         );
  INV_X4 u4_sll_454_U282 ( .A(u4_sll_454_ML_int_7__61_), .ZN(u4_sll_454_n50)
         );
  INV_X4 u4_sll_454_U281 ( .A(u4_sll_454_ML_int_7__62_), .ZN(u4_sll_454_n49)
         );
  INV_X4 u4_sll_454_U280 ( .A(u4_sll_454_ML_int_7__63_), .ZN(u4_sll_454_n48)
         );
  INV_X4 u4_sll_454_U279 ( .A(u4_sll_454_ML_int_7__64_), .ZN(u4_sll_454_n47)
         );
  INV_X4 u4_sll_454_U278 ( .A(u4_sll_454_ML_int_7__65_), .ZN(u4_sll_454_n46)
         );
  INV_X4 u4_sll_454_U277 ( .A(u4_sll_454_ML_int_7__66_), .ZN(u4_sll_454_n45)
         );
  INV_X4 u4_sll_454_U276 ( .A(u4_sll_454_ML_int_7__67_), .ZN(u4_sll_454_n44)
         );
  INV_X4 u4_sll_454_U275 ( .A(u4_sll_454_ML_int_7__68_), .ZN(u4_sll_454_n43)
         );
  INV_X4 u4_sll_454_U274 ( .A(u4_sll_454_ML_int_7__69_), .ZN(u4_sll_454_n42)
         );
  INV_X4 u4_sll_454_U273 ( .A(u4_sll_454_ML_int_7__70_), .ZN(u4_sll_454_n41)
         );
  INV_X4 u4_sll_454_U272 ( .A(u4_sll_454_ML_int_7__71_), .ZN(u4_sll_454_n40)
         );
  INV_X4 u4_sll_454_U271 ( .A(u4_sll_454_ML_int_7__72_), .ZN(u4_sll_454_n39)
         );
  INV_X4 u4_sll_454_U270 ( .A(u4_sll_454_ML_int_7__73_), .ZN(u4_sll_454_n38)
         );
  INV_X4 u4_sll_454_U269 ( .A(u4_sll_454_ML_int_7__74_), .ZN(u4_sll_454_n37)
         );
  INV_X4 u4_sll_454_U268 ( .A(u4_sll_454_ML_int_7__75_), .ZN(u4_sll_454_n36)
         );
  INV_X4 u4_sll_454_U267 ( .A(u4_sll_454_ML_int_7__76_), .ZN(u4_sll_454_n35)
         );
  INV_X4 u4_sll_454_U266 ( .A(u4_sll_454_ML_int_7__77_), .ZN(u4_sll_454_n34)
         );
  INV_X4 u4_sll_454_U265 ( .A(u4_sll_454_ML_int_7__78_), .ZN(u4_sll_454_n33)
         );
  INV_X4 u4_sll_454_U264 ( .A(u4_sll_454_ML_int_7__79_), .ZN(u4_sll_454_n32)
         );
  INV_X4 u4_sll_454_U263 ( .A(u4_sll_454_ML_int_7__80_), .ZN(u4_sll_454_n31)
         );
  INV_X4 u4_sll_454_U262 ( .A(u4_sll_454_ML_int_7__81_), .ZN(u4_sll_454_n30)
         );
  INV_X4 u4_sll_454_U261 ( .A(u4_sll_454_ML_int_7__82_), .ZN(u4_sll_454_n29)
         );
  INV_X4 u4_sll_454_U260 ( .A(u4_sll_454_ML_int_7__83_), .ZN(u4_sll_454_n28)
         );
  INV_X4 u4_sll_454_U259 ( .A(u4_sll_454_ML_int_7__84_), .ZN(u4_sll_454_n27)
         );
  INV_X4 u4_sll_454_U258 ( .A(u4_sll_454_ML_int_7__85_), .ZN(u4_sll_454_n26)
         );
  INV_X4 u4_sll_454_U257 ( .A(u4_sll_454_ML_int_7__86_), .ZN(u4_sll_454_n25)
         );
  INV_X4 u4_sll_454_U256 ( .A(u4_sll_454_ML_int_7__87_), .ZN(u4_sll_454_n24)
         );
  INV_X4 u4_sll_454_U255 ( .A(u4_sll_454_ML_int_7__88_), .ZN(u4_sll_454_n23)
         );
  INV_X4 u4_sll_454_U254 ( .A(u4_sll_454_ML_int_7__89_), .ZN(u4_sll_454_n22)
         );
  INV_X4 u4_sll_454_U253 ( .A(u4_sll_454_ML_int_7__90_), .ZN(u4_sll_454_n21)
         );
  INV_X4 u4_sll_454_U252 ( .A(u4_sll_454_ML_int_7__91_), .ZN(u4_sll_454_n20)
         );
  INV_X4 u4_sll_454_U251 ( .A(u4_sll_454_ML_int_7__92_), .ZN(u4_sll_454_n19)
         );
  INV_X4 u4_sll_454_U250 ( .A(u4_sll_454_ML_int_7__93_), .ZN(u4_sll_454_n18)
         );
  INV_X4 u4_sll_454_U249 ( .A(u4_sll_454_ML_int_7__94_), .ZN(u4_sll_454_n17)
         );
  INV_X4 u4_sll_454_U248 ( .A(u4_sll_454_ML_int_7__95_), .ZN(u4_sll_454_n16)
         );
  INV_X4 u4_sll_454_U247 ( .A(u4_sll_454_ML_int_7__96_), .ZN(u4_sll_454_n15)
         );
  INV_X4 u4_sll_454_U246 ( .A(u4_sll_454_ML_int_7__97_), .ZN(u4_sll_454_n14)
         );
  INV_X4 u4_sll_454_U245 ( .A(u4_sll_454_ML_int_7__98_), .ZN(u4_sll_454_n13)
         );
  INV_X4 u4_sll_454_U244 ( .A(u4_sll_454_ML_int_7__99_), .ZN(u4_sll_454_n12)
         );
  INV_X4 u4_sll_454_U243 ( .A(u4_sll_454_ML_int_7__100_), .ZN(u4_sll_454_n11)
         );
  INV_X4 u4_sll_454_U242 ( .A(u4_sll_454_ML_int_7__101_), .ZN(u4_sll_454_n10)
         );
  INV_X4 u4_sll_454_U241 ( .A(u4_sll_454_ML_int_7__102_), .ZN(u4_sll_454_n9)
         );
  INV_X4 u4_sll_454_U240 ( .A(u4_sll_454_ML_int_7__103_), .ZN(u4_sll_454_n8)
         );
  INV_X4 u4_sll_454_U239 ( .A(u4_sll_454_ML_int_7__104_), .ZN(u4_sll_454_n7)
         );
  INV_X4 u4_sll_454_U238 ( .A(u4_sll_454_ML_int_7__105_), .ZN(u4_sll_454_n6)
         );
  OAI21_X1 u4_sll_454_U237 ( .B1(u4_shift_left[6]), .B2(u4_sll_454_net61032), 
        .A(u4_sll_454_net61030), .ZN(u4_sll_454_SHMAG_6_) );
  NOR2_X4 u4_sll_454_U236 ( .A1(u4_sll_454_net61028), .A2(u4_sll_454_n1), .ZN(
        u4_sll_454_temp_int_SH_0_) );
  INV_X8 u4_sll_454_U235 ( .A(u4_sll_454_temp_int_SH_0_), .ZN(
        u4_sll_454_net66387) );
  INV_X32 u4_sll_454_U234 ( .A(u4_sll_454_net66379), .ZN(u4_sll_454_net66361)
         );
  INV_X32 u4_sll_454_U233 ( .A(u4_sll_454_net66377), .ZN(u4_sll_454_net66359)
         );
  INV_X32 u4_sll_454_U232 ( .A(u4_sll_454_net66383), .ZN(u4_sll_454_net66379)
         );
  INV_X4 u4_sll_454_U231 ( .A(u4_shift_left[1]), .ZN(u4_sll_454_net61037) );
  NAND2_X2 u4_sll_454_U230 ( .A1(u4_sll_454_net63273), .A2(u4_sll_454_net61037), .ZN(u4_sll_454_n5) );
  NAND3_X1 u4_sll_454_U229 ( .A1(u4_sll_454_net61034), .A2(u4_sll_454_n5), 
        .A3(u4_sll_454_net61030), .ZN(u4_sll_454_SHMAG_1_) );
  OAI21_X1 u4_sll_454_U228 ( .B1(u4_shift_left[4]), .B2(u4_sll_454_net61032), 
        .A(u4_sll_454_net61030), .ZN(u4_sll_454_SHMAG_4_) );
  INV_X32 u4_sll_454_U227 ( .A(u4_sll_454_net66593), .ZN(u4_sll_454_net66591)
         );
  INV_X32 u4_sll_454_U226 ( .A(u4_sll_454_net66593), .ZN(u4_sll_454_net66589)
         );
  INV_X32 u4_sll_454_U225 ( .A(u4_sll_454_net66585), .ZN(u4_sll_454_net66563)
         );
  INV_X32 u4_sll_454_U224 ( .A(u4_sll_454_net66677), .ZN(u4_sll_454_net66659)
         );
  OAI21_X1 u4_sll_454_U223 ( .B1(u4_shift_left[3]), .B2(u4_sll_454_net61032), 
        .A(u4_sll_454_net61030), .ZN(u4_sll_454_SHMAG_3_) );
  INV_X32 u4_sll_454_U222 ( .A(u4_sll_454_net66621), .ZN(u4_sll_454_net66603)
         );
  INV_X32 u4_sll_454_U221 ( .A(u4_sll_454_net66621), .ZN(u4_sll_454_net66601)
         );
  INV_X32 u4_sll_454_U220 ( .A(u4_sll_454_net66621), .ZN(u4_sll_454_net66599)
         );
  OAI21_X1 u4_sll_454_U219 ( .B1(u4_shift_left[2]), .B2(u4_sll_454_net61032), 
        .A(u4_sll_454_net61030), .ZN(u4_sll_454_SHMAG_2_) );
  INV_X32 u4_sll_454_U218 ( .A(u4_sll_454_net66589), .ZN(u4_sll_454_net66585)
         );
  INV_X32 u4_sll_454_U217 ( .A(u4_sll_454_net66565), .ZN(u4_sll_454_net66545)
         );
  INV_X32 u4_sll_454_U216 ( .A(u4_sll_454_net66585), .ZN(u4_sll_454_net66565)
         );
  INV_X32 u4_sll_454_U215 ( .A(u4_sll_454_net66565), .ZN(u4_sll_454_net66547)
         );
  NOR2_X4 u4_sll_454_U214 ( .A1(u4_sll_454_net63267), .A2(
        u4_sll_454__UDW__90347_net74043), .ZN(u4_N6058) );
  INV_X32 u4_sll_454_U213 ( .A(u4_sll_454_net66455), .ZN(u4_sll_454_net66433)
         );
  INV_X32 u4_sll_454_U212 ( .A(u4_sll_454_net66455), .ZN(u4_sll_454_net66431)
         );
  INV_X32 u4_sll_454_U211 ( .A(u4_sll_454_net66451), .ZN(u4_sll_454_net66435)
         );
  INV_X32 u4_sll_454_U210 ( .A(u4_sll_454_n3), .ZN(u4_sll_454_net63277) );
  INV_X32 u4_sll_454_U209 ( .A(u4_sll_454_net63277), .ZN(u4_sll_454_net63271)
         );
  AOI21_X2 u4_sll_454_U208 ( .B1(u4_sll_454_n2), .B2(u4_sll_454_net63277), .A(
        u4_shift_left[0]), .ZN(u4_sll_454_net61028) );
  NAND2_X2 u4_sll_454_U207 ( .A1(u4_sll_454_n2), .A2(u4_sll_454_net63277), 
        .ZN(u4_sll_454_net61033) );
  INV_X4 u4_sll_454_U206 ( .A(u4_sll_454_net61033), .ZN(u4_sll_454_net61032)
         );
  OAI21_X1 u4_sll_454_U205 ( .B1(u4_shift_left[5]), .B2(u4_sll_454_net61032), 
        .A(u4_sll_454_net61030), .ZN(u4_sll_454_SHMAG_5_) );
  INV_X32 u4_sll_454_U204 ( .A(u4_sll_454_net66509), .ZN(u4_sll_454_net66489)
         );
  INV_X32 u4_sll_454_U203 ( .A(u4_sll_454_net66509), .ZN(u4_sll_454_net66487)
         );
  INV_X32 u4_sll_454_U202 ( .A(u4_sll_454_net66537), .ZN(u4_sll_454_net66509)
         );
  INV_X32 u4_sll_454_U201 ( .A(u4_sll_454_net66509), .ZN(u4_sll_454_net66491)
         );
  INV_X4 u4_sll_454_U200 ( .A(u4_sll_454_ML_int_6__44_), .ZN(
        u4_sll_454__UDW__90155_net73403) );
  NOR2_X4 u4_sll_454_U199 ( .A1(u4_sll_454_net66435), .A2(
        u4_sll_454__UDW__90155_net73403), .ZN(u4_sll_454_ML_int_7__44_) );
  INV_X8 u4_sll_454_U198 ( .A(u4_shift_left[7]), .ZN(u4_sll_454_net61036) );
  INV_X16 u4_sll_454_U197 ( .A(u4_sll_454_net66379), .ZN(u4_sll_454_net66373)
         );
  INV_X16 u4_sll_454_U196 ( .A(u4_sll_454_net66379), .ZN(u4_sll_454_net66363)
         );
  INV_X16 u4_sll_454_U195 ( .A(u4_sll_454_net66377), .ZN(u4_sll_454_net66365)
         );
  INV_X16 u4_sll_454_U194 ( .A(u4_sll_454_net66379), .ZN(u4_sll_454_net66367)
         );
  INV_X16 u4_sll_454_U193 ( .A(u4_sll_454_net66383), .ZN(u4_sll_454_net66377)
         );
  INV_X16 u4_sll_454_U192 ( .A(u4_sll_454_net66379), .ZN(u4_sll_454_net66369)
         );
  INV_X16 u4_sll_454_U191 ( .A(u4_sll_454_net66377), .ZN(u4_sll_454_net66371)
         );
  INV_X2 u4_sll_454_U190 ( .A(u4_sll_454_ML_int_6__33_), .ZN(u4_sll_454_n140)
         );
  INV_X8 u4_sll_454_U189 ( .A(u4_sll_454_net66387), .ZN(u4_sll_454_net66385)
         );
  NOR2_X2 u4_sll_454_U188 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n47), 
        .ZN(u4_N6078) );
  INV_X8 u4_sll_454_U187 ( .A(u4_shift_left[8]), .ZN(u4_sll_454_n4) );
  INV_X8 u4_sll_454_U186 ( .A(u4_sll_454_ML_int_7__44_), .ZN(
        u4_sll_454__UDW__90347_net74043) );
  INV_X16 u4_sll_454_U185 ( .A(u4_sll_454_n4), .ZN(u4_sll_454_n3) );
  INV_X4 u4_sll_454_U184 ( .A(u4_sll_454_net63277), .ZN(u4_sll_454_net63267)
         );
  INV_X4 u4_sll_454_U183 ( .A(u4_sll_454_net63277), .ZN(u4_sll_454_net63265)
         );
  INV_X8 u4_sll_454_U182 ( .A(u4_sll_454_n4), .ZN(u4_sll_454_net63261) );
  INV_X4 u4_sll_454_U181 ( .A(u4_sll_454_net63277), .ZN(u4_sll_454_net63269)
         );
  INV_X16 u4_sll_454_U180 ( .A(u4_sll_454_net66647), .ZN(u4_sll_454_net66613)
         );
  INV_X16 u4_sll_454_U179 ( .A(u4_sll_454_net66757), .ZN(u4_sll_454_net66719)
         );
  INV_X16 u4_sll_454_U178 ( .A(u4_sll_454_net66757), .ZN(u4_sll_454_net66717)
         );
  INV_X4 u4_sll_454_U177 ( .A(u4_sll_454_SHMAG_5_), .ZN(u4_sll_454_net66537)
         );
  INV_X4 u4_sll_454_U176 ( .A(u4_sll_454_net66705), .ZN(u4_sll_454_net66701)
         );
  INV_X2 u4_sll_454_U175 ( .A(u4_sll_454_SHMAG_2_), .ZN(u4_sll_454_net66705)
         );
  INV_X16 u4_sll_454_U174 ( .A(u4_sll_454_net66591), .ZN(u4_sll_454_net66555)
         );
  INV_X4 u4_sll_454_U173 ( .A(u4_sll_454_SHMAG_6_), .ZN(u4_sll_454_net66481)
         );
  INV_X8 u4_sll_454_U172 ( .A(u4_sll_454_net66675), .ZN(u4_sll_454_net66661)
         );
  INV_X16 u4_sll_454_U171 ( .A(u4_sll_454_net66701), .ZN(u4_sll_454_net66699)
         );
  INV_X16 u4_sll_454_U170 ( .A(u4_sll_454_net66481), .ZN(u4_sll_454_net66455)
         );
  INV_X16 u4_sll_454_U169 ( .A(u4_sll_454_net66481), .ZN(u4_sll_454_net66451)
         );
  INV_X16 u4_sll_454_U168 ( .A(u4_sll_454_net66757), .ZN(u4_sll_454_net66721)
         );
  INV_X4 u4_sll_454_U167 ( .A(u4_sll_454_SHMAG_1_), .ZN(u4_sll_454_net66761)
         );
  INV_X8 u4_sll_454_U166 ( .A(u4_sll_454_net66761), .ZN(u4_sll_454_net66757)
         );
  INV_X16 u4_sll_454_U165 ( .A(u4_sll_454_net66697), .ZN(u4_sll_454_net66677)
         );
  INV_X16 u4_sll_454_U164 ( .A(u4_sll_454_net66701), .ZN(u4_sll_454_net66697)
         );
  INV_X8 u4_sll_454_U163 ( .A(u4_sll_454_net66647), .ZN(u4_sll_454_net66611)
         );
  INV_X4 u4_sll_454_U162 ( .A(u4_sll_454_SHMAG_3_), .ZN(u4_sll_454_net66649)
         );
  INV_X16 u4_sll_454_U161 ( .A(u4_sll_454_net66733), .ZN(u4_sll_454_net66715)
         );
  INV_X16 u4_sll_454_U160 ( .A(u4_sll_454_net66733), .ZN(u4_sll_454_net66711)
         );
  INV_X4 u4_sll_454_U159 ( .A(u4_sll_454_net66761), .ZN(u4_sll_454_net66733)
         );
  NOR2_X2 u4_sll_454_U158 ( .A1(u4_sll_454_net63259), .A2(u4_sll_454_n19), 
        .ZN(u4_N6106) );
  NOR2_X2 u4_sll_454_U157 ( .A1(u4_sll_454_net63261), .A2(u4_sll_454_n21), 
        .ZN(u4_N6104) );
  NOR2_X2 u4_sll_454_U156 ( .A1(u4_sll_454_net63261), .A2(u4_sll_454_n22), 
        .ZN(u4_N6103) );
  NOR2_X2 u4_sll_454_U155 ( .A1(u4_sll_454_net63261), .A2(u4_sll_454_n23), 
        .ZN(u4_N6102) );
  NOR2_X2 u4_sll_454_U154 ( .A1(u4_sll_454_net63259), .A2(u4_sll_454_n16), 
        .ZN(u4_N6109) );
  NOR2_X2 u4_sll_454_U153 ( .A1(u4_sll_454_net63259), .A2(u4_sll_454_n15), 
        .ZN(u4_N6110) );
  NOR2_X2 u4_sll_454_U152 ( .A1(u4_sll_454_net63259), .A2(u4_sll_454_n14), 
        .ZN(u4_N6111) );
  NOR2_X2 u4_sll_454_U151 ( .A1(u4_sll_454_net63259), .A2(u4_sll_454_n13), 
        .ZN(u4_N6112) );
  NOR2_X2 u4_sll_454_U150 ( .A1(u4_sll_454_net63259), .A2(u4_sll_454_n18), 
        .ZN(u4_N6107) );
  NOR2_X2 u4_sll_454_U149 ( .A1(u4_sll_454_net63259), .A2(u4_sll_454_n17), 
        .ZN(u4_N6108) );
  NOR2_X2 u4_sll_454_U148 ( .A1(u4_sll_454_net66441), .A2(u4_sll_454_n117), 
        .ZN(u4_sll_454_ML_int_7__57_) );
  NOR2_X2 u4_sll_454_U147 ( .A1(u4_sll_454_net63265), .A2(u4_sll_454_n54), 
        .ZN(u4_N6071) );
  NOR2_X2 u4_sll_454_U146 ( .A1(u4_sll_454_net63259), .A2(u4_sll_454_n8), .ZN(
        u4_N6117) );
  NOR2_X2 u4_sll_454_U145 ( .A1(u4_sll_454_net66441), .A2(u4_sll_454_n116), 
        .ZN(u4_sll_454_ML_int_7__58_) );
  NOR2_X2 u4_sll_454_U144 ( .A1(u4_sll_454_net63265), .A2(u4_sll_454_n53), 
        .ZN(u4_N6072) );
  NOR2_X2 u4_sll_454_U143 ( .A1(u4_sll_454_net63259), .A2(u4_sll_454_n9), .ZN(
        u4_N6116) );
  NOR2_X2 u4_sll_454_U142 ( .A1(u4_sll_454_net63259), .A2(u4_sll_454_n12), 
        .ZN(u4_N6113) );
  NOR2_X2 u4_sll_454_U141 ( .A1(u4_sll_454_net63259), .A2(u4_sll_454_n10), 
        .ZN(u4_N6115) );
  NOR2_X2 u4_sll_454_U140 ( .A1(u4_sll_454_net63259), .A2(u4_sll_454_n11), 
        .ZN(u4_N6114) );
  NOR2_X2 u4_sll_454_U139 ( .A1(u4_sll_454_net66441), .A2(u4_sll_454_n114), 
        .ZN(u4_sll_454_ML_int_7__60_) );
  NOR2_X2 u4_sll_454_U138 ( .A1(u4_sll_454_net63265), .A2(u4_sll_454_n51), 
        .ZN(u4_N6074) );
  NOR2_X2 u4_sll_454_U137 ( .A1(u4_sll_454_net66441), .A2(u4_sll_454_n113), 
        .ZN(u4_sll_454_ML_int_7__61_) );
  NOR2_X2 u4_sll_454_U136 ( .A1(u4_sll_454_net63265), .A2(u4_sll_454_n50), 
        .ZN(u4_N6075) );
  NOR2_X2 u4_sll_454_U135 ( .A1(u4_sll_454_net66441), .A2(u4_sll_454_n112), 
        .ZN(u4_sll_454_ML_int_7__62_) );
  NOR2_X2 u4_sll_454_U134 ( .A1(u4_sll_454_net63265), .A2(u4_sll_454_n49), 
        .ZN(u4_N6076) );
  NOR2_X2 u4_sll_454_U133 ( .A1(u4_sll_454_net66441), .A2(u4_sll_454_n111), 
        .ZN(u4_sll_454_ML_int_7__63_) );
  NOR2_X2 u4_sll_454_U132 ( .A1(u4_sll_454_net63265), .A2(u4_sll_454_n48), 
        .ZN(u4_N6077) );
  NOR2_X2 u4_sll_454_U131 ( .A1(u4_sll_454_net63259), .A2(u4_sll_454_n7), .ZN(
        u4_N6118) );
  NOR2_X2 u4_sll_454_U130 ( .A1(u4_sll_454_net66441), .A2(u4_sll_454_n115), 
        .ZN(u4_sll_454_ML_int_7__59_) );
  NOR2_X2 u4_sll_454_U129 ( .A1(u4_sll_454_net63265), .A2(u4_sll_454_n52), 
        .ZN(u4_N6073) );
  NOR2_X2 u4_sll_454_U128 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n44), 
        .ZN(u4_N6081) );
  NOR2_X2 u4_sll_454_U127 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n43), 
        .ZN(u4_N6082) );
  NOR2_X2 u4_sll_454_U126 ( .A1(u4_sll_454_net66435), .A2(u4_sll_454_n120), 
        .ZN(u4_sll_454_ML_int_7__54_) );
  NOR2_X2 u4_sll_454_U125 ( .A1(u4_sll_454_net63265), .A2(u4_sll_454_n57), 
        .ZN(u4_N6068) );
  NOR2_X2 u4_sll_454_U124 ( .A1(u4_sll_454_net63261), .A2(u4_sll_454_n46), 
        .ZN(u4_N6079) );
  NOR2_X2 u4_sll_454_U123 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n39), 
        .ZN(u4_N6086) );
  NOR2_X2 u4_sll_454_U122 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n38), 
        .ZN(u4_N6087) );
  NOR2_X2 u4_sll_454_U121 ( .A1(u4_sll_454_net66441), .A2(u4_sll_454_n119), 
        .ZN(u4_sll_454_ML_int_7__55_) );
  NOR2_X2 u4_sll_454_U120 ( .A1(u4_sll_454_net63265), .A2(u4_sll_454_n56), 
        .ZN(u4_N6069) );
  NOR2_X2 u4_sll_454_U119 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n37), 
        .ZN(u4_N6088) );
  NOR2_X2 u4_sll_454_U118 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n42), 
        .ZN(u4_N6083) );
  NOR2_X2 u4_sll_454_U117 ( .A1(u4_sll_454_net63261), .A2(u4_sll_454_n40), 
        .ZN(u4_N6085) );
  NOR2_X2 u4_sll_454_U116 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n41), 
        .ZN(u4_N6084) );
  NOR2_X2 u4_sll_454_U115 ( .A1(u4_sll_454_net63261), .A2(u4_sll_454_n32), 
        .ZN(u4_N6093) );
  NOR2_X2 u4_sll_454_U114 ( .A1(u4_sll_454_net63261), .A2(u4_sll_454_n31), 
        .ZN(u4_N6094) );
  NOR2_X2 u4_sll_454_U113 ( .A1(u4_sll_454_net63261), .A2(u4_sll_454_n33), 
        .ZN(u4_N6092) );
  NOR2_X2 u4_sll_454_U112 ( .A1(u4_sll_454_net63261), .A2(u4_sll_454_n36), 
        .ZN(u4_N6089) );
  NOR2_X2 u4_sll_454_U111 ( .A1(u4_sll_454_net63261), .A2(u4_sll_454_n34), 
        .ZN(u4_N6091) );
  NOR2_X2 u4_sll_454_U110 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n35), 
        .ZN(u4_N6090) );
  NOR2_X2 u4_sll_454_U109 ( .A1(u4_sll_454_net66441), .A2(u4_sll_454_n118), 
        .ZN(u4_sll_454_ML_int_7__56_) );
  NOR2_X2 u4_sll_454_U108 ( .A1(u4_sll_454_net63265), .A2(u4_sll_454_n55), 
        .ZN(u4_N6070) );
  NOR2_X2 u4_sll_454_U107 ( .A1(u4_sll_454_net63261), .A2(u4_sll_454_n27), 
        .ZN(u4_N6098) );
  NOR2_X2 u4_sll_454_U106 ( .A1(u4_sll_454_net63261), .A2(u4_sll_454_n26), 
        .ZN(u4_N6099) );
  NOR2_X2 u4_sll_454_U105 ( .A1(u4_sll_454_net63261), .A2(u4_sll_454_n25), 
        .ZN(u4_N6100) );
  NOR2_X2 u4_sll_454_U104 ( .A1(u4_sll_454_net63261), .A2(u4_sll_454_n28), 
        .ZN(u4_N6097) );
  NOR2_X2 u4_sll_454_U103 ( .A1(u4_sll_454_net63261), .A2(u4_sll_454_n29), 
        .ZN(u4_N6096) );
  NOR2_X2 u4_sll_454_U102 ( .A1(u4_sll_454_net66435), .A2(u4_sll_454_n121), 
        .ZN(u4_sll_454_ML_int_7__53_) );
  NOR2_X2 u4_sll_454_U101 ( .A1(u4_sll_454_net63265), .A2(u4_sll_454_n58), 
        .ZN(u4_N6067) );
  NOR2_X2 u4_sll_454_U100 ( .A1(u4_sll_454_net63261), .A2(u4_sll_454_n30), 
        .ZN(u4_N6095) );
  NOR2_X2 u4_sll_454_U99 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n45), .ZN(
        u4_N6080) );
  NOR2_X2 u4_sll_454_U98 ( .A1(u4_sll_454_net63261), .A2(u4_sll_454_n20), .ZN(
        u4_N6105) );
  NOR2_X2 u4_sll_454_U97 ( .A1(u4_sll_454_net63261), .A2(u4_sll_454_n24), .ZN(
        u4_N6101) );
  NOR2_X2 u4_sll_454_U96 ( .A1(u4_sll_454_net63265), .A2(u4_sll_454_n6), .ZN(
        u4_N6119) );
  INV_X16 u4_sll_454_U95 ( .A(u4_sll_454_net66697), .ZN(u4_sll_454_net66675)
         );
  INV_X16 u4_sll_454_U94 ( .A(u4_sll_454_net66387), .ZN(u4_sll_454_net66383)
         );
  INV_X16 u4_sll_454_U93 ( .A(u4_sll_454_net66757), .ZN(u4_sll_454_net66727)
         );
  NOR2_X2 u4_sll_454_U92 ( .A1(u4_sll_454_net63271), .A2(u4_sll_454_n98), .ZN(
        u4_N6026) );
  NOR2_X2 u4_sll_454_U91 ( .A1(u4_sll_454_net66445), .A2(u4_sll_454_n166), 
        .ZN(u4_sll_454_ML_int_7__7_) );
  NOR2_X2 u4_sll_454_U90 ( .A1(u4_sll_454_net63273), .A2(u4_sll_454_n103), 
        .ZN(u4_N6021) );
  NOR2_X2 u4_sll_454_U89 ( .A1(u4_sll_454_net66445), .A2(u4_sll_454_n165), 
        .ZN(u4_sll_454_ML_int_7__8_) );
  NOR2_X2 u4_sll_454_U88 ( .A1(u4_sll_454_net63273), .A2(u4_sll_454_n102), 
        .ZN(u4_N6022) );
  NOR2_X2 u4_sll_454_U87 ( .A1(u4_sll_454_net66429), .A2(u4_sll_454_n160), 
        .ZN(u4_sll_454_ML_int_7__13_) );
  NOR2_X2 u4_sll_454_U86 ( .A1(u4_sll_454_net63271), .A2(u4_sll_454_n97), .ZN(
        u4_N6027) );
  NOR2_X2 u4_sll_454_U85 ( .A1(u4_sll_454_net66445), .A2(u4_sll_454_n163), 
        .ZN(u4_sll_454_ML_int_7__10_) );
  NOR2_X2 u4_sll_454_U84 ( .A1(u4_sll_454_net63271), .A2(u4_sll_454_n100), 
        .ZN(u4_N6024) );
  NOR2_X2 u4_sll_454_U83 ( .A1(u4_sll_454_net66445), .A2(u4_sll_454_n164), 
        .ZN(u4_sll_454_ML_int_7__9_) );
  NOR2_X2 u4_sll_454_U82 ( .A1(u4_sll_454_net66429), .A2(u4_sll_454_n154), 
        .ZN(u4_sll_454_ML_int_7__19_) );
  NOR2_X2 u4_sll_454_U81 ( .A1(u4_sll_454_net66431), .A2(u4_sll_454_n150), 
        .ZN(u4_sll_454_ML_int_7__23_) );
  NOR2_X2 u4_sll_454_U80 ( .A1(u4_sll_454_net66431), .A2(u4_sll_454_n151), 
        .ZN(u4_sll_454_ML_int_7__22_) );
  NOR2_X2 u4_sll_454_U79 ( .A1(u4_sll_454_net66429), .A2(u4_sll_454_n159), 
        .ZN(u4_sll_454_ML_int_7__14_) );
  NOR2_X2 u4_sll_454_U78 ( .A1(u4_sll_454_net63271), .A2(u4_sll_454_n96), .ZN(
        u4_N6028) );
  NOR2_X2 u4_sll_454_U77 ( .A1(u4_sll_454_net66429), .A2(u4_sll_454_n156), 
        .ZN(u4_sll_454_ML_int_7__17_) );
  NOR2_X2 u4_sll_454_U76 ( .A1(u4_sll_454_net63271), .A2(u4_sll_454_n93), .ZN(
        u4_N6031) );
  NOR2_X2 u4_sll_454_U75 ( .A1(u4_sll_454_net66429), .A2(u4_sll_454_n158), 
        .ZN(u4_sll_454_ML_int_7__15_) );
  NOR2_X2 u4_sll_454_U74 ( .A1(u4_sll_454_net63271), .A2(u4_sll_454_n95), .ZN(
        u4_N6029) );
  NOR2_X2 u4_sll_454_U73 ( .A1(u4_sll_454_net66429), .A2(u4_sll_454_n157), 
        .ZN(u4_sll_454_ML_int_7__16_) );
  NOR2_X2 u4_sll_454_U72 ( .A1(u4_sll_454_net63271), .A2(u4_sll_454_n94), .ZN(
        u4_N6030) );
  NOR2_X2 u4_sll_454_U71 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n82), .ZN(
        u4_N6042) );
  NOR2_X2 u4_sll_454_U70 ( .A1(u4_sll_454_net66433), .A2(u4_sll_454_n140), 
        .ZN(u4_sll_454_ML_int_7__33_) );
  NOR2_X2 u4_sll_454_U69 ( .A1(u4_sll_454_net66431), .A2(u4_sll_454_n147), 
        .ZN(u4_sll_454_ML_int_7__26_) );
  NOR2_X2 u4_sll_454_U68 ( .A1(u4_sll_454_net66431), .A2(u4_sll_454_n149), 
        .ZN(u4_sll_454_ML_int_7__24_) );
  NOR2_X2 u4_sll_454_U67 ( .A1(u4_sll_454_net66431), .A2(u4_sll_454_n148), 
        .ZN(u4_sll_454_ML_int_7__25_) );
  NOR2_X2 u4_sll_454_U66 ( .A1(u4_sll_454_net66431), .A2(u4_sll_454_n142), 
        .ZN(u4_sll_454_ML_int_7__31_) );
  NOR2_X2 u4_sll_454_U65 ( .A1(u4_sll_454_net66431), .A2(u4_sll_454_n141), 
        .ZN(u4_sll_454_ML_int_7__32_) );
  NOR2_X2 u4_sll_454_U64 ( .A1(u4_sll_454_net66433), .A2(u4_sll_454_n133), 
        .ZN(u4_sll_454_ML_int_7__40_) );
  NOR2_X2 u4_sll_454_U63 ( .A1(u4_sll_454_net66433), .A2(u4_sll_454_n132), 
        .ZN(u4_sll_454_ML_int_7__41_) );
  NOR2_X2 u4_sll_454_U62 ( .A1(u4_sll_454_net63267), .A2(u4_sll_454_n69), .ZN(
        u4_N6055) );
  NOR2_X2 u4_sll_454_U61 ( .A1(u4_sll_454_net66433), .A2(u4_sll_454_n130), 
        .ZN(u4_sll_454_ML_int_7__43_) );
  NOR2_X2 u4_sll_454_U60 ( .A1(u4_sll_454_net63267), .A2(u4_sll_454_n67), .ZN(
        u4_N6057) );
  INV_X4 u4_sll_454_U59 ( .A(u4_sll_454_net66649), .ZN(u4_sll_454_net66647) );
  NOR2_X2 u4_sll_454_U58 ( .A1(u4_sll_454_net66611), .A2(u4_sll_454_n226), 
        .ZN(u4_sll_454_ML_int_4__0_) );
  NOR2_X2 u4_sll_454_U57 ( .A1(u4_sll_454_net66611), .A2(u4_sll_454_n225), 
        .ZN(u4_sll_454_ML_int_4__1_) );
  INV_X16 u4_sll_454_U56 ( .A(u4_sll_454_net66611), .ZN(u4_sll_454_net66619)
         );
  INV_X16 u4_sll_454_U55 ( .A(u4_sll_454_net66649), .ZN(u4_sll_454_net66621)
         );
  INV_X16 u4_sll_454_U54 ( .A(u4_sll_454_net66677), .ZN(u4_sll_454_net66655)
         );
  NOR2_X2 u4_sll_454_U53 ( .A1(u4_sll_454_net63273), .A2(u4_sll_454_n106), 
        .ZN(u4_N6018) );
  NOR2_X2 u4_sll_454_U52 ( .A1(u4_sll_454_net63273), .A2(u4_sll_454_n105), 
        .ZN(u4_N6019) );
  NOR2_X2 u4_sll_454_U51 ( .A1(u4_sll_454_net66429), .A2(u4_sll_454_n171), 
        .ZN(u4_sll_454_ML_int_7__2_) );
  NOR2_X2 u4_sll_454_U50 ( .A1(u4_sll_454_net63273), .A2(u4_sll_454_n108), 
        .ZN(u4_N6016) );
  NOR2_X2 u4_sll_454_U49 ( .A1(u4_sll_454_net66429), .A2(u4_sll_454_n170), 
        .ZN(u4_sll_454_ML_int_7__3_) );
  NOR2_X2 u4_sll_454_U48 ( .A1(u4_sll_454_net63273), .A2(u4_sll_454_n107), 
        .ZN(u4_N6017) );
  NOR2_X2 u4_sll_454_U47 ( .A1(u4_sll_454_net66429), .A2(u4_sll_454_n167), 
        .ZN(u4_sll_454_ML_int_7__6_) );
  NOR2_X2 u4_sll_454_U46 ( .A1(u4_sll_454_net63273), .A2(u4_sll_454_n104), 
        .ZN(u4_N6020) );
  NOR2_X2 u4_sll_454_U45 ( .A1(u4_sll_454_net66429), .A2(u4_sll_454_n161), 
        .ZN(u4_sll_454_ML_int_7__12_) );
  NOR2_X2 u4_sll_454_U44 ( .A1(u4_sll_454_net66433), .A2(u4_sll_454_n136), 
        .ZN(u4_sll_454_ML_int_7__37_) );
  NOR2_X2 u4_sll_454_U43 ( .A1(u4_sll_454_net63267), .A2(u4_sll_454_n73), .ZN(
        u4_N6051) );
  NOR2_X2 u4_sll_454_U42 ( .A1(u4_sll_454_net66433), .A2(u4_sll_454_n135), 
        .ZN(u4_sll_454_ML_int_7__38_) );
  NOR2_X2 u4_sll_454_U41 ( .A1(u4_sll_454_net63267), .A2(u4_sll_454_n72), .ZN(
        u4_N6052) );
  NOR2_X2 u4_sll_454_U40 ( .A1(u4_sll_454_net66433), .A2(u4_sll_454_n134), 
        .ZN(u4_sll_454_ML_int_7__39_) );
  NOR2_X2 u4_sll_454_U39 ( .A1(u4_sll_454_net63267), .A2(u4_sll_454_n71), .ZN(
        u4_N6053) );
  NOR2_X2 u4_sll_454_U38 ( .A1(u4_sll_454_net66433), .A2(u4_sll_454_n139), 
        .ZN(u4_sll_454_ML_int_7__34_) );
  NOR2_X2 u4_sll_454_U37 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n76), .ZN(
        u4_N6048) );
  NOR2_X2 u4_sll_454_U36 ( .A1(u4_sll_454_net66433), .A2(u4_sll_454_n138), 
        .ZN(u4_sll_454_ML_int_7__35_) );
  NOR2_X2 u4_sll_454_U35 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n75), .ZN(
        u4_N6049) );
  NOR2_X2 u4_sll_454_U34 ( .A1(u4_sll_454_net66433), .A2(u4_sll_454_n137), 
        .ZN(u4_sll_454_ML_int_7__36_) );
  NOR2_X2 u4_sll_454_U33 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n74), .ZN(
        u4_N6050) );
  NOR2_X2 u4_sll_454_U32 ( .A1(u4_sll_454_net66431), .A2(u4_sll_454_n146), 
        .ZN(u4_sll_454_ML_int_7__27_) );
  NOR2_X2 u4_sll_454_U31 ( .A1(u4_sll_454_net66431), .A2(u4_sll_454_n143), 
        .ZN(u4_sll_454_ML_int_7__30_) );
  NOR2_X2 u4_sll_454_U30 ( .A1(u4_sll_454_net63269), .A2(u4_sll_454_n80), .ZN(
        u4_N6044) );
  NOR2_X2 u4_sll_454_U29 ( .A1(u4_sll_454_net66431), .A2(u4_sll_454_n144), 
        .ZN(u4_sll_454_ML_int_7__29_) );
  NOR2_X2 u4_sll_454_U28 ( .A1(u4_sll_454_net66431), .A2(u4_sll_454_n145), 
        .ZN(u4_sll_454_ML_int_7__28_) );
  NOR2_X2 u4_sll_454_U27 ( .A1(u4_sll_454_net66435), .A2(u4_sll_454_n124), 
        .ZN(u4_sll_454_ML_int_7__50_) );
  NOR2_X2 u4_sll_454_U26 ( .A1(u4_sll_454_net63267), .A2(u4_sll_454_n61), .ZN(
        u4_N6064) );
  NOR2_X2 u4_sll_454_U25 ( .A1(u4_sll_454_net66435), .A2(u4_sll_454_n123), 
        .ZN(u4_sll_454_ML_int_7__51_) );
  NOR2_X2 u4_sll_454_U24 ( .A1(u4_sll_454_net63265), .A2(u4_sll_454_n60), .ZN(
        u4_N6065) );
  NOR2_X2 u4_sll_454_U23 ( .A1(u4_sll_454_net66435), .A2(u4_sll_454_n122), 
        .ZN(u4_sll_454_ML_int_7__52_) );
  NOR2_X2 u4_sll_454_U22 ( .A1(u4_sll_454_net63265), .A2(u4_sll_454_n59), .ZN(
        u4_N6066) );
  NOR2_X2 u4_sll_454_U21 ( .A1(u4_sll_454_net66435), .A2(u4_sll_454_n127), 
        .ZN(u4_sll_454_ML_int_7__47_) );
  NOR2_X2 u4_sll_454_U20 ( .A1(u4_sll_454_net63267), .A2(u4_sll_454_n64), .ZN(
        u4_N6061) );
  NOR2_X2 u4_sll_454_U19 ( .A1(u4_sll_454_net66667), .A2(u4_sll_454_n230), 
        .ZN(u4_sll_454_ML_int_3__0_) );
  NOR2_X2 u4_sll_454_U18 ( .A1(u4_sll_454_net66727), .A2(u4_sll_454_n231), 
        .ZN(u4_sll_454_ML_int_2__1_) );
  NOR2_X2 u4_sll_454_U17 ( .A1(u4_sll_454_net66727), .A2(u4_sll_454_n232), 
        .ZN(u4_sll_454_ML_int_2__0_) );
  NOR2_X2 u4_sll_454_U16 ( .A1(u4_sll_454_net66429), .A2(u4_sll_454_n169), 
        .ZN(u4_sll_454_ML_int_7__4_) );
  NOR2_X2 u4_sll_454_U15 ( .A1(u4_sll_454_net66429), .A2(u4_sll_454_n168), 
        .ZN(u4_sll_454_ML_int_7__5_) );
  NOR2_X2 u4_sll_454_U14 ( .A1(u4_sll_454_net66435), .A2(u4_sll_454_n126), 
        .ZN(u4_sll_454_ML_int_7__48_) );
  NOR2_X2 u4_sll_454_U13 ( .A1(u4_sll_454_net63267), .A2(u4_sll_454_n63), .ZN(
        u4_N6062) );
  NOR2_X2 u4_sll_454_U12 ( .A1(u4_sll_454_net66435), .A2(u4_sll_454_n125), 
        .ZN(u4_sll_454_ML_int_7__49_) );
  NOR2_X2 u4_sll_454_U11 ( .A1(u4_sll_454_net63267), .A2(u4_sll_454_n62), .ZN(
        u4_N6063) );
  INV_X4 u4_sll_454_U10 ( .A(u4_sll_454_SHMAG_4_), .ZN(u4_sll_454_net66593) );
  MUX2_X2 u4_sll_454_U9 ( .A(u4_sll_454_ML_int_4__28_), .B(
        u4_sll_454_ML_int_4__44_), .S(u4_sll_454_net66565), .Z(
        u4_sll_454_ML_int_5__44_) );
  INV_X16 u4_sll_454_U8 ( .A(u4_sll_454_net63277), .ZN(u4_sll_454_net63273) );
  INV_X4 u4_sll_454_U7 ( .A(u4_sll_454_n1), .ZN(u4_sll_454_net61030) );
  NOR2_X4 u4_sll_454_U6 ( .A1(u4_shift_left[7]), .A2(u4_sll_454_net63277), 
        .ZN(u4_sll_454_n1) );
  INV_X16 u4_sll_454_U5 ( .A(u4_sll_454_net66379), .ZN(u4_sll_454_net66357) );
  NAND2_X2 u4_sll_454_U4 ( .A1(u4_sll_454_net61036), .A2(u4_sll_454_net61037), 
        .ZN(u4_sll_454_net61034) );
  INV_X4 u4_sll_454_U3 ( .A(u4_sll_454_net61036), .ZN(u4_sll_454_n2) );
  MUX2_X2 u4_sll_454_M1_5_44 ( .A(u4_sll_454_ML_int_5__44_), .B(
        u4_sll_454_ML_int_5__12_), .S(u4_sll_454_net66491), .Z(
        u4_sll_454_ML_int_6__44_) );
  MUX2_X2 u4_sll_454_M1_5_76 ( .A(u4_sll_454_ML_int_5__76_), .B(
        u4_sll_454_ML_int_5__44_), .S(u4_sll_454_net66495), .Z(
        u4_sll_454_ML_int_6__76_) );
  MUX2_X2 u4_sll_454_M1_2_20 ( .A(u4_sll_454_ML_int_2__20_), .B(
        u4_sll_454_ML_int_2__16_), .S(u4_sll_454_net66699), .Z(
        u4_sll_454_ML_int_3__20_) );
  MUX2_X2 u4_sll_454_M1_3_20 ( .A(u4_sll_454_ML_int_3__20_), .B(
        u4_sll_454_ML_int_3__12_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__20_) );
  MUX2_X2 u4_sll_454_M1_3_28 ( .A(u4_sll_454_ML_int_3__28_), .B(
        u4_sll_454_ML_int_3__20_), .S(u4_sll_454_net66599), .Z(
        u4_sll_454_ML_int_4__28_) );
  MUX2_X2 u4_sll_454_M1_1_20 ( .A(u4_sll_454_ML_int_1__20_), .B(
        u4_sll_454_ML_int_1__18_), .S(u4_sll_454_net66717), .Z(
        u4_sll_454_ML_int_2__20_) );
  MUX2_X2 u4_sll_454_M1_2_24 ( .A(u4_sll_454_ML_int_2__24_), .B(
        u4_sll_454_ML_int_2__20_), .S(u4_sll_454_net66655), .Z(
        u4_sll_454_ML_int_3__24_) );
  MUX2_X2 u4_sll_454_M1_4_28 ( .A(u4_sll_454_ML_int_4__28_), .B(
        u4_sll_454_ML_int_4__12_), .S(u4_sll_454_net66555), .Z(
        u4_sll_454_ML_int_5__28_) );
  MUX2_X2 u4_sll_454_M1_2_28 ( .A(u4_sll_454_ML_int_2__28_), .B(
        u4_sll_454_ML_int_2__24_), .S(u4_sll_454_net66655), .Z(
        u4_sll_454_ML_int_3__28_) );
  MUX2_X2 u4_sll_454_M1_3_36 ( .A(u4_sll_454_ML_int_3__36_), .B(
        u4_sll_454_ML_int_3__28_), .S(u4_sll_454_net66601), .Z(
        u4_sll_454_ML_int_4__36_) );
  MUX2_X2 u4_sll_454_M1_3_44 ( .A(u4_sll_454_ML_int_3__44_), .B(
        u4_sll_454_ML_int_3__36_), .S(u4_sll_454_net66603), .Z(
        u4_sll_454_ML_int_4__44_) );
  MUX2_X2 u4_sll_454_M1_4_60 ( .A(u4_sll_454_ML_int_4__60_), .B(
        u4_sll_454_ML_int_4__44_), .S(u4_sll_454_net66549), .Z(
        u4_sll_454_ML_int_5__60_) );
  MUX2_X2 u4_sll_454_M1_1_16 ( .A(u4_sll_454_ML_int_1__16_), .B(
        u4_sll_454_ML_int_1__14_), .S(u4_sll_454_net66721), .Z(
        u4_sll_454_ML_int_2__16_) );
  MUX2_X2 u4_sll_454_M1_2_16 ( .A(u4_sll_454_ML_int_2__16_), .B(
        u4_sll_454_ML_int_2__12_), .S(u4_sll_454_net66699), .Z(
        u4_sll_454_ML_int_3__16_) );
  MUX2_X2 u4_sll_454_M1_0_16 ( .A(n8516), .B(n8517), .S(u4_sll_454_net66357), 
        .Z(u4_sll_454_ML_int_1__16_) );
  MUX2_X2 u4_sll_454_M1_1_18 ( .A(u4_sll_454_ML_int_1__18_), .B(
        u4_sll_454_ML_int_1__16_), .S(u4_sll_454_net66721), .Z(
        u4_sll_454_ML_int_2__18_) );
  MUX2_X2 u4_sll_454_M1_0_14 ( .A(net33577), .B(net33578), .S(
        u4_sll_454_net66357), .Z(u4_sll_454_ML_int_1__14_) );
  MUX2_X2 u4_sll_454_M1_1_14 ( .A(u4_sll_454_ML_int_1__14_), .B(
        u4_sll_454_ML_int_1__12_), .S(u4_sll_454_net66721), .Z(
        u4_sll_454_ML_int_2__14_) );
  MUX2_X2 u4_sll_454_M1_0_15 ( .A(n8517), .B(net33577), .S(u4_sll_454_net66357), .Z(u4_sll_454_ML_int_1__15_) );
  MUX2_X2 u4_sll_454_M1_0_13 ( .A(net33578), .B(net33579), .S(
        u4_sll_454_net66357), .Z(u4_sll_454_ML_int_1__13_) );
  MUX2_X2 u4_sll_454_M1_0_1 ( .A(net33648), .B(net33546), .S(
        u4_sll_454_net66369), .Z(u4_sll_454_ML_int_1__1_) );
  MUX2_X2 u4_sll_454_M1_0_2 ( .A(net33647), .B(net33648), .S(
        u4_sll_454_net66385), .Z(u4_sll_454_ML_int_1__2_) );
  MUX2_X2 u4_sll_454_M1_0_3 ( .A(n8511), .B(net33647), .S(u4_sll_454_net66385), 
        .Z(u4_sll_454_ML_int_1__3_) );
  MUX2_X2 u4_sll_454_M1_0_4 ( .A(n8512), .B(n8511), .S(u4_sll_454_net66385), 
        .Z(u4_sll_454_ML_int_1__4_) );
  MUX2_X2 u4_sll_454_M1_0_5 ( .A(n8513), .B(n8512), .S(u4_sll_454_net66385), 
        .Z(u4_sll_454_ML_int_1__5_) );
  MUX2_X2 u4_sll_454_M1_0_6 ( .A(n8514), .B(n8513), .S(u4_sll_454_net66385), 
        .Z(u4_sll_454_ML_int_1__6_) );
  MUX2_X2 u4_sll_454_M1_0_7 ( .A(net33642), .B(n8514), .S(u4_sll_454_net66385), 
        .Z(u4_sll_454_ML_int_1__7_) );
  MUX2_X2 u4_sll_454_M1_0_8 ( .A(net33641), .B(net33642), .S(
        u4_sll_454_net66385), .Z(u4_sll_454_ML_int_1__8_) );
  MUX2_X2 u4_sll_454_M1_0_9 ( .A(net33548), .B(net33641), .S(
        u4_sll_454_net66385), .Z(u4_sll_454_ML_int_1__9_) );
  MUX2_X2 u4_sll_454_M1_0_10 ( .A(net33549), .B(net33548), .S(
        u4_sll_454_net66385), .Z(u4_sll_454_ML_int_1__10_) );
  MUX2_X2 u4_sll_454_M1_0_11 ( .A(net33581), .B(net33549), .S(
        u4_sll_454_net66357), .Z(u4_sll_454_ML_int_1__11_) );
  MUX2_X2 u4_sll_454_M1_0_12 ( .A(net33579), .B(net33581), .S(
        u4_sll_454_net66357), .Z(u4_sll_454_ML_int_1__12_) );
  MUX2_X2 u4_sll_454_M1_0_17 ( .A(net33575), .B(n8516), .S(u4_sll_454_net66357), .Z(u4_sll_454_ML_int_1__17_) );
  MUX2_X2 u4_sll_454_M1_0_18 ( .A(net33550), .B(net33575), .S(
        u4_sll_454_net66357), .Z(u4_sll_454_ML_int_1__18_) );
  MUX2_X2 u4_sll_454_M1_0_19 ( .A(net33573), .B(net33550), .S(
        u4_sll_454_net66357), .Z(u4_sll_454_ML_int_1__19_) );
  MUX2_X2 u4_sll_454_M1_0_20 ( .A(net33572), .B(net33573), .S(
        u4_sll_454_net66357), .Z(u4_sll_454_ML_int_1__20_) );
  MUX2_X2 u4_sll_454_M1_0_21 ( .A(n8518), .B(net33572), .S(u4_sll_454_net66357), .Z(u4_sll_454_ML_int_1__21_) );
  MUX2_X2 u4_sll_454_M1_0_22 ( .A(n8519), .B(n8518), .S(u4_sll_454_net66359), 
        .Z(u4_sll_454_ML_int_1__22_) );
  MUX2_X2 u4_sll_454_M1_0_23 ( .A(n8520), .B(n8519), .S(u4_sll_454_net66359), 
        .Z(u4_sll_454_ML_int_1__23_) );
  MUX2_X2 u4_sll_454_M1_0_24 ( .A(net33569), .B(n8520), .S(u4_sll_454_net66359), .Z(u4_sll_454_ML_int_1__24_) );
  MUX2_X2 u4_sll_454_M1_0_25 ( .A(net33568), .B(net33569), .S(
        u4_sll_454_net66359), .Z(u4_sll_454_ML_int_1__25_) );
  MUX2_X2 u4_sll_454_M1_0_26 ( .A(net33551), .B(net33568), .S(
        u4_sll_454_net66359), .Z(u4_sll_454_ML_int_1__26_) );
  MUX2_X2 u4_sll_454_M1_0_27 ( .A(net33566), .B(net33551), .S(
        u4_sll_454_net66359), .Z(u4_sll_454_ML_int_1__27_) );
  MUX2_X2 u4_sll_454_M1_0_28 ( .A(net33565), .B(net33566), .S(
        u4_sll_454_net66359), .Z(u4_sll_454_ML_int_1__28_) );
  MUX2_X2 u4_sll_454_M1_0_29 ( .A(net33564), .B(net33565), .S(
        u4_sll_454_net66359), .Z(u4_sll_454_ML_int_1__29_) );
  MUX2_X2 u4_sll_454_M1_0_30 ( .A(net33563), .B(net33564), .S(
        u4_sll_454_net66359), .Z(u4_sll_454_ML_int_1__30_) );
  MUX2_X2 u4_sll_454_M1_0_31 ( .A(n8521), .B(net33563), .S(u4_sll_454_net66359), .Z(u4_sll_454_ML_int_1__31_) );
  MUX2_X2 u4_sll_454_M1_0_32 ( .A(net33562), .B(n8521), .S(u4_sll_454_net66359), .Z(u4_sll_454_ML_int_1__32_) );
  MUX2_X2 u4_sll_454_M1_0_33 ( .A(net33561), .B(net33562), .S(
        u4_sll_454_net66361), .Z(u4_sll_454_ML_int_1__33_) );
  MUX2_X2 u4_sll_454_M1_0_34 ( .A(net33552), .B(net33561), .S(
        u4_sll_454_net66361), .Z(u4_sll_454_ML_int_1__34_) );
  MUX2_X2 u4_sll_454_M1_0_35 ( .A(net33559), .B(net33552), .S(
        u4_sll_454_net66361), .Z(u4_sll_454_ML_int_1__35_) );
  MUX2_X2 u4_sll_454_M1_0_36 ( .A(net33558), .B(net33559), .S(
        u4_sll_454_net66361), .Z(u4_sll_454_ML_int_1__36_) );
  MUX2_X2 u4_sll_454_M1_0_37 ( .A(n8522), .B(net33558), .S(u4_sll_454_net66361), .Z(u4_sll_454_ML_int_1__37_) );
  MUX2_X2 u4_sll_454_M1_0_38 ( .A(n8523), .B(n8522), .S(u4_sll_454_net66361), 
        .Z(u4_sll_454_ML_int_1__38_) );
  MUX2_X2 u4_sll_454_M1_0_39 ( .A(n8525), .B(n8523), .S(u4_sll_454_net66361), 
        .Z(u4_sll_454_ML_int_1__39_) );
  MUX2_X2 u4_sll_454_M1_0_40 ( .A(n8524), .B(n8525), .S(u4_sll_454_net66361), 
        .Z(u4_sll_454_ML_int_1__40_) );
  MUX2_X2 u4_sll_454_M1_0_41 ( .A(net33554), .B(n8524), .S(u4_sll_454_net66361), .Z(u4_sll_454_ML_int_1__41_) );
  MUX2_X2 u4_sll_454_M1_0_42 ( .A(net33547), .B(net33554), .S(
        u4_sll_454_net66361), .Z(u4_sll_454_ML_int_1__42_) );
  MUX2_X2 u4_sll_454_M1_0_43 ( .A(net33587), .B(net33547), .S(
        u4_sll_454_net66361), .Z(u4_sll_454_ML_int_1__43_) );
  MUX2_X2 u4_sll_454_M1_0_44 ( .A(net33586), .B(net33587), .S(
        u4_sll_454_net66363), .Z(u4_sll_454_ML_int_1__44_) );
  MUX2_X2 u4_sll_454_M1_0_45 ( .A(net33585), .B(net33586), .S(
        u4_sll_454_net66363), .Z(u4_sll_454_ML_int_1__45_) );
  MUX2_X2 u4_sll_454_M1_0_46 ( .A(net33584), .B(net33585), .S(
        u4_sll_454_net66363), .Z(u4_sll_454_ML_int_1__46_) );
  MUX2_X2 u4_sll_454_M1_0_47 ( .A(n8515), .B(net33584), .S(u4_sll_454_net66363), .Z(u4_sll_454_ML_int_1__47_) );
  MUX2_X2 u4_sll_454_M1_0_48 ( .A(net33583), .B(n8515), .S(u4_sll_454_net66363), .Z(u4_sll_454_ML_int_1__48_) );
  MUX2_X2 u4_sll_454_M1_0_49 ( .A(net33625), .B(net33583), .S(
        u4_sll_454_net66363), .Z(u4_sll_454_ML_int_1__49_) );
  MUX2_X2 u4_sll_454_M1_0_50 ( .A(fract_denorm[50]), .B(net33625), .S(
        u4_sll_454_net66363), .Z(u4_sll_454_ML_int_1__50_) );
  MUX2_X2 u4_sll_454_M1_0_51 ( .A(fract_denorm[51]), .B(fract_denorm[50]), .S(
        u4_sll_454_net66363), .Z(u4_sll_454_ML_int_1__51_) );
  MUX2_X2 u4_sll_454_M1_0_52 ( .A(fract_denorm[52]), .B(fract_denorm[51]), .S(
        u4_sll_454_net66363), .Z(u4_sll_454_ML_int_1__52_) );
  MUX2_X2 u4_sll_454_M1_0_53 ( .A(fract_denorm[53]), .B(fract_denorm[52]), .S(
        u4_sll_454_net66363), .Z(u4_sll_454_ML_int_1__53_) );
  MUX2_X2 u4_sll_454_M1_0_54 ( .A(fract_denorm[54]), .B(fract_denorm[53]), .S(
        u4_sll_454_net66363), .Z(u4_sll_454_ML_int_1__54_) );
  MUX2_X2 u4_sll_454_M1_0_55 ( .A(fract_denorm[55]), .B(fract_denorm[54]), .S(
        u4_sll_454_net66365), .Z(u4_sll_454_ML_int_1__55_) );
  MUX2_X2 u4_sll_454_M1_0_56 ( .A(fract_denorm[56]), .B(fract_denorm[55]), .S(
        u4_sll_454_net66365), .Z(u4_sll_454_ML_int_1__56_) );
  MUX2_X2 u4_sll_454_M1_0_57 ( .A(fract_denorm[57]), .B(fract_denorm[56]), .S(
        u4_sll_454_net66365), .Z(u4_sll_454_ML_int_1__57_) );
  MUX2_X2 u4_sll_454_M1_0_58 ( .A(fract_denorm[58]), .B(fract_denorm[57]), .S(
        u4_sll_454_net66365), .Z(u4_sll_454_ML_int_1__58_) );
  MUX2_X2 u4_sll_454_M1_0_59 ( .A(fract_denorm[59]), .B(fract_denorm[58]), .S(
        u4_sll_454_net66365), .Z(u4_sll_454_ML_int_1__59_) );
  MUX2_X2 u4_sll_454_M1_0_60 ( .A(fract_denorm[60]), .B(fract_denorm[59]), .S(
        u4_sll_454_net66365), .Z(u4_sll_454_ML_int_1__60_) );
  MUX2_X2 u4_sll_454_M1_0_61 ( .A(fract_denorm[61]), .B(fract_denorm[60]), .S(
        u4_sll_454_net66365), .Z(u4_sll_454_ML_int_1__61_) );
  MUX2_X2 u4_sll_454_M1_0_62 ( .A(fract_denorm[62]), .B(fract_denorm[61]), .S(
        u4_sll_454_net66365), .Z(u4_sll_454_ML_int_1__62_) );
  MUX2_X2 u4_sll_454_M1_0_63 ( .A(fract_denorm[63]), .B(fract_denorm[62]), .S(
        u4_sll_454_net66365), .Z(u4_sll_454_ML_int_1__63_) );
  MUX2_X2 u4_sll_454_M1_0_64 ( .A(fract_denorm[64]), .B(fract_denorm[63]), .S(
        u4_sll_454_net66365), .Z(u4_sll_454_ML_int_1__64_) );
  MUX2_X2 u4_sll_454_M1_0_65 ( .A(fract_denorm[65]), .B(fract_denorm[64]), .S(
        u4_sll_454_net66365), .Z(u4_sll_454_ML_int_1__65_) );
  MUX2_X2 u4_sll_454_M1_0_66 ( .A(fract_denorm[66]), .B(fract_denorm[65]), .S(
        u4_sll_454_net66367), .Z(u4_sll_454_ML_int_1__66_) );
  MUX2_X2 u4_sll_454_M1_0_67 ( .A(fract_denorm[67]), .B(fract_denorm[66]), .S(
        u4_sll_454_net66367), .Z(u4_sll_454_ML_int_1__67_) );
  MUX2_X2 u4_sll_454_M1_0_68 ( .A(fract_denorm[68]), .B(fract_denorm[67]), .S(
        u4_sll_454_net66367), .Z(u4_sll_454_ML_int_1__68_) );
  MUX2_X2 u4_sll_454_M1_0_69 ( .A(fract_denorm[69]), .B(fract_denorm[68]), .S(
        u4_sll_454_net66367), .Z(u4_sll_454_ML_int_1__69_) );
  MUX2_X2 u4_sll_454_M1_0_70 ( .A(fract_denorm[70]), .B(fract_denorm[69]), .S(
        u4_sll_454_net66367), .Z(u4_sll_454_ML_int_1__70_) );
  MUX2_X2 u4_sll_454_M1_0_71 ( .A(fract_denorm[71]), .B(fract_denorm[70]), .S(
        u4_sll_454_net66367), .Z(u4_sll_454_ML_int_1__71_) );
  MUX2_X2 u4_sll_454_M1_0_72 ( .A(fract_denorm[72]), .B(fract_denorm[71]), .S(
        u4_sll_454_net66367), .Z(u4_sll_454_ML_int_1__72_) );
  MUX2_X2 u4_sll_454_M1_0_73 ( .A(fract_denorm[73]), .B(fract_denorm[72]), .S(
        u4_sll_454_net66367), .Z(u4_sll_454_ML_int_1__73_) );
  MUX2_X2 u4_sll_454_M1_0_74 ( .A(fract_denorm[74]), .B(fract_denorm[73]), .S(
        u4_sll_454_net66367), .Z(u4_sll_454_ML_int_1__74_) );
  MUX2_X2 u4_sll_454_M1_0_75 ( .A(fract_denorm[75]), .B(fract_denorm[74]), .S(
        u4_sll_454_net66367), .Z(u4_sll_454_ML_int_1__75_) );
  MUX2_X2 u4_sll_454_M1_0_76 ( .A(fract_denorm[76]), .B(fract_denorm[75]), .S(
        u4_sll_454_net66367), .Z(u4_sll_454_ML_int_1__76_) );
  MUX2_X2 u4_sll_454_M1_0_77 ( .A(fract_denorm[77]), .B(fract_denorm[76]), .S(
        u4_sll_454_net66369), .Z(u4_sll_454_ML_int_1__77_) );
  MUX2_X2 u4_sll_454_M1_0_78 ( .A(fract_denorm[78]), .B(fract_denorm[77]), .S(
        u4_sll_454_net66369), .Z(u4_sll_454_ML_int_1__78_) );
  MUX2_X2 u4_sll_454_M1_0_79 ( .A(fract_denorm[79]), .B(fract_denorm[78]), .S(
        u4_sll_454_net66369), .Z(u4_sll_454_ML_int_1__79_) );
  MUX2_X2 u4_sll_454_M1_0_80 ( .A(fract_denorm[80]), .B(fract_denorm[79]), .S(
        u4_sll_454_net66369), .Z(u4_sll_454_ML_int_1__80_) );
  MUX2_X2 u4_sll_454_M1_0_81 ( .A(fract_denorm[81]), .B(fract_denorm[80]), .S(
        u4_sll_454_net66369), .Z(u4_sll_454_ML_int_1__81_) );
  MUX2_X2 u4_sll_454_M1_0_82 ( .A(fract_denorm[82]), .B(fract_denorm[81]), .S(
        u4_sll_454_net66369), .Z(u4_sll_454_ML_int_1__82_) );
  MUX2_X2 u4_sll_454_M1_0_83 ( .A(fract_denorm[83]), .B(fract_denorm[82]), .S(
        u4_sll_454_net66369), .Z(u4_sll_454_ML_int_1__83_) );
  MUX2_X2 u4_sll_454_M1_0_84 ( .A(fract_denorm[84]), .B(fract_denorm[83]), .S(
        u4_sll_454_net66369), .Z(u4_sll_454_ML_int_1__84_) );
  MUX2_X2 u4_sll_454_M1_0_85 ( .A(fract_denorm[85]), .B(fract_denorm[84]), .S(
        u4_sll_454_net66369), .Z(u4_sll_454_ML_int_1__85_) );
  MUX2_X2 u4_sll_454_M1_0_86 ( .A(fract_denorm[86]), .B(fract_denorm[85]), .S(
        u4_sll_454_net66369), .Z(u4_sll_454_ML_int_1__86_) );
  MUX2_X2 u4_sll_454_M1_0_87 ( .A(fract_denorm[87]), .B(fract_denorm[86]), .S(
        u4_sll_454_net66369), .Z(u4_sll_454_ML_int_1__87_) );
  MUX2_X2 u4_sll_454_M1_0_88 ( .A(fract_denorm[88]), .B(fract_denorm[87]), .S(
        u4_sll_454_net66371), .Z(u4_sll_454_ML_int_1__88_) );
  MUX2_X2 u4_sll_454_M1_0_89 ( .A(fract_denorm[89]), .B(fract_denorm[88]), .S(
        u4_sll_454_net66371), .Z(u4_sll_454_ML_int_1__89_) );
  MUX2_X2 u4_sll_454_M1_0_90 ( .A(fract_denorm[90]), .B(fract_denorm[89]), .S(
        u4_sll_454_net66371), .Z(u4_sll_454_ML_int_1__90_) );
  MUX2_X2 u4_sll_454_M1_0_91 ( .A(fract_denorm[91]), .B(fract_denorm[90]), .S(
        u4_sll_454_net66371), .Z(u4_sll_454_ML_int_1__91_) );
  MUX2_X2 u4_sll_454_M1_0_92 ( .A(fract_denorm[92]), .B(fract_denorm[91]), .S(
        u4_sll_454_net66371), .Z(u4_sll_454_ML_int_1__92_) );
  MUX2_X2 u4_sll_454_M1_0_93 ( .A(fract_denorm[93]), .B(fract_denorm[92]), .S(
        u4_sll_454_net66371), .Z(u4_sll_454_ML_int_1__93_) );
  MUX2_X2 u4_sll_454_M1_0_94 ( .A(fract_denorm[94]), .B(fract_denorm[93]), .S(
        u4_sll_454_net66371), .Z(u4_sll_454_ML_int_1__94_) );
  MUX2_X2 u4_sll_454_M1_0_95 ( .A(fract_denorm[95]), .B(fract_denorm[94]), .S(
        u4_sll_454_net66371), .Z(u4_sll_454_ML_int_1__95_) );
  MUX2_X2 u4_sll_454_M1_0_96 ( .A(fract_denorm[96]), .B(fract_denorm[95]), .S(
        u4_sll_454_net66371), .Z(u4_sll_454_ML_int_1__96_) );
  MUX2_X2 u4_sll_454_M1_0_97 ( .A(fract_denorm[97]), .B(fract_denorm[96]), .S(
        u4_sll_454_net66371), .Z(u4_sll_454_ML_int_1__97_) );
  MUX2_X2 u4_sll_454_M1_0_98 ( .A(fract_denorm[98]), .B(fract_denorm[97]), .S(
        u4_sll_454_net66371), .Z(u4_sll_454_ML_int_1__98_) );
  MUX2_X2 u4_sll_454_M1_0_99 ( .A(fract_denorm[99]), .B(fract_denorm[98]), .S(
        u4_sll_454_net66373), .Z(u4_sll_454_ML_int_1__99_) );
  MUX2_X2 u4_sll_454_M1_0_100 ( .A(fract_denorm[100]), .B(fract_denorm[99]), 
        .S(u4_sll_454_net66373), .Z(u4_sll_454_ML_int_1__100_) );
  MUX2_X2 u4_sll_454_M1_0_101 ( .A(fract_denorm[101]), .B(fract_denorm[100]), 
        .S(u4_sll_454_net66373), .Z(u4_sll_454_ML_int_1__101_) );
  MUX2_X2 u4_sll_454_M1_0_102 ( .A(fract_denorm[102]), .B(fract_denorm[101]), 
        .S(u4_sll_454_net66373), .Z(u4_sll_454_ML_int_1__102_) );
  MUX2_X2 u4_sll_454_M1_0_103 ( .A(fract_denorm[103]), .B(fract_denorm[102]), 
        .S(u4_sll_454_net66373), .Z(u4_sll_454_ML_int_1__103_) );
  MUX2_X2 u4_sll_454_M1_0_104 ( .A(fract_denorm[104]), .B(fract_denorm[103]), 
        .S(u4_sll_454_net66373), .Z(u4_sll_454_ML_int_1__104_) );
  MUX2_X2 u4_sll_454_M1_0_105 ( .A(net63217), .B(fract_denorm[104]), .S(
        u4_sll_454_net66373), .Z(u4_sll_454_ML_int_1__105_) );
  MUX2_X2 u4_sll_454_M1_1_2 ( .A(u4_sll_454_ML_int_1__2_), .B(
        u4_sll_454_ML_int_1__0_), .S(u4_sll_454_net66727), .Z(
        u4_sll_454_ML_int_2__2_) );
  MUX2_X2 u4_sll_454_M1_1_3 ( .A(u4_sll_454_ML_int_1__3_), .B(
        u4_sll_454_ML_int_1__1_), .S(u4_sll_454_net66727), .Z(
        u4_sll_454_ML_int_2__3_) );
  MUX2_X2 u4_sll_454_M1_1_4 ( .A(u4_sll_454_ML_int_1__4_), .B(
        u4_sll_454_ML_int_1__2_), .S(u4_sll_454_net66727), .Z(
        u4_sll_454_ML_int_2__4_) );
  MUX2_X2 u4_sll_454_M1_1_5 ( .A(u4_sll_454_ML_int_1__5_), .B(
        u4_sll_454_ML_int_1__3_), .S(u4_sll_454_net66727), .Z(
        u4_sll_454_ML_int_2__5_) );
  MUX2_X2 u4_sll_454_M1_1_6 ( .A(u4_sll_454_ML_int_1__6_), .B(
        u4_sll_454_ML_int_1__4_), .S(u4_sll_454_net66727), .Z(
        u4_sll_454_ML_int_2__6_) );
  MUX2_X2 u4_sll_454_M1_1_7 ( .A(u4_sll_454_ML_int_1__7_), .B(
        u4_sll_454_ML_int_1__5_), .S(u4_sll_454_net66723), .Z(
        u4_sll_454_ML_int_2__7_) );
  MUX2_X2 u4_sll_454_M1_1_8 ( .A(u4_sll_454_ML_int_1__8_), .B(
        u4_sll_454_ML_int_1__6_), .S(u4_sll_454_net66723), .Z(
        u4_sll_454_ML_int_2__8_) );
  MUX2_X2 u4_sll_454_M1_1_9 ( .A(u4_sll_454_ML_int_1__9_), .B(
        u4_sll_454_ML_int_1__7_), .S(u4_sll_454_net66717), .Z(
        u4_sll_454_ML_int_2__9_) );
  MUX2_X2 u4_sll_454_M1_1_10 ( .A(u4_sll_454_ML_int_1__10_), .B(
        u4_sll_454_ML_int_1__8_), .S(u4_sll_454_net66719), .Z(
        u4_sll_454_ML_int_2__10_) );
  MUX2_X2 u4_sll_454_M1_1_11 ( .A(u4_sll_454_ML_int_1__11_), .B(
        u4_sll_454_ML_int_1__9_), .S(u4_sll_454_net66723), .Z(
        u4_sll_454_ML_int_2__11_) );
  MUX2_X2 u4_sll_454_M1_1_12 ( .A(u4_sll_454_ML_int_1__12_), .B(
        u4_sll_454_ML_int_1__10_), .S(u4_sll_454_net66721), .Z(
        u4_sll_454_ML_int_2__12_) );
  MUX2_X2 u4_sll_454_M1_1_13 ( .A(u4_sll_454_ML_int_1__13_), .B(
        u4_sll_454_ML_int_1__11_), .S(u4_sll_454_net66721), .Z(
        u4_sll_454_ML_int_2__13_) );
  MUX2_X2 u4_sll_454_M1_1_15 ( .A(u4_sll_454_ML_int_1__15_), .B(
        u4_sll_454_ML_int_1__13_), .S(u4_sll_454_net66721), .Z(
        u4_sll_454_ML_int_2__15_) );
  MUX2_X2 u4_sll_454_M1_1_17 ( .A(u4_sll_454_ML_int_1__17_), .B(
        u4_sll_454_ML_int_1__15_), .S(u4_sll_454_net66711), .Z(
        u4_sll_454_ML_int_2__17_) );
  MUX2_X2 u4_sll_454_M1_1_19 ( .A(u4_sll_454_ML_int_1__19_), .B(
        u4_sll_454_ML_int_1__17_), .S(u4_sll_454_net66719), .Z(
        u4_sll_454_ML_int_2__19_) );
  MUX2_X2 u4_sll_454_M1_1_21 ( .A(u4_sll_454_ML_int_1__21_), .B(
        u4_sll_454_ML_int_1__19_), .S(u4_sll_454_net66715), .Z(
        u4_sll_454_ML_int_2__21_) );
  MUX2_X2 u4_sll_454_M1_1_22 ( .A(u4_sll_454_ML_int_1__22_), .B(
        u4_sll_454_ML_int_1__20_), .S(u4_sll_454_net66711), .Z(
        u4_sll_454_ML_int_2__22_) );
  MUX2_X2 u4_sll_454_M1_1_23 ( .A(u4_sll_454_ML_int_1__23_), .B(
        u4_sll_454_ML_int_1__21_), .S(u4_sll_454_net66711), .Z(
        u4_sll_454_ML_int_2__23_) );
  MUX2_X2 u4_sll_454_M1_1_24 ( .A(u4_sll_454_ML_int_1__24_), .B(
        u4_sll_454_ML_int_1__22_), .S(u4_sll_454_net66711), .Z(
        u4_sll_454_ML_int_2__24_) );
  MUX2_X2 u4_sll_454_M1_1_25 ( .A(u4_sll_454_ML_int_1__25_), .B(
        u4_sll_454_ML_int_1__23_), .S(u4_sll_454_net66711), .Z(
        u4_sll_454_ML_int_2__25_) );
  MUX2_X2 u4_sll_454_M1_1_26 ( .A(u4_sll_454_ML_int_1__26_), .B(
        u4_sll_454_ML_int_1__24_), .S(u4_sll_454_net66711), .Z(
        u4_sll_454_ML_int_2__26_) );
  MUX2_X2 u4_sll_454_M1_1_27 ( .A(u4_sll_454_ML_int_1__27_), .B(
        u4_sll_454_ML_int_1__25_), .S(u4_sll_454_net66711), .Z(
        u4_sll_454_ML_int_2__27_) );
  MUX2_X2 u4_sll_454_M1_1_28 ( .A(u4_sll_454_ML_int_1__28_), .B(
        u4_sll_454_ML_int_1__26_), .S(u4_sll_454_net66711), .Z(
        u4_sll_454_ML_int_2__28_) );
  MUX2_X2 u4_sll_454_M1_1_29 ( .A(u4_sll_454_ML_int_1__29_), .B(
        u4_sll_454_ML_int_1__27_), .S(u4_sll_454_net66711), .Z(
        u4_sll_454_ML_int_2__29_) );
  MUX2_X2 u4_sll_454_M1_1_30 ( .A(u4_sll_454_ML_int_1__30_), .B(
        u4_sll_454_ML_int_1__28_), .S(u4_sll_454_net66711), .Z(
        u4_sll_454_ML_int_2__30_) );
  MUX2_X2 u4_sll_454_M1_1_31 ( .A(u4_sll_454_ML_int_1__31_), .B(
        u4_sll_454_ML_int_1__29_), .S(u4_sll_454_net66711), .Z(
        u4_sll_454_ML_int_2__31_) );
  MUX2_X2 u4_sll_454_M1_1_32 ( .A(u4_sll_454_ML_int_1__32_), .B(
        u4_sll_454_ML_int_1__30_), .S(u4_sll_454_net66711), .Z(
        u4_sll_454_ML_int_2__32_) );
  MUX2_X2 u4_sll_454_M1_1_33 ( .A(u4_sll_454_ML_int_1__33_), .B(
        u4_sll_454_ML_int_1__31_), .S(u4_sll_454_net66715), .Z(
        u4_sll_454_ML_int_2__33_) );
  MUX2_X2 u4_sll_454_M1_1_34 ( .A(u4_sll_454_ML_int_1__34_), .B(
        u4_sll_454_ML_int_1__32_), .S(u4_sll_454_net66715), .Z(
        u4_sll_454_ML_int_2__34_) );
  MUX2_X2 u4_sll_454_M1_1_35 ( .A(u4_sll_454_ML_int_1__35_), .B(
        u4_sll_454_ML_int_1__33_), .S(u4_sll_454_net66711), .Z(
        u4_sll_454_ML_int_2__35_) );
  MUX2_X2 u4_sll_454_M1_1_36 ( .A(u4_sll_454_ML_int_1__36_), .B(
        u4_sll_454_ML_int_1__34_), .S(u4_sll_454_net66711), .Z(
        u4_sll_454_ML_int_2__36_) );
  MUX2_X2 u4_sll_454_M1_1_37 ( .A(u4_sll_454_ML_int_1__37_), .B(
        u4_sll_454_ML_int_1__35_), .S(u4_sll_454_net66711), .Z(
        u4_sll_454_ML_int_2__37_) );
  MUX2_X2 u4_sll_454_M1_1_38 ( .A(u4_sll_454_ML_int_1__38_), .B(
        u4_sll_454_ML_int_1__36_), .S(u4_sll_454_net66715), .Z(
        u4_sll_454_ML_int_2__38_) );
  MUX2_X2 u4_sll_454_M1_1_39 ( .A(u4_sll_454_ML_int_1__39_), .B(
        u4_sll_454_ML_int_1__37_), .S(u4_sll_454_net66715), .Z(
        u4_sll_454_ML_int_2__39_) );
  MUX2_X2 u4_sll_454_M1_1_40 ( .A(u4_sll_454_ML_int_1__40_), .B(
        u4_sll_454_ML_int_1__38_), .S(u4_sll_454_net66715), .Z(
        u4_sll_454_ML_int_2__40_) );
  MUX2_X2 u4_sll_454_M1_1_41 ( .A(u4_sll_454_ML_int_1__41_), .B(
        u4_sll_454_ML_int_1__39_), .S(u4_sll_454_net66711), .Z(
        u4_sll_454_ML_int_2__41_) );
  MUX2_X2 u4_sll_454_M1_1_42 ( .A(u4_sll_454_ML_int_1__42_), .B(
        u4_sll_454_ML_int_1__40_), .S(u4_sll_454_net66715), .Z(
        u4_sll_454_ML_int_2__42_) );
  MUX2_X2 u4_sll_454_M1_1_43 ( .A(u4_sll_454_ML_int_1__43_), .B(
        u4_sll_454_ML_int_1__41_), .S(u4_sll_454_net66711), .Z(
        u4_sll_454_ML_int_2__43_) );
  MUX2_X2 u4_sll_454_M1_1_44 ( .A(u4_sll_454_ML_int_1__44_), .B(
        u4_sll_454_ML_int_1__42_), .S(u4_sll_454_net66715), .Z(
        u4_sll_454_ML_int_2__44_) );
  MUX2_X2 u4_sll_454_M1_1_45 ( .A(u4_sll_454_ML_int_1__45_), .B(
        u4_sll_454_ML_int_1__43_), .S(u4_sll_454_net66715), .Z(
        u4_sll_454_ML_int_2__45_) );
  MUX2_X2 u4_sll_454_M1_1_46 ( .A(u4_sll_454_ML_int_1__46_), .B(
        u4_sll_454_ML_int_1__44_), .S(u4_sll_454_net66715), .Z(
        u4_sll_454_ML_int_2__46_) );
  MUX2_X2 u4_sll_454_M1_1_47 ( .A(u4_sll_454_ML_int_1__47_), .B(
        u4_sll_454_ML_int_1__45_), .S(u4_sll_454_net66715), .Z(
        u4_sll_454_ML_int_2__47_) );
  MUX2_X2 u4_sll_454_M1_1_48 ( .A(u4_sll_454_ML_int_1__48_), .B(
        u4_sll_454_ML_int_1__46_), .S(u4_sll_454_net66715), .Z(
        u4_sll_454_ML_int_2__48_) );
  MUX2_X2 u4_sll_454_M1_1_49 ( .A(u4_sll_454_ML_int_1__49_), .B(
        u4_sll_454_ML_int_1__47_), .S(u4_sll_454_net66715), .Z(
        u4_sll_454_ML_int_2__49_) );
  MUX2_X2 u4_sll_454_M1_1_50 ( .A(u4_sll_454_ML_int_1__50_), .B(
        u4_sll_454_ML_int_1__48_), .S(u4_sll_454_net66715), .Z(
        u4_sll_454_ML_int_2__50_) );
  MUX2_X2 u4_sll_454_M1_1_51 ( .A(u4_sll_454_ML_int_1__51_), .B(
        u4_sll_454_ML_int_1__49_), .S(u4_sll_454_net66715), .Z(
        u4_sll_454_ML_int_2__51_) );
  MUX2_X2 u4_sll_454_M1_1_52 ( .A(u4_sll_454_ML_int_1__52_), .B(
        u4_sll_454_ML_int_1__50_), .S(u4_sll_454_net66715), .Z(
        u4_sll_454_ML_int_2__52_) );
  MUX2_X2 u4_sll_454_M1_1_53 ( .A(u4_sll_454_ML_int_1__53_), .B(
        u4_sll_454_ML_int_1__51_), .S(u4_sll_454_net66715), .Z(
        u4_sll_454_ML_int_2__53_) );
  MUX2_X2 u4_sll_454_M1_1_54 ( .A(u4_sll_454_ML_int_1__54_), .B(
        u4_sll_454_ML_int_1__52_), .S(u4_sll_454_net66715), .Z(
        u4_sll_454_ML_int_2__54_) );
  MUX2_X2 u4_sll_454_M1_1_55 ( .A(u4_sll_454_ML_int_1__55_), .B(
        u4_sll_454_ML_int_1__53_), .S(u4_sll_454_net66717), .Z(
        u4_sll_454_ML_int_2__55_) );
  MUX2_X2 u4_sll_454_M1_1_56 ( .A(u4_sll_454_ML_int_1__56_), .B(
        u4_sll_454_ML_int_1__54_), .S(u4_sll_454_net66717), .Z(
        u4_sll_454_ML_int_2__56_) );
  MUX2_X2 u4_sll_454_M1_1_57 ( .A(u4_sll_454_ML_int_1__57_), .B(
        u4_sll_454_ML_int_1__55_), .S(u4_sll_454_net66717), .Z(
        u4_sll_454_ML_int_2__57_) );
  MUX2_X2 u4_sll_454_M1_1_58 ( .A(u4_sll_454_ML_int_1__58_), .B(
        u4_sll_454_ML_int_1__56_), .S(u4_sll_454_net66717), .Z(
        u4_sll_454_ML_int_2__58_) );
  MUX2_X2 u4_sll_454_M1_1_59 ( .A(u4_sll_454_ML_int_1__59_), .B(
        u4_sll_454_ML_int_1__57_), .S(u4_sll_454_net66717), .Z(
        u4_sll_454_ML_int_2__59_) );
  MUX2_X2 u4_sll_454_M1_1_60 ( .A(u4_sll_454_ML_int_1__60_), .B(
        u4_sll_454_ML_int_1__58_), .S(u4_sll_454_net66717), .Z(
        u4_sll_454_ML_int_2__60_) );
  MUX2_X2 u4_sll_454_M1_1_61 ( .A(u4_sll_454_ML_int_1__61_), .B(
        u4_sll_454_ML_int_1__59_), .S(u4_sll_454_net66717), .Z(
        u4_sll_454_ML_int_2__61_) );
  MUX2_X2 u4_sll_454_M1_1_62 ( .A(u4_sll_454_ML_int_1__62_), .B(
        u4_sll_454_ML_int_1__60_), .S(u4_sll_454_net66717), .Z(
        u4_sll_454_ML_int_2__62_) );
  MUX2_X2 u4_sll_454_M1_1_63 ( .A(u4_sll_454_ML_int_1__63_), .B(
        u4_sll_454_ML_int_1__61_), .S(u4_sll_454_net66717), .Z(
        u4_sll_454_ML_int_2__63_) );
  MUX2_X2 u4_sll_454_M1_1_64 ( .A(u4_sll_454_ML_int_1__64_), .B(
        u4_sll_454_ML_int_1__62_), .S(u4_sll_454_net66717), .Z(
        u4_sll_454_ML_int_2__64_) );
  MUX2_X2 u4_sll_454_M1_1_65 ( .A(u4_sll_454_ML_int_1__65_), .B(
        u4_sll_454_ML_int_1__63_), .S(u4_sll_454_net66717), .Z(
        u4_sll_454_ML_int_2__65_) );
  MUX2_X2 u4_sll_454_M1_1_66 ( .A(u4_sll_454_ML_int_1__66_), .B(
        u4_sll_454_ML_int_1__64_), .S(u4_sll_454_net66719), .Z(
        u4_sll_454_ML_int_2__66_) );
  MUX2_X2 u4_sll_454_M1_1_67 ( .A(u4_sll_454_ML_int_1__67_), .B(
        u4_sll_454_ML_int_1__65_), .S(u4_sll_454_net66719), .Z(
        u4_sll_454_ML_int_2__67_) );
  MUX2_X2 u4_sll_454_M1_1_68 ( .A(u4_sll_454_ML_int_1__68_), .B(
        u4_sll_454_ML_int_1__66_), .S(u4_sll_454_net66719), .Z(
        u4_sll_454_ML_int_2__68_) );
  MUX2_X2 u4_sll_454_M1_1_69 ( .A(u4_sll_454_ML_int_1__69_), .B(
        u4_sll_454_ML_int_1__67_), .S(u4_sll_454_net66719), .Z(
        u4_sll_454_ML_int_2__69_) );
  MUX2_X2 u4_sll_454_M1_1_70 ( .A(u4_sll_454_ML_int_1__70_), .B(
        u4_sll_454_ML_int_1__68_), .S(u4_sll_454_net66719), .Z(
        u4_sll_454_ML_int_2__70_) );
  MUX2_X2 u4_sll_454_M1_1_71 ( .A(u4_sll_454_ML_int_1__71_), .B(
        u4_sll_454_ML_int_1__69_), .S(u4_sll_454_net66719), .Z(
        u4_sll_454_ML_int_2__71_) );
  MUX2_X2 u4_sll_454_M1_1_72 ( .A(u4_sll_454_ML_int_1__72_), .B(
        u4_sll_454_ML_int_1__70_), .S(u4_sll_454_net66719), .Z(
        u4_sll_454_ML_int_2__72_) );
  MUX2_X2 u4_sll_454_M1_1_73 ( .A(u4_sll_454_ML_int_1__73_), .B(
        u4_sll_454_ML_int_1__71_), .S(u4_sll_454_net66719), .Z(
        u4_sll_454_ML_int_2__73_) );
  MUX2_X2 u4_sll_454_M1_1_74 ( .A(u4_sll_454_ML_int_1__74_), .B(
        u4_sll_454_ML_int_1__72_), .S(u4_sll_454_net66719), .Z(
        u4_sll_454_ML_int_2__74_) );
  MUX2_X2 u4_sll_454_M1_1_75 ( .A(u4_sll_454_ML_int_1__75_), .B(
        u4_sll_454_ML_int_1__73_), .S(u4_sll_454_net66719), .Z(
        u4_sll_454_ML_int_2__75_) );
  MUX2_X2 u4_sll_454_M1_1_76 ( .A(u4_sll_454_ML_int_1__76_), .B(
        u4_sll_454_ML_int_1__74_), .S(u4_sll_454_net66719), .Z(
        u4_sll_454_ML_int_2__76_) );
  MUX2_X2 u4_sll_454_M1_1_77 ( .A(u4_sll_454_ML_int_1__77_), .B(
        u4_sll_454_ML_int_1__75_), .S(u4_sll_454_net66721), .Z(
        u4_sll_454_ML_int_2__77_) );
  MUX2_X2 u4_sll_454_M1_1_78 ( .A(u4_sll_454_ML_int_1__78_), .B(
        u4_sll_454_ML_int_1__76_), .S(u4_sll_454_net66721), .Z(
        u4_sll_454_ML_int_2__78_) );
  MUX2_X2 u4_sll_454_M1_1_79 ( .A(u4_sll_454_ML_int_1__79_), .B(
        u4_sll_454_ML_int_1__77_), .S(u4_sll_454_net66721), .Z(
        u4_sll_454_ML_int_2__79_) );
  MUX2_X2 u4_sll_454_M1_1_80 ( .A(u4_sll_454_ML_int_1__80_), .B(
        u4_sll_454_ML_int_1__78_), .S(u4_sll_454_net66721), .Z(
        u4_sll_454_ML_int_2__80_) );
  MUX2_X2 u4_sll_454_M1_1_81 ( .A(u4_sll_454_ML_int_1__81_), .B(
        u4_sll_454_ML_int_1__79_), .S(u4_sll_454_net66721), .Z(
        u4_sll_454_ML_int_2__81_) );
  MUX2_X2 u4_sll_454_M1_1_82 ( .A(u4_sll_454_ML_int_1__82_), .B(
        u4_sll_454_ML_int_1__80_), .S(u4_sll_454_net66721), .Z(
        u4_sll_454_ML_int_2__82_) );
  MUX2_X2 u4_sll_454_M1_1_83 ( .A(u4_sll_454_ML_int_1__83_), .B(
        u4_sll_454_ML_int_1__81_), .S(u4_sll_454_net66721), .Z(
        u4_sll_454_ML_int_2__83_) );
  MUX2_X2 u4_sll_454_M1_1_84 ( .A(u4_sll_454_ML_int_1__84_), .B(
        u4_sll_454_ML_int_1__82_), .S(u4_sll_454_net66721), .Z(
        u4_sll_454_ML_int_2__84_) );
  MUX2_X2 u4_sll_454_M1_1_85 ( .A(u4_sll_454_ML_int_1__85_), .B(
        u4_sll_454_ML_int_1__83_), .S(u4_sll_454_net66721), .Z(
        u4_sll_454_ML_int_2__85_) );
  MUX2_X2 u4_sll_454_M1_1_86 ( .A(u4_sll_454_ML_int_1__86_), .B(
        u4_sll_454_ML_int_1__84_), .S(u4_sll_454_net66721), .Z(
        u4_sll_454_ML_int_2__86_) );
  MUX2_X2 u4_sll_454_M1_1_87 ( .A(u4_sll_454_ML_int_1__87_), .B(
        u4_sll_454_ML_int_1__85_), .S(u4_sll_454_net66721), .Z(
        u4_sll_454_ML_int_2__87_) );
  MUX2_X2 u4_sll_454_M1_1_88 ( .A(u4_sll_454_ML_int_1__88_), .B(
        u4_sll_454_ML_int_1__86_), .S(u4_sll_454_net66723), .Z(
        u4_sll_454_ML_int_2__88_) );
  MUX2_X2 u4_sll_454_M1_1_89 ( .A(u4_sll_454_ML_int_1__89_), .B(
        u4_sll_454_ML_int_1__87_), .S(u4_sll_454_net66723), .Z(
        u4_sll_454_ML_int_2__89_) );
  MUX2_X2 u4_sll_454_M1_1_90 ( .A(u4_sll_454_ML_int_1__90_), .B(
        u4_sll_454_ML_int_1__88_), .S(u4_sll_454_net66723), .Z(
        u4_sll_454_ML_int_2__90_) );
  MUX2_X2 u4_sll_454_M1_1_91 ( .A(u4_sll_454_ML_int_1__91_), .B(
        u4_sll_454_ML_int_1__89_), .S(u4_sll_454_net66723), .Z(
        u4_sll_454_ML_int_2__91_) );
  MUX2_X2 u4_sll_454_M1_1_92 ( .A(u4_sll_454_ML_int_1__92_), .B(
        u4_sll_454_ML_int_1__90_), .S(u4_sll_454_net66723), .Z(
        u4_sll_454_ML_int_2__92_) );
  MUX2_X2 u4_sll_454_M1_1_93 ( .A(u4_sll_454_ML_int_1__93_), .B(
        u4_sll_454_ML_int_1__91_), .S(u4_sll_454_net66723), .Z(
        u4_sll_454_ML_int_2__93_) );
  MUX2_X2 u4_sll_454_M1_1_94 ( .A(u4_sll_454_ML_int_1__94_), .B(
        u4_sll_454_ML_int_1__92_), .S(u4_sll_454_net66723), .Z(
        u4_sll_454_ML_int_2__94_) );
  MUX2_X2 u4_sll_454_M1_1_95 ( .A(u4_sll_454_ML_int_1__95_), .B(
        u4_sll_454_ML_int_1__93_), .S(u4_sll_454_net66723), .Z(
        u4_sll_454_ML_int_2__95_) );
  MUX2_X2 u4_sll_454_M1_1_96 ( .A(u4_sll_454_ML_int_1__96_), .B(
        u4_sll_454_ML_int_1__94_), .S(u4_sll_454_net66723), .Z(
        u4_sll_454_ML_int_2__96_) );
  MUX2_X2 u4_sll_454_M1_1_97 ( .A(u4_sll_454_ML_int_1__97_), .B(
        u4_sll_454_ML_int_1__95_), .S(u4_sll_454_net66723), .Z(
        u4_sll_454_ML_int_2__97_) );
  MUX2_X2 u4_sll_454_M1_1_98 ( .A(u4_sll_454_ML_int_1__98_), .B(
        u4_sll_454_ML_int_1__96_), .S(u4_sll_454_net66723), .Z(
        u4_sll_454_ML_int_2__98_) );
  MUX2_X2 u4_sll_454_M1_1_99 ( .A(u4_sll_454_ML_int_1__99_), .B(
        u4_sll_454_ML_int_1__97_), .S(u4_sll_454_net66723), .Z(
        u4_sll_454_ML_int_2__99_) );
  MUX2_X2 u4_sll_454_M1_1_100 ( .A(u4_sll_454_ML_int_1__100_), .B(
        u4_sll_454_ML_int_1__98_), .S(u4_sll_454_net66715), .Z(
        u4_sll_454_ML_int_2__100_) );
  MUX2_X2 u4_sll_454_M1_1_101 ( .A(u4_sll_454_ML_int_1__101_), .B(
        u4_sll_454_ML_int_1__99_), .S(u4_sll_454_net66711), .Z(
        u4_sll_454_ML_int_2__101_) );
  MUX2_X2 u4_sll_454_M1_1_102 ( .A(u4_sll_454_ML_int_1__102_), .B(
        u4_sll_454_ML_int_1__100_), .S(u4_sll_454_net66717), .Z(
        u4_sll_454_ML_int_2__102_) );
  MUX2_X2 u4_sll_454_M1_1_103 ( .A(u4_sll_454_ML_int_1__103_), .B(
        u4_sll_454_ML_int_1__101_), .S(u4_sll_454_net66719), .Z(
        u4_sll_454_ML_int_2__103_) );
  MUX2_X2 u4_sll_454_M1_1_104 ( .A(u4_sll_454_ML_int_1__104_), .B(
        u4_sll_454_ML_int_1__102_), .S(u4_sll_454_net66723), .Z(
        u4_sll_454_ML_int_2__104_) );
  MUX2_X2 u4_sll_454_M1_1_105 ( .A(u4_sll_454_ML_int_1__105_), .B(
        u4_sll_454_ML_int_1__103_), .S(u4_sll_454_net66715), .Z(
        u4_sll_454_ML_int_2__105_) );
  MUX2_X2 u4_sll_454_M1_2_4 ( .A(u4_sll_454_ML_int_2__4_), .B(
        u4_sll_454_ML_int_2__0_), .S(u4_sll_454_net66667), .Z(
        u4_sll_454_ML_int_3__4_) );
  MUX2_X2 u4_sll_454_M1_2_5 ( .A(u4_sll_454_ML_int_2__5_), .B(
        u4_sll_454_ML_int_2__1_), .S(u4_sll_454_net66667), .Z(
        u4_sll_454_ML_int_3__5_) );
  MUX2_X2 u4_sll_454_M1_2_6 ( .A(u4_sll_454_ML_int_2__6_), .B(
        u4_sll_454_ML_int_2__2_), .S(u4_sll_454_net66667), .Z(
        u4_sll_454_ML_int_3__6_) );
  MUX2_X2 u4_sll_454_M1_2_7 ( .A(u4_sll_454_ML_int_2__7_), .B(
        u4_sll_454_ML_int_2__3_), .S(u4_sll_454_net66667), .Z(
        u4_sll_454_ML_int_3__7_) );
  MUX2_X2 u4_sll_454_M1_2_8 ( .A(u4_sll_454_ML_int_2__8_), .B(
        u4_sll_454_ML_int_2__4_), .S(u4_sll_454_net66699), .Z(
        u4_sll_454_ML_int_3__8_) );
  MUX2_X2 u4_sll_454_M1_2_9 ( .A(u4_sll_454_ML_int_2__9_), .B(
        u4_sll_454_ML_int_2__5_), .S(u4_sll_454_net66699), .Z(
        u4_sll_454_ML_int_3__9_) );
  MUX2_X2 u4_sll_454_M1_2_10 ( .A(u4_sll_454_ML_int_2__10_), .B(
        u4_sll_454_ML_int_2__6_), .S(u4_sll_454_net66699), .Z(
        u4_sll_454_ML_int_3__10_) );
  MUX2_X2 u4_sll_454_M1_2_11 ( .A(u4_sll_454_ML_int_2__11_), .B(
        u4_sll_454_ML_int_2__7_), .S(u4_sll_454_net66699), .Z(
        u4_sll_454_ML_int_3__11_) );
  MUX2_X2 u4_sll_454_M1_2_12 ( .A(u4_sll_454_ML_int_2__12_), .B(
        u4_sll_454_ML_int_2__8_), .S(u4_sll_454_net66699), .Z(
        u4_sll_454_ML_int_3__12_) );
  MUX2_X2 u4_sll_454_M1_2_13 ( .A(u4_sll_454_ML_int_2__13_), .B(
        u4_sll_454_ML_int_2__9_), .S(u4_sll_454_net66699), .Z(
        u4_sll_454_ML_int_3__13_) );
  MUX2_X2 u4_sll_454_M1_2_14 ( .A(u4_sll_454_ML_int_2__14_), .B(
        u4_sll_454_ML_int_2__10_), .S(u4_sll_454_net66699), .Z(
        u4_sll_454_ML_int_3__14_) );
  MUX2_X2 u4_sll_454_M1_2_15 ( .A(u4_sll_454_ML_int_2__15_), .B(
        u4_sll_454_ML_int_2__11_), .S(u4_sll_454_net66699), .Z(
        u4_sll_454_ML_int_3__15_) );
  MUX2_X2 u4_sll_454_M1_2_17 ( .A(u4_sll_454_ML_int_2__17_), .B(
        u4_sll_454_ML_int_2__13_), .S(u4_sll_454_net66699), .Z(
        u4_sll_454_ML_int_3__17_) );
  MUX2_X2 u4_sll_454_M1_2_18 ( .A(u4_sll_454_ML_int_2__18_), .B(
        u4_sll_454_ML_int_2__14_), .S(u4_sll_454_net66699), .Z(
        u4_sll_454_ML_int_3__18_) );
  MUX2_X2 u4_sll_454_M1_2_19 ( .A(u4_sll_454_ML_int_2__19_), .B(
        u4_sll_454_ML_int_2__15_), .S(u4_sll_454_net66661), .Z(
        u4_sll_454_ML_int_3__19_) );
  MUX2_X2 u4_sll_454_M1_2_21 ( .A(u4_sll_454_ML_int_2__21_), .B(
        u4_sll_454_ML_int_2__17_), .S(u4_sll_454_net66699), .Z(
        u4_sll_454_ML_int_3__21_) );
  MUX2_X2 u4_sll_454_M1_2_22 ( .A(u4_sll_454_ML_int_2__22_), .B(
        u4_sll_454_ML_int_2__18_), .S(u4_sll_454_net66655), .Z(
        u4_sll_454_ML_int_3__22_) );
  MUX2_X2 u4_sll_454_M1_2_23 ( .A(u4_sll_454_ML_int_2__23_), .B(
        u4_sll_454_ML_int_2__19_), .S(u4_sll_454_net66655), .Z(
        u4_sll_454_ML_int_3__23_) );
  MUX2_X2 u4_sll_454_M1_2_25 ( .A(u4_sll_454_ML_int_2__25_), .B(
        u4_sll_454_ML_int_2__21_), .S(u4_sll_454_net66655), .Z(
        u4_sll_454_ML_int_3__25_) );
  MUX2_X2 u4_sll_454_M1_2_26 ( .A(u4_sll_454_ML_int_2__26_), .B(
        u4_sll_454_ML_int_2__22_), .S(u4_sll_454_net66655), .Z(
        u4_sll_454_ML_int_3__26_) );
  MUX2_X2 u4_sll_454_M1_2_27 ( .A(u4_sll_454_ML_int_2__27_), .B(
        u4_sll_454_ML_int_2__23_), .S(u4_sll_454_net66655), .Z(
        u4_sll_454_ML_int_3__27_) );
  MUX2_X2 u4_sll_454_M1_2_29 ( .A(u4_sll_454_ML_int_2__29_), .B(
        u4_sll_454_ML_int_2__25_), .S(u4_sll_454_net66655), .Z(
        u4_sll_454_ML_int_3__29_) );
  MUX2_X2 u4_sll_454_M1_2_30 ( .A(u4_sll_454_ML_int_2__30_), .B(
        u4_sll_454_ML_int_2__26_), .S(u4_sll_454_net66655), .Z(
        u4_sll_454_ML_int_3__30_) );
  MUX2_X2 u4_sll_454_M1_2_31 ( .A(u4_sll_454_ML_int_2__31_), .B(
        u4_sll_454_ML_int_2__27_), .S(u4_sll_454_net66655), .Z(
        u4_sll_454_ML_int_3__31_) );
  MUX2_X2 u4_sll_454_M1_2_32 ( .A(u4_sll_454_ML_int_2__32_), .B(
        u4_sll_454_ML_int_2__28_), .S(u4_sll_454_net66655), .Z(
        u4_sll_454_ML_int_3__32_) );
  MUX2_X2 u4_sll_454_M1_2_33 ( .A(u4_sll_454_ML_int_2__33_), .B(
        u4_sll_454_ML_int_2__29_), .S(u4_sll_454_net66661), .Z(
        u4_sll_454_ML_int_3__33_) );
  MUX2_X2 u4_sll_454_M1_2_34 ( .A(u4_sll_454_ML_int_2__34_), .B(
        u4_sll_454_ML_int_2__30_), .S(u4_sll_454_net66697), .Z(
        u4_sll_454_ML_int_3__34_) );
  MUX2_X2 u4_sll_454_M1_2_35 ( .A(u4_sll_454_ML_int_2__35_), .B(
        u4_sll_454_ML_int_2__31_), .S(u4_sll_454_net66659), .Z(
        u4_sll_454_ML_int_3__35_) );
  MUX2_X2 u4_sll_454_M1_2_36 ( .A(u4_sll_454_ML_int_2__36_), .B(
        u4_sll_454_ML_int_2__32_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__36_) );
  MUX2_X2 u4_sll_454_M1_2_37 ( .A(u4_sll_454_ML_int_2__37_), .B(
        u4_sll_454_ML_int_2__33_), .S(u4_sll_454_net66659), .Z(
        u4_sll_454_ML_int_3__37_) );
  MUX2_X2 u4_sll_454_M1_2_38 ( .A(u4_sll_454_ML_int_2__38_), .B(
        u4_sll_454_ML_int_2__34_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__38_) );
  MUX2_X2 u4_sll_454_M1_2_39 ( .A(u4_sll_454_ML_int_2__39_), .B(
        u4_sll_454_ML_int_2__35_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__39_) );
  MUX2_X2 u4_sll_454_M1_2_40 ( .A(u4_sll_454_ML_int_2__40_), .B(
        u4_sll_454_ML_int_2__36_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__40_) );
  MUX2_X2 u4_sll_454_M1_2_41 ( .A(u4_sll_454_ML_int_2__41_), .B(
        u4_sll_454_ML_int_2__37_), .S(u4_sll_454_net66659), .Z(
        u4_sll_454_ML_int_3__41_) );
  MUX2_X2 u4_sll_454_M1_2_42 ( .A(u4_sll_454_ML_int_2__42_), .B(
        u4_sll_454_ML_int_2__38_), .S(u4_sll_454_net66659), .Z(
        u4_sll_454_ML_int_3__42_) );
  MUX2_X2 u4_sll_454_M1_2_43 ( .A(u4_sll_454_ML_int_2__43_), .B(
        u4_sll_454_ML_int_2__39_), .S(u4_sll_454_net66659), .Z(
        u4_sll_454_ML_int_3__43_) );
  MUX2_X2 u4_sll_454_M1_2_44 ( .A(u4_sll_454_ML_int_2__44_), .B(
        u4_sll_454_ML_int_2__40_), .S(u4_sll_454_net66659), .Z(
        u4_sll_454_ML_int_3__44_) );
  MUX2_X2 u4_sll_454_M1_2_45 ( .A(u4_sll_454_ML_int_2__45_), .B(
        u4_sll_454_ML_int_2__41_), .S(u4_sll_454_net66659), .Z(
        u4_sll_454_ML_int_3__45_) );
  MUX2_X2 u4_sll_454_M1_2_46 ( .A(u4_sll_454_ML_int_2__46_), .B(
        u4_sll_454_ML_int_2__42_), .S(u4_sll_454_net66659), .Z(
        u4_sll_454_ML_int_3__46_) );
  MUX2_X2 u4_sll_454_M1_2_47 ( .A(u4_sll_454_ML_int_2__47_), .B(
        u4_sll_454_ML_int_2__43_), .S(u4_sll_454_net66659), .Z(
        u4_sll_454_ML_int_3__47_) );
  MUX2_X2 u4_sll_454_M1_2_48 ( .A(u4_sll_454_ML_int_2__48_), .B(
        u4_sll_454_ML_int_2__44_), .S(u4_sll_454_net66659), .Z(
        u4_sll_454_ML_int_3__48_) );
  MUX2_X2 u4_sll_454_M1_2_49 ( .A(u4_sll_454_ML_int_2__49_), .B(
        u4_sll_454_ML_int_2__45_), .S(u4_sll_454_net66659), .Z(
        u4_sll_454_ML_int_3__49_) );
  MUX2_X2 u4_sll_454_M1_2_50 ( .A(u4_sll_454_ML_int_2__50_), .B(
        u4_sll_454_ML_int_2__46_), .S(u4_sll_454_net66659), .Z(
        u4_sll_454_ML_int_3__50_) );
  MUX2_X2 u4_sll_454_M1_2_51 ( .A(u4_sll_454_ML_int_2__51_), .B(
        u4_sll_454_ML_int_2__47_), .S(u4_sll_454_net66659), .Z(
        u4_sll_454_ML_int_3__51_) );
  MUX2_X2 u4_sll_454_M1_2_52 ( .A(u4_sll_454_ML_int_2__52_), .B(
        u4_sll_454_ML_int_2__48_), .S(u4_sll_454_net66659), .Z(
        u4_sll_454_ML_int_3__52_) );
  MUX2_X2 u4_sll_454_M1_2_53 ( .A(u4_sll_454_ML_int_2__53_), .B(
        u4_sll_454_ML_int_2__49_), .S(u4_sll_454_net66659), .Z(
        u4_sll_454_ML_int_3__53_) );
  MUX2_X2 u4_sll_454_M1_2_54 ( .A(u4_sll_454_ML_int_2__54_), .B(
        u4_sll_454_ML_int_2__50_), .S(u4_sll_454_net66659), .Z(
        u4_sll_454_ML_int_3__54_) );
  MUX2_X2 u4_sll_454_M1_2_55 ( .A(u4_sll_454_ML_int_2__55_), .B(
        u4_sll_454_ML_int_2__51_), .S(u4_sll_454_net66661), .Z(
        u4_sll_454_ML_int_3__55_) );
  MUX2_X2 u4_sll_454_M1_2_56 ( .A(u4_sll_454_ML_int_2__56_), .B(
        u4_sll_454_ML_int_2__52_), .S(u4_sll_454_net66661), .Z(
        u4_sll_454_ML_int_3__56_) );
  MUX2_X2 u4_sll_454_M1_2_57 ( .A(u4_sll_454_ML_int_2__57_), .B(
        u4_sll_454_ML_int_2__53_), .S(u4_sll_454_net66661), .Z(
        u4_sll_454_ML_int_3__57_) );
  MUX2_X2 u4_sll_454_M1_2_58 ( .A(u4_sll_454_ML_int_2__58_), .B(
        u4_sll_454_ML_int_2__54_), .S(u4_sll_454_net66661), .Z(
        u4_sll_454_ML_int_3__58_) );
  MUX2_X2 u4_sll_454_M1_2_59 ( .A(u4_sll_454_ML_int_2__59_), .B(
        u4_sll_454_ML_int_2__55_), .S(u4_sll_454_net66661), .Z(
        u4_sll_454_ML_int_3__59_) );
  MUX2_X2 u4_sll_454_M1_2_60 ( .A(u4_sll_454_ML_int_2__60_), .B(
        u4_sll_454_ML_int_2__56_), .S(u4_sll_454_net66661), .Z(
        u4_sll_454_ML_int_3__60_) );
  MUX2_X2 u4_sll_454_M1_2_61 ( .A(u4_sll_454_ML_int_2__61_), .B(
        u4_sll_454_ML_int_2__57_), .S(u4_sll_454_net66661), .Z(
        u4_sll_454_ML_int_3__61_) );
  MUX2_X2 u4_sll_454_M1_2_62 ( .A(u4_sll_454_ML_int_2__62_), .B(
        u4_sll_454_ML_int_2__58_), .S(u4_sll_454_net66661), .Z(
        u4_sll_454_ML_int_3__62_) );
  MUX2_X2 u4_sll_454_M1_2_63 ( .A(u4_sll_454_ML_int_2__63_), .B(
        u4_sll_454_ML_int_2__59_), .S(u4_sll_454_net66661), .Z(
        u4_sll_454_ML_int_3__63_) );
  MUX2_X2 u4_sll_454_M1_2_64 ( .A(u4_sll_454_ML_int_2__64_), .B(
        u4_sll_454_ML_int_2__60_), .S(u4_sll_454_net66661), .Z(
        u4_sll_454_ML_int_3__64_) );
  MUX2_X2 u4_sll_454_M1_2_65 ( .A(u4_sll_454_ML_int_2__65_), .B(
        u4_sll_454_ML_int_2__61_), .S(u4_sll_454_net66661), .Z(
        u4_sll_454_ML_int_3__65_) );
  MUX2_X2 u4_sll_454_M1_2_66 ( .A(u4_sll_454_ML_int_2__66_), .B(
        u4_sll_454_ML_int_2__62_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__66_) );
  MUX2_X2 u4_sll_454_M1_2_67 ( .A(u4_sll_454_ML_int_2__67_), .B(
        u4_sll_454_ML_int_2__63_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__67_) );
  MUX2_X2 u4_sll_454_M1_2_68 ( .A(u4_sll_454_ML_int_2__68_), .B(
        u4_sll_454_ML_int_2__64_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__68_) );
  MUX2_X2 u4_sll_454_M1_2_69 ( .A(u4_sll_454_ML_int_2__69_), .B(
        u4_sll_454_ML_int_2__65_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__69_) );
  MUX2_X2 u4_sll_454_M1_2_70 ( .A(u4_sll_454_ML_int_2__70_), .B(
        u4_sll_454_ML_int_2__66_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__70_) );
  MUX2_X2 u4_sll_454_M1_2_71 ( .A(u4_sll_454_ML_int_2__71_), .B(
        u4_sll_454_ML_int_2__67_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__71_) );
  MUX2_X2 u4_sll_454_M1_2_72 ( .A(u4_sll_454_ML_int_2__72_), .B(
        u4_sll_454_ML_int_2__68_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__72_) );
  MUX2_X2 u4_sll_454_M1_2_73 ( .A(u4_sll_454_ML_int_2__73_), .B(
        u4_sll_454_ML_int_2__69_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__73_) );
  MUX2_X2 u4_sll_454_M1_2_74 ( .A(u4_sll_454_ML_int_2__74_), .B(
        u4_sll_454_ML_int_2__70_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__74_) );
  MUX2_X2 u4_sll_454_M1_2_75 ( .A(u4_sll_454_ML_int_2__75_), .B(
        u4_sll_454_ML_int_2__71_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__75_) );
  MUX2_X2 u4_sll_454_M1_2_76 ( .A(u4_sll_454_ML_int_2__76_), .B(
        u4_sll_454_ML_int_2__72_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__76_) );
  MUX2_X2 u4_sll_454_M1_2_77 ( .A(u4_sll_454_ML_int_2__77_), .B(
        u4_sll_454_ML_int_2__73_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__77_) );
  MUX2_X2 u4_sll_454_M1_2_78 ( .A(u4_sll_454_ML_int_2__78_), .B(
        u4_sll_454_ML_int_2__74_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__78_) );
  MUX2_X2 u4_sll_454_M1_2_79 ( .A(u4_sll_454_ML_int_2__79_), .B(
        u4_sll_454_ML_int_2__75_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__79_) );
  MUX2_X2 u4_sll_454_M1_2_80 ( .A(u4_sll_454_ML_int_2__80_), .B(
        u4_sll_454_ML_int_2__76_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__80_) );
  MUX2_X2 u4_sll_454_M1_2_81 ( .A(u4_sll_454_ML_int_2__81_), .B(
        u4_sll_454_ML_int_2__77_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__81_) );
  MUX2_X2 u4_sll_454_M1_2_82 ( .A(u4_sll_454_ML_int_2__82_), .B(
        u4_sll_454_ML_int_2__78_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__82_) );
  MUX2_X2 u4_sll_454_M1_2_83 ( .A(u4_sll_454_ML_int_2__83_), .B(
        u4_sll_454_ML_int_2__79_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__83_) );
  MUX2_X2 u4_sll_454_M1_2_84 ( .A(u4_sll_454_ML_int_2__84_), .B(
        u4_sll_454_ML_int_2__80_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__84_) );
  MUX2_X2 u4_sll_454_M1_2_85 ( .A(u4_sll_454_ML_int_2__85_), .B(
        u4_sll_454_ML_int_2__81_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__85_) );
  MUX2_X2 u4_sll_454_M1_2_86 ( .A(u4_sll_454_ML_int_2__86_), .B(
        u4_sll_454_ML_int_2__82_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__86_) );
  MUX2_X2 u4_sll_454_M1_2_87 ( .A(u4_sll_454_ML_int_2__87_), .B(
        u4_sll_454_ML_int_2__83_), .S(u4_sll_454_net66663), .Z(
        u4_sll_454_ML_int_3__87_) );
  MUX2_X2 u4_sll_454_M1_2_88 ( .A(u4_sll_454_ML_int_2__88_), .B(
        u4_sll_454_ML_int_2__84_), .S(u4_sll_454_net66667), .Z(
        u4_sll_454_ML_int_3__88_) );
  MUX2_X2 u4_sll_454_M1_2_89 ( .A(u4_sll_454_ML_int_2__89_), .B(
        u4_sll_454_ML_int_2__85_), .S(u4_sll_454_net66667), .Z(
        u4_sll_454_ML_int_3__89_) );
  MUX2_X2 u4_sll_454_M1_2_90 ( .A(u4_sll_454_ML_int_2__90_), .B(
        u4_sll_454_ML_int_2__86_), .S(u4_sll_454_net66667), .Z(
        u4_sll_454_ML_int_3__90_) );
  MUX2_X2 u4_sll_454_M1_2_91 ( .A(u4_sll_454_ML_int_2__91_), .B(
        u4_sll_454_ML_int_2__87_), .S(u4_sll_454_net66667), .Z(
        u4_sll_454_ML_int_3__91_) );
  MUX2_X2 u4_sll_454_M1_2_92 ( .A(u4_sll_454_ML_int_2__92_), .B(
        u4_sll_454_ML_int_2__88_), .S(u4_sll_454_net66667), .Z(
        u4_sll_454_ML_int_3__92_) );
  MUX2_X2 u4_sll_454_M1_2_93 ( .A(u4_sll_454_ML_int_2__93_), .B(
        u4_sll_454_ML_int_2__89_), .S(u4_sll_454_net66667), .Z(
        u4_sll_454_ML_int_3__93_) );
  MUX2_X2 u4_sll_454_M1_2_94 ( .A(u4_sll_454_ML_int_2__94_), .B(
        u4_sll_454_ML_int_2__90_), .S(u4_sll_454_net66667), .Z(
        u4_sll_454_ML_int_3__94_) );
  MUX2_X2 u4_sll_454_M1_2_95 ( .A(u4_sll_454_ML_int_2__95_), .B(
        u4_sll_454_ML_int_2__91_), .S(u4_sll_454_net66667), .Z(
        u4_sll_454_ML_int_3__95_) );
  MUX2_X2 u4_sll_454_M1_2_96 ( .A(u4_sll_454_ML_int_2__96_), .B(
        u4_sll_454_ML_int_2__92_), .S(u4_sll_454_net66667), .Z(
        u4_sll_454_ML_int_3__96_) );
  MUX2_X2 u4_sll_454_M1_2_97 ( .A(u4_sll_454_ML_int_2__97_), .B(
        u4_sll_454_ML_int_2__93_), .S(u4_sll_454_net66667), .Z(
        u4_sll_454_ML_int_3__97_) );
  MUX2_X2 u4_sll_454_M1_2_98 ( .A(u4_sll_454_ML_int_2__98_), .B(
        u4_sll_454_ML_int_2__94_), .S(u4_sll_454_net66667), .Z(
        u4_sll_454_ML_int_3__98_) );
  MUX2_X2 u4_sll_454_M1_2_99 ( .A(u4_sll_454_ML_int_2__99_), .B(
        u4_sll_454_ML_int_2__95_), .S(u4_sll_454_net66667), .Z(
        u4_sll_454_ML_int_3__99_) );
  MUX2_X2 u4_sll_454_M1_2_100 ( .A(u4_sll_454_ML_int_2__100_), .B(
        u4_sll_454_ML_int_2__96_), .S(u4_sll_454_net66667), .Z(
        u4_sll_454_ML_int_3__100_) );
  MUX2_X2 u4_sll_454_M1_2_101 ( .A(u4_sll_454_ML_int_2__101_), .B(
        u4_sll_454_ML_int_2__97_), .S(u4_sll_454_net66667), .Z(
        u4_sll_454_ML_int_3__101_) );
  MUX2_X2 u4_sll_454_M1_2_102 ( .A(u4_sll_454_ML_int_2__102_), .B(
        u4_sll_454_ML_int_2__98_), .S(u4_sll_454_net66667), .Z(
        u4_sll_454_ML_int_3__102_) );
  MUX2_X2 u4_sll_454_M1_2_103 ( .A(u4_sll_454_ML_int_2__103_), .B(
        u4_sll_454_ML_int_2__99_), .S(u4_sll_454_net66667), .Z(
        u4_sll_454_ML_int_3__103_) );
  MUX2_X2 u4_sll_454_M1_2_104 ( .A(u4_sll_454_ML_int_2__104_), .B(
        u4_sll_454_ML_int_2__100_), .S(u4_sll_454_net66667), .Z(
        u4_sll_454_ML_int_3__104_) );
  MUX2_X2 u4_sll_454_M1_2_105 ( .A(u4_sll_454_ML_int_2__105_), .B(
        u4_sll_454_ML_int_2__101_), .S(u4_sll_454_net66667), .Z(
        u4_sll_454_ML_int_3__105_) );
  MUX2_X2 u4_sll_454_M1_3_8 ( .A(u4_sll_454_ML_int_3__8_), .B(
        u4_sll_454_ML_int_3__0_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__8_) );
  MUX2_X2 u4_sll_454_M1_3_9 ( .A(u4_sll_454_ML_int_3__9_), .B(
        u4_sll_454_ML_int_3__1_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__9_) );
  MUX2_X2 u4_sll_454_M1_3_10 ( .A(u4_sll_454_ML_int_3__10_), .B(
        u4_sll_454_ML_int_3__2_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__10_) );
  MUX2_X2 u4_sll_454_M1_3_11 ( .A(u4_sll_454_ML_int_3__11_), .B(
        u4_sll_454_ML_int_3__3_), .S(u4_sll_454_net66611), .Z(
        u4_sll_454_ML_int_4__11_) );
  MUX2_X2 u4_sll_454_M1_3_12 ( .A(u4_sll_454_ML_int_3__12_), .B(
        u4_sll_454_ML_int_3__4_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__12_) );
  MUX2_X2 u4_sll_454_M1_3_13 ( .A(u4_sll_454_ML_int_3__13_), .B(
        u4_sll_454_ML_int_3__5_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__13_) );
  MUX2_X2 u4_sll_454_M1_3_14 ( .A(u4_sll_454_ML_int_3__14_), .B(
        u4_sll_454_ML_int_3__6_), .S(u4_sll_454_net66611), .Z(
        u4_sll_454_ML_int_4__14_) );
  MUX2_X2 u4_sll_454_M1_3_15 ( .A(u4_sll_454_ML_int_3__15_), .B(
        u4_sll_454_ML_int_3__7_), .S(u4_sll_454_net66611), .Z(
        u4_sll_454_ML_int_4__15_) );
  MUX2_X2 u4_sll_454_M1_3_16 ( .A(u4_sll_454_ML_int_3__16_), .B(
        u4_sll_454_ML_int_3__8_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__16_) );
  MUX2_X2 u4_sll_454_M1_3_17 ( .A(u4_sll_454_ML_int_3__17_), .B(
        u4_sll_454_ML_int_3__9_), .S(u4_sll_454_net66611), .Z(
        u4_sll_454_ML_int_4__17_) );
  MUX2_X2 u4_sll_454_M1_3_18 ( .A(u4_sll_454_ML_int_3__18_), .B(
        u4_sll_454_ML_int_3__10_), .S(u4_sll_454_net66611), .Z(
        u4_sll_454_ML_int_4__18_) );
  MUX2_X2 u4_sll_454_M1_3_19 ( .A(u4_sll_454_ML_int_3__19_), .B(
        u4_sll_454_ML_int_3__11_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__19_) );
  MUX2_X2 u4_sll_454_M1_3_21 ( .A(u4_sll_454_ML_int_3__21_), .B(
        u4_sll_454_ML_int_3__13_), .S(u4_sll_454_net66611), .Z(
        u4_sll_454_ML_int_4__21_) );
  MUX2_X2 u4_sll_454_M1_3_22 ( .A(u4_sll_454_ML_int_3__22_), .B(
        u4_sll_454_ML_int_3__14_), .S(u4_sll_454_net66599), .Z(
        u4_sll_454_ML_int_4__22_) );
  MUX2_X2 u4_sll_454_M1_3_23 ( .A(u4_sll_454_ML_int_3__23_), .B(
        u4_sll_454_ML_int_3__15_), .S(u4_sll_454_net66599), .Z(
        u4_sll_454_ML_int_4__23_) );
  MUX2_X2 u4_sll_454_M1_3_24 ( .A(u4_sll_454_ML_int_3__24_), .B(
        u4_sll_454_ML_int_3__16_), .S(u4_sll_454_net66599), .Z(
        u4_sll_454_ML_int_4__24_) );
  MUX2_X2 u4_sll_454_M1_3_25 ( .A(u4_sll_454_ML_int_3__25_), .B(
        u4_sll_454_ML_int_3__17_), .S(u4_sll_454_net66599), .Z(
        u4_sll_454_ML_int_4__25_) );
  MUX2_X2 u4_sll_454_M1_3_26 ( .A(u4_sll_454_ML_int_3__26_), .B(
        u4_sll_454_ML_int_3__18_), .S(u4_sll_454_net66599), .Z(
        u4_sll_454_ML_int_4__26_) );
  MUX2_X2 u4_sll_454_M1_3_27 ( .A(u4_sll_454_ML_int_3__27_), .B(
        u4_sll_454_ML_int_3__19_), .S(u4_sll_454_net66599), .Z(
        u4_sll_454_ML_int_4__27_) );
  MUX2_X2 u4_sll_454_M1_3_29 ( .A(u4_sll_454_ML_int_3__29_), .B(
        u4_sll_454_ML_int_3__21_), .S(u4_sll_454_net66599), .Z(
        u4_sll_454_ML_int_4__29_) );
  MUX2_X2 u4_sll_454_M1_3_30 ( .A(u4_sll_454_ML_int_3__30_), .B(
        u4_sll_454_ML_int_3__22_), .S(u4_sll_454_net66599), .Z(
        u4_sll_454_ML_int_4__30_) );
  MUX2_X2 u4_sll_454_M1_3_31 ( .A(u4_sll_454_ML_int_3__31_), .B(
        u4_sll_454_ML_int_3__23_), .S(u4_sll_454_net66599), .Z(
        u4_sll_454_ML_int_4__31_) );
  MUX2_X2 u4_sll_454_M1_3_32 ( .A(u4_sll_454_ML_int_3__32_), .B(
        u4_sll_454_ML_int_3__24_), .S(u4_sll_454_net66599), .Z(
        u4_sll_454_ML_int_4__32_) );
  MUX2_X2 u4_sll_454_M1_3_33 ( .A(u4_sll_454_ML_int_3__33_), .B(
        u4_sll_454_ML_int_3__25_), .S(u4_sll_454_net66601), .Z(
        u4_sll_454_ML_int_4__33_) );
  MUX2_X2 u4_sll_454_M1_3_34 ( .A(u4_sll_454_ML_int_3__34_), .B(
        u4_sll_454_ML_int_3__26_), .S(u4_sll_454_net66601), .Z(
        u4_sll_454_ML_int_4__34_) );
  MUX2_X2 u4_sll_454_M1_3_35 ( .A(u4_sll_454_ML_int_3__35_), .B(
        u4_sll_454_ML_int_3__27_), .S(u4_sll_454_net66601), .Z(
        u4_sll_454_ML_int_4__35_) );
  MUX2_X2 u4_sll_454_M1_3_37 ( .A(u4_sll_454_ML_int_3__37_), .B(
        u4_sll_454_ML_int_3__29_), .S(u4_sll_454_net66601), .Z(
        u4_sll_454_ML_int_4__37_) );
  MUX2_X2 u4_sll_454_M1_3_38 ( .A(u4_sll_454_ML_int_3__38_), .B(
        u4_sll_454_ML_int_3__30_), .S(u4_sll_454_net66601), .Z(
        u4_sll_454_ML_int_4__38_) );
  MUX2_X2 u4_sll_454_M1_3_39 ( .A(u4_sll_454_ML_int_3__39_), .B(
        u4_sll_454_ML_int_3__31_), .S(u4_sll_454_net66601), .Z(
        u4_sll_454_ML_int_4__39_) );
  MUX2_X2 u4_sll_454_M1_3_40 ( .A(u4_sll_454_ML_int_3__40_), .B(
        u4_sll_454_ML_int_3__32_), .S(u4_sll_454_net66601), .Z(
        u4_sll_454_ML_int_4__40_) );
  MUX2_X2 u4_sll_454_M1_3_41 ( .A(u4_sll_454_ML_int_3__41_), .B(
        u4_sll_454_ML_int_3__33_), .S(u4_sll_454_net66601), .Z(
        u4_sll_454_ML_int_4__41_) );
  MUX2_X2 u4_sll_454_M1_3_42 ( .A(u4_sll_454_ML_int_3__42_), .B(
        u4_sll_454_ML_int_3__34_), .S(u4_sll_454_net66601), .Z(
        u4_sll_454_ML_int_4__42_) );
  MUX2_X2 u4_sll_454_M1_3_43 ( .A(u4_sll_454_ML_int_3__43_), .B(
        u4_sll_454_ML_int_3__35_), .S(u4_sll_454_net66601), .Z(
        u4_sll_454_ML_int_4__43_) );
  MUX2_X2 u4_sll_454_M1_3_45 ( .A(u4_sll_454_ML_int_3__45_), .B(
        u4_sll_454_ML_int_3__37_), .S(u4_sll_454_net66603), .Z(
        u4_sll_454_ML_int_4__45_) );
  MUX2_X2 u4_sll_454_M1_3_46 ( .A(u4_sll_454_ML_int_3__46_), .B(
        u4_sll_454_ML_int_3__38_), .S(u4_sll_454_net66603), .Z(
        u4_sll_454_ML_int_4__46_) );
  MUX2_X2 u4_sll_454_M1_3_47 ( .A(u4_sll_454_ML_int_3__47_), .B(
        u4_sll_454_ML_int_3__39_), .S(u4_sll_454_net66603), .Z(
        u4_sll_454_ML_int_4__47_) );
  MUX2_X2 u4_sll_454_M1_3_48 ( .A(u4_sll_454_ML_int_3__48_), .B(
        u4_sll_454_ML_int_3__40_), .S(u4_sll_454_net66603), .Z(
        u4_sll_454_ML_int_4__48_) );
  MUX2_X2 u4_sll_454_M1_3_49 ( .A(u4_sll_454_ML_int_3__49_), .B(
        u4_sll_454_ML_int_3__41_), .S(u4_sll_454_net66603), .Z(
        u4_sll_454_ML_int_4__49_) );
  MUX2_X2 u4_sll_454_M1_3_50 ( .A(u4_sll_454_ML_int_3__50_), .B(
        u4_sll_454_ML_int_3__42_), .S(u4_sll_454_net66603), .Z(
        u4_sll_454_ML_int_4__50_) );
  MUX2_X2 u4_sll_454_M1_3_51 ( .A(u4_sll_454_ML_int_3__51_), .B(
        u4_sll_454_ML_int_3__43_), .S(u4_sll_454_net66603), .Z(
        u4_sll_454_ML_int_4__51_) );
  MUX2_X2 u4_sll_454_M1_3_52 ( .A(u4_sll_454_ML_int_3__52_), .B(
        u4_sll_454_ML_int_3__44_), .S(u4_sll_454_net66603), .Z(
        u4_sll_454_ML_int_4__52_) );
  MUX2_X2 u4_sll_454_M1_3_53 ( .A(u4_sll_454_ML_int_3__53_), .B(
        u4_sll_454_ML_int_3__45_), .S(u4_sll_454_net66603), .Z(
        u4_sll_454_ML_int_4__53_) );
  MUX2_X2 u4_sll_454_M1_3_54 ( .A(u4_sll_454_ML_int_3__54_), .B(
        u4_sll_454_ML_int_3__46_), .S(u4_sll_454_net66603), .Z(
        u4_sll_454_ML_int_4__54_) );
  MUX2_X2 u4_sll_454_M1_3_55 ( .A(u4_sll_454_ML_int_3__55_), .B(
        u4_sll_454_ML_int_3__47_), .S(u4_sll_454_net66611), .Z(
        u4_sll_454_ML_int_4__55_) );
  MUX2_X2 u4_sll_454_M1_3_56 ( .A(u4_sll_454_ML_int_3__56_), .B(
        u4_sll_454_ML_int_3__48_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__56_) );
  MUX2_X2 u4_sll_454_M1_3_57 ( .A(u4_sll_454_ML_int_3__57_), .B(
        u4_sll_454_ML_int_3__49_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__57_) );
  MUX2_X2 u4_sll_454_M1_3_58 ( .A(u4_sll_454_ML_int_3__58_), .B(
        u4_sll_454_ML_int_3__50_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__58_) );
  MUX2_X2 u4_sll_454_M1_3_59 ( .A(u4_sll_454_ML_int_3__59_), .B(
        u4_sll_454_ML_int_3__51_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__59_) );
  MUX2_X2 u4_sll_454_M1_3_60 ( .A(u4_sll_454_ML_int_3__60_), .B(
        u4_sll_454_ML_int_3__52_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__60_) );
  MUX2_X2 u4_sll_454_M1_3_61 ( .A(u4_sll_454_ML_int_3__61_), .B(
        u4_sll_454_ML_int_3__53_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__61_) );
  MUX2_X2 u4_sll_454_M1_3_62 ( .A(u4_sll_454_ML_int_3__62_), .B(
        u4_sll_454_ML_int_3__54_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__62_) );
  MUX2_X2 u4_sll_454_M1_3_63 ( .A(u4_sll_454_ML_int_3__63_), .B(
        u4_sll_454_ML_int_3__55_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__63_) );
  MUX2_X2 u4_sll_454_M1_3_64 ( .A(u4_sll_454_ML_int_3__64_), .B(
        u4_sll_454_ML_int_3__56_), .S(u4_sll_454_net66609), .Z(
        u4_sll_454_ML_int_4__64_) );
  MUX2_X2 u4_sll_454_M1_3_65 ( .A(u4_sll_454_ML_int_3__65_), .B(
        u4_sll_454_ML_int_3__57_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__65_) );
  MUX2_X2 u4_sll_454_M1_3_66 ( .A(u4_sll_454_ML_int_3__66_), .B(
        u4_sll_454_ML_int_3__58_), .S(u4_sll_454_net66607), .Z(
        u4_sll_454_ML_int_4__66_) );
  MUX2_X2 u4_sll_454_M1_3_67 ( .A(u4_sll_454_ML_int_3__67_), .B(
        u4_sll_454_ML_int_3__59_), .S(u4_sll_454_net66607), .Z(
        u4_sll_454_ML_int_4__67_) );
  MUX2_X2 u4_sll_454_M1_3_68 ( .A(u4_sll_454_ML_int_3__68_), .B(
        u4_sll_454_ML_int_3__60_), .S(u4_sll_454_net66607), .Z(
        u4_sll_454_ML_int_4__68_) );
  MUX2_X2 u4_sll_454_M1_3_69 ( .A(u4_sll_454_ML_int_3__69_), .B(
        u4_sll_454_ML_int_3__61_), .S(u4_sll_454_net66607), .Z(
        u4_sll_454_ML_int_4__69_) );
  MUX2_X2 u4_sll_454_M1_3_70 ( .A(u4_sll_454_ML_int_3__70_), .B(
        u4_sll_454_ML_int_3__62_), .S(u4_sll_454_net66607), .Z(
        u4_sll_454_ML_int_4__70_) );
  MUX2_X2 u4_sll_454_M1_3_71 ( .A(u4_sll_454_ML_int_3__71_), .B(
        u4_sll_454_ML_int_3__63_), .S(u4_sll_454_net66607), .Z(
        u4_sll_454_ML_int_4__71_) );
  MUX2_X2 u4_sll_454_M1_3_72 ( .A(u4_sll_454_ML_int_3__72_), .B(
        u4_sll_454_ML_int_3__64_), .S(u4_sll_454_net66607), .Z(
        u4_sll_454_ML_int_4__72_) );
  MUX2_X2 u4_sll_454_M1_3_73 ( .A(u4_sll_454_ML_int_3__73_), .B(
        u4_sll_454_ML_int_3__65_), .S(u4_sll_454_net66607), .Z(
        u4_sll_454_ML_int_4__73_) );
  MUX2_X2 u4_sll_454_M1_3_74 ( .A(u4_sll_454_ML_int_3__74_), .B(
        u4_sll_454_ML_int_3__66_), .S(u4_sll_454_net66607), .Z(
        u4_sll_454_ML_int_4__74_) );
  MUX2_X2 u4_sll_454_M1_3_75 ( .A(u4_sll_454_ML_int_3__75_), .B(
        u4_sll_454_ML_int_3__67_), .S(u4_sll_454_net66607), .Z(
        u4_sll_454_ML_int_4__75_) );
  MUX2_X2 u4_sll_454_M1_3_76 ( .A(u4_sll_454_ML_int_3__76_), .B(
        u4_sll_454_ML_int_3__68_), .S(u4_sll_454_net66607), .Z(
        u4_sll_454_ML_int_4__76_) );
  MUX2_X2 u4_sll_454_M1_3_77 ( .A(u4_sll_454_ML_int_3__77_), .B(
        u4_sll_454_ML_int_3__69_), .S(u4_sll_454_net66609), .Z(
        u4_sll_454_ML_int_4__77_) );
  MUX2_X2 u4_sll_454_M1_3_78 ( .A(u4_sll_454_ML_int_3__78_), .B(
        u4_sll_454_ML_int_3__70_), .S(u4_sll_454_net66609), .Z(
        u4_sll_454_ML_int_4__78_) );
  MUX2_X2 u4_sll_454_M1_3_79 ( .A(u4_sll_454_ML_int_3__79_), .B(
        u4_sll_454_ML_int_3__71_), .S(u4_sll_454_net66609), .Z(
        u4_sll_454_ML_int_4__79_) );
  MUX2_X2 u4_sll_454_M1_3_80 ( .A(u4_sll_454_ML_int_3__80_), .B(
        u4_sll_454_ML_int_3__72_), .S(u4_sll_454_net66609), .Z(
        u4_sll_454_ML_int_4__80_) );
  MUX2_X2 u4_sll_454_M1_3_81 ( .A(u4_sll_454_ML_int_3__81_), .B(
        u4_sll_454_ML_int_3__73_), .S(u4_sll_454_net66609), .Z(
        u4_sll_454_ML_int_4__81_) );
  MUX2_X2 u4_sll_454_M1_3_82 ( .A(u4_sll_454_ML_int_3__82_), .B(
        u4_sll_454_ML_int_3__74_), .S(u4_sll_454_net66609), .Z(
        u4_sll_454_ML_int_4__82_) );
  MUX2_X2 u4_sll_454_M1_3_83 ( .A(u4_sll_454_ML_int_3__83_), .B(
        u4_sll_454_ML_int_3__75_), .S(u4_sll_454_net66609), .Z(
        u4_sll_454_ML_int_4__83_) );
  MUX2_X2 u4_sll_454_M1_3_84 ( .A(u4_sll_454_ML_int_3__84_), .B(
        u4_sll_454_ML_int_3__76_), .S(u4_sll_454_net66609), .Z(
        u4_sll_454_ML_int_4__84_) );
  MUX2_X2 u4_sll_454_M1_3_85 ( .A(u4_sll_454_ML_int_3__85_), .B(
        u4_sll_454_ML_int_3__77_), .S(u4_sll_454_net66609), .Z(
        u4_sll_454_ML_int_4__85_) );
  MUX2_X2 u4_sll_454_M1_3_86 ( .A(u4_sll_454_ML_int_3__86_), .B(
        u4_sll_454_ML_int_3__78_), .S(u4_sll_454_net66609), .Z(
        u4_sll_454_ML_int_4__86_) );
  MUX2_X2 u4_sll_454_M1_3_87 ( .A(u4_sll_454_ML_int_3__87_), .B(
        u4_sll_454_ML_int_3__79_), .S(u4_sll_454_net66609), .Z(
        u4_sll_454_ML_int_4__87_) );
  MUX2_X2 u4_sll_454_M1_3_88 ( .A(u4_sll_454_ML_int_3__88_), .B(
        u4_sll_454_ML_int_3__80_), .S(u4_sll_454_net66611), .Z(
        u4_sll_454_ML_int_4__88_) );
  MUX2_X2 u4_sll_454_M1_3_89 ( .A(u4_sll_454_ML_int_3__89_), .B(
        u4_sll_454_ML_int_3__81_), .S(u4_sll_454_net66611), .Z(
        u4_sll_454_ML_int_4__89_) );
  MUX2_X2 u4_sll_454_M1_3_90 ( .A(u4_sll_454_ML_int_3__90_), .B(
        u4_sll_454_ML_int_3__82_), .S(u4_sll_454_net66611), .Z(
        u4_sll_454_ML_int_4__90_) );
  MUX2_X2 u4_sll_454_M1_3_91 ( .A(u4_sll_454_ML_int_3__91_), .B(
        u4_sll_454_ML_int_3__83_), .S(u4_sll_454_net66611), .Z(
        u4_sll_454_ML_int_4__91_) );
  MUX2_X2 u4_sll_454_M1_3_92 ( .A(u4_sll_454_ML_int_3__92_), .B(
        u4_sll_454_ML_int_3__84_), .S(u4_sll_454_net66611), .Z(
        u4_sll_454_ML_int_4__92_) );
  MUX2_X2 u4_sll_454_M1_3_93 ( .A(u4_sll_454_ML_int_3__93_), .B(
        u4_sll_454_ML_int_3__85_), .S(u4_sll_454_net66611), .Z(
        u4_sll_454_ML_int_4__93_) );
  MUX2_X2 u4_sll_454_M1_3_94 ( .A(u4_sll_454_ML_int_3__94_), .B(
        u4_sll_454_ML_int_3__86_), .S(u4_sll_454_net66611), .Z(
        u4_sll_454_ML_int_4__94_) );
  MUX2_X2 u4_sll_454_M1_3_95 ( .A(u4_sll_454_ML_int_3__95_), .B(
        u4_sll_454_ML_int_3__87_), .S(u4_sll_454_net66611), .Z(
        u4_sll_454_ML_int_4__95_) );
  MUX2_X2 u4_sll_454_M1_3_96 ( .A(u4_sll_454_ML_int_3__96_), .B(
        u4_sll_454_ML_int_3__88_), .S(u4_sll_454_net66611), .Z(
        u4_sll_454_ML_int_4__96_) );
  MUX2_X2 u4_sll_454_M1_3_97 ( .A(u4_sll_454_ML_int_3__97_), .B(
        u4_sll_454_ML_int_3__89_), .S(u4_sll_454_net66611), .Z(
        u4_sll_454_ML_int_4__97_) );
  MUX2_X2 u4_sll_454_M1_3_98 ( .A(u4_sll_454_ML_int_3__98_), .B(
        u4_sll_454_ML_int_3__90_), .S(u4_sll_454_net66611), .Z(
        u4_sll_454_ML_int_4__98_) );
  MUX2_X2 u4_sll_454_M1_3_99 ( .A(u4_sll_454_ML_int_3__99_), .B(
        u4_sll_454_ML_int_3__91_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__99_) );
  MUX2_X2 u4_sll_454_M1_3_100 ( .A(u4_sll_454_ML_int_3__100_), .B(
        u4_sll_454_ML_int_3__92_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__100_) );
  MUX2_X2 u4_sll_454_M1_3_101 ( .A(u4_sll_454_ML_int_3__101_), .B(
        u4_sll_454_ML_int_3__93_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__101_) );
  MUX2_X2 u4_sll_454_M1_3_102 ( .A(u4_sll_454_ML_int_3__102_), .B(
        u4_sll_454_ML_int_3__94_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__102_) );
  MUX2_X2 u4_sll_454_M1_3_103 ( .A(u4_sll_454_ML_int_3__103_), .B(
        u4_sll_454_ML_int_3__95_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__103_) );
  MUX2_X2 u4_sll_454_M1_3_104 ( .A(u4_sll_454_ML_int_3__104_), .B(
        u4_sll_454_ML_int_3__96_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__104_) );
  MUX2_X2 u4_sll_454_M1_3_105 ( .A(u4_sll_454_ML_int_3__105_), .B(
        u4_sll_454_ML_int_3__97_), .S(u4_sll_454_net66613), .Z(
        u4_sll_454_ML_int_4__105_) );
  MUX2_X2 u4_sll_454_M1_4_16 ( .A(u4_sll_454_ML_int_4__16_), .B(
        u4_sll_454_ML_int_4__0_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__16_) );
  MUX2_X2 u4_sll_454_M1_4_17 ( .A(u4_sll_454_ML_int_4__17_), .B(
        u4_sll_454_ML_int_4__1_), .S(u4_sll_454_net66555), .Z(
        u4_sll_454_ML_int_5__17_) );
  MUX2_X2 u4_sll_454_M1_4_18 ( .A(u4_sll_454_ML_int_4__18_), .B(
        u4_sll_454_ML_int_4__2_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__18_) );
  MUX2_X2 u4_sll_454_M1_4_19 ( .A(u4_sll_454_ML_int_4__19_), .B(
        u4_sll_454_ML_int_4__3_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__19_) );
  MUX2_X2 u4_sll_454_M1_4_20 ( .A(u4_sll_454_ML_int_4__20_), .B(
        u4_sll_454_ML_int_4__4_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__20_) );
  MUX2_X2 u4_sll_454_M1_4_21 ( .A(u4_sll_454_ML_int_4__21_), .B(
        u4_sll_454_ML_int_4__5_), .S(u4_sll_454_net66551), .Z(
        u4_sll_454_ML_int_5__21_) );
  MUX2_X2 u4_sll_454_M1_4_22 ( .A(u4_sll_454_ML_int_4__22_), .B(
        u4_sll_454_ML_int_4__6_), .S(u4_sll_454_net66555), .Z(
        u4_sll_454_ML_int_5__22_) );
  MUX2_X2 u4_sll_454_M1_4_23 ( .A(u4_sll_454_ML_int_4__23_), .B(
        u4_sll_454_ML_int_4__7_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__23_) );
  MUX2_X2 u4_sll_454_M1_4_24 ( .A(u4_sll_454_ML_int_4__24_), .B(
        u4_sll_454_ML_int_4__8_), .S(u4_sll_454_net66555), .Z(
        u4_sll_454_ML_int_5__24_) );
  MUX2_X2 u4_sll_454_M1_4_25 ( .A(u4_sll_454_ML_int_4__25_), .B(
        u4_sll_454_ML_int_4__9_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__25_) );
  MUX2_X2 u4_sll_454_M1_4_26 ( .A(u4_sll_454_ML_int_4__26_), .B(
        u4_sll_454_ML_int_4__10_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__26_) );
  MUX2_X2 u4_sll_454_M1_4_27 ( .A(u4_sll_454_ML_int_4__27_), .B(
        u4_sll_454_ML_int_4__11_), .S(u4_sll_454_net66555), .Z(
        u4_sll_454_ML_int_5__27_) );
  MUX2_X2 u4_sll_454_M1_4_29 ( .A(u4_sll_454_ML_int_4__29_), .B(
        u4_sll_454_ML_int_4__13_), .S(u4_sll_454_net66555), .Z(
        u4_sll_454_ML_int_5__29_) );
  MUX2_X2 u4_sll_454_M1_4_30 ( .A(u4_sll_454_ML_int_4__30_), .B(
        u4_sll_454_ML_int_4__14_), .S(u4_sll_454_net66555), .Z(
        u4_sll_454_ML_int_5__30_) );
  MUX2_X2 u4_sll_454_M1_4_31 ( .A(u4_sll_454_ML_int_4__31_), .B(
        u4_sll_454_ML_int_4__15_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__31_) );
  MUX2_X2 u4_sll_454_M1_4_32 ( .A(u4_sll_454_ML_int_4__32_), .B(
        u4_sll_454_ML_int_4__16_), .S(u4_sll_454_net66555), .Z(
        u4_sll_454_ML_int_5__32_) );
  MUX2_X2 u4_sll_454_M1_4_33 ( .A(u4_sll_454_ML_int_4__33_), .B(
        u4_sll_454_ML_int_4__17_), .S(u4_sll_454_net66545), .Z(
        u4_sll_454_ML_int_5__33_) );
  MUX2_X2 u4_sll_454_M1_4_34 ( .A(u4_sll_454_ML_int_4__34_), .B(
        u4_sll_454_ML_int_4__18_), .S(u4_sll_454_net66545), .Z(
        u4_sll_454_ML_int_5__34_) );
  MUX2_X2 u4_sll_454_M1_4_35 ( .A(u4_sll_454_ML_int_4__35_), .B(
        u4_sll_454_ML_int_4__19_), .S(u4_sll_454_net66545), .Z(
        u4_sll_454_ML_int_5__35_) );
  MUX2_X2 u4_sll_454_M1_4_36 ( .A(u4_sll_454_ML_int_4__36_), .B(
        u4_sll_454_ML_int_4__20_), .S(u4_sll_454_net66545), .Z(
        u4_sll_454_ML_int_5__36_) );
  MUX2_X2 u4_sll_454_M1_4_37 ( .A(u4_sll_454_ML_int_4__37_), .B(
        u4_sll_454_ML_int_4__21_), .S(u4_sll_454_net66545), .Z(
        u4_sll_454_ML_int_5__37_) );
  MUX2_X2 u4_sll_454_M1_4_38 ( .A(u4_sll_454_ML_int_4__38_), .B(
        u4_sll_454_ML_int_4__22_), .S(u4_sll_454_net66545), .Z(
        u4_sll_454_ML_int_5__38_) );
  MUX2_X2 u4_sll_454_M1_4_39 ( .A(u4_sll_454_ML_int_4__39_), .B(
        u4_sll_454_ML_int_4__23_), .S(u4_sll_454_net66545), .Z(
        u4_sll_454_ML_int_5__39_) );
  MUX2_X2 u4_sll_454_M1_4_40 ( .A(u4_sll_454_ML_int_4__40_), .B(
        u4_sll_454_ML_int_4__24_), .S(u4_sll_454_net66545), .Z(
        u4_sll_454_ML_int_5__40_) );
  MUX2_X2 u4_sll_454_M1_4_41 ( .A(u4_sll_454_ML_int_4__41_), .B(
        u4_sll_454_ML_int_4__25_), .S(u4_sll_454_net66545), .Z(
        u4_sll_454_ML_int_5__41_) );
  MUX2_X2 u4_sll_454_M1_4_42 ( .A(u4_sll_454_ML_int_4__42_), .B(
        u4_sll_454_ML_int_4__26_), .S(u4_sll_454_net66545), .Z(
        u4_sll_454_ML_int_5__42_) );
  MUX2_X2 u4_sll_454_M1_4_43 ( .A(u4_sll_454_ML_int_4__43_), .B(
        u4_sll_454_ML_int_4__27_), .S(u4_sll_454_net66545), .Z(
        u4_sll_454_ML_int_5__43_) );
  MUX2_X2 u4_sll_454_M1_4_45 ( .A(u4_sll_454_ML_int_4__45_), .B(
        u4_sll_454_ML_int_4__29_), .S(u4_sll_454_net66547), .Z(
        u4_sll_454_ML_int_5__45_) );
  MUX2_X2 u4_sll_454_M1_4_46 ( .A(u4_sll_454_ML_int_4__46_), .B(
        u4_sll_454_ML_int_4__30_), .S(u4_sll_454_net66547), .Z(
        u4_sll_454_ML_int_5__46_) );
  MUX2_X2 u4_sll_454_M1_4_47 ( .A(u4_sll_454_ML_int_4__47_), .B(
        u4_sll_454_ML_int_4__31_), .S(u4_sll_454_net66547), .Z(
        u4_sll_454_ML_int_5__47_) );
  MUX2_X2 u4_sll_454_M1_4_48 ( .A(u4_sll_454_ML_int_4__48_), .B(
        u4_sll_454_ML_int_4__32_), .S(u4_sll_454_net66547), .Z(
        u4_sll_454_ML_int_5__48_) );
  MUX2_X2 u4_sll_454_M1_4_49 ( .A(u4_sll_454_ML_int_4__49_), .B(
        u4_sll_454_ML_int_4__33_), .S(u4_sll_454_net66547), .Z(
        u4_sll_454_ML_int_5__49_) );
  MUX2_X2 u4_sll_454_M1_4_50 ( .A(u4_sll_454_ML_int_4__50_), .B(
        u4_sll_454_ML_int_4__34_), .S(u4_sll_454_net66547), .Z(
        u4_sll_454_ML_int_5__50_) );
  MUX2_X2 u4_sll_454_M1_4_51 ( .A(u4_sll_454_ML_int_4__51_), .B(
        u4_sll_454_ML_int_4__35_), .S(u4_sll_454_net66547), .Z(
        u4_sll_454_ML_int_5__51_) );
  MUX2_X2 u4_sll_454_M1_4_52 ( .A(u4_sll_454_ML_int_4__52_), .B(
        u4_sll_454_ML_int_4__36_), .S(u4_sll_454_net66547), .Z(
        u4_sll_454_ML_int_5__52_) );
  MUX2_X2 u4_sll_454_M1_4_53 ( .A(u4_sll_454_ML_int_4__53_), .B(
        u4_sll_454_ML_int_4__37_), .S(u4_sll_454_net66547), .Z(
        u4_sll_454_ML_int_5__53_) );
  MUX2_X2 u4_sll_454_M1_4_54 ( .A(u4_sll_454_ML_int_4__54_), .B(
        u4_sll_454_ML_int_4__38_), .S(u4_sll_454_net66547), .Z(
        u4_sll_454_ML_int_5__54_) );
  MUX2_X2 u4_sll_454_M1_4_55 ( .A(u4_sll_454_ML_int_4__55_), .B(
        u4_sll_454_ML_int_4__39_), .S(u4_sll_454_net66549), .Z(
        u4_sll_454_ML_int_5__55_) );
  MUX2_X2 u4_sll_454_M1_4_56 ( .A(u4_sll_454_ML_int_4__56_), .B(
        u4_sll_454_ML_int_4__40_), .S(u4_sll_454_net66549), .Z(
        u4_sll_454_ML_int_5__56_) );
  MUX2_X2 u4_sll_454_M1_4_57 ( .A(u4_sll_454_ML_int_4__57_), .B(
        u4_sll_454_ML_int_4__41_), .S(u4_sll_454_net66549), .Z(
        u4_sll_454_ML_int_5__57_) );
  MUX2_X2 u4_sll_454_M1_4_58 ( .A(u4_sll_454_ML_int_4__58_), .B(
        u4_sll_454_ML_int_4__42_), .S(u4_sll_454_net66549), .Z(
        u4_sll_454_ML_int_5__58_) );
  MUX2_X2 u4_sll_454_M1_4_59 ( .A(u4_sll_454_ML_int_4__59_), .B(
        u4_sll_454_ML_int_4__43_), .S(u4_sll_454_net66549), .Z(
        u4_sll_454_ML_int_5__59_) );
  MUX2_X2 u4_sll_454_M1_4_61 ( .A(u4_sll_454_ML_int_4__61_), .B(
        u4_sll_454_ML_int_4__45_), .S(u4_sll_454_net66549), .Z(
        u4_sll_454_ML_int_5__61_) );
  MUX2_X2 u4_sll_454_M1_4_62 ( .A(u4_sll_454_ML_int_4__62_), .B(
        u4_sll_454_ML_int_4__46_), .S(u4_sll_454_net66549), .Z(
        u4_sll_454_ML_int_5__62_) );
  MUX2_X2 u4_sll_454_M1_4_63 ( .A(u4_sll_454_ML_int_4__63_), .B(
        u4_sll_454_ML_int_4__47_), .S(u4_sll_454_net66549), .Z(
        u4_sll_454_ML_int_5__63_) );
  MUX2_X2 u4_sll_454_M1_4_64 ( .A(u4_sll_454_ML_int_4__64_), .B(
        u4_sll_454_ML_int_4__48_), .S(u4_sll_454_net66549), .Z(
        u4_sll_454_ML_int_5__64_) );
  MUX2_X2 u4_sll_454_M1_4_65 ( .A(u4_sll_454_ML_int_4__65_), .B(
        u4_sll_454_ML_int_4__49_), .S(u4_sll_454_net66549), .Z(
        u4_sll_454_ML_int_5__65_) );
  MUX2_X2 u4_sll_454_M1_4_66 ( .A(u4_sll_454_ML_int_4__66_), .B(
        u4_sll_454_ML_int_4__50_), .S(u4_sll_454_net66551), .Z(
        u4_sll_454_ML_int_5__66_) );
  MUX2_X2 u4_sll_454_M1_4_67 ( .A(u4_sll_454_ML_int_4__67_), .B(
        u4_sll_454_ML_int_4__51_), .S(u4_sll_454_net66551), .Z(
        u4_sll_454_ML_int_5__67_) );
  MUX2_X2 u4_sll_454_M1_4_68 ( .A(u4_sll_454_ML_int_4__68_), .B(
        u4_sll_454_ML_int_4__52_), .S(u4_sll_454_net66551), .Z(
        u4_sll_454_ML_int_5__68_) );
  MUX2_X2 u4_sll_454_M1_4_69 ( .A(u4_sll_454_ML_int_4__69_), .B(
        u4_sll_454_ML_int_4__53_), .S(u4_sll_454_net66551), .Z(
        u4_sll_454_ML_int_5__69_) );
  MUX2_X2 u4_sll_454_M1_4_70 ( .A(u4_sll_454_ML_int_4__70_), .B(
        u4_sll_454_ML_int_4__54_), .S(u4_sll_454_net66551), .Z(
        u4_sll_454_ML_int_5__70_) );
  MUX2_X2 u4_sll_454_M1_4_71 ( .A(u4_sll_454_ML_int_4__71_), .B(
        u4_sll_454_ML_int_4__55_), .S(u4_sll_454_net66551), .Z(
        u4_sll_454_ML_int_5__71_) );
  MUX2_X2 u4_sll_454_M1_4_72 ( .A(u4_sll_454_ML_int_4__72_), .B(
        u4_sll_454_ML_int_4__56_), .S(u4_sll_454_net66551), .Z(
        u4_sll_454_ML_int_5__72_) );
  MUX2_X2 u4_sll_454_M1_4_73 ( .A(u4_sll_454_ML_int_4__73_), .B(
        u4_sll_454_ML_int_4__57_), .S(u4_sll_454_net66551), .Z(
        u4_sll_454_ML_int_5__73_) );
  MUX2_X2 u4_sll_454_M1_4_74 ( .A(u4_sll_454_ML_int_4__74_), .B(
        u4_sll_454_ML_int_4__58_), .S(u4_sll_454_net66551), .Z(
        u4_sll_454_ML_int_5__74_) );
  MUX2_X2 u4_sll_454_M1_4_75 ( .A(u4_sll_454_ML_int_4__75_), .B(
        u4_sll_454_ML_int_4__59_), .S(u4_sll_454_net66551), .Z(
        u4_sll_454_ML_int_5__75_) );
  MUX2_X2 u4_sll_454_M1_4_76 ( .A(u4_sll_454_ML_int_4__76_), .B(
        u4_sll_454_ML_int_4__60_), .S(u4_sll_454_net66551), .Z(
        u4_sll_454_ML_int_5__76_) );
  MUX2_X2 u4_sll_454_M1_4_77 ( .A(u4_sll_454_ML_int_4__77_), .B(
        u4_sll_454_ML_int_4__61_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__77_) );
  MUX2_X2 u4_sll_454_M1_4_78 ( .A(u4_sll_454_ML_int_4__78_), .B(
        u4_sll_454_ML_int_4__62_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__78_) );
  MUX2_X2 u4_sll_454_M1_4_79 ( .A(u4_sll_454_ML_int_4__79_), .B(
        u4_sll_454_ML_int_4__63_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__79_) );
  MUX2_X2 u4_sll_454_M1_4_80 ( .A(u4_sll_454_ML_int_4__80_), .B(
        u4_sll_454_ML_int_4__64_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__80_) );
  MUX2_X2 u4_sll_454_M1_4_81 ( .A(u4_sll_454_ML_int_4__81_), .B(
        u4_sll_454_ML_int_4__65_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__81_) );
  MUX2_X2 u4_sll_454_M1_4_82 ( .A(u4_sll_454_ML_int_4__82_), .B(
        u4_sll_454_ML_int_4__66_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__82_) );
  MUX2_X2 u4_sll_454_M1_4_83 ( .A(u4_sll_454_ML_int_4__83_), .B(
        u4_sll_454_ML_int_4__67_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__83_) );
  MUX2_X2 u4_sll_454_M1_4_84 ( .A(u4_sll_454_ML_int_4__84_), .B(
        u4_sll_454_ML_int_4__68_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__84_) );
  MUX2_X2 u4_sll_454_M1_4_85 ( .A(u4_sll_454_ML_int_4__85_), .B(
        u4_sll_454_ML_int_4__69_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__85_) );
  MUX2_X2 u4_sll_454_M1_4_86 ( .A(u4_sll_454_ML_int_4__86_), .B(
        u4_sll_454_ML_int_4__70_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__86_) );
  MUX2_X2 u4_sll_454_M1_4_87 ( .A(u4_sll_454_ML_int_4__87_), .B(
        u4_sll_454_ML_int_4__71_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__87_) );
  MUX2_X2 u4_sll_454_M1_4_88 ( .A(u4_sll_454_ML_int_4__88_), .B(
        u4_sll_454_ML_int_4__72_), .S(u4_sll_454_net66555), .Z(
        u4_sll_454_ML_int_5__88_) );
  MUX2_X2 u4_sll_454_M1_4_89 ( .A(u4_sll_454_ML_int_4__89_), .B(
        u4_sll_454_ML_int_4__73_), .S(u4_sll_454_net66555), .Z(
        u4_sll_454_ML_int_5__89_) );
  MUX2_X2 u4_sll_454_M1_4_90 ( .A(u4_sll_454_ML_int_4__90_), .B(
        u4_sll_454_ML_int_4__74_), .S(u4_sll_454_net66555), .Z(
        u4_sll_454_ML_int_5__90_) );
  MUX2_X2 u4_sll_454_M1_4_91 ( .A(u4_sll_454_ML_int_4__91_), .B(
        u4_sll_454_ML_int_4__75_), .S(u4_sll_454_net66555), .Z(
        u4_sll_454_ML_int_5__91_) );
  MUX2_X2 u4_sll_454_M1_4_92 ( .A(u4_sll_454_ML_int_4__92_), .B(
        u4_sll_454_ML_int_4__76_), .S(u4_sll_454_net66555), .Z(
        u4_sll_454_ML_int_5__92_) );
  MUX2_X2 u4_sll_454_M1_4_93 ( .A(u4_sll_454_ML_int_4__93_), .B(
        u4_sll_454_ML_int_4__77_), .S(u4_sll_454_net66555), .Z(
        u4_sll_454_ML_int_5__93_) );
  MUX2_X2 u4_sll_454_M1_4_94 ( .A(u4_sll_454_ML_int_4__94_), .B(
        u4_sll_454_ML_int_4__78_), .S(u4_sll_454_net66555), .Z(
        u4_sll_454_ML_int_5__94_) );
  MUX2_X2 u4_sll_454_M1_4_95 ( .A(u4_sll_454_ML_int_4__95_), .B(
        u4_sll_454_ML_int_4__79_), .S(u4_sll_454_net66555), .Z(
        u4_sll_454_ML_int_5__95_) );
  MUX2_X2 u4_sll_454_M1_4_96 ( .A(u4_sll_454_ML_int_4__96_), .B(
        u4_sll_454_ML_int_4__80_), .S(u4_sll_454_net66555), .Z(
        u4_sll_454_ML_int_5__96_) );
  MUX2_X2 u4_sll_454_M1_4_97 ( .A(u4_sll_454_ML_int_4__97_), .B(
        u4_sll_454_ML_int_4__81_), .S(u4_sll_454_net66555), .Z(
        u4_sll_454_ML_int_5__97_) );
  MUX2_X2 u4_sll_454_M1_4_98 ( .A(u4_sll_454_ML_int_4__98_), .B(
        u4_sll_454_ML_int_4__82_), .S(u4_sll_454_net66555), .Z(
        u4_sll_454_ML_int_5__98_) );
  MUX2_X2 u4_sll_454_M1_4_99 ( .A(u4_sll_454_ML_int_4__99_), .B(
        u4_sll_454_ML_int_4__83_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__99_) );
  MUX2_X2 u4_sll_454_M1_4_100 ( .A(u4_sll_454_ML_int_4__100_), .B(
        u4_sll_454_ML_int_4__84_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__100_) );
  MUX2_X2 u4_sll_454_M1_4_101 ( .A(u4_sll_454_ML_int_4__101_), .B(
        u4_sll_454_ML_int_4__85_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__101_) );
  MUX2_X2 u4_sll_454_M1_4_102 ( .A(u4_sll_454_ML_int_4__102_), .B(
        u4_sll_454_ML_int_4__86_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__102_) );
  MUX2_X2 u4_sll_454_M1_4_103 ( .A(u4_sll_454_ML_int_4__103_), .B(
        u4_sll_454_ML_int_4__87_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__103_) );
  MUX2_X2 u4_sll_454_M1_4_104 ( .A(u4_sll_454_ML_int_4__104_), .B(
        u4_sll_454_ML_int_4__88_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__104_) );
  MUX2_X2 u4_sll_454_M1_4_105 ( .A(u4_sll_454_ML_int_4__105_), .B(
        u4_sll_454_ML_int_4__89_), .S(u4_sll_454_net66557), .Z(
        u4_sll_454_ML_int_5__105_) );
  MUX2_X2 u4_sll_454_M1_5_32 ( .A(u4_sll_454_ML_int_5__32_), .B(
        u4_sll_454_ML_int_5__0_), .S(u4_sll_454_net66487), .Z(
        u4_sll_454_ML_int_6__32_) );
  MUX2_X2 u4_sll_454_M1_5_33 ( .A(u4_sll_454_ML_int_5__33_), .B(
        u4_sll_454_ML_int_5__1_), .S(u4_sll_454_net66489), .Z(
        u4_sll_454_ML_int_6__33_) );
  MUX2_X2 u4_sll_454_M1_5_34 ( .A(u4_sll_454_ML_int_5__34_), .B(
        u4_sll_454_ML_int_5__2_), .S(u4_sll_454_net66489), .Z(
        u4_sll_454_ML_int_6__34_) );
  MUX2_X2 u4_sll_454_M1_5_35 ( .A(u4_sll_454_ML_int_5__35_), .B(
        u4_sll_454_ML_int_5__3_), .S(u4_sll_454_net66489), .Z(
        u4_sll_454_ML_int_6__35_) );
  MUX2_X2 u4_sll_454_M1_5_36 ( .A(u4_sll_454_ML_int_5__36_), .B(
        u4_sll_454_ML_int_5__4_), .S(u4_sll_454_net66489), .Z(
        u4_sll_454_ML_int_6__36_) );
  MUX2_X2 u4_sll_454_M1_5_37 ( .A(u4_sll_454_ML_int_5__37_), .B(
        u4_sll_454_ML_int_5__5_), .S(u4_sll_454_net66489), .Z(
        u4_sll_454_ML_int_6__37_) );
  MUX2_X2 u4_sll_454_M1_5_38 ( .A(u4_sll_454_ML_int_5__38_), .B(
        u4_sll_454_ML_int_5__6_), .S(u4_sll_454_net66489), .Z(
        u4_sll_454_ML_int_6__38_) );
  MUX2_X2 u4_sll_454_M1_5_39 ( .A(u4_sll_454_ML_int_5__39_), .B(
        u4_sll_454_ML_int_5__7_), .S(u4_sll_454_net66489), .Z(
        u4_sll_454_ML_int_6__39_) );
  MUX2_X2 u4_sll_454_M1_5_40 ( .A(u4_sll_454_ML_int_5__40_), .B(
        u4_sll_454_ML_int_5__8_), .S(u4_sll_454_net66489), .Z(
        u4_sll_454_ML_int_6__40_) );
  MUX2_X2 u4_sll_454_M1_5_41 ( .A(u4_sll_454_ML_int_5__41_), .B(
        u4_sll_454_ML_int_5__9_), .S(u4_sll_454_net66489), .Z(
        u4_sll_454_ML_int_6__41_) );
  MUX2_X2 u4_sll_454_M1_5_42 ( .A(u4_sll_454_ML_int_5__42_), .B(
        u4_sll_454_ML_int_5__10_), .S(u4_sll_454_net66489), .Z(
        u4_sll_454_ML_int_6__42_) );
  MUX2_X2 u4_sll_454_M1_5_43 ( .A(u4_sll_454_ML_int_5__43_), .B(
        u4_sll_454_ML_int_5__11_), .S(u4_sll_454_net66489), .Z(
        u4_sll_454_ML_int_6__43_) );
  MUX2_X2 u4_sll_454_M1_5_45 ( .A(u4_sll_454_ML_int_5__45_), .B(
        u4_sll_454_ML_int_5__13_), .S(u4_sll_454_net66491), .Z(
        u4_sll_454_ML_int_6__45_) );
  MUX2_X2 u4_sll_454_M1_5_46 ( .A(u4_sll_454_ML_int_5__46_), .B(
        u4_sll_454_ML_int_5__14_), .S(u4_sll_454_net66491), .Z(
        u4_sll_454_ML_int_6__46_) );
  MUX2_X2 u4_sll_454_M1_5_47 ( .A(u4_sll_454_ML_int_5__47_), .B(
        u4_sll_454_ML_int_5__15_), .S(u4_sll_454_net66491), .Z(
        u4_sll_454_ML_int_6__47_) );
  MUX2_X2 u4_sll_454_M1_5_48 ( .A(u4_sll_454_ML_int_5__48_), .B(
        u4_sll_454_ML_int_5__16_), .S(u4_sll_454_net66491), .Z(
        u4_sll_454_ML_int_6__48_) );
  MUX2_X2 u4_sll_454_M1_5_49 ( .A(u4_sll_454_ML_int_5__49_), .B(
        u4_sll_454_ML_int_5__17_), .S(u4_sll_454_net66491), .Z(
        u4_sll_454_ML_int_6__49_) );
  MUX2_X2 u4_sll_454_M1_5_50 ( .A(u4_sll_454_ML_int_5__50_), .B(
        u4_sll_454_ML_int_5__18_), .S(u4_sll_454_net66491), .Z(
        u4_sll_454_ML_int_6__50_) );
  MUX2_X2 u4_sll_454_M1_5_51 ( .A(u4_sll_454_ML_int_5__51_), .B(
        u4_sll_454_ML_int_5__19_), .S(u4_sll_454_net66491), .Z(
        u4_sll_454_ML_int_6__51_) );
  MUX2_X2 u4_sll_454_M1_5_52 ( .A(u4_sll_454_ML_int_5__52_), .B(
        u4_sll_454_ML_int_5__20_), .S(u4_sll_454_net66491), .Z(
        u4_sll_454_ML_int_6__52_) );
  MUX2_X2 u4_sll_454_M1_5_53 ( .A(u4_sll_454_ML_int_5__53_), .B(
        u4_sll_454_ML_int_5__21_), .S(u4_sll_454_net66491), .Z(
        u4_sll_454_ML_int_6__53_) );
  MUX2_X2 u4_sll_454_M1_5_54 ( .A(u4_sll_454_ML_int_5__54_), .B(
        u4_sll_454_ML_int_5__22_), .S(u4_sll_454_net66491), .Z(
        u4_sll_454_ML_int_6__54_) );
  MUX2_X2 u4_sll_454_M1_5_55 ( .A(u4_sll_454_ML_int_5__55_), .B(
        u4_sll_454_ML_int_5__23_), .S(u4_sll_454_net66493), .Z(
        u4_sll_454_ML_int_6__55_) );
  MUX2_X2 u4_sll_454_M1_5_56 ( .A(u4_sll_454_ML_int_5__56_), .B(
        u4_sll_454_ML_int_5__24_), .S(u4_sll_454_net66493), .Z(
        u4_sll_454_ML_int_6__56_) );
  MUX2_X2 u4_sll_454_M1_5_57 ( .A(u4_sll_454_ML_int_5__57_), .B(
        u4_sll_454_ML_int_5__25_), .S(u4_sll_454_net66493), .Z(
        u4_sll_454_ML_int_6__57_) );
  MUX2_X2 u4_sll_454_M1_5_58 ( .A(u4_sll_454_ML_int_5__58_), .B(
        u4_sll_454_ML_int_5__26_), .S(u4_sll_454_net66493), .Z(
        u4_sll_454_ML_int_6__58_) );
  MUX2_X2 u4_sll_454_M1_5_59 ( .A(u4_sll_454_ML_int_5__59_), .B(
        u4_sll_454_ML_int_5__27_), .S(u4_sll_454_net66493), .Z(
        u4_sll_454_ML_int_6__59_) );
  MUX2_X2 u4_sll_454_M1_5_60 ( .A(u4_sll_454_ML_int_5__60_), .B(
        u4_sll_454_ML_int_5__28_), .S(u4_sll_454_net66493), .Z(
        u4_sll_454_ML_int_6__60_) );
  MUX2_X2 u4_sll_454_M1_5_61 ( .A(u4_sll_454_ML_int_5__61_), .B(
        u4_sll_454_ML_int_5__29_), .S(u4_sll_454_net66493), .Z(
        u4_sll_454_ML_int_6__61_) );
  MUX2_X2 u4_sll_454_M1_5_62 ( .A(u4_sll_454_ML_int_5__62_), .B(
        u4_sll_454_ML_int_5__30_), .S(u4_sll_454_net66493), .Z(
        u4_sll_454_ML_int_6__62_) );
  MUX2_X2 u4_sll_454_M1_5_63 ( .A(u4_sll_454_ML_int_5__63_), .B(
        u4_sll_454_ML_int_5__31_), .S(u4_sll_454_net66493), .Z(
        u4_sll_454_ML_int_6__63_) );
  MUX2_X2 u4_sll_454_M1_5_64 ( .A(u4_sll_454_ML_int_5__64_), .B(
        u4_sll_454_ML_int_5__32_), .S(u4_sll_454_net66493), .Z(
        u4_sll_454_ML_int_6__64_) );
  MUX2_X2 u4_sll_454_M1_5_65 ( .A(u4_sll_454_ML_int_5__65_), .B(
        u4_sll_454_ML_int_5__33_), .S(u4_sll_454_net66493), .Z(
        u4_sll_454_ML_int_6__65_) );
  MUX2_X2 u4_sll_454_M1_5_66 ( .A(u4_sll_454_ML_int_5__66_), .B(
        u4_sll_454_ML_int_5__34_), .S(u4_sll_454_net66495), .Z(
        u4_sll_454_ML_int_6__66_) );
  MUX2_X2 u4_sll_454_M1_5_67 ( .A(u4_sll_454_ML_int_5__67_), .B(
        u4_sll_454_ML_int_5__35_), .S(u4_sll_454_net66495), .Z(
        u4_sll_454_ML_int_6__67_) );
  MUX2_X2 u4_sll_454_M1_5_68 ( .A(u4_sll_454_ML_int_5__68_), .B(
        u4_sll_454_ML_int_5__36_), .S(u4_sll_454_net66495), .Z(
        u4_sll_454_ML_int_6__68_) );
  MUX2_X2 u4_sll_454_M1_5_69 ( .A(u4_sll_454_ML_int_5__69_), .B(
        u4_sll_454_ML_int_5__37_), .S(u4_sll_454_net66495), .Z(
        u4_sll_454_ML_int_6__69_) );
  MUX2_X2 u4_sll_454_M1_5_70 ( .A(u4_sll_454_ML_int_5__70_), .B(
        u4_sll_454_ML_int_5__38_), .S(u4_sll_454_net66495), .Z(
        u4_sll_454_ML_int_6__70_) );
  MUX2_X2 u4_sll_454_M1_5_71 ( .A(u4_sll_454_ML_int_5__71_), .B(
        u4_sll_454_ML_int_5__39_), .S(u4_sll_454_net66495), .Z(
        u4_sll_454_ML_int_6__71_) );
  MUX2_X2 u4_sll_454_M1_5_72 ( .A(u4_sll_454_ML_int_5__72_), .B(
        u4_sll_454_ML_int_5__40_), .S(u4_sll_454_net66495), .Z(
        u4_sll_454_ML_int_6__72_) );
  MUX2_X2 u4_sll_454_M1_5_73 ( .A(u4_sll_454_ML_int_5__73_), .B(
        u4_sll_454_ML_int_5__41_), .S(u4_sll_454_net66495), .Z(
        u4_sll_454_ML_int_6__73_) );
  MUX2_X2 u4_sll_454_M1_5_74 ( .A(u4_sll_454_ML_int_5__74_), .B(
        u4_sll_454_ML_int_5__42_), .S(u4_sll_454_net66495), .Z(
        u4_sll_454_ML_int_6__74_) );
  MUX2_X2 u4_sll_454_M1_5_75 ( .A(u4_sll_454_ML_int_5__75_), .B(
        u4_sll_454_ML_int_5__43_), .S(u4_sll_454_net66495), .Z(
        u4_sll_454_ML_int_6__75_) );
  MUX2_X2 u4_sll_454_M1_5_77 ( .A(u4_sll_454_ML_int_5__77_), .B(
        u4_sll_454_ML_int_5__45_), .S(u4_sll_454_net66497), .Z(
        u4_sll_454_ML_int_6__77_) );
  MUX2_X2 u4_sll_454_M1_5_78 ( .A(u4_sll_454_ML_int_5__78_), .B(
        u4_sll_454_ML_int_5__46_), .S(u4_sll_454_net66497), .Z(
        u4_sll_454_ML_int_6__78_) );
  MUX2_X2 u4_sll_454_M1_5_79 ( .A(u4_sll_454_ML_int_5__79_), .B(
        u4_sll_454_ML_int_5__47_), .S(u4_sll_454_net66497), .Z(
        u4_sll_454_ML_int_6__79_) );
  MUX2_X2 u4_sll_454_M1_5_80 ( .A(u4_sll_454_ML_int_5__80_), .B(
        u4_sll_454_ML_int_5__48_), .S(u4_sll_454_net66497), .Z(
        u4_sll_454_ML_int_6__80_) );
  MUX2_X2 u4_sll_454_M1_5_81 ( .A(u4_sll_454_ML_int_5__81_), .B(
        u4_sll_454_ML_int_5__49_), .S(u4_sll_454_net66497), .Z(
        u4_sll_454_ML_int_6__81_) );
  MUX2_X2 u4_sll_454_M1_5_82 ( .A(u4_sll_454_ML_int_5__82_), .B(
        u4_sll_454_ML_int_5__50_), .S(u4_sll_454_net66497), .Z(
        u4_sll_454_ML_int_6__82_) );
  MUX2_X2 u4_sll_454_M1_5_83 ( .A(u4_sll_454_ML_int_5__83_), .B(
        u4_sll_454_ML_int_5__51_), .S(u4_sll_454_net66497), .Z(
        u4_sll_454_ML_int_6__83_) );
  MUX2_X2 u4_sll_454_M1_5_84 ( .A(u4_sll_454_ML_int_5__84_), .B(
        u4_sll_454_ML_int_5__52_), .S(u4_sll_454_net66497), .Z(
        u4_sll_454_ML_int_6__84_) );
  MUX2_X2 u4_sll_454_M1_5_85 ( .A(u4_sll_454_ML_int_5__85_), .B(
        u4_sll_454_ML_int_5__53_), .S(u4_sll_454_net66497), .Z(
        u4_sll_454_ML_int_6__85_) );
  MUX2_X2 u4_sll_454_M1_5_86 ( .A(u4_sll_454_ML_int_5__86_), .B(
        u4_sll_454_ML_int_5__54_), .S(u4_sll_454_net66497), .Z(
        u4_sll_454_ML_int_6__86_) );
  MUX2_X2 u4_sll_454_M1_5_87 ( .A(u4_sll_454_ML_int_5__87_), .B(
        u4_sll_454_ML_int_5__55_), .S(u4_sll_454_net66497), .Z(
        u4_sll_454_ML_int_6__87_) );
  MUX2_X2 u4_sll_454_M1_5_88 ( .A(u4_sll_454_ML_int_5__88_), .B(
        u4_sll_454_ML_int_5__56_), .S(u4_sll_454_net66499), .Z(
        u4_sll_454_ML_int_6__88_) );
  MUX2_X2 u4_sll_454_M1_5_89 ( .A(u4_sll_454_ML_int_5__89_), .B(
        u4_sll_454_ML_int_5__57_), .S(u4_sll_454_net66499), .Z(
        u4_sll_454_ML_int_6__89_) );
  MUX2_X2 u4_sll_454_M1_5_90 ( .A(u4_sll_454_ML_int_5__90_), .B(
        u4_sll_454_ML_int_5__58_), .S(u4_sll_454_net66499), .Z(
        u4_sll_454_ML_int_6__90_) );
  MUX2_X2 u4_sll_454_M1_5_91 ( .A(u4_sll_454_ML_int_5__91_), .B(
        u4_sll_454_ML_int_5__59_), .S(u4_sll_454_net66499), .Z(
        u4_sll_454_ML_int_6__91_) );
  MUX2_X2 u4_sll_454_M1_5_92 ( .A(u4_sll_454_ML_int_5__92_), .B(
        u4_sll_454_ML_int_5__60_), .S(u4_sll_454_net66499), .Z(
        u4_sll_454_ML_int_6__92_) );
  MUX2_X2 u4_sll_454_M1_5_93 ( .A(u4_sll_454_ML_int_5__93_), .B(
        u4_sll_454_ML_int_5__61_), .S(u4_sll_454_net66499), .Z(
        u4_sll_454_ML_int_6__93_) );
  MUX2_X2 u4_sll_454_M1_5_94 ( .A(u4_sll_454_ML_int_5__94_), .B(
        u4_sll_454_ML_int_5__62_), .S(u4_sll_454_net66499), .Z(
        u4_sll_454_ML_int_6__94_) );
  MUX2_X2 u4_sll_454_M1_5_95 ( .A(u4_sll_454_ML_int_5__95_), .B(
        u4_sll_454_ML_int_5__63_), .S(u4_sll_454_net66499), .Z(
        u4_sll_454_ML_int_6__95_) );
  MUX2_X2 u4_sll_454_M1_5_96 ( .A(u4_sll_454_ML_int_5__96_), .B(
        u4_sll_454_ML_int_5__64_), .S(u4_sll_454_net66499), .Z(
        u4_sll_454_ML_int_6__96_) );
  MUX2_X2 u4_sll_454_M1_5_97 ( .A(u4_sll_454_ML_int_5__97_), .B(
        u4_sll_454_ML_int_5__65_), .S(u4_sll_454_net66499), .Z(
        u4_sll_454_ML_int_6__97_) );
  MUX2_X2 u4_sll_454_M1_5_98 ( .A(u4_sll_454_ML_int_5__98_), .B(
        u4_sll_454_ML_int_5__66_), .S(u4_sll_454_net66499), .Z(
        u4_sll_454_ML_int_6__98_) );
  MUX2_X2 u4_sll_454_M1_5_99 ( .A(u4_sll_454_ML_int_5__99_), .B(
        u4_sll_454_ML_int_5__67_), .S(u4_sll_454_net66501), .Z(
        u4_sll_454_ML_int_6__99_) );
  MUX2_X2 u4_sll_454_M1_5_100 ( .A(u4_sll_454_ML_int_5__100_), .B(
        u4_sll_454_ML_int_5__68_), .S(u4_sll_454_net66501), .Z(
        u4_sll_454_ML_int_6__100_) );
  MUX2_X2 u4_sll_454_M1_5_101 ( .A(u4_sll_454_ML_int_5__101_), .B(
        u4_sll_454_ML_int_5__69_), .S(u4_sll_454_net66501), .Z(
        u4_sll_454_ML_int_6__101_) );
  MUX2_X2 u4_sll_454_M1_5_102 ( .A(u4_sll_454_ML_int_5__102_), .B(
        u4_sll_454_ML_int_5__70_), .S(u4_sll_454_net66501), .Z(
        u4_sll_454_ML_int_6__102_) );
  MUX2_X2 u4_sll_454_M1_5_103 ( .A(u4_sll_454_ML_int_5__103_), .B(
        u4_sll_454_ML_int_5__71_), .S(u4_sll_454_net66501), .Z(
        u4_sll_454_ML_int_6__103_) );
  MUX2_X2 u4_sll_454_M1_5_104 ( .A(u4_sll_454_ML_int_5__104_), .B(
        u4_sll_454_ML_int_5__72_), .S(u4_sll_454_net66501), .Z(
        u4_sll_454_ML_int_6__104_) );
  MUX2_X2 u4_sll_454_M1_5_105 ( .A(u4_sll_454_ML_int_5__105_), .B(
        u4_sll_454_ML_int_5__73_), .S(u4_sll_454_net66501), .Z(
        u4_sll_454_ML_int_6__105_) );
  MUX2_X2 u4_sll_454_M1_6_64 ( .A(u4_sll_454_ML_int_6__64_), .B(
        u4_sll_454_ML_int_6__0_), .S(u4_sll_454_net66441), .Z(
        u4_sll_454_ML_int_7__64_) );
  MUX2_X2 u4_sll_454_M1_6_65 ( .A(u4_sll_454_ML_int_6__65_), .B(
        u4_sll_454_ML_int_6__1_), .S(u4_sll_454_net66441), .Z(
        u4_sll_454_ML_int_7__65_) );
  MUX2_X2 u4_sll_454_M1_6_66 ( .A(u4_sll_454_ML_int_6__66_), .B(
        u4_sll_454_ML_int_6__2_), .S(u4_sll_454_net66439), .Z(
        u4_sll_454_ML_int_7__66_) );
  MUX2_X2 u4_sll_454_M1_6_67 ( .A(u4_sll_454_ML_int_6__67_), .B(
        u4_sll_454_ML_int_6__3_), .S(u4_sll_454_net66439), .Z(
        u4_sll_454_ML_int_7__67_) );
  MUX2_X2 u4_sll_454_M1_6_68 ( .A(u4_sll_454_ML_int_6__68_), .B(
        u4_sll_454_ML_int_6__4_), .S(u4_sll_454_net66439), .Z(
        u4_sll_454_ML_int_7__68_) );
  MUX2_X2 u4_sll_454_M1_6_69 ( .A(u4_sll_454_ML_int_6__69_), .B(
        u4_sll_454_ML_int_6__5_), .S(u4_sll_454_net66439), .Z(
        u4_sll_454_ML_int_7__69_) );
  MUX2_X2 u4_sll_454_M1_6_70 ( .A(u4_sll_454_ML_int_6__70_), .B(
        u4_sll_454_ML_int_6__6_), .S(u4_sll_454_net66439), .Z(
        u4_sll_454_ML_int_7__70_) );
  MUX2_X2 u4_sll_454_M1_6_71 ( .A(u4_sll_454_ML_int_6__71_), .B(
        u4_sll_454_ML_int_6__7_), .S(u4_sll_454_net66439), .Z(
        u4_sll_454_ML_int_7__71_) );
  MUX2_X2 u4_sll_454_M1_6_72 ( .A(u4_sll_454_ML_int_6__72_), .B(
        u4_sll_454_ML_int_6__8_), .S(u4_sll_454_net66439), .Z(
        u4_sll_454_ML_int_7__72_) );
  MUX2_X2 u4_sll_454_M1_6_73 ( .A(u4_sll_454_ML_int_6__73_), .B(
        u4_sll_454_ML_int_6__9_), .S(u4_sll_454_net66439), .Z(
        u4_sll_454_ML_int_7__73_) );
  MUX2_X2 u4_sll_454_M1_6_74 ( .A(u4_sll_454_ML_int_6__74_), .B(
        u4_sll_454_ML_int_6__10_), .S(u4_sll_454_net66439), .Z(
        u4_sll_454_ML_int_7__74_) );
  MUX2_X2 u4_sll_454_M1_6_75 ( .A(u4_sll_454_ML_int_6__75_), .B(
        u4_sll_454_ML_int_6__11_), .S(u4_sll_454_net66439), .Z(
        u4_sll_454_ML_int_7__75_) );
  MUX2_X2 u4_sll_454_M1_6_76 ( .A(u4_sll_454_ML_int_6__76_), .B(
        u4_sll_454_ML_int_6__12_), .S(u4_sll_454_net66439), .Z(
        u4_sll_454_ML_int_7__76_) );
  MUX2_X2 u4_sll_454_M1_6_77 ( .A(u4_sll_454_ML_int_6__77_), .B(
        u4_sll_454_ML_int_6__13_), .S(u4_sll_454_net66441), .Z(
        u4_sll_454_ML_int_7__77_) );
  MUX2_X2 u4_sll_454_M1_6_78 ( .A(u4_sll_454_ML_int_6__78_), .B(
        u4_sll_454_ML_int_6__14_), .S(u4_sll_454_net66441), .Z(
        u4_sll_454_ML_int_7__78_) );
  MUX2_X2 u4_sll_454_M1_6_79 ( .A(u4_sll_454_ML_int_6__79_), .B(
        u4_sll_454_ML_int_6__15_), .S(u4_sll_454_net66441), .Z(
        u4_sll_454_ML_int_7__79_) );
  MUX2_X2 u4_sll_454_M1_6_80 ( .A(u4_sll_454_ML_int_6__80_), .B(
        u4_sll_454_ML_int_6__16_), .S(u4_sll_454_net66441), .Z(
        u4_sll_454_ML_int_7__80_) );
  MUX2_X2 u4_sll_454_M1_6_81 ( .A(u4_sll_454_ML_int_6__81_), .B(
        u4_sll_454_ML_int_6__17_), .S(u4_sll_454_net66441), .Z(
        u4_sll_454_ML_int_7__81_) );
  MUX2_X2 u4_sll_454_M1_6_82 ( .A(u4_sll_454_ML_int_6__82_), .B(
        u4_sll_454_ML_int_6__18_), .S(u4_sll_454_net66441), .Z(
        u4_sll_454_ML_int_7__82_) );
  MUX2_X2 u4_sll_454_M1_6_83 ( .A(u4_sll_454_ML_int_6__83_), .B(
        u4_sll_454_ML_int_6__19_), .S(u4_sll_454_net66441), .Z(
        u4_sll_454_ML_int_7__83_) );
  MUX2_X2 u4_sll_454_M1_6_84 ( .A(u4_sll_454_ML_int_6__84_), .B(
        u4_sll_454_ML_int_6__20_), .S(u4_sll_454_net66441), .Z(
        u4_sll_454_ML_int_7__84_) );
  MUX2_X2 u4_sll_454_M1_6_85 ( .A(u4_sll_454_ML_int_6__85_), .B(
        u4_sll_454_ML_int_6__21_), .S(u4_sll_454_net66441), .Z(
        u4_sll_454_ML_int_7__85_) );
  MUX2_X2 u4_sll_454_M1_6_86 ( .A(u4_sll_454_ML_int_6__86_), .B(
        u4_sll_454_ML_int_6__22_), .S(u4_sll_454_net66441), .Z(
        u4_sll_454_ML_int_7__86_) );
  MUX2_X2 u4_sll_454_M1_6_87 ( .A(u4_sll_454_ML_int_6__87_), .B(
        u4_sll_454_ML_int_6__23_), .S(u4_sll_454_net66441), .Z(
        u4_sll_454_ML_int_7__87_) );
  MUX2_X2 u4_sll_454_M1_6_88 ( .A(u4_sll_454_ML_int_6__88_), .B(
        u4_sll_454_ML_int_6__24_), .S(u4_sll_454_net66443), .Z(
        u4_sll_454_ML_int_7__88_) );
  MUX2_X2 u4_sll_454_M1_6_89 ( .A(u4_sll_454_ML_int_6__89_), .B(
        u4_sll_454_ML_int_6__25_), .S(u4_sll_454_net66443), .Z(
        u4_sll_454_ML_int_7__89_) );
  MUX2_X2 u4_sll_454_M1_6_90 ( .A(u4_sll_454_ML_int_6__90_), .B(
        u4_sll_454_ML_int_6__26_), .S(u4_sll_454_net66443), .Z(
        u4_sll_454_ML_int_7__90_) );
  MUX2_X2 u4_sll_454_M1_6_91 ( .A(u4_sll_454_ML_int_6__91_), .B(
        u4_sll_454_ML_int_6__27_), .S(u4_sll_454_net66443), .Z(
        u4_sll_454_ML_int_7__91_) );
  MUX2_X2 u4_sll_454_M1_6_92 ( .A(u4_sll_454_ML_int_6__92_), .B(
        u4_sll_454_ML_int_6__28_), .S(u4_sll_454_net66443), .Z(
        u4_sll_454_ML_int_7__92_) );
  MUX2_X2 u4_sll_454_M1_6_93 ( .A(u4_sll_454_ML_int_6__93_), .B(
        u4_sll_454_ML_int_6__29_), .S(u4_sll_454_net66443), .Z(
        u4_sll_454_ML_int_7__93_) );
  MUX2_X2 u4_sll_454_M1_6_94 ( .A(u4_sll_454_ML_int_6__94_), .B(
        u4_sll_454_ML_int_6__30_), .S(u4_sll_454_net66443), .Z(
        u4_sll_454_ML_int_7__94_) );
  MUX2_X2 u4_sll_454_M1_6_95 ( .A(u4_sll_454_ML_int_6__95_), .B(
        u4_sll_454_ML_int_6__31_), .S(u4_sll_454_net66443), .Z(
        u4_sll_454_ML_int_7__95_) );
  MUX2_X2 u4_sll_454_M1_6_96 ( .A(u4_sll_454_ML_int_6__96_), .B(
        u4_sll_454_ML_int_6__32_), .S(u4_sll_454_net66443), .Z(
        u4_sll_454_ML_int_7__96_) );
  MUX2_X2 u4_sll_454_M1_6_97 ( .A(u4_sll_454_ML_int_6__97_), .B(
        u4_sll_454_ML_int_6__33_), .S(u4_sll_454_net66443), .Z(
        u4_sll_454_ML_int_7__97_) );
  MUX2_X2 u4_sll_454_M1_6_98 ( .A(u4_sll_454_ML_int_6__98_), .B(
        u4_sll_454_ML_int_6__34_), .S(u4_sll_454_net66443), .Z(
        u4_sll_454_ML_int_7__98_) );
  MUX2_X2 u4_sll_454_M1_6_99 ( .A(u4_sll_454_ML_int_6__99_), .B(
        u4_sll_454_ML_int_6__35_), .S(u4_sll_454_net66445), .Z(
        u4_sll_454_ML_int_7__99_) );
  MUX2_X2 u4_sll_454_M1_6_100 ( .A(u4_sll_454_ML_int_6__100_), .B(
        u4_sll_454_ML_int_6__36_), .S(u4_sll_454_net66445), .Z(
        u4_sll_454_ML_int_7__100_) );
  MUX2_X2 u4_sll_454_M1_6_101 ( .A(u4_sll_454_ML_int_6__101_), .B(
        u4_sll_454_ML_int_6__37_), .S(u4_sll_454_net66445), .Z(
        u4_sll_454_ML_int_7__101_) );
  MUX2_X2 u4_sll_454_M1_6_102 ( .A(u4_sll_454_ML_int_6__102_), .B(
        u4_sll_454_ML_int_6__38_), .S(u4_sll_454_net66445), .Z(
        u4_sll_454_ML_int_7__102_) );
  MUX2_X2 u4_sll_454_M1_6_103 ( .A(u4_sll_454_ML_int_6__103_), .B(
        u4_sll_454_ML_int_6__39_), .S(u4_sll_454_net66445), .Z(
        u4_sll_454_ML_int_7__103_) );
  MUX2_X2 u4_sll_454_M1_6_104 ( .A(u4_sll_454_ML_int_6__104_), .B(
        u4_sll_454_ML_int_6__40_), .S(u4_sll_454_net66445), .Z(
        u4_sll_454_ML_int_7__104_) );
  MUX2_X2 u4_sll_454_M1_6_105 ( .A(u4_sll_454_ML_int_6__105_), .B(
        u4_sll_454_ML_int_6__41_), .S(u4_sll_454_net66445), .Z(
        u4_sll_454_ML_int_7__105_) );
endmodule

