
module fpu ( clk, rmode, fpu_op, opa, opb, out, inf, snan, qnan, ine, overflow, 
        underflow, zero, div_by_zero );
  input [1:0] rmode;
  input [2:0] fpu_op;
  input [63:0] opa;
  input [63:0] opb;
  output [63:0] out;
  input clk;
  output inf, snan, qnan, ine, overflow, underflow, zero, div_by_zero;
  wire   inf_d, qnan_d, snan_d, opa_nan, opb_nan, opa_00, opb_00, opa_inf,
         opb_inf, opb_dn, sign_fasu, nan_sign_d, result_zero_sign_d, fasu_op,
         sign_fasu_r, sign_mul, sign_exe, inf_mul, sign_mul_r, sign_exe_r,
         inf_mul_r, exp_ovf_r_1_, N261, N262, N263, N264, N265, N266, N267,
         N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278,
         N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289,
         N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300,
         N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311,
         N312, N313, N342, N347, N348, N349, N350, N351, N352, N353, N354,
         N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365,
         N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376,
         N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387,
         N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398,
         N399, N400, N505, N506, N507, N508, N509, N510, N511, N512, N513,
         N514, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524,
         N525, N526, N527, N528, N529, N530, N531, N532, N533, N534, N535,
         N536, N537, N538, N539, N540, N541, N542, N543, N544, N545, N546,
         N547, N548, N549, N550, N551, N552, N553, N554, N555, N556, N557,
         N558, N559, N560, N561, N608, N609, N610, N611, N612, N613, N614,
         N615, N616, N617, N618, N619, N620, N621, N622, N623, N624, N625,
         N626, N627, N628, N629, N630, N631, N632, N633, N634, N635, N636,
         N637, N638, N639, N640, N641, N642, N643, N644, N645, N646, N647,
         N648, N649, N650, N651, N652, N653, N654, N655, N656, N657, N658,
         N659, N660, N661, N662, N663, N664, N665, N666, N667, N686, N689,
         N692, N694, N697, N698, N699, N700, N704, N705, N709, N710, N711,
         N712, N715, N716, N717, N721, N722, N723, N724, N727, N728, N729,
         N730, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743,
         N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754,
         N755, N756, N757, N758, N759, N760, N761, N762, N763, N764, N765,
         N766, N767, N768, N769, N770, N771, N772, N773, N774, N775, N776,
         N777, N778, N779, N780, N781, N782, N783, N784, N785, N786, N787,
         N788, N789, N790, N791, opas_r1, opas_r2, sign, N794, fasu_op_r1,
         fasu_op_r2, inf_mul2, N798, N799, N800, N801, N802, N803, N804, N805,
         N806, N807, N808, N809, N810, N811, N812, N813, N814, N815, N816,
         N817, N818, N819, N820, N821, N822, N823, N824, N825, N826, N827,
         N828, N829, N830, N831, N832, N833, N834, N835, N836, N837, N838,
         N839, N840, N841, N842, N843, N844, N845, N846, N847, N848, N849,
         N850, N851, N852, N853, N854, N855, N856, N857, N858, N859, N860,
         N880, N894, N904, N907, N909, N911, N916, N917, opa_nan_r, N918, N928,
         u0_N17, u0_N16, u0_fractb_00, u0_fracta_00, u0_expb_00, u0_expa_00,
         u0_N11, u0_N10, u0_N7, u0_N6, u0_snan_r_b, u0_N5, u0_qnan_r_b,
         u0_snan_r_a, u0_N4, u0_qnan_r_a, u0_infb_f_r, u0_infa_f_r, u0_expb_ff,
         u0_expa_ff, u1_N334, u1_fracta_eq_fractb, u1_N325,
         u1_fracta_lt_fractb, u1_N324, u1_add_r, u1_signa_r, u1_sign_d,
         u1_fractb_lt_fracta, u1_N296, u1_N295, u1_sticky,
         u1_adj_op_out_sft_0_, u1_adj_op_out_sft_1_, u1_adj_op_out_sft_2_,
         u1_adj_op_out_sft_3_, u1_adj_op_out_sft_4_, u1_adj_op_out_sft_5_,
         u1_adj_op_out_sft_6_, u1_adj_op_out_sft_7_, u1_adj_op_out_sft_8_,
         u1_adj_op_out_sft_9_, u1_adj_op_out_sft_10_, u1_adj_op_out_sft_11_,
         u1_adj_op_out_sft_12_, u1_adj_op_out_sft_13_, u1_adj_op_out_sft_14_,
         u1_adj_op_out_sft_15_, u1_adj_op_out_sft_16_, u1_adj_op_out_sft_17_,
         u1_adj_op_out_sft_18_, u1_adj_op_out_sft_19_, u1_adj_op_out_sft_20_,
         u1_adj_op_out_sft_21_, u1_adj_op_out_sft_22_, u1_adj_op_out_sft_23_,
         u1_adj_op_out_sft_24_, u1_adj_op_out_sft_25_, u1_adj_op_out_sft_26_,
         u1_adj_op_out_sft_27_, u1_adj_op_out_sft_28_, u1_adj_op_out_sft_29_,
         u1_adj_op_out_sft_30_, u1_adj_op_out_sft_31_, u1_adj_op_out_sft_32_,
         u1_adj_op_out_sft_33_, u1_adj_op_out_sft_34_, u1_adj_op_out_sft_35_,
         u1_adj_op_out_sft_36_, u1_adj_op_out_sft_37_, u1_adj_op_out_sft_38_,
         u1_adj_op_out_sft_39_, u1_adj_op_out_sft_40_, u1_adj_op_out_sft_41_,
         u1_adj_op_out_sft_42_, u1_adj_op_out_sft_43_, u1_adj_op_out_sft_44_,
         u1_adj_op_out_sft_45_, u1_adj_op_out_sft_46_, u1_adj_op_out_sft_47_,
         u1_adj_op_out_sft_48_, u1_adj_op_out_sft_49_, u1_adj_op_out_sft_50_,
         u1_adj_op_out_sft_51_, u1_adj_op_out_sft_52_, u1_adj_op_out_sft_53_,
         u1_adj_op_out_sft_54_, u1_adj_op_out_sft_55_, u1_exp_diff_sft_0_,
         u1_exp_lt_27, u1_adj_op_29_, u1_adj_op_36_, u1_N88, u1_N87, u1_N86,
         u1_N85, u1_N84, u1_N83, u1_N82, u1_N81, u1_N80, u1_N79, u1_N78,
         u1_N75, u1_exp_diff_0_, u1_exp_diff_1_, u1_exp_diff_2_,
         u1_exp_diff_3_, u1_exp_diff_4_, u1_exp_diff_5_, u1_exp_diff_6_,
         u1_exp_diff_7_, u1_exp_diff_8_, u1_exp_diff_9_, u1_exp_diff_10_,
         u1_expa_lt_expb, u2_N157, u2_N121, u2_sign_d, u2_N114, u2_N113,
         u2_N111, u2_exp_ovf_d_0_, u2_exp_ovf_d_1_, u2_N86, u2_N85, u2_N84,
         u2_N83, u2_N82, u2_N81, u2_N80, u2_N79, u2_N78, u2_N77, u2_N76,
         u2_N75, u2_N74, u2_N73, u2_N72, u2_N71, u2_N70, u2_N69, u2_N68,
         u2_N67, u2_N66, u2_N64, u2_N63, u2_N62, u2_N61, u2_N60, u2_N59,
         u2_N58, u2_N57, u2_N56, u2_N55, u2_N54, u2_exp_tmp4_1_,
         u2_exp_tmp4_2_, u2_exp_tmp4_3_, u2_exp_tmp4_4_, u2_exp_tmp4_10_,
         u2_exp_tmp3_0_, u2_exp_tmp3_1_, u2_exp_tmp3_2_, u2_exp_tmp3_3_,
         u2_exp_tmp3_4_, u2_exp_tmp3_5_, u2_exp_tmp3_6_, u2_exp_tmp3_7_,
         u2_exp_tmp3_8_, u2_exp_tmp3_9_, u2_exp_tmp3_10_, u2_N53, u2_N52,
         u2_N51, u2_N50, u2_N49, u2_N48, u2_N47, u2_N46, u2_N45, u2_N44,
         u2_N43, u2_N41, u2_N40, u2_N39, u2_N38, u2_N37, u2_N36, u2_N35,
         u2_N34, u2_N33, u2_N32, u2_N31, u2_exp_tmp1_1_, u2_exp_tmp1_2_,
         u2_exp_tmp1_3_, u2_N29, u2_N28, u2_N27, u2_N26, u2_N25, u2_N24,
         u2_N23, u2_N22, u2_N21, u2_N20, u2_N19, u2_N18, u2_N17, u2_N16,
         u2_N15, u2_N14, u2_N13, u2_N12, u2_N11, u2_N10, u2_N9, u2_N8, u2_N7,
         u2_N6, u3_N116, u3_N115, u3_N114, u3_N113, u3_N112, u3_N111, u3_N110,
         u3_N109, u3_N108, u3_N107, u3_N106, u3_N105, u3_N104, u3_N103,
         u3_N102, u3_N101, u3_N100, u3_N99, u3_N98, u3_N97, u3_N96, u3_N95,
         u3_N94, u3_N93, u3_N92, u3_N91, u3_N90, u3_N89, u3_N88, u3_N87,
         u3_N86, u3_N85, u3_N84, u3_N83, u3_N82, u3_N81, u3_N80, u3_N79,
         u3_N78, u3_N77, u3_N76, u3_N75, u3_N74, u3_N73, u3_N72, u3_N71,
         u3_N70, u3_N69, u3_N68, u3_N67, u3_N66, u3_N65, u3_N64, u3_N63,
         u3_N62, u3_N61, u3_N60, u3_N59, u3_N58, u3_N57, u3_N56, u3_N55,
         u3_N54, u3_N53, u3_N52, u3_N51, u3_N50, u3_N49, u3_N48, u3_N47,
         u3_N46, u3_N45, u3_N44, u3_N43, u3_N42, u3_N41, u3_N40, u3_N39,
         u3_N38, u3_N37, u3_N36, u3_N35, u3_N34, u3_N33, u3_N32, u3_N31,
         u3_N30, u3_N29, u3_N28, u3_N27, u3_N26, u3_N25, u3_N24, u3_N23,
         u3_N22, u3_N21, u3_N20, u3_N19, u3_N18, u3_N17, u3_N16, u3_N15,
         u3_N14, u3_N13, u3_N12, u3_N11, u3_N10, u3_N9, u3_N8, u3_N7, u3_N6,
         u3_N5, u3_N4, u3_N3, u5_N105, u5_N104, u5_N103, u5_N102, u5_N101,
         u5_N100, u5_N99, u5_N98, u5_N97, u5_N96, u5_N95, u5_N94, u5_N93,
         u5_N92, u5_N91, u5_N90, u5_N89, u5_N88, u5_N87, u5_N86, u5_N85,
         u5_N84, u5_N83, u5_N82, u5_N81, u5_N80, u5_N79, u5_N78, u5_N77,
         u5_N76, u5_N75, u5_N74, u5_N73, u5_N72, u5_N71, u5_N70, u5_N69,
         u5_N68, u5_N67, u5_N66, u5_N65, u5_N64, u5_N63, u5_N62, u5_N61,
         u5_N60, u5_N59, u5_N58, u5_N57, u5_N56, u5_N55, u5_N54, u5_N53,
         u5_N52, u5_N51, u5_N50, u5_N49, u5_N48, u5_N47, u5_N46, u5_N45,
         u5_N44, u5_N43, u5_N42, u5_N41, u5_N40, u5_N39, u5_N38, u5_N37,
         u5_N36, u5_N35, u5_N34, u5_N33, u5_N32, u5_N31, u5_N30, u5_N29,
         u5_N28, u5_N27, u5_N26, u5_N25, u5_N24, u5_N23, u5_N22, u5_N21,
         u5_N20, u5_N19, u5_N18, u5_N17, u5_N16, u5_N15, u5_N14, u5_N13,
         u5_N12, u5_N11, u5_N10, u5_N9, u5_N8, u5_N7, u5_N6, u5_N5, u5_N4,
         u5_N3, u5_N2, u5_N1, u5_N0, u6_N107, u6_N106, u6_N105, u6_N104,
         u6_N103, u6_N102, u6_N101, u6_N100, u6_N99, u6_N98, u6_N97, u6_N96,
         u6_N95, u6_N94, u6_N93, u6_N92, u6_N91, u6_N90, u6_N89, u6_N88,
         u6_N87, u6_N86, u6_N85, u6_N84, u6_N83, u6_N82, u6_N81, u6_N80,
         u6_N79, u6_N78, u6_N77, u6_N76, u6_N75, u6_N74, u6_N73, u6_N72,
         u6_N71, u6_N70, u6_N69, u6_N68, u6_N67, u6_N66, u6_N65, u6_N64,
         u6_N63, u6_N62, u6_N61, u6_N60, u6_N59, u6_N58, u6_N57, u6_N56,
         u6_N55, u6_N52, u6_N51, u6_N50, u6_N49, u6_N48, u6_N47, u6_N46,
         u6_N45, u6_N44, u6_N43, u6_N42, u6_N41, u6_N40, u6_N39, u6_N38,
         u6_N37, u6_N36, u6_N35, u6_N34, u6_N33, u6_N32, u6_N31, u6_N30,
         u6_N29, u6_N28, u6_N27, u6_N26, u6_N25, u6_N24, u6_N23, u6_N22,
         u6_N21, u6_N20, u6_N19, u6_N18, u6_N17, u6_N16, u6_N15, u6_N14,
         u6_N13, u6_N12, u6_N11, u6_N10, u6_N9, u6_N8, u6_N7, u6_N6, u6_N5,
         u6_N4, u6_N3, u6_N2, u6_N1, u6_N0, u4_N6893, u4_N6892, u4_N6891,
         u4_N6440, u4_N6439, u4_N6438, u4_N6437, u4_N6436, u4_N6435, u4_N6434,
         u4_N6433, u4_N6432, u4_N6431, u4_N6275, u4_N6273, u4_N6272, u4_N6269,
         u4_N6268, u4_N6267, u4_N6240, u4_N6238, u4_N6188, u4_N6179, u4_N6159,
         u4_N6158, u4_div_exp2_0_, u4_div_exp2_1_, u4_div_exp2_2_,
         u4_div_exp2_3_, u4_div_exp2_4_, u4_div_exp2_5_, u4_div_exp2_6_,
         u4_div_exp2_7_, u4_div_exp2_8_, u4_div_exp2_9_, u4_div_exp2_10_,
         u4_div_exp1_0_, u4_div_exp1_1_, u4_div_exp1_2_, u4_div_exp1_3_,
         u4_div_exp1_4_, u4_div_exp1_5_, u4_div_exp1_6_, u4_div_exp1_7_,
         u4_div_exp1_8_, u4_div_exp1_9_, u4_div_exp1_10_, u4_fi_ldz_2a_0_,
         u4_fi_ldz_2a_1_, u4_fi_ldz_2a_2_, u4_fi_ldz_2a_3_, u4_fi_ldz_2a_4_,
         u4_fi_ldz_2a_5_, u4_fi_ldz_2a_6_, u4_ldz_all_0_, u4_ldz_all_1_,
         u4_ldz_all_2_, u4_ldz_all_3_, u4_ldz_all_4_, u4_ldz_all_5_,
         u4_ldz_all_6_, u4_N6137, u4_N6136, u4_N6135, u4_N6134, u4_N6133,
         u4_N6132, u4_N6131, u4_exp_out1_1_, u4_exp_out_pl1_0_,
         u4_exp_out_pl1_1_, u4_exp_out_pl1_2_, u4_exp_out_pl1_3_,
         u4_exp_out_pl1_4_, u4_exp_out_pl1_5_, u4_exp_out_pl1_6_,
         u4_exp_out_pl1_7_, u4_exp_out_pl1_8_, u4_exp_out_pl1_9_,
         u4_exp_out_pl1_10_, u4_fi_ldz_mi1_0_, u4_fi_ldz_mi1_1_,
         u4_fi_ldz_mi1_2_, u4_fi_ldz_mi1_3_, u4_fi_ldz_mi1_4_,
         u4_fi_ldz_mi1_5_, u4_fi_ldz_mi1_6_, u4_N6113, u4_N6112, u4_N6111,
         u4_N6110, u4_N6109, u4_N6108, u4_N6107, u4_N6106, u4_N6105, u4_N6104,
         u4_N6103, u4_N6102, u4_N6101, u4_N6100, u4_N6099, u4_N6098, u4_N6097,
         u4_N6096, u4_N6095, u4_N6094, u4_N6093, u4_N6092, u4_N6091, u4_N6090,
         u4_N6089, u4_N6088, u4_N6087, u4_N6086, u4_N6085, u4_N6084, u4_N6083,
         u4_N6082, u4_N6081, u4_N6080, u4_N6079, u4_N6078, u4_N6077, u4_N6076,
         u4_N6075, u4_N6074, u4_N6073, u4_N6072, u4_N6071, u4_N6070, u4_N6069,
         u4_N6068, u4_N6067, u4_N6066, u4_N6065, u4_N6064, u4_N6063, u4_N6062,
         u4_N6061, u4_N6060, u4_N6059, u4_N6058, u4_N6057, u4_N6056, u4_N6055,
         u4_N6054, u4_N6053, u4_N6052, u4_N6051, u4_N6050, u4_N6049, u4_N6048,
         u4_N6047, u4_N6046, u4_N6045, u4_N6044, u4_N6043, u4_N6042, u4_N6041,
         u4_N6040, u4_N6039, u4_N6038, u4_N6037, u4_N6036, u4_N6035, u4_N6034,
         u4_N6033, u4_N6032, u4_N6031, u4_N6030, u4_N6029, u4_N6028, u4_N6027,
         u4_N6026, u4_N6025, u4_N6024, u4_N6023, u4_N6022, u4_N6021, u4_N6020,
         u4_N6019, u4_N6018, u4_N6017, u4_N6016, u4_N6015, u4_N6014, u4_N6013,
         u4_N6012, u4_N6011, u4_N6010, u4_N6009, u4_N6008, u4_N6005, u4_N6004,
         u4_N6003, u4_N6002, u4_N6001, u4_N6000, u4_N5999, u4_N5998, u4_N5997,
         u4_N5996, u4_N5995, u4_N5994, u4_N5993, u4_N5992, u4_N5991, u4_N5990,
         u4_N5989, u4_N5988, u4_N5987, u4_N5986, u4_N5985, u4_N5984, u4_N5983,
         u4_N5982, u4_N5981, u4_N5980, u4_N5979, u4_N5978, u4_N5977, u4_N5976,
         u4_N5975, u4_N5974, u4_N5973, u4_N5972, u4_N5971, u4_N5970, u4_N5969,
         u4_N5968, u4_N5967, u4_N5966, u4_N5965, u4_N5964, u4_N5963, u4_N5962,
         u4_N5961, u4_N5960, u4_N5959, u4_N5958, u4_N5957, u4_N5956, u4_N5955,
         u4_N5954, u4_N5953, u4_N5952, u4_N5951, u4_N5950, u4_N5949, u4_N5948,
         u4_N5947, u4_N5946, u4_N5945, u4_N5944, u4_N5943, u4_N5942, u4_N5941,
         u4_N5940, u4_N5939, u4_N5938, u4_N5937, u4_N5936, u4_N5935, u4_N5934,
         u4_N5933, u4_N5932, u4_N5931, u4_N5930, u4_N5929, u4_N5928, u4_N5927,
         u4_N5926, u4_N5925, u4_N5924, u4_N5923, u4_N5922, u4_N5921, u4_N5920,
         u4_N5919, u4_N5918, u4_N5917, u4_N5916, u4_N5915, u4_N5914, u4_N5913,
         u4_N5912, u4_N5911, u4_N5910, u4_N5909, u4_N5908, u4_N5907, u4_N5906,
         u4_N5905, u4_N5904, u4_N5903, u4_N5902, u4_N5901, u4_N5900, u4_N5898,
         u4_exp_in_pl1_0_, u4_exp_in_pl1_1_, u4_exp_in_pl1_2_,
         u4_exp_in_pl1_3_, u4_exp_in_pl1_4_, u4_exp_in_pl1_5_,
         u4_exp_in_pl1_6_, u4_exp_in_pl1_7_, u4_exp_in_pl1_8_,
         u4_exp_in_pl1_9_, u4_exp_in_pl1_10_, u4_exp_in_pl1_11_,
         u4_f2i_shft_1_, u4_f2i_shft_2_, u4_f2i_shft_3_, u4_f2i_shft_4_,
         u4_f2i_shft_5_, u4_f2i_shft_6_, u4_f2i_shft_7_, u4_f2i_shft_8_,
         u4_f2i_shft_9_, u4_f2i_shft_10_, u4_N5837, u4_div_shft3_0_,
         u4_div_shft3_1_, u4_div_shft3_2_, u4_div_shft3_3_, u4_div_shft3_4_,
         u4_div_shft3_5_, u4_div_shft3_6_, u4_div_shft3_7_, u4_div_shft3_8_,
         u4_div_shft3_9_, u4_div_shft3_10_, u4_exp_in_mi1_1_, u4_exp_in_mi1_2_,
         u4_exp_in_mi1_3_, u4_exp_in_mi1_4_, u4_exp_in_mi1_5_,
         u4_exp_in_mi1_6_, u4_exp_in_mi1_7_, u4_exp_in_mi1_8_,
         u4_exp_in_mi1_9_, u4_exp_in_mi1_10_, u4_exp_in_mi1_11_, u4_N5831,
         u4_N5830, u4_fract_out_pl1_0_, u4_fract_out_pl1_1_,
         u4_fract_out_pl1_2_, u4_fract_out_pl1_3_, u4_fract_out_pl1_4_,
         u4_fract_out_pl1_5_, u4_fract_out_pl1_6_, u4_fract_out_pl1_7_,
         u4_fract_out_pl1_8_, u4_fract_out_pl1_9_, u4_fract_out_pl1_10_,
         u4_fract_out_pl1_11_, u4_fract_out_pl1_12_, u4_fract_out_pl1_13_,
         u4_fract_out_pl1_14_, u4_fract_out_pl1_15_, u4_fract_out_pl1_16_,
         u4_fract_out_pl1_17_, u4_fract_out_pl1_18_, u4_fract_out_pl1_19_,
         u4_fract_out_pl1_20_, u4_fract_out_pl1_21_, u4_fract_out_pl1_22_,
         u4_fract_out_pl1_23_, u4_fract_out_pl1_24_, u4_fract_out_pl1_25_,
         u4_fract_out_pl1_26_, u4_fract_out_pl1_27_, u4_fract_out_pl1_28_,
         u4_fract_out_pl1_29_, u4_fract_out_pl1_30_, u4_fract_out_pl1_31_,
         u4_fract_out_pl1_32_, u4_fract_out_pl1_33_, u4_fract_out_pl1_34_,
         u4_fract_out_pl1_35_, u4_fract_out_pl1_36_, u4_fract_out_pl1_37_,
         u4_fract_out_pl1_38_, u4_fract_out_pl1_39_, u4_fract_out_pl1_40_,
         u4_fract_out_pl1_41_, u4_fract_out_pl1_42_, u4_fract_out_pl1_43_,
         u4_fract_out_pl1_44_, u4_fract_out_pl1_45_, u4_fract_out_pl1_46_,
         u4_fract_out_pl1_47_, u4_fract_out_pl1_48_, u4_fract_out_pl1_49_,
         u4_fract_out_pl1_50_, u4_fract_out_pl1_51_, u4_fract_out_pl1_52_,
         u4_exp_next_mi_0_, u4_exp_next_mi_1_, u4_exp_next_mi_2_,
         u4_exp_next_mi_3_, u4_exp_next_mi_4_, u4_exp_next_mi_5_,
         u4_exp_next_mi_6_, u4_exp_next_mi_7_, u4_exp_next_mi_8_,
         u4_exp_next_mi_9_, u4_exp_next_mi_10_, u4_exp_next_mi_11_,
         u4_fract_out_0_, u4_fract_out_1_, u4_fract_out_2_, u4_fract_out_3_,
         u4_fract_out_4_, u4_fract_out_5_, u4_fract_out_6_, u4_fract_out_7_,
         u4_fract_out_8_, u4_fract_out_9_, u4_fract_out_10_, u4_fract_out_11_,
         u4_fract_out_12_, u4_fract_out_13_, u4_fract_out_14_,
         u4_fract_out_15_, u4_fract_out_16_, u4_fract_out_17_,
         u4_fract_out_18_, u4_fract_out_19_, u4_fract_out_20_,
         u4_fract_out_21_, u4_fract_out_22_, u4_fract_out_23_,
         u4_fract_out_24_, u4_fract_out_25_, u4_fract_out_26_,
         u4_fract_out_27_, u4_fract_out_28_, u4_fract_out_29_,
         u4_fract_out_30_, u4_fract_out_31_, u4_fract_out_32_,
         u4_fract_out_33_, u4_fract_out_34_, u4_fract_out_35_,
         u4_fract_out_36_, u4_fract_out_37_, u4_fract_out_38_,
         u4_fract_out_39_, u4_fract_out_40_, u4_fract_out_41_,
         u4_fract_out_42_, u4_fract_out_43_, u4_fract_out_44_,
         u4_fract_out_45_, u4_fract_out_46_, u4_fract_out_47_,
         u4_fract_out_48_, u4_fract_out_49_, u4_fract_out_50_,
         u4_fract_out_51_, u4_exp_out_0_, u4_exp_out_1_, u4_exp_out_2_,
         u4_exp_out_3_, u4_exp_out_4_, u4_exp_out_5_, u4_exp_out_6_,
         u4_exp_out_7_, u4_exp_out_8_, u4_exp_out_9_, u4_exp_out_10_,
         u4_fi_ldz_1_, u4_fi_ldz_2_, u4_fi_ldz_3_, u4_fi_ldz_4_, u4_fi_ldz_5_,
         u4_fi_ldz_6_, n205, n206, n207, n208, n209, n211, n212, n214, n215,
         n216, n217, n218, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n244, n246, n247, n249, n251, n252, n253,
         n255, n257, n258, n259, n260, n261, n262, n263, n264, n266, n267,
         n268, n270, n271, n273, n274, n275, n276, n277, n279, n281, n282,
         n283, n286, n287, n288, n289, n290, n291, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n312, n313, n315, n318, n319, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n341, n342, n343, n345, n346, n348, n349, n350,
         n351, n352, n353, n354, n357, n358, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n374, n375, n376,
         n382, n383, n384, n385, n386, n387, n390, n391, n392, n393, n394,
         n396, n397, n400, n401, n403, n404, n405, n406, n408, n409, n411,
         n412, n413, n416, n417, n418, n419, n420, n421, n424, n425, n426,
         n427, n431, n432, n433, n437, n438, n439, n440, n441, n443, n447,
         n448, n450, n454, n455, n456, n457, n459, n461, n462, n465, n466,
         n467, n471, n472, n478, n480, n481, n482, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n496, n497, n504, n505, n507, n508,
         n510, n511, n512, n513, n514, n515, n518, n519, n523, n524, n525,
         n527, n529, n532, n533, n535, n536, n537, n540, n544, n545, n546,
         n547, n548, n549, n550, n553, n554, n555, n560, n561, n563, n564,
         n566, n567, n568, n572, n573, n576, n579, n581, n583, n584, n585,
         n586, n587, n588, n591, n595, n600, n601, n602, n605, n606, n608,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n638, n639, n640, n642, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n773, n774, n775, n776, n777, n779, n780, n790, n792, n793, n796,
         n798, n799, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n815, n816, n817, n818, n819, n820, n821,
         n823, n825, n827, n828, n829, n830, n831, n833, n834, n835, n836,
         n838, n839, n840, n841, n842, n844, n845, n847, n849, n851, n852,
         n853, n855, n856, n857, n858, n859, n860, n862, n863, n864, n865,
         n866, n868, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n921, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n934, n935, n936, n937, n938,
         n939, n940, n941, n943, n944, n946, n947, n948, n949, n950, n951,
         n952, n955, n960, n965, n971, n974, n986, n993, n994, n1001, n1004,
         n1009, n1012, n1013, n1016, n1019, n1022, n1033, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1048, n1049,
         n1050, n1051, n1052, n1054, n1056, n1057, n1062, n1064, n1066, n1071,
         n1075, n1078, n1079, n1081, n1083, n1084, n1085, n1086, n1087, n1088,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1138, n1140, n1144,
         n1147, n1150, n1153, n1156, n1159, n1162, n1165, n1168, n1171, n1174,
         n1177, n1180, n1183, n1186, n1189, n1192, n1195, n1198, n1201, n1204,
         n1207, n1210, n1211, n1212, n1213, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1310,
         n1312, n1313, n1314, n1317, n1320, n1323, n1326, n1329, n1332, n1335,
         n1338, n1341, n1344, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1364, n1365, n1366, n1367, n1369, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1381, n1382, n1384, n1385, n1386, n1387,
         n1388, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1402, n1404, n1406, n1407, n1408, n1409, n1410, n1412,
         n1413, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1425,
         n1426, n1427, n1428, n1430, n1431, n1432, n1433, n1435, n1436, n1438,
         n1439, n1440, n1441, n1442, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1454, n1455, n1456, n1457, n1460, n1464, n1465, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1475, n1476, n1477, n1480,
         n1481, n1482, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1526, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1541, n1545, n1550, n1554, n1555, n1556, n1557, n1558, n1563,
         n1568, n1573, n1577, n1578, n1579, n1580, n1581, n1586, n1590, n1595,
         n1599, n1600, n1601, n1602, n1603, n1608, n1613, n1618, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1653, n1654,
         n1655, n1656, n1659, n1661, n1662, n1663, n1664, n1666, n1667, n1668,
         n1669, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1698, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1735, n1736, n1737, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1749, n1750, n1751, n1752, n1755, n1756, n1757, n1759,
         n1760, n1761, n1763, n1764, n1766, n1767, n1768, n1769, n1771, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1842, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1923, n1924, n1925, n1926, n1927, n1928,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1981, n1982, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2032, n2033, n2034, n2035,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2071, n2072, n2073, n2075, n2076, n2078, n2079, n2080, n2081,
         n2082, n2083, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2099, n2100, n2101, n2102, n2103,
         n2104, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2122, n2123, n2124, n2126, n2127,
         n2128, n2129, n2130, n2131, n2133, n2134, n2135, n2136, n2138, n2142,
         n2143, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2162, n2163, n2164, n2165, n2166, n2168, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2327, n2328, n2329, n2330,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2341, n2342, n2344,
         n2346, n2348, n2351, n2354, n2356, n2357, n2359, n2361, n2364, n2367,
         n2370, n2372, n2374, n2376, n2378, n2381, n2384, n2386, n2388, n2390,
         n2392, n2395, n2398, n2401, n2403, n2405, n2408, n2411, n2414, n2416,
         n2418, n2420, n2422, n2425, n2428, n2430, n2432, n2434, n2437, n2440,
         n2443, n2445, n2447, n2449, n2451, n2454, n2457, n2459, n2461, n2463,
         n2466, n2469, n2472, n2474, n2476, n2478, n2481, n2483, n2485, n2487,
         n2489, n2491, n2493, n2495, n2497, n2499, n2501, n2503, n2505, n2507,
         n2509, n2511, n2513, n2515, n2517, n2519, n2521, n2523, n2525, n2527,
         n2529, n2532, n2533, n2633, n2636, n2639, n2642, n2645, n2648, n2651,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n3953, n4070, n4123, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4166, n4170, n4173, n4174, n4175, n4177, n4179, n4180, n4181, n4185,
         n4186, n4190, n4193, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4348, n4349, n4350,
         u4_ldz_dif_7_, u4_ldz_dif_6_, u4_ldz_dif_5_, u4_ldz_dif_4_,
         u4_ldz_dif_3_, u4_ldz_dif_2_, u4_ldz_dif_1_, u4_ldz_dif_0_, r482_B_0_,
         u2_lt_131_A_0_, u2_lt_131_A_4_, u2_lt_131_A_5_, u2_lt_131_A_6_,
         u2_lt_131_A_7_, u2_lt_131_A_8_, u2_lt_131_A_9_, u2_gt_141_B_11_,
         u4_sub_461_carry_2_, u4_sub_461_carry_3_, u4_sub_461_carry_4_,
         u4_sub_461_carry_5_, u4_sub_461_carry_6_, u4_sub_466_A_0_,
         u4_sub_466_A_2_, u4_sub_466_A_3_, u4_sub_466_A_4_, u4_sub_466_A_5_,
         u4_sub_466_A_6_, u4_sub_466_A_7_, u4_sub_466_A_8_, u4_sub_466_A_9_,
         u4_sub_466_A_10_, u4_sub_415_carry_2_, u4_sub_415_carry_3_,
         u4_sub_415_carry_4_, u4_sub_415_carry_5_, u4_sub_415_carry_6_,
         u4_sub_415_carry_7_, u4_sub_415_carry_8_, u4_sub_415_carry_9_,
         u4_sub_415_carry_10_, u2_sub_112_carry_2_, u2_sub_112_carry_3_,
         u2_sub_112_carry_4_, u2_sub_112_carry_5_, u2_sub_112_carry_6_,
         u2_sub_112_carry_7_, u2_sub_112_carry_8_, u2_sub_112_carry_9_,
         u2_sub_112_carry_10_, u2_sub_112_carry_11_, u2_add_112_carry_2_,
         u2_add_112_carry_3_, u2_add_112_carry_4_, u2_add_112_carry_5_,
         u2_add_112_carry_6_, u2_add_112_carry_7_, u2_add_112_carry_8_,
         u2_add_112_carry_9_, u2_add_112_carry_10_, u2_add_112_carry_11_,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, u4_sub_471_n14, u4_sub_471_n13,
         u4_sub_471_n12, u4_sub_471_n11, u4_sub_471_n10, u4_sub_471_n9,
         u4_sub_471_n8, u4_sub_471_n7, u4_sub_471_n6, u4_sub_471_n5,
         u4_sub_471_n4, u4_sub_471_n3, u4_sub_471_n2, u4_sub_471_n1,
         u4_sub_471_carry_1_, u4_sub_471_carry_2_, u4_sub_471_carry_3_,
         u4_sub_471_carry_4_, u4_sub_471_carry_5_, u4_sub_471_carry_6_,
         u4_sub_471_carry_7_, u4_sub_471_carry_8_, u4_sub_471_carry_9_,
         u4_sub_471_carry_10_, u4_sub_470_n14, u4_sub_470_n13, u4_sub_470_n12,
         u4_sub_470_n11, u4_sub_470_n10, u4_sub_470_n9, u4_sub_470_n8,
         u4_sub_470_n7, u4_sub_470_n6, u4_sub_470_n5, u4_sub_470_n4,
         u4_sub_470_n3, u4_sub_470_n2, u4_sub_470_n1, u4_sub_470_carry_1_,
         u4_sub_470_carry_2_, u4_sub_470_carry_3_, u4_sub_470_carry_4_,
         u4_sub_470_carry_5_, u4_sub_470_carry_6_, u4_sub_470_carry_7_,
         u4_sub_470_carry_8_, u4_sub_470_carry_9_, u4_sub_470_carry_10_,
         u4_sll_452_n91, u4_sll_452_n90, u4_sll_452_n89, u4_sll_452_n88,
         u4_sll_452_n87, u4_sll_452_n86, u4_sll_452_n85, u4_sll_452_n84,
         u4_sll_452_n83, u4_sll_452_n82, u4_sll_452_n81, u4_sll_452_n80,
         u4_sll_452_n79, u4_sll_452_n78, u4_sll_452_n77, u4_sll_452_n76,
         u4_sll_452_n75, u4_sll_452_n74, u4_sll_452_n73, u4_sll_452_n72,
         u4_sll_452_n71, u4_sll_452_n70, u4_sll_452_n69, u4_sll_452_n68,
         u4_sll_452_n67, u4_sll_452_n66, u4_sll_452_n65, u4_sll_452_n64,
         u4_sll_452_n63, u4_sll_452_n62, u4_sll_452_n61, u4_sll_452_n60,
         u4_sll_452_n59, u4_sll_452_n58, u4_sll_452_n57, u4_sll_452_n56,
         u4_sll_452_n55, u4_sll_452_n54, u4_sll_452_n53, u4_sll_452_n52,
         u4_sll_452_n51, u4_sll_452_n50, u4_sll_452_n49, u4_sll_452_n48,
         u4_sll_452_n47, u4_sll_452_n46, u4_sll_452_n45, u4_sll_452_n44,
         u4_sll_452_n43, u4_sll_452_n42, u4_sll_452_n41, u4_sll_452_n40,
         u4_sll_452_n39, u4_sll_452_n38, u4_sll_452_n37, u4_sll_452_n36,
         u4_sll_452_n35, u4_sll_452_n34, u4_sll_452_n33, u4_sll_452_n32,
         u4_sll_452_n31, u4_sll_452_n30, u4_sll_452_n29, u4_sll_452_n28,
         u4_sll_452_n27, u4_sll_452_n26, u4_sll_452_n25, u4_sll_452_n24,
         u4_sll_452_n23, u4_sll_452_n22, u4_sll_452_n21, u4_sll_452_n20,
         u4_sll_452_n19, u4_sll_452_n18, u4_sll_452_n17, u4_sll_452_n16,
         u4_sll_452_n15, u4_sll_452_n14, u4_sll_452_n13, u4_sll_452_n12,
         u4_sll_452_n11, u4_sll_452_n10, u4_sll_452_n9, u4_sll_452_n8,
         u4_sll_452_n7, u4_sll_452_n6, u4_sll_452_n5, u4_sll_452_n4,
         u4_sll_452_n3, u4_sll_452_n2, u4_sll_452_n1, u4_sll_452_ML_int_7__64_,
         u4_sll_452_ML_int_7__65_, u4_sll_452_ML_int_7__66_,
         u4_sll_452_ML_int_7__67_, u4_sll_452_ML_int_7__68_,
         u4_sll_452_ML_int_7__69_, u4_sll_452_ML_int_7__70_,
         u4_sll_452_ML_int_7__71_, u4_sll_452_ML_int_7__72_,
         u4_sll_452_ML_int_7__73_, u4_sll_452_ML_int_7__74_,
         u4_sll_452_ML_int_7__75_, u4_sll_452_ML_int_7__76_,
         u4_sll_452_ML_int_7__77_, u4_sll_452_ML_int_7__78_,
         u4_sll_452_ML_int_7__79_, u4_sll_452_ML_int_7__80_,
         u4_sll_452_ML_int_7__81_, u4_sll_452_ML_int_7__82_,
         u4_sll_452_ML_int_7__83_, u4_sll_452_ML_int_7__84_,
         u4_sll_452_ML_int_7__85_, u4_sll_452_ML_int_7__86_,
         u4_sll_452_ML_int_7__87_, u4_sll_452_ML_int_7__88_,
         u4_sll_452_ML_int_7__89_, u4_sll_452_ML_int_7__90_,
         u4_sll_452_ML_int_7__91_, u4_sll_452_ML_int_7__92_,
         u4_sll_452_ML_int_7__93_, u4_sll_452_ML_int_7__94_,
         u4_sll_452_ML_int_7__95_, u4_sll_452_ML_int_7__96_,
         u4_sll_452_ML_int_7__97_, u4_sll_452_ML_int_7__98_,
         u4_sll_452_ML_int_7__99_, u4_sll_452_ML_int_7__100_,
         u4_sll_452_ML_int_7__101_, u4_sll_452_ML_int_7__102_,
         u4_sll_452_ML_int_7__103_, u4_sll_452_ML_int_7__104_,
         u4_sll_452_ML_int_7__105_, u4_sll_452_ML_int_6__0_,
         u4_sll_452_ML_int_6__1_, u4_sll_452_ML_int_6__2_,
         u4_sll_452_ML_int_6__3_, u4_sll_452_ML_int_6__4_,
         u4_sll_452_ML_int_6__5_, u4_sll_452_ML_int_6__6_,
         u4_sll_452_ML_int_6__7_, u4_sll_452_ML_int_6__8_,
         u4_sll_452_ML_int_6__9_, u4_sll_452_ML_int_6__10_,
         u4_sll_452_ML_int_6__11_, u4_sll_452_ML_int_6__12_,
         u4_sll_452_ML_int_6__13_, u4_sll_452_ML_int_6__14_,
         u4_sll_452_ML_int_6__15_, u4_sll_452_ML_int_6__16_,
         u4_sll_452_ML_int_6__17_, u4_sll_452_ML_int_6__18_,
         u4_sll_452_ML_int_6__19_, u4_sll_452_ML_int_6__20_,
         u4_sll_452_ML_int_6__21_, u4_sll_452_ML_int_6__22_,
         u4_sll_452_ML_int_6__23_, u4_sll_452_ML_int_6__24_,
         u4_sll_452_ML_int_6__25_, u4_sll_452_ML_int_6__26_,
         u4_sll_452_ML_int_6__27_, u4_sll_452_ML_int_6__28_,
         u4_sll_452_ML_int_6__29_, u4_sll_452_ML_int_6__30_,
         u4_sll_452_ML_int_6__31_, u4_sll_452_ML_int_6__32_,
         u4_sll_452_ML_int_6__33_, u4_sll_452_ML_int_6__34_,
         u4_sll_452_ML_int_6__35_, u4_sll_452_ML_int_6__36_,
         u4_sll_452_ML_int_6__37_, u4_sll_452_ML_int_6__38_,
         u4_sll_452_ML_int_6__39_, u4_sll_452_ML_int_6__40_,
         u4_sll_452_ML_int_6__41_, u4_sll_452_ML_int_6__42_,
         u4_sll_452_ML_int_6__43_, u4_sll_452_ML_int_6__44_,
         u4_sll_452_ML_int_6__45_, u4_sll_452_ML_int_6__46_,
         u4_sll_452_ML_int_6__47_, u4_sll_452_ML_int_6__48_,
         u4_sll_452_ML_int_6__49_, u4_sll_452_ML_int_6__50_,
         u4_sll_452_ML_int_6__51_, u4_sll_452_ML_int_6__52_,
         u4_sll_452_ML_int_6__53_, u4_sll_452_ML_int_6__54_,
         u4_sll_452_ML_int_6__55_, u4_sll_452_ML_int_6__56_,
         u4_sll_452_ML_int_6__57_, u4_sll_452_ML_int_6__58_,
         u4_sll_452_ML_int_6__59_, u4_sll_452_ML_int_6__60_,
         u4_sll_452_ML_int_6__61_, u4_sll_452_ML_int_6__62_,
         u4_sll_452_ML_int_6__63_, u4_sll_452_ML_int_6__64_,
         u4_sll_452_ML_int_6__65_, u4_sll_452_ML_int_6__66_,
         u4_sll_452_ML_int_6__67_, u4_sll_452_ML_int_6__68_,
         u4_sll_452_ML_int_6__69_, u4_sll_452_ML_int_6__70_,
         u4_sll_452_ML_int_6__71_, u4_sll_452_ML_int_6__72_,
         u4_sll_452_ML_int_6__73_, u4_sll_452_ML_int_6__74_,
         u4_sll_452_ML_int_6__75_, u4_sll_452_ML_int_6__76_,
         u4_sll_452_ML_int_6__77_, u4_sll_452_ML_int_6__78_,
         u4_sll_452_ML_int_6__79_, u4_sll_452_ML_int_6__80_,
         u4_sll_452_ML_int_6__81_, u4_sll_452_ML_int_6__82_,
         u4_sll_452_ML_int_6__83_, u4_sll_452_ML_int_6__84_,
         u4_sll_452_ML_int_6__85_, u4_sll_452_ML_int_6__86_,
         u4_sll_452_ML_int_6__87_, u4_sll_452_ML_int_6__88_,
         u4_sll_452_ML_int_6__89_, u4_sll_452_ML_int_6__90_,
         u4_sll_452_ML_int_6__91_, u4_sll_452_ML_int_6__92_,
         u4_sll_452_ML_int_6__93_, u4_sll_452_ML_int_6__94_,
         u4_sll_452_ML_int_6__95_, u4_sll_452_ML_int_6__96_,
         u4_sll_452_ML_int_6__97_, u4_sll_452_ML_int_6__98_,
         u4_sll_452_ML_int_6__99_, u4_sll_452_ML_int_6__100_,
         u4_sll_452_ML_int_6__101_, u4_sll_452_ML_int_6__102_,
         u4_sll_452_ML_int_6__103_, u4_sll_452_ML_int_6__104_,
         u4_sll_452_ML_int_6__105_, u4_sll_452_ML_int_5__0_,
         u4_sll_452_ML_int_5__1_, u4_sll_452_ML_int_5__2_,
         u4_sll_452_ML_int_5__3_, u4_sll_452_ML_int_5__4_,
         u4_sll_452_ML_int_5__5_, u4_sll_452_ML_int_5__6_,
         u4_sll_452_ML_int_5__7_, u4_sll_452_ML_int_5__8_,
         u4_sll_452_ML_int_5__9_, u4_sll_452_ML_int_5__10_,
         u4_sll_452_ML_int_5__11_, u4_sll_452_ML_int_5__12_,
         u4_sll_452_ML_int_5__13_, u4_sll_452_ML_int_5__14_,
         u4_sll_452_ML_int_5__15_, u4_sll_452_ML_int_5__16_,
         u4_sll_452_ML_int_5__17_, u4_sll_452_ML_int_5__18_,
         u4_sll_452_ML_int_5__19_, u4_sll_452_ML_int_5__20_,
         u4_sll_452_ML_int_5__21_, u4_sll_452_ML_int_5__22_,
         u4_sll_452_ML_int_5__23_, u4_sll_452_ML_int_5__24_,
         u4_sll_452_ML_int_5__25_, u4_sll_452_ML_int_5__26_,
         u4_sll_452_ML_int_5__27_, u4_sll_452_ML_int_5__28_,
         u4_sll_452_ML_int_5__29_, u4_sll_452_ML_int_5__30_,
         u4_sll_452_ML_int_5__31_, u4_sll_452_ML_int_5__32_,
         u4_sll_452_ML_int_5__33_, u4_sll_452_ML_int_5__34_,
         u4_sll_452_ML_int_5__35_, u4_sll_452_ML_int_5__36_,
         u4_sll_452_ML_int_5__37_, u4_sll_452_ML_int_5__38_,
         u4_sll_452_ML_int_5__39_, u4_sll_452_ML_int_5__40_,
         u4_sll_452_ML_int_5__41_, u4_sll_452_ML_int_5__42_,
         u4_sll_452_ML_int_5__43_, u4_sll_452_ML_int_5__44_,
         u4_sll_452_ML_int_5__45_, u4_sll_452_ML_int_5__46_,
         u4_sll_452_ML_int_5__47_, u4_sll_452_ML_int_5__48_,
         u4_sll_452_ML_int_5__49_, u4_sll_452_ML_int_5__50_,
         u4_sll_452_ML_int_5__51_, u4_sll_452_ML_int_5__52_,
         u4_sll_452_ML_int_5__53_, u4_sll_452_ML_int_5__54_,
         u4_sll_452_ML_int_5__55_, u4_sll_452_ML_int_5__56_,
         u4_sll_452_ML_int_5__57_, u4_sll_452_ML_int_5__58_,
         u4_sll_452_ML_int_5__59_, u4_sll_452_ML_int_5__60_,
         u4_sll_452_ML_int_5__61_, u4_sll_452_ML_int_5__62_,
         u4_sll_452_ML_int_5__63_, u4_sll_452_ML_int_5__64_,
         u4_sll_452_ML_int_5__65_, u4_sll_452_ML_int_5__66_,
         u4_sll_452_ML_int_5__67_, u4_sll_452_ML_int_5__68_,
         u4_sll_452_ML_int_5__69_, u4_sll_452_ML_int_5__70_,
         u4_sll_452_ML_int_5__71_, u4_sll_452_ML_int_5__72_,
         u4_sll_452_ML_int_5__73_, u4_sll_452_ML_int_5__74_,
         u4_sll_452_ML_int_5__75_, u4_sll_452_ML_int_5__76_,
         u4_sll_452_ML_int_5__77_, u4_sll_452_ML_int_5__78_,
         u4_sll_452_ML_int_5__79_, u4_sll_452_ML_int_5__80_,
         u4_sll_452_ML_int_5__81_, u4_sll_452_ML_int_5__82_,
         u4_sll_452_ML_int_5__83_, u4_sll_452_ML_int_5__84_,
         u4_sll_452_ML_int_5__85_, u4_sll_452_ML_int_5__86_,
         u4_sll_452_ML_int_5__87_, u4_sll_452_ML_int_5__88_,
         u4_sll_452_ML_int_5__89_, u4_sll_452_ML_int_5__90_,
         u4_sll_452_ML_int_5__91_, u4_sll_452_ML_int_5__92_,
         u4_sll_452_ML_int_5__93_, u4_sll_452_ML_int_5__94_,
         u4_sll_452_ML_int_5__95_, u4_sll_452_ML_int_5__96_,
         u4_sll_452_ML_int_5__97_, u4_sll_452_ML_int_5__98_,
         u4_sll_452_ML_int_5__99_, u4_sll_452_ML_int_5__100_,
         u4_sll_452_ML_int_5__101_, u4_sll_452_ML_int_5__102_,
         u4_sll_452_ML_int_5__103_, u4_sll_452_ML_int_5__104_,
         u4_sll_452_ML_int_5__105_, u4_sll_452_ML_int_4__0_,
         u4_sll_452_ML_int_4__1_, u4_sll_452_ML_int_4__2_,
         u4_sll_452_ML_int_4__3_, u4_sll_452_ML_int_4__4_,
         u4_sll_452_ML_int_4__5_, u4_sll_452_ML_int_4__6_,
         u4_sll_452_ML_int_4__7_, u4_sll_452_ML_int_4__8_,
         u4_sll_452_ML_int_4__9_, u4_sll_452_ML_int_4__10_,
         u4_sll_452_ML_int_4__11_, u4_sll_452_ML_int_4__12_,
         u4_sll_452_ML_int_4__13_, u4_sll_452_ML_int_4__14_,
         u4_sll_452_ML_int_4__15_, u4_sll_452_ML_int_4__16_,
         u4_sll_452_ML_int_4__17_, u4_sll_452_ML_int_4__18_,
         u4_sll_452_ML_int_4__19_, u4_sll_452_ML_int_4__20_,
         u4_sll_452_ML_int_4__21_, u4_sll_452_ML_int_4__22_,
         u4_sll_452_ML_int_4__23_, u4_sll_452_ML_int_4__24_,
         u4_sll_452_ML_int_4__25_, u4_sll_452_ML_int_4__26_,
         u4_sll_452_ML_int_4__27_, u4_sll_452_ML_int_4__28_,
         u4_sll_452_ML_int_4__29_, u4_sll_452_ML_int_4__30_,
         u4_sll_452_ML_int_4__31_, u4_sll_452_ML_int_4__32_,
         u4_sll_452_ML_int_4__33_, u4_sll_452_ML_int_4__34_,
         u4_sll_452_ML_int_4__35_, u4_sll_452_ML_int_4__36_,
         u4_sll_452_ML_int_4__37_, u4_sll_452_ML_int_4__38_,
         u4_sll_452_ML_int_4__39_, u4_sll_452_ML_int_4__40_,
         u4_sll_452_ML_int_4__41_, u4_sll_452_ML_int_4__42_,
         u4_sll_452_ML_int_4__43_, u4_sll_452_ML_int_4__44_,
         u4_sll_452_ML_int_4__45_, u4_sll_452_ML_int_4__46_,
         u4_sll_452_ML_int_4__47_, u4_sll_452_ML_int_4__48_,
         u4_sll_452_ML_int_4__49_, u4_sll_452_ML_int_4__50_,
         u4_sll_452_ML_int_4__51_, u4_sll_452_ML_int_4__52_,
         u4_sll_452_ML_int_4__53_, u4_sll_452_ML_int_4__54_,
         u4_sll_452_ML_int_4__55_, u4_sll_452_ML_int_4__56_,
         u4_sll_452_ML_int_4__57_, u4_sll_452_ML_int_4__58_,
         u4_sll_452_ML_int_4__59_, u4_sll_452_ML_int_4__60_,
         u4_sll_452_ML_int_4__61_, u4_sll_452_ML_int_4__62_,
         u4_sll_452_ML_int_4__63_, u4_sll_452_ML_int_4__64_,
         u4_sll_452_ML_int_4__65_, u4_sll_452_ML_int_4__66_,
         u4_sll_452_ML_int_4__67_, u4_sll_452_ML_int_4__68_,
         u4_sll_452_ML_int_4__69_, u4_sll_452_ML_int_4__70_,
         u4_sll_452_ML_int_4__71_, u4_sll_452_ML_int_4__72_,
         u4_sll_452_ML_int_4__73_, u4_sll_452_ML_int_4__74_,
         u4_sll_452_ML_int_4__75_, u4_sll_452_ML_int_4__76_,
         u4_sll_452_ML_int_4__77_, u4_sll_452_ML_int_4__78_,
         u4_sll_452_ML_int_4__79_, u4_sll_452_ML_int_4__80_,
         u4_sll_452_ML_int_4__81_, u4_sll_452_ML_int_4__82_,
         u4_sll_452_ML_int_4__83_, u4_sll_452_ML_int_4__84_,
         u4_sll_452_ML_int_4__85_, u4_sll_452_ML_int_4__86_,
         u4_sll_452_ML_int_4__87_, u4_sll_452_ML_int_4__88_,
         u4_sll_452_ML_int_4__89_, u4_sll_452_ML_int_4__90_,
         u4_sll_452_ML_int_4__91_, u4_sll_452_ML_int_4__92_,
         u4_sll_452_ML_int_4__93_, u4_sll_452_ML_int_4__94_,
         u4_sll_452_ML_int_4__95_, u4_sll_452_ML_int_4__96_,
         u4_sll_452_ML_int_4__97_, u4_sll_452_ML_int_4__98_,
         u4_sll_452_ML_int_4__99_, u4_sll_452_ML_int_4__100_,
         u4_sll_452_ML_int_4__101_, u4_sll_452_ML_int_4__102_,
         u4_sll_452_ML_int_4__103_, u4_sll_452_ML_int_4__104_,
         u4_sll_452_ML_int_4__105_, u4_sll_452_ML_int_3__0_,
         u4_sll_452_ML_int_3__1_, u4_sll_452_ML_int_3__2_,
         u4_sll_452_ML_int_3__3_, u4_sll_452_ML_int_3__4_,
         u4_sll_452_ML_int_3__5_, u4_sll_452_ML_int_3__6_,
         u4_sll_452_ML_int_3__7_, u4_sll_452_ML_int_3__8_,
         u4_sll_452_ML_int_3__9_, u4_sll_452_ML_int_3__10_,
         u4_sll_452_ML_int_3__11_, u4_sll_452_ML_int_3__12_,
         u4_sll_452_ML_int_3__13_, u4_sll_452_ML_int_3__14_,
         u4_sll_452_ML_int_3__15_, u4_sll_452_ML_int_3__16_,
         u4_sll_452_ML_int_3__17_, u4_sll_452_ML_int_3__18_,
         u4_sll_452_ML_int_3__19_, u4_sll_452_ML_int_3__20_,
         u4_sll_452_ML_int_3__21_, u4_sll_452_ML_int_3__22_,
         u4_sll_452_ML_int_3__23_, u4_sll_452_ML_int_3__24_,
         u4_sll_452_ML_int_3__25_, u4_sll_452_ML_int_3__26_,
         u4_sll_452_ML_int_3__27_, u4_sll_452_ML_int_3__28_,
         u4_sll_452_ML_int_3__29_, u4_sll_452_ML_int_3__30_,
         u4_sll_452_ML_int_3__31_, u4_sll_452_ML_int_3__32_,
         u4_sll_452_ML_int_3__33_, u4_sll_452_ML_int_3__34_,
         u4_sll_452_ML_int_3__35_, u4_sll_452_ML_int_3__36_,
         u4_sll_452_ML_int_3__37_, u4_sll_452_ML_int_3__38_,
         u4_sll_452_ML_int_3__39_, u4_sll_452_ML_int_3__40_,
         u4_sll_452_ML_int_3__41_, u4_sll_452_ML_int_3__42_,
         u4_sll_452_ML_int_3__43_, u4_sll_452_ML_int_3__44_,
         u4_sll_452_ML_int_3__45_, u4_sll_452_ML_int_3__46_,
         u4_sll_452_ML_int_3__47_, u4_sll_452_ML_int_3__48_,
         u4_sll_452_ML_int_3__49_, u4_sll_452_ML_int_3__50_,
         u4_sll_452_ML_int_3__51_, u4_sll_452_ML_int_3__52_,
         u4_sll_452_ML_int_3__53_, u4_sll_452_ML_int_3__54_,
         u4_sll_452_ML_int_3__55_, u4_sll_452_ML_int_3__56_,
         u4_sll_452_ML_int_3__57_, u4_sll_452_ML_int_3__58_,
         u4_sll_452_ML_int_3__59_, u4_sll_452_ML_int_3__60_,
         u4_sll_452_ML_int_3__61_, u4_sll_452_ML_int_3__62_,
         u4_sll_452_ML_int_3__63_, u4_sll_452_ML_int_3__64_,
         u4_sll_452_ML_int_3__65_, u4_sll_452_ML_int_3__66_,
         u4_sll_452_ML_int_3__67_, u4_sll_452_ML_int_3__68_,
         u4_sll_452_ML_int_3__69_, u4_sll_452_ML_int_3__70_,
         u4_sll_452_ML_int_3__71_, u4_sll_452_ML_int_3__72_,
         u4_sll_452_ML_int_3__73_, u4_sll_452_ML_int_3__74_,
         u4_sll_452_ML_int_3__75_, u4_sll_452_ML_int_3__76_,
         u4_sll_452_ML_int_3__77_, u4_sll_452_ML_int_3__78_,
         u4_sll_452_ML_int_3__79_, u4_sll_452_ML_int_3__80_,
         u4_sll_452_ML_int_3__81_, u4_sll_452_ML_int_3__82_,
         u4_sll_452_ML_int_3__83_, u4_sll_452_ML_int_3__84_,
         u4_sll_452_ML_int_3__85_, u4_sll_452_ML_int_3__86_,
         u4_sll_452_ML_int_3__87_, u4_sll_452_ML_int_3__88_,
         u4_sll_452_ML_int_3__89_, u4_sll_452_ML_int_3__90_,
         u4_sll_452_ML_int_3__91_, u4_sll_452_ML_int_3__92_,
         u4_sll_452_ML_int_3__93_, u4_sll_452_ML_int_3__94_,
         u4_sll_452_ML_int_3__95_, u4_sll_452_ML_int_3__96_,
         u4_sll_452_ML_int_3__97_, u4_sll_452_ML_int_3__98_,
         u4_sll_452_ML_int_3__99_, u4_sll_452_ML_int_3__100_,
         u4_sll_452_ML_int_3__101_, u4_sll_452_ML_int_3__102_,
         u4_sll_452_ML_int_3__103_, u4_sll_452_ML_int_3__104_,
         u4_sll_452_ML_int_3__105_, u4_sll_452_ML_int_2__0_,
         u4_sll_452_ML_int_2__1_, u4_sll_452_ML_int_2__2_,
         u4_sll_452_ML_int_2__3_, u4_sll_452_ML_int_2__4_,
         u4_sll_452_ML_int_2__5_, u4_sll_452_ML_int_2__6_,
         u4_sll_452_ML_int_2__7_, u4_sll_452_ML_int_2__8_,
         u4_sll_452_ML_int_2__9_, u4_sll_452_ML_int_2__10_,
         u4_sll_452_ML_int_2__11_, u4_sll_452_ML_int_2__12_,
         u4_sll_452_ML_int_2__13_, u4_sll_452_ML_int_2__14_,
         u4_sll_452_ML_int_2__15_, u4_sll_452_ML_int_2__16_,
         u4_sll_452_ML_int_2__17_, u4_sll_452_ML_int_2__18_,
         u4_sll_452_ML_int_2__19_, u4_sll_452_ML_int_2__20_,
         u4_sll_452_ML_int_2__21_, u4_sll_452_ML_int_2__22_,
         u4_sll_452_ML_int_2__23_, u4_sll_452_ML_int_2__24_,
         u4_sll_452_ML_int_2__25_, u4_sll_452_ML_int_2__26_,
         u4_sll_452_ML_int_2__27_, u4_sll_452_ML_int_2__28_,
         u4_sll_452_ML_int_2__29_, u4_sll_452_ML_int_2__30_,
         u4_sll_452_ML_int_2__31_, u4_sll_452_ML_int_2__32_,
         u4_sll_452_ML_int_2__33_, u4_sll_452_ML_int_2__34_,
         u4_sll_452_ML_int_2__35_, u4_sll_452_ML_int_2__36_,
         u4_sll_452_ML_int_2__37_, u4_sll_452_ML_int_2__38_,
         u4_sll_452_ML_int_2__39_, u4_sll_452_ML_int_2__40_,
         u4_sll_452_ML_int_2__41_, u4_sll_452_ML_int_2__42_,
         u4_sll_452_ML_int_2__43_, u4_sll_452_ML_int_2__44_,
         u4_sll_452_ML_int_2__45_, u4_sll_452_ML_int_2__46_,
         u4_sll_452_ML_int_2__47_, u4_sll_452_ML_int_2__48_,
         u4_sll_452_ML_int_2__49_, u4_sll_452_ML_int_2__50_,
         u4_sll_452_ML_int_2__51_, u4_sll_452_ML_int_2__52_,
         u4_sll_452_ML_int_2__53_, u4_sll_452_ML_int_2__54_,
         u4_sll_452_ML_int_2__55_, u4_sll_452_ML_int_2__56_,
         u4_sll_452_ML_int_2__57_, u4_sll_452_ML_int_2__58_,
         u4_sll_452_ML_int_2__59_, u4_sll_452_ML_int_2__60_,
         u4_sll_452_ML_int_2__61_, u4_sll_452_ML_int_2__62_,
         u4_sll_452_ML_int_2__63_, u4_sll_452_ML_int_2__64_,
         u4_sll_452_ML_int_2__65_, u4_sll_452_ML_int_2__66_,
         u4_sll_452_ML_int_2__67_, u4_sll_452_ML_int_2__68_,
         u4_sll_452_ML_int_2__69_, u4_sll_452_ML_int_2__70_,
         u4_sll_452_ML_int_2__71_, u4_sll_452_ML_int_2__72_,
         u4_sll_452_ML_int_2__73_, u4_sll_452_ML_int_2__74_,
         u4_sll_452_ML_int_2__75_, u4_sll_452_ML_int_2__76_,
         u4_sll_452_ML_int_2__77_, u4_sll_452_ML_int_2__78_,
         u4_sll_452_ML_int_2__79_, u4_sll_452_ML_int_2__80_,
         u4_sll_452_ML_int_2__81_, u4_sll_452_ML_int_2__82_,
         u4_sll_452_ML_int_2__83_, u4_sll_452_ML_int_2__84_,
         u4_sll_452_ML_int_2__85_, u4_sll_452_ML_int_2__86_,
         u4_sll_452_ML_int_2__87_, u4_sll_452_ML_int_2__88_,
         u4_sll_452_ML_int_2__89_, u4_sll_452_ML_int_2__90_,
         u4_sll_452_ML_int_2__91_, u4_sll_452_ML_int_2__92_,
         u4_sll_452_ML_int_2__93_, u4_sll_452_ML_int_2__94_,
         u4_sll_452_ML_int_2__95_, u4_sll_452_ML_int_2__96_,
         u4_sll_452_ML_int_2__97_, u4_sll_452_ML_int_2__98_,
         u4_sll_452_ML_int_2__99_, u4_sll_452_ML_int_2__100_,
         u4_sll_452_ML_int_2__101_, u4_sll_452_ML_int_2__102_,
         u4_sll_452_ML_int_2__103_, u4_sll_452_ML_int_2__104_,
         u4_sll_452_ML_int_2__105_, u4_sll_452_ML_int_1__0_,
         u4_sll_452_ML_int_1__1_, u4_sll_452_ML_int_1__2_,
         u4_sll_452_ML_int_1__3_, u4_sll_452_ML_int_1__4_,
         u4_sll_452_ML_int_1__5_, u4_sll_452_ML_int_1__6_,
         u4_sll_452_ML_int_1__7_, u4_sll_452_ML_int_1__8_,
         u4_sll_452_ML_int_1__9_, u4_sll_452_ML_int_1__10_,
         u4_sll_452_ML_int_1__11_, u4_sll_452_ML_int_1__12_,
         u4_sll_452_ML_int_1__13_, u4_sll_452_ML_int_1__14_,
         u4_sll_452_ML_int_1__15_, u4_sll_452_ML_int_1__16_,
         u4_sll_452_ML_int_1__17_, u4_sll_452_ML_int_1__18_,
         u4_sll_452_ML_int_1__19_, u4_sll_452_ML_int_1__20_,
         u4_sll_452_ML_int_1__21_, u4_sll_452_ML_int_1__22_,
         u4_sll_452_ML_int_1__23_, u4_sll_452_ML_int_1__24_,
         u4_sll_452_ML_int_1__25_, u4_sll_452_ML_int_1__26_,
         u4_sll_452_ML_int_1__27_, u4_sll_452_ML_int_1__28_,
         u4_sll_452_ML_int_1__29_, u4_sll_452_ML_int_1__30_,
         u4_sll_452_ML_int_1__31_, u4_sll_452_ML_int_1__32_,
         u4_sll_452_ML_int_1__33_, u4_sll_452_ML_int_1__34_,
         u4_sll_452_ML_int_1__35_, u4_sll_452_ML_int_1__36_,
         u4_sll_452_ML_int_1__37_, u4_sll_452_ML_int_1__38_,
         u4_sll_452_ML_int_1__39_, u4_sll_452_ML_int_1__40_,
         u4_sll_452_ML_int_1__41_, u4_sll_452_ML_int_1__42_,
         u4_sll_452_ML_int_1__43_, u4_sll_452_ML_int_1__44_,
         u4_sll_452_ML_int_1__45_, u4_sll_452_ML_int_1__46_,
         u4_sll_452_ML_int_1__47_, u4_sll_452_ML_int_1__48_,
         u4_sll_452_ML_int_1__49_, u4_sll_452_ML_int_1__50_,
         u4_sll_452_ML_int_1__51_, u4_sll_452_ML_int_1__52_,
         u4_sll_452_ML_int_1__53_, u4_sll_452_ML_int_1__54_,
         u4_sll_452_ML_int_1__55_, u4_sll_452_ML_int_1__56_,
         u4_sll_452_ML_int_1__57_, u4_sll_452_ML_int_1__58_,
         u4_sll_452_ML_int_1__59_, u4_sll_452_ML_int_1__60_,
         u4_sll_452_ML_int_1__61_, u4_sll_452_ML_int_1__62_,
         u4_sll_452_ML_int_1__63_, u4_sll_452_ML_int_1__64_,
         u4_sll_452_ML_int_1__65_, u4_sll_452_ML_int_1__66_,
         u4_sll_452_ML_int_1__67_, u4_sll_452_ML_int_1__68_,
         u4_sll_452_ML_int_1__69_, u4_sll_452_ML_int_1__70_,
         u4_sll_452_ML_int_1__71_, u4_sll_452_ML_int_1__72_,
         u4_sll_452_ML_int_1__73_, u4_sll_452_ML_int_1__74_,
         u4_sll_452_ML_int_1__75_, u4_sll_452_ML_int_1__76_,
         u4_sll_452_ML_int_1__77_, u4_sll_452_ML_int_1__78_,
         u4_sll_452_ML_int_1__79_, u4_sll_452_ML_int_1__80_,
         u4_sll_452_ML_int_1__81_, u4_sll_452_ML_int_1__82_,
         u4_sll_452_ML_int_1__83_, u4_sll_452_ML_int_1__84_,
         u4_sll_452_ML_int_1__85_, u4_sll_452_ML_int_1__86_,
         u4_sll_452_ML_int_1__87_, u4_sll_452_ML_int_1__88_,
         u4_sll_452_ML_int_1__89_, u4_sll_452_ML_int_1__90_,
         u4_sll_452_ML_int_1__91_, u4_sll_452_ML_int_1__92_,
         u4_sll_452_ML_int_1__93_, u4_sll_452_ML_int_1__94_,
         u4_sll_452_ML_int_1__95_, u4_sll_452_ML_int_1__96_,
         u4_sll_452_ML_int_1__97_, u4_sll_452_ML_int_1__98_,
         u4_sll_452_ML_int_1__99_, u4_sll_452_ML_int_1__100_,
         u4_sll_452_ML_int_1__101_, u4_sll_452_ML_int_1__102_,
         u4_sll_452_ML_int_1__103_, u4_sll_452_ML_int_1__104_,
         u4_sll_452_ML_int_1__105_, u4_sll_452_SHMAG_0_, u4_sll_452_SHMAG_1_,
         u4_sll_452_SHMAG_2_, u4_sll_452_SHMAG_3_, u4_sll_452_SHMAG_4_,
         u4_sll_452_SHMAG_6_, u4_sll_452_temp_int_SH_5_, u4_srl_451_n883,
         u4_srl_451_n882, u4_srl_451_n881, u4_srl_451_n880, u4_srl_451_n879,
         u4_srl_451_n878, u4_srl_451_n877, u4_srl_451_n876, u4_srl_451_n875,
         u4_srl_451_n874, u4_srl_451_n873, u4_srl_451_n872, u4_srl_451_n871,
         u4_srl_451_n870, u4_srl_451_n869, u4_srl_451_n868, u4_srl_451_n867,
         u4_srl_451_n866, u4_srl_451_n865, u4_srl_451_n864, u4_srl_451_n863,
         u4_srl_451_n862, u4_srl_451_n861, u4_srl_451_n860, u4_srl_451_n859,
         u4_srl_451_n858, u4_srl_451_n857, u4_srl_451_n856, u4_srl_451_n855,
         u4_srl_451_n854, u4_srl_451_n853, u4_srl_451_n852, u4_srl_451_n851,
         u4_srl_451_n850, u4_srl_451_n849, u4_srl_451_n848, u4_srl_451_n847,
         u4_srl_451_n846, u4_srl_451_n845, u4_srl_451_n844, u4_srl_451_n843,
         u4_srl_451_n842, u4_srl_451_n841, u4_srl_451_n840, u4_srl_451_n839,
         u4_srl_451_n838, u4_srl_451_n837, u4_srl_451_n836, u4_srl_451_n835,
         u4_srl_451_n834, u4_srl_451_n833, u4_srl_451_n832, u4_srl_451_n831,
         u4_srl_451_n830, u4_srl_451_n829, u4_srl_451_n828, u4_srl_451_n827,
         u4_srl_451_n826, u4_srl_451_n825, u4_srl_451_n824, u4_srl_451_n823,
         u4_srl_451_n822, u4_srl_451_n821, u4_srl_451_n820, u4_srl_451_n819,
         u4_srl_451_n818, u4_srl_451_n817, u4_srl_451_n816, u4_srl_451_n815,
         u4_srl_451_n814, u4_srl_451_n813, u4_srl_451_n812, u4_srl_451_n811,
         u4_srl_451_n810, u4_srl_451_n809, u4_srl_451_n808, u4_srl_451_n807,
         u4_srl_451_n806, u4_srl_451_n805, u4_srl_451_n804, u4_srl_451_n803,
         u4_srl_451_n802, u4_srl_451_n801, u4_srl_451_n800, u4_srl_451_n799,
         u4_srl_451_n798, u4_srl_451_n797, u4_srl_451_n796, u4_srl_451_n795,
         u4_srl_451_n794, u4_srl_451_n793, u4_srl_451_n792, u4_srl_451_n791,
         u4_srl_451_n790, u4_srl_451_n789, u4_srl_451_n788, u4_srl_451_n787,
         u4_srl_451_n786, u4_srl_451_n785, u4_srl_451_n784, u4_srl_451_n783,
         u4_srl_451_n782, u4_srl_451_n781, u4_srl_451_n780, u4_srl_451_n779,
         u4_srl_451_n778, u4_srl_451_n777, u4_srl_451_n776, u4_srl_451_n775,
         u4_srl_451_n774, u4_srl_451_n773, u4_srl_451_n772, u4_srl_451_n771,
         u4_srl_451_n770, u4_srl_451_n769, u4_srl_451_n768, u4_srl_451_n767,
         u4_srl_451_n766, u4_srl_451_n765, u4_srl_451_n764, u4_srl_451_n763,
         u4_srl_451_n762, u4_srl_451_n761, u4_srl_451_n760, u4_srl_451_n759,
         u4_srl_451_n758, u4_srl_451_n757, u4_srl_451_n756, u4_srl_451_n755,
         u4_srl_451_n754, u4_srl_451_n753, u4_srl_451_n752, u4_srl_451_n751,
         u4_srl_451_n750, u4_srl_451_n749, u4_srl_451_n748, u4_srl_451_n747,
         u4_srl_451_n746, u4_srl_451_n745, u4_srl_451_n744, u4_srl_451_n743,
         u4_srl_451_n742, u4_srl_451_n741, u4_srl_451_n740, u4_srl_451_n739,
         u4_srl_451_n738, u4_srl_451_n737, u4_srl_451_n736, u4_srl_451_n735,
         u4_srl_451_n734, u4_srl_451_n733, u4_srl_451_n732, u4_srl_451_n731,
         u4_srl_451_n730, u4_srl_451_n729, u4_srl_451_n728, u4_srl_451_n727,
         u4_srl_451_n726, u4_srl_451_n725, u4_srl_451_n724, u4_srl_451_n723,
         u4_srl_451_n722, u4_srl_451_n721, u4_srl_451_n720, u4_srl_451_n719,
         u4_srl_451_n718, u4_srl_451_n717, u4_srl_451_n716, u4_srl_451_n715,
         u4_srl_451_n714, u4_srl_451_n713, u4_srl_451_n712, u4_srl_451_n711,
         u4_srl_451_n710, u4_srl_451_n709, u4_srl_451_n708, u4_srl_451_n707,
         u4_srl_451_n706, u4_srl_451_n705, u4_srl_451_n704, u4_srl_451_n703,
         u4_srl_451_n702, u4_srl_451_n701, u4_srl_451_n700, u4_srl_451_n699,
         u4_srl_451_n698, u4_srl_451_n697, u4_srl_451_n696, u4_srl_451_n695,
         u4_srl_451_n694, u4_srl_451_n693, u4_srl_451_n692, u4_srl_451_n691,
         u4_srl_451_n690, u4_srl_451_n689, u4_srl_451_n688, u4_srl_451_n687,
         u4_srl_451_n686, u4_srl_451_n685, u4_srl_451_n684, u4_srl_451_n683,
         u4_srl_451_n682, u4_srl_451_n681, u4_srl_451_n680, u4_srl_451_n679,
         u4_srl_451_n678, u4_srl_451_n677, u4_srl_451_n676, u4_srl_451_n675,
         u4_srl_451_n674, u4_srl_451_n673, u4_srl_451_n672, u4_srl_451_n671,
         u4_srl_451_n670, u4_srl_451_n669, u4_srl_451_n668, u4_srl_451_n667,
         u4_srl_451_n666, u4_srl_451_n665, u4_srl_451_n664, u4_srl_451_n663,
         u4_srl_451_n662, u4_srl_451_n661, u4_srl_451_n660, u4_srl_451_n659,
         u4_srl_451_n658, u4_srl_451_n657, u4_srl_451_n656, u4_srl_451_n655,
         u4_srl_451_n654, u4_srl_451_n653, u4_srl_451_n652, u4_srl_451_n651,
         u4_srl_451_n650, u4_srl_451_n649, u4_srl_451_n648, u4_srl_451_n647,
         u4_srl_451_n646, u4_srl_451_n645, u4_srl_451_n644, u4_srl_451_n643,
         u4_srl_451_n642, u4_srl_451_n641, u4_srl_451_n640, u4_srl_451_n639,
         u4_srl_451_n638, u4_srl_451_n637, u4_srl_451_n636, u4_srl_451_n635,
         u4_srl_451_n634, u4_srl_451_n633, u4_srl_451_n632, u4_srl_451_n631,
         u4_srl_451_n630, u4_srl_451_n629, u4_srl_451_n628, u4_srl_451_n627,
         u4_srl_451_n626, u4_srl_451_n625, u4_srl_451_n624, u4_srl_451_n623,
         u4_srl_451_n622, u4_srl_451_n621, u4_srl_451_n620, u4_srl_451_n619,
         u4_srl_451_n618, u4_srl_451_n617, u4_srl_451_n616, u4_srl_451_n615,
         u4_srl_451_n614, u4_srl_451_n613, u4_srl_451_n612, u4_srl_451_n611,
         u4_srl_451_n610, u4_srl_451_n609, u4_srl_451_n608, u4_srl_451_n607,
         u4_srl_451_n606, u4_srl_451_n605, u4_srl_451_n604, u4_srl_451_n603,
         u4_srl_451_n602, u4_srl_451_n601, u4_srl_451_n600, u4_srl_451_n599,
         u4_srl_451_n598, u4_srl_451_n597, u4_srl_451_n596, u4_srl_451_n595,
         u4_srl_451_n594, u4_srl_451_n593, u4_srl_451_n592, u4_srl_451_n591,
         u4_srl_451_n590, u4_srl_451_n589, u4_srl_451_n588, u4_srl_451_n587,
         u4_srl_451_n586, u4_srl_451_n585, u4_srl_451_n584, u4_srl_451_n583,
         u4_srl_451_n582, u4_srl_451_n581, u4_srl_451_n580, u4_srl_451_n579,
         u4_srl_451_n578, u4_srl_451_n577, u4_srl_451_n576, u4_srl_451_n575,
         u4_srl_451_n574, u4_srl_451_n573, u4_srl_451_n572, u4_srl_451_n571,
         u4_srl_451_n570, u4_srl_451_n569, u4_srl_451_n568, u4_srl_451_n567,
         u4_srl_451_n566, u4_srl_451_n565, u4_srl_451_n564, u4_srl_451_n563,
         u4_srl_451_n562, u4_srl_451_n561, u4_srl_451_n560, u4_srl_451_n559,
         u4_srl_451_n558, u4_srl_451_n557, u4_srl_451_n556, u4_srl_451_n555,
         u4_srl_451_n554, u4_srl_451_n553, u4_srl_451_n552, u4_srl_451_n551,
         u4_srl_451_n550, u4_srl_451_n549, u4_srl_451_n548, u4_srl_451_n547,
         u4_srl_451_n546, u4_srl_451_n545, u4_srl_451_n544, u4_srl_451_n543,
         u4_srl_451_n542, u4_srl_451_n541, u4_srl_451_n540, u4_srl_451_n539,
         u4_srl_451_n538, u4_srl_451_n537, u4_srl_451_n536, u4_srl_451_n535,
         u4_srl_451_n534, u4_srl_451_n533, u4_srl_451_n532, u4_srl_451_n531,
         u4_srl_451_n530, u4_srl_451_n529, u4_srl_451_n528, u4_srl_451_n527,
         u4_srl_451_n526, u4_srl_451_n525, u4_srl_451_n524, u4_srl_451_n523,
         u4_srl_451_n522, u4_srl_451_n521, u4_srl_451_n520, u4_srl_451_n519,
         u4_srl_451_n518, u4_srl_451_n517, u4_srl_451_n516, u4_srl_451_n515,
         u4_srl_451_n514, u4_srl_451_n513, u4_srl_451_n512, u4_srl_451_n511,
         u4_srl_451_n510, u4_srl_451_n509, u4_srl_451_n508, u4_srl_451_n507,
         u4_srl_451_n506, u4_srl_451_n505, u4_srl_451_n504, u4_srl_451_n503,
         u4_srl_451_n502, u4_srl_451_n501, u4_srl_451_n500, u4_srl_451_n499,
         u4_srl_451_n498, u4_srl_451_n497, u4_srl_451_n496, u4_srl_451_n495,
         u4_srl_451_n494, u4_srl_451_n493, u4_srl_451_n492, u4_srl_451_n491,
         u4_srl_451_n490, u4_srl_451_n489, u4_srl_451_n488, u4_srl_451_n487,
         u4_srl_451_n486, u4_srl_451_n485, u4_srl_451_n484, u4_srl_451_n483,
         u4_srl_451_n482, u4_srl_451_n481, u4_srl_451_n480, u4_srl_451_n479,
         u4_srl_451_n478, u4_srl_451_n477, u4_srl_451_n476, u4_srl_451_n475,
         u4_srl_451_n474, u4_srl_451_n473, u4_srl_451_n472, u4_srl_451_n471,
         u4_srl_451_n470, u4_srl_451_n469, u4_srl_451_n468, u4_srl_451_n467,
         u4_srl_451_n466, u4_srl_451_n465, u4_srl_451_n464, u4_srl_451_n463,
         u4_srl_451_n462, u4_srl_451_n461, u4_srl_451_n460, u4_srl_451_n459,
         u4_srl_451_n458, u4_srl_451_n457, u4_srl_451_n456, u4_srl_451_n455,
         u4_srl_451_n454, u4_srl_451_n453, u4_srl_451_n452, u4_srl_451_n451,
         u4_srl_451_n450, u4_srl_451_n449, u4_srl_451_n448, u4_srl_451_n447,
         u4_srl_451_n446, u4_srl_451_n445, u4_srl_451_n444, u4_srl_451_n443,
         u4_srl_451_n442, u4_srl_451_n441, u4_srl_451_n440, u4_srl_451_n439,
         u4_srl_451_n438, u4_srl_451_n437, u4_srl_451_n436, u4_srl_451_n435,
         u4_srl_451_n434, u4_srl_451_n433, u4_srl_451_n432, u4_srl_451_n431,
         u4_srl_451_n430, u4_srl_451_n429, u4_srl_451_n428, u4_srl_451_n427,
         u4_srl_451_n426, u4_srl_451_n425, u4_srl_451_n424, u4_srl_451_n423,
         u4_srl_451_n422, u4_srl_451_n421, u4_srl_451_n420, u4_srl_451_n419,
         u4_srl_451_n418, u4_srl_451_n417, u4_srl_451_n416, u4_srl_451_n415,
         u4_srl_451_n414, u4_srl_451_n413, u4_srl_451_n412, u4_srl_451_n411,
         u4_srl_451_n410, u4_srl_451_n409, u4_srl_451_n408, u4_srl_451_n407,
         u4_srl_451_n406, u4_srl_451_n405, u4_srl_451_n404, u4_srl_451_n403,
         u4_srl_451_n402, u4_srl_451_n401, u4_srl_451_n400, u4_srl_451_n399,
         u4_srl_451_n398, u4_srl_451_n397, u4_srl_451_n396, u4_srl_451_n395,
         u4_srl_451_n394, u4_srl_451_n393, u4_srl_451_n392, u4_srl_451_n391,
         u4_srl_451_n390, u4_srl_451_n389, u4_srl_451_n388, u4_srl_451_n387,
         u4_srl_451_n386, u4_srl_451_n385, u4_srl_451_n384, u4_srl_451_n383,
         u4_srl_451_n382, u4_srl_451_n381, u4_srl_451_n380, u4_srl_451_n379,
         u4_srl_451_n378, u4_srl_451_n377, u4_srl_451_n376, u4_srl_451_n375,
         u4_srl_451_n374, u4_srl_451_n373, u4_srl_451_n372, u4_srl_451_n371,
         u4_srl_451_n370, u4_srl_451_n369, u4_srl_451_n368, u4_srl_451_n367,
         u4_srl_451_n366, u4_srl_451_n365, u4_srl_451_n364, u4_srl_451_n363,
         u4_srl_451_n362, u4_srl_451_n361, u4_srl_451_n360, u4_srl_451_n359,
         u4_srl_451_n358, u4_srl_451_n357, u4_srl_451_n356, u4_srl_451_n355,
         u4_srl_451_n354, u4_srl_451_n353, u4_srl_451_n352, u4_srl_451_n351,
         u4_srl_451_n350, u4_srl_451_n349, u4_srl_451_n348, u4_srl_451_n347,
         u4_srl_451_n346, u4_srl_451_n345, u4_srl_451_n344, u4_srl_451_n343,
         u4_srl_451_n342, u4_srl_451_n341, u4_srl_451_n340, u4_srl_451_n339,
         u4_srl_451_n338, u4_srl_451_n337, u4_srl_451_n336, u4_srl_451_n335,
         u4_srl_451_n334, u4_srl_451_n333, u4_srl_451_n332, u4_srl_451_n331,
         u4_srl_451_n330, u4_srl_451_n329, u4_srl_451_n328, u4_srl_451_n327,
         u4_srl_451_n326, u4_srl_451_n325, u4_srl_451_n324, u4_srl_451_n323,
         u4_srl_451_n322, u4_srl_451_n321, u4_srl_451_n320, u4_srl_451_n319,
         u4_srl_451_n318, u4_srl_451_n317, u4_srl_451_n316, u4_srl_451_n315,
         u4_srl_451_n314, u4_srl_451_n313, u4_srl_451_n312, u4_srl_451_n311,
         u4_srl_451_n310, u4_srl_451_n309, u4_srl_451_n308, u4_srl_451_n307,
         u4_srl_451_n306, u4_srl_451_n305, u4_srl_451_n304, u4_srl_451_n303,
         u4_srl_451_n302, u4_srl_451_n301, u4_srl_451_n300, u4_srl_451_n299,
         u4_srl_451_n298, u4_srl_451_n297, u4_srl_451_n296, u4_srl_451_n295,
         u4_srl_451_n294, u4_srl_451_n293, u4_srl_451_n292, u4_srl_451_n291,
         u4_srl_451_n290, u4_srl_451_n289, u4_srl_451_n288, u4_srl_451_n287,
         u4_srl_451_n286, u4_srl_451_n285, u4_srl_451_n284, u4_srl_451_n283,
         u4_srl_451_n282, u4_srl_451_n281, u4_srl_451_n280, u4_srl_451_n279,
         u4_srl_451_n278, u4_srl_451_n277, u4_srl_451_n276, u4_srl_451_n275,
         u4_srl_451_n274, u4_srl_451_n273, u4_srl_451_n272, u4_srl_451_n271,
         u4_srl_451_n270, u4_srl_451_n269, u4_srl_451_n268, u4_srl_451_n267,
         u4_srl_451_n266, u4_srl_451_n265, u4_srl_451_n264, u4_srl_451_n263,
         u4_srl_451_n262, u4_srl_451_n261, u4_srl_451_n260, u4_srl_451_n259,
         u4_srl_451_n258, u4_srl_451_n257, u4_srl_451_n256, u4_srl_451_n255,
         u4_srl_451_n254, u4_srl_451_n253, u4_srl_451_n252, u4_srl_451_n251,
         u4_srl_451_n250, u4_srl_451_n249, u4_srl_451_n248, u4_srl_451_n247,
         u4_srl_451_n246, u4_srl_451_n245, u4_srl_451_n244, u4_srl_451_n243,
         u4_srl_451_n242, u4_srl_451_n241, u4_srl_451_n240, u4_srl_451_n239,
         u4_srl_451_n238, u4_srl_451_n237, u4_srl_451_n236, u4_srl_451_n235,
         u4_srl_451_n234, u4_srl_451_n233, u4_srl_451_n232, u4_srl_451_n231,
         u4_srl_451_n230, u4_srl_451_n229, u4_srl_451_n228, u4_srl_451_n227,
         u4_srl_451_n226, u4_srl_451_n225, u4_srl_451_n224, u4_srl_451_n223,
         u4_srl_451_n222, u4_srl_451_n221, u4_srl_451_n220, u4_srl_451_n219,
         u4_srl_451_n218, u4_srl_451_n217, u4_srl_451_n216, u4_srl_451_n215,
         u4_srl_451_n214, u4_srl_451_n213, u4_srl_451_n212, u4_srl_451_n211,
         u4_srl_451_n210, u4_srl_451_n209, u4_srl_451_n208, u4_srl_451_n207,
         u4_srl_451_n206, u4_srl_451_n205, u4_srl_451_n204, u4_srl_451_n203,
         u4_srl_451_n202, u4_srl_451_n201, u4_srl_451_n200, u4_srl_451_n199,
         u4_srl_451_n198, u4_srl_451_n197, u4_srl_451_n196, u4_srl_451_n195,
         u4_srl_451_n194, u4_srl_451_n193, u4_srl_451_n192, u4_srl_451_n191,
         u4_srl_451_n190, u4_srl_451_n189, u4_srl_451_n188, u4_srl_451_n187,
         u4_srl_451_n186, u4_srl_451_n185, u4_srl_451_n184, u4_srl_451_n183,
         u4_srl_451_n182, u4_srl_451_n181, u4_srl_451_n180, u4_srl_451_n179,
         u4_srl_451_n178, u4_srl_451_n177, u4_srl_451_n176, u4_srl_451_n175,
         u4_srl_451_n174, u4_srl_451_n173, u4_srl_451_n172, u4_srl_451_n171,
         u4_srl_451_n170, u4_srl_451_n169, u4_srl_451_n168, u4_srl_451_n167,
         u4_srl_451_n166, u4_srl_451_n165, u4_srl_451_n164, u4_srl_451_n163,
         u4_srl_451_n162, u4_srl_451_n161, u4_srl_451_n160, u4_srl_451_n159,
         u4_srl_451_n158, u4_srl_451_n157, u4_srl_451_n156, u4_srl_451_n155,
         u4_srl_451_n154, u4_srl_451_n153, u4_srl_451_n152, u4_srl_451_n151,
         u4_srl_451_n150, u4_srl_451_n149, u4_srl_451_n148, u4_srl_451_n147,
         u4_srl_451_n146, u4_srl_451_n145, u4_srl_451_n144, u4_srl_451_n143,
         u4_srl_451_n142, u4_srl_451_n141, u4_srl_451_n140, u4_srl_451_n139,
         u4_srl_451_n138, u4_srl_451_n137, u4_srl_451_n136, u4_srl_451_n135,
         u4_srl_451_n134, u4_srl_451_n133, u4_srl_451_n132, u4_srl_451_n131,
         u4_srl_451_n130, u4_srl_451_n129, u4_srl_451_n128, u4_srl_451_n127,
         u4_srl_451_n126, u4_srl_451_n125, u4_srl_451_n124, u4_srl_451_n123,
         u4_srl_451_n122, u4_srl_451_n121, u4_srl_451_n120, u4_srl_451_n119,
         u4_srl_451_n118, u4_srl_451_n117, u4_srl_451_n116, u4_srl_451_n115,
         u4_srl_451_n114, u4_srl_451_n113, u4_srl_451_n112, u4_srl_451_n111,
         u4_srl_451_n110, u4_srl_451_n109, u4_srl_451_n108, u4_srl_451_n107,
         u4_srl_451_n106, u4_srl_451_n105, u4_srl_451_n104, u4_srl_451_n103,
         u4_srl_451_n102, u4_srl_451_n101, u4_srl_451_n100, u4_srl_451_n99,
         u4_srl_451_n98, u4_srl_451_n97, u4_srl_451_n96, u4_srl_451_n95,
         u4_srl_451_n94, u4_srl_451_n93, u4_srl_451_n92, u4_srl_451_n91,
         u4_srl_451_n90, u4_srl_451_n89, u4_srl_451_n88, u4_srl_451_n87,
         u4_srl_451_n86, u4_srl_451_n85, u4_srl_451_n84, u4_srl_451_n83,
         u4_srl_451_n82, u4_srl_451_n81, u4_srl_451_n80, u4_srl_451_n79,
         u4_srl_451_n78, u4_srl_451_n77, u4_srl_451_n76, u4_srl_451_n75,
         u4_srl_451_n74, u4_srl_451_n73, u4_srl_451_n72, u4_srl_451_n71,
         u4_srl_451_n70, u4_srl_451_n69, u4_srl_451_n68, u4_srl_451_n67,
         u4_srl_451_n66, u4_srl_451_n65, u4_srl_451_n64, u4_srl_451_n63,
         u4_srl_451_n62, u4_srl_451_n61, u4_srl_451_n60, u4_srl_451_n59,
         u4_srl_451_n58, u4_srl_451_n57, u4_srl_451_n56, u4_srl_451_n55,
         u4_srl_451_n54, u4_srl_451_n53, u4_srl_451_n52, u4_srl_451_n51,
         u4_srl_451_n50, u4_srl_451_n49, u4_srl_451_n48, u4_srl_451_n47,
         u4_srl_451_n46, u4_srl_451_n45, u4_srl_451_n44, u4_srl_451_n43,
         u4_srl_451_n42, u4_srl_451_n41, u4_srl_451_n40, u4_srl_451_n39,
         u4_srl_451_n38, u4_srl_451_n37, u4_srl_451_n36, u4_srl_451_n35,
         u4_srl_451_n34, u4_srl_451_n33, u4_srl_451_n32, u4_srl_451_n31,
         u4_srl_451_n30, u4_srl_451_n29, u4_srl_451_n28, u4_srl_451_n27,
         u4_srl_451_n26, u4_srl_451_n25, u4_srl_451_n24, u4_srl_451_n23,
         u4_srl_451_n22, u4_srl_451_n21, u4_srl_451_n20, u4_srl_451_n19,
         u4_srl_451_n18, u4_srl_451_n17, u4_srl_451_n16, u4_srl_451_n15,
         u4_srl_451_n14, u4_srl_451_n13, u4_srl_451_n12, u4_srl_451_n11,
         u4_srl_451_n10, u4_srl_451_n9, u4_srl_451_n8, u4_srl_451_n7,
         u4_srl_451_n6, u4_srl_451_n5, u4_srl_451_n4, u4_srl_451_n3,
         u4_srl_451_n2, u4_srl_451_n1, u4_sll_480_n58, u4_sll_480_n57,
         u4_sll_480_n56, u4_sll_480_n55, u4_sll_480_n54, u4_sll_480_n53,
         u4_sll_480_n52, u4_sll_480_n51, u4_sll_480_n50, u4_sll_480_n49,
         u4_sll_480_n48, u4_sll_480_n47, u4_sll_480_n46, u4_sll_480_n45,
         u4_sll_480_n44, u4_sll_480_n43, u4_sll_480_n42, u4_sll_480_n41,
         u4_sll_480_n40, u4_sll_480_n39, u4_sll_480_n38, u4_sll_480_n37,
         u4_sll_480_n36, u4_sll_480_n35, u4_sll_480_n34, u4_sll_480_n33,
         u4_sll_480_n32, u4_sll_480_n31, u4_sll_480_n30, u4_sll_480_n29,
         u4_sll_480_n28, u4_sll_480_n27, u4_sll_480_n26, u4_sll_480_n25,
         u4_sll_480_n24, u4_sll_480_n23, u4_sll_480_n22, u4_sll_480_n21,
         u4_sll_480_n20, u4_sll_480_n19, u4_sll_480_n18, u4_sll_480_n17,
         u4_sll_480_n16, u4_sll_480_n15, u4_sll_480_n14, u4_sll_480_n13,
         u4_sll_480_n12, u4_sll_480_n11, u4_sll_480_n10, u4_sll_480_n9,
         u4_sll_480_n8, u4_sll_480_n7, u4_sll_480_n6, u4_sll_480_n5,
         u4_sll_480_n4, u4_sll_480_n3, u4_sll_480_n2, u4_sll_480_n1,
         u4_sll_480_ML_int_7__107_, u4_sll_480_ML_int_7__108_,
         u4_sll_480_ML_int_7__109_, u4_sll_480_ML_int_7__110_,
         u4_sll_480_ML_int_7__111_, u4_sll_480_ML_int_7__112_,
         u4_sll_480_ML_int_7__113_, u4_sll_480_ML_int_7__114_,
         u4_sll_480_ML_int_7__115_, u4_sll_480_ML_int_7__116_,
         u4_sll_480_ML_int_7__117_, u4_sll_480_ML_int_6__43_,
         u4_sll_480_ML_int_6__44_, u4_sll_480_ML_int_6__45_,
         u4_sll_480_ML_int_6__46_, u4_sll_480_ML_int_6__47_,
         u4_sll_480_ML_int_6__48_, u4_sll_480_ML_int_6__49_,
         u4_sll_480_ML_int_6__50_, u4_sll_480_ML_int_6__51_,
         u4_sll_480_ML_int_6__52_, u4_sll_480_ML_int_6__53_,
         u4_sll_480_ML_int_6__107_, u4_sll_480_ML_int_6__108_,
         u4_sll_480_ML_int_6__109_, u4_sll_480_ML_int_6__110_,
         u4_sll_480_ML_int_6__111_, u4_sll_480_ML_int_6__112_,
         u4_sll_480_ML_int_6__113_, u4_sll_480_ML_int_6__114_,
         u4_sll_480_ML_int_6__115_, u4_sll_480_ML_int_6__116_,
         u4_sll_480_ML_int_6__117_, u4_sll_480_ML_int_5__11_,
         u4_sll_480_ML_int_5__12_, u4_sll_480_ML_int_5__13_,
         u4_sll_480_ML_int_5__14_, u4_sll_480_ML_int_5__15_,
         u4_sll_480_ML_int_5__16_, u4_sll_480_ML_int_5__17_,
         u4_sll_480_ML_int_5__18_, u4_sll_480_ML_int_5__19_,
         u4_sll_480_ML_int_5__20_, u4_sll_480_ML_int_5__21_,
         u4_sll_480_ML_int_5__43_, u4_sll_480_ML_int_5__44_,
         u4_sll_480_ML_int_5__45_, u4_sll_480_ML_int_5__46_,
         u4_sll_480_ML_int_5__47_, u4_sll_480_ML_int_5__48_,
         u4_sll_480_ML_int_5__49_, u4_sll_480_ML_int_5__50_,
         u4_sll_480_ML_int_5__51_, u4_sll_480_ML_int_5__52_,
         u4_sll_480_ML_int_5__53_, u4_sll_480_ML_int_5__75_,
         u4_sll_480_ML_int_5__76_, u4_sll_480_ML_int_5__77_,
         u4_sll_480_ML_int_5__78_, u4_sll_480_ML_int_5__79_,
         u4_sll_480_ML_int_5__80_, u4_sll_480_ML_int_5__81_,
         u4_sll_480_ML_int_5__82_, u4_sll_480_ML_int_5__83_,
         u4_sll_480_ML_int_5__84_, u4_sll_480_ML_int_5__85_,
         u4_sll_480_ML_int_5__107_, u4_sll_480_ML_int_5__108_,
         u4_sll_480_ML_int_5__109_, u4_sll_480_ML_int_5__110_,
         u4_sll_480_ML_int_5__111_, u4_sll_480_ML_int_5__112_,
         u4_sll_480_ML_int_5__113_, u4_sll_480_ML_int_5__114_,
         u4_sll_480_ML_int_5__115_, u4_sll_480_ML_int_5__116_,
         u4_sll_480_ML_int_5__117_, u4_sll_480_ML_int_4__0_,
         u4_sll_480_ML_int_4__1_, u4_sll_480_ML_int_4__2_,
         u4_sll_480_ML_int_4__3_, u4_sll_480_ML_int_4__4_,
         u4_sll_480_ML_int_4__5_, u4_sll_480_ML_int_4__11_,
         u4_sll_480_ML_int_4__12_, u4_sll_480_ML_int_4__13_,
         u4_sll_480_ML_int_4__14_, u4_sll_480_ML_int_4__15_,
         u4_sll_480_ML_int_4__16_, u4_sll_480_ML_int_4__17_,
         u4_sll_480_ML_int_4__18_, u4_sll_480_ML_int_4__19_,
         u4_sll_480_ML_int_4__20_, u4_sll_480_ML_int_4__21_,
         u4_sll_480_ML_int_4__27_, u4_sll_480_ML_int_4__28_,
         u4_sll_480_ML_int_4__29_, u4_sll_480_ML_int_4__30_,
         u4_sll_480_ML_int_4__31_, u4_sll_480_ML_int_4__32_,
         u4_sll_480_ML_int_4__33_, u4_sll_480_ML_int_4__34_,
         u4_sll_480_ML_int_4__35_, u4_sll_480_ML_int_4__36_,
         u4_sll_480_ML_int_4__37_, u4_sll_480_ML_int_4__43_,
         u4_sll_480_ML_int_4__44_, u4_sll_480_ML_int_4__45_,
         u4_sll_480_ML_int_4__46_, u4_sll_480_ML_int_4__47_,
         u4_sll_480_ML_int_4__48_, u4_sll_480_ML_int_4__49_,
         u4_sll_480_ML_int_4__50_, u4_sll_480_ML_int_4__51_,
         u4_sll_480_ML_int_4__52_, u4_sll_480_ML_int_4__53_,
         u4_sll_480_ML_int_4__59_, u4_sll_480_ML_int_4__60_,
         u4_sll_480_ML_int_4__61_, u4_sll_480_ML_int_4__62_,
         u4_sll_480_ML_int_4__63_, u4_sll_480_ML_int_4__64_,
         u4_sll_480_ML_int_4__65_, u4_sll_480_ML_int_4__66_,
         u4_sll_480_ML_int_4__67_, u4_sll_480_ML_int_4__68_,
         u4_sll_480_ML_int_4__69_, u4_sll_480_ML_int_4__75_,
         u4_sll_480_ML_int_4__76_, u4_sll_480_ML_int_4__77_,
         u4_sll_480_ML_int_4__78_, u4_sll_480_ML_int_4__79_,
         u4_sll_480_ML_int_4__80_, u4_sll_480_ML_int_4__81_,
         u4_sll_480_ML_int_4__82_, u4_sll_480_ML_int_4__83_,
         u4_sll_480_ML_int_4__84_, u4_sll_480_ML_int_4__85_,
         u4_sll_480_ML_int_4__91_, u4_sll_480_ML_int_4__92_,
         u4_sll_480_ML_int_4__93_, u4_sll_480_ML_int_4__94_,
         u4_sll_480_ML_int_4__95_, u4_sll_480_ML_int_4__96_,
         u4_sll_480_ML_int_4__97_, u4_sll_480_ML_int_4__98_,
         u4_sll_480_ML_int_4__99_, u4_sll_480_ML_int_4__100_,
         u4_sll_480_ML_int_4__101_, u4_sll_480_ML_int_4__107_,
         u4_sll_480_ML_int_4__108_, u4_sll_480_ML_int_4__109_,
         u4_sll_480_ML_int_4__110_, u4_sll_480_ML_int_4__111_,
         u4_sll_480_ML_int_4__112_, u4_sll_480_ML_int_4__113_,
         u4_sll_480_ML_int_4__114_, u4_sll_480_ML_int_4__115_,
         u4_sll_480_ML_int_4__116_, u4_sll_480_ML_int_4__117_,
         u4_sll_480_ML_int_3__4_, u4_sll_480_ML_int_3__5_,
         u4_sll_480_ML_int_3__6_, u4_sll_480_ML_int_3__7_,
         u4_sll_480_ML_int_3__8_, u4_sll_480_ML_int_3__9_,
         u4_sll_480_ML_int_3__10_, u4_sll_480_ML_int_3__11_,
         u4_sll_480_ML_int_3__12_, u4_sll_480_ML_int_3__13_,
         u4_sll_480_ML_int_3__14_, u4_sll_480_ML_int_3__15_,
         u4_sll_480_ML_int_3__16_, u4_sll_480_ML_int_3__17_,
         u4_sll_480_ML_int_3__18_, u4_sll_480_ML_int_3__19_,
         u4_sll_480_ML_int_3__20_, u4_sll_480_ML_int_3__21_,
         u4_sll_480_ML_int_3__22_, u4_sll_480_ML_int_3__23_,
         u4_sll_480_ML_int_3__24_, u4_sll_480_ML_int_3__25_,
         u4_sll_480_ML_int_3__26_, u4_sll_480_ML_int_3__27_,
         u4_sll_480_ML_int_3__28_, u4_sll_480_ML_int_3__29_,
         u4_sll_480_ML_int_3__30_, u4_sll_480_ML_int_3__31_,
         u4_sll_480_ML_int_3__32_, u4_sll_480_ML_int_3__33_,
         u4_sll_480_ML_int_3__34_, u4_sll_480_ML_int_3__35_,
         u4_sll_480_ML_int_3__36_, u4_sll_480_ML_int_3__37_,
         u4_sll_480_ML_int_3__38_, u4_sll_480_ML_int_3__39_,
         u4_sll_480_ML_int_3__40_, u4_sll_480_ML_int_3__41_,
         u4_sll_480_ML_int_3__42_, u4_sll_480_ML_int_3__43_,
         u4_sll_480_ML_int_3__44_, u4_sll_480_ML_int_3__45_,
         u4_sll_480_ML_int_3__46_, u4_sll_480_ML_int_3__47_,
         u4_sll_480_ML_int_3__48_, u4_sll_480_ML_int_3__49_,
         u4_sll_480_ML_int_3__50_, u4_sll_480_ML_int_3__51_,
         u4_sll_480_ML_int_3__52_, u4_sll_480_ML_int_3__53_,
         u4_sll_480_ML_int_3__54_, u4_sll_480_ML_int_3__55_,
         u4_sll_480_ML_int_3__56_, u4_sll_480_ML_int_3__57_,
         u4_sll_480_ML_int_3__58_, u4_sll_480_ML_int_3__59_,
         u4_sll_480_ML_int_3__60_, u4_sll_480_ML_int_3__61_,
         u4_sll_480_ML_int_3__62_, u4_sll_480_ML_int_3__63_,
         u4_sll_480_ML_int_3__64_, u4_sll_480_ML_int_3__65_,
         u4_sll_480_ML_int_3__66_, u4_sll_480_ML_int_3__67_,
         u4_sll_480_ML_int_3__68_, u4_sll_480_ML_int_3__69_,
         u4_sll_480_ML_int_3__70_, u4_sll_480_ML_int_3__71_,
         u4_sll_480_ML_int_3__72_, u4_sll_480_ML_int_3__73_,
         u4_sll_480_ML_int_3__74_, u4_sll_480_ML_int_3__75_,
         u4_sll_480_ML_int_3__76_, u4_sll_480_ML_int_3__77_,
         u4_sll_480_ML_int_3__78_, u4_sll_480_ML_int_3__79_,
         u4_sll_480_ML_int_3__80_, u4_sll_480_ML_int_3__81_,
         u4_sll_480_ML_int_3__82_, u4_sll_480_ML_int_3__83_,
         u4_sll_480_ML_int_3__84_, u4_sll_480_ML_int_3__85_,
         u4_sll_480_ML_int_3__86_, u4_sll_480_ML_int_3__87_,
         u4_sll_480_ML_int_3__88_, u4_sll_480_ML_int_3__89_,
         u4_sll_480_ML_int_3__90_, u4_sll_480_ML_int_3__91_,
         u4_sll_480_ML_int_3__92_, u4_sll_480_ML_int_3__93_,
         u4_sll_480_ML_int_3__94_, u4_sll_480_ML_int_3__95_,
         u4_sll_480_ML_int_3__96_, u4_sll_480_ML_int_3__97_,
         u4_sll_480_ML_int_3__98_, u4_sll_480_ML_int_3__99_,
         u4_sll_480_ML_int_3__100_, u4_sll_480_ML_int_3__101_,
         u4_sll_480_ML_int_3__102_, u4_sll_480_ML_int_3__103_,
         u4_sll_480_ML_int_3__104_, u4_sll_480_ML_int_3__105_,
         u4_sll_480_ML_int_3__106_, u4_sll_480_ML_int_3__107_,
         u4_sll_480_ML_int_3__108_, u4_sll_480_ML_int_3__109_,
         u4_sll_480_ML_int_3__110_, u4_sll_480_ML_int_3__111_,
         u4_sll_480_ML_int_3__112_, u4_sll_480_ML_int_3__113_,
         u4_sll_480_ML_int_3__114_, u4_sll_480_ML_int_3__115_,
         u4_sll_480_ML_int_3__116_, u4_sll_480_ML_int_2__2_,
         u4_sll_480_ML_int_2__3_, u4_sll_480_ML_int_2__4_,
         u4_sll_480_ML_int_2__5_, u4_sll_480_ML_int_2__6_,
         u4_sll_480_ML_int_2__7_, u4_sll_480_ML_int_2__8_,
         u4_sll_480_ML_int_2__9_, u4_sll_480_ML_int_2__10_,
         u4_sll_480_ML_int_2__11_, u4_sll_480_ML_int_2__12_,
         u4_sll_480_ML_int_2__13_, u4_sll_480_ML_int_2__14_,
         u4_sll_480_ML_int_2__15_, u4_sll_480_ML_int_2__16_,
         u4_sll_480_ML_int_2__17_, u4_sll_480_ML_int_2__18_,
         u4_sll_480_ML_int_2__19_, u4_sll_480_ML_int_2__20_,
         u4_sll_480_ML_int_2__21_, u4_sll_480_ML_int_2__22_,
         u4_sll_480_ML_int_2__23_, u4_sll_480_ML_int_2__24_,
         u4_sll_480_ML_int_2__25_, u4_sll_480_ML_int_2__26_,
         u4_sll_480_ML_int_2__27_, u4_sll_480_ML_int_2__28_,
         u4_sll_480_ML_int_2__29_, u4_sll_480_ML_int_2__30_,
         u4_sll_480_ML_int_2__31_, u4_sll_480_ML_int_2__32_,
         u4_sll_480_ML_int_2__33_, u4_sll_480_ML_int_2__34_,
         u4_sll_480_ML_int_2__35_, u4_sll_480_ML_int_2__36_,
         u4_sll_480_ML_int_2__37_, u4_sll_480_ML_int_2__38_,
         u4_sll_480_ML_int_2__39_, u4_sll_480_ML_int_2__40_,
         u4_sll_480_ML_int_2__41_, u4_sll_480_ML_int_2__42_,
         u4_sll_480_ML_int_2__43_, u4_sll_480_ML_int_2__44_,
         u4_sll_480_ML_int_2__45_, u4_sll_480_ML_int_2__46_,
         u4_sll_480_ML_int_2__47_, u4_sll_480_ML_int_2__48_,
         u4_sll_480_ML_int_2__49_, u4_sll_480_ML_int_2__50_,
         u4_sll_480_ML_int_2__51_, u4_sll_480_ML_int_2__52_,
         u4_sll_480_ML_int_2__53_, u4_sll_480_ML_int_2__54_,
         u4_sll_480_ML_int_2__55_, u4_sll_480_ML_int_2__56_,
         u4_sll_480_ML_int_2__57_, u4_sll_480_ML_int_2__58_,
         u4_sll_480_ML_int_2__59_, u4_sll_480_ML_int_2__60_,
         u4_sll_480_ML_int_2__61_, u4_sll_480_ML_int_2__62_,
         u4_sll_480_ML_int_2__63_, u4_sll_480_ML_int_2__64_,
         u4_sll_480_ML_int_2__65_, u4_sll_480_ML_int_2__66_,
         u4_sll_480_ML_int_2__67_, u4_sll_480_ML_int_2__68_,
         u4_sll_480_ML_int_2__69_, u4_sll_480_ML_int_2__70_,
         u4_sll_480_ML_int_2__71_, u4_sll_480_ML_int_2__72_,
         u4_sll_480_ML_int_2__73_, u4_sll_480_ML_int_2__74_,
         u4_sll_480_ML_int_2__75_, u4_sll_480_ML_int_2__76_,
         u4_sll_480_ML_int_2__77_, u4_sll_480_ML_int_2__78_,
         u4_sll_480_ML_int_2__79_, u4_sll_480_ML_int_2__80_,
         u4_sll_480_ML_int_2__81_, u4_sll_480_ML_int_2__82_,
         u4_sll_480_ML_int_2__83_, u4_sll_480_ML_int_2__84_,
         u4_sll_480_ML_int_2__85_, u4_sll_480_ML_int_2__86_,
         u4_sll_480_ML_int_2__87_, u4_sll_480_ML_int_2__88_,
         u4_sll_480_ML_int_2__89_, u4_sll_480_ML_int_2__90_,
         u4_sll_480_ML_int_2__91_, u4_sll_480_ML_int_2__92_,
         u4_sll_480_ML_int_2__93_, u4_sll_480_ML_int_2__94_,
         u4_sll_480_ML_int_2__95_, u4_sll_480_ML_int_2__96_,
         u4_sll_480_ML_int_2__97_, u4_sll_480_ML_int_2__98_,
         u4_sll_480_ML_int_2__99_, u4_sll_480_ML_int_2__100_,
         u4_sll_480_ML_int_2__101_, u4_sll_480_ML_int_2__102_,
         u4_sll_480_ML_int_2__103_, u4_sll_480_ML_int_2__104_,
         u4_sll_480_ML_int_2__105_, u4_sll_480_ML_int_2__106_,
         u4_sll_480_ML_int_2__107_, u4_sll_480_ML_int_2__108_,
         u4_sll_480_ML_int_2__109_, u4_sll_480_ML_int_2__110_,
         u4_sll_480_ML_int_2__111_, u4_sll_480_ML_int_2__112_,
         u4_sll_480_ML_int_2__113_, u4_sll_480_ML_int_2__114_,
         u4_sll_480_ML_int_1__0_, u4_sll_480_ML_int_1__1_,
         u4_sll_480_ML_int_1__2_, u4_sll_480_ML_int_1__3_,
         u4_sll_480_ML_int_1__4_, u4_sll_480_ML_int_1__5_,
         u4_sll_480_ML_int_1__6_, u4_sll_480_ML_int_1__7_,
         u4_sll_480_ML_int_1__8_, u4_sll_480_ML_int_1__9_,
         u4_sll_480_ML_int_1__10_, u4_sll_480_ML_int_1__11_,
         u4_sll_480_ML_int_1__12_, u4_sll_480_ML_int_1__13_,
         u4_sll_480_ML_int_1__14_, u4_sll_480_ML_int_1__15_,
         u4_sll_480_ML_int_1__16_, u4_sll_480_ML_int_1__17_,
         u4_sll_480_ML_int_1__18_, u4_sll_480_ML_int_1__19_,
         u4_sll_480_ML_int_1__20_, u4_sll_480_ML_int_1__21_,
         u4_sll_480_ML_int_1__22_, u4_sll_480_ML_int_1__23_,
         u4_sll_480_ML_int_1__24_, u4_sll_480_ML_int_1__25_,
         u4_sll_480_ML_int_1__26_, u4_sll_480_ML_int_1__27_,
         u4_sll_480_ML_int_1__28_, u4_sll_480_ML_int_1__29_,
         u4_sll_480_ML_int_1__30_, u4_sll_480_ML_int_1__31_,
         u4_sll_480_ML_int_1__32_, u4_sll_480_ML_int_1__33_,
         u4_sll_480_ML_int_1__34_, u4_sll_480_ML_int_1__35_,
         u4_sll_480_ML_int_1__36_, u4_sll_480_ML_int_1__37_,
         u4_sll_480_ML_int_1__38_, u4_sll_480_ML_int_1__39_,
         u4_sll_480_ML_int_1__40_, u4_sll_480_ML_int_1__41_,
         u4_sll_480_ML_int_1__42_, u4_sll_480_ML_int_1__43_,
         u4_sll_480_ML_int_1__44_, u4_sll_480_ML_int_1__45_,
         u4_sll_480_ML_int_1__46_, u4_sll_480_ML_int_1__47_,
         u4_sll_480_ML_int_1__48_, u4_sll_480_ML_int_1__49_,
         u4_sll_480_ML_int_1__50_, u4_sll_480_ML_int_1__51_,
         u4_sll_480_ML_int_1__52_, u4_sll_480_ML_int_1__53_,
         u4_sll_480_ML_int_1__54_, u4_sll_480_ML_int_1__55_,
         u4_sll_480_ML_int_1__56_, u4_sll_480_ML_int_1__57_,
         u4_sll_480_ML_int_1__58_, u4_sll_480_ML_int_1__59_,
         u4_sll_480_ML_int_1__60_, u4_sll_480_ML_int_1__61_,
         u4_sll_480_ML_int_1__62_, u4_sll_480_ML_int_1__63_,
         u4_sll_480_ML_int_1__64_, u4_sll_480_ML_int_1__65_,
         u4_sll_480_ML_int_1__66_, u4_sll_480_ML_int_1__67_,
         u4_sll_480_ML_int_1__68_, u4_sll_480_ML_int_1__69_,
         u4_sll_480_ML_int_1__70_, u4_sll_480_ML_int_1__71_,
         u4_sll_480_ML_int_1__72_, u4_sll_480_ML_int_1__73_,
         u4_sll_480_ML_int_1__74_, u4_sll_480_ML_int_1__75_,
         u4_sll_480_ML_int_1__76_, u4_sll_480_ML_int_1__77_,
         u4_sll_480_ML_int_1__78_, u4_sll_480_ML_int_1__79_,
         u4_sll_480_ML_int_1__80_, u4_sll_480_ML_int_1__81_,
         u4_sll_480_ML_int_1__82_, u4_sll_480_ML_int_1__83_,
         u4_sll_480_ML_int_1__84_, u4_sll_480_ML_int_1__85_,
         u4_sll_480_ML_int_1__86_, u4_sll_480_ML_int_1__87_,
         u4_sll_480_ML_int_1__88_, u4_sll_480_ML_int_1__89_,
         u4_sll_480_ML_int_1__90_, u4_sll_480_ML_int_1__91_,
         u4_sll_480_ML_int_1__92_, u4_sll_480_ML_int_1__93_,
         u4_sll_480_ML_int_1__94_, u4_sll_480_ML_int_1__95_,
         u4_sll_480_ML_int_1__96_, u4_sll_480_ML_int_1__97_,
         u4_sll_480_ML_int_1__98_, u4_sll_480_ML_int_1__99_,
         u4_sll_480_ML_int_1__100_, u4_sll_480_ML_int_1__101_,
         u4_sll_480_ML_int_1__102_, u4_sll_480_ML_int_1__103_,
         u4_sll_480_ML_int_1__104_, u4_sll_480_ML_int_1__105_,
         u4_sll_480_ML_int_1__106_, u4_sll_480_ML_int_1__107_,
         u4_sll_480_ML_int_1__108_, u4_sll_480_ML_int_1__109_,
         u4_sll_480_ML_int_1__110_, u4_sll_480_ML_int_1__111_,
         u4_sll_480_ML_int_1__112_, u4_sll_480_ML_int_1__113_,
         u4_sll_480_MR_int_1__113_, u4_sll_480_temp_int_SH_0_,
         u4_sll_480_temp_int_SH_3_, u4_sll_480_temp_int_SH_4_, u4_sub_468_n16,
         u4_sub_468_n15, u4_sub_468_n14, u4_sub_468_n13, u4_sub_468_n12,
         u4_sub_468_n11, u4_sub_468_n10, u4_sub_468_n9, u4_sub_468_n8,
         u4_sub_468_n7, u4_sub_468_n6, u4_sub_468_n5, u4_sub_468_n4,
         u4_sub_468_n3, u4_sub_468_n2, u4_sub_468_n1, u4_sub_468_carry_1_,
         u4_sub_468_carry_2_, u4_sub_468_carry_3_, u4_sub_468_carry_4_,
         u4_sub_468_carry_5_, u4_sub_468_carry_6_, u4_sub_468_carry_7_,
         u4_sub_468_carry_8_, u4_sub_468_carry_9_, u4_sub_468_carry_10_,
         u4_sub_468_carry_11_, u4_sub_494_n14, u4_sub_494_n13, u4_sub_494_n12,
         u4_sub_494_n11, u4_sub_494_n10, u4_sub_494_n9, u4_sub_494_n8,
         u4_sub_494_n7, u4_sub_494_n6, u4_sub_494_n5, u4_sub_494_n4,
         u4_sub_494_n3, u4_sub_494_n2, u4_sub_494_n1, u4_sub_494_carry_1_,
         u4_sub_494_carry_2_, u4_sub_494_carry_3_, u4_sub_494_carry_4_,
         u4_sub_494_carry_5_, u4_sub_494_carry_6_, u4_sub_494_carry_7_,
         u4_sub_494_carry_8_, u4_sub_494_carry_9_, u4_sub_494_carry_10_,
         u4_add_487_n5, u4_add_487_n4, u4_add_487_carry_2_,
         u4_add_487_carry_3_, u4_add_487_carry_4_, u4_add_487_carry_5_,
         u4_add_492_n6, u4_add_492_n4, u4_add_492_n3, u4_add_492_carry_2_,
         u4_add_492_carry_3_, u4_add_492_carry_4_, u4_add_492_carry_5_,
         u4_add_492_carry_6_, u4_add_492_carry_7_, u4_add_492_carry_8_,
         u3_sub_61_n58, u3_sub_61_n57, u3_sub_61_n56, u3_sub_61_n55,
         u3_sub_61_n54, u3_sub_61_n53, u3_sub_61_n52, u3_sub_61_n51,
         u3_sub_61_n50, u3_sub_61_n49, u3_sub_61_n48, u3_sub_61_n47,
         u3_sub_61_n46, u3_sub_61_n45, u3_sub_61_n44, u3_sub_61_n43,
         u3_sub_61_n42, u3_sub_61_n41, u3_sub_61_n40, u3_sub_61_n39,
         u3_sub_61_n38, u3_sub_61_n37, u3_sub_61_n36, u3_sub_61_n35,
         u3_sub_61_n34, u3_sub_61_n33, u3_sub_61_n32, u3_sub_61_n31,
         u3_sub_61_n30, u3_sub_61_n29, u3_sub_61_n28, u3_sub_61_n27,
         u3_sub_61_n26, u3_sub_61_n25, u3_sub_61_n24, u3_sub_61_n23,
         u3_sub_61_n22, u3_sub_61_n21, u3_sub_61_n20, u3_sub_61_n19,
         u3_sub_61_n18, u3_sub_61_n17, u3_sub_61_n16, u3_sub_61_n15,
         u3_sub_61_n14, u3_sub_61_n13, u3_sub_61_n12, u3_sub_61_n11,
         u3_sub_61_n10, u3_sub_61_n9, u3_sub_61_n8, u3_sub_61_n7, u3_sub_61_n6,
         u3_sub_61_n5, u3_sub_61_n4, u3_sub_61_n3, u3_sub_61_n1, u3_add_61_n1,
         u2_add_111_n2, u2_sub_111_n13, u2_sub_111_n12, u2_sub_111_n11,
         u2_sub_111_n10, u2_sub_111_n9, u2_sub_111_n8, u2_sub_111_n7,
         u2_sub_111_n6, u2_sub_111_n5, u2_sub_111_n4, u2_sub_111_n3,
         u2_sub_111_n1, u1_gt_226_n167, u1_gt_226_n166, u1_gt_226_n165,
         u1_gt_226_n164, u1_gt_226_n163, u1_gt_226_n162, u1_gt_226_n161,
         u1_gt_226_n160, u1_gt_226_n159, u1_gt_226_n158, u1_gt_226_n157,
         u1_gt_226_n156, u1_gt_226_n155, u1_gt_226_n154, u1_gt_226_n153,
         u1_gt_226_n152, u1_gt_226_n151, u1_gt_226_n150, u1_gt_226_n149,
         u1_gt_226_n148, u1_gt_226_n147, u1_gt_226_n146, u1_gt_226_n145,
         u1_gt_226_n144, u1_gt_226_n143, u1_gt_226_n142, u1_gt_226_n141,
         u1_gt_226_n140, u1_gt_226_n139, u1_gt_226_n138, u1_gt_226_n137,
         u1_gt_226_n136, u1_gt_226_n135, u1_gt_226_n134, u1_gt_226_n133,
         u1_gt_226_n132, u1_gt_226_n131, u1_gt_226_n130, u1_gt_226_n129,
         u1_gt_226_n128, u1_gt_226_n127, u1_gt_226_n126, u1_gt_226_n125,
         u1_gt_226_n124, u1_gt_226_n123, u1_gt_226_n122, u1_gt_226_n121,
         u1_gt_226_n120, u1_gt_226_n119, u1_gt_226_n118, u1_gt_226_n117,
         u1_gt_226_n116, u1_gt_226_n115, u1_gt_226_n114, u1_gt_226_n113,
         u1_gt_226_n112, u1_gt_226_n111, u1_gt_226_n110, u1_gt_226_n109,
         u1_gt_226_n108, u1_gt_226_n107, u1_gt_226_n106, u1_gt_226_n105,
         u1_gt_226_n104, u1_gt_226_n103, u1_gt_226_n102, u1_gt_226_n101,
         u1_gt_226_n100, u1_gt_226_n99, u1_gt_226_n98, u1_gt_226_n97,
         u1_gt_226_n96, u1_gt_226_n95, u1_gt_226_n94, u1_gt_226_n93,
         u1_gt_226_n92, u1_gt_226_n91, u1_gt_226_n90, u1_gt_226_n89,
         u1_gt_226_n88, u1_gt_226_n87, u1_gt_226_n86, u1_gt_226_n85,
         u1_gt_226_n84, u1_gt_226_n83, u1_gt_226_n82, u1_gt_226_n81,
         u1_gt_226_n80, u1_gt_226_n79, u1_gt_226_n78, u1_gt_226_n77,
         u1_gt_226_n76, u1_gt_226_n75, u1_gt_226_n74, u1_gt_226_n73,
         u1_gt_226_n72, u1_gt_226_n71, u1_gt_226_n70, u1_gt_226_n69,
         u1_gt_226_n68, u1_gt_226_n67, u1_gt_226_n66, u1_gt_226_n65,
         u1_gt_226_n64, u1_gt_226_n63, u1_gt_226_n62, u1_gt_226_n61,
         u1_gt_226_n60, u1_gt_226_n59, u1_gt_226_n58, u1_gt_226_n57,
         u1_gt_226_n56, u1_gt_226_n55, u1_gt_226_n54, u1_gt_226_n53,
         u1_gt_226_n52, u1_gt_226_n51, u1_gt_226_n50, u1_gt_226_n49,
         u1_gt_226_n48, u1_gt_226_n47, u1_gt_226_n46, u1_gt_226_n45,
         u1_gt_226_n44, u1_gt_226_n43, u1_gt_226_n42, u1_gt_226_n41,
         u1_gt_226_n40, u1_gt_226_n39, u1_gt_226_n38, u1_gt_226_n37,
         u1_gt_226_n36, u1_gt_226_n35, u1_gt_226_n34, u1_gt_226_n33,
         u1_gt_226_n32, u1_gt_226_n31, u1_gt_226_n30, u1_gt_226_n29,
         u1_gt_226_n28, u1_gt_226_n27, u1_gt_226_n26, u1_gt_226_n25,
         u1_gt_226_n24, u1_gt_226_n23, u1_gt_226_n22, u1_gt_226_n21,
         u1_gt_226_n20, u1_gt_226_n19, u1_gt_226_n18, u1_gt_226_n17,
         u1_gt_226_n16, u1_gt_226_n15, u1_gt_226_n14, u1_gt_226_n13,
         u1_gt_226_n12, u1_gt_226_n11, u1_gt_226_n10, u1_gt_226_n9,
         u1_gt_226_n8, u1_gt_226_n7, u1_gt_226_n6, u1_gt_226_n5, u1_gt_226_n4,
         u1_gt_226_n3, u1_gt_226_n2, u1_gt_226_n1, u1_srl_148_n360,
         u1_srl_148_n359, u1_srl_148_n358, u1_srl_148_n357, u1_srl_148_n356,
         u1_srl_148_n355, u1_srl_148_n354, u1_srl_148_n353, u1_srl_148_n352,
         u1_srl_148_n351, u1_srl_148_n350, u1_srl_148_n349, u1_srl_148_n348,
         u1_srl_148_n347, u1_srl_148_n346, u1_srl_148_n345, u1_srl_148_n344,
         u1_srl_148_n343, u1_srl_148_n342, u1_srl_148_n341, u1_srl_148_n340,
         u1_srl_148_n339, u1_srl_148_n338, u1_srl_148_n337, u1_srl_148_n336,
         u1_srl_148_n335, u1_srl_148_n334, u1_srl_148_n333, u1_srl_148_n332,
         u1_srl_148_n331, u1_srl_148_n330, u1_srl_148_n329, u1_srl_148_n328,
         u1_srl_148_n327, u1_srl_148_n326, u1_srl_148_n325, u1_srl_148_n324,
         u1_srl_148_n323, u1_srl_148_n322, u1_srl_148_n321, u1_srl_148_n320,
         u1_srl_148_n319, u1_srl_148_n318, u1_srl_148_n317, u1_srl_148_n316,
         u1_srl_148_n315, u1_srl_148_n314, u1_srl_148_n313, u1_srl_148_n312,
         u1_srl_148_n311, u1_srl_148_n310, u1_srl_148_n309, u1_srl_148_n308,
         u1_srl_148_n307, u1_srl_148_n306, u1_srl_148_n305, u1_srl_148_n304,
         u1_srl_148_n303, u1_srl_148_n302, u1_srl_148_n301, u1_srl_148_n300,
         u1_srl_148_n299, u1_srl_148_n298, u1_srl_148_n297, u1_srl_148_n296,
         u1_srl_148_n295, u1_srl_148_n294, u1_srl_148_n293, u1_srl_148_n292,
         u1_srl_148_n291, u1_srl_148_n290, u1_srl_148_n289, u1_srl_148_n288,
         u1_srl_148_n287, u1_srl_148_n286, u1_srl_148_n285, u1_srl_148_n284,
         u1_srl_148_n283, u1_srl_148_n282, u1_srl_148_n281, u1_srl_148_n280,
         u1_srl_148_n279, u1_srl_148_n278, u1_srl_148_n277, u1_srl_148_n276,
         u1_srl_148_n275, u1_srl_148_n274, u1_srl_148_n273, u1_srl_148_n272,
         u1_srl_148_n271, u1_srl_148_n270, u1_srl_148_n269, u1_srl_148_n268,
         u1_srl_148_n267, u1_srl_148_n266, u1_srl_148_n265, u1_srl_148_n264,
         u1_srl_148_n263, u1_srl_148_n262, u1_srl_148_n261, u1_srl_148_n260,
         u1_srl_148_n259, u1_srl_148_n258, u1_srl_148_n257, u1_srl_148_n256,
         u1_srl_148_n255, u1_srl_148_n254, u1_srl_148_n253, u1_srl_148_n252,
         u1_srl_148_n251, u1_srl_148_n250, u1_srl_148_n249, u1_srl_148_n248,
         u1_srl_148_n247, u1_srl_148_n246, u1_srl_148_n245, u1_srl_148_n244,
         u1_srl_148_n243, u1_srl_148_n242, u1_srl_148_n241, u1_srl_148_n240,
         u1_srl_148_n239, u1_srl_148_n238, u1_srl_148_n237, u1_srl_148_n236,
         u1_srl_148_n235, u1_srl_148_n234, u1_srl_148_n233, u1_srl_148_n232,
         u1_srl_148_n231, u1_srl_148_n230, u1_srl_148_n229, u1_srl_148_n228,
         u1_srl_148_n227, u1_srl_148_n226, u1_srl_148_n225, u1_srl_148_n224,
         u1_srl_148_n223, u1_srl_148_n222, u1_srl_148_n221, u1_srl_148_n220,
         u1_srl_148_n219, u1_srl_148_n218, u1_srl_148_n217, u1_srl_148_n216,
         u1_srl_148_n215, u1_srl_148_n214, u1_srl_148_n213, u1_srl_148_n212,
         u1_srl_148_n211, u1_srl_148_n210, u1_srl_148_n209, u1_srl_148_n208,
         u1_srl_148_n207, u1_srl_148_n206, u1_srl_148_n205, u1_srl_148_n204,
         u1_srl_148_n203, u1_srl_148_n202, u1_srl_148_n201, u1_srl_148_n200,
         u1_srl_148_n199, u1_srl_148_n198, u1_srl_148_n197, u1_srl_148_n196,
         u1_srl_148_n195, u1_srl_148_n194, u1_srl_148_n193, u1_srl_148_n192,
         u1_srl_148_n191, u1_srl_148_n190, u1_srl_148_n189, u1_srl_148_n188,
         u1_srl_148_n187, u1_srl_148_n186, u1_srl_148_n185, u1_srl_148_n184,
         u1_srl_148_n183, u1_srl_148_n182, u1_srl_148_n181, u1_srl_148_n180,
         u1_srl_148_n179, u1_srl_148_n178, u1_srl_148_n177, u1_srl_148_n176,
         u1_srl_148_n175, u1_srl_148_n174, u1_srl_148_n173, u1_srl_148_n172,
         u1_srl_148_n171, u1_srl_148_n170, u1_srl_148_n169, u1_srl_148_n168,
         u1_srl_148_n167, u1_srl_148_n166, u1_srl_148_n165, u1_srl_148_n164,
         u1_srl_148_n163, u1_srl_148_n162, u1_srl_148_n161, u1_srl_148_n160,
         u1_srl_148_n159, u1_srl_148_n158, u1_srl_148_n157, u1_srl_148_n156,
         u1_srl_148_n155, u1_srl_148_n154, u1_srl_148_n153, u1_srl_148_n152,
         u1_srl_148_n151, u1_srl_148_n150, u1_srl_148_n149, u1_srl_148_n148,
         u1_srl_148_n147, u1_srl_148_n146, u1_srl_148_n145, u1_srl_148_n144,
         u1_srl_148_n143, u1_srl_148_n142, u1_srl_148_n141, u1_srl_148_n140,
         u1_srl_148_n139, u1_srl_148_n138, u1_srl_148_n137, u1_srl_148_n136,
         u1_srl_148_n135, u1_srl_148_n134, u1_srl_148_n133, u1_srl_148_n132,
         u1_srl_148_n131, u1_srl_148_n130, u1_srl_148_n129, u1_srl_148_n128,
         u1_srl_148_n127, u1_srl_148_n126, u1_srl_148_n125, u1_srl_148_n124,
         u1_srl_148_n123, u1_srl_148_n122, u1_srl_148_n121, u1_srl_148_n120,
         u1_srl_148_n119, u1_srl_148_n118, u1_srl_148_n117, u1_srl_148_n116,
         u1_srl_148_n115, u1_srl_148_n114, u1_srl_148_n113, u1_srl_148_n112,
         u1_srl_148_n111, u1_srl_148_n110, u1_srl_148_n109, u1_srl_148_n108,
         u1_srl_148_n107, u1_srl_148_n106, u1_srl_148_n105, u1_srl_148_n104,
         u1_srl_148_n103, u1_srl_148_n102, u1_srl_148_n101, u1_srl_148_n100,
         u1_srl_148_n99, u1_srl_148_n98, u1_srl_148_n97, u1_srl_148_n96,
         u1_srl_148_n95, u1_srl_148_n94, u1_srl_148_n93, u1_srl_148_n92,
         u1_srl_148_n91, u1_srl_148_n90, u1_srl_148_n89, u1_srl_148_n88,
         u1_srl_148_n87, u1_srl_148_n86, u1_srl_148_n85, u1_srl_148_n84,
         u1_srl_148_n83, u1_srl_148_n82, u1_srl_148_n81, u1_srl_148_n80,
         u1_srl_148_n79, u1_srl_148_n78, u1_srl_148_n77, u1_srl_148_n76,
         u1_srl_148_n75, u1_srl_148_n74, u1_srl_148_n73, u1_srl_148_n72,
         u1_srl_148_n71, u1_srl_148_n70, u1_srl_148_n69, u1_srl_148_n68,
         u1_srl_148_n67, u1_srl_148_n66, u1_srl_148_n65, u1_srl_148_n64,
         u1_srl_148_n63, u1_srl_148_n62, u1_srl_148_n61, u1_srl_148_n60,
         u1_srl_148_n59, u1_srl_148_n58, u1_srl_148_n57, u1_srl_148_n56,
         u1_srl_148_n55, u1_srl_148_n54, u1_srl_148_n53, u1_srl_148_n52,
         u1_srl_148_n51, u1_srl_148_n50, u1_srl_148_n49, u1_srl_148_n48,
         u1_srl_148_n47, u1_srl_148_n46, u1_srl_148_n45, u1_srl_148_n44,
         u1_srl_148_n43, u1_srl_148_n42, u1_srl_148_n41, u1_srl_148_n40,
         u1_srl_148_n39, u1_srl_148_n38, u1_srl_148_n37, u1_srl_148_n36,
         u1_srl_148_n35, u1_srl_148_n34, u1_srl_148_n33, u1_srl_148_n32,
         u1_srl_148_n31, u1_srl_148_n30, u1_srl_148_n29, u1_srl_148_n28,
         u1_srl_148_n27, u1_srl_148_n26, u1_srl_148_n25, u1_srl_148_n24,
         u1_srl_148_n23, u1_srl_148_n22, u1_srl_148_n21, u1_srl_148_n20,
         u1_srl_148_n19, u1_srl_148_n18, u1_srl_148_n17, u1_srl_148_n16,
         u1_srl_148_n15, u1_srl_148_n14, u1_srl_148_n13, u1_srl_148_n12,
         u1_srl_148_n11, u1_srl_148_n10, u1_srl_148_n9, u1_srl_148_n8,
         u1_srl_148_n7, u1_srl_148_n6, u1_srl_148_n5, u1_srl_148_n4,
         u1_srl_148_n3, u1_srl_148_n2, u1_srl_148_n1,
         sub_1_root_u1_sub_130_aco_n12, sub_1_root_u1_sub_130_aco_n11,
         sub_1_root_u1_sub_130_aco_n10, sub_1_root_u1_sub_130_aco_n9,
         sub_1_root_u1_sub_130_aco_n8, sub_1_root_u1_sub_130_aco_n7,
         sub_1_root_u1_sub_130_aco_n6, sub_1_root_u1_sub_130_aco_n5,
         sub_1_root_u1_sub_130_aco_n4, sub_1_root_u1_sub_130_aco_n3,
         sub_1_root_u1_sub_130_aco_n2, sub_1_root_u1_sub_130_aco_n1,
         sub_430_3_n171, sub_430_3_n170, sub_430_3_n169, sub_430_3_n168,
         sub_430_3_n167, sub_430_3_n166, sub_430_3_n165, sub_430_3_n164,
         sub_430_3_n163, sub_430_3_n162, sub_430_3_n161, sub_430_3_n160,
         sub_430_3_n159, sub_430_3_n158, sub_430_3_n157, sub_430_3_n156,
         sub_430_3_n155, sub_430_3_n154, sub_430_3_n153, sub_430_3_n152,
         sub_430_3_n151, sub_430_3_n150, sub_430_3_n149, sub_430_3_n148,
         sub_430_3_n147, sub_430_3_n146, sub_430_3_n145, sub_430_3_n144,
         sub_430_3_n143, sub_430_3_n142, sub_430_3_n141, sub_430_3_n140,
         sub_430_3_n139, sub_430_3_n138, sub_430_3_n137, sub_430_3_n136,
         sub_430_3_n135, sub_430_3_n134, sub_430_3_n133, sub_430_3_n132,
         sub_430_3_n131, sub_430_3_n130, sub_430_3_n129, sub_430_3_n128,
         sub_430_3_n127, sub_430_3_n126, sub_430_3_n125, sub_430_3_n124,
         sub_430_3_n123, sub_430_3_n122, sub_430_3_n121, sub_430_3_n120,
         sub_430_3_n119, sub_430_3_n118, sub_430_3_n117, sub_430_3_n116,
         sub_430_3_n115, sub_430_3_n114, sub_430_3_n102, sub_430_3_n101,
         sub_430_3_n100, sub_430_3_n99, sub_430_3_n98, sub_430_3_n97,
         sub_430_3_n96, sub_430_3_n95, sub_430_3_n94, sub_430_3_n93,
         sub_430_3_n92, sub_430_3_n91, sub_430_3_n90, sub_430_3_n89,
         sub_430_3_n88, sub_430_3_n87, sub_430_3_n86, sub_430_3_n85,
         sub_430_3_n84, sub_430_3_n83, sub_430_3_n82, sub_430_3_n81,
         sub_430_3_n80, sub_430_3_n79, sub_430_3_n46, sub_430_3_n45,
         sub_430_3_n44, sub_430_3_n43, sub_430_3_n42, sub_430_3_n41,
         sub_430_3_n40, sub_430_3_n39, sub_430_3_n38, sub_430_3_n37,
         sub_430_3_n36, sub_430_3_n35, sub_430_3_n31, sub_430_3_n30,
         sub_430_3_n29, sub_430_3_n28, sub_430_3_n27, sub_430_3_n26,
         sub_430_3_n25, sub_430_3_n24, sub_430_3_n23, sub_430_3_n22,
         sub_430_3_n21, sub_430_3_n20, sub_430_3_n19, sub_430_3_n18,
         sub_430_3_n17, sub_430_3_n16, sub_430_3_n15, sub_430_3_n14,
         sub_430_3_n13, sub_430_3_n12, sub_430_b0_n157, sub_430_b0_n156,
         sub_430_b0_n155, sub_430_b0_n154, sub_430_b0_n153, sub_430_b0_n152,
         sub_430_b0_n151, sub_430_b0_n150, sub_430_b0_n149, sub_430_b0_n148,
         sub_430_b0_n147, sub_430_b0_n146, sub_430_b0_n145, sub_430_b0_n144,
         sub_430_b0_n143, sub_430_b0_n142, sub_430_b0_n141, sub_430_b0_n140,
         sub_430_b0_n139, sub_430_b0_n138, sub_430_b0_n137, sub_430_b0_n136,
         sub_430_b0_n135, sub_430_b0_n134, sub_430_b0_n133, sub_430_b0_n132,
         sub_430_b0_n131, sub_430_b0_n130, sub_430_b0_n129, sub_430_b0_n128,
         sub_430_b0_n127, sub_430_b0_n126, sub_430_b0_n125, sub_430_b0_n124,
         sub_430_b0_n123, sub_430_b0_n122, sub_430_b0_n121, sub_430_b0_n120,
         sub_430_b0_n119, sub_430_b0_n118, sub_430_b0_n117, sub_430_b0_n116,
         sub_430_b0_n115, sub_430_b0_n114, sub_430_b0_n113, sub_430_b0_n112,
         sub_430_b0_n111, sub_430_b0_n110, sub_430_b0_n109, sub_430_b0_n108,
         sub_430_b0_n107, sub_430_b0_n106, sub_430_b0_n105, sub_430_b0_n68,
         sub_430_b0_n67, sub_430_b0_n66, sub_430_b0_n65, sub_430_b0_n64,
         sub_430_b0_n63, sub_430_b0_n62, sub_430_b0_n61, sub_430_b0_n60,
         sub_430_b0_n59, sub_430_b0_n58, sub_430_b0_n57, sub_430_b0_n56,
         sub_430_b0_n55, sub_430_b0_n54, sub_430_b0_n53, sub_430_b0_n52,
         sub_430_b0_n51, sub_430_b0_n50, sub_430_b0_n49, sub_430_b0_n48,
         sub_430_b0_n47, sub_430_b0_n46, sub_430_b0_n45, sub_430_b0_n44,
         sub_430_b0_n43, sub_430_b0_n25, sub_430_b0_n24, sub_430_b0_n23,
         sub_430_b0_n22, sub_430_b0_n21, sub_430_b0_n20, sub_430_b0_n19,
         sub_430_b0_n18, sub_430_b0_n17, sub_430_b0_n16, sub_430_b0_n15,
         sub_430_b0_n14, sub_430_b0_n13, sub_430_b0_n12, sub_430_b0_n11,
         sub_430_b0_n10, sub_430_b0_n9, sub_430_b0_n8, sub_430_b0_n7,
         sub_430_b0_n6, sub_430_b0_n5, sub_430_b0_n4, sub_430_b0_n3,
         sub_430_b0_n2, sub_430_b0_n1, sll_381_n30, sll_381_n29, sll_381_n28,
         sll_381_n27, sll_381_n26, sll_381_n25, sll_381_n24, sll_381_n23,
         sll_381_n22, sll_381_n21, sll_381_n20, sll_381_n19, sll_381_n18,
         sll_381_n17, sll_381_n16, sll_381_n15, sll_381_n14, sll_381_n13,
         sll_381_n12, sll_381_n11, sll_381_n10, sll_381_n9, sll_381_n8,
         sll_381_n7, sll_381_n6, sll_381_n5, sll_381_n4, sll_381_n3,
         sll_381_n2, sll_381_n1, sll_381_ML_int_4__8_, sll_381_ML_int_4__9_,
         sll_381_ML_int_4__10_, sll_381_ML_int_4__11_, sll_381_ML_int_4__12_,
         sll_381_ML_int_4__13_, sll_381_ML_int_4__14_, sll_381_ML_int_4__15_,
         sll_381_ML_int_4__16_, sll_381_ML_int_4__17_, sll_381_ML_int_4__18_,
         sll_381_ML_int_4__19_, sll_381_ML_int_4__20_, sll_381_ML_int_4__21_,
         sll_381_ML_int_4__22_, sll_381_ML_int_4__23_, sll_381_ML_int_4__24_,
         sll_381_ML_int_4__25_, sll_381_ML_int_4__26_, sll_381_ML_int_4__27_,
         sll_381_ML_int_4__28_, sll_381_ML_int_4__29_, sll_381_ML_int_4__30_,
         sll_381_ML_int_4__31_, sll_381_ML_int_4__32_, sll_381_ML_int_4__33_,
         sll_381_ML_int_4__34_, sll_381_ML_int_4__35_, sll_381_ML_int_4__36_,
         sll_381_ML_int_4__37_, sll_381_ML_int_4__38_, sll_381_ML_int_4__39_,
         sll_381_ML_int_4__40_, sll_381_ML_int_4__41_, sll_381_ML_int_4__42_,
         sll_381_ML_int_4__43_, sll_381_ML_int_4__44_, sll_381_ML_int_4__45_,
         sll_381_ML_int_4__46_, sll_381_ML_int_4__47_, sll_381_ML_int_4__48_,
         sll_381_ML_int_4__49_, sll_381_ML_int_4__50_, sll_381_ML_int_4__51_,
         sll_381_ML_int_4__52_, sll_381_ML_int_3__0_, sll_381_ML_int_3__1_,
         sll_381_ML_int_3__2_, sll_381_ML_int_3__3_, sll_381_ML_int_3__4_,
         sll_381_ML_int_3__5_, sll_381_ML_int_3__6_, sll_381_ML_int_3__7_,
         sll_381_ML_int_3__8_, sll_381_ML_int_3__9_, sll_381_ML_int_3__10_,
         sll_381_ML_int_3__11_, sll_381_ML_int_3__12_, sll_381_ML_int_3__13_,
         sll_381_ML_int_3__14_, sll_381_ML_int_3__15_, sll_381_ML_int_3__16_,
         sll_381_ML_int_3__17_, sll_381_ML_int_3__18_, sll_381_ML_int_3__19_,
         sll_381_ML_int_3__20_, sll_381_ML_int_3__21_, sll_381_ML_int_3__22_,
         sll_381_ML_int_3__23_, sll_381_ML_int_3__24_, sll_381_ML_int_3__25_,
         sll_381_ML_int_3__26_, sll_381_ML_int_3__27_, sll_381_ML_int_3__28_,
         sll_381_ML_int_3__29_, sll_381_ML_int_3__30_, sll_381_ML_int_3__31_,
         sll_381_ML_int_3__32_, sll_381_ML_int_3__33_, sll_381_ML_int_3__34_,
         sll_381_ML_int_3__35_, sll_381_ML_int_3__36_, sll_381_ML_int_3__37_,
         sll_381_ML_int_3__38_, sll_381_ML_int_3__39_, sll_381_ML_int_3__40_,
         sll_381_ML_int_3__41_, sll_381_ML_int_3__42_, sll_381_ML_int_3__43_,
         sll_381_ML_int_3__44_, sll_381_ML_int_3__45_, sll_381_ML_int_3__46_,
         sll_381_ML_int_3__47_, sll_381_ML_int_3__48_, sll_381_ML_int_3__49_,
         sll_381_ML_int_3__50_, sll_381_ML_int_3__51_, sll_381_ML_int_3__52_,
         sll_381_ML_int_2__0_, sll_381_ML_int_2__1_, sll_381_ML_int_2__2_,
         sll_381_ML_int_2__3_, sll_381_ML_int_2__4_, sll_381_ML_int_2__5_,
         sll_381_ML_int_2__6_, sll_381_ML_int_2__7_, sll_381_ML_int_2__8_,
         sll_381_ML_int_2__9_, sll_381_ML_int_2__10_, sll_381_ML_int_2__11_,
         sll_381_ML_int_2__12_, sll_381_ML_int_2__13_, sll_381_ML_int_2__14_,
         sll_381_ML_int_2__15_, sll_381_ML_int_2__16_, sll_381_ML_int_2__17_,
         sll_381_ML_int_2__18_, sll_381_ML_int_2__19_, sll_381_ML_int_2__20_,
         sll_381_ML_int_2__21_, sll_381_ML_int_2__22_, sll_381_ML_int_2__23_,
         sll_381_ML_int_2__24_, sll_381_ML_int_2__25_, sll_381_ML_int_2__26_,
         sll_381_ML_int_2__27_, sll_381_ML_int_2__28_, sll_381_ML_int_2__29_,
         sll_381_ML_int_2__30_, sll_381_ML_int_2__31_, sll_381_ML_int_2__32_,
         sll_381_ML_int_2__33_, sll_381_ML_int_2__34_, sll_381_ML_int_2__35_,
         sll_381_ML_int_2__36_, sll_381_ML_int_2__37_, sll_381_ML_int_2__38_,
         sll_381_ML_int_2__39_, sll_381_ML_int_2__40_, sll_381_ML_int_2__41_,
         sll_381_ML_int_2__42_, sll_381_ML_int_2__43_, sll_381_ML_int_2__44_,
         sll_381_ML_int_2__45_, sll_381_ML_int_2__46_, sll_381_ML_int_2__47_,
         sll_381_ML_int_2__48_, sll_381_ML_int_2__49_, sll_381_ML_int_2__50_,
         sll_381_ML_int_2__51_, sll_381_ML_int_2__52_, sll_381_ML_int_1__0_,
         sll_381_ML_int_1__1_, sll_381_ML_int_1__2_, sll_381_ML_int_1__3_,
         sll_381_ML_int_1__4_, sll_381_ML_int_1__5_, sll_381_ML_int_1__6_,
         sll_381_ML_int_1__7_, sll_381_ML_int_1__8_, sll_381_ML_int_1__9_,
         sll_381_ML_int_1__10_, sll_381_ML_int_1__11_, sll_381_ML_int_1__12_,
         sll_381_ML_int_1__13_, sll_381_ML_int_1__14_, sll_381_ML_int_1__15_,
         sll_381_ML_int_1__16_, sll_381_ML_int_1__17_, sll_381_ML_int_1__18_,
         sll_381_ML_int_1__19_, sll_381_ML_int_1__20_, sll_381_ML_int_1__21_,
         sll_381_ML_int_1__22_, sll_381_ML_int_1__23_, sll_381_ML_int_1__24_,
         sll_381_ML_int_1__25_, sll_381_ML_int_1__26_, sll_381_ML_int_1__27_,
         sll_381_ML_int_1__28_, sll_381_ML_int_1__29_, sll_381_ML_int_1__30_,
         sll_381_ML_int_1__31_, sll_381_ML_int_1__32_, sll_381_ML_int_1__33_,
         sll_381_ML_int_1__34_, sll_381_ML_int_1__35_, sll_381_ML_int_1__36_,
         sll_381_ML_int_1__37_, sll_381_ML_int_1__38_, sll_381_ML_int_1__39_,
         sll_381_ML_int_1__40_, sll_381_ML_int_1__41_, sll_381_ML_int_1__42_,
         sll_381_ML_int_1__43_, sll_381_ML_int_1__44_, sll_381_ML_int_1__45_,
         sll_381_ML_int_1__46_, sll_381_ML_int_1__47_, sll_381_ML_int_1__48_,
         sll_381_ML_int_1__49_, sll_381_ML_int_1__50_, sll_381_ML_int_1__51_,
         sll_381_ML_int_1__52_, r466_n178, r466_n177, r466_n176, r466_n175,
         r466_n174, r466_n173, r466_n172, r466_n171, r466_n170, r466_n169,
         r466_n168, r466_n167, r466_n166, r466_n165, r466_n164, r466_n163,
         r466_n162, r466_n161, r466_n160, r466_n159, r466_n158, r466_n157,
         r466_n156, r466_n155, r466_n154, r466_n153, r466_n152, r466_n151,
         r466_n150, r466_n149, r466_n148, r466_n147, r466_n146, r466_n145,
         r466_n144, r466_n143, r466_n142, r466_n141, r466_n140, r466_n139,
         r466_n138, r466_n137, r466_n136, r466_n135, r466_n134, r466_n133,
         r466_n132, r466_n131, r466_n130, r466_n129, r466_n128, r466_n127,
         r466_n126, r466_n125, r466_n124, r466_n123, r466_n122, r466_n121,
         r466_n120, r466_n119, r466_n118, r466_n117, r466_n116, r466_n115,
         r466_n114, r466_n113, r466_n112, r466_n111, r466_n110, r466_n109,
         r466_n108, r466_n107, r466_n106, r466_n105, r466_n104, r466_n103,
         r466_n102, r466_n101, r466_n100, r466_n99, r466_n98, r466_n97,
         r466_n96, r466_n95, r466_n94, r466_n93, r466_n92, r466_n91, r466_n90,
         r466_n89, r466_n88, r466_n87, r466_n86, r466_n85, r466_n84, r466_n83,
         r466_n82, r466_n81, r466_n80, r466_n79, r466_n78, r466_n77, r466_n76,
         r466_n75, r466_n74, r466_n73, r466_n72, r466_n71, r466_n70, r466_n69,
         r466_n68, r466_n67, r466_n66, r466_n65, r466_n64, r466_n63, r466_n62,
         r466_n61, r466_n60, r466_n59, r466_n58, r466_n57, r466_n56, r466_n55,
         r466_n54, r466_n53, r466_n52, r466_n51, r466_n50, r466_n49, r466_n48,
         r466_n47, r466_n46, r466_n45, r466_n44, r466_n43, r466_n42, r466_n41,
         r466_n40, r466_n39, r466_n38, r466_n37, r466_n36, r466_n35, r466_n34,
         r466_n33, r466_n32, r466_n31, r466_n30, r466_n29, r466_n28, r466_n27,
         r466_n26, r466_n25, r466_n24, r466_n23, r466_n22, r466_n21, r466_n20,
         r466_n19, r466_n18, r466_n17, r466_n16, r466_n15, r466_n14, r466_n13,
         r466_n12, r466_n11, r466_n10, r466_n9, r466_n8, r466_n7, r466_n6,
         r466_n5, r466_n4, r466_n3, r466_n2, r466_n1,
         add_0_root_sub_0_root_u4_add_495_n1, u5_mult_87_n482, u5_mult_87_n481,
         u5_mult_87_n480, u5_mult_87_n479, u5_mult_87_n478, u5_mult_87_n477,
         u5_mult_87_n476, u5_mult_87_n475, u5_mult_87_n474, u5_mult_87_n473,
         u5_mult_87_n472, u5_mult_87_n471, u5_mult_87_n470, u5_mult_87_n469,
         u5_mult_87_n468, u5_mult_87_n467, u5_mult_87_n466, u5_mult_87_n465,
         u5_mult_87_n464, u5_mult_87_n463, u5_mult_87_n462, u5_mult_87_n461,
         u5_mult_87_n460, u5_mult_87_n459, u5_mult_87_n458, u5_mult_87_n457,
         u5_mult_87_n456, u5_mult_87_n455, u5_mult_87_n454, u5_mult_87_n453,
         u5_mult_87_n452, u5_mult_87_n451, u5_mult_87_n450, u5_mult_87_n449,
         u5_mult_87_n448, u5_mult_87_n447, u5_mult_87_n446, u5_mult_87_n445,
         u5_mult_87_n444, u5_mult_87_n443, u5_mult_87_n442, u5_mult_87_n441,
         u5_mult_87_n440, u5_mult_87_n439, u5_mult_87_n438, u5_mult_87_n437,
         u5_mult_87_n436, u5_mult_87_n435, u5_mult_87_n434, u5_mult_87_n433,
         u5_mult_87_n432, u5_mult_87_n431, u5_mult_87_n430, u5_mult_87_n429,
         u5_mult_87_n428, u5_mult_87_n427, u5_mult_87_n426, u5_mult_87_n425,
         u5_mult_87_n424, u5_mult_87_n423, u5_mult_87_n422, u5_mult_87_n421,
         u5_mult_87_n420, u5_mult_87_n419, u5_mult_87_n418, u5_mult_87_n417,
         u5_mult_87_n416, u5_mult_87_n415, u5_mult_87_n414, u5_mult_87_n413,
         u5_mult_87_n412, u5_mult_87_n411, u5_mult_87_n410, u5_mult_87_n409,
         u5_mult_87_n408, u5_mult_87_n407, u5_mult_87_n406, u5_mult_87_n405,
         u5_mult_87_n404, u5_mult_87_n403, u5_mult_87_n402, u5_mult_87_n401,
         u5_mult_87_n400, u5_mult_87_n399, u5_mult_87_n398, u5_mult_87_n397,
         u5_mult_87_n396, u5_mult_87_n395, u5_mult_87_n394, u5_mult_87_n393,
         u5_mult_87_n392, u5_mult_87_n391, u5_mult_87_n390, u5_mult_87_n389,
         u5_mult_87_n388, u5_mult_87_n387, u5_mult_87_n386, u5_mult_87_n385,
         u5_mult_87_n384, u5_mult_87_n383, u5_mult_87_n382, u5_mult_87_n381,
         u5_mult_87_n380, u5_mult_87_n379, u5_mult_87_n378, u5_mult_87_n377,
         u5_mult_87_n376, u5_mult_87_n375, u5_mult_87_n374, u5_mult_87_n373,
         u5_mult_87_n372, u5_mult_87_n371, u5_mult_87_n370, u5_mult_87_n369,
         u5_mult_87_n368, u5_mult_87_n367, u5_mult_87_n366, u5_mult_87_n365,
         u5_mult_87_n364, u5_mult_87_n363, u5_mult_87_n362, u5_mult_87_n361,
         u5_mult_87_n360, u5_mult_87_n359, u5_mult_87_n358, u5_mult_87_n357,
         u5_mult_87_n356, u5_mult_87_n355, u5_mult_87_n354, u5_mult_87_n353,
         u5_mult_87_n352, u5_mult_87_n351, u5_mult_87_n350, u5_mult_87_n349,
         u5_mult_87_n348, u5_mult_87_n347, u5_mult_87_n346, u5_mult_87_n345,
         u5_mult_87_n344, u5_mult_87_n343, u5_mult_87_n342, u5_mult_87_n341,
         u5_mult_87_n340, u5_mult_87_n339, u5_mult_87_n338, u5_mult_87_n337,
         u5_mult_87_n336, u5_mult_87_n335, u5_mult_87_n334, u5_mult_87_n333,
         u5_mult_87_n332, u5_mult_87_n331, u5_mult_87_n330, u5_mult_87_n329,
         u5_mult_87_n328, u5_mult_87_n327, u5_mult_87_n326, u5_mult_87_n325,
         u5_mult_87_n324, u5_mult_87_n323, u5_mult_87_n322, u5_mult_87_n321,
         u5_mult_87_n320, u5_mult_87_n319, u5_mult_87_n318, u5_mult_87_n317,
         u5_mult_87_n316, u5_mult_87_n315, u5_mult_87_n314, u5_mult_87_n313,
         u5_mult_87_n312, u5_mult_87_n311, u5_mult_87_n310, u5_mult_87_n309,
         u5_mult_87_n308, u5_mult_87_n307, u5_mult_87_n306, u5_mult_87_n305,
         u5_mult_87_n304, u5_mult_87_n303, u5_mult_87_n302, u5_mult_87_n301,
         u5_mult_87_n300, u5_mult_87_n299, u5_mult_87_n298, u5_mult_87_n297,
         u5_mult_87_n296, u5_mult_87_n295, u5_mult_87_n294, u5_mult_87_n293,
         u5_mult_87_n292, u5_mult_87_n291, u5_mult_87_n290, u5_mult_87_n289,
         u5_mult_87_n288, u5_mult_87_n287, u5_mult_87_n286, u5_mult_87_n285,
         u5_mult_87_n284, u5_mult_87_n283, u5_mult_87_n282, u5_mult_87_n281,
         u5_mult_87_n280, u5_mult_87_n279, u5_mult_87_n278, u5_mult_87_n277,
         u5_mult_87_n276, u5_mult_87_n275, u5_mult_87_n274, u5_mult_87_n273,
         u5_mult_87_n272, u5_mult_87_n271, u5_mult_87_n270, u5_mult_87_n269,
         u5_mult_87_n268, u5_mult_87_n267, u5_mult_87_n266, u5_mult_87_n265,
         u5_mult_87_n264, u5_mult_87_n263, u5_mult_87_n262, u5_mult_87_n261,
         u5_mult_87_n260, u5_mult_87_n259, u5_mult_87_n258, u5_mult_87_n257,
         u5_mult_87_n256, u5_mult_87_n255, u5_mult_87_n254, u5_mult_87_n253,
         u5_mult_87_n252, u5_mult_87_n251, u5_mult_87_n250, u5_mult_87_n249,
         u5_mult_87_n248, u5_mult_87_n247, u5_mult_87_n246, u5_mult_87_n245,
         u5_mult_87_n244, u5_mult_87_n243, u5_mult_87_n242, u5_mult_87_n241,
         u5_mult_87_n240, u5_mult_87_n239, u5_mult_87_n238, u5_mult_87_n237,
         u5_mult_87_n236, u5_mult_87_n235, u5_mult_87_n234, u5_mult_87_n233,
         u5_mult_87_n232, u5_mult_87_n231, u5_mult_87_n230, u5_mult_87_n229,
         u5_mult_87_n228, u5_mult_87_n227, u5_mult_87_n226, u5_mult_87_n225,
         u5_mult_87_n224, u5_mult_87_n223, u5_mult_87_n222, u5_mult_87_n221,
         u5_mult_87_n220, u5_mult_87_n219, u5_mult_87_n218, u5_mult_87_n217,
         u5_mult_87_n216, u5_mult_87_n215, u5_mult_87_n214, u5_mult_87_n213,
         u5_mult_87_n212, u5_mult_87_n211, u5_mult_87_n210, u5_mult_87_n208,
         u5_mult_87_n206, u5_mult_87_n205, u5_mult_87_n204, u5_mult_87_n203,
         u5_mult_87_n202, u5_mult_87_n201, u5_mult_87_n200, u5_mult_87_n199,
         u5_mult_87_n198, u5_mult_87_n197, u5_mult_87_n196, u5_mult_87_n195,
         u5_mult_87_n194, u5_mult_87_n193, u5_mult_87_n192, u5_mult_87_n191,
         u5_mult_87_n190, u5_mult_87_n189, u5_mult_87_n188, u5_mult_87_n187,
         u5_mult_87_n186, u5_mult_87_n185, u5_mult_87_n184, u5_mult_87_n183,
         u5_mult_87_n182, u5_mult_87_n181, u5_mult_87_n180, u5_mult_87_n179,
         u5_mult_87_n178, u5_mult_87_n177, u5_mult_87_n176, u5_mult_87_n175,
         u5_mult_87_n174, u5_mult_87_n173, u5_mult_87_n172, u5_mult_87_n171,
         u5_mult_87_n170, u5_mult_87_n169, u5_mult_87_n168, u5_mult_87_n167,
         u5_mult_87_n166, u5_mult_87_n165, u5_mult_87_n164, u5_mult_87_n163,
         u5_mult_87_n162, u5_mult_87_n161, u5_mult_87_n160, u5_mult_87_n159,
         u5_mult_87_n158, u5_mult_87_n157, u5_mult_87_n156, u5_mult_87_n155,
         u5_mult_87_n154, u5_mult_87_n153, u5_mult_87_n152, u5_mult_87_n151,
         u5_mult_87_n150, u5_mult_87_n149, u5_mult_87_n148, u5_mult_87_n147,
         u5_mult_87_n146, u5_mult_87_n145, u5_mult_87_n144, u5_mult_87_n143,
         u5_mult_87_n142, u5_mult_87_n141, u5_mult_87_n140, u5_mult_87_n139,
         u5_mult_87_n138, u5_mult_87_n137, u5_mult_87_n136, u5_mult_87_n135,
         u5_mult_87_n134, u5_mult_87_n133, u5_mult_87_n132, u5_mult_87_n131,
         u5_mult_87_n130, u5_mult_87_n129, u5_mult_87_n128, u5_mult_87_n127,
         u5_mult_87_n126, u5_mult_87_n125, u5_mult_87_n124, u5_mult_87_n123,
         u5_mult_87_n122, u5_mult_87_n121, u5_mult_87_n120, u5_mult_87_n119,
         u5_mult_87_n118, u5_mult_87_n117, u5_mult_87_n116, u5_mult_87_n115,
         u5_mult_87_n114, u5_mult_87_n113, u5_mult_87_n112, u5_mult_87_n111,
         u5_mult_87_n110, u5_mult_87_n109, u5_mult_87_n108, u5_mult_87_n107,
         u5_mult_87_n106, u5_mult_87_n105, u5_mult_87_n104, u5_mult_87_n103,
         u5_mult_87_n102, u5_mult_87_n101, u5_mult_87_n100, u5_mult_87_n99,
         u5_mult_87_n98, u5_mult_87_n97, u5_mult_87_n96, u5_mult_87_n95,
         u5_mult_87_n94, u5_mult_87_n93, u5_mult_87_n92, u5_mult_87_n91,
         u5_mult_87_n90, u5_mult_87_n89, u5_mult_87_n88, u5_mult_87_n87,
         u5_mult_87_n86, u5_mult_87_n85, u5_mult_87_n84, u5_mult_87_n83,
         u5_mult_87_n82, u5_mult_87_n81, u5_mult_87_n80, u5_mult_87_n79,
         u5_mult_87_n78, u5_mult_87_n77, u5_mult_87_n76, u5_mult_87_n75,
         u5_mult_87_n74, u5_mult_87_n73, u5_mult_87_n72, u5_mult_87_n71,
         u5_mult_87_n70, u5_mult_87_n69, u5_mult_87_n68, u5_mult_87_n67,
         u5_mult_87_n66, u5_mult_87_n65, u5_mult_87_n64, u5_mult_87_n63,
         u5_mult_87_n62, u5_mult_87_n61, u5_mult_87_n60, u5_mult_87_n59,
         u5_mult_87_n58, u5_mult_87_n57, u5_mult_87_n56, u5_mult_87_n55,
         u5_mult_87_n54, u5_mult_87_n53, u5_mult_87_n52, u5_mult_87_n51,
         u5_mult_87_n50, u5_mult_87_n49, u5_mult_87_n48, u5_mult_87_n47,
         u5_mult_87_n46, u5_mult_87_n45, u5_mult_87_n44, u5_mult_87_n43,
         u5_mult_87_n42, u5_mult_87_n41, u5_mult_87_n40, u5_mult_87_n39,
         u5_mult_87_n38, u5_mult_87_n37, u5_mult_87_n36, u5_mult_87_n35,
         u5_mult_87_n34, u5_mult_87_n33, u5_mult_87_n32, u5_mult_87_n31,
         u5_mult_87_n30, u5_mult_87_n29, u5_mult_87_n28, u5_mult_87_n27,
         u5_mult_87_n26, u5_mult_87_n25, u5_mult_87_n24, u5_mult_87_n23,
         u5_mult_87_n22, u5_mult_87_n21, u5_mult_87_n20, u5_mult_87_n19,
         u5_mult_87_n18, u5_mult_87_n17, u5_mult_87_n16, u5_mult_87_n15,
         u5_mult_87_n14, u5_mult_87_n13, u5_mult_87_n12, u5_mult_87_n11,
         u5_mult_87_n10, u5_mult_87_n9, u5_mult_87_n8, u5_mult_87_n7,
         u5_mult_87_n6, u5_mult_87_n5, u5_mult_87_n4, u5_mult_87_n3,
         u5_mult_87_n2, u5_mult_87_SUMB_43__18_, u5_mult_87_SUMB_43__19_,
         u5_mult_87_SUMB_43__20_, u5_mult_87_SUMB_43__21_,
         u5_mult_87_SUMB_43__22_, u5_mult_87_SUMB_43__23_,
         u5_mult_87_SUMB_43__24_, u5_mult_87_SUMB_43__25_,
         u5_mult_87_SUMB_43__26_, u5_mult_87_SUMB_43__27_,
         u5_mult_87_SUMB_43__28_, u5_mult_87_SUMB_43__29_,
         u5_mult_87_SUMB_43__30_, u5_mult_87_SUMB_43__31_,
         u5_mult_87_SUMB_43__32_, u5_mult_87_SUMB_43__33_,
         u5_mult_87_SUMB_43__34_, u5_mult_87_SUMB_43__35_,
         u5_mult_87_SUMB_43__36_, u5_mult_87_SUMB_43__37_,
         u5_mult_87_SUMB_43__38_, u5_mult_87_SUMB_43__39_,
         u5_mult_87_SUMB_43__40_, u5_mult_87_SUMB_43__41_,
         u5_mult_87_SUMB_43__42_, u5_mult_87_SUMB_43__43_,
         u5_mult_87_SUMB_43__44_, u5_mult_87_SUMB_43__45_,
         u5_mult_87_SUMB_43__46_, u5_mult_87_SUMB_43__47_,
         u5_mult_87_SUMB_43__48_, u5_mult_87_SUMB_43__49_,
         u5_mult_87_SUMB_43__50_, u5_mult_87_SUMB_43__51_,
         u5_mult_87_SUMB_44__1_, u5_mult_87_SUMB_44__2_,
         u5_mult_87_SUMB_44__3_, u5_mult_87_SUMB_44__4_,
         u5_mult_87_SUMB_44__5_, u5_mult_87_SUMB_44__6_,
         u5_mult_87_SUMB_44__7_, u5_mult_87_SUMB_44__8_,
         u5_mult_87_SUMB_44__9_, u5_mult_87_SUMB_44__10_,
         u5_mult_87_SUMB_44__11_, u5_mult_87_SUMB_44__12_,
         u5_mult_87_SUMB_44__13_, u5_mult_87_SUMB_44__14_,
         u5_mult_87_SUMB_44__15_, u5_mult_87_SUMB_44__16_,
         u5_mult_87_SUMB_44__17_, u5_mult_87_SUMB_44__18_,
         u5_mult_87_SUMB_44__19_, u5_mult_87_SUMB_44__20_,
         u5_mult_87_SUMB_44__21_, u5_mult_87_SUMB_44__22_,
         u5_mult_87_SUMB_44__23_, u5_mult_87_SUMB_44__24_,
         u5_mult_87_SUMB_44__25_, u5_mult_87_SUMB_44__26_,
         u5_mult_87_SUMB_44__27_, u5_mult_87_SUMB_44__28_,
         u5_mult_87_SUMB_44__29_, u5_mult_87_SUMB_44__30_,
         u5_mult_87_SUMB_44__31_, u5_mult_87_SUMB_44__32_,
         u5_mult_87_SUMB_44__33_, u5_mult_87_SUMB_44__34_,
         u5_mult_87_SUMB_44__35_, u5_mult_87_SUMB_44__36_,
         u5_mult_87_SUMB_44__37_, u5_mult_87_SUMB_44__38_,
         u5_mult_87_SUMB_44__39_, u5_mult_87_SUMB_44__40_,
         u5_mult_87_SUMB_44__41_, u5_mult_87_SUMB_44__42_,
         u5_mult_87_SUMB_44__43_, u5_mult_87_SUMB_44__44_,
         u5_mult_87_SUMB_44__45_, u5_mult_87_SUMB_44__46_,
         u5_mult_87_SUMB_44__47_, u5_mult_87_SUMB_44__48_,
         u5_mult_87_SUMB_44__49_, u5_mult_87_SUMB_44__50_,
         u5_mult_87_SUMB_44__51_, u5_mult_87_SUMB_45__1_,
         u5_mult_87_SUMB_45__2_, u5_mult_87_SUMB_45__3_,
         u5_mult_87_SUMB_45__4_, u5_mult_87_SUMB_45__5_,
         u5_mult_87_SUMB_45__6_, u5_mult_87_SUMB_45__7_,
         u5_mult_87_SUMB_45__8_, u5_mult_87_SUMB_45__9_,
         u5_mult_87_SUMB_45__10_, u5_mult_87_SUMB_45__11_,
         u5_mult_87_SUMB_45__12_, u5_mult_87_SUMB_45__13_,
         u5_mult_87_SUMB_45__14_, u5_mult_87_SUMB_45__15_,
         u5_mult_87_SUMB_45__16_, u5_mult_87_SUMB_45__17_,
         u5_mult_87_SUMB_45__18_, u5_mult_87_SUMB_45__19_,
         u5_mult_87_SUMB_45__20_, u5_mult_87_SUMB_45__21_,
         u5_mult_87_SUMB_45__22_, u5_mult_87_SUMB_45__23_,
         u5_mult_87_SUMB_45__24_, u5_mult_87_SUMB_45__25_,
         u5_mult_87_SUMB_45__26_, u5_mult_87_SUMB_45__27_,
         u5_mult_87_SUMB_45__28_, u5_mult_87_SUMB_45__29_,
         u5_mult_87_SUMB_45__30_, u5_mult_87_SUMB_45__31_,
         u5_mult_87_SUMB_45__32_, u5_mult_87_SUMB_45__33_,
         u5_mult_87_SUMB_45__34_, u5_mult_87_SUMB_45__35_,
         u5_mult_87_SUMB_45__36_, u5_mult_87_SUMB_45__37_,
         u5_mult_87_SUMB_45__38_, u5_mult_87_SUMB_45__39_,
         u5_mult_87_SUMB_45__40_, u5_mult_87_SUMB_45__41_,
         u5_mult_87_SUMB_45__42_, u5_mult_87_SUMB_45__43_,
         u5_mult_87_SUMB_45__44_, u5_mult_87_SUMB_45__45_,
         u5_mult_87_SUMB_45__46_, u5_mult_87_SUMB_45__47_,
         u5_mult_87_SUMB_45__48_, u5_mult_87_SUMB_45__49_,
         u5_mult_87_SUMB_45__50_, u5_mult_87_SUMB_45__51_,
         u5_mult_87_SUMB_46__1_, u5_mult_87_SUMB_46__2_,
         u5_mult_87_SUMB_46__3_, u5_mult_87_SUMB_46__4_,
         u5_mult_87_SUMB_46__5_, u5_mult_87_SUMB_46__6_,
         u5_mult_87_SUMB_46__7_, u5_mult_87_SUMB_46__8_,
         u5_mult_87_SUMB_46__9_, u5_mult_87_SUMB_46__10_,
         u5_mult_87_SUMB_46__11_, u5_mult_87_SUMB_46__12_,
         u5_mult_87_SUMB_46__13_, u5_mult_87_SUMB_46__14_,
         u5_mult_87_SUMB_46__15_, u5_mult_87_SUMB_46__16_,
         u5_mult_87_SUMB_46__17_, u5_mult_87_SUMB_46__18_,
         u5_mult_87_SUMB_46__19_, u5_mult_87_SUMB_46__20_,
         u5_mult_87_SUMB_46__21_, u5_mult_87_SUMB_46__22_,
         u5_mult_87_SUMB_46__23_, u5_mult_87_SUMB_46__24_,
         u5_mult_87_SUMB_46__25_, u5_mult_87_SUMB_46__26_,
         u5_mult_87_SUMB_46__27_, u5_mult_87_SUMB_46__28_,
         u5_mult_87_SUMB_46__29_, u5_mult_87_SUMB_46__30_,
         u5_mult_87_SUMB_46__31_, u5_mult_87_SUMB_46__32_,
         u5_mult_87_SUMB_46__33_, u5_mult_87_SUMB_46__34_,
         u5_mult_87_SUMB_46__35_, u5_mult_87_SUMB_46__36_,
         u5_mult_87_SUMB_46__37_, u5_mult_87_SUMB_46__38_,
         u5_mult_87_SUMB_46__39_, u5_mult_87_SUMB_46__40_,
         u5_mult_87_SUMB_46__41_, u5_mult_87_SUMB_46__42_,
         u5_mult_87_SUMB_46__43_, u5_mult_87_SUMB_46__44_,
         u5_mult_87_SUMB_46__45_, u5_mult_87_SUMB_46__46_,
         u5_mult_87_SUMB_46__47_, u5_mult_87_SUMB_46__48_,
         u5_mult_87_SUMB_46__49_, u5_mult_87_SUMB_46__50_,
         u5_mult_87_SUMB_46__51_, u5_mult_87_SUMB_47__1_,
         u5_mult_87_SUMB_47__2_, u5_mult_87_SUMB_47__3_,
         u5_mult_87_SUMB_47__4_, u5_mult_87_SUMB_47__5_,
         u5_mult_87_SUMB_47__6_, u5_mult_87_SUMB_47__7_,
         u5_mult_87_SUMB_47__8_, u5_mult_87_SUMB_47__9_,
         u5_mult_87_SUMB_47__10_, u5_mult_87_SUMB_47__11_,
         u5_mult_87_SUMB_47__12_, u5_mult_87_SUMB_47__13_,
         u5_mult_87_SUMB_47__14_, u5_mult_87_SUMB_47__15_,
         u5_mult_87_SUMB_47__16_, u5_mult_87_SUMB_47__17_,
         u5_mult_87_SUMB_47__18_, u5_mult_87_SUMB_47__19_,
         u5_mult_87_SUMB_47__20_, u5_mult_87_SUMB_47__21_,
         u5_mult_87_SUMB_47__22_, u5_mult_87_SUMB_47__23_,
         u5_mult_87_SUMB_47__24_, u5_mult_87_SUMB_47__25_,
         u5_mult_87_SUMB_47__26_, u5_mult_87_SUMB_47__27_,
         u5_mult_87_SUMB_47__28_, u5_mult_87_SUMB_47__29_,
         u5_mult_87_SUMB_47__30_, u5_mult_87_SUMB_47__31_,
         u5_mult_87_SUMB_47__32_, u5_mult_87_SUMB_47__33_,
         u5_mult_87_SUMB_47__34_, u5_mult_87_SUMB_47__35_,
         u5_mult_87_SUMB_47__36_, u5_mult_87_SUMB_47__37_,
         u5_mult_87_SUMB_47__38_, u5_mult_87_SUMB_47__39_,
         u5_mult_87_SUMB_47__40_, u5_mult_87_SUMB_47__41_,
         u5_mult_87_SUMB_47__42_, u5_mult_87_SUMB_47__43_,
         u5_mult_87_SUMB_47__44_, u5_mult_87_SUMB_47__45_,
         u5_mult_87_SUMB_47__46_, u5_mult_87_SUMB_47__47_,
         u5_mult_87_SUMB_47__48_, u5_mult_87_SUMB_47__49_,
         u5_mult_87_SUMB_47__50_, u5_mult_87_SUMB_47__51_,
         u5_mult_87_SUMB_48__1_, u5_mult_87_SUMB_48__2_,
         u5_mult_87_SUMB_48__3_, u5_mult_87_SUMB_48__4_,
         u5_mult_87_SUMB_48__5_, u5_mult_87_SUMB_48__6_,
         u5_mult_87_SUMB_48__7_, u5_mult_87_SUMB_48__8_,
         u5_mult_87_SUMB_48__9_, u5_mult_87_SUMB_48__10_,
         u5_mult_87_SUMB_48__11_, u5_mult_87_SUMB_48__12_,
         u5_mult_87_SUMB_48__13_, u5_mult_87_SUMB_48__14_,
         u5_mult_87_SUMB_48__15_, u5_mult_87_SUMB_48__16_,
         u5_mult_87_SUMB_48__17_, u5_mult_87_SUMB_48__18_,
         u5_mult_87_SUMB_48__19_, u5_mult_87_SUMB_48__20_,
         u5_mult_87_SUMB_48__21_, u5_mult_87_SUMB_48__22_,
         u5_mult_87_SUMB_48__23_, u5_mult_87_SUMB_48__24_,
         u5_mult_87_SUMB_48__25_, u5_mult_87_SUMB_48__26_,
         u5_mult_87_SUMB_48__27_, u5_mult_87_SUMB_48__28_,
         u5_mult_87_SUMB_48__29_, u5_mult_87_SUMB_48__30_,
         u5_mult_87_SUMB_48__31_, u5_mult_87_SUMB_48__32_,
         u5_mult_87_SUMB_48__33_, u5_mult_87_SUMB_48__34_,
         u5_mult_87_SUMB_48__35_, u5_mult_87_SUMB_48__36_,
         u5_mult_87_SUMB_48__37_, u5_mult_87_SUMB_48__38_,
         u5_mult_87_SUMB_48__39_, u5_mult_87_SUMB_48__40_,
         u5_mult_87_SUMB_48__41_, u5_mult_87_SUMB_48__42_,
         u5_mult_87_SUMB_48__43_, u5_mult_87_SUMB_48__44_,
         u5_mult_87_SUMB_48__45_, u5_mult_87_SUMB_48__46_,
         u5_mult_87_SUMB_48__47_, u5_mult_87_SUMB_48__48_,
         u5_mult_87_SUMB_48__49_, u5_mult_87_SUMB_48__50_,
         u5_mult_87_SUMB_48__51_, u5_mult_87_SUMB_49__1_,
         u5_mult_87_SUMB_49__2_, u5_mult_87_SUMB_49__3_,
         u5_mult_87_SUMB_49__4_, u5_mult_87_SUMB_49__5_,
         u5_mult_87_SUMB_49__6_, u5_mult_87_SUMB_49__7_,
         u5_mult_87_SUMB_49__8_, u5_mult_87_SUMB_49__9_,
         u5_mult_87_SUMB_49__10_, u5_mult_87_SUMB_49__11_,
         u5_mult_87_SUMB_49__12_, u5_mult_87_SUMB_49__13_,
         u5_mult_87_SUMB_49__14_, u5_mult_87_SUMB_49__15_,
         u5_mult_87_SUMB_49__16_, u5_mult_87_SUMB_49__17_,
         u5_mult_87_SUMB_49__18_, u5_mult_87_SUMB_49__19_,
         u5_mult_87_SUMB_49__20_, u5_mult_87_SUMB_49__21_,
         u5_mult_87_SUMB_49__22_, u5_mult_87_SUMB_49__23_,
         u5_mult_87_SUMB_49__24_, u5_mult_87_SUMB_49__25_,
         u5_mult_87_SUMB_49__26_, u5_mult_87_SUMB_49__27_,
         u5_mult_87_SUMB_49__28_, u5_mult_87_SUMB_49__29_,
         u5_mult_87_SUMB_49__30_, u5_mult_87_SUMB_49__31_,
         u5_mult_87_SUMB_49__32_, u5_mult_87_SUMB_49__33_,
         u5_mult_87_SUMB_49__34_, u5_mult_87_SUMB_49__35_,
         u5_mult_87_SUMB_49__36_, u5_mult_87_SUMB_49__37_,
         u5_mult_87_SUMB_49__38_, u5_mult_87_SUMB_49__39_,
         u5_mult_87_SUMB_49__40_, u5_mult_87_SUMB_49__41_,
         u5_mult_87_SUMB_49__42_, u5_mult_87_SUMB_49__43_,
         u5_mult_87_SUMB_49__44_, u5_mult_87_SUMB_49__45_,
         u5_mult_87_SUMB_49__46_, u5_mult_87_SUMB_49__47_,
         u5_mult_87_SUMB_49__48_, u5_mult_87_SUMB_49__49_,
         u5_mult_87_SUMB_49__50_, u5_mult_87_SUMB_49__51_,
         u5_mult_87_SUMB_50__1_, u5_mult_87_SUMB_50__2_,
         u5_mult_87_SUMB_50__3_, u5_mult_87_SUMB_50__4_,
         u5_mult_87_SUMB_50__5_, u5_mult_87_SUMB_50__6_,
         u5_mult_87_SUMB_50__7_, u5_mult_87_SUMB_50__8_,
         u5_mult_87_SUMB_50__9_, u5_mult_87_SUMB_50__10_,
         u5_mult_87_SUMB_50__11_, u5_mult_87_SUMB_50__12_,
         u5_mult_87_SUMB_50__13_, u5_mult_87_SUMB_50__14_,
         u5_mult_87_SUMB_50__15_, u5_mult_87_SUMB_50__16_,
         u5_mult_87_SUMB_50__17_, u5_mult_87_SUMB_50__18_,
         u5_mult_87_SUMB_50__19_, u5_mult_87_SUMB_50__20_,
         u5_mult_87_SUMB_50__21_, u5_mult_87_SUMB_50__22_,
         u5_mult_87_SUMB_50__23_, u5_mult_87_SUMB_50__24_,
         u5_mult_87_SUMB_50__25_, u5_mult_87_SUMB_50__26_,
         u5_mult_87_SUMB_50__27_, u5_mult_87_SUMB_50__28_,
         u5_mult_87_SUMB_50__29_, u5_mult_87_SUMB_50__30_,
         u5_mult_87_SUMB_50__31_, u5_mult_87_SUMB_50__32_,
         u5_mult_87_SUMB_50__33_, u5_mult_87_SUMB_50__34_,
         u5_mult_87_SUMB_50__35_, u5_mult_87_SUMB_50__36_,
         u5_mult_87_SUMB_50__37_, u5_mult_87_SUMB_50__38_,
         u5_mult_87_SUMB_50__39_, u5_mult_87_SUMB_50__40_,
         u5_mult_87_SUMB_50__41_, u5_mult_87_SUMB_50__42_,
         u5_mult_87_SUMB_50__43_, u5_mult_87_SUMB_50__44_,
         u5_mult_87_SUMB_50__45_, u5_mult_87_SUMB_50__46_,
         u5_mult_87_SUMB_50__47_, u5_mult_87_SUMB_50__48_,
         u5_mult_87_SUMB_50__49_, u5_mult_87_SUMB_50__50_,
         u5_mult_87_SUMB_50__51_, u5_mult_87_SUMB_51__1_,
         u5_mult_87_SUMB_51__2_, u5_mult_87_SUMB_51__3_,
         u5_mult_87_SUMB_51__4_, u5_mult_87_SUMB_51__5_,
         u5_mult_87_SUMB_51__6_, u5_mult_87_SUMB_51__7_,
         u5_mult_87_SUMB_51__8_, u5_mult_87_SUMB_51__9_,
         u5_mult_87_SUMB_51__10_, u5_mult_87_SUMB_51__11_,
         u5_mult_87_SUMB_51__12_, u5_mult_87_SUMB_51__13_,
         u5_mult_87_SUMB_51__14_, u5_mult_87_SUMB_51__15_,
         u5_mult_87_SUMB_51__16_, u5_mult_87_SUMB_51__17_,
         u5_mult_87_SUMB_51__18_, u5_mult_87_SUMB_51__19_,
         u5_mult_87_SUMB_51__20_, u5_mult_87_SUMB_51__21_,
         u5_mult_87_SUMB_51__22_, u5_mult_87_SUMB_51__23_,
         u5_mult_87_SUMB_51__24_, u5_mult_87_SUMB_51__25_,
         u5_mult_87_SUMB_51__26_, u5_mult_87_SUMB_51__27_,
         u5_mult_87_SUMB_51__28_, u5_mult_87_SUMB_51__29_,
         u5_mult_87_SUMB_51__30_, u5_mult_87_SUMB_51__31_,
         u5_mult_87_SUMB_51__32_, u5_mult_87_SUMB_51__33_,
         u5_mult_87_SUMB_51__34_, u5_mult_87_SUMB_51__35_,
         u5_mult_87_SUMB_51__36_, u5_mult_87_SUMB_51__37_,
         u5_mult_87_SUMB_51__38_, u5_mult_87_SUMB_51__39_,
         u5_mult_87_SUMB_51__40_, u5_mult_87_SUMB_51__41_,
         u5_mult_87_SUMB_51__42_, u5_mult_87_SUMB_51__43_,
         u5_mult_87_SUMB_51__44_, u5_mult_87_SUMB_51__45_,
         u5_mult_87_SUMB_51__46_, u5_mult_87_SUMB_51__47_,
         u5_mult_87_SUMB_51__48_, u5_mult_87_SUMB_51__49_,
         u5_mult_87_SUMB_51__50_, u5_mult_87_SUMB_51__51_,
         u5_mult_87_SUMB_52__1_, u5_mult_87_SUMB_52__2_,
         u5_mult_87_SUMB_52__3_, u5_mult_87_SUMB_52__4_,
         u5_mult_87_SUMB_52__5_, u5_mult_87_SUMB_52__6_,
         u5_mult_87_SUMB_52__7_, u5_mult_87_SUMB_52__8_,
         u5_mult_87_SUMB_52__9_, u5_mult_87_SUMB_52__10_,
         u5_mult_87_SUMB_52__11_, u5_mult_87_SUMB_52__12_,
         u5_mult_87_SUMB_52__13_, u5_mult_87_SUMB_52__14_,
         u5_mult_87_SUMB_52__15_, u5_mult_87_SUMB_52__16_,
         u5_mult_87_SUMB_52__17_, u5_mult_87_SUMB_52__18_,
         u5_mult_87_SUMB_52__19_, u5_mult_87_SUMB_52__20_,
         u5_mult_87_SUMB_52__21_, u5_mult_87_SUMB_52__22_,
         u5_mult_87_SUMB_52__23_, u5_mult_87_SUMB_52__24_,
         u5_mult_87_SUMB_52__25_, u5_mult_87_SUMB_52__26_,
         u5_mult_87_SUMB_52__27_, u5_mult_87_SUMB_52__28_,
         u5_mult_87_SUMB_52__29_, u5_mult_87_SUMB_52__30_,
         u5_mult_87_SUMB_52__31_, u5_mult_87_SUMB_52__32_,
         u5_mult_87_SUMB_52__33_, u5_mult_87_SUMB_52__34_,
         u5_mult_87_SUMB_52__35_, u5_mult_87_SUMB_52__36_,
         u5_mult_87_SUMB_52__37_, u5_mult_87_SUMB_52__38_,
         u5_mult_87_SUMB_52__39_, u5_mult_87_SUMB_52__40_,
         u5_mult_87_SUMB_52__41_, u5_mult_87_SUMB_52__42_,
         u5_mult_87_SUMB_52__43_, u5_mult_87_SUMB_52__44_,
         u5_mult_87_SUMB_52__45_, u5_mult_87_SUMB_52__46_,
         u5_mult_87_SUMB_52__47_, u5_mult_87_SUMB_52__48_,
         u5_mult_87_SUMB_52__49_, u5_mult_87_SUMB_52__50_,
         u5_mult_87_SUMB_52__51_, u5_mult_87_CARRYB_43__18_,
         u5_mult_87_CARRYB_43__19_, u5_mult_87_CARRYB_43__20_,
         u5_mult_87_CARRYB_43__21_, u5_mult_87_CARRYB_43__22_,
         u5_mult_87_CARRYB_43__23_, u5_mult_87_CARRYB_43__24_,
         u5_mult_87_CARRYB_43__25_, u5_mult_87_CARRYB_43__26_,
         u5_mult_87_CARRYB_43__27_, u5_mult_87_CARRYB_43__28_,
         u5_mult_87_CARRYB_43__29_, u5_mult_87_CARRYB_43__30_,
         u5_mult_87_CARRYB_43__31_, u5_mult_87_CARRYB_43__32_,
         u5_mult_87_CARRYB_43__33_, u5_mult_87_CARRYB_43__34_,
         u5_mult_87_CARRYB_43__35_, u5_mult_87_CARRYB_43__36_,
         u5_mult_87_CARRYB_43__37_, u5_mult_87_CARRYB_43__38_,
         u5_mult_87_CARRYB_43__39_, u5_mult_87_CARRYB_43__40_,
         u5_mult_87_CARRYB_43__41_, u5_mult_87_CARRYB_43__42_,
         u5_mult_87_CARRYB_43__43_, u5_mult_87_CARRYB_43__44_,
         u5_mult_87_CARRYB_43__45_, u5_mult_87_CARRYB_43__46_,
         u5_mult_87_CARRYB_43__47_, u5_mult_87_CARRYB_43__48_,
         u5_mult_87_CARRYB_43__49_, u5_mult_87_CARRYB_43__50_,
         u5_mult_87_CARRYB_43__51_, u5_mult_87_CARRYB_44__0_,
         u5_mult_87_CARRYB_44__1_, u5_mult_87_CARRYB_44__2_,
         u5_mult_87_CARRYB_44__3_, u5_mult_87_CARRYB_44__4_,
         u5_mult_87_CARRYB_44__5_, u5_mult_87_CARRYB_44__6_,
         u5_mult_87_CARRYB_44__7_, u5_mult_87_CARRYB_44__8_,
         u5_mult_87_CARRYB_44__9_, u5_mult_87_CARRYB_44__10_,
         u5_mult_87_CARRYB_44__11_, u5_mult_87_CARRYB_44__12_,
         u5_mult_87_CARRYB_44__13_, u5_mult_87_CARRYB_44__14_,
         u5_mult_87_CARRYB_44__15_, u5_mult_87_CARRYB_44__16_,
         u5_mult_87_CARRYB_44__17_, u5_mult_87_CARRYB_44__18_,
         u5_mult_87_CARRYB_44__19_, u5_mult_87_CARRYB_44__20_,
         u5_mult_87_CARRYB_44__21_, u5_mult_87_CARRYB_44__22_,
         u5_mult_87_CARRYB_44__23_, u5_mult_87_CARRYB_44__24_,
         u5_mult_87_CARRYB_44__25_, u5_mult_87_CARRYB_44__26_,
         u5_mult_87_CARRYB_44__27_, u5_mult_87_CARRYB_44__28_,
         u5_mult_87_CARRYB_44__29_, u5_mult_87_CARRYB_44__30_,
         u5_mult_87_CARRYB_44__31_, u5_mult_87_CARRYB_44__32_,
         u5_mult_87_CARRYB_44__33_, u5_mult_87_CARRYB_44__34_,
         u5_mult_87_CARRYB_44__35_, u5_mult_87_CARRYB_44__36_,
         u5_mult_87_CARRYB_44__37_, u5_mult_87_CARRYB_44__38_,
         u5_mult_87_CARRYB_44__39_, u5_mult_87_CARRYB_44__40_,
         u5_mult_87_CARRYB_44__41_, u5_mult_87_CARRYB_44__42_,
         u5_mult_87_CARRYB_44__43_, u5_mult_87_CARRYB_44__44_,
         u5_mult_87_CARRYB_44__45_, u5_mult_87_CARRYB_44__46_,
         u5_mult_87_CARRYB_44__47_, u5_mult_87_CARRYB_44__48_,
         u5_mult_87_CARRYB_44__49_, u5_mult_87_CARRYB_44__50_,
         u5_mult_87_CARRYB_44__51_, u5_mult_87_CARRYB_45__0_,
         u5_mult_87_CARRYB_45__1_, u5_mult_87_CARRYB_45__2_,
         u5_mult_87_CARRYB_45__3_, u5_mult_87_CARRYB_45__4_,
         u5_mult_87_CARRYB_45__5_, u5_mult_87_CARRYB_45__6_,
         u5_mult_87_CARRYB_45__7_, u5_mult_87_CARRYB_45__8_,
         u5_mult_87_CARRYB_45__9_, u5_mult_87_CARRYB_45__10_,
         u5_mult_87_CARRYB_45__11_, u5_mult_87_CARRYB_45__12_,
         u5_mult_87_CARRYB_45__13_, u5_mult_87_CARRYB_45__14_,
         u5_mult_87_CARRYB_45__15_, u5_mult_87_CARRYB_45__16_,
         u5_mult_87_CARRYB_45__17_, u5_mult_87_CARRYB_45__18_,
         u5_mult_87_CARRYB_45__19_, u5_mult_87_CARRYB_45__20_,
         u5_mult_87_CARRYB_45__21_, u5_mult_87_CARRYB_45__22_,
         u5_mult_87_CARRYB_45__23_, u5_mult_87_CARRYB_45__24_,
         u5_mult_87_CARRYB_45__25_, u5_mult_87_CARRYB_45__26_,
         u5_mult_87_CARRYB_45__27_, u5_mult_87_CARRYB_45__28_,
         u5_mult_87_CARRYB_45__29_, u5_mult_87_CARRYB_45__30_,
         u5_mult_87_CARRYB_45__31_, u5_mult_87_CARRYB_45__32_,
         u5_mult_87_CARRYB_45__33_, u5_mult_87_CARRYB_45__34_,
         u5_mult_87_CARRYB_45__35_, u5_mult_87_CARRYB_45__36_,
         u5_mult_87_CARRYB_45__37_, u5_mult_87_CARRYB_45__38_,
         u5_mult_87_CARRYB_45__39_, u5_mult_87_CARRYB_45__40_,
         u5_mult_87_CARRYB_45__41_, u5_mult_87_CARRYB_45__42_,
         u5_mult_87_CARRYB_45__43_, u5_mult_87_CARRYB_45__44_,
         u5_mult_87_CARRYB_45__45_, u5_mult_87_CARRYB_45__46_,
         u5_mult_87_CARRYB_45__47_, u5_mult_87_CARRYB_45__48_,
         u5_mult_87_CARRYB_45__49_, u5_mult_87_CARRYB_45__50_,
         u5_mult_87_CARRYB_45__51_, u5_mult_87_CARRYB_46__0_,
         u5_mult_87_CARRYB_46__1_, u5_mult_87_CARRYB_46__2_,
         u5_mult_87_CARRYB_46__3_, u5_mult_87_CARRYB_46__4_,
         u5_mult_87_CARRYB_46__5_, u5_mult_87_CARRYB_46__6_,
         u5_mult_87_CARRYB_46__7_, u5_mult_87_CARRYB_46__8_,
         u5_mult_87_CARRYB_46__9_, u5_mult_87_CARRYB_46__10_,
         u5_mult_87_CARRYB_46__11_, u5_mult_87_CARRYB_46__12_,
         u5_mult_87_CARRYB_46__13_, u5_mult_87_CARRYB_46__14_,
         u5_mult_87_CARRYB_46__15_, u5_mult_87_CARRYB_46__16_,
         u5_mult_87_CARRYB_46__17_, u5_mult_87_CARRYB_46__18_,
         u5_mult_87_CARRYB_46__19_, u5_mult_87_CARRYB_46__20_,
         u5_mult_87_CARRYB_46__21_, u5_mult_87_CARRYB_46__22_,
         u5_mult_87_CARRYB_46__23_, u5_mult_87_CARRYB_46__24_,
         u5_mult_87_CARRYB_46__25_, u5_mult_87_CARRYB_46__26_,
         u5_mult_87_CARRYB_46__27_, u5_mult_87_CARRYB_46__28_,
         u5_mult_87_CARRYB_46__29_, u5_mult_87_CARRYB_46__30_,
         u5_mult_87_CARRYB_46__31_, u5_mult_87_CARRYB_46__32_,
         u5_mult_87_CARRYB_46__33_, u5_mult_87_CARRYB_46__34_,
         u5_mult_87_CARRYB_46__35_, u5_mult_87_CARRYB_46__36_,
         u5_mult_87_CARRYB_46__37_, u5_mult_87_CARRYB_46__38_,
         u5_mult_87_CARRYB_46__39_, u5_mult_87_CARRYB_46__40_,
         u5_mult_87_CARRYB_46__41_, u5_mult_87_CARRYB_46__42_,
         u5_mult_87_CARRYB_46__43_, u5_mult_87_CARRYB_46__44_,
         u5_mult_87_CARRYB_46__45_, u5_mult_87_CARRYB_46__46_,
         u5_mult_87_CARRYB_46__47_, u5_mult_87_CARRYB_46__48_,
         u5_mult_87_CARRYB_46__49_, u5_mult_87_CARRYB_46__50_,
         u5_mult_87_CARRYB_46__51_, u5_mult_87_CARRYB_47__0_,
         u5_mult_87_CARRYB_47__1_, u5_mult_87_CARRYB_47__2_,
         u5_mult_87_CARRYB_47__3_, u5_mult_87_CARRYB_47__4_,
         u5_mult_87_CARRYB_47__5_, u5_mult_87_CARRYB_47__6_,
         u5_mult_87_CARRYB_47__7_, u5_mult_87_CARRYB_47__8_,
         u5_mult_87_CARRYB_47__9_, u5_mult_87_CARRYB_47__10_,
         u5_mult_87_CARRYB_47__11_, u5_mult_87_CARRYB_47__12_,
         u5_mult_87_CARRYB_47__13_, u5_mult_87_CARRYB_47__14_,
         u5_mult_87_CARRYB_47__15_, u5_mult_87_CARRYB_47__16_,
         u5_mult_87_CARRYB_47__17_, u5_mult_87_CARRYB_47__18_,
         u5_mult_87_CARRYB_47__19_, u5_mult_87_CARRYB_47__20_,
         u5_mult_87_CARRYB_47__21_, u5_mult_87_CARRYB_47__22_,
         u5_mult_87_CARRYB_47__23_, u5_mult_87_CARRYB_47__24_,
         u5_mult_87_CARRYB_47__25_, u5_mult_87_CARRYB_47__26_,
         u5_mult_87_CARRYB_47__27_, u5_mult_87_CARRYB_47__28_,
         u5_mult_87_CARRYB_47__29_, u5_mult_87_CARRYB_47__30_,
         u5_mult_87_CARRYB_47__31_, u5_mult_87_CARRYB_47__32_,
         u5_mult_87_CARRYB_47__33_, u5_mult_87_CARRYB_47__34_,
         u5_mult_87_CARRYB_47__35_, u5_mult_87_CARRYB_47__36_,
         u5_mult_87_CARRYB_47__37_, u5_mult_87_CARRYB_47__38_,
         u5_mult_87_CARRYB_47__39_, u5_mult_87_CARRYB_47__40_,
         u5_mult_87_CARRYB_47__41_, u5_mult_87_CARRYB_47__42_,
         u5_mult_87_CARRYB_47__43_, u5_mult_87_CARRYB_47__44_,
         u5_mult_87_CARRYB_47__45_, u5_mult_87_CARRYB_47__46_,
         u5_mult_87_CARRYB_47__47_, u5_mult_87_CARRYB_47__48_,
         u5_mult_87_CARRYB_47__49_, u5_mult_87_CARRYB_47__50_,
         u5_mult_87_CARRYB_47__51_, u5_mult_87_CARRYB_48__0_,
         u5_mult_87_CARRYB_48__1_, u5_mult_87_CARRYB_48__2_,
         u5_mult_87_CARRYB_48__3_, u5_mult_87_CARRYB_48__4_,
         u5_mult_87_CARRYB_48__5_, u5_mult_87_CARRYB_48__6_,
         u5_mult_87_CARRYB_48__7_, u5_mult_87_CARRYB_48__8_,
         u5_mult_87_CARRYB_48__9_, u5_mult_87_CARRYB_48__10_,
         u5_mult_87_CARRYB_48__11_, u5_mult_87_CARRYB_48__12_,
         u5_mult_87_CARRYB_48__13_, u5_mult_87_CARRYB_48__14_,
         u5_mult_87_CARRYB_48__15_, u5_mult_87_CARRYB_48__16_,
         u5_mult_87_CARRYB_48__17_, u5_mult_87_CARRYB_48__18_,
         u5_mult_87_CARRYB_48__19_, u5_mult_87_CARRYB_48__20_,
         u5_mult_87_CARRYB_48__21_, u5_mult_87_CARRYB_48__22_,
         u5_mult_87_CARRYB_48__23_, u5_mult_87_CARRYB_48__24_,
         u5_mult_87_CARRYB_48__25_, u5_mult_87_CARRYB_48__26_,
         u5_mult_87_CARRYB_48__27_, u5_mult_87_CARRYB_48__28_,
         u5_mult_87_CARRYB_48__29_, u5_mult_87_CARRYB_48__30_,
         u5_mult_87_CARRYB_48__31_, u5_mult_87_CARRYB_48__32_,
         u5_mult_87_CARRYB_48__33_, u5_mult_87_CARRYB_48__34_,
         u5_mult_87_CARRYB_48__35_, u5_mult_87_CARRYB_48__36_,
         u5_mult_87_CARRYB_48__37_, u5_mult_87_CARRYB_48__38_,
         u5_mult_87_CARRYB_48__39_, u5_mult_87_CARRYB_48__40_,
         u5_mult_87_CARRYB_48__41_, u5_mult_87_CARRYB_48__42_,
         u5_mult_87_CARRYB_48__43_, u5_mult_87_CARRYB_48__44_,
         u5_mult_87_CARRYB_48__45_, u5_mult_87_CARRYB_48__46_,
         u5_mult_87_CARRYB_48__47_, u5_mult_87_CARRYB_48__48_,
         u5_mult_87_CARRYB_48__49_, u5_mult_87_CARRYB_48__50_,
         u5_mult_87_CARRYB_48__51_, u5_mult_87_CARRYB_49__0_,
         u5_mult_87_CARRYB_49__1_, u5_mult_87_CARRYB_49__2_,
         u5_mult_87_CARRYB_49__3_, u5_mult_87_CARRYB_49__4_,
         u5_mult_87_CARRYB_49__5_, u5_mult_87_CARRYB_49__6_,
         u5_mult_87_CARRYB_49__7_, u5_mult_87_CARRYB_49__8_,
         u5_mult_87_CARRYB_49__9_, u5_mult_87_CARRYB_49__10_,
         u5_mult_87_CARRYB_49__11_, u5_mult_87_CARRYB_49__12_,
         u5_mult_87_CARRYB_49__13_, u5_mult_87_CARRYB_49__14_,
         u5_mult_87_CARRYB_49__15_, u5_mult_87_CARRYB_49__16_,
         u5_mult_87_CARRYB_49__17_, u5_mult_87_CARRYB_49__18_,
         u5_mult_87_CARRYB_49__19_, u5_mult_87_CARRYB_49__20_,
         u5_mult_87_CARRYB_49__21_, u5_mult_87_CARRYB_49__22_,
         u5_mult_87_CARRYB_49__23_, u5_mult_87_CARRYB_49__24_,
         u5_mult_87_CARRYB_49__25_, u5_mult_87_CARRYB_49__26_,
         u5_mult_87_CARRYB_49__27_, u5_mult_87_CARRYB_49__28_,
         u5_mult_87_CARRYB_49__29_, u5_mult_87_CARRYB_49__30_,
         u5_mult_87_CARRYB_49__31_, u5_mult_87_CARRYB_49__32_,
         u5_mult_87_CARRYB_49__33_, u5_mult_87_CARRYB_49__34_,
         u5_mult_87_CARRYB_49__35_, u5_mult_87_CARRYB_49__36_,
         u5_mult_87_CARRYB_49__37_, u5_mult_87_CARRYB_49__38_,
         u5_mult_87_CARRYB_49__39_, u5_mult_87_CARRYB_49__40_,
         u5_mult_87_CARRYB_49__41_, u5_mult_87_CARRYB_49__42_,
         u5_mult_87_CARRYB_49__43_, u5_mult_87_CARRYB_49__44_,
         u5_mult_87_CARRYB_49__45_, u5_mult_87_CARRYB_49__46_,
         u5_mult_87_CARRYB_49__47_, u5_mult_87_CARRYB_49__48_,
         u5_mult_87_CARRYB_49__49_, u5_mult_87_CARRYB_49__50_,
         u5_mult_87_CARRYB_49__51_, u5_mult_87_CARRYB_50__0_,
         u5_mult_87_CARRYB_50__1_, u5_mult_87_CARRYB_50__2_,
         u5_mult_87_CARRYB_50__3_, u5_mult_87_CARRYB_50__4_,
         u5_mult_87_CARRYB_50__5_, u5_mult_87_CARRYB_50__6_,
         u5_mult_87_CARRYB_50__7_, u5_mult_87_CARRYB_50__8_,
         u5_mult_87_CARRYB_50__9_, u5_mult_87_CARRYB_50__10_,
         u5_mult_87_CARRYB_50__11_, u5_mult_87_CARRYB_50__12_,
         u5_mult_87_CARRYB_50__13_, u5_mult_87_CARRYB_50__14_,
         u5_mult_87_CARRYB_50__15_, u5_mult_87_CARRYB_50__16_,
         u5_mult_87_CARRYB_50__17_, u5_mult_87_CARRYB_50__18_,
         u5_mult_87_CARRYB_50__19_, u5_mult_87_CARRYB_50__20_,
         u5_mult_87_CARRYB_50__21_, u5_mult_87_CARRYB_50__22_,
         u5_mult_87_CARRYB_50__23_, u5_mult_87_CARRYB_50__24_,
         u5_mult_87_CARRYB_50__25_, u5_mult_87_CARRYB_50__26_,
         u5_mult_87_CARRYB_50__27_, u5_mult_87_CARRYB_50__28_,
         u5_mult_87_CARRYB_50__29_, u5_mult_87_CARRYB_50__30_,
         u5_mult_87_CARRYB_50__31_, u5_mult_87_CARRYB_50__32_,
         u5_mult_87_CARRYB_50__33_, u5_mult_87_CARRYB_50__34_,
         u5_mult_87_CARRYB_50__35_, u5_mult_87_CARRYB_50__36_,
         u5_mult_87_CARRYB_50__37_, u5_mult_87_CARRYB_50__38_,
         u5_mult_87_CARRYB_50__39_, u5_mult_87_CARRYB_50__40_,
         u5_mult_87_CARRYB_50__41_, u5_mult_87_CARRYB_50__42_,
         u5_mult_87_CARRYB_50__43_, u5_mult_87_CARRYB_50__44_,
         u5_mult_87_CARRYB_50__45_, u5_mult_87_CARRYB_50__46_,
         u5_mult_87_CARRYB_50__47_, u5_mult_87_CARRYB_50__48_,
         u5_mult_87_CARRYB_50__49_, u5_mult_87_CARRYB_50__50_,
         u5_mult_87_CARRYB_50__51_, u5_mult_87_CARRYB_51__0_,
         u5_mult_87_CARRYB_51__1_, u5_mult_87_CARRYB_51__2_,
         u5_mult_87_CARRYB_51__3_, u5_mult_87_CARRYB_51__4_,
         u5_mult_87_CARRYB_51__5_, u5_mult_87_CARRYB_51__6_,
         u5_mult_87_CARRYB_51__7_, u5_mult_87_CARRYB_51__8_,
         u5_mult_87_CARRYB_51__9_, u5_mult_87_CARRYB_51__10_,
         u5_mult_87_CARRYB_51__11_, u5_mult_87_CARRYB_51__12_,
         u5_mult_87_CARRYB_51__13_, u5_mult_87_CARRYB_51__14_,
         u5_mult_87_CARRYB_51__15_, u5_mult_87_CARRYB_51__16_,
         u5_mult_87_CARRYB_51__17_, u5_mult_87_CARRYB_51__18_,
         u5_mult_87_CARRYB_51__19_, u5_mult_87_CARRYB_51__20_,
         u5_mult_87_CARRYB_51__21_, u5_mult_87_CARRYB_51__22_,
         u5_mult_87_CARRYB_51__23_, u5_mult_87_CARRYB_51__24_,
         u5_mult_87_CARRYB_51__25_, u5_mult_87_CARRYB_51__26_,
         u5_mult_87_CARRYB_51__27_, u5_mult_87_CARRYB_51__28_,
         u5_mult_87_CARRYB_51__29_, u5_mult_87_CARRYB_51__30_,
         u5_mult_87_CARRYB_51__31_, u5_mult_87_CARRYB_51__32_,
         u5_mult_87_CARRYB_51__33_, u5_mult_87_CARRYB_51__34_,
         u5_mult_87_CARRYB_51__35_, u5_mult_87_CARRYB_51__36_,
         u5_mult_87_CARRYB_51__37_, u5_mult_87_CARRYB_51__38_,
         u5_mult_87_CARRYB_51__39_, u5_mult_87_CARRYB_51__40_,
         u5_mult_87_CARRYB_51__41_, u5_mult_87_CARRYB_51__42_,
         u5_mult_87_CARRYB_51__43_, u5_mult_87_CARRYB_51__44_,
         u5_mult_87_CARRYB_51__45_, u5_mult_87_CARRYB_51__46_,
         u5_mult_87_CARRYB_51__47_, u5_mult_87_CARRYB_51__48_,
         u5_mult_87_CARRYB_51__49_, u5_mult_87_CARRYB_51__50_,
         u5_mult_87_CARRYB_51__51_, u5_mult_87_CARRYB_52__0_,
         u5_mult_87_CARRYB_52__1_, u5_mult_87_CARRYB_52__2_,
         u5_mult_87_CARRYB_52__3_, u5_mult_87_CARRYB_52__4_,
         u5_mult_87_CARRYB_52__5_, u5_mult_87_CARRYB_52__6_,
         u5_mult_87_CARRYB_52__7_, u5_mult_87_CARRYB_52__8_,
         u5_mult_87_CARRYB_52__9_, u5_mult_87_CARRYB_52__10_,
         u5_mult_87_CARRYB_52__11_, u5_mult_87_CARRYB_52__12_,
         u5_mult_87_CARRYB_52__13_, u5_mult_87_CARRYB_52__14_,
         u5_mult_87_CARRYB_52__15_, u5_mult_87_CARRYB_52__16_,
         u5_mult_87_CARRYB_52__17_, u5_mult_87_CARRYB_52__18_,
         u5_mult_87_CARRYB_52__19_, u5_mult_87_CARRYB_52__20_,
         u5_mult_87_CARRYB_52__21_, u5_mult_87_CARRYB_52__22_,
         u5_mult_87_CARRYB_52__23_, u5_mult_87_CARRYB_52__24_,
         u5_mult_87_CARRYB_52__25_, u5_mult_87_CARRYB_52__26_,
         u5_mult_87_CARRYB_52__27_, u5_mult_87_CARRYB_52__28_,
         u5_mult_87_CARRYB_52__29_, u5_mult_87_CARRYB_52__30_,
         u5_mult_87_CARRYB_52__31_, u5_mult_87_CARRYB_52__32_,
         u5_mult_87_CARRYB_52__33_, u5_mult_87_CARRYB_52__34_,
         u5_mult_87_CARRYB_52__35_, u5_mult_87_CARRYB_52__36_,
         u5_mult_87_CARRYB_52__37_, u5_mult_87_CARRYB_52__38_,
         u5_mult_87_CARRYB_52__39_, u5_mult_87_CARRYB_52__40_,
         u5_mult_87_CARRYB_52__41_, u5_mult_87_CARRYB_52__42_,
         u5_mult_87_CARRYB_52__43_, u5_mult_87_CARRYB_52__44_,
         u5_mult_87_CARRYB_52__45_, u5_mult_87_CARRYB_52__46_,
         u5_mult_87_CARRYB_52__47_, u5_mult_87_CARRYB_52__48_,
         u5_mult_87_CARRYB_52__49_, u5_mult_87_CARRYB_52__50_,
         u5_mult_87_CARRYB_52__51_, u5_mult_87_SUMB_33__36_,
         u5_mult_87_SUMB_33__37_, u5_mult_87_SUMB_33__38_,
         u5_mult_87_SUMB_33__39_, u5_mult_87_SUMB_33__40_,
         u5_mult_87_SUMB_33__41_, u5_mult_87_SUMB_33__42_,
         u5_mult_87_SUMB_33__43_, u5_mult_87_SUMB_33__44_,
         u5_mult_87_SUMB_33__45_, u5_mult_87_SUMB_33__46_,
         u5_mult_87_SUMB_33__47_, u5_mult_87_SUMB_33__48_,
         u5_mult_87_SUMB_33__49_, u5_mult_87_SUMB_33__50_,
         u5_mult_87_SUMB_33__51_, u5_mult_87_SUMB_34__1_,
         u5_mult_87_SUMB_34__2_, u5_mult_87_SUMB_34__3_,
         u5_mult_87_SUMB_34__4_, u5_mult_87_SUMB_34__5_,
         u5_mult_87_SUMB_34__6_, u5_mult_87_SUMB_34__7_,
         u5_mult_87_SUMB_34__8_, u5_mult_87_SUMB_34__9_,
         u5_mult_87_SUMB_34__10_, u5_mult_87_SUMB_34__11_,
         u5_mult_87_SUMB_34__12_, u5_mult_87_SUMB_34__13_,
         u5_mult_87_SUMB_34__14_, u5_mult_87_SUMB_34__15_,
         u5_mult_87_SUMB_34__16_, u5_mult_87_SUMB_34__17_,
         u5_mult_87_SUMB_34__18_, u5_mult_87_SUMB_34__19_,
         u5_mult_87_SUMB_34__20_, u5_mult_87_SUMB_34__21_,
         u5_mult_87_SUMB_34__22_, u5_mult_87_SUMB_34__23_,
         u5_mult_87_SUMB_34__24_, u5_mult_87_SUMB_34__25_,
         u5_mult_87_SUMB_34__26_, u5_mult_87_SUMB_34__27_,
         u5_mult_87_SUMB_34__28_, u5_mult_87_SUMB_34__29_,
         u5_mult_87_SUMB_34__30_, u5_mult_87_SUMB_34__31_,
         u5_mult_87_SUMB_34__32_, u5_mult_87_SUMB_34__33_,
         u5_mult_87_SUMB_34__34_, u5_mult_87_SUMB_34__35_,
         u5_mult_87_SUMB_34__36_, u5_mult_87_SUMB_34__37_,
         u5_mult_87_SUMB_34__38_, u5_mult_87_SUMB_34__39_,
         u5_mult_87_SUMB_34__40_, u5_mult_87_SUMB_34__41_,
         u5_mult_87_SUMB_34__42_, u5_mult_87_SUMB_34__43_,
         u5_mult_87_SUMB_34__44_, u5_mult_87_SUMB_34__45_,
         u5_mult_87_SUMB_34__46_, u5_mult_87_SUMB_34__47_,
         u5_mult_87_SUMB_34__48_, u5_mult_87_SUMB_34__49_,
         u5_mult_87_SUMB_34__50_, u5_mult_87_SUMB_34__51_,
         u5_mult_87_SUMB_35__1_, u5_mult_87_SUMB_35__2_,
         u5_mult_87_SUMB_35__3_, u5_mult_87_SUMB_35__4_,
         u5_mult_87_SUMB_35__5_, u5_mult_87_SUMB_35__6_,
         u5_mult_87_SUMB_35__7_, u5_mult_87_SUMB_35__8_,
         u5_mult_87_SUMB_35__9_, u5_mult_87_SUMB_35__10_,
         u5_mult_87_SUMB_35__11_, u5_mult_87_SUMB_35__12_,
         u5_mult_87_SUMB_35__13_, u5_mult_87_SUMB_35__14_,
         u5_mult_87_SUMB_35__15_, u5_mult_87_SUMB_35__16_,
         u5_mult_87_SUMB_35__17_, u5_mult_87_SUMB_35__18_,
         u5_mult_87_SUMB_35__19_, u5_mult_87_SUMB_35__20_,
         u5_mult_87_SUMB_35__21_, u5_mult_87_SUMB_35__22_,
         u5_mult_87_SUMB_35__23_, u5_mult_87_SUMB_35__24_,
         u5_mult_87_SUMB_35__25_, u5_mult_87_SUMB_35__26_,
         u5_mult_87_SUMB_35__27_, u5_mult_87_SUMB_35__28_,
         u5_mult_87_SUMB_35__29_, u5_mult_87_SUMB_35__30_,
         u5_mult_87_SUMB_35__31_, u5_mult_87_SUMB_35__32_,
         u5_mult_87_SUMB_35__33_, u5_mult_87_SUMB_35__34_,
         u5_mult_87_SUMB_35__35_, u5_mult_87_SUMB_35__36_,
         u5_mult_87_SUMB_35__37_, u5_mult_87_SUMB_35__38_,
         u5_mult_87_SUMB_35__39_, u5_mult_87_SUMB_35__40_,
         u5_mult_87_SUMB_35__41_, u5_mult_87_SUMB_35__42_,
         u5_mult_87_SUMB_35__43_, u5_mult_87_SUMB_35__44_,
         u5_mult_87_SUMB_35__45_, u5_mult_87_SUMB_35__46_,
         u5_mult_87_SUMB_35__47_, u5_mult_87_SUMB_35__48_,
         u5_mult_87_SUMB_35__49_, u5_mult_87_SUMB_35__50_,
         u5_mult_87_SUMB_35__51_, u5_mult_87_SUMB_36__1_,
         u5_mult_87_SUMB_36__2_, u5_mult_87_SUMB_36__3_,
         u5_mult_87_SUMB_36__4_, u5_mult_87_SUMB_36__5_,
         u5_mult_87_SUMB_36__6_, u5_mult_87_SUMB_36__7_,
         u5_mult_87_SUMB_36__8_, u5_mult_87_SUMB_36__9_,
         u5_mult_87_SUMB_36__10_, u5_mult_87_SUMB_36__11_,
         u5_mult_87_SUMB_36__12_, u5_mult_87_SUMB_36__13_,
         u5_mult_87_SUMB_36__14_, u5_mult_87_SUMB_36__15_,
         u5_mult_87_SUMB_36__16_, u5_mult_87_SUMB_36__17_,
         u5_mult_87_SUMB_36__18_, u5_mult_87_SUMB_36__19_,
         u5_mult_87_SUMB_36__20_, u5_mult_87_SUMB_36__21_,
         u5_mult_87_SUMB_36__22_, u5_mult_87_SUMB_36__23_,
         u5_mult_87_SUMB_36__24_, u5_mult_87_SUMB_36__25_,
         u5_mult_87_SUMB_36__26_, u5_mult_87_SUMB_36__27_,
         u5_mult_87_SUMB_36__28_, u5_mult_87_SUMB_36__29_,
         u5_mult_87_SUMB_36__30_, u5_mult_87_SUMB_36__31_,
         u5_mult_87_SUMB_36__32_, u5_mult_87_SUMB_36__33_,
         u5_mult_87_SUMB_36__34_, u5_mult_87_SUMB_36__35_,
         u5_mult_87_SUMB_36__36_, u5_mult_87_SUMB_36__37_,
         u5_mult_87_SUMB_36__38_, u5_mult_87_SUMB_36__39_,
         u5_mult_87_SUMB_36__40_, u5_mult_87_SUMB_36__41_,
         u5_mult_87_SUMB_36__42_, u5_mult_87_SUMB_36__43_,
         u5_mult_87_SUMB_36__44_, u5_mult_87_SUMB_36__45_,
         u5_mult_87_SUMB_36__46_, u5_mult_87_SUMB_36__47_,
         u5_mult_87_SUMB_36__48_, u5_mult_87_SUMB_36__49_,
         u5_mult_87_SUMB_36__50_, u5_mult_87_SUMB_36__51_,
         u5_mult_87_SUMB_37__1_, u5_mult_87_SUMB_37__2_,
         u5_mult_87_SUMB_37__3_, u5_mult_87_SUMB_37__4_,
         u5_mult_87_SUMB_37__5_, u5_mult_87_SUMB_37__6_,
         u5_mult_87_SUMB_37__7_, u5_mult_87_SUMB_37__8_,
         u5_mult_87_SUMB_37__9_, u5_mult_87_SUMB_37__10_,
         u5_mult_87_SUMB_37__11_, u5_mult_87_SUMB_37__12_,
         u5_mult_87_SUMB_37__13_, u5_mult_87_SUMB_37__14_,
         u5_mult_87_SUMB_37__15_, u5_mult_87_SUMB_37__16_,
         u5_mult_87_SUMB_37__17_, u5_mult_87_SUMB_37__18_,
         u5_mult_87_SUMB_37__19_, u5_mult_87_SUMB_37__20_,
         u5_mult_87_SUMB_37__21_, u5_mult_87_SUMB_37__22_,
         u5_mult_87_SUMB_37__23_, u5_mult_87_SUMB_37__24_,
         u5_mult_87_SUMB_37__25_, u5_mult_87_SUMB_37__26_,
         u5_mult_87_SUMB_37__27_, u5_mult_87_SUMB_37__28_,
         u5_mult_87_SUMB_37__29_, u5_mult_87_SUMB_37__30_,
         u5_mult_87_SUMB_37__31_, u5_mult_87_SUMB_37__32_,
         u5_mult_87_SUMB_37__33_, u5_mult_87_SUMB_37__34_,
         u5_mult_87_SUMB_37__35_, u5_mult_87_SUMB_37__36_,
         u5_mult_87_SUMB_37__37_, u5_mult_87_SUMB_37__38_,
         u5_mult_87_SUMB_37__39_, u5_mult_87_SUMB_37__40_,
         u5_mult_87_SUMB_37__41_, u5_mult_87_SUMB_37__42_,
         u5_mult_87_SUMB_37__43_, u5_mult_87_SUMB_37__44_,
         u5_mult_87_SUMB_37__45_, u5_mult_87_SUMB_37__46_,
         u5_mult_87_SUMB_37__47_, u5_mult_87_SUMB_37__48_,
         u5_mult_87_SUMB_37__49_, u5_mult_87_SUMB_37__50_,
         u5_mult_87_SUMB_37__51_, u5_mult_87_SUMB_38__1_,
         u5_mult_87_SUMB_38__2_, u5_mult_87_SUMB_38__3_,
         u5_mult_87_SUMB_38__4_, u5_mult_87_SUMB_38__5_,
         u5_mult_87_SUMB_38__6_, u5_mult_87_SUMB_38__7_,
         u5_mult_87_SUMB_38__8_, u5_mult_87_SUMB_38__9_,
         u5_mult_87_SUMB_38__10_, u5_mult_87_SUMB_38__11_,
         u5_mult_87_SUMB_38__12_, u5_mult_87_SUMB_38__13_,
         u5_mult_87_SUMB_38__14_, u5_mult_87_SUMB_38__15_,
         u5_mult_87_SUMB_38__16_, u5_mult_87_SUMB_38__17_,
         u5_mult_87_SUMB_38__18_, u5_mult_87_SUMB_38__19_,
         u5_mult_87_SUMB_38__20_, u5_mult_87_SUMB_38__21_,
         u5_mult_87_SUMB_38__22_, u5_mult_87_SUMB_38__23_,
         u5_mult_87_SUMB_38__24_, u5_mult_87_SUMB_38__25_,
         u5_mult_87_SUMB_38__26_, u5_mult_87_SUMB_38__27_,
         u5_mult_87_SUMB_38__28_, u5_mult_87_SUMB_38__29_,
         u5_mult_87_SUMB_38__30_, u5_mult_87_SUMB_38__31_,
         u5_mult_87_SUMB_38__32_, u5_mult_87_SUMB_38__33_,
         u5_mult_87_SUMB_38__34_, u5_mult_87_SUMB_38__35_,
         u5_mult_87_SUMB_38__36_, u5_mult_87_SUMB_38__37_,
         u5_mult_87_SUMB_38__38_, u5_mult_87_SUMB_38__39_,
         u5_mult_87_SUMB_38__40_, u5_mult_87_SUMB_38__41_,
         u5_mult_87_SUMB_38__42_, u5_mult_87_SUMB_38__43_,
         u5_mult_87_SUMB_38__44_, u5_mult_87_SUMB_38__45_,
         u5_mult_87_SUMB_38__46_, u5_mult_87_SUMB_38__47_,
         u5_mult_87_SUMB_38__48_, u5_mult_87_SUMB_38__49_,
         u5_mult_87_SUMB_38__50_, u5_mult_87_SUMB_38__51_,
         u5_mult_87_SUMB_39__1_, u5_mult_87_SUMB_39__2_,
         u5_mult_87_SUMB_39__3_, u5_mult_87_SUMB_39__4_,
         u5_mult_87_SUMB_39__5_, u5_mult_87_SUMB_39__6_,
         u5_mult_87_SUMB_39__7_, u5_mult_87_SUMB_39__8_,
         u5_mult_87_SUMB_39__9_, u5_mult_87_SUMB_39__10_,
         u5_mult_87_SUMB_39__11_, u5_mult_87_SUMB_39__12_,
         u5_mult_87_SUMB_39__13_, u5_mult_87_SUMB_39__14_,
         u5_mult_87_SUMB_39__15_, u5_mult_87_SUMB_39__16_,
         u5_mult_87_SUMB_39__17_, u5_mult_87_SUMB_39__18_,
         u5_mult_87_SUMB_39__19_, u5_mult_87_SUMB_39__20_,
         u5_mult_87_SUMB_39__21_, u5_mult_87_SUMB_39__22_,
         u5_mult_87_SUMB_39__23_, u5_mult_87_SUMB_39__24_,
         u5_mult_87_SUMB_39__25_, u5_mult_87_SUMB_39__26_,
         u5_mult_87_SUMB_39__27_, u5_mult_87_SUMB_39__28_,
         u5_mult_87_SUMB_39__29_, u5_mult_87_SUMB_39__30_,
         u5_mult_87_SUMB_39__31_, u5_mult_87_SUMB_39__32_,
         u5_mult_87_SUMB_39__33_, u5_mult_87_SUMB_39__34_,
         u5_mult_87_SUMB_39__35_, u5_mult_87_SUMB_39__36_,
         u5_mult_87_SUMB_39__37_, u5_mult_87_SUMB_39__38_,
         u5_mult_87_SUMB_39__39_, u5_mult_87_SUMB_39__40_,
         u5_mult_87_SUMB_39__41_, u5_mult_87_SUMB_39__42_,
         u5_mult_87_SUMB_39__43_, u5_mult_87_SUMB_39__44_,
         u5_mult_87_SUMB_39__45_, u5_mult_87_SUMB_39__46_,
         u5_mult_87_SUMB_39__47_, u5_mult_87_SUMB_39__48_,
         u5_mult_87_SUMB_39__49_, u5_mult_87_SUMB_39__50_,
         u5_mult_87_SUMB_39__51_, u5_mult_87_SUMB_40__1_,
         u5_mult_87_SUMB_40__2_, u5_mult_87_SUMB_40__3_,
         u5_mult_87_SUMB_40__4_, u5_mult_87_SUMB_40__5_,
         u5_mult_87_SUMB_40__6_, u5_mult_87_SUMB_40__7_,
         u5_mult_87_SUMB_40__8_, u5_mult_87_SUMB_40__9_,
         u5_mult_87_SUMB_40__10_, u5_mult_87_SUMB_40__11_,
         u5_mult_87_SUMB_40__12_, u5_mult_87_SUMB_40__13_,
         u5_mult_87_SUMB_40__14_, u5_mult_87_SUMB_40__15_,
         u5_mult_87_SUMB_40__16_, u5_mult_87_SUMB_40__17_,
         u5_mult_87_SUMB_40__18_, u5_mult_87_SUMB_40__19_,
         u5_mult_87_SUMB_40__20_, u5_mult_87_SUMB_40__21_,
         u5_mult_87_SUMB_40__22_, u5_mult_87_SUMB_40__23_,
         u5_mult_87_SUMB_40__24_, u5_mult_87_SUMB_40__25_,
         u5_mult_87_SUMB_40__26_, u5_mult_87_SUMB_40__27_,
         u5_mult_87_SUMB_40__28_, u5_mult_87_SUMB_40__29_,
         u5_mult_87_SUMB_40__30_, u5_mult_87_SUMB_40__31_,
         u5_mult_87_SUMB_40__32_, u5_mult_87_SUMB_40__33_,
         u5_mult_87_SUMB_40__34_, u5_mult_87_SUMB_40__35_,
         u5_mult_87_SUMB_40__36_, u5_mult_87_SUMB_40__37_,
         u5_mult_87_SUMB_40__38_, u5_mult_87_SUMB_40__39_,
         u5_mult_87_SUMB_40__40_, u5_mult_87_SUMB_40__41_,
         u5_mult_87_SUMB_40__42_, u5_mult_87_SUMB_40__43_,
         u5_mult_87_SUMB_40__44_, u5_mult_87_SUMB_40__45_,
         u5_mult_87_SUMB_40__46_, u5_mult_87_SUMB_40__47_,
         u5_mult_87_SUMB_40__48_, u5_mult_87_SUMB_40__49_,
         u5_mult_87_SUMB_40__50_, u5_mult_87_SUMB_40__51_,
         u5_mult_87_SUMB_41__1_, u5_mult_87_SUMB_41__2_,
         u5_mult_87_SUMB_41__3_, u5_mult_87_SUMB_41__4_,
         u5_mult_87_SUMB_41__5_, u5_mult_87_SUMB_41__6_,
         u5_mult_87_SUMB_41__7_, u5_mult_87_SUMB_41__8_,
         u5_mult_87_SUMB_41__9_, u5_mult_87_SUMB_41__10_,
         u5_mult_87_SUMB_41__11_, u5_mult_87_SUMB_41__12_,
         u5_mult_87_SUMB_41__13_, u5_mult_87_SUMB_41__14_,
         u5_mult_87_SUMB_41__15_, u5_mult_87_SUMB_41__16_,
         u5_mult_87_SUMB_41__17_, u5_mult_87_SUMB_41__18_,
         u5_mult_87_SUMB_41__19_, u5_mult_87_SUMB_41__20_,
         u5_mult_87_SUMB_41__21_, u5_mult_87_SUMB_41__22_,
         u5_mult_87_SUMB_41__23_, u5_mult_87_SUMB_41__24_,
         u5_mult_87_SUMB_41__25_, u5_mult_87_SUMB_41__26_,
         u5_mult_87_SUMB_41__27_, u5_mult_87_SUMB_41__28_,
         u5_mult_87_SUMB_41__29_, u5_mult_87_SUMB_41__30_,
         u5_mult_87_SUMB_41__31_, u5_mult_87_SUMB_41__32_,
         u5_mult_87_SUMB_41__33_, u5_mult_87_SUMB_41__34_,
         u5_mult_87_SUMB_41__35_, u5_mult_87_SUMB_41__36_,
         u5_mult_87_SUMB_41__37_, u5_mult_87_SUMB_41__38_,
         u5_mult_87_SUMB_41__39_, u5_mult_87_SUMB_41__40_,
         u5_mult_87_SUMB_41__41_, u5_mult_87_SUMB_41__42_,
         u5_mult_87_SUMB_41__43_, u5_mult_87_SUMB_41__44_,
         u5_mult_87_SUMB_41__45_, u5_mult_87_SUMB_41__46_,
         u5_mult_87_SUMB_41__47_, u5_mult_87_SUMB_41__48_,
         u5_mult_87_SUMB_41__49_, u5_mult_87_SUMB_41__50_,
         u5_mult_87_SUMB_41__51_, u5_mult_87_SUMB_42__1_,
         u5_mult_87_SUMB_42__2_, u5_mult_87_SUMB_42__3_,
         u5_mult_87_SUMB_42__4_, u5_mult_87_SUMB_42__5_,
         u5_mult_87_SUMB_42__6_, u5_mult_87_SUMB_42__7_,
         u5_mult_87_SUMB_42__8_, u5_mult_87_SUMB_42__9_,
         u5_mult_87_SUMB_42__10_, u5_mult_87_SUMB_42__11_,
         u5_mult_87_SUMB_42__12_, u5_mult_87_SUMB_42__13_,
         u5_mult_87_SUMB_42__14_, u5_mult_87_SUMB_42__15_,
         u5_mult_87_SUMB_42__16_, u5_mult_87_SUMB_42__17_,
         u5_mult_87_SUMB_42__18_, u5_mult_87_SUMB_42__19_,
         u5_mult_87_SUMB_42__20_, u5_mult_87_SUMB_42__21_,
         u5_mult_87_SUMB_42__22_, u5_mult_87_SUMB_42__23_,
         u5_mult_87_SUMB_42__24_, u5_mult_87_SUMB_42__25_,
         u5_mult_87_SUMB_42__26_, u5_mult_87_SUMB_42__27_,
         u5_mult_87_SUMB_42__28_, u5_mult_87_SUMB_42__29_,
         u5_mult_87_SUMB_42__30_, u5_mult_87_SUMB_42__31_,
         u5_mult_87_SUMB_42__32_, u5_mult_87_SUMB_42__33_,
         u5_mult_87_SUMB_42__34_, u5_mult_87_SUMB_42__35_,
         u5_mult_87_SUMB_42__36_, u5_mult_87_SUMB_42__37_,
         u5_mult_87_SUMB_42__38_, u5_mult_87_SUMB_42__39_,
         u5_mult_87_SUMB_42__40_, u5_mult_87_SUMB_42__41_,
         u5_mult_87_SUMB_42__42_, u5_mult_87_SUMB_42__43_,
         u5_mult_87_SUMB_42__44_, u5_mult_87_SUMB_42__45_,
         u5_mult_87_SUMB_42__46_, u5_mult_87_SUMB_42__47_,
         u5_mult_87_SUMB_42__48_, u5_mult_87_SUMB_42__49_,
         u5_mult_87_SUMB_42__50_, u5_mult_87_SUMB_42__51_,
         u5_mult_87_SUMB_43__1_, u5_mult_87_SUMB_43__2_,
         u5_mult_87_SUMB_43__3_, u5_mult_87_SUMB_43__4_,
         u5_mult_87_SUMB_43__5_, u5_mult_87_SUMB_43__6_,
         u5_mult_87_SUMB_43__7_, u5_mult_87_SUMB_43__8_,
         u5_mult_87_SUMB_43__9_, u5_mult_87_SUMB_43__10_,
         u5_mult_87_SUMB_43__11_, u5_mult_87_SUMB_43__12_,
         u5_mult_87_SUMB_43__13_, u5_mult_87_SUMB_43__14_,
         u5_mult_87_SUMB_43__15_, u5_mult_87_SUMB_43__16_,
         u5_mult_87_SUMB_43__17_, u5_mult_87_CARRYB_33__36_,
         u5_mult_87_CARRYB_33__37_, u5_mult_87_CARRYB_33__38_,
         u5_mult_87_CARRYB_33__39_, u5_mult_87_CARRYB_33__40_,
         u5_mult_87_CARRYB_33__41_, u5_mult_87_CARRYB_33__42_,
         u5_mult_87_CARRYB_33__43_, u5_mult_87_CARRYB_33__44_,
         u5_mult_87_CARRYB_33__45_, u5_mult_87_CARRYB_33__46_,
         u5_mult_87_CARRYB_33__47_, u5_mult_87_CARRYB_33__48_,
         u5_mult_87_CARRYB_33__49_, u5_mult_87_CARRYB_33__50_,
         u5_mult_87_CARRYB_33__51_, u5_mult_87_CARRYB_34__0_,
         u5_mult_87_CARRYB_34__1_, u5_mult_87_CARRYB_34__2_,
         u5_mult_87_CARRYB_34__3_, u5_mult_87_CARRYB_34__4_,
         u5_mult_87_CARRYB_34__5_, u5_mult_87_CARRYB_34__6_,
         u5_mult_87_CARRYB_34__7_, u5_mult_87_CARRYB_34__8_,
         u5_mult_87_CARRYB_34__9_, u5_mult_87_CARRYB_34__10_,
         u5_mult_87_CARRYB_34__11_, u5_mult_87_CARRYB_34__12_,
         u5_mult_87_CARRYB_34__13_, u5_mult_87_CARRYB_34__14_,
         u5_mult_87_CARRYB_34__15_, u5_mult_87_CARRYB_34__16_,
         u5_mult_87_CARRYB_34__17_, u5_mult_87_CARRYB_34__18_,
         u5_mult_87_CARRYB_34__19_, u5_mult_87_CARRYB_34__20_,
         u5_mult_87_CARRYB_34__21_, u5_mult_87_CARRYB_34__22_,
         u5_mult_87_CARRYB_34__23_, u5_mult_87_CARRYB_34__24_,
         u5_mult_87_CARRYB_34__25_, u5_mult_87_CARRYB_34__26_,
         u5_mult_87_CARRYB_34__27_, u5_mult_87_CARRYB_34__28_,
         u5_mult_87_CARRYB_34__29_, u5_mult_87_CARRYB_34__30_,
         u5_mult_87_CARRYB_34__31_, u5_mult_87_CARRYB_34__32_,
         u5_mult_87_CARRYB_34__33_, u5_mult_87_CARRYB_34__34_,
         u5_mult_87_CARRYB_34__35_, u5_mult_87_CARRYB_34__36_,
         u5_mult_87_CARRYB_34__37_, u5_mult_87_CARRYB_34__38_,
         u5_mult_87_CARRYB_34__39_, u5_mult_87_CARRYB_34__40_,
         u5_mult_87_CARRYB_34__41_, u5_mult_87_CARRYB_34__42_,
         u5_mult_87_CARRYB_34__43_, u5_mult_87_CARRYB_34__44_,
         u5_mult_87_CARRYB_34__45_, u5_mult_87_CARRYB_34__46_,
         u5_mult_87_CARRYB_34__47_, u5_mult_87_CARRYB_34__48_,
         u5_mult_87_CARRYB_34__49_, u5_mult_87_CARRYB_34__50_,
         u5_mult_87_CARRYB_34__51_, u5_mult_87_CARRYB_35__0_,
         u5_mult_87_CARRYB_35__1_, u5_mult_87_CARRYB_35__2_,
         u5_mult_87_CARRYB_35__3_, u5_mult_87_CARRYB_35__4_,
         u5_mult_87_CARRYB_35__5_, u5_mult_87_CARRYB_35__6_,
         u5_mult_87_CARRYB_35__7_, u5_mult_87_CARRYB_35__8_,
         u5_mult_87_CARRYB_35__9_, u5_mult_87_CARRYB_35__10_,
         u5_mult_87_CARRYB_35__11_, u5_mult_87_CARRYB_35__12_,
         u5_mult_87_CARRYB_35__13_, u5_mult_87_CARRYB_35__14_,
         u5_mult_87_CARRYB_35__15_, u5_mult_87_CARRYB_35__16_,
         u5_mult_87_CARRYB_35__17_, u5_mult_87_CARRYB_35__18_,
         u5_mult_87_CARRYB_35__19_, u5_mult_87_CARRYB_35__20_,
         u5_mult_87_CARRYB_35__21_, u5_mult_87_CARRYB_35__22_,
         u5_mult_87_CARRYB_35__23_, u5_mult_87_CARRYB_35__24_,
         u5_mult_87_CARRYB_35__25_, u5_mult_87_CARRYB_35__26_,
         u5_mult_87_CARRYB_35__27_, u5_mult_87_CARRYB_35__28_,
         u5_mult_87_CARRYB_35__29_, u5_mult_87_CARRYB_35__30_,
         u5_mult_87_CARRYB_35__31_, u5_mult_87_CARRYB_35__32_,
         u5_mult_87_CARRYB_35__33_, u5_mult_87_CARRYB_35__34_,
         u5_mult_87_CARRYB_35__35_, u5_mult_87_CARRYB_35__36_,
         u5_mult_87_CARRYB_35__37_, u5_mult_87_CARRYB_35__38_,
         u5_mult_87_CARRYB_35__39_, u5_mult_87_CARRYB_35__40_,
         u5_mult_87_CARRYB_35__41_, u5_mult_87_CARRYB_35__42_,
         u5_mult_87_CARRYB_35__43_, u5_mult_87_CARRYB_35__44_,
         u5_mult_87_CARRYB_35__45_, u5_mult_87_CARRYB_35__46_,
         u5_mult_87_CARRYB_35__47_, u5_mult_87_CARRYB_35__48_,
         u5_mult_87_CARRYB_35__49_, u5_mult_87_CARRYB_35__50_,
         u5_mult_87_CARRYB_35__51_, u5_mult_87_CARRYB_36__0_,
         u5_mult_87_CARRYB_36__1_, u5_mult_87_CARRYB_36__2_,
         u5_mult_87_CARRYB_36__3_, u5_mult_87_CARRYB_36__4_,
         u5_mult_87_CARRYB_36__5_, u5_mult_87_CARRYB_36__6_,
         u5_mult_87_CARRYB_36__7_, u5_mult_87_CARRYB_36__8_,
         u5_mult_87_CARRYB_36__9_, u5_mult_87_CARRYB_36__10_,
         u5_mult_87_CARRYB_36__11_, u5_mult_87_CARRYB_36__12_,
         u5_mult_87_CARRYB_36__13_, u5_mult_87_CARRYB_36__14_,
         u5_mult_87_CARRYB_36__15_, u5_mult_87_CARRYB_36__16_,
         u5_mult_87_CARRYB_36__17_, u5_mult_87_CARRYB_36__18_,
         u5_mult_87_CARRYB_36__19_, u5_mult_87_CARRYB_36__20_,
         u5_mult_87_CARRYB_36__21_, u5_mult_87_CARRYB_36__22_,
         u5_mult_87_CARRYB_36__23_, u5_mult_87_CARRYB_36__24_,
         u5_mult_87_CARRYB_36__25_, u5_mult_87_CARRYB_36__26_,
         u5_mult_87_CARRYB_36__27_, u5_mult_87_CARRYB_36__28_,
         u5_mult_87_CARRYB_36__29_, u5_mult_87_CARRYB_36__30_,
         u5_mult_87_CARRYB_36__31_, u5_mult_87_CARRYB_36__32_,
         u5_mult_87_CARRYB_36__33_, u5_mult_87_CARRYB_36__34_,
         u5_mult_87_CARRYB_36__35_, u5_mult_87_CARRYB_36__36_,
         u5_mult_87_CARRYB_36__37_, u5_mult_87_CARRYB_36__38_,
         u5_mult_87_CARRYB_36__39_, u5_mult_87_CARRYB_36__40_,
         u5_mult_87_CARRYB_36__41_, u5_mult_87_CARRYB_36__42_,
         u5_mult_87_CARRYB_36__43_, u5_mult_87_CARRYB_36__44_,
         u5_mult_87_CARRYB_36__45_, u5_mult_87_CARRYB_36__46_,
         u5_mult_87_CARRYB_36__47_, u5_mult_87_CARRYB_36__48_,
         u5_mult_87_CARRYB_36__49_, u5_mult_87_CARRYB_36__50_,
         u5_mult_87_CARRYB_36__51_, u5_mult_87_CARRYB_37__0_,
         u5_mult_87_CARRYB_37__1_, u5_mult_87_CARRYB_37__2_,
         u5_mult_87_CARRYB_37__3_, u5_mult_87_CARRYB_37__4_,
         u5_mult_87_CARRYB_37__5_, u5_mult_87_CARRYB_37__6_,
         u5_mult_87_CARRYB_37__7_, u5_mult_87_CARRYB_37__8_,
         u5_mult_87_CARRYB_37__9_, u5_mult_87_CARRYB_37__10_,
         u5_mult_87_CARRYB_37__11_, u5_mult_87_CARRYB_37__12_,
         u5_mult_87_CARRYB_37__13_, u5_mult_87_CARRYB_37__14_,
         u5_mult_87_CARRYB_37__15_, u5_mult_87_CARRYB_37__16_,
         u5_mult_87_CARRYB_37__17_, u5_mult_87_CARRYB_37__18_,
         u5_mult_87_CARRYB_37__19_, u5_mult_87_CARRYB_37__20_,
         u5_mult_87_CARRYB_37__21_, u5_mult_87_CARRYB_37__22_,
         u5_mult_87_CARRYB_37__23_, u5_mult_87_CARRYB_37__24_,
         u5_mult_87_CARRYB_37__25_, u5_mult_87_CARRYB_37__26_,
         u5_mult_87_CARRYB_37__27_, u5_mult_87_CARRYB_37__28_,
         u5_mult_87_CARRYB_37__29_, u5_mult_87_CARRYB_37__30_,
         u5_mult_87_CARRYB_37__31_, u5_mult_87_CARRYB_37__32_,
         u5_mult_87_CARRYB_37__33_, u5_mult_87_CARRYB_37__34_,
         u5_mult_87_CARRYB_37__35_, u5_mult_87_CARRYB_37__36_,
         u5_mult_87_CARRYB_37__37_, u5_mult_87_CARRYB_37__38_,
         u5_mult_87_CARRYB_37__39_, u5_mult_87_CARRYB_37__40_,
         u5_mult_87_CARRYB_37__41_, u5_mult_87_CARRYB_37__42_,
         u5_mult_87_CARRYB_37__43_, u5_mult_87_CARRYB_37__44_,
         u5_mult_87_CARRYB_37__45_, u5_mult_87_CARRYB_37__46_,
         u5_mult_87_CARRYB_37__47_, u5_mult_87_CARRYB_37__48_,
         u5_mult_87_CARRYB_37__49_, u5_mult_87_CARRYB_37__50_,
         u5_mult_87_CARRYB_37__51_, u5_mult_87_CARRYB_38__0_,
         u5_mult_87_CARRYB_38__1_, u5_mult_87_CARRYB_38__2_,
         u5_mult_87_CARRYB_38__3_, u5_mult_87_CARRYB_38__4_,
         u5_mult_87_CARRYB_38__5_, u5_mult_87_CARRYB_38__6_,
         u5_mult_87_CARRYB_38__7_, u5_mult_87_CARRYB_38__8_,
         u5_mult_87_CARRYB_38__9_, u5_mult_87_CARRYB_38__10_,
         u5_mult_87_CARRYB_38__11_, u5_mult_87_CARRYB_38__12_,
         u5_mult_87_CARRYB_38__13_, u5_mult_87_CARRYB_38__14_,
         u5_mult_87_CARRYB_38__15_, u5_mult_87_CARRYB_38__16_,
         u5_mult_87_CARRYB_38__17_, u5_mult_87_CARRYB_38__18_,
         u5_mult_87_CARRYB_38__19_, u5_mult_87_CARRYB_38__20_,
         u5_mult_87_CARRYB_38__21_, u5_mult_87_CARRYB_38__22_,
         u5_mult_87_CARRYB_38__23_, u5_mult_87_CARRYB_38__24_,
         u5_mult_87_CARRYB_38__25_, u5_mult_87_CARRYB_38__26_,
         u5_mult_87_CARRYB_38__27_, u5_mult_87_CARRYB_38__28_,
         u5_mult_87_CARRYB_38__29_, u5_mult_87_CARRYB_38__30_,
         u5_mult_87_CARRYB_38__31_, u5_mult_87_CARRYB_38__32_,
         u5_mult_87_CARRYB_38__33_, u5_mult_87_CARRYB_38__34_,
         u5_mult_87_CARRYB_38__35_, u5_mult_87_CARRYB_38__36_,
         u5_mult_87_CARRYB_38__37_, u5_mult_87_CARRYB_38__38_,
         u5_mult_87_CARRYB_38__39_, u5_mult_87_CARRYB_38__40_,
         u5_mult_87_CARRYB_38__41_, u5_mult_87_CARRYB_38__42_,
         u5_mult_87_CARRYB_38__43_, u5_mult_87_CARRYB_38__44_,
         u5_mult_87_CARRYB_38__45_, u5_mult_87_CARRYB_38__46_,
         u5_mult_87_CARRYB_38__47_, u5_mult_87_CARRYB_38__48_,
         u5_mult_87_CARRYB_38__49_, u5_mult_87_CARRYB_38__50_,
         u5_mult_87_CARRYB_38__51_, u5_mult_87_CARRYB_39__0_,
         u5_mult_87_CARRYB_39__1_, u5_mult_87_CARRYB_39__2_,
         u5_mult_87_CARRYB_39__3_, u5_mult_87_CARRYB_39__4_,
         u5_mult_87_CARRYB_39__5_, u5_mult_87_CARRYB_39__6_,
         u5_mult_87_CARRYB_39__7_, u5_mult_87_CARRYB_39__8_,
         u5_mult_87_CARRYB_39__9_, u5_mult_87_CARRYB_39__10_,
         u5_mult_87_CARRYB_39__11_, u5_mult_87_CARRYB_39__12_,
         u5_mult_87_CARRYB_39__13_, u5_mult_87_CARRYB_39__14_,
         u5_mult_87_CARRYB_39__15_, u5_mult_87_CARRYB_39__16_,
         u5_mult_87_CARRYB_39__17_, u5_mult_87_CARRYB_39__18_,
         u5_mult_87_CARRYB_39__19_, u5_mult_87_CARRYB_39__20_,
         u5_mult_87_CARRYB_39__21_, u5_mult_87_CARRYB_39__22_,
         u5_mult_87_CARRYB_39__23_, u5_mult_87_CARRYB_39__24_,
         u5_mult_87_CARRYB_39__25_, u5_mult_87_CARRYB_39__26_,
         u5_mult_87_CARRYB_39__27_, u5_mult_87_CARRYB_39__28_,
         u5_mult_87_CARRYB_39__29_, u5_mult_87_CARRYB_39__30_,
         u5_mult_87_CARRYB_39__31_, u5_mult_87_CARRYB_39__32_,
         u5_mult_87_CARRYB_39__33_, u5_mult_87_CARRYB_39__34_,
         u5_mult_87_CARRYB_39__35_, u5_mult_87_CARRYB_39__36_,
         u5_mult_87_CARRYB_39__37_, u5_mult_87_CARRYB_39__38_,
         u5_mult_87_CARRYB_39__39_, u5_mult_87_CARRYB_39__40_,
         u5_mult_87_CARRYB_39__41_, u5_mult_87_CARRYB_39__42_,
         u5_mult_87_CARRYB_39__43_, u5_mult_87_CARRYB_39__44_,
         u5_mult_87_CARRYB_39__45_, u5_mult_87_CARRYB_39__46_,
         u5_mult_87_CARRYB_39__47_, u5_mult_87_CARRYB_39__48_,
         u5_mult_87_CARRYB_39__49_, u5_mult_87_CARRYB_39__50_,
         u5_mult_87_CARRYB_39__51_, u5_mult_87_CARRYB_40__0_,
         u5_mult_87_CARRYB_40__1_, u5_mult_87_CARRYB_40__2_,
         u5_mult_87_CARRYB_40__3_, u5_mult_87_CARRYB_40__4_,
         u5_mult_87_CARRYB_40__5_, u5_mult_87_CARRYB_40__6_,
         u5_mult_87_CARRYB_40__7_, u5_mult_87_CARRYB_40__8_,
         u5_mult_87_CARRYB_40__9_, u5_mult_87_CARRYB_40__10_,
         u5_mult_87_CARRYB_40__11_, u5_mult_87_CARRYB_40__12_,
         u5_mult_87_CARRYB_40__13_, u5_mult_87_CARRYB_40__14_,
         u5_mult_87_CARRYB_40__15_, u5_mult_87_CARRYB_40__16_,
         u5_mult_87_CARRYB_40__17_, u5_mult_87_CARRYB_40__18_,
         u5_mult_87_CARRYB_40__19_, u5_mult_87_CARRYB_40__20_,
         u5_mult_87_CARRYB_40__21_, u5_mult_87_CARRYB_40__22_,
         u5_mult_87_CARRYB_40__23_, u5_mult_87_CARRYB_40__24_,
         u5_mult_87_CARRYB_40__25_, u5_mult_87_CARRYB_40__26_,
         u5_mult_87_CARRYB_40__27_, u5_mult_87_CARRYB_40__28_,
         u5_mult_87_CARRYB_40__29_, u5_mult_87_CARRYB_40__30_,
         u5_mult_87_CARRYB_40__31_, u5_mult_87_CARRYB_40__32_,
         u5_mult_87_CARRYB_40__33_, u5_mult_87_CARRYB_40__34_,
         u5_mult_87_CARRYB_40__35_, u5_mult_87_CARRYB_40__36_,
         u5_mult_87_CARRYB_40__37_, u5_mult_87_CARRYB_40__38_,
         u5_mult_87_CARRYB_40__39_, u5_mult_87_CARRYB_40__40_,
         u5_mult_87_CARRYB_40__41_, u5_mult_87_CARRYB_40__42_,
         u5_mult_87_CARRYB_40__43_, u5_mult_87_CARRYB_40__44_,
         u5_mult_87_CARRYB_40__45_, u5_mult_87_CARRYB_40__46_,
         u5_mult_87_CARRYB_40__47_, u5_mult_87_CARRYB_40__48_,
         u5_mult_87_CARRYB_40__49_, u5_mult_87_CARRYB_40__50_,
         u5_mult_87_CARRYB_40__51_, u5_mult_87_CARRYB_41__0_,
         u5_mult_87_CARRYB_41__1_, u5_mult_87_CARRYB_41__2_,
         u5_mult_87_CARRYB_41__3_, u5_mult_87_CARRYB_41__4_,
         u5_mult_87_CARRYB_41__5_, u5_mult_87_CARRYB_41__6_,
         u5_mult_87_CARRYB_41__7_, u5_mult_87_CARRYB_41__8_,
         u5_mult_87_CARRYB_41__9_, u5_mult_87_CARRYB_41__10_,
         u5_mult_87_CARRYB_41__11_, u5_mult_87_CARRYB_41__12_,
         u5_mult_87_CARRYB_41__13_, u5_mult_87_CARRYB_41__14_,
         u5_mult_87_CARRYB_41__15_, u5_mult_87_CARRYB_41__16_,
         u5_mult_87_CARRYB_41__17_, u5_mult_87_CARRYB_41__18_,
         u5_mult_87_CARRYB_41__19_, u5_mult_87_CARRYB_41__20_,
         u5_mult_87_CARRYB_41__21_, u5_mult_87_CARRYB_41__22_,
         u5_mult_87_CARRYB_41__23_, u5_mult_87_CARRYB_41__24_,
         u5_mult_87_CARRYB_41__25_, u5_mult_87_CARRYB_41__26_,
         u5_mult_87_CARRYB_41__27_, u5_mult_87_CARRYB_41__28_,
         u5_mult_87_CARRYB_41__29_, u5_mult_87_CARRYB_41__30_,
         u5_mult_87_CARRYB_41__31_, u5_mult_87_CARRYB_41__32_,
         u5_mult_87_CARRYB_41__33_, u5_mult_87_CARRYB_41__34_,
         u5_mult_87_CARRYB_41__35_, u5_mult_87_CARRYB_41__36_,
         u5_mult_87_CARRYB_41__37_, u5_mult_87_CARRYB_41__38_,
         u5_mult_87_CARRYB_41__39_, u5_mult_87_CARRYB_41__40_,
         u5_mult_87_CARRYB_41__41_, u5_mult_87_CARRYB_41__42_,
         u5_mult_87_CARRYB_41__43_, u5_mult_87_CARRYB_41__44_,
         u5_mult_87_CARRYB_41__45_, u5_mult_87_CARRYB_41__46_,
         u5_mult_87_CARRYB_41__47_, u5_mult_87_CARRYB_41__48_,
         u5_mult_87_CARRYB_41__49_, u5_mult_87_CARRYB_41__50_,
         u5_mult_87_CARRYB_41__51_, u5_mult_87_CARRYB_42__0_,
         u5_mult_87_CARRYB_42__1_, u5_mult_87_CARRYB_42__2_,
         u5_mult_87_CARRYB_42__3_, u5_mult_87_CARRYB_42__4_,
         u5_mult_87_CARRYB_42__5_, u5_mult_87_CARRYB_42__6_,
         u5_mult_87_CARRYB_42__7_, u5_mult_87_CARRYB_42__8_,
         u5_mult_87_CARRYB_42__9_, u5_mult_87_CARRYB_42__10_,
         u5_mult_87_CARRYB_42__11_, u5_mult_87_CARRYB_42__12_,
         u5_mult_87_CARRYB_42__13_, u5_mult_87_CARRYB_42__14_,
         u5_mult_87_CARRYB_42__15_, u5_mult_87_CARRYB_42__16_,
         u5_mult_87_CARRYB_42__17_, u5_mult_87_CARRYB_42__18_,
         u5_mult_87_CARRYB_42__19_, u5_mult_87_CARRYB_42__20_,
         u5_mult_87_CARRYB_42__21_, u5_mult_87_CARRYB_42__22_,
         u5_mult_87_CARRYB_42__23_, u5_mult_87_CARRYB_42__24_,
         u5_mult_87_CARRYB_42__25_, u5_mult_87_CARRYB_42__26_,
         u5_mult_87_CARRYB_42__27_, u5_mult_87_CARRYB_42__28_,
         u5_mult_87_CARRYB_42__29_, u5_mult_87_CARRYB_42__30_,
         u5_mult_87_CARRYB_42__31_, u5_mult_87_CARRYB_42__32_,
         u5_mult_87_CARRYB_42__33_, u5_mult_87_CARRYB_42__34_,
         u5_mult_87_CARRYB_42__35_, u5_mult_87_CARRYB_42__36_,
         u5_mult_87_CARRYB_42__37_, u5_mult_87_CARRYB_42__38_,
         u5_mult_87_CARRYB_42__39_, u5_mult_87_CARRYB_42__40_,
         u5_mult_87_CARRYB_42__41_, u5_mult_87_CARRYB_42__42_,
         u5_mult_87_CARRYB_42__43_, u5_mult_87_CARRYB_42__44_,
         u5_mult_87_CARRYB_42__45_, u5_mult_87_CARRYB_42__46_,
         u5_mult_87_CARRYB_42__47_, u5_mult_87_CARRYB_42__48_,
         u5_mult_87_CARRYB_42__49_, u5_mult_87_CARRYB_42__50_,
         u5_mult_87_CARRYB_42__51_, u5_mult_87_CARRYB_43__0_,
         u5_mult_87_CARRYB_43__1_, u5_mult_87_CARRYB_43__2_,
         u5_mult_87_CARRYB_43__3_, u5_mult_87_CARRYB_43__4_,
         u5_mult_87_CARRYB_43__5_, u5_mult_87_CARRYB_43__6_,
         u5_mult_87_CARRYB_43__7_, u5_mult_87_CARRYB_43__8_,
         u5_mult_87_CARRYB_43__9_, u5_mult_87_CARRYB_43__10_,
         u5_mult_87_CARRYB_43__11_, u5_mult_87_CARRYB_43__12_,
         u5_mult_87_CARRYB_43__13_, u5_mult_87_CARRYB_43__14_,
         u5_mult_87_CARRYB_43__15_, u5_mult_87_CARRYB_43__16_,
         u5_mult_87_CARRYB_43__17_, u5_mult_87_SUMB_24__1_,
         u5_mult_87_SUMB_24__2_, u5_mult_87_SUMB_24__3_,
         u5_mult_87_SUMB_24__4_, u5_mult_87_SUMB_24__5_,
         u5_mult_87_SUMB_24__6_, u5_mult_87_SUMB_24__7_,
         u5_mult_87_SUMB_24__8_, u5_mult_87_SUMB_24__9_,
         u5_mult_87_SUMB_24__10_, u5_mult_87_SUMB_24__11_,
         u5_mult_87_SUMB_24__12_, u5_mult_87_SUMB_24__13_,
         u5_mult_87_SUMB_24__14_, u5_mult_87_SUMB_24__15_,
         u5_mult_87_SUMB_24__16_, u5_mult_87_SUMB_24__17_,
         u5_mult_87_SUMB_24__18_, u5_mult_87_SUMB_24__19_,
         u5_mult_87_SUMB_24__20_, u5_mult_87_SUMB_24__21_,
         u5_mult_87_SUMB_24__22_, u5_mult_87_SUMB_24__23_,
         u5_mult_87_SUMB_24__24_, u5_mult_87_SUMB_24__25_,
         u5_mult_87_SUMB_24__26_, u5_mult_87_SUMB_24__27_,
         u5_mult_87_SUMB_24__28_, u5_mult_87_SUMB_24__29_,
         u5_mult_87_SUMB_24__30_, u5_mult_87_SUMB_24__31_,
         u5_mult_87_SUMB_24__32_, u5_mult_87_SUMB_24__33_,
         u5_mult_87_SUMB_24__34_, u5_mult_87_SUMB_24__35_,
         u5_mult_87_SUMB_24__36_, u5_mult_87_SUMB_24__37_,
         u5_mult_87_SUMB_24__38_, u5_mult_87_SUMB_24__39_,
         u5_mult_87_SUMB_24__40_, u5_mult_87_SUMB_24__41_,
         u5_mult_87_SUMB_24__42_, u5_mult_87_SUMB_24__43_,
         u5_mult_87_SUMB_24__44_, u5_mult_87_SUMB_24__45_,
         u5_mult_87_SUMB_24__46_, u5_mult_87_SUMB_24__47_,
         u5_mult_87_SUMB_24__48_, u5_mult_87_SUMB_24__49_,
         u5_mult_87_SUMB_24__50_, u5_mult_87_SUMB_24__51_,
         u5_mult_87_SUMB_25__1_, u5_mult_87_SUMB_25__2_,
         u5_mult_87_SUMB_25__3_, u5_mult_87_SUMB_25__4_,
         u5_mult_87_SUMB_25__5_, u5_mult_87_SUMB_25__6_,
         u5_mult_87_SUMB_25__7_, u5_mult_87_SUMB_25__8_,
         u5_mult_87_SUMB_25__9_, u5_mult_87_SUMB_25__10_,
         u5_mult_87_SUMB_25__11_, u5_mult_87_SUMB_25__12_,
         u5_mult_87_SUMB_25__13_, u5_mult_87_SUMB_25__14_,
         u5_mult_87_SUMB_25__15_, u5_mult_87_SUMB_25__16_,
         u5_mult_87_SUMB_25__17_, u5_mult_87_SUMB_25__18_,
         u5_mult_87_SUMB_25__19_, u5_mult_87_SUMB_25__20_,
         u5_mult_87_SUMB_25__21_, u5_mult_87_SUMB_25__22_,
         u5_mult_87_SUMB_25__23_, u5_mult_87_SUMB_25__24_,
         u5_mult_87_SUMB_25__25_, u5_mult_87_SUMB_25__26_,
         u5_mult_87_SUMB_25__27_, u5_mult_87_SUMB_25__28_,
         u5_mult_87_SUMB_25__29_, u5_mult_87_SUMB_25__30_,
         u5_mult_87_SUMB_25__31_, u5_mult_87_SUMB_25__32_,
         u5_mult_87_SUMB_25__33_, u5_mult_87_SUMB_25__34_,
         u5_mult_87_SUMB_25__35_, u5_mult_87_SUMB_25__36_,
         u5_mult_87_SUMB_25__37_, u5_mult_87_SUMB_25__38_,
         u5_mult_87_SUMB_25__39_, u5_mult_87_SUMB_25__40_,
         u5_mult_87_SUMB_25__41_, u5_mult_87_SUMB_25__42_,
         u5_mult_87_SUMB_25__43_, u5_mult_87_SUMB_25__44_,
         u5_mult_87_SUMB_25__45_, u5_mult_87_SUMB_25__46_,
         u5_mult_87_SUMB_25__47_, u5_mult_87_SUMB_25__48_,
         u5_mult_87_SUMB_25__49_, u5_mult_87_SUMB_25__50_,
         u5_mult_87_SUMB_25__51_, u5_mult_87_SUMB_26__1_,
         u5_mult_87_SUMB_26__2_, u5_mult_87_SUMB_26__3_,
         u5_mult_87_SUMB_26__4_, u5_mult_87_SUMB_26__5_,
         u5_mult_87_SUMB_26__6_, u5_mult_87_SUMB_26__7_,
         u5_mult_87_SUMB_26__8_, u5_mult_87_SUMB_26__9_,
         u5_mult_87_SUMB_26__10_, u5_mult_87_SUMB_26__11_,
         u5_mult_87_SUMB_26__12_, u5_mult_87_SUMB_26__13_,
         u5_mult_87_SUMB_26__14_, u5_mult_87_SUMB_26__15_,
         u5_mult_87_SUMB_26__16_, u5_mult_87_SUMB_26__17_,
         u5_mult_87_SUMB_26__18_, u5_mult_87_SUMB_26__19_,
         u5_mult_87_SUMB_26__20_, u5_mult_87_SUMB_26__21_,
         u5_mult_87_SUMB_26__22_, u5_mult_87_SUMB_26__23_,
         u5_mult_87_SUMB_26__24_, u5_mult_87_SUMB_26__25_,
         u5_mult_87_SUMB_26__26_, u5_mult_87_SUMB_26__27_,
         u5_mult_87_SUMB_26__28_, u5_mult_87_SUMB_26__29_,
         u5_mult_87_SUMB_26__30_, u5_mult_87_SUMB_26__31_,
         u5_mult_87_SUMB_26__32_, u5_mult_87_SUMB_26__33_,
         u5_mult_87_SUMB_26__34_, u5_mult_87_SUMB_26__35_,
         u5_mult_87_SUMB_26__36_, u5_mult_87_SUMB_26__37_,
         u5_mult_87_SUMB_26__38_, u5_mult_87_SUMB_26__39_,
         u5_mult_87_SUMB_26__40_, u5_mult_87_SUMB_26__41_,
         u5_mult_87_SUMB_26__42_, u5_mult_87_SUMB_26__43_,
         u5_mult_87_SUMB_26__44_, u5_mult_87_SUMB_26__45_,
         u5_mult_87_SUMB_26__46_, u5_mult_87_SUMB_26__47_,
         u5_mult_87_SUMB_26__48_, u5_mult_87_SUMB_26__49_,
         u5_mult_87_SUMB_26__50_, u5_mult_87_SUMB_26__51_,
         u5_mult_87_SUMB_27__1_, u5_mult_87_SUMB_27__2_,
         u5_mult_87_SUMB_27__3_, u5_mult_87_SUMB_27__4_,
         u5_mult_87_SUMB_27__5_, u5_mult_87_SUMB_27__6_,
         u5_mult_87_SUMB_27__7_, u5_mult_87_SUMB_27__8_,
         u5_mult_87_SUMB_27__9_, u5_mult_87_SUMB_27__10_,
         u5_mult_87_SUMB_27__11_, u5_mult_87_SUMB_27__12_,
         u5_mult_87_SUMB_27__13_, u5_mult_87_SUMB_27__14_,
         u5_mult_87_SUMB_27__15_, u5_mult_87_SUMB_27__16_,
         u5_mult_87_SUMB_27__17_, u5_mult_87_SUMB_27__18_,
         u5_mult_87_SUMB_27__19_, u5_mult_87_SUMB_27__20_,
         u5_mult_87_SUMB_27__21_, u5_mult_87_SUMB_27__22_,
         u5_mult_87_SUMB_27__23_, u5_mult_87_SUMB_27__24_,
         u5_mult_87_SUMB_27__25_, u5_mult_87_SUMB_27__26_,
         u5_mult_87_SUMB_27__27_, u5_mult_87_SUMB_27__28_,
         u5_mult_87_SUMB_27__29_, u5_mult_87_SUMB_27__30_,
         u5_mult_87_SUMB_27__31_, u5_mult_87_SUMB_27__32_,
         u5_mult_87_SUMB_27__33_, u5_mult_87_SUMB_27__34_,
         u5_mult_87_SUMB_27__35_, u5_mult_87_SUMB_27__36_,
         u5_mult_87_SUMB_27__37_, u5_mult_87_SUMB_27__38_,
         u5_mult_87_SUMB_27__39_, u5_mult_87_SUMB_27__40_,
         u5_mult_87_SUMB_27__41_, u5_mult_87_SUMB_27__42_,
         u5_mult_87_SUMB_27__43_, u5_mult_87_SUMB_27__44_,
         u5_mult_87_SUMB_27__45_, u5_mult_87_SUMB_27__46_,
         u5_mult_87_SUMB_27__47_, u5_mult_87_SUMB_27__48_,
         u5_mult_87_SUMB_27__49_, u5_mult_87_SUMB_27__50_,
         u5_mult_87_SUMB_27__51_, u5_mult_87_SUMB_28__1_,
         u5_mult_87_SUMB_28__2_, u5_mult_87_SUMB_28__3_,
         u5_mult_87_SUMB_28__4_, u5_mult_87_SUMB_28__5_,
         u5_mult_87_SUMB_28__6_, u5_mult_87_SUMB_28__7_,
         u5_mult_87_SUMB_28__8_, u5_mult_87_SUMB_28__9_,
         u5_mult_87_SUMB_28__10_, u5_mult_87_SUMB_28__11_,
         u5_mult_87_SUMB_28__12_, u5_mult_87_SUMB_28__13_,
         u5_mult_87_SUMB_28__14_, u5_mult_87_SUMB_28__15_,
         u5_mult_87_SUMB_28__16_, u5_mult_87_SUMB_28__17_,
         u5_mult_87_SUMB_28__18_, u5_mult_87_SUMB_28__19_,
         u5_mult_87_SUMB_28__20_, u5_mult_87_SUMB_28__21_,
         u5_mult_87_SUMB_28__22_, u5_mult_87_SUMB_28__23_,
         u5_mult_87_SUMB_28__24_, u5_mult_87_SUMB_28__25_,
         u5_mult_87_SUMB_28__26_, u5_mult_87_SUMB_28__27_,
         u5_mult_87_SUMB_28__28_, u5_mult_87_SUMB_28__29_,
         u5_mult_87_SUMB_28__30_, u5_mult_87_SUMB_28__31_,
         u5_mult_87_SUMB_28__32_, u5_mult_87_SUMB_28__33_,
         u5_mult_87_SUMB_28__34_, u5_mult_87_SUMB_28__35_,
         u5_mult_87_SUMB_28__36_, u5_mult_87_SUMB_28__37_,
         u5_mult_87_SUMB_28__38_, u5_mult_87_SUMB_28__39_,
         u5_mult_87_SUMB_28__40_, u5_mult_87_SUMB_28__41_,
         u5_mult_87_SUMB_28__42_, u5_mult_87_SUMB_28__43_,
         u5_mult_87_SUMB_28__44_, u5_mult_87_SUMB_28__45_,
         u5_mult_87_SUMB_28__46_, u5_mult_87_SUMB_28__47_,
         u5_mult_87_SUMB_28__48_, u5_mult_87_SUMB_28__49_,
         u5_mult_87_SUMB_28__50_, u5_mult_87_SUMB_28__51_,
         u5_mult_87_SUMB_29__1_, u5_mult_87_SUMB_29__2_,
         u5_mult_87_SUMB_29__3_, u5_mult_87_SUMB_29__4_,
         u5_mult_87_SUMB_29__5_, u5_mult_87_SUMB_29__6_,
         u5_mult_87_SUMB_29__7_, u5_mult_87_SUMB_29__8_,
         u5_mult_87_SUMB_29__9_, u5_mult_87_SUMB_29__10_,
         u5_mult_87_SUMB_29__11_, u5_mult_87_SUMB_29__12_,
         u5_mult_87_SUMB_29__13_, u5_mult_87_SUMB_29__14_,
         u5_mult_87_SUMB_29__15_, u5_mult_87_SUMB_29__16_,
         u5_mult_87_SUMB_29__17_, u5_mult_87_SUMB_29__18_,
         u5_mult_87_SUMB_29__19_, u5_mult_87_SUMB_29__20_,
         u5_mult_87_SUMB_29__21_, u5_mult_87_SUMB_29__22_,
         u5_mult_87_SUMB_29__23_, u5_mult_87_SUMB_29__24_,
         u5_mult_87_SUMB_29__25_, u5_mult_87_SUMB_29__26_,
         u5_mult_87_SUMB_29__27_, u5_mult_87_SUMB_29__28_,
         u5_mult_87_SUMB_29__29_, u5_mult_87_SUMB_29__30_,
         u5_mult_87_SUMB_29__31_, u5_mult_87_SUMB_29__32_,
         u5_mult_87_SUMB_29__33_, u5_mult_87_SUMB_29__34_,
         u5_mult_87_SUMB_29__35_, u5_mult_87_SUMB_29__36_,
         u5_mult_87_SUMB_29__37_, u5_mult_87_SUMB_29__38_,
         u5_mult_87_SUMB_29__39_, u5_mult_87_SUMB_29__40_,
         u5_mult_87_SUMB_29__41_, u5_mult_87_SUMB_29__42_,
         u5_mult_87_SUMB_29__43_, u5_mult_87_SUMB_29__44_,
         u5_mult_87_SUMB_29__45_, u5_mult_87_SUMB_29__46_,
         u5_mult_87_SUMB_29__47_, u5_mult_87_SUMB_29__48_,
         u5_mult_87_SUMB_29__49_, u5_mult_87_SUMB_29__50_,
         u5_mult_87_SUMB_29__51_, u5_mult_87_SUMB_30__1_,
         u5_mult_87_SUMB_30__2_, u5_mult_87_SUMB_30__3_,
         u5_mult_87_SUMB_30__4_, u5_mult_87_SUMB_30__5_,
         u5_mult_87_SUMB_30__6_, u5_mult_87_SUMB_30__7_,
         u5_mult_87_SUMB_30__8_, u5_mult_87_SUMB_30__9_,
         u5_mult_87_SUMB_30__10_, u5_mult_87_SUMB_30__11_,
         u5_mult_87_SUMB_30__12_, u5_mult_87_SUMB_30__13_,
         u5_mult_87_SUMB_30__14_, u5_mult_87_SUMB_30__15_,
         u5_mult_87_SUMB_30__16_, u5_mult_87_SUMB_30__17_,
         u5_mult_87_SUMB_30__18_, u5_mult_87_SUMB_30__19_,
         u5_mult_87_SUMB_30__20_, u5_mult_87_SUMB_30__21_,
         u5_mult_87_SUMB_30__22_, u5_mult_87_SUMB_30__23_,
         u5_mult_87_SUMB_30__24_, u5_mult_87_SUMB_30__25_,
         u5_mult_87_SUMB_30__26_, u5_mult_87_SUMB_30__27_,
         u5_mult_87_SUMB_30__28_, u5_mult_87_SUMB_30__29_,
         u5_mult_87_SUMB_30__30_, u5_mult_87_SUMB_30__31_,
         u5_mult_87_SUMB_30__32_, u5_mult_87_SUMB_30__33_,
         u5_mult_87_SUMB_30__34_, u5_mult_87_SUMB_30__35_,
         u5_mult_87_SUMB_30__36_, u5_mult_87_SUMB_30__37_,
         u5_mult_87_SUMB_30__38_, u5_mult_87_SUMB_30__39_,
         u5_mult_87_SUMB_30__40_, u5_mult_87_SUMB_30__41_,
         u5_mult_87_SUMB_30__42_, u5_mult_87_SUMB_30__43_,
         u5_mult_87_SUMB_30__44_, u5_mult_87_SUMB_30__45_,
         u5_mult_87_SUMB_30__46_, u5_mult_87_SUMB_30__47_,
         u5_mult_87_SUMB_30__48_, u5_mult_87_SUMB_30__49_,
         u5_mult_87_SUMB_30__50_, u5_mult_87_SUMB_30__51_,
         u5_mult_87_SUMB_31__1_, u5_mult_87_SUMB_31__2_,
         u5_mult_87_SUMB_31__3_, u5_mult_87_SUMB_31__4_,
         u5_mult_87_SUMB_31__5_, u5_mult_87_SUMB_31__6_,
         u5_mult_87_SUMB_31__7_, u5_mult_87_SUMB_31__8_,
         u5_mult_87_SUMB_31__9_, u5_mult_87_SUMB_31__10_,
         u5_mult_87_SUMB_31__11_, u5_mult_87_SUMB_31__12_,
         u5_mult_87_SUMB_31__13_, u5_mult_87_SUMB_31__14_,
         u5_mult_87_SUMB_31__15_, u5_mult_87_SUMB_31__16_,
         u5_mult_87_SUMB_31__17_, u5_mult_87_SUMB_31__18_,
         u5_mult_87_SUMB_31__19_, u5_mult_87_SUMB_31__20_,
         u5_mult_87_SUMB_31__21_, u5_mult_87_SUMB_31__22_,
         u5_mult_87_SUMB_31__23_, u5_mult_87_SUMB_31__24_,
         u5_mult_87_SUMB_31__25_, u5_mult_87_SUMB_31__26_,
         u5_mult_87_SUMB_31__27_, u5_mult_87_SUMB_31__28_,
         u5_mult_87_SUMB_31__29_, u5_mult_87_SUMB_31__30_,
         u5_mult_87_SUMB_31__31_, u5_mult_87_SUMB_31__32_,
         u5_mult_87_SUMB_31__33_, u5_mult_87_SUMB_31__34_,
         u5_mult_87_SUMB_31__35_, u5_mult_87_SUMB_31__36_,
         u5_mult_87_SUMB_31__37_, u5_mult_87_SUMB_31__38_,
         u5_mult_87_SUMB_31__39_, u5_mult_87_SUMB_31__40_,
         u5_mult_87_SUMB_31__41_, u5_mult_87_SUMB_31__42_,
         u5_mult_87_SUMB_31__43_, u5_mult_87_SUMB_31__44_,
         u5_mult_87_SUMB_31__45_, u5_mult_87_SUMB_31__46_,
         u5_mult_87_SUMB_31__47_, u5_mult_87_SUMB_31__48_,
         u5_mult_87_SUMB_31__49_, u5_mult_87_SUMB_31__50_,
         u5_mult_87_SUMB_31__51_, u5_mult_87_SUMB_32__1_,
         u5_mult_87_SUMB_32__2_, u5_mult_87_SUMB_32__3_,
         u5_mult_87_SUMB_32__4_, u5_mult_87_SUMB_32__5_,
         u5_mult_87_SUMB_32__6_, u5_mult_87_SUMB_32__7_,
         u5_mult_87_SUMB_32__8_, u5_mult_87_SUMB_32__9_,
         u5_mult_87_SUMB_32__10_, u5_mult_87_SUMB_32__11_,
         u5_mult_87_SUMB_32__12_, u5_mult_87_SUMB_32__13_,
         u5_mult_87_SUMB_32__14_, u5_mult_87_SUMB_32__15_,
         u5_mult_87_SUMB_32__16_, u5_mult_87_SUMB_32__17_,
         u5_mult_87_SUMB_32__18_, u5_mult_87_SUMB_32__19_,
         u5_mult_87_SUMB_32__20_, u5_mult_87_SUMB_32__21_,
         u5_mult_87_SUMB_32__22_, u5_mult_87_SUMB_32__23_,
         u5_mult_87_SUMB_32__24_, u5_mult_87_SUMB_32__25_,
         u5_mult_87_SUMB_32__26_, u5_mult_87_SUMB_32__27_,
         u5_mult_87_SUMB_32__28_, u5_mult_87_SUMB_32__29_,
         u5_mult_87_SUMB_32__30_, u5_mult_87_SUMB_32__31_,
         u5_mult_87_SUMB_32__32_, u5_mult_87_SUMB_32__33_,
         u5_mult_87_SUMB_32__34_, u5_mult_87_SUMB_32__35_,
         u5_mult_87_SUMB_32__36_, u5_mult_87_SUMB_32__37_,
         u5_mult_87_SUMB_32__38_, u5_mult_87_SUMB_32__39_,
         u5_mult_87_SUMB_32__40_, u5_mult_87_SUMB_32__41_,
         u5_mult_87_SUMB_32__42_, u5_mult_87_SUMB_32__43_,
         u5_mult_87_SUMB_32__44_, u5_mult_87_SUMB_32__45_,
         u5_mult_87_SUMB_32__46_, u5_mult_87_SUMB_32__47_,
         u5_mult_87_SUMB_32__48_, u5_mult_87_SUMB_32__49_,
         u5_mult_87_SUMB_32__50_, u5_mult_87_SUMB_32__51_,
         u5_mult_87_SUMB_33__1_, u5_mult_87_SUMB_33__2_,
         u5_mult_87_SUMB_33__3_, u5_mult_87_SUMB_33__4_,
         u5_mult_87_SUMB_33__5_, u5_mult_87_SUMB_33__6_,
         u5_mult_87_SUMB_33__7_, u5_mult_87_SUMB_33__8_,
         u5_mult_87_SUMB_33__9_, u5_mult_87_SUMB_33__10_,
         u5_mult_87_SUMB_33__11_, u5_mult_87_SUMB_33__12_,
         u5_mult_87_SUMB_33__13_, u5_mult_87_SUMB_33__14_,
         u5_mult_87_SUMB_33__15_, u5_mult_87_SUMB_33__16_,
         u5_mult_87_SUMB_33__17_, u5_mult_87_SUMB_33__18_,
         u5_mult_87_SUMB_33__19_, u5_mult_87_SUMB_33__20_,
         u5_mult_87_SUMB_33__21_, u5_mult_87_SUMB_33__22_,
         u5_mult_87_SUMB_33__23_, u5_mult_87_SUMB_33__24_,
         u5_mult_87_SUMB_33__25_, u5_mult_87_SUMB_33__26_,
         u5_mult_87_SUMB_33__27_, u5_mult_87_SUMB_33__28_,
         u5_mult_87_SUMB_33__29_, u5_mult_87_SUMB_33__30_,
         u5_mult_87_SUMB_33__31_, u5_mult_87_SUMB_33__32_,
         u5_mult_87_SUMB_33__33_, u5_mult_87_SUMB_33__34_,
         u5_mult_87_SUMB_33__35_, u5_mult_87_CARRYB_24__1_,
         u5_mult_87_CARRYB_24__2_, u5_mult_87_CARRYB_24__3_,
         u5_mult_87_CARRYB_24__4_, u5_mult_87_CARRYB_24__5_,
         u5_mult_87_CARRYB_24__6_, u5_mult_87_CARRYB_24__7_,
         u5_mult_87_CARRYB_24__8_, u5_mult_87_CARRYB_24__9_,
         u5_mult_87_CARRYB_24__10_, u5_mult_87_CARRYB_24__11_,
         u5_mult_87_CARRYB_24__12_, u5_mult_87_CARRYB_24__13_,
         u5_mult_87_CARRYB_24__14_, u5_mult_87_CARRYB_24__15_,
         u5_mult_87_CARRYB_24__16_, u5_mult_87_CARRYB_24__17_,
         u5_mult_87_CARRYB_24__18_, u5_mult_87_CARRYB_24__19_,
         u5_mult_87_CARRYB_24__20_, u5_mult_87_CARRYB_24__21_,
         u5_mult_87_CARRYB_24__22_, u5_mult_87_CARRYB_24__23_,
         u5_mult_87_CARRYB_24__24_, u5_mult_87_CARRYB_24__25_,
         u5_mult_87_CARRYB_24__26_, u5_mult_87_CARRYB_24__27_,
         u5_mult_87_CARRYB_24__28_, u5_mult_87_CARRYB_24__29_,
         u5_mult_87_CARRYB_24__30_, u5_mult_87_CARRYB_24__31_,
         u5_mult_87_CARRYB_24__32_, u5_mult_87_CARRYB_24__33_,
         u5_mult_87_CARRYB_24__34_, u5_mult_87_CARRYB_24__35_,
         u5_mult_87_CARRYB_24__36_, u5_mult_87_CARRYB_24__37_,
         u5_mult_87_CARRYB_24__38_, u5_mult_87_CARRYB_24__39_,
         u5_mult_87_CARRYB_24__40_, u5_mult_87_CARRYB_24__41_,
         u5_mult_87_CARRYB_24__42_, u5_mult_87_CARRYB_24__43_,
         u5_mult_87_CARRYB_24__44_, u5_mult_87_CARRYB_24__45_,
         u5_mult_87_CARRYB_24__46_, u5_mult_87_CARRYB_24__47_,
         u5_mult_87_CARRYB_24__48_, u5_mult_87_CARRYB_24__49_,
         u5_mult_87_CARRYB_24__50_, u5_mult_87_CARRYB_24__51_,
         u5_mult_87_CARRYB_25__0_, u5_mult_87_CARRYB_25__1_,
         u5_mult_87_CARRYB_25__2_, u5_mult_87_CARRYB_25__3_,
         u5_mult_87_CARRYB_25__4_, u5_mult_87_CARRYB_25__5_,
         u5_mult_87_CARRYB_25__6_, u5_mult_87_CARRYB_25__7_,
         u5_mult_87_CARRYB_25__8_, u5_mult_87_CARRYB_25__9_,
         u5_mult_87_CARRYB_25__10_, u5_mult_87_CARRYB_25__11_,
         u5_mult_87_CARRYB_25__12_, u5_mult_87_CARRYB_25__13_,
         u5_mult_87_CARRYB_25__14_, u5_mult_87_CARRYB_25__15_,
         u5_mult_87_CARRYB_25__16_, u5_mult_87_CARRYB_25__17_,
         u5_mult_87_CARRYB_25__18_, u5_mult_87_CARRYB_25__19_,
         u5_mult_87_CARRYB_25__20_, u5_mult_87_CARRYB_25__21_,
         u5_mult_87_CARRYB_25__22_, u5_mult_87_CARRYB_25__23_,
         u5_mult_87_CARRYB_25__24_, u5_mult_87_CARRYB_25__25_,
         u5_mult_87_CARRYB_25__26_, u5_mult_87_CARRYB_25__27_,
         u5_mult_87_CARRYB_25__28_, u5_mult_87_CARRYB_25__29_,
         u5_mult_87_CARRYB_25__30_, u5_mult_87_CARRYB_25__31_,
         u5_mult_87_CARRYB_25__32_, u5_mult_87_CARRYB_25__33_,
         u5_mult_87_CARRYB_25__34_, u5_mult_87_CARRYB_25__35_,
         u5_mult_87_CARRYB_25__36_, u5_mult_87_CARRYB_25__37_,
         u5_mult_87_CARRYB_25__38_, u5_mult_87_CARRYB_25__39_,
         u5_mult_87_CARRYB_25__40_, u5_mult_87_CARRYB_25__41_,
         u5_mult_87_CARRYB_25__42_, u5_mult_87_CARRYB_25__43_,
         u5_mult_87_CARRYB_25__44_, u5_mult_87_CARRYB_25__45_,
         u5_mult_87_CARRYB_25__46_, u5_mult_87_CARRYB_25__47_,
         u5_mult_87_CARRYB_25__48_, u5_mult_87_CARRYB_25__49_,
         u5_mult_87_CARRYB_25__50_, u5_mult_87_CARRYB_25__51_,
         u5_mult_87_CARRYB_26__0_, u5_mult_87_CARRYB_26__1_,
         u5_mult_87_CARRYB_26__2_, u5_mult_87_CARRYB_26__3_,
         u5_mult_87_CARRYB_26__4_, u5_mult_87_CARRYB_26__5_,
         u5_mult_87_CARRYB_26__6_, u5_mult_87_CARRYB_26__7_,
         u5_mult_87_CARRYB_26__8_, u5_mult_87_CARRYB_26__9_,
         u5_mult_87_CARRYB_26__10_, u5_mult_87_CARRYB_26__11_,
         u5_mult_87_CARRYB_26__12_, u5_mult_87_CARRYB_26__13_,
         u5_mult_87_CARRYB_26__14_, u5_mult_87_CARRYB_26__15_,
         u5_mult_87_CARRYB_26__16_, u5_mult_87_CARRYB_26__17_,
         u5_mult_87_CARRYB_26__18_, u5_mult_87_CARRYB_26__19_,
         u5_mult_87_CARRYB_26__20_, u5_mult_87_CARRYB_26__21_,
         u5_mult_87_CARRYB_26__22_, u5_mult_87_CARRYB_26__23_,
         u5_mult_87_CARRYB_26__24_, u5_mult_87_CARRYB_26__25_,
         u5_mult_87_CARRYB_26__26_, u5_mult_87_CARRYB_26__27_,
         u5_mult_87_CARRYB_26__28_, u5_mult_87_CARRYB_26__29_,
         u5_mult_87_CARRYB_26__30_, u5_mult_87_CARRYB_26__31_,
         u5_mult_87_CARRYB_26__32_, u5_mult_87_CARRYB_26__33_,
         u5_mult_87_CARRYB_26__34_, u5_mult_87_CARRYB_26__35_,
         u5_mult_87_CARRYB_26__36_, u5_mult_87_CARRYB_26__37_,
         u5_mult_87_CARRYB_26__38_, u5_mult_87_CARRYB_26__39_,
         u5_mult_87_CARRYB_26__40_, u5_mult_87_CARRYB_26__41_,
         u5_mult_87_CARRYB_26__42_, u5_mult_87_CARRYB_26__43_,
         u5_mult_87_CARRYB_26__44_, u5_mult_87_CARRYB_26__45_,
         u5_mult_87_CARRYB_26__46_, u5_mult_87_CARRYB_26__47_,
         u5_mult_87_CARRYB_26__48_, u5_mult_87_CARRYB_26__49_,
         u5_mult_87_CARRYB_26__50_, u5_mult_87_CARRYB_26__51_,
         u5_mult_87_CARRYB_27__0_, u5_mult_87_CARRYB_27__1_,
         u5_mult_87_CARRYB_27__2_, u5_mult_87_CARRYB_27__3_,
         u5_mult_87_CARRYB_27__4_, u5_mult_87_CARRYB_27__5_,
         u5_mult_87_CARRYB_27__6_, u5_mult_87_CARRYB_27__7_,
         u5_mult_87_CARRYB_27__8_, u5_mult_87_CARRYB_27__9_,
         u5_mult_87_CARRYB_27__10_, u5_mult_87_CARRYB_27__11_,
         u5_mult_87_CARRYB_27__12_, u5_mult_87_CARRYB_27__13_,
         u5_mult_87_CARRYB_27__14_, u5_mult_87_CARRYB_27__15_,
         u5_mult_87_CARRYB_27__16_, u5_mult_87_CARRYB_27__17_,
         u5_mult_87_CARRYB_27__18_, u5_mult_87_CARRYB_27__19_,
         u5_mult_87_CARRYB_27__20_, u5_mult_87_CARRYB_27__21_,
         u5_mult_87_CARRYB_27__22_, u5_mult_87_CARRYB_27__23_,
         u5_mult_87_CARRYB_27__24_, u5_mult_87_CARRYB_27__25_,
         u5_mult_87_CARRYB_27__26_, u5_mult_87_CARRYB_27__27_,
         u5_mult_87_CARRYB_27__28_, u5_mult_87_CARRYB_27__29_,
         u5_mult_87_CARRYB_27__30_, u5_mult_87_CARRYB_27__31_,
         u5_mult_87_CARRYB_27__32_, u5_mult_87_CARRYB_27__33_,
         u5_mult_87_CARRYB_27__34_, u5_mult_87_CARRYB_27__35_,
         u5_mult_87_CARRYB_27__36_, u5_mult_87_CARRYB_27__37_,
         u5_mult_87_CARRYB_27__38_, u5_mult_87_CARRYB_27__39_,
         u5_mult_87_CARRYB_27__40_, u5_mult_87_CARRYB_27__41_,
         u5_mult_87_CARRYB_27__42_, u5_mult_87_CARRYB_27__43_,
         u5_mult_87_CARRYB_27__44_, u5_mult_87_CARRYB_27__45_,
         u5_mult_87_CARRYB_27__46_, u5_mult_87_CARRYB_27__47_,
         u5_mult_87_CARRYB_27__48_, u5_mult_87_CARRYB_27__49_,
         u5_mult_87_CARRYB_27__50_, u5_mult_87_CARRYB_27__51_,
         u5_mult_87_CARRYB_28__0_, u5_mult_87_CARRYB_28__1_,
         u5_mult_87_CARRYB_28__2_, u5_mult_87_CARRYB_28__3_,
         u5_mult_87_CARRYB_28__4_, u5_mult_87_CARRYB_28__5_,
         u5_mult_87_CARRYB_28__6_, u5_mult_87_CARRYB_28__7_,
         u5_mult_87_CARRYB_28__8_, u5_mult_87_CARRYB_28__9_,
         u5_mult_87_CARRYB_28__10_, u5_mult_87_CARRYB_28__11_,
         u5_mult_87_CARRYB_28__12_, u5_mult_87_CARRYB_28__13_,
         u5_mult_87_CARRYB_28__14_, u5_mult_87_CARRYB_28__15_,
         u5_mult_87_CARRYB_28__16_, u5_mult_87_CARRYB_28__17_,
         u5_mult_87_CARRYB_28__18_, u5_mult_87_CARRYB_28__19_,
         u5_mult_87_CARRYB_28__20_, u5_mult_87_CARRYB_28__21_,
         u5_mult_87_CARRYB_28__22_, u5_mult_87_CARRYB_28__23_,
         u5_mult_87_CARRYB_28__24_, u5_mult_87_CARRYB_28__25_,
         u5_mult_87_CARRYB_28__26_, u5_mult_87_CARRYB_28__27_,
         u5_mult_87_CARRYB_28__28_, u5_mult_87_CARRYB_28__29_,
         u5_mult_87_CARRYB_28__30_, u5_mult_87_CARRYB_28__31_,
         u5_mult_87_CARRYB_28__32_, u5_mult_87_CARRYB_28__33_,
         u5_mult_87_CARRYB_28__34_, u5_mult_87_CARRYB_28__35_,
         u5_mult_87_CARRYB_28__36_, u5_mult_87_CARRYB_28__37_,
         u5_mult_87_CARRYB_28__38_, u5_mult_87_CARRYB_28__39_,
         u5_mult_87_CARRYB_28__40_, u5_mult_87_CARRYB_28__41_,
         u5_mult_87_CARRYB_28__42_, u5_mult_87_CARRYB_28__43_,
         u5_mult_87_CARRYB_28__44_, u5_mult_87_CARRYB_28__45_,
         u5_mult_87_CARRYB_28__46_, u5_mult_87_CARRYB_28__47_,
         u5_mult_87_CARRYB_28__48_, u5_mult_87_CARRYB_28__49_,
         u5_mult_87_CARRYB_28__50_, u5_mult_87_CARRYB_28__51_,
         u5_mult_87_CARRYB_29__0_, u5_mult_87_CARRYB_29__1_,
         u5_mult_87_CARRYB_29__2_, u5_mult_87_CARRYB_29__3_,
         u5_mult_87_CARRYB_29__4_, u5_mult_87_CARRYB_29__5_,
         u5_mult_87_CARRYB_29__6_, u5_mult_87_CARRYB_29__7_,
         u5_mult_87_CARRYB_29__8_, u5_mult_87_CARRYB_29__9_,
         u5_mult_87_CARRYB_29__10_, u5_mult_87_CARRYB_29__11_,
         u5_mult_87_CARRYB_29__12_, u5_mult_87_CARRYB_29__13_,
         u5_mult_87_CARRYB_29__14_, u5_mult_87_CARRYB_29__15_,
         u5_mult_87_CARRYB_29__16_, u5_mult_87_CARRYB_29__17_,
         u5_mult_87_CARRYB_29__18_, u5_mult_87_CARRYB_29__19_,
         u5_mult_87_CARRYB_29__20_, u5_mult_87_CARRYB_29__21_,
         u5_mult_87_CARRYB_29__22_, u5_mult_87_CARRYB_29__23_,
         u5_mult_87_CARRYB_29__24_, u5_mult_87_CARRYB_29__25_,
         u5_mult_87_CARRYB_29__26_, u5_mult_87_CARRYB_29__27_,
         u5_mult_87_CARRYB_29__28_, u5_mult_87_CARRYB_29__29_,
         u5_mult_87_CARRYB_29__30_, u5_mult_87_CARRYB_29__31_,
         u5_mult_87_CARRYB_29__32_, u5_mult_87_CARRYB_29__33_,
         u5_mult_87_CARRYB_29__34_, u5_mult_87_CARRYB_29__35_,
         u5_mult_87_CARRYB_29__36_, u5_mult_87_CARRYB_29__37_,
         u5_mult_87_CARRYB_29__38_, u5_mult_87_CARRYB_29__39_,
         u5_mult_87_CARRYB_29__40_, u5_mult_87_CARRYB_29__41_,
         u5_mult_87_CARRYB_29__42_, u5_mult_87_CARRYB_29__43_,
         u5_mult_87_CARRYB_29__44_, u5_mult_87_CARRYB_29__45_,
         u5_mult_87_CARRYB_29__46_, u5_mult_87_CARRYB_29__47_,
         u5_mult_87_CARRYB_29__48_, u5_mult_87_CARRYB_29__49_,
         u5_mult_87_CARRYB_29__50_, u5_mult_87_CARRYB_29__51_,
         u5_mult_87_CARRYB_30__0_, u5_mult_87_CARRYB_30__1_,
         u5_mult_87_CARRYB_30__2_, u5_mult_87_CARRYB_30__3_,
         u5_mult_87_CARRYB_30__4_, u5_mult_87_CARRYB_30__5_,
         u5_mult_87_CARRYB_30__6_, u5_mult_87_CARRYB_30__7_,
         u5_mult_87_CARRYB_30__8_, u5_mult_87_CARRYB_30__9_,
         u5_mult_87_CARRYB_30__10_, u5_mult_87_CARRYB_30__11_,
         u5_mult_87_CARRYB_30__12_, u5_mult_87_CARRYB_30__13_,
         u5_mult_87_CARRYB_30__14_, u5_mult_87_CARRYB_30__15_,
         u5_mult_87_CARRYB_30__16_, u5_mult_87_CARRYB_30__17_,
         u5_mult_87_CARRYB_30__18_, u5_mult_87_CARRYB_30__19_,
         u5_mult_87_CARRYB_30__20_, u5_mult_87_CARRYB_30__21_,
         u5_mult_87_CARRYB_30__22_, u5_mult_87_CARRYB_30__23_,
         u5_mult_87_CARRYB_30__24_, u5_mult_87_CARRYB_30__25_,
         u5_mult_87_CARRYB_30__26_, u5_mult_87_CARRYB_30__27_,
         u5_mult_87_CARRYB_30__28_, u5_mult_87_CARRYB_30__29_,
         u5_mult_87_CARRYB_30__30_, u5_mult_87_CARRYB_30__31_,
         u5_mult_87_CARRYB_30__32_, u5_mult_87_CARRYB_30__33_,
         u5_mult_87_CARRYB_30__34_, u5_mult_87_CARRYB_30__35_,
         u5_mult_87_CARRYB_30__36_, u5_mult_87_CARRYB_30__37_,
         u5_mult_87_CARRYB_30__38_, u5_mult_87_CARRYB_30__39_,
         u5_mult_87_CARRYB_30__40_, u5_mult_87_CARRYB_30__41_,
         u5_mult_87_CARRYB_30__42_, u5_mult_87_CARRYB_30__43_,
         u5_mult_87_CARRYB_30__44_, u5_mult_87_CARRYB_30__45_,
         u5_mult_87_CARRYB_30__46_, u5_mult_87_CARRYB_30__47_,
         u5_mult_87_CARRYB_30__48_, u5_mult_87_CARRYB_30__49_,
         u5_mult_87_CARRYB_30__50_, u5_mult_87_CARRYB_30__51_,
         u5_mult_87_CARRYB_31__0_, u5_mult_87_CARRYB_31__1_,
         u5_mult_87_CARRYB_31__2_, u5_mult_87_CARRYB_31__3_,
         u5_mult_87_CARRYB_31__4_, u5_mult_87_CARRYB_31__5_,
         u5_mult_87_CARRYB_31__6_, u5_mult_87_CARRYB_31__7_,
         u5_mult_87_CARRYB_31__8_, u5_mult_87_CARRYB_31__9_,
         u5_mult_87_CARRYB_31__10_, u5_mult_87_CARRYB_31__11_,
         u5_mult_87_CARRYB_31__12_, u5_mult_87_CARRYB_31__13_,
         u5_mult_87_CARRYB_31__14_, u5_mult_87_CARRYB_31__15_,
         u5_mult_87_CARRYB_31__16_, u5_mult_87_CARRYB_31__17_,
         u5_mult_87_CARRYB_31__18_, u5_mult_87_CARRYB_31__19_,
         u5_mult_87_CARRYB_31__20_, u5_mult_87_CARRYB_31__21_,
         u5_mult_87_CARRYB_31__22_, u5_mult_87_CARRYB_31__23_,
         u5_mult_87_CARRYB_31__24_, u5_mult_87_CARRYB_31__25_,
         u5_mult_87_CARRYB_31__26_, u5_mult_87_CARRYB_31__27_,
         u5_mult_87_CARRYB_31__28_, u5_mult_87_CARRYB_31__29_,
         u5_mult_87_CARRYB_31__30_, u5_mult_87_CARRYB_31__31_,
         u5_mult_87_CARRYB_31__32_, u5_mult_87_CARRYB_31__33_,
         u5_mult_87_CARRYB_31__34_, u5_mult_87_CARRYB_31__35_,
         u5_mult_87_CARRYB_31__36_, u5_mult_87_CARRYB_31__37_,
         u5_mult_87_CARRYB_31__38_, u5_mult_87_CARRYB_31__39_,
         u5_mult_87_CARRYB_31__40_, u5_mult_87_CARRYB_31__41_,
         u5_mult_87_CARRYB_31__42_, u5_mult_87_CARRYB_31__43_,
         u5_mult_87_CARRYB_31__44_, u5_mult_87_CARRYB_31__45_,
         u5_mult_87_CARRYB_31__46_, u5_mult_87_CARRYB_31__47_,
         u5_mult_87_CARRYB_31__48_, u5_mult_87_CARRYB_31__49_,
         u5_mult_87_CARRYB_31__50_, u5_mult_87_CARRYB_31__51_,
         u5_mult_87_CARRYB_32__0_, u5_mult_87_CARRYB_32__1_,
         u5_mult_87_CARRYB_32__2_, u5_mult_87_CARRYB_32__3_,
         u5_mult_87_CARRYB_32__4_, u5_mult_87_CARRYB_32__5_,
         u5_mult_87_CARRYB_32__6_, u5_mult_87_CARRYB_32__7_,
         u5_mult_87_CARRYB_32__8_, u5_mult_87_CARRYB_32__9_,
         u5_mult_87_CARRYB_32__10_, u5_mult_87_CARRYB_32__11_,
         u5_mult_87_CARRYB_32__12_, u5_mult_87_CARRYB_32__13_,
         u5_mult_87_CARRYB_32__14_, u5_mult_87_CARRYB_32__15_,
         u5_mult_87_CARRYB_32__16_, u5_mult_87_CARRYB_32__17_,
         u5_mult_87_CARRYB_32__18_, u5_mult_87_CARRYB_32__19_,
         u5_mult_87_CARRYB_32__20_, u5_mult_87_CARRYB_32__21_,
         u5_mult_87_CARRYB_32__22_, u5_mult_87_CARRYB_32__23_,
         u5_mult_87_CARRYB_32__24_, u5_mult_87_CARRYB_32__25_,
         u5_mult_87_CARRYB_32__26_, u5_mult_87_CARRYB_32__27_,
         u5_mult_87_CARRYB_32__28_, u5_mult_87_CARRYB_32__29_,
         u5_mult_87_CARRYB_32__30_, u5_mult_87_CARRYB_32__31_,
         u5_mult_87_CARRYB_32__32_, u5_mult_87_CARRYB_32__33_,
         u5_mult_87_CARRYB_32__34_, u5_mult_87_CARRYB_32__35_,
         u5_mult_87_CARRYB_32__36_, u5_mult_87_CARRYB_32__37_,
         u5_mult_87_CARRYB_32__38_, u5_mult_87_CARRYB_32__39_,
         u5_mult_87_CARRYB_32__40_, u5_mult_87_CARRYB_32__41_,
         u5_mult_87_CARRYB_32__42_, u5_mult_87_CARRYB_32__43_,
         u5_mult_87_CARRYB_32__44_, u5_mult_87_CARRYB_32__45_,
         u5_mult_87_CARRYB_32__46_, u5_mult_87_CARRYB_32__47_,
         u5_mult_87_CARRYB_32__48_, u5_mult_87_CARRYB_32__49_,
         u5_mult_87_CARRYB_32__50_, u5_mult_87_CARRYB_32__51_,
         u5_mult_87_CARRYB_33__0_, u5_mult_87_CARRYB_33__1_,
         u5_mult_87_CARRYB_33__2_, u5_mult_87_CARRYB_33__3_,
         u5_mult_87_CARRYB_33__4_, u5_mult_87_CARRYB_33__5_,
         u5_mult_87_CARRYB_33__6_, u5_mult_87_CARRYB_33__7_,
         u5_mult_87_CARRYB_33__8_, u5_mult_87_CARRYB_33__9_,
         u5_mult_87_CARRYB_33__10_, u5_mult_87_CARRYB_33__11_,
         u5_mult_87_CARRYB_33__12_, u5_mult_87_CARRYB_33__13_,
         u5_mult_87_CARRYB_33__14_, u5_mult_87_CARRYB_33__15_,
         u5_mult_87_CARRYB_33__16_, u5_mult_87_CARRYB_33__17_,
         u5_mult_87_CARRYB_33__18_, u5_mult_87_CARRYB_33__19_,
         u5_mult_87_CARRYB_33__20_, u5_mult_87_CARRYB_33__21_,
         u5_mult_87_CARRYB_33__22_, u5_mult_87_CARRYB_33__23_,
         u5_mult_87_CARRYB_33__24_, u5_mult_87_CARRYB_33__25_,
         u5_mult_87_CARRYB_33__26_, u5_mult_87_CARRYB_33__27_,
         u5_mult_87_CARRYB_33__28_, u5_mult_87_CARRYB_33__29_,
         u5_mult_87_CARRYB_33__30_, u5_mult_87_CARRYB_33__31_,
         u5_mult_87_CARRYB_33__32_, u5_mult_87_CARRYB_33__33_,
         u5_mult_87_CARRYB_33__34_, u5_mult_87_CARRYB_33__35_,
         u5_mult_87_SUMB_14__19_, u5_mult_87_SUMB_14__20_,
         u5_mult_87_SUMB_14__21_, u5_mult_87_SUMB_14__22_,
         u5_mult_87_SUMB_14__23_, u5_mult_87_SUMB_14__24_,
         u5_mult_87_SUMB_14__25_, u5_mult_87_SUMB_14__26_,
         u5_mult_87_SUMB_14__27_, u5_mult_87_SUMB_14__28_,
         u5_mult_87_SUMB_14__29_, u5_mult_87_SUMB_14__30_,
         u5_mult_87_SUMB_14__31_, u5_mult_87_SUMB_14__32_,
         u5_mult_87_SUMB_14__33_, u5_mult_87_SUMB_14__34_,
         u5_mult_87_SUMB_14__35_, u5_mult_87_SUMB_14__36_,
         u5_mult_87_SUMB_14__37_, u5_mult_87_SUMB_14__38_,
         u5_mult_87_SUMB_14__39_, u5_mult_87_SUMB_14__40_,
         u5_mult_87_SUMB_14__41_, u5_mult_87_SUMB_14__42_,
         u5_mult_87_SUMB_14__43_, u5_mult_87_SUMB_14__44_,
         u5_mult_87_SUMB_14__45_, u5_mult_87_SUMB_14__46_,
         u5_mult_87_SUMB_14__47_, u5_mult_87_SUMB_14__48_,
         u5_mult_87_SUMB_14__49_, u5_mult_87_SUMB_14__50_,
         u5_mult_87_SUMB_14__51_, u5_mult_87_SUMB_15__1_,
         u5_mult_87_SUMB_15__2_, u5_mult_87_SUMB_15__3_,
         u5_mult_87_SUMB_15__4_, u5_mult_87_SUMB_15__5_,
         u5_mult_87_SUMB_15__6_, u5_mult_87_SUMB_15__7_,
         u5_mult_87_SUMB_15__8_, u5_mult_87_SUMB_15__9_,
         u5_mult_87_SUMB_15__10_, u5_mult_87_SUMB_15__11_,
         u5_mult_87_SUMB_15__12_, u5_mult_87_SUMB_15__13_,
         u5_mult_87_SUMB_15__14_, u5_mult_87_SUMB_15__15_,
         u5_mult_87_SUMB_15__16_, u5_mult_87_SUMB_15__17_,
         u5_mult_87_SUMB_15__18_, u5_mult_87_SUMB_15__19_,
         u5_mult_87_SUMB_15__20_, u5_mult_87_SUMB_15__21_,
         u5_mult_87_SUMB_15__22_, u5_mult_87_SUMB_15__23_,
         u5_mult_87_SUMB_15__24_, u5_mult_87_SUMB_15__25_,
         u5_mult_87_SUMB_15__26_, u5_mult_87_SUMB_15__27_,
         u5_mult_87_SUMB_15__28_, u5_mult_87_SUMB_15__29_,
         u5_mult_87_SUMB_15__30_, u5_mult_87_SUMB_15__31_,
         u5_mult_87_SUMB_15__32_, u5_mult_87_SUMB_15__33_,
         u5_mult_87_SUMB_15__34_, u5_mult_87_SUMB_15__35_,
         u5_mult_87_SUMB_15__36_, u5_mult_87_SUMB_15__37_,
         u5_mult_87_SUMB_15__38_, u5_mult_87_SUMB_15__39_,
         u5_mult_87_SUMB_15__40_, u5_mult_87_SUMB_15__41_,
         u5_mult_87_SUMB_15__42_, u5_mult_87_SUMB_15__43_,
         u5_mult_87_SUMB_15__44_, u5_mult_87_SUMB_15__45_,
         u5_mult_87_SUMB_15__46_, u5_mult_87_SUMB_15__47_,
         u5_mult_87_SUMB_15__48_, u5_mult_87_SUMB_15__49_,
         u5_mult_87_SUMB_15__50_, u5_mult_87_SUMB_15__51_,
         u5_mult_87_SUMB_16__1_, u5_mult_87_SUMB_16__2_,
         u5_mult_87_SUMB_16__3_, u5_mult_87_SUMB_16__4_,
         u5_mult_87_SUMB_16__5_, u5_mult_87_SUMB_16__6_,
         u5_mult_87_SUMB_16__7_, u5_mult_87_SUMB_16__8_,
         u5_mult_87_SUMB_16__9_, u5_mult_87_SUMB_16__10_,
         u5_mult_87_SUMB_16__11_, u5_mult_87_SUMB_16__12_,
         u5_mult_87_SUMB_16__13_, u5_mult_87_SUMB_16__14_,
         u5_mult_87_SUMB_16__15_, u5_mult_87_SUMB_16__16_,
         u5_mult_87_SUMB_16__17_, u5_mult_87_SUMB_16__18_,
         u5_mult_87_SUMB_16__19_, u5_mult_87_SUMB_16__20_,
         u5_mult_87_SUMB_16__21_, u5_mult_87_SUMB_16__22_,
         u5_mult_87_SUMB_16__23_, u5_mult_87_SUMB_16__24_,
         u5_mult_87_SUMB_16__25_, u5_mult_87_SUMB_16__26_,
         u5_mult_87_SUMB_16__27_, u5_mult_87_SUMB_16__28_,
         u5_mult_87_SUMB_16__29_, u5_mult_87_SUMB_16__30_,
         u5_mult_87_SUMB_16__31_, u5_mult_87_SUMB_16__32_,
         u5_mult_87_SUMB_16__33_, u5_mult_87_SUMB_16__34_,
         u5_mult_87_SUMB_16__35_, u5_mult_87_SUMB_16__36_,
         u5_mult_87_SUMB_16__37_, u5_mult_87_SUMB_16__38_,
         u5_mult_87_SUMB_16__39_, u5_mult_87_SUMB_16__40_,
         u5_mult_87_SUMB_16__41_, u5_mult_87_SUMB_16__42_,
         u5_mult_87_SUMB_16__43_, u5_mult_87_SUMB_16__44_,
         u5_mult_87_SUMB_16__45_, u5_mult_87_SUMB_16__46_,
         u5_mult_87_SUMB_16__47_, u5_mult_87_SUMB_16__48_,
         u5_mult_87_SUMB_16__49_, u5_mult_87_SUMB_16__50_,
         u5_mult_87_SUMB_16__51_, u5_mult_87_SUMB_17__1_,
         u5_mult_87_SUMB_17__2_, u5_mult_87_SUMB_17__3_,
         u5_mult_87_SUMB_17__4_, u5_mult_87_SUMB_17__5_,
         u5_mult_87_SUMB_17__6_, u5_mult_87_SUMB_17__7_,
         u5_mult_87_SUMB_17__8_, u5_mult_87_SUMB_17__9_,
         u5_mult_87_SUMB_17__10_, u5_mult_87_SUMB_17__11_,
         u5_mult_87_SUMB_17__12_, u5_mult_87_SUMB_17__13_,
         u5_mult_87_SUMB_17__14_, u5_mult_87_SUMB_17__15_,
         u5_mult_87_SUMB_17__16_, u5_mult_87_SUMB_17__17_,
         u5_mult_87_SUMB_17__18_, u5_mult_87_SUMB_17__19_,
         u5_mult_87_SUMB_17__20_, u5_mult_87_SUMB_17__21_,
         u5_mult_87_SUMB_17__22_, u5_mult_87_SUMB_17__23_,
         u5_mult_87_SUMB_17__24_, u5_mult_87_SUMB_17__25_,
         u5_mult_87_SUMB_17__26_, u5_mult_87_SUMB_17__27_,
         u5_mult_87_SUMB_17__28_, u5_mult_87_SUMB_17__29_,
         u5_mult_87_SUMB_17__30_, u5_mult_87_SUMB_17__31_,
         u5_mult_87_SUMB_17__32_, u5_mult_87_SUMB_17__33_,
         u5_mult_87_SUMB_17__34_, u5_mult_87_SUMB_17__35_,
         u5_mult_87_SUMB_17__36_, u5_mult_87_SUMB_17__37_,
         u5_mult_87_SUMB_17__38_, u5_mult_87_SUMB_17__39_,
         u5_mult_87_SUMB_17__40_, u5_mult_87_SUMB_17__41_,
         u5_mult_87_SUMB_17__42_, u5_mult_87_SUMB_17__43_,
         u5_mult_87_SUMB_17__44_, u5_mult_87_SUMB_17__45_,
         u5_mult_87_SUMB_17__46_, u5_mult_87_SUMB_17__47_,
         u5_mult_87_SUMB_17__48_, u5_mult_87_SUMB_17__49_,
         u5_mult_87_SUMB_17__50_, u5_mult_87_SUMB_17__51_,
         u5_mult_87_SUMB_18__1_, u5_mult_87_SUMB_18__2_,
         u5_mult_87_SUMB_18__3_, u5_mult_87_SUMB_18__4_,
         u5_mult_87_SUMB_18__5_, u5_mult_87_SUMB_18__6_,
         u5_mult_87_SUMB_18__7_, u5_mult_87_SUMB_18__8_,
         u5_mult_87_SUMB_18__9_, u5_mult_87_SUMB_18__10_,
         u5_mult_87_SUMB_18__11_, u5_mult_87_SUMB_18__12_,
         u5_mult_87_SUMB_18__13_, u5_mult_87_SUMB_18__14_,
         u5_mult_87_SUMB_18__15_, u5_mult_87_SUMB_18__16_,
         u5_mult_87_SUMB_18__17_, u5_mult_87_SUMB_18__18_,
         u5_mult_87_SUMB_18__19_, u5_mult_87_SUMB_18__20_,
         u5_mult_87_SUMB_18__21_, u5_mult_87_SUMB_18__22_,
         u5_mult_87_SUMB_18__23_, u5_mult_87_SUMB_18__24_,
         u5_mult_87_SUMB_18__25_, u5_mult_87_SUMB_18__26_,
         u5_mult_87_SUMB_18__27_, u5_mult_87_SUMB_18__28_,
         u5_mult_87_SUMB_18__29_, u5_mult_87_SUMB_18__30_,
         u5_mult_87_SUMB_18__31_, u5_mult_87_SUMB_18__32_,
         u5_mult_87_SUMB_18__33_, u5_mult_87_SUMB_18__34_,
         u5_mult_87_SUMB_18__35_, u5_mult_87_SUMB_18__36_,
         u5_mult_87_SUMB_18__37_, u5_mult_87_SUMB_18__38_,
         u5_mult_87_SUMB_18__39_, u5_mult_87_SUMB_18__40_,
         u5_mult_87_SUMB_18__41_, u5_mult_87_SUMB_18__42_,
         u5_mult_87_SUMB_18__43_, u5_mult_87_SUMB_18__44_,
         u5_mult_87_SUMB_18__45_, u5_mult_87_SUMB_18__46_,
         u5_mult_87_SUMB_18__47_, u5_mult_87_SUMB_18__48_,
         u5_mult_87_SUMB_18__49_, u5_mult_87_SUMB_18__50_,
         u5_mult_87_SUMB_18__51_, u5_mult_87_SUMB_19__1_,
         u5_mult_87_SUMB_19__2_, u5_mult_87_SUMB_19__3_,
         u5_mult_87_SUMB_19__4_, u5_mult_87_SUMB_19__5_,
         u5_mult_87_SUMB_19__6_, u5_mult_87_SUMB_19__7_,
         u5_mult_87_SUMB_19__8_, u5_mult_87_SUMB_19__9_,
         u5_mult_87_SUMB_19__10_, u5_mult_87_SUMB_19__11_,
         u5_mult_87_SUMB_19__12_, u5_mult_87_SUMB_19__13_,
         u5_mult_87_SUMB_19__14_, u5_mult_87_SUMB_19__15_,
         u5_mult_87_SUMB_19__16_, u5_mult_87_SUMB_19__17_,
         u5_mult_87_SUMB_19__18_, u5_mult_87_SUMB_19__19_,
         u5_mult_87_SUMB_19__20_, u5_mult_87_SUMB_19__21_,
         u5_mult_87_SUMB_19__22_, u5_mult_87_SUMB_19__23_,
         u5_mult_87_SUMB_19__24_, u5_mult_87_SUMB_19__25_,
         u5_mult_87_SUMB_19__26_, u5_mult_87_SUMB_19__27_,
         u5_mult_87_SUMB_19__28_, u5_mult_87_SUMB_19__29_,
         u5_mult_87_SUMB_19__30_, u5_mult_87_SUMB_19__31_,
         u5_mult_87_SUMB_19__32_, u5_mult_87_SUMB_19__33_,
         u5_mult_87_SUMB_19__34_, u5_mult_87_SUMB_19__35_,
         u5_mult_87_SUMB_19__36_, u5_mult_87_SUMB_19__37_,
         u5_mult_87_SUMB_19__38_, u5_mult_87_SUMB_19__39_,
         u5_mult_87_SUMB_19__40_, u5_mult_87_SUMB_19__41_,
         u5_mult_87_SUMB_19__42_, u5_mult_87_SUMB_19__43_,
         u5_mult_87_SUMB_19__44_, u5_mult_87_SUMB_19__45_,
         u5_mult_87_SUMB_19__46_, u5_mult_87_SUMB_19__47_,
         u5_mult_87_SUMB_19__48_, u5_mult_87_SUMB_19__49_,
         u5_mult_87_SUMB_19__50_, u5_mult_87_SUMB_19__51_,
         u5_mult_87_SUMB_20__1_, u5_mult_87_SUMB_20__2_,
         u5_mult_87_SUMB_20__3_, u5_mult_87_SUMB_20__4_,
         u5_mult_87_SUMB_20__5_, u5_mult_87_SUMB_20__6_,
         u5_mult_87_SUMB_20__7_, u5_mult_87_SUMB_20__8_,
         u5_mult_87_SUMB_20__9_, u5_mult_87_SUMB_20__10_,
         u5_mult_87_SUMB_20__11_, u5_mult_87_SUMB_20__12_,
         u5_mult_87_SUMB_20__13_, u5_mult_87_SUMB_20__14_,
         u5_mult_87_SUMB_20__15_, u5_mult_87_SUMB_20__16_,
         u5_mult_87_SUMB_20__17_, u5_mult_87_SUMB_20__18_,
         u5_mult_87_SUMB_20__19_, u5_mult_87_SUMB_20__20_,
         u5_mult_87_SUMB_20__21_, u5_mult_87_SUMB_20__22_,
         u5_mult_87_SUMB_20__23_, u5_mult_87_SUMB_20__24_,
         u5_mult_87_SUMB_20__25_, u5_mult_87_SUMB_20__26_,
         u5_mult_87_SUMB_20__27_, u5_mult_87_SUMB_20__28_,
         u5_mult_87_SUMB_20__29_, u5_mult_87_SUMB_20__30_,
         u5_mult_87_SUMB_20__31_, u5_mult_87_SUMB_20__32_,
         u5_mult_87_SUMB_20__33_, u5_mult_87_SUMB_20__34_,
         u5_mult_87_SUMB_20__35_, u5_mult_87_SUMB_20__36_,
         u5_mult_87_SUMB_20__37_, u5_mult_87_SUMB_20__38_,
         u5_mult_87_SUMB_20__39_, u5_mult_87_SUMB_20__40_,
         u5_mult_87_SUMB_20__41_, u5_mult_87_SUMB_20__42_,
         u5_mult_87_SUMB_20__43_, u5_mult_87_SUMB_20__44_,
         u5_mult_87_SUMB_20__45_, u5_mult_87_SUMB_20__46_,
         u5_mult_87_SUMB_20__47_, u5_mult_87_SUMB_20__48_,
         u5_mult_87_SUMB_20__49_, u5_mult_87_SUMB_20__50_,
         u5_mult_87_SUMB_20__51_, u5_mult_87_SUMB_21__1_,
         u5_mult_87_SUMB_21__2_, u5_mult_87_SUMB_21__3_,
         u5_mult_87_SUMB_21__4_, u5_mult_87_SUMB_21__5_,
         u5_mult_87_SUMB_21__6_, u5_mult_87_SUMB_21__7_,
         u5_mult_87_SUMB_21__8_, u5_mult_87_SUMB_21__9_,
         u5_mult_87_SUMB_21__10_, u5_mult_87_SUMB_21__11_,
         u5_mult_87_SUMB_21__12_, u5_mult_87_SUMB_21__13_,
         u5_mult_87_SUMB_21__14_, u5_mult_87_SUMB_21__15_,
         u5_mult_87_SUMB_21__16_, u5_mult_87_SUMB_21__17_,
         u5_mult_87_SUMB_21__18_, u5_mult_87_SUMB_21__19_,
         u5_mult_87_SUMB_21__20_, u5_mult_87_SUMB_21__21_,
         u5_mult_87_SUMB_21__22_, u5_mult_87_SUMB_21__23_,
         u5_mult_87_SUMB_21__24_, u5_mult_87_SUMB_21__25_,
         u5_mult_87_SUMB_21__26_, u5_mult_87_SUMB_21__27_,
         u5_mult_87_SUMB_21__28_, u5_mult_87_SUMB_21__29_,
         u5_mult_87_SUMB_21__30_, u5_mult_87_SUMB_21__31_,
         u5_mult_87_SUMB_21__32_, u5_mult_87_SUMB_21__33_,
         u5_mult_87_SUMB_21__34_, u5_mult_87_SUMB_21__35_,
         u5_mult_87_SUMB_21__36_, u5_mult_87_SUMB_21__37_,
         u5_mult_87_SUMB_21__38_, u5_mult_87_SUMB_21__39_,
         u5_mult_87_SUMB_21__40_, u5_mult_87_SUMB_21__41_,
         u5_mult_87_SUMB_21__42_, u5_mult_87_SUMB_21__43_,
         u5_mult_87_SUMB_21__44_, u5_mult_87_SUMB_21__45_,
         u5_mult_87_SUMB_21__46_, u5_mult_87_SUMB_21__47_,
         u5_mult_87_SUMB_21__48_, u5_mult_87_SUMB_21__49_,
         u5_mult_87_SUMB_21__50_, u5_mult_87_SUMB_21__51_,
         u5_mult_87_SUMB_22__1_, u5_mult_87_SUMB_22__2_,
         u5_mult_87_SUMB_22__3_, u5_mult_87_SUMB_22__4_,
         u5_mult_87_SUMB_22__5_, u5_mult_87_SUMB_22__6_,
         u5_mult_87_SUMB_22__7_, u5_mult_87_SUMB_22__8_,
         u5_mult_87_SUMB_22__9_, u5_mult_87_SUMB_22__10_,
         u5_mult_87_SUMB_22__11_, u5_mult_87_SUMB_22__12_,
         u5_mult_87_SUMB_22__13_, u5_mult_87_SUMB_22__14_,
         u5_mult_87_SUMB_22__15_, u5_mult_87_SUMB_22__16_,
         u5_mult_87_SUMB_22__17_, u5_mult_87_SUMB_22__18_,
         u5_mult_87_SUMB_22__19_, u5_mult_87_SUMB_22__20_,
         u5_mult_87_SUMB_22__21_, u5_mult_87_SUMB_22__22_,
         u5_mult_87_SUMB_22__23_, u5_mult_87_SUMB_22__24_,
         u5_mult_87_SUMB_22__25_, u5_mult_87_SUMB_22__26_,
         u5_mult_87_SUMB_22__27_, u5_mult_87_SUMB_22__28_,
         u5_mult_87_SUMB_22__29_, u5_mult_87_SUMB_22__30_,
         u5_mult_87_SUMB_22__31_, u5_mult_87_SUMB_22__32_,
         u5_mult_87_SUMB_22__33_, u5_mult_87_SUMB_22__34_,
         u5_mult_87_SUMB_22__35_, u5_mult_87_SUMB_22__36_,
         u5_mult_87_SUMB_22__37_, u5_mult_87_SUMB_22__38_,
         u5_mult_87_SUMB_22__39_, u5_mult_87_SUMB_22__40_,
         u5_mult_87_SUMB_22__41_, u5_mult_87_SUMB_22__42_,
         u5_mult_87_SUMB_22__43_, u5_mult_87_SUMB_22__44_,
         u5_mult_87_SUMB_22__45_, u5_mult_87_SUMB_22__46_,
         u5_mult_87_SUMB_22__47_, u5_mult_87_SUMB_22__48_,
         u5_mult_87_SUMB_22__49_, u5_mult_87_SUMB_22__50_,
         u5_mult_87_SUMB_22__51_, u5_mult_87_SUMB_23__1_,
         u5_mult_87_SUMB_23__2_, u5_mult_87_SUMB_23__3_,
         u5_mult_87_SUMB_23__4_, u5_mult_87_SUMB_23__5_,
         u5_mult_87_SUMB_23__6_, u5_mult_87_SUMB_23__7_,
         u5_mult_87_SUMB_23__8_, u5_mult_87_SUMB_23__9_,
         u5_mult_87_SUMB_23__10_, u5_mult_87_SUMB_23__11_,
         u5_mult_87_SUMB_23__12_, u5_mult_87_SUMB_23__13_,
         u5_mult_87_SUMB_23__14_, u5_mult_87_SUMB_23__15_,
         u5_mult_87_SUMB_23__16_, u5_mult_87_SUMB_23__17_,
         u5_mult_87_SUMB_23__18_, u5_mult_87_SUMB_23__19_,
         u5_mult_87_SUMB_23__20_, u5_mult_87_SUMB_23__21_,
         u5_mult_87_SUMB_23__22_, u5_mult_87_SUMB_23__23_,
         u5_mult_87_SUMB_23__24_, u5_mult_87_SUMB_23__25_,
         u5_mult_87_SUMB_23__26_, u5_mult_87_SUMB_23__27_,
         u5_mult_87_SUMB_23__28_, u5_mult_87_SUMB_23__29_,
         u5_mult_87_SUMB_23__30_, u5_mult_87_SUMB_23__31_,
         u5_mult_87_SUMB_23__32_, u5_mult_87_SUMB_23__33_,
         u5_mult_87_SUMB_23__34_, u5_mult_87_SUMB_23__35_,
         u5_mult_87_SUMB_23__36_, u5_mult_87_SUMB_23__37_,
         u5_mult_87_SUMB_23__38_, u5_mult_87_SUMB_23__39_,
         u5_mult_87_SUMB_23__40_, u5_mult_87_SUMB_23__41_,
         u5_mult_87_SUMB_23__42_, u5_mult_87_SUMB_23__43_,
         u5_mult_87_SUMB_23__44_, u5_mult_87_SUMB_23__45_,
         u5_mult_87_SUMB_23__46_, u5_mult_87_SUMB_23__47_,
         u5_mult_87_SUMB_23__48_, u5_mult_87_SUMB_23__49_,
         u5_mult_87_SUMB_23__50_, u5_mult_87_SUMB_23__51_,
         u5_mult_87_CARRYB_14__19_, u5_mult_87_CARRYB_14__20_,
         u5_mult_87_CARRYB_14__21_, u5_mult_87_CARRYB_14__22_,
         u5_mult_87_CARRYB_14__23_, u5_mult_87_CARRYB_14__24_,
         u5_mult_87_CARRYB_14__25_, u5_mult_87_CARRYB_14__26_,
         u5_mult_87_CARRYB_14__27_, u5_mult_87_CARRYB_14__28_,
         u5_mult_87_CARRYB_14__29_, u5_mult_87_CARRYB_14__30_,
         u5_mult_87_CARRYB_14__31_, u5_mult_87_CARRYB_14__32_,
         u5_mult_87_CARRYB_14__33_, u5_mult_87_CARRYB_14__34_,
         u5_mult_87_CARRYB_14__35_, u5_mult_87_CARRYB_14__36_,
         u5_mult_87_CARRYB_14__37_, u5_mult_87_CARRYB_14__38_,
         u5_mult_87_CARRYB_14__39_, u5_mult_87_CARRYB_14__40_,
         u5_mult_87_CARRYB_14__41_, u5_mult_87_CARRYB_14__42_,
         u5_mult_87_CARRYB_14__43_, u5_mult_87_CARRYB_14__44_,
         u5_mult_87_CARRYB_14__45_, u5_mult_87_CARRYB_14__46_,
         u5_mult_87_CARRYB_14__47_, u5_mult_87_CARRYB_14__48_,
         u5_mult_87_CARRYB_14__49_, u5_mult_87_CARRYB_14__50_,
         u5_mult_87_CARRYB_14__51_, u5_mult_87_CARRYB_15__0_,
         u5_mult_87_CARRYB_15__1_, u5_mult_87_CARRYB_15__2_,
         u5_mult_87_CARRYB_15__3_, u5_mult_87_CARRYB_15__4_,
         u5_mult_87_CARRYB_15__5_, u5_mult_87_CARRYB_15__6_,
         u5_mult_87_CARRYB_15__7_, u5_mult_87_CARRYB_15__8_,
         u5_mult_87_CARRYB_15__9_, u5_mult_87_CARRYB_15__10_,
         u5_mult_87_CARRYB_15__11_, u5_mult_87_CARRYB_15__12_,
         u5_mult_87_CARRYB_15__13_, u5_mult_87_CARRYB_15__14_,
         u5_mult_87_CARRYB_15__15_, u5_mult_87_CARRYB_15__16_,
         u5_mult_87_CARRYB_15__17_, u5_mult_87_CARRYB_15__18_,
         u5_mult_87_CARRYB_15__19_, u5_mult_87_CARRYB_15__20_,
         u5_mult_87_CARRYB_15__21_, u5_mult_87_CARRYB_15__22_,
         u5_mult_87_CARRYB_15__23_, u5_mult_87_CARRYB_15__24_,
         u5_mult_87_CARRYB_15__25_, u5_mult_87_CARRYB_15__26_,
         u5_mult_87_CARRYB_15__27_, u5_mult_87_CARRYB_15__28_,
         u5_mult_87_CARRYB_15__29_, u5_mult_87_CARRYB_15__30_,
         u5_mult_87_CARRYB_15__31_, u5_mult_87_CARRYB_15__32_,
         u5_mult_87_CARRYB_15__33_, u5_mult_87_CARRYB_15__34_,
         u5_mult_87_CARRYB_15__35_, u5_mult_87_CARRYB_15__36_,
         u5_mult_87_CARRYB_15__37_, u5_mult_87_CARRYB_15__38_,
         u5_mult_87_CARRYB_15__39_, u5_mult_87_CARRYB_15__40_,
         u5_mult_87_CARRYB_15__41_, u5_mult_87_CARRYB_15__42_,
         u5_mult_87_CARRYB_15__43_, u5_mult_87_CARRYB_15__44_,
         u5_mult_87_CARRYB_15__45_, u5_mult_87_CARRYB_15__46_,
         u5_mult_87_CARRYB_15__47_, u5_mult_87_CARRYB_15__48_,
         u5_mult_87_CARRYB_15__49_, u5_mult_87_CARRYB_15__50_,
         u5_mult_87_CARRYB_15__51_, u5_mult_87_CARRYB_16__0_,
         u5_mult_87_CARRYB_16__1_, u5_mult_87_CARRYB_16__2_,
         u5_mult_87_CARRYB_16__3_, u5_mult_87_CARRYB_16__4_,
         u5_mult_87_CARRYB_16__5_, u5_mult_87_CARRYB_16__6_,
         u5_mult_87_CARRYB_16__7_, u5_mult_87_CARRYB_16__8_,
         u5_mult_87_CARRYB_16__9_, u5_mult_87_CARRYB_16__10_,
         u5_mult_87_CARRYB_16__11_, u5_mult_87_CARRYB_16__12_,
         u5_mult_87_CARRYB_16__13_, u5_mult_87_CARRYB_16__14_,
         u5_mult_87_CARRYB_16__15_, u5_mult_87_CARRYB_16__16_,
         u5_mult_87_CARRYB_16__17_, u5_mult_87_CARRYB_16__18_,
         u5_mult_87_CARRYB_16__19_, u5_mult_87_CARRYB_16__20_,
         u5_mult_87_CARRYB_16__21_, u5_mult_87_CARRYB_16__22_,
         u5_mult_87_CARRYB_16__23_, u5_mult_87_CARRYB_16__24_,
         u5_mult_87_CARRYB_16__25_, u5_mult_87_CARRYB_16__26_,
         u5_mult_87_CARRYB_16__27_, u5_mult_87_CARRYB_16__28_,
         u5_mult_87_CARRYB_16__29_, u5_mult_87_CARRYB_16__30_,
         u5_mult_87_CARRYB_16__31_, u5_mult_87_CARRYB_16__32_,
         u5_mult_87_CARRYB_16__33_, u5_mult_87_CARRYB_16__34_,
         u5_mult_87_CARRYB_16__35_, u5_mult_87_CARRYB_16__36_,
         u5_mult_87_CARRYB_16__37_, u5_mult_87_CARRYB_16__38_,
         u5_mult_87_CARRYB_16__39_, u5_mult_87_CARRYB_16__40_,
         u5_mult_87_CARRYB_16__41_, u5_mult_87_CARRYB_16__42_,
         u5_mult_87_CARRYB_16__43_, u5_mult_87_CARRYB_16__44_,
         u5_mult_87_CARRYB_16__45_, u5_mult_87_CARRYB_16__46_,
         u5_mult_87_CARRYB_16__47_, u5_mult_87_CARRYB_16__48_,
         u5_mult_87_CARRYB_16__49_, u5_mult_87_CARRYB_16__50_,
         u5_mult_87_CARRYB_16__51_, u5_mult_87_CARRYB_17__0_,
         u5_mult_87_CARRYB_17__1_, u5_mult_87_CARRYB_17__2_,
         u5_mult_87_CARRYB_17__3_, u5_mult_87_CARRYB_17__4_,
         u5_mult_87_CARRYB_17__5_, u5_mult_87_CARRYB_17__6_,
         u5_mult_87_CARRYB_17__7_, u5_mult_87_CARRYB_17__8_,
         u5_mult_87_CARRYB_17__9_, u5_mult_87_CARRYB_17__10_,
         u5_mult_87_CARRYB_17__11_, u5_mult_87_CARRYB_17__12_,
         u5_mult_87_CARRYB_17__13_, u5_mult_87_CARRYB_17__14_,
         u5_mult_87_CARRYB_17__15_, u5_mult_87_CARRYB_17__16_,
         u5_mult_87_CARRYB_17__17_, u5_mult_87_CARRYB_17__18_,
         u5_mult_87_CARRYB_17__19_, u5_mult_87_CARRYB_17__20_,
         u5_mult_87_CARRYB_17__21_, u5_mult_87_CARRYB_17__22_,
         u5_mult_87_CARRYB_17__23_, u5_mult_87_CARRYB_17__24_,
         u5_mult_87_CARRYB_17__25_, u5_mult_87_CARRYB_17__26_,
         u5_mult_87_CARRYB_17__27_, u5_mult_87_CARRYB_17__28_,
         u5_mult_87_CARRYB_17__29_, u5_mult_87_CARRYB_17__30_,
         u5_mult_87_CARRYB_17__31_, u5_mult_87_CARRYB_17__32_,
         u5_mult_87_CARRYB_17__33_, u5_mult_87_CARRYB_17__34_,
         u5_mult_87_CARRYB_17__35_, u5_mult_87_CARRYB_17__36_,
         u5_mult_87_CARRYB_17__37_, u5_mult_87_CARRYB_17__38_,
         u5_mult_87_CARRYB_17__39_, u5_mult_87_CARRYB_17__40_,
         u5_mult_87_CARRYB_17__41_, u5_mult_87_CARRYB_17__42_,
         u5_mult_87_CARRYB_17__43_, u5_mult_87_CARRYB_17__44_,
         u5_mult_87_CARRYB_17__45_, u5_mult_87_CARRYB_17__46_,
         u5_mult_87_CARRYB_17__47_, u5_mult_87_CARRYB_17__48_,
         u5_mult_87_CARRYB_17__49_, u5_mult_87_CARRYB_17__50_,
         u5_mult_87_CARRYB_17__51_, u5_mult_87_CARRYB_18__0_,
         u5_mult_87_CARRYB_18__1_, u5_mult_87_CARRYB_18__2_,
         u5_mult_87_CARRYB_18__3_, u5_mult_87_CARRYB_18__4_,
         u5_mult_87_CARRYB_18__5_, u5_mult_87_CARRYB_18__6_,
         u5_mult_87_CARRYB_18__7_, u5_mult_87_CARRYB_18__8_,
         u5_mult_87_CARRYB_18__9_, u5_mult_87_CARRYB_18__10_,
         u5_mult_87_CARRYB_18__11_, u5_mult_87_CARRYB_18__12_,
         u5_mult_87_CARRYB_18__13_, u5_mult_87_CARRYB_18__14_,
         u5_mult_87_CARRYB_18__15_, u5_mult_87_CARRYB_18__16_,
         u5_mult_87_CARRYB_18__17_, u5_mult_87_CARRYB_18__18_,
         u5_mult_87_CARRYB_18__19_, u5_mult_87_CARRYB_18__20_,
         u5_mult_87_CARRYB_18__21_, u5_mult_87_CARRYB_18__22_,
         u5_mult_87_CARRYB_18__23_, u5_mult_87_CARRYB_18__24_,
         u5_mult_87_CARRYB_18__25_, u5_mult_87_CARRYB_18__26_,
         u5_mult_87_CARRYB_18__27_, u5_mult_87_CARRYB_18__28_,
         u5_mult_87_CARRYB_18__29_, u5_mult_87_CARRYB_18__30_,
         u5_mult_87_CARRYB_18__31_, u5_mult_87_CARRYB_18__32_,
         u5_mult_87_CARRYB_18__33_, u5_mult_87_CARRYB_18__34_,
         u5_mult_87_CARRYB_18__35_, u5_mult_87_CARRYB_18__36_,
         u5_mult_87_CARRYB_18__37_, u5_mult_87_CARRYB_18__38_,
         u5_mult_87_CARRYB_18__39_, u5_mult_87_CARRYB_18__40_,
         u5_mult_87_CARRYB_18__41_, u5_mult_87_CARRYB_18__42_,
         u5_mult_87_CARRYB_18__43_, u5_mult_87_CARRYB_18__44_,
         u5_mult_87_CARRYB_18__45_, u5_mult_87_CARRYB_18__46_,
         u5_mult_87_CARRYB_18__47_, u5_mult_87_CARRYB_18__48_,
         u5_mult_87_CARRYB_18__49_, u5_mult_87_CARRYB_18__50_,
         u5_mult_87_CARRYB_18__51_, u5_mult_87_CARRYB_19__0_,
         u5_mult_87_CARRYB_19__1_, u5_mult_87_CARRYB_19__2_,
         u5_mult_87_CARRYB_19__3_, u5_mult_87_CARRYB_19__4_,
         u5_mult_87_CARRYB_19__5_, u5_mult_87_CARRYB_19__6_,
         u5_mult_87_CARRYB_19__7_, u5_mult_87_CARRYB_19__8_,
         u5_mult_87_CARRYB_19__9_, u5_mult_87_CARRYB_19__10_,
         u5_mult_87_CARRYB_19__11_, u5_mult_87_CARRYB_19__12_,
         u5_mult_87_CARRYB_19__13_, u5_mult_87_CARRYB_19__14_,
         u5_mult_87_CARRYB_19__15_, u5_mult_87_CARRYB_19__16_,
         u5_mult_87_CARRYB_19__17_, u5_mult_87_CARRYB_19__18_,
         u5_mult_87_CARRYB_19__19_, u5_mult_87_CARRYB_19__20_,
         u5_mult_87_CARRYB_19__21_, u5_mult_87_CARRYB_19__22_,
         u5_mult_87_CARRYB_19__23_, u5_mult_87_CARRYB_19__24_,
         u5_mult_87_CARRYB_19__25_, u5_mult_87_CARRYB_19__26_,
         u5_mult_87_CARRYB_19__27_, u5_mult_87_CARRYB_19__28_,
         u5_mult_87_CARRYB_19__29_, u5_mult_87_CARRYB_19__30_,
         u5_mult_87_CARRYB_19__31_, u5_mult_87_CARRYB_19__32_,
         u5_mult_87_CARRYB_19__33_, u5_mult_87_CARRYB_19__34_,
         u5_mult_87_CARRYB_19__35_, u5_mult_87_CARRYB_19__36_,
         u5_mult_87_CARRYB_19__37_, u5_mult_87_CARRYB_19__38_,
         u5_mult_87_CARRYB_19__39_, u5_mult_87_CARRYB_19__40_,
         u5_mult_87_CARRYB_19__41_, u5_mult_87_CARRYB_19__42_,
         u5_mult_87_CARRYB_19__43_, u5_mult_87_CARRYB_19__44_,
         u5_mult_87_CARRYB_19__45_, u5_mult_87_CARRYB_19__46_,
         u5_mult_87_CARRYB_19__47_, u5_mult_87_CARRYB_19__48_,
         u5_mult_87_CARRYB_19__49_, u5_mult_87_CARRYB_19__50_,
         u5_mult_87_CARRYB_19__51_, u5_mult_87_CARRYB_20__0_,
         u5_mult_87_CARRYB_20__1_, u5_mult_87_CARRYB_20__2_,
         u5_mult_87_CARRYB_20__3_, u5_mult_87_CARRYB_20__4_,
         u5_mult_87_CARRYB_20__5_, u5_mult_87_CARRYB_20__6_,
         u5_mult_87_CARRYB_20__7_, u5_mult_87_CARRYB_20__8_,
         u5_mult_87_CARRYB_20__9_, u5_mult_87_CARRYB_20__10_,
         u5_mult_87_CARRYB_20__11_, u5_mult_87_CARRYB_20__12_,
         u5_mult_87_CARRYB_20__13_, u5_mult_87_CARRYB_20__14_,
         u5_mult_87_CARRYB_20__15_, u5_mult_87_CARRYB_20__16_,
         u5_mult_87_CARRYB_20__17_, u5_mult_87_CARRYB_20__18_,
         u5_mult_87_CARRYB_20__19_, u5_mult_87_CARRYB_20__20_,
         u5_mult_87_CARRYB_20__21_, u5_mult_87_CARRYB_20__22_,
         u5_mult_87_CARRYB_20__23_, u5_mult_87_CARRYB_20__24_,
         u5_mult_87_CARRYB_20__25_, u5_mult_87_CARRYB_20__26_,
         u5_mult_87_CARRYB_20__27_, u5_mult_87_CARRYB_20__28_,
         u5_mult_87_CARRYB_20__29_, u5_mult_87_CARRYB_20__30_,
         u5_mult_87_CARRYB_20__31_, u5_mult_87_CARRYB_20__32_,
         u5_mult_87_CARRYB_20__33_, u5_mult_87_CARRYB_20__34_,
         u5_mult_87_CARRYB_20__35_, u5_mult_87_CARRYB_20__36_,
         u5_mult_87_CARRYB_20__37_, u5_mult_87_CARRYB_20__38_,
         u5_mult_87_CARRYB_20__39_, u5_mult_87_CARRYB_20__40_,
         u5_mult_87_CARRYB_20__41_, u5_mult_87_CARRYB_20__42_,
         u5_mult_87_CARRYB_20__43_, u5_mult_87_CARRYB_20__44_,
         u5_mult_87_CARRYB_20__45_, u5_mult_87_CARRYB_20__46_,
         u5_mult_87_CARRYB_20__47_, u5_mult_87_CARRYB_20__48_,
         u5_mult_87_CARRYB_20__49_, u5_mult_87_CARRYB_20__50_,
         u5_mult_87_CARRYB_20__51_, u5_mult_87_CARRYB_21__0_,
         u5_mult_87_CARRYB_21__1_, u5_mult_87_CARRYB_21__2_,
         u5_mult_87_CARRYB_21__3_, u5_mult_87_CARRYB_21__4_,
         u5_mult_87_CARRYB_21__5_, u5_mult_87_CARRYB_21__6_,
         u5_mult_87_CARRYB_21__7_, u5_mult_87_CARRYB_21__8_,
         u5_mult_87_CARRYB_21__9_, u5_mult_87_CARRYB_21__10_,
         u5_mult_87_CARRYB_21__11_, u5_mult_87_CARRYB_21__12_,
         u5_mult_87_CARRYB_21__13_, u5_mult_87_CARRYB_21__14_,
         u5_mult_87_CARRYB_21__15_, u5_mult_87_CARRYB_21__16_,
         u5_mult_87_CARRYB_21__17_, u5_mult_87_CARRYB_21__18_,
         u5_mult_87_CARRYB_21__19_, u5_mult_87_CARRYB_21__20_,
         u5_mult_87_CARRYB_21__21_, u5_mult_87_CARRYB_21__22_,
         u5_mult_87_CARRYB_21__23_, u5_mult_87_CARRYB_21__24_,
         u5_mult_87_CARRYB_21__25_, u5_mult_87_CARRYB_21__26_,
         u5_mult_87_CARRYB_21__27_, u5_mult_87_CARRYB_21__28_,
         u5_mult_87_CARRYB_21__29_, u5_mult_87_CARRYB_21__30_,
         u5_mult_87_CARRYB_21__31_, u5_mult_87_CARRYB_21__32_,
         u5_mult_87_CARRYB_21__33_, u5_mult_87_CARRYB_21__34_,
         u5_mult_87_CARRYB_21__35_, u5_mult_87_CARRYB_21__36_,
         u5_mult_87_CARRYB_21__37_, u5_mult_87_CARRYB_21__38_,
         u5_mult_87_CARRYB_21__39_, u5_mult_87_CARRYB_21__40_,
         u5_mult_87_CARRYB_21__41_, u5_mult_87_CARRYB_21__42_,
         u5_mult_87_CARRYB_21__43_, u5_mult_87_CARRYB_21__44_,
         u5_mult_87_CARRYB_21__45_, u5_mult_87_CARRYB_21__46_,
         u5_mult_87_CARRYB_21__47_, u5_mult_87_CARRYB_21__48_,
         u5_mult_87_CARRYB_21__49_, u5_mult_87_CARRYB_21__50_,
         u5_mult_87_CARRYB_21__51_, u5_mult_87_CARRYB_22__0_,
         u5_mult_87_CARRYB_22__1_, u5_mult_87_CARRYB_22__2_,
         u5_mult_87_CARRYB_22__3_, u5_mult_87_CARRYB_22__4_,
         u5_mult_87_CARRYB_22__5_, u5_mult_87_CARRYB_22__6_,
         u5_mult_87_CARRYB_22__7_, u5_mult_87_CARRYB_22__8_,
         u5_mult_87_CARRYB_22__9_, u5_mult_87_CARRYB_22__10_,
         u5_mult_87_CARRYB_22__11_, u5_mult_87_CARRYB_22__12_,
         u5_mult_87_CARRYB_22__13_, u5_mult_87_CARRYB_22__14_,
         u5_mult_87_CARRYB_22__15_, u5_mult_87_CARRYB_22__16_,
         u5_mult_87_CARRYB_22__17_, u5_mult_87_CARRYB_22__18_,
         u5_mult_87_CARRYB_22__19_, u5_mult_87_CARRYB_22__20_,
         u5_mult_87_CARRYB_22__21_, u5_mult_87_CARRYB_22__22_,
         u5_mult_87_CARRYB_22__23_, u5_mult_87_CARRYB_22__24_,
         u5_mult_87_CARRYB_22__25_, u5_mult_87_CARRYB_22__26_,
         u5_mult_87_CARRYB_22__27_, u5_mult_87_CARRYB_22__28_,
         u5_mult_87_CARRYB_22__29_, u5_mult_87_CARRYB_22__30_,
         u5_mult_87_CARRYB_22__31_, u5_mult_87_CARRYB_22__32_,
         u5_mult_87_CARRYB_22__33_, u5_mult_87_CARRYB_22__34_,
         u5_mult_87_CARRYB_22__35_, u5_mult_87_CARRYB_22__36_,
         u5_mult_87_CARRYB_22__37_, u5_mult_87_CARRYB_22__38_,
         u5_mult_87_CARRYB_22__39_, u5_mult_87_CARRYB_22__40_,
         u5_mult_87_CARRYB_22__41_, u5_mult_87_CARRYB_22__42_,
         u5_mult_87_CARRYB_22__43_, u5_mult_87_CARRYB_22__44_,
         u5_mult_87_CARRYB_22__45_, u5_mult_87_CARRYB_22__46_,
         u5_mult_87_CARRYB_22__47_, u5_mult_87_CARRYB_22__48_,
         u5_mult_87_CARRYB_22__49_, u5_mult_87_CARRYB_22__50_,
         u5_mult_87_CARRYB_22__51_, u5_mult_87_CARRYB_23__0_,
         u5_mult_87_CARRYB_23__1_, u5_mult_87_CARRYB_23__2_,
         u5_mult_87_CARRYB_23__3_, u5_mult_87_CARRYB_23__4_,
         u5_mult_87_CARRYB_23__5_, u5_mult_87_CARRYB_23__6_,
         u5_mult_87_CARRYB_23__7_, u5_mult_87_CARRYB_23__8_,
         u5_mult_87_CARRYB_23__9_, u5_mult_87_CARRYB_23__10_,
         u5_mult_87_CARRYB_23__11_, u5_mult_87_CARRYB_23__12_,
         u5_mult_87_CARRYB_23__13_, u5_mult_87_CARRYB_23__14_,
         u5_mult_87_CARRYB_23__15_, u5_mult_87_CARRYB_23__16_,
         u5_mult_87_CARRYB_23__17_, u5_mult_87_CARRYB_23__18_,
         u5_mult_87_CARRYB_23__19_, u5_mult_87_CARRYB_23__20_,
         u5_mult_87_CARRYB_23__21_, u5_mult_87_CARRYB_23__22_,
         u5_mult_87_CARRYB_23__23_, u5_mult_87_CARRYB_23__24_,
         u5_mult_87_CARRYB_23__25_, u5_mult_87_CARRYB_23__26_,
         u5_mult_87_CARRYB_23__27_, u5_mult_87_CARRYB_23__28_,
         u5_mult_87_CARRYB_23__29_, u5_mult_87_CARRYB_23__30_,
         u5_mult_87_CARRYB_23__31_, u5_mult_87_CARRYB_23__32_,
         u5_mult_87_CARRYB_23__33_, u5_mult_87_CARRYB_23__34_,
         u5_mult_87_CARRYB_23__35_, u5_mult_87_CARRYB_23__36_,
         u5_mult_87_CARRYB_23__37_, u5_mult_87_CARRYB_23__38_,
         u5_mult_87_CARRYB_23__39_, u5_mult_87_CARRYB_23__40_,
         u5_mult_87_CARRYB_23__41_, u5_mult_87_CARRYB_23__42_,
         u5_mult_87_CARRYB_23__43_, u5_mult_87_CARRYB_23__44_,
         u5_mult_87_CARRYB_23__45_, u5_mult_87_CARRYB_23__46_,
         u5_mult_87_CARRYB_23__47_, u5_mult_87_CARRYB_23__48_,
         u5_mult_87_CARRYB_23__49_, u5_mult_87_CARRYB_23__50_,
         u5_mult_87_CARRYB_23__51_, u5_mult_87_CARRYB_24__0_,
         u5_mult_87_SUMB_4__37_, u5_mult_87_SUMB_4__38_,
         u5_mult_87_SUMB_4__39_, u5_mult_87_SUMB_4__40_,
         u5_mult_87_SUMB_4__41_, u5_mult_87_SUMB_4__42_,
         u5_mult_87_SUMB_4__43_, u5_mult_87_SUMB_4__44_,
         u5_mult_87_SUMB_4__45_, u5_mult_87_SUMB_4__46_,
         u5_mult_87_SUMB_4__47_, u5_mult_87_SUMB_4__48_,
         u5_mult_87_SUMB_4__49_, u5_mult_87_SUMB_4__50_,
         u5_mult_87_SUMB_4__51_, u5_mult_87_SUMB_5__1_, u5_mult_87_SUMB_5__2_,
         u5_mult_87_SUMB_5__3_, u5_mult_87_SUMB_5__4_, u5_mult_87_SUMB_5__5_,
         u5_mult_87_SUMB_5__6_, u5_mult_87_SUMB_5__7_, u5_mult_87_SUMB_5__8_,
         u5_mult_87_SUMB_5__9_, u5_mult_87_SUMB_5__10_, u5_mult_87_SUMB_5__11_,
         u5_mult_87_SUMB_5__12_, u5_mult_87_SUMB_5__13_,
         u5_mult_87_SUMB_5__14_, u5_mult_87_SUMB_5__15_,
         u5_mult_87_SUMB_5__16_, u5_mult_87_SUMB_5__17_,
         u5_mult_87_SUMB_5__18_, u5_mult_87_SUMB_5__19_,
         u5_mult_87_SUMB_5__20_, u5_mult_87_SUMB_5__21_,
         u5_mult_87_SUMB_5__22_, u5_mult_87_SUMB_5__23_,
         u5_mult_87_SUMB_5__24_, u5_mult_87_SUMB_5__25_,
         u5_mult_87_SUMB_5__26_, u5_mult_87_SUMB_5__27_,
         u5_mult_87_SUMB_5__28_, u5_mult_87_SUMB_5__29_,
         u5_mult_87_SUMB_5__30_, u5_mult_87_SUMB_5__31_,
         u5_mult_87_SUMB_5__32_, u5_mult_87_SUMB_5__33_,
         u5_mult_87_SUMB_5__34_, u5_mult_87_SUMB_5__35_,
         u5_mult_87_SUMB_5__36_, u5_mult_87_SUMB_5__37_,
         u5_mult_87_SUMB_5__38_, u5_mult_87_SUMB_5__39_,
         u5_mult_87_SUMB_5__40_, u5_mult_87_SUMB_5__41_,
         u5_mult_87_SUMB_5__42_, u5_mult_87_SUMB_5__43_,
         u5_mult_87_SUMB_5__44_, u5_mult_87_SUMB_5__45_,
         u5_mult_87_SUMB_5__46_, u5_mult_87_SUMB_5__47_,
         u5_mult_87_SUMB_5__48_, u5_mult_87_SUMB_5__49_,
         u5_mult_87_SUMB_5__50_, u5_mult_87_SUMB_5__51_, u5_mult_87_SUMB_6__1_,
         u5_mult_87_SUMB_6__2_, u5_mult_87_SUMB_6__3_, u5_mult_87_SUMB_6__4_,
         u5_mult_87_SUMB_6__5_, u5_mult_87_SUMB_6__6_, u5_mult_87_SUMB_6__7_,
         u5_mult_87_SUMB_6__8_, u5_mult_87_SUMB_6__9_, u5_mult_87_SUMB_6__10_,
         u5_mult_87_SUMB_6__11_, u5_mult_87_SUMB_6__12_,
         u5_mult_87_SUMB_6__13_, u5_mult_87_SUMB_6__14_,
         u5_mult_87_SUMB_6__15_, u5_mult_87_SUMB_6__16_,
         u5_mult_87_SUMB_6__17_, u5_mult_87_SUMB_6__18_,
         u5_mult_87_SUMB_6__19_, u5_mult_87_SUMB_6__20_,
         u5_mult_87_SUMB_6__21_, u5_mult_87_SUMB_6__22_,
         u5_mult_87_SUMB_6__23_, u5_mult_87_SUMB_6__24_,
         u5_mult_87_SUMB_6__25_, u5_mult_87_SUMB_6__26_,
         u5_mult_87_SUMB_6__27_, u5_mult_87_SUMB_6__28_,
         u5_mult_87_SUMB_6__29_, u5_mult_87_SUMB_6__30_,
         u5_mult_87_SUMB_6__31_, u5_mult_87_SUMB_6__32_,
         u5_mult_87_SUMB_6__33_, u5_mult_87_SUMB_6__34_,
         u5_mult_87_SUMB_6__35_, u5_mult_87_SUMB_6__36_,
         u5_mult_87_SUMB_6__37_, u5_mult_87_SUMB_6__38_,
         u5_mult_87_SUMB_6__39_, u5_mult_87_SUMB_6__40_,
         u5_mult_87_SUMB_6__41_, u5_mult_87_SUMB_6__42_,
         u5_mult_87_SUMB_6__43_, u5_mult_87_SUMB_6__44_,
         u5_mult_87_SUMB_6__45_, u5_mult_87_SUMB_6__46_,
         u5_mult_87_SUMB_6__47_, u5_mult_87_SUMB_6__48_,
         u5_mult_87_SUMB_6__49_, u5_mult_87_SUMB_6__50_,
         u5_mult_87_SUMB_6__51_, u5_mult_87_SUMB_7__1_, u5_mult_87_SUMB_7__2_,
         u5_mult_87_SUMB_7__3_, u5_mult_87_SUMB_7__4_, u5_mult_87_SUMB_7__5_,
         u5_mult_87_SUMB_7__6_, u5_mult_87_SUMB_7__7_, u5_mult_87_SUMB_7__8_,
         u5_mult_87_SUMB_7__9_, u5_mult_87_SUMB_7__10_, u5_mult_87_SUMB_7__11_,
         u5_mult_87_SUMB_7__12_, u5_mult_87_SUMB_7__13_,
         u5_mult_87_SUMB_7__14_, u5_mult_87_SUMB_7__15_,
         u5_mult_87_SUMB_7__16_, u5_mult_87_SUMB_7__17_,
         u5_mult_87_SUMB_7__18_, u5_mult_87_SUMB_7__19_,
         u5_mult_87_SUMB_7__20_, u5_mult_87_SUMB_7__21_,
         u5_mult_87_SUMB_7__22_, u5_mult_87_SUMB_7__23_,
         u5_mult_87_SUMB_7__24_, u5_mult_87_SUMB_7__25_,
         u5_mult_87_SUMB_7__26_, u5_mult_87_SUMB_7__27_,
         u5_mult_87_SUMB_7__28_, u5_mult_87_SUMB_7__29_,
         u5_mult_87_SUMB_7__30_, u5_mult_87_SUMB_7__31_,
         u5_mult_87_SUMB_7__32_, u5_mult_87_SUMB_7__33_,
         u5_mult_87_SUMB_7__34_, u5_mult_87_SUMB_7__35_,
         u5_mult_87_SUMB_7__36_, u5_mult_87_SUMB_7__37_,
         u5_mult_87_SUMB_7__38_, u5_mult_87_SUMB_7__39_,
         u5_mult_87_SUMB_7__40_, u5_mult_87_SUMB_7__41_,
         u5_mult_87_SUMB_7__42_, u5_mult_87_SUMB_7__43_,
         u5_mult_87_SUMB_7__44_, u5_mult_87_SUMB_7__45_,
         u5_mult_87_SUMB_7__46_, u5_mult_87_SUMB_7__47_,
         u5_mult_87_SUMB_7__48_, u5_mult_87_SUMB_7__49_,
         u5_mult_87_SUMB_7__50_, u5_mult_87_SUMB_7__51_, u5_mult_87_SUMB_8__1_,
         u5_mult_87_SUMB_8__2_, u5_mult_87_SUMB_8__3_, u5_mult_87_SUMB_8__4_,
         u5_mult_87_SUMB_8__5_, u5_mult_87_SUMB_8__6_, u5_mult_87_SUMB_8__7_,
         u5_mult_87_SUMB_8__8_, u5_mult_87_SUMB_8__9_, u5_mult_87_SUMB_8__10_,
         u5_mult_87_SUMB_8__11_, u5_mult_87_SUMB_8__12_,
         u5_mult_87_SUMB_8__13_, u5_mult_87_SUMB_8__14_,
         u5_mult_87_SUMB_8__15_, u5_mult_87_SUMB_8__16_,
         u5_mult_87_SUMB_8__17_, u5_mult_87_SUMB_8__18_,
         u5_mult_87_SUMB_8__19_, u5_mult_87_SUMB_8__20_,
         u5_mult_87_SUMB_8__21_, u5_mult_87_SUMB_8__22_,
         u5_mult_87_SUMB_8__23_, u5_mult_87_SUMB_8__24_,
         u5_mult_87_SUMB_8__25_, u5_mult_87_SUMB_8__26_,
         u5_mult_87_SUMB_8__27_, u5_mult_87_SUMB_8__28_,
         u5_mult_87_SUMB_8__29_, u5_mult_87_SUMB_8__30_,
         u5_mult_87_SUMB_8__31_, u5_mult_87_SUMB_8__32_,
         u5_mult_87_SUMB_8__33_, u5_mult_87_SUMB_8__34_,
         u5_mult_87_SUMB_8__35_, u5_mult_87_SUMB_8__36_,
         u5_mult_87_SUMB_8__37_, u5_mult_87_SUMB_8__38_,
         u5_mult_87_SUMB_8__39_, u5_mult_87_SUMB_8__40_,
         u5_mult_87_SUMB_8__41_, u5_mult_87_SUMB_8__42_,
         u5_mult_87_SUMB_8__43_, u5_mult_87_SUMB_8__44_,
         u5_mult_87_SUMB_8__45_, u5_mult_87_SUMB_8__46_,
         u5_mult_87_SUMB_8__47_, u5_mult_87_SUMB_8__48_,
         u5_mult_87_SUMB_8__49_, u5_mult_87_SUMB_8__50_,
         u5_mult_87_SUMB_8__51_, u5_mult_87_SUMB_9__1_, u5_mult_87_SUMB_9__2_,
         u5_mult_87_SUMB_9__3_, u5_mult_87_SUMB_9__4_, u5_mult_87_SUMB_9__5_,
         u5_mult_87_SUMB_9__6_, u5_mult_87_SUMB_9__7_, u5_mult_87_SUMB_9__8_,
         u5_mult_87_SUMB_9__9_, u5_mult_87_SUMB_9__10_, u5_mult_87_SUMB_9__11_,
         u5_mult_87_SUMB_9__12_, u5_mult_87_SUMB_9__13_,
         u5_mult_87_SUMB_9__14_, u5_mult_87_SUMB_9__15_,
         u5_mult_87_SUMB_9__16_, u5_mult_87_SUMB_9__17_,
         u5_mult_87_SUMB_9__18_, u5_mult_87_SUMB_9__19_,
         u5_mult_87_SUMB_9__20_, u5_mult_87_SUMB_9__21_,
         u5_mult_87_SUMB_9__22_, u5_mult_87_SUMB_9__23_,
         u5_mult_87_SUMB_9__24_, u5_mult_87_SUMB_9__25_,
         u5_mult_87_SUMB_9__26_, u5_mult_87_SUMB_9__27_,
         u5_mult_87_SUMB_9__28_, u5_mult_87_SUMB_9__29_,
         u5_mult_87_SUMB_9__30_, u5_mult_87_SUMB_9__31_,
         u5_mult_87_SUMB_9__32_, u5_mult_87_SUMB_9__33_,
         u5_mult_87_SUMB_9__34_, u5_mult_87_SUMB_9__35_,
         u5_mult_87_SUMB_9__36_, u5_mult_87_SUMB_9__37_,
         u5_mult_87_SUMB_9__38_, u5_mult_87_SUMB_9__39_,
         u5_mult_87_SUMB_9__40_, u5_mult_87_SUMB_9__41_,
         u5_mult_87_SUMB_9__42_, u5_mult_87_SUMB_9__43_,
         u5_mult_87_SUMB_9__44_, u5_mult_87_SUMB_9__45_,
         u5_mult_87_SUMB_9__46_, u5_mult_87_SUMB_9__47_,
         u5_mult_87_SUMB_9__48_, u5_mult_87_SUMB_9__49_,
         u5_mult_87_SUMB_9__50_, u5_mult_87_SUMB_9__51_,
         u5_mult_87_SUMB_10__1_, u5_mult_87_SUMB_10__2_,
         u5_mult_87_SUMB_10__3_, u5_mult_87_SUMB_10__4_,
         u5_mult_87_SUMB_10__5_, u5_mult_87_SUMB_10__6_,
         u5_mult_87_SUMB_10__7_, u5_mult_87_SUMB_10__8_,
         u5_mult_87_SUMB_10__9_, u5_mult_87_SUMB_10__10_,
         u5_mult_87_SUMB_10__11_, u5_mult_87_SUMB_10__12_,
         u5_mult_87_SUMB_10__13_, u5_mult_87_SUMB_10__14_,
         u5_mult_87_SUMB_10__15_, u5_mult_87_SUMB_10__16_,
         u5_mult_87_SUMB_10__17_, u5_mult_87_SUMB_10__18_,
         u5_mult_87_SUMB_10__19_, u5_mult_87_SUMB_10__20_,
         u5_mult_87_SUMB_10__21_, u5_mult_87_SUMB_10__22_,
         u5_mult_87_SUMB_10__23_, u5_mult_87_SUMB_10__24_,
         u5_mult_87_SUMB_10__25_, u5_mult_87_SUMB_10__26_,
         u5_mult_87_SUMB_10__27_, u5_mult_87_SUMB_10__28_,
         u5_mult_87_SUMB_10__29_, u5_mult_87_SUMB_10__30_,
         u5_mult_87_SUMB_10__31_, u5_mult_87_SUMB_10__32_,
         u5_mult_87_SUMB_10__33_, u5_mult_87_SUMB_10__34_,
         u5_mult_87_SUMB_10__35_, u5_mult_87_SUMB_10__36_,
         u5_mult_87_SUMB_10__37_, u5_mult_87_SUMB_10__38_,
         u5_mult_87_SUMB_10__39_, u5_mult_87_SUMB_10__40_,
         u5_mult_87_SUMB_10__41_, u5_mult_87_SUMB_10__42_,
         u5_mult_87_SUMB_10__43_, u5_mult_87_SUMB_10__44_,
         u5_mult_87_SUMB_10__45_, u5_mult_87_SUMB_10__46_,
         u5_mult_87_SUMB_10__47_, u5_mult_87_SUMB_10__48_,
         u5_mult_87_SUMB_10__49_, u5_mult_87_SUMB_10__50_,
         u5_mult_87_SUMB_10__51_, u5_mult_87_SUMB_11__1_,
         u5_mult_87_SUMB_11__2_, u5_mult_87_SUMB_11__3_,
         u5_mult_87_SUMB_11__4_, u5_mult_87_SUMB_11__5_,
         u5_mult_87_SUMB_11__6_, u5_mult_87_SUMB_11__7_,
         u5_mult_87_SUMB_11__8_, u5_mult_87_SUMB_11__9_,
         u5_mult_87_SUMB_11__10_, u5_mult_87_SUMB_11__11_,
         u5_mult_87_SUMB_11__12_, u5_mult_87_SUMB_11__13_,
         u5_mult_87_SUMB_11__14_, u5_mult_87_SUMB_11__15_,
         u5_mult_87_SUMB_11__16_, u5_mult_87_SUMB_11__17_,
         u5_mult_87_SUMB_11__18_, u5_mult_87_SUMB_11__19_,
         u5_mult_87_SUMB_11__20_, u5_mult_87_SUMB_11__21_,
         u5_mult_87_SUMB_11__22_, u5_mult_87_SUMB_11__23_,
         u5_mult_87_SUMB_11__24_, u5_mult_87_SUMB_11__25_,
         u5_mult_87_SUMB_11__26_, u5_mult_87_SUMB_11__27_,
         u5_mult_87_SUMB_11__28_, u5_mult_87_SUMB_11__29_,
         u5_mult_87_SUMB_11__30_, u5_mult_87_SUMB_11__31_,
         u5_mult_87_SUMB_11__32_, u5_mult_87_SUMB_11__33_,
         u5_mult_87_SUMB_11__34_, u5_mult_87_SUMB_11__35_,
         u5_mult_87_SUMB_11__36_, u5_mult_87_SUMB_11__37_,
         u5_mult_87_SUMB_11__38_, u5_mult_87_SUMB_11__39_,
         u5_mult_87_SUMB_11__40_, u5_mult_87_SUMB_11__41_,
         u5_mult_87_SUMB_11__42_, u5_mult_87_SUMB_11__43_,
         u5_mult_87_SUMB_11__44_, u5_mult_87_SUMB_11__45_,
         u5_mult_87_SUMB_11__46_, u5_mult_87_SUMB_11__47_,
         u5_mult_87_SUMB_11__48_, u5_mult_87_SUMB_11__49_,
         u5_mult_87_SUMB_11__50_, u5_mult_87_SUMB_11__51_,
         u5_mult_87_SUMB_12__1_, u5_mult_87_SUMB_12__2_,
         u5_mult_87_SUMB_12__3_, u5_mult_87_SUMB_12__4_,
         u5_mult_87_SUMB_12__5_, u5_mult_87_SUMB_12__6_,
         u5_mult_87_SUMB_12__7_, u5_mult_87_SUMB_12__8_,
         u5_mult_87_SUMB_12__9_, u5_mult_87_SUMB_12__10_,
         u5_mult_87_SUMB_12__11_, u5_mult_87_SUMB_12__12_,
         u5_mult_87_SUMB_12__13_, u5_mult_87_SUMB_12__14_,
         u5_mult_87_SUMB_12__15_, u5_mult_87_SUMB_12__16_,
         u5_mult_87_SUMB_12__17_, u5_mult_87_SUMB_12__18_,
         u5_mult_87_SUMB_12__19_, u5_mult_87_SUMB_12__20_,
         u5_mult_87_SUMB_12__21_, u5_mult_87_SUMB_12__22_,
         u5_mult_87_SUMB_12__23_, u5_mult_87_SUMB_12__24_,
         u5_mult_87_SUMB_12__25_, u5_mult_87_SUMB_12__26_,
         u5_mult_87_SUMB_12__27_, u5_mult_87_SUMB_12__28_,
         u5_mult_87_SUMB_12__29_, u5_mult_87_SUMB_12__30_,
         u5_mult_87_SUMB_12__31_, u5_mult_87_SUMB_12__32_,
         u5_mult_87_SUMB_12__33_, u5_mult_87_SUMB_12__34_,
         u5_mult_87_SUMB_12__35_, u5_mult_87_SUMB_12__36_,
         u5_mult_87_SUMB_12__37_, u5_mult_87_SUMB_12__38_,
         u5_mult_87_SUMB_12__39_, u5_mult_87_SUMB_12__40_,
         u5_mult_87_SUMB_12__41_, u5_mult_87_SUMB_12__42_,
         u5_mult_87_SUMB_12__43_, u5_mult_87_SUMB_12__44_,
         u5_mult_87_SUMB_12__45_, u5_mult_87_SUMB_12__46_,
         u5_mult_87_SUMB_12__47_, u5_mult_87_SUMB_12__48_,
         u5_mult_87_SUMB_12__49_, u5_mult_87_SUMB_12__50_,
         u5_mult_87_SUMB_12__51_, u5_mult_87_SUMB_13__1_,
         u5_mult_87_SUMB_13__2_, u5_mult_87_SUMB_13__3_,
         u5_mult_87_SUMB_13__4_, u5_mult_87_SUMB_13__5_,
         u5_mult_87_SUMB_13__6_, u5_mult_87_SUMB_13__7_,
         u5_mult_87_SUMB_13__8_, u5_mult_87_SUMB_13__9_,
         u5_mult_87_SUMB_13__10_, u5_mult_87_SUMB_13__11_,
         u5_mult_87_SUMB_13__12_, u5_mult_87_SUMB_13__13_,
         u5_mult_87_SUMB_13__14_, u5_mult_87_SUMB_13__15_,
         u5_mult_87_SUMB_13__16_, u5_mult_87_SUMB_13__17_,
         u5_mult_87_SUMB_13__18_, u5_mult_87_SUMB_13__19_,
         u5_mult_87_SUMB_13__20_, u5_mult_87_SUMB_13__21_,
         u5_mult_87_SUMB_13__22_, u5_mult_87_SUMB_13__23_,
         u5_mult_87_SUMB_13__24_, u5_mult_87_SUMB_13__25_,
         u5_mult_87_SUMB_13__26_, u5_mult_87_SUMB_13__27_,
         u5_mult_87_SUMB_13__28_, u5_mult_87_SUMB_13__29_,
         u5_mult_87_SUMB_13__30_, u5_mult_87_SUMB_13__31_,
         u5_mult_87_SUMB_13__32_, u5_mult_87_SUMB_13__33_,
         u5_mult_87_SUMB_13__34_, u5_mult_87_SUMB_13__35_,
         u5_mult_87_SUMB_13__36_, u5_mult_87_SUMB_13__37_,
         u5_mult_87_SUMB_13__38_, u5_mult_87_SUMB_13__39_,
         u5_mult_87_SUMB_13__40_, u5_mult_87_SUMB_13__41_,
         u5_mult_87_SUMB_13__42_, u5_mult_87_SUMB_13__43_,
         u5_mult_87_SUMB_13__44_, u5_mult_87_SUMB_13__45_,
         u5_mult_87_SUMB_13__46_, u5_mult_87_SUMB_13__47_,
         u5_mult_87_SUMB_13__48_, u5_mult_87_SUMB_13__49_,
         u5_mult_87_SUMB_13__50_, u5_mult_87_SUMB_13__51_,
         u5_mult_87_SUMB_14__1_, u5_mult_87_SUMB_14__2_,
         u5_mult_87_SUMB_14__3_, u5_mult_87_SUMB_14__4_,
         u5_mult_87_SUMB_14__5_, u5_mult_87_SUMB_14__6_,
         u5_mult_87_SUMB_14__7_, u5_mult_87_SUMB_14__8_,
         u5_mult_87_SUMB_14__9_, u5_mult_87_SUMB_14__10_,
         u5_mult_87_SUMB_14__11_, u5_mult_87_SUMB_14__12_,
         u5_mult_87_SUMB_14__13_, u5_mult_87_SUMB_14__14_,
         u5_mult_87_SUMB_14__15_, u5_mult_87_SUMB_14__16_,
         u5_mult_87_SUMB_14__17_, u5_mult_87_SUMB_14__18_,
         u5_mult_87_CARRYB_4__37_, u5_mult_87_CARRYB_4__38_,
         u5_mult_87_CARRYB_4__39_, u5_mult_87_CARRYB_4__40_,
         u5_mult_87_CARRYB_4__41_, u5_mult_87_CARRYB_4__42_,
         u5_mult_87_CARRYB_4__43_, u5_mult_87_CARRYB_4__44_,
         u5_mult_87_CARRYB_4__45_, u5_mult_87_CARRYB_4__46_,
         u5_mult_87_CARRYB_4__47_, u5_mult_87_CARRYB_4__48_,
         u5_mult_87_CARRYB_4__49_, u5_mult_87_CARRYB_4__50_,
         u5_mult_87_CARRYB_4__51_, u5_mult_87_CARRYB_5__0_,
         u5_mult_87_CARRYB_5__1_, u5_mult_87_CARRYB_5__2_,
         u5_mult_87_CARRYB_5__3_, u5_mult_87_CARRYB_5__4_,
         u5_mult_87_CARRYB_5__5_, u5_mult_87_CARRYB_5__6_,
         u5_mult_87_CARRYB_5__7_, u5_mult_87_CARRYB_5__8_,
         u5_mult_87_CARRYB_5__9_, u5_mult_87_CARRYB_5__10_,
         u5_mult_87_CARRYB_5__11_, u5_mult_87_CARRYB_5__12_,
         u5_mult_87_CARRYB_5__13_, u5_mult_87_CARRYB_5__14_,
         u5_mult_87_CARRYB_5__15_, u5_mult_87_CARRYB_5__16_,
         u5_mult_87_CARRYB_5__17_, u5_mult_87_CARRYB_5__18_,
         u5_mult_87_CARRYB_5__19_, u5_mult_87_CARRYB_5__20_,
         u5_mult_87_CARRYB_5__21_, u5_mult_87_CARRYB_5__22_,
         u5_mult_87_CARRYB_5__23_, u5_mult_87_CARRYB_5__24_,
         u5_mult_87_CARRYB_5__25_, u5_mult_87_CARRYB_5__26_,
         u5_mult_87_CARRYB_5__27_, u5_mult_87_CARRYB_5__28_,
         u5_mult_87_CARRYB_5__29_, u5_mult_87_CARRYB_5__30_,
         u5_mult_87_CARRYB_5__31_, u5_mult_87_CARRYB_5__32_,
         u5_mult_87_CARRYB_5__33_, u5_mult_87_CARRYB_5__34_,
         u5_mult_87_CARRYB_5__35_, u5_mult_87_CARRYB_5__36_,
         u5_mult_87_CARRYB_5__37_, u5_mult_87_CARRYB_5__38_,
         u5_mult_87_CARRYB_5__39_, u5_mult_87_CARRYB_5__40_,
         u5_mult_87_CARRYB_5__41_, u5_mult_87_CARRYB_5__42_,
         u5_mult_87_CARRYB_5__43_, u5_mult_87_CARRYB_5__44_,
         u5_mult_87_CARRYB_5__45_, u5_mult_87_CARRYB_5__46_,
         u5_mult_87_CARRYB_5__47_, u5_mult_87_CARRYB_5__48_,
         u5_mult_87_CARRYB_5__49_, u5_mult_87_CARRYB_5__50_,
         u5_mult_87_CARRYB_5__51_, u5_mult_87_CARRYB_6__0_,
         u5_mult_87_CARRYB_6__1_, u5_mult_87_CARRYB_6__2_,
         u5_mult_87_CARRYB_6__3_, u5_mult_87_CARRYB_6__4_,
         u5_mult_87_CARRYB_6__5_, u5_mult_87_CARRYB_6__6_,
         u5_mult_87_CARRYB_6__7_, u5_mult_87_CARRYB_6__8_,
         u5_mult_87_CARRYB_6__9_, u5_mult_87_CARRYB_6__10_,
         u5_mult_87_CARRYB_6__11_, u5_mult_87_CARRYB_6__12_,
         u5_mult_87_CARRYB_6__13_, u5_mult_87_CARRYB_6__14_,
         u5_mult_87_CARRYB_6__15_, u5_mult_87_CARRYB_6__16_,
         u5_mult_87_CARRYB_6__17_, u5_mult_87_CARRYB_6__18_,
         u5_mult_87_CARRYB_6__19_, u5_mult_87_CARRYB_6__20_,
         u5_mult_87_CARRYB_6__21_, u5_mult_87_CARRYB_6__22_,
         u5_mult_87_CARRYB_6__23_, u5_mult_87_CARRYB_6__24_,
         u5_mult_87_CARRYB_6__25_, u5_mult_87_CARRYB_6__26_,
         u5_mult_87_CARRYB_6__27_, u5_mult_87_CARRYB_6__28_,
         u5_mult_87_CARRYB_6__29_, u5_mult_87_CARRYB_6__30_,
         u5_mult_87_CARRYB_6__31_, u5_mult_87_CARRYB_6__32_,
         u5_mult_87_CARRYB_6__33_, u5_mult_87_CARRYB_6__34_,
         u5_mult_87_CARRYB_6__35_, u5_mult_87_CARRYB_6__36_,
         u5_mult_87_CARRYB_6__37_, u5_mult_87_CARRYB_6__38_,
         u5_mult_87_CARRYB_6__39_, u5_mult_87_CARRYB_6__40_,
         u5_mult_87_CARRYB_6__41_, u5_mult_87_CARRYB_6__42_,
         u5_mult_87_CARRYB_6__43_, u5_mult_87_CARRYB_6__44_,
         u5_mult_87_CARRYB_6__45_, u5_mult_87_CARRYB_6__46_,
         u5_mult_87_CARRYB_6__47_, u5_mult_87_CARRYB_6__48_,
         u5_mult_87_CARRYB_6__49_, u5_mult_87_CARRYB_6__50_,
         u5_mult_87_CARRYB_6__51_, u5_mult_87_CARRYB_7__0_,
         u5_mult_87_CARRYB_7__1_, u5_mult_87_CARRYB_7__2_,
         u5_mult_87_CARRYB_7__3_, u5_mult_87_CARRYB_7__4_,
         u5_mult_87_CARRYB_7__5_, u5_mult_87_CARRYB_7__6_,
         u5_mult_87_CARRYB_7__7_, u5_mult_87_CARRYB_7__8_,
         u5_mult_87_CARRYB_7__9_, u5_mult_87_CARRYB_7__10_,
         u5_mult_87_CARRYB_7__11_, u5_mult_87_CARRYB_7__12_,
         u5_mult_87_CARRYB_7__13_, u5_mult_87_CARRYB_7__14_,
         u5_mult_87_CARRYB_7__15_, u5_mult_87_CARRYB_7__16_,
         u5_mult_87_CARRYB_7__17_, u5_mult_87_CARRYB_7__18_,
         u5_mult_87_CARRYB_7__19_, u5_mult_87_CARRYB_7__20_,
         u5_mult_87_CARRYB_7__21_, u5_mult_87_CARRYB_7__22_,
         u5_mult_87_CARRYB_7__23_, u5_mult_87_CARRYB_7__24_,
         u5_mult_87_CARRYB_7__25_, u5_mult_87_CARRYB_7__26_,
         u5_mult_87_CARRYB_7__27_, u5_mult_87_CARRYB_7__28_,
         u5_mult_87_CARRYB_7__29_, u5_mult_87_CARRYB_7__30_,
         u5_mult_87_CARRYB_7__31_, u5_mult_87_CARRYB_7__32_,
         u5_mult_87_CARRYB_7__33_, u5_mult_87_CARRYB_7__34_,
         u5_mult_87_CARRYB_7__35_, u5_mult_87_CARRYB_7__36_,
         u5_mult_87_CARRYB_7__37_, u5_mult_87_CARRYB_7__38_,
         u5_mult_87_CARRYB_7__39_, u5_mult_87_CARRYB_7__40_,
         u5_mult_87_CARRYB_7__41_, u5_mult_87_CARRYB_7__42_,
         u5_mult_87_CARRYB_7__43_, u5_mult_87_CARRYB_7__44_,
         u5_mult_87_CARRYB_7__45_, u5_mult_87_CARRYB_7__46_,
         u5_mult_87_CARRYB_7__47_, u5_mult_87_CARRYB_7__48_,
         u5_mult_87_CARRYB_7__49_, u5_mult_87_CARRYB_7__50_,
         u5_mult_87_CARRYB_7__51_, u5_mult_87_CARRYB_8__0_,
         u5_mult_87_CARRYB_8__1_, u5_mult_87_CARRYB_8__2_,
         u5_mult_87_CARRYB_8__3_, u5_mult_87_CARRYB_8__4_,
         u5_mult_87_CARRYB_8__5_, u5_mult_87_CARRYB_8__6_,
         u5_mult_87_CARRYB_8__7_, u5_mult_87_CARRYB_8__8_,
         u5_mult_87_CARRYB_8__9_, u5_mult_87_CARRYB_8__10_,
         u5_mult_87_CARRYB_8__11_, u5_mult_87_CARRYB_8__12_,
         u5_mult_87_CARRYB_8__13_, u5_mult_87_CARRYB_8__14_,
         u5_mult_87_CARRYB_8__15_, u5_mult_87_CARRYB_8__16_,
         u5_mult_87_CARRYB_8__17_, u5_mult_87_CARRYB_8__18_,
         u5_mult_87_CARRYB_8__19_, u5_mult_87_CARRYB_8__20_,
         u5_mult_87_CARRYB_8__21_, u5_mult_87_CARRYB_8__22_,
         u5_mult_87_CARRYB_8__23_, u5_mult_87_CARRYB_8__24_,
         u5_mult_87_CARRYB_8__25_, u5_mult_87_CARRYB_8__26_,
         u5_mult_87_CARRYB_8__27_, u5_mult_87_CARRYB_8__28_,
         u5_mult_87_CARRYB_8__29_, u5_mult_87_CARRYB_8__30_,
         u5_mult_87_CARRYB_8__31_, u5_mult_87_CARRYB_8__32_,
         u5_mult_87_CARRYB_8__33_, u5_mult_87_CARRYB_8__34_,
         u5_mult_87_CARRYB_8__35_, u5_mult_87_CARRYB_8__36_,
         u5_mult_87_CARRYB_8__37_, u5_mult_87_CARRYB_8__38_,
         u5_mult_87_CARRYB_8__39_, u5_mult_87_CARRYB_8__40_,
         u5_mult_87_CARRYB_8__41_, u5_mult_87_CARRYB_8__42_,
         u5_mult_87_CARRYB_8__43_, u5_mult_87_CARRYB_8__44_,
         u5_mult_87_CARRYB_8__45_, u5_mult_87_CARRYB_8__46_,
         u5_mult_87_CARRYB_8__47_, u5_mult_87_CARRYB_8__48_,
         u5_mult_87_CARRYB_8__49_, u5_mult_87_CARRYB_8__50_,
         u5_mult_87_CARRYB_8__51_, u5_mult_87_CARRYB_9__0_,
         u5_mult_87_CARRYB_9__1_, u5_mult_87_CARRYB_9__2_,
         u5_mult_87_CARRYB_9__3_, u5_mult_87_CARRYB_9__4_,
         u5_mult_87_CARRYB_9__5_, u5_mult_87_CARRYB_9__6_,
         u5_mult_87_CARRYB_9__7_, u5_mult_87_CARRYB_9__8_,
         u5_mult_87_CARRYB_9__9_, u5_mult_87_CARRYB_9__10_,
         u5_mult_87_CARRYB_9__11_, u5_mult_87_CARRYB_9__12_,
         u5_mult_87_CARRYB_9__13_, u5_mult_87_CARRYB_9__14_,
         u5_mult_87_CARRYB_9__15_, u5_mult_87_CARRYB_9__16_,
         u5_mult_87_CARRYB_9__17_, u5_mult_87_CARRYB_9__18_,
         u5_mult_87_CARRYB_9__19_, u5_mult_87_CARRYB_9__20_,
         u5_mult_87_CARRYB_9__21_, u5_mult_87_CARRYB_9__22_,
         u5_mult_87_CARRYB_9__23_, u5_mult_87_CARRYB_9__24_,
         u5_mult_87_CARRYB_9__25_, u5_mult_87_CARRYB_9__26_,
         u5_mult_87_CARRYB_9__27_, u5_mult_87_CARRYB_9__28_,
         u5_mult_87_CARRYB_9__29_, u5_mult_87_CARRYB_9__30_,
         u5_mult_87_CARRYB_9__31_, u5_mult_87_CARRYB_9__32_,
         u5_mult_87_CARRYB_9__33_, u5_mult_87_CARRYB_9__34_,
         u5_mult_87_CARRYB_9__35_, u5_mult_87_CARRYB_9__36_,
         u5_mult_87_CARRYB_9__37_, u5_mult_87_CARRYB_9__38_,
         u5_mult_87_CARRYB_9__39_, u5_mult_87_CARRYB_9__40_,
         u5_mult_87_CARRYB_9__41_, u5_mult_87_CARRYB_9__42_,
         u5_mult_87_CARRYB_9__43_, u5_mult_87_CARRYB_9__44_,
         u5_mult_87_CARRYB_9__45_, u5_mult_87_CARRYB_9__46_,
         u5_mult_87_CARRYB_9__47_, u5_mult_87_CARRYB_9__48_,
         u5_mult_87_CARRYB_9__49_, u5_mult_87_CARRYB_9__50_,
         u5_mult_87_CARRYB_9__51_, u5_mult_87_CARRYB_10__0_,
         u5_mult_87_CARRYB_10__1_, u5_mult_87_CARRYB_10__2_,
         u5_mult_87_CARRYB_10__3_, u5_mult_87_CARRYB_10__4_,
         u5_mult_87_CARRYB_10__5_, u5_mult_87_CARRYB_10__6_,
         u5_mult_87_CARRYB_10__7_, u5_mult_87_CARRYB_10__8_,
         u5_mult_87_CARRYB_10__9_, u5_mult_87_CARRYB_10__10_,
         u5_mult_87_CARRYB_10__11_, u5_mult_87_CARRYB_10__12_,
         u5_mult_87_CARRYB_10__13_, u5_mult_87_CARRYB_10__14_,
         u5_mult_87_CARRYB_10__15_, u5_mult_87_CARRYB_10__16_,
         u5_mult_87_CARRYB_10__17_, u5_mult_87_CARRYB_10__18_,
         u5_mult_87_CARRYB_10__19_, u5_mult_87_CARRYB_10__20_,
         u5_mult_87_CARRYB_10__21_, u5_mult_87_CARRYB_10__22_,
         u5_mult_87_CARRYB_10__23_, u5_mult_87_CARRYB_10__24_,
         u5_mult_87_CARRYB_10__25_, u5_mult_87_CARRYB_10__26_,
         u5_mult_87_CARRYB_10__27_, u5_mult_87_CARRYB_10__28_,
         u5_mult_87_CARRYB_10__29_, u5_mult_87_CARRYB_10__30_,
         u5_mult_87_CARRYB_10__31_, u5_mult_87_CARRYB_10__32_,
         u5_mult_87_CARRYB_10__33_, u5_mult_87_CARRYB_10__34_,
         u5_mult_87_CARRYB_10__35_, u5_mult_87_CARRYB_10__36_,
         u5_mult_87_CARRYB_10__37_, u5_mult_87_CARRYB_10__38_,
         u5_mult_87_CARRYB_10__39_, u5_mult_87_CARRYB_10__40_,
         u5_mult_87_CARRYB_10__41_, u5_mult_87_CARRYB_10__42_,
         u5_mult_87_CARRYB_10__43_, u5_mult_87_CARRYB_10__44_,
         u5_mult_87_CARRYB_10__45_, u5_mult_87_CARRYB_10__46_,
         u5_mult_87_CARRYB_10__47_, u5_mult_87_CARRYB_10__48_,
         u5_mult_87_CARRYB_10__49_, u5_mult_87_CARRYB_10__50_,
         u5_mult_87_CARRYB_10__51_, u5_mult_87_CARRYB_11__0_,
         u5_mult_87_CARRYB_11__1_, u5_mult_87_CARRYB_11__2_,
         u5_mult_87_CARRYB_11__3_, u5_mult_87_CARRYB_11__4_,
         u5_mult_87_CARRYB_11__5_, u5_mult_87_CARRYB_11__6_,
         u5_mult_87_CARRYB_11__7_, u5_mult_87_CARRYB_11__8_,
         u5_mult_87_CARRYB_11__9_, u5_mult_87_CARRYB_11__10_,
         u5_mult_87_CARRYB_11__11_, u5_mult_87_CARRYB_11__12_,
         u5_mult_87_CARRYB_11__13_, u5_mult_87_CARRYB_11__14_,
         u5_mult_87_CARRYB_11__15_, u5_mult_87_CARRYB_11__16_,
         u5_mult_87_CARRYB_11__17_, u5_mult_87_CARRYB_11__18_,
         u5_mult_87_CARRYB_11__19_, u5_mult_87_CARRYB_11__20_,
         u5_mult_87_CARRYB_11__21_, u5_mult_87_CARRYB_11__22_,
         u5_mult_87_CARRYB_11__23_, u5_mult_87_CARRYB_11__24_,
         u5_mult_87_CARRYB_11__25_, u5_mult_87_CARRYB_11__26_,
         u5_mult_87_CARRYB_11__27_, u5_mult_87_CARRYB_11__28_,
         u5_mult_87_CARRYB_11__29_, u5_mult_87_CARRYB_11__30_,
         u5_mult_87_CARRYB_11__31_, u5_mult_87_CARRYB_11__32_,
         u5_mult_87_CARRYB_11__33_, u5_mult_87_CARRYB_11__34_,
         u5_mult_87_CARRYB_11__35_, u5_mult_87_CARRYB_11__36_,
         u5_mult_87_CARRYB_11__37_, u5_mult_87_CARRYB_11__38_,
         u5_mult_87_CARRYB_11__39_, u5_mult_87_CARRYB_11__40_,
         u5_mult_87_CARRYB_11__41_, u5_mult_87_CARRYB_11__42_,
         u5_mult_87_CARRYB_11__43_, u5_mult_87_CARRYB_11__44_,
         u5_mult_87_CARRYB_11__45_, u5_mult_87_CARRYB_11__46_,
         u5_mult_87_CARRYB_11__47_, u5_mult_87_CARRYB_11__48_,
         u5_mult_87_CARRYB_11__49_, u5_mult_87_CARRYB_11__50_,
         u5_mult_87_CARRYB_11__51_, u5_mult_87_CARRYB_12__0_,
         u5_mult_87_CARRYB_12__1_, u5_mult_87_CARRYB_12__2_,
         u5_mult_87_CARRYB_12__3_, u5_mult_87_CARRYB_12__4_,
         u5_mult_87_CARRYB_12__5_, u5_mult_87_CARRYB_12__6_,
         u5_mult_87_CARRYB_12__7_, u5_mult_87_CARRYB_12__8_,
         u5_mult_87_CARRYB_12__9_, u5_mult_87_CARRYB_12__10_,
         u5_mult_87_CARRYB_12__11_, u5_mult_87_CARRYB_12__12_,
         u5_mult_87_CARRYB_12__13_, u5_mult_87_CARRYB_12__14_,
         u5_mult_87_CARRYB_12__15_, u5_mult_87_CARRYB_12__16_,
         u5_mult_87_CARRYB_12__17_, u5_mult_87_CARRYB_12__18_,
         u5_mult_87_CARRYB_12__19_, u5_mult_87_CARRYB_12__20_,
         u5_mult_87_CARRYB_12__21_, u5_mult_87_CARRYB_12__22_,
         u5_mult_87_CARRYB_12__23_, u5_mult_87_CARRYB_12__24_,
         u5_mult_87_CARRYB_12__25_, u5_mult_87_CARRYB_12__26_,
         u5_mult_87_CARRYB_12__27_, u5_mult_87_CARRYB_12__28_,
         u5_mult_87_CARRYB_12__29_, u5_mult_87_CARRYB_12__30_,
         u5_mult_87_CARRYB_12__31_, u5_mult_87_CARRYB_12__32_,
         u5_mult_87_CARRYB_12__33_, u5_mult_87_CARRYB_12__34_,
         u5_mult_87_CARRYB_12__35_, u5_mult_87_CARRYB_12__36_,
         u5_mult_87_CARRYB_12__37_, u5_mult_87_CARRYB_12__38_,
         u5_mult_87_CARRYB_12__39_, u5_mult_87_CARRYB_12__40_,
         u5_mult_87_CARRYB_12__41_, u5_mult_87_CARRYB_12__42_,
         u5_mult_87_CARRYB_12__43_, u5_mult_87_CARRYB_12__44_,
         u5_mult_87_CARRYB_12__45_, u5_mult_87_CARRYB_12__46_,
         u5_mult_87_CARRYB_12__47_, u5_mult_87_CARRYB_12__48_,
         u5_mult_87_CARRYB_12__49_, u5_mult_87_CARRYB_12__50_,
         u5_mult_87_CARRYB_12__51_, u5_mult_87_CARRYB_13__0_,
         u5_mult_87_CARRYB_13__1_, u5_mult_87_CARRYB_13__2_,
         u5_mult_87_CARRYB_13__3_, u5_mult_87_CARRYB_13__4_,
         u5_mult_87_CARRYB_13__5_, u5_mult_87_CARRYB_13__6_,
         u5_mult_87_CARRYB_13__7_, u5_mult_87_CARRYB_13__8_,
         u5_mult_87_CARRYB_13__9_, u5_mult_87_CARRYB_13__10_,
         u5_mult_87_CARRYB_13__11_, u5_mult_87_CARRYB_13__12_,
         u5_mult_87_CARRYB_13__13_, u5_mult_87_CARRYB_13__14_,
         u5_mult_87_CARRYB_13__15_, u5_mult_87_CARRYB_13__16_,
         u5_mult_87_CARRYB_13__17_, u5_mult_87_CARRYB_13__18_,
         u5_mult_87_CARRYB_13__19_, u5_mult_87_CARRYB_13__20_,
         u5_mult_87_CARRYB_13__21_, u5_mult_87_CARRYB_13__22_,
         u5_mult_87_CARRYB_13__23_, u5_mult_87_CARRYB_13__24_,
         u5_mult_87_CARRYB_13__25_, u5_mult_87_CARRYB_13__26_,
         u5_mult_87_CARRYB_13__27_, u5_mult_87_CARRYB_13__28_,
         u5_mult_87_CARRYB_13__29_, u5_mult_87_CARRYB_13__30_,
         u5_mult_87_CARRYB_13__31_, u5_mult_87_CARRYB_13__32_,
         u5_mult_87_CARRYB_13__33_, u5_mult_87_CARRYB_13__34_,
         u5_mult_87_CARRYB_13__35_, u5_mult_87_CARRYB_13__36_,
         u5_mult_87_CARRYB_13__37_, u5_mult_87_CARRYB_13__38_,
         u5_mult_87_CARRYB_13__39_, u5_mult_87_CARRYB_13__40_,
         u5_mult_87_CARRYB_13__41_, u5_mult_87_CARRYB_13__42_,
         u5_mult_87_CARRYB_13__43_, u5_mult_87_CARRYB_13__44_,
         u5_mult_87_CARRYB_13__45_, u5_mult_87_CARRYB_13__46_,
         u5_mult_87_CARRYB_13__47_, u5_mult_87_CARRYB_13__48_,
         u5_mult_87_CARRYB_13__49_, u5_mult_87_CARRYB_13__50_,
         u5_mult_87_CARRYB_13__51_, u5_mult_87_CARRYB_14__0_,
         u5_mult_87_CARRYB_14__1_, u5_mult_87_CARRYB_14__2_,
         u5_mult_87_CARRYB_14__3_, u5_mult_87_CARRYB_14__4_,
         u5_mult_87_CARRYB_14__5_, u5_mult_87_CARRYB_14__6_,
         u5_mult_87_CARRYB_14__7_, u5_mult_87_CARRYB_14__8_,
         u5_mult_87_CARRYB_14__9_, u5_mult_87_CARRYB_14__10_,
         u5_mult_87_CARRYB_14__11_, u5_mult_87_CARRYB_14__12_,
         u5_mult_87_CARRYB_14__13_, u5_mult_87_CARRYB_14__14_,
         u5_mult_87_CARRYB_14__15_, u5_mult_87_CARRYB_14__16_,
         u5_mult_87_CARRYB_14__17_, u5_mult_87_CARRYB_14__18_,
         u5_mult_87_SUMB_2__1_, u5_mult_87_SUMB_2__2_, u5_mult_87_SUMB_2__3_,
         u5_mult_87_SUMB_2__4_, u5_mult_87_SUMB_2__5_, u5_mult_87_SUMB_2__6_,
         u5_mult_87_SUMB_2__7_, u5_mult_87_SUMB_2__8_, u5_mult_87_SUMB_2__9_,
         u5_mult_87_SUMB_2__10_, u5_mult_87_SUMB_2__11_,
         u5_mult_87_SUMB_2__12_, u5_mult_87_SUMB_2__13_,
         u5_mult_87_SUMB_2__14_, u5_mult_87_SUMB_2__15_,
         u5_mult_87_SUMB_2__16_, u5_mult_87_SUMB_2__17_,
         u5_mult_87_SUMB_2__18_, u5_mult_87_SUMB_2__19_,
         u5_mult_87_SUMB_2__20_, u5_mult_87_SUMB_2__21_,
         u5_mult_87_SUMB_2__22_, u5_mult_87_SUMB_2__23_,
         u5_mult_87_SUMB_2__24_, u5_mult_87_SUMB_2__25_,
         u5_mult_87_SUMB_2__26_, u5_mult_87_SUMB_2__27_,
         u5_mult_87_SUMB_2__28_, u5_mult_87_SUMB_2__29_,
         u5_mult_87_SUMB_2__30_, u5_mult_87_SUMB_2__31_,
         u5_mult_87_SUMB_2__32_, u5_mult_87_SUMB_2__33_,
         u5_mult_87_SUMB_2__34_, u5_mult_87_SUMB_2__35_,
         u5_mult_87_SUMB_2__36_, u5_mult_87_SUMB_2__37_,
         u5_mult_87_SUMB_2__38_, u5_mult_87_SUMB_2__39_,
         u5_mult_87_SUMB_2__40_, u5_mult_87_SUMB_2__41_,
         u5_mult_87_SUMB_2__42_, u5_mult_87_SUMB_2__43_,
         u5_mult_87_SUMB_2__44_, u5_mult_87_SUMB_2__45_,
         u5_mult_87_SUMB_2__46_, u5_mult_87_SUMB_2__47_,
         u5_mult_87_SUMB_2__48_, u5_mult_87_SUMB_2__49_,
         u5_mult_87_SUMB_2__50_, u5_mult_87_SUMB_2__51_, u5_mult_87_SUMB_3__1_,
         u5_mult_87_SUMB_3__2_, u5_mult_87_SUMB_3__3_, u5_mult_87_SUMB_3__4_,
         u5_mult_87_SUMB_3__5_, u5_mult_87_SUMB_3__6_, u5_mult_87_SUMB_3__7_,
         u5_mult_87_SUMB_3__8_, u5_mult_87_SUMB_3__9_, u5_mult_87_SUMB_3__10_,
         u5_mult_87_SUMB_3__11_, u5_mult_87_SUMB_3__12_,
         u5_mult_87_SUMB_3__13_, u5_mult_87_SUMB_3__14_,
         u5_mult_87_SUMB_3__15_, u5_mult_87_SUMB_3__16_,
         u5_mult_87_SUMB_3__17_, u5_mult_87_SUMB_3__18_,
         u5_mult_87_SUMB_3__19_, u5_mult_87_SUMB_3__20_,
         u5_mult_87_SUMB_3__21_, u5_mult_87_SUMB_3__22_,
         u5_mult_87_SUMB_3__23_, u5_mult_87_SUMB_3__24_,
         u5_mult_87_SUMB_3__25_, u5_mult_87_SUMB_3__26_,
         u5_mult_87_SUMB_3__27_, u5_mult_87_SUMB_3__28_,
         u5_mult_87_SUMB_3__29_, u5_mult_87_SUMB_3__30_,
         u5_mult_87_SUMB_3__31_, u5_mult_87_SUMB_3__32_,
         u5_mult_87_SUMB_3__33_, u5_mult_87_SUMB_3__34_,
         u5_mult_87_SUMB_3__35_, u5_mult_87_SUMB_3__36_,
         u5_mult_87_SUMB_3__37_, u5_mult_87_SUMB_3__38_,
         u5_mult_87_SUMB_3__39_, u5_mult_87_SUMB_3__40_,
         u5_mult_87_SUMB_3__41_, u5_mult_87_SUMB_3__42_,
         u5_mult_87_SUMB_3__43_, u5_mult_87_SUMB_3__44_,
         u5_mult_87_SUMB_3__45_, u5_mult_87_SUMB_3__46_,
         u5_mult_87_SUMB_3__47_, u5_mult_87_SUMB_3__48_,
         u5_mult_87_SUMB_3__49_, u5_mult_87_SUMB_3__50_,
         u5_mult_87_SUMB_3__51_, u5_mult_87_SUMB_4__1_, u5_mult_87_SUMB_4__2_,
         u5_mult_87_SUMB_4__3_, u5_mult_87_SUMB_4__4_, u5_mult_87_SUMB_4__5_,
         u5_mult_87_SUMB_4__6_, u5_mult_87_SUMB_4__7_, u5_mult_87_SUMB_4__8_,
         u5_mult_87_SUMB_4__9_, u5_mult_87_SUMB_4__10_, u5_mult_87_SUMB_4__11_,
         u5_mult_87_SUMB_4__12_, u5_mult_87_SUMB_4__13_,
         u5_mult_87_SUMB_4__14_, u5_mult_87_SUMB_4__15_,
         u5_mult_87_SUMB_4__16_, u5_mult_87_SUMB_4__17_,
         u5_mult_87_SUMB_4__18_, u5_mult_87_SUMB_4__19_,
         u5_mult_87_SUMB_4__20_, u5_mult_87_SUMB_4__21_,
         u5_mult_87_SUMB_4__22_, u5_mult_87_SUMB_4__23_,
         u5_mult_87_SUMB_4__24_, u5_mult_87_SUMB_4__25_,
         u5_mult_87_SUMB_4__26_, u5_mult_87_SUMB_4__27_,
         u5_mult_87_SUMB_4__28_, u5_mult_87_SUMB_4__29_,
         u5_mult_87_SUMB_4__30_, u5_mult_87_SUMB_4__31_,
         u5_mult_87_SUMB_4__32_, u5_mult_87_SUMB_4__33_,
         u5_mult_87_SUMB_4__34_, u5_mult_87_SUMB_4__35_,
         u5_mult_87_SUMB_4__36_, u5_mult_87_CARRYB_2__0_,
         u5_mult_87_CARRYB_2__1_, u5_mult_87_CARRYB_2__2_,
         u5_mult_87_CARRYB_2__3_, u5_mult_87_CARRYB_2__4_,
         u5_mult_87_CARRYB_2__5_, u5_mult_87_CARRYB_2__6_,
         u5_mult_87_CARRYB_2__7_, u5_mult_87_CARRYB_2__8_,
         u5_mult_87_CARRYB_2__9_, u5_mult_87_CARRYB_2__10_,
         u5_mult_87_CARRYB_2__11_, u5_mult_87_CARRYB_2__12_,
         u5_mult_87_CARRYB_2__13_, u5_mult_87_CARRYB_2__14_,
         u5_mult_87_CARRYB_2__15_, u5_mult_87_CARRYB_2__16_,
         u5_mult_87_CARRYB_2__17_, u5_mult_87_CARRYB_2__18_,
         u5_mult_87_CARRYB_2__19_, u5_mult_87_CARRYB_2__20_,
         u5_mult_87_CARRYB_2__21_, u5_mult_87_CARRYB_2__22_,
         u5_mult_87_CARRYB_2__23_, u5_mult_87_CARRYB_2__24_,
         u5_mult_87_CARRYB_2__25_, u5_mult_87_CARRYB_2__26_,
         u5_mult_87_CARRYB_2__27_, u5_mult_87_CARRYB_2__28_,
         u5_mult_87_CARRYB_2__29_, u5_mult_87_CARRYB_2__30_,
         u5_mult_87_CARRYB_2__31_, u5_mult_87_CARRYB_2__32_,
         u5_mult_87_CARRYB_2__33_, u5_mult_87_CARRYB_2__34_,
         u5_mult_87_CARRYB_2__35_, u5_mult_87_CARRYB_2__36_,
         u5_mult_87_CARRYB_2__37_, u5_mult_87_CARRYB_2__38_,
         u5_mult_87_CARRYB_2__39_, u5_mult_87_CARRYB_2__40_,
         u5_mult_87_CARRYB_2__41_, u5_mult_87_CARRYB_2__42_,
         u5_mult_87_CARRYB_2__43_, u5_mult_87_CARRYB_2__44_,
         u5_mult_87_CARRYB_2__45_, u5_mult_87_CARRYB_2__46_,
         u5_mult_87_CARRYB_2__47_, u5_mult_87_CARRYB_2__48_,
         u5_mult_87_CARRYB_2__49_, u5_mult_87_CARRYB_2__50_,
         u5_mult_87_CARRYB_2__51_, u5_mult_87_CARRYB_3__0_,
         u5_mult_87_CARRYB_3__1_, u5_mult_87_CARRYB_3__2_,
         u5_mult_87_CARRYB_3__3_, u5_mult_87_CARRYB_3__4_,
         u5_mult_87_CARRYB_3__5_, u5_mult_87_CARRYB_3__6_,
         u5_mult_87_CARRYB_3__7_, u5_mult_87_CARRYB_3__8_,
         u5_mult_87_CARRYB_3__9_, u5_mult_87_CARRYB_3__10_,
         u5_mult_87_CARRYB_3__11_, u5_mult_87_CARRYB_3__12_,
         u5_mult_87_CARRYB_3__13_, u5_mult_87_CARRYB_3__14_,
         u5_mult_87_CARRYB_3__15_, u5_mult_87_CARRYB_3__16_,
         u5_mult_87_CARRYB_3__17_, u5_mult_87_CARRYB_3__18_,
         u5_mult_87_CARRYB_3__19_, u5_mult_87_CARRYB_3__20_,
         u5_mult_87_CARRYB_3__21_, u5_mult_87_CARRYB_3__22_,
         u5_mult_87_CARRYB_3__23_, u5_mult_87_CARRYB_3__24_,
         u5_mult_87_CARRYB_3__25_, u5_mult_87_CARRYB_3__26_,
         u5_mult_87_CARRYB_3__27_, u5_mult_87_CARRYB_3__28_,
         u5_mult_87_CARRYB_3__29_, u5_mult_87_CARRYB_3__30_,
         u5_mult_87_CARRYB_3__31_, u5_mult_87_CARRYB_3__32_,
         u5_mult_87_CARRYB_3__33_, u5_mult_87_CARRYB_3__34_,
         u5_mult_87_CARRYB_3__35_, u5_mult_87_CARRYB_3__36_,
         u5_mult_87_CARRYB_3__37_, u5_mult_87_CARRYB_3__38_,
         u5_mult_87_CARRYB_3__39_, u5_mult_87_CARRYB_3__40_,
         u5_mult_87_CARRYB_3__41_, u5_mult_87_CARRYB_3__42_,
         u5_mult_87_CARRYB_3__43_, u5_mult_87_CARRYB_3__44_,
         u5_mult_87_CARRYB_3__45_, u5_mult_87_CARRYB_3__46_,
         u5_mult_87_CARRYB_3__47_, u5_mult_87_CARRYB_3__48_,
         u5_mult_87_CARRYB_3__49_, u5_mult_87_CARRYB_3__50_,
         u5_mult_87_CARRYB_3__51_, u5_mult_87_CARRYB_4__0_,
         u5_mult_87_CARRYB_4__1_, u5_mult_87_CARRYB_4__2_,
         u5_mult_87_CARRYB_4__3_, u5_mult_87_CARRYB_4__4_,
         u5_mult_87_CARRYB_4__5_, u5_mult_87_CARRYB_4__6_,
         u5_mult_87_CARRYB_4__7_, u5_mult_87_CARRYB_4__8_,
         u5_mult_87_CARRYB_4__9_, u5_mult_87_CARRYB_4__10_,
         u5_mult_87_CARRYB_4__11_, u5_mult_87_CARRYB_4__12_,
         u5_mult_87_CARRYB_4__13_, u5_mult_87_CARRYB_4__14_,
         u5_mult_87_CARRYB_4__15_, u5_mult_87_CARRYB_4__16_,
         u5_mult_87_CARRYB_4__17_, u5_mult_87_CARRYB_4__18_,
         u5_mult_87_CARRYB_4__19_, u5_mult_87_CARRYB_4__20_,
         u5_mult_87_CARRYB_4__21_, u5_mult_87_CARRYB_4__22_,
         u5_mult_87_CARRYB_4__23_, u5_mult_87_CARRYB_4__24_,
         u5_mult_87_CARRYB_4__25_, u5_mult_87_CARRYB_4__26_,
         u5_mult_87_CARRYB_4__27_, u5_mult_87_CARRYB_4__28_,
         u5_mult_87_CARRYB_4__29_, u5_mult_87_CARRYB_4__30_,
         u5_mult_87_CARRYB_4__31_, u5_mult_87_CARRYB_4__32_,
         u5_mult_87_CARRYB_4__33_, u5_mult_87_CARRYB_4__34_,
         u5_mult_87_CARRYB_4__35_, u5_mult_87_CARRYB_4__36_,
         u5_mult_87_ab_0__1_, u5_mult_87_ab_0__2_, u5_mult_87_ab_0__3_,
         u5_mult_87_ab_0__4_, u5_mult_87_ab_0__5_, u5_mult_87_ab_0__6_,
         u5_mult_87_ab_0__7_, u5_mult_87_ab_0__8_, u5_mult_87_ab_0__9_,
         u5_mult_87_ab_0__10_, u5_mult_87_ab_0__11_, u5_mult_87_ab_0__12_,
         u5_mult_87_ab_0__13_, u5_mult_87_ab_0__14_, u5_mult_87_ab_0__15_,
         u5_mult_87_ab_0__16_, u5_mult_87_ab_0__17_, u5_mult_87_ab_0__18_,
         u5_mult_87_ab_0__19_, u5_mult_87_ab_0__20_, u5_mult_87_ab_0__21_,
         u5_mult_87_ab_0__22_, u5_mult_87_ab_0__23_, u5_mult_87_ab_0__24_,
         u5_mult_87_ab_0__25_, u5_mult_87_ab_0__26_, u5_mult_87_ab_0__27_,
         u5_mult_87_ab_0__28_, u5_mult_87_ab_0__29_, u5_mult_87_ab_0__30_,
         u5_mult_87_ab_0__31_, u5_mult_87_ab_0__32_, u5_mult_87_ab_0__33_,
         u5_mult_87_ab_0__34_, u5_mult_87_ab_0__35_, u5_mult_87_ab_0__36_,
         u5_mult_87_ab_0__37_, u5_mult_87_ab_0__38_, u5_mult_87_ab_0__39_,
         u5_mult_87_ab_0__40_, u5_mult_87_ab_0__41_, u5_mult_87_ab_0__42_,
         u5_mult_87_ab_0__43_, u5_mult_87_ab_0__44_, u5_mult_87_ab_0__45_,
         u5_mult_87_ab_0__46_, u5_mult_87_ab_0__47_, u5_mult_87_ab_0__48_,
         u5_mult_87_ab_0__49_, u5_mult_87_ab_0__50_, u5_mult_87_ab_0__51_,
         u5_mult_87_ab_0__52_, u5_mult_87_ab_1__0_, u5_mult_87_ab_1__1_,
         u5_mult_87_ab_1__2_, u5_mult_87_ab_1__3_, u5_mult_87_ab_1__4_,
         u5_mult_87_ab_1__5_, u5_mult_87_ab_1__6_, u5_mult_87_ab_1__7_,
         u5_mult_87_ab_1__8_, u5_mult_87_ab_1__9_, u5_mult_87_ab_1__10_,
         u5_mult_87_ab_1__11_, u5_mult_87_ab_1__12_, u5_mult_87_ab_1__13_,
         u5_mult_87_ab_1__14_, u5_mult_87_ab_1__15_, u5_mult_87_ab_1__16_,
         u5_mult_87_ab_1__17_, u5_mult_87_ab_1__18_, u5_mult_87_ab_1__19_,
         u5_mult_87_ab_1__20_, u5_mult_87_ab_1__21_, u5_mult_87_ab_1__22_,
         u5_mult_87_ab_1__23_, u5_mult_87_ab_1__24_, u5_mult_87_ab_1__25_,
         u5_mult_87_ab_1__26_, u5_mult_87_ab_1__27_, u5_mult_87_ab_1__28_,
         u5_mult_87_ab_1__29_, u5_mult_87_ab_1__30_, u5_mult_87_ab_1__31_,
         u5_mult_87_ab_1__32_, u5_mult_87_ab_1__33_, u5_mult_87_ab_1__34_,
         u5_mult_87_ab_1__35_, u5_mult_87_ab_1__36_, u5_mult_87_ab_1__37_,
         u5_mult_87_ab_1__38_, u5_mult_87_ab_1__39_, u5_mult_87_ab_1__40_,
         u5_mult_87_ab_1__41_, u5_mult_87_ab_1__42_, u5_mult_87_ab_1__43_,
         u5_mult_87_ab_1__44_, u5_mult_87_ab_1__45_, u5_mult_87_ab_1__46_,
         u5_mult_87_ab_1__47_, u5_mult_87_ab_1__48_, u5_mult_87_ab_1__49_,
         u5_mult_87_ab_1__50_, u5_mult_87_ab_1__51_, u5_mult_87_ab_1__52_,
         u5_mult_87_ab_2__0_, u5_mult_87_ab_2__1_, u5_mult_87_ab_2__2_,
         u5_mult_87_ab_2__3_, u5_mult_87_ab_2__4_, u5_mult_87_ab_2__5_,
         u5_mult_87_ab_2__6_, u5_mult_87_ab_2__7_, u5_mult_87_ab_2__8_,
         u5_mult_87_ab_2__9_, u5_mult_87_ab_2__10_, u5_mult_87_ab_2__11_,
         u5_mult_87_ab_2__12_, u5_mult_87_ab_2__13_, u5_mult_87_ab_2__14_,
         u5_mult_87_ab_2__15_, u5_mult_87_ab_2__16_, u5_mult_87_ab_2__17_,
         u5_mult_87_ab_2__18_, u5_mult_87_ab_2__19_, u5_mult_87_ab_2__20_,
         u5_mult_87_ab_2__21_, u5_mult_87_ab_2__22_, u5_mult_87_ab_2__23_,
         u5_mult_87_ab_2__24_, u5_mult_87_ab_2__25_, u5_mult_87_ab_2__26_,
         u5_mult_87_ab_2__27_, u5_mult_87_ab_2__28_, u5_mult_87_ab_2__29_,
         u5_mult_87_ab_2__30_, u5_mult_87_ab_2__31_, u5_mult_87_ab_2__32_,
         u5_mult_87_ab_2__33_, u5_mult_87_ab_2__34_, u5_mult_87_ab_2__35_,
         u5_mult_87_ab_2__36_, u5_mult_87_ab_2__37_, u5_mult_87_ab_2__38_,
         u5_mult_87_ab_2__39_, u5_mult_87_ab_2__40_, u5_mult_87_ab_2__41_,
         u5_mult_87_ab_2__42_, u5_mult_87_ab_2__43_, u5_mult_87_ab_2__44_,
         u5_mult_87_ab_2__45_, u5_mult_87_ab_2__46_, u5_mult_87_ab_2__47_,
         u5_mult_87_ab_2__48_, u5_mult_87_ab_2__49_, u5_mult_87_ab_2__50_,
         u5_mult_87_ab_2__51_, u5_mult_87_ab_2__52_, u5_mult_87_ab_3__0_,
         u5_mult_87_ab_3__1_, u5_mult_87_ab_3__2_, u5_mult_87_ab_3__3_,
         u5_mult_87_ab_3__4_, u5_mult_87_ab_3__5_, u5_mult_87_ab_3__6_,
         u5_mult_87_ab_3__7_, u5_mult_87_ab_3__8_, u5_mult_87_ab_3__9_,
         u5_mult_87_ab_3__10_, u5_mult_87_ab_3__11_, u5_mult_87_ab_3__12_,
         u5_mult_87_ab_3__13_, u5_mult_87_ab_3__14_, u5_mult_87_ab_3__15_,
         u5_mult_87_ab_3__16_, u5_mult_87_ab_3__17_, u5_mult_87_ab_3__18_,
         u5_mult_87_ab_3__19_, u5_mult_87_ab_3__20_, u5_mult_87_ab_3__21_,
         u5_mult_87_ab_3__22_, u5_mult_87_ab_3__23_, u5_mult_87_ab_3__24_,
         u5_mult_87_ab_3__25_, u5_mult_87_ab_3__26_, u5_mult_87_ab_3__27_,
         u5_mult_87_ab_3__28_, u5_mult_87_ab_3__29_, u5_mult_87_ab_3__30_,
         u5_mult_87_ab_3__31_, u5_mult_87_ab_3__32_, u5_mult_87_ab_3__33_,
         u5_mult_87_ab_3__34_, u5_mult_87_ab_3__35_, u5_mult_87_ab_3__36_,
         u5_mult_87_ab_3__37_, u5_mult_87_ab_3__38_, u5_mult_87_ab_3__39_,
         u5_mult_87_ab_3__40_, u5_mult_87_ab_3__41_, u5_mult_87_ab_3__42_,
         u5_mult_87_ab_3__43_, u5_mult_87_ab_3__44_, u5_mult_87_ab_3__45_,
         u5_mult_87_ab_3__46_, u5_mult_87_ab_3__47_, u5_mult_87_ab_3__48_,
         u5_mult_87_ab_3__49_, u5_mult_87_ab_3__50_, u5_mult_87_ab_3__51_,
         u5_mult_87_ab_3__52_, u5_mult_87_ab_4__0_, u5_mult_87_ab_4__1_,
         u5_mult_87_ab_4__2_, u5_mult_87_ab_4__3_, u5_mult_87_ab_4__4_,
         u5_mult_87_ab_4__5_, u5_mult_87_ab_4__6_, u5_mult_87_ab_4__7_,
         u5_mult_87_ab_4__8_, u5_mult_87_ab_4__9_, u5_mult_87_ab_4__10_,
         u5_mult_87_ab_4__11_, u5_mult_87_ab_4__12_, u5_mult_87_ab_4__13_,
         u5_mult_87_ab_4__14_, u5_mult_87_ab_4__15_, u5_mult_87_ab_4__16_,
         u5_mult_87_ab_4__17_, u5_mult_87_ab_4__18_, u5_mult_87_ab_4__19_,
         u5_mult_87_ab_4__20_, u5_mult_87_ab_4__21_, u5_mult_87_ab_4__22_,
         u5_mult_87_ab_4__23_, u5_mult_87_ab_4__24_, u5_mult_87_ab_4__25_,
         u5_mult_87_ab_4__26_, u5_mult_87_ab_4__27_, u5_mult_87_ab_4__28_,
         u5_mult_87_ab_4__29_, u5_mult_87_ab_4__30_, u5_mult_87_ab_4__31_,
         u5_mult_87_ab_4__32_, u5_mult_87_ab_4__33_, u5_mult_87_ab_4__34_,
         u5_mult_87_ab_4__35_, u5_mult_87_ab_4__36_, u5_mult_87_ab_4__37_,
         u5_mult_87_ab_4__38_, u5_mult_87_ab_4__39_, u5_mult_87_ab_4__40_,
         u5_mult_87_ab_4__41_, u5_mult_87_ab_4__42_, u5_mult_87_ab_4__43_,
         u5_mult_87_ab_4__44_, u5_mult_87_ab_4__45_, u5_mult_87_ab_4__46_,
         u5_mult_87_ab_4__47_, u5_mult_87_ab_4__48_, u5_mult_87_ab_4__49_,
         u5_mult_87_ab_4__50_, u5_mult_87_ab_4__51_, u5_mult_87_ab_4__52_,
         u5_mult_87_ab_5__0_, u5_mult_87_ab_5__1_, u5_mult_87_ab_5__2_,
         u5_mult_87_ab_5__3_, u5_mult_87_ab_5__4_, u5_mult_87_ab_5__5_,
         u5_mult_87_ab_5__6_, u5_mult_87_ab_5__7_, u5_mult_87_ab_5__8_,
         u5_mult_87_ab_5__9_, u5_mult_87_ab_5__10_, u5_mult_87_ab_5__11_,
         u5_mult_87_ab_5__12_, u5_mult_87_ab_5__13_, u5_mult_87_ab_5__14_,
         u5_mult_87_ab_5__15_, u5_mult_87_ab_5__16_, u5_mult_87_ab_5__17_,
         u5_mult_87_ab_5__18_, u5_mult_87_ab_5__19_, u5_mult_87_ab_5__20_,
         u5_mult_87_ab_5__21_, u5_mult_87_ab_5__22_, u5_mult_87_ab_5__23_,
         u5_mult_87_ab_5__24_, u5_mult_87_ab_5__25_, u5_mult_87_ab_5__26_,
         u5_mult_87_ab_5__27_, u5_mult_87_ab_5__28_, u5_mult_87_ab_5__29_,
         u5_mult_87_ab_5__30_, u5_mult_87_ab_5__31_, u5_mult_87_ab_5__32_,
         u5_mult_87_ab_5__33_, u5_mult_87_ab_5__34_, u5_mult_87_ab_5__35_,
         u5_mult_87_ab_5__36_, u5_mult_87_ab_5__37_, u5_mult_87_ab_5__38_,
         u5_mult_87_ab_5__39_, u5_mult_87_ab_5__40_, u5_mult_87_ab_5__41_,
         u5_mult_87_ab_5__42_, u5_mult_87_ab_5__43_, u5_mult_87_ab_5__44_,
         u5_mult_87_ab_5__45_, u5_mult_87_ab_5__46_, u5_mult_87_ab_5__47_,
         u5_mult_87_ab_5__48_, u5_mult_87_ab_5__49_, u5_mult_87_ab_5__50_,
         u5_mult_87_ab_5__51_, u5_mult_87_ab_5__52_, u5_mult_87_ab_6__0_,
         u5_mult_87_ab_6__1_, u5_mult_87_ab_6__2_, u5_mult_87_ab_6__3_,
         u5_mult_87_ab_6__4_, u5_mult_87_ab_6__5_, u5_mult_87_ab_6__6_,
         u5_mult_87_ab_6__7_, u5_mult_87_ab_6__8_, u5_mult_87_ab_6__9_,
         u5_mult_87_ab_6__10_, u5_mult_87_ab_6__11_, u5_mult_87_ab_6__12_,
         u5_mult_87_ab_6__13_, u5_mult_87_ab_6__14_, u5_mult_87_ab_6__15_,
         u5_mult_87_ab_6__16_, u5_mult_87_ab_6__17_, u5_mult_87_ab_6__18_,
         u5_mult_87_ab_6__19_, u5_mult_87_ab_6__20_, u5_mult_87_ab_6__21_,
         u5_mult_87_ab_6__22_, u5_mult_87_ab_6__23_, u5_mult_87_ab_6__24_,
         u5_mult_87_ab_6__25_, u5_mult_87_ab_6__26_, u5_mult_87_ab_6__27_,
         u5_mult_87_ab_6__28_, u5_mult_87_ab_6__29_, u5_mult_87_ab_6__30_,
         u5_mult_87_ab_6__31_, u5_mult_87_ab_6__32_, u5_mult_87_ab_6__33_,
         u5_mult_87_ab_6__34_, u5_mult_87_ab_6__35_, u5_mult_87_ab_6__36_,
         u5_mult_87_ab_6__37_, u5_mult_87_ab_6__38_, u5_mult_87_ab_6__39_,
         u5_mult_87_ab_6__40_, u5_mult_87_ab_6__41_, u5_mult_87_ab_6__42_,
         u5_mult_87_ab_6__43_, u5_mult_87_ab_6__44_, u5_mult_87_ab_6__45_,
         u5_mult_87_ab_6__46_, u5_mult_87_ab_6__47_, u5_mult_87_ab_6__48_,
         u5_mult_87_ab_6__49_, u5_mult_87_ab_6__50_, u5_mult_87_ab_6__51_,
         u5_mult_87_ab_6__52_, u5_mult_87_ab_7__0_, u5_mult_87_ab_7__1_,
         u5_mult_87_ab_7__2_, u5_mult_87_ab_7__3_, u5_mult_87_ab_7__4_,
         u5_mult_87_ab_7__5_, u5_mult_87_ab_7__6_, u5_mult_87_ab_7__7_,
         u5_mult_87_ab_7__8_, u5_mult_87_ab_7__9_, u5_mult_87_ab_7__10_,
         u5_mult_87_ab_7__11_, u5_mult_87_ab_7__12_, u5_mult_87_ab_7__13_,
         u5_mult_87_ab_7__14_, u5_mult_87_ab_7__15_, u5_mult_87_ab_7__16_,
         u5_mult_87_ab_7__17_, u5_mult_87_ab_7__18_, u5_mult_87_ab_7__19_,
         u5_mult_87_ab_7__20_, u5_mult_87_ab_7__21_, u5_mult_87_ab_7__22_,
         u5_mult_87_ab_7__23_, u5_mult_87_ab_7__24_, u5_mult_87_ab_7__25_,
         u5_mult_87_ab_7__26_, u5_mult_87_ab_7__27_, u5_mult_87_ab_7__28_,
         u5_mult_87_ab_7__29_, u5_mult_87_ab_7__30_, u5_mult_87_ab_7__31_,
         u5_mult_87_ab_7__32_, u5_mult_87_ab_7__33_, u5_mult_87_ab_7__34_,
         u5_mult_87_ab_7__35_, u5_mult_87_ab_7__36_, u5_mult_87_ab_7__37_,
         u5_mult_87_ab_7__38_, u5_mult_87_ab_7__39_, u5_mult_87_ab_7__40_,
         u5_mult_87_ab_7__41_, u5_mult_87_ab_7__42_, u5_mult_87_ab_7__43_,
         u5_mult_87_ab_7__44_, u5_mult_87_ab_7__45_, u5_mult_87_ab_7__46_,
         u5_mult_87_ab_7__47_, u5_mult_87_ab_7__48_, u5_mult_87_ab_7__49_,
         u5_mult_87_ab_7__50_, u5_mult_87_ab_7__51_, u5_mult_87_ab_7__52_,
         u5_mult_87_ab_8__0_, u5_mult_87_ab_8__1_, u5_mult_87_ab_8__2_,
         u5_mult_87_ab_8__3_, u5_mult_87_ab_8__4_, u5_mult_87_ab_8__5_,
         u5_mult_87_ab_8__6_, u5_mult_87_ab_8__7_, u5_mult_87_ab_8__8_,
         u5_mult_87_ab_8__9_, u5_mult_87_ab_8__10_, u5_mult_87_ab_8__11_,
         u5_mult_87_ab_8__12_, u5_mult_87_ab_8__13_, u5_mult_87_ab_8__14_,
         u5_mult_87_ab_8__15_, u5_mult_87_ab_8__16_, u5_mult_87_ab_8__17_,
         u5_mult_87_ab_8__18_, u5_mult_87_ab_8__19_, u5_mult_87_ab_8__20_,
         u5_mult_87_ab_8__21_, u5_mult_87_ab_8__22_, u5_mult_87_ab_8__23_,
         u5_mult_87_ab_8__24_, u5_mult_87_ab_8__25_, u5_mult_87_ab_8__26_,
         u5_mult_87_ab_8__27_, u5_mult_87_ab_8__28_, u5_mult_87_ab_8__29_,
         u5_mult_87_ab_8__30_, u5_mult_87_ab_8__31_, u5_mult_87_ab_8__32_,
         u5_mult_87_ab_8__33_, u5_mult_87_ab_8__34_, u5_mult_87_ab_8__35_,
         u5_mult_87_ab_8__36_, u5_mult_87_ab_8__37_, u5_mult_87_ab_8__38_,
         u5_mult_87_ab_8__39_, u5_mult_87_ab_8__40_, u5_mult_87_ab_8__41_,
         u5_mult_87_ab_8__42_, u5_mult_87_ab_8__43_, u5_mult_87_ab_8__44_,
         u5_mult_87_ab_8__45_, u5_mult_87_ab_8__46_, u5_mult_87_ab_8__47_,
         u5_mult_87_ab_8__48_, u5_mult_87_ab_8__49_, u5_mult_87_ab_8__50_,
         u5_mult_87_ab_8__51_, u5_mult_87_ab_8__52_, u5_mult_87_ab_9__0_,
         u5_mult_87_ab_9__1_, u5_mult_87_ab_9__2_, u5_mult_87_ab_9__3_,
         u5_mult_87_ab_9__4_, u5_mult_87_ab_9__5_, u5_mult_87_ab_9__6_,
         u5_mult_87_ab_9__7_, u5_mult_87_ab_9__8_, u5_mult_87_ab_9__9_,
         u5_mult_87_ab_9__10_, u5_mult_87_ab_9__11_, u5_mult_87_ab_9__12_,
         u5_mult_87_ab_9__13_, u5_mult_87_ab_9__14_, u5_mult_87_ab_9__15_,
         u5_mult_87_ab_9__16_, u5_mult_87_ab_9__17_, u5_mult_87_ab_9__18_,
         u5_mult_87_ab_9__19_, u5_mult_87_ab_9__20_, u5_mult_87_ab_9__21_,
         u5_mult_87_ab_9__22_, u5_mult_87_ab_9__23_, u5_mult_87_ab_9__24_,
         u5_mult_87_ab_9__25_, u5_mult_87_ab_9__26_, u5_mult_87_ab_9__27_,
         u5_mult_87_ab_9__28_, u5_mult_87_ab_9__29_, u5_mult_87_ab_9__30_,
         u5_mult_87_ab_9__31_, u5_mult_87_ab_9__32_, u5_mult_87_ab_9__33_,
         u5_mult_87_ab_9__34_, u5_mult_87_ab_9__35_, u5_mult_87_ab_9__36_,
         u5_mult_87_ab_9__37_, u5_mult_87_ab_9__38_, u5_mult_87_ab_9__39_,
         u5_mult_87_ab_9__40_, u5_mult_87_ab_9__41_, u5_mult_87_ab_9__42_,
         u5_mult_87_ab_9__43_, u5_mult_87_ab_9__44_, u5_mult_87_ab_9__45_,
         u5_mult_87_ab_9__46_, u5_mult_87_ab_9__47_, u5_mult_87_ab_9__48_,
         u5_mult_87_ab_9__49_, u5_mult_87_ab_9__50_, u5_mult_87_ab_9__51_,
         u5_mult_87_ab_9__52_, u5_mult_87_ab_10__0_, u5_mult_87_ab_10__1_,
         u5_mult_87_ab_10__2_, u5_mult_87_ab_10__3_, u5_mult_87_ab_10__4_,
         u5_mult_87_ab_10__5_, u5_mult_87_ab_10__6_, u5_mult_87_ab_10__7_,
         u5_mult_87_ab_10__8_, u5_mult_87_ab_10__9_, u5_mult_87_ab_10__10_,
         u5_mult_87_ab_10__11_, u5_mult_87_ab_10__12_, u5_mult_87_ab_10__13_,
         u5_mult_87_ab_10__14_, u5_mult_87_ab_10__15_, u5_mult_87_ab_10__16_,
         u5_mult_87_ab_10__17_, u5_mult_87_ab_10__18_, u5_mult_87_ab_10__19_,
         u5_mult_87_ab_10__20_, u5_mult_87_ab_10__21_, u5_mult_87_ab_10__22_,
         u5_mult_87_ab_10__23_, u5_mult_87_ab_10__24_, u5_mult_87_ab_10__25_,
         u5_mult_87_ab_10__26_, u5_mult_87_ab_10__27_, u5_mult_87_ab_10__28_,
         u5_mult_87_ab_10__29_, u5_mult_87_ab_10__30_, u5_mult_87_ab_10__31_,
         u5_mult_87_ab_10__32_, u5_mult_87_ab_10__33_, u5_mult_87_ab_10__34_,
         u5_mult_87_ab_10__35_, u5_mult_87_ab_10__36_, u5_mult_87_ab_10__37_,
         u5_mult_87_ab_10__38_, u5_mult_87_ab_10__39_, u5_mult_87_ab_10__40_,
         u5_mult_87_ab_10__41_, u5_mult_87_ab_10__42_, u5_mult_87_ab_10__43_,
         u5_mult_87_ab_10__44_, u5_mult_87_ab_10__45_, u5_mult_87_ab_10__46_,
         u5_mult_87_ab_10__47_, u5_mult_87_ab_10__48_, u5_mult_87_ab_10__49_,
         u5_mult_87_ab_10__50_, u5_mult_87_ab_10__51_, u5_mult_87_ab_10__52_,
         u5_mult_87_ab_11__0_, u5_mult_87_ab_11__1_, u5_mult_87_ab_11__2_,
         u5_mult_87_ab_11__3_, u5_mult_87_ab_11__4_, u5_mult_87_ab_11__5_,
         u5_mult_87_ab_11__6_, u5_mult_87_ab_11__7_, u5_mult_87_ab_11__8_,
         u5_mult_87_ab_11__9_, u5_mult_87_ab_11__10_, u5_mult_87_ab_11__11_,
         u5_mult_87_ab_11__12_, u5_mult_87_ab_11__13_, u5_mult_87_ab_11__14_,
         u5_mult_87_ab_11__15_, u5_mult_87_ab_11__16_, u5_mult_87_ab_11__17_,
         u5_mult_87_ab_11__18_, u5_mult_87_ab_11__19_, u5_mult_87_ab_11__20_,
         u5_mult_87_ab_11__21_, u5_mult_87_ab_11__22_, u5_mult_87_ab_11__23_,
         u5_mult_87_ab_11__24_, u5_mult_87_ab_11__25_, u5_mult_87_ab_11__26_,
         u5_mult_87_ab_11__27_, u5_mult_87_ab_11__28_, u5_mult_87_ab_11__29_,
         u5_mult_87_ab_11__30_, u5_mult_87_ab_11__31_, u5_mult_87_ab_11__32_,
         u5_mult_87_ab_11__33_, u5_mult_87_ab_11__34_, u5_mult_87_ab_11__35_,
         u5_mult_87_ab_11__36_, u5_mult_87_ab_11__37_, u5_mult_87_ab_11__38_,
         u5_mult_87_ab_11__39_, u5_mult_87_ab_11__40_, u5_mult_87_ab_11__41_,
         u5_mult_87_ab_11__42_, u5_mult_87_ab_11__43_, u5_mult_87_ab_11__44_,
         u5_mult_87_ab_11__45_, u5_mult_87_ab_11__46_, u5_mult_87_ab_11__47_,
         u5_mult_87_ab_11__48_, u5_mult_87_ab_11__49_, u5_mult_87_ab_11__50_,
         u5_mult_87_ab_11__51_, u5_mult_87_ab_11__52_, u5_mult_87_ab_12__0_,
         u5_mult_87_ab_12__1_, u5_mult_87_ab_12__2_, u5_mult_87_ab_12__3_,
         u5_mult_87_ab_12__4_, u5_mult_87_ab_12__5_, u5_mult_87_ab_12__6_,
         u5_mult_87_ab_12__7_, u5_mult_87_ab_12__8_, u5_mult_87_ab_12__9_,
         u5_mult_87_ab_12__10_, u5_mult_87_ab_12__11_, u5_mult_87_ab_12__12_,
         u5_mult_87_ab_12__13_, u5_mult_87_ab_12__14_, u5_mult_87_ab_12__15_,
         u5_mult_87_ab_12__16_, u5_mult_87_ab_12__17_, u5_mult_87_ab_12__18_,
         u5_mult_87_ab_12__19_, u5_mult_87_ab_12__20_, u5_mult_87_ab_12__21_,
         u5_mult_87_ab_12__22_, u5_mult_87_ab_12__23_, u5_mult_87_ab_12__24_,
         u5_mult_87_ab_12__25_, u5_mult_87_ab_12__26_, u5_mult_87_ab_12__27_,
         u5_mult_87_ab_12__28_, u5_mult_87_ab_12__29_, u5_mult_87_ab_12__30_,
         u5_mult_87_ab_12__31_, u5_mult_87_ab_12__32_, u5_mult_87_ab_12__33_,
         u5_mult_87_ab_12__34_, u5_mult_87_ab_12__35_, u5_mult_87_ab_12__36_,
         u5_mult_87_ab_12__37_, u5_mult_87_ab_12__38_, u5_mult_87_ab_12__39_,
         u5_mult_87_ab_12__40_, u5_mult_87_ab_12__41_, u5_mult_87_ab_12__42_,
         u5_mult_87_ab_12__43_, u5_mult_87_ab_12__44_, u5_mult_87_ab_12__45_,
         u5_mult_87_ab_12__46_, u5_mult_87_ab_12__47_, u5_mult_87_ab_12__48_,
         u5_mult_87_ab_12__49_, u5_mult_87_ab_12__50_, u5_mult_87_ab_12__51_,
         u5_mult_87_ab_12__52_, u5_mult_87_ab_13__0_, u5_mult_87_ab_13__1_,
         u5_mult_87_ab_13__2_, u5_mult_87_ab_13__3_, u5_mult_87_ab_13__4_,
         u5_mult_87_ab_13__5_, u5_mult_87_ab_13__6_, u5_mult_87_ab_13__7_,
         u5_mult_87_ab_13__8_, u5_mult_87_ab_13__9_, u5_mult_87_ab_13__10_,
         u5_mult_87_ab_13__11_, u5_mult_87_ab_13__12_, u5_mult_87_ab_13__13_,
         u5_mult_87_ab_13__14_, u5_mult_87_ab_13__15_, u5_mult_87_ab_13__16_,
         u5_mult_87_ab_13__17_, u5_mult_87_ab_13__18_, u5_mult_87_ab_13__19_,
         u5_mult_87_ab_13__20_, u5_mult_87_ab_13__21_, u5_mult_87_ab_13__22_,
         u5_mult_87_ab_13__23_, u5_mult_87_ab_13__24_, u5_mult_87_ab_13__25_,
         u5_mult_87_ab_13__26_, u5_mult_87_ab_13__27_, u5_mult_87_ab_13__28_,
         u5_mult_87_ab_13__29_, u5_mult_87_ab_13__30_, u5_mult_87_ab_13__31_,
         u5_mult_87_ab_13__32_, u5_mult_87_ab_13__33_, u5_mult_87_ab_13__34_,
         u5_mult_87_ab_13__35_, u5_mult_87_ab_13__36_, u5_mult_87_ab_13__37_,
         u5_mult_87_ab_13__38_, u5_mult_87_ab_13__39_, u5_mult_87_ab_13__40_,
         u5_mult_87_ab_13__41_, u5_mult_87_ab_13__42_, u5_mult_87_ab_13__43_,
         u5_mult_87_ab_13__44_, u5_mult_87_ab_13__45_, u5_mult_87_ab_13__46_,
         u5_mult_87_ab_13__47_, u5_mult_87_ab_13__48_, u5_mult_87_ab_13__49_,
         u5_mult_87_ab_13__50_, u5_mult_87_ab_13__51_, u5_mult_87_ab_13__52_,
         u5_mult_87_ab_14__0_, u5_mult_87_ab_14__1_, u5_mult_87_ab_14__2_,
         u5_mult_87_ab_14__3_, u5_mult_87_ab_14__4_, u5_mult_87_ab_14__5_,
         u5_mult_87_ab_14__6_, u5_mult_87_ab_14__7_, u5_mult_87_ab_14__8_,
         u5_mult_87_ab_14__9_, u5_mult_87_ab_14__10_, u5_mult_87_ab_14__11_,
         u5_mult_87_ab_14__12_, u5_mult_87_ab_14__13_, u5_mult_87_ab_14__14_,
         u5_mult_87_ab_14__15_, u5_mult_87_ab_14__16_, u5_mult_87_ab_14__17_,
         u5_mult_87_ab_14__18_, u5_mult_87_ab_14__19_, u5_mult_87_ab_14__20_,
         u5_mult_87_ab_14__21_, u5_mult_87_ab_14__22_, u5_mult_87_ab_14__23_,
         u5_mult_87_ab_14__24_, u5_mult_87_ab_14__25_, u5_mult_87_ab_14__26_,
         u5_mult_87_ab_14__27_, u5_mult_87_ab_14__28_, u5_mult_87_ab_14__29_,
         u5_mult_87_ab_14__30_, u5_mult_87_ab_14__31_, u5_mult_87_ab_14__32_,
         u5_mult_87_ab_14__33_, u5_mult_87_ab_14__34_, u5_mult_87_ab_14__35_,
         u5_mult_87_ab_14__36_, u5_mult_87_ab_14__37_, u5_mult_87_ab_14__38_,
         u5_mult_87_ab_14__39_, u5_mult_87_ab_14__40_, u5_mult_87_ab_14__41_,
         u5_mult_87_ab_14__42_, u5_mult_87_ab_14__43_, u5_mult_87_ab_14__44_,
         u5_mult_87_ab_14__45_, u5_mult_87_ab_14__46_, u5_mult_87_ab_14__47_,
         u5_mult_87_ab_14__48_, u5_mult_87_ab_14__49_, u5_mult_87_ab_14__50_,
         u5_mult_87_ab_14__51_, u5_mult_87_ab_14__52_, u5_mult_87_ab_15__0_,
         u5_mult_87_ab_15__1_, u5_mult_87_ab_15__2_, u5_mult_87_ab_15__3_,
         u5_mult_87_ab_15__4_, u5_mult_87_ab_15__5_, u5_mult_87_ab_15__6_,
         u5_mult_87_ab_15__7_, u5_mult_87_ab_15__8_, u5_mult_87_ab_15__9_,
         u5_mult_87_ab_15__10_, u5_mult_87_ab_15__11_, u5_mult_87_ab_15__12_,
         u5_mult_87_ab_15__13_, u5_mult_87_ab_15__14_, u5_mult_87_ab_15__15_,
         u5_mult_87_ab_15__16_, u5_mult_87_ab_15__17_, u5_mult_87_ab_15__18_,
         u5_mult_87_ab_15__19_, u5_mult_87_ab_15__20_, u5_mult_87_ab_15__21_,
         u5_mult_87_ab_15__22_, u5_mult_87_ab_15__23_, u5_mult_87_ab_15__24_,
         u5_mult_87_ab_15__25_, u5_mult_87_ab_15__26_, u5_mult_87_ab_15__27_,
         u5_mult_87_ab_15__28_, u5_mult_87_ab_15__29_, u5_mult_87_ab_15__30_,
         u5_mult_87_ab_15__31_, u5_mult_87_ab_15__32_, u5_mult_87_ab_15__33_,
         u5_mult_87_ab_15__34_, u5_mult_87_ab_15__35_, u5_mult_87_ab_15__36_,
         u5_mult_87_ab_15__37_, u5_mult_87_ab_15__38_, u5_mult_87_ab_15__39_,
         u5_mult_87_ab_15__40_, u5_mult_87_ab_15__41_, u5_mult_87_ab_15__42_,
         u5_mult_87_ab_15__43_, u5_mult_87_ab_15__44_, u5_mult_87_ab_15__45_,
         u5_mult_87_ab_15__46_, u5_mult_87_ab_15__47_, u5_mult_87_ab_15__48_,
         u5_mult_87_ab_15__49_, u5_mult_87_ab_15__50_, u5_mult_87_ab_15__51_,
         u5_mult_87_ab_15__52_, u5_mult_87_ab_16__0_, u5_mult_87_ab_16__1_,
         u5_mult_87_ab_16__2_, u5_mult_87_ab_16__3_, u5_mult_87_ab_16__4_,
         u5_mult_87_ab_16__5_, u5_mult_87_ab_16__6_, u5_mult_87_ab_16__7_,
         u5_mult_87_ab_16__8_, u5_mult_87_ab_16__9_, u5_mult_87_ab_16__10_,
         u5_mult_87_ab_16__11_, u5_mult_87_ab_16__12_, u5_mult_87_ab_16__13_,
         u5_mult_87_ab_16__14_, u5_mult_87_ab_16__15_, u5_mult_87_ab_16__16_,
         u5_mult_87_ab_16__17_, u5_mult_87_ab_16__18_, u5_mult_87_ab_16__19_,
         u5_mult_87_ab_16__20_, u5_mult_87_ab_16__21_, u5_mult_87_ab_16__22_,
         u5_mult_87_ab_16__23_, u5_mult_87_ab_16__24_, u5_mult_87_ab_16__25_,
         u5_mult_87_ab_16__26_, u5_mult_87_ab_16__27_, u5_mult_87_ab_16__28_,
         u5_mult_87_ab_16__29_, u5_mult_87_ab_16__30_, u5_mult_87_ab_16__31_,
         u5_mult_87_ab_16__32_, u5_mult_87_ab_16__33_, u5_mult_87_ab_16__34_,
         u5_mult_87_ab_16__35_, u5_mult_87_ab_16__36_, u5_mult_87_ab_16__37_,
         u5_mult_87_ab_16__38_, u5_mult_87_ab_16__39_, u5_mult_87_ab_16__40_,
         u5_mult_87_ab_16__41_, u5_mult_87_ab_16__42_, u5_mult_87_ab_16__43_,
         u5_mult_87_ab_16__44_, u5_mult_87_ab_16__45_, u5_mult_87_ab_16__46_,
         u5_mult_87_ab_16__47_, u5_mult_87_ab_16__48_, u5_mult_87_ab_16__49_,
         u5_mult_87_ab_16__50_, u5_mult_87_ab_16__51_, u5_mult_87_ab_16__52_,
         u5_mult_87_ab_17__0_, u5_mult_87_ab_17__1_, u5_mult_87_ab_17__2_,
         u5_mult_87_ab_17__3_, u5_mult_87_ab_17__4_, u5_mult_87_ab_17__5_,
         u5_mult_87_ab_17__6_, u5_mult_87_ab_17__7_, u5_mult_87_ab_17__8_,
         u5_mult_87_ab_17__9_, u5_mult_87_ab_17__10_, u5_mult_87_ab_17__11_,
         u5_mult_87_ab_17__12_, u5_mult_87_ab_17__13_, u5_mult_87_ab_17__14_,
         u5_mult_87_ab_17__15_, u5_mult_87_ab_17__16_, u5_mult_87_ab_17__17_,
         u5_mult_87_ab_17__18_, u5_mult_87_ab_17__19_, u5_mult_87_ab_17__20_,
         u5_mult_87_ab_17__21_, u5_mult_87_ab_17__22_, u5_mult_87_ab_17__23_,
         u5_mult_87_ab_17__24_, u5_mult_87_ab_17__25_, u5_mult_87_ab_17__26_,
         u5_mult_87_ab_17__27_, u5_mult_87_ab_17__28_, u5_mult_87_ab_17__29_,
         u5_mult_87_ab_17__30_, u5_mult_87_ab_17__31_, u5_mult_87_ab_17__32_,
         u5_mult_87_ab_17__33_, u5_mult_87_ab_17__34_, u5_mult_87_ab_17__35_,
         u5_mult_87_ab_17__36_, u5_mult_87_ab_17__37_, u5_mult_87_ab_17__38_,
         u5_mult_87_ab_17__39_, u5_mult_87_ab_17__40_, u5_mult_87_ab_17__41_,
         u5_mult_87_ab_17__42_, u5_mult_87_ab_17__43_, u5_mult_87_ab_17__44_,
         u5_mult_87_ab_17__45_, u5_mult_87_ab_17__46_, u5_mult_87_ab_17__47_,
         u5_mult_87_ab_17__48_, u5_mult_87_ab_17__49_, u5_mult_87_ab_17__50_,
         u5_mult_87_ab_17__51_, u5_mult_87_ab_17__52_, u5_mult_87_ab_18__0_,
         u5_mult_87_ab_18__1_, u5_mult_87_ab_18__2_, u5_mult_87_ab_18__3_,
         u5_mult_87_ab_18__4_, u5_mult_87_ab_18__5_, u5_mult_87_ab_18__6_,
         u5_mult_87_ab_18__7_, u5_mult_87_ab_18__8_, u5_mult_87_ab_18__9_,
         u5_mult_87_ab_18__10_, u5_mult_87_ab_18__11_, u5_mult_87_ab_18__12_,
         u5_mult_87_ab_18__13_, u5_mult_87_ab_18__14_, u5_mult_87_ab_18__15_,
         u5_mult_87_ab_18__16_, u5_mult_87_ab_18__17_, u5_mult_87_ab_18__18_,
         u5_mult_87_ab_18__19_, u5_mult_87_ab_18__20_, u5_mult_87_ab_18__21_,
         u5_mult_87_ab_18__22_, u5_mult_87_ab_18__23_, u5_mult_87_ab_18__24_,
         u5_mult_87_ab_18__25_, u5_mult_87_ab_18__26_, u5_mult_87_ab_18__27_,
         u5_mult_87_ab_18__28_, u5_mult_87_ab_18__29_, u5_mult_87_ab_18__30_,
         u5_mult_87_ab_18__31_, u5_mult_87_ab_18__32_, u5_mult_87_ab_18__33_,
         u5_mult_87_ab_18__34_, u5_mult_87_ab_18__35_, u5_mult_87_ab_18__36_,
         u5_mult_87_ab_18__37_, u5_mult_87_ab_18__38_, u5_mult_87_ab_18__39_,
         u5_mult_87_ab_18__40_, u5_mult_87_ab_18__41_, u5_mult_87_ab_18__42_,
         u5_mult_87_ab_18__43_, u5_mult_87_ab_18__44_, u5_mult_87_ab_18__45_,
         u5_mult_87_ab_18__46_, u5_mult_87_ab_18__47_, u5_mult_87_ab_18__48_,
         u5_mult_87_ab_18__49_, u5_mult_87_ab_18__50_, u5_mult_87_ab_18__51_,
         u5_mult_87_ab_18__52_, u5_mult_87_ab_19__0_, u5_mult_87_ab_19__1_,
         u5_mult_87_ab_19__2_, u5_mult_87_ab_19__3_, u5_mult_87_ab_19__4_,
         u5_mult_87_ab_19__5_, u5_mult_87_ab_19__6_, u5_mult_87_ab_19__7_,
         u5_mult_87_ab_19__8_, u5_mult_87_ab_19__9_, u5_mult_87_ab_19__10_,
         u5_mult_87_ab_19__11_, u5_mult_87_ab_19__12_, u5_mult_87_ab_19__13_,
         u5_mult_87_ab_19__14_, u5_mult_87_ab_19__15_, u5_mult_87_ab_19__16_,
         u5_mult_87_ab_19__17_, u5_mult_87_ab_19__18_, u5_mult_87_ab_19__19_,
         u5_mult_87_ab_19__20_, u5_mult_87_ab_19__21_, u5_mult_87_ab_19__22_,
         u5_mult_87_ab_19__23_, u5_mult_87_ab_19__24_, u5_mult_87_ab_19__25_,
         u5_mult_87_ab_19__26_, u5_mult_87_ab_19__27_, u5_mult_87_ab_19__28_,
         u5_mult_87_ab_19__29_, u5_mult_87_ab_19__30_, u5_mult_87_ab_19__31_,
         u5_mult_87_ab_19__32_, u5_mult_87_ab_19__33_, u5_mult_87_ab_19__34_,
         u5_mult_87_ab_19__35_, u5_mult_87_ab_19__36_, u5_mult_87_ab_19__37_,
         u5_mult_87_ab_19__38_, u5_mult_87_ab_19__39_, u5_mult_87_ab_19__40_,
         u5_mult_87_ab_19__41_, u5_mult_87_ab_19__42_, u5_mult_87_ab_19__43_,
         u5_mult_87_ab_19__44_, u5_mult_87_ab_19__45_, u5_mult_87_ab_19__46_,
         u5_mult_87_ab_19__47_, u5_mult_87_ab_19__48_, u5_mult_87_ab_19__49_,
         u5_mult_87_ab_19__50_, u5_mult_87_ab_19__51_, u5_mult_87_ab_19__52_,
         u5_mult_87_ab_20__0_, u5_mult_87_ab_20__1_, u5_mult_87_ab_20__2_,
         u5_mult_87_ab_20__3_, u5_mult_87_ab_20__4_, u5_mult_87_ab_20__5_,
         u5_mult_87_ab_20__6_, u5_mult_87_ab_20__7_, u5_mult_87_ab_20__8_,
         u5_mult_87_ab_20__9_, u5_mult_87_ab_20__10_, u5_mult_87_ab_20__11_,
         u5_mult_87_ab_20__12_, u5_mult_87_ab_20__13_, u5_mult_87_ab_20__14_,
         u5_mult_87_ab_20__15_, u5_mult_87_ab_20__16_, u5_mult_87_ab_20__17_,
         u5_mult_87_ab_20__18_, u5_mult_87_ab_20__19_, u5_mult_87_ab_20__20_,
         u5_mult_87_ab_20__21_, u5_mult_87_ab_20__22_, u5_mult_87_ab_20__23_,
         u5_mult_87_ab_20__24_, u5_mult_87_ab_20__25_, u5_mult_87_ab_20__26_,
         u5_mult_87_ab_20__27_, u5_mult_87_ab_20__28_, u5_mult_87_ab_20__29_,
         u5_mult_87_ab_20__30_, u5_mult_87_ab_20__31_, u5_mult_87_ab_20__32_,
         u5_mult_87_ab_20__33_, u5_mult_87_ab_20__34_, u5_mult_87_ab_20__35_,
         u5_mult_87_ab_20__36_, u5_mult_87_ab_20__37_, u5_mult_87_ab_20__38_,
         u5_mult_87_ab_20__39_, u5_mult_87_ab_20__40_, u5_mult_87_ab_20__41_,
         u5_mult_87_ab_20__42_, u5_mult_87_ab_20__43_, u5_mult_87_ab_20__44_,
         u5_mult_87_ab_20__45_, u5_mult_87_ab_20__46_, u5_mult_87_ab_20__47_,
         u5_mult_87_ab_20__48_, u5_mult_87_ab_20__49_, u5_mult_87_ab_20__50_,
         u5_mult_87_ab_20__51_, u5_mult_87_ab_20__52_, u5_mult_87_ab_21__0_,
         u5_mult_87_ab_21__1_, u5_mult_87_ab_21__2_, u5_mult_87_ab_21__3_,
         u5_mult_87_ab_21__4_, u5_mult_87_ab_21__5_, u5_mult_87_ab_21__6_,
         u5_mult_87_ab_21__7_, u5_mult_87_ab_21__8_, u5_mult_87_ab_21__9_,
         u5_mult_87_ab_21__10_, u5_mult_87_ab_21__11_, u5_mult_87_ab_21__12_,
         u5_mult_87_ab_21__13_, u5_mult_87_ab_21__14_, u5_mult_87_ab_21__15_,
         u5_mult_87_ab_21__16_, u5_mult_87_ab_21__17_, u5_mult_87_ab_21__18_,
         u5_mult_87_ab_21__19_, u5_mult_87_ab_21__20_, u5_mult_87_ab_21__21_,
         u5_mult_87_ab_21__22_, u5_mult_87_ab_21__23_, u5_mult_87_ab_21__24_,
         u5_mult_87_ab_21__25_, u5_mult_87_ab_21__26_, u5_mult_87_ab_21__27_,
         u5_mult_87_ab_21__28_, u5_mult_87_ab_21__29_, u5_mult_87_ab_21__30_,
         u5_mult_87_ab_21__31_, u5_mult_87_ab_21__32_, u5_mult_87_ab_21__33_,
         u5_mult_87_ab_21__34_, u5_mult_87_ab_21__35_, u5_mult_87_ab_21__36_,
         u5_mult_87_ab_21__37_, u5_mult_87_ab_21__38_, u5_mult_87_ab_21__39_,
         u5_mult_87_ab_21__40_, u5_mult_87_ab_21__41_, u5_mult_87_ab_21__42_,
         u5_mult_87_ab_21__43_, u5_mult_87_ab_21__44_, u5_mult_87_ab_21__45_,
         u5_mult_87_ab_21__46_, u5_mult_87_ab_21__47_, u5_mult_87_ab_21__48_,
         u5_mult_87_ab_21__49_, u5_mult_87_ab_21__50_, u5_mult_87_ab_21__51_,
         u5_mult_87_ab_21__52_, u5_mult_87_ab_22__0_, u5_mult_87_ab_22__1_,
         u5_mult_87_ab_22__2_, u5_mult_87_ab_22__3_, u5_mult_87_ab_22__4_,
         u5_mult_87_ab_22__5_, u5_mult_87_ab_22__6_, u5_mult_87_ab_22__7_,
         u5_mult_87_ab_22__8_, u5_mult_87_ab_22__9_, u5_mult_87_ab_22__10_,
         u5_mult_87_ab_22__11_, u5_mult_87_ab_22__12_, u5_mult_87_ab_22__13_,
         u5_mult_87_ab_22__14_, u5_mult_87_ab_22__15_, u5_mult_87_ab_22__16_,
         u5_mult_87_ab_22__17_, u5_mult_87_ab_22__18_, u5_mult_87_ab_22__19_,
         u5_mult_87_ab_22__20_, u5_mult_87_ab_22__21_, u5_mult_87_ab_22__22_,
         u5_mult_87_ab_22__23_, u5_mult_87_ab_22__24_, u5_mult_87_ab_22__25_,
         u5_mult_87_ab_22__26_, u5_mult_87_ab_22__27_, u5_mult_87_ab_22__28_,
         u5_mult_87_ab_22__29_, u5_mult_87_ab_22__30_, u5_mult_87_ab_22__31_,
         u5_mult_87_ab_22__32_, u5_mult_87_ab_22__33_, u5_mult_87_ab_22__34_,
         u5_mult_87_ab_22__35_, u5_mult_87_ab_22__36_, u5_mult_87_ab_22__37_,
         u5_mult_87_ab_22__38_, u5_mult_87_ab_22__39_, u5_mult_87_ab_22__40_,
         u5_mult_87_ab_22__41_, u5_mult_87_ab_22__42_, u5_mult_87_ab_22__43_,
         u5_mult_87_ab_22__44_, u5_mult_87_ab_22__45_, u5_mult_87_ab_22__46_,
         u5_mult_87_ab_22__47_, u5_mult_87_ab_22__48_, u5_mult_87_ab_22__49_,
         u5_mult_87_ab_22__50_, u5_mult_87_ab_22__51_, u5_mult_87_ab_22__52_,
         u5_mult_87_ab_23__0_, u5_mult_87_ab_23__1_, u5_mult_87_ab_23__2_,
         u5_mult_87_ab_23__3_, u5_mult_87_ab_23__4_, u5_mult_87_ab_23__5_,
         u5_mult_87_ab_23__6_, u5_mult_87_ab_23__7_, u5_mult_87_ab_23__8_,
         u5_mult_87_ab_23__9_, u5_mult_87_ab_23__10_, u5_mult_87_ab_23__11_,
         u5_mult_87_ab_23__12_, u5_mult_87_ab_23__13_, u5_mult_87_ab_23__14_,
         u5_mult_87_ab_23__15_, u5_mult_87_ab_23__16_, u5_mult_87_ab_23__17_,
         u5_mult_87_ab_23__18_, u5_mult_87_ab_23__19_, u5_mult_87_ab_23__20_,
         u5_mult_87_ab_23__21_, u5_mult_87_ab_23__22_, u5_mult_87_ab_23__23_,
         u5_mult_87_ab_23__24_, u5_mult_87_ab_23__25_, u5_mult_87_ab_23__26_,
         u5_mult_87_ab_23__27_, u5_mult_87_ab_23__28_, u5_mult_87_ab_23__29_,
         u5_mult_87_ab_23__30_, u5_mult_87_ab_23__31_, u5_mult_87_ab_23__32_,
         u5_mult_87_ab_23__33_, u5_mult_87_ab_23__34_, u5_mult_87_ab_23__35_,
         u5_mult_87_ab_23__36_, u5_mult_87_ab_23__37_, u5_mult_87_ab_23__38_,
         u5_mult_87_ab_23__39_, u5_mult_87_ab_23__40_, u5_mult_87_ab_23__41_,
         u5_mult_87_ab_23__42_, u5_mult_87_ab_23__43_, u5_mult_87_ab_23__44_,
         u5_mult_87_ab_23__45_, u5_mult_87_ab_23__46_, u5_mult_87_ab_23__47_,
         u5_mult_87_ab_23__48_, u5_mult_87_ab_23__49_, u5_mult_87_ab_23__50_,
         u5_mult_87_ab_23__51_, u5_mult_87_ab_23__52_, u5_mult_87_ab_24__0_,
         u5_mult_87_ab_24__1_, u5_mult_87_ab_24__2_, u5_mult_87_ab_24__3_,
         u5_mult_87_ab_24__4_, u5_mult_87_ab_24__5_, u5_mult_87_ab_24__6_,
         u5_mult_87_ab_24__7_, u5_mult_87_ab_24__8_, u5_mult_87_ab_24__9_,
         u5_mult_87_ab_24__10_, u5_mult_87_ab_24__11_, u5_mult_87_ab_24__12_,
         u5_mult_87_ab_24__13_, u5_mult_87_ab_24__14_, u5_mult_87_ab_24__15_,
         u5_mult_87_ab_24__16_, u5_mult_87_ab_24__17_, u5_mult_87_ab_24__18_,
         u5_mult_87_ab_24__19_, u5_mult_87_ab_24__20_, u5_mult_87_ab_24__21_,
         u5_mult_87_ab_24__22_, u5_mult_87_ab_24__23_, u5_mult_87_ab_24__24_,
         u5_mult_87_ab_24__25_, u5_mult_87_ab_24__26_, u5_mult_87_ab_24__27_,
         u5_mult_87_ab_24__28_, u5_mult_87_ab_24__29_, u5_mult_87_ab_24__30_,
         u5_mult_87_ab_24__31_, u5_mult_87_ab_24__32_, u5_mult_87_ab_24__33_,
         u5_mult_87_ab_24__34_, u5_mult_87_ab_24__35_, u5_mult_87_ab_24__36_,
         u5_mult_87_ab_24__37_, u5_mult_87_ab_24__38_, u5_mult_87_ab_24__39_,
         u5_mult_87_ab_24__40_, u5_mult_87_ab_24__41_, u5_mult_87_ab_24__42_,
         u5_mult_87_ab_24__43_, u5_mult_87_ab_24__44_, u5_mult_87_ab_24__45_,
         u5_mult_87_ab_24__46_, u5_mult_87_ab_24__47_, u5_mult_87_ab_24__48_,
         u5_mult_87_ab_24__49_, u5_mult_87_ab_24__50_, u5_mult_87_ab_24__51_,
         u5_mult_87_ab_24__52_, u5_mult_87_ab_25__0_, u5_mult_87_ab_25__1_,
         u5_mult_87_ab_25__2_, u5_mult_87_ab_25__3_, u5_mult_87_ab_25__4_,
         u5_mult_87_ab_25__5_, u5_mult_87_ab_25__6_, u5_mult_87_ab_25__7_,
         u5_mult_87_ab_25__8_, u5_mult_87_ab_25__9_, u5_mult_87_ab_25__10_,
         u5_mult_87_ab_25__11_, u5_mult_87_ab_25__12_, u5_mult_87_ab_25__13_,
         u5_mult_87_ab_25__14_, u5_mult_87_ab_25__15_, u5_mult_87_ab_25__16_,
         u5_mult_87_ab_25__17_, u5_mult_87_ab_25__18_, u5_mult_87_ab_25__19_,
         u5_mult_87_ab_25__20_, u5_mult_87_ab_25__21_, u5_mult_87_ab_25__22_,
         u5_mult_87_ab_25__23_, u5_mult_87_ab_25__24_, u5_mult_87_ab_25__25_,
         u5_mult_87_ab_25__26_, u5_mult_87_ab_25__27_, u5_mult_87_ab_25__28_,
         u5_mult_87_ab_25__29_, u5_mult_87_ab_25__30_, u5_mult_87_ab_25__31_,
         u5_mult_87_ab_25__32_, u5_mult_87_ab_25__33_, u5_mult_87_ab_25__34_,
         u5_mult_87_ab_25__35_, u5_mult_87_ab_25__36_, u5_mult_87_ab_25__37_,
         u5_mult_87_ab_25__38_, u5_mult_87_ab_25__39_, u5_mult_87_ab_25__40_,
         u5_mult_87_ab_25__41_, u5_mult_87_ab_25__42_, u5_mult_87_ab_25__43_,
         u5_mult_87_ab_25__44_, u5_mult_87_ab_25__45_, u5_mult_87_ab_25__46_,
         u5_mult_87_ab_25__47_, u5_mult_87_ab_25__48_, u5_mult_87_ab_25__49_,
         u5_mult_87_ab_25__50_, u5_mult_87_ab_25__51_, u5_mult_87_ab_25__52_,
         u5_mult_87_ab_26__0_, u5_mult_87_ab_26__1_, u5_mult_87_ab_26__2_,
         u5_mult_87_ab_26__3_, u5_mult_87_ab_26__4_, u5_mult_87_ab_26__5_,
         u5_mult_87_ab_26__6_, u5_mult_87_ab_26__7_, u5_mult_87_ab_26__8_,
         u5_mult_87_ab_26__9_, u5_mult_87_ab_26__10_, u5_mult_87_ab_26__11_,
         u5_mult_87_ab_26__12_, u5_mult_87_ab_26__13_, u5_mult_87_ab_26__14_,
         u5_mult_87_ab_26__15_, u5_mult_87_ab_26__16_, u5_mult_87_ab_26__17_,
         u5_mult_87_ab_26__18_, u5_mult_87_ab_26__19_, u5_mult_87_ab_26__20_,
         u5_mult_87_ab_26__21_, u5_mult_87_ab_26__22_, u5_mult_87_ab_26__23_,
         u5_mult_87_ab_26__24_, u5_mult_87_ab_26__25_, u5_mult_87_ab_26__26_,
         u5_mult_87_ab_26__27_, u5_mult_87_ab_26__28_, u5_mult_87_ab_26__29_,
         u5_mult_87_ab_26__30_, u5_mult_87_ab_26__31_, u5_mult_87_ab_26__32_,
         u5_mult_87_ab_26__33_, u5_mult_87_ab_26__34_, u5_mult_87_ab_26__35_,
         u5_mult_87_ab_26__36_, u5_mult_87_ab_26__37_, u5_mult_87_ab_26__38_,
         u5_mult_87_ab_26__39_, u5_mult_87_ab_26__40_, u5_mult_87_ab_26__41_,
         u5_mult_87_ab_26__42_, u5_mult_87_ab_26__43_, u5_mult_87_ab_26__44_,
         u5_mult_87_ab_26__45_, u5_mult_87_ab_26__46_, u5_mult_87_ab_26__47_,
         u5_mult_87_ab_26__48_, u5_mult_87_ab_26__49_, u5_mult_87_ab_26__50_,
         u5_mult_87_ab_26__51_, u5_mult_87_ab_26__52_, u5_mult_87_ab_27__0_,
         u5_mult_87_ab_27__1_, u5_mult_87_ab_27__2_, u5_mult_87_ab_27__3_,
         u5_mult_87_ab_27__4_, u5_mult_87_ab_27__5_, u5_mult_87_ab_27__6_,
         u5_mult_87_ab_27__7_, u5_mult_87_ab_27__8_, u5_mult_87_ab_27__9_,
         u5_mult_87_ab_27__10_, u5_mult_87_ab_27__11_, u5_mult_87_ab_27__12_,
         u5_mult_87_ab_27__13_, u5_mult_87_ab_27__14_, u5_mult_87_ab_27__15_,
         u5_mult_87_ab_27__16_, u5_mult_87_ab_27__17_, u5_mult_87_ab_27__18_,
         u5_mult_87_ab_27__19_, u5_mult_87_ab_27__20_, u5_mult_87_ab_27__21_,
         u5_mult_87_ab_27__22_, u5_mult_87_ab_27__23_, u5_mult_87_ab_27__24_,
         u5_mult_87_ab_27__25_, u5_mult_87_ab_27__26_, u5_mult_87_ab_27__27_,
         u5_mult_87_ab_27__28_, u5_mult_87_ab_27__29_, u5_mult_87_ab_27__30_,
         u5_mult_87_ab_27__31_, u5_mult_87_ab_27__32_, u5_mult_87_ab_27__33_,
         u5_mult_87_ab_27__34_, u5_mult_87_ab_27__35_, u5_mult_87_ab_27__36_,
         u5_mult_87_ab_27__37_, u5_mult_87_ab_27__38_, u5_mult_87_ab_27__39_,
         u5_mult_87_ab_27__40_, u5_mult_87_ab_27__41_, u5_mult_87_ab_27__42_,
         u5_mult_87_ab_27__43_, u5_mult_87_ab_27__44_, u5_mult_87_ab_27__45_,
         u5_mult_87_ab_27__46_, u5_mult_87_ab_27__47_, u5_mult_87_ab_27__48_,
         u5_mult_87_ab_27__49_, u5_mult_87_ab_27__50_, u5_mult_87_ab_27__51_,
         u5_mult_87_ab_27__52_, u5_mult_87_ab_28__0_, u5_mult_87_ab_28__1_,
         u5_mult_87_ab_28__2_, u5_mult_87_ab_28__3_, u5_mult_87_ab_28__4_,
         u5_mult_87_ab_28__5_, u5_mult_87_ab_28__6_, u5_mult_87_ab_28__7_,
         u5_mult_87_ab_28__8_, u5_mult_87_ab_28__9_, u5_mult_87_ab_28__10_,
         u5_mult_87_ab_28__11_, u5_mult_87_ab_28__12_, u5_mult_87_ab_28__13_,
         u5_mult_87_ab_28__14_, u5_mult_87_ab_28__15_, u5_mult_87_ab_28__16_,
         u5_mult_87_ab_28__17_, u5_mult_87_ab_28__18_, u5_mult_87_ab_28__19_,
         u5_mult_87_ab_28__20_, u5_mult_87_ab_28__21_, u5_mult_87_ab_28__22_,
         u5_mult_87_ab_28__23_, u5_mult_87_ab_28__24_, u5_mult_87_ab_28__25_,
         u5_mult_87_ab_28__26_, u5_mult_87_ab_28__27_, u5_mult_87_ab_28__28_,
         u5_mult_87_ab_28__29_, u5_mult_87_ab_28__30_, u5_mult_87_ab_28__31_,
         u5_mult_87_ab_28__32_, u5_mult_87_ab_28__33_, u5_mult_87_ab_28__34_,
         u5_mult_87_ab_28__35_, u5_mult_87_ab_28__36_, u5_mult_87_ab_28__37_,
         u5_mult_87_ab_28__38_, u5_mult_87_ab_28__39_, u5_mult_87_ab_28__40_,
         u5_mult_87_ab_28__41_, u5_mult_87_ab_28__42_, u5_mult_87_ab_28__43_,
         u5_mult_87_ab_28__44_, u5_mult_87_ab_28__45_, u5_mult_87_ab_28__46_,
         u5_mult_87_ab_28__47_, u5_mult_87_ab_28__48_, u5_mult_87_ab_28__49_,
         u5_mult_87_ab_28__50_, u5_mult_87_ab_28__51_, u5_mult_87_ab_28__52_,
         u5_mult_87_ab_29__0_, u5_mult_87_ab_29__1_, u5_mult_87_ab_29__2_,
         u5_mult_87_ab_29__3_, u5_mult_87_ab_29__4_, u5_mult_87_ab_29__5_,
         u5_mult_87_ab_29__6_, u5_mult_87_ab_29__7_, u5_mult_87_ab_29__8_,
         u5_mult_87_ab_29__9_, u5_mult_87_ab_29__10_, u5_mult_87_ab_29__11_,
         u5_mult_87_ab_29__12_, u5_mult_87_ab_29__13_, u5_mult_87_ab_29__14_,
         u5_mult_87_ab_29__15_, u5_mult_87_ab_29__16_, u5_mult_87_ab_29__17_,
         u5_mult_87_ab_29__18_, u5_mult_87_ab_29__19_, u5_mult_87_ab_29__20_,
         u5_mult_87_ab_29__21_, u5_mult_87_ab_29__22_, u5_mult_87_ab_29__23_,
         u5_mult_87_ab_29__24_, u5_mult_87_ab_29__25_, u5_mult_87_ab_29__26_,
         u5_mult_87_ab_29__27_, u5_mult_87_ab_29__28_, u5_mult_87_ab_29__29_,
         u5_mult_87_ab_29__30_, u5_mult_87_ab_29__31_, u5_mult_87_ab_29__32_,
         u5_mult_87_ab_29__33_, u5_mult_87_ab_29__34_, u5_mult_87_ab_29__35_,
         u5_mult_87_ab_29__36_, u5_mult_87_ab_29__37_, u5_mult_87_ab_29__38_,
         u5_mult_87_ab_29__39_, u5_mult_87_ab_29__40_, u5_mult_87_ab_29__41_,
         u5_mult_87_ab_29__42_, u5_mult_87_ab_29__43_, u5_mult_87_ab_29__44_,
         u5_mult_87_ab_29__45_, u5_mult_87_ab_29__46_, u5_mult_87_ab_29__47_,
         u5_mult_87_ab_29__48_, u5_mult_87_ab_29__49_, u5_mult_87_ab_29__50_,
         u5_mult_87_ab_29__51_, u5_mult_87_ab_29__52_, u5_mult_87_ab_30__0_,
         u5_mult_87_ab_30__1_, u5_mult_87_ab_30__2_, u5_mult_87_ab_30__3_,
         u5_mult_87_ab_30__4_, u5_mult_87_ab_30__5_, u5_mult_87_ab_30__6_,
         u5_mult_87_ab_30__7_, u5_mult_87_ab_30__8_, u5_mult_87_ab_30__9_,
         u5_mult_87_ab_30__10_, u5_mult_87_ab_30__11_, u5_mult_87_ab_30__12_,
         u5_mult_87_ab_30__13_, u5_mult_87_ab_30__14_, u5_mult_87_ab_30__15_,
         u5_mult_87_ab_30__16_, u5_mult_87_ab_30__17_, u5_mult_87_ab_30__18_,
         u5_mult_87_ab_30__19_, u5_mult_87_ab_30__20_, u5_mult_87_ab_30__21_,
         u5_mult_87_ab_30__22_, u5_mult_87_ab_30__23_, u5_mult_87_ab_30__24_,
         u5_mult_87_ab_30__25_, u5_mult_87_ab_30__26_, u5_mult_87_ab_30__27_,
         u5_mult_87_ab_30__28_, u5_mult_87_ab_30__29_, u5_mult_87_ab_30__30_,
         u5_mult_87_ab_30__31_, u5_mult_87_ab_30__32_, u5_mult_87_ab_30__33_,
         u5_mult_87_ab_30__34_, u5_mult_87_ab_30__35_, u5_mult_87_ab_30__36_,
         u5_mult_87_ab_30__37_, u5_mult_87_ab_30__38_, u5_mult_87_ab_30__39_,
         u5_mult_87_ab_30__40_, u5_mult_87_ab_30__41_, u5_mult_87_ab_30__42_,
         u5_mult_87_ab_30__43_, u5_mult_87_ab_30__44_, u5_mult_87_ab_30__45_,
         u5_mult_87_ab_30__46_, u5_mult_87_ab_30__47_, u5_mult_87_ab_30__48_,
         u5_mult_87_ab_30__49_, u5_mult_87_ab_30__50_, u5_mult_87_ab_30__51_,
         u5_mult_87_ab_30__52_, u5_mult_87_ab_31__0_, u5_mult_87_ab_31__1_,
         u5_mult_87_ab_31__2_, u5_mult_87_ab_31__3_, u5_mult_87_ab_31__4_,
         u5_mult_87_ab_31__5_, u5_mult_87_ab_31__6_, u5_mult_87_ab_31__7_,
         u5_mult_87_ab_31__8_, u5_mult_87_ab_31__9_, u5_mult_87_ab_31__10_,
         u5_mult_87_ab_31__11_, u5_mult_87_ab_31__12_, u5_mult_87_ab_31__13_,
         u5_mult_87_ab_31__14_, u5_mult_87_ab_31__15_, u5_mult_87_ab_31__16_,
         u5_mult_87_ab_31__17_, u5_mult_87_ab_31__18_, u5_mult_87_ab_31__19_,
         u5_mult_87_ab_31__20_, u5_mult_87_ab_31__21_, u5_mult_87_ab_31__22_,
         u5_mult_87_ab_31__23_, u5_mult_87_ab_31__24_, u5_mult_87_ab_31__25_,
         u5_mult_87_ab_31__26_, u5_mult_87_ab_31__27_, u5_mult_87_ab_31__28_,
         u5_mult_87_ab_31__29_, u5_mult_87_ab_31__30_, u5_mult_87_ab_31__31_,
         u5_mult_87_ab_31__32_, u5_mult_87_ab_31__33_, u5_mult_87_ab_31__34_,
         u5_mult_87_ab_31__35_, u5_mult_87_ab_31__36_, u5_mult_87_ab_31__37_,
         u5_mult_87_ab_31__38_, u5_mult_87_ab_31__39_, u5_mult_87_ab_31__40_,
         u5_mult_87_ab_31__41_, u5_mult_87_ab_31__42_, u5_mult_87_ab_31__43_,
         u5_mult_87_ab_31__44_, u5_mult_87_ab_31__45_, u5_mult_87_ab_31__46_,
         u5_mult_87_ab_31__47_, u5_mult_87_ab_31__48_, u5_mult_87_ab_31__49_,
         u5_mult_87_ab_31__50_, u5_mult_87_ab_31__51_, u5_mult_87_ab_31__52_,
         u5_mult_87_ab_32__0_, u5_mult_87_ab_32__1_, u5_mult_87_ab_32__2_,
         u5_mult_87_ab_32__3_, u5_mult_87_ab_32__4_, u5_mult_87_ab_32__5_,
         u5_mult_87_ab_32__6_, u5_mult_87_ab_32__7_, u5_mult_87_ab_32__8_,
         u5_mult_87_ab_32__9_, u5_mult_87_ab_32__10_, u5_mult_87_ab_32__11_,
         u5_mult_87_ab_32__12_, u5_mult_87_ab_32__13_, u5_mult_87_ab_32__14_,
         u5_mult_87_ab_32__15_, u5_mult_87_ab_32__16_, u5_mult_87_ab_32__17_,
         u5_mult_87_ab_32__18_, u5_mult_87_ab_32__19_, u5_mult_87_ab_32__20_,
         u5_mult_87_ab_32__21_, u5_mult_87_ab_32__22_, u5_mult_87_ab_32__23_,
         u5_mult_87_ab_32__24_, u5_mult_87_ab_32__25_, u5_mult_87_ab_32__26_,
         u5_mult_87_ab_32__27_, u5_mult_87_ab_32__28_, u5_mult_87_ab_32__29_,
         u5_mult_87_ab_32__30_, u5_mult_87_ab_32__31_, u5_mult_87_ab_32__32_,
         u5_mult_87_ab_32__33_, u5_mult_87_ab_32__34_, u5_mult_87_ab_32__35_,
         u5_mult_87_ab_32__36_, u5_mult_87_ab_32__37_, u5_mult_87_ab_32__38_,
         u5_mult_87_ab_32__39_, u5_mult_87_ab_32__40_, u5_mult_87_ab_32__41_,
         u5_mult_87_ab_32__42_, u5_mult_87_ab_32__43_, u5_mult_87_ab_32__44_,
         u5_mult_87_ab_32__45_, u5_mult_87_ab_32__46_, u5_mult_87_ab_32__47_,
         u5_mult_87_ab_32__48_, u5_mult_87_ab_32__49_, u5_mult_87_ab_32__50_,
         u5_mult_87_ab_32__51_, u5_mult_87_ab_32__52_, u5_mult_87_ab_33__0_,
         u5_mult_87_ab_33__1_, u5_mult_87_ab_33__2_, u5_mult_87_ab_33__3_,
         u5_mult_87_ab_33__4_, u5_mult_87_ab_33__5_, u5_mult_87_ab_33__6_,
         u5_mult_87_ab_33__7_, u5_mult_87_ab_33__8_, u5_mult_87_ab_33__9_,
         u5_mult_87_ab_33__10_, u5_mult_87_ab_33__11_, u5_mult_87_ab_33__12_,
         u5_mult_87_ab_33__13_, u5_mult_87_ab_33__14_, u5_mult_87_ab_33__15_,
         u5_mult_87_ab_33__16_, u5_mult_87_ab_33__17_, u5_mult_87_ab_33__18_,
         u5_mult_87_ab_33__19_, u5_mult_87_ab_33__20_, u5_mult_87_ab_33__21_,
         u5_mult_87_ab_33__22_, u5_mult_87_ab_33__23_, u5_mult_87_ab_33__24_,
         u5_mult_87_ab_33__25_, u5_mult_87_ab_33__26_, u5_mult_87_ab_33__27_,
         u5_mult_87_ab_33__28_, u5_mult_87_ab_33__29_, u5_mult_87_ab_33__30_,
         u5_mult_87_ab_33__31_, u5_mult_87_ab_33__32_, u5_mult_87_ab_33__33_,
         u5_mult_87_ab_33__34_, u5_mult_87_ab_33__35_, u5_mult_87_ab_33__36_,
         u5_mult_87_ab_33__37_, u5_mult_87_ab_33__38_, u5_mult_87_ab_33__39_,
         u5_mult_87_ab_33__40_, u5_mult_87_ab_33__41_, u5_mult_87_ab_33__42_,
         u5_mult_87_ab_33__43_, u5_mult_87_ab_33__44_, u5_mult_87_ab_33__45_,
         u5_mult_87_ab_33__46_, u5_mult_87_ab_33__47_, u5_mult_87_ab_33__48_,
         u5_mult_87_ab_33__49_, u5_mult_87_ab_33__50_, u5_mult_87_ab_33__51_,
         u5_mult_87_ab_33__52_, u5_mult_87_ab_34__0_, u5_mult_87_ab_34__1_,
         u5_mult_87_ab_34__2_, u5_mult_87_ab_34__3_, u5_mult_87_ab_34__4_,
         u5_mult_87_ab_34__5_, u5_mult_87_ab_34__6_, u5_mult_87_ab_34__7_,
         u5_mult_87_ab_34__8_, u5_mult_87_ab_34__9_, u5_mult_87_ab_34__10_,
         u5_mult_87_ab_34__11_, u5_mult_87_ab_34__12_, u5_mult_87_ab_34__13_,
         u5_mult_87_ab_34__14_, u5_mult_87_ab_34__15_, u5_mult_87_ab_34__16_,
         u5_mult_87_ab_34__17_, u5_mult_87_ab_34__18_, u5_mult_87_ab_34__19_,
         u5_mult_87_ab_34__20_, u5_mult_87_ab_34__21_, u5_mult_87_ab_34__22_,
         u5_mult_87_ab_34__23_, u5_mult_87_ab_34__24_, u5_mult_87_ab_34__25_,
         u5_mult_87_ab_34__26_, u5_mult_87_ab_34__27_, u5_mult_87_ab_34__28_,
         u5_mult_87_ab_34__29_, u5_mult_87_ab_34__30_, u5_mult_87_ab_34__31_,
         u5_mult_87_ab_34__32_, u5_mult_87_ab_34__33_, u5_mult_87_ab_34__34_,
         u5_mult_87_ab_34__35_, u5_mult_87_ab_34__36_, u5_mult_87_ab_34__37_,
         u5_mult_87_ab_34__38_, u5_mult_87_ab_34__39_, u5_mult_87_ab_34__40_,
         u5_mult_87_ab_34__41_, u5_mult_87_ab_34__42_, u5_mult_87_ab_34__43_,
         u5_mult_87_ab_34__44_, u5_mult_87_ab_34__45_, u5_mult_87_ab_34__46_,
         u5_mult_87_ab_34__47_, u5_mult_87_ab_34__48_, u5_mult_87_ab_34__49_,
         u5_mult_87_ab_34__50_, u5_mult_87_ab_34__51_, u5_mult_87_ab_34__52_,
         u5_mult_87_ab_35__0_, u5_mult_87_ab_35__1_, u5_mult_87_ab_35__2_,
         u5_mult_87_ab_35__3_, u5_mult_87_ab_35__4_, u5_mult_87_ab_35__5_,
         u5_mult_87_ab_35__6_, u5_mult_87_ab_35__7_, u5_mult_87_ab_35__8_,
         u5_mult_87_ab_35__9_, u5_mult_87_ab_35__10_, u5_mult_87_ab_35__11_,
         u5_mult_87_ab_35__12_, u5_mult_87_ab_35__13_, u5_mult_87_ab_35__14_,
         u5_mult_87_ab_35__15_, u5_mult_87_ab_35__16_, u5_mult_87_ab_35__17_,
         u5_mult_87_ab_35__18_, u5_mult_87_ab_35__19_, u5_mult_87_ab_35__20_,
         u5_mult_87_ab_35__21_, u5_mult_87_ab_35__22_, u5_mult_87_ab_35__23_,
         u5_mult_87_ab_35__24_, u5_mult_87_ab_35__25_, u5_mult_87_ab_35__26_,
         u5_mult_87_ab_35__27_, u5_mult_87_ab_35__28_, u5_mult_87_ab_35__29_,
         u5_mult_87_ab_35__30_, u5_mult_87_ab_35__31_, u5_mult_87_ab_35__32_,
         u5_mult_87_ab_35__33_, u5_mult_87_ab_35__34_, u5_mult_87_ab_35__35_,
         u5_mult_87_ab_35__36_, u5_mult_87_ab_35__37_, u5_mult_87_ab_35__38_,
         u5_mult_87_ab_35__39_, u5_mult_87_ab_35__40_, u5_mult_87_ab_35__41_,
         u5_mult_87_ab_35__42_, u5_mult_87_ab_35__43_, u5_mult_87_ab_35__44_,
         u5_mult_87_ab_35__45_, u5_mult_87_ab_35__46_, u5_mult_87_ab_35__47_,
         u5_mult_87_ab_35__48_, u5_mult_87_ab_35__49_, u5_mult_87_ab_35__50_,
         u5_mult_87_ab_35__51_, u5_mult_87_ab_35__52_, u5_mult_87_ab_36__0_,
         u5_mult_87_ab_36__1_, u5_mult_87_ab_36__2_, u5_mult_87_ab_36__3_,
         u5_mult_87_ab_36__4_, u5_mult_87_ab_36__5_, u5_mult_87_ab_36__6_,
         u5_mult_87_ab_36__7_, u5_mult_87_ab_36__8_, u5_mult_87_ab_36__9_,
         u5_mult_87_ab_36__10_, u5_mult_87_ab_36__11_, u5_mult_87_ab_36__12_,
         u5_mult_87_ab_36__13_, u5_mult_87_ab_36__14_, u5_mult_87_ab_36__15_,
         u5_mult_87_ab_36__16_, u5_mult_87_ab_36__17_, u5_mult_87_ab_36__18_,
         u5_mult_87_ab_36__19_, u5_mult_87_ab_36__20_, u5_mult_87_ab_36__21_,
         u5_mult_87_ab_36__22_, u5_mult_87_ab_36__23_, u5_mult_87_ab_36__24_,
         u5_mult_87_ab_36__25_, u5_mult_87_ab_36__26_, u5_mult_87_ab_36__27_,
         u5_mult_87_ab_36__28_, u5_mult_87_ab_36__29_, u5_mult_87_ab_36__30_,
         u5_mult_87_ab_36__31_, u5_mult_87_ab_36__32_, u5_mult_87_ab_36__33_,
         u5_mult_87_ab_36__34_, u5_mult_87_ab_36__35_, u5_mult_87_ab_36__36_,
         u5_mult_87_ab_36__37_, u5_mult_87_ab_36__38_, u5_mult_87_ab_36__39_,
         u5_mult_87_ab_36__40_, u5_mult_87_ab_36__41_, u5_mult_87_ab_36__42_,
         u5_mult_87_ab_36__43_, u5_mult_87_ab_36__44_, u5_mult_87_ab_36__45_,
         u5_mult_87_ab_36__46_, u5_mult_87_ab_36__47_, u5_mult_87_ab_36__48_,
         u5_mult_87_ab_36__49_, u5_mult_87_ab_36__50_, u5_mult_87_ab_36__51_,
         u5_mult_87_ab_36__52_, u5_mult_87_ab_37__0_, u5_mult_87_ab_37__1_,
         u5_mult_87_ab_37__2_, u5_mult_87_ab_37__3_, u5_mult_87_ab_37__4_,
         u5_mult_87_ab_37__5_, u5_mult_87_ab_37__6_, u5_mult_87_ab_37__7_,
         u5_mult_87_ab_37__8_, u5_mult_87_ab_37__9_, u5_mult_87_ab_37__10_,
         u5_mult_87_ab_37__11_, u5_mult_87_ab_37__12_, u5_mult_87_ab_37__13_,
         u5_mult_87_ab_37__14_, u5_mult_87_ab_37__15_, u5_mult_87_ab_37__16_,
         u5_mult_87_ab_37__17_, u5_mult_87_ab_37__18_, u5_mult_87_ab_37__19_,
         u5_mult_87_ab_37__20_, u5_mult_87_ab_37__21_, u5_mult_87_ab_37__22_,
         u5_mult_87_ab_37__23_, u5_mult_87_ab_37__24_, u5_mult_87_ab_37__25_,
         u5_mult_87_ab_37__26_, u5_mult_87_ab_37__27_, u5_mult_87_ab_37__28_,
         u5_mult_87_ab_37__29_, u5_mult_87_ab_37__30_, u5_mult_87_ab_37__31_,
         u5_mult_87_ab_37__32_, u5_mult_87_ab_37__33_, u5_mult_87_ab_37__34_,
         u5_mult_87_ab_37__35_, u5_mult_87_ab_37__36_, u5_mult_87_ab_37__37_,
         u5_mult_87_ab_37__38_, u5_mult_87_ab_37__39_, u5_mult_87_ab_37__40_,
         u5_mult_87_ab_37__41_, u5_mult_87_ab_37__42_, u5_mult_87_ab_37__43_,
         u5_mult_87_ab_37__44_, u5_mult_87_ab_37__45_, u5_mult_87_ab_37__46_,
         u5_mult_87_ab_37__47_, u5_mult_87_ab_37__48_, u5_mult_87_ab_37__49_,
         u5_mult_87_ab_37__50_, u5_mult_87_ab_37__51_, u5_mult_87_ab_37__52_,
         u5_mult_87_ab_38__0_, u5_mult_87_ab_38__1_, u5_mult_87_ab_38__2_,
         u5_mult_87_ab_38__3_, u5_mult_87_ab_38__4_, u5_mult_87_ab_38__5_,
         u5_mult_87_ab_38__6_, u5_mult_87_ab_38__7_, u5_mult_87_ab_38__8_,
         u5_mult_87_ab_38__9_, u5_mult_87_ab_38__10_, u5_mult_87_ab_38__11_,
         u5_mult_87_ab_38__12_, u5_mult_87_ab_38__13_, u5_mult_87_ab_38__14_,
         u5_mult_87_ab_38__15_, u5_mult_87_ab_38__16_, u5_mult_87_ab_38__17_,
         u5_mult_87_ab_38__18_, u5_mult_87_ab_38__19_, u5_mult_87_ab_38__20_,
         u5_mult_87_ab_38__21_, u5_mult_87_ab_38__22_, u5_mult_87_ab_38__23_,
         u5_mult_87_ab_38__24_, u5_mult_87_ab_38__25_, u5_mult_87_ab_38__26_,
         u5_mult_87_ab_38__27_, u5_mult_87_ab_38__28_, u5_mult_87_ab_38__29_,
         u5_mult_87_ab_38__30_, u5_mult_87_ab_38__31_, u5_mult_87_ab_38__32_,
         u5_mult_87_ab_38__33_, u5_mult_87_ab_38__34_, u5_mult_87_ab_38__35_,
         u5_mult_87_ab_38__36_, u5_mult_87_ab_38__37_, u5_mult_87_ab_38__38_,
         u5_mult_87_ab_38__39_, u5_mult_87_ab_38__40_, u5_mult_87_ab_38__41_,
         u5_mult_87_ab_38__42_, u5_mult_87_ab_38__43_, u5_mult_87_ab_38__44_,
         u5_mult_87_ab_38__45_, u5_mult_87_ab_38__46_, u5_mult_87_ab_38__47_,
         u5_mult_87_ab_38__48_, u5_mult_87_ab_38__49_, u5_mult_87_ab_38__50_,
         u5_mult_87_ab_38__51_, u5_mult_87_ab_38__52_, u5_mult_87_ab_39__0_,
         u5_mult_87_ab_39__1_, u5_mult_87_ab_39__2_, u5_mult_87_ab_39__3_,
         u5_mult_87_ab_39__4_, u5_mult_87_ab_39__5_, u5_mult_87_ab_39__6_,
         u5_mult_87_ab_39__7_, u5_mult_87_ab_39__8_, u5_mult_87_ab_39__9_,
         u5_mult_87_ab_39__10_, u5_mult_87_ab_39__11_, u5_mult_87_ab_39__12_,
         u5_mult_87_ab_39__13_, u5_mult_87_ab_39__14_, u5_mult_87_ab_39__15_,
         u5_mult_87_ab_39__16_, u5_mult_87_ab_39__17_, u5_mult_87_ab_39__18_,
         u5_mult_87_ab_39__19_, u5_mult_87_ab_39__20_, u5_mult_87_ab_39__21_,
         u5_mult_87_ab_39__22_, u5_mult_87_ab_39__23_, u5_mult_87_ab_39__24_,
         u5_mult_87_ab_39__25_, u5_mult_87_ab_39__26_, u5_mult_87_ab_39__27_,
         u5_mult_87_ab_39__28_, u5_mult_87_ab_39__29_, u5_mult_87_ab_39__30_,
         u5_mult_87_ab_39__31_, u5_mult_87_ab_39__32_, u5_mult_87_ab_39__33_,
         u5_mult_87_ab_39__34_, u5_mult_87_ab_39__35_, u5_mult_87_ab_39__36_,
         u5_mult_87_ab_39__37_, u5_mult_87_ab_39__38_, u5_mult_87_ab_39__39_,
         u5_mult_87_ab_39__40_, u5_mult_87_ab_39__41_, u5_mult_87_ab_39__42_,
         u5_mult_87_ab_39__43_, u5_mult_87_ab_39__44_, u5_mult_87_ab_39__45_,
         u5_mult_87_ab_39__46_, u5_mult_87_ab_39__47_, u5_mult_87_ab_39__48_,
         u5_mult_87_ab_39__49_, u5_mult_87_ab_39__50_, u5_mult_87_ab_39__51_,
         u5_mult_87_ab_39__52_, u5_mult_87_ab_40__0_, u5_mult_87_ab_40__1_,
         u5_mult_87_ab_40__2_, u5_mult_87_ab_40__3_, u5_mult_87_ab_40__4_,
         u5_mult_87_ab_40__5_, u5_mult_87_ab_40__6_, u5_mult_87_ab_40__7_,
         u5_mult_87_ab_40__8_, u5_mult_87_ab_40__9_, u5_mult_87_ab_40__10_,
         u5_mult_87_ab_40__11_, u5_mult_87_ab_40__12_, u5_mult_87_ab_40__13_,
         u5_mult_87_ab_40__14_, u5_mult_87_ab_40__15_, u5_mult_87_ab_40__16_,
         u5_mult_87_ab_40__17_, u5_mult_87_ab_40__18_, u5_mult_87_ab_40__19_,
         u5_mult_87_ab_40__20_, u5_mult_87_ab_40__21_, u5_mult_87_ab_40__22_,
         u5_mult_87_ab_40__23_, u5_mult_87_ab_40__24_, u5_mult_87_ab_40__25_,
         u5_mult_87_ab_40__26_, u5_mult_87_ab_40__27_, u5_mult_87_ab_40__28_,
         u5_mult_87_ab_40__29_, u5_mult_87_ab_40__30_, u5_mult_87_ab_40__31_,
         u5_mult_87_ab_40__32_, u5_mult_87_ab_40__33_, u5_mult_87_ab_40__34_,
         u5_mult_87_ab_40__35_, u5_mult_87_ab_40__36_, u5_mult_87_ab_40__37_,
         u5_mult_87_ab_40__38_, u5_mult_87_ab_40__39_, u5_mult_87_ab_40__40_,
         u5_mult_87_ab_40__41_, u5_mult_87_ab_40__42_, u5_mult_87_ab_40__43_,
         u5_mult_87_ab_40__44_, u5_mult_87_ab_40__45_, u5_mult_87_ab_40__46_,
         u5_mult_87_ab_40__47_, u5_mult_87_ab_40__48_, u5_mult_87_ab_40__49_,
         u5_mult_87_ab_40__50_, u5_mult_87_ab_40__51_, u5_mult_87_ab_40__52_,
         u5_mult_87_ab_41__0_, u5_mult_87_ab_41__1_, u5_mult_87_ab_41__2_,
         u5_mult_87_ab_41__3_, u5_mult_87_ab_41__4_, u5_mult_87_ab_41__5_,
         u5_mult_87_ab_41__6_, u5_mult_87_ab_41__7_, u5_mult_87_ab_41__8_,
         u5_mult_87_ab_41__9_, u5_mult_87_ab_41__10_, u5_mult_87_ab_41__11_,
         u5_mult_87_ab_41__12_, u5_mult_87_ab_41__13_, u5_mult_87_ab_41__14_,
         u5_mult_87_ab_41__15_, u5_mult_87_ab_41__16_, u5_mult_87_ab_41__17_,
         u5_mult_87_ab_41__18_, u5_mult_87_ab_41__19_, u5_mult_87_ab_41__20_,
         u5_mult_87_ab_41__21_, u5_mult_87_ab_41__22_, u5_mult_87_ab_41__23_,
         u5_mult_87_ab_41__24_, u5_mult_87_ab_41__25_, u5_mult_87_ab_41__26_,
         u5_mult_87_ab_41__27_, u5_mult_87_ab_41__28_, u5_mult_87_ab_41__29_,
         u5_mult_87_ab_41__30_, u5_mult_87_ab_41__31_, u5_mult_87_ab_41__32_,
         u5_mult_87_ab_41__33_, u5_mult_87_ab_41__34_, u5_mult_87_ab_41__35_,
         u5_mult_87_ab_41__36_, u5_mult_87_ab_41__37_, u5_mult_87_ab_41__38_,
         u5_mult_87_ab_41__39_, u5_mult_87_ab_41__40_, u5_mult_87_ab_41__41_,
         u5_mult_87_ab_41__42_, u5_mult_87_ab_41__43_, u5_mult_87_ab_41__44_,
         u5_mult_87_ab_41__45_, u5_mult_87_ab_41__46_, u5_mult_87_ab_41__47_,
         u5_mult_87_ab_41__48_, u5_mult_87_ab_41__49_, u5_mult_87_ab_41__50_,
         u5_mult_87_ab_41__51_, u5_mult_87_ab_41__52_, u5_mult_87_ab_42__0_,
         u5_mult_87_ab_42__1_, u5_mult_87_ab_42__2_, u5_mult_87_ab_42__3_,
         u5_mult_87_ab_42__4_, u5_mult_87_ab_42__5_, u5_mult_87_ab_42__6_,
         u5_mult_87_ab_42__7_, u5_mult_87_ab_42__8_, u5_mult_87_ab_42__9_,
         u5_mult_87_ab_42__10_, u5_mult_87_ab_42__11_, u5_mult_87_ab_42__12_,
         u5_mult_87_ab_42__13_, u5_mult_87_ab_42__14_, u5_mult_87_ab_42__15_,
         u5_mult_87_ab_42__16_, u5_mult_87_ab_42__17_, u5_mult_87_ab_42__18_,
         u5_mult_87_ab_42__19_, u5_mult_87_ab_42__20_, u5_mult_87_ab_42__21_,
         u5_mult_87_ab_42__22_, u5_mult_87_ab_42__23_, u5_mult_87_ab_42__24_,
         u5_mult_87_ab_42__25_, u5_mult_87_ab_42__26_, u5_mult_87_ab_42__27_,
         u5_mult_87_ab_42__28_, u5_mult_87_ab_42__29_, u5_mult_87_ab_42__30_,
         u5_mult_87_ab_42__31_, u5_mult_87_ab_42__32_, u5_mult_87_ab_42__33_,
         u5_mult_87_ab_42__34_, u5_mult_87_ab_42__35_, u5_mult_87_ab_42__36_,
         u5_mult_87_ab_42__37_, u5_mult_87_ab_42__38_, u5_mult_87_ab_42__39_,
         u5_mult_87_ab_42__40_, u5_mult_87_ab_42__41_, u5_mult_87_ab_42__42_,
         u5_mult_87_ab_42__43_, u5_mult_87_ab_42__44_, u5_mult_87_ab_42__45_,
         u5_mult_87_ab_42__46_, u5_mult_87_ab_42__47_, u5_mult_87_ab_42__48_,
         u5_mult_87_ab_42__49_, u5_mult_87_ab_42__50_, u5_mult_87_ab_42__51_,
         u5_mult_87_ab_42__52_, u5_mult_87_ab_43__0_, u5_mult_87_ab_43__1_,
         u5_mult_87_ab_43__2_, u5_mult_87_ab_43__3_, u5_mult_87_ab_43__4_,
         u5_mult_87_ab_43__5_, u5_mult_87_ab_43__6_, u5_mult_87_ab_43__7_,
         u5_mult_87_ab_43__8_, u5_mult_87_ab_43__9_, u5_mult_87_ab_43__10_,
         u5_mult_87_ab_43__11_, u5_mult_87_ab_43__12_, u5_mult_87_ab_43__13_,
         u5_mult_87_ab_43__14_, u5_mult_87_ab_43__15_, u5_mult_87_ab_43__16_,
         u5_mult_87_ab_43__17_, u5_mult_87_ab_43__18_, u5_mult_87_ab_43__19_,
         u5_mult_87_ab_43__20_, u5_mult_87_ab_43__21_, u5_mult_87_ab_43__22_,
         u5_mult_87_ab_43__23_, u5_mult_87_ab_43__24_, u5_mult_87_ab_43__25_,
         u5_mult_87_ab_43__26_, u5_mult_87_ab_43__27_, u5_mult_87_ab_43__28_,
         u5_mult_87_ab_43__29_, u5_mult_87_ab_43__30_, u5_mult_87_ab_43__31_,
         u5_mult_87_ab_43__32_, u5_mult_87_ab_43__33_, u5_mult_87_ab_43__34_,
         u5_mult_87_ab_43__35_, u5_mult_87_ab_43__36_, u5_mult_87_ab_43__37_,
         u5_mult_87_ab_43__38_, u5_mult_87_ab_43__39_, u5_mult_87_ab_43__40_,
         u5_mult_87_ab_43__41_, u5_mult_87_ab_43__42_, u5_mult_87_ab_43__43_,
         u5_mult_87_ab_43__44_, u5_mult_87_ab_43__45_, u5_mult_87_ab_43__46_,
         u5_mult_87_ab_43__47_, u5_mult_87_ab_43__48_, u5_mult_87_ab_43__49_,
         u5_mult_87_ab_43__50_, u5_mult_87_ab_43__51_, u5_mult_87_ab_43__52_,
         u5_mult_87_ab_44__0_, u5_mult_87_ab_44__1_, u5_mult_87_ab_44__2_,
         u5_mult_87_ab_44__3_, u5_mult_87_ab_44__4_, u5_mult_87_ab_44__5_,
         u5_mult_87_ab_44__6_, u5_mult_87_ab_44__7_, u5_mult_87_ab_44__8_,
         u5_mult_87_ab_44__9_, u5_mult_87_ab_44__10_, u5_mult_87_ab_44__11_,
         u5_mult_87_ab_44__12_, u5_mult_87_ab_44__13_, u5_mult_87_ab_44__14_,
         u5_mult_87_ab_44__15_, u5_mult_87_ab_44__16_, u5_mult_87_ab_44__17_,
         u5_mult_87_ab_44__18_, u5_mult_87_ab_44__19_, u5_mult_87_ab_44__20_,
         u5_mult_87_ab_44__21_, u5_mult_87_ab_44__22_, u5_mult_87_ab_44__23_,
         u5_mult_87_ab_44__24_, u5_mult_87_ab_44__25_, u5_mult_87_ab_44__26_,
         u5_mult_87_ab_44__27_, u5_mult_87_ab_44__28_, u5_mult_87_ab_44__29_,
         u5_mult_87_ab_44__30_, u5_mult_87_ab_44__31_, u5_mult_87_ab_44__32_,
         u5_mult_87_ab_44__33_, u5_mult_87_ab_44__34_, u5_mult_87_ab_44__35_,
         u5_mult_87_ab_44__36_, u5_mult_87_ab_44__37_, u5_mult_87_ab_44__38_,
         u5_mult_87_ab_44__39_, u5_mult_87_ab_44__40_, u5_mult_87_ab_44__41_,
         u5_mult_87_ab_44__42_, u5_mult_87_ab_44__43_, u5_mult_87_ab_44__44_,
         u5_mult_87_ab_44__45_, u5_mult_87_ab_44__46_, u5_mult_87_ab_44__47_,
         u5_mult_87_ab_44__48_, u5_mult_87_ab_44__49_, u5_mult_87_ab_44__50_,
         u5_mult_87_ab_44__51_, u5_mult_87_ab_44__52_, u5_mult_87_ab_45__0_,
         u5_mult_87_ab_45__1_, u5_mult_87_ab_45__2_, u5_mult_87_ab_45__3_,
         u5_mult_87_ab_45__4_, u5_mult_87_ab_45__5_, u5_mult_87_ab_45__6_,
         u5_mult_87_ab_45__7_, u5_mult_87_ab_45__8_, u5_mult_87_ab_45__9_,
         u5_mult_87_ab_45__10_, u5_mult_87_ab_45__11_, u5_mult_87_ab_45__12_,
         u5_mult_87_ab_45__13_, u5_mult_87_ab_45__14_, u5_mult_87_ab_45__15_,
         u5_mult_87_ab_45__16_, u5_mult_87_ab_45__17_, u5_mult_87_ab_45__18_,
         u5_mult_87_ab_45__19_, u5_mult_87_ab_45__20_, u5_mult_87_ab_45__21_,
         u5_mult_87_ab_45__22_, u5_mult_87_ab_45__23_, u5_mult_87_ab_45__24_,
         u5_mult_87_ab_45__25_, u5_mult_87_ab_45__26_, u5_mult_87_ab_45__27_,
         u5_mult_87_ab_45__28_, u5_mult_87_ab_45__29_, u5_mult_87_ab_45__30_,
         u5_mult_87_ab_45__31_, u5_mult_87_ab_45__32_, u5_mult_87_ab_45__33_,
         u5_mult_87_ab_45__34_, u5_mult_87_ab_45__35_, u5_mult_87_ab_45__36_,
         u5_mult_87_ab_45__37_, u5_mult_87_ab_45__38_, u5_mult_87_ab_45__39_,
         u5_mult_87_ab_45__40_, u5_mult_87_ab_45__41_, u5_mult_87_ab_45__42_,
         u5_mult_87_ab_45__43_, u5_mult_87_ab_45__44_, u5_mult_87_ab_45__45_,
         u5_mult_87_ab_45__46_, u5_mult_87_ab_45__47_, u5_mult_87_ab_45__48_,
         u5_mult_87_ab_45__49_, u5_mult_87_ab_45__50_, u5_mult_87_ab_45__51_,
         u5_mult_87_ab_45__52_, u5_mult_87_ab_46__0_, u5_mult_87_ab_46__1_,
         u5_mult_87_ab_46__2_, u5_mult_87_ab_46__3_, u5_mult_87_ab_46__4_,
         u5_mult_87_ab_46__5_, u5_mult_87_ab_46__6_, u5_mult_87_ab_46__7_,
         u5_mult_87_ab_46__8_, u5_mult_87_ab_46__9_, u5_mult_87_ab_46__10_,
         u5_mult_87_ab_46__11_, u5_mult_87_ab_46__12_, u5_mult_87_ab_46__13_,
         u5_mult_87_ab_46__14_, u5_mult_87_ab_46__15_, u5_mult_87_ab_46__16_,
         u5_mult_87_ab_46__17_, u5_mult_87_ab_46__18_, u5_mult_87_ab_46__19_,
         u5_mult_87_ab_46__20_, u5_mult_87_ab_46__21_, u5_mult_87_ab_46__22_,
         u5_mult_87_ab_46__23_, u5_mult_87_ab_46__24_, u5_mult_87_ab_46__25_,
         u5_mult_87_ab_46__26_, u5_mult_87_ab_46__27_, u5_mult_87_ab_46__28_,
         u5_mult_87_ab_46__29_, u5_mult_87_ab_46__30_, u5_mult_87_ab_46__31_,
         u5_mult_87_ab_46__32_, u5_mult_87_ab_46__33_, u5_mult_87_ab_46__34_,
         u5_mult_87_ab_46__35_, u5_mult_87_ab_46__36_, u5_mult_87_ab_46__37_,
         u5_mult_87_ab_46__38_, u5_mult_87_ab_46__39_, u5_mult_87_ab_46__40_,
         u5_mult_87_ab_46__41_, u5_mult_87_ab_46__42_, u5_mult_87_ab_46__43_,
         u5_mult_87_ab_46__44_, u5_mult_87_ab_46__45_, u5_mult_87_ab_46__46_,
         u5_mult_87_ab_46__47_, u5_mult_87_ab_46__48_, u5_mult_87_ab_46__49_,
         u5_mult_87_ab_46__50_, u5_mult_87_ab_46__51_, u5_mult_87_ab_46__52_,
         u5_mult_87_ab_47__0_, u5_mult_87_ab_47__1_, u5_mult_87_ab_47__2_,
         u5_mult_87_ab_47__3_, u5_mult_87_ab_47__4_, u5_mult_87_ab_47__5_,
         u5_mult_87_ab_47__6_, u5_mult_87_ab_47__7_, u5_mult_87_ab_47__8_,
         u5_mult_87_ab_47__9_, u5_mult_87_ab_47__10_, u5_mult_87_ab_47__11_,
         u5_mult_87_ab_47__12_, u5_mult_87_ab_47__13_, u5_mult_87_ab_47__14_,
         u5_mult_87_ab_47__15_, u5_mult_87_ab_47__16_, u5_mult_87_ab_47__17_,
         u5_mult_87_ab_47__18_, u5_mult_87_ab_47__19_, u5_mult_87_ab_47__20_,
         u5_mult_87_ab_47__21_, u5_mult_87_ab_47__22_, u5_mult_87_ab_47__23_,
         u5_mult_87_ab_47__24_, u5_mult_87_ab_47__25_, u5_mult_87_ab_47__26_,
         u5_mult_87_ab_47__27_, u5_mult_87_ab_47__28_, u5_mult_87_ab_47__29_,
         u5_mult_87_ab_47__30_, u5_mult_87_ab_47__31_, u5_mult_87_ab_47__32_,
         u5_mult_87_ab_47__33_, u5_mult_87_ab_47__34_, u5_mult_87_ab_47__35_,
         u5_mult_87_ab_47__36_, u5_mult_87_ab_47__37_, u5_mult_87_ab_47__38_,
         u5_mult_87_ab_47__39_, u5_mult_87_ab_47__40_, u5_mult_87_ab_47__41_,
         u5_mult_87_ab_47__42_, u5_mult_87_ab_47__43_, u5_mult_87_ab_47__44_,
         u5_mult_87_ab_47__45_, u5_mult_87_ab_47__46_, u5_mult_87_ab_47__47_,
         u5_mult_87_ab_47__48_, u5_mult_87_ab_47__49_, u5_mult_87_ab_47__50_,
         u5_mult_87_ab_47__51_, u5_mult_87_ab_47__52_, u5_mult_87_ab_48__0_,
         u5_mult_87_ab_48__1_, u5_mult_87_ab_48__2_, u5_mult_87_ab_48__3_,
         u5_mult_87_ab_48__4_, u5_mult_87_ab_48__5_, u5_mult_87_ab_48__6_,
         u5_mult_87_ab_48__7_, u5_mult_87_ab_48__8_, u5_mult_87_ab_48__9_,
         u5_mult_87_ab_48__10_, u5_mult_87_ab_48__11_, u5_mult_87_ab_48__12_,
         u5_mult_87_ab_48__13_, u5_mult_87_ab_48__14_, u5_mult_87_ab_48__15_,
         u5_mult_87_ab_48__16_, u5_mult_87_ab_48__17_, u5_mult_87_ab_48__18_,
         u5_mult_87_ab_48__19_, u5_mult_87_ab_48__20_, u5_mult_87_ab_48__21_,
         u5_mult_87_ab_48__22_, u5_mult_87_ab_48__23_, u5_mult_87_ab_48__24_,
         u5_mult_87_ab_48__25_, u5_mult_87_ab_48__26_, u5_mult_87_ab_48__27_,
         u5_mult_87_ab_48__28_, u5_mult_87_ab_48__29_, u5_mult_87_ab_48__30_,
         u5_mult_87_ab_48__31_, u5_mult_87_ab_48__32_, u5_mult_87_ab_48__33_,
         u5_mult_87_ab_48__34_, u5_mult_87_ab_48__35_, u5_mult_87_ab_48__36_,
         u5_mult_87_ab_48__37_, u5_mult_87_ab_48__38_, u5_mult_87_ab_48__39_,
         u5_mult_87_ab_48__40_, u5_mult_87_ab_48__41_, u5_mult_87_ab_48__42_,
         u5_mult_87_ab_48__43_, u5_mult_87_ab_48__44_, u5_mult_87_ab_48__45_,
         u5_mult_87_ab_48__46_, u5_mult_87_ab_48__47_, u5_mult_87_ab_48__48_,
         u5_mult_87_ab_48__49_, u5_mult_87_ab_48__50_, u5_mult_87_ab_48__51_,
         u5_mult_87_ab_48__52_, u5_mult_87_ab_49__0_, u5_mult_87_ab_49__1_,
         u5_mult_87_ab_49__2_, u5_mult_87_ab_49__3_, u5_mult_87_ab_49__4_,
         u5_mult_87_ab_49__5_, u5_mult_87_ab_49__6_, u5_mult_87_ab_49__7_,
         u5_mult_87_ab_49__8_, u5_mult_87_ab_49__9_, u5_mult_87_ab_49__10_,
         u5_mult_87_ab_49__11_, u5_mult_87_ab_49__12_, u5_mult_87_ab_49__13_,
         u5_mult_87_ab_49__14_, u5_mult_87_ab_49__15_, u5_mult_87_ab_49__16_,
         u5_mult_87_ab_49__17_, u5_mult_87_ab_49__18_, u5_mult_87_ab_49__19_,
         u5_mult_87_ab_49__20_, u5_mult_87_ab_49__21_, u5_mult_87_ab_49__22_,
         u5_mult_87_ab_49__23_, u5_mult_87_ab_49__24_, u5_mult_87_ab_49__25_,
         u5_mult_87_ab_49__26_, u5_mult_87_ab_49__27_, u5_mult_87_ab_49__28_,
         u5_mult_87_ab_49__29_, u5_mult_87_ab_49__30_, u5_mult_87_ab_49__31_,
         u5_mult_87_ab_49__32_, u5_mult_87_ab_49__33_, u5_mult_87_ab_49__34_,
         u5_mult_87_ab_49__35_, u5_mult_87_ab_49__36_, u5_mult_87_ab_49__37_,
         u5_mult_87_ab_49__38_, u5_mult_87_ab_49__39_, u5_mult_87_ab_49__40_,
         u5_mult_87_ab_49__41_, u5_mult_87_ab_49__42_, u5_mult_87_ab_49__43_,
         u5_mult_87_ab_49__44_, u5_mult_87_ab_49__45_, u5_mult_87_ab_49__46_,
         u5_mult_87_ab_49__47_, u5_mult_87_ab_49__48_, u5_mult_87_ab_49__49_,
         u5_mult_87_ab_49__50_, u5_mult_87_ab_49__51_, u5_mult_87_ab_49__52_,
         u5_mult_87_ab_50__0_, u5_mult_87_ab_50__1_, u5_mult_87_ab_50__2_,
         u5_mult_87_ab_50__3_, u5_mult_87_ab_50__4_, u5_mult_87_ab_50__5_,
         u5_mult_87_ab_50__6_, u5_mult_87_ab_50__7_, u5_mult_87_ab_50__8_,
         u5_mult_87_ab_50__9_, u5_mult_87_ab_50__10_, u5_mult_87_ab_50__11_,
         u5_mult_87_ab_50__12_, u5_mult_87_ab_50__13_, u5_mult_87_ab_50__14_,
         u5_mult_87_ab_50__15_, u5_mult_87_ab_50__16_, u5_mult_87_ab_50__17_,
         u5_mult_87_ab_50__18_, u5_mult_87_ab_50__19_, u5_mult_87_ab_50__20_,
         u5_mult_87_ab_50__21_, u5_mult_87_ab_50__22_, u5_mult_87_ab_50__23_,
         u5_mult_87_ab_50__24_, u5_mult_87_ab_50__25_, u5_mult_87_ab_50__26_,
         u5_mult_87_ab_50__27_, u5_mult_87_ab_50__28_, u5_mult_87_ab_50__29_,
         u5_mult_87_ab_50__30_, u5_mult_87_ab_50__31_, u5_mult_87_ab_50__32_,
         u5_mult_87_ab_50__33_, u5_mult_87_ab_50__34_, u5_mult_87_ab_50__35_,
         u5_mult_87_ab_50__36_, u5_mult_87_ab_50__37_, u5_mult_87_ab_50__38_,
         u5_mult_87_ab_50__39_, u5_mult_87_ab_50__40_, u5_mult_87_ab_50__41_,
         u5_mult_87_ab_50__42_, u5_mult_87_ab_50__43_, u5_mult_87_ab_50__44_,
         u5_mult_87_ab_50__45_, u5_mult_87_ab_50__46_, u5_mult_87_ab_50__47_,
         u5_mult_87_ab_50__48_, u5_mult_87_ab_50__49_, u5_mult_87_ab_50__50_,
         u5_mult_87_ab_50__51_, u5_mult_87_ab_50__52_, u5_mult_87_ab_51__0_,
         u5_mult_87_ab_51__1_, u5_mult_87_ab_51__2_, u5_mult_87_ab_51__3_,
         u5_mult_87_ab_51__4_, u5_mult_87_ab_51__5_, u5_mult_87_ab_51__6_,
         u5_mult_87_ab_51__7_, u5_mult_87_ab_51__8_, u5_mult_87_ab_51__9_,
         u5_mult_87_ab_51__10_, u5_mult_87_ab_51__11_, u5_mult_87_ab_51__12_,
         u5_mult_87_ab_51__13_, u5_mult_87_ab_51__14_, u5_mult_87_ab_51__15_,
         u5_mult_87_ab_51__16_, u5_mult_87_ab_51__17_, u5_mult_87_ab_51__18_,
         u5_mult_87_ab_51__19_, u5_mult_87_ab_51__20_, u5_mult_87_ab_51__21_,
         u5_mult_87_ab_51__22_, u5_mult_87_ab_51__23_, u5_mult_87_ab_51__24_,
         u5_mult_87_ab_51__25_, u5_mult_87_ab_51__26_, u5_mult_87_ab_51__27_,
         u5_mult_87_ab_51__28_, u5_mult_87_ab_51__29_, u5_mult_87_ab_51__30_,
         u5_mult_87_ab_51__31_, u5_mult_87_ab_51__32_, u5_mult_87_ab_51__33_,
         u5_mult_87_ab_51__34_, u5_mult_87_ab_51__35_, u5_mult_87_ab_51__36_,
         u5_mult_87_ab_51__37_, u5_mult_87_ab_51__38_, u5_mult_87_ab_51__39_,
         u5_mult_87_ab_51__40_, u5_mult_87_ab_51__41_, u5_mult_87_ab_51__42_,
         u5_mult_87_ab_51__43_, u5_mult_87_ab_51__44_, u5_mult_87_ab_51__45_,
         u5_mult_87_ab_51__46_, u5_mult_87_ab_51__47_, u5_mult_87_ab_51__48_,
         u5_mult_87_ab_51__49_, u5_mult_87_ab_51__50_, u5_mult_87_ab_51__51_,
         u5_mult_87_ab_51__52_, u5_mult_87_ab_52__0_, u5_mult_87_ab_52__1_,
         u5_mult_87_ab_52__2_, u5_mult_87_ab_52__3_, u5_mult_87_ab_52__4_,
         u5_mult_87_ab_52__5_, u5_mult_87_ab_52__6_, u5_mult_87_ab_52__7_,
         u5_mult_87_ab_52__8_, u5_mult_87_ab_52__9_, u5_mult_87_ab_52__10_,
         u5_mult_87_ab_52__11_, u5_mult_87_ab_52__12_, u5_mult_87_ab_52__13_,
         u5_mult_87_ab_52__14_, u5_mult_87_ab_52__15_, u5_mult_87_ab_52__16_,
         u5_mult_87_ab_52__17_, u5_mult_87_ab_52__18_, u5_mult_87_ab_52__19_,
         u5_mult_87_ab_52__20_, u5_mult_87_ab_52__21_, u5_mult_87_ab_52__22_,
         u5_mult_87_ab_52__23_, u5_mult_87_ab_52__24_, u5_mult_87_ab_52__25_,
         u5_mult_87_ab_52__26_, u5_mult_87_ab_52__27_, u5_mult_87_ab_52__28_,
         u5_mult_87_ab_52__29_, u5_mult_87_ab_52__30_, u5_mult_87_ab_52__31_,
         u5_mult_87_ab_52__32_, u5_mult_87_ab_52__33_, u5_mult_87_ab_52__34_,
         u5_mult_87_ab_52__35_, u5_mult_87_ab_52__36_, u5_mult_87_ab_52__37_,
         u5_mult_87_ab_52__38_, u5_mult_87_ab_52__39_, u5_mult_87_ab_52__40_,
         u5_mult_87_ab_52__41_, u5_mult_87_ab_52__42_, u5_mult_87_ab_52__43_,
         u5_mult_87_ab_52__44_, u5_mult_87_ab_52__45_, u5_mult_87_ab_52__46_,
         u5_mult_87_ab_52__47_, u5_mult_87_ab_52__48_, u5_mult_87_ab_52__49_,
         u5_mult_87_ab_52__50_, u5_mult_87_ab_52__51_, u5_mult_87_ab_52__52_,
         u5_mult_87_FS_1_n331, u5_mult_87_FS_1_n330, u5_mult_87_FS_1_n329,
         u5_mult_87_FS_1_n328, u5_mult_87_FS_1_n327, u5_mult_87_FS_1_n326,
         u5_mult_87_FS_1_n325, u5_mult_87_FS_1_n324, u5_mult_87_FS_1_n323,
         u5_mult_87_FS_1_n322, u5_mult_87_FS_1_n321, u5_mult_87_FS_1_n320,
         u5_mult_87_FS_1_n319, u5_mult_87_FS_1_n318, u5_mult_87_FS_1_n317,
         u5_mult_87_FS_1_n316, u5_mult_87_FS_1_n315, u5_mult_87_FS_1_n314,
         u5_mult_87_FS_1_n313, u5_mult_87_FS_1_n312, u5_mult_87_FS_1_n311,
         u5_mult_87_FS_1_n310, u5_mult_87_FS_1_n309, u5_mult_87_FS_1_n308,
         u5_mult_87_FS_1_n307, u5_mult_87_FS_1_n306, u5_mult_87_FS_1_n305,
         u5_mult_87_FS_1_n304, u5_mult_87_FS_1_n303, u5_mult_87_FS_1_n302,
         u5_mult_87_FS_1_n301, u5_mult_87_FS_1_n300, u5_mult_87_FS_1_n299,
         u5_mult_87_FS_1_n298, u5_mult_87_FS_1_n297, u5_mult_87_FS_1_n296,
         u5_mult_87_FS_1_n295, u5_mult_87_FS_1_n294, u5_mult_87_FS_1_n293,
         u5_mult_87_FS_1_n292, u5_mult_87_FS_1_n291, u5_mult_87_FS_1_n290,
         u5_mult_87_FS_1_n289, u5_mult_87_FS_1_n288, u5_mult_87_FS_1_n287,
         u5_mult_87_FS_1_n286, u5_mult_87_FS_1_n285, u5_mult_87_FS_1_n284,
         u5_mult_87_FS_1_n283, u5_mult_87_FS_1_n282, u5_mult_87_FS_1_n281,
         u5_mult_87_FS_1_n280, u5_mult_87_FS_1_n279, u5_mult_87_FS_1_n278,
         u5_mult_87_FS_1_n277, u5_mult_87_FS_1_n276, u5_mult_87_FS_1_n275,
         u5_mult_87_FS_1_n274, u5_mult_87_FS_1_n273, u5_mult_87_FS_1_n272,
         u5_mult_87_FS_1_n271, u5_mult_87_FS_1_n270, u5_mult_87_FS_1_n269,
         u5_mult_87_FS_1_n268, u5_mult_87_FS_1_n267, u5_mult_87_FS_1_n266,
         u5_mult_87_FS_1_n265, u5_mult_87_FS_1_n264, u5_mult_87_FS_1_n263,
         u5_mult_87_FS_1_n262, u5_mult_87_FS_1_n261, u5_mult_87_FS_1_n260,
         u5_mult_87_FS_1_n259, u5_mult_87_FS_1_n258, u5_mult_87_FS_1_n257,
         u5_mult_87_FS_1_n256, u5_mult_87_FS_1_n255, u5_mult_87_FS_1_n254,
         u5_mult_87_FS_1_n253, u5_mult_87_FS_1_n252, u5_mult_87_FS_1_n251,
         u5_mult_87_FS_1_n250, u5_mult_87_FS_1_n249, u5_mult_87_FS_1_n248,
         u5_mult_87_FS_1_n247, u5_mult_87_FS_1_n246, u5_mult_87_FS_1_n245,
         u5_mult_87_FS_1_n244, u5_mult_87_FS_1_n243, u5_mult_87_FS_1_n242,
         u5_mult_87_FS_1_n241, u5_mult_87_FS_1_n240, u5_mult_87_FS_1_n239,
         u5_mult_87_FS_1_n238, u5_mult_87_FS_1_n237, u5_mult_87_FS_1_n236,
         u5_mult_87_FS_1_n235, u5_mult_87_FS_1_n234, u5_mult_87_FS_1_n233,
         u5_mult_87_FS_1_n232, u5_mult_87_FS_1_n231, u5_mult_87_FS_1_n230,
         u5_mult_87_FS_1_n229, u5_mult_87_FS_1_n228, u5_mult_87_FS_1_n227,
         u5_mult_87_FS_1_n226, u5_mult_87_FS_1_n225, u5_mult_87_FS_1_n224,
         u5_mult_87_FS_1_n223, u5_mult_87_FS_1_n222, u5_mult_87_FS_1_n221,
         u5_mult_87_FS_1_n220, u5_mult_87_FS_1_n219, u5_mult_87_FS_1_n218,
         u5_mult_87_FS_1_n217, u5_mult_87_FS_1_n216, u5_mult_87_FS_1_n215,
         u5_mult_87_FS_1_n214, u5_mult_87_FS_1_n213, u5_mult_87_FS_1_n212,
         u5_mult_87_FS_1_n211, u5_mult_87_FS_1_n210, u5_mult_87_FS_1_n209,
         u5_mult_87_FS_1_n208, u5_mult_87_FS_1_n207, u5_mult_87_FS_1_n206,
         u5_mult_87_FS_1_n205, u5_mult_87_FS_1_n204, u5_mult_87_FS_1_n203,
         u5_mult_87_FS_1_n202, u5_mult_87_FS_1_n201, u5_mult_87_FS_1_n200,
         u5_mult_87_FS_1_n199, u5_mult_87_FS_1_n198, u5_mult_87_FS_1_n197,
         u5_mult_87_FS_1_n196, u5_mult_87_FS_1_n195, u5_mult_87_FS_1_n194,
         u5_mult_87_FS_1_n193, u5_mult_87_FS_1_n192, u5_mult_87_FS_1_n191,
         u5_mult_87_FS_1_n190, u5_mult_87_FS_1_n189, u5_mult_87_FS_1_n188,
         u5_mult_87_FS_1_n187, u5_mult_87_FS_1_n186, u5_mult_87_FS_1_n185,
         u5_mult_87_FS_1_n184, u5_mult_87_FS_1_n183, u5_mult_87_FS_1_n182,
         u5_mult_87_FS_1_n181, u5_mult_87_FS_1_n180, u5_mult_87_FS_1_n179,
         u5_mult_87_FS_1_n178, u5_mult_87_FS_1_n177, u5_mult_87_FS_1_n176,
         u5_mult_87_FS_1_n175, u5_mult_87_FS_1_n174, u5_mult_87_FS_1_n173,
         u5_mult_87_FS_1_n172, u5_mult_87_FS_1_n171, u5_mult_87_FS_1_n170,
         u5_mult_87_FS_1_n169, u5_mult_87_FS_1_n168, u5_mult_87_FS_1_n167,
         u5_mult_87_FS_1_n166, u5_mult_87_FS_1_n165, u5_mult_87_FS_1_n164,
         u5_mult_87_FS_1_n163, u5_mult_87_FS_1_n162, u5_mult_87_FS_1_n161,
         u5_mult_87_FS_1_n160, u5_mult_87_FS_1_n159, u5_mult_87_FS_1_n158,
         u5_mult_87_FS_1_n157, u5_mult_87_FS_1_n156, u5_mult_87_FS_1_n155,
         u5_mult_87_FS_1_n154, u5_mult_87_FS_1_n153, u5_mult_87_FS_1_n152,
         u5_mult_87_FS_1_n151, u5_mult_87_FS_1_n150, u5_mult_87_FS_1_n149,
         u5_mult_87_FS_1_n148, u5_mult_87_FS_1_n147, u5_mult_87_FS_1_n146,
         u5_mult_87_FS_1_n145, u5_mult_87_FS_1_n144, u5_mult_87_FS_1_n143,
         u5_mult_87_FS_1_n142, u5_mult_87_FS_1_n141, u5_mult_87_FS_1_n140,
         u5_mult_87_FS_1_n139, u5_mult_87_FS_1_n138, u5_mult_87_FS_1_n137,
         u5_mult_87_FS_1_n136, u5_mult_87_FS_1_n135, u5_mult_87_FS_1_n134,
         u5_mult_87_FS_1_n133, u5_mult_87_FS_1_n132, u5_mult_87_FS_1_n131,
         u5_mult_87_FS_1_n130, u5_mult_87_FS_1_n129, u5_mult_87_FS_1_n128,
         u5_mult_87_FS_1_n127, u5_mult_87_FS_1_n126, u5_mult_87_FS_1_n125,
         u5_mult_87_FS_1_n124, u5_mult_87_FS_1_n123, u5_mult_87_FS_1_n122,
         u5_mult_87_FS_1_n121, u5_mult_87_FS_1_n120, u5_mult_87_FS_1_n119,
         u5_mult_87_FS_1_n118, u5_mult_87_FS_1_n117, u5_mult_87_FS_1_n116,
         u5_mult_87_FS_1_n115, u5_mult_87_FS_1_n114, u5_mult_87_FS_1_n113,
         u5_mult_87_FS_1_n112, u5_mult_87_FS_1_n111, u5_mult_87_FS_1_n110,
         u5_mult_87_FS_1_n109, u5_mult_87_FS_1_n108, u5_mult_87_FS_1_n107,
         u5_mult_87_FS_1_n106, u5_mult_87_FS_1_n105, u5_mult_87_FS_1_n104,
         u5_mult_87_FS_1_n103, u5_mult_87_FS_1_n102, u5_mult_87_FS_1_n101,
         u5_mult_87_FS_1_n100, u5_mult_87_FS_1_n99, u5_mult_87_FS_1_n98,
         u5_mult_87_FS_1_n97, u5_mult_87_FS_1_n96, u5_mult_87_FS_1_n95,
         u5_mult_87_FS_1_n94, u5_mult_87_FS_1_n93, u5_mult_87_FS_1_n92,
         u5_mult_87_FS_1_n91, u5_mult_87_FS_1_n90, u5_mult_87_FS_1_n89,
         u5_mult_87_FS_1_n88, u5_mult_87_FS_1_n87, u5_mult_87_FS_1_n86,
         u5_mult_87_FS_1_n85, u5_mult_87_FS_1_n84, u5_mult_87_FS_1_n83,
         u5_mult_87_FS_1_n82, u5_mult_87_FS_1_n81, u5_mult_87_FS_1_n80,
         u5_mult_87_FS_1_n79, u5_mult_87_FS_1_n78, u5_mult_87_FS_1_n77,
         u5_mult_87_FS_1_n76, u5_mult_87_FS_1_n75, u5_mult_87_FS_1_n74,
         u5_mult_87_FS_1_n73, u5_mult_87_FS_1_n72, u5_mult_87_FS_1_n71,
         u5_mult_87_FS_1_n70, u5_mult_87_FS_1_n69, u5_mult_87_FS_1_n68,
         u5_mult_87_FS_1_n67, u5_mult_87_FS_1_n66, u5_mult_87_FS_1_n65,
         u5_mult_87_FS_1_n64, u5_mult_87_FS_1_n63, u5_mult_87_FS_1_n62,
         u5_mult_87_FS_1_n61, u5_mult_87_FS_1_n60, u5_mult_87_FS_1_n59,
         u5_mult_87_FS_1_n58, u5_mult_87_FS_1_n57, u5_mult_87_FS_1_n56,
         u5_mult_87_FS_1_n55, u5_mult_87_FS_1_n54, u5_mult_87_FS_1_n53,
         u5_mult_87_FS_1_n52, u5_mult_87_FS_1_n51, u5_mult_87_FS_1_n50,
         u5_mult_87_FS_1_n49, u5_mult_87_FS_1_n48, u5_mult_87_FS_1_n47,
         u5_mult_87_FS_1_n46, u5_mult_87_FS_1_n45, u5_mult_87_FS_1_n44,
         u5_mult_87_FS_1_n43, u5_mult_87_FS_1_n42, u5_mult_87_FS_1_n41,
         u5_mult_87_FS_1_n40, u5_mult_87_FS_1_n39, u5_mult_87_FS_1_n38,
         u5_mult_87_FS_1_n37, u5_mult_87_FS_1_n36, u5_mult_87_FS_1_n35,
         u5_mult_87_FS_1_n34, u5_mult_87_FS_1_n33, u5_mult_87_FS_1_n32,
         u5_mult_87_FS_1_n31, u5_mult_87_FS_1_n30, u5_mult_87_FS_1_n29,
         u5_mult_87_FS_1_n28, u5_mult_87_FS_1_n27, u5_mult_87_FS_1_n26,
         u5_mult_87_FS_1_n25, u5_mult_87_FS_1_n24, u5_mult_87_FS_1_n23,
         u5_mult_87_FS_1_n22, u5_mult_87_FS_1_n21, u5_mult_87_FS_1_n20,
         u5_mult_87_FS_1_n19, u5_mult_87_FS_1_n18, u5_mult_87_FS_1_n17,
         u5_mult_87_FS_1_n16, u5_mult_87_FS_1_n15, u5_mult_87_FS_1_n14,
         u5_mult_87_FS_1_n13, u5_mult_87_FS_1_n12, u5_mult_87_FS_1_n11,
         u5_mult_87_FS_1_n10, u5_mult_87_FS_1_n9, u5_mult_87_FS_1_n8,
         u5_mult_87_FS_1_n7, u5_mult_87_FS_1_n6, u5_mult_87_FS_1_n5,
         u5_mult_87_FS_1_n4, u5_mult_87_FS_1_n3, u5_mult_87_FS_1_n2;
  wire   [63:52] opa_r;
  wire   [63:52] opb_r;
  wire   [1:0] rmode_r1;
  wire   [1:0] rmode_r2;
  wire   [1:0] rmode_r3;
  wire   [2:0] fpu_op_r1;
  wire   [2:0] fpu_op_r2;
  wire   [2:0] fpu_op_r3;
  wire   [55:0] fracta;
  wire   [55:0] fractb;
  wire   [10:0] exp_fasu;
  wire   [51:0] fracta_mul;
  wire   [10:0] exp_mul;
  wire   [1:0] exp_ovf;
  wire   [2:0] underflow_fmul_d;
  wire   [56:0] fract_out_q;
  wire   [105:0] prod;
  wire   [4:0] div_opa_ldz_d;
  wire   [55:0] quo;
  wire   [107:0] remainder;
  wire   [4:0] div_opa_ldz_r1;
  wire   [4:0] div_opa_ldz_r2;
  wire   [10:2] exp_r;
  wire   [59:1] opa_r1;
  wire   [105:0] fract_i2f;
  wire   [105:0] fract_denorm;
  wire   [2:0] underflow_fmul_r;
  wire   [55:0] u1_fractb_s;
  wire   [55:0] u1_fracta_s;
  wire   [10:0] u1_exp_diff2;
  wire   [10:0] u1_exp_small;
  wire   [2:0] u2_underflow_d;
  wire   [105:0] u5_prod1;
  wire   [107:0] u6_remainder;
  wire   [107:0] u6_quo1;
  wire   [10:0] u4_div_exp3;
  wire   [117:107] u4_exp_f2i_1;
  wire   [10:0] u4_exp_fix_divb;
  wire   [10:0] u4_exp_fix_diva;
  wire   [10:0] u4_exp_out1_mi1;
  wire   [10:0] u4_exp_out_mi1;
  wire   [6:1] u4_fi_ldz_mi22;
  wire   [8:0] u4_shift_left;
  wire   [10:0] u4_shift_right;
  wire   [10:0] u4_div_shft4;
  wire   [10:2] u4_div_shft2;
  wire   [10:0] u4_div_scht1a;
  wire   [6:2] u4_sub_479_carry;
  wire   [10:1] u4_sub_410_carry;
  wire   [10:1] u4_add_409_carry;
  wire   [10:3] u4_add_408_carry;
  wire   [10:1] u4_sub_407_carry;
  wire   [6:2] u4_sub_489_carry;
  wire   [7:1] sub_1_root_sub_0_root_u4_add_495_carry;
  wire   [10:2] u4_add_462_carry;
  wire   [6:5] u4_sll_480_SHMAG;
  wire   [10:2] u4_add_464_carry;
  wire   [51:2] u4_add_394_carry;
  wire   [56:1] u3_sub_61_carry;
  wire   [55:2] u3_add_61_carry;
  wire   [10:2] u2_add_116_carry;
  wire   [10:2] u2_add_114_carry;
  wire   [10:2] u2_add_111_carry;
  wire   [11:1] u2_sub_111_carry;
  wire   [10:1] sub_1_root_u1_sub_130_aco_carry;
  wire   [10:2] add_0_root_sub_0_root_u4_add_495_carry;

  OR2_X2 u4_C19002 ( .A1(u4_N6439), .A2(u4_exp_out_0_), .ZN(u4_N6440) );
  OR2_X2 u4_C19003 ( .A1(u4_N6438), .A2(u4_exp_out_1_), .ZN(u4_N6439) );
  OR2_X2 u4_C19004 ( .A1(u4_N6437), .A2(u4_exp_out_2_), .ZN(u4_N6438) );
  OR2_X2 u4_C19005 ( .A1(u4_N6436), .A2(u4_exp_out_3_), .ZN(u4_N6437) );
  OR2_X2 u4_C19006 ( .A1(u4_N6435), .A2(u4_exp_out_4_), .ZN(u4_N6436) );
  OR2_X2 u4_C19007 ( .A1(u4_N6434), .A2(u4_exp_out_5_), .ZN(u4_N6435) );
  OR2_X2 u4_C19008 ( .A1(u4_N6433), .A2(u4_exp_out_6_), .ZN(u4_N6434) );
  OR2_X2 u4_C19009 ( .A1(u4_N6432), .A2(u4_exp_out_7_), .ZN(u4_N6433) );
  OR2_X2 u4_C19010 ( .A1(u4_N6431), .A2(u4_exp_out_8_), .ZN(u4_N6432) );
  OR2_X2 u4_C19011 ( .A1(u4_exp_out_10_), .A2(u4_exp_out_9_), .ZN(u4_N6431) );
  OR2_X2 u4_C19431 ( .A1(u4_shift_right[10]), .A2(u4_shift_right[9]), .ZN(
        u4_N5898) );
  OR2_X2 u4_C19692 ( .A1(u4_N6891), .A2(u4_N6892), .ZN(u4_N6893) );
  AND2_X2 u4_C19694 ( .A1(u4_exp_out_10_), .A2(1'b1), .ZN(u4_N6892) );
  OAI33_X1 U122 ( .A1(n6526), .A2(n279), .A3(n4819), .B1(n281), .B2(n282), 
        .B3(n283), .ZN(n277) );
  OAI33_X1 U180 ( .A1(n418), .A2(fract_denorm[104]), .A3(fract_denorm[103]), 
        .B1(n6468), .B2(fract_denorm[55]), .B3(n419), .ZN(n417) );
  OAI33_X1 U189 ( .A1(n6493), .A2(fract_denorm[79]), .A3(n351), .B1(n6476), 
        .B2(fract_denorm[63]), .B3(n310), .ZN(n433) );
  OAI33_X1 U196 ( .A1(n6450), .A2(fract_denorm[41]), .A3(n443), .B1(n6435), 
        .B2(fract_denorm[25]), .B3(n331), .ZN(n441) );
  OAI33_X1 U201 ( .A1(n6516), .A2(fract_denorm[102]), .A3(fract_denorm[101]), 
        .B1(n6486), .B2(fract_denorm[73]), .B3(n6488), .ZN(n450) );
  OAI33_X1 U209 ( .A1(n6442), .A2(fract_denorm[33]), .A3(n461), .B1(n462), 
        .B2(n387), .B3(n6426), .ZN(n459) );
  OAI33_X1 U240 ( .A1(n6501), .A2(fract_denorm[86]), .A3(n6503), .B1(n6482), 
        .B2(fract_denorm[70]), .B3(n6485), .ZN(n497) );
  OAI33_X1 U244 ( .A1(n6431), .A2(fract_denorm[22]), .A3(n420), .B1(n6410), 
        .B2(n6411), .B3(n504), .ZN(n491) );
  OAI33_X1 U262 ( .A1(n6489), .A2(fract_denorm[76]), .A3(n312), .B1(n6473), 
        .B2(fract_denorm[60]), .B3(n376), .ZN(n519) );
  OAI33_X1 U311 ( .A1(n6496), .A2(fract_denorm[82]), .A3(n400), .B1(n6512), 
        .B2(fract_denorm[98]), .B3(n394), .ZN(n568) );
  OAI33_X1 U318 ( .A1(n6445), .A2(fract_denorm[36]), .A3(n6446), .B1(n6415), 
        .B2(fract_denorm[10]), .B3(n296), .ZN(n573) );
  OAI33_X1 U1654 ( .A1(n6363), .A2(fracta_mul[43]), .A3(n4375), .B1(n6361), 
        .B2(fracta_mul[35]), .B3(n1395), .ZN(n1409) );
  OAI33_X1 U1710 ( .A1(n6363), .A2(n1284), .A3(n4618), .B1(n1449), .B2(n6371), 
        .B3(n1450), .ZN(n1448) );
  OAI33_X1 U1780 ( .A1(n1470), .A2(opb_inf), .A3(n1471), .B1(n1472), .B2(n1473), .B3(n4432), .ZN(n1469) );
  OAI33_X1 U1798 ( .A1(n1517), .A2(n1518), .A3(n1519), .B1(n1480), .B2(
        inf_mul_r), .B3(n1520), .ZN(N907) );
  OAI33_X1 U2227 ( .A1(n1974), .A2(r482_B_0_), .A3(n4821), .B1(n4427), .B2(
        sign), .B3(n1975), .ZN(n1681) );
  DFF_X2 opa_r_reg_63_ ( .D(opa[63]), .CK(clk), .Q(opa_r[63]), .QN(n4666) );
  DFF_X2 opa_r_reg_62_ ( .D(opa[62]), .CK(clk), .Q(opa_r[62]), .QN(n4592) );
  DFF_X2 opa_r_reg_61_ ( .D(opa[61]), .CK(clk), .Q(opa_r[61]), .QN(n4482) );
  DFF_X2 opa_r_reg_60_ ( .D(opa[60]), .CK(clk), .Q(opa_r[60]), .QN(n4580) );
  DFF_X2 opa_r_reg_59_ ( .D(opa[59]), .CK(clk), .Q(opa_r[59]), .QN(n4582) );
  DFF_X2 opa_r_reg_58_ ( .D(opa[58]), .CK(clk), .Q(opa_r[58]), .QN(n4575) );
  DFF_X2 opa_r_reg_57_ ( .D(opa[57]), .CK(clk), .Q(opa_r[57]), .QN(n4586) );
  DFF_X2 opa_r_reg_56_ ( .D(opa[56]), .CK(clk), .Q(opa_r[56]), .QN(n4589) );
  DFF_X2 opa_r_reg_55_ ( .D(opa[55]), .CK(clk), .Q(opa_r[55]), .QN(n4485) );
  DFF_X2 opa_r_reg_54_ ( .D(opa[54]), .CK(clk), .Q(opa_r[54]), .QN(n4583) );
  DFF_X2 opa_r_reg_53_ ( .D(opa[53]), .CK(clk), .Q(opa_r[53]), .QN(n4584) );
  DFF_X2 opa_r_reg_52_ ( .D(opa[52]), .CK(clk), .Q(opa_r[52]), .QN(n4585) );
  DFF_X2 opa_r_reg_51_ ( .D(opa[51]), .CK(clk), .Q(fracta_mul[51]), .QN(n4354)
         );
  DFF_X2 opa_r_reg_50_ ( .D(opa[50]), .CK(clk), .Q(fracta_mul[50]), .QN(n4352)
         );
  DFF_X2 opa_r_reg_49_ ( .D(opa[49]), .CK(clk), .Q(fracta_mul[49]), .QN(n4355)
         );
  DFF_X2 opa_r_reg_48_ ( .D(opa[48]), .CK(clk), .Q(fracta_mul[48]), .QN(n4366)
         );
  DFF_X2 opa_r_reg_47_ ( .D(opa[47]), .CK(clk), .Q(fracta_mul[47]), .QN(n4362)
         );
  DFF_X2 opa_r_reg_46_ ( .D(opa[46]), .CK(clk), .Q(fracta_mul[46]) );
  DFF_X2 opa_r_reg_45_ ( .D(opa[45]), .CK(clk), .Q(fracta_mul[45]), .QN(n4499)
         );
  DFF_X2 opa_r_reg_44_ ( .D(opa[44]), .CK(clk), .Q(fracta_mul[44]), .QN(n4611)
         );
  DFF_X2 opa_r_reg_43_ ( .D(opa[43]), .CK(clk), .Q(fracta_mul[43]) );
  DFF_X2 opa_r_reg_42_ ( .D(opa[42]), .CK(clk), .Q(fracta_mul[42]), .QN(n4375)
         );
  DFF_X2 opa_r_reg_41_ ( .D(opa[41]), .CK(clk), .Q(fracta_mul[41]), .QN(n4617)
         );
  DFF_X2 opa_r_reg_40_ ( .D(opa[40]), .CK(clk), .Q(fracta_mul[40]) );
  DFF_X2 opa_r_reg_39_ ( .D(opa[39]), .CK(clk), .Q(fracta_mul[39]), .QN(n4618)
         );
  DFF_X2 opa_r_reg_38_ ( .D(opa[38]), .CK(clk), .Q(fracta_mul[38]), .QN(n4374)
         );
  DFF_X2 opa_r_reg_37_ ( .D(opa[37]), .CK(clk), .Q(fracta_mul[37]) );
  DFF_X2 opa_r_reg_36_ ( .D(opa[36]), .CK(clk), .Q(fracta_mul[36]), .QN(n4365)
         );
  DFF_X2 opa_r_reg_35_ ( .D(opa[35]), .CK(clk), .Q(fracta_mul[35]), .QN(n4614)
         );
  DFF_X2 opa_r_reg_34_ ( .D(opa[34]), .CK(clk), .Q(fracta_mul[34]), .QN(n4613)
         );
  DFF_X2 opa_r_reg_33_ ( .D(opa[33]), .CK(clk), .Q(fracta_mul[33]) );
  DFF_X2 opa_r_reg_32_ ( .D(opa[32]), .CK(clk), .Q(fracta_mul[32]), .QN(n4372)
         );
  DFF_X2 opa_r_reg_31_ ( .D(opa[31]), .CK(clk), .Q(fracta_mul[31]) );
  DFF_X2 opa_r_reg_30_ ( .D(opa[30]), .CK(clk), .Q(fracta_mul[30]), .QN(n4612)
         );
  DFF_X2 opa_r_reg_29_ ( .D(opa[29]), .CK(clk), .Q(fracta_mul[29]), .QN(n4373)
         );
  DFF_X2 opa_r_reg_28_ ( .D(opa[28]), .CK(clk), .Q(fracta_mul[28]), .QN(n4363)
         );
  DFF_X2 opa_r_reg_27_ ( .D(opa[27]), .CK(clk), .Q(fracta_mul[27]), .QN(n4364)
         );
  DFF_X2 opa_r_reg_26_ ( .D(opa[26]), .CK(clk), .Q(fracta_mul[26]), .QN(n4615)
         );
  DFF_X2 opa_r_reg_25_ ( .D(opa[25]), .CK(clk), .Q(fracta_mul[25]), .QN(n4376)
         );
  DFF_X2 opa_r_reg_24_ ( .D(opa[24]), .CK(clk), .Q(fracta_mul[24]) );
  DFF_X2 opa_r_reg_23_ ( .D(opa[23]), .CK(clk), .Q(fracta_mul[23]), .QN(n4356)
         );
  DFF_X2 opa_r_reg_22_ ( .D(opa[22]), .CK(clk), .Q(fracta_mul[22]), .QN(n4367)
         );
  DFF_X2 opa_r_reg_21_ ( .D(opa[21]), .CK(clk), .Q(fracta_mul[21]), .QN(n4377)
         );
  DFF_X2 opa_r_reg_20_ ( .D(opa[20]), .CK(clk), .Q(fracta_mul[20]) );
  DFF_X2 opa_r_reg_19_ ( .D(opa[19]), .CK(clk), .Q(fracta_mul[19]) );
  DFF_X2 opa_r_reg_18_ ( .D(opa[18]), .CK(clk), .Q(fracta_mul[18]), .QN(n4616)
         );
  DFF_X2 opa_r_reg_17_ ( .D(opa[17]), .CK(clk), .Q(fracta_mul[17]), .QN(n4488)
         );
  DFF_X2 opa_r_reg_16_ ( .D(opa[16]), .CK(clk), .Q(fracta_mul[16]), .QN(n4489)
         );
  DFF_X2 opa_r_reg_15_ ( .D(opa[15]), .CK(clk), .Q(fracta_mul[15]) );
  DFF_X2 opa_r_reg_14_ ( .D(opa[14]), .CK(clk), .Q(fracta_mul[14]), .QN(n4496)
         );
  DFF_X2 opa_r_reg_13_ ( .D(opa[13]), .CK(clk), .Q(fracta_mul[13]) );
  DFF_X2 opa_r_reg_12_ ( .D(opa[12]), .CK(clk), .Q(fracta_mul[12]), .QN(n4491)
         );
  DFF_X2 opa_r_reg_11_ ( .D(opa[11]), .CK(clk), .Q(fracta_mul[11]), .QN(n4495)
         );
  DFF_X2 opa_r_reg_10_ ( .D(opa[10]), .CK(clk), .Q(fracta_mul[10]) );
  DFF_X2 opa_r_reg_9_ ( .D(opa[9]), .CK(clk), .Q(fracta_mul[9]), .QN(n4492) );
  DFF_X2 opa_r_reg_8_ ( .D(opa[8]), .CK(clk), .Q(fracta_mul[8]) );
  DFF_X2 opa_r_reg_7_ ( .D(opa[7]), .CK(clk), .Q(fracta_mul[7]) );
  DFF_X2 opa_r_reg_6_ ( .D(opa[6]), .CK(clk), .Q(fracta_mul[6]) );
  DFF_X2 opa_r_reg_5_ ( .D(opa[5]), .CK(clk), .Q(fracta_mul[5]), .QN(n4498) );
  DFF_X2 opa_r_reg_4_ ( .D(opa[4]), .CK(clk), .Q(fracta_mul[4]) );
  DFF_X2 opa_r_reg_3_ ( .D(opa[3]), .CK(clk), .Q(fracta_mul[3]), .QN(n4500) );
  DFF_X2 opa_r_reg_2_ ( .D(opa[2]), .CK(clk), .Q(fracta_mul[2]) );
  DFF_X2 opa_r_reg_1_ ( .D(opa[1]), .CK(clk), .Q(fracta_mul[1]), .QN(n4497) );
  DFF_X2 opa_r_reg_0_ ( .D(opa[0]), .CK(clk), .Q(fracta_mul[0]) );
  DFF_X2 opb_r_reg_63_ ( .D(opb[63]), .CK(clk), .Q(opb_r[63]) );
  DFF_X2 opb_r_reg_62_ ( .D(opb[62]), .CK(clk), .Q(opb_r[62]), .QN(n4487) );
  DFF_X2 opb_r_reg_61_ ( .D(opb[61]), .CK(clk), .Q(opb_r[61]) );
  DFF_X2 opb_r_reg_60_ ( .D(opb[60]), .CK(clk), .Q(opb_r[60]) );
  DFF_X2 opb_r_reg_59_ ( .D(opb[59]), .CK(clk), .Q(opb_r[59]), .QN(n4569) );
  DFF_X2 opb_r_reg_58_ ( .D(opb[58]), .CK(clk), .Q(opb_r[58]), .QN(n4471) );
  DFF_X2 opb_r_reg_57_ ( .D(opb[57]), .CK(clk), .Q(opb_r[57]), .QN(n4398) );
  DFF_X2 opb_r_reg_56_ ( .D(opb[56]), .CK(clk), .Q(opb_r[56]), .QN(n4486) );
  DFF_X2 opb_r_reg_55_ ( .D(opb[55]), .CK(clk), .Q(opb_r[55]), .QN(n4591) );
  DFF_X2 opb_r_reg_54_ ( .D(opb[54]), .CK(clk), .Q(opb_r[54]), .QN(n4590) );
  DFF_X2 opb_r_reg_53_ ( .D(opb[53]), .CK(clk), .Q(opb_r[53]), .QN(n4360) );
  DFF_X2 opb_r_reg_52_ ( .D(opb[52]), .CK(clk), .Q(opb_r[52]), .QN(n4371) );
  DFF_X2 opb_r_reg_51_ ( .D(opb[51]), .CK(clk), .Q(u6_N51), .QN(n4594) );
  DFF_X2 opb_r_reg_50_ ( .D(opb[50]), .CK(clk), .Q(u6_N50), .QN(n4597) );
  DFF_X2 opb_r_reg_49_ ( .D(opb[49]), .CK(clk), .Q(u6_N49), .QN(n4490) );
  DFF_X2 opb_r_reg_48_ ( .D(opb[48]), .CK(clk), .Q(u6_N48), .QN(n4431) );
  DFF_X2 opb_r_reg_47_ ( .D(opb[47]), .CK(clk), .Q(u6_N47), .QN(n4593) );
  DFF_X2 opb_r_reg_46_ ( .D(opb[46]), .CK(clk), .Q(u6_N46) );
  DFF_X2 opb_r_reg_45_ ( .D(opb[45]), .CK(clk), .Q(u6_N45) );
  DFF_X2 opb_r_reg_44_ ( .D(opb[44]), .CK(clk), .Q(u6_N44) );
  DFF_X2 opb_r_reg_43_ ( .D(opb[43]), .CK(clk), .Q(u6_N43) );
  DFF_X2 opb_r_reg_42_ ( .D(opb[42]), .CK(clk), .Q(u6_N42), .QN(n4600) );
  DFF_X2 opb_r_reg_41_ ( .D(opb[41]), .CK(clk), .Q(u6_N41) );
  DFF_X2 opb_r_reg_40_ ( .D(opb[40]), .CK(clk), .Q(u6_N40) );
  DFF_X2 opb_r_reg_39_ ( .D(opb[39]), .CK(clk), .Q(u6_N39) );
  DFF_X2 opb_r_reg_38_ ( .D(opb[38]), .CK(clk), .Q(u6_N38), .QN(n4596) );
  DFF_X2 opb_r_reg_37_ ( .D(opb[37]), .CK(clk), .Q(u6_N37) );
  DFF_X2 opb_r_reg_36_ ( .D(opb[36]), .CK(clk), .Q(u6_N36), .QN(n4604) );
  DFF_X2 opb_r_reg_35_ ( .D(opb[35]), .CK(clk), .Q(u6_N35) );
  DFF_X2 opb_r_reg_34_ ( .D(opb[34]), .CK(clk), .Q(u6_N34) );
  DFF_X2 opb_r_reg_33_ ( .D(opb[33]), .CK(clk), .Q(u6_N33) );
  DFF_X2 opb_r_reg_32_ ( .D(opb[32]), .CK(clk), .Q(u6_N32), .QN(n4595) );
  DFF_X2 opb_r_reg_31_ ( .D(opb[31]), .CK(clk), .Q(u6_N31) );
  DFF_X2 opb_r_reg_30_ ( .D(opb[30]), .CK(clk), .Q(u6_N30) );
  DFF_X2 opb_r_reg_29_ ( .D(opb[29]), .CK(clk), .Q(u6_N29), .QN(n4599) );
  DFF_X2 opb_r_reg_28_ ( .D(opb[28]), .CK(clk), .Q(u6_N28), .QN(n4603) );
  DFF_X2 opb_r_reg_27_ ( .D(opb[27]), .CK(clk), .Q(u6_N27), .QN(n4607) );
  DFF_X2 opb_r_reg_26_ ( .D(opb[26]), .CK(clk), .Q(u6_N26) );
  DFF_X2 opb_r_reg_25_ ( .D(opb[25]), .CK(clk), .Q(u6_N25), .QN(n4605) );
  DFF_X2 opb_r_reg_24_ ( .D(opb[24]), .CK(clk), .Q(u6_N24) );
  DFF_X2 opb_r_reg_23_ ( .D(opb[23]), .CK(clk), .Q(u6_N23), .QN(n4610) );
  DFF_X2 opb_r_reg_22_ ( .D(opb[22]), .CK(clk), .Q(u6_N22), .QN(n4602) );
  DFF_X2 opb_r_reg_21_ ( .D(opb[21]), .CK(clk), .Q(u6_N21), .QN(n4606) );
  DFF_X2 opb_r_reg_20_ ( .D(opb[20]), .CK(clk), .Q(u6_N20) );
  DFF_X2 opb_r_reg_19_ ( .D(opb[19]), .CK(clk), .Q(u6_N19) );
  DFF_X2 opb_r_reg_18_ ( .D(opb[18]), .CK(clk), .Q(u6_N18) );
  DFF_X2 opb_r_reg_17_ ( .D(opb[17]), .CK(clk), .Q(u6_N17), .QN(n4601) );
  DFF_X2 opb_r_reg_16_ ( .D(opb[16]), .CK(clk), .Q(u6_N16), .QN(n4598) );
  DFF_X2 opb_r_reg_15_ ( .D(opb[15]), .CK(clk), .Q(u6_N15) );
  DFF_X2 opb_r_reg_14_ ( .D(opb[14]), .CK(clk), .Q(u6_N14) );
  DFF_X2 opb_r_reg_13_ ( .D(opb[13]), .CK(clk), .Q(u6_N13) );
  DFF_X2 opb_r_reg_12_ ( .D(opb[12]), .CK(clk), .Q(u6_N12), .QN(n4609) );
  DFF_X2 opb_r_reg_11_ ( .D(opb[11]), .CK(clk), .Q(u6_N11) );
  DFF_X2 opb_r_reg_10_ ( .D(opb[10]), .CK(clk), .Q(u6_N10) );
  DFF_X2 opb_r_reg_9_ ( .D(opb[9]), .CK(clk), .Q(u6_N9), .QN(n4608) );
  DFF_X2 opb_r_reg_8_ ( .D(opb[8]), .CK(clk), .Q(u6_N8) );
  DFF_X2 opb_r_reg_7_ ( .D(opb[7]), .CK(clk), .Q(u6_N7) );
  DFF_X2 opb_r_reg_6_ ( .D(opb[6]), .CK(clk), .Q(u6_N6) );
  DFF_X2 opb_r_reg_5_ ( .D(opb[5]), .CK(clk), .Q(u6_N5) );
  DFF_X2 opb_r_reg_4_ ( .D(opb[4]), .CK(clk), .Q(u6_N4) );
  DFF_X2 opb_r_reg_3_ ( .D(opb[3]), .CK(clk), .Q(u6_N3) );
  DFF_X2 opb_r_reg_2_ ( .D(opb[2]), .CK(clk), .Q(u6_N2) );
  DFF_X2 opb_r_reg_1_ ( .D(opb[1]), .CK(clk), .Q(u6_N1) );
  DFF_X2 opb_r_reg_0_ ( .D(opb[0]), .CK(clk), .Q(u6_N0) );
  DFF_X2 rmode_r1_reg_1_ ( .D(rmode[1]), .CK(clk), .Q(rmode_r1[1]) );
  DFF_X2 rmode_r1_reg_0_ ( .D(rmode[0]), .CK(clk), .Q(rmode_r1[0]) );
  DFF_X2 rmode_r2_reg_1_ ( .D(rmode_r1[1]), .CK(clk), .Q(rmode_r2[1]) );
  DFF_X2 rmode_r2_reg_0_ ( .D(rmode_r1[0]), .CK(clk), .Q(rmode_r2[0]) );
  DFF_X2 rmode_r3_reg_1_ ( .D(rmode_r2[1]), .CK(clk), .Q(rmode_r3[1]), .QN(
        n4427) );
  DFF_X2 rmode_r3_reg_0_ ( .D(rmode_r2[0]), .CK(clk), .Q(rmode_r3[0]), .QN(
        n4483) );
  DFF_X2 fpu_op_r1_reg_2_ ( .D(fpu_op[2]), .CK(clk), .Q(fpu_op_r1[2]), .QN(
        n4501) );
  DFF_X2 fpu_op_r1_reg_1_ ( .D(fpu_op[1]), .CK(clk), .Q(fpu_op_r1[1]) );
  DFF_X2 fpu_op_r1_reg_0_ ( .D(fpu_op[0]), .CK(clk), .Q(fpu_op_r1[0]), .QN(
        n4620) );
  DFF_X2 fpu_op_r2_reg_2_ ( .D(fpu_op_r1[2]), .CK(clk), .Q(fpu_op_r2[2]) );
  DFF_X2 fpu_op_r2_reg_1_ ( .D(fpu_op_r1[1]), .CK(clk), .Q(fpu_op_r2[1]), .QN(
        n4505) );
  DFF_X2 fpu_op_r2_reg_0_ ( .D(fpu_op_r1[0]), .CK(clk), .Q(fpu_op_r2[0]), .QN(
        n4634) );
  DFF_X2 fpu_op_r3_reg_2_ ( .D(fpu_op_r2[2]), .CK(clk), .Q(fpu_op_r3[2]), .QN(
        n4351) );
  DFF_X2 fpu_op_r3_reg_1_ ( .D(fpu_op_r2[1]), .CK(clk), .Q(fpu_op_r3[1]), .QN(
        n4353) );
  DFF_X2 fpu_op_r3_reg_0_ ( .D(fpu_op_r2[0]), .CK(clk), .Q(fpu_op_r3[0]), .QN(
        n4481) );
  DFF_X2 div_opa_ldz_r1_reg_4_ ( .D(div_opa_ldz_d[4]), .CK(clk), .Q(
        div_opa_ldz_r1[4]) );
  DFF_X2 div_opa_ldz_r1_reg_3_ ( .D(div_opa_ldz_d[3]), .CK(clk), .Q(
        div_opa_ldz_r1[3]) );
  DFF_X2 div_opa_ldz_r1_reg_2_ ( .D(div_opa_ldz_d[2]), .CK(clk), .Q(
        div_opa_ldz_r1[2]) );
  DFF_X2 div_opa_ldz_r1_reg_1_ ( .D(div_opa_ldz_d[1]), .CK(clk), .Q(
        div_opa_ldz_r1[1]) );
  DFF_X2 div_opa_ldz_r1_reg_0_ ( .D(div_opa_ldz_d[0]), .CK(clk), .Q(
        div_opa_ldz_r1[0]) );
  DFF_X2 div_opa_ldz_r2_reg_4_ ( .D(div_opa_ldz_r1[4]), .CK(clk), .Q(
        div_opa_ldz_r2[4]), .QN(n4581) );
  DFF_X2 div_opa_ldz_r2_reg_3_ ( .D(div_opa_ldz_r1[3]), .CK(clk), .Q(
        div_opa_ldz_r2[3]), .QN(n4576) );
  DFF_X2 div_opa_ldz_r2_reg_2_ ( .D(div_opa_ldz_r1[2]), .CK(clk), .Q(
        div_opa_ldz_r2[2]), .QN(n4577) );
  DFF_X2 div_opa_ldz_r2_reg_1_ ( .D(div_opa_ldz_r1[1]), .CK(clk), .Q(
        div_opa_ldz_r2[1]), .QN(n4578) );
  DFF_X2 div_opa_ldz_r2_reg_0_ ( .D(div_opa_ldz_r1[0]), .CK(clk), .Q(
        div_opa_ldz_r2[0]), .QN(n4570) );
  DFF_X2 opa_r1_reg_62_ ( .D(opa_r[62]), .CK(clk), .QN(n4508) );
  DFF_X2 opa_r1_reg_61_ ( .D(opa_r[61]), .CK(clk), .QN(n4623) );
  DFF_X2 opa_r1_reg_60_ ( .D(opa_r[60]), .CK(clk), .QN(n4433) );
  DFF_X2 opa_r1_reg_59_ ( .D(opa_r[59]), .CK(clk), .Q(opa_r1[59]), .QN(n4629)
         );
  DFF_X2 opa_r1_reg_58_ ( .D(opa_r[58]), .CK(clk), .Q(opa_r1[58]), .QN(n4410)
         );
  DFF_X2 opa_r1_reg_57_ ( .D(opa_r[57]), .CK(clk), .Q(opa_r1[57]), .QN(n4409)
         );
  DFF_X2 opa_r1_reg_56_ ( .D(opa_r[56]), .CK(clk), .Q(opa_r1[56]), .QN(n4408)
         );
  DFF_X2 opa_r1_reg_55_ ( .D(opa_r[55]), .CK(clk), .Q(opa_r1[55]), .QN(n4407)
         );
  DFF_X2 opa_r1_reg_54_ ( .D(opa_r[54]), .CK(clk), .Q(opa_r1[54]), .QN(n4625)
         );
  DFF_X2 opa_r1_reg_53_ ( .D(opa_r[53]), .CK(clk), .Q(opa_r1[53]), .QN(n4622)
         );
  DFF_X2 opa_r1_reg_52_ ( .D(opa_r[52]), .CK(clk), .Q(opa_r1[52]), .QN(n4509)
         );
  DFF_X2 opa_r1_reg_51_ ( .D(fracta_mul[51]), .CK(clk), .Q(opa_r1[51]), .QN(
        n4419) );
  DFF_X2 opa_r1_reg_50_ ( .D(fracta_mul[50]), .CK(clk), .Q(opa_r1[50]), .QN(
        n4418) );
  DFF_X2 opa_r1_reg_49_ ( .D(fracta_mul[49]), .CK(clk), .Q(opa_r1[49]), .QN(
        n4417) );
  DFF_X2 opa_r1_reg_48_ ( .D(fracta_mul[48]), .CK(clk), .Q(opa_r1[48]), .QN(
        n4450) );
  DFF_X2 opa_r1_reg_47_ ( .D(fracta_mul[47]), .CK(clk), .Q(opa_r1[47]), .QN(
        n4449) );
  DFF_X2 opa_r1_reg_46_ ( .D(fracta_mul[46]), .CK(clk), .Q(opa_r1[46]), .QN(
        n4448) );
  DFF_X2 opa_r1_reg_45_ ( .D(fracta_mul[45]), .CK(clk), .Q(opa_r1[45]), .QN(
        n4665) );
  DFF_X2 opa_r1_reg_44_ ( .D(fracta_mul[44]), .CK(clk), .Q(opa_r1[44]), .QN(
        n4664) );
  DFF_X2 opa_r1_reg_43_ ( .D(fracta_mul[43]), .CK(clk), .Q(opa_r1[43]), .QN(
        n4663) );
  DFF_X2 opa_r1_reg_42_ ( .D(fracta_mul[42]), .CK(clk), .Q(opa_r1[42]), .QN(
        n4662) );
  DFF_X2 opa_r1_reg_41_ ( .D(fracta_mul[41]), .CK(clk), .Q(opa_r1[41]), .QN(
        n4661) );
  DFF_X2 opa_r1_reg_40_ ( .D(fracta_mul[40]), .CK(clk), .Q(opa_r1[40]), .QN(
        n4660) );
  DFF_X2 opa_r1_reg_39_ ( .D(fracta_mul[39]), .CK(clk), .Q(opa_r1[39]), .QN(
        n4659) );
  DFF_X2 opa_r1_reg_38_ ( .D(fracta_mul[38]), .CK(clk), .Q(opa_r1[38]), .QN(
        n4658) );
  DFF_X2 opa_r1_reg_37_ ( .D(fracta_mul[37]), .CK(clk), .Q(opa_r1[37]), .QN(
        n4657) );
  DFF_X2 opa_r1_reg_36_ ( .D(fracta_mul[36]), .CK(clk), .Q(opa_r1[36]), .QN(
        n4656) );
  DFF_X2 opa_r1_reg_35_ ( .D(fracta_mul[35]), .CK(clk), .Q(opa_r1[35]), .QN(
        n4655) );
  DFF_X2 opa_r1_reg_34_ ( .D(fracta_mul[34]), .CK(clk), .Q(opa_r1[34]), .QN(
        n4654) );
  DFF_X2 opa_r1_reg_33_ ( .D(fracta_mul[33]), .CK(clk), .Q(opa_r1[33]), .QN(
        n4653) );
  DFF_X2 opa_r1_reg_32_ ( .D(fracta_mul[32]), .CK(clk), .Q(opa_r1[32]), .QN(
        n4652) );
  DFF_X2 opa_r1_reg_31_ ( .D(fracta_mul[31]), .CK(clk), .Q(opa_r1[31]), .QN(
        n4651) );
  DFF_X2 opa_r1_reg_30_ ( .D(fracta_mul[30]), .CK(clk), .Q(opa_r1[30]), .QN(
        n4650) );
  DFF_X2 opa_r1_reg_29_ ( .D(fracta_mul[29]), .CK(clk), .Q(opa_r1[29]), .QN(
        n4649) );
  DFF_X2 opa_r1_reg_28_ ( .D(fracta_mul[28]), .CK(clk), .Q(opa_r1[28]), .QN(
        n4648) );
  DFF_X2 opa_r1_reg_27_ ( .D(fracta_mul[27]), .CK(clk), .Q(opa_r1[27]), .QN(
        n4647) );
  DFF_X2 opa_r1_reg_26_ ( .D(fracta_mul[26]), .CK(clk), .Q(opa_r1[26]), .QN(
        n4646) );
  DFF_X2 opa_r1_reg_25_ ( .D(fracta_mul[25]), .CK(clk), .Q(opa_r1[25]), .QN(
        n4645) );
  DFF_X2 opa_r1_reg_24_ ( .D(fracta_mul[24]), .CK(clk), .Q(opa_r1[24]), .QN(
        n4644) );
  DFF_X2 opa_r1_reg_23_ ( .D(fracta_mul[23]), .CK(clk), .Q(opa_r1[23]), .QN(
        n4643) );
  DFF_X2 opa_r1_reg_22_ ( .D(fracta_mul[22]), .CK(clk), .Q(opa_r1[22]), .QN(
        n4642) );
  DFF_X2 opa_r1_reg_21_ ( .D(fracta_mul[21]), .CK(clk), .Q(opa_r1[21]), .QN(
        n4641) );
  DFF_X2 opa_r1_reg_20_ ( .D(fracta_mul[20]), .CK(clk), .Q(opa_r1[20]), .QN(
        n4640) );
  DFF_X2 opa_r1_reg_19_ ( .D(fracta_mul[19]), .CK(clk), .Q(opa_r1[19]), .QN(
        n4639) );
  DFF_X2 opa_r1_reg_18_ ( .D(fracta_mul[18]), .CK(clk), .Q(opa_r1[18]), .QN(
        n4638) );
  DFF_X2 opa_r1_reg_17_ ( .D(fracta_mul[17]), .CK(clk), .Q(opa_r1[17]), .QN(
        n4637) );
  DFF_X2 opa_r1_reg_16_ ( .D(fracta_mul[16]), .CK(clk), .Q(opa_r1[16]), .QN(
        n4636) );
  DFF_X2 opa_r1_reg_15_ ( .D(fracta_mul[15]), .CK(clk), .Q(opa_r1[15]), .QN(
        n4635) );
  DFF_X2 opa_r1_reg_14_ ( .D(fracta_mul[14]), .CK(clk), .Q(opa_r1[14]), .QN(
        n4524) );
  DFF_X2 opa_r1_reg_13_ ( .D(fracta_mul[13]), .CK(clk), .Q(opa_r1[13]), .QN(
        n4460) );
  DFF_X2 opa_r1_reg_12_ ( .D(fracta_mul[12]), .CK(clk), .Q(opa_r1[12]), .QN(
        n4459) );
  DFF_X2 opa_r1_reg_11_ ( .D(fracta_mul[11]), .CK(clk), .Q(opa_r1[11]), .QN(
        n4458) );
  DFF_X2 opa_r1_reg_10_ ( .D(fracta_mul[10]), .CK(clk), .Q(opa_r1[10]), .QN(
        n4457) );
  DFF_X2 opa_r1_reg_9_ ( .D(fracta_mul[9]), .CK(clk), .Q(opa_r1[9]), .QN(n4456) );
  DFF_X2 opa_r1_reg_8_ ( .D(fracta_mul[8]), .CK(clk), .Q(opa_r1[8]), .QN(n4455) );
  DFF_X2 opa_r1_reg_7_ ( .D(fracta_mul[7]), .CK(clk), .Q(opa_r1[7]), .QN(n4454) );
  DFF_X2 opa_r1_reg_6_ ( .D(fracta_mul[6]), .CK(clk), .Q(opa_r1[6]), .QN(n4453) );
  DFF_X2 opa_r1_reg_5_ ( .D(fracta_mul[5]), .CK(clk), .Q(opa_r1[5]), .QN(n4452) );
  DFF_X2 opa_r1_reg_4_ ( .D(fracta_mul[4]), .CK(clk), .Q(opa_r1[4]), .QN(n4421) );
  DFF_X2 opa_r1_reg_3_ ( .D(fracta_mul[3]), .CK(clk), .Q(opa_r1[3]), .QN(n4420) );
  DFF_X2 opa_r1_reg_2_ ( .D(fracta_mul[2]), .CK(clk), .Q(opa_r1[2]), .QN(n4451) );
  DFF_X2 opa_r1_reg_1_ ( .D(fracta_mul[1]), .CK(clk), .Q(opa_r1[1]), .QN(n4627) );
  DFF_X2 opa_r1_reg_0_ ( .D(fracta_mul[0]), .CK(clk), .Q(N347), .QN(n4402) );
  DFF_X2 opas_r1_reg ( .D(opa_r[63]), .CK(clk), .Q(opas_r1) );
  DFF_X2 opas_r2_reg ( .D(opas_r1), .CK(clk), .Q(opas_r2), .QN(n4574) );
  DFF_X2 u0_fractb_00_reg ( .D(n4350), .CK(clk), .Q(u0_fractb_00) );
  DFF_X2 u0_fracta_00_reg ( .D(n4349), .CK(clk), .Q(u0_fracta_00) );
  DFF_X2 u0_expb_00_reg ( .D(n6373), .CK(clk), .Q(u0_expb_00) );
  DFF_X2 u0_opb_dn_reg ( .D(u0_expb_00), .CK(clk), .Q(opb_dn), .QN(n4479) );
  DFF_X2 u0_opb_00_reg ( .D(u0_N17), .CK(clk), .Q(opb_00), .QN(n4504) );
  DFF_X2 u0_expa_00_reg ( .D(n4824), .CK(clk), .Q(u0_expa_00) );
  DFF_X2 u0_opa_dn_reg ( .D(u0_expa_00), .CK(clk), .QN(n4426) );
  DFF_X2 u0_opa_00_reg ( .D(u0_N16), .CK(clk), .Q(opa_00), .QN(n4493) );
  DFF_X2 u0_opb_nan_reg ( .D(u0_N11), .CK(clk), .Q(opb_nan), .QN(n4633) );
  DFF_X2 u0_opa_nan_reg ( .D(u0_N10), .CK(clk), .Q(opa_nan), .QN(n4628) );
  DFF_X2 opa_nan_r_reg ( .D(N917), .CK(clk), .Q(opa_nan_r) );
  DFF_X2 u0_snan_r_b_reg ( .D(u0_N5), .CK(clk), .Q(u0_snan_r_b) );
  DFF_X2 u0_qnan_r_b_reg ( .D(u6_N51), .CK(clk), .Q(u0_qnan_r_b) );
  DFF_X2 u0_snan_r_a_reg ( .D(u0_N4), .CK(clk), .Q(u0_snan_r_a) );
  DFF_X2 u0_qnan_r_a_reg ( .D(fracta_mul[51]), .CK(clk), .Q(u0_qnan_r_a) );
  DFF_X2 u0_infb_f_r_reg ( .D(n4350), .CK(clk), .Q(u0_infb_f_r) );
  DFF_X2 u0_infa_f_r_reg ( .D(n4349), .CK(clk), .Q(u0_infa_f_r) );
  DFF_X2 u0_expb_ff_reg ( .D(n6372), .CK(clk), .Q(u0_expb_ff) );
  DFF_X2 u0_opb_inf_reg ( .D(n6395), .CK(clk), .Q(opb_inf), .QN(n4432) );
  DFF_X2 u0_expa_ff_reg ( .D(n6350), .CK(clk), .Q(u0_expa_ff) );
  DFF_X2 u0_snan_reg ( .D(n6393), .CK(clk), .Q(snan_d) );
  DFF_X2 snan_reg ( .D(snan_d), .CK(clk), .Q(snan) );
  DFF_X2 u0_qnan_reg ( .D(n6394), .CK(clk), .Q(qnan_d) );
  DFF_X2 u0_opa_inf_reg ( .D(n6396), .CK(clk), .Q(opa_inf), .QN(n4619) );
  DFF_X2 div_by_zero_reg ( .D(N918), .CK(clk), .Q(div_by_zero) );
  DFF_X2 u0_inf_reg ( .D(u0_N7), .CK(clk), .Q(inf_d), .QN(n4621) );
  DFF_X2 u0_ind_reg ( .D(u0_N6), .CK(clk), .QN(n4626) );
  DFF_X2 u1_fasu_op_reg ( .D(n3953), .CK(clk), .Q(fasu_op), .QN(n4422) );
  DFF_X2 fasu_op_r1_reg ( .D(n4879), .CK(clk), .Q(fasu_op_r1) );
  DFF_X2 fasu_op_r2_reg ( .D(fasu_op_r1), .CK(clk), .Q(fasu_op_r2) );
  DFF_X2 qnan_reg ( .D(N909), .CK(clk), .Q(qnan) );
  DFF_X2 u1_fracta_eq_fractb_reg ( .D(u1_N325), .CK(clk), .Q(
        u1_fracta_eq_fractb) );
  DFF_X2 u1_fracta_lt_fractb_reg ( .D(u1_N324), .CK(clk), .Q(
        u1_fracta_lt_fractb), .QN(n4632) );
  DFF_X2 u1_add_r_reg ( .D(n4620), .CK(clk), .Q(u1_add_r) );
  DFF_X2 u1_signb_r_reg ( .D(opb_r[63]), .CK(clk), .QN(n4624) );
  DFF_X2 u1_signa_r_reg ( .D(opa_r[63]), .CK(clk), .Q(u1_signa_r) );
  DFF_X2 u1_result_zero_sign_reg ( .D(n6374), .CK(clk), .Q(result_zero_sign_d)
         );
  DFF_X2 u1_nan_sign_reg ( .D(u1_N334), .CK(clk), .Q(nan_sign_d) );
  DLH_X2 u1_sticky_reg ( .G(u1_N295), .D(u1_N296), .Q(u1_sticky) );
  DFF_X2 u1_sign_reg ( .D(u1_sign_d), .CK(clk), .Q(sign_fasu) );
  DFF_X2 sign_fasu_r_reg ( .D(sign_fasu), .CK(clk), .Q(sign_fasu_r) );
  DFF_X2 u1_fractb_out_reg_9_ ( .D(u1_fractb_s[9]), .CK(clk), .Q(fractb[9]) );
  DFF_X2 u1_fractb_out_reg_8_ ( .D(u1_fractb_s[8]), .CK(clk), .Q(fractb[8]) );
  DFF_X2 u1_fractb_out_reg_7_ ( .D(u1_fractb_s[7]), .CK(clk), .Q(fractb[7]) );
  DFF_X2 u1_fractb_out_reg_6_ ( .D(u1_fractb_s[6]), .CK(clk), .Q(fractb[6]) );
  DFF_X2 u1_fractb_out_reg_5_ ( .D(u1_fractb_s[5]), .CK(clk), .Q(fractb[5]) );
  DFF_X2 u1_fractb_out_reg_55_ ( .D(u1_fractb_s[55]), .CK(clk), .Q(fractb[55])
         );
  DFF_X2 u1_fractb_out_reg_54_ ( .D(u1_fractb_s[54]), .CK(clk), .Q(fractb[54])
         );
  DFF_X2 u1_fractb_out_reg_53_ ( .D(u1_fractb_s[53]), .CK(clk), .Q(fractb[53])
         );
  DFF_X2 u1_fractb_out_reg_52_ ( .D(u1_fractb_s[52]), .CK(clk), .Q(fractb[52])
         );
  DFF_X2 u1_fractb_out_reg_51_ ( .D(u1_fractb_s[51]), .CK(clk), .Q(fractb[51])
         );
  DFF_X2 u1_fractb_out_reg_50_ ( .D(u1_fractb_s[50]), .CK(clk), .Q(fractb[50])
         );
  DFF_X2 u1_fractb_out_reg_4_ ( .D(u1_fractb_s[4]), .CK(clk), .Q(fractb[4]) );
  DFF_X2 u1_fractb_out_reg_49_ ( .D(u1_fractb_s[49]), .CK(clk), .Q(fractb[49])
         );
  DFF_X2 u1_fractb_out_reg_48_ ( .D(u1_fractb_s[48]), .CK(clk), .Q(fractb[48])
         );
  DFF_X2 u1_fractb_out_reg_47_ ( .D(u1_fractb_s[47]), .CK(clk), .Q(fractb[47])
         );
  DFF_X2 u1_fractb_out_reg_46_ ( .D(u1_fractb_s[46]), .CK(clk), .Q(fractb[46])
         );
  DFF_X2 u1_fractb_out_reg_45_ ( .D(u1_fractb_s[45]), .CK(clk), .Q(fractb[45])
         );
  DFF_X2 u1_fractb_out_reg_44_ ( .D(u1_fractb_s[44]), .CK(clk), .Q(fractb[44])
         );
  DFF_X2 u1_fractb_out_reg_43_ ( .D(u1_fractb_s[43]), .CK(clk), .Q(fractb[43])
         );
  DFF_X2 u1_fractb_out_reg_42_ ( .D(u1_fractb_s[42]), .CK(clk), .Q(fractb[42])
         );
  DFF_X2 u1_fractb_out_reg_41_ ( .D(u1_fractb_s[41]), .CK(clk), .Q(fractb[41])
         );
  DFF_X2 u1_fractb_out_reg_40_ ( .D(u1_fractb_s[40]), .CK(clk), .Q(fractb[40])
         );
  DFF_X2 u1_fractb_out_reg_3_ ( .D(u1_fractb_s[3]), .CK(clk), .Q(fractb[3]) );
  DFF_X2 u1_fractb_out_reg_39_ ( .D(u1_fractb_s[39]), .CK(clk), .Q(fractb[39])
         );
  DFF_X2 u1_fractb_out_reg_38_ ( .D(u1_fractb_s[38]), .CK(clk), .Q(fractb[38])
         );
  DFF_X2 u1_fractb_out_reg_37_ ( .D(u1_fractb_s[37]), .CK(clk), .Q(fractb[37])
         );
  DFF_X2 u1_fractb_out_reg_36_ ( .D(u1_fractb_s[36]), .CK(clk), .Q(fractb[36])
         );
  DFF_X2 u1_fractb_out_reg_35_ ( .D(u1_fractb_s[35]), .CK(clk), .Q(fractb[35])
         );
  DFF_X2 u1_fractb_out_reg_34_ ( .D(u1_fractb_s[34]), .CK(clk), .Q(fractb[34])
         );
  DFF_X2 u1_fractb_out_reg_33_ ( .D(u1_fractb_s[33]), .CK(clk), .Q(fractb[33])
         );
  DFF_X2 u1_fractb_out_reg_32_ ( .D(u1_fractb_s[32]), .CK(clk), .Q(fractb[32])
         );
  DFF_X2 u1_fractb_out_reg_31_ ( .D(u1_fractb_s[31]), .CK(clk), .Q(fractb[31])
         );
  DFF_X2 u1_fractb_out_reg_30_ ( .D(u1_fractb_s[30]), .CK(clk), .Q(fractb[30])
         );
  DFF_X2 u1_fractb_out_reg_2_ ( .D(u1_fractb_s[2]), .CK(clk), .Q(fractb[2]) );
  DFF_X2 u1_fractb_out_reg_29_ ( .D(u1_fractb_s[29]), .CK(clk), .Q(fractb[29])
         );
  DFF_X2 u1_fractb_out_reg_28_ ( .D(u1_fractb_s[28]), .CK(clk), .Q(fractb[28])
         );
  DFF_X2 u1_fractb_out_reg_27_ ( .D(u1_fractb_s[27]), .CK(clk), .Q(fractb[27])
         );
  DFF_X2 u1_fractb_out_reg_26_ ( .D(u1_fractb_s[26]), .CK(clk), .Q(fractb[26])
         );
  DFF_X2 u1_fractb_out_reg_25_ ( .D(u1_fractb_s[25]), .CK(clk), .Q(fractb[25])
         );
  DFF_X2 u1_fractb_out_reg_24_ ( .D(u1_fractb_s[24]), .CK(clk), .Q(fractb[24])
         );
  DFF_X2 u1_fractb_out_reg_23_ ( .D(u1_fractb_s[23]), .CK(clk), .Q(fractb[23])
         );
  DFF_X2 u1_fractb_out_reg_22_ ( .D(u1_fractb_s[22]), .CK(clk), .Q(fractb[22])
         );
  DFF_X2 u1_fractb_out_reg_21_ ( .D(u1_fractb_s[21]), .CK(clk), .Q(fractb[21])
         );
  DFF_X2 u1_fractb_out_reg_20_ ( .D(u1_fractb_s[20]), .CK(clk), .Q(fractb[20])
         );
  DFF_X2 u1_fractb_out_reg_1_ ( .D(u1_fractb_s[1]), .CK(clk), .Q(fractb[1]) );
  DFF_X2 u1_fractb_out_reg_19_ ( .D(u1_fractb_s[19]), .CK(clk), .Q(fractb[19])
         );
  DFF_X2 u1_fractb_out_reg_18_ ( .D(u1_fractb_s[18]), .CK(clk), .Q(fractb[18])
         );
  DFF_X2 u1_fractb_out_reg_17_ ( .D(u1_fractb_s[17]), .CK(clk), .Q(fractb[17])
         );
  DFF_X2 u1_fractb_out_reg_16_ ( .D(u1_fractb_s[16]), .CK(clk), .Q(fractb[16])
         );
  DFF_X2 u1_fractb_out_reg_15_ ( .D(u1_fractb_s[15]), .CK(clk), .Q(fractb[15])
         );
  DFF_X2 u1_fractb_out_reg_14_ ( .D(u1_fractb_s[14]), .CK(clk), .Q(fractb[14])
         );
  DFF_X2 u1_fractb_out_reg_13_ ( .D(u1_fractb_s[13]), .CK(clk), .Q(fractb[13])
         );
  DFF_X2 u1_fractb_out_reg_12_ ( .D(u1_fractb_s[12]), .CK(clk), .Q(fractb[12])
         );
  DFF_X2 u1_fractb_out_reg_11_ ( .D(u1_fractb_s[11]), .CK(clk), .Q(fractb[11])
         );
  DFF_X2 u1_fractb_out_reg_10_ ( .D(u1_fractb_s[10]), .CK(clk), .Q(fractb[10])
         );
  DFF_X2 u1_fracta_out_reg_9_ ( .D(u1_fracta_s[9]), .CK(clk), .Q(fracta[9]) );
  DFF_X2 u1_fracta_out_reg_8_ ( .D(u1_fracta_s[8]), .CK(clk), .Q(fracta[8]) );
  DFF_X2 u1_fracta_out_reg_7_ ( .D(u1_fracta_s[7]), .CK(clk), .Q(fracta[7]) );
  DFF_X2 u1_fracta_out_reg_6_ ( .D(u1_fracta_s[6]), .CK(clk), .Q(fracta[6]) );
  DFF_X2 u1_fracta_out_reg_5_ ( .D(u1_fracta_s[5]), .CK(clk), .Q(fracta[5]) );
  DFF_X2 u1_fracta_out_reg_55_ ( .D(u1_fracta_s[55]), .CK(clk), .Q(fracta[55])
         );
  DFF_X2 u1_fracta_out_reg_54_ ( .D(u1_fracta_s[54]), .CK(clk), .Q(fracta[54])
         );
  DFF_X2 u1_fracta_out_reg_53_ ( .D(u1_fracta_s[53]), .CK(clk), .Q(fracta[53])
         );
  DFF_X2 u1_fracta_out_reg_52_ ( .D(u1_fracta_s[52]), .CK(clk), .Q(fracta[52])
         );
  DFF_X2 u1_fracta_out_reg_51_ ( .D(u1_fracta_s[51]), .CK(clk), .Q(fracta[51])
         );
  DFF_X2 u1_fracta_out_reg_50_ ( .D(u1_fracta_s[50]), .CK(clk), .Q(fracta[50])
         );
  DFF_X2 u1_fracta_out_reg_4_ ( .D(u1_fracta_s[4]), .CK(clk), .Q(fracta[4]) );
  DFF_X2 u1_fracta_out_reg_49_ ( .D(u1_fracta_s[49]), .CK(clk), .Q(fracta[49])
         );
  DFF_X2 u1_fracta_out_reg_48_ ( .D(u1_fracta_s[48]), .CK(clk), .Q(fracta[48])
         );
  DFF_X2 u1_fracta_out_reg_47_ ( .D(u1_fracta_s[47]), .CK(clk), .Q(fracta[47])
         );
  DFF_X2 u1_fracta_out_reg_46_ ( .D(u1_fracta_s[46]), .CK(clk), .Q(fracta[46])
         );
  DFF_X2 u1_fracta_out_reg_45_ ( .D(u1_fracta_s[45]), .CK(clk), .Q(fracta[45])
         );
  DFF_X2 u1_fracta_out_reg_44_ ( .D(u1_fracta_s[44]), .CK(clk), .Q(fracta[44])
         );
  DFF_X2 u1_fracta_out_reg_43_ ( .D(u1_fracta_s[43]), .CK(clk), .Q(fracta[43])
         );
  DFF_X2 u1_fracta_out_reg_42_ ( .D(u1_fracta_s[42]), .CK(clk), .Q(fracta[42])
         );
  DFF_X2 u1_fracta_out_reg_41_ ( .D(u1_fracta_s[41]), .CK(clk), .Q(fracta[41])
         );
  DFF_X2 u1_fracta_out_reg_40_ ( .D(u1_fracta_s[40]), .CK(clk), .Q(fracta[40])
         );
  DFF_X2 u1_fracta_out_reg_3_ ( .D(u1_fracta_s[3]), .CK(clk), .Q(fracta[3]) );
  DFF_X2 u1_fracta_out_reg_39_ ( .D(u1_fracta_s[39]), .CK(clk), .Q(fracta[39])
         );
  DFF_X2 u1_fracta_out_reg_38_ ( .D(u1_fracta_s[38]), .CK(clk), .Q(fracta[38])
         );
  DFF_X2 u1_fracta_out_reg_37_ ( .D(u1_fracta_s[37]), .CK(clk), .Q(fracta[37])
         );
  DFF_X2 u1_fracta_out_reg_36_ ( .D(u1_fracta_s[36]), .CK(clk), .Q(fracta[36])
         );
  DFF_X2 u1_fracta_out_reg_35_ ( .D(u1_fracta_s[35]), .CK(clk), .Q(fracta[35])
         );
  DFF_X2 u1_fracta_out_reg_34_ ( .D(u1_fracta_s[34]), .CK(clk), .Q(fracta[34])
         );
  DFF_X2 u1_fracta_out_reg_33_ ( .D(u1_fracta_s[33]), .CK(clk), .Q(fracta[33])
         );
  DFF_X2 u1_fracta_out_reg_32_ ( .D(u1_fracta_s[32]), .CK(clk), .Q(fracta[32])
         );
  DFF_X2 u1_fracta_out_reg_31_ ( .D(u1_fracta_s[31]), .CK(clk), .Q(fracta[31])
         );
  DFF_X2 u1_fracta_out_reg_30_ ( .D(u1_fracta_s[30]), .CK(clk), .Q(fracta[30])
         );
  DFF_X2 u1_fracta_out_reg_2_ ( .D(u1_fracta_s[2]), .CK(clk), .Q(fracta[2]) );
  DFF_X2 u1_fracta_out_reg_29_ ( .D(u1_fracta_s[29]), .CK(clk), .Q(fracta[29])
         );
  DFF_X2 u1_fracta_out_reg_28_ ( .D(u1_fracta_s[28]), .CK(clk), .Q(fracta[28])
         );
  DFF_X2 u1_fracta_out_reg_27_ ( .D(u1_fracta_s[27]), .CK(clk), .Q(fracta[27])
         );
  DFF_X2 u1_fracta_out_reg_26_ ( .D(u1_fracta_s[26]), .CK(clk), .Q(fracta[26])
         );
  DFF_X2 u1_fracta_out_reg_25_ ( .D(u1_fracta_s[25]), .CK(clk), .Q(fracta[25])
         );
  DFF_X2 u1_fracta_out_reg_24_ ( .D(u1_fracta_s[24]), .CK(clk), .Q(fracta[24])
         );
  DFF_X2 u1_fracta_out_reg_23_ ( .D(u1_fracta_s[23]), .CK(clk), .Q(fracta[23])
         );
  DFF_X2 u1_fracta_out_reg_22_ ( .D(u1_fracta_s[22]), .CK(clk), .Q(fracta[22])
         );
  DFF_X2 u1_fracta_out_reg_21_ ( .D(u1_fracta_s[21]), .CK(clk), .Q(fracta[21])
         );
  DFF_X2 u1_fracta_out_reg_20_ ( .D(u1_fracta_s[20]), .CK(clk), .Q(fracta[20])
         );
  DFF_X2 u1_fracta_out_reg_1_ ( .D(u1_fracta_s[1]), .CK(clk), .Q(fracta[1]) );
  DFF_X2 u1_fracta_out_reg_19_ ( .D(u1_fracta_s[19]), .CK(clk), .Q(fracta[19])
         );
  DFF_X2 u1_fracta_out_reg_18_ ( .D(u1_fracta_s[18]), .CK(clk), .Q(fracta[18])
         );
  DFF_X2 u1_fracta_out_reg_17_ ( .D(u1_fracta_s[17]), .CK(clk), .Q(fracta[17])
         );
  DFF_X2 u1_fracta_out_reg_16_ ( .D(u1_fracta_s[16]), .CK(clk), .Q(fracta[16])
         );
  DFF_X2 u1_fracta_out_reg_15_ ( .D(u1_fracta_s[15]), .CK(clk), .Q(fracta[15])
         );
  DFF_X2 u1_fracta_out_reg_14_ ( .D(u1_fracta_s[14]), .CK(clk), .Q(fracta[14])
         );
  DFF_X2 u1_fracta_out_reg_13_ ( .D(u1_fracta_s[13]), .CK(clk), .Q(fracta[13])
         );
  DFF_X2 u1_fracta_out_reg_12_ ( .D(u1_fracta_s[12]), .CK(clk), .Q(fracta[12])
         );
  DFF_X2 u1_fracta_out_reg_11_ ( .D(u1_fracta_s[11]), .CK(clk), .Q(fracta[11])
         );
  DFF_X2 u1_fracta_out_reg_10_ ( .D(u1_fracta_s[10]), .CK(clk), .Q(fracta[10])
         );
  DFF_X2 u1_fractb_out_reg_0_ ( .D(u1_fractb_s[0]), .CK(clk), .Q(fractb[0]) );
  DFF_X2 u1_fracta_out_reg_0_ ( .D(u1_fracta_s[0]), .CK(clk), .Q(fracta[0]) );
  DFF_X2 fract_out_q_reg_0_ ( .D(n6160), .CK(clk), .Q(fract_out_q[0]) );
  DFF_X2 fract_out_q_reg_1_ ( .D(n6159), .CK(clk), .Q(fract_out_q[1]) );
  DFF_X2 fract_out_q_reg_2_ ( .D(n6158), .CK(clk), .Q(fract_out_q[2]) );
  DFF_X2 fract_out_q_reg_3_ ( .D(n6157), .CK(clk), .Q(fract_out_q[3]) );
  DFF_X2 fract_out_q_reg_4_ ( .D(n6156), .CK(clk), .Q(fract_out_q[4]) );
  DFF_X2 fract_out_q_reg_5_ ( .D(n6155), .CK(clk), .Q(fract_out_q[5]) );
  DFF_X2 fract_out_q_reg_6_ ( .D(n6154), .CK(clk), .Q(fract_out_q[6]) );
  DFF_X2 fract_out_q_reg_7_ ( .D(n6153), .CK(clk), .Q(fract_out_q[7]) );
  DFF_X2 fract_out_q_reg_8_ ( .D(n6152), .CK(clk), .Q(fract_out_q[8]) );
  DFF_X2 fract_out_q_reg_9_ ( .D(n6151), .CK(clk), .Q(fract_out_q[9]) );
  DFF_X2 fract_out_q_reg_10_ ( .D(n6150), .CK(clk), .Q(fract_out_q[10]) );
  DFF_X2 fract_out_q_reg_11_ ( .D(n6149), .CK(clk), .Q(fract_out_q[11]) );
  DFF_X2 fract_out_q_reg_12_ ( .D(n6148), .CK(clk), .Q(fract_out_q[12]) );
  DFF_X2 fract_out_q_reg_13_ ( .D(n6147), .CK(clk), .Q(fract_out_q[13]) );
  DFF_X2 fract_out_q_reg_14_ ( .D(n6146), .CK(clk), .Q(fract_out_q[14]) );
  DFF_X2 fract_out_q_reg_15_ ( .D(n6145), .CK(clk), .Q(fract_out_q[15]) );
  DFF_X2 fract_out_q_reg_16_ ( .D(n6144), .CK(clk), .Q(fract_out_q[16]) );
  DFF_X2 fract_out_q_reg_17_ ( .D(n6143), .CK(clk), .Q(fract_out_q[17]) );
  DFF_X2 fract_out_q_reg_18_ ( .D(n6142), .CK(clk), .Q(fract_out_q[18]) );
  DFF_X2 fract_out_q_reg_19_ ( .D(n6141), .CK(clk), .Q(fract_out_q[19]) );
  DFF_X2 fract_out_q_reg_20_ ( .D(n6140), .CK(clk), .Q(fract_out_q[20]) );
  DFF_X2 fract_out_q_reg_21_ ( .D(n6139), .CK(clk), .Q(fract_out_q[21]) );
  DFF_X2 fract_out_q_reg_22_ ( .D(n6138), .CK(clk), .Q(fract_out_q[22]) );
  DFF_X2 fract_out_q_reg_23_ ( .D(n6137), .CK(clk), .Q(fract_out_q[23]) );
  DFF_X2 fract_out_q_reg_24_ ( .D(n6136), .CK(clk), .Q(fract_out_q[24]) );
  DFF_X2 fract_out_q_reg_25_ ( .D(n6135), .CK(clk), .Q(fract_out_q[25]) );
  DFF_X2 fract_out_q_reg_26_ ( .D(n6134), .CK(clk), .Q(fract_out_q[26]) );
  DFF_X2 fract_out_q_reg_27_ ( .D(n6133), .CK(clk), .Q(fract_out_q[27]) );
  DFF_X2 fract_out_q_reg_28_ ( .D(n6132), .CK(clk), .Q(fract_out_q[28]) );
  DFF_X2 fract_out_q_reg_29_ ( .D(n6131), .CK(clk), .Q(fract_out_q[29]) );
  DFF_X2 fract_out_q_reg_30_ ( .D(n6130), .CK(clk), .Q(fract_out_q[30]) );
  DFF_X2 fract_out_q_reg_31_ ( .D(n6129), .CK(clk), .Q(fract_out_q[31]) );
  DFF_X2 fract_out_q_reg_32_ ( .D(n6128), .CK(clk), .Q(fract_out_q[32]) );
  DFF_X2 fract_out_q_reg_33_ ( .D(n6127), .CK(clk), .Q(fract_out_q[33]) );
  DFF_X2 fract_out_q_reg_34_ ( .D(n6126), .CK(clk), .Q(fract_out_q[34]) );
  DFF_X2 fract_out_q_reg_35_ ( .D(n6125), .CK(clk), .Q(fract_out_q[35]) );
  DFF_X2 fract_out_q_reg_36_ ( .D(n6124), .CK(clk), .Q(fract_out_q[36]) );
  DFF_X2 fract_out_q_reg_37_ ( .D(n6123), .CK(clk), .Q(fract_out_q[37]) );
  DFF_X2 fract_out_q_reg_38_ ( .D(n6122), .CK(clk), .Q(fract_out_q[38]) );
  DFF_X2 fract_out_q_reg_39_ ( .D(n6121), .CK(clk), .Q(fract_out_q[39]) );
  DFF_X2 fract_out_q_reg_40_ ( .D(n6120), .CK(clk), .Q(fract_out_q[40]) );
  DFF_X2 fract_out_q_reg_41_ ( .D(n6119), .CK(clk), .Q(fract_out_q[41]) );
  DFF_X2 fract_out_q_reg_42_ ( .D(n6118), .CK(clk), .Q(fract_out_q[42]) );
  DFF_X2 fract_out_q_reg_43_ ( .D(n6117), .CK(clk), .Q(fract_out_q[43]) );
  DFF_X2 fract_out_q_reg_44_ ( .D(n6116), .CK(clk), .Q(fract_out_q[44]) );
  DFF_X2 fract_out_q_reg_45_ ( .D(n6115), .CK(clk), .Q(fract_out_q[45]) );
  DFF_X2 fract_out_q_reg_46_ ( .D(n6114), .CK(clk), .Q(fract_out_q[46]) );
  DFF_X2 fract_out_q_reg_47_ ( .D(n6113), .CK(clk), .Q(fract_out_q[47]) );
  DFF_X2 fract_out_q_reg_48_ ( .D(n6112), .CK(clk), .Q(fract_out_q[48]) );
  DFF_X2 fract_out_q_reg_49_ ( .D(n6111), .CK(clk), .Q(fract_out_q[49]) );
  DFF_X2 fract_out_q_reg_50_ ( .D(n6110), .CK(clk), .Q(fract_out_q[50]) );
  DFF_X2 fract_out_q_reg_51_ ( .D(n6109), .CK(clk), .Q(fract_out_q[51]) );
  DFF_X2 fract_out_q_reg_52_ ( .D(n6108), .CK(clk), .Q(fract_out_q[52]) );
  DFF_X2 fract_out_q_reg_53_ ( .D(n6107), .CK(clk), .Q(fract_out_q[53]) );
  DFF_X2 fract_out_q_reg_54_ ( .D(n6106), .CK(clk), .Q(fract_out_q[54]) );
  DFF_X2 fract_out_q_reg_55_ ( .D(n6105), .CK(clk), .Q(fract_out_q[55]) );
  DFF_X2 fract_out_q_reg_56_ ( .D(n6104), .CK(clk), .Q(fract_out_q[56]) );
  DFF_X2 u1_exp_dn_out_reg_0_ ( .D(u1_N78), .CK(clk), .Q(exp_fasu[0]) );
  DFF_X2 u1_exp_dn_out_reg_1_ ( .D(u1_N79), .CK(clk), .Q(exp_fasu[1]) );
  DFF_X2 u1_exp_dn_out_reg_2_ ( .D(u1_N80), .CK(clk), .Q(exp_fasu[2]) );
  DFF_X2 u1_exp_dn_out_reg_3_ ( .D(u1_N81), .CK(clk), .Q(exp_fasu[3]) );
  DFF_X2 u1_exp_dn_out_reg_4_ ( .D(u1_N82), .CK(clk), .Q(exp_fasu[4]) );
  DFF_X2 u1_exp_dn_out_reg_5_ ( .D(u1_N83), .CK(clk), .Q(exp_fasu[5]) );
  DFF_X2 u1_exp_dn_out_reg_6_ ( .D(u1_N84), .CK(clk), .Q(exp_fasu[6]) );
  DFF_X2 u1_exp_dn_out_reg_7_ ( .D(u1_N85), .CK(clk), .Q(exp_fasu[7]) );
  DFF_X2 u1_exp_dn_out_reg_8_ ( .D(u1_N86), .CK(clk), .Q(exp_fasu[8]) );
  DFF_X2 u1_exp_dn_out_reg_9_ ( .D(u1_N87), .CK(clk), .Q(exp_fasu[9]) );
  DFF_X2 u1_exp_dn_out_reg_10_ ( .D(u1_N88), .CK(clk), .Q(exp_fasu[10]) );
  DFF_X2 u2_sign_exe_reg ( .D(u2_N121), .CK(clk), .Q(sign_exe) );
  DFF_X2 sign_exe_r_reg ( .D(sign_exe), .CK(clk), .Q(sign_exe_r), .QN(n4630)
         );
  DFF_X2 u2_sign_reg ( .D(u2_sign_d), .CK(clk), .Q(sign_mul) );
  DFF_X2 sign_mul_r_reg ( .D(sign_mul), .CK(clk), .Q(sign_mul_r), .QN(n4667)
         );
  DFF_X2 sign_reg ( .D(N794), .CK(clk), .Q(sign), .QN(n4494) );
  DFF_X2 fract_i2f_reg_105_ ( .D(N667), .CK(clk), .Q(fract_i2f[105]) );
  DFF_X2 fract_i2f_reg_104_ ( .D(N666), .CK(clk), .Q(fract_i2f[104]) );
  DFF_X2 fract_i2f_reg_103_ ( .D(N665), .CK(clk), .Q(fract_i2f[103]) );
  DFF_X2 fract_i2f_reg_102_ ( .D(N664), .CK(clk), .Q(fract_i2f[102]) );
  DFF_X2 fract_i2f_reg_101_ ( .D(N663), .CK(clk), .Q(fract_i2f[101]) );
  DFF_X2 fract_i2f_reg_100_ ( .D(N662), .CK(clk), .Q(fract_i2f[100]) );
  DFF_X2 fract_i2f_reg_99_ ( .D(N661), .CK(clk), .Q(fract_i2f[99]) );
  DFF_X2 fract_i2f_reg_98_ ( .D(N660), .CK(clk), .Q(fract_i2f[98]) );
  DFF_X2 fract_i2f_reg_97_ ( .D(N659), .CK(clk), .Q(fract_i2f[97]) );
  DFF_X2 fract_i2f_reg_96_ ( .D(N658), .CK(clk), .Q(fract_i2f[96]) );
  DFF_X2 fract_i2f_reg_95_ ( .D(N657), .CK(clk), .Q(fract_i2f[95]) );
  DFF_X2 fract_i2f_reg_94_ ( .D(N656), .CK(clk), .Q(fract_i2f[94]) );
  DFF_X2 fract_i2f_reg_93_ ( .D(N655), .CK(clk), .Q(fract_i2f[93]) );
  DFF_X2 fract_i2f_reg_92_ ( .D(N654), .CK(clk), .Q(fract_i2f[92]) );
  DFF_X2 fract_i2f_reg_91_ ( .D(N653), .CK(clk), .Q(fract_i2f[91]) );
  DFF_X2 fract_i2f_reg_90_ ( .D(N652), .CK(clk), .Q(fract_i2f[90]) );
  DFF_X2 fract_i2f_reg_89_ ( .D(N651), .CK(clk), .Q(fract_i2f[89]) );
  DFF_X2 fract_i2f_reg_88_ ( .D(N650), .CK(clk), .Q(fract_i2f[88]) );
  DFF_X2 fract_i2f_reg_87_ ( .D(N649), .CK(clk), .Q(fract_i2f[87]) );
  DFF_X2 fract_i2f_reg_86_ ( .D(N648), .CK(clk), .Q(fract_i2f[86]) );
  DFF_X2 fract_i2f_reg_85_ ( .D(N647), .CK(clk), .Q(fract_i2f[85]) );
  DFF_X2 fract_i2f_reg_84_ ( .D(N646), .CK(clk), .Q(fract_i2f[84]) );
  DFF_X2 fract_i2f_reg_83_ ( .D(N645), .CK(clk), .Q(fract_i2f[83]) );
  DFF_X2 fract_i2f_reg_82_ ( .D(N644), .CK(clk), .Q(fract_i2f[82]) );
  DFF_X2 fract_i2f_reg_81_ ( .D(N643), .CK(clk), .Q(fract_i2f[81]) );
  DFF_X2 fract_i2f_reg_80_ ( .D(N642), .CK(clk), .Q(fract_i2f[80]) );
  DFF_X2 fract_i2f_reg_79_ ( .D(N641), .CK(clk), .Q(fract_i2f[79]) );
  DFF_X2 fract_i2f_reg_78_ ( .D(N640), .CK(clk), .Q(fract_i2f[78]) );
  DFF_X2 fract_i2f_reg_77_ ( .D(N639), .CK(clk), .Q(fract_i2f[77]) );
  DFF_X2 fract_i2f_reg_76_ ( .D(N638), .CK(clk), .Q(fract_i2f[76]) );
  DFF_X2 fract_i2f_reg_75_ ( .D(N637), .CK(clk), .Q(fract_i2f[75]) );
  DFF_X2 fract_i2f_reg_74_ ( .D(N636), .CK(clk), .Q(fract_i2f[74]) );
  DFF_X2 fract_i2f_reg_73_ ( .D(N635), .CK(clk), .Q(fract_i2f[73]) );
  DFF_X2 fract_i2f_reg_72_ ( .D(N634), .CK(clk), .Q(fract_i2f[72]) );
  DFF_X2 fract_i2f_reg_71_ ( .D(N633), .CK(clk), .Q(fract_i2f[71]) );
  DFF_X2 fract_i2f_reg_70_ ( .D(N632), .CK(clk), .Q(fract_i2f[70]) );
  DFF_X2 fract_i2f_reg_69_ ( .D(N631), .CK(clk), .Q(fract_i2f[69]) );
  DFF_X2 fract_i2f_reg_68_ ( .D(N630), .CK(clk), .Q(fract_i2f[68]) );
  DFF_X2 fract_i2f_reg_67_ ( .D(N629), .CK(clk), .Q(fract_i2f[67]) );
  DFF_X2 fract_i2f_reg_66_ ( .D(N628), .CK(clk), .Q(fract_i2f[66]) );
  DFF_X2 fract_i2f_reg_65_ ( .D(N627), .CK(clk), .Q(fract_i2f[65]) );
  DFF_X2 fract_i2f_reg_64_ ( .D(N626), .CK(clk), .Q(fract_i2f[64]) );
  DFF_X2 fract_i2f_reg_63_ ( .D(N625), .CK(clk), .Q(fract_i2f[63]) );
  DFF_X2 fract_i2f_reg_62_ ( .D(N624), .CK(clk), .Q(fract_i2f[62]) );
  DFF_X2 fract_i2f_reg_61_ ( .D(N623), .CK(clk), .Q(fract_i2f[61]) );
  DFF_X2 fract_i2f_reg_60_ ( .D(N622), .CK(clk), .Q(fract_i2f[60]) );
  DFF_X2 fract_i2f_reg_59_ ( .D(N621), .CK(clk), .Q(fract_i2f[59]) );
  DFF_X2 fract_i2f_reg_58_ ( .D(N620), .CK(clk), .Q(fract_i2f[58]) );
  DFF_X2 fract_i2f_reg_57_ ( .D(N619), .CK(clk), .Q(fract_i2f[57]) );
  DFF_X2 fract_i2f_reg_56_ ( .D(N618), .CK(clk), .Q(fract_i2f[56]) );
  DFF_X2 fract_i2f_reg_55_ ( .D(N617), .CK(clk), .Q(fract_i2f[55]) );
  DFF_X2 fract_i2f_reg_54_ ( .D(N616), .CK(clk), .Q(fract_i2f[54]) );
  DFF_X2 fract_i2f_reg_53_ ( .D(N615), .CK(clk), .Q(fract_i2f[53]) );
  DFF_X2 fract_i2f_reg_52_ ( .D(N614), .CK(clk), .Q(fract_i2f[52]) );
  DFF_X2 fract_i2f_reg_51_ ( .D(N613), .CK(clk), .Q(fract_i2f[51]) );
  DFF_X2 fract_i2f_reg_50_ ( .D(N612), .CK(clk), .Q(fract_i2f[50]) );
  DFF_X2 fract_i2f_reg_49_ ( .D(N611), .CK(clk), .Q(fract_i2f[49]) );
  DFF_X2 fract_i2f_reg_48_ ( .D(N610), .CK(clk), .Q(fract_i2f[48]) );
  DFF_X2 fract_i2f_reg_47_ ( .D(N609), .CK(clk), .Q(fract_i2f[47]) );
  DFF_X2 fract_i2f_reg_46_ ( .D(N608), .CK(clk), .Q(fract_i2f[46]) );
  DFF_X2 fract_i2f_reg_45_ ( .D(n5980), .CK(clk), .Q(fract_i2f[45]) );
  DFF_X2 fract_i2f_reg_44_ ( .D(n5981), .CK(clk), .Q(fract_i2f[44]) );
  DFF_X2 fract_i2f_reg_43_ ( .D(n5982), .CK(clk), .Q(fract_i2f[43]) );
  DFF_X2 fract_i2f_reg_42_ ( .D(n5983), .CK(clk), .Q(fract_i2f[42]) );
  DFF_X2 fract_i2f_reg_41_ ( .D(n5984), .CK(clk), .Q(fract_i2f[41]) );
  DFF_X2 fract_i2f_reg_40_ ( .D(n5985), .CK(clk), .Q(fract_i2f[40]) );
  DFF_X2 fract_i2f_reg_39_ ( .D(n5986), .CK(clk), .Q(fract_i2f[39]) );
  DFF_X2 fract_i2f_reg_38_ ( .D(n5987), .CK(clk), .Q(fract_i2f[38]) );
  DFF_X2 fract_i2f_reg_37_ ( .D(n5988), .CK(clk), .Q(fract_i2f[37]) );
  DFF_X2 fract_i2f_reg_36_ ( .D(n5989), .CK(clk), .Q(fract_i2f[36]) );
  DFF_X2 fract_i2f_reg_35_ ( .D(n5990), .CK(clk), .Q(fract_i2f[35]) );
  DFF_X2 fract_i2f_reg_34_ ( .D(n5991), .CK(clk), .Q(fract_i2f[34]) );
  DFF_X2 fract_i2f_reg_33_ ( .D(n5992), .CK(clk), .Q(fract_i2f[33]) );
  DFF_X2 fract_i2f_reg_32_ ( .D(n5993), .CK(clk), .Q(fract_i2f[32]) );
  DFF_X2 fract_i2f_reg_31_ ( .D(n5994), .CK(clk), .Q(fract_i2f[31]) );
  DFF_X2 fract_i2f_reg_30_ ( .D(n5995), .CK(clk), .Q(fract_i2f[30]) );
  DFF_X2 fract_i2f_reg_29_ ( .D(n5996), .CK(clk), .Q(fract_i2f[29]) );
  DFF_X2 fract_i2f_reg_28_ ( .D(n5997), .CK(clk), .Q(fract_i2f[28]) );
  DFF_X2 fract_i2f_reg_27_ ( .D(n5998), .CK(clk), .Q(fract_i2f[27]) );
  DFF_X2 fract_i2f_reg_26_ ( .D(n5999), .CK(clk), .Q(fract_i2f[26]) );
  DFF_X2 fract_i2f_reg_25_ ( .D(n6000), .CK(clk), .Q(fract_i2f[25]) );
  DFF_X2 fract_i2f_reg_24_ ( .D(n6001), .CK(clk), .Q(fract_i2f[24]) );
  DFF_X2 fract_i2f_reg_23_ ( .D(n6002), .CK(clk), .Q(fract_i2f[23]) );
  DFF_X2 fract_i2f_reg_22_ ( .D(n6003), .CK(clk), .Q(fract_i2f[22]) );
  DFF_X2 fract_i2f_reg_21_ ( .D(n6004), .CK(clk), .Q(fract_i2f[21]) );
  DFF_X2 fract_i2f_reg_20_ ( .D(n6005), .CK(clk), .Q(fract_i2f[20]) );
  DFF_X2 fract_i2f_reg_19_ ( .D(n6006), .CK(clk), .Q(fract_i2f[19]) );
  DFF_X2 fract_i2f_reg_18_ ( .D(n6007), .CK(clk), .Q(fract_i2f[18]) );
  DFF_X2 fract_i2f_reg_17_ ( .D(n6008), .CK(clk), .Q(fract_i2f[17]) );
  DFF_X2 fract_i2f_reg_16_ ( .D(n6009), .CK(clk), .Q(fract_i2f[16]) );
  DFF_X2 fract_i2f_reg_15_ ( .D(n6010), .CK(clk), .Q(fract_i2f[15]) );
  DFF_X2 fract_i2f_reg_14_ ( .D(n6011), .CK(clk), .Q(fract_i2f[14]) );
  DFF_X2 fract_i2f_reg_13_ ( .D(n6012), .CK(clk), .Q(fract_i2f[13]) );
  DFF_X2 fract_i2f_reg_12_ ( .D(n6013), .CK(clk), .Q(fract_i2f[12]) );
  DFF_X2 fract_i2f_reg_11_ ( .D(n6014), .CK(clk), .Q(fract_i2f[11]) );
  DFF_X2 fract_i2f_reg_10_ ( .D(n6015), .CK(clk), .Q(fract_i2f[10]) );
  DFF_X2 fract_i2f_reg_9_ ( .D(n6016), .CK(clk), .Q(fract_i2f[9]) );
  DFF_X2 fract_i2f_reg_8_ ( .D(n6017), .CK(clk), .Q(fract_i2f[8]) );
  DFF_X2 fract_i2f_reg_7_ ( .D(n6018), .CK(clk), .Q(fract_i2f[7]) );
  DFF_X2 fract_i2f_reg_6_ ( .D(n6019), .CK(clk), .Q(fract_i2f[6]) );
  DFF_X2 fract_i2f_reg_5_ ( .D(n6020), .CK(clk), .Q(fract_i2f[5]) );
  DFF_X2 fract_i2f_reg_4_ ( .D(n6021), .CK(clk), .Q(fract_i2f[4]) );
  DFF_X2 fract_i2f_reg_3_ ( .D(n6022), .CK(clk), .Q(fract_i2f[3]) );
  DFF_X2 fract_i2f_reg_2_ ( .D(n6023), .CK(clk), .Q(fract_i2f[2]) );
  DFF_X2 fract_i2f_reg_1_ ( .D(n6024), .CK(clk), .Q(fract_i2f[1]) );
  DFF_X2 fract_i2f_reg_0_ ( .D(n6380), .CK(clk), .Q(fract_i2f[0]) );
  DFF_X2 u2_inf_reg ( .D(u2_N114), .CK(clk), .Q(inf_mul) );
  DFF_X2 inf_mul_r_reg ( .D(inf_mul), .CK(clk), .Q(inf_mul_r) );
  DFF_X2 u2_underflow_reg_0_ ( .D(u2_underflow_d[0]), .CK(clk), .Q(
        underflow_fmul_d[0]) );
  DFF_X2 underflow_fmul_r_reg_0_ ( .D(underflow_fmul_d[0]), .CK(clk), .Q(
        underflow_fmul_r[0]) );
  DFF_X2 u2_underflow_reg_1_ ( .D(u2_underflow_d[1]), .CK(clk), .Q(
        underflow_fmul_d[1]) );
  DFF_X2 underflow_fmul_r_reg_1_ ( .D(underflow_fmul_d[1]), .CK(clk), .Q(
        underflow_fmul_r[1]) );
  DFF_X2 u2_underflow_reg_2_ ( .D(u2_underflow_d[2]), .CK(clk), .Q(
        underflow_fmul_d[2]) );
  DFF_X2 underflow_fmul_r_reg_2_ ( .D(underflow_fmul_d[2]), .CK(clk), .Q(
        underflow_fmul_r[2]) );
  DFF_X2 u2_exp_ovf_reg_0_ ( .D(u2_exp_ovf_d_0_), .CK(clk), .Q(exp_ovf[0]) );
  DFF_X2 exp_ovf_r_reg_0_ ( .D(exp_ovf[0]), .CK(clk), .Q(n4430), .QN(n4579) );
  DFF_X2 u2_exp_ovf_reg_1_ ( .D(u2_exp_ovf_d_1_), .CK(clk), .Q(exp_ovf[1]) );
  DFF_X2 exp_ovf_r_reg_1_ ( .D(exp_ovf[1]), .CK(clk), .Q(exp_ovf_r_1_), .QN(
        n4401) );
  DFF_X2 u2_exp_out_reg_0_ ( .D(u2_N76), .CK(clk), .Q(exp_mul[0]), .QN(n4525)
         );
  DFF_X2 u2_exp_out_reg_1_ ( .D(u2_N77), .CK(clk), .Q(exp_mul[1]) );
  DFF_X2 u2_exp_out_reg_2_ ( .D(u2_N78), .CK(clk), .Q(exp_mul[2]) );
  DFF_X2 u2_exp_out_reg_3_ ( .D(u2_N79), .CK(clk), .Q(exp_mul[3]) );
  DFF_X2 u2_exp_out_reg_4_ ( .D(u2_N80), .CK(clk), .Q(exp_mul[4]) );
  DFF_X2 u2_exp_out_reg_5_ ( .D(u2_N81), .CK(clk), .Q(exp_mul[5]) );
  DFF_X2 u2_exp_out_reg_6_ ( .D(u2_N82), .CK(clk), .Q(exp_mul[6]) );
  DFF_X2 u2_exp_out_reg_7_ ( .D(u2_N83), .CK(clk), .Q(exp_mul[7]) );
  DFF_X2 u2_exp_out_reg_8_ ( .D(u2_N84), .CK(clk), .Q(exp_mul[8]) );
  DFF_X2 u2_exp_out_reg_9_ ( .D(u2_N85), .CK(clk), .Q(exp_mul[9]) );
  DFF_X2 u2_exp_out_reg_10_ ( .D(u2_N86), .CK(clk), .Q(exp_mul[10]), .QN(n4668) );
  DFF_X2 inf_mul2_reg ( .D(N928), .CK(clk), .Q(inf_mul2) );
  DFF_X2 u5_prod1_reg_0_ ( .D(u5_N0), .CK(clk), .Q(u5_prod1[0]) );
  DFF_X2 u5_prod_reg_0_ ( .D(u5_prod1[0]), .CK(clk), .Q(prod[0]), .QN(n4714)
         );
  DFF_X2 u5_prod1_reg_1_ ( .D(u5_N1), .CK(clk), .Q(u5_prod1[1]) );
  DFF_X2 u5_prod_reg_1_ ( .D(u5_prod1[1]), .CK(clk), .QN(n4438) );
  DFF_X2 u5_prod1_reg_2_ ( .D(u5_N2), .CK(clk), .Q(u5_prod1[2]) );
  DFF_X2 u5_prod_reg_2_ ( .D(u5_prod1[2]), .CK(clk), .Q(prod[2]), .QN(n4705)
         );
  DFF_X2 u5_prod1_reg_3_ ( .D(u5_N3), .CK(clk), .Q(u5_prod1[3]) );
  DFF_X2 u5_prod_reg_3_ ( .D(u5_prod1[3]), .CK(clk), .Q(prod[3]), .QN(n4713)
         );
  DFF_X2 u5_prod1_reg_4_ ( .D(u5_N4), .CK(clk), .Q(u5_prod1[4]) );
  DFF_X2 u5_prod_reg_4_ ( .D(u5_prod1[4]), .CK(clk), .QN(n4446) );
  DFF_X2 u5_prod1_reg_5_ ( .D(u5_N5), .CK(clk), .Q(u5_prod1[5]) );
  DFF_X2 u5_prod_reg_5_ ( .D(u5_prod1[5]), .CK(clk), .Q(prod[5]), .QN(n4704)
         );
  DFF_X2 u5_prod1_reg_6_ ( .D(u5_N6), .CK(clk), .Q(u5_prod1[6]) );
  DFF_X2 u5_prod_reg_6_ ( .D(u5_prod1[6]), .CK(clk), .Q(prod[6]), .QN(n4712)
         );
  DFF_X2 u5_prod1_reg_7_ ( .D(u5_N7), .CK(clk), .Q(u5_prod1[7]) );
  DFF_X2 u5_prod_reg_7_ ( .D(u5_prod1[7]), .CK(clk), .QN(n4437) );
  DFF_X2 u5_prod1_reg_8_ ( .D(u5_N8), .CK(clk), .Q(u5_prod1[8]) );
  DFF_X2 u5_prod_reg_8_ ( .D(u5_prod1[8]), .CK(clk), .Q(prod[8]), .QN(n4703)
         );
  DFF_X2 u5_prod1_reg_9_ ( .D(u5_N9), .CK(clk), .Q(u5_prod1[9]) );
  DFF_X2 u5_prod_reg_9_ ( .D(u5_prod1[9]), .CK(clk), .QN(n4390) );
  DFF_X2 u5_prod1_reg_10_ ( .D(u5_N10), .CK(clk), .Q(u5_prod1[10]) );
  DFF_X2 u5_prod_reg_10_ ( .D(u5_prod1[10]), .CK(clk), .Q(prod[10]), .QN(n4696) );
  DFF_X2 u5_prod1_reg_11_ ( .D(u5_N11), .CK(clk), .Q(u5_prod1[11]) );
  DFF_X2 u5_prod_reg_11_ ( .D(u5_prod1[11]), .CK(clk), .Q(prod[11]), .QN(n4702) );
  DFF_X2 u5_prod1_reg_12_ ( .D(u5_N12), .CK(clk), .Q(u5_prod1[12]) );
  DFF_X2 u5_prod_reg_12_ ( .D(u5_prod1[12]), .CK(clk), .QN(n4416) );
  DFF_X2 u5_prod1_reg_13_ ( .D(u5_N13), .CK(clk), .Q(u5_prod1[13]) );
  DFF_X2 u5_prod_reg_13_ ( .D(u5_prod1[13]), .CK(clk), .QN(n4447) );
  DFF_X2 u5_prod1_reg_14_ ( .D(u5_N14), .CK(clk), .Q(u5_prod1[14]) );
  DFF_X2 u5_prod_reg_14_ ( .D(u5_prod1[14]), .CK(clk), .QN(n4396) );
  DFF_X2 u5_prod1_reg_15_ ( .D(u5_N15), .CK(clk), .Q(u5_prod1[15]) );
  DFF_X2 u5_prod_reg_15_ ( .D(u5_prod1[15]), .CK(clk), .QN(n4514) );
  DFF_X2 u5_prod1_reg_16_ ( .D(u5_N16), .CK(clk), .Q(u5_prod1[16]) );
  DFF_X2 u5_prod_reg_16_ ( .D(u5_prod1[16]), .CK(clk), .Q(prod[16]), .QN(n4711) );
  DFF_X2 u5_prod1_reg_17_ ( .D(u5_N17), .CK(clk), .Q(u5_prod1[17]) );
  DFF_X2 u5_prod_reg_17_ ( .D(u5_prod1[17]), .CK(clk), .Q(prod[17]), .QN(n4695) );
  DFF_X2 u5_prod1_reg_18_ ( .D(u5_N18), .CK(clk), .Q(u5_prod1[18]) );
  DFF_X2 u5_prod_reg_18_ ( .D(u5_prod1[18]), .CK(clk), .Q(prod[18]), .QN(n4701) );
  DFF_X2 u5_prod1_reg_19_ ( .D(u5_N19), .CK(clk), .Q(u5_prod1[19]) );
  DFF_X2 u5_prod_reg_19_ ( .D(u5_prod1[19]), .CK(clk), .QN(n4406) );
  DFF_X2 u5_prod1_reg_20_ ( .D(u5_N20), .CK(clk), .Q(u5_prod1[20]) );
  DFF_X2 u5_prod_reg_20_ ( .D(u5_prod1[20]), .CK(clk), .QN(n4507) );
  DFF_X2 u5_prod1_reg_21_ ( .D(u5_N21), .CK(clk), .Q(u5_prod1[21]) );
  DFF_X2 u5_prod_reg_21_ ( .D(u5_prod1[21]), .CK(clk), .Q(prod[21]), .QN(n4710) );
  DFF_X2 u5_prod1_reg_22_ ( .D(u5_N22), .CK(clk), .Q(u5_prod1[22]) );
  DFF_X2 u5_prod_reg_22_ ( .D(u5_prod1[22]), .CK(clk), .Q(prod[22]), .QN(n4694) );
  DFF_X2 u5_prod1_reg_23_ ( .D(u5_N23), .CK(clk), .Q(u5_prod1[23]) );
  DFF_X2 u5_prod_reg_23_ ( .D(u5_prod1[23]), .CK(clk), .Q(prod[23]), .QN(n4700) );
  DFF_X2 u5_prod1_reg_24_ ( .D(u5_N24), .CK(clk), .Q(u5_prod1[24]) );
  DFF_X2 u5_prod_reg_24_ ( .D(u5_prod1[24]), .CK(clk), .QN(n4445) );
  DFF_X2 u5_prod1_reg_25_ ( .D(u5_N25), .CK(clk), .Q(u5_prod1[25]) );
  DFF_X2 u5_prod_reg_25_ ( .D(u5_prod1[25]), .CK(clk), .QN(n4523) );
  DFF_X2 u5_prod1_reg_26_ ( .D(u5_N26), .CK(clk), .Q(u5_prod1[26]) );
  DFF_X2 u5_prod_reg_26_ ( .D(u5_prod1[26]), .CK(clk), .QN(n4397) );
  DFF_X2 u5_prod1_reg_27_ ( .D(u5_N27), .CK(clk), .Q(u5_prod1[27]) );
  DFF_X2 u5_prod_reg_27_ ( .D(u5_prod1[27]), .CK(clk), .QN(n4381) );
  DFF_X2 u5_prod1_reg_28_ ( .D(u5_N28), .CK(clk), .Q(u5_prod1[28]) );
  DFF_X2 u5_prod_reg_28_ ( .D(u5_prod1[28]), .CK(clk), .Q(prod[28]), .QN(n4709) );
  DFF_X2 u5_prod1_reg_29_ ( .D(u5_N29), .CK(clk), .Q(u5_prod1[29]) );
  DFF_X2 u5_prod_reg_29_ ( .D(u5_prod1[29]), .CK(clk), .Q(prod[29]), .QN(n4693) );
  DFF_X2 u5_prod1_reg_30_ ( .D(u5_N30), .CK(clk), .Q(u5_prod1[30]) );
  DFF_X2 u5_prod_reg_30_ ( .D(u5_prod1[30]), .CK(clk), .QN(n4386) );
  DFF_X2 u5_prod1_reg_31_ ( .D(u5_N31), .CK(clk), .Q(u5_prod1[31]) );
  DFF_X2 u5_prod_reg_31_ ( .D(u5_prod1[31]), .CK(clk), .QN(n4512) );
  DFF_X2 u5_prod1_reg_32_ ( .D(u5_N32), .CK(clk), .Q(u5_prod1[32]) );
  DFF_X2 u5_prod_reg_32_ ( .D(u5_prod1[32]), .CK(clk), .QN(n4435) );
  DFF_X2 u5_prod1_reg_33_ ( .D(u5_N33), .CK(clk), .Q(u5_prod1[33]) );
  DFF_X2 u5_prod_reg_33_ ( .D(u5_prod1[33]), .CK(clk), .Q(prod[33]), .QN(n4708) );
  DFF_X2 u5_prod1_reg_34_ ( .D(u5_N34), .CK(clk), .Q(u5_prod1[34]) );
  DFF_X2 u5_prod_reg_34_ ( .D(u5_prod1[34]), .CK(clk), .Q(prod[34]), .QN(n4692) );
  DFF_X2 u5_prod1_reg_35_ ( .D(u5_N35), .CK(clk), .Q(u5_prod1[35]) );
  DFF_X2 u5_prod_reg_35_ ( .D(u5_prod1[35]), .CK(clk), .Q(prod[35]), .QN(n4699) );
  DFF_X2 u5_prod1_reg_36_ ( .D(u5_N36), .CK(clk), .Q(u5_prod1[36]) );
  DFF_X2 u5_prod_reg_36_ ( .D(u5_prod1[36]), .CK(clk), .QN(n4443) );
  DFF_X2 u5_prod1_reg_37_ ( .D(u5_N37), .CK(clk), .Q(u5_prod1[37]) );
  DFF_X2 u5_prod_reg_37_ ( .D(u5_prod1[37]), .CK(clk), .QN(n4521) );
  DFF_X2 u5_prod1_reg_38_ ( .D(u5_N38), .CK(clk), .Q(u5_prod1[38]) );
  DFF_X2 u5_prod_reg_38_ ( .D(u5_prod1[38]), .CK(clk), .QN(n4393) );
  DFF_X2 u5_prod1_reg_39_ ( .D(u5_N39), .CK(clk), .Q(u5_prod1[39]) );
  DFF_X2 u5_prod_reg_39_ ( .D(u5_prod1[39]), .CK(clk), .QN(n4379) );
  DFF_X2 u5_prod1_reg_40_ ( .D(u5_N40), .CK(clk), .Q(u5_prod1[40]) );
  DFF_X2 u5_prod_reg_40_ ( .D(u5_prod1[40]), .CK(clk), .Q(prod[40]), .QN(n4691) );
  DFF_X2 u5_prod1_reg_41_ ( .D(u5_N41), .CK(clk), .Q(u5_prod1[41]) );
  DFF_X2 u5_prod_reg_41_ ( .D(u5_prod1[41]), .CK(clk), .Q(prod[41]), .QN(n4698) );
  DFF_X2 u5_prod1_reg_42_ ( .D(u5_N42), .CK(clk), .Q(u5_prod1[42]) );
  DFF_X2 u5_prod_reg_42_ ( .D(u5_prod1[42]), .CK(clk), .QN(n4444) );
  DFF_X2 u5_prod1_reg_43_ ( .D(u5_N43), .CK(clk), .Q(u5_prod1[43]) );
  DFF_X2 u5_prod_reg_43_ ( .D(u5_prod1[43]), .CK(clk), .QN(n4522) );
  DFF_X2 u5_prod1_reg_44_ ( .D(u5_N44), .CK(clk), .Q(u5_prod1[44]) );
  DFF_X2 u5_prod_reg_44_ ( .D(u5_prod1[44]), .CK(clk), .QN(n4394) );
  DFF_X2 u5_prod1_reg_45_ ( .D(u5_N45), .CK(clk), .Q(u5_prod1[45]) );
  DFF_X2 u5_prod_reg_45_ ( .D(u5_prod1[45]), .CK(clk), .QN(n4380) );
  DFF_X2 u5_prod1_reg_46_ ( .D(u5_N46), .CK(clk), .Q(u5_prod1[46]) );
  DFF_X2 u5_prod_reg_46_ ( .D(u5_prod1[46]), .CK(clk), .Q(prod[46]), .QN(n4707) );
  DFF_X2 u5_prod1_reg_47_ ( .D(u5_N47), .CK(clk), .Q(u5_prod1[47]) );
  DFF_X2 u5_prod_reg_47_ ( .D(u5_prod1[47]), .CK(clk), .Q(prod[47]), .QN(n4690) );
  DFF_X2 u5_prod1_reg_48_ ( .D(u5_N48), .CK(clk), .Q(u5_prod1[48]) );
  DFF_X2 u5_prod_reg_48_ ( .D(u5_prod1[48]), .CK(clk), .Q(prod[48]), .QN(n4697) );
  DFF_X2 u5_prod1_reg_49_ ( .D(u5_N49), .CK(clk), .Q(u5_prod1[49]) );
  DFF_X2 u5_prod_reg_49_ ( .D(u5_prod1[49]), .CK(clk), .QN(n4515) );
  DFF_X2 u5_prod1_reg_50_ ( .D(u5_N50), .CK(clk), .Q(u5_prod1[50]) );
  DFF_X2 u5_prod_reg_50_ ( .D(u5_prod1[50]), .CK(clk), .QN(n4395) );
  DFF_X2 u5_prod1_reg_51_ ( .D(u5_N51), .CK(clk), .Q(u5_prod1[51]) );
  DFF_X2 u5_prod_reg_51_ ( .D(u5_prod1[51]), .CK(clk), .QN(n4631) );
  DFF_X2 u5_prod1_reg_52_ ( .D(u5_N52), .CK(clk), .Q(u5_prod1[52]) );
  DFF_X2 u5_prod_reg_52_ ( .D(u5_prod1[52]), .CK(clk), .Q(prod[52]), .QN(n4706) );
  DFF_X2 u5_prod1_reg_53_ ( .D(u5_N53), .CK(clk), .Q(u5_prod1[53]) );
  DFF_X2 u5_prod_reg_53_ ( .D(u5_prod1[53]), .CK(clk), .Q(prod[53]), .QN(n4689) );
  DFF_X2 u5_prod1_reg_54_ ( .D(u5_N54), .CK(clk), .Q(u5_prod1[54]) );
  DFF_X2 u5_prod_reg_54_ ( .D(u5_prod1[54]), .CK(clk), .Q(prod[54]), .QN(n4555) );
  DFF_X2 u5_prod1_reg_55_ ( .D(u5_N55), .CK(clk), .Q(u5_prod1[55]) );
  DFF_X2 u5_prod_reg_55_ ( .D(u5_prod1[55]), .CK(clk), .QN(n4403) );
  DFF_X2 u5_prod1_reg_56_ ( .D(u5_N56), .CK(clk), .Q(u5_prod1[56]) );
  DFF_X2 u5_prod_reg_56_ ( .D(u5_prod1[56]), .CK(clk), .QN(n4510) );
  DFF_X2 u5_prod1_reg_57_ ( .D(u5_N57), .CK(clk), .Q(u5_prod1[57]) );
  DFF_X2 u5_prod_reg_57_ ( .D(u5_prod1[57]), .CK(clk), .QN(n4387) );
  DFF_X2 u5_prod1_reg_58_ ( .D(u5_N58), .CK(clk), .Q(u5_prod1[58]) );
  DFF_X2 u5_prod_reg_58_ ( .D(u5_prod1[58]), .CK(clk), .Q(prod[58]), .QN(n4562) );
  DFF_X2 u5_prod1_reg_59_ ( .D(u5_N59), .CK(clk), .Q(u5_prod1[59]) );
  DFF_X2 u5_prod_reg_59_ ( .D(u5_prod1[59]), .CK(clk), .Q(prod[59]), .QN(n4547) );
  DFF_X2 u5_prod1_reg_60_ ( .D(u5_N60), .CK(clk), .Q(u5_prod1[60]) );
  DFF_X2 u5_prod_reg_60_ ( .D(u5_prod1[60]), .CK(clk), .QN(n4415) );
  DFF_X2 u5_prod1_reg_61_ ( .D(u5_N61), .CK(clk), .Q(u5_prod1[61]) );
  DFF_X2 u5_prod_reg_61_ ( .D(u5_prod1[61]), .CK(clk), .QN(n4519) );
  DFF_X2 u5_prod1_reg_62_ ( .D(u5_N62), .CK(clk), .Q(u5_prod1[62]) );
  DFF_X2 u5_prod_reg_62_ ( .D(u5_prod1[62]), .CK(clk), .QN(n4392) );
  DFF_X2 u5_prod1_reg_63_ ( .D(u5_N63), .CK(clk), .Q(u5_prod1[63]) );
  DFF_X2 u5_prod_reg_63_ ( .D(u5_prod1[63]), .CK(clk), .QN(n4378) );
  DFF_X2 u5_prod1_reg_64_ ( .D(u5_N64), .CK(clk), .Q(u5_prod1[64]) );
  DFF_X2 u5_prod_reg_64_ ( .D(u5_prod1[64]), .CK(clk), .Q(prod[64]), .QN(n4563) );
  DFF_X2 u5_prod1_reg_65_ ( .D(u5_N65), .CK(clk), .Q(u5_prod1[65]) );
  DFF_X2 u5_prod_reg_65_ ( .D(u5_prod1[65]), .CK(clk), .Q(prod[65]), .QN(n4548) );
  DFF_X2 u5_prod1_reg_66_ ( .D(u5_N66), .CK(clk), .Q(u5_prod1[66]) );
  DFF_X2 u5_prod_reg_66_ ( .D(u5_prod1[66]), .CK(clk), .Q(prod[66]), .QN(n4556) );
  DFF_X2 u5_prod1_reg_67_ ( .D(u5_N67), .CK(clk), .Q(u5_prod1[67]) );
  DFF_X2 u5_prod_reg_67_ ( .D(u5_prod1[67]), .CK(clk), .QN(n4404) );
  DFF_X2 u5_prod1_reg_68_ ( .D(u5_N68), .CK(clk), .Q(u5_prod1[68]) );
  DFF_X2 u5_prod_reg_68_ ( .D(u5_prod1[68]), .CK(clk), .QN(n4511) );
  DFF_X2 u5_prod1_reg_69_ ( .D(u5_N69), .CK(clk), .Q(u5_prod1[69]) );
  DFF_X2 u5_prod_reg_69_ ( .D(u5_prod1[69]), .CK(clk), .QN(n4434) );
  DFF_X2 u5_prod1_reg_70_ ( .D(u5_N70), .CK(clk), .Q(u5_prod1[70]) );
  DFF_X2 u5_prod_reg_70_ ( .D(u5_prod1[70]), .CK(clk), .Q(prod[70]), .QN(n4549) );
  DFF_X2 u5_prod1_reg_71_ ( .D(u5_N71), .CK(clk), .Q(u5_prod1[71]) );
  DFF_X2 u5_prod_reg_71_ ( .D(u5_prod1[71]), .CK(clk), .Q(prod[71]), .QN(n4557) );
  DFF_X2 u5_prod1_reg_72_ ( .D(u5_N72), .CK(clk), .Q(u5_prod1[72]) );
  DFF_X2 u5_prod_reg_72_ ( .D(u5_prod1[72]), .CK(clk), .QN(n4442) );
  DFF_X2 u5_prod1_reg_73_ ( .D(u5_N73), .CK(clk), .Q(u5_prod1[73]) );
  DFF_X2 u5_prod_reg_73_ ( .D(u5_prod1[73]), .CK(clk), .QN(n4520) );
  DFF_X2 u5_prod1_reg_74_ ( .D(u5_N74), .CK(clk), .Q(u5_prod1[74]) );
  DFF_X2 u5_prod_reg_74_ ( .D(u5_prod1[74]), .CK(clk), .QN(n4413) );
  DFF_X2 u5_prod1_reg_75_ ( .D(u5_N75), .CK(clk), .Q(u5_prod1[75]) );
  DFF_X2 u5_prod_reg_75_ ( .D(u5_prod1[75]), .CK(clk), .QN(n4391) );
  DFF_X2 u5_prod1_reg_76_ ( .D(u5_N76), .CK(clk), .Q(u5_prod1[76]) );
  DFF_X2 u5_prod_reg_76_ ( .D(u5_prod1[76]), .CK(clk), .Q(prod[76]), .QN(n4564) );
  DFF_X2 u5_prod1_reg_77_ ( .D(u5_N77), .CK(clk), .Q(u5_prod1[77]) );
  DFF_X2 u5_prod_reg_77_ ( .D(u5_prod1[77]), .CK(clk), .Q(prod[77]), .QN(n4550) );
  DFF_X2 u5_prod1_reg_78_ ( .D(u5_N78), .CK(clk), .Q(u5_prod1[78]) );
  DFF_X2 u5_prod_reg_78_ ( .D(u5_prod1[78]), .CK(clk), .Q(prod[78]), .QN(n4558) );
  DFF_X2 u5_prod1_reg_79_ ( .D(u5_N79), .CK(clk), .Q(u5_prod1[79]) );
  DFF_X2 u5_prod_reg_79_ ( .D(u5_prod1[79]), .CK(clk), .QN(n4385) );
  DFF_X2 u5_prod1_reg_80_ ( .D(u5_N80), .CK(clk), .Q(u5_prod1[80]) );
  DFF_X2 u5_prod_reg_80_ ( .D(u5_prod1[80]), .CK(clk), .QN(n4506) );
  DFF_X2 u5_prod1_reg_81_ ( .D(u5_N81), .CK(clk), .Q(u5_prod1[81]) );
  DFF_X2 u5_prod_reg_81_ ( .D(u5_prod1[81]), .CK(clk), .Q(prod[81]), .QN(n4565) );
  DFF_X2 u5_prod1_reg_82_ ( .D(u5_N82), .CK(clk), .Q(u5_prod1[82]) );
  DFF_X2 u5_prod_reg_82_ ( .D(u5_prod1[82]), .CK(clk), .Q(prod[82]), .QN(n4551) );
  DFF_X2 u5_prod1_reg_83_ ( .D(u5_N83), .CK(clk), .Q(u5_prod1[83]) );
  DFF_X2 u5_prod_reg_83_ ( .D(u5_prod1[83]), .CK(clk), .Q(prod[83]), .QN(n4559) );
  DFF_X2 u5_prod1_reg_84_ ( .D(u5_N84), .CK(clk), .Q(u5_prod1[84]) );
  DFF_X2 u5_prod_reg_84_ ( .D(u5_prod1[84]), .CK(clk), .QN(n4414) );
  DFF_X2 u5_prod1_reg_85_ ( .D(u5_N85), .CK(clk), .Q(u5_prod1[85]) );
  DFF_X2 u5_prod_reg_85_ ( .D(u5_prod1[85]), .CK(clk), .QN(n4516) );
  DFF_X2 u5_prod1_reg_86_ ( .D(u5_N86), .CK(clk), .Q(u5_prod1[86]) );
  DFF_X2 u5_prod_reg_86_ ( .D(u5_prod1[86]), .CK(clk), .QN(n4439) );
  DFF_X2 u5_prod1_reg_87_ ( .D(u5_N87), .CK(clk), .Q(u5_prod1[87]) );
  DFF_X2 u5_prod_reg_87_ ( .D(u5_prod1[87]), .CK(clk), .QN(n4388) );
  DFF_X2 u5_prod1_reg_88_ ( .D(u5_N88), .CK(clk), .Q(u5_prod1[88]) );
  DFF_X2 u5_prod_reg_88_ ( .D(u5_prod1[88]), .CK(clk), .Q(prod[88]), .QN(n4566) );
  DFF_X2 u5_prod1_reg_89_ ( .D(u5_N89), .CK(clk), .Q(u5_prod1[89]) );
  DFF_X2 u5_prod_reg_89_ ( .D(u5_prod1[89]), .CK(clk), .Q(prod[89]), .QN(n4552) );
  DFF_X2 u5_prod1_reg_90_ ( .D(u5_N90), .CK(clk), .Q(u5_prod1[90]) );
  DFF_X2 u5_prod_reg_90_ ( .D(u5_prod1[90]), .CK(clk), .QN(n4440) );
  DFF_X2 u5_prod1_reg_91_ ( .D(u5_N91), .CK(clk), .Q(u5_prod1[91]) );
  DFF_X2 u5_prod_reg_91_ ( .D(u5_prod1[91]), .CK(clk), .QN(n4517) );
  DFF_X2 u5_prod1_reg_92_ ( .D(u5_N92), .CK(clk), .Q(u5_prod1[92]) );
  DFF_X2 u5_prod_reg_92_ ( .D(u5_prod1[92]), .CK(clk), .QN(n4411) );
  DFF_X2 u5_prod1_reg_93_ ( .D(u5_N93), .CK(clk), .Q(u5_prod1[93]) );
  DFF_X2 u5_prod_reg_93_ ( .D(u5_prod1[93]), .CK(clk), .QN(n4389) );
  DFF_X2 u5_prod1_reg_94_ ( .D(u5_N94), .CK(clk), .Q(u5_prod1[94]) );
  DFF_X2 u5_prod_reg_94_ ( .D(u5_prod1[94]), .CK(clk), .Q(prod[94]), .QN(n4567) );
  DFF_X2 u5_prod1_reg_95_ ( .D(u5_N95), .CK(clk), .Q(u5_prod1[95]) );
  DFF_X2 u5_prod_reg_95_ ( .D(u5_prod1[95]), .CK(clk), .Q(prod[95]), .QN(n4553) );
  DFF_X2 u5_prod1_reg_96_ ( .D(u5_N96), .CK(clk), .Q(u5_prod1[96]) );
  DFF_X2 u5_prod_reg_96_ ( .D(u5_prod1[96]), .CK(clk), .Q(prod[96]), .QN(n4560) );
  DFF_X2 u5_prod1_reg_97_ ( .D(u5_N97), .CK(clk), .Q(u5_prod1[97]) );
  DFF_X2 u5_prod_reg_97_ ( .D(u5_prod1[97]), .CK(clk), .QN(n4441) );
  DFF_X2 u5_prod1_reg_98_ ( .D(u5_N98), .CK(clk), .Q(u5_prod1[98]) );
  DFF_X2 u5_prod_reg_98_ ( .D(u5_prod1[98]), .CK(clk), .QN(n4518) );
  DFF_X2 u5_prod1_reg_99_ ( .D(u5_N99), .CK(clk), .Q(u5_prod1[99]) );
  DFF_X2 u5_prod_reg_99_ ( .D(u5_prod1[99]), .CK(clk), .QN(n4412) );
  DFF_X2 u5_prod1_reg_100_ ( .D(u5_N100), .CK(clk), .Q(u5_prod1[100]) );
  DFF_X2 u5_prod_reg_100_ ( .D(u5_prod1[100]), .CK(clk), .Q(prod[100]), .QN(
        n4554) );
  DFF_X2 u5_prod1_reg_101_ ( .D(u5_N101), .CK(clk), .Q(u5_prod1[101]) );
  DFF_X2 u5_prod_reg_101_ ( .D(u5_prod1[101]), .CK(clk), .Q(prod[101]), .QN(
        n4561) );
  DFF_X2 u5_prod1_reg_102_ ( .D(u5_N102), .CK(clk), .Q(u5_prod1[102]) );
  DFF_X2 u5_prod_reg_102_ ( .D(u5_prod1[102]), .CK(clk), .QN(n4405) );
  DFF_X2 u5_prod1_reg_103_ ( .D(u5_N103), .CK(clk), .Q(u5_prod1[103]) );
  DFF_X2 u5_prod_reg_103_ ( .D(u5_prod1[103]), .CK(clk), .QN(n4513) );
  DFF_X2 u5_prod1_reg_104_ ( .D(u5_N104), .CK(clk), .Q(u5_prod1[104]) );
  DFF_X2 u5_prod_reg_104_ ( .D(u5_prod1[104]), .CK(clk), .QN(n4436) );
  DFF_X2 u5_prod1_reg_105_ ( .D(u5_N105), .CK(clk), .Q(u5_prod1[105]) );
  DFF_X2 u5_prod_reg_105_ ( .D(u5_prod1[105]), .CK(clk), .Q(prod[105]), .QN(
        n4568) );
  DFF_X2 u6_remainder_reg_0_ ( .D(u6_N0), .CK(clk), .Q(u6_remainder[0]) );
  DFF_X2 u6_rem_reg_0_ ( .D(u6_remainder[0]), .CK(clk), .Q(remainder[0]) );
  DFF_X2 u6_remainder_reg_1_ ( .D(u6_N1), .CK(clk), .Q(u6_remainder[1]) );
  DFF_X2 u6_rem_reg_1_ ( .D(u6_remainder[1]), .CK(clk), .Q(remainder[1]) );
  DFF_X2 u6_remainder_reg_2_ ( .D(u6_N2), .CK(clk), .Q(u6_remainder[2]) );
  DFF_X2 u6_rem_reg_2_ ( .D(u6_remainder[2]), .CK(clk), .Q(remainder[2]) );
  DFF_X2 u6_remainder_reg_3_ ( .D(u6_N3), .CK(clk), .Q(u6_remainder[3]) );
  DFF_X2 u6_rem_reg_3_ ( .D(u6_remainder[3]), .CK(clk), .Q(remainder[3]) );
  DFF_X2 u6_remainder_reg_4_ ( .D(u6_N4), .CK(clk), .Q(u6_remainder[4]) );
  DFF_X2 u6_rem_reg_4_ ( .D(u6_remainder[4]), .CK(clk), .Q(remainder[4]) );
  DFF_X2 u6_remainder_reg_5_ ( .D(u6_N5), .CK(clk), .Q(u6_remainder[5]) );
  DFF_X2 u6_rem_reg_5_ ( .D(u6_remainder[5]), .CK(clk), .Q(remainder[5]) );
  DFF_X2 u6_remainder_reg_6_ ( .D(u6_N6), .CK(clk), .Q(u6_remainder[6]) );
  DFF_X2 u6_rem_reg_6_ ( .D(u6_remainder[6]), .CK(clk), .Q(remainder[6]) );
  DFF_X2 u6_remainder_reg_7_ ( .D(u6_N7), .CK(clk), .Q(u6_remainder[7]) );
  DFF_X2 u6_rem_reg_7_ ( .D(u6_remainder[7]), .CK(clk), .Q(remainder[7]) );
  DFF_X2 u6_remainder_reg_8_ ( .D(u6_N8), .CK(clk), .Q(u6_remainder[8]) );
  DFF_X2 u6_rem_reg_8_ ( .D(u6_remainder[8]), .CK(clk), .Q(remainder[8]) );
  DFF_X2 u6_remainder_reg_9_ ( .D(u6_N9), .CK(clk), .Q(u6_remainder[9]) );
  DFF_X2 u6_rem_reg_9_ ( .D(u6_remainder[9]), .CK(clk), .Q(remainder[9]) );
  DFF_X2 u6_remainder_reg_10_ ( .D(u6_N10), .CK(clk), .Q(u6_remainder[10]) );
  DFF_X2 u6_rem_reg_10_ ( .D(u6_remainder[10]), .CK(clk), .Q(remainder[10]) );
  DFF_X2 u6_remainder_reg_11_ ( .D(u6_N11), .CK(clk), .Q(u6_remainder[11]) );
  DFF_X2 u6_rem_reg_11_ ( .D(u6_remainder[11]), .CK(clk), .Q(remainder[11]) );
  DFF_X2 u6_remainder_reg_12_ ( .D(u6_N12), .CK(clk), .Q(u6_remainder[12]) );
  DFF_X2 u6_rem_reg_12_ ( .D(u6_remainder[12]), .CK(clk), .Q(remainder[12]) );
  DFF_X2 u6_remainder_reg_13_ ( .D(u6_N13), .CK(clk), .Q(u6_remainder[13]) );
  DFF_X2 u6_rem_reg_13_ ( .D(u6_remainder[13]), .CK(clk), .Q(remainder[13]) );
  DFF_X2 u6_remainder_reg_14_ ( .D(u6_N14), .CK(clk), .Q(u6_remainder[14]) );
  DFF_X2 u6_rem_reg_14_ ( .D(u6_remainder[14]), .CK(clk), .Q(remainder[14]) );
  DFF_X2 u6_remainder_reg_15_ ( .D(u6_N15), .CK(clk), .Q(u6_remainder[15]) );
  DFF_X2 u6_rem_reg_15_ ( .D(u6_remainder[15]), .CK(clk), .Q(remainder[15]) );
  DFF_X2 u6_remainder_reg_16_ ( .D(u6_N16), .CK(clk), .Q(u6_remainder[16]) );
  DFF_X2 u6_rem_reg_16_ ( .D(u6_remainder[16]), .CK(clk), .Q(remainder[16]) );
  DFF_X2 u6_remainder_reg_17_ ( .D(u6_N17), .CK(clk), .Q(u6_remainder[17]) );
  DFF_X2 u6_rem_reg_17_ ( .D(u6_remainder[17]), .CK(clk), .Q(remainder[17]) );
  DFF_X2 u6_remainder_reg_18_ ( .D(u6_N18), .CK(clk), .Q(u6_remainder[18]) );
  DFF_X2 u6_rem_reg_18_ ( .D(u6_remainder[18]), .CK(clk), .Q(remainder[18]) );
  DFF_X2 u6_remainder_reg_19_ ( .D(u6_N19), .CK(clk), .Q(u6_remainder[19]) );
  DFF_X2 u6_rem_reg_19_ ( .D(u6_remainder[19]), .CK(clk), .Q(remainder[19]) );
  DFF_X2 u6_remainder_reg_20_ ( .D(u6_N20), .CK(clk), .Q(u6_remainder[20]) );
  DFF_X2 u6_rem_reg_20_ ( .D(u6_remainder[20]), .CK(clk), .Q(remainder[20]) );
  DFF_X2 u6_remainder_reg_21_ ( .D(u6_N21), .CK(clk), .Q(u6_remainder[21]) );
  DFF_X2 u6_rem_reg_21_ ( .D(u6_remainder[21]), .CK(clk), .Q(remainder[21]) );
  DFF_X2 u6_remainder_reg_22_ ( .D(u6_N22), .CK(clk), .Q(u6_remainder[22]) );
  DFF_X2 u6_rem_reg_22_ ( .D(u6_remainder[22]), .CK(clk), .Q(remainder[22]) );
  DFF_X2 u6_remainder_reg_23_ ( .D(u6_N23), .CK(clk), .Q(u6_remainder[23]) );
  DFF_X2 u6_rem_reg_23_ ( .D(u6_remainder[23]), .CK(clk), .Q(remainder[23]) );
  DFF_X2 u6_remainder_reg_24_ ( .D(u6_N24), .CK(clk), .Q(u6_remainder[24]) );
  DFF_X2 u6_rem_reg_24_ ( .D(u6_remainder[24]), .CK(clk), .Q(remainder[24]) );
  DFF_X2 u6_remainder_reg_25_ ( .D(u6_N25), .CK(clk), .Q(u6_remainder[25]) );
  DFF_X2 u6_rem_reg_25_ ( .D(u6_remainder[25]), .CK(clk), .Q(remainder[25]) );
  DFF_X2 u6_remainder_reg_26_ ( .D(u6_N26), .CK(clk), .Q(u6_remainder[26]) );
  DFF_X2 u6_rem_reg_26_ ( .D(u6_remainder[26]), .CK(clk), .Q(remainder[26]) );
  DFF_X2 u6_remainder_reg_27_ ( .D(u6_N27), .CK(clk), .Q(u6_remainder[27]) );
  DFF_X2 u6_rem_reg_27_ ( .D(u6_remainder[27]), .CK(clk), .Q(remainder[27]) );
  DFF_X2 u6_remainder_reg_28_ ( .D(u6_N28), .CK(clk), .Q(u6_remainder[28]) );
  DFF_X2 u6_rem_reg_28_ ( .D(u6_remainder[28]), .CK(clk), .Q(remainder[28]) );
  DFF_X2 u6_remainder_reg_29_ ( .D(u6_N29), .CK(clk), .Q(u6_remainder[29]) );
  DFF_X2 u6_rem_reg_29_ ( .D(u6_remainder[29]), .CK(clk), .Q(remainder[29]) );
  DFF_X2 u6_remainder_reg_30_ ( .D(u6_N30), .CK(clk), .Q(u6_remainder[30]) );
  DFF_X2 u6_rem_reg_30_ ( .D(u6_remainder[30]), .CK(clk), .Q(remainder[30]) );
  DFF_X2 u6_remainder_reg_31_ ( .D(u6_N31), .CK(clk), .Q(u6_remainder[31]) );
  DFF_X2 u6_rem_reg_31_ ( .D(u6_remainder[31]), .CK(clk), .Q(remainder[31]) );
  DFF_X2 u6_remainder_reg_32_ ( .D(u6_N32), .CK(clk), .Q(u6_remainder[32]) );
  DFF_X2 u6_rem_reg_32_ ( .D(u6_remainder[32]), .CK(clk), .Q(remainder[32]) );
  DFF_X2 u6_remainder_reg_33_ ( .D(u6_N33), .CK(clk), .Q(u6_remainder[33]) );
  DFF_X2 u6_rem_reg_33_ ( .D(u6_remainder[33]), .CK(clk), .Q(remainder[33]) );
  DFF_X2 u6_remainder_reg_34_ ( .D(u6_N34), .CK(clk), .Q(u6_remainder[34]) );
  DFF_X2 u6_rem_reg_34_ ( .D(u6_remainder[34]), .CK(clk), .Q(remainder[34]) );
  DFF_X2 u6_remainder_reg_35_ ( .D(u6_N35), .CK(clk), .Q(u6_remainder[35]) );
  DFF_X2 u6_rem_reg_35_ ( .D(u6_remainder[35]), .CK(clk), .Q(remainder[35]) );
  DFF_X2 u6_remainder_reg_36_ ( .D(u6_N36), .CK(clk), .Q(u6_remainder[36]) );
  DFF_X2 u6_rem_reg_36_ ( .D(u6_remainder[36]), .CK(clk), .Q(remainder[36]) );
  DFF_X2 u6_remainder_reg_37_ ( .D(u6_N37), .CK(clk), .Q(u6_remainder[37]) );
  DFF_X2 u6_rem_reg_37_ ( .D(u6_remainder[37]), .CK(clk), .Q(remainder[37]) );
  DFF_X2 u6_remainder_reg_38_ ( .D(u6_N38), .CK(clk), .Q(u6_remainder[38]) );
  DFF_X2 u6_rem_reg_38_ ( .D(u6_remainder[38]), .CK(clk), .Q(remainder[38]) );
  DFF_X2 u6_remainder_reg_39_ ( .D(u6_N39), .CK(clk), .Q(u6_remainder[39]) );
  DFF_X2 u6_rem_reg_39_ ( .D(u6_remainder[39]), .CK(clk), .Q(remainder[39]) );
  DFF_X2 u6_remainder_reg_40_ ( .D(u6_N40), .CK(clk), .Q(u6_remainder[40]) );
  DFF_X2 u6_rem_reg_40_ ( .D(u6_remainder[40]), .CK(clk), .Q(remainder[40]) );
  DFF_X2 u6_remainder_reg_41_ ( .D(u6_N41), .CK(clk), .Q(u6_remainder[41]) );
  DFF_X2 u6_rem_reg_41_ ( .D(u6_remainder[41]), .CK(clk), .Q(remainder[41]) );
  DFF_X2 u6_remainder_reg_42_ ( .D(u6_N42), .CK(clk), .Q(u6_remainder[42]) );
  DFF_X2 u6_rem_reg_42_ ( .D(u6_remainder[42]), .CK(clk), .Q(remainder[42]) );
  DFF_X2 u6_remainder_reg_43_ ( .D(u6_N43), .CK(clk), .Q(u6_remainder[43]) );
  DFF_X2 u6_rem_reg_43_ ( .D(u6_remainder[43]), .CK(clk), .Q(remainder[43]) );
  DFF_X2 u6_remainder_reg_44_ ( .D(u6_N44), .CK(clk), .Q(u6_remainder[44]) );
  DFF_X2 u6_rem_reg_44_ ( .D(u6_remainder[44]), .CK(clk), .Q(remainder[44]) );
  DFF_X2 u6_remainder_reg_45_ ( .D(u6_N45), .CK(clk), .Q(u6_remainder[45]) );
  DFF_X2 u6_rem_reg_45_ ( .D(u6_remainder[45]), .CK(clk), .Q(remainder[45]) );
  DFF_X2 u6_remainder_reg_46_ ( .D(u6_N46), .CK(clk), .Q(u6_remainder[46]) );
  DFF_X2 u6_rem_reg_46_ ( .D(u6_remainder[46]), .CK(clk), .Q(remainder[46]) );
  DFF_X2 u6_remainder_reg_47_ ( .D(u6_N47), .CK(clk), .Q(u6_remainder[47]) );
  DFF_X2 u6_rem_reg_47_ ( .D(u6_remainder[47]), .CK(clk), .Q(remainder[47]) );
  DFF_X2 u6_remainder_reg_48_ ( .D(u6_N48), .CK(clk), .Q(u6_remainder[48]) );
  DFF_X2 u6_rem_reg_48_ ( .D(u6_remainder[48]), .CK(clk), .Q(remainder[48]) );
  DFF_X2 u6_remainder_reg_49_ ( .D(u6_N49), .CK(clk), .Q(u6_remainder[49]) );
  DFF_X2 u6_rem_reg_49_ ( .D(u6_remainder[49]), .CK(clk), .Q(remainder[49]) );
  DFF_X2 u6_remainder_reg_50_ ( .D(u6_N50), .CK(clk), .Q(u6_remainder[50]) );
  DFF_X2 u6_rem_reg_50_ ( .D(u6_remainder[50]), .CK(clk), .Q(remainder[50]) );
  DFF_X2 u6_remainder_reg_51_ ( .D(u6_N51), .CK(clk), .Q(u6_remainder[51]) );
  DFF_X2 u6_rem_reg_51_ ( .D(u6_remainder[51]), .CK(clk), .Q(remainder[51]) );
  DFF_X2 u6_remainder_reg_52_ ( .D(u6_N52), .CK(clk), .Q(u6_remainder[52]) );
  DFF_X2 u6_rem_reg_52_ ( .D(u6_remainder[52]), .CK(clk), .Q(remainder[52]) );
  DFF_X2 u6_remainder_reg_55_ ( .D(u6_N55), .CK(clk), .Q(u6_remainder[55]) );
  DFF_X2 u6_rem_reg_55_ ( .D(u6_remainder[55]), .CK(clk), .Q(remainder[55]) );
  DFF_X2 u6_remainder_reg_56_ ( .D(u6_N56), .CK(clk), .Q(u6_remainder[56]) );
  DFF_X2 u6_rem_reg_56_ ( .D(u6_remainder[56]), .CK(clk), .Q(remainder[56]) );
  DFF_X2 u6_remainder_reg_57_ ( .D(u6_N57), .CK(clk), .Q(u6_remainder[57]) );
  DFF_X2 u6_rem_reg_57_ ( .D(u6_remainder[57]), .CK(clk), .Q(remainder[57]) );
  DFF_X2 u6_remainder_reg_58_ ( .D(u6_N58), .CK(clk), .Q(u6_remainder[58]) );
  DFF_X2 u6_rem_reg_58_ ( .D(u6_remainder[58]), .CK(clk), .Q(remainder[58]) );
  DFF_X2 u6_remainder_reg_59_ ( .D(u6_N59), .CK(clk), .Q(u6_remainder[59]) );
  DFF_X2 u6_rem_reg_59_ ( .D(u6_remainder[59]), .CK(clk), .Q(remainder[59]) );
  DFF_X2 u6_remainder_reg_60_ ( .D(u6_N60), .CK(clk), .Q(u6_remainder[60]) );
  DFF_X2 u6_rem_reg_60_ ( .D(u6_remainder[60]), .CK(clk), .Q(remainder[60]) );
  DFF_X2 u6_remainder_reg_61_ ( .D(u6_N61), .CK(clk), .Q(u6_remainder[61]) );
  DFF_X2 u6_rem_reg_61_ ( .D(u6_remainder[61]), .CK(clk), .Q(remainder[61]) );
  DFF_X2 u6_remainder_reg_62_ ( .D(u6_N62), .CK(clk), .Q(u6_remainder[62]) );
  DFF_X2 u6_rem_reg_62_ ( .D(u6_remainder[62]), .CK(clk), .Q(remainder[62]) );
  DFF_X2 u6_remainder_reg_63_ ( .D(u6_N63), .CK(clk), .Q(u6_remainder[63]) );
  DFF_X2 u6_rem_reg_63_ ( .D(u6_remainder[63]), .CK(clk), .Q(remainder[63]) );
  DFF_X2 u6_remainder_reg_64_ ( .D(u6_N64), .CK(clk), .Q(u6_remainder[64]) );
  DFF_X2 u6_rem_reg_64_ ( .D(u6_remainder[64]), .CK(clk), .Q(remainder[64]) );
  DFF_X2 u6_remainder_reg_65_ ( .D(u6_N65), .CK(clk), .Q(u6_remainder[65]) );
  DFF_X2 u6_rem_reg_65_ ( .D(u6_remainder[65]), .CK(clk), .Q(remainder[65]) );
  DFF_X2 u6_remainder_reg_66_ ( .D(u6_N66), .CK(clk), .Q(u6_remainder[66]) );
  DFF_X2 u6_rem_reg_66_ ( .D(u6_remainder[66]), .CK(clk), .Q(remainder[66]) );
  DFF_X2 u6_remainder_reg_67_ ( .D(u6_N67), .CK(clk), .Q(u6_remainder[67]) );
  DFF_X2 u6_rem_reg_67_ ( .D(u6_remainder[67]), .CK(clk), .Q(remainder[67]) );
  DFF_X2 u6_remainder_reg_68_ ( .D(u6_N68), .CK(clk), .Q(u6_remainder[68]) );
  DFF_X2 u6_rem_reg_68_ ( .D(u6_remainder[68]), .CK(clk), .Q(remainder[68]) );
  DFF_X2 u6_remainder_reg_69_ ( .D(u6_N69), .CK(clk), .Q(u6_remainder[69]) );
  DFF_X2 u6_rem_reg_69_ ( .D(u6_remainder[69]), .CK(clk), .Q(remainder[69]) );
  DFF_X2 u6_remainder_reg_70_ ( .D(u6_N70), .CK(clk), .Q(u6_remainder[70]) );
  DFF_X2 u6_rem_reg_70_ ( .D(u6_remainder[70]), .CK(clk), .Q(remainder[70]) );
  DFF_X2 u6_remainder_reg_71_ ( .D(u6_N71), .CK(clk), .Q(u6_remainder[71]) );
  DFF_X2 u6_rem_reg_71_ ( .D(u6_remainder[71]), .CK(clk), .Q(remainder[71]) );
  DFF_X2 u6_remainder_reg_72_ ( .D(u6_N72), .CK(clk), .Q(u6_remainder[72]) );
  DFF_X2 u6_rem_reg_72_ ( .D(u6_remainder[72]), .CK(clk), .Q(remainder[72]) );
  DFF_X2 u6_remainder_reg_73_ ( .D(u6_N73), .CK(clk), .Q(u6_remainder[73]) );
  DFF_X2 u6_rem_reg_73_ ( .D(u6_remainder[73]), .CK(clk), .Q(remainder[73]) );
  DFF_X2 u6_remainder_reg_74_ ( .D(u6_N74), .CK(clk), .Q(u6_remainder[74]) );
  DFF_X2 u6_rem_reg_74_ ( .D(u6_remainder[74]), .CK(clk), .Q(remainder[74]) );
  DFF_X2 u6_remainder_reg_75_ ( .D(u6_N75), .CK(clk), .Q(u6_remainder[75]) );
  DFF_X2 u6_rem_reg_75_ ( .D(u6_remainder[75]), .CK(clk), .Q(remainder[75]) );
  DFF_X2 u6_remainder_reg_76_ ( .D(u6_N76), .CK(clk), .Q(u6_remainder[76]) );
  DFF_X2 u6_rem_reg_76_ ( .D(u6_remainder[76]), .CK(clk), .Q(remainder[76]) );
  DFF_X2 u6_remainder_reg_77_ ( .D(u6_N77), .CK(clk), .Q(u6_remainder[77]) );
  DFF_X2 u6_rem_reg_77_ ( .D(u6_remainder[77]), .CK(clk), .Q(remainder[77]) );
  DFF_X2 u6_remainder_reg_78_ ( .D(u6_N78), .CK(clk), .Q(u6_remainder[78]) );
  DFF_X2 u6_rem_reg_78_ ( .D(u6_remainder[78]), .CK(clk), .Q(remainder[78]) );
  DFF_X2 u6_remainder_reg_79_ ( .D(u6_N79), .CK(clk), .Q(u6_remainder[79]) );
  DFF_X2 u6_rem_reg_79_ ( .D(u6_remainder[79]), .CK(clk), .Q(remainder[79]) );
  DFF_X2 u6_remainder_reg_80_ ( .D(u6_N80), .CK(clk), .Q(u6_remainder[80]) );
  DFF_X2 u6_rem_reg_80_ ( .D(u6_remainder[80]), .CK(clk), .Q(remainder[80]) );
  DFF_X2 u6_remainder_reg_81_ ( .D(u6_N81), .CK(clk), .Q(u6_remainder[81]) );
  DFF_X2 u6_rem_reg_81_ ( .D(u6_remainder[81]), .CK(clk), .Q(remainder[81]) );
  DFF_X2 u6_remainder_reg_82_ ( .D(u6_N82), .CK(clk), .Q(u6_remainder[82]) );
  DFF_X2 u6_rem_reg_82_ ( .D(u6_remainder[82]), .CK(clk), .Q(remainder[82]) );
  DFF_X2 u6_remainder_reg_83_ ( .D(u6_N83), .CK(clk), .Q(u6_remainder[83]) );
  DFF_X2 u6_rem_reg_83_ ( .D(u6_remainder[83]), .CK(clk), .Q(remainder[83]) );
  DFF_X2 u6_remainder_reg_84_ ( .D(u6_N84), .CK(clk), .Q(u6_remainder[84]) );
  DFF_X2 u6_rem_reg_84_ ( .D(u6_remainder[84]), .CK(clk), .Q(remainder[84]) );
  DFF_X2 u6_remainder_reg_85_ ( .D(u6_N85), .CK(clk), .Q(u6_remainder[85]) );
  DFF_X2 u6_rem_reg_85_ ( .D(u6_remainder[85]), .CK(clk), .Q(remainder[85]) );
  DFF_X2 u6_remainder_reg_86_ ( .D(u6_N86), .CK(clk), .Q(u6_remainder[86]) );
  DFF_X2 u6_rem_reg_86_ ( .D(u6_remainder[86]), .CK(clk), .Q(remainder[86]) );
  DFF_X2 u6_remainder_reg_87_ ( .D(u6_N87), .CK(clk), .Q(u6_remainder[87]) );
  DFF_X2 u6_rem_reg_87_ ( .D(u6_remainder[87]), .CK(clk), .Q(remainder[87]) );
  DFF_X2 u6_remainder_reg_88_ ( .D(u6_N88), .CK(clk), .Q(u6_remainder[88]) );
  DFF_X2 u6_rem_reg_88_ ( .D(u6_remainder[88]), .CK(clk), .Q(remainder[88]) );
  DFF_X2 u6_remainder_reg_89_ ( .D(u6_N89), .CK(clk), .Q(u6_remainder[89]) );
  DFF_X2 u6_rem_reg_89_ ( .D(u6_remainder[89]), .CK(clk), .Q(remainder[89]) );
  DFF_X2 u6_remainder_reg_90_ ( .D(u6_N90), .CK(clk), .Q(u6_remainder[90]) );
  DFF_X2 u6_rem_reg_90_ ( .D(u6_remainder[90]), .CK(clk), .Q(remainder[90]) );
  DFF_X2 u6_remainder_reg_91_ ( .D(u6_N91), .CK(clk), .Q(u6_remainder[91]) );
  DFF_X2 u6_rem_reg_91_ ( .D(u6_remainder[91]), .CK(clk), .Q(remainder[91]) );
  DFF_X2 u6_remainder_reg_92_ ( .D(u6_N92), .CK(clk), .Q(u6_remainder[92]) );
  DFF_X2 u6_rem_reg_92_ ( .D(u6_remainder[92]), .CK(clk), .Q(remainder[92]) );
  DFF_X2 u6_remainder_reg_93_ ( .D(u6_N93), .CK(clk), .Q(u6_remainder[93]) );
  DFF_X2 u6_rem_reg_93_ ( .D(u6_remainder[93]), .CK(clk), .Q(remainder[93]) );
  DFF_X2 u6_remainder_reg_94_ ( .D(u6_N94), .CK(clk), .Q(u6_remainder[94]) );
  DFF_X2 u6_rem_reg_94_ ( .D(u6_remainder[94]), .CK(clk), .Q(remainder[94]) );
  DFF_X2 u6_remainder_reg_95_ ( .D(u6_N95), .CK(clk), .Q(u6_remainder[95]) );
  DFF_X2 u6_rem_reg_95_ ( .D(u6_remainder[95]), .CK(clk), .Q(remainder[95]) );
  DFF_X2 u6_remainder_reg_96_ ( .D(u6_N96), .CK(clk), .Q(u6_remainder[96]) );
  DFF_X2 u6_rem_reg_96_ ( .D(u6_remainder[96]), .CK(clk), .Q(remainder[96]) );
  DFF_X2 u6_remainder_reg_97_ ( .D(u6_N97), .CK(clk), .Q(u6_remainder[97]) );
  DFF_X2 u6_rem_reg_97_ ( .D(u6_remainder[97]), .CK(clk), .Q(remainder[97]) );
  DFF_X2 u6_remainder_reg_98_ ( .D(u6_N98), .CK(clk), .Q(u6_remainder[98]) );
  DFF_X2 u6_rem_reg_98_ ( .D(u6_remainder[98]), .CK(clk), .Q(remainder[98]) );
  DFF_X2 u6_remainder_reg_99_ ( .D(u6_N99), .CK(clk), .Q(u6_remainder[99]) );
  DFF_X2 u6_rem_reg_99_ ( .D(u6_remainder[99]), .CK(clk), .Q(remainder[99]) );
  DFF_X2 u6_remainder_reg_100_ ( .D(u6_N100), .CK(clk), .Q(u6_remainder[100])
         );
  DFF_X2 u6_rem_reg_100_ ( .D(u6_remainder[100]), .CK(clk), .Q(remainder[100])
         );
  DFF_X2 u6_remainder_reg_101_ ( .D(u6_N101), .CK(clk), .Q(u6_remainder[101])
         );
  DFF_X2 u6_rem_reg_101_ ( .D(u6_remainder[101]), .CK(clk), .Q(remainder[101])
         );
  DFF_X2 u6_remainder_reg_102_ ( .D(u6_N102), .CK(clk), .Q(u6_remainder[102])
         );
  DFF_X2 u6_rem_reg_102_ ( .D(u6_remainder[102]), .CK(clk), .Q(remainder[102])
         );
  DFF_X2 u6_remainder_reg_103_ ( .D(u6_N103), .CK(clk), .Q(u6_remainder[103])
         );
  DFF_X2 u6_rem_reg_103_ ( .D(u6_remainder[103]), .CK(clk), .Q(remainder[103])
         );
  DFF_X2 u6_remainder_reg_104_ ( .D(u6_N104), .CK(clk), .Q(u6_remainder[104])
         );
  DFF_X2 u6_rem_reg_104_ ( .D(u6_remainder[104]), .CK(clk), .Q(remainder[104])
         );
  DFF_X2 u6_remainder_reg_105_ ( .D(u6_N105), .CK(clk), .Q(u6_remainder[105])
         );
  DFF_X2 u6_rem_reg_105_ ( .D(u6_remainder[105]), .CK(clk), .Q(remainder[105])
         );
  DFF_X2 u6_remainder_reg_106_ ( .D(u6_N106), .CK(clk), .Q(u6_remainder[106])
         );
  DFF_X2 u6_rem_reg_106_ ( .D(u6_remainder[106]), .CK(clk), .Q(remainder[106])
         );
  DFF_X2 u6_remainder_reg_107_ ( .D(u6_N107), .CK(clk), .Q(u6_remainder[107])
         );
  DFF_X2 u6_rem_reg_107_ ( .D(u6_remainder[107]), .CK(clk), .Q(remainder[107])
         );
  DFF_X2 u6_quo1_reg_0_ ( .D(u6_N0), .CK(clk), .Q(u6_quo1[0]) );
  DFF_X2 u6_quo_reg_0_ ( .D(u6_quo1[0]), .CK(clk), .Q(quo[0]) );
  DFF_X2 u6_quo1_reg_1_ ( .D(u6_N1), .CK(clk), .Q(u6_quo1[1]) );
  DFF_X2 u6_quo_reg_1_ ( .D(u6_quo1[1]), .CK(clk), .Q(quo[1]) );
  DFF_X2 u6_quo1_reg_2_ ( .D(u6_N2), .CK(clk), .Q(u6_quo1[2]) );
  DFF_X2 u6_quo_reg_2_ ( .D(u6_quo1[2]), .CK(clk), .Q(quo[2]), .QN(n4538) );
  DLH_X2 fract_denorm_reg_0_ ( .G(n4870), .D(n4252), .Q(fract_denorm[0]) );
  DFF_X2 u6_quo1_reg_3_ ( .D(u6_N3), .CK(clk), .Q(u6_quo1[3]) );
  DFF_X2 u6_quo_reg_3_ ( .D(u6_quo1[3]), .CK(clk), .Q(quo[3]), .QN(n4539) );
  DLH_X2 fract_denorm_reg_1_ ( .G(N784), .D(N686), .Q(fract_denorm[1]) );
  DFF_X2 u6_quo1_reg_4_ ( .D(u6_N4), .CK(clk), .Q(u6_quo1[4]) );
  DFF_X2 u6_quo_reg_4_ ( .D(u6_quo1[4]), .CK(clk), .Q(quo[4]), .QN(n4537) );
  DLH_X2 fract_denorm_reg_2_ ( .G(n4870), .D(n4253), .Q(fract_denorm[2]) );
  DFF_X2 u6_quo1_reg_5_ ( .D(u6_N5), .CK(clk), .Q(u6_quo1[5]) );
  DFF_X2 u6_quo_reg_5_ ( .D(u6_quo1[5]), .CK(clk), .Q(quo[5]), .QN(n4536) );
  DLH_X2 fract_denorm_reg_3_ ( .G(n4869), .D(n4254), .Q(fract_denorm[3]) );
  DFF_X2 u6_quo1_reg_6_ ( .D(u6_N6), .CK(clk), .Q(u6_quo1[6]) );
  DFF_X2 u6_quo_reg_6_ ( .D(u6_quo1[6]), .CK(clk), .Q(quo[6]), .QN(n4540) );
  DLH_X2 fract_denorm_reg_4_ ( .G(N784), .D(N689), .Q(fract_denorm[4]) );
  DFF_X2 u6_quo1_reg_7_ ( .D(u6_N7), .CK(clk), .Q(u6_quo1[7]) );
  DFF_X2 u6_quo_reg_7_ ( .D(u6_quo1[7]), .CK(clk), .Q(quo[7]), .QN(n4535) );
  DLH_X2 fract_denorm_reg_5_ ( .G(n4870), .D(n4255), .Q(fract_denorm[5]) );
  DFF_X2 u6_quo1_reg_8_ ( .D(u6_N8), .CK(clk), .Q(u6_quo1[8]) );
  DFF_X2 u6_quo_reg_8_ ( .D(u6_quo1[8]), .CK(clk), .Q(quo[8]), .QN(n4534) );
  DLH_X2 fract_denorm_reg_6_ ( .G(n4869), .D(n4256), .Q(fract_denorm[6]) );
  DFF_X2 u6_quo1_reg_9_ ( .D(u6_N9), .CK(clk), .Q(u6_quo1[9]) );
  DFF_X2 u6_quo_reg_9_ ( .D(u6_quo1[9]), .CK(clk), .Q(quo[9]), .QN(n4541) );
  DLH_X2 fract_denorm_reg_7_ ( .G(N784), .D(N692), .Q(fract_denorm[7]) );
  DFF_X2 u6_quo1_reg_10_ ( .D(u6_N10), .CK(clk), .Q(u6_quo1[10]) );
  DFF_X2 u6_quo_reg_10_ ( .D(u6_quo1[10]), .CK(clk), .Q(quo[10]), .QN(n4533)
         );
  DLH_X2 fract_denorm_reg_8_ ( .G(n4870), .D(n4257), .Q(fract_denorm[8]) );
  DFF_X2 u6_quo1_reg_11_ ( .D(u6_N11), .CK(clk), .Q(u6_quo1[11]) );
  DFF_X2 u6_quo_reg_11_ ( .D(u6_quo1[11]), .CK(clk), .Q(quo[11]), .QN(n4542)
         );
  DLH_X2 fract_denorm_reg_9_ ( .G(n4869), .D(N694), .Q(fract_denorm[9]) );
  DFF_X2 u6_quo1_reg_12_ ( .D(u6_N12), .CK(clk), .Q(u6_quo1[12]) );
  DFF_X2 u6_quo_reg_12_ ( .D(u6_quo1[12]), .CK(clk), .Q(quo[12]), .QN(n4532)
         );
  DLH_X2 fract_denorm_reg_10_ ( .G(N784), .D(n4258), .Q(fract_denorm[10]) );
  DFF_X2 u6_quo1_reg_13_ ( .D(u6_N13), .CK(clk), .Q(u6_quo1[13]) );
  DFF_X2 u6_quo_reg_13_ ( .D(u6_quo1[13]), .CK(clk), .Q(quo[13]), .QN(n4531)
         );
  DLH_X2 fract_denorm_reg_11_ ( .G(n4870), .D(n4259), .Q(fract_denorm[11]) );
  DFF_X2 u6_quo1_reg_14_ ( .D(u6_N14), .CK(clk), .Q(u6_quo1[14]) );
  DFF_X2 u6_quo_reg_14_ ( .D(u6_quo1[14]), .CK(clk), .Q(quo[14]), .QN(n4543)
         );
  DLH_X2 fract_denorm_reg_12_ ( .G(n4869), .D(N697), .Q(fract_denorm[12]) );
  DFF_X2 u6_quo1_reg_15_ ( .D(u6_N15), .CK(clk), .Q(u6_quo1[15]) );
  DFF_X2 u6_quo_reg_15_ ( .D(u6_quo1[15]), .CK(clk), .Q(quo[15]), .QN(n4544)
         );
  DLH_X2 fract_denorm_reg_13_ ( .G(n4870), .D(N698), .Q(fract_denorm[13]) );
  DFF_X2 u6_quo1_reg_16_ ( .D(u6_N16), .CK(clk), .Q(u6_quo1[16]) );
  DFF_X2 u6_quo_reg_16_ ( .D(u6_quo1[16]), .CK(clk), .Q(quo[16]), .QN(n4545)
         );
  DLH_X2 fract_denorm_reg_14_ ( .G(N784), .D(N699), .Q(fract_denorm[14]) );
  DFF_X2 u6_quo1_reg_17_ ( .D(u6_N17), .CK(clk), .Q(u6_quo1[17]) );
  DFF_X2 u6_quo_reg_17_ ( .D(u6_quo1[17]), .CK(clk), .Q(quo[17]), .QN(n4669)
         );
  DLH_X2 fract_denorm_reg_15_ ( .G(n4869), .D(N700), .Q(fract_denorm[15]) );
  DFF_X2 u6_quo1_reg_18_ ( .D(u6_N18), .CK(clk), .Q(u6_quo1[18]) );
  DFF_X2 u6_quo_reg_18_ ( .D(u6_quo1[18]), .CK(clk), .Q(quo[18]), .QN(n4530)
         );
  DLH_X2 fract_denorm_reg_16_ ( .G(n4872), .D(n4260), .Q(fract_denorm[16]) );
  DFF_X2 u6_quo1_reg_19_ ( .D(u6_N19), .CK(clk), .Q(u6_quo1[19]) );
  DFF_X2 u6_quo_reg_19_ ( .D(u6_quo1[19]), .CK(clk), .Q(quo[19]), .QN(n4529)
         );
  DLH_X2 fract_denorm_reg_17_ ( .G(n4869), .D(n4261), .Q(fract_denorm[17]) );
  DFF_X2 u6_quo1_reg_20_ ( .D(u6_N20), .CK(clk), .Q(u6_quo1[20]) );
  DFF_X2 u6_quo_reg_20_ ( .D(u6_quo1[20]), .CK(clk), .Q(quo[20]), .QN(n4528)
         );
  DLH_X2 fract_denorm_reg_18_ ( .G(n4870), .D(n4262), .Q(fract_denorm[18]) );
  DFF_X2 u6_quo1_reg_21_ ( .D(u6_N21), .CK(clk), .Q(u6_quo1[21]) );
  DFF_X2 u6_quo_reg_21_ ( .D(u6_quo1[21]), .CK(clk), .Q(quo[21]), .QN(n4670)
         );
  DLH_X2 fract_denorm_reg_19_ ( .G(n4869), .D(N704), .Q(fract_denorm[19]) );
  DFF_X2 u6_quo1_reg_22_ ( .D(u6_N22), .CK(clk), .Q(u6_quo1[22]) );
  DFF_X2 u6_quo_reg_22_ ( .D(u6_quo1[22]), .CK(clk), .Q(quo[22]), .QN(n4671)
         );
  DLH_X2 fract_denorm_reg_20_ ( .G(N784), .D(N705), .Q(fract_denorm[20]) );
  DFF_X2 u6_quo1_reg_23_ ( .D(u6_N23), .CK(clk), .Q(u6_quo1[23]) );
  DFF_X2 u6_quo_reg_23_ ( .D(u6_quo1[23]), .CK(clk), .Q(quo[23]), .QN(n4470)
         );
  DLH_X2 fract_denorm_reg_21_ ( .G(n4870), .D(n4263), .Q(fract_denorm[21]) );
  DFF_X2 u6_quo1_reg_24_ ( .D(u6_N24), .CK(clk), .Q(u6_quo1[24]) );
  DFF_X2 u6_quo_reg_24_ ( .D(u6_quo1[24]), .CK(clk), .Q(quo[24]), .QN(n4469)
         );
  DLH_X2 fract_denorm_reg_22_ ( .G(N784), .D(n4264), .Q(fract_denorm[22]) );
  DFF_X2 u6_quo1_reg_25_ ( .D(u6_N25), .CK(clk), .Q(u6_quo1[25]) );
  DFF_X2 u6_quo_reg_25_ ( .D(u6_quo1[25]), .CK(clk), .Q(quo[25]), .QN(n4468)
         );
  DLH_X2 fract_denorm_reg_23_ ( .G(n4869), .D(n4265), .Q(fract_denorm[23]) );
  DFF_X2 u6_quo1_reg_26_ ( .D(u6_N26), .CK(clk), .Q(u6_quo1[26]) );
  DFF_X2 u6_quo_reg_26_ ( .D(u6_quo1[26]), .CK(clk), .Q(quo[26]), .QN(n4672)
         );
  DLH_X2 fract_denorm_reg_24_ ( .G(n4870), .D(N709), .Q(fract_denorm[24]) );
  DFF_X2 u6_quo1_reg_27_ ( .D(u6_N27), .CK(clk), .Q(u6_quo1[27]) );
  DFF_X2 u6_quo_reg_27_ ( .D(u6_quo1[27]), .CK(clk), .Q(quo[27]), .QN(n4673)
         );
  DLH_X2 fract_denorm_reg_25_ ( .G(N784), .D(N710), .Q(fract_denorm[25]) );
  DFF_X2 u6_quo1_reg_28_ ( .D(u6_N28), .CK(clk), .Q(u6_quo1[28]) );
  DFF_X2 u6_quo_reg_28_ ( .D(u6_quo1[28]), .CK(clk), .Q(quo[28]), .QN(n4674)
         );
  DLH_X2 fract_denorm_reg_26_ ( .G(n4869), .D(N711), .Q(fract_denorm[26]) );
  DFF_X2 u6_quo1_reg_29_ ( .D(u6_N29), .CK(clk), .Q(u6_quo1[29]) );
  DFF_X2 u6_quo_reg_29_ ( .D(u6_quo1[29]), .CK(clk), .Q(quo[29]), .QN(n4675)
         );
  DLH_X2 fract_denorm_reg_27_ ( .G(n4870), .D(N712), .Q(fract_denorm[27]) );
  DFF_X2 u6_quo1_reg_30_ ( .D(u6_N30), .CK(clk), .Q(u6_quo1[30]) );
  DFF_X2 u6_quo_reg_30_ ( .D(u6_quo1[30]), .CK(clk), .Q(quo[30]), .QN(n4467)
         );
  DLH_X2 fract_denorm_reg_28_ ( .G(n4872), .D(n4266), .Q(fract_denorm[28]) );
  DFF_X2 u6_quo1_reg_31_ ( .D(u6_N31), .CK(clk), .Q(u6_quo1[31]) );
  DFF_X2 u6_quo_reg_31_ ( .D(u6_quo1[31]), .CK(clk), .Q(quo[31]), .QN(n4423)
         );
  DLH_X2 fract_denorm_reg_29_ ( .G(n4869), .D(n4267), .Q(fract_denorm[29]) );
  DFF_X2 u6_quo1_reg_32_ ( .D(u6_N32), .CK(clk), .Q(u6_quo1[32]) );
  DFF_X2 u6_quo_reg_32_ ( .D(u6_quo1[32]), .CK(clk), .Q(quo[32]), .QN(n4676)
         );
  DLH_X2 fract_denorm_reg_30_ ( .G(N784), .D(N715), .Q(fract_denorm[30]) );
  DFF_X2 u6_quo1_reg_33_ ( .D(u6_N33), .CK(clk), .Q(u6_quo1[33]) );
  DFF_X2 u6_quo_reg_33_ ( .D(u6_quo1[33]), .CK(clk), .Q(quo[33]), .QN(n4677)
         );
  DLH_X2 fract_denorm_reg_31_ ( .G(n4872), .D(N716), .Q(fract_denorm[31]) );
  DFF_X2 u6_quo1_reg_34_ ( .D(u6_N34), .CK(clk), .Q(u6_quo1[34]) );
  DFF_X2 u6_quo_reg_34_ ( .D(u6_quo1[34]), .CK(clk), .Q(quo[34]), .QN(n4678)
         );
  DLH_X2 fract_denorm_reg_32_ ( .G(n4869), .D(N717), .Q(fract_denorm[32]) );
  DFF_X2 u6_quo1_reg_35_ ( .D(u6_N35), .CK(clk), .Q(u6_quo1[35]) );
  DFF_X2 u6_quo_reg_35_ ( .D(u6_quo1[35]), .CK(clk), .Q(quo[35]), .QN(n4466)
         );
  DLH_X2 fract_denorm_reg_33_ ( .G(n4870), .D(n4268), .Q(fract_denorm[33]) );
  DFF_X2 u6_quo1_reg_36_ ( .D(u6_N36), .CK(clk), .Q(u6_quo1[36]) );
  DFF_X2 u6_quo_reg_36_ ( .D(u6_quo1[36]), .CK(clk), .Q(quo[36]), .QN(n4465)
         );
  DLH_X2 fract_denorm_reg_34_ ( .G(n4872), .D(n4269), .Q(fract_denorm[34]) );
  DFF_X2 u6_quo1_reg_37_ ( .D(u6_N37), .CK(clk), .Q(u6_quo1[37]) );
  DFF_X2 u6_quo_reg_37_ ( .D(u6_quo1[37]), .CK(clk), .Q(quo[37]), .QN(n4464)
         );
  DLH_X2 fract_denorm_reg_35_ ( .G(n4872), .D(n4270), .Q(fract_denorm[35]) );
  DFF_X2 u6_quo1_reg_38_ ( .D(u6_N38), .CK(clk), .Q(u6_quo1[38]) );
  DFF_X2 u6_quo_reg_38_ ( .D(u6_quo1[38]), .CK(clk), .Q(quo[38]), .QN(n4679)
         );
  DLH_X2 fract_denorm_reg_36_ ( .G(n4869), .D(N721), .Q(fract_denorm[36]) );
  DFF_X2 u6_quo1_reg_39_ ( .D(u6_N39), .CK(clk), .Q(u6_quo1[39]) );
  DFF_X2 u6_quo_reg_39_ ( .D(u6_quo1[39]), .CK(clk), .Q(quo[39]), .QN(n4680)
         );
  DLH_X2 fract_denorm_reg_37_ ( .G(n4869), .D(N722), .Q(fract_denorm[37]) );
  DFF_X2 u6_quo1_reg_40_ ( .D(u6_N40), .CK(clk), .Q(u6_quo1[40]) );
  DFF_X2 u6_quo_reg_40_ ( .D(u6_quo1[40]), .CK(clk), .Q(quo[40]), .QN(n4681)
         );
  DLH_X2 fract_denorm_reg_38_ ( .G(N784), .D(N723), .Q(fract_denorm[38]) );
  DFF_X2 u6_quo1_reg_41_ ( .D(u6_N41), .CK(clk), .Q(u6_quo1[41]) );
  DFF_X2 u6_quo_reg_41_ ( .D(u6_quo1[41]), .CK(clk), .Q(quo[41]), .QN(n4682)
         );
  DLH_X2 fract_denorm_reg_39_ ( .G(n4869), .D(N724), .Q(fract_denorm[39]) );
  DFF_X2 u6_quo1_reg_42_ ( .D(u6_N42), .CK(clk), .Q(u6_quo1[42]) );
  DFF_X2 u6_quo_reg_42_ ( .D(u6_quo1[42]), .CK(clk), .Q(quo[42]), .QN(n4463)
         );
  DLH_X2 fract_denorm_reg_40_ ( .G(n4870), .D(n4271), .Q(fract_denorm[40]) );
  DFF_X2 u6_quo1_reg_43_ ( .D(u6_N43), .CK(clk), .Q(u6_quo1[43]) );
  DFF_X2 u6_quo_reg_43_ ( .D(u6_quo1[43]), .CK(clk), .Q(quo[43]), .QN(n4462)
         );
  DLH_X2 fract_denorm_reg_41_ ( .G(n4872), .D(n4272), .Q(fract_denorm[41]) );
  DFF_X2 u6_quo1_reg_44_ ( .D(u6_N44), .CK(clk), .Q(u6_quo1[44]) );
  DFF_X2 u6_quo_reg_44_ ( .D(u6_quo1[44]), .CK(clk), .Q(quo[44]), .QN(n4683)
         );
  DLH_X2 fract_denorm_reg_42_ ( .G(N784), .D(N727), .Q(fract_denorm[42]) );
  DFF_X2 u6_quo1_reg_45_ ( .D(u6_N45), .CK(clk), .Q(u6_quo1[45]) );
  DFF_X2 u6_quo_reg_45_ ( .D(u6_quo1[45]), .CK(clk), .Q(quo[45]), .QN(n4684)
         );
  DLH_X2 fract_denorm_reg_43_ ( .G(n4869), .D(N728), .Q(fract_denorm[43]) );
  DFF_X2 u6_quo1_reg_46_ ( .D(u6_N46), .CK(clk), .Q(u6_quo1[46]) );
  DFF_X2 u6_quo_reg_46_ ( .D(u6_quo1[46]), .CK(clk), .Q(quo[46]), .QN(n4685)
         );
  DLH_X2 fract_denorm_reg_44_ ( .G(N784), .D(N729), .Q(fract_denorm[44]) );
  DFF_X2 u6_quo1_reg_47_ ( .D(u6_N47), .CK(clk), .Q(u6_quo1[47]) );
  DFF_X2 u6_quo_reg_47_ ( .D(u6_quo1[47]), .CK(clk), .Q(quo[47]), .QN(n4686)
         );
  DLH_X2 fract_denorm_reg_45_ ( .G(n4870), .D(N730), .Q(fract_denorm[45]) );
  DFF_X2 u6_quo1_reg_48_ ( .D(u6_N48), .CK(clk), .Q(u6_quo1[48]) );
  DFF_X2 u6_quo_reg_48_ ( .D(u6_quo1[48]), .CK(clk), .Q(quo[48]), .QN(n4461)
         );
  DLH_X2 fract_denorm_reg_46_ ( .G(n4869), .D(n4273), .Q(fract_denorm[46]) );
  DFF_X2 u6_quo1_reg_49_ ( .D(u6_N49), .CK(clk), .Q(u6_quo1[49]) );
  DFF_X2 u6_quo_reg_49_ ( .D(u6_quo1[49]), .CK(clk), .Q(quo[49]), .QN(n4527)
         );
  DLH_X2 fract_denorm_reg_47_ ( .G(n4870), .D(n4274), .Q(fract_denorm[47]) );
  DFF_X2 u6_quo1_reg_50_ ( .D(u6_N50), .CK(clk), .Q(u6_quo1[50]) );
  DFF_X2 u6_quo_reg_50_ ( .D(u6_quo1[50]), .CK(clk), .Q(quo[50]), .QN(n4526)
         );
  DLH_X2 fract_denorm_reg_48_ ( .G(n4869), .D(n4275), .Q(fract_denorm[48]) );
  DFF_X2 u6_quo1_reg_51_ ( .D(u6_N51), .CK(clk), .Q(u6_quo1[51]) );
  DFF_X2 u6_quo_reg_51_ ( .D(u6_quo1[51]), .CK(clk), .Q(quo[51]), .QN(n4687)
         );
  DLH_X2 fract_denorm_reg_49_ ( .G(n4870), .D(N734), .Q(fract_denorm[49]) );
  DFF_X2 u6_quo1_reg_52_ ( .D(u6_N52), .CK(clk), .Q(u6_quo1[52]) );
  DFF_X2 u6_quo_reg_52_ ( .D(u6_quo1[52]), .CK(clk), .Q(quo[52]), .QN(n4688)
         );
  DLH_X2 fract_denorm_reg_50_ ( .G(n4869), .D(N735), .Q(fract_denorm[50]) );
  DLH_X2 fract_denorm_reg_51_ ( .G(n4872), .D(N736), .Q(fract_denorm[51]) );
  DLH_X2 fract_denorm_reg_52_ ( .G(n4870), .D(N737), .Q(fract_denorm[52]) );
  DFF_X2 u6_quo1_reg_55_ ( .D(u6_N55), .CK(clk), .Q(u6_quo1[55]) );
  DFF_X2 u6_quo_reg_55_ ( .D(u6_quo1[55]), .CK(clk), .Q(quo[55]), .QN(n4546)
         );
  DLH_X2 fract_denorm_reg_53_ ( .G(n4872), .D(N738), .Q(fract_denorm[53]) );
  DFF_X2 u6_quo1_reg_56_ ( .D(u6_N56), .CK(clk), .Q(u6_quo1[56]) );
  DFF_X2 u6_quo_reg_56_ ( .D(u6_quo1[56]), .CK(clk), .QN(n4715) );
  DLH_X2 fract_denorm_reg_54_ ( .G(N784), .D(N739), .Q(fract_denorm[54]) );
  DFF_X2 u6_quo1_reg_57_ ( .D(u6_N57), .CK(clk), .Q(u6_quo1[57]) );
  DFF_X2 u6_quo_reg_57_ ( .D(u6_quo1[57]), .CK(clk), .QN(n4716) );
  DLH_X2 fract_denorm_reg_55_ ( .G(n4872), .D(N740), .Q(fract_denorm[55]) );
  DFF_X2 u6_quo1_reg_58_ ( .D(u6_N58), .CK(clk), .Q(u6_quo1[58]) );
  DFF_X2 u6_quo_reg_58_ ( .D(u6_quo1[58]), .CK(clk), .QN(n4717) );
  DLH_X2 fract_denorm_reg_56_ ( .G(n4872), .D(N741), .Q(fract_denorm[56]) );
  DFF_X2 u6_quo1_reg_59_ ( .D(u6_N59), .CK(clk), .Q(u6_quo1[59]) );
  DFF_X2 u6_quo_reg_59_ ( .D(u6_quo1[59]), .CK(clk), .QN(n4718) );
  DLH_X2 fract_denorm_reg_57_ ( .G(n4872), .D(N742), .Q(fract_denorm[57]) );
  DFF_X2 u6_quo1_reg_60_ ( .D(u6_N60), .CK(clk), .Q(u6_quo1[60]) );
  DFF_X2 u6_quo_reg_60_ ( .D(u6_quo1[60]), .CK(clk), .QN(n4719) );
  DLH_X2 fract_denorm_reg_58_ ( .G(n4872), .D(N743), .Q(fract_denorm[58]) );
  DFF_X2 u6_quo1_reg_61_ ( .D(u6_N61), .CK(clk), .Q(u6_quo1[61]) );
  DFF_X2 u6_quo_reg_61_ ( .D(u6_quo1[61]), .CK(clk), .QN(n4720) );
  DLH_X2 fract_denorm_reg_59_ ( .G(n4872), .D(N744), .Q(fract_denorm[59]) );
  DFF_X2 u6_quo1_reg_62_ ( .D(u6_N62), .CK(clk), .Q(u6_quo1[62]) );
  DFF_X2 u6_quo_reg_62_ ( .D(u6_quo1[62]), .CK(clk), .QN(n4721) );
  DLH_X2 fract_denorm_reg_60_ ( .G(n4872), .D(N745), .Q(fract_denorm[60]) );
  DFF_X2 u6_quo1_reg_63_ ( .D(u6_N63), .CK(clk), .Q(u6_quo1[63]) );
  DFF_X2 u6_quo_reg_63_ ( .D(u6_quo1[63]), .CK(clk), .QN(n4722) );
  DLH_X2 fract_denorm_reg_61_ ( .G(n4872), .D(N746), .Q(fract_denorm[61]) );
  DFF_X2 u6_quo1_reg_64_ ( .D(u6_N64), .CK(clk), .Q(u6_quo1[64]) );
  DFF_X2 u6_quo_reg_64_ ( .D(u6_quo1[64]), .CK(clk), .QN(n4723) );
  DLH_X2 fract_denorm_reg_62_ ( .G(n4872), .D(N747), .Q(fract_denorm[62]) );
  DFF_X2 u6_quo1_reg_65_ ( .D(u6_N65), .CK(clk), .Q(u6_quo1[65]) );
  DFF_X2 u6_quo_reg_65_ ( .D(u6_quo1[65]), .CK(clk), .QN(n4724) );
  DLH_X2 fract_denorm_reg_63_ ( .G(n4872), .D(N748), .Q(fract_denorm[63]) );
  DFF_X2 u6_quo1_reg_66_ ( .D(u6_N66), .CK(clk), .Q(u6_quo1[66]) );
  DFF_X2 u6_quo_reg_66_ ( .D(u6_quo1[66]), .CK(clk), .QN(n4725) );
  DLH_X2 fract_denorm_reg_64_ ( .G(n4872), .D(N749), .Q(fract_denorm[64]) );
  DFF_X2 u6_quo1_reg_67_ ( .D(u6_N67), .CK(clk), .Q(u6_quo1[67]) );
  DFF_X2 u6_quo_reg_67_ ( .D(u6_quo1[67]), .CK(clk), .QN(n4726) );
  DLH_X2 fract_denorm_reg_65_ ( .G(n4872), .D(N750), .Q(fract_denorm[65]) );
  DFF_X2 u6_quo1_reg_68_ ( .D(u6_N68), .CK(clk), .Q(u6_quo1[68]) );
  DFF_X2 u6_quo_reg_68_ ( .D(u6_quo1[68]), .CK(clk), .QN(n4727) );
  DLH_X2 fract_denorm_reg_66_ ( .G(N784), .D(N751), .Q(fract_denorm[66]) );
  DFF_X2 u6_quo1_reg_69_ ( .D(u6_N69), .CK(clk), .Q(u6_quo1[69]) );
  DFF_X2 u6_quo_reg_69_ ( .D(u6_quo1[69]), .CK(clk), .QN(n4728) );
  DLH_X2 fract_denorm_reg_67_ ( .G(n4872), .D(N752), .Q(fract_denorm[67]) );
  DFF_X2 u6_quo1_reg_70_ ( .D(u6_N70), .CK(clk), .Q(u6_quo1[70]) );
  DFF_X2 u6_quo_reg_70_ ( .D(u6_quo1[70]), .CK(clk), .QN(n4729) );
  DLH_X2 fract_denorm_reg_68_ ( .G(n4870), .D(N753), .Q(fract_denorm[68]) );
  DFF_X2 u6_quo1_reg_71_ ( .D(u6_N71), .CK(clk), .Q(u6_quo1[71]) );
  DFF_X2 u6_quo_reg_71_ ( .D(u6_quo1[71]), .CK(clk), .QN(n4730) );
  DLH_X2 fract_denorm_reg_69_ ( .G(n4869), .D(N754), .Q(fract_denorm[69]) );
  DFF_X2 u6_quo1_reg_72_ ( .D(u6_N72), .CK(clk), .Q(u6_quo1[72]) );
  DFF_X2 u6_quo_reg_72_ ( .D(u6_quo1[72]), .CK(clk), .QN(n4731) );
  DLH_X2 fract_denorm_reg_70_ ( .G(N784), .D(N755), .Q(fract_denorm[70]) );
  DFF_X2 u6_quo1_reg_73_ ( .D(u6_N73), .CK(clk), .Q(u6_quo1[73]) );
  DFF_X2 u6_quo_reg_73_ ( .D(u6_quo1[73]), .CK(clk), .QN(n4732) );
  DLH_X2 fract_denorm_reg_71_ ( .G(n4872), .D(N756), .Q(fract_denorm[71]) );
  DFF_X2 u6_quo1_reg_74_ ( .D(u6_N74), .CK(clk), .Q(u6_quo1[74]) );
  DFF_X2 u6_quo_reg_74_ ( .D(u6_quo1[74]), .CK(clk), .QN(n4733) );
  DLH_X2 fract_denorm_reg_72_ ( .G(n4870), .D(N757), .Q(fract_denorm[72]) );
  DFF_X2 u6_quo1_reg_75_ ( .D(u6_N75), .CK(clk), .Q(u6_quo1[75]) );
  DFF_X2 u6_quo_reg_75_ ( .D(u6_quo1[75]), .CK(clk), .QN(n4734) );
  DLH_X2 fract_denorm_reg_73_ ( .G(n4870), .D(N758), .Q(fract_denorm[73]) );
  DFF_X2 u6_quo1_reg_76_ ( .D(u6_N76), .CK(clk), .Q(u6_quo1[76]) );
  DFF_X2 u6_quo_reg_76_ ( .D(u6_quo1[76]), .CK(clk), .QN(n4735) );
  DLH_X2 fract_denorm_reg_74_ ( .G(n4869), .D(N759), .Q(fract_denorm[74]) );
  DFF_X2 u6_quo1_reg_77_ ( .D(u6_N77), .CK(clk), .Q(u6_quo1[77]) );
  DFF_X2 u6_quo_reg_77_ ( .D(u6_quo1[77]), .CK(clk), .QN(n4736) );
  DLH_X2 fract_denorm_reg_75_ ( .G(N784), .D(N760), .Q(fract_denorm[75]) );
  DFF_X2 u6_quo1_reg_78_ ( .D(u6_N78), .CK(clk), .Q(u6_quo1[78]) );
  DFF_X2 u6_quo_reg_78_ ( .D(u6_quo1[78]), .CK(clk), .QN(n4737) );
  DLH_X2 fract_denorm_reg_76_ ( .G(n4872), .D(N761), .Q(fract_denorm[76]) );
  DFF_X2 u6_quo1_reg_79_ ( .D(u6_N79), .CK(clk), .Q(u6_quo1[79]) );
  DFF_X2 u6_quo_reg_79_ ( .D(u6_quo1[79]), .CK(clk), .QN(n4738) );
  DLH_X2 fract_denorm_reg_77_ ( .G(n4869), .D(N762), .Q(fract_denorm[77]) );
  DFF_X2 u6_quo1_reg_80_ ( .D(u6_N80), .CK(clk), .Q(u6_quo1[80]) );
  DFF_X2 u6_quo_reg_80_ ( .D(u6_quo1[80]), .CK(clk), .QN(n4739) );
  DLH_X2 fract_denorm_reg_78_ ( .G(N784), .D(N763), .Q(fract_denorm[78]) );
  DFF_X2 u6_quo1_reg_81_ ( .D(u6_N81), .CK(clk), .Q(u6_quo1[81]) );
  DFF_X2 u6_quo_reg_81_ ( .D(u6_quo1[81]), .CK(clk), .QN(n4740) );
  DLH_X2 fract_denorm_reg_79_ ( .G(n4870), .D(N764), .Q(fract_denorm[79]) );
  DFF_X2 u6_quo1_reg_82_ ( .D(u6_N82), .CK(clk), .Q(u6_quo1[82]) );
  DFF_X2 u6_quo_reg_82_ ( .D(u6_quo1[82]), .CK(clk), .QN(n4741) );
  DLH_X2 fract_denorm_reg_80_ ( .G(n4872), .D(N765), .Q(fract_denorm[80]) );
  DFF_X2 u6_quo1_reg_83_ ( .D(u6_N83), .CK(clk), .Q(u6_quo1[83]) );
  DFF_X2 u6_quo_reg_83_ ( .D(u6_quo1[83]), .CK(clk), .QN(n4742) );
  DLH_X2 fract_denorm_reg_81_ ( .G(N784), .D(N766), .Q(fract_denorm[81]) );
  DFF_X2 u6_quo1_reg_84_ ( .D(u6_N84), .CK(clk), .Q(u6_quo1[84]) );
  DFF_X2 u6_quo_reg_84_ ( .D(u6_quo1[84]), .CK(clk), .QN(n4743) );
  DLH_X2 fract_denorm_reg_82_ ( .G(n4869), .D(N767), .Q(fract_denorm[82]) );
  DFF_X2 u6_quo1_reg_85_ ( .D(u6_N85), .CK(clk), .Q(u6_quo1[85]) );
  DFF_X2 u6_quo_reg_85_ ( .D(u6_quo1[85]), .CK(clk), .QN(n4744) );
  DLH_X2 fract_denorm_reg_83_ ( .G(n4869), .D(N768), .Q(fract_denorm[83]) );
  DFF_X2 u6_quo1_reg_86_ ( .D(u6_N86), .CK(clk), .Q(u6_quo1[86]) );
  DFF_X2 u6_quo_reg_86_ ( .D(u6_quo1[86]), .CK(clk), .QN(n4745) );
  DLH_X2 fract_denorm_reg_84_ ( .G(n4869), .D(N769), .Q(fract_denorm[84]) );
  DFF_X2 u6_quo1_reg_87_ ( .D(u6_N87), .CK(clk), .Q(u6_quo1[87]) );
  DFF_X2 u6_quo_reg_87_ ( .D(u6_quo1[87]), .CK(clk), .QN(n4746) );
  DLH_X2 fract_denorm_reg_85_ ( .G(n4870), .D(N770), .Q(fract_denorm[85]) );
  DFF_X2 u6_quo1_reg_88_ ( .D(u6_N88), .CK(clk), .Q(u6_quo1[88]) );
  DFF_X2 u6_quo_reg_88_ ( .D(u6_quo1[88]), .CK(clk), .QN(n4747) );
  DLH_X2 fract_denorm_reg_86_ ( .G(n4872), .D(N771), .Q(fract_denorm[86]) );
  DFF_X2 u6_quo1_reg_89_ ( .D(u6_N89), .CK(clk), .Q(u6_quo1[89]) );
  DFF_X2 u6_quo_reg_89_ ( .D(u6_quo1[89]), .CK(clk), .QN(n4748) );
  DLH_X2 fract_denorm_reg_87_ ( .G(N784), .D(N772), .Q(fract_denorm[87]) );
  DFF_X2 u6_quo1_reg_90_ ( .D(u6_N90), .CK(clk), .Q(u6_quo1[90]) );
  DFF_X2 u6_quo_reg_90_ ( .D(u6_quo1[90]), .CK(clk), .QN(n4749) );
  DLH_X2 fract_denorm_reg_88_ ( .G(n4870), .D(N773), .Q(fract_denorm[88]) );
  DFF_X2 u6_quo1_reg_91_ ( .D(u6_N91), .CK(clk), .Q(u6_quo1[91]) );
  DFF_X2 u6_quo_reg_91_ ( .D(u6_quo1[91]), .CK(clk), .QN(n4750) );
  DLH_X2 fract_denorm_reg_89_ ( .G(n4872), .D(N774), .Q(fract_denorm[89]) );
  DFF_X2 u6_quo1_reg_92_ ( .D(u6_N92), .CK(clk), .Q(u6_quo1[92]) );
  DFF_X2 u6_quo_reg_92_ ( .D(u6_quo1[92]), .CK(clk), .QN(n4751) );
  DLH_X2 fract_denorm_reg_90_ ( .G(n4869), .D(N775), .Q(fract_denorm[90]) );
  DFF_X2 u6_quo1_reg_93_ ( .D(u6_N93), .CK(clk), .Q(u6_quo1[93]) );
  DFF_X2 u6_quo_reg_93_ ( .D(u6_quo1[93]), .CK(clk), .QN(n4752) );
  DLH_X2 fract_denorm_reg_91_ ( .G(N784), .D(N776), .Q(fract_denorm[91]) );
  DFF_X2 u6_quo1_reg_94_ ( .D(u6_N94), .CK(clk), .Q(u6_quo1[94]) );
  DFF_X2 u6_quo_reg_94_ ( .D(u6_quo1[94]), .CK(clk), .QN(n4753) );
  DLH_X2 fract_denorm_reg_92_ ( .G(n4870), .D(N777), .Q(fract_denorm[92]) );
  DFF_X2 u6_quo1_reg_95_ ( .D(u6_N95), .CK(clk), .Q(u6_quo1[95]) );
  DFF_X2 u6_quo_reg_95_ ( .D(u6_quo1[95]), .CK(clk), .QN(n4754) );
  DLH_X2 fract_denorm_reg_93_ ( .G(n4872), .D(N778), .Q(fract_denorm[93]) );
  DFF_X2 u6_quo1_reg_96_ ( .D(u6_N96), .CK(clk), .Q(u6_quo1[96]) );
  DFF_X2 u6_quo_reg_96_ ( .D(u6_quo1[96]), .CK(clk), .QN(n4755) );
  DLH_X2 fract_denorm_reg_94_ ( .G(n4869), .D(N779), .Q(fract_denorm[94]) );
  DFF_X2 u6_quo1_reg_97_ ( .D(u6_N97), .CK(clk), .Q(u6_quo1[97]) );
  DFF_X2 u6_quo_reg_97_ ( .D(u6_quo1[97]), .CK(clk), .QN(n4756) );
  DLH_X2 fract_denorm_reg_95_ ( .G(n4870), .D(N780), .Q(fract_denorm[95]) );
  DFF_X2 u6_quo1_reg_98_ ( .D(u6_N98), .CK(clk), .Q(u6_quo1[98]) );
  DFF_X2 u6_quo_reg_98_ ( .D(u6_quo1[98]), .CK(clk), .QN(n4757) );
  DLH_X2 fract_denorm_reg_96_ ( .G(n4872), .D(N781), .Q(fract_denorm[96]) );
  DFF_X2 u6_quo1_reg_99_ ( .D(u6_N99), .CK(clk), .Q(u6_quo1[99]) );
  DFF_X2 u6_quo_reg_99_ ( .D(u6_quo1[99]), .CK(clk), .QN(n4758) );
  DLH_X2 fract_denorm_reg_97_ ( .G(n4869), .D(N782), .Q(fract_denorm[97]) );
  DFF_X2 u6_quo1_reg_100_ ( .D(u6_N100), .CK(clk), .Q(u6_quo1[100]) );
  DFF_X2 u6_quo_reg_100_ ( .D(u6_quo1[100]), .CK(clk), .QN(n4759) );
  DLH_X2 fract_denorm_reg_98_ ( .G(N784), .D(N783), .Q(fract_denorm[98]) );
  DFF_X2 u6_quo1_reg_101_ ( .D(u6_N101), .CK(clk), .Q(u6_quo1[101]) );
  DFF_X2 u6_quo_reg_101_ ( .D(u6_quo1[101]), .CK(clk), .QN(n4760) );
  DLH_X2 fract_denorm_reg_99_ ( .G(N784), .D(N785), .Q(fract_denorm[99]) );
  DFF_X2 u6_quo1_reg_102_ ( .D(u6_N102), .CK(clk), .Q(u6_quo1[102]) );
  DFF_X2 u6_quo_reg_102_ ( .D(u6_quo1[102]), .CK(clk), .QN(n4761) );
  DLH_X2 fract_denorm_reg_100_ ( .G(n4870), .D(N786), .Q(fract_denorm[100]) );
  DFF_X2 u6_quo1_reg_103_ ( .D(u6_N103), .CK(clk), .Q(u6_quo1[103]) );
  DFF_X2 u6_quo_reg_103_ ( .D(u6_quo1[103]), .CK(clk), .QN(n4762) );
  DLH_X2 fract_denorm_reg_101_ ( .G(N784), .D(N787), .Q(fract_denorm[101]) );
  DFF_X2 u6_quo1_reg_104_ ( .D(u6_N104), .CK(clk), .Q(u6_quo1[104]) );
  DFF_X2 u6_quo_reg_104_ ( .D(u6_quo1[104]), .CK(clk), .QN(n4763) );
  DLH_X2 fract_denorm_reg_102_ ( .G(n4870), .D(N788), .Q(fract_denorm[102]) );
  DFF_X2 u6_quo1_reg_105_ ( .D(u6_N105), .CK(clk), .Q(u6_quo1[105]) );
  DFF_X2 u6_quo_reg_105_ ( .D(u6_quo1[105]), .CK(clk), .QN(n4764) );
  DLH_X2 fract_denorm_reg_103_ ( .G(N784), .D(N789), .Q(fract_denorm[103]) );
  DFF_X2 u6_quo1_reg_106_ ( .D(u6_N106), .CK(clk), .Q(u6_quo1[106]) );
  DFF_X2 u6_quo_reg_106_ ( .D(u6_quo1[106]), .CK(clk), .QN(n4765) );
  DLH_X2 fract_denorm_reg_104_ ( .G(n4870), .D(N790), .Q(fract_denorm[104]) );
  DFF_X2 u6_quo1_reg_107_ ( .D(u6_N107), .CK(clk), .Q(u6_quo1[107]) );
  DFF_X2 u6_quo_reg_107_ ( .D(u6_quo1[107]), .CK(clk), .QN(n4766) );
  DLH_X2 fract_denorm_reg_105_ ( .G(N784), .D(N791), .Q(fract_denorm[105]) );
  DFF_X2 out_reg_52_ ( .D(N850), .CK(clk), .Q(out[52]) );
  DFF_X2 out_reg_55_ ( .D(N853), .CK(clk), .Q(out[55]) );
  DFF_X2 out_reg_56_ ( .D(N854), .CK(clk), .Q(out[56]) );
  DFF_X2 out_reg_54_ ( .D(N852), .CK(clk), .Q(out[54]) );
  DFF_X2 out_reg_57_ ( .D(N855), .CK(clk), .Q(out[57]) );
  DFF_X2 out_reg_59_ ( .D(N857), .CK(clk), .Q(out[59]) );
  DFF_X2 out_reg_58_ ( .D(N856), .CK(clk), .Q(out[58]) );
  DFF_X2 out_reg_53_ ( .D(N851), .CK(clk), .Q(out[53]) );
  DFF_X2 out_reg_62_ ( .D(N860), .CK(clk), .Q(out[62]) );
  DFF_X2 out_reg_61_ ( .D(N859), .CK(clk), .Q(out[61]) );
  DFF_X2 out_reg_60_ ( .D(N858), .CK(clk), .Q(out[60]) );
  DFF_X2 overflow_reg ( .D(N904), .CK(clk), .Q(overflow) );
  DFF_X2 out_reg_51_ ( .D(N849), .CK(clk), .Q(out[51]) );
  DFF_X2 out_reg_50_ ( .D(N848), .CK(clk), .Q(out[50]) );
  DFF_X2 out_reg_49_ ( .D(N847), .CK(clk), .Q(out[49]) );
  DFF_X2 out_reg_48_ ( .D(N846), .CK(clk), .Q(out[48]) );
  DFF_X2 out_reg_47_ ( .D(N845), .CK(clk), .Q(out[47]) );
  DFF_X2 out_reg_46_ ( .D(N844), .CK(clk), .Q(out[46]) );
  DFF_X2 out_reg_45_ ( .D(N843), .CK(clk), .Q(out[45]) );
  DFF_X2 out_reg_44_ ( .D(N842), .CK(clk), .Q(out[44]) );
  DFF_X2 out_reg_43_ ( .D(N841), .CK(clk), .Q(out[43]) );
  DFF_X2 out_reg_42_ ( .D(N840), .CK(clk), .Q(out[42]) );
  DFF_X2 out_reg_41_ ( .D(N839), .CK(clk), .Q(out[41]) );
  DFF_X2 out_reg_40_ ( .D(N838), .CK(clk), .Q(out[40]) );
  DFF_X2 out_reg_39_ ( .D(N837), .CK(clk), .Q(out[39]) );
  DFF_X2 out_reg_38_ ( .D(N836), .CK(clk), .Q(out[38]) );
  DFF_X2 out_reg_37_ ( .D(N835), .CK(clk), .Q(out[37]) );
  DFF_X2 out_reg_36_ ( .D(N834), .CK(clk), .Q(out[36]) );
  DFF_X2 out_reg_35_ ( .D(N833), .CK(clk), .Q(out[35]) );
  DFF_X2 out_reg_34_ ( .D(N832), .CK(clk), .Q(out[34]) );
  DFF_X2 out_reg_33_ ( .D(N831), .CK(clk), .Q(out[33]) );
  DFF_X2 out_reg_32_ ( .D(N830), .CK(clk), .Q(out[32]) );
  DFF_X2 out_reg_31_ ( .D(N829), .CK(clk), .Q(out[31]) );
  DFF_X2 out_reg_30_ ( .D(N828), .CK(clk), .Q(out[30]) );
  DFF_X2 out_reg_29_ ( .D(N827), .CK(clk), .Q(out[29]) );
  DFF_X2 out_reg_28_ ( .D(N826), .CK(clk), .Q(out[28]) );
  DFF_X2 out_reg_27_ ( .D(N825), .CK(clk), .Q(out[27]) );
  DFF_X2 out_reg_26_ ( .D(N824), .CK(clk), .Q(out[26]) );
  DFF_X2 out_reg_25_ ( .D(N823), .CK(clk), .Q(out[25]) );
  DFF_X2 out_reg_24_ ( .D(N822), .CK(clk), .Q(out[24]) );
  DFF_X2 out_reg_23_ ( .D(N821), .CK(clk), .Q(out[23]) );
  DFF_X2 out_reg_22_ ( .D(N820), .CK(clk), .Q(out[22]) );
  DFF_X2 out_reg_21_ ( .D(N819), .CK(clk), .Q(out[21]) );
  DFF_X2 out_reg_20_ ( .D(N818), .CK(clk), .Q(out[20]) );
  DFF_X2 out_reg_19_ ( .D(N817), .CK(clk), .Q(out[19]) );
  DFF_X2 out_reg_18_ ( .D(N816), .CK(clk), .Q(out[18]) );
  DFF_X2 out_reg_17_ ( .D(N815), .CK(clk), .Q(out[17]) );
  DFF_X2 out_reg_16_ ( .D(N814), .CK(clk), .Q(out[16]) );
  DFF_X2 out_reg_15_ ( .D(N813), .CK(clk), .Q(out[15]) );
  DFF_X2 out_reg_14_ ( .D(N812), .CK(clk), .Q(out[14]) );
  DFF_X2 out_reg_13_ ( .D(N811), .CK(clk), .Q(out[13]) );
  DFF_X2 out_reg_12_ ( .D(N810), .CK(clk), .Q(out[12]) );
  DFF_X2 out_reg_11_ ( .D(N809), .CK(clk), .Q(out[11]) );
  DFF_X2 out_reg_10_ ( .D(N808), .CK(clk), .Q(out[10]) );
  DFF_X2 out_reg_9_ ( .D(N807), .CK(clk), .Q(out[9]) );
  DFF_X2 out_reg_8_ ( .D(N806), .CK(clk), .Q(out[8]) );
  DFF_X2 out_reg_7_ ( .D(N805), .CK(clk), .Q(out[7]) );
  DFF_X2 out_reg_6_ ( .D(N804), .CK(clk), .Q(out[6]) );
  DFF_X2 out_reg_5_ ( .D(N803), .CK(clk), .Q(out[5]) );
  DFF_X2 out_reg_4_ ( .D(N802), .CK(clk), .Q(out[4]) );
  DFF_X2 out_reg_3_ ( .D(N801), .CK(clk), .Q(out[3]) );
  DFF_X2 out_reg_2_ ( .D(N800), .CK(clk), .Q(out[2]) );
  DFF_X2 out_reg_1_ ( .D(N799), .CK(clk), .Q(out[1]) );
  DFF_X2 ine_reg ( .D(N894), .CK(clk), .Q(ine) );
  DFF_X2 zero_reg ( .D(N916), .CK(clk), .Q(zero) );
  DFF_X2 out_reg_63_ ( .D(N880), .CK(clk), .Q(out[63]) );
  DFF_X2 inf_reg ( .D(N911), .CK(clk), .Q(inf) );
  DFF_X2 underflow_reg ( .D(N907), .CK(clk), .Q(underflow) );
  DFF_X2 out_reg_0_ ( .D(N798), .CK(clk), .Q(out[0]) );
  DFF_X2 exp_r_reg_0_ ( .D(n2666), .CK(clk), .QN(n4400) );
  DFF_X2 exp_r_reg_1_ ( .D(n2665), .CK(clk), .Q(n4368), .QN(n4588) );
  DFF_X2 exp_r_reg_2_ ( .D(n2664), .CK(clk), .Q(exp_r[2]), .QN(n4425) );
  DFF_X2 exp_r_reg_3_ ( .D(n2663), .CK(clk), .Q(exp_r[3]), .QN(n4473) );
  DFF_X2 exp_r_reg_4_ ( .D(n2662), .CK(clk), .Q(n4399), .QN(n4424) );
  DFF_X2 exp_r_reg_5_ ( .D(n2661), .CK(clk), .Q(n4370), .QN(n4477) );
  DFF_X2 exp_r_reg_6_ ( .D(n2660), .CK(clk), .Q(n4382), .QN(n4571) );
  DFF_X2 exp_r_reg_7_ ( .D(n2659), .CK(clk), .Q(n4359), .QN(n4475) );
  DFF_X2 exp_r_reg_8_ ( .D(n2658), .CK(clk), .Q(n4369), .QN(n4474) );
  DFF_X2 exp_r_reg_9_ ( .D(n2657), .CK(clk), .Q(n4428), .QN(n4476) );
  DFF_X2 exp_r_reg_10_ ( .D(n2656), .CK(clk), .Q(exp_r[10]), .QN(n4587) );
  OAI211_X2 U3 ( .C1(n205), .C2(n206), .A(n207), .B(n208), .ZN(
        u4_shift_right[9]) );
  AOI22_X2 U4 ( .A1(u4_div_shft2[9]), .A2(n209), .B1(u4_exp_in_mi1_9_), .B2(
        n6387), .ZN(n208) );
  AOI22_X2 U5 ( .A1(u4_div_shft3_9_), .A2(n211), .B1(u4_div_shft4[9]), .B2(
        n212), .ZN(n207) );
  OAI211_X2 U6 ( .C1(n4949), .C2(n206), .A(n214), .B(n215), .ZN(
        u4_shift_right[8]) );
  AOI22_X2 U7 ( .A1(u4_div_shft2[8]), .A2(n209), .B1(u4_exp_in_mi1_8_), .B2(
        n6387), .ZN(n215) );
  AOI22_X2 U8 ( .A1(u4_div_shft3_8_), .A2(n211), .B1(u4_div_shft4[8]), .B2(
        n212), .ZN(n214) );
  OAI211_X2 U9 ( .C1(n216), .C2(n206), .A(n217), .B(n218), .ZN(
        u4_shift_right[7]) );
  AOI22_X2 U10 ( .A1(u4_div_shft2[7]), .A2(n209), .B1(u4_exp_in_mi1_7_), .B2(
        n6387), .ZN(n218) );
  AOI22_X2 U11 ( .A1(u4_div_shft3_7_), .A2(n211), .B1(u4_div_shft4[7]), .B2(
        n212), .ZN(n217) );
  OAI211_X2 U12 ( .C1(n4945), .C2(n206), .A(n220), .B(n221), .ZN(
        u4_shift_right[6]) );
  AOI22_X2 U13 ( .A1(u4_div_shft2[6]), .A2(n209), .B1(u4_exp_in_mi1_6_), .B2(
        n6387), .ZN(n221) );
  AOI22_X2 U14 ( .A1(u4_div_shft3_6_), .A2(n211), .B1(u4_div_shft4[6]), .B2(
        n212), .ZN(n220) );
  OAI211_X2 U15 ( .C1(n222), .C2(n206), .A(n223), .B(n224), .ZN(
        u4_shift_right[5]) );
  AOI22_X2 U16 ( .A1(u4_div_shft2[5]), .A2(n209), .B1(u4_exp_in_mi1_5_), .B2(
        n6387), .ZN(n224) );
  AOI22_X2 U17 ( .A1(u4_div_shft3_5_), .A2(n211), .B1(u4_div_shft4[5]), .B2(
        n212), .ZN(n223) );
  OAI211_X2 U18 ( .C1(n225), .C2(n206), .A(n226), .B(n227), .ZN(
        u4_shift_right[4]) );
  AOI22_X2 U19 ( .A1(u4_div_shft2[4]), .A2(n209), .B1(u4_exp_in_mi1_4_), .B2(
        n6387), .ZN(n227) );
  AOI22_X2 U20 ( .A1(u4_div_shft3_4_), .A2(n211), .B1(u4_div_shft4[4]), .B2(
        n212), .ZN(n226) );
  OAI211_X2 U21 ( .C1(n228), .C2(n206), .A(n229), .B(n230), .ZN(
        u4_shift_right[3]) );
  AOI22_X2 U22 ( .A1(u4_div_shft2[3]), .A2(n209), .B1(u4_exp_in_mi1_3_), .B2(
        n6387), .ZN(n230) );
  AOI22_X2 U23 ( .A1(u4_div_shft3_3_), .A2(n211), .B1(u4_div_shft4[3]), .B2(
        n212), .ZN(n229) );
  INV_X4 U24 ( .A(u4_exp_out_3_), .ZN(n228) );
  OAI211_X2 U25 ( .C1(n231), .C2(n206), .A(n232), .B(n233), .ZN(
        u4_shift_right[2]) );
  AOI22_X2 U26 ( .A1(u4_div_shft2[2]), .A2(n209), .B1(u4_exp_in_mi1_2_), .B2(
        n6387), .ZN(n233) );
  AOI22_X2 U27 ( .A1(u4_div_shft3_2_), .A2(n211), .B1(u4_div_shft4[2]), .B2(
        n212), .ZN(n232) );
  INV_X4 U28 ( .A(u4_exp_out_2_), .ZN(n231) );
  OAI211_X2 U29 ( .C1(n234), .C2(n206), .A(n235), .B(n236), .ZN(
        u4_shift_right[1]) );
  AOI22_X2 U30 ( .A1(n4588), .A2(n209), .B1(u4_exp_in_mi1_1_), .B2(n6387), 
        .ZN(n236) );
  AOI22_X2 U31 ( .A1(u4_div_shft3_1_), .A2(n211), .B1(u4_div_shft4[1]), .B2(
        n212), .ZN(n235) );
  INV_X4 U32 ( .A(u4_exp_out_1_), .ZN(n234) );
  OAI211_X2 U33 ( .C1(u4_N6891), .C2(n206), .A(n237), .B(n238), .ZN(
        u4_shift_right[10]) );
  AOI22_X2 U34 ( .A1(u4_div_shft2[10]), .A2(n209), .B1(u4_exp_in_mi1_10_), 
        .B2(n6387), .ZN(n238) );
  AOI22_X2 U35 ( .A1(u4_div_shft3_10_), .A2(n211), .B1(u4_div_shft4[10]), .B2(
        n212), .ZN(n237) );
  OAI211_X2 U36 ( .C1(u4_exp_out_mi1[0]), .C2(n206), .A(n239), .B(n240), .ZN(
        u4_shift_right[0]) );
  AOI22_X2 U37 ( .A1(n4823), .A2(n209), .B1(n4400), .B2(n6387), .ZN(n240) );
  AOI22_X2 U95 ( .A1(u4_div_shft3_0_), .A2(n211), .B1(u4_div_shft4[0]), .B2(
        n212), .ZN(n239) );
  OAI211_X2 U99 ( .C1(n249), .C2(n6521), .A(n251), .B(n252), .ZN(
        u4_shift_left[8]) );
  AOI22_X2 U100 ( .A1(n4369), .A2(n253), .B1(u4_f2i_shft_8_), .B2(n6390), .ZN(
        n252) );
  NAND2_X2 U101 ( .A1(u4_div_scht1a[8]), .A2(n255), .ZN(n251) );
  OAI211_X2 U102 ( .C1(n249), .C2(n6522), .A(n257), .B(n258), .ZN(
        u4_shift_left[7]) );
  AOI22_X2 U103 ( .A1(n4359), .A2(n253), .B1(u4_f2i_shft_7_), .B2(n6390), .ZN(
        n258) );
  NAND2_X2 U104 ( .A1(u4_div_scht1a[7]), .A2(n255), .ZN(n257) );
  NAND2_X2 U105 ( .A1(n259), .A2(n260), .ZN(u4_shift_left[6]) );
  AOI22_X2 U107 ( .A1(n4382), .A2(n253), .B1(u4_f2i_shft_6_), .B2(n6390), .ZN(
        n259) );
  NAND2_X2 U108 ( .A1(n263), .A2(n264), .ZN(u4_shift_left[5]) );
  AOI22_X2 U110 ( .A1(n4370), .A2(n253), .B1(u4_f2i_shft_5_), .B2(n6390), .ZN(
        n263) );
  OAI211_X2 U111 ( .C1(n249), .C2(n6523), .A(n266), .B(n267), .ZN(
        u4_shift_left[4]) );
  AOI22_X2 U113 ( .A1(div_opa_ldz_r2[4]), .A2(n268), .B1(u4_fi_ldz_4_), .B2(
        n261), .ZN(n266) );
  OAI211_X2 U114 ( .C1(n249), .C2(n6524), .A(n270), .B(n271), .ZN(
        u4_shift_left[3]) );
  AOI22_X2 U116 ( .A1(div_opa_ldz_r2[3]), .A2(n268), .B1(u4_fi_ldz_3_), .B2(
        n261), .ZN(n270) );
  OAI211_X2 U117 ( .C1(n249), .C2(n6525), .A(n273), .B(n274), .ZN(
        u4_shift_left[2]) );
  AOI22_X2 U119 ( .A1(div_opa_ldz_r2[2]), .A2(n268), .B1(u4_fi_ldz_2_), .B2(
        n261), .ZN(n273) );
  NAND2_X2 U120 ( .A1(n275), .A2(n276), .ZN(u4_shift_left[1]) );
  AOI221_X2 U121 ( .B1(div_opa_ldz_r2[1]), .B2(n268), .C1(u4_fi_ldz_1_), .C2(
        n261), .A(n277), .ZN(n276) );
  OAI211_X2 U125 ( .C1(n249), .C2(n4823), .A(n286), .B(n287), .ZN(
        u4_shift_left[0]) );
  AOI22_X2 U128 ( .A1(div_opa_ldz_r2[0]), .A2(n268), .B1(u4_fi_ldz_2a_0_), 
        .B2(n261), .ZN(n286) );
  OAI221_X2 U129 ( .B1(n4818), .B2(n289), .C1(n281), .C2(n290), .A(n291), .ZN(
        n261) );
  AND3_X2 U132 ( .A1(n6527), .A2(n4822), .A3(n295), .ZN(n268) );
  INV_X4 U133 ( .A(n262), .ZN(n249) );
  AOI221_X2 U137 ( .B1(n304), .B2(fract_denorm[74]), .C1(fract_denorm[67]), 
        .C2(n305), .A(n306), .ZN(n303) );
  OAI22_X2 U138 ( .A1(n307), .A2(n308), .B1(n309), .B2(n310), .ZN(n306) );
  NOR4_X2 U143 ( .A1(n324), .A2(n325), .A3(n326), .A4(n327), .ZN(n323) );
  OAI221_X2 U144 ( .B1(n328), .B2(n329), .C1(n330), .C2(n331), .A(n332), .ZN(
        n324) );
  OAI222_X2 U149 ( .A1(n345), .A2(n312), .B1(n346), .B2(n6503), .C1(n348), 
        .C2(n349), .ZN(n343) );
  OAI211_X2 U150 ( .C1(n350), .C2(n351), .A(n352), .B(n353), .ZN(n342) );
  NAND4_X2 U151 ( .A1(fract_denorm[90]), .A2(n354), .A3(n6506), .A4(n6507), 
        .ZN(n353) );
  OAI211_X2 U155 ( .C1(fract_denorm[105]), .C2(n358), .A(n6455), .B(n360), 
        .ZN(n301) );
  NOR4_X2 U156 ( .A1(n361), .A2(n362), .A3(n363), .A4(n364), .ZN(n360) );
  OAI22_X2 U158 ( .A1(n366), .A2(n367), .B1(n368), .B2(n369), .ZN(n365) );
  AOI221_X2 U159 ( .B1(n370), .B2(n371), .C1(n372), .C2(fract_denorm[58]), .A(
        n6464), .ZN(n358) );
  OAI221_X2 U166 ( .B1(n387), .B2(n6428), .C1(n6409), .C2(n390), .A(n391), 
        .ZN(n385) );
  OAI211_X2 U168 ( .C1(n394), .C2(n6514), .A(n396), .B(n397), .ZN(n384) );
  AOI22_X2 U169 ( .A1(fract_denorm[82]), .A2(n6497), .B1(fract_denorm[66]), 
        .B2(n6479), .ZN(n397) );
  AOI221_X2 U175 ( .B1(fract_denorm[22]), .B2(n6434), .C1(fract_denorm[38]), 
        .C2(n6448), .A(n411), .ZN(n409) );
  AOI221_X2 U179 ( .B1(fract_denorm[70]), .B2(n315), .C1(fract_denorm[86]), 
        .C2(n416), .A(n417), .ZN(n412) );
  OAI211_X2 U184 ( .C1(n421), .C2(n6440), .A(n6420), .B(n424), .ZN(n386) );
  AND4_X2 U186 ( .A1(n6460), .A2(n6459), .A3(n6461), .A4(fract_denorm[46]), 
        .ZN(n427) );
  NAND4_X2 U194 ( .A1(n406), .A2(n6405), .A3(n437), .A4(n438), .ZN(
        u4_fi_ldz_1_) );
  AOI221_X2 U195 ( .B1(fract_denorm[8]), .B2(n439), .C1(n440), .C2(n4874), .A(
        n441), .ZN(n438) );
  NAND4_X2 U199 ( .A1(n6518), .A2(n6519), .A3(n447), .A4(n448), .ZN(n440) );
  OAI221_X2 U207 ( .B1(fract_denorm[105]), .B2(n455), .C1(n368), .C2(n6460), 
        .A(n456), .ZN(n405) );
  NAND2_X2 U210 ( .A1(n6427), .A2(n6428), .ZN(n462) );
  NOR4_X2 U213 ( .A1(fract_denorm[66]), .A2(fract_denorm[65]), .A3(n308), .A4(
        n6477), .ZN(n467) );
  NOR4_X2 U215 ( .A1(fract_denorm[82]), .A2(fract_denorm[81]), .A3(n400), .A4(
        n6494), .ZN(n466) );
  NOR4_X2 U217 ( .A1(n6416), .A2(n404), .A3(n471), .A4(n472), .ZN(n406) );
  OR4_X2 U218 ( .A1(n6481), .A2(n364), .A3(n327), .A4(n325), .ZN(n472) );
  AND4_X2 U220 ( .A1(fract_denorm[84]), .A2(n416), .A3(n346), .A4(n4874), .ZN(
        n327) );
  NOR4_X2 U221 ( .A1(n6467), .A2(n6469), .A3(fract_denorm[105]), .A4(
        fract_denorm[53]), .ZN(n364) );
  NAND4_X2 U223 ( .A1(fract_denorm[68]), .A2(n319), .A3(n315), .A4(n4874), 
        .ZN(n298) );
  OAI22_X2 U224 ( .A1(n6446), .A2(n393), .B1(n390), .B2(n478), .ZN(n471) );
  OAI221_X2 U225 ( .B1(n6456), .B2(n480), .C1(fract_denorm[105]), .C2(n481), 
        .A(n482), .ZN(n404) );
  AOI22_X2 U226 ( .A1(fract_denorm[12]), .A2(n337), .B1(fract_denorm[28]), 
        .B2(n333), .ZN(n482) );
  NAND2_X2 U230 ( .A1(n6458), .A2(n6457), .ZN(n480) );
  AND4_X2 U233 ( .A1(n490), .A2(n437), .A3(n486), .A4(n408), .ZN(n489) );
  AND3_X2 U250 ( .A1(n401), .A2(n4874), .A3(fract_denorm[51]), .ZN(n362) );
  OAI211_X2 U251 ( .C1(n349), .C2(n6498), .A(n510), .B(n511), .ZN(n508) );
  NAND4_X2 U252 ( .A1(fract_denorm[99]), .A2(n418), .A3(n6518), .A4(n6519), 
        .ZN(n511) );
  NAND4_X2 U254 ( .A1(n512), .A2(n513), .A3(n514), .A4(n515), .ZN(n403) );
  NAND4_X2 U255 ( .A1(fract_denorm[43]), .A2(n6458), .A3(n6456), .A4(n6457), 
        .ZN(n515) );
  AND4_X2 U267 ( .A1(n523), .A2(n524), .A3(n6423), .A4(n525), .ZN(n437) );
  NOR4_X2 U268 ( .A1(n363), .A2(n326), .A3(n6484), .A4(n527), .ZN(n525) );
  NOR4_X2 U269 ( .A1(fract_denorm[25]), .A2(fract_denorm[24]), .A3(n331), .A4(
        n6433), .ZN(n527) );
  NAND4_X2 U272 ( .A1(fract_denorm[71]), .A2(n313), .A3(n529), .A4(n4874), 
        .ZN(n297) );
  NOR4_X2 U273 ( .A1(n6502), .A2(n454), .A3(fract_denorm[105]), .A4(
        fract_denorm[88]), .ZN(n326) );
  OAI221_X2 U278 ( .B1(fract_denorm[105]), .B2(n533), .C1(n329), .C2(n6424), 
        .A(n535), .ZN(n532) );
  AOI221_X2 U282 ( .B1(fract_denorm[79]), .B2(n6495), .C1(fract_denorm[63]), 
        .C2(n6478), .A(n540), .ZN(n533) );
  NAND2_X2 U286 ( .A1(fract_denorm[7]), .A2(n6413), .ZN(n523) );
  AND3_X2 U287 ( .A1(n6408), .A2(n6420), .A3(n545), .ZN(n490) );
  AOI22_X2 U288 ( .A1(fract_denorm[73]), .A2(n313), .B1(fract_denorm[89]), 
        .B2(n357), .ZN(n545) );
  OAI221_X2 U290 ( .B1(fract_denorm[105]), .B2(n547), .C1(n366), .C2(n6457), 
        .A(n548), .ZN(n546) );
  NOR4_X2 U294 ( .A1(fract_denorm[15]), .A2(fract_denorm[14]), .A3(n329), .A4(
        n6421), .ZN(n549) );
  NOR4_X2 U298 ( .A1(fract_denorm[79]), .A2(fract_denorm[78]), .A3(n351), .A4(
        n6491), .ZN(n555) );
  NOR4_X2 U300 ( .A1(fract_denorm[63]), .A2(fract_denorm[62]), .A3(n310), .A4(
        n6474), .ZN(n554) );
  OAI221_X2 U305 ( .B1(fract_denorm[105]), .B2(n561), .C1(n461), .C2(n6443), 
        .A(n563), .ZN(n560) );
  NAND2_X2 U308 ( .A1(n335), .A2(n6429), .ZN(n387) );
  AND2_X2 U309 ( .A1(fract_denorm[49]), .A2(n566), .ZN(n361) );
  NAND2_X2 U313 ( .A1(n6499), .A2(n6498), .ZN(n400) );
  AOI221_X2 U323 ( .B1(n576), .B2(n6519), .C1(fract_denorm[25]), .C2(n6436), 
        .A(n6451), .ZN(n487) );
  AOI22_X2 U325 ( .A1(n370), .A2(fract_denorm[57]), .B1(n6452), .B2(
        fract_denorm[41]), .ZN(n579) );
  AOI22_X2 U330 ( .A1(n584), .A2(n585), .B1(n586), .B2(n587), .ZN(n581) );
  NOR4_X2 U331 ( .A1(n588), .A2(n6091), .A3(u2_N16), .A4(n4815), .ZN(n587) );
  NOR4_X2 U333 ( .A1(n591), .A2(n6093), .A3(n6097), .A4(n6095), .ZN(n586) );
  NOR4_X2 U335 ( .A1(n595), .A2(n6101), .A3(n6103), .A4(n6102), .ZN(n585) );
  AND4_X2 U337 ( .A1(n600), .A2(u2_N27), .A3(u2_N25), .A4(u2_N26), .ZN(n584)
         );
  AND3_X2 U338 ( .A1(u2_N23), .A2(u2_N22), .A3(u2_N24), .ZN(n600) );
  OAI221_X2 U339 ( .B1(u6_N52), .B2(n4350), .C1(n4825), .C2(n4349), .A(n601), 
        .ZN(u2_underflow_d[1]) );
  AOI22_X2 U341 ( .A1(n6373), .A2(n4350), .B1(n4826), .B2(n4349), .ZN(n583) );
  AND3_X2 U342 ( .A1(n602), .A2(n6352), .A3(u2_N111), .ZN(u2_underflow_d[0])
         );
  OAI22_X2 U343 ( .A1(n4815), .A2(n6093), .B1(n4817), .B2(n6101), .ZN(
        u2_exp_tmp1_3_) );
  OAI22_X2 U346 ( .A1(n4815), .A2(n6095), .B1(n4817), .B2(n6102), .ZN(
        u2_exp_tmp1_2_) );
  OAI22_X2 U349 ( .A1(n4815), .A2(n6097), .B1(n4817), .B2(n6103), .ZN(
        u2_exp_tmp1_1_) );
  OR3_X2 U353 ( .A1(n608), .A2(n4817), .A3(n4487), .ZN(n606) );
  NAND2_X2 U354 ( .A1(n4817), .A2(n4487), .ZN(n605) );
  NAND2_X2 U355 ( .A1(n610), .A2(n611), .ZN(u2_N86) );
  AOI22_X2 U357 ( .A1(u2_N64), .A2(n615), .B1(n616), .B2(n6083), .ZN(n610) );
  NAND2_X2 U358 ( .A1(n617), .A2(n618), .ZN(u2_N85) );
  AOI22_X2 U360 ( .A1(u2_N63), .A2(n615), .B1(n616), .B2(n6085), .ZN(n617) );
  NAND2_X2 U361 ( .A1(n619), .A2(n620), .ZN(u2_N84) );
  AOI22_X2 U363 ( .A1(u2_N62), .A2(n615), .B1(n616), .B2(n6086), .ZN(n619) );
  NAND2_X2 U364 ( .A1(n621), .A2(n622), .ZN(u2_N83) );
  AOI22_X2 U366 ( .A1(u2_N61), .A2(n615), .B1(n616), .B2(n6087), .ZN(n621) );
  NAND2_X2 U367 ( .A1(n623), .A2(n624), .ZN(u2_N82) );
  AOI22_X2 U369 ( .A1(u2_N60), .A2(n615), .B1(n616), .B2(n6088), .ZN(n623) );
  NAND2_X2 U370 ( .A1(n625), .A2(n626), .ZN(u2_N81) );
  AOI22_X2 U372 ( .A1(u2_N59), .A2(n615), .B1(n616), .B2(n6089), .ZN(n625) );
  NAND2_X2 U373 ( .A1(n627), .A2(n628), .ZN(u2_N80) );
  AOI22_X2 U375 ( .A1(u2_N58), .A2(n615), .B1(n616), .B2(n6090), .ZN(n627) );
  NAND2_X2 U376 ( .A1(n629), .A2(n630), .ZN(u2_N79) );
  AOI22_X2 U378 ( .A1(u2_N57), .A2(n615), .B1(n616), .B2(n6092), .ZN(n629) );
  NAND2_X2 U379 ( .A1(n631), .A2(n632), .ZN(u2_N78) );
  AOI22_X2 U381 ( .A1(u2_N56), .A2(n615), .B1(n616), .B2(n6094), .ZN(n631) );
  NAND2_X2 U382 ( .A1(n633), .A2(n634), .ZN(u2_N77) );
  AOI22_X2 U384 ( .A1(u2_N55), .A2(n615), .B1(n616), .B2(n6096), .ZN(n633) );
  NAND2_X2 U385 ( .A1(n635), .A2(n636), .ZN(u2_N76) );
  AOI22_X2 U391 ( .A1(u2_N54), .A2(n615), .B1(n616), .B2(n6098), .ZN(n635) );
  NAND2_X2 U393 ( .A1(n608), .A2(n638), .ZN(u2_exp_ovf_d_1_) );
  NAND4_X2 U394 ( .A1(n6083), .A2(n4815), .A3(n4592), .A4(n4487), .ZN(n638) );
  OAI22_X2 U396 ( .A1(u2_N41), .A2(n4815), .B1(u2_N53), .B2(n4817), .ZN(n608)
         );
  AND2_X2 U398 ( .A1(opb_r[63]), .A2(opa_r[63]), .ZN(u2_N121) );
  NAND2_X2 U400 ( .A1(u2_N113), .A2(n4815), .ZN(n640) );
  NAND2_X2 U401 ( .A1(n6373), .A2(n4592), .ZN(n639) );
  OAI22_X2 U402 ( .A1(n4856), .A2(n4666), .B1(n642), .B2(n4861), .ZN(u1_sign_d) );
  XOR2_X2 U403 ( .A(opb_r[63]), .B(n4620), .Z(n642) );
  OAI22_X2 U405 ( .A1(n4861), .A2(n644), .B1(n4867), .B2(n645), .ZN(
        u1_fractb_s[9]) );
  OAI22_X2 U406 ( .A1(n4861), .A2(n646), .B1(n4867), .B2(n647), .ZN(
        u1_fractb_s[8]) );
  OAI22_X2 U407 ( .A1(n4861), .A2(n648), .B1(n4867), .B2(n649), .ZN(
        u1_fractb_s[7]) );
  OAI22_X2 U408 ( .A1(n4861), .A2(n650), .B1(n4857), .B2(n651), .ZN(
        u1_fractb_s[6]) );
  OAI22_X2 U409 ( .A1(n4861), .A2(n652), .B1(n4857), .B2(n653), .ZN(
        u1_fractb_s[5]) );
  OAI22_X2 U410 ( .A1(n4861), .A2(n654), .B1(n4857), .B2(n655), .ZN(
        u1_fractb_s[55]) );
  OAI22_X2 U411 ( .A1(n4861), .A2(n656), .B1(n4857), .B2(n657), .ZN(
        u1_fractb_s[54]) );
  OAI22_X2 U412 ( .A1(n4861), .A2(n658), .B1(n4857), .B2(n659), .ZN(
        u1_fractb_s[53]) );
  OAI22_X2 U413 ( .A1(n4860), .A2(n660), .B1(n4857), .B2(n661), .ZN(
        u1_fractb_s[52]) );
  OAI22_X2 U414 ( .A1(n4861), .A2(n662), .B1(n4857), .B2(n663), .ZN(
        u1_fractb_s[51]) );
  OAI22_X2 U415 ( .A1(n4860), .A2(n664), .B1(n4857), .B2(n665), .ZN(
        u1_fractb_s[50]) );
  OAI22_X2 U416 ( .A1(n4860), .A2(n666), .B1(n4857), .B2(n667), .ZN(
        u1_fractb_s[4]) );
  OAI22_X2 U417 ( .A1(n4860), .A2(n668), .B1(n4857), .B2(n669), .ZN(
        u1_fractb_s[49]) );
  OAI22_X2 U418 ( .A1(n4860), .A2(n670), .B1(n4856), .B2(n671), .ZN(
        u1_fractb_s[48]) );
  OAI22_X2 U419 ( .A1(n4860), .A2(n672), .B1(n4856), .B2(n673), .ZN(
        u1_fractb_s[47]) );
  OAI22_X2 U420 ( .A1(n4860), .A2(n674), .B1(n4856), .B2(n675), .ZN(
        u1_fractb_s[46]) );
  OAI22_X2 U421 ( .A1(n4860), .A2(n676), .B1(n4856), .B2(n677), .ZN(
        u1_fractb_s[45]) );
  OAI22_X2 U422 ( .A1(n4860), .A2(n678), .B1(n4856), .B2(n679), .ZN(
        u1_fractb_s[44]) );
  OAI22_X2 U423 ( .A1(n4860), .A2(n680), .B1(n4856), .B2(n681), .ZN(
        u1_fractb_s[43]) );
  OAI22_X2 U424 ( .A1(n4860), .A2(n682), .B1(n4856), .B2(n683), .ZN(
        u1_fractb_s[42]) );
  OAI22_X2 U425 ( .A1(n4860), .A2(n684), .B1(n4856), .B2(n685), .ZN(
        u1_fractb_s[41]) );
  OAI22_X2 U426 ( .A1(n4860), .A2(n686), .B1(n4856), .B2(n687), .ZN(
        u1_fractb_s[40]) );
  OAI22_X2 U427 ( .A1(n4860), .A2(n688), .B1(n4856), .B2(n689), .ZN(
        u1_fractb_s[3]) );
  OAI22_X2 U428 ( .A1(n4860), .A2(n690), .B1(n4866), .B2(n691), .ZN(
        u1_fractb_s[39]) );
  OAI22_X2 U429 ( .A1(n4860), .A2(n692), .B1(n4866), .B2(n693), .ZN(
        u1_fractb_s[38]) );
  OAI22_X2 U430 ( .A1(n4860), .A2(n694), .B1(n4866), .B2(n695), .ZN(
        u1_fractb_s[37]) );
  OAI22_X2 U431 ( .A1(n4860), .A2(n696), .B1(n4866), .B2(n697), .ZN(
        u1_fractb_s[36]) );
  OAI22_X2 U432 ( .A1(n4860), .A2(n698), .B1(n4866), .B2(n699), .ZN(
        u1_fractb_s[35]) );
  OAI22_X2 U433 ( .A1(n4859), .A2(n700), .B1(n4866), .B2(n701), .ZN(
        u1_fractb_s[34]) );
  OAI22_X2 U434 ( .A1(n4859), .A2(n702), .B1(n4866), .B2(n703), .ZN(
        u1_fractb_s[33]) );
  OAI22_X2 U435 ( .A1(n4859), .A2(n704), .B1(n4866), .B2(n705), .ZN(
        u1_fractb_s[32]) );
  OAI22_X2 U436 ( .A1(n4859), .A2(n706), .B1(n4866), .B2(n707), .ZN(
        u1_fractb_s[31]) );
  OAI22_X2 U437 ( .A1(n4859), .A2(n708), .B1(n4866), .B2(n709), .ZN(
        u1_fractb_s[30]) );
  OAI22_X2 U438 ( .A1(n4855), .A2(n710), .B1(n4861), .B2(n711), .ZN(
        u1_fractb_s[2]) );
  OAI22_X2 U439 ( .A1(n4859), .A2(n712), .B1(n4867), .B2(n713), .ZN(
        u1_fractb_s[29]) );
  OAI22_X2 U440 ( .A1(n4859), .A2(n714), .B1(n4867), .B2(n715), .ZN(
        u1_fractb_s[28]) );
  OAI22_X2 U441 ( .A1(n4859), .A2(n716), .B1(n4867), .B2(n717), .ZN(
        u1_fractb_s[27]) );
  OAI22_X2 U442 ( .A1(n4859), .A2(n718), .B1(n4867), .B2(n719), .ZN(
        u1_fractb_s[26]) );
  OAI22_X2 U443 ( .A1(n4859), .A2(n720), .B1(n4866), .B2(n721), .ZN(
        u1_fractb_s[25]) );
  OAI22_X2 U444 ( .A1(n4859), .A2(n722), .B1(n4867), .B2(n723), .ZN(
        u1_fractb_s[24]) );
  OAI22_X2 U445 ( .A1(n4859), .A2(n724), .B1(n4867), .B2(n725), .ZN(
        u1_fractb_s[23]) );
  OAI22_X2 U446 ( .A1(n4859), .A2(n726), .B1(n4867), .B2(n727), .ZN(
        u1_fractb_s[22]) );
  OAI22_X2 U447 ( .A1(n4859), .A2(n728), .B1(n4867), .B2(n729), .ZN(
        u1_fractb_s[21]) );
  OAI22_X2 U448 ( .A1(n4859), .A2(n730), .B1(n4867), .B2(n731), .ZN(
        u1_fractb_s[20]) );
  OAI22_X2 U449 ( .A1(n4854), .A2(n732), .B1(n4861), .B2(n733), .ZN(
        u1_fractb_s[1]) );
  OAI22_X2 U450 ( .A1(n4859), .A2(n734), .B1(n4867), .B2(n735), .ZN(
        u1_fractb_s[19]) );
  OAI22_X2 U451 ( .A1(n4859), .A2(n736), .B1(n4867), .B2(n737), .ZN(
        u1_fractb_s[18]) );
  OAI22_X2 U452 ( .A1(n4859), .A2(n738), .B1(n4867), .B2(n739), .ZN(
        u1_fractb_s[17]) );
  OAI22_X2 U453 ( .A1(n4859), .A2(n740), .B1(n4867), .B2(n741), .ZN(
        u1_fractb_s[16]) );
  OAI22_X2 U454 ( .A1(n4859), .A2(n742), .B1(n4867), .B2(n743), .ZN(
        u1_fractb_s[15]) );
  OAI22_X2 U455 ( .A1(n4858), .A2(n744), .B1(n4867), .B2(n745), .ZN(
        u1_fractb_s[14]) );
  OAI22_X2 U456 ( .A1(n4858), .A2(n746), .B1(n4867), .B2(n747), .ZN(
        u1_fractb_s[13]) );
  OAI22_X2 U457 ( .A1(n4858), .A2(n748), .B1(n4867), .B2(n749), .ZN(
        u1_fractb_s[12]) );
  OAI22_X2 U458 ( .A1(n4858), .A2(n750), .B1(n4854), .B2(n751), .ZN(
        u1_fractb_s[11]) );
  OAI22_X2 U459 ( .A1(n4858), .A2(n752), .B1(n4855), .B2(n753), .ZN(
        u1_fractb_s[10]) );
  OAI22_X2 U460 ( .A1(n4865), .A2(n754), .B1(n4861), .B2(n755), .ZN(
        u1_fractb_s[0]) );
  OAI22_X2 U461 ( .A1(n4865), .A2(n644), .B1(n4861), .B2(n645), .ZN(
        u1_fracta_s[9]) );
  OAI22_X2 U462 ( .A1(n4865), .A2(n646), .B1(n4861), .B2(n647), .ZN(
        u1_fracta_s[8]) );
  OAI22_X2 U463 ( .A1(n4865), .A2(n648), .B1(n4861), .B2(n649), .ZN(
        u1_fracta_s[7]) );
  OAI22_X2 U464 ( .A1(n4865), .A2(n650), .B1(n4861), .B2(n651), .ZN(
        u1_fracta_s[6]) );
  OAI22_X2 U465 ( .A1(n4865), .A2(n652), .B1(n4861), .B2(n653), .ZN(
        u1_fracta_s[5]) );
  OAI22_X2 U466 ( .A1(n4865), .A2(n654), .B1(n4861), .B2(n655), .ZN(
        u1_fracta_s[55]) );
  OAI22_X2 U467 ( .A1(n4865), .A2(n656), .B1(n4861), .B2(n657), .ZN(
        u1_fracta_s[54]) );
  OAI22_X2 U468 ( .A1(n4865), .A2(n658), .B1(n4862), .B2(n659), .ZN(
        u1_fracta_s[53]) );
  OAI22_X2 U469 ( .A1(n4865), .A2(n660), .B1(n4862), .B2(n661), .ZN(
        u1_fracta_s[52]) );
  OAI22_X2 U470 ( .A1(n4865), .A2(n662), .B1(n4862), .B2(n663), .ZN(
        u1_fracta_s[51]) );
  OAI22_X2 U471 ( .A1(n4855), .A2(n664), .B1(n4862), .B2(n665), .ZN(
        u1_fracta_s[50]) );
  OAI22_X2 U472 ( .A1(n4855), .A2(n666), .B1(n4862), .B2(n667), .ZN(
        u1_fracta_s[4]) );
  OAI22_X2 U473 ( .A1(n4855), .A2(n668), .B1(n4862), .B2(n669), .ZN(
        u1_fracta_s[49]) );
  OAI22_X2 U474 ( .A1(n4855), .A2(n670), .B1(n4862), .B2(n671), .ZN(
        u1_fracta_s[48]) );
  OAI22_X2 U475 ( .A1(n4855), .A2(n672), .B1(n4862), .B2(n673), .ZN(
        u1_fracta_s[47]) );
  OAI22_X2 U476 ( .A1(n4855), .A2(n674), .B1(n4862), .B2(n675), .ZN(
        u1_fracta_s[46]) );
  OAI22_X2 U477 ( .A1(n4855), .A2(n676), .B1(n4862), .B2(n677), .ZN(
        u1_fracta_s[45]) );
  OAI22_X2 U478 ( .A1(n4855), .A2(n678), .B1(n4862), .B2(n679), .ZN(
        u1_fracta_s[44]) );
  OAI22_X2 U479 ( .A1(n4855), .A2(n680), .B1(n4862), .B2(n681), .ZN(
        u1_fracta_s[43]) );
  OAI22_X2 U480 ( .A1(n4855), .A2(n682), .B1(n4862), .B2(n683), .ZN(
        u1_fracta_s[42]) );
  OAI22_X2 U481 ( .A1(n4855), .A2(n684), .B1(n4862), .B2(n685), .ZN(
        u1_fracta_s[41]) );
  OAI22_X2 U482 ( .A1(n4854), .A2(n686), .B1(n4862), .B2(n687), .ZN(
        u1_fracta_s[40]) );
  OAI22_X2 U483 ( .A1(n4854), .A2(n688), .B1(n4862), .B2(n689), .ZN(
        u1_fracta_s[3]) );
  OAI22_X2 U484 ( .A1(n4854), .A2(n690), .B1(n4862), .B2(n691), .ZN(
        u1_fracta_s[39]) );
  OAI22_X2 U485 ( .A1(n4854), .A2(n692), .B1(n4862), .B2(n693), .ZN(
        u1_fracta_s[38]) );
  OAI22_X2 U486 ( .A1(n4854), .A2(n694), .B1(n4862), .B2(n695), .ZN(
        u1_fracta_s[37]) );
  OAI22_X2 U487 ( .A1(n4854), .A2(n696), .B1(n4862), .B2(n697), .ZN(
        u1_fracta_s[36]) );
  OAI22_X2 U488 ( .A1(n4854), .A2(n698), .B1(n4862), .B2(n699), .ZN(
        u1_fracta_s[35]) );
  OAI22_X2 U489 ( .A1(n4854), .A2(n700), .B1(n4863), .B2(n701), .ZN(
        u1_fracta_s[34]) );
  OAI22_X2 U490 ( .A1(n4854), .A2(n702), .B1(n4863), .B2(n703), .ZN(
        u1_fracta_s[33]) );
  OAI22_X2 U491 ( .A1(n4854), .A2(n704), .B1(n4863), .B2(n705), .ZN(
        u1_fracta_s[32]) );
  OAI22_X2 U492 ( .A1(n4854), .A2(n706), .B1(n4863), .B2(n707), .ZN(
        u1_fracta_s[31]) );
  OAI22_X2 U493 ( .A1(n4853), .A2(n708), .B1(n4863), .B2(n709), .ZN(
        u1_fracta_s[30]) );
  OAI22_X2 U494 ( .A1(n4858), .A2(n710), .B1(n4856), .B2(n711), .ZN(
        u1_fracta_s[2]) );
  OAI22_X2 U495 ( .A1(n4853), .A2(n712), .B1(n4863), .B2(n713), .ZN(
        u1_fracta_s[29]) );
  OAI22_X2 U496 ( .A1(n4853), .A2(n714), .B1(n4863), .B2(n715), .ZN(
        u1_fracta_s[28]) );
  OAI22_X2 U497 ( .A1(n4853), .A2(n716), .B1(n4863), .B2(n717), .ZN(
        u1_fracta_s[27]) );
  OAI22_X2 U498 ( .A1(n4853), .A2(n718), .B1(n4863), .B2(n719), .ZN(
        u1_fracta_s[26]) );
  OAI22_X2 U499 ( .A1(n4853), .A2(n720), .B1(n4863), .B2(n721), .ZN(
        u1_fracta_s[25]) );
  OAI22_X2 U500 ( .A1(n4853), .A2(n722), .B1(n4863), .B2(n723), .ZN(
        u1_fracta_s[24]) );
  OAI22_X2 U501 ( .A1(n4853), .A2(n724), .B1(n4863), .B2(n725), .ZN(
        u1_fracta_s[23]) );
  OAI22_X2 U502 ( .A1(n4853), .A2(n726), .B1(n4863), .B2(n727), .ZN(
        u1_fracta_s[22]) );
  OAI22_X2 U503 ( .A1(n4853), .A2(n728), .B1(n4863), .B2(n729), .ZN(
        u1_fracta_s[21]) );
  OAI22_X2 U504 ( .A1(n4853), .A2(n730), .B1(n4863), .B2(n731), .ZN(
        u1_fracta_s[20]) );
  OAI22_X2 U505 ( .A1(n4858), .A2(n732), .B1(n4857), .B2(n733), .ZN(
        u1_fracta_s[1]) );
  OAI22_X2 U506 ( .A1(n4856), .A2(n734), .B1(n4863), .B2(n735), .ZN(
        u1_fracta_s[19]) );
  OAI22_X2 U507 ( .A1(n4853), .A2(n736), .B1(n4863), .B2(n737), .ZN(
        u1_fracta_s[18]) );
  OAI22_X2 U508 ( .A1(n4857), .A2(n738), .B1(n4863), .B2(n739), .ZN(
        u1_fracta_s[17]) );
  OAI22_X2 U509 ( .A1(n4857), .A2(n740), .B1(n4863), .B2(n741), .ZN(
        u1_fracta_s[16]) );
  OAI22_X2 U510 ( .A1(n4853), .A2(n742), .B1(n4863), .B2(n743), .ZN(
        u1_fracta_s[15]) );
  OAI22_X2 U511 ( .A1(n4856), .A2(n744), .B1(n4868), .B2(n745), .ZN(
        u1_fracta_s[14]) );
  OAI22_X2 U512 ( .A1(n4857), .A2(n746), .B1(n4868), .B2(n747), .ZN(
        u1_fracta_s[13]) );
  OAI22_X2 U513 ( .A1(n4853), .A2(n748), .B1(n4868), .B2(n749), .ZN(
        u1_fracta_s[12]) );
  OAI22_X2 U514 ( .A1(n4853), .A2(n750), .B1(n4868), .B2(n751), .ZN(
        u1_fracta_s[11]) );
  OAI22_X2 U515 ( .A1(n4856), .A2(n752), .B1(n4863), .B2(n753), .ZN(
        u1_fracta_s[10]) );
  OAI22_X2 U516 ( .A1(n4860), .A2(n754), .B1(n4854), .B2(n755), .ZN(
        u1_fracta_s[0]) );
  OAI22_X2 U518 ( .A1(n4841), .A2(n4569), .B1(n4832), .B2(n4582), .ZN(
        u1_exp_small[7]) );
  OAI22_X2 U519 ( .A1(n4840), .A2(n4471), .B1(n4833), .B2(n4575), .ZN(
        u1_exp_small[6]) );
  OAI22_X2 U520 ( .A1(n4841), .A2(n4398), .B1(n4834), .B2(n4586), .ZN(
        u1_exp_small[5]) );
  OAI22_X2 U521 ( .A1(n4841), .A2(n4486), .B1(n4834), .B2(n4589), .ZN(
        u1_exp_small[4]) );
  OAI22_X2 U522 ( .A1(n4841), .A2(n4591), .B1(n4833), .B2(n4485), .ZN(
        u1_exp_small[3]) );
  OAI22_X2 U523 ( .A1(n4841), .A2(n4590), .B1(n4833), .B2(n4583), .ZN(
        u1_exp_small[2]) );
  OAI22_X2 U524 ( .A1(n4841), .A2(n4360), .B1(n4833), .B2(n4584), .ZN(
        u1_exp_small[1]) );
  OAI22_X2 U525 ( .A1(n4487), .A2(n4843), .B1(n4833), .B2(n4592), .ZN(
        u1_exp_small[10]) );
  OAI22_X2 U526 ( .A1(n4841), .A2(n4371), .B1(n4833), .B2(n4585), .ZN(
        u1_exp_small[0]) );
  AND2_X2 U527 ( .A1(u1_exp_diff2[9]), .A2(n773), .ZN(u1_exp_diff_9_) );
  AND2_X2 U528 ( .A1(u1_exp_diff2[8]), .A2(n773), .ZN(u1_exp_diff_8_) );
  AND2_X2 U529 ( .A1(u1_exp_diff2[7]), .A2(n773), .ZN(u1_exp_diff_7_) );
  AND2_X2 U530 ( .A1(u1_exp_diff2[6]), .A2(n773), .ZN(u1_exp_diff_6_) );
  AND2_X2 U531 ( .A1(u1_exp_diff2[10]), .A2(n773), .ZN(u1_exp_diff_10_) );
  OAI211_X2 U568 ( .C1(u1_signa_r), .C2(n799), .A(rmode_r2[0]), .B(rmode_r2[1]), .ZN(n801) );
  XOR2_X2 U569 ( .A(n4624), .B(u1_add_r), .Z(n799) );
  OAI221_X2 U571 ( .B1(n802), .B2(n803), .C1(n804), .C2(n805), .A(n806), .ZN(
        u1_N296) );
  OAI221_X2 U573 ( .B1(n809), .B2(n810), .C1(n811), .C2(n812), .A(n813), .ZN(
        n808) );
  OAI221_X2 U575 ( .B1(n817), .B2(n818), .C1(n819), .C2(n820), .A(n821), .ZN(
        n807) );
  AND4_X2 U577 ( .A1(n828), .A2(n829), .A3(n830), .A4(n831), .ZN(n804) );
  OAI22_X2 U581 ( .A1(n839), .A2(n840), .B1(n841), .B2(n842), .ZN(n834) );
  AOI221_X2 U584 ( .B1(n6287), .B2(n855), .C1(n6298), .C2(n856), .A(n857), 
        .ZN(n828) );
  NOR4_X2 U585 ( .A1(n858), .A2(n859), .A3(n860), .A4(n6286), .ZN(n802) );
  AOI221_X2 U587 ( .B1(n4180), .B2(n852), .C1(n4158), .C2(n6297), .A(n816), 
        .ZN(n862) );
  OAI211_X2 U588 ( .C1(n863), .C2(n864), .A(n865), .B(n866), .ZN(n816) );
  AOI221_X2 U589 ( .B1(n6344), .B2(n6294), .C1(n6347), .C2(n868), .A(n857), 
        .ZN(n866) );
  OAI22_X2 U590 ( .A1(n6295), .A2(n870), .B1(n871), .B2(n872), .ZN(n857) );
  AOI22_X2 U592 ( .A1(n6297), .A2(n873), .B1(n852), .B2(n874), .ZN(n865) );
  OAI221_X2 U593 ( .B1(n875), .B2(n876), .C1(n872), .C2(n877), .A(n878), .ZN(
        n860) );
  AOI22_X2 U594 ( .A1(n868), .A2(n6308), .B1(n6296), .B2(n6335), .ZN(n878) );
  OAI221_X2 U596 ( .B1(n880), .B2(n818), .C1(n881), .C2(n820), .A(n882), .ZN(
        n859) );
  AOI22_X2 U597 ( .A1(n6299), .A2(n883), .B1(n6287), .B2(n884), .ZN(n882) );
  OAI221_X2 U598 ( .B1(n885), .B2(n840), .C1(n886), .C2(n887), .A(n888), .ZN(
        n858) );
  AOI22_X2 U599 ( .A1(u1_exp_diff_sft_0_), .A2(n889), .B1(n6288), .B2(n890), 
        .ZN(n888) );
  NAND4_X2 U600 ( .A1(n891), .A2(n892), .A3(n893), .A4(n894), .ZN(n889) );
  AOI221_X2 U601 ( .B1(n6288), .B2(n895), .C1(n6291), .C2(n896), .A(n897), 
        .ZN(n894) );
  OAI22_X2 U602 ( .A1(n836), .A2(n898), .B1(n899), .B2(n840), .ZN(n897) );
  OR2_X2 U604 ( .A1(n833), .A2(n4159), .ZN(n873) );
  OR2_X2 U605 ( .A1(n895), .A2(n4160), .ZN(n833) );
  OR2_X2 U606 ( .A1(n890), .A2(n4161), .ZN(n895) );
  OR2_X2 U607 ( .A1(n825), .A2(n6322), .ZN(n890) );
  NAND2_X2 U608 ( .A1(n841), .A2(n900), .ZN(n825) );
  AND2_X2 U609 ( .A1(n899), .A2(n901), .ZN(n841) );
  AND2_X2 U610 ( .A1(n885), .A2(n902), .ZN(n899) );
  NAND2_X2 U615 ( .A1(n908), .A2(n903), .ZN(n820) );
  NAND2_X2 U622 ( .A1(n839), .A2(n916), .ZN(n827) );
  NAND2_X2 U624 ( .A1(n886), .A2(n917), .ZN(n896) );
  OR2_X2 U626 ( .A1(n845), .A2(n6304), .ZN(n823) );
  AOI22_X2 U628 ( .A1(n4846), .A2(u6_N37), .B1(n4839), .B2(fracta_mul[37]), 
        .ZN(n918) );
  OR2_X2 U629 ( .A1(n906), .A2(u1_adj_op_36_), .ZN(n845) );
  OAI22_X2 U630 ( .A1(n4841), .A2(n4604), .B1(n4833), .B2(n4365), .ZN(
        u1_adj_op_36_) );
  NAND2_X2 U632 ( .A1(n880), .A2(n774), .ZN(n906) );
  AOI22_X2 U633 ( .A1(n4829), .A2(u6_N35), .B1(n4839), .B2(fracta_mul[35]), 
        .ZN(n774) );
  AND2_X2 U634 ( .A1(n817), .A2(n921), .ZN(n880) );
  OR2_X2 U636 ( .A1(n907), .A2(n4173), .ZN(n847) );
  NAND2_X2 U637 ( .A1(n881), .A2(n775), .ZN(n907) );
  AOI22_X2 U638 ( .A1(n4846), .A2(u6_N31), .B1(n4839), .B2(fracta_mul[31]), 
        .ZN(n775) );
  AND2_X2 U639 ( .A1(n819), .A2(n776), .ZN(n881) );
  AOI22_X2 U640 ( .A1(n4829), .A2(u6_N30), .B1(n4839), .B2(fracta_mul[30]), 
        .ZN(n776) );
  OAI22_X2 U642 ( .A1(n4841), .A2(n4599), .B1(n4833), .B2(n4373), .ZN(
        u1_adj_op_29_) );
  OR2_X2 U644 ( .A1(n905), .A2(n4174), .ZN(n844) );
  OR2_X2 U645 ( .A1(n883), .A2(n4175), .ZN(n905) );
  NAND2_X2 U646 ( .A1(n809), .A2(n924), .ZN(n883) );
  OR2_X2 U648 ( .A1(n910), .A2(n6332), .ZN(n851) );
  OR3_X2 U649 ( .A1(n4180), .A2(n4179), .A3(n874), .ZN(n910) );
  OR2_X2 U650 ( .A1(n853), .A2(n4181), .ZN(n874) );
  OR2_X2 U651 ( .A1(n911), .A2(n6333), .ZN(n853) );
  OR2_X2 U654 ( .A1(n909), .A2(n4186), .ZN(n849) );
  OR2_X2 U655 ( .A1(n884), .A2(n6336), .ZN(n909) );
  NAND2_X2 U656 ( .A1(n811), .A2(n927), .ZN(n884) );
  OR2_X2 U658 ( .A1(n914), .A2(n4190), .ZN(n855) );
  NAND2_X2 U659 ( .A1(n875), .A2(n928), .ZN(n914) );
  OR2_X2 U661 ( .A1(n856), .A2(n4193), .ZN(n815) );
  OR2_X2 U662 ( .A1(n915), .A2(n6341), .ZN(n856) );
  NAND4_X2 U663 ( .A1(n871), .A2(n877), .A3(n929), .A4(n930), .ZN(n915) );
  NAND4_X2 U665 ( .A1(n931), .A2(n870), .A3(n932), .A4(n879), .ZN(n913) );
  AOI22_X2 U666 ( .A1(n4829), .A2(u6_N2), .B1(n4839), .B2(fracta_mul[2]), .ZN(
        n879) );
  NAND4_X2 U667 ( .A1(n6284), .A2(n934), .A3(n935), .A4(n936), .ZN(u1_N295) );
  NAND2_X2 U670 ( .A1(n937), .A2(n6303), .ZN(n810) );
  NAND2_X2 U672 ( .A1(n908), .A2(n6301), .ZN(n887) );
  NAND4_X2 U675 ( .A1(n6293), .A2(n6302), .A3(n938), .A4(n903), .ZN(n818) );
  NAND4_X2 U678 ( .A1(n6293), .A2(n6301), .A3(n6302), .A4(n938), .ZN(n840) );
  NAND2_X2 U680 ( .A1(n937), .A2(n938), .ZN(n876) );
  NAND2_X2 U683 ( .A1(n940), .A2(n6302), .ZN(n898) );
  NAND2_X2 U686 ( .A1(n940), .A2(n912), .ZN(n864) );
  AND3_X2 U688 ( .A1(n6301), .A2(n912), .A3(n904), .ZN(n852) );
  NOR4_X2 U689 ( .A1(n939), .A2(n6303), .A3(n6302), .A4(n6301), .ZN(n868) );
  OAI221_X2 U691 ( .B1(n6293), .B2(n6301), .C1(n805), .C2(n838), .A(n872), 
        .ZN(n941) );
  NAND4_X2 U692 ( .A1(n939), .A2(n6301), .A3(n938), .A4(n912), .ZN(n872) );
  OR2_X2 U695 ( .A1(n6285), .A2(u1_exp_diff_sft_0_), .ZN(n805) );
  AND2_X2 U696 ( .A1(u1_exp_diff_0_), .A2(n6300), .ZN(u1_exp_diff_sft_0_) );
  AND2_X2 U697 ( .A1(u1_exp_diff2[0]), .A2(n773), .ZN(u1_exp_diff_0_) );
  NAND2_X2 U699 ( .A1(u1_exp_diff_1_), .A2(n6300), .ZN(n803) );
  AND2_X2 U700 ( .A1(u1_exp_diff2[1]), .A2(n773), .ZN(u1_exp_diff_1_) );
  NAND2_X2 U701 ( .A1(n943), .A2(n944), .ZN(u0_N7) );
  AND2_X2 U703 ( .A1(n4594), .A2(n946), .ZN(u0_N5) );
  AND2_X2 U705 ( .A1(u0_fractb_00), .A2(u0_expb_00), .ZN(u0_N17) );
  AND2_X2 U706 ( .A1(u0_fracta_00), .A2(u0_expa_00), .ZN(u0_N16) );
  XOR2_X2 U709 ( .A(n4620), .B(u2_sign_d), .Z(n3953) );
  XOR2_X2 U710 ( .A(opa_r[63]), .B(opb_r[63]), .Z(u2_sign_d) );
  OAI22_X2 U712 ( .A1(u1_adj_op_out_sft_55_), .A2(n4842), .B1(n4833), .B2(
        u6_N52), .ZN(n655) );
  OAI22_X2 U714 ( .A1(n4832), .A2(u1_adj_op_out_sft_55_), .B1(n4825), .B2(
        n4842), .ZN(n654) );
  OAI22_X2 U716 ( .A1(u1_adj_op_out_sft_54_), .A2(n4843), .B1(n4833), .B2(
        u6_N51), .ZN(n657) );
  OAI22_X2 U718 ( .A1(n4832), .A2(u1_adj_op_out_sft_54_), .B1(fracta_mul[51]), 
        .B2(n4842), .ZN(n656) );
  OAI22_X2 U720 ( .A1(u1_adj_op_out_sft_53_), .A2(n4843), .B1(n4833), .B2(
        u6_N50), .ZN(n659) );
  OAI22_X2 U722 ( .A1(n4831), .A2(u1_adj_op_out_sft_53_), .B1(fracta_mul[50]), 
        .B2(n4842), .ZN(n658) );
  OAI22_X2 U724 ( .A1(u1_adj_op_out_sft_52_), .A2(n4843), .B1(n4833), .B2(
        u6_N49), .ZN(n661) );
  OAI22_X2 U726 ( .A1(n4829), .A2(u1_adj_op_out_sft_52_), .B1(fracta_mul[49]), 
        .B2(n4842), .ZN(n660) );
  OAI22_X2 U728 ( .A1(u1_adj_op_out_sft_51_), .A2(n4843), .B1(n4833), .B2(
        u6_N48), .ZN(n663) );
  OAI22_X2 U730 ( .A1(n4846), .A2(u1_adj_op_out_sft_51_), .B1(fracta_mul[48]), 
        .B2(n4842), .ZN(n662) );
  OAI22_X2 U732 ( .A1(u1_adj_op_out_sft_50_), .A2(n4843), .B1(n4829), .B2(
        u6_N47), .ZN(n665) );
  OAI22_X2 U734 ( .A1(n4832), .A2(u1_adj_op_out_sft_50_), .B1(fracta_mul[47]), 
        .B2(n4842), .ZN(n664) );
  OAI22_X2 U736 ( .A1(u1_adj_op_out_sft_49_), .A2(n4843), .B1(n4833), .B2(
        u6_N46), .ZN(n669) );
  OAI22_X2 U738 ( .A1(n4832), .A2(u1_adj_op_out_sft_49_), .B1(fracta_mul[46]), 
        .B2(n4842), .ZN(n668) );
  OAI22_X2 U740 ( .A1(u1_adj_op_out_sft_48_), .A2(n4843), .B1(n4833), .B2(
        u6_N45), .ZN(n671) );
  OAI22_X2 U742 ( .A1(n4829), .A2(u1_adj_op_out_sft_48_), .B1(fracta_mul[45]), 
        .B2(n4842), .ZN(n670) );
  OAI22_X2 U744 ( .A1(u1_adj_op_out_sft_47_), .A2(n4843), .B1(n4829), .B2(
        u6_N44), .ZN(n673) );
  OAI22_X2 U746 ( .A1(n4832), .A2(u1_adj_op_out_sft_47_), .B1(fracta_mul[44]), 
        .B2(n4842), .ZN(n672) );
  OAI22_X2 U748 ( .A1(u1_adj_op_out_sft_46_), .A2(n4843), .B1(n4846), .B2(
        u6_N43), .ZN(n675) );
  OAI22_X2 U750 ( .A1(n4829), .A2(u1_adj_op_out_sft_46_), .B1(fracta_mul[43]), 
        .B2(n4842), .ZN(n674) );
  OAI22_X2 U752 ( .A1(u1_adj_op_out_sft_45_), .A2(n4843), .B1(n4829), .B2(
        u6_N42), .ZN(n677) );
  OAI22_X2 U754 ( .A1(n4829), .A2(u1_adj_op_out_sft_45_), .B1(fracta_mul[42]), 
        .B2(n4842), .ZN(n676) );
  OAI22_X2 U756 ( .A1(u1_adj_op_out_sft_44_), .A2(n4843), .B1(n4829), .B2(
        u6_N41), .ZN(n679) );
  OAI22_X2 U758 ( .A1(n4829), .A2(u1_adj_op_out_sft_44_), .B1(fracta_mul[41]), 
        .B2(n4842), .ZN(n678) );
  OAI22_X2 U760 ( .A1(u1_adj_op_out_sft_43_), .A2(n4843), .B1(n4829), .B2(
        u6_N40), .ZN(n681) );
  OAI22_X2 U762 ( .A1(n4846), .A2(u1_adj_op_out_sft_43_), .B1(fracta_mul[40]), 
        .B2(n4842), .ZN(n680) );
  OAI22_X2 U764 ( .A1(u1_adj_op_out_sft_42_), .A2(n4843), .B1(n4829), .B2(
        u6_N39), .ZN(n683) );
  OAI22_X2 U766 ( .A1(n4829), .A2(u1_adj_op_out_sft_42_), .B1(fracta_mul[39]), 
        .B2(n4842), .ZN(n682) );
  OAI22_X2 U768 ( .A1(u1_adj_op_out_sft_41_), .A2(n4843), .B1(n4846), .B2(
        u6_N38), .ZN(n685) );
  OAI22_X2 U770 ( .A1(n4829), .A2(u1_adj_op_out_sft_41_), .B1(fracta_mul[38]), 
        .B2(n4842), .ZN(n684) );
  OAI22_X2 U772 ( .A1(u1_adj_op_out_sft_40_), .A2(n4843), .B1(n4829), .B2(
        u6_N37), .ZN(n687) );
  OAI22_X2 U774 ( .A1(n4829), .A2(u1_adj_op_out_sft_40_), .B1(fracta_mul[37]), 
        .B2(n4842), .ZN(n686) );
  OAI22_X2 U776 ( .A1(u1_adj_op_out_sft_39_), .A2(n4843), .B1(n4829), .B2(
        u6_N36), .ZN(n691) );
  OAI22_X2 U778 ( .A1(n4829), .A2(u1_adj_op_out_sft_39_), .B1(fracta_mul[36]), 
        .B2(n4842), .ZN(n690) );
  OAI22_X2 U780 ( .A1(u1_adj_op_out_sft_38_), .A2(n4843), .B1(n4829), .B2(
        u6_N35), .ZN(n693) );
  OAI22_X2 U782 ( .A1(n4846), .A2(u1_adj_op_out_sft_38_), .B1(fracta_mul[35]), 
        .B2(n4842), .ZN(n692) );
  OAI22_X2 U784 ( .A1(u1_adj_op_out_sft_37_), .A2(n4843), .B1(n4829), .B2(
        u6_N34), .ZN(n695) );
  OAI22_X2 U786 ( .A1(n4829), .A2(u1_adj_op_out_sft_37_), .B1(fracta_mul[34]), 
        .B2(n4842), .ZN(n694) );
  OAI22_X2 U788 ( .A1(u1_adj_op_out_sft_36_), .A2(n4842), .B1(n4846), .B2(
        u6_N33), .ZN(n697) );
  OAI22_X2 U790 ( .A1(n4829), .A2(u1_adj_op_out_sft_36_), .B1(fracta_mul[33]), 
        .B2(n4842), .ZN(n696) );
  OAI22_X2 U792 ( .A1(u1_adj_op_out_sft_35_), .A2(n4843), .B1(n4829), .B2(
        u6_N32), .ZN(n699) );
  OAI22_X2 U794 ( .A1(n4829), .A2(u1_adj_op_out_sft_35_), .B1(fracta_mul[32]), 
        .B2(n4842), .ZN(n698) );
  OAI22_X2 U796 ( .A1(u1_adj_op_out_sft_34_), .A2(n4843), .B1(n4829), .B2(
        u6_N31), .ZN(n701) );
  OAI22_X2 U798 ( .A1(n4831), .A2(u1_adj_op_out_sft_34_), .B1(fracta_mul[31]), 
        .B2(n4842), .ZN(n700) );
  OAI22_X2 U800 ( .A1(u1_adj_op_out_sft_33_), .A2(n4843), .B1(n4829), .B2(
        u6_N30), .ZN(n703) );
  OAI22_X2 U802 ( .A1(n4831), .A2(u1_adj_op_out_sft_33_), .B1(fracta_mul[30]), 
        .B2(n4842), .ZN(n702) );
  OAI22_X2 U804 ( .A1(u1_adj_op_out_sft_32_), .A2(n4843), .B1(n4846), .B2(
        u6_N29), .ZN(n705) );
  OAI22_X2 U806 ( .A1(n4831), .A2(u1_adj_op_out_sft_32_), .B1(fracta_mul[29]), 
        .B2(n4842), .ZN(n704) );
  OAI22_X2 U808 ( .A1(u1_adj_op_out_sft_31_), .A2(n4843), .B1(n4829), .B2(
        u6_N28), .ZN(n707) );
  OAI22_X2 U810 ( .A1(n4831), .A2(u1_adj_op_out_sft_31_), .B1(fracta_mul[28]), 
        .B2(n4842), .ZN(n706) );
  OAI22_X2 U812 ( .A1(u1_adj_op_out_sft_30_), .A2(n4843), .B1(n4829), .B2(
        u6_N27), .ZN(n709) );
  OAI22_X2 U814 ( .A1(n4831), .A2(u1_adj_op_out_sft_30_), .B1(fracta_mul[27]), 
        .B2(n4842), .ZN(n708) );
  OAI22_X2 U816 ( .A1(u1_adj_op_out_sft_29_), .A2(n4843), .B1(n4829), .B2(
        u6_N26), .ZN(n713) );
  OAI22_X2 U818 ( .A1(n4831), .A2(u1_adj_op_out_sft_29_), .B1(fracta_mul[26]), 
        .B2(n4842), .ZN(n712) );
  OAI22_X2 U820 ( .A1(u1_adj_op_out_sft_28_), .A2(n4843), .B1(n4829), .B2(
        u6_N25), .ZN(n715) );
  OAI22_X2 U822 ( .A1(n4831), .A2(u1_adj_op_out_sft_28_), .B1(fracta_mul[25]), 
        .B2(n4842), .ZN(n714) );
  OAI22_X2 U824 ( .A1(u1_adj_op_out_sft_27_), .A2(n4843), .B1(n4846), .B2(
        u6_N24), .ZN(n717) );
  OAI22_X2 U826 ( .A1(n4831), .A2(u1_adj_op_out_sft_27_), .B1(fracta_mul[24]), 
        .B2(n4842), .ZN(n716) );
  OAI22_X2 U828 ( .A1(u1_adj_op_out_sft_26_), .A2(n4842), .B1(n4829), .B2(
        u6_N23), .ZN(n719) );
  OAI22_X2 U830 ( .A1(n4831), .A2(u1_adj_op_out_sft_26_), .B1(fracta_mul[23]), 
        .B2(n4842), .ZN(n718) );
  OAI22_X2 U832 ( .A1(u1_adj_op_out_sft_25_), .A2(n4842), .B1(n4829), .B2(
        u6_N22), .ZN(n721) );
  OAI22_X2 U834 ( .A1(n4831), .A2(u1_adj_op_out_sft_25_), .B1(fracta_mul[22]), 
        .B2(n4842), .ZN(n720) );
  OAI22_X2 U836 ( .A1(u1_adj_op_out_sft_24_), .A2(n4842), .B1(n4829), .B2(
        u6_N21), .ZN(n723) );
  OAI22_X2 U838 ( .A1(n4831), .A2(u1_adj_op_out_sft_24_), .B1(fracta_mul[21]), 
        .B2(n4842), .ZN(n722) );
  OAI22_X2 U840 ( .A1(u1_adj_op_out_sft_23_), .A2(n4842), .B1(n4829), .B2(
        u6_N20), .ZN(n725) );
  OAI22_X2 U842 ( .A1(n4831), .A2(u1_adj_op_out_sft_23_), .B1(fracta_mul[20]), 
        .B2(n4843), .ZN(n724) );
  OAI22_X2 U844 ( .A1(u1_adj_op_out_sft_22_), .A2(n4843), .B1(n4846), .B2(
        u6_N19), .ZN(n727) );
  OAI22_X2 U846 ( .A1(n4830), .A2(u1_adj_op_out_sft_22_), .B1(fracta_mul[19]), 
        .B2(n4842), .ZN(n726) );
  OAI22_X2 U848 ( .A1(u1_adj_op_out_sft_21_), .A2(n4843), .B1(n4829), .B2(
        u6_N18), .ZN(n729) );
  OAI22_X2 U850 ( .A1(n4830), .A2(u1_adj_op_out_sft_21_), .B1(fracta_mul[18]), 
        .B2(n4842), .ZN(n728) );
  OAI22_X2 U852 ( .A1(u1_adj_op_out_sft_20_), .A2(n4843), .B1(n4829), .B2(
        u6_N17), .ZN(n731) );
  OAI22_X2 U854 ( .A1(n4830), .A2(u1_adj_op_out_sft_20_), .B1(fracta_mul[17]), 
        .B2(n4842), .ZN(n730) );
  OAI22_X2 U856 ( .A1(u1_adj_op_out_sft_19_), .A2(n4843), .B1(n4829), .B2(
        u6_N16), .ZN(n735) );
  OAI22_X2 U858 ( .A1(n4830), .A2(u1_adj_op_out_sft_19_), .B1(fracta_mul[16]), 
        .B2(n4842), .ZN(n734) );
  OAI22_X2 U860 ( .A1(u1_adj_op_out_sft_18_), .A2(n4842), .B1(n4829), .B2(
        u6_N15), .ZN(n737) );
  OAI22_X2 U862 ( .A1(n4830), .A2(u1_adj_op_out_sft_18_), .B1(fracta_mul[15]), 
        .B2(n4842), .ZN(n736) );
  OAI22_X2 U864 ( .A1(u1_adj_op_out_sft_17_), .A2(n4842), .B1(n4846), .B2(
        u6_N14), .ZN(n739) );
  OAI22_X2 U866 ( .A1(n4830), .A2(u1_adj_op_out_sft_17_), .B1(fracta_mul[14]), 
        .B2(n4842), .ZN(n738) );
  OAI22_X2 U868 ( .A1(u1_adj_op_out_sft_16_), .A2(n4843), .B1(n4829), .B2(
        u6_N13), .ZN(n741) );
  OAI22_X2 U870 ( .A1(n4829), .A2(u1_adj_op_out_sft_16_), .B1(fracta_mul[13]), 
        .B2(n4842), .ZN(n740) );
  OAI22_X2 U872 ( .A1(u1_adj_op_out_sft_15_), .A2(n4842), .B1(n4829), .B2(
        u6_N12), .ZN(n743) );
  OAI22_X2 U874 ( .A1(n4829), .A2(u1_adj_op_out_sft_15_), .B1(fracta_mul[12]), 
        .B2(n4842), .ZN(n742) );
  OAI22_X2 U876 ( .A1(u1_adj_op_out_sft_14_), .A2(n4842), .B1(n4829), .B2(
        u6_N11), .ZN(n745) );
  OAI22_X2 U878 ( .A1(n4829), .A2(u1_adj_op_out_sft_14_), .B1(fracta_mul[11]), 
        .B2(n4839), .ZN(n744) );
  OAI22_X2 U880 ( .A1(u1_adj_op_out_sft_13_), .A2(n4842), .B1(n4829), .B2(
        u6_N10), .ZN(n747) );
  OAI22_X2 U882 ( .A1(n4829), .A2(u1_adj_op_out_sft_13_), .B1(fracta_mul[10]), 
        .B2(n4839), .ZN(n746) );
  OAI22_X2 U884 ( .A1(u1_adj_op_out_sft_12_), .A2(n4842), .B1(n4846), .B2(
        u6_N9), .ZN(n749) );
  OAI22_X2 U886 ( .A1(n4830), .A2(u1_adj_op_out_sft_12_), .B1(fracta_mul[9]), 
        .B2(n4839), .ZN(n748) );
  OAI22_X2 U888 ( .A1(u1_adj_op_out_sft_11_), .A2(n4843), .B1(n4829), .B2(
        u6_N8), .ZN(n751) );
  OAI22_X2 U890 ( .A1(n4829), .A2(u1_adj_op_out_sft_11_), .B1(fracta_mul[8]), 
        .B2(n4839), .ZN(n750) );
  OAI22_X2 U892 ( .A1(u1_adj_op_out_sft_10_), .A2(n4843), .B1(n4829), .B2(
        u6_N7), .ZN(n753) );
  OAI22_X2 U894 ( .A1(n4829), .A2(u1_adj_op_out_sft_10_), .B1(fracta_mul[7]), 
        .B2(n4839), .ZN(n752) );
  OAI22_X2 U896 ( .A1(u1_adj_op_out_sft_9_), .A2(n4843), .B1(n4829), .B2(u6_N6), .ZN(n645) );
  OAI22_X2 U898 ( .A1(n4829), .A2(u1_adj_op_out_sft_9_), .B1(fracta_mul[6]), 
        .B2(n4843), .ZN(n644) );
  OAI22_X2 U900 ( .A1(u1_adj_op_out_sft_8_), .A2(n4843), .B1(n4829), .B2(u6_N5), .ZN(n647) );
  OAI22_X2 U902 ( .A1(n4829), .A2(u1_adj_op_out_sft_8_), .B1(fracta_mul[5]), 
        .B2(n4839), .ZN(n646) );
  OAI22_X2 U904 ( .A1(u1_adj_op_out_sft_7_), .A2(n4843), .B1(n4846), .B2(u6_N4), .ZN(n649) );
  OAI22_X2 U906 ( .A1(n4829), .A2(u1_adj_op_out_sft_7_), .B1(fracta_mul[4]), 
        .B2(n4839), .ZN(n648) );
  OAI22_X2 U908 ( .A1(u1_adj_op_out_sft_6_), .A2(n4843), .B1(n4829), .B2(u6_N3), .ZN(n651) );
  OAI22_X2 U910 ( .A1(n4829), .A2(u1_adj_op_out_sft_6_), .B1(fracta_mul[3]), 
        .B2(n4843), .ZN(n650) );
  OAI22_X2 U912 ( .A1(u1_adj_op_out_sft_5_), .A2(n4843), .B1(n4829), .B2(u6_N2), .ZN(n653) );
  OAI22_X2 U914 ( .A1(n4829), .A2(u1_adj_op_out_sft_5_), .B1(fracta_mul[2]), 
        .B2(n4839), .ZN(n652) );
  OAI22_X2 U916 ( .A1(u1_adj_op_out_sft_4_), .A2(n4843), .B1(n4829), .B2(u6_N1), .ZN(n667) );
  OAI22_X2 U918 ( .A1(n4831), .A2(u1_adj_op_out_sft_4_), .B1(fracta_mul[1]), 
        .B2(n4839), .ZN(n666) );
  OAI22_X2 U920 ( .A1(u1_adj_op_out_sft_3_), .A2(n4843), .B1(n4832), .B2(u6_N0), .ZN(n689) );
  OAI22_X2 U922 ( .A1(n4830), .A2(u1_adj_op_out_sft_3_), .B1(fracta_mul[0]), 
        .B2(n4843), .ZN(n688) );
  NAND2_X2 U924 ( .A1(u1_adj_op_out_sft_2_), .A2(n4834), .ZN(n710) );
  NAND2_X2 U926 ( .A1(u1_adj_op_out_sft_2_), .A2(n4844), .ZN(n711) );
  NAND2_X2 U928 ( .A1(u1_adj_op_out_sft_1_), .A2(n4834), .ZN(n732) );
  NAND2_X2 U930 ( .A1(u1_adj_op_out_sft_1_), .A2(n4844), .ZN(n733) );
  AND2_X2 U937 ( .A1(u1_exp_diff2[3]), .A2(n773), .ZN(u1_exp_diff_3_) );
  AND2_X2 U940 ( .A1(u1_exp_diff2[5]), .A2(n773), .ZN(u1_exp_diff_5_) );
  AND2_X2 U943 ( .A1(u1_exp_diff2[4]), .A2(n773), .ZN(u1_exp_diff_4_) );
  NAND2_X2 U945 ( .A1(u1_exp_diff_2_), .A2(n6300), .ZN(n939) );
  AND2_X2 U947 ( .A1(u1_exp_diff2[2]), .A2(n773), .ZN(u1_exp_diff_2_) );
  OAI22_X2 U949 ( .A1(n4830), .A2(n4487), .B1(n4592), .B2(n4843), .ZN(n4070)
         );
  NAND4_X2 U953 ( .A1(opa_r[60]), .A2(opa_r[61]), .A3(n950), .A4(n951), .ZN(
        n949) );
  NOR4_X2 U954 ( .A1(n952), .A2(n4485), .A3(n4586), .A4(n4589), .ZN(n951) );
  OAI22_X2 U957 ( .A1(n4824), .A2(n4611), .B1(n4825), .B2(n5951), .ZN(u6_N99)
         );
  AOI22_X2 U960 ( .A1(n4825), .A2(fracta_mul[43]), .B1(n4826), .B2(N304), .ZN(
        n955) );
  OAI22_X2 U961 ( .A1(n4824), .A2(n4375), .B1(n4825), .B2(n5952), .ZN(u6_N97)
         );
  OAI22_X2 U963 ( .A1(n4824), .A2(n4617), .B1(n4825), .B2(n5953), .ZN(u6_N96)
         );
  AOI22_X2 U966 ( .A1(n4825), .A2(fracta_mul[40]), .B1(n4826), .B2(N301), .ZN(
        n960) );
  OAI22_X2 U967 ( .A1(n4824), .A2(n4618), .B1(n4825), .B2(n5954), .ZN(u6_N94)
         );
  OAI22_X2 U969 ( .A1(n4824), .A2(n4374), .B1(n4825), .B2(n5955), .ZN(u6_N93)
         );
  AOI22_X2 U972 ( .A1(n4825), .A2(fracta_mul[37]), .B1(n4826), .B2(N298), .ZN(
        n965) );
  OAI22_X2 U973 ( .A1(n4824), .A2(n4365), .B1(n4825), .B2(n5956), .ZN(u6_N91)
         );
  OAI22_X2 U975 ( .A1(n4824), .A2(n4614), .B1(n4825), .B2(n5957), .ZN(u6_N90)
         );
  OAI22_X2 U977 ( .A1(n4824), .A2(n4613), .B1(n4825), .B2(n5958), .ZN(u6_N89)
         );
  AOI22_X2 U980 ( .A1(n4825), .A2(fracta_mul[33]), .B1(n4826), .B2(N294), .ZN(
        n971) );
  OAI22_X2 U981 ( .A1(n4824), .A2(n4372), .B1(n4825), .B2(n5959), .ZN(u6_N87)
         );
  AOI22_X2 U984 ( .A1(n4825), .A2(fracta_mul[31]), .B1(n4826), .B2(N292), .ZN(
        n974) );
  OAI22_X2 U985 ( .A1(n4824), .A2(n4612), .B1(n4825), .B2(n5960), .ZN(u6_N85)
         );
  OAI22_X2 U987 ( .A1(n4824), .A2(n4373), .B1(n4825), .B2(n5961), .ZN(u6_N84)
         );
  OAI22_X2 U989 ( .A1(n4824), .A2(n4363), .B1(n4825), .B2(n5962), .ZN(u6_N83)
         );
  OAI22_X2 U991 ( .A1(n4824), .A2(n4364), .B1(n4825), .B2(n5963), .ZN(u6_N82)
         );
  OAI22_X2 U993 ( .A1(n4824), .A2(n4615), .B1(n4825), .B2(n5964), .ZN(u6_N81)
         );
  OAI22_X2 U995 ( .A1(n4824), .A2(n4376), .B1(n4825), .B2(n5965), .ZN(u6_N80)
         );
  AOI22_X2 U998 ( .A1(n4825), .A2(fracta_mul[24]), .B1(n4824), .B2(N285), .ZN(
        n986) );
  OAI22_X2 U999 ( .A1(n4824), .A2(n4356), .B1(n4825), .B2(n5966), .ZN(u6_N78)
         );
  OAI22_X2 U1001 ( .A1(n4824), .A2(n4367), .B1(n4825), .B2(n5967), .ZN(u6_N77)
         );
  OAI22_X2 U1003 ( .A1(n4824), .A2(n4377), .B1(n4825), .B2(n5968), .ZN(u6_N76)
         );
  AOI22_X2 U1006 ( .A1(n4825), .A2(fracta_mul[20]), .B1(n4826), .B2(N281), 
        .ZN(n993) );
  AOI22_X2 U1008 ( .A1(n4825), .A2(fracta_mul[19]), .B1(n4826), .B2(N280), 
        .ZN(n994) );
  OAI22_X2 U1009 ( .A1(n4824), .A2(n4616), .B1(n4825), .B2(n5969), .ZN(u6_N73)
         );
  OAI22_X2 U1011 ( .A1(n4824), .A2(n4488), .B1(n4825), .B2(n5970), .ZN(u6_N72)
         );
  OAI22_X2 U1013 ( .A1(n4824), .A2(n4489), .B1(n4825), .B2(n5971), .ZN(u6_N71)
         );
  AOI22_X2 U1016 ( .A1(n4825), .A2(fracta_mul[15]), .B1(n4826), .B2(N276), 
        .ZN(n1001) );
  OAI22_X2 U1017 ( .A1(n4824), .A2(n4496), .B1(n4825), .B2(n5972), .ZN(u6_N69)
         );
  AOI22_X2 U1020 ( .A1(n4825), .A2(fracta_mul[13]), .B1(n4826), .B2(N274), 
        .ZN(n1004) );
  OAI22_X2 U1021 ( .A1(n4824), .A2(n4491), .B1(n4825), .B2(n5973), .ZN(u6_N67)
         );
  OAI22_X2 U1023 ( .A1(n4824), .A2(n4495), .B1(n4825), .B2(n5974), .ZN(u6_N66)
         );
  AOI22_X2 U1026 ( .A1(n4825), .A2(fracta_mul[10]), .B1(n4826), .B2(N271), 
        .ZN(n1009) );
  OAI22_X2 U1027 ( .A1(n4824), .A2(n4492), .B1(n4825), .B2(n5975), .ZN(u6_N64)
         );
  AOI22_X2 U1030 ( .A1(n4825), .A2(fracta_mul[8]), .B1(n4826), .B2(N269), .ZN(
        n1012) );
  AOI22_X2 U1032 ( .A1(n4825), .A2(fracta_mul[7]), .B1(n4826), .B2(N268), .ZN(
        n1013) );
  OAI22_X2 U1033 ( .A1(n4824), .A2(n4498), .B1(n4825), .B2(n5976), .ZN(u6_N60)
         );
  AOI22_X2 U1036 ( .A1(n4825), .A2(fracta_mul[4]), .B1(n4826), .B2(N265), .ZN(
        n1016) );
  OAI22_X2 U1037 ( .A1(n4824), .A2(n4500), .B1(n4825), .B2(n5977), .ZN(u6_N58)
         );
  AOI22_X2 U1040 ( .A1(n4825), .A2(fracta_mul[2]), .B1(n4826), .B2(N263), .ZN(
        n1019) );
  OAI22_X2 U1041 ( .A1(n4824), .A2(n4497), .B1(n4825), .B2(n5978), .ZN(u6_N56)
         );
  AOI22_X2 U1044 ( .A1(n4825), .A2(fracta_mul[0]), .B1(n4826), .B2(N261), .ZN(
        n1022) );
  OAI22_X2 U1045 ( .A1(n4824), .A2(n4354), .B1(n4825), .B2(n5945), .ZN(u6_N106) );
  OAI22_X2 U1047 ( .A1(n4824), .A2(n4352), .B1(n4825), .B2(n5946), .ZN(u6_N105) );
  OAI22_X2 U1049 ( .A1(n4824), .A2(n4355), .B1(n4825), .B2(n5947), .ZN(u6_N104) );
  OAI22_X2 U1051 ( .A1(n4824), .A2(n4366), .B1(n4825), .B2(n5948), .ZN(u6_N103) );
  OAI22_X2 U1053 ( .A1(n4824), .A2(n4362), .B1(n4825), .B2(n5949), .ZN(u6_N102) );
  AOI22_X2 U1056 ( .A1(n4825), .A2(fracta_mul[46]), .B1(n4826), .B2(N307), 
        .ZN(n1033) );
  OAI22_X2 U1057 ( .A1(n4824), .A2(n4499), .B1(n4825), .B2(n5950), .ZN(u6_N100) );
  NAND2_X2 U1059 ( .A1(u6_N52), .A2(n4825), .ZN(n4123) );
  OAI22_X2 U1061 ( .A1(u2_N40), .A2(n4815), .B1(u2_N52), .B2(n4817), .ZN(n1036) );
  AOI22_X2 U1063 ( .A1(u2_N51), .A2(n4815), .B1(u2_N39), .B2(n4817), .ZN(n1037) );
  AOI22_X2 U1065 ( .A1(u2_N50), .A2(n4815), .B1(u2_N38), .B2(n4817), .ZN(n1038) );
  AOI22_X2 U1067 ( .A1(u2_N49), .A2(n4815), .B1(u2_N37), .B2(n4817), .ZN(n1039) );
  AOI22_X2 U1069 ( .A1(u2_N48), .A2(n4815), .B1(u2_N36), .B2(n4817), .ZN(n1040) );
  AOI22_X2 U1071 ( .A1(u2_N47), .A2(n4815), .B1(u2_N35), .B2(n4817), .ZN(n1041) );
  AOI22_X2 U1073 ( .A1(u2_N46), .A2(n4815), .B1(u2_N34), .B2(n4817), .ZN(n1042) );
  AOI22_X2 U1075 ( .A1(u2_N45), .A2(n4815), .B1(u2_N33), .B2(n4817), .ZN(n1043) );
  AOI22_X2 U1077 ( .A1(u2_N44), .A2(n4815), .B1(u2_N32), .B2(n4817), .ZN(n1044) );
  AOI22_X2 U1079 ( .A1(u2_N43), .A2(n4815), .B1(u2_N31), .B2(n4817), .ZN(n1045) );
  AOI22_X2 U1081 ( .A1(n1054), .A2(n4815), .B1(n1054), .B2(n4817), .ZN(n1046)
         );
  AOI22_X2 U1083 ( .A1(u2_N29), .A2(n4815), .B1(u2_N17), .B2(n4817), .ZN(n602)
         );
  AOI22_X2 U1088 ( .A1(n4816), .A2(u2_N15), .B1(n4815), .B2(u2_N27), .ZN(n1048) );
  AOI22_X2 U1090 ( .A1(n4816), .A2(u2_N14), .B1(n4815), .B2(u2_N26), .ZN(n1049) );
  AOI22_X2 U1092 ( .A1(n4816), .A2(u2_N13), .B1(n4815), .B2(u2_N25), .ZN(n1050) );
  AOI22_X2 U1094 ( .A1(n4816), .A2(u2_N12), .B1(n4815), .B2(u2_N24), .ZN(n1051) );
  AOI22_X2 U1096 ( .A1(n4816), .A2(u2_N11), .B1(n4815), .B2(u2_N23), .ZN(n1052) );
  OAI22_X2 U1097 ( .A1(n4815), .A2(n6091), .B1(n4817), .B2(n6100), .ZN(
        u2_lt_131_A_4_) );
  AOI22_X2 U1101 ( .A1(n4817), .A2(u2_N6), .B1(n4815), .B2(u2_N18), .ZN(n1054)
         );
  AOI22_X2 U1106 ( .A1(n4846), .A2(opb_r[61]), .B1(n4840), .B2(opa_r[61]), 
        .ZN(n1056) );
  AOI22_X2 U1108 ( .A1(n4846), .A2(opb_r[60]), .B1(n4840), .B2(opa_r[60]), 
        .ZN(n1057) );
  AOI22_X2 U1110 ( .A1(n4839), .A2(opb_r[61]), .B1(n4829), .B2(opa_r[61]), 
        .ZN(n779) );
  AOI22_X2 U1112 ( .A1(n4839), .A2(opb_r[60]), .B1(n4829), .B2(opa_r[60]), 
        .ZN(n780) );
  OAI22_X2 U1113 ( .A1(n4829), .A2(n4569), .B1(n4844), .B2(n4582), .ZN(n4149)
         );
  OAI22_X2 U1114 ( .A1(n4830), .A2(n4471), .B1(n4844), .B2(n4575), .ZN(n4150)
         );
  OAI22_X2 U1115 ( .A1(n4831), .A2(n4398), .B1(n4844), .B2(n4586), .ZN(n4151)
         );
  OAI22_X2 U1116 ( .A1(n4830), .A2(n4486), .B1(n4844), .B2(n4589), .ZN(n4152)
         );
  OAI22_X2 U1118 ( .A1(n4830), .A2(n4591), .B1(n4844), .B2(n4485), .ZN(n4153)
         );
  OAI22_X2 U1120 ( .A1(n4830), .A2(n4590), .B1(n4844), .B2(n4583), .ZN(n4154)
         );
  OAI22_X2 U1122 ( .A1(n4830), .A2(n4360), .B1(n4844), .B2(n4584), .ZN(n4155)
         );
  OAI22_X2 U1123 ( .A1(n4830), .A2(n4371), .B1(n4844), .B2(n4585), .ZN(n4156)
         );
  OAI22_X2 U1124 ( .A1(n4843), .A2(n4594), .B1(n4829), .B2(n4354), .ZN(n4157)
         );
  OAI22_X2 U1126 ( .A1(n4843), .A2(n4597), .B1(n4846), .B2(n4352), .ZN(n4158)
         );
  OAI22_X2 U1128 ( .A1(n4843), .A2(n4490), .B1(n4846), .B2(n4355), .ZN(n4159)
         );
  OAI22_X2 U1129 ( .A1(n4843), .A2(n4431), .B1(n4846), .B2(n4366), .ZN(n4160)
         );
  OAI22_X2 U1130 ( .A1(n4841), .A2(n4593), .B1(n4829), .B2(n4362), .ZN(n4161)
         );
  AOI22_X2 U1132 ( .A1(n4846), .A2(u6_N46), .B1(n4840), .B2(fracta_mul[46]), 
        .ZN(n1062) );
  AOI22_X2 U1134 ( .A1(n4846), .A2(u6_N45), .B1(n4840), .B2(fracta_mul[45]), 
        .ZN(n900) );
  AOI22_X2 U1136 ( .A1(n4846), .A2(u6_N44), .B1(n4840), .B2(fracta_mul[44]), 
        .ZN(n901) );
  AOI22_X2 U1138 ( .A1(n4846), .A2(u6_N43), .B1(n4840), .B2(fracta_mul[43]), 
        .ZN(n902) );
  OAI22_X2 U1139 ( .A1(n4841), .A2(n4600), .B1(n4846), .B2(n4375), .ZN(n4166)
         );
  AOI22_X2 U1142 ( .A1(n4829), .A2(u6_N41), .B1(n4840), .B2(fracta_mul[41]), 
        .ZN(n916) );
  AOI22_X2 U1144 ( .A1(n4846), .A2(u6_N40), .B1(n4840), .B2(fracta_mul[40]), 
        .ZN(n1064) );
  AOI22_X2 U1146 ( .A1(n4846), .A2(u6_N39), .B1(n4840), .B2(fracta_mul[39]), 
        .ZN(n917) );
  OAI22_X2 U1147 ( .A1(n4843), .A2(n4596), .B1(n4846), .B2(n4374), .ZN(n4170)
         );
  AOI22_X2 U1150 ( .A1(n4829), .A2(u6_N34), .B1(n4840), .B2(fracta_mul[34]), 
        .ZN(n921) );
  AOI22_X2 U1152 ( .A1(n4846), .A2(u6_N33), .B1(n4840), .B2(fracta_mul[33]), 
        .ZN(n1066) );
  OAI22_X2 U1153 ( .A1(n4841), .A2(n4595), .B1(n4829), .B2(n4372), .ZN(n4173)
         );
  OAI22_X2 U1155 ( .A1(n4839), .A2(n4603), .B1(n4832), .B2(n4363), .ZN(n4174)
         );
  OAI22_X2 U1157 ( .A1(n4841), .A2(n4607), .B1(n4832), .B2(n4364), .ZN(n4175)
         );
  AOI22_X2 U1160 ( .A1(n4829), .A2(u6_N26), .B1(n4840), .B2(fracta_mul[26]), 
        .ZN(n924) );
  OAI22_X2 U1161 ( .A1(n4841), .A2(n4605), .B1(n4829), .B2(n4376), .ZN(n4177)
         );
  AOI22_X2 U1164 ( .A1(n4829), .A2(u6_N24), .B1(n4840), .B2(fracta_mul[24]), 
        .ZN(n1071) );
  OAI22_X2 U1165 ( .A1(n4841), .A2(n4610), .B1(n4832), .B2(n4356), .ZN(n4179)
         );
  OAI22_X2 U1167 ( .A1(n4843), .A2(n4602), .B1(n4829), .B2(n4367), .ZN(n4180)
         );
  OAI22_X2 U1169 ( .A1(n4841), .A2(n4606), .B1(n4832), .B2(n4377), .ZN(n4181)
         );
  AOI22_X2 U1172 ( .A1(n4846), .A2(u6_N20), .B1(n4840), .B2(fracta_mul[20]), 
        .ZN(n1075) );
  AOI22_X2 U1174 ( .A1(n4846), .A2(u6_N19), .B1(n4840), .B2(fracta_mul[19]), 
        .ZN(n926) );
  AOI22_X2 U1176 ( .A1(n4846), .A2(u6_N18), .B1(n4840), .B2(fracta_mul[18]), 
        .ZN(n925) );
  OAI22_X2 U1177 ( .A1(n4841), .A2(n4601), .B1(n4832), .B2(n4488), .ZN(n4185)
         );
  OAI22_X2 U1179 ( .A1(n4841), .A2(n4598), .B1(n4832), .B2(n4489), .ZN(n4186)
         );
  AOI22_X2 U1182 ( .A1(n4829), .A2(u6_N15), .B1(n4840), .B2(fracta_mul[15]), 
        .ZN(n1078) );
  AOI22_X2 U1184 ( .A1(n4846), .A2(u6_N14), .B1(n4839), .B2(fracta_mul[14]), 
        .ZN(n927) );
  AOI22_X2 U1186 ( .A1(n4846), .A2(u6_N13), .B1(n4839), .B2(fracta_mul[13]), 
        .ZN(n1079) );
  OAI22_X2 U1187 ( .A1(n4841), .A2(n4609), .B1(n4832), .B2(n4491), .ZN(n4190)
         );
  AOI22_X2 U1190 ( .A1(n4829), .A2(u6_N11), .B1(n4840), .B2(fracta_mul[11]), 
        .ZN(n928) );
  AOI22_X2 U1192 ( .A1(n4829), .A2(u6_N10), .B1(n4839), .B2(fracta_mul[10]), 
        .ZN(n1081) );
  OAI22_X2 U1193 ( .A1(n4841), .A2(n4608), .B1(n4832), .B2(n4492), .ZN(n4193)
         );
  AOI22_X2 U1196 ( .A1(n4829), .A2(u6_N8), .B1(n4840), .B2(fracta_mul[8]), 
        .ZN(n1083) );
  AOI22_X2 U1198 ( .A1(n4829), .A2(u6_N7), .B1(n4839), .B2(fracta_mul[7]), 
        .ZN(n930) );
  OAI22_X2 U1200 ( .A1(u6_N6), .A2(n4843), .B1(n4832), .B2(fracta_mul[6]), 
        .ZN(n877) );
  OAI22_X2 U1202 ( .A1(u6_N5), .A2(n4842), .B1(n4832), .B2(fracta_mul[5]), 
        .ZN(n929) );
  AOI22_X2 U1204 ( .A1(n4846), .A2(u6_N4), .B1(n4839), .B2(fracta_mul[4]), 
        .ZN(n1084) );
  AOI22_X2 U1206 ( .A1(n4846), .A2(u6_N3), .B1(n4839), .B2(fracta_mul[3]), 
        .ZN(n932) );
  OAI22_X2 U1208 ( .A1(u6_N1), .A2(n4842), .B1(n4832), .B2(fracta_mul[1]), 
        .ZN(n931) );
  OAI22_X2 U1210 ( .A1(u6_N0), .A2(n4842), .B1(n4832), .B2(fracta_mul[0]), 
        .ZN(n870) );
  NAND4_X2 U1212 ( .A1(opb_r[60]), .A2(opb_r[61]), .A3(n1085), .A4(n1086), 
        .ZN(n948) );
  NOR4_X2 U1213 ( .A1(n1087), .A2(n4591), .A3(n4398), .A4(n4486), .ZN(n1086)
         );
  OAI221_X2 U1312 ( .B1(n4818), .B2(n4714), .C1(n1138), .C2(n4538), .A(n1140), 
        .ZN(n4252) );
  NAND2_X2 U1313 ( .A1(fract_i2f[0]), .A2(n4775), .ZN(n1140) );
  OAI221_X2 U1316 ( .B1(n4819), .B2(n4705), .C1(n4804), .C2(n4537), .A(n1144), 
        .ZN(n4253) );
  NAND2_X2 U1317 ( .A1(fract_i2f[2]), .A2(n4778), .ZN(n1144) );
  OAI221_X2 U1320 ( .B1(n4819), .B2(n4713), .C1(n4803), .C2(n4536), .A(n1147), 
        .ZN(n4254) );
  NAND2_X2 U1321 ( .A1(fract_i2f[3]), .A2(n4777), .ZN(n1147) );
  OAI221_X2 U1324 ( .B1(n4818), .B2(n4704), .C1(n1138), .C2(n4535), .A(n1150), 
        .ZN(n4255) );
  NAND2_X2 U1325 ( .A1(fract_i2f[5]), .A2(n4775), .ZN(n1150) );
  OAI221_X2 U1328 ( .B1(n4818), .B2(n4712), .C1(n4804), .C2(n4534), .A(n1153), 
        .ZN(n4256) );
  NAND2_X2 U1329 ( .A1(fract_i2f[6]), .A2(n4776), .ZN(n1153) );
  OAI221_X2 U1332 ( .B1(n4819), .B2(n4703), .C1(n4803), .C2(n4533), .A(n1156), 
        .ZN(n4257) );
  NAND2_X2 U1333 ( .A1(fract_i2f[8]), .A2(n4778), .ZN(n1156) );
  OAI221_X2 U1336 ( .B1(n4818), .B2(n4696), .C1(n1138), .C2(n4532), .A(n1159), 
        .ZN(n4258) );
  NAND2_X2 U1337 ( .A1(fract_i2f[10]), .A2(n4777), .ZN(n1159) );
  OAI221_X2 U1340 ( .B1(n4819), .B2(n4702), .C1(n4804), .C2(n4531), .A(n1162), 
        .ZN(n4259) );
  NAND2_X2 U1341 ( .A1(fract_i2f[11]), .A2(n4776), .ZN(n1162) );
  OAI221_X2 U1344 ( .B1(n4819), .B2(n4711), .C1(n4803), .C2(n4530), .A(n1165), 
        .ZN(n4260) );
  NAND2_X2 U1345 ( .A1(fract_i2f[16]), .A2(n4775), .ZN(n1165) );
  OAI221_X2 U1348 ( .B1(n4819), .B2(n4695), .C1(n1138), .C2(n4529), .A(n1168), 
        .ZN(n4261) );
  NAND2_X2 U1349 ( .A1(fract_i2f[17]), .A2(n4778), .ZN(n1168) );
  OAI221_X2 U1352 ( .B1(n4818), .B2(n4701), .C1(n4804), .C2(n4528), .A(n1171), 
        .ZN(n4262) );
  NAND2_X2 U1353 ( .A1(fract_i2f[18]), .A2(n4777), .ZN(n1171) );
  OAI221_X2 U1356 ( .B1(n4819), .B2(n4710), .C1(n4803), .C2(n4470), .A(n1174), 
        .ZN(n4263) );
  NAND2_X2 U1357 ( .A1(fract_i2f[21]), .A2(n4776), .ZN(n1174) );
  OAI221_X2 U1360 ( .B1(n4819), .B2(n4694), .C1(n4804), .C2(n4469), .A(n1177), 
        .ZN(n4264) );
  NAND2_X2 U1361 ( .A1(fract_i2f[22]), .A2(n4775), .ZN(n1177) );
  OAI221_X2 U1364 ( .B1(n4819), .B2(n4700), .C1(n4803), .C2(n4468), .A(n1180), 
        .ZN(n4265) );
  NAND2_X2 U1365 ( .A1(fract_i2f[23]), .A2(n4778), .ZN(n1180) );
  OAI221_X2 U1368 ( .B1(n4819), .B2(n4709), .C1(n4806), .C2(n4467), .A(n1183), 
        .ZN(n4266) );
  NAND2_X2 U1369 ( .A1(fract_i2f[28]), .A2(n4777), .ZN(n1183) );
  OAI221_X2 U1372 ( .B1(n4819), .B2(n4693), .C1(n4803), .C2(n4423), .A(n1186), 
        .ZN(n4267) );
  NAND2_X2 U1373 ( .A1(fract_i2f[29]), .A2(n4776), .ZN(n1186) );
  OAI221_X2 U1376 ( .B1(n4819), .B2(n4708), .C1(n1138), .C2(n4466), .A(n1189), 
        .ZN(n4268) );
  NAND2_X2 U1377 ( .A1(fract_i2f[33]), .A2(n4775), .ZN(n1189) );
  OAI221_X2 U1380 ( .B1(n4819), .B2(n4692), .C1(n4804), .C2(n4465), .A(n1192), 
        .ZN(n4269) );
  NAND2_X2 U1381 ( .A1(fract_i2f[34]), .A2(n4778), .ZN(n1192) );
  OAI221_X2 U1384 ( .B1(n4819), .B2(n4699), .C1(n4803), .C2(n4464), .A(n1195), 
        .ZN(n4270) );
  NAND2_X2 U1385 ( .A1(fract_i2f[35]), .A2(n4777), .ZN(n1195) );
  OAI221_X2 U1388 ( .B1(n4819), .B2(n4691), .C1(n4804), .C2(n4463), .A(n1198), 
        .ZN(n4271) );
  NAND2_X2 U1389 ( .A1(fract_i2f[40]), .A2(n4776), .ZN(n1198) );
  OAI221_X2 U1392 ( .B1(n4819), .B2(n4698), .C1(n1138), .C2(n4462), .A(n1201), 
        .ZN(n4272) );
  NAND2_X2 U1393 ( .A1(fract_i2f[41]), .A2(n4775), .ZN(n1201) );
  OAI221_X2 U1396 ( .B1(n4819), .B2(n4707), .C1(n4804), .C2(n4461), .A(n1204), 
        .ZN(n4273) );
  NAND2_X2 U1397 ( .A1(fract_i2f[46]), .A2(n4778), .ZN(n1204) );
  OAI221_X2 U1400 ( .B1(n4819), .B2(n4690), .C1(n4803), .C2(n4527), .A(n1207), 
        .ZN(n4274) );
  NAND2_X2 U1401 ( .A1(fract_i2f[47]), .A2(n4777), .ZN(n1207) );
  OAI221_X2 U1404 ( .B1(n4819), .B2(n4697), .C1(n4806), .C2(n4526), .A(n1210), 
        .ZN(n4275) );
  NAND2_X2 U1405 ( .A1(fract_i2f[48]), .A2(n4776), .ZN(n1210) );
  AOI22_X2 U1409 ( .A1(u0_snan_r_a), .A2(u0_expa_ff), .B1(u0_snan_r_b), .B2(
        u0_expb_ff), .ZN(n1211) );
  AOI22_X2 U1411 ( .A1(u0_qnan_r_a), .A2(u0_expa_ff), .B1(u0_qnan_r_b), .B2(
        u0_expb_ff), .ZN(n1212) );
  NAND2_X2 U1413 ( .A1(u0_infb_f_r), .A2(u0_expb_ff), .ZN(n943) );
  NAND2_X2 U1415 ( .A1(u0_infa_f_r), .A2(u0_expa_ff), .ZN(n944) );
  AOI22_X2 U1417 ( .A1(u3_N69), .A2(n4878), .B1(u3_N12), .B2(n4879), .ZN(n1213) );
  AOI22_X2 U1419 ( .A1(u3_N68), .A2(n4878), .B1(u3_N11), .B2(n4879), .ZN(n1215) );
  AOI22_X2 U1421 ( .A1(u3_N67), .A2(n4878), .B1(u3_N10), .B2(n4877), .ZN(n1216) );
  AOI22_X2 U1423 ( .A1(u3_N66), .A2(n4878), .B1(u3_N9), .B2(n4877), .ZN(n1217)
         );
  AOI22_X2 U1425 ( .A1(u3_N65), .A2(n4878), .B1(u3_N8), .B2(n4876), .ZN(n1218)
         );
  AOI22_X2 U1427 ( .A1(u3_N115), .A2(n4878), .B1(u3_N58), .B2(n4877), .ZN(
        n1219) );
  AOI22_X2 U1429 ( .A1(u3_N114), .A2(n4878), .B1(u3_N57), .B2(n4876), .ZN(
        n1220) );
  AOI22_X2 U1431 ( .A1(u3_N113), .A2(n4878), .B1(u3_N56), .B2(n4877), .ZN(
        n1221) );
  AOI22_X2 U1433 ( .A1(u3_N112), .A2(n4878), .B1(u3_N55), .B2(n4876), .ZN(
        n1222) );
  AOI22_X2 U1435 ( .A1(u3_N111), .A2(n4878), .B1(u3_N54), .B2(n4877), .ZN(
        n1223) );
  AOI22_X2 U1437 ( .A1(u3_N110), .A2(n4878), .B1(u3_N53), .B2(n4876), .ZN(
        n1224) );
  AOI22_X2 U1439 ( .A1(u3_N64), .A2(n4878), .B1(u3_N7), .B2(n4877), .ZN(n1225)
         );
  AOI22_X2 U1441 ( .A1(u3_N109), .A2(n4878), .B1(u3_N52), .B2(n4876), .ZN(
        n1226) );
  AOI22_X2 U1443 ( .A1(u3_N108), .A2(n4878), .B1(u3_N51), .B2(fasu_op), .ZN(
        n1227) );
  AOI22_X2 U1445 ( .A1(u3_N107), .A2(n4878), .B1(u3_N50), .B2(fasu_op), .ZN(
        n1228) );
  AOI22_X2 U1447 ( .A1(u3_N106), .A2(n4878), .B1(u3_N49), .B2(fasu_op), .ZN(
        n1229) );
  AOI22_X2 U1449 ( .A1(u3_N105), .A2(n4878), .B1(u3_N48), .B2(fasu_op), .ZN(
        n1230) );
  AOI22_X2 U1451 ( .A1(u3_N104), .A2(n4878), .B1(u3_N47), .B2(fasu_op), .ZN(
        n1231) );
  AOI22_X2 U1453 ( .A1(u3_N103), .A2(n4878), .B1(u3_N46), .B2(fasu_op), .ZN(
        n1232) );
  AOI22_X2 U1455 ( .A1(u3_N102), .A2(n4878), .B1(u3_N45), .B2(fasu_op), .ZN(
        n1233) );
  AOI22_X2 U1457 ( .A1(u3_N101), .A2(n4422), .B1(u3_N44), .B2(fasu_op), .ZN(
        n1234) );
  AOI22_X2 U1459 ( .A1(u3_N100), .A2(n4422), .B1(u3_N43), .B2(fasu_op), .ZN(
        n1235) );
  AOI22_X2 U1461 ( .A1(u3_N63), .A2(n4422), .B1(u3_N6), .B2(fasu_op), .ZN(
        n1236) );
  AOI22_X2 U1463 ( .A1(u3_N99), .A2(n4878), .B1(u3_N42), .B2(fasu_op), .ZN(
        n1237) );
  AOI22_X2 U1465 ( .A1(u3_N98), .A2(n4878), .B1(u3_N41), .B2(n4876), .ZN(n1238) );
  AOI22_X2 U1467 ( .A1(u3_N97), .A2(n4878), .B1(u3_N40), .B2(n4877), .ZN(n1239) );
  AOI22_X2 U1469 ( .A1(u3_N96), .A2(n4422), .B1(u3_N39), .B2(n4876), .ZN(n1240) );
  AOI22_X2 U1471 ( .A1(u3_N95), .A2(n4422), .B1(u3_N38), .B2(n4877), .ZN(n1241) );
  AOI22_X2 U1473 ( .A1(u3_N94), .A2(n4422), .B1(u3_N37), .B2(n4876), .ZN(n1242) );
  AOI22_X2 U1475 ( .A1(u3_N93), .A2(n4422), .B1(u3_N36), .B2(n4877), .ZN(n1243) );
  AOI22_X2 U1477 ( .A1(u3_N92), .A2(n4422), .B1(u3_N35), .B2(n4876), .ZN(n1244) );
  AOI22_X2 U1479 ( .A1(u3_N91), .A2(n4422), .B1(u3_N34), .B2(n4877), .ZN(n1245) );
  AOI22_X2 U1481 ( .A1(u3_N90), .A2(n4422), .B1(u3_N33), .B2(n4876), .ZN(n1246) );
  AOI22_X2 U1483 ( .A1(u3_N62), .A2(n4422), .B1(u3_N5), .B2(n4877), .ZN(n1247)
         );
  AOI22_X2 U1485 ( .A1(u3_N89), .A2(n4422), .B1(u3_N32), .B2(n4876), .ZN(n1248) );
  AOI22_X2 U1487 ( .A1(u3_N88), .A2(n4422), .B1(u3_N31), .B2(n4877), .ZN(n1249) );
  AOI22_X2 U1489 ( .A1(u3_N87), .A2(n4422), .B1(u3_N30), .B2(n4877), .ZN(n1250) );
  AOI22_X2 U1491 ( .A1(u3_N86), .A2(n4422), .B1(u3_N29), .B2(n4877), .ZN(n1251) );
  AOI22_X2 U1493 ( .A1(u3_N85), .A2(n4422), .B1(u3_N28), .B2(n4877), .ZN(n1252) );
  AOI22_X2 U1495 ( .A1(u3_N84), .A2(n4422), .B1(u3_N27), .B2(n4877), .ZN(n1253) );
  AOI22_X2 U1497 ( .A1(u3_N83), .A2(n4878), .B1(u3_N26), .B2(n4877), .ZN(n1254) );
  AOI22_X2 U1499 ( .A1(u3_N82), .A2(n4422), .B1(u3_N25), .B2(n4877), .ZN(n1255) );
  AOI22_X2 U1501 ( .A1(u3_N81), .A2(n4878), .B1(u3_N24), .B2(n4877), .ZN(n1256) );
  AOI22_X2 U1503 ( .A1(u3_N80), .A2(n4422), .B1(u3_N23), .B2(n4877), .ZN(n1257) );
  AOI22_X2 U1505 ( .A1(u3_N61), .A2(n4878), .B1(u3_N4), .B2(n4877), .ZN(n1258)
         );
  AOI22_X2 U1507 ( .A1(u3_N79), .A2(n4422), .B1(u3_N22), .B2(n4877), .ZN(n1259) );
  AOI22_X2 U1509 ( .A1(u3_N78), .A2(n4878), .B1(u3_N21), .B2(n4876), .ZN(n1260) );
  AOI22_X2 U1511 ( .A1(u3_N77), .A2(n4422), .B1(u3_N20), .B2(n4876), .ZN(n1261) );
  AOI22_X2 U1513 ( .A1(u3_N76), .A2(n4878), .B1(u3_N19), .B2(n4876), .ZN(n1262) );
  AOI22_X2 U1515 ( .A1(u3_N75), .A2(n4422), .B1(u3_N18), .B2(n4876), .ZN(n1263) );
  AOI22_X2 U1517 ( .A1(u3_N74), .A2(n4878), .B1(u3_N17), .B2(n4876), .ZN(n1264) );
  AOI22_X2 U1519 ( .A1(u3_N73), .A2(n4422), .B1(u3_N16), .B2(n4876), .ZN(n1265) );
  AOI22_X2 U1521 ( .A1(u3_N72), .A2(n4878), .B1(u3_N15), .B2(n4876), .ZN(n1266) );
  AOI22_X2 U1523 ( .A1(u3_N71), .A2(n4422), .B1(u3_N14), .B2(n4876), .ZN(n1267) );
  AOI22_X2 U1525 ( .A1(u3_N70), .A2(n4878), .B1(u3_N13), .B2(n4876), .ZN(n1268) );
  AOI22_X2 U1527 ( .A1(u3_N60), .A2(n4422), .B1(u3_N3), .B2(n4876), .ZN(n1269)
         );
  AOI22_X2 U1529 ( .A1(u3_N116), .A2(n4878), .B1(u3_N59), .B2(n4876), .ZN(
        n1270) );
  OAI22_X2 U1531 ( .A1(n6373), .A2(n4843), .B1(n4832), .B2(n4826), .ZN(n4348)
         );
  NAND4_X2 U1534 ( .A1(n4371), .A2(n4360), .A3(n1271), .A4(n1272), .ZN(u6_N52)
         );
  NOR4_X2 U1535 ( .A1(n1273), .A2(opb_r[60]), .A3(opb_r[62]), .A4(opb_r[61]), 
        .ZN(n1272) );
  AND2_X2 U1543 ( .A1(n947), .A2(n4354), .ZN(n4349) );
  AND4_X2 U1544 ( .A1(n1274), .A2(n1275), .A3(n1276), .A4(n1277), .ZN(n947) );
  NOR4_X2 U1545 ( .A1(n1278), .A2(n1279), .A3(fracta_mul[30]), .A4(
        fracta_mul[29]), .ZN(n1277) );
  OR3_X2 U1546 ( .A1(fracta_mul[36]), .A2(fracta_mul[37]), .A3(fracta_mul[31]), 
        .ZN(n1279) );
  NAND4_X2 U1547 ( .A1(n4355), .A2(n4352), .A3(n4366), .A4(n1280), .ZN(n1278)
         );
  NOR4_X2 U1549 ( .A1(n1281), .A2(n1282), .A3(n1283), .A4(n1284), .ZN(n1276)
         );
  NAND4_X2 U1553 ( .A1(n1286), .A2(n1287), .A3(n1288), .A4(n1289), .ZN(n946)
         );
  NOR4_X2 U1554 ( .A1(n1290), .A2(n1291), .A3(n1292), .A4(n1293), .ZN(n1289)
         );
  OR4_X2 U1555 ( .A1(u6_N10), .A2(u6_N11), .A3(u6_N0), .A4(n1294), .ZN(n1293)
         );
  OR3_X2 U1556 ( .A1(u6_N12), .A2(u6_N14), .A3(u6_N13), .ZN(n1294) );
  OR4_X2 U1557 ( .A1(u6_N16), .A2(u6_N17), .A3(u6_N15), .A4(n1295), .ZN(n1292)
         );
  OR3_X2 U1558 ( .A1(u6_N18), .A2(u6_N1), .A3(u6_N19), .ZN(n1295) );
  OR4_X2 U1559 ( .A1(u6_N21), .A2(u6_N22), .A3(u6_N20), .A4(n1296), .ZN(n1291)
         );
  OR3_X2 U1560 ( .A1(u6_N23), .A2(u6_N25), .A3(u6_N24), .ZN(n1296) );
  OR4_X2 U1561 ( .A1(u6_N27), .A2(u6_N28), .A3(u6_N26), .A4(n1297), .ZN(n1290)
         );
  OR4_X2 U1562 ( .A1(u6_N31), .A2(u6_N30), .A3(u6_N2), .A4(u6_N29), .ZN(n1297)
         );
  OR3_X2 U1564 ( .A1(u6_N50), .A2(u6_N5), .A3(u6_N4), .ZN(n1300) );
  OR4_X2 U1565 ( .A1(u6_N6), .A2(u6_N7), .A3(u6_N8), .A4(u6_N9), .ZN(n1299) );
  OR4_X2 U1566 ( .A1(u6_N45), .A2(u6_N46), .A3(u6_N44), .A4(n1301), .ZN(n1298)
         );
  NOR4_X2 U1571 ( .A1(n1302), .A2(u6_N38), .A3(u6_N3), .A4(u6_N39), .ZN(n1287)
         );
  OR4_X2 U1572 ( .A1(u6_N40), .A2(u6_N41), .A3(u6_N42), .A4(u6_N43), .ZN(n1302) );
  NOR4_X2 U1573 ( .A1(n1303), .A2(u6_N32), .A3(u6_N34), .A4(u6_N33), .ZN(n1286) );
  OR3_X2 U1574 ( .A1(u6_N36), .A2(u6_N37), .A3(u6_N35), .ZN(n1303) );
  AOI22_X2 U1576 ( .A1(n4825), .A2(fracta_mul[6]), .B1(n4826), .B2(N267), .ZN(
        n1304) );
  OR2_X2 U1578 ( .A1(N313), .A2(n4825), .ZN(u6_N107) );
  NAND4_X2 U1579 ( .A1(n4585), .A2(n4584), .A3(n1305), .A4(n1306), .ZN(u2_N157) );
  NOR4_X2 U1580 ( .A1(n1307), .A2(opa_r[60]), .A3(opa_r[62]), .A4(opa_r[61]), 
        .ZN(n1306) );
  OAI221_X2 U1588 ( .B1(n1308), .B2(n4623), .C1(n1310), .C2(n4476), .A(n1312), 
        .ZN(n2657) );
  AOI22_X2 U1589 ( .A1(exp_fasu[9]), .A2(n1313), .B1(exp_mul[9]), .B2(n1314), 
        .ZN(n1312) );
  OAI221_X2 U1590 ( .B1(n1308), .B2(n4433), .C1(n4474), .C2(n1310), .A(n1317), 
        .ZN(n2658) );
  AOI22_X2 U1591 ( .A1(exp_fasu[8]), .A2(n1313), .B1(exp_mul[8]), .B2(n1314), 
        .ZN(n1317) );
  OAI221_X2 U1593 ( .B1(n1308), .B2(n4629), .C1(n4475), .C2(n1310), .A(n1320), 
        .ZN(n2659) );
  AOI22_X2 U1594 ( .A1(exp_fasu[7]), .A2(n1313), .B1(exp_mul[7]), .B2(n1314), 
        .ZN(n1320) );
  OAI221_X2 U1596 ( .B1(n1308), .B2(n4410), .C1(n4571), .C2(n1310), .A(n1323), 
        .ZN(n2660) );
  AOI22_X2 U1597 ( .A1(exp_fasu[6]), .A2(n1313), .B1(exp_mul[6]), .B2(n1314), 
        .ZN(n1323) );
  OAI221_X2 U1598 ( .B1(n1308), .B2(n4409), .C1(n4477), .C2(n1310), .A(n1326), 
        .ZN(n2661) );
  AOI22_X2 U1599 ( .A1(exp_fasu[5]), .A2(n1313), .B1(exp_mul[5]), .B2(n1314), 
        .ZN(n1326) );
  OAI221_X2 U1600 ( .B1(n1308), .B2(n4408), .C1(n4424), .C2(n1310), .A(n1329), 
        .ZN(n2662) );
  AOI22_X2 U1601 ( .A1(exp_fasu[4]), .A2(n1313), .B1(exp_mul[4]), .B2(n1314), 
        .ZN(n1329) );
  OAI221_X2 U1602 ( .B1(n1308), .B2(n4407), .C1(n4473), .C2(n1310), .A(n1332), 
        .ZN(n2663) );
  AOI22_X2 U1603 ( .A1(exp_fasu[3]), .A2(n1313), .B1(exp_mul[3]), .B2(n1314), 
        .ZN(n1332) );
  OAI221_X2 U1604 ( .B1(n1308), .B2(n4625), .C1(n4425), .C2(n1310), .A(n1335), 
        .ZN(n2664) );
  AOI22_X2 U1605 ( .A1(exp_fasu[2]), .A2(n1313), .B1(exp_mul[2]), .B2(n1314), 
        .ZN(n1335) );
  OAI221_X2 U1606 ( .B1(n1308), .B2(n4622), .C1(n4588), .C2(n1310), .A(n1338), 
        .ZN(n2665) );
  AOI22_X2 U1607 ( .A1(exp_fasu[1]), .A2(n1313), .B1(exp_mul[1]), .B2(n1314), 
        .ZN(n1338) );
  OAI221_X2 U1608 ( .B1(n1308), .B2(n4508), .C1(n4587), .C2(n1310), .A(n1341), 
        .ZN(n2656) );
  AOI22_X2 U1609 ( .A1(exp_fasu[10]), .A2(n1313), .B1(exp_mul[10]), .B2(n1314), 
        .ZN(n1341) );
  OAI221_X2 U1610 ( .B1(n1308), .B2(n4509), .C1(n4400), .C2(n1310), .A(n1344), 
        .ZN(n2666) );
  AOI22_X2 U1611 ( .A1(exp_fasu[0]), .A2(n1313), .B1(exp_mul[0]), .B2(n1314), 
        .ZN(n1344) );
  NAND4_X2 U1615 ( .A1(n1346), .A2(n1347), .A3(n1348), .A4(n1349), .ZN(
        div_opa_ldz_d[4]) );
  NOR4_X2 U1616 ( .A1(n1350), .A2(n1351), .A3(n1352), .A4(n1353), .ZN(n1349)
         );
  NAND4_X2 U1621 ( .A1(n1358), .A2(n1347), .A3(n1359), .A4(n1360), .ZN(
        div_opa_ldz_d[3]) );
  AOI221_X2 U1622 ( .B1(n1361), .B2(n1362), .C1(n6357), .C2(fracta_mul[27]), 
        .A(n1364), .ZN(n1360) );
  NAND4_X2 U1625 ( .A1(n6353), .A2(fracta_mul[44]), .A3(n1371), .A4(n4362), 
        .ZN(n1366) );
  NAND4_X2 U1626 ( .A1(n1372), .A2(fracta_mul[28]), .A3(n4373), .A4(n4612), 
        .ZN(n1365) );
  OAI221_X2 U1627 ( .B1(n4491), .B2(n1373), .C1(n1374), .C2(n1375), .A(n1376), 
        .ZN(n1362) );
  NAND2_X2 U1628 ( .A1(n1377), .A2(n1378), .ZN(n1373) );
  AND2_X2 U1629 ( .A1(n1379), .A2(n6354), .ZN(n1359) );
  NAND4_X2 U1631 ( .A1(n1384), .A2(n1385), .A3(n1386), .A4(n1387), .ZN(
        div_opa_ldz_d[2]) );
  NOR4_X2 U1632 ( .A1(n1388), .A2(n6362), .A3(n1352), .A4(n1390), .ZN(n1387)
         );
  NAND4_X2 U1635 ( .A1(n1355), .A2(fracta_mul[32]), .A3(n1395), .A4(n4614), 
        .ZN(n1394) );
  NAND4_X2 U1636 ( .A1(n1369), .A2(fracta_mul[40]), .A3(n1396), .A4(n4617), 
        .ZN(n1392) );
  AND3_X2 U1639 ( .A1(fracta_mul[24]), .A2(n4376), .A3(n1399), .ZN(n1381) );
  OAI211_X2 U1641 ( .C1(n1400), .C2(n4489), .A(n1285), .B(n6367), .ZN(n1397)
         );
  OAI22_X2 U1643 ( .A1(n1376), .A2(n6371), .B1(n4496), .B2(n1404), .ZN(n1402)
         );
  OR3_X2 U1646 ( .A1(fracta_mul[1]), .A2(fracta_mul[2]), .A3(n1406), .ZN(n1285) );
  NAND2_X2 U1648 ( .A1(n6353), .A2(fracta_mul[46]), .ZN(n1385) );
  NAND4_X2 U1649 ( .A1(n1379), .A2(n1358), .A3(n1407), .A4(n1408), .ZN(
        div_opa_ldz_d[1]) );
  NOR4_X2 U1650 ( .A1(n1409), .A2(n1410), .A3(n6359), .A4(n1352), .ZN(n1408)
         );
  AND2_X2 U1651 ( .A1(n1372), .A2(fracta_mul[30]), .ZN(n1352) );
  AOI221_X2 U1656 ( .B1(n1416), .B2(n4354), .C1(n1361), .C2(n1417), .A(n6356), 
        .ZN(n1407) );
  AND4_X2 U1659 ( .A1(n6357), .A2(fracta_mul[22]), .A3(n1420), .A4(n4356), 
        .ZN(n1390) );
  OAI211_X2 U1660 ( .C1(n1421), .C2(n1406), .A(n1422), .B(n1423), .ZN(n1417)
         );
  NAND2_X2 U1669 ( .A1(n4352), .A2(n4355), .ZN(n1416) );
  AND4_X2 U1671 ( .A1(n1393), .A2(n1391), .A3(n1426), .A4(n1427), .ZN(n1358)
         );
  NAND2_X2 U1672 ( .A1(n1428), .A2(fracta_mul[38]), .ZN(n1391) );
  NAND4_X2 U1675 ( .A1(n1384), .A2(n1346), .A3(n1431), .A4(n1432), .ZN(
        div_opa_ldz_d[0]) );
  NOR4_X2 U1676 ( .A1(n1433), .A2(n6364), .A3(fracta_mul[51]), .A4(n1419), 
        .ZN(n1432) );
  AND3_X2 U1677 ( .A1(fracta_mul[25]), .A2(n4615), .A3(n1399), .ZN(n1419) );
  NAND4_X2 U1683 ( .A1(n1361), .A2(fracta_mul[9]), .A3(n6369), .A4(n1374), 
        .ZN(n1426) );
  AOI221_X2 U1684 ( .B1(fracta_mul[17]), .B2(n4616), .C1(fracta_mul[11]), .C2(
        n6369), .A(fracta_mul[19]), .ZN(n1436) );
  AOI22_X2 U1686 ( .A1(n1369), .A2(fracta_mul[43]), .B1(fracta_mul[49]), .B2(
        n4352), .ZN(n1431) );
  OAI22_X2 U1689 ( .A1(n6361), .A2(n1441), .B1(n1435), .B2(n4364), .ZN(n1440)
         );
  NOR4_X2 U1693 ( .A1(n6358), .A2(n4497), .A3(n1406), .A4(fracta_mul[2]), .ZN(
        n1439) );
  OR4_X2 U1694 ( .A1(n1442), .A2(fracta_mul[3]), .A3(fracta_mul[4]), .A4(
        fracta_mul[5]), .ZN(n1406) );
  AND4_X2 U1699 ( .A1(n1379), .A2(n6360), .A3(n6354), .A4(n1444), .ZN(n1384)
         );
  AOI221_X2 U1700 ( .B1(n6353), .B2(n1445), .C1(n1446), .C2(n1361), .A(n1382), 
        .ZN(n1444) );
  AND3_X2 U1701 ( .A1(fracta_mul[23]), .A2(n1420), .A3(n6357), .ZN(n1382) );
  OR2_X2 U1711 ( .A1(fracta_mul[8]), .A2(fracta_mul[9]), .ZN(n1450) );
  NAND2_X2 U1716 ( .A1(n1412), .A2(n1451), .ZN(n1357) );
  NAND4_X2 U1726 ( .A1(n1372), .A2(n4363), .A3(n4373), .A4(n4612), .ZN(n1435)
         );
  NOR4_X2 U1738 ( .A1(fracta_mul[24]), .A2(fracta_mul[25]), .A3(fracta_mul[26]), .A4(fracta_mul[27]), .ZN(n1420) );
  OR2_X2 U1741 ( .A1(n1430), .A2(fracta_mul[6]), .ZN(n1442) );
  OR2_X2 U1748 ( .A1(n1400), .A2(fracta_mul[16]), .ZN(n1404) );
  OR3_X2 U1749 ( .A1(fracta_mul[18]), .A2(fracta_mul[19]), .A3(fracta_mul[17]), 
        .ZN(n1400) );
  NAND2_X2 U1754 ( .A1(n1428), .A2(n4374), .ZN(n1354) );
  NAND2_X2 U1763 ( .A1(n1398), .A2(n4366), .ZN(n1413) );
  OR3_X2 U1766 ( .A1(fracta_mul[40]), .A2(fracta_mul[41]), .A3(n6365), .ZN(
        n1284) );
  NOR4_X2 U1769 ( .A1(n1456), .A2(n1457), .A3(n4668), .A4(n4525), .ZN(N928) );
  NAND4_X2 U1773 ( .A1(exp_mul[5]), .A2(exp_mul[6]), .A3(exp_mul[4]), .A4(
        n1460), .ZN(n1456) );
  AND3_X2 U1774 ( .A1(exp_mul[7]), .A2(exp_mul[9]), .A3(exp_mul[8]), .ZN(n1460) );
  AND4_X2 U1775 ( .A1(opb_00), .A2(opa_nan_r), .A3(n4493), .A4(n4619), .ZN(
        N918) );
  NOR4_X2 U1776 ( .A1(opa_nan), .A2(fpu_op_r2[2]), .A3(n4634), .A4(n4505), 
        .ZN(N917) );
  INV_X4 U1778 ( .A(n1464), .ZN(N916) );
  AOI221_X2 U1779 ( .B1(n1465), .B2(n6384), .C1(n1467), .C2(n1468), .A(n1469), 
        .ZN(n1464) );
  NAND2_X2 U1781 ( .A1(n1475), .A2(n4619), .ZN(n1472) );
  AOI22_X2 U1782 ( .A1(n1476), .A2(n1477), .B1(n6382), .B2(n4504), .ZN(n1471)
         );
  NAND4_X2 U1785 ( .A1(inf_d), .A2(n4773), .A3(n1468), .A4(n6398), .ZN(n1482)
         );
  AOI22_X2 U1787 ( .A1(n6382), .A2(n1486), .B1(n1468), .B2(n1487), .ZN(n1481)
         );
  NAND4_X2 U1789 ( .A1(n1491), .A2(n1492), .A3(n1493), .A4(n1494), .ZN(n1489)
         );
  NOR4_X2 U1790 ( .A1(n1495), .A2(n1496), .A3(n1497), .A4(n1498), .ZN(n1494)
         );
  NAND4_X2 U1792 ( .A1(n1502), .A2(n1503), .A3(n1504), .A4(n1505), .ZN(n1488)
         );
  NOR4_X2 U1793 ( .A1(n1506), .A2(n1507), .A3(n1508), .A4(n1509), .ZN(n1505)
         );
  OAI22_X2 U1796 ( .A1(opb_inf), .A2(n4619), .B1(opa_00), .B2(n4504), .ZN(
        n1486) );
  AOI221_X2 U1799 ( .B1(underflow_fmul_r[2]), .B2(n1521), .C1(
        underflow_fmul_r[1]), .C2(n1522), .A(n1523), .ZN(n1520) );
  OR2_X2 U1800 ( .A1(underflow_fmul_r[0]), .A2(n1524), .ZN(n1523) );
  NOR4_X2 U1801 ( .A1(n4429), .A2(n1526), .A3(n4494), .A4(n1470), .ZN(n1524)
         );
  NOR4_X2 U1802 ( .A1(n1528), .A2(n1529), .A3(n1530), .A4(n1531), .ZN(n1526)
         );
  NAND4_X2 U1803 ( .A1(n1532), .A2(n1533), .A3(n1534), .A4(n1535), .ZN(n1531)
         );
  NOR4_X2 U1804 ( .A1(n1536), .A2(prod[21]), .A3(prod[23]), .A4(prod[22]), 
        .ZN(n1535) );
  NAND4_X2 U1805 ( .A1(n4445), .A2(n4523), .A3(n4397), .A4(n4381), .ZN(n1536)
         );
  NOR4_X2 U1806 ( .A1(n1541), .A2(prod[16]), .A3(prod[18]), .A4(prod[17]), 
        .ZN(n1534) );
  NOR4_X2 U1808 ( .A1(n1545), .A2(prod[105]), .A3(prod[11]), .A4(prod[10]), 
        .ZN(n1533) );
  NAND4_X2 U1809 ( .A1(n4416), .A2(n4447), .A3(n4396), .A4(n4514), .ZN(n1545)
         );
  NOR4_X2 U1810 ( .A1(n1550), .A2(prod[0]), .A3(prod[101]), .A4(prod[100]), 
        .ZN(n1532) );
  NAND4_X2 U1812 ( .A1(n1554), .A2(n1555), .A3(n1556), .A4(n1557), .ZN(n1530)
         );
  NOR4_X2 U1813 ( .A1(n1558), .A2(prod[46]), .A3(prod[48]), .A4(prod[47]), 
        .ZN(n1557) );
  NAND4_X2 U1814 ( .A1(n4515), .A2(n4446), .A3(n4395), .A4(n4631), .ZN(n1558)
         );
  NOR4_X2 U1815 ( .A1(n1563), .A2(prod[3]), .A3(prod[41]), .A4(prod[40]), .ZN(
        n1556) );
  NAND4_X2 U1816 ( .A1(n4444), .A2(n4522), .A3(n4394), .A4(n4380), .ZN(n1563)
         );
  NOR4_X2 U1817 ( .A1(n1568), .A2(prod[33]), .A3(prod[35]), .A4(prod[34]), 
        .ZN(n1555) );
  NAND4_X2 U1818 ( .A1(n4443), .A2(n4521), .A3(n4393), .A4(n4379), .ZN(n1568)
         );
  NOR4_X2 U1819 ( .A1(n1573), .A2(prod[28]), .A3(prod[2]), .A4(prod[29]), .ZN(
        n1554) );
  NAND4_X2 U1821 ( .A1(n1577), .A2(n1578), .A3(n1579), .A4(n1580), .ZN(n1529)
         );
  NOR4_X2 U1822 ( .A1(n1581), .A2(prod[6]), .A3(prod[71]), .A4(prod[70]), .ZN(
        n1580) );
  NAND4_X2 U1823 ( .A1(n4442), .A2(n4520), .A3(n4413), .A4(n4391), .ZN(n1581)
         );
  NOR4_X2 U1824 ( .A1(n1586), .A2(prod[64]), .A3(prod[66]), .A4(prod[65]), 
        .ZN(n1579) );
  NOR4_X2 U1826 ( .A1(n1590), .A2(prod[58]), .A3(prod[5]), .A4(prod[59]), .ZN(
        n1578) );
  NAND4_X2 U1827 ( .A1(n4415), .A2(n4519), .A3(n4392), .A4(n4378), .ZN(n1590)
         );
  NOR4_X2 U1828 ( .A1(n1595), .A2(prod[52]), .A3(prod[54]), .A4(prod[53]), 
        .ZN(n1577) );
  NAND4_X2 U1830 ( .A1(n1599), .A2(n1600), .A3(n1601), .A4(n1602), .ZN(n1528)
         );
  NOR4_X2 U1831 ( .A1(n1603), .A2(prod[94]), .A3(prod[96]), .A4(prod[95]), 
        .ZN(n1602) );
  NAND4_X2 U1832 ( .A1(n4441), .A2(n4518), .A3(n4412), .A4(n4390), .ZN(n1603)
         );
  NOR4_X2 U1833 ( .A1(n1608), .A2(prod[88]), .A3(prod[8]), .A4(prod[89]), .ZN(
        n1601) );
  NAND4_X2 U1834 ( .A1(n4440), .A2(n4517), .A3(n4411), .A4(n4389), .ZN(n1608)
         );
  NOR4_X2 U1835 ( .A1(n1613), .A2(prod[81]), .A3(prod[83]), .A4(prod[82]), 
        .ZN(n1600) );
  NAND4_X2 U1836 ( .A1(n4414), .A2(n4516), .A3(n4439), .A4(n4388), .ZN(n1613)
         );
  NOR4_X2 U1837 ( .A1(n1618), .A2(prod[76]), .A3(prod[78]), .A4(prod[77]), 
        .ZN(n1599) );
  NAND4_X2 U1840 ( .A1(n1625), .A2(n1626), .A3(n1627), .A4(n1628), .ZN(n1624)
         );
  NOR4_X2 U1841 ( .A1(n1629), .A2(n1630), .A3(n1631), .A4(n1632), .ZN(n1628)
         );
  NAND4_X2 U1844 ( .A1(n1491), .A2(n1492), .A3(n1493), .A4(n1639), .ZN(n1623)
         );
  NAND4_X2 U1848 ( .A1(n1500), .A2(n1502), .A3(n1645), .A4(n1646), .ZN(n1622)
         );
  NOR4_X2 U1849 ( .A1(n1647), .A2(n1648), .A3(n1509), .A4(n1507), .ZN(n1646)
         );
  INV_X4 U1854 ( .A(n1522), .ZN(n1518) );
  NAND2_X2 U1858 ( .A1(n4820), .A2(n6399), .ZN(n1653) );
  OAI211_X2 U1859 ( .C1(n1659), .C2(n4351), .A(n1661), .B(n1662), .ZN(N894) );
  OR3_X2 U1860 ( .A1(n1517), .A2(n1663), .A3(n1664), .ZN(n1662) );
  OAI211_X2 U1863 ( .C1(n1668), .C2(n1669), .A(n4493), .B(n6388), .ZN(n1667)
         );
  NAND2_X2 U1865 ( .A1(n1490), .A2(n1470), .ZN(n1668) );
  INV_X4 U1869 ( .A(n1659), .ZN(n1675) );
  NAND4_X2 U1875 ( .A1(n1687), .A2(n1688), .A3(n1689), .A4(n1690), .ZN(n1522)
         );
  NAND4_X2 U1876 ( .A1(n1691), .A2(n1692), .A3(n1685), .A4(n1693), .ZN(n1690)
         );
  NAND4_X2 U1884 ( .A1(n294), .A2(n4587), .A3(u4_N6275), .A4(n1709), .ZN(n1707) );
  NAND4_X2 U1886 ( .A1(n4477), .A2(n4571), .A3(n4424), .A4(n1710), .ZN(n1706)
         );
  XOR2_X2 U1890 ( .A(n4875), .B(n1715), .Z(n1714) );
  AND4_X2 U1891 ( .A1(n1716), .A2(n1717), .A3(n1718), .A4(n1719), .ZN(n1713)
         );
  AND4_X2 U1892 ( .A1(n1720), .A2(n1721), .A3(n1722), .A4(n6527), .ZN(n1712)
         );
  NAND4_X2 U1896 ( .A1(n1625), .A2(n1725), .A3(n1726), .A4(n1727), .ZN(n1691)
         );
  NOR4_X2 U1897 ( .A1(n1728), .A2(n1635), .A3(n1729), .A4(n1730), .ZN(n1727)
         );
  NAND4_X2 U1900 ( .A1(n4820), .A2(n1732), .A3(n1696), .A4(n1733), .ZN(n1689)
         );
  NAND4_X2 U1901 ( .A1(n4401), .A2(n6520), .A3(n1735), .A4(n1736), .ZN(n1733)
         );
  NAND4_X2 U1903 ( .A1(n6386), .A2(n1737), .A3(n1739), .A4(n6459), .ZN(n1688)
         );
  INV_X4 U1905 ( .A(n1743), .ZN(n1742) );
  OAI222_X2 U1907 ( .A1(n1745), .A2(n1746), .B1(n4821), .B2(n6402), .C1(n6161), 
        .C2(n1749), .ZN(n1744) );
  AND3_X2 U1908 ( .A1(n1750), .A2(n1751), .A3(n1752), .ZN(n1746) );
  INV_X4 U1909 ( .A(n1696), .ZN(n1752) );
  NAND4_X2 U1910 ( .A1(rmode_r3[1]), .A2(rmode_r3[0]), .A3(n6377), .A4(n4587), 
        .ZN(n1751) );
  OAI211_X2 U1911 ( .C1(n4574), .C2(n4587), .A(n1755), .B(n1741), .ZN(n1750)
         );
  NAND4_X2 U1913 ( .A1(n1467), .A2(n1468), .A3(opas_r2), .A4(n6376), .ZN(n1757) );
  AOI22_X2 U1914 ( .A1(n1759), .A2(n1480), .B1(n6388), .B2(n1760), .ZN(n1756)
         );
  XOR2_X2 U1915 ( .A(sign_mul_r), .B(n1761), .Z(n1760) );
  AOI22_X2 U1918 ( .A1(opb_00), .A2(opa_inf), .B1(opa_00), .B2(opb_inf), .ZN(
        n1673) );
  NAND2_X2 U1920 ( .A1(n1468), .A2(n4820), .ZN(n1480) );
  OAI22_X2 U1921 ( .A1(n1763), .A2(n1473), .B1(n6382), .B2(n1764), .ZN(n1759)
         );
  AOI22_X2 U1922 ( .A1(n6397), .A2(n1766), .B1(nan_sign_d), .B2(n1767), .ZN(
        n1764) );
  INV_X4 U1923 ( .A(n1768), .ZN(n1766) );
  AOI22_X2 U1924 ( .A1(sign_fasu_r), .A2(n1769), .B1(result_zero_sign_d), .B2(
        n1465), .ZN(n1768) );
  INV_X4 U1925 ( .A(n1465), .ZN(n1769) );
  NAND2_X2 U1927 ( .A1(n1468), .A2(n4621), .ZN(n1517) );
  NAND2_X2 U1930 ( .A1(n1468), .A2(n4626), .ZN(n1767) );
  NAND2_X2 U1932 ( .A1(n1468), .A2(n4822), .ZN(n1473) );
  AOI22_X2 U1933 ( .A1(n1771), .A2(n4667), .B1(sign_mul_r), .B2(n1773), .ZN(
        n1763) );
  NAND2_X2 U1935 ( .A1(n1773), .A2(n1475), .ZN(n1771) );
  NAND4_X2 U1938 ( .A1(n1774), .A2(n1775), .A3(n1776), .A4(n1777), .ZN(n1470)
         );
  NOR4_X2 U1939 ( .A1(n1778), .A2(n1779), .A3(n1780), .A4(n1781), .ZN(n1777)
         );
  NAND4_X2 U1940 ( .A1(n1625), .A2(n1626), .A3(n1491), .A4(n1725), .ZN(n1781)
         );
  AND4_X2 U1941 ( .A1(n1782), .A2(n1783), .A3(n1784), .A4(n1785), .ZN(n1491)
         );
  NOR4_X2 U1942 ( .A1(n1786), .A2(n1787), .A3(n1788), .A4(n1789), .ZN(n1785)
         );
  NAND4_X2 U1943 ( .A1(n1790), .A2(n1791), .A3(n1792), .A4(n1729), .ZN(n1780)
         );
  NAND4_X2 U1944 ( .A1(n1730), .A2(n1492), .A3(n1793), .A4(n1794), .ZN(n1779)
         );
  NAND4_X2 U1945 ( .A1(n1795), .A2(n1796), .A3(n1797), .A4(n1641), .ZN(n1778)
         );
  NOR4_X2 U1946 ( .A1(n1798), .A2(n1799), .A3(n1800), .A4(n1509), .ZN(n1776)
         );
  NAND4_X2 U1947 ( .A1(n1801), .A2(n1802), .A3(n1803), .A4(n1804), .ZN(n1509)
         );
  NOR4_X2 U1948 ( .A1(n1805), .A2(n1806), .A3(n1807), .A4(n1808), .ZN(n1804)
         );
  NAND4_X2 U1949 ( .A1(n1809), .A2(n1810), .A3(n1811), .A4(n1812), .ZN(n1805)
         );
  NOR4_X2 U1950 ( .A1(n1813), .A2(n1814), .A3(n1815), .A4(n1816), .ZN(n1803)
         );
  NOR4_X2 U1952 ( .A1(n1820), .A2(n1821), .A3(n1822), .A4(n1823), .ZN(n1802)
         );
  NAND4_X2 U1953 ( .A1(n1824), .A2(n1825), .A3(n1826), .A4(n1827), .ZN(n1820)
         );
  NOR4_X2 U1954 ( .A1(n1828), .A2(n1829), .A3(n1830), .A4(n1831), .ZN(n1801)
         );
  NAND2_X2 U1956 ( .A1(n1633), .A2(n1634), .ZN(n1799) );
  NAND4_X2 U1957 ( .A1(n1512), .A2(n1510), .A3(n1511), .A4(n1835), .ZN(n1798)
         );
  NOR4_X2 U1958 ( .A1(n1514), .A2(n1515), .A3(n1513), .A4(n1650), .ZN(n1775)
         );
  NOR4_X2 U1959 ( .A1(n1836), .A2(n1837), .A3(n1838), .A4(n1839), .ZN(n1774)
         );
  NAND2_X2 U1960 ( .A1(n1625), .A2(n1840), .ZN(N860) );
  NAND2_X2 U1961 ( .A1(n1790), .A2(n1840), .ZN(N859) );
  INV_X4 U1962 ( .A(n1638), .ZN(n1790) );
  NAND2_X2 U1963 ( .A1(n1725), .A2(n1840), .ZN(N858) );
  NAND2_X2 U1964 ( .A1(n1840), .A2(n1633), .ZN(N857) );
  NAND2_X2 U1965 ( .A1(n1840), .A2(n1634), .ZN(N856) );
  NAND2_X2 U1966 ( .A1(n1840), .A2(n1635), .ZN(N855) );
  NAND2_X2 U1967 ( .A1(n1729), .A2(n1840), .ZN(N854) );
  INV_X4 U1968 ( .A(n1632), .ZN(n1729) );
  NAND2_X2 U1969 ( .A1(n1730), .A2(n1840), .ZN(N853) );
  INV_X4 U1970 ( .A(n1631), .ZN(n1730) );
  NAND2_X2 U1971 ( .A1(n1792), .A2(n1840), .ZN(N852) );
  INV_X4 U1972 ( .A(n1630), .ZN(n1792) );
  NAND2_X2 U1973 ( .A1(n1791), .A2(n1840), .ZN(N851) );
  INV_X4 U1974 ( .A(n1637), .ZN(n1791) );
  NAND2_X2 U1975 ( .A1(n1626), .A2(n1840), .ZN(N850) );
  AND2_X2 U1977 ( .A1(n1842), .A2(n4797), .ZN(n1812) );
  AOI22_X2 U1978 ( .A1(n4796), .A2(u4_fract_out_51_), .B1(u4_fract_out_pl1_51_), .B2(n4793), .ZN(n1842) );
  INV_X4 U1979 ( .A(n1846), .ZN(u4_fract_out_51_) );
  AND2_X2 U1981 ( .A1(n1847), .A2(n4799), .ZN(n1811) );
  AOI22_X2 U1982 ( .A1(n4796), .A2(u4_fract_out_50_), .B1(u4_fract_out_pl1_50_), .B2(n4793), .ZN(n1847) );
  INV_X4 U1983 ( .A(n1848), .ZN(u4_fract_out_50_) );
  AND2_X2 U1985 ( .A1(n1849), .A2(n4799), .ZN(n1810) );
  AOI22_X2 U1986 ( .A1(n4796), .A2(u4_fract_out_49_), .B1(u4_fract_out_pl1_49_), .B2(n4793), .ZN(n1849) );
  AND2_X2 U1988 ( .A1(n1850), .A2(n4799), .ZN(n1809) );
  AOI22_X2 U1989 ( .A1(n4796), .A2(u4_fract_out_48_), .B1(u4_fract_out_pl1_48_), .B2(n4793), .ZN(n1850) );
  AND2_X2 U1990 ( .A1(n1807), .A2(n1840), .ZN(N845) );
  NAND2_X2 U1991 ( .A1(n1851), .A2(n4799), .ZN(n1807) );
  AOI22_X2 U1992 ( .A1(n4795), .A2(u4_fract_out_47_), .B1(u4_fract_out_pl1_47_), .B2(n4793), .ZN(n1851) );
  INV_X4 U1993 ( .A(n1852), .ZN(u4_fract_out_47_) );
  AND2_X2 U1994 ( .A1(n1808), .A2(n4801), .ZN(N844) );
  NAND2_X2 U1995 ( .A1(n1853), .A2(n4799), .ZN(n1808) );
  AOI22_X2 U1996 ( .A1(n4795), .A2(u4_fract_out_46_), .B1(u4_fract_out_pl1_46_), .B2(n4793), .ZN(n1853) );
  INV_X4 U1997 ( .A(n1854), .ZN(u4_fract_out_46_) );
  AND2_X2 U1998 ( .A1(n1806), .A2(n4801), .ZN(N843) );
  NAND2_X2 U1999 ( .A1(n1855), .A2(n4799), .ZN(n1806) );
  AOI22_X2 U2000 ( .A1(n4796), .A2(u4_fract_out_45_), .B1(u4_fract_out_pl1_45_), .B2(n4793), .ZN(n1855) );
  INV_X4 U2001 ( .A(n1856), .ZN(u4_fract_out_45_) );
  AND2_X2 U2003 ( .A1(n1857), .A2(n4798), .ZN(n1818) );
  AOI22_X2 U2004 ( .A1(n4795), .A2(u4_fract_out_44_), .B1(u4_fract_out_pl1_44_), .B2(n4793), .ZN(n1857) );
  AND2_X2 U2006 ( .A1(n1858), .A2(n4798), .ZN(n1817) );
  AOI22_X2 U2007 ( .A1(n4795), .A2(u4_fract_out_43_), .B1(u4_fract_out_pl1_43_), .B2(n4793), .ZN(n1858) );
  AND2_X2 U2009 ( .A1(n1859), .A2(n4798), .ZN(n1819) );
  AOI22_X2 U2010 ( .A1(n4795), .A2(u4_fract_out_42_), .B1(u4_fract_out_pl1_42_), .B2(n4793), .ZN(n1859) );
  AND2_X2 U2011 ( .A1(n1815), .A2(n4801), .ZN(N839) );
  NAND2_X2 U2012 ( .A1(n1860), .A2(n4799), .ZN(n1815) );
  AOI22_X2 U2013 ( .A1(n4796), .A2(u4_fract_out_41_), .B1(u4_fract_out_pl1_41_), .B2(n4793), .ZN(n1860) );
  AND2_X2 U2014 ( .A1(n1816), .A2(n4801), .ZN(N838) );
  NAND2_X2 U2015 ( .A1(n1861), .A2(n4799), .ZN(n1816) );
  AOI22_X2 U2016 ( .A1(n4795), .A2(u4_fract_out_40_), .B1(u4_fract_out_pl1_40_), .B2(n4793), .ZN(n1861) );
  INV_X4 U2017 ( .A(n1862), .ZN(u4_fract_out_40_) );
  AND2_X2 U2018 ( .A1(n1814), .A2(n4801), .ZN(N837) );
  NAND2_X2 U2019 ( .A1(n1863), .A2(n4799), .ZN(n1814) );
  AOI22_X2 U2020 ( .A1(n4795), .A2(u4_fract_out_39_), .B1(u4_fract_out_pl1_39_), .B2(n4793), .ZN(n1863) );
  INV_X4 U2021 ( .A(n1864), .ZN(u4_fract_out_39_) );
  AND2_X2 U2023 ( .A1(n1865), .A2(n4798), .ZN(n1827) );
  AOI22_X2 U2024 ( .A1(n4795), .A2(u4_fract_out_38_), .B1(u4_fract_out_pl1_38_), .B2(n4793), .ZN(n1865) );
  AND2_X2 U2026 ( .A1(n1866), .A2(n4798), .ZN(n1826) );
  AOI22_X2 U2027 ( .A1(n4795), .A2(u4_fract_out_37_), .B1(u4_fract_out_pl1_37_), .B2(n4793), .ZN(n1866) );
  AND2_X2 U2029 ( .A1(n1867), .A2(n4798), .ZN(n1825) );
  AOI22_X2 U2030 ( .A1(n4795), .A2(u4_fract_out_36_), .B1(u4_fract_out_pl1_36_), .B2(n4793), .ZN(n1867) );
  AND2_X2 U2032 ( .A1(n1868), .A2(n4798), .ZN(n1824) );
  AOI22_X2 U2033 ( .A1(n4795), .A2(u4_fract_out_35_), .B1(u4_fract_out_pl1_35_), .B2(n4793), .ZN(n1868) );
  INV_X4 U2034 ( .A(n1869), .ZN(u4_fract_out_35_) );
  AND2_X2 U2035 ( .A1(n1822), .A2(n4801), .ZN(N832) );
  NAND2_X2 U2036 ( .A1(n1870), .A2(n4799), .ZN(n1822) );
  AOI22_X2 U2037 ( .A1(n4795), .A2(u4_fract_out_34_), .B1(u4_fract_out_pl1_34_), .B2(n4793), .ZN(n1870) );
  INV_X4 U2038 ( .A(n1871), .ZN(u4_fract_out_34_) );
  AND2_X2 U2039 ( .A1(n1823), .A2(n1840), .ZN(N831) );
  NAND2_X2 U2040 ( .A1(n1872), .A2(n4799), .ZN(n1823) );
  AOI22_X2 U2041 ( .A1(n4795), .A2(u4_fract_out_33_), .B1(u4_fract_out_pl1_33_), .B2(n4793), .ZN(n1872) );
  INV_X4 U2042 ( .A(n1873), .ZN(u4_fract_out_33_) );
  AND2_X2 U2043 ( .A1(n1821), .A2(n1840), .ZN(N830) );
  NAND2_X2 U2044 ( .A1(n1874), .A2(n4799), .ZN(n1821) );
  AOI22_X2 U2045 ( .A1(n4795), .A2(u4_fract_out_32_), .B1(u4_fract_out_pl1_32_), .B2(n4793), .ZN(n1874) );
  AND2_X2 U2047 ( .A1(n1875), .A2(n4798), .ZN(n1833) );
  AOI22_X2 U2048 ( .A1(n4795), .A2(u4_fract_out_31_), .B1(u4_fract_out_pl1_31_), .B2(n4793), .ZN(n1875) );
  AND2_X2 U2050 ( .A1(n1876), .A2(n4799), .ZN(n1832) );
  AOI22_X2 U2051 ( .A1(n4795), .A2(u4_fract_out_30_), .B1(u4_fract_out_pl1_30_), .B2(n4793), .ZN(n1876) );
  AND2_X2 U2053 ( .A1(n1877), .A2(n4798), .ZN(n1834) );
  AOI22_X2 U2054 ( .A1(n4795), .A2(u4_fract_out_29_), .B1(u4_fract_out_pl1_29_), .B2(n4794), .ZN(n1877) );
  INV_X4 U2055 ( .A(n1878), .ZN(u4_fract_out_29_) );
  AND2_X2 U2056 ( .A1(n1830), .A2(n1840), .ZN(N826) );
  NAND2_X2 U2057 ( .A1(n1879), .A2(n4798), .ZN(n1830) );
  AOI22_X2 U2058 ( .A1(n4795), .A2(u4_fract_out_28_), .B1(u4_fract_out_pl1_28_), .B2(n4794), .ZN(n1879) );
  INV_X4 U2059 ( .A(n1880), .ZN(u4_fract_out_28_) );
  AND2_X2 U2060 ( .A1(n1831), .A2(n1840), .ZN(N825) );
  NAND2_X2 U2061 ( .A1(n1881), .A2(n4798), .ZN(n1831) );
  AOI22_X2 U2062 ( .A1(n4795), .A2(u4_fract_out_27_), .B1(u4_fract_out_pl1_27_), .B2(n4794), .ZN(n1881) );
  INV_X4 U2063 ( .A(n1882), .ZN(u4_fract_out_27_) );
  AND2_X2 U2064 ( .A1(n1829), .A2(n1840), .ZN(N824) );
  NAND2_X2 U2065 ( .A1(n1883), .A2(n4798), .ZN(n1829) );
  AOI22_X2 U2066 ( .A1(n4795), .A2(u4_fract_out_26_), .B1(u4_fract_out_pl1_26_), .B2(n4794), .ZN(n1883) );
  INV_X4 U2068 ( .A(n1507), .ZN(n1835) );
  NAND2_X2 U2069 ( .A1(n1884), .A2(n4798), .ZN(n1507) );
  AOI22_X2 U2070 ( .A1(n4795), .A2(u4_fract_out_25_), .B1(u4_fract_out_pl1_25_), .B2(n4794), .ZN(n1884) );
  INV_X4 U2072 ( .A(n1648), .ZN(n1511) );
  NAND2_X2 U2073 ( .A1(n1885), .A2(n4798), .ZN(n1648) );
  AOI22_X2 U2074 ( .A1(n4795), .A2(u4_fract_out_24_), .B1(u4_fract_out_pl1_24_), .B2(n4794), .ZN(n1885) );
  AND2_X2 U2076 ( .A1(n1886), .A2(n4799), .ZN(n1510) );
  AOI22_X2 U2077 ( .A1(n4795), .A2(u4_fract_out_23_), .B1(u4_fract_out_pl1_23_), .B2(n4794), .ZN(n1886) );
  INV_X4 U2078 ( .A(n1887), .ZN(u4_fract_out_23_) );
  AND2_X2 U2080 ( .A1(n1888), .A2(n4798), .ZN(n1512) );
  AOI22_X2 U2081 ( .A1(n4795), .A2(u4_fract_out_22_), .B1(u4_fract_out_pl1_22_), .B2(n4794), .ZN(n1888) );
  INV_X4 U2082 ( .A(n1889), .ZN(u4_fract_out_22_) );
  INV_X4 U2084 ( .A(n1514), .ZN(n1649) );
  NAND2_X2 U2085 ( .A1(n1890), .A2(n4798), .ZN(n1514) );
  AOI22_X2 U2086 ( .A1(n4795), .A2(u4_fract_out_21_), .B1(u4_fract_out_pl1_21_), .B2(n4794), .ZN(n1890) );
  INV_X4 U2087 ( .A(n1891), .ZN(u4_fract_out_21_) );
  AND2_X2 U2088 ( .A1(n1515), .A2(n1840), .ZN(N818) );
  NAND2_X2 U2089 ( .A1(n1892), .A2(n4798), .ZN(n1515) );
  AOI22_X2 U2090 ( .A1(n4796), .A2(u4_fract_out_20_), .B1(u4_fract_out_pl1_20_), .B2(n4794), .ZN(n1892) );
  AND2_X2 U2091 ( .A1(n1786), .A2(n1840), .ZN(N817) );
  NAND2_X2 U2092 ( .A1(n1893), .A2(n4798), .ZN(n1786) );
  AOI22_X2 U2093 ( .A1(n4795), .A2(u4_fract_out_19_), .B1(u4_fract_out_pl1_19_), .B2(n4794), .ZN(n1893) );
  AND2_X2 U2094 ( .A1(n1787), .A2(n1840), .ZN(N816) );
  NAND2_X2 U2095 ( .A1(n1894), .A2(n4798), .ZN(n1787) );
  AOI22_X2 U2096 ( .A1(n4796), .A2(u4_fract_out_18_), .B1(u4_fract_out_pl1_18_), .B2(n4794), .ZN(n1894) );
  AND2_X2 U2097 ( .A1(n1788), .A2(n1840), .ZN(N815) );
  NAND2_X2 U2098 ( .A1(n1895), .A2(n4798), .ZN(n1788) );
  AOI22_X2 U2099 ( .A1(n4796), .A2(u4_fract_out_17_), .B1(u4_fract_out_pl1_17_), .B2(n4794), .ZN(n1895) );
  INV_X4 U2100 ( .A(n1896), .ZN(u4_fract_out_17_) );
  AND2_X2 U2101 ( .A1(n1789), .A2(n1840), .ZN(N814) );
  NAND2_X2 U2102 ( .A1(n1897), .A2(n4798), .ZN(n1789) );
  AOI22_X2 U2103 ( .A1(n4796), .A2(u4_fract_out_16_), .B1(u4_fract_out_pl1_16_), .B2(n4794), .ZN(n1897) );
  INV_X4 U2104 ( .A(n1898), .ZN(u4_fract_out_16_) );
  AND2_X2 U2106 ( .A1(n1899), .A2(n4798), .ZN(n1783) );
  AOI22_X2 U2107 ( .A1(n4796), .A2(u4_fract_out_15_), .B1(u4_fract_out_pl1_15_), .B2(n4794), .ZN(n1899) );
  INV_X4 U2108 ( .A(n1900), .ZN(u4_fract_out_15_) );
  AND2_X2 U2110 ( .A1(n1901), .A2(n4798), .ZN(n1782) );
  AOI22_X2 U2111 ( .A1(n4796), .A2(u4_fract_out_14_), .B1(u4_fract_out_pl1_14_), .B2(n4794), .ZN(n1901) );
  AND2_X2 U2113 ( .A1(n1902), .A2(n4798), .ZN(n1784) );
  AOI22_X2 U2114 ( .A1(n4796), .A2(u4_fract_out_13_), .B1(u4_fract_out_pl1_13_), .B2(n4794), .ZN(n1902) );
  AND2_X2 U2115 ( .A1(n1513), .A2(n1840), .ZN(N810) );
  NAND2_X2 U2116 ( .A1(n1903), .A2(n4799), .ZN(n1513) );
  AOI22_X2 U2117 ( .A1(n4796), .A2(u4_fract_out_12_), .B1(u4_fract_out_pl1_12_), .B2(n4794), .ZN(n1903) );
  INV_X4 U2119 ( .A(n1650), .ZN(n1503) );
  NAND2_X2 U2120 ( .A1(n1904), .A2(n4797), .ZN(n1650) );
  AOI22_X2 U2121 ( .A1(n4796), .A2(u4_fract_out_11_), .B1(u4_fract_out_pl1_11_), .B2(n4794), .ZN(n1904) );
  INV_X4 U2122 ( .A(n1905), .ZN(u4_fract_out_11_) );
  INV_X4 U2124 ( .A(n1836), .ZN(n1502) );
  NAND2_X2 U2125 ( .A1(n1906), .A2(n4797), .ZN(n1836) );
  AOI22_X2 U2126 ( .A1(n4796), .A2(u4_fract_out_10_), .B1(u4_fract_out_pl1_10_), .B2(n4794), .ZN(n1906) );
  INV_X4 U2127 ( .A(n1907), .ZN(u4_fract_out_10_) );
  INV_X4 U2129 ( .A(n1837), .ZN(n1500) );
  NAND2_X2 U2130 ( .A1(n1908), .A2(n4797), .ZN(n1837) );
  AOI22_X2 U2131 ( .A1(n4796), .A2(u4_fract_out_9_), .B1(u4_fract_out_pl1_9_), 
        .B2(n4793), .ZN(n1908) );
  INV_X4 U2133 ( .A(n1838), .ZN(n1499) );
  NAND2_X2 U2134 ( .A1(n1909), .A2(n4797), .ZN(n1838) );
  AOI22_X2 U2135 ( .A1(n4796), .A2(u4_fract_out_8_), .B1(u4_fract_out_pl1_8_), 
        .B2(n4794), .ZN(n1909) );
  INV_X4 U2137 ( .A(n1839), .ZN(n1501) );
  NAND2_X2 U2138 ( .A1(n1910), .A2(n4797), .ZN(n1839) );
  AOI22_X2 U2139 ( .A1(n4796), .A2(u4_fract_out_7_), .B1(u4_fract_out_pl1_7_), 
        .B2(n4793), .ZN(n1910) );
  INV_X4 U2141 ( .A(n1497), .ZN(n1641) );
  NAND2_X2 U2142 ( .A1(n1911), .A2(n4797), .ZN(n1497) );
  AOI22_X2 U2143 ( .A1(n4796), .A2(u4_fract_out_6_), .B1(u4_fract_out_pl1_6_), 
        .B2(n4794), .ZN(n1911) );
  INV_X4 U2145 ( .A(n1498), .ZN(n1797) );
  NAND2_X2 U2146 ( .A1(n1912), .A2(n4797), .ZN(n1498) );
  AOI22_X2 U2147 ( .A1(n4796), .A2(u4_fract_out_5_), .B1(u4_fract_out_pl1_5_), 
        .B2(n4793), .ZN(n1912) );
  INV_X4 U2148 ( .A(n1913), .ZN(u4_fract_out_5_) );
  INV_X4 U2150 ( .A(n1496), .ZN(n1796) );
  NAND2_X2 U2151 ( .A1(n1914), .A2(n4797), .ZN(n1496) );
  AOI22_X2 U2152 ( .A1(n4796), .A2(u4_fract_out_4_), .B1(u4_fract_out_pl1_4_), 
        .B2(n4793), .ZN(n1914) );
  INV_X4 U2154 ( .A(n1643), .ZN(n1795) );
  NAND2_X2 U2155 ( .A1(n1915), .A2(n4797), .ZN(n1643) );
  AOI22_X2 U2156 ( .A1(n4796), .A2(u4_fract_out_3_), .B1(u4_fract_out_pl1_3_), 
        .B2(n4794), .ZN(n1915) );
  INV_X4 U2157 ( .A(n1916), .ZN(u4_fract_out_3_) );
  INV_X4 U2159 ( .A(n1644), .ZN(n1794) );
  NAND2_X2 U2160 ( .A1(n1917), .A2(n4797), .ZN(n1644) );
  AOI22_X2 U2161 ( .A1(n4796), .A2(u4_fract_out_2_), .B1(u4_fract_out_pl1_2_), 
        .B2(n4793), .ZN(n1917) );
  INV_X4 U2163 ( .A(n1642), .ZN(n1793) );
  NAND2_X2 U2164 ( .A1(n1918), .A2(n4797), .ZN(n1642) );
  AOI22_X2 U2165 ( .A1(n4796), .A2(u4_fract_out_1_), .B1(u4_fract_out_pl1_1_), 
        .B2(n4793), .ZN(n1918) );
  OAI22_X2 U2166 ( .A1(n1492), .A2(n4802), .B1(n6383), .B2(n4801), .ZN(N798)
         );
  OAI211_X2 U2168 ( .C1(n4619), .C2(n1920), .A(n1468), .B(n1921), .ZN(n1919)
         );
  AOI221_X2 U2169 ( .B1(n6392), .B2(n4822), .C1(n1923), .C2(opb_inf), .A(n1485), .ZN(n1921) );
  NAND2_X2 U2174 ( .A1(opa_00), .A2(opb_00), .ZN(n1475) );
  NAND2_X2 U2176 ( .A1(n1924), .A2(n1925), .ZN(n1840) );
  OAI211_X2 U2177 ( .C1(n4819), .C2(n1674), .A(n1468), .B(n1926), .ZN(n1924)
         );
  NAND2_X2 U2184 ( .A1(n6399), .A2(n5046), .ZN(n1674) );
  AND2_X2 U2187 ( .A1(n1930), .A2(n4798), .ZN(n1492) );
  INV_X4 U2192 ( .A(n1938), .ZN(n1934) );
  AOI22_X2 U2194 ( .A1(n4796), .A2(u4_fract_out_0_), .B1(u4_fract_out_pl1_0_), 
        .B2(n4793), .ZN(n1930) );
  OAI221_X2 U2198 ( .B1(r482_B_0_), .B2(n1944), .C1(n4427), .C2(n1946), .A(
        n1671), .ZN(n1943) );
  OR4_X2 U2201 ( .A1(n1634), .A2(n1633), .A3(n1948), .A4(n1949), .ZN(n1508) );
  OR4_X2 U2202 ( .A1(n1950), .A2(n1725), .A3(n1625), .A4(n1626), .ZN(n1949) );
  INV_X4 U2203 ( .A(n1731), .ZN(n1626) );
  INV_X4 U2205 ( .A(n1954), .ZN(n1625) );
  INV_X4 U2207 ( .A(n1636), .ZN(n1725) );
  INV_X4 U2209 ( .A(n1957), .ZN(n1956) );
  NAND2_X2 U2213 ( .A1(n1962), .A2(n1963), .ZN(n1952) );
  INV_X4 U2214 ( .A(n1964), .ZN(n1961) );
  INV_X4 U2219 ( .A(n1968), .ZN(n1960) );
  INV_X4 U2220 ( .A(n1635), .ZN(n1800) );
  NAND2_X2 U2225 ( .A1(n1972), .A2(n1963), .ZN(n1953) );
  OR3_X2 U2226 ( .A1(n1973), .A2(n1939), .A3(n1681), .ZN(n1972) );
  AOI22_X2 U2228 ( .A1(n4822), .A2(n1976), .B1(n1977), .B2(n1978), .ZN(n1975)
         );
  NAND2_X2 U2231 ( .A1(n1981), .A2(n1982), .ZN(n1976) );
  NAND4_X2 U2232 ( .A1(u4_N6238), .A2(n6528), .A3(n1984), .A4(n4767), .ZN(
        n1982) );
  NAND4_X2 U2233 ( .A1(n1955), .A2(n1951), .A3(n1985), .A4(n1986), .ZN(n1984)
         );
  NOR4_X2 U2234 ( .A1(n1987), .A2(n1966), .A3(n1958), .A4(n1967), .ZN(n1986)
         );
  AND3_X2 U2235 ( .A1(n1988), .A2(n1989), .A3(n1990), .ZN(n1967) );
  AOI22_X2 U2237 ( .A1(u4_exp_out_pl1_4_), .A2(n1994), .B1(u4_exp_out_mi1[4]), 
        .B2(n1995), .ZN(n1989) );
  AOI22_X2 U2238 ( .A1(u4_exp_out_4_), .A2(n1996), .B1(n1997), .B2(n4399), 
        .ZN(n1988) );
  AND3_X2 U2239 ( .A1(n1998), .A2(n1999), .A3(n2000), .ZN(n1958) );
  AOI22_X2 U2241 ( .A1(u4_exp_out_pl1_2_), .A2(n1994), .B1(u4_exp_out_mi1[2]), 
        .B2(n1995), .ZN(n1999) );
  AOI22_X2 U2242 ( .A1(u4_exp_out_2_), .A2(n1996), .B1(n1997), .B2(exp_r[2]), 
        .ZN(n1998) );
  AND3_X2 U2243 ( .A1(n2001), .A2(n2002), .A3(n2003), .ZN(n1966) );
  AOI22_X2 U2245 ( .A1(u4_exp_out_pl1_3_), .A2(n1994), .B1(u4_exp_out_mi1[3]), 
        .B2(n1995), .ZN(n2002) );
  AOI22_X2 U2246 ( .A1(u4_exp_out_3_), .A2(n1996), .B1(n1997), .B2(exp_r[3]), 
        .ZN(n2001) );
  AOI22_X2 U2250 ( .A1(n1996), .A2(u4_exp_out_5_), .B1(u4_exp_out_pl1_5_), 
        .B2(n1994), .ZN(n2005) );
  AOI22_X2 U2251 ( .A1(n1991), .A2(u4_exp_next_mi_5_), .B1(u4_exp_fix_diva[5]), 
        .B2(n1993), .ZN(n2004) );
  AOI22_X2 U2254 ( .A1(n1996), .A2(u4_exp_out_6_), .B1(u4_exp_out_pl1_6_), 
        .B2(n1994), .ZN(n2008) );
  AOI22_X2 U2255 ( .A1(n1991), .A2(u4_exp_next_mi_6_), .B1(u4_exp_fix_diva[6]), 
        .B2(n1993), .ZN(n2007) );
  AOI22_X2 U2258 ( .A1(n1996), .A2(u4_exp_out_7_), .B1(u4_exp_out_pl1_7_), 
        .B2(n1994), .ZN(n2011) );
  AOI22_X2 U2259 ( .A1(n1991), .A2(u4_exp_next_mi_7_), .B1(u4_exp_fix_diva[7]), 
        .B2(n1993), .ZN(n2010) );
  AOI22_X2 U2263 ( .A1(u4_exp_out_pl1_8_), .A2(n1994), .B1(n1991), .B2(
        u4_exp_next_mi_8_), .ZN(n2014) );
  AOI22_X2 U2264 ( .A1(n2016), .A2(u4_exp_out_8_), .B1(u4_exp_fix_diva[8]), 
        .B2(n1993), .ZN(n2013) );
  AND3_X2 U2265 ( .A1(n2017), .A2(n2018), .A3(n2019), .ZN(n1965) );
  AOI22_X2 U2267 ( .A1(n1996), .A2(u4_exp_out_1_), .B1(u4_exp_out_pl1_1_), 
        .B2(n1994), .ZN(n2018) );
  NAND2_X2 U2268 ( .A1(n2020), .A2(n2021), .ZN(n1996) );
  AOI22_X2 U2270 ( .A1(n1991), .A2(u4_exp_next_mi_1_), .B1(u4_exp_fix_diva[1]), 
        .B2(n1993), .ZN(n2017) );
  AOI22_X2 U2273 ( .A1(u4_exp_out_pl1_9_), .A2(n1994), .B1(n1991), .B2(
        u4_exp_next_mi_9_), .ZN(n2025) );
  AOI22_X2 U2274 ( .A1(n2016), .A2(u4_exp_out_9_), .B1(u4_exp_fix_diva[9]), 
        .B2(n1993), .ZN(n2024) );
  AND3_X2 U2275 ( .A1(n2027), .A2(n2028), .A3(n2029), .ZN(n1951) );
  AOI22_X2 U2277 ( .A1(u4_exp_out_pl1_0_), .A2(n1994), .B1(n1991), .B2(
        u4_exp_next_mi_0_), .ZN(n2028) );
  AOI22_X2 U2278 ( .A1(n2016), .A2(u4_exp_out_0_), .B1(u4_exp_fix_diva[0]), 
        .B2(n1993), .ZN(n2027) );
  INV_X4 U2283 ( .A(n1682), .ZN(n1962) );
  OAI221_X2 U2284 ( .B1(n2033), .B2(n1974), .C1(exp_ovf_r_1_), .C2(n2034), .A(
        n2035), .ZN(n1682) );
  NAND2_X2 U2287 ( .A1(n4430), .A2(exp_ovf_r_1_), .ZN(n1685) );
  AND4_X2 U2289 ( .A1(sign), .A2(rmode_r3[1]), .A3(n4822), .A4(n2039), .ZN(
        n2038) );
  OAI221_X2 U2290 ( .B1(n2040), .B2(n1735), .C1(n2041), .C2(n6459), .A(n2042), 
        .ZN(n2039) );
  NAND4_X2 U2291 ( .A1(n1955), .A2(n4875), .A3(n2043), .A4(n2044), .ZN(n2042)
         );
  NAND4_X2 U2292 ( .A1(n2045), .A2(u4_exp_out_0_), .A3(u4_exp_out_8_), .A4(
        u4_exp_out_9_), .ZN(n2043) );
  AND3_X2 U2293 ( .A1(n2046), .A2(n2047), .A3(n2048), .ZN(n1955) );
  AOI22_X2 U2298 ( .A1(u4_exp_out_pl1_10_), .A2(n1994), .B1(n1991), .B2(
        u4_exp_next_mi_10_), .ZN(n2047) );
  INV_X4 U2302 ( .A(n1941), .ZN(n1944) );
  AOI22_X2 U2303 ( .A1(n2016), .A2(u4_exp_out_10_), .B1(u4_exp_fix_diva[10]), 
        .B2(n1993), .ZN(n2046) );
  INV_X4 U2307 ( .A(n2055), .ZN(n2020) );
  NAND2_X2 U2311 ( .A1(n1938), .A2(n2049), .ZN(n2056) );
  NAND4_X2 U2312 ( .A1(n6528), .A2(n2059), .A3(n2058), .A4(u4_fract_out_0_), 
        .ZN(n2049) );
  INV_X4 U2313 ( .A(n2060), .ZN(u4_fract_out_0_) );
  OAI22_X2 U2314 ( .A1(n2022), .A2(n2023), .B1(n1938), .B2(n4494), .ZN(n2054)
         );
  NAND2_X2 U2316 ( .A1(n1678), .A2(n1745), .ZN(n1938) );
  INV_X4 U2317 ( .A(n1946), .ZN(n2022) );
  NOR4_X2 U2322 ( .A1(n2061), .A2(n5046), .A3(n4430), .A4(n6386), .ZN(n2037)
         );
  NAND2_X2 U2324 ( .A1(n4483), .A2(n4427), .ZN(r482_B_0_) );
  NAND4_X2 U2326 ( .A1(n2045), .A2(u4_exp_out_mi1[0]), .A3(n4949), .A4(n205), 
        .ZN(n2063) );
  AND2_X2 U2328 ( .A1(n2064), .A2(u4_N6891), .ZN(n2045) );
  NAND4_X2 U2330 ( .A1(n4428), .A2(n4823), .A3(n2065), .A4(n2066), .ZN(n1732)
         );
  NOR4_X2 U2331 ( .A1(n2067), .A2(n4424), .A3(n4571), .A4(n4477), .ZN(n2066)
         );
  INV_X4 U2337 ( .A(n1684), .ZN(n1678) );
  AOI22_X2 U2342 ( .A1(u4_exp_f2i_1[115]), .A2(n2072), .B1(n2073), .B2(
        u4_sub_466_A_8_), .ZN(n2071) );
  OAI22_X2 U2343 ( .A1(n4874), .A2(n6521), .B1(n4873), .B2(n6164), .ZN(
        u4_sub_466_A_8_) );
  AOI221_X2 U2346 ( .B1(u4_div_exp2_8_), .B2(n2075), .C1(u4_exp_out1_mi1[8]), 
        .C2(n2076), .A(n5943), .ZN(n2069) );
  AOI22_X2 U2348 ( .A1(u4_div_exp1_8_), .A2(n2079), .B1(u4_div_exp3[8]), .B2(
        n2080), .ZN(n2078) );
  INV_X4 U2349 ( .A(u4_exp_out_9_), .ZN(n205) );
  AOI22_X2 U2351 ( .A1(u4_exp_f2i_1[116]), .A2(n2072), .B1(n2073), .B2(
        u4_sub_466_A_9_), .ZN(n2082) );
  AOI22_X2 U2353 ( .A1(fract_denorm[105]), .A2(u4_exp_in_pl1_9_), .B1(n4874), 
        .B2(u4_exp_next_mi_9_), .ZN(n2083) );
  AOI221_X2 U2354 ( .B1(u4_div_exp2_9_), .B2(n2075), .C1(u4_exp_out1_mi1[9]), 
        .C2(n2076), .A(n5942), .ZN(n2081) );
  AOI22_X2 U2356 ( .A1(u4_div_exp1_9_), .A2(n2079), .B1(u4_div_exp3[9]), .B2(
        n2080), .ZN(n2085) );
  INV_X4 U2357 ( .A(u4_exp_out_10_), .ZN(u4_N6891) );
  AOI22_X2 U2359 ( .A1(u4_exp_f2i_1[117]), .A2(n2072), .B1(n2073), .B2(
        u4_sub_466_A_10_), .ZN(n2086) );
  AOI22_X2 U2361 ( .A1(fract_denorm[105]), .A2(u4_exp_in_pl1_10_), .B1(n4874), 
        .B2(u4_exp_next_mi_10_), .ZN(n2087) );
  AND2_X2 U2363 ( .A1(n2089), .A2(n2090), .ZN(n1715) );
  AOI22_X2 U2364 ( .A1(u4_div_exp2_10_), .A2(n2075), .B1(u4_div_exp3[10]), 
        .B2(n2080), .ZN(n2090) );
  AOI22_X2 U2365 ( .A1(u4_div_exp1_10_), .A2(n2079), .B1(u4_exp_out1_mi1[10]), 
        .B2(n2076), .ZN(n2089) );
  NAND2_X2 U2366 ( .A1(n2091), .A2(n2092), .ZN(u4_exp_out_0_) );
  AOI221_X2 U2367 ( .B1(u4_exp_f2i_1[107]), .B2(n2072), .C1(n2093), .C2(
        fract_denorm[104]), .A(n2094), .ZN(n2092) );
  AOI22_X2 U2369 ( .A1(u4_div_exp2_0_), .A2(n2075), .B1(u4_exp_out1_mi1[0]), 
        .B2(n2076), .ZN(n2096) );
  AOI22_X2 U2370 ( .A1(u4_div_exp1_0_), .A2(n2079), .B1(u4_div_exp3[0]), .B2(
        n2080), .ZN(n2095) );
  AOI22_X2 U2372 ( .A1(n2073), .A2(u4_sub_466_A_0_), .B1(u4_fi_ldz_2a_0_), 
        .B2(n2088), .ZN(n2091) );
  OAI22_X2 U2373 ( .A1(n4874), .A2(n4823), .B1(n4873), .B2(n6170), .ZN(
        u4_sub_466_A_0_) );
  AND4_X2 U2376 ( .A1(u4_exp_out_2_), .A2(u4_exp_out_3_), .A3(u4_exp_out_1_), 
        .A4(n2099), .ZN(n2064) );
  NOR4_X2 U2377 ( .A1(n216), .A2(n4945), .A3(n222), .A4(n225), .ZN(n2099) );
  INV_X4 U2378 ( .A(u4_exp_out_4_), .ZN(n225) );
  NAND2_X2 U2379 ( .A1(n2100), .A2(n2101), .ZN(u4_exp_out_4_) );
  AOI221_X2 U2380 ( .B1(u4_exp_f2i_1[111]), .B2(n2072), .C1(n4822), .C2(n1722), 
        .A(n2102), .ZN(n2101) );
  NAND2_X2 U2381 ( .A1(n2103), .A2(n2104), .ZN(n1722) );
  AOI22_X2 U2382 ( .A1(u4_div_exp2_4_), .A2(n2075), .B1(u4_exp_out1_mi1[4]), 
        .B2(n2076), .ZN(n2104) );
  AOI22_X2 U2383 ( .A1(u4_div_exp1_4_), .A2(n2079), .B1(u4_div_exp3[4]), .B2(
        n2080), .ZN(n2103) );
  AOI22_X2 U2384 ( .A1(n2073), .A2(u4_sub_466_A_4_), .B1(u4_N6134), .B2(n2088), 
        .ZN(n2100) );
  OAI22_X2 U2385 ( .A1(n4874), .A2(n6523), .B1(n4873), .B2(n6166), .ZN(
        u4_sub_466_A_4_) );
  INV_X4 U2388 ( .A(u4_exp_out_5_), .ZN(n222) );
  NAND2_X2 U2389 ( .A1(n2106), .A2(n2107), .ZN(u4_exp_out_5_) );
  AOI22_X2 U2390 ( .A1(n4822), .A2(n1719), .B1(u4_exp_f2i_1[112]), .B2(n2072), 
        .ZN(n2107) );
  NAND2_X2 U2391 ( .A1(n2108), .A2(n2109), .ZN(n1719) );
  AOI22_X2 U2392 ( .A1(u4_div_exp2_5_), .A2(n2075), .B1(u4_div_exp3[5]), .B2(
        n2080), .ZN(n2109) );
  AOI22_X2 U2393 ( .A1(u4_div_exp1_5_), .A2(n2079), .B1(u4_exp_out1_mi1[5]), 
        .B2(n2076), .ZN(n2108) );
  AOI22_X2 U2394 ( .A1(n2073), .A2(u4_sub_466_A_5_), .B1(u4_N6135), .B2(n2088), 
        .ZN(n2106) );
  AOI22_X2 U2396 ( .A1(fract_denorm[105]), .A2(u4_exp_in_pl1_5_), .B1(n4874), 
        .B2(u4_exp_next_mi_5_), .ZN(n2110) );
  NAND2_X2 U2398 ( .A1(n2111), .A2(n2112), .ZN(u4_exp_out_6_) );
  AOI22_X2 U2399 ( .A1(n4822), .A2(n1720), .B1(u4_exp_f2i_1[113]), .B2(n2072), 
        .ZN(n2112) );
  NAND2_X2 U2400 ( .A1(n2113), .A2(n2114), .ZN(n1720) );
  AOI22_X2 U2401 ( .A1(u4_div_exp2_6_), .A2(n2075), .B1(u4_div_exp3[6]), .B2(
        n2080), .ZN(n2114) );
  AOI22_X2 U2402 ( .A1(u4_div_exp1_6_), .A2(n2079), .B1(u4_exp_out1_mi1[6]), 
        .B2(n2076), .ZN(n2113) );
  AOI22_X2 U2403 ( .A1(n2073), .A2(u4_sub_466_A_6_), .B1(u4_N6136), .B2(n2088), 
        .ZN(n2111) );
  AOI22_X2 U2405 ( .A1(fract_denorm[105]), .A2(u4_exp_in_pl1_6_), .B1(n4874), 
        .B2(u4_exp_next_mi_6_), .ZN(n2115) );
  INV_X4 U2406 ( .A(u4_exp_out_7_), .ZN(n216) );
  NAND2_X2 U2407 ( .A1(n2116), .A2(n2117), .ZN(u4_exp_out_7_) );
  AOI221_X2 U2408 ( .B1(u4_exp_f2i_1[114]), .B2(n2072), .C1(n4822), .C2(n1721), 
        .A(n2102), .ZN(n2117) );
  NAND2_X2 U2409 ( .A1(n2118), .A2(n2119), .ZN(n1721) );
  AOI22_X2 U2410 ( .A1(u4_div_exp2_7_), .A2(n2075), .B1(u4_exp_out1_mi1[7]), 
        .B2(n2076), .ZN(n2119) );
  AOI22_X2 U2411 ( .A1(u4_div_exp1_7_), .A2(n2079), .B1(u4_div_exp3[7]), .B2(
        n2080), .ZN(n2118) );
  AOI22_X2 U2412 ( .A1(n2073), .A2(u4_sub_466_A_7_), .B1(u4_N6137), .B2(n2088), 
        .ZN(n2116) );
  OAI22_X2 U2413 ( .A1(n4874), .A2(n6522), .B1(fract_denorm[105]), .B2(n6165), 
        .ZN(u4_sub_466_A_7_) );
  OAI211_X2 U2416 ( .C1(n5944), .C2(n4821), .A(n2122), .B(n2123), .ZN(
        u4_exp_out_1_) );
  AOI221_X2 U2417 ( .B1(u4_exp_f2i_1[108]), .B2(n2072), .C1(n2124), .C2(n6161), 
        .A(n2102), .ZN(n2123) );
  NOR2_X4 U2418 ( .A1(n4874), .A2(n2097), .ZN(n2124) );
  AOI22_X2 U2419 ( .A1(n2073), .A2(u4_exp_out1_1_), .B1(u4_N6131), .B2(n2088), 
        .ZN(n2122) );
  OAI22_X2 U2420 ( .A1(n4874), .A2(n6526), .B1(n4873), .B2(n6169), .ZN(
        u4_exp_out1_1_) );
  NAND2_X2 U2424 ( .A1(n2126), .A2(n2127), .ZN(n1716) );
  AOI22_X2 U2425 ( .A1(u4_div_exp2_1_), .A2(n2075), .B1(u4_div_exp3[1]), .B2(
        n2080), .ZN(n2127) );
  AOI22_X2 U2426 ( .A1(u4_div_exp1_1_), .A2(n2079), .B1(u4_exp_out1_mi1[1]), 
        .B2(n2076), .ZN(n2126) );
  NAND2_X2 U2427 ( .A1(n2128), .A2(n2129), .ZN(u4_exp_out_3_) );
  AOI221_X2 U2428 ( .B1(u4_exp_f2i_1[110]), .B2(n2072), .C1(n4822), .C2(n1718), 
        .A(n2102), .ZN(n2129) );
  NAND2_X2 U2429 ( .A1(n2130), .A2(n2131), .ZN(n1718) );
  AOI22_X2 U2430 ( .A1(u4_div_exp2_3_), .A2(n2075), .B1(u4_div_exp3[3]), .B2(
        n2080), .ZN(n2131) );
  AOI22_X2 U2431 ( .A1(u4_div_exp1_3_), .A2(n2079), .B1(u4_exp_out1_mi1[3]), 
        .B2(n2076), .ZN(n2130) );
  AOI22_X2 U2432 ( .A1(n2073), .A2(u4_sub_466_A_3_), .B1(u4_N6133), .B2(n2088), 
        .ZN(n2128) );
  OAI22_X2 U2433 ( .A1(n4874), .A2(n6524), .B1(fract_denorm[105]), .B2(n6167), 
        .ZN(u4_sub_466_A_3_) );
  NAND2_X2 U2436 ( .A1(n2133), .A2(n2134), .ZN(u4_exp_out_2_) );
  AOI221_X2 U2437 ( .B1(u4_exp_f2i_1[109]), .B2(n2072), .C1(n4822), .C2(n1717), 
        .A(n2102), .ZN(n2134) );
  NAND2_X2 U2439 ( .A1(n2135), .A2(n2136), .ZN(n1717) );
  AOI22_X2 U2440 ( .A1(u4_div_exp2_2_), .A2(n2075), .B1(u4_div_exp3[2]), .B2(
        n2080), .ZN(n2136) );
  AOI22_X2 U2442 ( .A1(u4_div_exp1_2_), .A2(n2079), .B1(u4_exp_out1_mi1[2]), 
        .B2(n2076), .ZN(n2135) );
  AOI22_X2 U2449 ( .A1(n4574), .A2(u4_N5831), .B1(u4_N5830), .B2(n2138), .ZN(
        n2032) );
  AOI22_X2 U2450 ( .A1(n2073), .A2(u4_sub_466_A_2_), .B1(u4_N6132), .B2(n2088), 
        .ZN(n2133) );
  OAI22_X2 U2452 ( .A1(n4874), .A2(n6525), .B1(fract_denorm[105]), .B2(n6168), 
        .ZN(u4_sub_466_A_2_) );
  OAI211_X2 U2457 ( .C1(n6162), .C2(n4819), .A(n2142), .B(n2143), .ZN(n2097)
         );
  INV_X4 U2461 ( .A(n2050), .ZN(n2051) );
  NAND2_X2 U2463 ( .A1(rmode_r3[1]), .A2(n1946), .ZN(n1942) );
  OAI211_X2 U2465 ( .C1(n2147), .C2(n1696), .A(n4483), .B(n6390), .ZN(n2146)
         );
  NAND2_X2 U2466 ( .A1(n2148), .A2(n2149), .ZN(n1696) );
  NOR4_X2 U2468 ( .A1(n2152), .A2(n2153), .A3(n2154), .A4(n2155), .ZN(n2151)
         );
  OR4_X2 U2469 ( .A1(fract_denorm[29]), .A2(fract_denorm[2]), .A3(
        fract_denorm[30]), .A4(fract_denorm[31]), .ZN(n2155) );
  NAND4_X2 U2470 ( .A1(n6442), .A2(n6443), .A3(n2156), .A4(n6444), .ZN(n2154)
         );
  NAND4_X2 U2474 ( .A1(n6449), .A2(n6453), .A3(n6462), .A4(n6463), .ZN(n2153)
         );
  NAND4_X2 U2475 ( .A1(n6465), .A2(n6467), .A3(n2162), .A4(n6410), .ZN(n2152)
         );
  NOR4_X2 U2478 ( .A1(n2163), .A2(n2164), .A3(n2165), .A4(n2166), .ZN(n2150)
         );
  NAND4_X2 U2479 ( .A1(n478), .A2(n505), .A3(n341), .A4(n328), .ZN(n2166) );
  NAND4_X2 U2480 ( .A1(n6425), .A2(n2168), .A3(n330), .A4(n334), .ZN(n2165) );
  NAND4_X2 U2481 ( .A1(n393), .A2(n544), .A3(n367), .A4(n369), .ZN(n2164) );
  NAND4_X2 U2482 ( .A1(n6430), .A2(n6437), .A3(n6407), .A4(n2170), .ZN(n2163)
         );
  AOI22_X2 U2485 ( .A1(n2171), .A2(u4_N6893), .B1(n2172), .B2(n1978), .ZN(
        n2145) );
  OAI221_X2 U2486 ( .B1(n1749), .B2(n2173), .C1(n6402), .C2(n4821), .A(n2174), 
        .ZN(n2172) );
  OAI211_X2 U2488 ( .C1(n4822), .C2(n4767), .A(n1743), .B(n1749), .ZN(n2175)
         );
  NAND2_X2 U2489 ( .A1(n2176), .A2(n2177), .ZN(n1743) );
  NOR4_X2 U2490 ( .A1(n2178), .A2(n2179), .A3(n2180), .A4(n2181), .ZN(n2177)
         );
  NAND4_X2 U2491 ( .A1(n1871), .A2(n1869), .A3(n1873), .A4(n2182), .ZN(n2181)
         );
  INV_X4 U2493 ( .A(n2183), .ZN(u4_fract_out_37_) );
  AOI22_X2 U2494 ( .A1(u4_N6099), .A2(n2184), .B1(u4_N5991), .B2(n4788), .ZN(
        n2183) );
  INV_X4 U2495 ( .A(n2186), .ZN(u4_fract_out_38_) );
  AOI22_X2 U2496 ( .A1(u4_N6100), .A2(n4790), .B1(u4_N5992), .B2(n4788), .ZN(
        n2186) );
  INV_X4 U2497 ( .A(n2187), .ZN(u4_fract_out_36_) );
  AOI22_X2 U2498 ( .A1(u4_N6098), .A2(n4790), .B1(u4_N5990), .B2(n4788), .ZN(
        n2187) );
  AOI22_X2 U2499 ( .A1(u4_N6095), .A2(n4790), .B1(u4_N5987), .B2(n4788), .ZN(
        n1873) );
  AOI22_X2 U2500 ( .A1(u4_N6097), .A2(n4790), .B1(u4_N5989), .B2(n4788), .ZN(
        n1869) );
  AOI22_X2 U2501 ( .A1(u4_N6096), .A2(n4790), .B1(u4_N5988), .B2(n4788), .ZN(
        n1871) );
  NAND4_X2 U2502 ( .A1(n1916), .A2(n1862), .A3(n1864), .A4(n2188), .ZN(n2180)
         );
  NOR4_X2 U2503 ( .A1(u4_fract_out_44_), .A2(u4_fract_out_43_), .A3(
        u4_fract_out_42_), .A4(u4_fract_out_41_), .ZN(n2188) );
  INV_X4 U2504 ( .A(n2189), .ZN(u4_fract_out_41_) );
  AOI22_X2 U2505 ( .A1(u4_N6103), .A2(n4790), .B1(u4_N5995), .B2(n4788), .ZN(
        n2189) );
  INV_X4 U2506 ( .A(n2190), .ZN(u4_fract_out_42_) );
  AOI22_X2 U2507 ( .A1(u4_N6104), .A2(n4790), .B1(u4_N5996), .B2(n4788), .ZN(
        n2190) );
  INV_X4 U2508 ( .A(n2191), .ZN(u4_fract_out_43_) );
  AOI22_X2 U2509 ( .A1(u4_N6105), .A2(n4790), .B1(u4_N5997), .B2(n4788), .ZN(
        n2191) );
  INV_X4 U2510 ( .A(n2192), .ZN(u4_fract_out_44_) );
  AOI22_X2 U2511 ( .A1(u4_N6106), .A2(n4790), .B1(u4_N5998), .B2(n4788), .ZN(
        n2192) );
  AOI22_X2 U2512 ( .A1(u4_N6101), .A2(n4790), .B1(u4_N5993), .B2(n4788), .ZN(
        n1864) );
  AOI22_X2 U2513 ( .A1(u4_N6102), .A2(n4791), .B1(u4_N5994), .B2(n4788), .ZN(
        n1862) );
  AOI22_X2 U2514 ( .A1(u4_N6065), .A2(n4791), .B1(u4_N5957), .B2(n4788), .ZN(
        n1916) );
  NAND4_X2 U2515 ( .A1(n1854), .A2(n1852), .A3(n1856), .A4(n2193), .ZN(n2179)
         );
  INV_X4 U2517 ( .A(n2194), .ZN(u4_fract_out_49_) );
  AOI22_X2 U2518 ( .A1(u4_N6111), .A2(n4791), .B1(u4_N6003), .B2(n4788), .ZN(
        n2194) );
  INV_X4 U2519 ( .A(n2195), .ZN(u4_fract_out_4_) );
  AOI22_X2 U2520 ( .A1(u4_N6066), .A2(n4791), .B1(u4_N5958), .B2(n4788), .ZN(
        n2195) );
  INV_X4 U2521 ( .A(n2196), .ZN(u4_fract_out_48_) );
  AOI22_X2 U2522 ( .A1(u4_N6110), .A2(n4791), .B1(u4_N6002), .B2(n4788), .ZN(
        n2196) );
  AOI22_X2 U2523 ( .A1(u4_N6107), .A2(n4791), .B1(u4_N5999), .B2(n4788), .ZN(
        n1856) );
  AOI22_X2 U2524 ( .A1(u4_N6109), .A2(n4791), .B1(u4_N6001), .B2(n4788), .ZN(
        n1852) );
  AOI22_X2 U2525 ( .A1(u4_N6108), .A2(n4791), .B1(u4_N6000), .B2(n4788), .ZN(
        n1854) );
  NAND4_X2 U2526 ( .A1(n1846), .A2(n1913), .A3(n1848), .A4(n2197), .ZN(n2178)
         );
  NOR4_X2 U2527 ( .A1(u4_fract_out_9_), .A2(u4_fract_out_8_), .A3(
        u4_fract_out_7_), .A4(u4_fract_out_6_), .ZN(n2197) );
  INV_X4 U2528 ( .A(n2198), .ZN(u4_fract_out_6_) );
  AOI22_X2 U2529 ( .A1(u4_N6068), .A2(n4791), .B1(u4_N5960), .B2(n4788), .ZN(
        n2198) );
  INV_X4 U2530 ( .A(n2199), .ZN(u4_fract_out_7_) );
  AOI22_X2 U2531 ( .A1(u4_N6069), .A2(n4791), .B1(u4_N5961), .B2(n4788), .ZN(
        n2199) );
  INV_X4 U2532 ( .A(n2200), .ZN(u4_fract_out_8_) );
  AOI22_X2 U2533 ( .A1(u4_N6070), .A2(n4791), .B1(u4_N5962), .B2(n4788), .ZN(
        n2200) );
  INV_X4 U2534 ( .A(n2201), .ZN(u4_fract_out_9_) );
  AOI22_X2 U2535 ( .A1(u4_N6071), .A2(n4790), .B1(u4_N5963), .B2(n4788), .ZN(
        n2201) );
  AOI22_X2 U2536 ( .A1(u4_N6112), .A2(n4790), .B1(u4_N6004), .B2(n4788), .ZN(
        n1848) );
  AOI22_X2 U2537 ( .A1(u4_N6067), .A2(n4790), .B1(u4_N5959), .B2(n4788), .ZN(
        n1913) );
  AOI22_X2 U2538 ( .A1(u4_N6113), .A2(n4790), .B1(u4_N6005), .B2(n4788), .ZN(
        n1846) );
  NOR4_X2 U2539 ( .A1(n2202), .A2(n2203), .A3(n2204), .A4(n2205), .ZN(n2176)
         );
  NAND4_X2 U2540 ( .A1(n1907), .A2(n1905), .A3(n2060), .A4(n2206), .ZN(n2205)
         );
  INV_X4 U2542 ( .A(n2207), .ZN(u4_fract_out_13_) );
  AOI22_X2 U2543 ( .A1(u4_N6075), .A2(n4790), .B1(u4_N5967), .B2(n4788), .ZN(
        n2207) );
  INV_X4 U2544 ( .A(n2208), .ZN(u4_fract_out_14_) );
  AOI22_X2 U2545 ( .A1(u4_N6076), .A2(n4790), .B1(u4_N5968), .B2(n4788), .ZN(
        n2208) );
  INV_X4 U2546 ( .A(n2209), .ZN(u4_fract_out_12_) );
  AOI22_X2 U2547 ( .A1(u4_N6074), .A2(n4790), .B1(u4_N5966), .B2(n4788), .ZN(
        n2209) );
  AOI22_X2 U2548 ( .A1(u4_N5954), .A2(n4789), .B1(u4_N6062), .B2(n2184), .ZN(
        n2060) );
  AOI22_X2 U2549 ( .A1(u4_N6073), .A2(n4790), .B1(u4_N5965), .B2(n4788), .ZN(
        n1905) );
  AOI22_X2 U2550 ( .A1(u4_N6072), .A2(n4790), .B1(u4_N5964), .B2(n4788), .ZN(
        n1907) );
  NAND4_X2 U2551 ( .A1(n1898), .A2(n1896), .A3(n1900), .A4(n2210), .ZN(n2204)
         );
  NOR4_X2 U2552 ( .A1(u4_fract_out_20_), .A2(u4_fract_out_1_), .A3(
        u4_fract_out_19_), .A4(u4_fract_out_18_), .ZN(n2210) );
  INV_X4 U2553 ( .A(n2211), .ZN(u4_fract_out_18_) );
  AOI22_X2 U2554 ( .A1(u4_N6080), .A2(n4790), .B1(u4_N5972), .B2(n4788), .ZN(
        n2211) );
  INV_X4 U2555 ( .A(n2212), .ZN(u4_fract_out_19_) );
  AOI22_X2 U2556 ( .A1(u4_N6081), .A2(n4790), .B1(u4_N5973), .B2(n4789), .ZN(
        n2212) );
  INV_X4 U2557 ( .A(n2213), .ZN(u4_fract_out_1_) );
  AOI22_X2 U2558 ( .A1(u4_N6063), .A2(n4791), .B1(u4_N5955), .B2(n4789), .ZN(
        n2213) );
  INV_X4 U2559 ( .A(n2214), .ZN(u4_fract_out_20_) );
  AOI22_X2 U2560 ( .A1(u4_N6082), .A2(n4790), .B1(u4_N5974), .B2(n4789), .ZN(
        n2214) );
  AOI22_X2 U2561 ( .A1(u4_N6077), .A2(n4790), .B1(u4_N5969), .B2(n4789), .ZN(
        n1900) );
  AOI22_X2 U2562 ( .A1(u4_N6079), .A2(n4790), .B1(u4_N5971), .B2(n4789), .ZN(
        n1896) );
  AOI22_X2 U2563 ( .A1(u4_N6078), .A2(n4790), .B1(u4_N5970), .B2(n4789), .ZN(
        n1898) );
  NAND4_X2 U2564 ( .A1(n1889), .A2(n1887), .A3(n1891), .A4(n2215), .ZN(n2203)
         );
  INV_X4 U2566 ( .A(n2216), .ZN(u4_fract_out_25_) );
  AOI22_X2 U2567 ( .A1(u4_N6087), .A2(n4790), .B1(u4_N5979), .B2(n4789), .ZN(
        n2216) );
  INV_X4 U2568 ( .A(n2217), .ZN(u4_fract_out_26_) );
  AOI22_X2 U2569 ( .A1(u4_N6088), .A2(n4790), .B1(u4_N5980), .B2(n4789), .ZN(
        n2217) );
  INV_X4 U2570 ( .A(n2218), .ZN(u4_fract_out_24_) );
  AOI22_X2 U2571 ( .A1(u4_N6086), .A2(n4790), .B1(u4_N5978), .B2(n4789), .ZN(
        n2218) );
  AOI22_X2 U2572 ( .A1(u4_N6083), .A2(n4790), .B1(u4_N5975), .B2(n4789), .ZN(
        n1891) );
  AOI22_X2 U2573 ( .A1(u4_N6085), .A2(n4790), .B1(u4_N5977), .B2(n4789), .ZN(
        n1887) );
  AOI22_X2 U2574 ( .A1(u4_N6084), .A2(n4790), .B1(u4_N5976), .B2(n4789), .ZN(
        n1889) );
  NAND4_X2 U2575 ( .A1(n1880), .A2(n1878), .A3(n1882), .A4(n2219), .ZN(n2202)
         );
  NOR4_X2 U2576 ( .A1(u4_fract_out_32_), .A2(u4_fract_out_31_), .A3(
        u4_fract_out_30_), .A4(u4_fract_out_2_), .ZN(n2219) );
  INV_X4 U2577 ( .A(n2220), .ZN(u4_fract_out_2_) );
  AOI22_X2 U2578 ( .A1(u4_N6064), .A2(n4790), .B1(u4_N5956), .B2(n4789), .ZN(
        n2220) );
  INV_X4 U2579 ( .A(n2221), .ZN(u4_fract_out_30_) );
  AOI22_X2 U2580 ( .A1(u4_N6092), .A2(n2184), .B1(u4_N5984), .B2(n4789), .ZN(
        n2221) );
  INV_X4 U2581 ( .A(n2222), .ZN(u4_fract_out_31_) );
  AOI22_X2 U2582 ( .A1(u4_N6093), .A2(n2184), .B1(u4_N5985), .B2(n4789), .ZN(
        n2222) );
  INV_X4 U2583 ( .A(n2223), .ZN(u4_fract_out_32_) );
  AOI22_X2 U2584 ( .A1(u4_N6094), .A2(n2184), .B1(u4_N5986), .B2(n4789), .ZN(
        n2223) );
  AOI22_X2 U2585 ( .A1(u4_N6089), .A2(n4791), .B1(u4_N5981), .B2(n4789), .ZN(
        n1882) );
  AOI22_X2 U2586 ( .A1(u4_N6091), .A2(n2184), .B1(u4_N5983), .B2(n4789), .ZN(
        n1878) );
  AOI22_X2 U2587 ( .A1(u4_N6090), .A2(n2184), .B1(u4_N5982), .B2(n4789), .ZN(
        n1880) );
  NAND2_X2 U2589 ( .A1(n2224), .A2(n2225), .ZN(n1705) );
  NOR4_X2 U2590 ( .A1(n2226), .A2(n2227), .A3(n2228), .A4(n2229), .ZN(n2225)
         );
  NAND4_X2 U2591 ( .A1(n2230), .A2(n2231), .A3(n2232), .A4(n2233), .ZN(n2229)
         );
  NOR4_X2 U2592 ( .A1(remainder[62]), .A2(remainder[61]), .A3(remainder[60]), 
        .A4(remainder[5]), .ZN(n2233) );
  NAND4_X2 U2596 ( .A1(n2234), .A2(n2235), .A3(n2236), .A4(n2237), .ZN(n2228)
         );
  NOR4_X2 U2597 ( .A1(remainder[75]), .A2(remainder[74]), .A3(remainder[73]), 
        .A4(remainder[72]), .ZN(n2237) );
  NOR4_X2 U2599 ( .A1(remainder[69]), .A2(remainder[68]), .A3(remainder[67]), 
        .A4(remainder[66]), .ZN(n2235) );
  NAND4_X2 U2601 ( .A1(n2238), .A2(n2239), .A3(n2240), .A4(n2241), .ZN(n2227)
         );
  NOR4_X2 U2602 ( .A1(remainder[87]), .A2(remainder[86]), .A3(remainder[85]), 
        .A4(remainder[84]), .ZN(n2241) );
  NAND4_X2 U2606 ( .A1(n2242), .A2(n2243), .A3(n2244), .A4(n2245), .ZN(n2226)
         );
  NOR4_X2 U2607 ( .A1(remainder[9]), .A2(remainder[99]), .A3(remainder[98]), 
        .A4(remainder[97]), .ZN(n2245) );
  NOR4_X2 U2609 ( .A1(remainder[93]), .A2(remainder[92]), .A3(remainder[91]), 
        .A4(remainder[90]), .ZN(n2243) );
  NOR4_X2 U2611 ( .A1(n2246), .A2(n2247), .A3(n2248), .A4(n2249), .ZN(n2224)
         );
  NAND4_X2 U2612 ( .A1(n2250), .A2(n2251), .A3(n2252), .A4(n2253), .ZN(n2249)
         );
  NOR4_X2 U2613 ( .A1(remainder[13]), .A2(remainder[12]), .A3(remainder[11]), 
        .A4(remainder[10]), .ZN(n2253) );
  NAND4_X2 U2617 ( .A1(n2254), .A2(n2255), .A3(n2256), .A4(n2257), .ZN(n2248)
         );
  NOR4_X2 U2618 ( .A1(remainder[26]), .A2(remainder[25]), .A3(remainder[24]), 
        .A4(remainder[23]), .ZN(n2257) );
  NOR4_X2 U2620 ( .A1(remainder[1]), .A2(remainder[19]), .A3(remainder[18]), 
        .A4(remainder[17]), .ZN(n2255) );
  NAND4_X2 U2622 ( .A1(n2258), .A2(n2259), .A3(n2260), .A4(n2261), .ZN(n2247)
         );
  NOR4_X2 U2623 ( .A1(remainder[38]), .A2(remainder[37]), .A3(remainder[36]), 
        .A4(remainder[35]), .ZN(n2261) );
  NAND4_X2 U2627 ( .A1(n2262), .A2(n2263), .A3(n2264), .A4(n2265), .ZN(n2246)
         );
  NOR4_X2 U2628 ( .A1(remainder[50]), .A2(remainder[4]), .A3(remainder[49]), 
        .A4(remainder[48]), .ZN(n2265) );
  NOR4_X2 U2630 ( .A1(remainder[44]), .A2(remainder[43]), .A3(remainder[42]), 
        .A4(remainder[41]), .ZN(n2263) );
  AOI221_X2 U2632 ( .B1(n1737), .B2(n4579), .C1(n2266), .C2(n4401), .A(n4822), 
        .ZN(n2173) );
  NAND2_X2 U2633 ( .A1(n4430), .A2(n2044), .ZN(n2266) );
  NAND2_X2 U2634 ( .A1(n4875), .A2(n2267), .ZN(n2044) );
  AND3_X2 U2638 ( .A1(n401), .A2(n211), .A3(u4_N5837), .ZN(n2269) );
  AOI22_X2 U2641 ( .A1(n2270), .A2(n2184), .B1(n2271), .B2(n4789), .ZN(n2149)
         );
  OR4_X2 U2642 ( .A1(n2272), .A2(n2273), .A3(n2274), .A4(n2275), .ZN(n2271) );
  NAND4_X2 U2643 ( .A1(n2276), .A2(n2277), .A3(n2278), .A4(n2279), .ZN(n2275)
         );
  NOR4_X2 U2644 ( .A1(u4_N5912), .A2(u4_N5911), .A3(u4_N5910), .A4(u4_N5909), 
        .ZN(n2279) );
  NAND4_X2 U2648 ( .A1(n2280), .A2(n2281), .A3(n2282), .A4(n2283), .ZN(n2274)
         );
  NOR4_X2 U2649 ( .A1(u4_N5925), .A2(u4_N5924), .A3(u4_N5923), .A4(u4_N5922), 
        .ZN(n2283) );
  NAND4_X2 U2653 ( .A1(n2284), .A2(n2285), .A3(n2286), .A4(n2287), .ZN(n2273)
         );
  NOR4_X2 U2654 ( .A1(u4_N5938), .A2(u4_N5937), .A3(u4_N5936), .A4(u4_N5935), 
        .ZN(n2287) );
  NAND4_X2 U2658 ( .A1(n2288), .A2(n2289), .A3(n2290), .A4(n2291), .ZN(n2272)
         );
  NOR4_X2 U2659 ( .A1(u4_N5952), .A2(u4_N5951), .A3(u4_N5950), .A4(u4_N5949), 
        .ZN(n2291) );
  NOR3_X4 U2660 ( .A1(u4_N5946), .A2(u4_N5948), .A3(u4_N5947), .ZN(n2290) );
  NOR4_X2 U2661 ( .A1(u4_N5945), .A2(u4_N5944), .A3(u4_N5943), .A4(u4_N5942), 
        .ZN(n2289) );
  NOR3_X4 U2662 ( .A1(u4_N5939), .A2(u4_N5941), .A3(u4_N5940), .ZN(n2288) );
  OR4_X2 U2663 ( .A1(n2292), .A2(n2293), .A3(n2294), .A4(n2295), .ZN(n2270) );
  NAND4_X2 U2664 ( .A1(n2296), .A2(n2297), .A3(n2298), .A4(n2299), .ZN(n2295)
         );
  NOR4_X2 U2665 ( .A1(u4_N6020), .A2(u4_N6019), .A3(u4_N6018), .A4(u4_N6017), 
        .ZN(n2299) );
  NAND4_X2 U2669 ( .A1(n2300), .A2(n2301), .A3(n2302), .A4(n2303), .ZN(n2294)
         );
  NOR4_X2 U2670 ( .A1(u4_N6033), .A2(u4_N6032), .A3(u4_N6031), .A4(u4_N6030), 
        .ZN(n2303) );
  NAND4_X2 U2674 ( .A1(n2304), .A2(n2305), .A3(n2306), .A4(n2307), .ZN(n2293)
         );
  NOR4_X2 U2675 ( .A1(u4_N6046), .A2(u4_N6045), .A3(u4_N6044), .A4(u4_N6043), 
        .ZN(n2307) );
  NAND4_X2 U2679 ( .A1(n2308), .A2(n2309), .A3(n2310), .A4(n2311), .ZN(n2292)
         );
  NOR4_X2 U2680 ( .A1(u4_N6060), .A2(u4_N6059), .A3(u4_N6058), .A4(u4_N6057), 
        .ZN(n2311) );
  NOR4_X2 U2682 ( .A1(u4_N6053), .A2(u4_N6052), .A3(u4_N6051), .A4(u4_N6050), 
        .ZN(n2309) );
  AOI22_X2 U2684 ( .A1(u4_N6061), .A2(n4790), .B1(u4_N5953), .B2(n4788), .ZN(
        n2148) );
  AND4_X2 U2686 ( .A1(n2313), .A2(n2312), .A3(n2314), .A4(n2315), .ZN(n2184)
         );
  NAND2_X2 U2689 ( .A1(n294), .A2(n4822), .ZN(n288) );
  NOR3_X4 U2690 ( .A1(exp_ovf_r_1_), .A2(u4_N6440), .A3(n4767), .ZN(n294) );
  OR3_X2 U2692 ( .A1(u4_f2i_shft_9_), .A2(u4_f2i_shft_10_), .A3(n1755), .ZN(
        n2316) );
  OAI22_X2 U2693 ( .A1(n4574), .A2(n6529), .B1(n2138), .B2(n6376), .ZN(n1755)
         );
  NOR4_X2 U2695 ( .A1(n4427), .A2(n4483), .A3(n4574), .A4(n6403), .ZN(n2138)
         );
  NAND2_X2 U2701 ( .A1(n439), .A2(n6414), .ZN(n504) );
  NAND2_X2 U2704 ( .A1(n337), .A2(n341), .ZN(n296) );
  NAND2_X2 U2709 ( .A1(n335), .A2(n6425), .ZN(n329) );
  NAND4_X2 U2711 ( .A1(n6426), .A2(n6427), .A3(n6428), .A4(n6429), .ZN(n336)
         );
  NAND2_X2 U2717 ( .A1(n6436), .A2(n330), .ZN(n420) );
  NAND2_X2 U2722 ( .A1(n536), .A2(n6441), .ZN(n421) );
  NAND2_X2 U2729 ( .A1(u4_fi_ldz_6_), .A2(n6453), .ZN(n443) );
  NAND2_X2 U2734 ( .A1(n6461), .A2(n369), .ZN(n366) );
  NAND2_X2 U2737 ( .A1(n566), .A2(n6462), .ZN(n368) );
  AND4_X2 U2739 ( .A1(n401), .A2(n4874), .A3(n6463), .A4(n6465), .ZN(n566) );
  NAND2_X2 U2748 ( .A1(n6478), .A2(n309), .ZN(n376) );
  NAND2_X2 U2751 ( .A1(n6479), .A2(n307), .ZN(n310) );
  NAND2_X2 U2760 ( .A1(n6495), .A2(n350), .ZN(n312) );
  NAND2_X2 U2763 ( .A1(n6499), .A2(n348), .ZN(n351) );
  NOR4_X2 U2764 ( .A1(fract_denorm[80]), .A2(fract_denorm[81]), .A3(
        fract_denorm[82]), .A4(fract_denorm[83]), .ZN(n348) );
  NAND2_X2 U2768 ( .A1(n357), .A2(n6505), .ZN(n454) );
  NOR4_X2 U2770 ( .A1(n6509), .A2(fract_denorm[90]), .A3(fract_denorm[91]), 
        .A4(fract_denorm[92]), .ZN(n357) );
  NAND4_X2 U2777 ( .A1(n418), .A2(n6518), .A3(n6519), .A4(n6515), .ZN(n394) );
  OR2_X2 U2790 ( .A1(fract_denorm[60]), .A2(fract_denorm[59]), .ZN(n318) );
  AOI21_X4 U2812 ( .B1(n2327), .B2(n247), .A(u4_N6440), .ZN(n295) );
  NAND2_X2 U2813 ( .A1(n4579), .A2(n4767), .ZN(n2327) );
  OAI221_X2 U2815 ( .B1(n241), .B2(n6520), .C1(n1740), .C2(n4822), .A(n2328), 
        .ZN(n2312) );
  AND2_X2 U2817 ( .A1(n247), .A2(n246), .ZN(n242) );
  NAND2_X2 U2819 ( .A1(exp_ovf_r_1_), .A2(n4767), .ZN(n247) );
  NAND2_X2 U2823 ( .A1(n1708), .A2(n4821), .ZN(n241) );
  OR3_X2 U2826 ( .A1(n282), .A2(n6527), .A3(n281), .ZN(n2329) );
  NAND2_X2 U2827 ( .A1(n6384), .A2(n1925), .ZN(n281) );
  NAND2_X2 U2828 ( .A1(n4778), .A2(n4481), .ZN(n1925) );
  NAND2_X2 U2830 ( .A1(n6386), .A2(n1745), .ZN(n2268) );
  INV_X4 U2831 ( .A(n290), .ZN(n282) );
  NAND2_X2 U2832 ( .A1(u4_N6440), .A2(n1739), .ZN(n290) );
  NAND2_X2 U2833 ( .A1(n6386), .A2(n2330), .ZN(n1739) );
  INV_X4 U2835 ( .A(n289), .ZN(n279) );
  INV_X4 U2838 ( .A(u4_N6440), .ZN(n1701) );
  NAND2_X2 U2840 ( .A1(n6527), .A2(n4401), .ZN(n1708) );
  NAND2_X2 U2842 ( .A1(n2267), .A2(n4587), .ZN(n1735) );
  AND4_X2 U2844 ( .A1(n4477), .A2(n4571), .A3(n1710), .A4(n2333), .ZN(n2267)
         );
  NOR4_X2 U2845 ( .A1(n2334), .A2(exp_r[2]), .A3(n4399), .A4(exp_r[3]), .ZN(
        n2333) );
  NAND2_X2 U2846 ( .A1(n4400), .A2(n4588), .ZN(n2334) );
  INV_X4 U2852 ( .A(u4_fract_out_pl1_52_), .ZN(n2023) );
  NAND2_X2 U2855 ( .A1(u4_exp_in_pl1_11_), .A2(n4873), .ZN(n2335) );
  NAND2_X2 U2860 ( .A1(n6379), .A2(n4822), .ZN(n2033) );
  NAND2_X2 U2866 ( .A1(n4778), .A2(fpu_op_r3[0]), .ZN(n1745) );
  NAND2_X2 U2868 ( .A1(rmode_r3[0]), .A2(n4427), .ZN(n1671) );
  OAI221_X2 U2870 ( .B1(n4821), .B2(n4432), .C1(n6386), .C2(n4493), .A(n1920), 
        .ZN(n1947) );
  NAND2_X2 U2871 ( .A1(opb_00), .A2(n4820), .ZN(n1920) );
  XOR2_X2 U2875 ( .A(n2337), .B(n2338), .Z(N794) );
  NAND2_X2 U2876 ( .A1(rmode_r2[1]), .A2(rmode_r2[0]), .ZN(n2338) );
  OAI221_X2 U2877 ( .B1(n4484), .B2(n4568), .C1(n1138), .C2(n4766), .A(n2341), 
        .ZN(N791) );
  OAI221_X2 U2881 ( .B1(n4819), .B2(n4436), .C1(n4803), .C2(n4765), .A(n2344), 
        .ZN(N790) );
  OAI221_X2 U2885 ( .B1(n4819), .B2(n4513), .C1(n4806), .C2(n4764), .A(n2346), 
        .ZN(N789) );
  OAI221_X2 U2889 ( .B1(n4819), .B2(n4405), .C1(n4804), .C2(n4763), .A(n2348), 
        .ZN(N788) );
  OAI221_X2 U2893 ( .B1(n4819), .B2(n4561), .C1(n4803), .C2(n4762), .A(n2351), 
        .ZN(N787) );
  OAI221_X2 U2897 ( .B1(n4818), .B2(n4554), .C1(n1138), .C2(n4761), .A(n2354), 
        .ZN(N786) );
  OAI221_X2 U2901 ( .B1(n4818), .B2(n4412), .C1(n4804), .C2(n4760), .A(n2356), 
        .ZN(N785) );
  NAND2_X2 U2907 ( .A1(n4484), .A2(n4821), .ZN(n1978) );
  OAI221_X2 U2908 ( .B1(n4484), .B2(n4518), .C1(n4803), .C2(n4759), .A(n2359), 
        .ZN(N783) );
  OAI221_X2 U2912 ( .B1(n4484), .B2(n4441), .C1(n1138), .C2(n4758), .A(n2361), 
        .ZN(N782) );
  OAI221_X2 U2916 ( .B1(n4484), .B2(n4560), .C1(n4803), .C2(n4757), .A(n2364), 
        .ZN(N781) );
  OAI221_X2 U2920 ( .B1(n4484), .B2(n4553), .C1(n1138), .C2(n4756), .A(n2367), 
        .ZN(N780) );
  OAI221_X2 U2924 ( .B1(n4484), .B2(n4567), .C1(n4806), .C2(n4755), .A(n2370), 
        .ZN(N779) );
  OAI221_X2 U2928 ( .B1(n4484), .B2(n4389), .C1(n4804), .C2(n4754), .A(n2372), 
        .ZN(N778) );
  OAI221_X2 U2932 ( .B1(n4484), .B2(n4411), .C1(n4803), .C2(n4753), .A(n2374), 
        .ZN(N777) );
  OAI221_X2 U2936 ( .B1(n4484), .B2(n4517), .C1(n1138), .C2(n4752), .A(n2376), 
        .ZN(N776) );
  OAI221_X2 U2940 ( .B1(n4484), .B2(n4440), .C1(n4803), .C2(n4751), .A(n2378), 
        .ZN(N775) );
  OAI221_X2 U2944 ( .B1(n4484), .B2(n4552), .C1(n4803), .C2(n4750), .A(n2381), 
        .ZN(N774) );
  OAI221_X2 U2948 ( .B1(n4484), .B2(n4566), .C1(n4806), .C2(n4749), .A(n2384), 
        .ZN(N773) );
  OAI221_X2 U2952 ( .B1(n4484), .B2(n4388), .C1(n4806), .C2(n4748), .A(n2386), 
        .ZN(N772) );
  OAI221_X2 U2956 ( .B1(n4484), .B2(n4439), .C1(n4804), .C2(n4747), .A(n2388), 
        .ZN(N771) );
  OAI221_X2 U2960 ( .B1(n4484), .B2(n4516), .C1(n4804), .C2(n4746), .A(n2390), 
        .ZN(N770) );
  OAI221_X2 U2964 ( .B1(n4818), .B2(n4414), .C1(n4806), .C2(n4745), .A(n2392), 
        .ZN(N769) );
  OAI221_X2 U2968 ( .B1(n4818), .B2(n4559), .C1(n4804), .C2(n4744), .A(n2395), 
        .ZN(N768) );
  OAI221_X2 U2972 ( .B1(n4818), .B2(n4551), .C1(n4806), .C2(n4743), .A(n2398), 
        .ZN(N767) );
  OAI221_X2 U2976 ( .B1(n4818), .B2(n4565), .C1(n1138), .C2(n4742), .A(n2401), 
        .ZN(N766) );
  OAI221_X2 U2980 ( .B1(n4818), .B2(n4506), .C1(n4803), .C2(n4741), .A(n2403), 
        .ZN(N765) );
  OAI221_X2 U2984 ( .B1(n4818), .B2(n4385), .C1(n4804), .C2(n4740), .A(n2405), 
        .ZN(N764) );
  OAI221_X2 U2988 ( .B1(n4818), .B2(n4558), .C1(n4804), .C2(n4739), .A(n2408), 
        .ZN(N763) );
  OAI221_X2 U2992 ( .B1(n4818), .B2(n4550), .C1(n1138), .C2(n4738), .A(n2411), 
        .ZN(N762) );
  OAI221_X2 U2996 ( .B1(n4818), .B2(n4564), .C1(n4803), .C2(n4737), .A(n2414), 
        .ZN(N761) );
  OAI221_X2 U3000 ( .B1(n4818), .B2(n4391), .C1(n4803), .C2(n4736), .A(n2416), 
        .ZN(N760) );
  OAI221_X2 U3004 ( .B1(n4818), .B2(n4413), .C1(n4806), .C2(n4735), .A(n2418), 
        .ZN(N759) );
  OAI221_X2 U3008 ( .B1(n4818), .B2(n4520), .C1(n4806), .C2(n4734), .A(n2420), 
        .ZN(N758) );
  OAI221_X2 U3012 ( .B1(n4818), .B2(n4442), .C1(n4806), .C2(n4733), .A(n2422), 
        .ZN(N757) );
  OAI221_X2 U3016 ( .B1(n4818), .B2(n4557), .C1(n4806), .C2(n4732), .A(n2425), 
        .ZN(N756) );
  OAI221_X2 U3020 ( .B1(n4818), .B2(n4549), .C1(n4806), .C2(n4731), .A(n2428), 
        .ZN(N755) );
  OAI221_X2 U3024 ( .B1(n4818), .B2(n4434), .C1(n4806), .C2(n4730), .A(n2430), 
        .ZN(N754) );
  OAI221_X2 U3028 ( .B1(n4818), .B2(n4511), .C1(n4806), .C2(n4729), .A(n2432), 
        .ZN(N753) );
  OAI221_X2 U3032 ( .B1(n4818), .B2(n4404), .C1(n4806), .C2(n4728), .A(n2434), 
        .ZN(N752) );
  OAI221_X2 U3036 ( .B1(n4819), .B2(n4556), .C1(n4806), .C2(n4727), .A(n2437), 
        .ZN(N751) );
  OAI221_X2 U3040 ( .B1(n4818), .B2(n4548), .C1(n4806), .C2(n4726), .A(n2440), 
        .ZN(N750) );
  OAI221_X2 U3044 ( .B1(n4818), .B2(n4563), .C1(n4806), .C2(n4725), .A(n2443), 
        .ZN(N749) );
  OAI221_X2 U3048 ( .B1(n4818), .B2(n4378), .C1(n4804), .C2(n4724), .A(n2445), 
        .ZN(N748) );
  OAI221_X2 U3052 ( .B1(n4819), .B2(n4392), .C1(n4803), .C2(n4723), .A(n2447), 
        .ZN(N747) );
  OAI221_X2 U3056 ( .B1(n4819), .B2(n4519), .C1(n1138), .C2(n4722), .A(n2449), 
        .ZN(N746) );
  OAI221_X2 U3060 ( .B1(n4818), .B2(n4415), .C1(n4806), .C2(n4721), .A(n2451), 
        .ZN(N745) );
  OAI221_X2 U3064 ( .B1(n4818), .B2(n4547), .C1(n1138), .C2(n4720), .A(n2454), 
        .ZN(N744) );
  OAI221_X2 U3068 ( .B1(n4819), .B2(n4562), .C1(n4806), .C2(n4719), .A(n2457), 
        .ZN(N743) );
  OAI221_X2 U3072 ( .B1(n4818), .B2(n4387), .C1(n4804), .C2(n4718), .A(n2459), 
        .ZN(N742) );
  OAI221_X2 U3076 ( .B1(n4818), .B2(n4510), .C1(n4803), .C2(n4717), .A(n2461), 
        .ZN(N741) );
  OAI221_X2 U3080 ( .B1(n4818), .B2(n4403), .C1(n1138), .C2(n4716), .A(n2463), 
        .ZN(N740) );
  OAI221_X2 U3084 ( .B1(n4819), .B2(n4555), .C1(n4806), .C2(n4715), .A(n2466), 
        .ZN(N739) );
  OAI221_X2 U3088 ( .B1(n4819), .B2(n4689), .C1(n4804), .C2(n4546), .A(n2469), 
        .ZN(N738) );
  OAI221_X2 U3100 ( .B1(n4819), .B2(n4395), .C1(n4806), .C2(n4688), .A(n2476), 
        .ZN(N735) );
  OAI221_X2 U3105 ( .B1(n4818), .B2(n4515), .C1(n1138), .C2(n4687), .A(n2478), 
        .ZN(N734) );
  AOI22_X2 U3106 ( .A1(fract_out_q[0]), .A2(n4772), .B1(fract_i2f[49]), .B2(
        n4777), .ZN(n2478) );
  NAND2_X2 U3108 ( .A1(n4353), .A2(n4351), .ZN(n1664) );
  OAI221_X2 U3111 ( .B1(n4819), .B2(n4380), .C1(n4803), .C2(n4686), .A(n2481), 
        .ZN(N730) );
  NAND2_X2 U3112 ( .A1(fract_i2f[45]), .A2(n4775), .ZN(n2481) );
  OAI221_X2 U3115 ( .B1(n4818), .B2(n4394), .C1(n1138), .C2(n4685), .A(n2483), 
        .ZN(N729) );
  NAND2_X2 U3116 ( .A1(fract_i2f[44]), .A2(n4778), .ZN(n2483) );
  OAI221_X2 U3119 ( .B1(n4819), .B2(n4522), .C1(n4804), .C2(n4684), .A(n2485), 
        .ZN(N728) );
  NAND2_X2 U3120 ( .A1(fract_i2f[43]), .A2(n4778), .ZN(n2485) );
  OAI221_X2 U3123 ( .B1(n4819), .B2(n4444), .C1(n4806), .C2(n4683), .A(n2487), 
        .ZN(N727) );
  NAND2_X2 U3124 ( .A1(fract_i2f[42]), .A2(n4778), .ZN(n2487) );
  OAI221_X2 U3127 ( .B1(n4819), .B2(n4379), .C1(n1138), .C2(n4682), .A(n2489), 
        .ZN(N724) );
  NAND2_X2 U3128 ( .A1(fract_i2f[39]), .A2(n4778), .ZN(n2489) );
  OAI221_X2 U3131 ( .B1(n4819), .B2(n4393), .C1(n4803), .C2(n4681), .A(n2491), 
        .ZN(N723) );
  NAND2_X2 U3132 ( .A1(fract_i2f[38]), .A2(n4778), .ZN(n2491) );
  OAI221_X2 U3135 ( .B1(n4818), .B2(n4521), .C1(n4803), .C2(n4680), .A(n2493), 
        .ZN(N722) );
  NAND2_X2 U3136 ( .A1(fract_i2f[37]), .A2(n4778), .ZN(n2493) );
  OAI221_X2 U3139 ( .B1(n4818), .B2(n4443), .C1(n4804), .C2(n4679), .A(n2495), 
        .ZN(N721) );
  NAND2_X2 U3140 ( .A1(fract_i2f[36]), .A2(n4778), .ZN(n2495) );
  OAI221_X2 U3143 ( .B1(n4818), .B2(n4435), .C1(n4806), .C2(n4678), .A(n2497), 
        .ZN(N717) );
  NAND2_X2 U3144 ( .A1(fract_i2f[32]), .A2(n4778), .ZN(n2497) );
  OAI221_X2 U3147 ( .B1(n4819), .B2(n4512), .C1(n4803), .C2(n4677), .A(n2499), 
        .ZN(N716) );
  NAND2_X2 U3148 ( .A1(fract_i2f[31]), .A2(n4778), .ZN(n2499) );
  OAI221_X2 U3151 ( .B1(n4819), .B2(n4386), .C1(n1138), .C2(n4676), .A(n2501), 
        .ZN(N715) );
  NAND2_X2 U3152 ( .A1(fract_i2f[30]), .A2(n4778), .ZN(n2501) );
  OAI221_X2 U3155 ( .B1(n4819), .B2(n4381), .C1(n4804), .C2(n4675), .A(n2503), 
        .ZN(N712) );
  NAND2_X2 U3156 ( .A1(fract_i2f[27]), .A2(n4778), .ZN(n2503) );
  OAI221_X2 U3159 ( .B1(n4818), .B2(n4397), .C1(n4806), .C2(n4674), .A(n2505), 
        .ZN(N711) );
  NAND2_X2 U3160 ( .A1(fract_i2f[26]), .A2(n4778), .ZN(n2505) );
  OAI221_X2 U3163 ( .B1(n4818), .B2(n4523), .C1(n4803), .C2(n4673), .A(n2507), 
        .ZN(N710) );
  NAND2_X2 U3164 ( .A1(fract_i2f[25]), .A2(n4778), .ZN(n2507) );
  OAI221_X2 U3167 ( .B1(n4819), .B2(n4445), .C1(n1138), .C2(n4672), .A(n2509), 
        .ZN(N709) );
  NAND2_X2 U3168 ( .A1(fract_i2f[24]), .A2(n4778), .ZN(n2509) );
  OAI221_X2 U3171 ( .B1(n4819), .B2(n4507), .C1(n4804), .C2(n4671), .A(n2511), 
        .ZN(N705) );
  NAND2_X2 U3172 ( .A1(fract_i2f[20]), .A2(n4778), .ZN(n2511) );
  OAI221_X2 U3175 ( .B1(n4819), .B2(n4406), .C1(n4806), .C2(n4670), .A(n2513), 
        .ZN(N704) );
  NAND2_X2 U3176 ( .A1(fract_i2f[19]), .A2(n4778), .ZN(n2513) );
  OAI221_X2 U3179 ( .B1(n4819), .B2(n4514), .C1(n4803), .C2(n4669), .A(n2515), 
        .ZN(N700) );
  NAND2_X2 U3180 ( .A1(fract_i2f[15]), .A2(n4778), .ZN(n2515) );
  OAI221_X2 U3183 ( .B1(n4819), .B2(n4396), .C1(n1138), .C2(n4545), .A(n2517), 
        .ZN(N699) );
  NAND2_X2 U3184 ( .A1(fract_i2f[14]), .A2(n4777), .ZN(n2517) );
  OAI221_X2 U3187 ( .B1(n4819), .B2(n4447), .C1(n4804), .C2(n4544), .A(n2519), 
        .ZN(N698) );
  NAND2_X2 U3188 ( .A1(fract_i2f[13]), .A2(n4778), .ZN(n2519) );
  OAI221_X2 U3191 ( .B1(n4819), .B2(n4416), .C1(n1138), .C2(n4543), .A(n2521), 
        .ZN(N697) );
  NAND2_X2 U3192 ( .A1(fract_i2f[12]), .A2(n4778), .ZN(n2521) );
  OAI221_X2 U3195 ( .B1(n4819), .B2(n4390), .C1(n4804), .C2(n4542), .A(n2523), 
        .ZN(N694) );
  NAND2_X2 U3196 ( .A1(fract_i2f[9]), .A2(n4776), .ZN(n2523) );
  OAI221_X2 U3199 ( .B1(n4818), .B2(n4437), .C1(n1138), .C2(n4541), .A(n2525), 
        .ZN(N692) );
  NAND2_X2 U3200 ( .A1(fract_i2f[7]), .A2(n4778), .ZN(n2525) );
  OAI221_X2 U3203 ( .B1(n4819), .B2(n4446), .C1(n4804), .C2(n4540), .A(n2527), 
        .ZN(N689) );
  NAND2_X2 U3204 ( .A1(fract_i2f[4]), .A2(n4778), .ZN(n2527) );
  OAI221_X2 U3207 ( .B1(n4819), .B2(n4438), .C1(n1138), .C2(n4539), .A(n2529), 
        .ZN(N686) );
  NAND2_X2 U3208 ( .A1(fract_i2f[1]), .A2(n4778), .ZN(n2529) );
  NAND2_X2 U3210 ( .A1(fpu_op_r3[2]), .A2(n4353), .ZN(n2357) );
  NAND2_X2 U3213 ( .A1(opb_dn), .A2(n4822), .ZN(n1138) );
  OAI221_X2 U3220 ( .B1(n4768), .B2(n6025), .C1(n4629), .C2(n2532), .A(n4779), 
        .ZN(N667) );
  OAI221_X2 U3223 ( .B1(n4769), .B2(n6026), .C1(n4410), .C2(n4782), .A(n4779), 
        .ZN(N666) );
  OAI221_X2 U3226 ( .B1(n4768), .B2(n6027), .C1(n4409), .C2(n4782), .A(n4779), 
        .ZN(N665) );
  OAI221_X2 U3229 ( .B1(n4769), .B2(n6028), .C1(n4408), .C2(n4782), .A(n4779), 
        .ZN(N664) );
  OAI221_X2 U3232 ( .B1(n4768), .B2(n6029), .C1(n4407), .C2(n4782), .A(n4779), 
        .ZN(N663) );
  OAI221_X2 U3235 ( .B1(n4769), .B2(n6030), .C1(n4625), .C2(n4784), .A(n4779), 
        .ZN(N662) );
  OAI221_X2 U3238 ( .B1(n4768), .B2(n6031), .C1(n4622), .C2(n4784), .A(n4779), 
        .ZN(N661) );
  OAI221_X2 U3240 ( .B1(n4769), .B2(n6032), .C1(n4509), .C2(n4784), .A(n4779), 
        .ZN(N660) );
  OAI221_X2 U3242 ( .B1(n4768), .B2(n6033), .C1(n2532), .C2(n4419), .A(n4779), 
        .ZN(N659) );
  OAI221_X2 U3245 ( .B1(n4769), .B2(n6034), .C1(n2532), .C2(n4418), .A(n4779), 
        .ZN(N658) );
  OAI221_X2 U3248 ( .B1(n4768), .B2(n6035), .C1(n2532), .C2(n4417), .A(n4779), 
        .ZN(N657) );
  OAI221_X2 U3251 ( .B1(n4768), .B2(n6036), .C1(n2532), .C2(n4450), .A(n4779), 
        .ZN(N656) );
  OAI221_X2 U3254 ( .B1(n4768), .B2(n6037), .C1(n2532), .C2(n4449), .A(n4779), 
        .ZN(N655) );
  OAI221_X2 U3257 ( .B1(n4768), .B2(n6038), .C1(n2532), .C2(n4448), .A(n4779), 
        .ZN(N654) );
  OAI221_X2 U3260 ( .B1(n4768), .B2(n6039), .C1(n4665), .C2(n4784), .A(n2533), 
        .ZN(N653) );
  OAI221_X2 U3263 ( .B1(n4768), .B2(n6040), .C1(n4664), .C2(n4784), .A(n2533), 
        .ZN(N652) );
  OAI221_X2 U3266 ( .B1(n4768), .B2(n6041), .C1(n4663), .C2(n4784), .A(n4779), 
        .ZN(N651) );
  OAI221_X2 U3269 ( .B1(n4768), .B2(n6042), .C1(n4662), .C2(n4784), .A(n4780), 
        .ZN(N650) );
  OAI221_X2 U3272 ( .B1(n4768), .B2(n6043), .C1(n4661), .C2(n4784), .A(n4780), 
        .ZN(N649) );
  OAI221_X2 U3275 ( .B1(n4768), .B2(n6044), .C1(n4660), .C2(n4784), .A(n4779), 
        .ZN(N648) );
  OAI221_X2 U3278 ( .B1(n4768), .B2(n6045), .C1(n4659), .C2(n4784), .A(n4779), 
        .ZN(N647) );
  OAI221_X2 U3281 ( .B1(n4768), .B2(n6046), .C1(n4658), .C2(n4784), .A(n4779), 
        .ZN(N646) );
  OAI221_X2 U3284 ( .B1(n4769), .B2(n6047), .C1(n4657), .C2(n4784), .A(n2533), 
        .ZN(N645) );
  OAI221_X2 U3287 ( .B1(n4769), .B2(n6048), .C1(n4656), .C2(n4784), .A(n2533), 
        .ZN(N644) );
  OAI221_X2 U3290 ( .B1(n4769), .B2(n6049), .C1(n4655), .C2(n4784), .A(n2533), 
        .ZN(N643) );
  OAI221_X2 U3293 ( .B1(n4769), .B2(n6050), .C1(n4654), .C2(n4784), .A(n2533), 
        .ZN(N642) );
  OAI221_X2 U3296 ( .B1(n4769), .B2(n6051), .C1(n4653), .C2(n4784), .A(n2533), 
        .ZN(N641) );
  OAI221_X2 U3299 ( .B1(n4769), .B2(n6052), .C1(n4652), .C2(n4784), .A(n2533), 
        .ZN(N640) );
  OAI221_X2 U3302 ( .B1(n4769), .B2(n6053), .C1(n4651), .C2(n4784), .A(n2533), 
        .ZN(N639) );
  OAI221_X2 U3305 ( .B1(n4769), .B2(n6054), .C1(n4650), .C2(n4784), .A(n2533), 
        .ZN(N638) );
  OAI221_X2 U3308 ( .B1(n4769), .B2(n6055), .C1(n4649), .C2(n4784), .A(n2533), 
        .ZN(N637) );
  OAI221_X2 U3311 ( .B1(n4769), .B2(n6056), .C1(n4648), .C2(n4784), .A(n4779), 
        .ZN(N636) );
  OAI221_X2 U3314 ( .B1(n4769), .B2(n6057), .C1(n4647), .C2(n4782), .A(n4780), 
        .ZN(N635) );
  OAI221_X2 U3317 ( .B1(n4770), .B2(n6058), .C1(n4646), .C2(n4782), .A(n4780), 
        .ZN(N634) );
  OAI221_X2 U3320 ( .B1(n4770), .B2(n6059), .C1(n4645), .C2(n4782), .A(n4780), 
        .ZN(N633) );
  OAI221_X2 U3323 ( .B1(n4770), .B2(n6060), .C1(n4644), .C2(n4782), .A(n4780), 
        .ZN(N632) );
  OAI221_X2 U3326 ( .B1(n4770), .B2(n6061), .C1(n4643), .C2(n4782), .A(n4780), 
        .ZN(N631) );
  OAI221_X2 U3329 ( .B1(n4770), .B2(n6062), .C1(n4642), .C2(n4782), .A(n4780), 
        .ZN(N630) );
  OAI221_X2 U3332 ( .B1(n4770), .B2(n6063), .C1(n4641), .C2(n4782), .A(n4780), 
        .ZN(N629) );
  OAI221_X2 U3335 ( .B1(n4770), .B2(n6064), .C1(n4640), .C2(n4782), .A(n4780), 
        .ZN(N628) );
  OAI221_X2 U3338 ( .B1(n4770), .B2(n6065), .C1(n4639), .C2(n4782), .A(n4780), 
        .ZN(N627) );
  OAI221_X2 U3341 ( .B1(n4770), .B2(n6066), .C1(n4638), .C2(n4782), .A(n4780), 
        .ZN(N626) );
  OAI221_X2 U3344 ( .B1(n4770), .B2(n6067), .C1(n4637), .C2(n2532), .A(n4780), 
        .ZN(N625) );
  OAI221_X2 U3347 ( .B1(n4770), .B2(n6068), .C1(n4636), .C2(n2532), .A(n4780), 
        .ZN(N624) );
  OAI221_X2 U3350 ( .B1(n4771), .B2(n6069), .C1(n4635), .C2(n2532), .A(n4780), 
        .ZN(N623) );
  OAI221_X2 U3353 ( .B1(n4771), .B2(n6070), .C1(n4524), .C2(n4782), .A(n4779), 
        .ZN(N622) );
  OAI221_X2 U3356 ( .B1(n4771), .B2(n6071), .C1(n4460), .C2(n2532), .A(n4780), 
        .ZN(N621) );
  OAI221_X2 U3359 ( .B1(n4771), .B2(n6072), .C1(n4459), .C2(n2532), .A(n4780), 
        .ZN(N620) );
  OAI221_X2 U3362 ( .B1(n4771), .B2(n6073), .C1(n4458), .C2(n2532), .A(n4780), 
        .ZN(N619) );
  OAI221_X2 U3365 ( .B1(n4771), .B2(n6074), .C1(n4457), .C2(n2532), .A(n4780), 
        .ZN(N618) );
  OAI221_X2 U3368 ( .B1(n4771), .B2(n6075), .C1(n4456), .C2(n2532), .A(n4780), 
        .ZN(N617) );
  OAI221_X2 U3371 ( .B1(n4771), .B2(n6076), .C1(n4455), .C2(n2532), .A(n4780), 
        .ZN(N616) );
  OAI221_X2 U3374 ( .B1(n4771), .B2(n6077), .C1(n4454), .C2(n2532), .A(n4780), 
        .ZN(N615) );
  NAND2_X2 U3375 ( .A1(N400), .A2(n1090), .ZN(n2533) );
  OAI221_X2 U3378 ( .B1(n4771), .B2(n6078), .C1(n4453), .C2(n2532), .A(n2633), 
        .ZN(N614) );
  AOI22_X2 U3379 ( .A1(N399), .A2(n4811), .B1(n1091), .B2(N342), .ZN(n2633) );
  OAI221_X2 U3382 ( .B1(n4771), .B2(n6079), .C1(n4452), .C2(n2532), .A(n2636), 
        .ZN(N613) );
  AOI22_X2 U3383 ( .A1(N398), .A2(n4813), .B1(opa_r1[51]), .B2(n1091), .ZN(
        n2636) );
  OAI221_X2 U3386 ( .B1(n4770), .B2(n6080), .C1(n4421), .C2(n2532), .A(n2639), 
        .ZN(N612) );
  AOI22_X2 U3387 ( .A1(N397), .A2(n4813), .B1(opa_r1[50]), .B2(n1091), .ZN(
        n2639) );
  OAI221_X2 U3390 ( .B1(n4771), .B2(n6081), .C1(n4420), .C2(n2532), .A(n2642), 
        .ZN(N611) );
  AOI22_X2 U3391 ( .A1(N396), .A2(n4812), .B1(opa_r1[49]), .B2(n1091), .ZN(
        n2642) );
  OAI221_X2 U3394 ( .B1(n4770), .B2(n4402), .C1(n4451), .C2(n2532), .A(n2645), 
        .ZN(N610) );
  AOI22_X2 U3395 ( .A1(N395), .A2(n4811), .B1(opa_r1[48]), .B2(n1091), .ZN(
        n2645) );
  AOI22_X2 U3399 ( .A1(N394), .A2(n4813), .B1(opa_r1[47]), .B2(n1091), .ZN(
        n2648) );
  AOI22_X2 U3403 ( .A1(N393), .A2(n4813), .B1(opa_r1[46]), .B2(n1091), .ZN(
        n2651) );
  AND2_X2 U3404 ( .A1(n6381), .A2(n2337), .ZN(n1091) );
  NAND2_X2 U3406 ( .A1(n2337), .A2(n1308), .ZN(n2532) );
  OAI22_X2 U3413 ( .A1(sign_mul), .A2(n4505), .B1(sign_fasu), .B2(fpu_op_r2[1]), .ZN(n2337) );
  NAND4_X2 U3415 ( .A1(n4509), .A2(n4622), .A3(n2653), .A4(n2654), .ZN(N342)
         );
  NOR4_X2 U3416 ( .A1(n2655), .A2(opa_r1[57]), .A3(opa_r1[59]), .A4(opa_r1[58]), .ZN(n2654) );
  FA_X1 u4_sub_410_U2_1 ( .A(div_opa_ldz_r2[1]), .B(n4588), .CI(
        u4_sub_410_carry[1]), .CO(u4_sub_410_carry[2]), .S(u4_div_shft4[1]) );
  FA_X1 u4_sub_410_U2_2 ( .A(div_opa_ldz_r2[2]), .B(n4425), .CI(
        u4_sub_410_carry[2]), .CO(u4_sub_410_carry[3]), .S(u4_div_shft4[2]) );
  FA_X1 u4_sub_410_U2_3 ( .A(div_opa_ldz_r2[3]), .B(n4473), .CI(
        u4_sub_410_carry[3]), .CO(u4_sub_410_carry[4]), .S(u4_div_shft4[3]) );
  FA_X1 u4_sub_410_U2_4 ( .A(div_opa_ldz_r2[4]), .B(n4424), .CI(
        u4_sub_410_carry[4]), .CO(u4_sub_410_carry[5]), .S(u4_div_shft4[4]) );
  FA_X1 u4_add_409_U1_1 ( .A(div_opa_ldz_r2[1]), .B(n4368), .CI(
        u4_add_409_carry[1]), .CO(u4_add_409_carry[2]), .S(u4_div_shft3_1_) );
  FA_X1 u4_add_409_U1_2 ( .A(div_opa_ldz_r2[2]), .B(exp_r[2]), .CI(
        u4_add_409_carry[2]), .CO(u4_add_409_carry[3]), .S(u4_div_shft3_2_) );
  FA_X1 u4_add_409_U1_3 ( .A(div_opa_ldz_r2[3]), .B(exp_r[3]), .CI(
        u4_add_409_carry[3]), .CO(u4_add_409_carry[4]), .S(u4_div_shft3_3_) );
  FA_X1 u4_add_409_U1_4 ( .A(div_opa_ldz_r2[4]), .B(n4399), .CI(
        u4_add_409_carry[4]), .CO(u4_add_409_carry[5]), .S(u4_div_shft3_4_) );
  FA_X1 u4_sub_407_U2_1 ( .A(n4368), .B(n4578), .CI(u4_sub_407_carry[1]), .CO(
        u4_sub_407_carry[2]), .S(u4_div_scht1a[1]) );
  FA_X1 u4_sub_407_U2_2 ( .A(exp_r[2]), .B(n4577), .CI(u4_sub_407_carry[2]), 
        .CO(u4_sub_407_carry[3]), .S(u4_div_scht1a[2]) );
  FA_X1 u4_sub_407_U2_3 ( .A(exp_r[3]), .B(n4576), .CI(u4_sub_407_carry[3]), 
        .CO(u4_sub_407_carry[4]), .S(u4_div_scht1a[3]) );
  FA_X1 u4_sub_407_U2_4 ( .A(n4399), .B(n4581), .CI(u4_sub_407_carry[4]), .CO(
        u4_sub_407_carry[5]), .S(u4_div_scht1a[4]) );
  FA_X1 sub_1_root_sub_0_root_u4_add_495_U2_1 ( .A(u4_fi_ldz_2a_1_), .B(n4578), 
        .CI(sub_1_root_sub_0_root_u4_add_495_carry[1]), .CO(
        sub_1_root_sub_0_root_u4_add_495_carry[2]), .S(u4_ldz_dif_1_) );
  FA_X1 sub_1_root_sub_0_root_u4_add_495_U2_2 ( .A(u4_fi_ldz_2a_2_), .B(n4577), 
        .CI(sub_1_root_sub_0_root_u4_add_495_carry[2]), .CO(
        sub_1_root_sub_0_root_u4_add_495_carry[3]), .S(u4_ldz_dif_2_) );
  FA_X1 sub_1_root_sub_0_root_u4_add_495_U2_3 ( .A(u4_fi_ldz_2a_3_), .B(n4576), 
        .CI(sub_1_root_sub_0_root_u4_add_495_carry[3]), .CO(
        sub_1_root_sub_0_root_u4_add_495_carry[4]), .S(u4_ldz_dif_3_) );
  FA_X1 sub_1_root_sub_0_root_u4_add_495_U2_4 ( .A(u4_fi_ldz_2a_4_), .B(n4581), 
        .CI(sub_1_root_sub_0_root_u4_add_495_carry[4]), .CO(
        sub_1_root_sub_0_root_u4_add_495_carry[5]), .S(u4_ldz_dif_4_) );
  OAI21_X4 U3425 ( .B1(n4818), .B2(n4706), .A(n2472), .ZN(N737) );
  OAI21_X4 U3426 ( .B1(n4818), .B2(n4631), .A(n2474), .ZN(N736) );
  AOI222_X1 U3427 ( .A1(fract_i2f[104]), .A2(n4776), .B1(1'b0), .B2(n4787), 
        .C1(fract_out_q[55]), .C2(n4772), .ZN(n2344) );
  AOI222_X1 U3428 ( .A1(fract_i2f[103]), .A2(n4775), .B1(1'b0), .B2(n2342), 
        .C1(fract_out_q[54]), .C2(n4773), .ZN(n2346) );
  NOR2_X4 U3429 ( .A1(remainder[56]), .A2(remainder[55]), .ZN(n2231) );
  NOR2_X4 U3430 ( .A1(remainder[51]), .A2(remainder[52]), .ZN(n2230) );
  NOR2_X2 U3431 ( .A1(fract_denorm[38]), .A2(fract_denorm[37]), .ZN(n2156) );
  NOR2_X2 U3432 ( .A1(fract_denorm[9]), .A2(fract_denorm[8]), .ZN(n2162) );
  NOR2_X2 U3433 ( .A1(fract_denorm[10]), .A2(fract_denorm[0]), .ZN(n2170) );
  NOR3_X2 U3434 ( .A1(fract_denorm[95]), .A2(fract_denorm[96]), .A3(n6513), 
        .ZN(n432) );
  NAND3_X2 U3435 ( .A1(n2175), .A2(n1741), .A3(exp_ovf_r_1_), .ZN(n2174) );
  NOR2_X2 U3436 ( .A1(n1749), .A2(n2268), .ZN(n2171) );
  NOR2_X2 U3437 ( .A1(fract_denorm[22]), .A2(fract_denorm[21]), .ZN(n2168) );
  NOR3_X2 U3438 ( .A1(fract_denorm[47]), .A2(fract_denorm[48]), .A3(
        fract_denorm[46]), .ZN(n369) );
  NOR2_X2 U3439 ( .A1(n6527), .A2(u4_exp_in_pl1_1_), .ZN(n283) );
  NOR3_X2 U3440 ( .A1(n4359), .A2(n4428), .A3(n4369), .ZN(n1710) );
  AOI222_X1 U3441 ( .A1(u4_div_scht1a[5]), .A2(n255), .B1(u4_fi_ldz_5_), .B2(
        n261), .C1(u4_exp_in_pl1_5_), .C2(n262), .ZN(n264) );
  NOR2_X2 U3442 ( .A1(n4873), .A2(n431), .ZN(n426) );
  AOI21_X2 U3443 ( .B1(fract_denorm[94]), .B2(n432), .A(n433), .ZN(n431) );
  NOR2_X2 U3444 ( .A1(fract_denorm[15]), .A2(n329), .ZN(n425) );
  NOR2_X2 U3445 ( .A1(fract_denorm[3]), .A2(fract_denorm[4]), .ZN(n478) );
  NOR2_X2 U3446 ( .A1(fract_denorm[35]), .A2(fract_denorm[36]), .ZN(n393) );
  NOR3_X2 U3447 ( .A1(fract_denorm[97]), .A2(fract_denorm[98]), .A3(n394), 
        .ZN(n465) );
  NOR3_X2 U3448 ( .A1(fract_denorm[65]), .A2(fract_denorm[66]), .A3(
        fract_denorm[64]), .ZN(n307) );
  NAND3_X2 U3449 ( .A1(n319), .A2(n6480), .A3(n305), .ZN(n308) );
  NOR3_X2 U3450 ( .A1(fract_denorm[62]), .A2(fract_denorm[63]), .A3(
        fract_denorm[61]), .ZN(n309) );
  NOR2_X2 U3451 ( .A1(fract_denorm[73]), .A2(fract_denorm[72]), .ZN(n529) );
  NOR3_X2 U3452 ( .A1(fract_denorm[14]), .A2(fract_denorm[15]), .A3(
        fract_denorm[13]), .ZN(n328) );
  NOR2_X2 U3453 ( .A1(fract_denorm[76]), .A2(fract_denorm[75]), .ZN(n345) );
  NOR3_X2 U3454 ( .A1(fract_denorm[78]), .A2(fract_denorm[79]), .A3(
        fract_denorm[77]), .ZN(n350) );
  NOR3_X2 U3455 ( .A1(fract_denorm[93]), .A2(fract_denorm[94]), .A3(n6511), 
        .ZN(n354) );
  NOR2_X2 U3456 ( .A1(n318), .A2(n376), .ZN(n372) );
  NAND3_X2 U3457 ( .A1(n6471), .A2(n6472), .A3(n6468), .ZN(n371) );
  OAI21_X2 U3458 ( .B1(fract_denorm[53]), .B2(fract_denorm[50]), .A(n375), 
        .ZN(n374) );
  NOR3_X2 U3459 ( .A1(u4_fract_out_12_), .A2(u4_fract_out_14_), .A3(
        u4_fract_out_13_), .ZN(n2206) );
  NOR3_X2 U3460 ( .A1(u4_fract_out_24_), .A2(u4_fract_out_26_), .A3(
        u4_fract_out_25_), .ZN(n2215) );
  NOR3_X2 U3461 ( .A1(u4_fract_out_48_), .A2(u4_fract_out_4_), .A3(
        u4_fract_out_49_), .ZN(n2193) );
  NOR3_X2 U3462 ( .A1(u4_fract_out_36_), .A2(u4_fract_out_38_), .A3(
        u4_fract_out_37_), .ZN(n2182) );
  NOR3_X2 U3463 ( .A1(n4368), .A2(exp_r[3]), .A3(exp_r[2]), .ZN(n1709) );
  AOI21_X2 U3464 ( .B1(u4_N6269), .B2(n1705), .A(u4_N6267), .ZN(n1723) );
  NAND3_X2 U3465 ( .A1(n4401), .A2(n1701), .A3(n4767), .ZN(n1724) );
  NOR2_X2 U3466 ( .A1(n1711), .A2(n4401), .ZN(n1703) );
  AOI222_X1 U3467 ( .A1(u4_N6273), .A2(u4_N6272), .B1(n1712), .B2(n1713), .C1(
        n1714), .C2(n1705), .ZN(n1711) );
  NOR3_X2 U3468 ( .A1(remainder[94]), .A2(remainder[96]), .A3(remainder[95]), 
        .ZN(n2244) );
  NOR3_X2 U3469 ( .A1(remainder[88]), .A2(remainder[8]), .A3(remainder[89]), 
        .ZN(n2242) );
  NOR3_X2 U3470 ( .A1(remainder[0]), .A2(remainder[101]), .A3(remainder[100]), 
        .ZN(n2250) );
  NOR3_X2 U3471 ( .A1(remainder[102]), .A2(remainder[104]), .A3(remainder[103]), .ZN(n2251) );
  NOR3_X2 U3472 ( .A1(remainder[105]), .A2(remainder[107]), .A3(remainder[106]), .ZN(n2252) );
  NOR3_X2 U3473 ( .A1(remainder[14]), .A2(remainder[16]), .A3(remainder[15]), 
        .ZN(n2254) );
  NOR3_X2 U3474 ( .A1(remainder[20]), .A2(remainder[22]), .A3(remainder[21]), 
        .ZN(n2256) );
  NOR3_X2 U3475 ( .A1(remainder[27]), .A2(remainder[29]), .A3(remainder[28]), 
        .ZN(n2258) );
  NOR3_X2 U3476 ( .A1(remainder[2]), .A2(remainder[31]), .A3(remainder[30]), 
        .ZN(n2259) );
  NOR3_X2 U3477 ( .A1(remainder[32]), .A2(remainder[34]), .A3(remainder[33]), 
        .ZN(n2260) );
  NOR3_X2 U3478 ( .A1(remainder[39]), .A2(remainder[40]), .A3(remainder[3]), 
        .ZN(n2262) );
  NOR3_X2 U3479 ( .A1(remainder[45]), .A2(remainder[47]), .A3(remainder[46]), 
        .ZN(n2264) );
  NOR3_X2 U3480 ( .A1(remainder[57]), .A2(remainder[59]), .A3(remainder[58]), 
        .ZN(n2232) );
  NOR3_X2 U3481 ( .A1(remainder[63]), .A2(remainder[65]), .A3(remainder[64]), 
        .ZN(n2234) );
  NOR3_X2 U3482 ( .A1(remainder[6]), .A2(remainder[71]), .A3(remainder[70]), 
        .ZN(n2236) );
  NOR3_X2 U3483 ( .A1(remainder[76]), .A2(remainder[78]), .A3(remainder[77]), 
        .ZN(n2238) );
  NOR3_X2 U3484 ( .A1(remainder[79]), .A2(remainder[80]), .A3(remainder[7]), 
        .ZN(n2239) );
  NOR3_X2 U3485 ( .A1(remainder[81]), .A2(remainder[83]), .A3(remainder[82]), 
        .ZN(n2240) );
  NOR3_X2 U3486 ( .A1(u4_N6014), .A2(u4_N6016), .A3(u4_N6015), .ZN(n2298) );
  NOR3_X2 U3487 ( .A1(u4_N6011), .A2(u4_N6013), .A3(u4_N6012), .ZN(n2297) );
  NOR3_X2 U3488 ( .A1(u4_N6008), .A2(u4_N6010), .A3(u4_N6009), .ZN(n2296) );
  NOR3_X2 U3489 ( .A1(u4_N6034), .A2(u4_N6036), .A3(u4_N6035), .ZN(n2304) );
  NOR3_X2 U3490 ( .A1(u4_N6037), .A2(u4_N6039), .A3(u4_N6038), .ZN(n2305) );
  NOR3_X2 U3491 ( .A1(u4_N6040), .A2(u4_N6042), .A3(u4_N6041), .ZN(n2306) );
  NOR3_X2 U3492 ( .A1(u4_N6047), .A2(u4_N6049), .A3(u4_N6048), .ZN(n2308) );
  NOR3_X2 U3493 ( .A1(u4_N6054), .A2(u4_N6056), .A3(u4_N6055), .ZN(n2310) );
  NOR3_X2 U3494 ( .A1(u4_N6021), .A2(u4_N6023), .A3(u4_N6022), .ZN(n2300) );
  NOR3_X2 U3495 ( .A1(u4_N6027), .A2(u4_N6029), .A3(u4_N6028), .ZN(n2302) );
  NOR3_X2 U3496 ( .A1(u4_N6024), .A2(u4_N6026), .A3(u4_N6025), .ZN(n2301) );
  AOI21_X2 U3497 ( .B1(sign), .B2(rmode_r3[1]), .A(n6379), .ZN(n1936) );
  OAI21_X2 U3498 ( .B1(sign), .B2(n2145), .A(n2146), .ZN(n1946) );
  AOI211_X2 U3499 ( .C1(n2150), .C2(n2151), .A(opas_r2), .B(n4875), .ZN(n2147)
         );
  OAI21_X2 U3500 ( .B1(u4_fract_out_0_), .B2(n2058), .A(n2059), .ZN(n1941) );
  NOR3_X2 U3501 ( .A1(n1947), .A2(n1679), .A3(n1681), .ZN(n1933) );
  NAND3_X2 U3502 ( .A1(n1970), .A2(n1971), .A3(n1969), .ZN(n1987) );
  NOR3_X2 U3503 ( .A1(n5012), .A2(u4_fi_ldz_2a_6_), .A3(u4_fi_ldz_2a_5_), .ZN(
        u4_N6240) );
  OAI21_X2 U3504 ( .B1(n1671), .B2(n2056), .A(n2057), .ZN(n2055) );
  OAI21_X2 U3505 ( .B1(n2023), .B2(n1941), .A(n5046), .ZN(n2057) );
  INV_X4 U3506 ( .A(n4828), .ZN(n4827) );
  INV_X4 U3507 ( .A(u1_expa_lt_expb), .ZN(n4828) );
  INV_X4 U3508 ( .A(n4827), .ZN(n4850) );
  INV_X4 U3509 ( .A(n4847), .ZN(n4840) );
  INV_X4 U3510 ( .A(n4847), .ZN(n4841) );
  NOR2_X2 U3511 ( .A1(fract_denorm[27]), .A2(fract_denorm[28]), .ZN(n334) );
  NOR3_X2 U3512 ( .A1(fract_denorm[37]), .A2(fract_denorm[38]), .A3(n496), 
        .ZN(n392) );
  NOR2_X2 U3513 ( .A1(fract_denorm[12]), .A2(fract_denorm[11]), .ZN(n341) );
  NOR3_X2 U3514 ( .A1(fract_denorm[52]), .A2(fract_denorm[53]), .A3(n6469), 
        .ZN(n401) );
  NOR2_X2 U3515 ( .A1(n329), .A2(n6422), .ZN(n337) );
  NOR3_X2 U3516 ( .A1(fract_denorm[29]), .A2(fract_denorm[30]), .A3(n421), 
        .ZN(n333) );
  OAI21_X2 U3517 ( .B1(n518), .B2(n519), .A(n4874), .ZN(n512) );
  NOR3_X2 U3518 ( .A1(n6506), .A2(fract_denorm[92]), .A3(n6509), .ZN(n518) );
  NOR3_X2 U3519 ( .A1(fract_denorm[101]), .A2(fract_denorm[102]), .A3(
        fract_denorm[100]), .ZN(n418) );
  NOR3_X2 U3520 ( .A1(fract_denorm[87]), .A2(fract_denorm[88]), .A3(n454), 
        .ZN(n416) );
  NOR2_X2 U3521 ( .A1(fract_denorm[86]), .A2(fract_denorm[85]), .ZN(n346) );
  NOR2_X2 U3522 ( .A1(fract_denorm[70]), .A2(fract_denorm[69]), .ZN(n319) );
  NOR2_X2 U3523 ( .A1(n6485), .A2(fract_denorm[68]), .ZN(n305) );
  NAND3_X2 U3524 ( .A1(n544), .A2(n6449), .A3(n6452), .ZN(n496) );
  NOR3_X2 U3525 ( .A1(fract_denorm[24]), .A2(fract_denorm[25]), .A3(
        fract_denorm[23]), .ZN(n330) );
  NOR2_X2 U3526 ( .A1(fract_denorm[6]), .A2(fract_denorm[7]), .ZN(n505) );
  NOR3_X2 U3527 ( .A1(fract_denorm[54]), .A2(fract_denorm[55]), .A3(n419), 
        .ZN(n375) );
  NOR3_X2 U3528 ( .A1(fract_denorm[32]), .A2(fract_denorm[33]), .A3(n461), 
        .ZN(n536) );
  NOR3_X2 U3529 ( .A1(n6459), .A2(fract_denorm[48]), .A3(n368), .ZN(n537) );
  NOR3_X2 U3530 ( .A1(n6510), .A2(fract_denorm[96]), .A3(n6513), .ZN(n540) );
  NAND3_X2 U3531 ( .A1(n6471), .A2(n6472), .A3(n370), .ZN(n419) );
  NOR3_X2 U3532 ( .A1(n6508), .A2(fract_denorm[94]), .A3(n6511), .ZN(n553) );
  NOR3_X2 U3533 ( .A1(n6439), .A2(fract_denorm[30]), .A3(n421), .ZN(n550) );
  NAND3_X2 U3534 ( .A1(n393), .A2(n6444), .A3(n392), .ZN(n461) );
  NOR3_X2 U3535 ( .A1(n6427), .A2(fract_denorm[18]), .A3(n387), .ZN(n564) );
  NOR2_X2 U3536 ( .A1(fract_denorm[66]), .A2(n308), .ZN(n567) );
  AOI222_X1 U3537 ( .A1(n4400), .A2(n6390), .B1(u4_div_scht1a[0]), .B2(n255), 
        .C1(n4823), .C2(n253), .ZN(n287) );
  AOI222_X1 U3538 ( .A1(u4_f2i_shft_1_), .A2(n6390), .B1(u4_div_scht1a[1]), 
        .B2(n255), .C1(n4368), .C2(n253), .ZN(n275) );
  AOI222_X1 U3539 ( .A1(u4_f2i_shft_2_), .A2(n6390), .B1(u4_div_scht1a[2]), 
        .B2(n255), .C1(exp_r[2]), .C2(n253), .ZN(n274) );
  AOI222_X1 U3540 ( .A1(u4_f2i_shft_4_), .A2(n6390), .B1(u4_div_scht1a[4]), 
        .B2(n255), .C1(n4399), .C2(n253), .ZN(n267) );
  NAND3_X2 U3541 ( .A1(n1708), .A2(n6520), .A3(n2332), .ZN(n289) );
  OAI21_X2 U3542 ( .B1(n1701), .B2(n1737), .A(n4401), .ZN(n2332) );
  AOI222_X1 U3543 ( .A1(u4_f2i_shft_3_), .A2(n6390), .B1(u4_div_scht1a[3]), 
        .B2(n255), .C1(exp_r[3]), .C2(n253), .ZN(n271) );
  NOR2_X2 U3544 ( .A1(n6389), .A2(n293), .ZN(n291) );
  NOR3_X2 U3545 ( .A1(n4821), .A2(n294), .A3(n295), .ZN(n293) );
  INV_X4 U3546 ( .A(n288), .ZN(n253) );
  NAND3_X2 U3547 ( .A1(n6413), .A2(n6412), .A3(fract_denorm[6]), .ZN(n413) );
  AOI222_X1 U3548 ( .A1(fract_denorm[92]), .A2(n354), .B1(fract_denorm[60]), 
        .B2(n6475), .C1(fract_denorm[76]), .C2(n6492), .ZN(n481) );
  NAND3_X2 U3549 ( .A1(n401), .A2(n6465), .A3(fract_denorm[50]), .ZN(n396) );
  NAND3_X2 U3550 ( .A1(n392), .A2(n393), .A3(fract_denorm[34]), .ZN(n391) );
  AOI211_X2 U3551 ( .C1(n425), .C2(fract_denorm[14]), .A(n426), .B(n427), .ZN(
        n424) );
  AOI21_X2 U3552 ( .B1(n457), .B2(n6407), .A(n459), .ZN(n456) );
  AOI211_X2 U3553 ( .C1(fract_denorm[96]), .C2(n465), .A(n466), .B(n467), .ZN(
        n455) );
  AOI21_X2 U3554 ( .B1(fract_denorm[88]), .B2(n6504), .A(n450), .ZN(n448) );
  NAND3_X2 U3555 ( .A1(n370), .A2(n6472), .A3(fract_denorm[56]), .ZN(n447) );
  NOR3_X2 U3556 ( .A1(fract_denorm[10]), .A2(fract_denorm[9]), .A3(n296), .ZN(
        n439) );
  NOR3_X2 U3557 ( .A1(fract_denorm[44]), .A2(fract_denorm[45]), .A3(
        fract_denorm[43]), .ZN(n367) );
  NOR3_X2 U3558 ( .A1(n6487), .A2(fract_denorm[71]), .A3(n6488), .ZN(n315) );
  NOR2_X2 U3559 ( .A1(n6490), .A2(n312), .ZN(n304) );
  NAND3_X2 U3560 ( .A1(n333), .A2(n334), .A3(fract_denorm[26]), .ZN(n332) );
  NOR3_X2 U3561 ( .A1(n420), .A2(n6432), .A3(n6430), .ZN(n325) );
  OAI21_X2 U3562 ( .B1(fract_denorm[88]), .B2(fract_denorm[89]), .A(n357), 
        .ZN(n352) );
  AOI222_X1 U3563 ( .A1(n335), .A2(n336), .B1(n337), .B2(n6417), .C1(n6434), 
        .C2(n6432), .ZN(n322) );
  NAND3_X2 U3564 ( .A1(n4438), .A2(n4507), .A3(n4406), .ZN(n1541) );
  NAND3_X2 U3565 ( .A1(n4513), .A2(n4436), .A3(n4405), .ZN(n1550) );
  NAND3_X2 U3566 ( .A1(n4512), .A2(n4435), .A3(n4386), .ZN(n1573) );
  NAND3_X2 U3567 ( .A1(n4511), .A2(n4434), .A3(n4404), .ZN(n1586) );
  NAND3_X2 U3568 ( .A1(n4510), .A2(n4387), .A3(n4403), .ZN(n1595) );
  NAND3_X2 U3569 ( .A1(n1637), .A2(n1731), .A3(n1630), .ZN(n1728) );
  NOR3_X2 U3570 ( .A1(n1638), .A2(n1633), .A3(n1634), .ZN(n1726) );
  NAND3_X2 U3571 ( .A1(n1696), .A2(n4479), .A3(n1698), .ZN(n1695) );
  NAND3_X2 U3572 ( .A1(n246), .A2(n4401), .A3(n1700), .ZN(n1698) );
  AOI21_X2 U3573 ( .B1(n4430), .B2(n4767), .A(n1701), .ZN(n1700) );
  AOI222_X1 U3574 ( .A1(u4_N6268), .A2(n1702), .B1(n1703), .B2(n4429), .C1(
        n1704), .C2(n1705), .ZN(n1694) );
  OAI21_X2 U3575 ( .B1(n1723), .B2(n247), .A(n1724), .ZN(n1702) );
  OAI21_X2 U3576 ( .B1(n1706), .B2(n1707), .A(n1708), .ZN(n1704) );
  NAND3_X2 U3577 ( .A1(n1832), .A2(n1833), .A3(n1834), .ZN(n1828) );
  NAND3_X2 U3578 ( .A1(n1817), .A2(n1818), .A3(n1819), .ZN(n1813) );
  OAI21_X2 U3579 ( .B1(n2148), .B2(n4821), .A(n2149), .ZN(n2058) );
  NOR2_X2 U3580 ( .A1(n2148), .A2(n2269), .ZN(n2059) );
  NAND3_X2 U3581 ( .A1(n1933), .A2(n1934), .A3(n1935), .ZN(n1932) );
  OAI21_X2 U3582 ( .B1(n1939), .B2(n1682), .A(n1933), .ZN(n1931) );
  NOR3_X2 U3583 ( .A1(n1936), .A2(n4822), .A3(n6161), .ZN(n1935) );
  OAI21_X2 U3584 ( .B1(r482_B_0_), .B2(n1941), .A(n1942), .ZN(n1940) );
  NAND3_X2 U3585 ( .A1(n1800), .A2(n1632), .A3(n1631), .ZN(n1948) );
  NAND3_X2 U3586 ( .A1(n1637), .A2(n1638), .A3(n1630), .ZN(n1950) );
  NOR3_X2 U3587 ( .A1(n1964), .A2(n1965), .A3(n1957), .ZN(n1985) );
  OAI21_X2 U3588 ( .B1(n2030), .B2(n6401), .A(n5979), .ZN(n1981) );
  NOR3_X2 U3589 ( .A1(n6528), .A2(exp_ovf_r_1_), .A3(n4430), .ZN(n2030) );
  OAI21_X2 U3590 ( .B1(n6527), .B2(n4875), .A(n6400), .ZN(n1979) );
  AOI21_X2 U3591 ( .B1(n6528), .B2(n4430), .A(n5979), .ZN(n2041) );
  AOI21_X2 U3592 ( .B1(u4_N6240), .B2(n1678), .A(n5979), .ZN(n2040) );
  NAND3_X2 U3593 ( .A1(n6528), .A2(n2063), .A3(u4_N6238), .ZN(n2061) );
  NAND3_X2 U3594 ( .A1(opb_dn), .A2(n4426), .A3(u4_N6179), .ZN(n1974) );
  NAND3_X2 U3595 ( .A1(n2013), .A2(n2014), .A3(n2015), .ZN(n1957) );
  AOI222_X1 U3596 ( .A1(u4_exp_out_mi1[8]), .A2(n1995), .B1(u4_exp_fix_divb[8]), .B2(n1992), .C1(n1997), .C2(n4369), .ZN(n2015) );
  NAND3_X2 U3597 ( .A1(n2024), .A2(n2025), .A3(n2026), .ZN(n1964) );
  AOI222_X1 U3598 ( .A1(u4_exp_out_mi1[9]), .A2(n1995), .B1(u4_exp_fix_divb[9]), .B2(n1992), .C1(n1997), .C2(n4428), .ZN(n2026) );
  OAI21_X2 U3599 ( .B1(n4427), .B2(n2054), .A(n2020), .ZN(n2016) );
  NOR2_X2 U3600 ( .A1(n1745), .A2(n2032), .ZN(n1939) );
  AOI222_X1 U3601 ( .A1(u4_exp_out_mi1[1]), .A2(n1995), .B1(u4_exp_fix_divb[1]), .B2(n1992), .C1(n1997), .C2(n4368), .ZN(n2019) );
  OAI21_X2 U3602 ( .B1(n2022), .B2(n2023), .A(rmode_r3[1]), .ZN(n2021) );
  OAI21_X2 U3603 ( .B1(n1740), .B2(n2051), .A(n2052), .ZN(n1994) );
  NAND3_X2 U3604 ( .A1(u4_fract_out_pl1_52_), .A2(n5046), .A3(n1944), .ZN(
        n2052) );
  AOI222_X1 U3605 ( .A1(n1991), .A2(u4_exp_next_mi_2_), .B1(u4_exp_fix_divb[2]), .B2(n1992), .C1(u4_exp_fix_diva[2]), .C2(n1993), .ZN(n2000) );
  AOI222_X1 U3606 ( .A1(n1991), .A2(u4_exp_next_mi_4_), .B1(u4_exp_fix_divb[4]), .B2(n1992), .C1(u4_exp_fix_diva[4]), .C2(n1993), .ZN(n1990) );
  AOI222_X1 U3607 ( .A1(n1991), .A2(u4_exp_next_mi_3_), .B1(u4_exp_fix_divb[3]), .B2(n1992), .C1(u4_exp_fix_diva[3]), .C2(n1993), .ZN(n2003) );
  AOI222_X1 U3608 ( .A1(u4_exp_out_mi1[0]), .A2(n1995), .B1(u4_exp_fix_divb[0]), .B2(n1992), .C1(n1997), .C2(n4823), .ZN(n2029) );
  INV_X4 U3609 ( .A(n4850), .ZN(n4849) );
  INV_X4 U3610 ( .A(n4827), .ZN(n4851) );
  INV_X4 U3611 ( .A(n4850), .ZN(n4848) );
  NOR2_X2 U3612 ( .A1(n849), .A2(n4185), .ZN(n863) );
  NOR2_X2 U3613 ( .A1(n913), .A2(n6345), .ZN(n871) );
  NAND2_X2 U3614 ( .A1(n4826), .A2(n6373), .ZN(n773) );
  NOR3_X2 U3615 ( .A1(n912), .A2(n6303), .A3(n6293), .ZN(n908) );
  NOR3_X2 U3616 ( .A1(n903), .A2(n6302), .A3(n939), .ZN(n937) );
  NOR3_X2 U3617 ( .A1(n938), .A2(n6301), .A3(n939), .ZN(n940) );
  NOR2_X2 U3618 ( .A1(u1_exp_diff_4_), .A2(u1_exp_lt_27), .ZN(n938) );
  NOR2_X2 U3619 ( .A1(u1_exp_diff_3_), .A2(u1_exp_lt_27), .ZN(n903) );
  NOR2_X2 U3620 ( .A1(u1_exp_diff_5_), .A2(u1_exp_lt_27), .ZN(n912) );
  NOR2_X2 U3621 ( .A1(n6293), .A2(n938), .ZN(n904) );
  NAND3_X2 U3622 ( .A1(n6369), .A2(n1374), .A3(n1455), .ZN(n1430) );
  NOR3_X2 U3623 ( .A1(fracta_mul[7]), .A2(fracta_mul[9]), .A3(fracta_mul[8]), 
        .ZN(n1455) );
  NOR3_X2 U3624 ( .A1(n1284), .A2(fracta_mul[39]), .A3(n6363), .ZN(n1428) );
  NOR3_X2 U3625 ( .A1(n6409), .A2(fract_denorm[2]), .A3(n390), .ZN(n457) );
  NAND3_X2 U3626 ( .A1(n334), .A2(n6437), .A3(n333), .ZN(n331) );
  NOR3_X2 U3627 ( .A1(n318), .A2(fract_denorm[58]), .A3(n376), .ZN(n370) );
  NAND3_X2 U3628 ( .A1(n505), .A2(n6410), .A3(n6413), .ZN(n390) );
  NAND3_X2 U3629 ( .A1(n337), .A2(n6418), .A3(fract_denorm[11]), .ZN(n514) );
  NAND3_X2 U3630 ( .A1(n333), .A2(n6438), .A3(fract_denorm[27]), .ZN(n513) );
  NOR3_X2 U3631 ( .A1(n6432), .A2(fract_denorm[20]), .A3(n420), .ZN(n335) );
  NAND3_X2 U3632 ( .A1(n346), .A2(n6500), .A3(n416), .ZN(n349) );
  NAND3_X2 U3633 ( .A1(n305), .A2(n319), .A3(fract_denorm[67]), .ZN(n510) );
  AOI21_X2 U3634 ( .B1(fract_denorm[53]), .B2(n375), .A(n497), .ZN(n493) );
  AOI21_X2 U3635 ( .B1(fract_denorm[31]), .B2(n536), .A(n537), .ZN(n535) );
  NOR3_X2 U3636 ( .A1(n419), .A2(n4873), .A3(n6470), .ZN(n363) );
  NOR2_X2 U3637 ( .A1(fract_denorm[40]), .A2(fract_denorm[41]), .ZN(n544) );
  NOR2_X2 U3638 ( .A1(n549), .A2(n550), .ZN(n548) );
  NOR3_X2 U3639 ( .A1(n553), .A2(n554), .A3(n555), .ZN(n547) );
  NOR3_X2 U3640 ( .A1(n6490), .A2(fract_denorm[74]), .A3(n312), .ZN(n313) );
  AOI21_X2 U3641 ( .B1(n567), .B2(fract_denorm[65]), .A(n568), .ZN(n561) );
  AOI211_X2 U3642 ( .C1(fract_denorm[1]), .C2(n457), .A(n361), .B(n564), .ZN(
        n563) );
  AOI222_X1 U3643 ( .A1(u4_div_scht1a[6]), .A2(n255), .B1(u4_fi_ldz_6_), .B2(
        n261), .C1(u4_exp_in_pl1_6_), .C2(n262), .ZN(n260) );
  OAI21_X2 U3644 ( .B1(n4873), .B2(n412), .A(n413), .ZN(n411) );
  NOR3_X2 U3645 ( .A1(n403), .A2(n404), .A3(n405), .ZN(n382) );
  AOI211_X2 U3646 ( .C1(n384), .C2(n4874), .A(n385), .B(n386), .ZN(n383) );
  NOR2_X2 U3647 ( .A1(n2023), .A2(n1942), .ZN(n2050) );
  NOR2_X2 U3648 ( .A1(n300), .A2(n301), .ZN(n299) );
  AOI21_X2 U3649 ( .B1(n302), .B2(n303), .A(fract_denorm[105]), .ZN(n300) );
  AOI222_X1 U3650 ( .A1(n313), .A2(n6487), .B1(n315), .B2(n6483), .C1(n6475), 
        .C2(n318), .ZN(n302) );
  OAI21_X2 U3651 ( .B1(n342), .B2(n343), .A(n4874), .ZN(n321) );
  NAND3_X2 U3652 ( .A1(n4437), .A2(n4506), .A3(n4385), .ZN(n1618) );
  NAND3_X2 U3653 ( .A1(n1512), .A2(n1510), .A3(n1649), .ZN(n1647) );
  NOR3_X2 U3654 ( .A1(n1650), .A2(n1515), .A3(n1513), .ZN(n1645) );
  NOR3_X2 U3655 ( .A1(n1640), .A2(n1498), .A3(n1496), .ZN(n1639) );
  NAND3_X2 U3656 ( .A1(n1501), .A2(n1499), .A3(n1641), .ZN(n1640) );
  NAND3_X2 U3657 ( .A1(n1633), .A2(n1634), .A3(n1635), .ZN(n1629) );
  NOR3_X2 U3658 ( .A1(n1636), .A2(n1637), .A3(n1638), .ZN(n1627) );
  NOR3_X2 U3659 ( .A1(n4588), .A2(n4473), .A3(n4425), .ZN(n2065) );
  NAND3_X2 U3660 ( .A1(n4369), .A2(n4875), .A3(n4359), .ZN(n2067) );
  NOR2_X2 U3661 ( .A1(n1701), .A2(n1737), .ZN(n1736) );
  OAI21_X2 U3662 ( .B1(n4430), .B2(n1694), .A(n1695), .ZN(n1692) );
  NOR3_X2 U3663 ( .A1(n1682), .A2(n244), .A3(n1681), .ZN(n1693) );
  NAND3_X2 U3664 ( .A1(n1499), .A2(n1500), .A3(n1501), .ZN(n1495) );
  NAND3_X2 U3665 ( .A1(n1510), .A2(n1511), .A3(n1512), .ZN(n1506) );
  NOR3_X2 U3666 ( .A1(n1513), .A2(n1514), .A3(n1515), .ZN(n1504) );
  NOR3_X2 U3667 ( .A1(n1642), .A2(n1643), .A3(n1644), .ZN(n1493) );
  NAND3_X2 U3668 ( .A1(opa_inf), .A2(opb_inf), .A3(sign_exe_r), .ZN(n1773) );
  NOR2_X2 U3669 ( .A1(n2058), .A2(n2059), .ZN(n1749) );
  NAND3_X2 U3670 ( .A1(n4820), .A2(n1672), .A3(n1673), .ZN(n1490) );
  NAND3_X2 U3671 ( .A1(n4619), .A2(n4432), .A3(n1674), .ZN(n1672) );
  NOR2_X2 U3672 ( .A1(inf_mul_r), .A2(inf_mul2), .ZN(n1477) );
  NAND3_X2 U3673 ( .A1(n2064), .A2(u4_exp_out_0_), .A3(n2068), .ZN(n1684) );
  NOR3_X2 U3674 ( .A1(u4_N6891), .A2(n205), .A3(n4949), .ZN(n2068) );
  AOI21_X2 U3675 ( .B1(n4875), .B2(n4767), .A(n4430), .ZN(n1683) );
  NOR3_X2 U3676 ( .A1(n6379), .A2(n6390), .A3(n1508), .ZN(n1679) );
  OAI21_X2 U3677 ( .B1(n4822), .B2(n1732), .A(n1979), .ZN(n1977) );
  NAND3_X2 U3678 ( .A1(r482_B_0_), .A2(n1978), .A3(n6400), .ZN(n2035) );
  AOI211_X2 U3679 ( .C1(n6378), .C2(n1678), .A(n2037), .B(n2038), .ZN(n2034)
         );
  OAI21_X2 U3680 ( .B1(n1956), .B2(n1952), .A(n1953), .ZN(n1636) );
  OAI21_X2 U3681 ( .B1(n1961), .B2(n1952), .A(n1953), .ZN(n1638) );
  AOI222_X1 U3682 ( .A1(u4_exp_out_mi1[10]), .A2(n1995), .B1(
        u4_exp_fix_divb[10]), .B2(n1992), .C1(n1997), .C2(n4875), .ZN(n2048)
         );
  NOR3_X2 U3683 ( .A1(n244), .A2(r482_B_0_), .A3(n1685), .ZN(n1973) );
  OAI21_X2 U3684 ( .B1(n6385), .B2(n1965), .A(n1960), .ZN(n1637) );
  NAND3_X2 U3685 ( .A1(n2007), .A2(n2008), .A3(n2009), .ZN(n1971) );
  AOI222_X1 U3686 ( .A1(u4_exp_out_mi1[6]), .A2(n1995), .B1(u4_exp_fix_divb[6]), .B2(n1992), .C1(n1997), .C2(n4382), .ZN(n2009) );
  NAND3_X2 U3687 ( .A1(n2010), .A2(n2011), .A3(n2012), .ZN(n1970) );
  AOI222_X1 U3688 ( .A1(u4_exp_out_mi1[7]), .A2(n1995), .B1(u4_exp_fix_divb[7]), .B2(n1992), .C1(n1997), .C2(n4359), .ZN(n2012) );
  NAND3_X2 U3689 ( .A1(n2004), .A2(n2005), .A3(n2006), .ZN(n1969) );
  AOI222_X1 U3690 ( .A1(u4_exp_out_mi1[5]), .A2(n1995), .B1(u4_exp_fix_divb[5]), .B2(n1992), .C1(n1997), .C2(n4370), .ZN(n2006) );
  OAI21_X2 U3691 ( .B1(n6385), .B2(n1962), .A(n1953), .ZN(n1968) );
  NOR2_X2 U3692 ( .A1(n1947), .A2(n2336), .ZN(n1963) );
  NOR3_X2 U3693 ( .A1(n4401), .A2(n4430), .A3(n244), .ZN(n2336) );
  OAI21_X2 U3694 ( .B1(n1958), .B2(n6385), .A(n1960), .ZN(n1630) );
  OAI21_X2 U3695 ( .B1(n1967), .B2(n6385), .A(n1960), .ZN(n1632) );
  OAI21_X2 U3696 ( .B1(n1966), .B2(n6385), .A(n1960), .ZN(n1631) );
  OAI21_X2 U3697 ( .B1(n1951), .B2(n1952), .A(n1953), .ZN(n1731) );
  AOI21_X2 U3698 ( .B1(n4504), .B2(n4619), .A(n4821), .ZN(n1928) );
  INV_X4 U3699 ( .A(n4845), .ZN(n4844) );
  INV_X4 U3700 ( .A(n4835), .ZN(n4834) );
  INV_X4 U3701 ( .A(n4838), .ZN(n4830) );
  INV_X4 U3702 ( .A(n4837), .ZN(n4831) );
  INV_X4 U3703 ( .A(n4835), .ZN(n4833) );
  NOR2_X2 U3704 ( .A1(n815), .A2(n6340), .ZN(n875) );
  NOR2_X2 U3705 ( .A1(n827), .A2(n4166), .ZN(n885) );
  NOR2_X2 U3706 ( .A1(n823), .A2(n4170), .ZN(n886) );
  NAND3_X2 U3707 ( .A1(n925), .A2(n926), .A3(n863), .ZN(n911) );
  AOI222_X1 U3708 ( .A1(n6299), .A2(n905), .B1(n6290), .B2(n906), .C1(n6292), 
        .C2(n907), .ZN(n893) );
  AOI222_X1 U3709 ( .A1(n868), .A2(n913), .B1(n6298), .B2(n914), .C1(n6294), 
        .C2(n915), .ZN(n891) );
  NOR2_X2 U3710 ( .A1(n844), .A2(u1_adj_op_29_), .ZN(n819) );
  NOR2_X2 U3711 ( .A1(n847), .A2(n6330), .ZN(n817) );
  NOR2_X2 U3712 ( .A1(n851), .A2(n4177), .ZN(n809) );
  NOR2_X2 U3713 ( .A1(n855), .A2(n6338), .ZN(n811) );
  NAND3_X2 U3714 ( .A1(n912), .A2(n903), .A3(n904), .ZN(n812) );
  NAND3_X2 U3715 ( .A1(n6302), .A2(n903), .A3(n904), .ZN(n842) );
  NOR2_X2 U3716 ( .A1(n896), .A2(n6327), .ZN(n839) );
  NOR3_X2 U3717 ( .A1(n4158), .A2(n4157), .A3(n873), .ZN(n836) );
  NAND3_X2 U3718 ( .A1(n6301), .A2(n6302), .A3(n904), .ZN(n838) );
  INV_X4 U3719 ( .A(n903), .ZN(n6301) );
  NOR2_X2 U3720 ( .A1(n4819), .A2(n4493), .ZN(n1923) );
  NOR2_X2 U3721 ( .A1(fracta_mul[39]), .A2(fracta_mul[38]), .ZN(n1280) );
  NOR2_X2 U3722 ( .A1(fracta_mul[0]), .A2(n1285), .ZN(n1274) );
  NAND3_X2 U3723 ( .A1(n4593), .A2(n4490), .A3(n4431), .ZN(n1301) );
  NAND3_X2 U3724 ( .A1(n4611), .A2(n4362), .A3(n1371), .ZN(n1281) );
  AOI21_X2 U3725 ( .B1(n4616), .B2(n4488), .A(fracta_mul[19]), .ZN(n1425) );
  NOR2_X2 U3726 ( .A1(fracta_mul[42]), .A2(fracta_mul[43]), .ZN(n1396) );
  NOR2_X2 U3727 ( .A1(fracta_mul[34]), .A2(fracta_mul[33]), .ZN(n1395) );
  NOR2_X2 U3728 ( .A1(n1435), .A2(fracta_mul[27]), .ZN(n1399) );
  NOR2_X2 U3729 ( .A1(n1447), .A2(n1404), .ZN(n1446) );
  AOI21_X2 U3730 ( .B1(fracta_mul[13]), .B2(n4496), .A(fracta_mul[15]), .ZN(
        n1447) );
  NOR2_X2 U3731 ( .A1(n1404), .A2(fracta_mul[15]), .ZN(n1377) );
  NOR2_X2 U3732 ( .A1(fracta_mul[14]), .A2(fracta_mul[13]), .ZN(n1378) );
  NAND3_X2 U3733 ( .A1(fracta_mul[6]), .A2(n6368), .A3(n1361), .ZN(n1393) );
  NAND3_X2 U3734 ( .A1(n4367), .A2(n4356), .A3(n1420), .ZN(n1282) );
  NOR3_X2 U3735 ( .A1(n1283), .A2(fracta_mul[31]), .A3(n6361), .ZN(n1372) );
  NAND3_X2 U3736 ( .A1(n4372), .A2(n4614), .A3(n1395), .ZN(n1283) );
  NAND3_X2 U3737 ( .A1(fracta_mul[29]), .A2(n4612), .A3(n1372), .ZN(n1412) );
  AOI21_X2 U3738 ( .B1(n4613), .B2(fracta_mul[33]), .A(fracta_mul[35]), .ZN(
        n1441) );
  NAND3_X2 U3739 ( .A1(n1735), .A2(n4767), .A3(n4573), .ZN(n246) );
  NAND3_X2 U3740 ( .A1(n6404), .A2(n6407), .A3(n457), .ZN(n1741) );
  NOR2_X2 U3741 ( .A1(n4479), .A2(n2080), .ZN(n2079) );
  OAI21_X2 U3742 ( .B1(fract_denorm[102]), .B2(n6517), .A(n6518), .ZN(n576) );
  NOR2_X2 U3743 ( .A1(fract_denorm[4]), .A2(n390), .ZN(n572) );
  AOI211_X2 U3744 ( .C1(n335), .C2(fract_denorm[19]), .A(n403), .B(n6466), 
        .ZN(n486) );
  AOI21_X2 U3745 ( .B1(n508), .B2(n4874), .A(n362), .ZN(n507) );
  NOR2_X2 U3746 ( .A1(n491), .A2(n492), .ZN(n408) );
  OAI21_X2 U3747 ( .B1(n4873), .B2(n493), .A(n494), .ZN(n492) );
  NAND3_X2 U3748 ( .A1(n6448), .A2(n6447), .A3(fract_denorm[37]), .ZN(n494) );
  NAND3_X2 U3749 ( .A1(n6452), .A2(n544), .A3(fract_denorm[39]), .ZN(n524) );
  OAI21_X2 U3750 ( .B1(n4873), .B2(n6163), .A(n1735), .ZN(n2330) );
  OAI21_X2 U3751 ( .B1(n4430), .B2(n242), .A(n4401), .ZN(n2328) );
  OAI21_X2 U3752 ( .B1(n279), .B2(n4818), .A(n2329), .ZN(n262) );
  AOI21_X2 U3753 ( .B1(n4476), .B2(n4587), .A(n288), .ZN(n2317) );
  NOR2_X2 U3754 ( .A1(n4819), .A2(n4401), .ZN(n1740) );
  OAI21_X2 U3755 ( .B1(n4873), .B2(n6163), .A(n2335), .ZN(n1737) );
  INV_X4 U3756 ( .A(n1745), .ZN(n6390) );
  INV_X4 U3757 ( .A(n4400), .ZN(n4823) );
  NAND3_X2 U3758 ( .A1(fpu_op_r2[2]), .A2(n4505), .A3(fpu_op_r2[0]), .ZN(n1308) );
  NOR2_X2 U3759 ( .A1(n4505), .A2(fpu_op_r2[2]), .ZN(n1314) );
  NOR2_X2 U3760 ( .A1(fpu_op_r2[1]), .A2(fpu_op_r2[2]), .ZN(n1313) );
  NAND2_X2 U3761 ( .A1(fpu_op_r2[1]), .A2(fpu_op_r2[2]), .ZN(n1310) );
  OAI21_X2 U3762 ( .B1(n1622), .B2(n1623), .A(n1624), .ZN(n1521) );
  NAND3_X2 U3763 ( .A1(n1740), .A2(n1741), .A3(n1742), .ZN(n1687) );
  NOR3_X2 U3764 ( .A1(n4481), .A2(opb_00), .A3(fpu_op_r3[2]), .ZN(n1651) );
  NOR2_X2 U3765 ( .A1(fasu_op_r2), .A2(n4626), .ZN(n1485) );
  OAI21_X2 U3766 ( .B1(n1488), .B2(n1489), .A(n1490), .ZN(n1487) );
  NOR2_X2 U3767 ( .A1(n1673), .A2(n4630), .ZN(n1761) );
  NOR2_X2 U3768 ( .A1(n1517), .A2(n1470), .ZN(n1465) );
  NOR2_X2 U3769 ( .A1(opa_inf), .A2(n1480), .ZN(n1476) );
  NOR2_X2 U3770 ( .A1(snan_d), .A2(qnan_d), .ZN(n1468) );
  NOR2_X2 U3771 ( .A1(n1470), .A2(n1745), .ZN(n1467) );
  AOI211_X2 U3772 ( .C1(n1696), .C2(n6389), .A(n1682), .B(n1744), .ZN(n1659)
         );
  OAI21_X2 U3773 ( .B1(n1477), .B2(n1671), .A(n1663), .ZN(n1669) );
  NOR3_X2 U3774 ( .A1(n1522), .A2(n1656), .A3(n1675), .ZN(n1663) );
  OAI21_X2 U3775 ( .B1(n1676), .B2(n244), .A(n1677), .ZN(n1656) );
  NOR3_X2 U3776 ( .A1(n1680), .A2(n1681), .A3(n1682), .ZN(n1676) );
  OAI21_X2 U3777 ( .B1(n1678), .B2(n1679), .A(n4821), .ZN(n1677) );
  OAI21_X2 U3778 ( .B1(n1683), .B2(n1684), .A(n1685), .ZN(n1680) );
  OAI21_X2 U3779 ( .B1(n1955), .B2(n1952), .A(n1953), .ZN(n1954) );
  OAI21_X2 U3780 ( .B1(n1968), .B2(n1971), .A(n1963), .ZN(n1634) );
  OAI21_X2 U3781 ( .B1(n1968), .B2(n1970), .A(n1963), .ZN(n1633) );
  OAI21_X2 U3782 ( .B1(n1968), .B2(n1969), .A(n1963), .ZN(n1635) );
  AOI21_X2 U3783 ( .B1(n1927), .B2(inf_d), .A(n1928), .ZN(n1926) );
  NOR2_X2 U3784 ( .A1(n4822), .A2(n6390), .ZN(n1927) );
  NOR2_X2 U3785 ( .A1(n4123), .A2(u2_exp_ovf_d_1_), .ZN(n616) );
  NOR3_X2 U3786 ( .A1(n4815), .A2(n6352), .A3(n608), .ZN(n615) );
  NAND3_X2 U3787 ( .A1(n4815), .A2(n6099), .A3(u2_N18), .ZN(n595) );
  NAND3_X2 U3788 ( .A1(u2_N12), .A2(u2_N11), .A3(u2_N13), .ZN(n588) );
  NAND3_X2 U3789 ( .A1(u2_N15), .A2(u2_N14), .A3(u2_N6), .ZN(n591) );
  OAI22_X2 U3790 ( .A1(n4815), .A2(n6084), .B1(n4817), .B2(n6099), .ZN(
        u2_exp_tmp4_10_) );
  NOR3_X2 U3791 ( .A1(opa_r1[54]), .A2(opa_r1[56]), .A3(opa_r1[55]), .ZN(n2653) );
  NAND3_X2 U3792 ( .A1(n4623), .A2(n4508), .A3(n4433), .ZN(n2655) );
  OAI21_X2 U3793 ( .B1(u1_sticky), .B2(u1_adj_op_out_sft_0_), .A(n4829), .ZN(
        n754) );
  OAI21_X2 U3794 ( .B1(u1_sticky), .B2(u1_adj_op_out_sft_0_), .A(n4839), .ZN(
        n755) );
  INV_X4 U3795 ( .A(n4865), .ZN(n4859) );
  INV_X4 U3796 ( .A(n4865), .ZN(n4860) );
  INV_X4 U3797 ( .A(n4865), .ZN(n4861) );
  AOI222_X1 U3798 ( .A1(n6287), .A2(n909), .B1(n852), .B2(n910), .C1(n6296), 
        .C2(n911), .ZN(n892) );
  AOI222_X1 U3799 ( .A1(n6291), .A2(n823), .B1(n6288), .B2(n825), .C1(n6289), 
        .C2(n827), .ZN(n821) );
  AOI21_X2 U3800 ( .B1(n6298), .B2(n815), .A(n816), .ZN(n813) );
  AOI222_X1 U3801 ( .A1(n6292), .A2(n844), .B1(n6291), .B2(n845), .C1(n6290), 
        .C2(n847), .ZN(n830) );
  AOI222_X1 U3802 ( .A1(n6296), .A2(n849), .B1(n6299), .B2(n851), .C1(n852), 
        .C2(n853), .ZN(n829) );
  AOI211_X2 U3803 ( .C1(n6297), .C2(n833), .A(n834), .B(n835), .ZN(n831) );
  AOI21_X2 U3804 ( .B1(n836), .B2(n6349), .A(n838), .ZN(n835) );
  NOR3_X2 U3805 ( .A1(n868), .A2(n852), .A3(n6296), .ZN(n934) );
  NOR3_X2 U3806 ( .A1(n4628), .A2(u1_fracta_lt_fractb), .A3(
        u1_fracta_eq_fractb), .ZN(n793) );
  NOR3_X2 U3807 ( .A1(n4585), .A2(n4583), .A3(n4584), .ZN(n950) );
  NAND3_X2 U3808 ( .A1(opa_r[59]), .A2(opa_r[62]), .A3(opa_r[58]), .ZN(n952)
         );
  NOR3_X2 U3809 ( .A1(n4371), .A2(n4590), .A3(n4360), .ZN(n1085) );
  NAND3_X2 U3810 ( .A1(opb_r[59]), .A2(opb_r[62]), .A3(opb_r[58]), .ZN(n1087)
         );
  NOR3_X2 U3811 ( .A1(opa_r[54]), .A2(opa_r[56]), .A3(opa_r[55]), .ZN(n1305)
         );
  NAND3_X2 U3812 ( .A1(n4575), .A2(n4582), .A3(n4586), .ZN(n1307) );
  NOR3_X2 U3813 ( .A1(fracta_mul[20]), .A2(fracta_mul[28]), .A3(fracta_mul[21]), .ZN(n1275) );
  NOR3_X2 U3814 ( .A1(n1298), .A2(n1299), .A3(n1300), .ZN(n1288) );
  NOR2_X2 U3815 ( .A1(n1413), .A2(n1281), .ZN(n1369) );
  NAND3_X2 U3816 ( .A1(fracta_mul[41]), .A2(n1396), .A3(n1369), .ZN(n1427) );
  OAI21_X2 U3817 ( .B1(n1436), .B2(n6358), .A(n1426), .ZN(n1433) );
  NOR2_X2 U3818 ( .A1(fracta_mul[46]), .A2(fracta_mul[45]), .ZN(n1371) );
  NOR2_X2 U3819 ( .A1(fracta_mul[1]), .A2(fracta_mul[2]), .ZN(n1421) );
  AOI21_X2 U3820 ( .B1(n1377), .B2(n6370), .A(n1425), .ZN(n1423) );
  NAND3_X2 U3821 ( .A1(n6369), .A2(n4495), .A3(fracta_mul[10]), .ZN(n1422) );
  AOI211_X2 U3822 ( .C1(fracta_mul[26]), .C2(n1399), .A(n1390), .B(n1419), 
        .ZN(n1418) );
  NAND3_X2 U3823 ( .A1(n1392), .A2(n1393), .A3(n1394), .ZN(n1388) );
  NOR3_X2 U3824 ( .A1(fracta_mul[50]), .A2(fracta_mul[51]), .A3(fracta_mul[49]), .ZN(n1398) );
  OAI21_X2 U3825 ( .B1(fracta_mul[46]), .B2(n4499), .A(n4362), .ZN(n1445) );
  NAND3_X2 U3826 ( .A1(n1378), .A2(n4491), .A3(n1377), .ZN(n1375) );
  NOR2_X2 U3827 ( .A1(fracta_mul[10]), .A2(fracta_mul[11]), .ZN(n1374) );
  NAND3_X2 U3828 ( .A1(n6369), .A2(n4492), .A3(fracta_mul[8]), .ZN(n1376) );
  NAND3_X2 U3829 ( .A1(fracta_mul[7]), .A2(n6369), .A3(n1361), .ZN(n1449) );
  NOR3_X2 U3830 ( .A1(n1282), .A2(fracta_mul[20]), .A3(n1435), .ZN(n1361) );
  NAND3_X2 U3831 ( .A1(n1365), .A2(n1366), .A3(n1367), .ZN(n1364) );
  OAI21_X2 U3832 ( .B1(fracta_mul[40]), .B2(n6365), .A(n1369), .ZN(n1367) );
  AOI211_X2 U3833 ( .C1(fracta_mul[37]), .C2(n6355), .A(n1454), .B(n1350), 
        .ZN(n1379) );
  NOR3_X2 U3834 ( .A1(n4498), .A2(n1442), .A3(n6358), .ZN(n1454) );
  NOR3_X2 U3835 ( .A1(n1442), .A2(fracta_mul[5]), .A3(n6358), .ZN(n1351) );
  NOR3_X2 U3836 ( .A1(n4377), .A2(n1282), .A3(n1435), .ZN(n1350) );
  NOR3_X2 U3837 ( .A1(n1354), .A2(fracta_mul[37]), .A3(n4365), .ZN(n1353) );
  NOR3_X2 U3838 ( .A1(fracta_mul[36]), .A2(fracta_mul[37]), .A3(n1354), .ZN(
        n1355) );
  NAND3_X2 U3839 ( .A1(fracta_mul[31]), .A2(n6366), .A3(n1355), .ZN(n1451) );
  AOI211_X2 U3840 ( .C1(n1351), .C2(n1438), .A(n1439), .B(n1440), .ZN(n1346)
         );
  NOR2_X2 U3841 ( .A1(n4500), .A2(fracta_mul[4]), .ZN(n1438) );
  NOR3_X2 U3842 ( .A1(n1381), .A2(n1382), .A3(n6356), .ZN(n1347) );
  INV_X4 U3843 ( .A(n241), .ZN(n6387) );
  NOR3_X2 U3844 ( .A1(n4821), .A2(n6391), .A3(n246), .ZN(n212) );
  NOR2_X2 U3845 ( .A1(n4821), .A2(n247), .ZN(n211) );
  NOR4_X2 U3846 ( .A1(opb_dn), .A2(n4426), .A3(u4_N6159), .A4(u4_N6158), .ZN(
        n2075) );
  NOR2_X2 U3847 ( .A1(n4767), .A2(n6401), .ZN(n2076) );
  NOR3_X2 U3848 ( .A1(n4574), .A2(n1925), .A3(n1741), .ZN(n2102) );
  AOI211_X2 U3849 ( .C1(n572), .C2(fract_denorm[3]), .A(n573), .B(n4873), .ZN(
        n488) );
  NOR2_X2 U3850 ( .A1(n2097), .A2(n1739), .ZN(n2093) );
  AOI21_X2 U3851 ( .B1(n6390), .B2(n2316), .A(n2317), .ZN(n2315) );
  OAI21_X2 U3852 ( .B1(u4_div_scht1a[10]), .B2(u4_div_scht1a[9]), .A(n255), 
        .ZN(n2314) );
  OAI21_X2 U3853 ( .B1(u4_exp_in_pl1_10_), .B2(u4_exp_in_pl1_9_), .A(n262), 
        .ZN(n2313) );
  NOR3_X2 U3854 ( .A1(n6389), .A2(n4822), .A3(n6390), .ZN(n2143) );
  NAND3_X2 U3855 ( .A1(n2051), .A2(n4579), .A3(n1740), .ZN(n2142) );
  NOR2_X2 U3856 ( .A1(n1925), .A2(n6403), .ZN(n2088) );
  NOR2_X2 U3857 ( .A1(n2097), .A2(n6161), .ZN(n2073) );
  NOR3_X2 U3858 ( .A1(n1755), .A2(n6377), .A3(n1745), .ZN(n2072) );
  NAND2_X2 U3859 ( .A1(n6401), .A2(n4821), .ZN(n206) );
  NOR2_X2 U3860 ( .A1(n1651), .A2(n4774), .ZN(n1519) );
  OAI21_X2 U3861 ( .B1(fpu_op_r3[2]), .B2(n1481), .A(n1482), .ZN(N911) );
  OAI21_X2 U3862 ( .B1(n1467), .B2(n1756), .A(n1757), .ZN(N880) );
  NAND3_X2 U3863 ( .A1(n4621), .A2(n4504), .A3(n1666), .ZN(n1661) );
  OAI21_X2 U3864 ( .B1(n1663), .B2(n1473), .A(n1667), .ZN(n1666) );
  NOR2_X2 U3865 ( .A1(n1793), .A2(n4800), .ZN(N799) );
  NOR2_X2 U3866 ( .A1(n1794), .A2(n4800), .ZN(N800) );
  NOR2_X2 U3867 ( .A1(n1795), .A2(n4800), .ZN(N801) );
  NOR2_X2 U3868 ( .A1(n1796), .A2(n4802), .ZN(N802) );
  NOR2_X2 U3869 ( .A1(n1797), .A2(n4800), .ZN(N803) );
  NOR2_X2 U3870 ( .A1(n1641), .A2(n4802), .ZN(N804) );
  NOR2_X2 U3871 ( .A1(n1501), .A2(n4800), .ZN(N805) );
  NOR2_X2 U3872 ( .A1(n1499), .A2(n4802), .ZN(N806) );
  NOR2_X2 U3873 ( .A1(n1500), .A2(n4800), .ZN(N807) );
  NOR2_X2 U3874 ( .A1(n1502), .A2(n4802), .ZN(N808) );
  NOR2_X2 U3875 ( .A1(n1503), .A2(n4802), .ZN(N809) );
  NOR2_X2 U3876 ( .A1(n1784), .A2(n4802), .ZN(N811) );
  NOR2_X2 U3877 ( .A1(n1782), .A2(n4802), .ZN(N812) );
  NOR2_X2 U3878 ( .A1(n1783), .A2(n4802), .ZN(N813) );
  NOR2_X2 U3879 ( .A1(n1649), .A2(n4802), .ZN(N819) );
  NOR2_X2 U3880 ( .A1(n1512), .A2(n4802), .ZN(N820) );
  NOR2_X2 U3881 ( .A1(n1510), .A2(n4802), .ZN(N821) );
  NOR2_X2 U3882 ( .A1(n1511), .A2(n4802), .ZN(N822) );
  NOR2_X2 U3883 ( .A1(n1835), .A2(n4802), .ZN(N823) );
  NOR2_X2 U3884 ( .A1(n1834), .A2(n4802), .ZN(N827) );
  NOR2_X2 U3885 ( .A1(n1832), .A2(n4802), .ZN(N828) );
  NOR2_X2 U3886 ( .A1(n1833), .A2(n4800), .ZN(N829) );
  NOR2_X2 U3887 ( .A1(n1824), .A2(n4800), .ZN(N833) );
  NOR2_X2 U3888 ( .A1(n1825), .A2(n4800), .ZN(N834) );
  NOR2_X2 U3889 ( .A1(n1826), .A2(n4800), .ZN(N835) );
  NOR2_X2 U3890 ( .A1(n1827), .A2(n4800), .ZN(N836) );
  NOR2_X2 U3891 ( .A1(n1819), .A2(n4800), .ZN(N840) );
  NOR2_X2 U3892 ( .A1(n1817), .A2(n4800), .ZN(N841) );
  NOR2_X2 U3893 ( .A1(n1818), .A2(n4800), .ZN(N842) );
  NOR2_X2 U3894 ( .A1(n1809), .A2(n4800), .ZN(N846) );
  NOR2_X2 U3895 ( .A1(n1810), .A2(n4800), .ZN(N847) );
  NOR2_X2 U3896 ( .A1(n1811), .A2(n4800), .ZN(N848) );
  NOR2_X2 U3897 ( .A1(n1812), .A2(n4800), .ZN(N849) );
  AOI21_X2 U3898 ( .B1(n1653), .B2(n1654), .A(n1517), .ZN(N904) );
  OAI21_X2 U3899 ( .B1(n1655), .B2(n4772), .A(n1656), .ZN(n1654) );
  AOI21_X2 U3900 ( .B1(opb_00), .B2(fpu_op_r3[0]), .A(fpu_op_r3[2]), .ZN(n1655) );
  AOI222_X1 U3901 ( .A1(fract_i2f[105]), .A2(n4775), .B1(quo[55]), .B2(n4786), 
        .C1(fract_out_q[56]), .C2(n4772), .ZN(n2341) );
  AOI222_X1 U3902 ( .A1(fract_i2f[102]), .A2(n4776), .B1(quo[52]), .B2(n2342), 
        .C1(fract_out_q[53]), .C2(n4772), .ZN(n2348) );
  AOI222_X1 U3903 ( .A1(fract_i2f[101]), .A2(n4776), .B1(quo[51]), .B2(n2342), 
        .C1(fract_out_q[52]), .C2(n4773), .ZN(n2351) );
  AOI222_X1 U3904 ( .A1(fract_i2f[100]), .A2(n4775), .B1(n2342), .B2(quo[50]), 
        .C1(fract_out_q[51]), .C2(n4772), .ZN(n2354) );
  AOI222_X1 U3905 ( .A1(fract_i2f[99]), .A2(n4776), .B1(n4786), .B2(quo[49]), 
        .C1(fract_out_q[50]), .C2(n4773), .ZN(n2356) );
  AOI222_X1 U3906 ( .A1(fract_i2f[98]), .A2(n4775), .B1(n2342), .B2(quo[48]), 
        .C1(fract_out_q[49]), .C2(n4772), .ZN(n2359) );
  AOI222_X1 U3907 ( .A1(fract_i2f[97]), .A2(n4775), .B1(quo[47]), .B2(n4786), 
        .C1(fract_out_q[48]), .C2(n4773), .ZN(n2361) );
  AOI222_X1 U3908 ( .A1(fract_i2f[96]), .A2(n4776), .B1(quo[46]), .B2(n2342), 
        .C1(fract_out_q[47]), .C2(n4774), .ZN(n2364) );
  AOI222_X1 U3909 ( .A1(fract_i2f[95]), .A2(n4778), .B1(quo[45]), .B2(n2342), 
        .C1(fract_out_q[46]), .C2(n4773), .ZN(n2367) );
  AOI222_X1 U3910 ( .A1(fract_i2f[94]), .A2(n4775), .B1(quo[44]), .B2(n4787), 
        .C1(fract_out_q[45]), .C2(n4772), .ZN(n2370) );
  AOI222_X1 U3911 ( .A1(fract_i2f[93]), .A2(n4775), .B1(n4787), .B2(quo[43]), 
        .C1(fract_out_q[44]), .C2(n4773), .ZN(n2372) );
  AOI222_X1 U3912 ( .A1(fract_i2f[92]), .A2(n4776), .B1(n4786), .B2(quo[42]), 
        .C1(fract_out_q[43]), .C2(n4774), .ZN(n2374) );
  AOI222_X1 U3913 ( .A1(fract_i2f[91]), .A2(n4775), .B1(quo[41]), .B2(n4787), 
        .C1(fract_out_q[42]), .C2(n4772), .ZN(n2376) );
  AOI222_X1 U3914 ( .A1(fract_i2f[90]), .A2(n4778), .B1(quo[40]), .B2(n4787), 
        .C1(fract_out_q[41]), .C2(n4773), .ZN(n2378) );
  AOI222_X1 U3915 ( .A1(fract_i2f[89]), .A2(n4777), .B1(quo[39]), .B2(n2342), 
        .C1(fract_out_q[40]), .C2(n4774), .ZN(n2381) );
  AOI222_X1 U3916 ( .A1(fract_i2f[88]), .A2(n4775), .B1(quo[38]), .B2(n4787), 
        .C1(fract_out_q[39]), .C2(n4772), .ZN(n2384) );
  AOI222_X1 U3917 ( .A1(fract_i2f[87]), .A2(n4776), .B1(n4786), .B2(quo[37]), 
        .C1(fract_out_q[38]), .C2(n4773), .ZN(n2386) );
  AOI222_X1 U3918 ( .A1(fract_i2f[86]), .A2(n4775), .B1(n4787), .B2(quo[36]), 
        .C1(fract_out_q[37]), .C2(n4774), .ZN(n2388) );
  AOI222_X1 U3919 ( .A1(fract_i2f[85]), .A2(n4776), .B1(n4786), .B2(quo[35]), 
        .C1(fract_out_q[36]), .C2(n4774), .ZN(n2390) );
  AOI222_X1 U3920 ( .A1(fract_i2f[84]), .A2(n4776), .B1(quo[34]), .B2(n4787), 
        .C1(fract_out_q[35]), .C2(n4774), .ZN(n2392) );
  AOI222_X1 U3921 ( .A1(fract_i2f[83]), .A2(n4777), .B1(quo[33]), .B2(n4787), 
        .C1(fract_out_q[34]), .C2(n4774), .ZN(n2395) );
  AOI222_X1 U3922 ( .A1(fract_i2f[82]), .A2(n4776), .B1(quo[32]), .B2(n4787), 
        .C1(fract_out_q[33]), .C2(n4774), .ZN(n2398) );
  AOI222_X1 U3923 ( .A1(fract_i2f[81]), .A2(n4775), .B1(n4787), .B2(quo[31]), 
        .C1(fract_out_q[32]), .C2(n4774), .ZN(n2401) );
  AOI222_X1 U3924 ( .A1(fract_i2f[80]), .A2(n4777), .B1(n4787), .B2(quo[30]), 
        .C1(fract_out_q[31]), .C2(n4774), .ZN(n2403) );
  AOI222_X1 U3925 ( .A1(fract_i2f[79]), .A2(n4776), .B1(quo[29]), .B2(n4787), 
        .C1(fract_out_q[30]), .C2(n4774), .ZN(n2405) );
  AOI222_X1 U3926 ( .A1(fract_i2f[78]), .A2(n4777), .B1(quo[28]), .B2(n4787), 
        .C1(fract_out_q[29]), .C2(n4774), .ZN(n2408) );
  AOI222_X1 U3927 ( .A1(fract_i2f[77]), .A2(n4776), .B1(quo[27]), .B2(n4787), 
        .C1(fract_out_q[28]), .C2(n4774), .ZN(n2411) );
  AOI222_X1 U3928 ( .A1(fract_i2f[76]), .A2(n4776), .B1(quo[26]), .B2(n4787), 
        .C1(fract_out_q[27]), .C2(n4774), .ZN(n2414) );
  AOI222_X1 U3929 ( .A1(fract_i2f[75]), .A2(n4777), .B1(n2342), .B2(quo[25]), 
        .C1(fract_out_q[26]), .C2(n4774), .ZN(n2416) );
  AOI222_X1 U3930 ( .A1(fract_i2f[74]), .A2(n4777), .B1(n2342), .B2(quo[24]), 
        .C1(fract_out_q[25]), .C2(n4773), .ZN(n2418) );
  AOI222_X1 U3931 ( .A1(fract_i2f[73]), .A2(n4776), .B1(n4786), .B2(quo[23]), 
        .C1(fract_out_q[24]), .C2(n4773), .ZN(n2420) );
  AOI222_X1 U3932 ( .A1(fract_i2f[72]), .A2(n4777), .B1(quo[22]), .B2(n4786), 
        .C1(fract_out_q[23]), .C2(n4773), .ZN(n2422) );
  AOI222_X1 U3933 ( .A1(fract_i2f[71]), .A2(n4777), .B1(quo[21]), .B2(n4786), 
        .C1(fract_out_q[22]), .C2(n4773), .ZN(n2425) );
  AOI222_X1 U3934 ( .A1(fract_i2f[70]), .A2(n4775), .B1(n4786), .B2(quo[20]), 
        .C1(fract_out_q[21]), .C2(n4773), .ZN(n2428) );
  AOI222_X1 U3935 ( .A1(fract_i2f[69]), .A2(n4777), .B1(n4787), .B2(quo[19]), 
        .C1(fract_out_q[20]), .C2(n4773), .ZN(n2430) );
  AOI222_X1 U3936 ( .A1(fract_i2f[68]), .A2(n4777), .B1(n2342), .B2(quo[18]), 
        .C1(fract_out_q[19]), .C2(n4773), .ZN(n2432) );
  AOI222_X1 U3937 ( .A1(fract_i2f[67]), .A2(n4777), .B1(quo[17]), .B2(n4786), 
        .C1(fract_out_q[18]), .C2(n4773), .ZN(n2434) );
  AOI222_X1 U3938 ( .A1(fract_i2f[66]), .A2(n4777), .B1(quo[16]), .B2(n4786), 
        .C1(fract_out_q[17]), .C2(n4773), .ZN(n2437) );
  AOI222_X1 U3939 ( .A1(fract_i2f[65]), .A2(n4775), .B1(quo[15]), .B2(n4786), 
        .C1(fract_out_q[16]), .C2(n4773), .ZN(n2440) );
  AOI222_X1 U3940 ( .A1(fract_i2f[64]), .A2(n4775), .B1(quo[14]), .B2(n4786), 
        .C1(fract_out_q[15]), .C2(n4773), .ZN(n2443) );
  AOI222_X1 U3941 ( .A1(fract_i2f[63]), .A2(n4778), .B1(n4787), .B2(quo[13]), 
        .C1(fract_out_q[14]), .C2(n4774), .ZN(n2445) );
  AOI222_X1 U3942 ( .A1(fract_i2f[62]), .A2(n4775), .B1(n2342), .B2(quo[12]), 
        .C1(fract_out_q[13]), .C2(n4773), .ZN(n2447) );
  AOI222_X1 U3943 ( .A1(fract_i2f[61]), .A2(n4775), .B1(quo[11]), .B2(n4786), 
        .C1(fract_out_q[12]), .C2(n4772), .ZN(n2449) );
  AOI222_X1 U3944 ( .A1(fract_i2f[60]), .A2(n4776), .B1(n4787), .B2(quo[10]), 
        .C1(fract_out_q[11]), .C2(n4772), .ZN(n2451) );
  AOI222_X1 U3945 ( .A1(fract_i2f[59]), .A2(n4777), .B1(quo[9]), .B2(n4786), 
        .C1(fract_out_q[10]), .C2(n4772), .ZN(n2454) );
  AOI222_X1 U3946 ( .A1(fract_i2f[58]), .A2(n4776), .B1(n4786), .B2(quo[8]), 
        .C1(fract_out_q[9]), .C2(n4772), .ZN(n2457) );
  AOI222_X1 U3947 ( .A1(fract_i2f[57]), .A2(n4775), .B1(n2342), .B2(quo[7]), 
        .C1(fract_out_q[8]), .C2(n4772), .ZN(n2459) );
  AOI222_X1 U3948 ( .A1(fract_i2f[56]), .A2(n4777), .B1(quo[6]), .B2(n4786), 
        .C1(fract_out_q[7]), .C2(n4772), .ZN(n2461) );
  AOI222_X1 U3949 ( .A1(fract_i2f[55]), .A2(n4777), .B1(n2342), .B2(quo[5]), 
        .C1(fract_out_q[6]), .C2(n4772), .ZN(n2463) );
  AOI222_X1 U3950 ( .A1(fract_i2f[54]), .A2(n4776), .B1(n2342), .B2(quo[4]), 
        .C1(fract_out_q[5]), .C2(n4772), .ZN(n2466) );
  AOI222_X1 U3951 ( .A1(fract_i2f[53]), .A2(n4777), .B1(quo[3]), .B2(n4786), 
        .C1(fract_out_q[4]), .C2(n4772), .ZN(n2469) );
  AOI222_X1 U3952 ( .A1(fract_i2f[52]), .A2(n4777), .B1(n2342), .B2(quo[2]), 
        .C1(fract_out_q[3]), .C2(n4772), .ZN(n2472) );
  AOI222_X1 U3953 ( .A1(fract_i2f[51]), .A2(n4775), .B1(quo[1]), .B2(n4786), 
        .C1(fract_out_q[2]), .C2(n4772), .ZN(n2474) );
  AOI222_X1 U3954 ( .A1(fract_i2f[50]), .A2(n4776), .B1(quo[0]), .B2(n4787), 
        .C1(fract_out_q[1]), .C2(n4772), .ZN(n2476) );
  NOR3_X2 U3955 ( .A1(opb_r[54]), .A2(opb_r[56]), .A3(opb_r[55]), .ZN(n1271)
         );
  NAND3_X2 U3956 ( .A1(n4471), .A2(n4569), .A3(n4398), .ZN(n1273) );
  NAND3_X2 U3957 ( .A1(exp_mul[2]), .A2(exp_mul[3]), .A3(exp_mul[1]), .ZN(
        n1457) );
  AOI222_X1 U3958 ( .A1(u2_N75), .A2(n612), .B1(u2_exp_tmp4_10_), .B2(n613), 
        .C1(u2_exp_tmp3_10_), .C2(n614), .ZN(n611) );
  AOI222_X1 U3959 ( .A1(u2_N74), .A2(n612), .B1(n1048), .B2(n613), .C1(
        u2_exp_tmp3_9_), .C2(n614), .ZN(n618) );
  AOI222_X1 U3960 ( .A1(u2_N73), .A2(n612), .B1(n1049), .B2(n613), .C1(
        u2_exp_tmp3_8_), .C2(n614), .ZN(n620) );
  AOI222_X1 U3961 ( .A1(u2_N72), .A2(n612), .B1(n1050), .B2(n613), .C1(
        u2_exp_tmp3_7_), .C2(n614), .ZN(n622) );
  AOI222_X1 U3962 ( .A1(u2_N71), .A2(n612), .B1(n1051), .B2(n613), .C1(
        u2_exp_tmp3_6_), .C2(n614), .ZN(n624) );
  AOI222_X1 U3963 ( .A1(u2_N70), .A2(n612), .B1(n1052), .B2(n613), .C1(
        u2_exp_tmp3_5_), .C2(n614), .ZN(n626) );
  AOI222_X1 U3964 ( .A1(u2_N69), .A2(n612), .B1(u2_exp_tmp4_4_), .B2(n613), 
        .C1(u2_exp_tmp3_4_), .C2(n614), .ZN(n628) );
  AOI222_X1 U3965 ( .A1(u2_N68), .A2(n612), .B1(u2_exp_tmp4_3_), .B2(n613), 
        .C1(u2_exp_tmp3_3_), .C2(n614), .ZN(n630) );
  AOI222_X1 U3966 ( .A1(u2_N67), .A2(n612), .B1(u2_exp_tmp4_2_), .B2(n613), 
        .C1(u2_exp_tmp3_2_), .C2(n614), .ZN(n632) );
  AOI222_X1 U3967 ( .A1(u2_N66), .A2(n612), .B1(u2_exp_tmp4_1_), .B2(n613), 
        .C1(u2_exp_tmp3_1_), .C2(n614), .ZN(n634) );
  AOI222_X1 U3968 ( .A1(u2_lt_131_A_0_), .A2(n612), .B1(n1054), .B2(n613), 
        .C1(u2_exp_tmp3_0_), .C2(n614), .ZN(n636) );
  AOI21_X2 U3969 ( .B1(n605), .B2(n606), .A(n4592), .ZN(u2_exp_ovf_d_0_) );
  NOR2_X2 U3970 ( .A1(n581), .A2(n6351), .ZN(u2_underflow_d[2]) );
  OAI21_X2 U3971 ( .B1(opa_r[62]), .B2(opb_r[62]), .A(n583), .ZN(n601) );
  OAI21_X2 U3972 ( .B1(n4815), .B2(n639), .A(n640), .ZN(u2_N114) );
  OAI21_X2 U3973 ( .B1(n4402), .B2(n2532), .A(n2651), .ZN(N608) );
  OAI21_X2 U3974 ( .B1(n4627), .B2(n2532), .A(n2648), .ZN(N609) );
  NOR2_X2 U3975 ( .A1(n777), .A2(n6309), .ZN(u1_N88) );
  NOR2_X2 U3976 ( .A1(n777), .A2(n779), .ZN(u1_N87) );
  NOR2_X2 U3977 ( .A1(n777), .A2(n780), .ZN(u1_N86) );
  NOR2_X2 U3978 ( .A1(n777), .A2(n6314), .ZN(u1_N85) );
  NOR2_X2 U3979 ( .A1(n777), .A2(n6315), .ZN(u1_N84) );
  NOR2_X2 U3980 ( .A1(n777), .A2(n6316), .ZN(u1_N83) );
  NOR2_X2 U3981 ( .A1(n777), .A2(n6317), .ZN(u1_N82) );
  NOR2_X2 U3982 ( .A1(n777), .A2(n6318), .ZN(u1_N81) );
  NOR2_X2 U3983 ( .A1(n777), .A2(n6319), .ZN(u1_N80) );
  NOR2_X2 U3984 ( .A1(n777), .A2(n6320), .ZN(u1_N79) );
  NOR2_X2 U3985 ( .A1(n777), .A2(n6321), .ZN(u1_N78) );
  OAI21_X2 U3986 ( .B1(n807), .B2(n808), .A(u1_exp_diff_sft_0_), .ZN(n806) );
  NOR3_X2 U3987 ( .A1(n6297), .A2(n6298), .A3(n6289), .ZN(n935) );
  NOR3_X2 U3988 ( .A1(n6290), .A2(n6291), .A3(n6299), .ZN(n936) );
  OAI21_X2 U3989 ( .B1(n790), .B2(n4624), .A(n792), .ZN(u1_N334) );
  AOI21_X2 U3990 ( .B1(opb_nan), .B2(n796), .A(u1_signa_r), .ZN(n790) );
  OAI21_X2 U3991 ( .B1(n793), .B2(n4633), .A(u1_signa_r), .ZN(n792) );
  OAI21_X2 U3992 ( .B1(u1_fracta_eq_fractb), .B2(n4632), .A(opa_nan), .ZN(n796) );
  AOI21_X2 U3993 ( .B1(u1_signa_r), .B2(n799), .A(n6375), .ZN(n798) );
  NOR2_X2 U3994 ( .A1(fpu_op_r3[2]), .A2(n6383), .ZN(N909) );
  NOR2_X2 U3995 ( .A1(n944), .A2(n943), .ZN(u0_N6) );
  NOR2_X2 U3996 ( .A1(fracta_mul[51]), .A2(n947), .ZN(u0_N4) );
  NOR2_X2 U3997 ( .A1(n4349), .A2(n949), .ZN(u0_N10) );
  NOR2_X2 U3998 ( .A1(n4350), .A2(n948), .ZN(u0_N11) );
  NOR2_X2 U3999 ( .A1(n946), .A2(u6_N51), .ZN(n4350) );
  NOR3_X2 U4000 ( .A1(n1413), .A2(fracta_mul[47]), .A3(n1371), .ZN(n1410) );
  AOI222_X1 U4001 ( .A1(n1361), .A2(n1397), .B1(n1398), .B2(fracta_mul[48]), 
        .C1(n1381), .C2(n4615), .ZN(n1386) );
  AOI21_X2 U4002 ( .B1(n1355), .B2(n1356), .A(n1357), .ZN(n1348) );
  NAND3_X2 U4003 ( .A1(n4372), .A2(n4613), .A3(n4363), .ZN(n1356) );
  OAI21_X2 U4004 ( .B1(n2081), .B2(n244), .A(n2082), .ZN(u4_exp_out_9_) );
  OAI21_X2 U4005 ( .B1(n1715), .B2(n244), .A(n2086), .ZN(u4_exp_out_10_) );
  AOI21_X2 U4006 ( .B1(n2095), .B2(n2096), .A(n244), .ZN(n2094) );
  NOR3_X2 U4007 ( .A1(u4_N5926), .A2(u4_N5928), .A3(u4_N5927), .ZN(n2284) );
  NOR3_X2 U4008 ( .A1(u4_N5929), .A2(u4_N5931), .A3(u4_N5930), .ZN(n2285) );
  NOR3_X2 U4009 ( .A1(u4_N5932), .A2(u4_N5934), .A3(u4_N5933), .ZN(n2286) );
  NOR3_X2 U4010 ( .A1(u4_N5913), .A2(u4_N5915), .A3(u4_N5914), .ZN(n2280) );
  NOR3_X2 U4011 ( .A1(u4_N5916), .A2(u4_N5918), .A3(u4_N5917), .ZN(n2281) );
  NOR3_X2 U4012 ( .A1(u4_N5919), .A2(u4_N5921), .A3(u4_N5920), .ZN(n2282) );
  NOR3_X2 U4013 ( .A1(u4_N5900), .A2(u4_N5902), .A3(u4_N5901), .ZN(n2276) );
  NOR3_X2 U4014 ( .A1(u4_N5903), .A2(u4_N5905), .A3(u4_N5904), .ZN(n2277) );
  NOR3_X2 U4015 ( .A1(u4_N5906), .A2(u4_N5908), .A3(u4_N5907), .ZN(n2278) );
  INV_X8 U4016 ( .A(n4838), .ZN(n4829) );
  INV_X4 U4017 ( .A(n4836), .ZN(n4832) );
  INV_X4 U4018 ( .A(n4858), .ZN(n4854) );
  INV_X4 U4019 ( .A(n4858), .ZN(n4855) );
  INV_X4 U4020 ( .A(n4850), .ZN(n4847) );
  INV_X4 U4021 ( .A(n4848), .ZN(n4839) );
  INV_X4 U4022 ( .A(n4879), .ZN(n4878) );
  NAND2_X2 U4023 ( .A1(n1933), .A2(n1940), .ZN(n4357) );
  NAND2_X2 U4024 ( .A1(n1933), .A2(n1943), .ZN(n4358) );
  OR2_X4 U4025 ( .A1(u4_N5898), .A2(n2312), .ZN(n4361) );
  INV_X4 U4026 ( .A(n4866), .ZN(n4858) );
  INV_X4 U4027 ( .A(n4858), .ZN(n4853) );
  INV_X4 U4028 ( .A(n4862), .ZN(n4856) );
  INV_X4 U4029 ( .A(n4863), .ZN(n4857) );
  INV_X4 U4030 ( .A(n4848), .ZN(n4838) );
  INV_X4 U4031 ( .A(n4358), .ZN(n4796) );
  INV_X4 U4032 ( .A(n4361), .ZN(n4789) );
  INV_X4 U4033 ( .A(n4868), .ZN(n4865) );
  NOR2_X2 U4034 ( .A1(n6082), .A2(n4123), .ZN(n613) );
  INV_X4 U4035 ( .A(n4805), .ZN(n4806) );
  INV_X4 U4036 ( .A(n4871), .ZN(n4872) );
  NAND2_X2 U4037 ( .A1(n1931), .A2(n1932), .ZN(n4383) );
  INV_X4 U4038 ( .A(n4851), .ZN(n4845) );
  INV_X4 U4039 ( .A(n4846), .ZN(n4843) );
  NOR2_X2 U4040 ( .A1(n2337), .A2(n6381), .ZN(n4384) );
  INV_X4 U4041 ( .A(n4814), .ZN(n4813) );
  INV_X4 U4042 ( .A(u1_fractb_lt_fracta), .ZN(n4852) );
  INV_X4 U4043 ( .A(n4849), .ZN(n4836) );
  INV_X4 U4044 ( .A(n2533), .ZN(n4781) );
  INV_X4 U4045 ( .A(n4781), .ZN(n4780) );
  INV_X4 U4046 ( .A(n4781), .ZN(n4779) );
  NOR3_X2 U4047 ( .A1(n6352), .A2(n4816), .A3(n6082), .ZN(n612) );
  INV_X4 U4048 ( .A(n4785), .ZN(n4786) );
  INV_X4 U4049 ( .A(n4785), .ZN(n4787) );
  INV_X4 U4050 ( .A(n2357), .ZN(n4777) );
  INV_X4 U4051 ( .A(n1138), .ZN(n4805) );
  INV_X4 U4052 ( .A(N784), .ZN(n4871) );
  INV_X4 U4053 ( .A(n4383), .ZN(n4798) );
  AND2_X4 U4054 ( .A1(n4426), .A2(n4479), .ZN(n4429) );
  NOR2_X2 U4055 ( .A1(n4479), .A2(n4426), .ZN(n2080) );
  INV_X4 U4056 ( .A(n4852), .ZN(n4866) );
  INV_X4 U4057 ( .A(u2_N157), .ZN(n4824) );
  INV_X8 U4058 ( .A(n4826), .ZN(n4825) );
  INV_X4 U4059 ( .A(u2_N157), .ZN(n4826) );
  NOR3_X2 U4060 ( .A1(n2033), .A2(u4_N6188), .A3(n2049), .ZN(n1992) );
  INV_X4 U4061 ( .A(n4851), .ZN(n4846) );
  INV_X4 U4062 ( .A(n4846), .ZN(n4842) );
  NOR2_X2 U4063 ( .A1(n6352), .A2(u2_exp_ovf_d_1_), .ZN(n614) );
  INV_X4 U4064 ( .A(n4801), .ZN(n4800) );
  INV_X4 U4065 ( .A(n4503), .ZN(n4816) );
  INV_X4 U4066 ( .A(n4816), .ZN(n4815) );
  INV_X4 U4067 ( .A(n4783), .ZN(n4784) );
  NOR2_X2 U4068 ( .A1(n1308), .A2(n2337), .ZN(n1090) );
  INV_X4 U4069 ( .A(n4384), .ZN(n4768) );
  INV_X4 U4070 ( .A(n4384), .ZN(n4769) );
  INV_X4 U4071 ( .A(n4820), .ZN(n4818) );
  INV_X4 U4072 ( .A(n4820), .ZN(n4819) );
  NAND3_X2 U4073 ( .A1(n487), .A2(n488), .A3(n489), .ZN(u4_fi_ldz_2a_0_) );
  INV_X4 U4074 ( .A(fract_denorm[105]), .ZN(n4874) );
  INV_X4 U4075 ( .A(n4874), .ZN(n4873) );
  INV_X4 U4076 ( .A(n4805), .ZN(n4803) );
  INV_X4 U4077 ( .A(n4871), .ZN(n4869) );
  INV_X4 U4078 ( .A(n244), .ZN(n4822) );
  OR2_X4 U4079 ( .A1(n4941), .A2(u4_exp_out_4_), .ZN(n4472) );
  OAI21_X2 U4080 ( .B1(n2069), .B2(n4821), .A(n2071), .ZN(u4_exp_out_8_) );
  OR2_X4 U4081 ( .A1(n4909), .A2(n4382), .ZN(n4478) );
  NOR2_X2 U4082 ( .A1(u4_fi_ldz_2a_6_), .A2(
        sub_1_root_sub_0_root_u4_add_495_carry[7]), .ZN(n4480) );
  INV_X4 U4083 ( .A(n4792), .ZN(n4791) );
  NAND3_X2 U4084 ( .A1(n4481), .A2(n4351), .A3(fpu_op_r3[1]), .ZN(n4484) );
  INV_X4 U4085 ( .A(n4587), .ZN(n4875) );
  INV_X4 U4086 ( .A(n4868), .ZN(n4864) );
  INV_X4 U4087 ( .A(n4864), .ZN(n4862) );
  INV_X4 U4088 ( .A(n4864), .ZN(n4863) );
  INV_X4 U4089 ( .A(u1_fractb_lt_fracta), .ZN(n4868) );
  NOR3_X2 U4090 ( .A1(n2049), .A2(n2033), .A3(n6406), .ZN(n1993) );
  INV_X4 U4091 ( .A(n4848), .ZN(n4837) );
  OR2_X4 U4092 ( .A1(n4896), .A2(u2_exp_tmp4_4_), .ZN(n4502) );
  NAND3_X2 U4093 ( .A1(fpu_op_r1[0]), .A2(n4501), .A3(fpu_op_r1[1]), .ZN(n4503) );
  INV_X4 U4094 ( .A(n4422), .ZN(n4876) );
  INV_X4 U4095 ( .A(n4422), .ZN(n4877) );
  INV_X4 U4096 ( .A(n4783), .ZN(n4782) );
  INV_X4 U4097 ( .A(n2532), .ZN(n4783) );
  INV_X4 U4098 ( .A(n1664), .ZN(n4772) );
  INV_X4 U4099 ( .A(n1664), .ZN(n4773) );
  INV_X4 U4100 ( .A(n1664), .ZN(n4774) );
  INV_X4 U4101 ( .A(n2342), .ZN(n4785) );
  OR2_X4 U4102 ( .A1(n4931), .A2(u4_sub_466_A_4_), .ZN(n4572) );
  NOR2_X2 U4103 ( .A1(n4875), .A2(u4_sub_407_carry[10]), .ZN(n4573) );
  INV_X4 U4104 ( .A(n4358), .ZN(n4795) );
  INV_X4 U4105 ( .A(n4357), .ZN(n4793) );
  INV_X4 U4106 ( .A(n4357), .ZN(n4794) );
  INV_X4 U4107 ( .A(n4383), .ZN(n4797) );
  INV_X4 U4108 ( .A(n4383), .ZN(n4799) );
  INV_X4 U4109 ( .A(n4822), .ZN(n4821) );
  NAND3_X2 U4110 ( .A1(fpu_op_r3[0]), .A2(n4351), .A3(fpu_op_r3[1]), .ZN(n244)
         );
  INV_X4 U4111 ( .A(n4868), .ZN(n4867) );
  INV_X4 U4112 ( .A(n4361), .ZN(n4788) );
  NOR3_X2 U4113 ( .A1(n1671), .A2(n4822), .A3(n2049), .ZN(n1991) );
  INV_X4 U4114 ( .A(n2184), .ZN(n4792) );
  INV_X4 U4115 ( .A(n4792), .ZN(n4790) );
  INV_X4 U4116 ( .A(n4849), .ZN(n4835) );
  INV_X4 U4117 ( .A(n4484), .ZN(n4820) );
  INV_X4 U4118 ( .A(n1054), .ZN(u2_lt_131_A_0_) );
  INV_X4 U4119 ( .A(n4429), .ZN(n4767) );
  INV_X4 U4120 ( .A(n4814), .ZN(n4811) );
  INV_X4 U4121 ( .A(n1090), .ZN(n4814) );
  INV_X4 U4122 ( .A(n4814), .ZN(n4812) );
  INV_X4 U4123 ( .A(n1840), .ZN(n4802) );
  INV_X4 U4124 ( .A(n4802), .ZN(n4801) );
  INV_X4 U4125 ( .A(n1091), .ZN(n4810) );
  INV_X4 U4126 ( .A(n4810), .ZN(n4808) );
  INV_X4 U4127 ( .A(n4810), .ZN(n4809) );
  INV_X4 U4128 ( .A(n4810), .ZN(n4807) );
  INV_X4 U4129 ( .A(n4384), .ZN(n4770) );
  INV_X4 U4130 ( .A(n4384), .ZN(n4771) );
  INV_X4 U4131 ( .A(n4422), .ZN(n4879) );
  INV_X4 U4132 ( .A(n4503), .ZN(n4817) );
  NAND4_X2 U4133 ( .A1(n296), .A2(n297), .A3(n298), .A4(n299), .ZN(
        u4_fi_ldz_5_) );
  NAND4_X2 U4134 ( .A1(n6408), .A2(n6423), .A3(n382), .A4(n383), .ZN(
        u4_fi_ldz_3_) );
  NAND4_X2 U4135 ( .A1(n406), .A2(n6419), .A3(n408), .A4(n409), .ZN(
        u4_fi_ldz_2_) );
  NAND4_X2 U4136 ( .A1(n6454), .A2(n321), .A3(n322), .A4(n323), .ZN(
        u4_fi_ldz_4_) );
  NOR2_X2 U4137 ( .A1(n244), .A2(opb_dn), .ZN(n2342) );
  INV_X4 U4138 ( .A(n4805), .ZN(n4804) );
  NAND3_X2 U4139 ( .A1(n1664), .A2(n2357), .A3(n6386), .ZN(N784) );
  INV_X4 U4140 ( .A(n4871), .ZN(n4870) );
  INV_X4 U4141 ( .A(n2357), .ZN(n4775) );
  INV_X4 U4142 ( .A(n2357), .ZN(n4776) );
  INV_X4 U4143 ( .A(n2357), .ZN(n4778) );
  OAI22_X2 U4144 ( .A1(u4_fi_ldz_2a_6_), .A2(n5035), .B1(u4_fi_ldz_2a_6_), 
        .B2(u4_fi_ldz_2a_5_), .ZN(u4_N6238) );
  XOR2_X2 U4147 ( .A(n4880), .B(u4_sub_489_carry[6]), .Z(u4_fi_ldz_2a_6_) );
  AND3_X4 U4148 ( .A1(n4822), .A2(n1735), .A3(n295), .ZN(n255) );
  AND2_X4 U4149 ( .A1(n6458), .A2(n367), .ZN(u4_fi_ldz_6_) );
  AND2_X4 U4150 ( .A1(n2050), .A2(n1740), .ZN(n1995) );
  AND3_X4 U4151 ( .A1(n1678), .A2(n2049), .A3(n6379), .ZN(n1997) );
  AND3_X4 U4152 ( .A1(u1_N325), .A2(n6171), .A3(u1_N75), .ZN(n777) );
  AND2_X4 U4153 ( .A1(n242), .A2(n4822), .ZN(n209) );
  XNOR2_X1 U4154 ( .A(u4_fi_ldz_6_), .B(u4_sub_461_carry_6_), .ZN(
        u4_fi_ldz_mi22[6]) );
  AND2_X1 U4155 ( .A1(u4_sub_461_carry_5_), .A2(u4_fi_ldz_5_), .ZN(
        u4_sub_461_carry_6_) );
  XOR2_X1 U4156 ( .A(u4_fi_ldz_5_), .B(u4_sub_461_carry_5_), .Z(
        u4_fi_ldz_mi22[5]) );
  AND2_X1 U4157 ( .A1(u4_sub_461_carry_4_), .A2(u4_fi_ldz_4_), .ZN(
        u4_sub_461_carry_5_) );
  XOR2_X1 U4158 ( .A(u4_fi_ldz_4_), .B(u4_sub_461_carry_4_), .Z(
        u4_fi_ldz_mi22[4]) );
  OR2_X1 U4159 ( .A1(u4_fi_ldz_3_), .A2(u4_sub_461_carry_3_), .ZN(
        u4_sub_461_carry_4_) );
  XNOR2_X1 U4160 ( .A(u4_sub_461_carry_3_), .B(u4_fi_ldz_3_), .ZN(
        u4_fi_ldz_mi22[3]) );
  OR2_X1 U4161 ( .A1(u4_fi_ldz_2_), .A2(u4_sub_461_carry_2_), .ZN(
        u4_sub_461_carry_3_) );
  XNOR2_X1 U4162 ( .A(u4_sub_461_carry_2_), .B(u4_fi_ldz_2_), .ZN(
        u4_fi_ldz_mi22[2]) );
  AND2_X1 U4163 ( .A1(u4_fi_ldz_2a_0_), .A2(u4_fi_ldz_1_), .ZN(
        u4_sub_461_carry_2_) );
  XOR2_X1 U4164 ( .A(u4_fi_ldz_1_), .B(u4_fi_ldz_2a_0_), .Z(u4_fi_ldz_mi22[1])
         );
  XOR2_X1 U4165 ( .A(n4875), .B(u4_add_408_carry[10]), .Z(u4_div_shft2[10]) );
  AND2_X1 U4166 ( .A1(n4428), .A2(u4_add_408_carry[9]), .ZN(
        u4_add_408_carry[10]) );
  XOR2_X1 U4167 ( .A(n4428), .B(u4_add_408_carry[9]), .Z(u4_div_shft2[9]) );
  XOR2_X1 U4168 ( .A(n4587), .B(u4_sub_410_carry[10]), .Z(u4_div_shft4[10]) );
  AND2_X1 U4169 ( .A1(u4_sub_410_carry[9]), .A2(n4476), .ZN(
        u4_sub_410_carry[10]) );
  XOR2_X1 U4170 ( .A(n4476), .B(u4_sub_410_carry[9]), .Z(u4_div_shft4[9]) );
  XOR2_X1 U4171 ( .A(n4875), .B(u4_add_409_carry[10]), .Z(u4_div_shft3_10_) );
  AND2_X1 U4172 ( .A1(n4428), .A2(u4_add_409_carry[9]), .ZN(
        u4_add_409_carry[10]) );
  XOR2_X1 U4173 ( .A(n4428), .B(u4_add_409_carry[9]), .Z(u4_div_shft3_9_) );
  AND2_X1 U4174 ( .A1(n4369), .A2(u4_add_408_carry[8]), .ZN(
        u4_add_408_carry[9]) );
  XOR2_X1 U4175 ( .A(n4369), .B(u4_add_408_carry[8]), .Z(u4_div_shft2[8]) );
  AND2_X1 U4176 ( .A1(u4_sub_410_carry[8]), .A2(n4474), .ZN(
        u4_sub_410_carry[9]) );
  XOR2_X1 U4177 ( .A(n4474), .B(u4_sub_410_carry[8]), .Z(u4_div_shft4[8]) );
  AND2_X1 U4178 ( .A1(n4369), .A2(u4_add_409_carry[8]), .ZN(
        u4_add_409_carry[9]) );
  XOR2_X1 U4179 ( .A(n4369), .B(u4_add_409_carry[8]), .Z(u4_div_shft3_8_) );
  AND2_X1 U4180 ( .A1(n4359), .A2(u4_add_408_carry[7]), .ZN(
        u4_add_408_carry[8]) );
  XOR2_X1 U4181 ( .A(n4359), .B(u4_add_408_carry[7]), .Z(u4_div_shft2[7]) );
  AND2_X1 U4182 ( .A1(u4_sub_410_carry[7]), .A2(n4475), .ZN(
        u4_sub_410_carry[8]) );
  XOR2_X1 U4183 ( .A(n4475), .B(u4_sub_410_carry[7]), .Z(u4_div_shft4[7]) );
  AND2_X1 U4184 ( .A1(n4359), .A2(u4_add_409_carry[7]), .ZN(
        u4_add_409_carry[8]) );
  XOR2_X1 U4185 ( .A(n4359), .B(u4_add_409_carry[7]), .Z(u4_div_shft3_7_) );
  AND2_X1 U4186 ( .A1(n4382), .A2(u4_add_408_carry[6]), .ZN(
        u4_add_408_carry[7]) );
  XOR2_X1 U4187 ( .A(n4382), .B(u4_add_408_carry[6]), .Z(u4_div_shft2[6]) );
  AND2_X1 U4188 ( .A1(n4370), .A2(u4_add_408_carry[5]), .ZN(
        u4_add_408_carry[6]) );
  XOR2_X1 U4189 ( .A(n4370), .B(u4_add_408_carry[5]), .Z(u4_div_shft2[5]) );
  AND2_X1 U4190 ( .A1(n4399), .A2(u4_add_408_carry[4]), .ZN(
        u4_add_408_carry[5]) );
  XOR2_X1 U4191 ( .A(n4399), .B(u4_add_408_carry[4]), .Z(u4_div_shft2[4]) );
  AND2_X1 U4192 ( .A1(exp_r[3]), .A2(u4_add_408_carry[3]), .ZN(
        u4_add_408_carry[4]) );
  XOR2_X1 U4193 ( .A(exp_r[3]), .B(u4_add_408_carry[3]), .Z(u4_div_shft2[3])
         );
  AND2_X1 U4194 ( .A1(exp_r[2]), .A2(n4368), .ZN(u4_add_408_carry[3]) );
  XOR2_X1 U4195 ( .A(exp_r[2]), .B(n4368), .Z(u4_div_shft2[2]) );
  AND2_X1 U4196 ( .A1(u4_sub_410_carry[6]), .A2(n4571), .ZN(
        u4_sub_410_carry[7]) );
  XOR2_X1 U4197 ( .A(n4571), .B(u4_sub_410_carry[6]), .Z(u4_div_shft4[6]) );
  AND2_X1 U4198 ( .A1(u4_sub_410_carry[5]), .A2(n4477), .ZN(
        u4_sub_410_carry[6]) );
  XOR2_X1 U4199 ( .A(n4477), .B(u4_sub_410_carry[5]), .Z(u4_div_shft4[5]) );
  OR2_X1 U4200 ( .A1(n4400), .A2(div_opa_ldz_r2[0]), .ZN(u4_sub_410_carry[1])
         );
  XNOR2_X1 U4201 ( .A(div_opa_ldz_r2[0]), .B(n4400), .ZN(u4_div_shft4[0]) );
  AND2_X1 U4202 ( .A1(n4382), .A2(u4_add_409_carry[6]), .ZN(
        u4_add_409_carry[7]) );
  XOR2_X1 U4203 ( .A(n4382), .B(u4_add_409_carry[6]), .Z(u4_div_shft3_6_) );
  AND2_X1 U4204 ( .A1(n4370), .A2(u4_add_409_carry[5]), .ZN(
        u4_add_409_carry[6]) );
  XOR2_X1 U4205 ( .A(n4370), .B(u4_add_409_carry[5]), .Z(u4_div_shft3_5_) );
  AND2_X1 U4206 ( .A1(n4823), .A2(div_opa_ldz_r2[0]), .ZN(u4_add_409_carry[1])
         );
  XOR2_X1 U4207 ( .A(n4823), .B(div_opa_ldz_r2[0]), .Z(u4_div_shft3_0_) );
  AND2_X1 U4208 ( .A1(u4_sub_479_carry[6]), .A2(n4880), .ZN(u4_N6137) );
  XOR2_X1 U4209 ( .A(n4880), .B(u4_sub_479_carry[6]), .Z(u4_N6136) );
  AND2_X1 U4210 ( .A1(u4_sub_479_carry[5]), .A2(n4881), .ZN(
        u4_sub_479_carry[6]) );
  XOR2_X1 U4211 ( .A(n4881), .B(u4_sub_479_carry[5]), .Z(u4_N6135) );
  OR2_X1 U4212 ( .A1(n4882), .A2(u4_sub_479_carry[4]), .ZN(u4_sub_479_carry[5]) );
  XNOR2_X1 U4213 ( .A(u4_sub_479_carry[4]), .B(n4882), .ZN(u4_N6134) );
  OR2_X1 U4214 ( .A1(n4935), .A2(u4_sub_479_carry[3]), .ZN(u4_sub_479_carry[4]) );
  XNOR2_X1 U4215 ( .A(u4_sub_479_carry[3]), .B(n4935), .ZN(u4_N6133) );
  OR2_X1 U4216 ( .A1(n4883), .A2(u4_sub_479_carry[2]), .ZN(u4_sub_479_carry[3]) );
  XNOR2_X1 U4217 ( .A(u4_sub_479_carry[2]), .B(n4883), .ZN(u4_N6132) );
  OR2_X1 U4218 ( .A1(n4936), .A2(u4_fi_ldz_mi1_0_), .ZN(u4_sub_479_carry[2])
         );
  XNOR2_X1 U4219 ( .A(u4_fi_ldz_mi1_0_), .B(n4936), .ZN(u4_N6131) );
  XNOR2_X1 U4220 ( .A(u4_sub_407_carry[10]), .B(n4875), .ZN(u4_div_scht1a[10])
         );
  OR2_X1 U4221 ( .A1(n4428), .A2(u4_sub_407_carry[9]), .ZN(
        u4_sub_407_carry[10]) );
  XNOR2_X1 U4222 ( .A(u4_sub_407_carry[9]), .B(n4428), .ZN(u4_div_scht1a[9])
         );
  OR2_X1 U4223 ( .A1(n4369), .A2(u4_sub_407_carry[8]), .ZN(u4_sub_407_carry[9]) );
  XNOR2_X1 U4224 ( .A(u4_sub_407_carry[8]), .B(n4369), .ZN(u4_div_scht1a[8])
         );
  OR2_X1 U4225 ( .A1(n4359), .A2(u4_sub_407_carry[7]), .ZN(u4_sub_407_carry[8]) );
  XNOR2_X1 U4226 ( .A(u4_sub_407_carry[7]), .B(n4359), .ZN(u4_div_scht1a[7])
         );
  OR2_X1 U4227 ( .A1(n4382), .A2(u4_sub_407_carry[6]), .ZN(u4_sub_407_carry[7]) );
  XNOR2_X1 U4228 ( .A(u4_sub_407_carry[6]), .B(n4382), .ZN(u4_div_scht1a[6])
         );
  OR2_X1 U4229 ( .A1(n4370), .A2(u4_sub_407_carry[5]), .ZN(u4_sub_407_carry[6]) );
  XNOR2_X1 U4230 ( .A(u4_sub_407_carry[5]), .B(n4370), .ZN(u4_div_scht1a[5])
         );
  OR2_X1 U4231 ( .A1(n4570), .A2(n4823), .ZN(u4_sub_407_carry[1]) );
  XNOR2_X1 U4232 ( .A(n4823), .B(n4570), .ZN(u4_div_scht1a[0]) );
  XNOR2_X1 U4233 ( .A(n4875), .B(u4_sub_415_carry_10_), .ZN(u4_f2i_shft_10_)
         );
  OR2_X1 U4234 ( .A1(n4428), .A2(u4_sub_415_carry_9_), .ZN(
        u4_sub_415_carry_10_) );
  XNOR2_X1 U4235 ( .A(u4_sub_415_carry_9_), .B(n4428), .ZN(u4_f2i_shft_9_) );
  OR2_X1 U4236 ( .A1(n4369), .A2(u4_sub_415_carry_8_), .ZN(u4_sub_415_carry_9_) );
  XNOR2_X1 U4237 ( .A(u4_sub_415_carry_8_), .B(n4369), .ZN(u4_f2i_shft_8_) );
  OR2_X1 U4238 ( .A1(n4359), .A2(u4_sub_415_carry_7_), .ZN(u4_sub_415_carry_8_) );
  XNOR2_X1 U4239 ( .A(u4_sub_415_carry_7_), .B(n4359), .ZN(u4_f2i_shft_7_) );
  AND2_X1 U4240 ( .A1(u4_sub_415_carry_6_), .A2(n4382), .ZN(
        u4_sub_415_carry_7_) );
  XOR2_X1 U4241 ( .A(n4382), .B(u4_sub_415_carry_6_), .Z(u4_f2i_shft_6_) );
  AND2_X1 U4242 ( .A1(u4_sub_415_carry_5_), .A2(n4370), .ZN(
        u4_sub_415_carry_6_) );
  XOR2_X1 U4243 ( .A(n4370), .B(u4_sub_415_carry_5_), .Z(u4_f2i_shft_5_) );
  AND2_X1 U4244 ( .A1(u4_sub_415_carry_4_), .A2(n4399), .ZN(
        u4_sub_415_carry_5_) );
  XOR2_X1 U4245 ( .A(n4399), .B(u4_sub_415_carry_4_), .Z(u4_f2i_shft_4_) );
  AND2_X1 U4246 ( .A1(u4_sub_415_carry_3_), .A2(exp_r[3]), .ZN(
        u4_sub_415_carry_4_) );
  XOR2_X1 U4247 ( .A(exp_r[3]), .B(u4_sub_415_carry_3_), .Z(u4_f2i_shft_3_) );
  AND2_X1 U4248 ( .A1(u4_sub_415_carry_2_), .A2(exp_r[2]), .ZN(
        u4_sub_415_carry_3_) );
  XOR2_X1 U4249 ( .A(exp_r[2]), .B(u4_sub_415_carry_2_), .Z(u4_f2i_shft_2_) );
  OR2_X1 U4250 ( .A1(n4368), .A2(n4823), .ZN(u4_sub_415_carry_2_) );
  XNOR2_X1 U4251 ( .A(n4823), .B(n4368), .ZN(u4_f2i_shft_1_) );
  XNOR2_X1 U4252 ( .A(sub_1_root_sub_0_root_u4_add_495_carry[7]), .B(
        u4_fi_ldz_2a_6_), .ZN(u4_ldz_dif_7_) );
  OR2_X1 U4253 ( .A1(u4_fi_ldz_2a_6_), .A2(
        sub_1_root_sub_0_root_u4_add_495_carry[6]), .ZN(
        sub_1_root_sub_0_root_u4_add_495_carry[7]) );
  XNOR2_X1 U4254 ( .A(sub_1_root_sub_0_root_u4_add_495_carry[6]), .B(
        u4_fi_ldz_2a_6_), .ZN(u4_ldz_dif_6_) );
  OR2_X1 U4255 ( .A1(u4_fi_ldz_2a_5_), .A2(
        sub_1_root_sub_0_root_u4_add_495_carry[5]), .ZN(
        sub_1_root_sub_0_root_u4_add_495_carry[6]) );
  XNOR2_X1 U4256 ( .A(sub_1_root_sub_0_root_u4_add_495_carry[5]), .B(
        u4_fi_ldz_2a_5_), .ZN(u4_ldz_dif_5_) );
  OR2_X1 U4257 ( .A1(n4570), .A2(u4_fi_ldz_2a_0_), .ZN(
        sub_1_root_sub_0_root_u4_add_495_carry[1]) );
  XNOR2_X1 U4258 ( .A(u4_fi_ldz_2a_0_), .B(n4570), .ZN(u4_ldz_dif_0_) );
  OR2_X1 U4259 ( .A1(n4881), .A2(u4_sub_489_carry[5]), .ZN(u4_sub_489_carry[6]) );
  XNOR2_X1 U4260 ( .A(u4_sub_489_carry[5]), .B(n4881), .ZN(u4_fi_ldz_2a_5_) );
  OR2_X1 U4261 ( .A1(n4882), .A2(u4_sub_489_carry[4]), .ZN(u4_sub_489_carry[5]) );
  XNOR2_X1 U4262 ( .A(u4_sub_489_carry[4]), .B(n4882), .ZN(u4_fi_ldz_2a_4_) );
  AND2_X1 U4263 ( .A1(u4_sub_489_carry[3]), .A2(n4935), .ZN(
        u4_sub_489_carry[4]) );
  XOR2_X1 U4264 ( .A(n4935), .B(u4_sub_489_carry[3]), .Z(u4_fi_ldz_2a_3_) );
  OR2_X1 U4265 ( .A1(n4883), .A2(u4_sub_489_carry[2]), .ZN(u4_sub_489_carry[3]) );
  XNOR2_X1 U4266 ( .A(u4_sub_489_carry[2]), .B(n4883), .ZN(u4_fi_ldz_2a_2_) );
  AND2_X1 U4267 ( .A1(u4_fi_ldz_mi1_0_), .A2(n4936), .ZN(u4_sub_489_carry[2])
         );
  XOR2_X1 U4268 ( .A(n4936), .B(u4_fi_ldz_mi1_0_), .Z(u4_fi_ldz_2a_1_) );
  XNOR2_X1 U4269 ( .A(u2_gt_141_B_11_), .B(u2_sub_112_carry_11_), .ZN(u2_N53)
         );
  OR2_X1 U4270 ( .A1(u2_exp_tmp4_10_), .A2(u2_sub_112_carry_10_), .ZN(
        u2_sub_112_carry_11_) );
  XNOR2_X1 U4271 ( .A(u2_sub_112_carry_10_), .B(u2_exp_tmp4_10_), .ZN(u2_N52)
         );
  AND2_X1 U4272 ( .A1(u2_sub_112_carry_9_), .A2(u2_lt_131_A_9_), .ZN(
        u2_sub_112_carry_10_) );
  XOR2_X1 U4273 ( .A(u2_lt_131_A_9_), .B(u2_sub_112_carry_9_), .Z(u2_N51) );
  AND2_X1 U4274 ( .A1(u2_sub_112_carry_8_), .A2(u2_lt_131_A_8_), .ZN(
        u2_sub_112_carry_9_) );
  XOR2_X1 U4275 ( .A(u2_lt_131_A_8_), .B(u2_sub_112_carry_8_), .Z(u2_N50) );
  AND2_X1 U4276 ( .A1(u2_sub_112_carry_7_), .A2(u2_lt_131_A_7_), .ZN(
        u2_sub_112_carry_8_) );
  XOR2_X1 U4277 ( .A(u2_lt_131_A_7_), .B(u2_sub_112_carry_7_), .Z(u2_N49) );
  AND2_X1 U4278 ( .A1(u2_sub_112_carry_6_), .A2(u2_lt_131_A_6_), .ZN(
        u2_sub_112_carry_7_) );
  XOR2_X1 U4279 ( .A(u2_lt_131_A_6_), .B(u2_sub_112_carry_6_), .Z(u2_N48) );
  AND2_X1 U4280 ( .A1(u2_sub_112_carry_5_), .A2(u2_lt_131_A_5_), .ZN(
        u2_sub_112_carry_6_) );
  XOR2_X1 U4281 ( .A(u2_lt_131_A_5_), .B(u2_sub_112_carry_5_), .Z(u2_N47) );
  AND2_X1 U4282 ( .A1(u2_sub_112_carry_4_), .A2(u2_lt_131_A_4_), .ZN(
        u2_sub_112_carry_5_) );
  XOR2_X1 U4283 ( .A(u2_lt_131_A_4_), .B(u2_sub_112_carry_4_), .Z(u2_N46) );
  AND2_X1 U4284 ( .A1(u2_sub_112_carry_3_), .A2(u2_exp_tmp1_3_), .ZN(
        u2_sub_112_carry_4_) );
  XOR2_X1 U4285 ( .A(u2_exp_tmp1_3_), .B(u2_sub_112_carry_3_), .Z(u2_N45) );
  AND2_X1 U4286 ( .A1(u2_sub_112_carry_2_), .A2(u2_exp_tmp1_2_), .ZN(
        u2_sub_112_carry_3_) );
  XOR2_X1 U4287 ( .A(u2_exp_tmp1_2_), .B(u2_sub_112_carry_2_), .Z(u2_N44) );
  AND2_X1 U4288 ( .A1(u2_lt_131_A_0_), .A2(u2_exp_tmp1_1_), .ZN(
        u2_sub_112_carry_2_) );
  XOR2_X1 U4289 ( .A(u2_exp_tmp1_1_), .B(u2_lt_131_A_0_), .Z(u2_N43) );
  XOR2_X1 U4290 ( .A(u2_gt_141_B_11_), .B(u2_add_112_carry_11_), .Z(u2_N41) );
  AND2_X1 U4291 ( .A1(u2_add_112_carry_10_), .A2(u2_exp_tmp4_10_), .ZN(
        u2_add_112_carry_11_) );
  XOR2_X1 U4292 ( .A(u2_exp_tmp4_10_), .B(u2_add_112_carry_10_), .Z(u2_N40) );
  OR2_X1 U4293 ( .A1(u2_lt_131_A_9_), .A2(u2_add_112_carry_9_), .ZN(
        u2_add_112_carry_10_) );
  XNOR2_X1 U4294 ( .A(u2_add_112_carry_9_), .B(u2_lt_131_A_9_), .ZN(u2_N39) );
  OR2_X1 U4295 ( .A1(u2_lt_131_A_8_), .A2(u2_add_112_carry_8_), .ZN(
        u2_add_112_carry_9_) );
  XNOR2_X1 U4296 ( .A(u2_add_112_carry_8_), .B(u2_lt_131_A_8_), .ZN(u2_N38) );
  OR2_X1 U4297 ( .A1(u2_lt_131_A_7_), .A2(u2_add_112_carry_7_), .ZN(
        u2_add_112_carry_8_) );
  XNOR2_X1 U4298 ( .A(u2_add_112_carry_7_), .B(u2_lt_131_A_7_), .ZN(u2_N37) );
  OR2_X1 U4299 ( .A1(u2_lt_131_A_6_), .A2(u2_add_112_carry_6_), .ZN(
        u2_add_112_carry_7_) );
  XNOR2_X1 U4300 ( .A(u2_add_112_carry_6_), .B(u2_lt_131_A_6_), .ZN(u2_N36) );
  OR2_X1 U4301 ( .A1(u2_lt_131_A_5_), .A2(u2_add_112_carry_5_), .ZN(
        u2_add_112_carry_6_) );
  XNOR2_X1 U4302 ( .A(u2_add_112_carry_5_), .B(u2_lt_131_A_5_), .ZN(u2_N35) );
  OR2_X1 U4303 ( .A1(u2_lt_131_A_4_), .A2(u2_add_112_carry_4_), .ZN(
        u2_add_112_carry_5_) );
  XNOR2_X1 U4304 ( .A(u2_add_112_carry_4_), .B(u2_lt_131_A_4_), .ZN(u2_N34) );
  OR2_X1 U4305 ( .A1(u2_exp_tmp1_3_), .A2(u2_add_112_carry_3_), .ZN(
        u2_add_112_carry_4_) );
  XNOR2_X1 U4306 ( .A(u2_add_112_carry_3_), .B(u2_exp_tmp1_3_), .ZN(u2_N33) );
  OR2_X1 U4307 ( .A1(u2_exp_tmp1_2_), .A2(u2_add_112_carry_2_), .ZN(
        u2_add_112_carry_3_) );
  XNOR2_X1 U4308 ( .A(u2_add_112_carry_2_), .B(u2_exp_tmp1_2_), .ZN(u2_N32) );
  OR2_X1 U4309 ( .A1(u2_exp_tmp1_1_), .A2(u2_lt_131_A_0_), .ZN(
        u2_add_112_carry_2_) );
  XNOR2_X1 U4310 ( .A(u2_lt_131_A_0_), .B(u2_exp_tmp1_1_), .ZN(u2_N31) );
  INV_X4 U4311 ( .A(u4_fi_ldz_6_), .ZN(n4880) );
  INV_X4 U4312 ( .A(u4_fi_ldz_5_), .ZN(n4881) );
  INV_X4 U4313 ( .A(u4_fi_ldz_4_), .ZN(n4882) );
  INV_X4 U4314 ( .A(u4_fi_ldz_2_), .ZN(n4883) );
  INV_X4 U4315 ( .A(u2_exp_tmp1_1_), .ZN(u2_exp_tmp4_1_) );
  INV_X4 U4316 ( .A(u2_exp_tmp1_2_), .ZN(u2_exp_tmp4_2_) );
  INV_X4 U4317 ( .A(u2_exp_tmp1_3_), .ZN(u2_exp_tmp4_3_) );
  INV_X4 U4318 ( .A(u2_lt_131_A_4_), .ZN(u2_exp_tmp4_4_) );
  NOR2_X1 U4319 ( .A1(u2_exp_tmp4_1_), .A2(n1054), .ZN(n4885) );
  NOR2_X1 U4320 ( .A1(n4894), .A2(u2_exp_tmp4_2_), .ZN(n4886) );
  NOR2_X1 U4321 ( .A1(n4895), .A2(u2_exp_tmp4_3_), .ZN(n4887) );
  NOR2_X1 U4322 ( .A1(n4502), .A2(n1052), .ZN(n4889) );
  NAND2_X1 U4323 ( .A1(n4889), .A2(u2_lt_131_A_6_), .ZN(n4890) );
  NOR2_X1 U4324 ( .A1(n4890), .A2(n1050), .ZN(n4892) );
  NAND2_X1 U4325 ( .A1(n4892), .A2(u2_lt_131_A_8_), .ZN(n4893) );
  NOR2_X1 U4326 ( .A1(n1048), .A2(n4893), .ZN(n4884) );
  XOR2_X1 U4327 ( .A(u2_exp_tmp4_10_), .B(n4884), .Z(u2_N75) );
  OAI21_X1 U4328 ( .B1(u2_lt_131_A_0_), .B2(u2_exp_tmp1_1_), .A(n4894), .ZN(
        u2_N66) );
  OAI21_X1 U4329 ( .B1(n4885), .B2(u2_exp_tmp1_2_), .A(n4895), .ZN(u2_N67) );
  OAI21_X1 U4330 ( .B1(n4886), .B2(u2_exp_tmp1_3_), .A(n4896), .ZN(u2_N68) );
  OAI21_X1 U4331 ( .B1(n4887), .B2(u2_lt_131_A_4_), .A(n4502), .ZN(u2_N69) );
  AOI21_X1 U4332 ( .B1(n4502), .B2(n1052), .A(n4889), .ZN(n4888) );
  OAI21_X1 U4333 ( .B1(n4889), .B2(u2_lt_131_A_6_), .A(n4890), .ZN(u2_N71) );
  AOI21_X1 U4334 ( .B1(n4890), .B2(n1050), .A(n4892), .ZN(n4891) );
  OAI21_X1 U4335 ( .B1(n4892), .B2(u2_lt_131_A_8_), .A(n4893), .ZN(u2_N73) );
  XNOR2_X1 U4336 ( .A(n1048), .B(n4893), .ZN(u2_N74) );
  INV_X4 U4337 ( .A(n4885), .ZN(n4894) );
  INV_X4 U4338 ( .A(n4886), .ZN(n4895) );
  INV_X4 U4339 ( .A(n4887), .ZN(n4896) );
  INV_X4 U4340 ( .A(n4888), .ZN(u2_N70) );
  INV_X4 U4341 ( .A(n4891), .ZN(u2_N72) );
  NOR2_X1 U4342 ( .A1(n4368), .A2(n4823), .ZN(n4898) );
  NOR2_X1 U4343 ( .A1(u4_sub_415_carry_2_), .A2(exp_r[2]), .ZN(n4899) );
  NOR2_X1 U4344 ( .A1(n4906), .A2(exp_r[3]), .ZN(n4900) );
  NOR2_X1 U4345 ( .A1(n4907), .A2(n4399), .ZN(n4901) );
  NOR2_X1 U4346 ( .A1(n4908), .A2(n4370), .ZN(n4902) );
  NOR2_X1 U4347 ( .A1(n4478), .A2(n4359), .ZN(n4904) );
  NAND2_X1 U4348 ( .A1(n4904), .A2(n4474), .ZN(n4905) );
  NOR3_X1 U4349 ( .A1(n4875), .A2(n4428), .A3(n4905), .ZN(u4_exp_in_mi1_11_)
         );
  OAI21_X1 U4350 ( .B1(n4428), .B2(n4905), .A(exp_r[10]), .ZN(n4897) );
  NAND2_X1 U4351 ( .A1(n6520), .A2(n4897), .ZN(u4_exp_in_mi1_10_) );
  OAI21_X1 U4352 ( .B1(n4400), .B2(n4588), .A(u4_sub_415_carry_2_), .ZN(
        u4_exp_in_mi1_1_) );
  OAI21_X1 U4353 ( .B1(n4898), .B2(n4425), .A(n4906), .ZN(u4_exp_in_mi1_2_) );
  OAI21_X1 U4354 ( .B1(n4899), .B2(n4473), .A(n4907), .ZN(u4_exp_in_mi1_3_) );
  OAI21_X1 U4355 ( .B1(n4900), .B2(n4424), .A(n4908), .ZN(u4_exp_in_mi1_4_) );
  OAI21_X1 U4356 ( .B1(n4901), .B2(n4477), .A(n4909), .ZN(u4_exp_in_mi1_5_) );
  OAI21_X1 U4357 ( .B1(n4902), .B2(n4571), .A(n4478), .ZN(u4_exp_in_mi1_6_) );
  AOI21_X1 U4358 ( .B1(n4478), .B2(n4359), .A(n4904), .ZN(n4903) );
  OAI21_X1 U4359 ( .B1(n4904), .B2(n4474), .A(n4905), .ZN(u4_exp_in_mi1_8_) );
  XNOR2_X1 U4360 ( .A(n4428), .B(n4905), .ZN(u4_exp_in_mi1_9_) );
  INV_X4 U4361 ( .A(n4899), .ZN(n4906) );
  INV_X4 U4362 ( .A(n4900), .ZN(n4907) );
  INV_X4 U4363 ( .A(n4901), .ZN(n4908) );
  INV_X4 U4364 ( .A(n4902), .ZN(n4909) );
  INV_X4 U4365 ( .A(n4903), .ZN(u4_exp_in_mi1_7_) );
  NOR2_X1 U4366 ( .A1(u4_fi_ldz_1_), .A2(u4_fi_ldz_2a_0_), .ZN(n4911) );
  AOI21_X1 U4367 ( .B1(u4_fi_ldz_2a_0_), .B2(u4_fi_ldz_1_), .A(n4911), .ZN(
        n4910) );
  NAND2_X1 U4368 ( .A1(n4911), .A2(n4883), .ZN(n4912) );
  OAI21_X1 U4369 ( .B1(n4911), .B2(n4883), .A(n4912), .ZN(u4_fi_ldz_mi1_2_) );
  NOR2_X1 U4370 ( .A1(n4912), .A2(u4_fi_ldz_3_), .ZN(n4914) );
  AOI21_X1 U4371 ( .B1(n4912), .B2(u4_fi_ldz_3_), .A(n4914), .ZN(n4913) );
  NAND2_X1 U4372 ( .A1(n4914), .A2(n4882), .ZN(n4915) );
  OAI21_X1 U4373 ( .B1(n4914), .B2(n4882), .A(n4915), .ZN(u4_fi_ldz_mi1_4_) );
  XNOR2_X1 U4374 ( .A(u4_fi_ldz_5_), .B(n4915), .ZN(u4_fi_ldz_mi1_5_) );
  NOR2_X1 U4375 ( .A1(u4_fi_ldz_5_), .A2(n4915), .ZN(n4916) );
  XOR2_X1 U4376 ( .A(u4_fi_ldz_6_), .B(n4916), .Z(u4_fi_ldz_mi1_6_) );
  INV_X4 U4377 ( .A(u4_fi_ldz_2a_0_), .ZN(u4_fi_ldz_mi1_0_) );
  INV_X4 U4378 ( .A(n4913), .ZN(u4_fi_ldz_mi1_3_) );
  INV_X4 U4379 ( .A(n4910), .ZN(u4_fi_ldz_mi1_1_) );
  NOR2_X1 U4380 ( .A1(u4_exp_out1_1_), .A2(u4_sub_466_A_0_), .ZN(n4918) );
  NOR2_X1 U4381 ( .A1(n4927), .A2(u4_sub_466_A_2_), .ZN(n4919) );
  NOR2_X1 U4382 ( .A1(n4929), .A2(u4_sub_466_A_3_), .ZN(n4920) );
  NOR2_X1 U4383 ( .A1(n4572), .A2(u4_sub_466_A_5_), .ZN(n4922) );
  NAND2_X1 U4384 ( .A1(n4922), .A2(n2115), .ZN(n4923) );
  NOR2_X1 U4385 ( .A1(n4923), .A2(u4_sub_466_A_7_), .ZN(n4925) );
  NAND2_X1 U4386 ( .A1(n4925), .A2(n4934), .ZN(n4926) );
  NOR2_X1 U4387 ( .A1(u4_sub_466_A_9_), .A2(n4926), .ZN(n4917) );
  XOR2_X1 U4388 ( .A(u4_sub_466_A_10_), .B(n4917), .Z(u4_exp_out1_mi1[10]) );
  OAI21_X1 U4389 ( .B1(u4_exp_out1_mi1[0]), .B2(n4928), .A(n4927), .ZN(
        u4_exp_out1_mi1[1]) );
  OAI21_X1 U4390 ( .B1(n4918), .B2(n4930), .A(n4929), .ZN(u4_exp_out1_mi1[2])
         );
  OAI21_X1 U4391 ( .B1(n4919), .B2(n4932), .A(n4931), .ZN(u4_exp_out1_mi1[3])
         );
  OAI21_X1 U4392 ( .B1(n4920), .B2(n4933), .A(n4572), .ZN(u4_exp_out1_mi1[4])
         );
  AOI21_X1 U4393 ( .B1(n4572), .B2(u4_sub_466_A_5_), .A(n4922), .ZN(n4921) );
  OAI21_X1 U4394 ( .B1(n4922), .B2(n2115), .A(n4923), .ZN(u4_exp_out1_mi1[6])
         );
  AOI21_X1 U4395 ( .B1(n4923), .B2(u4_sub_466_A_7_), .A(n4925), .ZN(n4924) );
  OAI21_X1 U4396 ( .B1(n4925), .B2(n4934), .A(n4926), .ZN(u4_exp_out1_mi1[8])
         );
  XNOR2_X1 U4397 ( .A(u4_sub_466_A_9_), .B(n4926), .ZN(u4_exp_out1_mi1[9]) );
  INV_X4 U4398 ( .A(u4_sub_466_A_0_), .ZN(u4_exp_out1_mi1[0]) );
  INV_X4 U4399 ( .A(n4918), .ZN(n4927) );
  INV_X4 U4400 ( .A(u4_exp_out1_1_), .ZN(n4928) );
  INV_X4 U4401 ( .A(n4919), .ZN(n4929) );
  INV_X4 U4402 ( .A(u4_sub_466_A_2_), .ZN(n4930) );
  INV_X4 U4403 ( .A(n4920), .ZN(n4931) );
  INV_X4 U4404 ( .A(u4_sub_466_A_3_), .ZN(n4932) );
  INV_X4 U4405 ( .A(u4_sub_466_A_4_), .ZN(n4933) );
  INV_X4 U4406 ( .A(n4921), .ZN(u4_exp_out1_mi1[5]) );
  INV_X4 U4407 ( .A(n4924), .ZN(u4_exp_out1_mi1[7]) );
  INV_X4 U4408 ( .A(u4_sub_466_A_8_), .ZN(n4934) );
  INV_X4 U4409 ( .A(u4_fi_ldz_3_), .ZN(n4935) );
  INV_X4 U4410 ( .A(u4_fi_ldz_1_), .ZN(n4936) );
  INV_X1 U4411 ( .A(u4_exp_out_0_), .ZN(u4_exp_out_mi1[0]) );
  NOR2_X1 U4412 ( .A1(u4_exp_out_1_), .A2(u4_exp_out_0_), .ZN(n4940) );
  INV_X1 U4413 ( .A(n4940), .ZN(n4938) );
  NOR2_X1 U4414 ( .A1(n4938), .A2(u4_exp_out_2_), .ZN(n4942) );
  INV_X1 U4415 ( .A(n4942), .ZN(n4939) );
  NOR2_X1 U4416 ( .A1(n4939), .A2(u4_exp_out_3_), .ZN(n4943) );
  INV_X1 U4417 ( .A(n4943), .ZN(n4941) );
  NOR2_X1 U4418 ( .A1(n4472), .A2(u4_exp_out_5_), .ZN(n4946) );
  INV_X1 U4419 ( .A(u4_exp_out_6_), .ZN(n4945) );
  NAND2_X1 U4420 ( .A1(n4946), .A2(n4945), .ZN(n4947) );
  NOR2_X1 U4421 ( .A1(n4947), .A2(u4_exp_out_7_), .ZN(n4950) );
  INV_X1 U4422 ( .A(u4_exp_out_8_), .ZN(n4949) );
  NAND2_X1 U4423 ( .A1(n4950), .A2(n4949), .ZN(n4951) );
  NOR2_X1 U4424 ( .A1(u4_exp_out_9_), .A2(n4951), .ZN(n4937) );
  XOR2_X1 U4425 ( .A(u4_exp_out_10_), .B(n4937), .Z(u4_exp_out_mi1[10]) );
  OAI21_X1 U4426 ( .B1(u4_exp_out_mi1[0]), .B2(n234), .A(n4938), .ZN(
        u4_exp_out_mi1[1]) );
  OAI21_X1 U4427 ( .B1(n4940), .B2(n231), .A(n4939), .ZN(u4_exp_out_mi1[2]) );
  OAI21_X1 U4428 ( .B1(n4942), .B2(n228), .A(n4941), .ZN(u4_exp_out_mi1[3]) );
  OAI21_X1 U4429 ( .B1(n4943), .B2(n225), .A(n4472), .ZN(u4_exp_out_mi1[4]) );
  AOI21_X1 U4430 ( .B1(n4472), .B2(u4_exp_out_5_), .A(n4946), .ZN(n4944) );
  INV_X1 U4431 ( .A(n4944), .ZN(u4_exp_out_mi1[5]) );
  OAI21_X1 U4432 ( .B1(n4946), .B2(n4945), .A(n4947), .ZN(u4_exp_out_mi1[6])
         );
  AOI21_X1 U4433 ( .B1(n4947), .B2(u4_exp_out_7_), .A(n4950), .ZN(n4948) );
  INV_X1 U4434 ( .A(n4948), .ZN(u4_exp_out_mi1[7]) );
  OAI21_X1 U4435 ( .B1(n4950), .B2(n4949), .A(n4951), .ZN(u4_exp_out_mi1[8])
         );
  XNOR2_X1 U4436 ( .A(u4_exp_out_9_), .B(n4951), .ZN(u4_exp_out_mi1[9]) );
  NAND2_X1 U4437 ( .A1(opb_r[54]), .A2(n4583), .ZN(n4968) );
  NAND2_X1 U4438 ( .A1(opb_r[59]), .A2(n4582), .ZN(n4970) );
  NAND2_X1 U4439 ( .A1(opb_r[60]), .A2(n4580), .ZN(n4971) );
  NAND2_X1 U4440 ( .A1(opb_r[57]), .A2(n4586), .ZN(n4965) );
  NAND2_X1 U4441 ( .A1(opb_r[58]), .A2(n4575), .ZN(n4963) );
  NAND2_X1 U4442 ( .A1(opb_r[55]), .A2(n4485), .ZN(n4964) );
  NAND2_X1 U4443 ( .A1(opb_r[56]), .A2(n4589), .ZN(n4967) );
  NOR2_X1 U4444 ( .A1(n4585), .A2(opb_r[52]), .ZN(n4953) );
  OAI21_X1 U4445 ( .B1(n4979), .B2(n4584), .A(opb_r[53]), .ZN(n4952) );
  OAI211_X1 U4446 ( .C1(opa_r[53]), .C2(n4953), .A(n4952), .B(n4968), .ZN(
        n4954) );
  OAI221_X1 U4447 ( .B1(opb_r[54]), .B2(n4583), .C1(opb_r[55]), .C2(n4485), 
        .A(n4954), .ZN(n4955) );
  NAND3_X1 U4448 ( .A1(n4964), .A2(n4967), .A3(n4955), .ZN(n4956) );
  OAI221_X1 U4449 ( .B1(opb_r[56]), .B2(n4589), .C1(opb_r[57]), .C2(n4586), 
        .A(n4956), .ZN(n4957) );
  NAND3_X1 U4450 ( .A1(n4965), .A2(n4963), .A3(n4957), .ZN(n4958) );
  OAI221_X1 U4451 ( .B1(opb_r[58]), .B2(n4575), .C1(opb_r[59]), .C2(n4582), 
        .A(n4958), .ZN(n4959) );
  NAND3_X1 U4452 ( .A1(n4970), .A2(n4971), .A3(n4959), .ZN(n4960) );
  OAI221_X1 U4453 ( .B1(opb_r[60]), .B2(n4580), .C1(opb_r[61]), .C2(n4482), 
        .A(n4960), .ZN(n4961) );
  NAND2_X1 U4454 ( .A1(opb_r[61]), .A2(n4482), .ZN(n4972) );
  OAI211_X1 U4455 ( .C1(opa_r[62]), .C2(n4978), .A(n4961), .B(n4972), .ZN(
        n4962) );
  AOI21_X1 U4456 ( .B1(n4978), .B2(opa_r[62]), .A(n4980), .ZN(n4977) );
  AND3_X1 U4457 ( .A1(n4965), .A2(n4964), .A3(n4963), .ZN(n4966) );
  NAND4_X1 U4458 ( .A1(n4968), .A2(n4977), .A3(n4967), .A4(n4966), .ZN(n4976)
         );
  AND2_X1 U4459 ( .A1(opb_r[52]), .A2(n4585), .ZN(n4969) );
  OAI22_X1 U4460 ( .A1(n4969), .A2(n4584), .B1(opb_r[53]), .B2(n4969), .ZN(
        n4974) );
  AND3_X1 U4461 ( .A1(n4972), .A2(n4971), .A3(n4970), .ZN(n4973) );
  OAI211_X1 U4462 ( .C1(opa_r[62]), .C2(n4978), .A(n4974), .B(n4973), .ZN(
        n4975) );
  NOR2_X1 U4463 ( .A1(n4976), .A2(n4975), .ZN(u1_N75) );
  INV_X4 U4464 ( .A(opb_r[62]), .ZN(n4978) );
  INV_X4 U4465 ( .A(n4953), .ZN(n4979) );
  INV_X4 U4466 ( .A(n4962), .ZN(n4980) );
  INV_X4 U4467 ( .A(n4977), .ZN(u1_expa_lt_expb) );
  NOR2_X1 U4468 ( .A1(u1_exp_diff_6_), .A2(u1_exp_diff_10_), .ZN(n4984) );
  OR3_X1 U4469 ( .A1(u1_exp_diff_2_), .A2(u1_exp_diff_1_), .A3(u1_exp_diff_0_), 
        .ZN(n4981) );
  NAND4_X1 U4470 ( .A1(u1_exp_diff_5_), .A2(u1_exp_diff_4_), .A3(
        u1_exp_diff_3_), .A4(n4981), .ZN(n4983) );
  NOR3_X1 U4471 ( .A1(u1_exp_diff_7_), .A2(u1_exp_diff_9_), .A3(u1_exp_diff_8_), .ZN(n4982) );
  NAND3_X1 U4472 ( .A1(n4984), .A2(n4983), .A3(n4982), .ZN(u1_exp_lt_27) );
  NOR2_X1 U4473 ( .A1(u4_div_shft3_6_), .A2(u4_div_shft3_10_), .ZN(n4987) );
  OAI211_X1 U4474 ( .C1(u4_div_shft3_2_), .C2(u4_div_shft3_3_), .A(
        u4_div_shft3_4_), .B(u4_div_shft3_5_), .ZN(n4986) );
  NOR3_X1 U4475 ( .A1(u4_div_shft3_7_), .A2(u4_div_shft3_9_), .A3(
        u4_div_shft3_8_), .ZN(n4985) );
  NAND3_X1 U4476 ( .A1(n4987), .A2(n4986), .A3(n4985), .ZN(u4_N5837) );
  NAND4_X1 U4477 ( .A1(u4_div_exp2_3_), .A2(u4_div_exp2_2_), .A3(
        u4_div_exp2_1_), .A4(u4_div_exp2_0_), .ZN(n4989) );
  NAND4_X1 U4478 ( .A1(u4_div_exp2_7_), .A2(u4_div_exp2_6_), .A3(
        u4_div_exp2_5_), .A4(u4_div_exp2_4_), .ZN(n4988) );
  NOR2_X1 U4479 ( .A1(n4989), .A2(n4988), .ZN(n4990) );
  OR4_X1 U4480 ( .A1(u4_div_exp2_10_), .A2(n4990), .A3(u4_div_exp2_9_), .A4(
        u4_div_exp2_8_), .ZN(u4_N6159) );
  NAND3_X1 U4481 ( .A1(u4_div_exp1_1_), .A2(u4_div_exp1_0_), .A3(
        u4_div_exp1_2_), .ZN(n4994) );
  NAND2_X1 U4482 ( .A1(u4_div_exp1_4_), .A2(u4_div_exp1_3_), .ZN(n4993) );
  NAND3_X1 U4483 ( .A1(u4_div_exp1_6_), .A2(u4_div_exp1_5_), .A3(
        u4_div_exp1_7_), .ZN(n4992) );
  NAND2_X1 U4484 ( .A1(u4_div_exp1_9_), .A2(u4_div_exp1_8_), .ZN(n4991) );
  NOR4_X1 U4485 ( .A1(n4994), .A2(n4993), .A3(n4992), .A4(n4991), .ZN(n4995)
         );
  NOR2_X1 U4486 ( .A1(u4_div_exp1_10_), .A2(n4995), .ZN(u4_N6179) );
  OAI211_X1 U4487 ( .C1(u4_ldz_all_3_), .C2(u4_ldz_all_2_), .A(u4_ldz_all_4_), 
        .B(u4_ldz_all_5_), .ZN(n4996) );
  NOR2_X1 U4488 ( .A1(u4_ldz_all_6_), .A2(n4997), .ZN(u4_N6275) );
  INV_X4 U4489 ( .A(n4996), .ZN(n4997) );
  OR3_X1 U4490 ( .A1(n4399), .A2(exp_r[3]), .A3(exp_r[2]), .ZN(n4998) );
  OR3_X1 U4491 ( .A1(n4368), .A2(n4823), .A3(n4998), .ZN(n4999) );
  AOI211_X1 U4492 ( .C1(n4370), .C2(n4999), .A(n4382), .B(exp_r[10]), .ZN(
        n5001) );
  NOR3_X1 U4493 ( .A1(n4359), .A2(n4428), .A3(n4369), .ZN(n5000) );
  NAND2_X1 U4494 ( .A1(n5001), .A2(n5000), .ZN(u4_N6273) );
  NAND4_X1 U4495 ( .A1(exp_r[3]), .A2(exp_r[2]), .A3(n4368), .A4(n4823), .ZN(
        n5003) );
  NAND3_X1 U4496 ( .A1(n4370), .A2(n4399), .A3(n4382), .ZN(n5002) );
  OAI21_X1 U4497 ( .B1(n5003), .B2(n5002), .A(n4587), .ZN(n5004) );
  NOR4_X1 U4498 ( .A1(n5004), .A2(n4359), .A3(n4428), .A4(n4369), .ZN(u4_N6272) );
  NOR2_X1 U4499 ( .A1(n4382), .A2(exp_r[10]), .ZN(n5006) );
  OAI211_X1 U4500 ( .C1(exp_r[3]), .C2(exp_r[2]), .A(n4399), .B(n4370), .ZN(
        n5005) );
  NAND2_X1 U4501 ( .A1(n5006), .A2(n5005), .ZN(n5007) );
  NOR4_X1 U4502 ( .A1(n5007), .A2(n4359), .A3(n4428), .A4(n4369), .ZN(u4_N6269) );
  NOR2_X1 U4503 ( .A1(n4370), .A2(exp_r[10]), .ZN(n5011) );
  AND3_X1 U4504 ( .A1(n4368), .A2(n4823), .A3(exp_r[2]), .ZN(n5008) );
  OAI21_X1 U4505 ( .B1(n5008), .B2(exp_r[3]), .A(n4399), .ZN(n5010) );
  NOR4_X1 U4506 ( .A1(n4428), .A2(n4369), .A3(n4359), .A4(n4382), .ZN(n5009)
         );
  NAND3_X1 U4507 ( .A1(n5011), .A2(n5010), .A3(n5009), .ZN(u4_N6267) );
  AND2_X1 U4508 ( .A1(u4_fi_ldz_2a_4_), .A2(u4_fi_ldz_2a_3_), .ZN(n5012) );
  OAI211_X1 U4509 ( .C1(u4_fi_ldz_2_), .C2(u4_fi_ldz_3_), .A(u4_fi_ldz_5_), 
        .B(u4_fi_ldz_4_), .ZN(n5013) );
  NAND2_X1 U4510 ( .A1(n4880), .A2(n5013), .ZN(u4_N6188) );
  OR4_X1 U4511 ( .A1(n4359), .A2(n4382), .A3(n4428), .A4(n4369), .ZN(n5020) );
  NOR2_X1 U4512 ( .A1(n4570), .A2(n4823), .ZN(n5014) );
  AOI21_X1 U4513 ( .B1(n5014), .B2(n4588), .A(div_opa_ldz_r2[1]), .ZN(n5015)
         );
  AOI221_X1 U4514 ( .B1(exp_r[2]), .B2(n4577), .C1(n4368), .C2(
        u4_sub_407_carry[1]), .A(n5015), .ZN(n5016) );
  AOI221_X1 U4515 ( .B1(div_opa_ldz_r2[3]), .B2(n4473), .C1(div_opa_ldz_r2[2]), 
        .C2(n4425), .A(n5016), .ZN(n5017) );
  AOI221_X1 U4516 ( .B1(n4399), .B2(n4581), .C1(exp_r[3]), .C2(n4576), .A(
        n5017), .ZN(n5018) );
  AOI21_X1 U4517 ( .B1(div_opa_ldz_r2[4]), .B2(n4424), .A(n5018), .ZN(n5019)
         );
  NOR4_X1 U4518 ( .A1(n5020), .A2(n5019), .A3(n4370), .A4(n4875), .ZN(u4_N6158) );
  NAND3_X1 U4519 ( .A1(u2_exp_tmp1_1_), .A2(u2_lt_131_A_0_), .A3(
        u2_exp_tmp1_2_), .ZN(n5024) );
  NAND2_X1 U4520 ( .A1(u2_lt_131_A_4_), .A2(u2_exp_tmp1_3_), .ZN(n5023) );
  NAND3_X1 U4521 ( .A1(u2_lt_131_A_6_), .A2(u2_lt_131_A_5_), .A3(
        u2_lt_131_A_7_), .ZN(n5022) );
  NAND2_X1 U4522 ( .A1(u2_lt_131_A_9_), .A2(u2_lt_131_A_8_), .ZN(n5021) );
  NOR4_X1 U4523 ( .A1(n5024), .A2(n5023), .A3(n5022), .A4(n5021), .ZN(n5025)
         );
  OAI21_X1 U4524 ( .B1(n5025), .B2(u2_exp_tmp4_10_), .A(u2_gt_141_B_11_), .ZN(
        n5026) );
  INV_X4 U4525 ( .A(n5026), .ZN(u2_N113) );
  NAND3_X1 U4526 ( .A1(u2_exp_tmp1_1_), .A2(u2_lt_131_A_0_), .A3(
        u2_exp_tmp1_2_), .ZN(n5030) );
  NAND2_X1 U4527 ( .A1(u2_lt_131_A_4_), .A2(u2_exp_tmp1_3_), .ZN(n5029) );
  NAND3_X1 U4528 ( .A1(u2_lt_131_A_6_), .A2(u2_lt_131_A_5_), .A3(
        u2_lt_131_A_7_), .ZN(n5028) );
  NAND2_X1 U4529 ( .A1(u2_lt_131_A_9_), .A2(u2_lt_131_A_8_), .ZN(n5027) );
  NOR4_X1 U4530 ( .A1(n5030), .A2(n5029), .A3(n5028), .A4(n5027), .ZN(n5031)
         );
  NOR2_X1 U4531 ( .A1(u2_exp_tmp4_10_), .A2(n5031), .ZN(u2_N111) );
  OAI211_X1 U4532 ( .C1(u4_fi_ldz_3_), .C2(u4_fi_ldz_2_), .A(u4_fi_ldz_4_), 
        .B(u4_fi_ldz_5_), .ZN(n5032) );
  NOR2_X1 U4533 ( .A1(u4_fi_ldz_6_), .A2(n5033), .ZN(u4_N6268) );
  INV_X4 U4534 ( .A(n5032), .ZN(n5033) );
  OAI21_X1 U4535 ( .B1(u4_fi_ldz_2a_1_), .B2(u4_fi_ldz_2a_0_), .A(
        u4_fi_ldz_2a_2_), .ZN(n5034) );
  AOI21_X1 U4536 ( .B1(n5034), .B2(n5036), .A(n5037), .ZN(n5035) );
  INV_X4 U4537 ( .A(u4_fi_ldz_2a_3_), .ZN(n5036) );
  INV_X4 U4538 ( .A(u4_fi_ldz_2a_4_), .ZN(n5037) );
  NOR2_X1 U4539 ( .A1(n4382), .A2(n4370), .ZN(n5039) );
  NAND4_X1 U4540 ( .A1(n4368), .A2(exp_r[2]), .A3(n4399), .A4(exp_r[3]), .ZN(
        n5038) );
  AOI21_X1 U4541 ( .B1(n5039), .B2(n5038), .A(n4475), .ZN(n5040) );
  OR4_X1 U4542 ( .A1(n4875), .A2(n5040), .A3(n4428), .A4(n4369), .ZN(u4_N5831)
         );
  OAI211_X1 U4543 ( .C1(n4823), .C2(n5046), .A(n4368), .B(exp_r[2]), .ZN(n5044) );
  NAND2_X1 U4544 ( .A1(n4399), .A2(exp_r[3]), .ZN(n5043) );
  NAND3_X1 U4545 ( .A1(n4382), .A2(n4370), .A3(n4359), .ZN(n5042) );
  NAND2_X1 U4546 ( .A1(n4428), .A2(n4369), .ZN(n5041) );
  NOR4_X1 U4547 ( .A1(n5044), .A2(n5043), .A3(n5042), .A4(n5041), .ZN(n5045)
         );
  NOR2_X1 U4548 ( .A1(n4875), .A2(n5045), .ZN(u4_N5830) );
  INV_X4 U4549 ( .A(r482_B_0_), .ZN(n5046) );
  AOI22_X2 U4550 ( .A1(N347), .A2(n4811), .B1(N347), .B2(n4808), .ZN(n1088) );
  AOI22_X2 U4551 ( .A1(N348), .A2(n4811), .B1(opa_r1[1]), .B2(n4809), .ZN(
        n1092) );
  AOI22_X2 U4552 ( .A1(N349), .A2(n4811), .B1(opa_r1[2]), .B2(n4807), .ZN(
        n1093) );
  AOI22_X2 U4553 ( .A1(N350), .A2(n4811), .B1(opa_r1[3]), .B2(n4809), .ZN(
        n1094) );
  AOI22_X2 U4554 ( .A1(N351), .A2(n4811), .B1(opa_r1[4]), .B2(n4807), .ZN(
        n1095) );
  AOI22_X2 U4555 ( .A1(N352), .A2(n4811), .B1(opa_r1[5]), .B2(n4808), .ZN(
        n1096) );
  AOI22_X2 U4556 ( .A1(N353), .A2(n4811), .B1(opa_r1[6]), .B2(n4809), .ZN(
        n1097) );
  AOI22_X2 U4557 ( .A1(N354), .A2(n4811), .B1(opa_r1[7]), .B2(n4807), .ZN(
        n1098) );
  AOI22_X2 U4558 ( .A1(N355), .A2(n4811), .B1(opa_r1[8]), .B2(n4808), .ZN(
        n1099) );
  AOI22_X2 U4559 ( .A1(N356), .A2(n4811), .B1(opa_r1[9]), .B2(n4809), .ZN(
        n1100) );
  AOI22_X2 U4560 ( .A1(N357), .A2(n4811), .B1(opa_r1[10]), .B2(n4809), .ZN(
        n1101) );
  AOI22_X2 U4561 ( .A1(N358), .A2(n4812), .B1(opa_r1[11]), .B2(n4809), .ZN(
        n1102) );
  AOI22_X2 U4562 ( .A1(N359), .A2(n4812), .B1(opa_r1[12]), .B2(n4809), .ZN(
        n1103) );
  AOI22_X2 U4563 ( .A1(N360), .A2(n4812), .B1(opa_r1[13]), .B2(n4809), .ZN(
        n1104) );
  AOI22_X2 U4564 ( .A1(N361), .A2(n4812), .B1(opa_r1[14]), .B2(n4809), .ZN(
        n1105) );
  AOI22_X2 U4565 ( .A1(N362), .A2(n4812), .B1(opa_r1[15]), .B2(n4809), .ZN(
        n1106) );
  AOI22_X2 U4566 ( .A1(N363), .A2(n4812), .B1(opa_r1[16]), .B2(n4809), .ZN(
        n1107) );
  AOI22_X2 U4567 ( .A1(N364), .A2(n4812), .B1(opa_r1[17]), .B2(n4809), .ZN(
        n1108) );
  AOI22_X2 U4568 ( .A1(N365), .A2(n4812), .B1(opa_r1[18]), .B2(n4809), .ZN(
        n1109) );
  AOI22_X2 U4569 ( .A1(N366), .A2(n4812), .B1(opa_r1[19]), .B2(n4809), .ZN(
        n1110) );
  AOI22_X2 U4570 ( .A1(N367), .A2(n4812), .B1(opa_r1[20]), .B2(n4808), .ZN(
        n1111) );
  AOI22_X2 U4571 ( .A1(N368), .A2(n4812), .B1(opa_r1[21]), .B2(n4808), .ZN(
        n1112) );
  AOI22_X2 U4572 ( .A1(N369), .A2(n4813), .B1(opa_r1[22]), .B2(n4808), .ZN(
        n1113) );
  AOI22_X2 U4573 ( .A1(N370), .A2(n4813), .B1(opa_r1[23]), .B2(n4808), .ZN(
        n1114) );
  AOI22_X2 U4574 ( .A1(N371), .A2(n4813), .B1(opa_r1[24]), .B2(n4808), .ZN(
        n1115) );
  AOI22_X2 U4575 ( .A1(N372), .A2(n4813), .B1(opa_r1[25]), .B2(n4808), .ZN(
        n1116) );
  AOI22_X2 U4576 ( .A1(N373), .A2(n4813), .B1(opa_r1[26]), .B2(n4808), .ZN(
        n1117) );
  AOI22_X2 U4577 ( .A1(N374), .A2(n4813), .B1(opa_r1[27]), .B2(n4808), .ZN(
        n1118) );
  AOI22_X2 U4578 ( .A1(N375), .A2(n4813), .B1(opa_r1[28]), .B2(n4808), .ZN(
        n1119) );
  AOI22_X2 U4579 ( .A1(N376), .A2(n4813), .B1(opa_r1[29]), .B2(n4808), .ZN(
        n1120) );
  AOI22_X2 U4580 ( .A1(N377), .A2(n4813), .B1(opa_r1[30]), .B2(n4808), .ZN(
        n1121) );
  AOI22_X2 U4581 ( .A1(N378), .A2(n4813), .B1(opa_r1[31]), .B2(n4807), .ZN(
        n1122) );
  AOI22_X2 U4582 ( .A1(N379), .A2(n4813), .B1(opa_r1[32]), .B2(n4807), .ZN(
        n1123) );
  AOI22_X2 U4583 ( .A1(N380), .A2(n4813), .B1(opa_r1[33]), .B2(n4807), .ZN(
        n1124) );
  AOI22_X2 U4584 ( .A1(N381), .A2(n4813), .B1(opa_r1[34]), .B2(n4807), .ZN(
        n1125) );
  AOI22_X2 U4585 ( .A1(N382), .A2(n4813), .B1(opa_r1[35]), .B2(n4807), .ZN(
        n1126) );
  AOI22_X2 U4586 ( .A1(N383), .A2(n4813), .B1(opa_r1[36]), .B2(n4807), .ZN(
        n1127) );
  AOI22_X2 U4587 ( .A1(N384), .A2(n4813), .B1(opa_r1[37]), .B2(n4807), .ZN(
        n1128) );
  AOI22_X2 U4588 ( .A1(N385), .A2(n4813), .B1(opa_r1[38]), .B2(n4807), .ZN(
        n1129) );
  AOI22_X2 U4589 ( .A1(N386), .A2(n4813), .B1(opa_r1[39]), .B2(n4807), .ZN(
        n1130) );
  AOI22_X2 U4590 ( .A1(N387), .A2(n4813), .B1(opa_r1[40]), .B2(n4807), .ZN(
        n1131) );
  AOI22_X2 U4591 ( .A1(N388), .A2(n4813), .B1(opa_r1[41]), .B2(n4807), .ZN(
        n1132) );
  AOI22_X2 U4592 ( .A1(N389), .A2(n4813), .B1(opa_r1[42]), .B2(n4807), .ZN(
        n1133) );
  AOI22_X2 U4593 ( .A1(N390), .A2(n4813), .B1(opa_r1[43]), .B2(n1091), .ZN(
        n1134) );
  AOI22_X2 U4594 ( .A1(N391), .A2(n4811), .B1(opa_r1[44]), .B2(n1091), .ZN(
        n1135) );
  AOI22_X2 U4595 ( .A1(N392), .A2(n4812), .B1(opa_r1[45]), .B2(n4807), .ZN(
        n1136) );
  INV_X4 U4596 ( .A(n2085), .ZN(n5942) );
  INV_X4 U4597 ( .A(n2078), .ZN(n5943) );
  INV_X4 U4598 ( .A(n1716), .ZN(n5944) );
  INV_X4 U4599 ( .A(N312), .ZN(n5945) );
  INV_X4 U4600 ( .A(N311), .ZN(n5946) );
  INV_X4 U4601 ( .A(N310), .ZN(n5947) );
  INV_X4 U4602 ( .A(N309), .ZN(n5948) );
  INV_X4 U4603 ( .A(N308), .ZN(n5949) );
  INV_X4 U4604 ( .A(n1033), .ZN(u6_N101) );
  INV_X4 U4605 ( .A(N306), .ZN(n5950) );
  INV_X4 U4606 ( .A(N305), .ZN(n5951) );
  INV_X4 U4607 ( .A(n955), .ZN(u6_N98) );
  INV_X4 U4608 ( .A(N303), .ZN(n5952) );
  INV_X4 U4609 ( .A(N302), .ZN(n5953) );
  INV_X4 U4610 ( .A(n960), .ZN(u6_N95) );
  INV_X4 U4611 ( .A(N300), .ZN(n5954) );
  INV_X4 U4612 ( .A(N299), .ZN(n5955) );
  INV_X4 U4613 ( .A(n965), .ZN(u6_N92) );
  INV_X4 U4614 ( .A(N297), .ZN(n5956) );
  INV_X4 U4615 ( .A(N296), .ZN(n5957) );
  INV_X4 U4616 ( .A(N295), .ZN(n5958) );
  INV_X4 U4617 ( .A(n971), .ZN(u6_N88) );
  INV_X4 U4618 ( .A(N293), .ZN(n5959) );
  INV_X4 U4619 ( .A(n974), .ZN(u6_N86) );
  INV_X4 U4620 ( .A(N291), .ZN(n5960) );
  INV_X4 U4621 ( .A(N290), .ZN(n5961) );
  INV_X4 U4622 ( .A(N289), .ZN(n5962) );
  INV_X4 U4623 ( .A(N288), .ZN(n5963) );
  INV_X4 U4624 ( .A(N287), .ZN(n5964) );
  INV_X4 U4625 ( .A(N286), .ZN(n5965) );
  INV_X4 U4626 ( .A(n986), .ZN(u6_N79) );
  INV_X4 U4627 ( .A(N284), .ZN(n5966) );
  INV_X4 U4628 ( .A(N283), .ZN(n5967) );
  INV_X4 U4629 ( .A(N282), .ZN(n5968) );
  INV_X4 U4630 ( .A(n993), .ZN(u6_N75) );
  INV_X4 U4631 ( .A(n994), .ZN(u6_N74) );
  INV_X4 U4632 ( .A(N279), .ZN(n5969) );
  INV_X4 U4633 ( .A(N278), .ZN(n5970) );
  INV_X4 U4634 ( .A(N277), .ZN(n5971) );
  INV_X4 U4635 ( .A(n1001), .ZN(u6_N70) );
  INV_X4 U4636 ( .A(N275), .ZN(n5972) );
  INV_X4 U4637 ( .A(n1004), .ZN(u6_N68) );
  INV_X4 U4638 ( .A(N273), .ZN(n5973) );
  INV_X4 U4639 ( .A(N272), .ZN(n5974) );
  INV_X4 U4640 ( .A(n1009), .ZN(u6_N65) );
  INV_X4 U4641 ( .A(N270), .ZN(n5975) );
  INV_X4 U4642 ( .A(n1012), .ZN(u6_N63) );
  INV_X4 U4643 ( .A(n1013), .ZN(u6_N62) );
  INV_X4 U4644 ( .A(n1304), .ZN(u6_N61) );
  INV_X4 U4645 ( .A(N266), .ZN(n5976) );
  INV_X4 U4646 ( .A(n1016), .ZN(u6_N59) );
  INV_X4 U4647 ( .A(N264), .ZN(n5977) );
  INV_X4 U4648 ( .A(n1019), .ZN(u6_N57) );
  INV_X4 U4649 ( .A(N262), .ZN(n5978) );
  INV_X4 U4650 ( .A(n1022), .ZN(u6_N55) );
  INV_X4 U4651 ( .A(n1974), .ZN(n5979) );
  INV_X4 U4652 ( .A(n1136), .ZN(n5980) );
  INV_X4 U4653 ( .A(n1135), .ZN(n5981) );
  INV_X4 U4654 ( .A(n1134), .ZN(n5982) );
  INV_X4 U4655 ( .A(n1133), .ZN(n5983) );
  INV_X4 U4656 ( .A(n1132), .ZN(n5984) );
  INV_X4 U4657 ( .A(n1131), .ZN(n5985) );
  INV_X4 U4658 ( .A(n1130), .ZN(n5986) );
  INV_X4 U4659 ( .A(n1129), .ZN(n5987) );
  INV_X4 U4660 ( .A(n1128), .ZN(n5988) );
  INV_X4 U4661 ( .A(n1127), .ZN(n5989) );
  INV_X4 U4662 ( .A(n1126), .ZN(n5990) );
  INV_X4 U4663 ( .A(n1125), .ZN(n5991) );
  INV_X4 U4664 ( .A(n1124), .ZN(n5992) );
  INV_X4 U4665 ( .A(n1123), .ZN(n5993) );
  INV_X4 U4666 ( .A(n1122), .ZN(n5994) );
  INV_X4 U4667 ( .A(n1121), .ZN(n5995) );
  INV_X4 U4668 ( .A(n1120), .ZN(n5996) );
  INV_X4 U4669 ( .A(n1119), .ZN(n5997) );
  INV_X4 U4670 ( .A(n1118), .ZN(n5998) );
  INV_X4 U4671 ( .A(n1117), .ZN(n5999) );
  INV_X4 U4672 ( .A(n1116), .ZN(n6000) );
  INV_X4 U4673 ( .A(n1115), .ZN(n6001) );
  INV_X4 U4674 ( .A(n1114), .ZN(n6002) );
  INV_X4 U4675 ( .A(n1113), .ZN(n6003) );
  INV_X4 U4676 ( .A(n1112), .ZN(n6004) );
  INV_X4 U4677 ( .A(n1111), .ZN(n6005) );
  INV_X4 U4678 ( .A(n1110), .ZN(n6006) );
  INV_X4 U4679 ( .A(n1109), .ZN(n6007) );
  INV_X4 U4680 ( .A(n1108), .ZN(n6008) );
  INV_X4 U4681 ( .A(n1107), .ZN(n6009) );
  INV_X4 U4682 ( .A(n1106), .ZN(n6010) );
  INV_X4 U4683 ( .A(n1105), .ZN(n6011) );
  INV_X4 U4684 ( .A(n1104), .ZN(n6012) );
  INV_X4 U4685 ( .A(n1103), .ZN(n6013) );
  INV_X4 U4686 ( .A(n1102), .ZN(n6014) );
  INV_X4 U4687 ( .A(n1101), .ZN(n6015) );
  INV_X4 U4688 ( .A(n1100), .ZN(n6016) );
  INV_X4 U4689 ( .A(n1099), .ZN(n6017) );
  INV_X4 U4690 ( .A(n1098), .ZN(n6018) );
  INV_X4 U4691 ( .A(n1097), .ZN(n6019) );
  INV_X4 U4692 ( .A(n1096), .ZN(n6020) );
  INV_X4 U4693 ( .A(n1095), .ZN(n6021) );
  INV_X4 U4694 ( .A(n1094), .ZN(n6022) );
  INV_X4 U4695 ( .A(n1093), .ZN(n6023) );
  INV_X4 U4696 ( .A(n1092), .ZN(n6024) );
  INV_X4 U4697 ( .A(N561), .ZN(n6025) );
  INV_X4 U4698 ( .A(N560), .ZN(n6026) );
  INV_X4 U4699 ( .A(N559), .ZN(n6027) );
  INV_X4 U4700 ( .A(N558), .ZN(n6028) );
  INV_X4 U4701 ( .A(N557), .ZN(n6029) );
  INV_X4 U4702 ( .A(N556), .ZN(n6030) );
  INV_X4 U4703 ( .A(N555), .ZN(n6031) );
  INV_X4 U4704 ( .A(N554), .ZN(n6032) );
  INV_X4 U4705 ( .A(N553), .ZN(n6033) );
  INV_X4 U4706 ( .A(N552), .ZN(n6034) );
  INV_X4 U4707 ( .A(N551), .ZN(n6035) );
  INV_X4 U4708 ( .A(N550), .ZN(n6036) );
  INV_X4 U4709 ( .A(N549), .ZN(n6037) );
  INV_X4 U4710 ( .A(N548), .ZN(n6038) );
  INV_X4 U4711 ( .A(N547), .ZN(n6039) );
  INV_X4 U4712 ( .A(N546), .ZN(n6040) );
  INV_X4 U4713 ( .A(N545), .ZN(n6041) );
  INV_X4 U4714 ( .A(N544), .ZN(n6042) );
  INV_X4 U4715 ( .A(N543), .ZN(n6043) );
  INV_X4 U4716 ( .A(N542), .ZN(n6044) );
  INV_X4 U4717 ( .A(N541), .ZN(n6045) );
  INV_X4 U4718 ( .A(N540), .ZN(n6046) );
  INV_X4 U4719 ( .A(N539), .ZN(n6047) );
  INV_X4 U4720 ( .A(N538), .ZN(n6048) );
  INV_X4 U4721 ( .A(N537), .ZN(n6049) );
  INV_X4 U4722 ( .A(N536), .ZN(n6050) );
  INV_X4 U4723 ( .A(N535), .ZN(n6051) );
  INV_X4 U4724 ( .A(N534), .ZN(n6052) );
  INV_X4 U4725 ( .A(N533), .ZN(n6053) );
  INV_X4 U4726 ( .A(N532), .ZN(n6054) );
  INV_X4 U4727 ( .A(N531), .ZN(n6055) );
  INV_X4 U4728 ( .A(N530), .ZN(n6056) );
  INV_X4 U4729 ( .A(N529), .ZN(n6057) );
  INV_X4 U4730 ( .A(N528), .ZN(n6058) );
  INV_X4 U4731 ( .A(N527), .ZN(n6059) );
  INV_X4 U4732 ( .A(N526), .ZN(n6060) );
  INV_X4 U4733 ( .A(N525), .ZN(n6061) );
  INV_X4 U4734 ( .A(N524), .ZN(n6062) );
  INV_X4 U4735 ( .A(N523), .ZN(n6063) );
  INV_X4 U4736 ( .A(N522), .ZN(n6064) );
  INV_X4 U4737 ( .A(N521), .ZN(n6065) );
  INV_X4 U4738 ( .A(N520), .ZN(n6066) );
  INV_X4 U4739 ( .A(N519), .ZN(n6067) );
  INV_X4 U4740 ( .A(N518), .ZN(n6068) );
  INV_X4 U4741 ( .A(N517), .ZN(n6069) );
  INV_X4 U4742 ( .A(N516), .ZN(n6070) );
  INV_X4 U4743 ( .A(N515), .ZN(n6071) );
  INV_X4 U4744 ( .A(N514), .ZN(n6072) );
  INV_X4 U4745 ( .A(N513), .ZN(n6073) );
  INV_X4 U4746 ( .A(N512), .ZN(n6074) );
  INV_X4 U4747 ( .A(N511), .ZN(n6075) );
  INV_X4 U4748 ( .A(N510), .ZN(n6076) );
  INV_X4 U4749 ( .A(N509), .ZN(n6077) );
  INV_X4 U4750 ( .A(N508), .ZN(n6078) );
  INV_X4 U4751 ( .A(N507), .ZN(n6079) );
  INV_X4 U4752 ( .A(N506), .ZN(n6080) );
  INV_X4 U4753 ( .A(N505), .ZN(n6081) );
  INV_X4 U4754 ( .A(u2_exp_ovf_d_1_), .ZN(n6082) );
  INV_X4 U4755 ( .A(n602), .ZN(u2_gt_141_B_11_) );
  INV_X4 U4756 ( .A(n1036), .ZN(n6083) );
  INV_X4 U4757 ( .A(u2_N16), .ZN(n6084) );
  INV_X4 U4758 ( .A(n1037), .ZN(n6085) );
  INV_X4 U4759 ( .A(n1048), .ZN(u2_lt_131_A_9_) );
  INV_X4 U4760 ( .A(n1038), .ZN(n6086) );
  INV_X4 U4761 ( .A(n1049), .ZN(u2_lt_131_A_8_) );
  INV_X4 U4762 ( .A(n1039), .ZN(n6087) );
  INV_X4 U4763 ( .A(n1050), .ZN(u2_lt_131_A_7_) );
  INV_X4 U4764 ( .A(n1040), .ZN(n6088) );
  INV_X4 U4765 ( .A(n1051), .ZN(u2_lt_131_A_6_) );
  INV_X4 U4766 ( .A(n1041), .ZN(n6089) );
  INV_X4 U4767 ( .A(n1052), .ZN(u2_lt_131_A_5_) );
  INV_X4 U4768 ( .A(n1042), .ZN(n6090) );
  INV_X4 U4769 ( .A(u2_N10), .ZN(n6091) );
  INV_X4 U4770 ( .A(n1043), .ZN(n6092) );
  INV_X4 U4771 ( .A(u2_N9), .ZN(n6093) );
  INV_X4 U4772 ( .A(n1044), .ZN(n6094) );
  INV_X4 U4773 ( .A(u2_N8), .ZN(n6095) );
  INV_X4 U4774 ( .A(n1045), .ZN(n6096) );
  INV_X4 U4775 ( .A(u2_N7), .ZN(n6097) );
  INV_X4 U4776 ( .A(n1046), .ZN(n6098) );
  INV_X4 U4777 ( .A(u2_N28), .ZN(n6099) );
  INV_X4 U4778 ( .A(u2_N22), .ZN(n6100) );
  INV_X4 U4779 ( .A(u2_N21), .ZN(n6101) );
  INV_X4 U4780 ( .A(u2_N20), .ZN(n6102) );
  INV_X4 U4781 ( .A(u2_N19), .ZN(n6103) );
  INV_X4 U4782 ( .A(n1270), .ZN(n6104) );
  INV_X4 U4783 ( .A(n1219), .ZN(n6105) );
  INV_X4 U4784 ( .A(n1220), .ZN(n6106) );
  INV_X4 U4785 ( .A(n1221), .ZN(n6107) );
  INV_X4 U4786 ( .A(n1222), .ZN(n6108) );
  INV_X4 U4787 ( .A(n1223), .ZN(n6109) );
  INV_X4 U4788 ( .A(n1224), .ZN(n6110) );
  INV_X4 U4789 ( .A(n1226), .ZN(n6111) );
  INV_X4 U4790 ( .A(n1227), .ZN(n6112) );
  INV_X4 U4791 ( .A(n1228), .ZN(n6113) );
  INV_X4 U4792 ( .A(n1229), .ZN(n6114) );
  INV_X4 U4793 ( .A(n1230), .ZN(n6115) );
  INV_X4 U4794 ( .A(n1231), .ZN(n6116) );
  INV_X4 U4795 ( .A(n1232), .ZN(n6117) );
  INV_X4 U4796 ( .A(n1233), .ZN(n6118) );
  INV_X4 U4797 ( .A(n1234), .ZN(n6119) );
  INV_X4 U4798 ( .A(n1235), .ZN(n6120) );
  INV_X4 U4799 ( .A(n1237), .ZN(n6121) );
  INV_X4 U4800 ( .A(n1238), .ZN(n6122) );
  INV_X4 U4801 ( .A(n1239), .ZN(n6123) );
  INV_X4 U4802 ( .A(n1240), .ZN(n6124) );
  INV_X4 U4803 ( .A(n1241), .ZN(n6125) );
  INV_X4 U4804 ( .A(n1242), .ZN(n6126) );
  INV_X4 U4805 ( .A(n1243), .ZN(n6127) );
  INV_X4 U4806 ( .A(n1244), .ZN(n6128) );
  INV_X4 U4807 ( .A(n1245), .ZN(n6129) );
  INV_X4 U4808 ( .A(n1246), .ZN(n6130) );
  INV_X4 U4809 ( .A(n1248), .ZN(n6131) );
  INV_X4 U4810 ( .A(n1249), .ZN(n6132) );
  INV_X4 U4811 ( .A(n1250), .ZN(n6133) );
  INV_X4 U4812 ( .A(n1251), .ZN(n6134) );
  INV_X4 U4813 ( .A(n1252), .ZN(n6135) );
  INV_X4 U4814 ( .A(n1253), .ZN(n6136) );
  INV_X4 U4815 ( .A(n1254), .ZN(n6137) );
  INV_X4 U4816 ( .A(n1255), .ZN(n6138) );
  INV_X4 U4817 ( .A(n1256), .ZN(n6139) );
  INV_X4 U4818 ( .A(n1257), .ZN(n6140) );
  INV_X4 U4819 ( .A(n1259), .ZN(n6141) );
  INV_X4 U4820 ( .A(n1260), .ZN(n6142) );
  INV_X4 U4821 ( .A(n1261), .ZN(n6143) );
  INV_X4 U4822 ( .A(n1262), .ZN(n6144) );
  INV_X4 U4823 ( .A(n1263), .ZN(n6145) );
  INV_X4 U4824 ( .A(n1264), .ZN(n6146) );
  INV_X4 U4825 ( .A(n1265), .ZN(n6147) );
  INV_X4 U4826 ( .A(n1266), .ZN(n6148) );
  INV_X4 U4827 ( .A(n1267), .ZN(n6149) );
  INV_X4 U4828 ( .A(n1268), .ZN(n6150) );
  INV_X4 U4829 ( .A(n1213), .ZN(n6151) );
  INV_X4 U4830 ( .A(n1215), .ZN(n6152) );
  INV_X4 U4831 ( .A(n1216), .ZN(n6153) );
  INV_X4 U4832 ( .A(n1217), .ZN(n6154) );
  INV_X4 U4833 ( .A(n1218), .ZN(n6155) );
  INV_X4 U4834 ( .A(n1225), .ZN(n6156) );
  INV_X4 U4835 ( .A(n1236), .ZN(n6157) );
  INV_X4 U4836 ( .A(n1247), .ZN(n6158) );
  INV_X4 U4837 ( .A(n1258), .ZN(n6159) );
  INV_X4 U4838 ( .A(n1269), .ZN(n6160) );
  INV_X4 U4839 ( .A(n1739), .ZN(n6161) );
  INV_X4 U4840 ( .A(n1737), .ZN(n6162) );
  INV_X4 U4841 ( .A(u4_exp_next_mi_11_), .ZN(n6163) );
  INV_X4 U4842 ( .A(n2087), .ZN(u4_sub_466_A_10_) );
  INV_X4 U4843 ( .A(n2083), .ZN(u4_sub_466_A_9_) );
  INV_X4 U4844 ( .A(u4_exp_next_mi_8_), .ZN(n6164) );
  INV_X4 U4845 ( .A(u4_exp_next_mi_7_), .ZN(n6165) );
  INV_X4 U4846 ( .A(n2115), .ZN(u4_sub_466_A_6_) );
  INV_X4 U4847 ( .A(n2110), .ZN(u4_sub_466_A_5_) );
  INV_X4 U4848 ( .A(u4_exp_next_mi_4_), .ZN(n6166) );
  INV_X4 U4849 ( .A(u4_exp_next_mi_3_), .ZN(n6167) );
  INV_X4 U4850 ( .A(u4_exp_next_mi_2_), .ZN(n6168) );
  INV_X4 U4851 ( .A(u4_exp_next_mi_1_), .ZN(n6169) );
  INV_X4 U4852 ( .A(u4_exp_next_mi_0_), .ZN(n6170) );
  INV_X4 U4853 ( .A(n3953), .ZN(n6171) );
  INV_X4 U4854 ( .A(n755), .ZN(n6172) );
  INV_X4 U4855 ( .A(n754), .ZN(n6173) );
  INV_X4 U4856 ( .A(n741), .ZN(n6174) );
  INV_X4 U4857 ( .A(n740), .ZN(n6175) );
  INV_X4 U4858 ( .A(n749), .ZN(n6176) );
  INV_X4 U4859 ( .A(n748), .ZN(n6177) );
  INV_X4 U4860 ( .A(n715), .ZN(n6178) );
  INV_X4 U4861 ( .A(n714), .ZN(n6179) );
  INV_X4 U4862 ( .A(n731), .ZN(n6180) );
  INV_X4 U4863 ( .A(n730), .ZN(n6181) );
  INV_X4 U4864 ( .A(n667), .ZN(n6182) );
  INV_X4 U4865 ( .A(n666), .ZN(n6183) );
  INV_X4 U4866 ( .A(n723), .ZN(n6184) );
  INV_X4 U4867 ( .A(n722), .ZN(n6185) );
  INV_X4 U4868 ( .A(n647), .ZN(n6186) );
  INV_X4 U4869 ( .A(n646), .ZN(n6187) );
  INV_X4 U4870 ( .A(n705), .ZN(n6188) );
  INV_X4 U4871 ( .A(n704), .ZN(n6189) );
  INV_X4 U4872 ( .A(n697), .ZN(n6190) );
  INV_X4 U4873 ( .A(n696), .ZN(n6191) );
  INV_X4 U4874 ( .A(n679), .ZN(n6192) );
  INV_X4 U4875 ( .A(n678), .ZN(n6193) );
  INV_X4 U4876 ( .A(n687), .ZN(n6194) );
  INV_X4 U4877 ( .A(n686), .ZN(n6195) );
  INV_X4 U4878 ( .A(n671), .ZN(n6196) );
  INV_X4 U4879 ( .A(n670), .ZN(n6197) );
  INV_X4 U4880 ( .A(n661), .ZN(n6198) );
  INV_X4 U4881 ( .A(n660), .ZN(n6199) );
  INV_X4 U4882 ( .A(n753), .ZN(n6200) );
  INV_X4 U4883 ( .A(n752), .ZN(n6201) );
  INV_X4 U4884 ( .A(n719), .ZN(n6202) );
  INV_X4 U4885 ( .A(n718), .ZN(n6203) );
  INV_X4 U4886 ( .A(n745), .ZN(n6204) );
  INV_X4 U4887 ( .A(n744), .ZN(n6205) );
  INV_X4 U4888 ( .A(n709), .ZN(n6206) );
  INV_X4 U4889 ( .A(n708), .ZN(n6207) );
  INV_X4 U4890 ( .A(n737), .ZN(n6208) );
  INV_X4 U4891 ( .A(n736), .ZN(n6209) );
  INV_X4 U4892 ( .A(n710), .ZN(n6210) );
  INV_X4 U4893 ( .A(n711), .ZN(n6211) );
  INV_X4 U4894 ( .A(n727), .ZN(n6212) );
  INV_X4 U4895 ( .A(n726), .ZN(n6213) );
  INV_X4 U4896 ( .A(n651), .ZN(n6214) );
  INV_X4 U4897 ( .A(n650), .ZN(n6215) );
  INV_X4 U4898 ( .A(n701), .ZN(n6216) );
  INV_X4 U4899 ( .A(n700), .ZN(n6217) );
  INV_X4 U4900 ( .A(n693), .ZN(n6218) );
  INV_X4 U4901 ( .A(n692), .ZN(n6219) );
  INV_X4 U4902 ( .A(n683), .ZN(n6220) );
  INV_X4 U4903 ( .A(n682), .ZN(n6221) );
  INV_X4 U4904 ( .A(n675), .ZN(n6222) );
  INV_X4 U4905 ( .A(n674), .ZN(n6223) );
  INV_X4 U4906 ( .A(n665), .ZN(n6224) );
  INV_X4 U4907 ( .A(n664), .ZN(n6225) );
  INV_X4 U4908 ( .A(n657), .ZN(n6226) );
  INV_X4 U4909 ( .A(n656), .ZN(n6227) );
  INV_X4 U4910 ( .A(n751), .ZN(n6228) );
  INV_X4 U4911 ( .A(n750), .ZN(n6229) );
  INV_X4 U4912 ( .A(n717), .ZN(n6230) );
  INV_X4 U4913 ( .A(n716), .ZN(n6231) );
  INV_X4 U4914 ( .A(n743), .ZN(n6232) );
  INV_X4 U4915 ( .A(n742), .ZN(n6233) );
  INV_X4 U4916 ( .A(n707), .ZN(n6234) );
  INV_X4 U4917 ( .A(n706), .ZN(n6235) );
  INV_X4 U4918 ( .A(n735), .ZN(n6236) );
  INV_X4 U4919 ( .A(n734), .ZN(n6237) );
  INV_X4 U4920 ( .A(n689), .ZN(n6238) );
  INV_X4 U4921 ( .A(n688), .ZN(n6239) );
  INV_X4 U4922 ( .A(n725), .ZN(n6240) );
  INV_X4 U4923 ( .A(n724), .ZN(n6241) );
  INV_X4 U4924 ( .A(n649), .ZN(n6242) );
  INV_X4 U4925 ( .A(n648), .ZN(n6243) );
  INV_X4 U4926 ( .A(n699), .ZN(n6244) );
  INV_X4 U4927 ( .A(n698), .ZN(n6245) );
  INV_X4 U4928 ( .A(n691), .ZN(n6246) );
  INV_X4 U4929 ( .A(n690), .ZN(n6247) );
  INV_X4 U4930 ( .A(n681), .ZN(n6248) );
  INV_X4 U4931 ( .A(n680), .ZN(n6249) );
  INV_X4 U4932 ( .A(n673), .ZN(n6250) );
  INV_X4 U4933 ( .A(n672), .ZN(n6251) );
  INV_X4 U4934 ( .A(n663), .ZN(n6252) );
  INV_X4 U4935 ( .A(n662), .ZN(n6253) );
  INV_X4 U4936 ( .A(n655), .ZN(n6254) );
  INV_X4 U4937 ( .A(n654), .ZN(n6255) );
  INV_X4 U4938 ( .A(n747), .ZN(n6256) );
  INV_X4 U4939 ( .A(n746), .ZN(n6257) );
  INV_X4 U4940 ( .A(n713), .ZN(n6258) );
  INV_X4 U4941 ( .A(n712), .ZN(n6259) );
  INV_X4 U4942 ( .A(n739), .ZN(n6260) );
  INV_X4 U4943 ( .A(n738), .ZN(n6261) );
  INV_X4 U4944 ( .A(n732), .ZN(n6262) );
  INV_X4 U4945 ( .A(n733), .ZN(n6263) );
  INV_X4 U4946 ( .A(n703), .ZN(n6264) );
  INV_X4 U4947 ( .A(n702), .ZN(n6265) );
  INV_X4 U4948 ( .A(n729), .ZN(n6266) );
  INV_X4 U4949 ( .A(n728), .ZN(n6267) );
  INV_X4 U4950 ( .A(n653), .ZN(n6268) );
  INV_X4 U4951 ( .A(n652), .ZN(n6269) );
  INV_X4 U4952 ( .A(n721), .ZN(n6270) );
  INV_X4 U4953 ( .A(n720), .ZN(n6271) );
  INV_X4 U4954 ( .A(n645), .ZN(n6272) );
  INV_X4 U4955 ( .A(n644), .ZN(n6273) );
  INV_X4 U4956 ( .A(n695), .ZN(n6274) );
  INV_X4 U4957 ( .A(n694), .ZN(n6275) );
  INV_X4 U4958 ( .A(n685), .ZN(n6276) );
  INV_X4 U4959 ( .A(n684), .ZN(n6277) );
  INV_X4 U4960 ( .A(n677), .ZN(n6278) );
  INV_X4 U4961 ( .A(n676), .ZN(n6279) );
  INV_X4 U4962 ( .A(n669), .ZN(n6280) );
  INV_X4 U4963 ( .A(n668), .ZN(n6281) );
  INV_X4 U4964 ( .A(n659), .ZN(n6282) );
  INV_X4 U4965 ( .A(n658), .ZN(n6283) );
  INV_X4 U4966 ( .A(n941), .ZN(n6284) );
  INV_X4 U4967 ( .A(n803), .ZN(n6285) );
  INV_X4 U4968 ( .A(n862), .ZN(n6286) );
  INV_X4 U4969 ( .A(n812), .ZN(n6287) );
  INV_X4 U4970 ( .A(n842), .ZN(n6288) );
  INV_X4 U4971 ( .A(n840), .ZN(n6289) );
  INV_X4 U4972 ( .A(n818), .ZN(n6290) );
  INV_X4 U4973 ( .A(n887), .ZN(n6291) );
  INV_X4 U4974 ( .A(n820), .ZN(n6292) );
  INV_X4 U4975 ( .A(n939), .ZN(n6293) );
  INV_X4 U4976 ( .A(n872), .ZN(n6294) );
  INV_X4 U4977 ( .A(n868), .ZN(n6295) );
  INV_X4 U4978 ( .A(n864), .ZN(n6296) );
  INV_X4 U4979 ( .A(n898), .ZN(n6297) );
  INV_X4 U4980 ( .A(n876), .ZN(n6298) );
  INV_X4 U4981 ( .A(n810), .ZN(n6299) );
  INV_X4 U4982 ( .A(u1_exp_lt_27), .ZN(n6300) );
  INV_X4 U4983 ( .A(n912), .ZN(n6302) );
  INV_X4 U4984 ( .A(n938), .ZN(n6303) );
  INV_X4 U4985 ( .A(n918), .ZN(n6304) );
  INV_X4 U4986 ( .A(n774), .ZN(n6305) );
  INV_X4 U4987 ( .A(n775), .ZN(n6306) );
  INV_X4 U4988 ( .A(n776), .ZN(n6307) );
  INV_X4 U4989 ( .A(n879), .ZN(n6308) );
  INV_X4 U4990 ( .A(n4070), .ZN(n6309) );
  INV_X4 U4991 ( .A(n1056), .ZN(n6310) );
  INV_X4 U4992 ( .A(n1057), .ZN(n6311) );
  INV_X4 U4993 ( .A(n779), .ZN(n6312) );
  INV_X4 U4994 ( .A(n780), .ZN(n6313) );
  INV_X4 U4995 ( .A(n4149), .ZN(n6314) );
  INV_X4 U4996 ( .A(n4150), .ZN(n6315) );
  INV_X4 U4997 ( .A(n4151), .ZN(n6316) );
  INV_X4 U4998 ( .A(n4152), .ZN(n6317) );
  INV_X4 U4999 ( .A(n4153), .ZN(n6318) );
  INV_X4 U5000 ( .A(n4154), .ZN(n6319) );
  INV_X4 U5001 ( .A(n4155), .ZN(n6320) );
  INV_X4 U5002 ( .A(n4156), .ZN(n6321) );
  INV_X4 U5003 ( .A(n1062), .ZN(n6322) );
  INV_X4 U5004 ( .A(n900), .ZN(n6323) );
  INV_X4 U5005 ( .A(n901), .ZN(n6324) );
  INV_X4 U5006 ( .A(n902), .ZN(n6325) );
  INV_X4 U5007 ( .A(n916), .ZN(n6326) );
  INV_X4 U5008 ( .A(n1064), .ZN(n6327) );
  INV_X4 U5009 ( .A(n917), .ZN(n6328) );
  INV_X4 U5010 ( .A(n921), .ZN(n6329) );
  INV_X4 U5011 ( .A(n1066), .ZN(n6330) );
  INV_X4 U5012 ( .A(n924), .ZN(n6331) );
  INV_X4 U5013 ( .A(n1071), .ZN(n6332) );
  INV_X4 U5014 ( .A(n1075), .ZN(n6333) );
  INV_X4 U5015 ( .A(n926), .ZN(n6334) );
  INV_X4 U5016 ( .A(n925), .ZN(n6335) );
  INV_X4 U5017 ( .A(n1078), .ZN(n6336) );
  INV_X4 U5018 ( .A(n927), .ZN(n6337) );
  INV_X4 U5019 ( .A(n1079), .ZN(n6338) );
  INV_X4 U5020 ( .A(n928), .ZN(n6339) );
  INV_X4 U5021 ( .A(n1081), .ZN(n6340) );
  INV_X4 U5022 ( .A(n1083), .ZN(n6341) );
  INV_X4 U5023 ( .A(n930), .ZN(n6342) );
  INV_X4 U5024 ( .A(n877), .ZN(n6343) );
  INV_X4 U5025 ( .A(n929), .ZN(n6344) );
  INV_X4 U5026 ( .A(n1084), .ZN(n6345) );
  INV_X4 U5027 ( .A(n932), .ZN(n6346) );
  INV_X4 U5028 ( .A(n931), .ZN(n6347) );
  INV_X4 U5029 ( .A(n870), .ZN(n6348) );
  INV_X4 U5030 ( .A(n4348), .ZN(n6349) );
  INV_X4 U5031 ( .A(n949), .ZN(n6350) );
  INV_X4 U5032 ( .A(n583), .ZN(n6351) );
  INV_X4 U5033 ( .A(n4123), .ZN(n6352) );
  INV_X4 U5034 ( .A(n1413), .ZN(n6353) );
  INV_X4 U5035 ( .A(n1448), .ZN(n6354) );
  INV_X4 U5036 ( .A(n1354), .ZN(n6355) );
  INV_X4 U5037 ( .A(n1418), .ZN(n6356) );
  INV_X4 U5038 ( .A(n1435), .ZN(n6357) );
  INV_X4 U5039 ( .A(n1361), .ZN(n6358) );
  INV_X4 U5040 ( .A(n1412), .ZN(n6359) );
  INV_X4 U5041 ( .A(n1357), .ZN(n6360) );
  INV_X4 U5042 ( .A(n1355), .ZN(n6361) );
  INV_X4 U5043 ( .A(n1391), .ZN(n6362) );
  INV_X4 U5044 ( .A(n1369), .ZN(n6363) );
  INV_X4 U5045 ( .A(n1427), .ZN(n6364) );
  INV_X4 U5046 ( .A(n1396), .ZN(n6365) );
  INV_X4 U5047 ( .A(n1283), .ZN(n6366) );
  INV_X4 U5048 ( .A(n1402), .ZN(n6367) );
  INV_X4 U5049 ( .A(n1430), .ZN(n6368) );
  INV_X4 U5050 ( .A(n1375), .ZN(n6369) );
  INV_X4 U5051 ( .A(n1378), .ZN(n6370) );
  INV_X4 U5052 ( .A(n1374), .ZN(n6371) );
  INV_X4 U5053 ( .A(n948), .ZN(n6372) );
  INV_X4 U5054 ( .A(u6_N52), .ZN(n6373) );
  INV_X4 U5055 ( .A(n798), .ZN(n6374) );
  INV_X4 U5056 ( .A(n801), .ZN(n6375) );
  INV_X4 U5057 ( .A(u4_N5830), .ZN(n6376) );
  INV_X4 U5058 ( .A(n2032), .ZN(n6377) );
  INV_X4 U5059 ( .A(n2033), .ZN(n6378) );
  INV_X4 U5060 ( .A(n1671), .ZN(n6379) );
  INV_X4 U5061 ( .A(n1088), .ZN(n6380) );
  INV_X4 U5062 ( .A(n1308), .ZN(n6381) );
  INV_X4 U5063 ( .A(n1473), .ZN(n6382) );
  INV_X4 U5064 ( .A(n1919), .ZN(n6383) );
  INV_X4 U5065 ( .A(n2268), .ZN(n6384) );
  INV_X4 U5066 ( .A(n1963), .ZN(n6385) );
  INV_X4 U5067 ( .A(n1978), .ZN(n6386) );
  INV_X4 U5068 ( .A(n1480), .ZN(n6388) );
  INV_X4 U5069 ( .A(n1925), .ZN(n6389) );
  INV_X4 U5070 ( .A(n247), .ZN(n6391) );
  INV_X4 U5071 ( .A(n1475), .ZN(n6392) );
  INV_X4 U5072 ( .A(n1211), .ZN(n6393) );
  INV_X4 U5073 ( .A(n1212), .ZN(n6394) );
  INV_X4 U5074 ( .A(n943), .ZN(n6395) );
  INV_X4 U5075 ( .A(n944), .ZN(n6396) );
  INV_X4 U5076 ( .A(n1767), .ZN(n6397) );
  INV_X4 U5077 ( .A(n1485), .ZN(n6398) );
  INV_X4 U5078 ( .A(n1477), .ZN(n6399) );
  INV_X4 U5079 ( .A(n1685), .ZN(n6400) );
  INV_X4 U5080 ( .A(n1708), .ZN(n6401) );
  INV_X4 U5081 ( .A(n1705), .ZN(n6402) );
  INV_X4 U5082 ( .A(n1741), .ZN(n6403) );
  INV_X4 U5083 ( .A(fract_denorm[0]), .ZN(n6404) );
  INV_X4 U5084 ( .A(n405), .ZN(n6405) );
  INV_X4 U5085 ( .A(u4_N6188), .ZN(n6406) );
  INV_X4 U5086 ( .A(fract_denorm[1]), .ZN(n6407) );
  INV_X4 U5087 ( .A(n560), .ZN(n6408) );
  INV_X4 U5088 ( .A(n478), .ZN(n6409) );
  INV_X4 U5089 ( .A(fract_denorm[5]), .ZN(n6410) );
  INV_X4 U5090 ( .A(n505), .ZN(n6411) );
  INV_X4 U5091 ( .A(fract_denorm[7]), .ZN(n6412) );
  INV_X4 U5092 ( .A(n504), .ZN(n6413) );
  INV_X4 U5093 ( .A(fract_denorm[8]), .ZN(n6414) );
  INV_X4 U5094 ( .A(fract_denorm[9]), .ZN(n6415) );
  INV_X4 U5095 ( .A(n486), .ZN(n6416) );
  INV_X4 U5096 ( .A(n341), .ZN(n6417) );
  INV_X4 U5097 ( .A(fract_denorm[12]), .ZN(n6418) );
  INV_X4 U5098 ( .A(n386), .ZN(n6419) );
  INV_X4 U5099 ( .A(n546), .ZN(n6420) );
  INV_X4 U5100 ( .A(fract_denorm[13]), .ZN(n6421) );
  INV_X4 U5101 ( .A(n328), .ZN(n6422) );
  INV_X4 U5102 ( .A(n532), .ZN(n6423) );
  INV_X4 U5103 ( .A(fract_denorm[15]), .ZN(n6424) );
  INV_X4 U5104 ( .A(n336), .ZN(n6425) );
  INV_X4 U5105 ( .A(fract_denorm[16]), .ZN(n6426) );
  INV_X4 U5106 ( .A(fract_denorm[17]), .ZN(n6427) );
  INV_X4 U5107 ( .A(fract_denorm[18]), .ZN(n6428) );
  INV_X4 U5108 ( .A(fract_denorm[19]), .ZN(n6429) );
  INV_X4 U5109 ( .A(fract_denorm[20]), .ZN(n6430) );
  INV_X4 U5110 ( .A(fract_denorm[21]), .ZN(n6431) );
  INV_X4 U5111 ( .A(n2168), .ZN(n6432) );
  INV_X4 U5112 ( .A(fract_denorm[23]), .ZN(n6433) );
  INV_X4 U5113 ( .A(n420), .ZN(n6434) );
  INV_X4 U5114 ( .A(fract_denorm[24]), .ZN(n6435) );
  INV_X4 U5115 ( .A(n331), .ZN(n6436) );
  INV_X4 U5116 ( .A(fract_denorm[26]), .ZN(n6437) );
  INV_X4 U5117 ( .A(fract_denorm[28]), .ZN(n6438) );
  INV_X4 U5118 ( .A(fract_denorm[29]), .ZN(n6439) );
  INV_X4 U5119 ( .A(fract_denorm[30]), .ZN(n6440) );
  INV_X4 U5120 ( .A(fract_denorm[31]), .ZN(n6441) );
  INV_X4 U5121 ( .A(fract_denorm[32]), .ZN(n6442) );
  INV_X4 U5122 ( .A(fract_denorm[33]), .ZN(n6443) );
  INV_X4 U5123 ( .A(fract_denorm[34]), .ZN(n6444) );
  INV_X4 U5124 ( .A(fract_denorm[35]), .ZN(n6445) );
  INV_X4 U5125 ( .A(n392), .ZN(n6446) );
  INV_X4 U5126 ( .A(fract_denorm[38]), .ZN(n6447) );
  INV_X4 U5127 ( .A(n496), .ZN(n6448) );
  INV_X4 U5128 ( .A(fract_denorm[39]), .ZN(n6449) );
  INV_X4 U5129 ( .A(fract_denorm[40]), .ZN(n6450) );
  INV_X4 U5130 ( .A(n579), .ZN(n6451) );
  INV_X4 U5131 ( .A(n443), .ZN(n6452) );
  INV_X4 U5132 ( .A(fract_denorm[42]), .ZN(n6453) );
  INV_X4 U5133 ( .A(n301), .ZN(n6454) );
  INV_X4 U5134 ( .A(n365), .ZN(n6455) );
  INV_X4 U5135 ( .A(fract_denorm[44]), .ZN(n6456) );
  INV_X4 U5136 ( .A(fract_denorm[45]), .ZN(n6457) );
  INV_X4 U5137 ( .A(n366), .ZN(n6458) );
  INV_X4 U5138 ( .A(fract_denorm[47]), .ZN(n6459) );
  INV_X4 U5139 ( .A(fract_denorm[48]), .ZN(n6460) );
  INV_X4 U5140 ( .A(n368), .ZN(n6461) );
  INV_X4 U5141 ( .A(fract_denorm[49]), .ZN(n6462) );
  INV_X4 U5142 ( .A(fract_denorm[50]), .ZN(n6463) );
  INV_X4 U5143 ( .A(n374), .ZN(n6464) );
  INV_X4 U5144 ( .A(fract_denorm[51]), .ZN(n6465) );
  INV_X4 U5145 ( .A(n507), .ZN(n6466) );
  INV_X4 U5146 ( .A(fract_denorm[52]), .ZN(n6467) );
  INV_X4 U5147 ( .A(fract_denorm[54]), .ZN(n6468) );
  INV_X4 U5148 ( .A(n375), .ZN(n6469) );
  INV_X4 U5149 ( .A(fract_denorm[55]), .ZN(n6470) );
  INV_X4 U5150 ( .A(fract_denorm[56]), .ZN(n6471) );
  INV_X4 U5151 ( .A(fract_denorm[57]), .ZN(n6472) );
  INV_X4 U5152 ( .A(fract_denorm[59]), .ZN(n6473) );
  INV_X4 U5153 ( .A(fract_denorm[61]), .ZN(n6474) );
  INV_X4 U5154 ( .A(n376), .ZN(n6475) );
  INV_X4 U5155 ( .A(fract_denorm[62]), .ZN(n6476) );
  INV_X4 U5156 ( .A(fract_denorm[64]), .ZN(n6477) );
  INV_X4 U5157 ( .A(n310), .ZN(n6478) );
  INV_X4 U5158 ( .A(n308), .ZN(n6479) );
  INV_X4 U5159 ( .A(fract_denorm[67]), .ZN(n6480) );
  INV_X4 U5160 ( .A(n298), .ZN(n6481) );
  INV_X4 U5161 ( .A(fract_denorm[69]), .ZN(n6482) );
  INV_X4 U5162 ( .A(n319), .ZN(n6483) );
  INV_X4 U5163 ( .A(n297), .ZN(n6484) );
  INV_X4 U5164 ( .A(n315), .ZN(n6485) );
  INV_X4 U5165 ( .A(fract_denorm[72]), .ZN(n6486) );
  INV_X4 U5166 ( .A(n529), .ZN(n6487) );
  INV_X4 U5167 ( .A(n313), .ZN(n6488) );
  INV_X4 U5168 ( .A(fract_denorm[75]), .ZN(n6489) );
  INV_X4 U5169 ( .A(n345), .ZN(n6490) );
  INV_X4 U5170 ( .A(fract_denorm[77]), .ZN(n6491) );
  INV_X4 U5171 ( .A(n312), .ZN(n6492) );
  INV_X4 U5172 ( .A(fract_denorm[78]), .ZN(n6493) );
  INV_X4 U5173 ( .A(fract_denorm[80]), .ZN(n6494) );
  INV_X4 U5174 ( .A(n351), .ZN(n6495) );
  INV_X4 U5175 ( .A(fract_denorm[81]), .ZN(n6496) );
  INV_X4 U5176 ( .A(n400), .ZN(n6497) );
  INV_X4 U5177 ( .A(fract_denorm[83]), .ZN(n6498) );
  INV_X4 U5178 ( .A(n349), .ZN(n6499) );
  INV_X4 U5179 ( .A(fract_denorm[84]), .ZN(n6500) );
  INV_X4 U5180 ( .A(fract_denorm[85]), .ZN(n6501) );
  INV_X4 U5181 ( .A(fract_denorm[87]), .ZN(n6502) );
  INV_X4 U5182 ( .A(n416), .ZN(n6503) );
  INV_X4 U5183 ( .A(n454), .ZN(n6504) );
  INV_X4 U5184 ( .A(fract_denorm[89]), .ZN(n6505) );
  INV_X4 U5185 ( .A(fract_denorm[91]), .ZN(n6506) );
  INV_X4 U5186 ( .A(fract_denorm[92]), .ZN(n6507) );
  INV_X4 U5187 ( .A(fract_denorm[93]), .ZN(n6508) );
  INV_X4 U5188 ( .A(n354), .ZN(n6509) );
  INV_X4 U5189 ( .A(fract_denorm[95]), .ZN(n6510) );
  INV_X4 U5190 ( .A(n432), .ZN(n6511) );
  INV_X4 U5191 ( .A(fract_denorm[97]), .ZN(n6512) );
  INV_X4 U5192 ( .A(n465), .ZN(n6513) );
  INV_X4 U5193 ( .A(fract_denorm[98]), .ZN(n6514) );
  INV_X4 U5194 ( .A(fract_denorm[99]), .ZN(n6515) );
  INV_X4 U5195 ( .A(fract_denorm[100]), .ZN(n6516) );
  INV_X4 U5196 ( .A(fract_denorm[101]), .ZN(n6517) );
  INV_X4 U5197 ( .A(fract_denorm[103]), .ZN(n6518) );
  INV_X4 U5198 ( .A(fract_denorm[104]), .ZN(n6519) );
  INV_X4 U5199 ( .A(u4_exp_in_mi1_11_), .ZN(n6520) );
  INV_X4 U5200 ( .A(u4_exp_in_pl1_8_), .ZN(n6521) );
  INV_X4 U5201 ( .A(u4_exp_in_pl1_7_), .ZN(n6522) );
  INV_X4 U5202 ( .A(u4_exp_in_pl1_4_), .ZN(n6523) );
  INV_X4 U5203 ( .A(u4_exp_in_pl1_3_), .ZN(n6524) );
  INV_X4 U5204 ( .A(u4_exp_in_pl1_2_), .ZN(n6525) );
  INV_X4 U5205 ( .A(u4_exp_in_pl1_1_), .ZN(n6526) );
  INV_X4 U5206 ( .A(n1735), .ZN(n6527) );
  INV_X4 U5207 ( .A(n1732), .ZN(n6528) );
  INV_X4 U5208 ( .A(u4_N5831), .ZN(n6529) );
  INV_X4 u4_sub_471_U23 ( .A(u4_fi_ldz_mi1_0_), .ZN(u4_sub_471_n14) );
  INV_X4 u4_sub_471_U22 ( .A(u4_fi_ldz_mi1_6_), .ZN(u4_sub_471_n13) );
  INV_X4 u4_sub_471_U21 ( .A(u4_fi_ldz_mi1_5_), .ZN(u4_sub_471_n12) );
  INV_X4 u4_sub_471_U20 ( .A(u4_fi_ldz_mi1_4_), .ZN(u4_sub_471_n11) );
  INV_X4 u4_sub_471_U19 ( .A(u4_fi_ldz_mi1_3_), .ZN(u4_sub_471_n10) );
  INV_X4 u4_sub_471_U18 ( .A(u4_fi_ldz_mi1_2_), .ZN(u4_sub_471_n9) );
  INV_X4 u4_sub_471_U17 ( .A(u4_fi_ldz_mi1_1_), .ZN(u4_sub_471_n8) );
  INV_X4 u4_sub_471_U16 ( .A(n4823), .ZN(u4_sub_471_n7) );
  XNOR2_X2 u4_sub_471_U15 ( .A(u4_sub_471_n14), .B(n4823), .ZN(
        u4_exp_fix_divb[0]) );
  NAND2_X2 u4_sub_471_U14 ( .A1(u4_fi_ldz_mi1_0_), .A2(u4_sub_471_n7), .ZN(
        u4_sub_471_carry_1_) );
  INV_X4 u4_sub_471_U13 ( .A(u4_sub_471_carry_9_), .ZN(u4_sub_471_n6) );
  INV_X4 u4_sub_471_U12 ( .A(n4428), .ZN(u4_sub_471_n5) );
  XNOR2_X2 u4_sub_471_U11 ( .A(n4428), .B(u4_sub_471_carry_9_), .ZN(
        u4_exp_fix_divb[9]) );
  NAND2_X2 u4_sub_471_U10 ( .A1(u4_sub_471_n5), .A2(u4_sub_471_n6), .ZN(
        u4_sub_471_carry_10_) );
  INV_X4 u4_sub_471_U9 ( .A(u4_sub_471_carry_8_), .ZN(u4_sub_471_n4) );
  INV_X4 u4_sub_471_U8 ( .A(n4369), .ZN(u4_sub_471_n3) );
  XNOR2_X2 u4_sub_471_U7 ( .A(n4369), .B(u4_sub_471_carry_8_), .ZN(
        u4_exp_fix_divb[8]) );
  NAND2_X2 u4_sub_471_U6 ( .A1(u4_sub_471_n3), .A2(u4_sub_471_n4), .ZN(
        u4_sub_471_carry_9_) );
  INV_X4 u4_sub_471_U5 ( .A(u4_sub_471_carry_7_), .ZN(u4_sub_471_n2) );
  INV_X4 u4_sub_471_U4 ( .A(n4359), .ZN(u4_sub_471_n1) );
  XNOR2_X2 u4_sub_471_U3 ( .A(n4359), .B(u4_sub_471_carry_7_), .ZN(
        u4_exp_fix_divb[7]) );
  NAND2_X2 u4_sub_471_U2 ( .A1(u4_sub_471_n1), .A2(u4_sub_471_n2), .ZN(
        u4_sub_471_carry_8_) );
  XNOR2_X2 u4_sub_471_U1 ( .A(n4875), .B(u4_sub_471_carry_10_), .ZN(
        u4_exp_fix_divb[10]) );
  FA_X1 u4_sub_471_U2_1 ( .A(n4368), .B(u4_sub_471_n8), .CI(
        u4_sub_471_carry_1_), .CO(u4_sub_471_carry_2_), .S(u4_exp_fix_divb[1])
         );
  FA_X1 u4_sub_471_U2_2 ( .A(exp_r[2]), .B(u4_sub_471_n9), .CI(
        u4_sub_471_carry_2_), .CO(u4_sub_471_carry_3_), .S(u4_exp_fix_divb[2])
         );
  FA_X1 u4_sub_471_U2_3 ( .A(exp_r[3]), .B(u4_sub_471_n10), .CI(
        u4_sub_471_carry_3_), .CO(u4_sub_471_carry_4_), .S(u4_exp_fix_divb[3])
         );
  FA_X1 u4_sub_471_U2_4 ( .A(n4399), .B(u4_sub_471_n11), .CI(
        u4_sub_471_carry_4_), .CO(u4_sub_471_carry_5_), .S(u4_exp_fix_divb[4])
         );
  FA_X1 u4_sub_471_U2_5 ( .A(n4370), .B(u4_sub_471_n12), .CI(
        u4_sub_471_carry_5_), .CO(u4_sub_471_carry_6_), .S(u4_exp_fix_divb[5])
         );
  FA_X1 u4_sub_471_U2_6 ( .A(n4382), .B(u4_sub_471_n13), .CI(
        u4_sub_471_carry_6_), .CO(u4_sub_471_carry_7_), .S(u4_exp_fix_divb[6])
         );
  INV_X4 u4_sub_470_U23 ( .A(u4_fi_ldz_mi1_0_), .ZN(u4_sub_470_n14) );
  INV_X4 u4_sub_470_U22 ( .A(u4_fi_ldz_mi22[1]), .ZN(u4_sub_470_n13) );
  INV_X4 u4_sub_470_U21 ( .A(u4_fi_ldz_mi22[2]), .ZN(u4_sub_470_n12) );
  INV_X4 u4_sub_470_U20 ( .A(u4_fi_ldz_mi22[3]), .ZN(u4_sub_470_n11) );
  INV_X4 u4_sub_470_U19 ( .A(u4_fi_ldz_mi22[4]), .ZN(u4_sub_470_n10) );
  INV_X4 u4_sub_470_U18 ( .A(u4_fi_ldz_mi22[5]), .ZN(u4_sub_470_n9) );
  INV_X4 u4_sub_470_U17 ( .A(u4_fi_ldz_mi22[6]), .ZN(u4_sub_470_n8) );
  INV_X4 u4_sub_470_U16 ( .A(n4823), .ZN(u4_sub_470_n7) );
  XNOR2_X2 u4_sub_470_U15 ( .A(u4_sub_470_n14), .B(n4823), .ZN(
        u4_exp_fix_diva[0]) );
  NAND2_X2 u4_sub_470_U14 ( .A1(u4_fi_ldz_mi1_0_), .A2(u4_sub_470_n7), .ZN(
        u4_sub_470_carry_1_) );
  INV_X4 u4_sub_470_U13 ( .A(u4_sub_470_carry_9_), .ZN(u4_sub_470_n6) );
  INV_X4 u4_sub_470_U12 ( .A(n4428), .ZN(u4_sub_470_n5) );
  XNOR2_X2 u4_sub_470_U11 ( .A(n4428), .B(u4_sub_470_carry_9_), .ZN(
        u4_exp_fix_diva[9]) );
  NAND2_X2 u4_sub_470_U10 ( .A1(u4_sub_470_n5), .A2(u4_sub_470_n6), .ZN(
        u4_sub_470_carry_10_) );
  INV_X4 u4_sub_470_U9 ( .A(u4_sub_470_carry_8_), .ZN(u4_sub_470_n4) );
  INV_X4 u4_sub_470_U8 ( .A(n4369), .ZN(u4_sub_470_n3) );
  XNOR2_X2 u4_sub_470_U7 ( .A(n4369), .B(u4_sub_470_carry_8_), .ZN(
        u4_exp_fix_diva[8]) );
  NAND2_X2 u4_sub_470_U6 ( .A1(u4_sub_470_n3), .A2(u4_sub_470_n4), .ZN(
        u4_sub_470_carry_9_) );
  INV_X4 u4_sub_470_U5 ( .A(u4_sub_470_carry_7_), .ZN(u4_sub_470_n2) );
  INV_X4 u4_sub_470_U4 ( .A(n4359), .ZN(u4_sub_470_n1) );
  XNOR2_X2 u4_sub_470_U3 ( .A(n4359), .B(u4_sub_470_carry_7_), .ZN(
        u4_exp_fix_diva[7]) );
  NAND2_X2 u4_sub_470_U2 ( .A1(u4_sub_470_n1), .A2(u4_sub_470_n2), .ZN(
        u4_sub_470_carry_8_) );
  XNOR2_X2 u4_sub_470_U1 ( .A(n4875), .B(u4_sub_470_carry_10_), .ZN(
        u4_exp_fix_diva[10]) );
  FA_X1 u4_sub_470_U2_1 ( .A(n4368), .B(u4_sub_470_n13), .CI(
        u4_sub_470_carry_1_), .CO(u4_sub_470_carry_2_), .S(u4_exp_fix_diva[1])
         );
  FA_X1 u4_sub_470_U2_2 ( .A(exp_r[2]), .B(u4_sub_470_n12), .CI(
        u4_sub_470_carry_2_), .CO(u4_sub_470_carry_3_), .S(u4_exp_fix_diva[2])
         );
  FA_X1 u4_sub_470_U2_3 ( .A(exp_r[3]), .B(u4_sub_470_n11), .CI(
        u4_sub_470_carry_3_), .CO(u4_sub_470_carry_4_), .S(u4_exp_fix_diva[3])
         );
  FA_X1 u4_sub_470_U2_4 ( .A(n4399), .B(u4_sub_470_n10), .CI(
        u4_sub_470_carry_4_), .CO(u4_sub_470_carry_5_), .S(u4_exp_fix_diva[4])
         );
  FA_X1 u4_sub_470_U2_5 ( .A(n4370), .B(u4_sub_470_n9), .CI(
        u4_sub_470_carry_5_), .CO(u4_sub_470_carry_6_), .S(u4_exp_fix_diva[5])
         );
  FA_X1 u4_sub_470_U2_6 ( .A(n4382), .B(u4_sub_470_n8), .CI(
        u4_sub_470_carry_6_), .CO(u4_sub_470_carry_7_), .S(u4_exp_fix_diva[6])
         );
  INV_X1 u4_add_462_U2 ( .A(u4_exp_out_0_), .ZN(u4_exp_out_pl1_0_) );
  XOR2_X1 u4_add_462_U1 ( .A(u4_add_462_carry[10]), .B(u4_exp_out_10_), .Z(
        u4_exp_out_pl1_10_) );
  HA_X1 u4_add_462_U1_1_1 ( .A(u4_exp_out_1_), .B(u4_exp_out_0_), .CO(
        u4_add_462_carry[2]), .S(u4_exp_out_pl1_1_) );
  HA_X1 u4_add_462_U1_1_2 ( .A(u4_exp_out_2_), .B(u4_add_462_carry[2]), .CO(
        u4_add_462_carry[3]), .S(u4_exp_out_pl1_2_) );
  HA_X1 u4_add_462_U1_1_3 ( .A(u4_exp_out_3_), .B(u4_add_462_carry[3]), .CO(
        u4_add_462_carry[4]), .S(u4_exp_out_pl1_3_) );
  HA_X1 u4_add_462_U1_1_4 ( .A(u4_exp_out_4_), .B(u4_add_462_carry[4]), .CO(
        u4_add_462_carry[5]), .S(u4_exp_out_pl1_4_) );
  HA_X1 u4_add_462_U1_1_5 ( .A(u4_exp_out_5_), .B(u4_add_462_carry[5]), .CO(
        u4_add_462_carry[6]), .S(u4_exp_out_pl1_5_) );
  HA_X1 u4_add_462_U1_1_6 ( .A(u4_exp_out_6_), .B(u4_add_462_carry[6]), .CO(
        u4_add_462_carry[7]), .S(u4_exp_out_pl1_6_) );
  HA_X1 u4_add_462_U1_1_7 ( .A(u4_exp_out_7_), .B(u4_add_462_carry[7]), .CO(
        u4_add_462_carry[8]), .S(u4_exp_out_pl1_7_) );
  HA_X1 u4_add_462_U1_1_8 ( .A(u4_exp_out_8_), .B(u4_add_462_carry[8]), .CO(
        u4_add_462_carry[9]), .S(u4_exp_out_pl1_8_) );
  HA_X1 u4_add_462_U1_1_9 ( .A(u4_exp_out_9_), .B(u4_add_462_carry[9]), .CO(
        u4_add_462_carry[10]), .S(u4_exp_out_pl1_9_) );
  INV_X1 u4_sll_452_U269 ( .A(u4_shift_left[8]), .ZN(u4_sll_452_n55) );
  OR2_X1 u4_sll_452_U268 ( .A1(u4_sll_452_n1), .A2(u4_shift_left[7]), .ZN(
        u4_sll_452_n88) );
  NAND2_X1 u4_sll_452_U267 ( .A1(u4_shift_left[7]), .A2(u4_sll_452_n1), .ZN(
        u4_sll_452_n90) );
  INV_X1 u4_sll_452_U266 ( .A(u4_sll_452_n90), .ZN(u4_sll_452_n89) );
  AOI21_X1 u4_sll_452_U265 ( .B1(u4_shift_left[0]), .B2(u4_sll_452_n88), .A(
        u4_sll_452_n89), .ZN(u4_sll_452_SHMAG_0_) );
  AND2_X1 u4_sll_452_U264 ( .A1(fract_denorm[0]), .A2(u4_sll_452_SHMAG_0_), 
        .ZN(u4_sll_452_ML_int_1__0_) );
  AOI21_X1 u4_sll_452_U263 ( .B1(u4_shift_left[1]), .B2(u4_sll_452_n88), .A(
        u4_sll_452_n89), .ZN(u4_sll_452_SHMAG_1_) );
  AND2_X1 u4_sll_452_U262 ( .A1(u4_sll_452_ML_int_1__0_), .A2(
        u4_sll_452_SHMAG_1_), .ZN(u4_sll_452_ML_int_2__0_) );
  AND2_X1 u4_sll_452_U261 ( .A1(u4_sll_452_ML_int_1__1_), .A2(
        u4_sll_452_SHMAG_1_), .ZN(u4_sll_452_ML_int_2__1_) );
  AOI21_X1 u4_sll_452_U260 ( .B1(u4_shift_left[2]), .B2(u4_sll_452_n88), .A(
        u4_sll_452_n89), .ZN(u4_sll_452_SHMAG_2_) );
  AND2_X1 u4_sll_452_U259 ( .A1(u4_sll_452_ML_int_2__0_), .A2(
        u4_sll_452_SHMAG_2_), .ZN(u4_sll_452_ML_int_3__0_) );
  AND2_X1 u4_sll_452_U258 ( .A1(u4_sll_452_ML_int_2__1_), .A2(
        u4_sll_452_SHMAG_2_), .ZN(u4_sll_452_ML_int_3__1_) );
  AND2_X1 u4_sll_452_U257 ( .A1(u4_sll_452_ML_int_2__2_), .A2(
        u4_sll_452_SHMAG_2_), .ZN(u4_sll_452_ML_int_3__2_) );
  AND2_X1 u4_sll_452_U256 ( .A1(u4_sll_452_ML_int_2__3_), .A2(
        u4_sll_452_SHMAG_2_), .ZN(u4_sll_452_ML_int_3__3_) );
  AOI21_X1 u4_sll_452_U255 ( .B1(u4_shift_left[3]), .B2(u4_sll_452_n88), .A(
        u4_sll_452_n89), .ZN(u4_sll_452_SHMAG_3_) );
  AND2_X1 u4_sll_452_U254 ( .A1(u4_sll_452_ML_int_3__0_), .A2(u4_sll_452_n18), 
        .ZN(u4_sll_452_ML_int_4__0_) );
  AND2_X1 u4_sll_452_U253 ( .A1(u4_sll_452_ML_int_3__1_), .A2(u4_sll_452_n18), 
        .ZN(u4_sll_452_ML_int_4__1_) );
  AND2_X1 u4_sll_452_U252 ( .A1(u4_sll_452_ML_int_3__2_), .A2(u4_sll_452_n18), 
        .ZN(u4_sll_452_ML_int_4__2_) );
  AND2_X1 u4_sll_452_U251 ( .A1(u4_sll_452_ML_int_3__3_), .A2(u4_sll_452_n18), 
        .ZN(u4_sll_452_ML_int_4__3_) );
  AND2_X1 u4_sll_452_U250 ( .A1(u4_sll_452_ML_int_3__4_), .A2(u4_sll_452_n18), 
        .ZN(u4_sll_452_ML_int_4__4_) );
  AND2_X1 u4_sll_452_U249 ( .A1(u4_sll_452_ML_int_3__5_), .A2(u4_sll_452_n18), 
        .ZN(u4_sll_452_ML_int_4__5_) );
  AND2_X1 u4_sll_452_U248 ( .A1(u4_sll_452_ML_int_3__6_), .A2(u4_sll_452_n25), 
        .ZN(u4_sll_452_ML_int_4__6_) );
  AND2_X1 u4_sll_452_U247 ( .A1(u4_sll_452_ML_int_3__7_), .A2(u4_sll_452_n18), 
        .ZN(u4_sll_452_ML_int_4__7_) );
  AOI21_X1 u4_sll_452_U246 ( .B1(u4_shift_left[4]), .B2(u4_sll_452_n88), .A(
        u4_sll_452_n89), .ZN(u4_sll_452_SHMAG_4_) );
  AND2_X1 u4_sll_452_U245 ( .A1(u4_sll_452_ML_int_4__0_), .A2(u4_sll_452_n37), 
        .ZN(u4_sll_452_ML_int_5__0_) );
  AND2_X1 u4_sll_452_U244 ( .A1(u4_sll_452_ML_int_4__10_), .A2(u4_sll_452_n27), 
        .ZN(u4_sll_452_ML_int_5__10_) );
  AND2_X1 u4_sll_452_U243 ( .A1(u4_sll_452_ML_int_4__11_), .A2(u4_sll_452_n27), 
        .ZN(u4_sll_452_ML_int_5__11_) );
  AND2_X1 u4_sll_452_U242 ( .A1(u4_sll_452_ML_int_4__12_), .A2(u4_sll_452_n27), 
        .ZN(u4_sll_452_ML_int_5__12_) );
  AND2_X1 u4_sll_452_U241 ( .A1(u4_sll_452_ML_int_4__13_), .A2(u4_sll_452_n27), 
        .ZN(u4_sll_452_ML_int_5__13_) );
  AND2_X1 u4_sll_452_U240 ( .A1(u4_sll_452_ML_int_4__14_), .A2(u4_sll_452_n27), 
        .ZN(u4_sll_452_ML_int_5__14_) );
  AND2_X1 u4_sll_452_U239 ( .A1(u4_sll_452_ML_int_4__15_), .A2(u4_sll_452_n27), 
        .ZN(u4_sll_452_ML_int_5__15_) );
  AND2_X1 u4_sll_452_U238 ( .A1(u4_sll_452_ML_int_4__1_), .A2(u4_sll_452_n28), 
        .ZN(u4_sll_452_ML_int_5__1_) );
  AND2_X1 u4_sll_452_U237 ( .A1(u4_sll_452_ML_int_4__2_), .A2(u4_sll_452_n28), 
        .ZN(u4_sll_452_ML_int_5__2_) );
  AND2_X1 u4_sll_452_U236 ( .A1(u4_sll_452_ML_int_4__3_), .A2(u4_sll_452_n27), 
        .ZN(u4_sll_452_ML_int_5__3_) );
  AND2_X1 u4_sll_452_U235 ( .A1(u4_sll_452_ML_int_4__4_), .A2(u4_sll_452_n27), 
        .ZN(u4_sll_452_ML_int_5__4_) );
  AND2_X1 u4_sll_452_U234 ( .A1(u4_sll_452_ML_int_4__5_), .A2(u4_sll_452_n27), 
        .ZN(u4_sll_452_ML_int_5__5_) );
  AND2_X1 u4_sll_452_U233 ( .A1(u4_sll_452_ML_int_4__6_), .A2(u4_sll_452_n27), 
        .ZN(u4_sll_452_ML_int_5__6_) );
  AND2_X1 u4_sll_452_U232 ( .A1(u4_sll_452_ML_int_4__7_), .A2(u4_sll_452_n28), 
        .ZN(u4_sll_452_ML_int_5__7_) );
  AND2_X1 u4_sll_452_U231 ( .A1(u4_sll_452_ML_int_4__8_), .A2(u4_sll_452_n27), 
        .ZN(u4_sll_452_ML_int_5__8_) );
  AND2_X1 u4_sll_452_U230 ( .A1(u4_sll_452_ML_int_4__9_), .A2(u4_sll_452_n28), 
        .ZN(u4_sll_452_ML_int_5__9_) );
  NAND2_X1 u4_sll_452_U229 ( .A1(u4_shift_left[5]), .A2(u4_sll_452_n88), .ZN(
        u4_sll_452_n91) );
  NAND2_X1 u4_sll_452_U228 ( .A1(u4_sll_452_n90), .A2(u4_sll_452_n91), .ZN(
        u4_sll_452_temp_int_SH_5_) );
  NAND2_X1 u4_sll_452_U227 ( .A1(u4_sll_452_ML_int_5__0_), .A2(u4_sll_452_n41), 
        .ZN(u4_sll_452_n87) );
  INV_X1 u4_sll_452_U226 ( .A(u4_sll_452_n87), .ZN(u4_sll_452_ML_int_6__0_) );
  NAND2_X1 u4_sll_452_U225 ( .A1(u4_sll_452_ML_int_5__10_), .A2(u4_sll_452_n42), .ZN(u4_sll_452_n86) );
  INV_X1 u4_sll_452_U224 ( .A(u4_sll_452_n86), .ZN(u4_sll_452_ML_int_6__10_)
         );
  NAND2_X1 u4_sll_452_U223 ( .A1(u4_sll_452_ML_int_5__11_), .A2(u4_sll_452_n42), .ZN(u4_sll_452_n85) );
  INV_X1 u4_sll_452_U222 ( .A(u4_sll_452_n85), .ZN(u4_sll_452_ML_int_6__11_)
         );
  NAND2_X1 u4_sll_452_U221 ( .A1(u4_sll_452_ML_int_5__12_), .A2(u4_sll_452_n42), .ZN(u4_sll_452_n84) );
  INV_X1 u4_sll_452_U220 ( .A(u4_sll_452_n84), .ZN(u4_sll_452_ML_int_6__12_)
         );
  NAND2_X1 u4_sll_452_U219 ( .A1(u4_sll_452_ML_int_5__13_), .A2(u4_sll_452_n42), .ZN(u4_sll_452_n83) );
  INV_X1 u4_sll_452_U218 ( .A(u4_sll_452_n83), .ZN(u4_sll_452_ML_int_6__13_)
         );
  NAND2_X1 u4_sll_452_U217 ( .A1(u4_sll_452_ML_int_5__14_), .A2(u4_sll_452_n42), .ZN(u4_sll_452_n82) );
  INV_X1 u4_sll_452_U216 ( .A(u4_sll_452_n82), .ZN(u4_sll_452_ML_int_6__14_)
         );
  NAND2_X1 u4_sll_452_U215 ( .A1(u4_sll_452_ML_int_5__15_), .A2(u4_sll_452_n42), .ZN(u4_sll_452_n81) );
  INV_X1 u4_sll_452_U214 ( .A(u4_sll_452_n81), .ZN(u4_sll_452_ML_int_6__15_)
         );
  NAND2_X1 u4_sll_452_U213 ( .A1(u4_sll_452_ML_int_5__16_), .A2(u4_sll_452_n42), .ZN(u4_sll_452_n80) );
  INV_X1 u4_sll_452_U212 ( .A(u4_sll_452_n80), .ZN(u4_sll_452_ML_int_6__16_)
         );
  NAND2_X1 u4_sll_452_U211 ( .A1(u4_sll_452_ML_int_5__17_), .A2(u4_sll_452_n42), .ZN(u4_sll_452_n79) );
  INV_X1 u4_sll_452_U210 ( .A(u4_sll_452_n79), .ZN(u4_sll_452_ML_int_6__17_)
         );
  NAND2_X1 u4_sll_452_U209 ( .A1(u4_sll_452_ML_int_5__18_), .A2(u4_sll_452_n42), .ZN(u4_sll_452_n78) );
  INV_X1 u4_sll_452_U208 ( .A(u4_sll_452_n78), .ZN(u4_sll_452_ML_int_6__18_)
         );
  NAND2_X1 u4_sll_452_U207 ( .A1(u4_sll_452_ML_int_5__19_), .A2(u4_sll_452_n42), .ZN(u4_sll_452_n77) );
  INV_X1 u4_sll_452_U206 ( .A(u4_sll_452_n77), .ZN(u4_sll_452_ML_int_6__19_)
         );
  NAND2_X1 u4_sll_452_U205 ( .A1(u4_sll_452_ML_int_5__1_), .A2(u4_sll_452_n43), 
        .ZN(u4_sll_452_n76) );
  INV_X1 u4_sll_452_U204 ( .A(u4_sll_452_n76), .ZN(u4_sll_452_ML_int_6__1_) );
  NAND2_X1 u4_sll_452_U203 ( .A1(u4_sll_452_ML_int_5__20_), .A2(u4_sll_452_n42), .ZN(u4_sll_452_n75) );
  INV_X1 u4_sll_452_U202 ( .A(u4_sll_452_n75), .ZN(u4_sll_452_ML_int_6__20_)
         );
  NAND2_X1 u4_sll_452_U201 ( .A1(u4_sll_452_ML_int_5__21_), .A2(u4_sll_452_n42), .ZN(u4_sll_452_n74) );
  INV_X1 u4_sll_452_U200 ( .A(u4_sll_452_n74), .ZN(u4_sll_452_ML_int_6__21_)
         );
  NAND2_X1 u4_sll_452_U199 ( .A1(u4_sll_452_ML_int_5__22_), .A2(u4_sll_452_n42), .ZN(u4_sll_452_n73) );
  INV_X1 u4_sll_452_U198 ( .A(u4_sll_452_n73), .ZN(u4_sll_452_ML_int_6__22_)
         );
  NAND2_X1 u4_sll_452_U197 ( .A1(u4_sll_452_ML_int_5__23_), .A2(u4_sll_452_n42), .ZN(u4_sll_452_n72) );
  INV_X1 u4_sll_452_U196 ( .A(u4_sll_452_n72), .ZN(u4_sll_452_ML_int_6__23_)
         );
  NAND2_X1 u4_sll_452_U195 ( .A1(u4_sll_452_ML_int_5__24_), .A2(u4_sll_452_n42), .ZN(u4_sll_452_n71) );
  INV_X1 u4_sll_452_U194 ( .A(u4_sll_452_n71), .ZN(u4_sll_452_ML_int_6__24_)
         );
  NAND2_X1 u4_sll_452_U193 ( .A1(u4_sll_452_ML_int_5__25_), .A2(u4_sll_452_n42), .ZN(u4_sll_452_n70) );
  INV_X1 u4_sll_452_U192 ( .A(u4_sll_452_n70), .ZN(u4_sll_452_ML_int_6__25_)
         );
  NAND2_X1 u4_sll_452_U191 ( .A1(u4_sll_452_ML_int_5__26_), .A2(u4_sll_452_n43), .ZN(u4_sll_452_n69) );
  INV_X1 u4_sll_452_U190 ( .A(u4_sll_452_n69), .ZN(u4_sll_452_ML_int_6__26_)
         );
  NAND2_X1 u4_sll_452_U189 ( .A1(u4_sll_452_ML_int_5__27_), .A2(u4_sll_452_n43), .ZN(u4_sll_452_n68) );
  INV_X1 u4_sll_452_U188 ( .A(u4_sll_452_n68), .ZN(u4_sll_452_ML_int_6__27_)
         );
  NAND2_X1 u4_sll_452_U187 ( .A1(u4_sll_452_ML_int_5__28_), .A2(u4_sll_452_n43), .ZN(u4_sll_452_n67) );
  INV_X1 u4_sll_452_U186 ( .A(u4_sll_452_n67), .ZN(u4_sll_452_ML_int_6__28_)
         );
  NAND2_X1 u4_sll_452_U185 ( .A1(u4_sll_452_ML_int_5__29_), .A2(u4_sll_452_n43), .ZN(u4_sll_452_n66) );
  INV_X1 u4_sll_452_U184 ( .A(u4_sll_452_n66), .ZN(u4_sll_452_ML_int_6__29_)
         );
  NAND2_X1 u4_sll_452_U183 ( .A1(u4_sll_452_ML_int_5__2_), .A2(u4_sll_452_n43), 
        .ZN(u4_sll_452_n65) );
  INV_X1 u4_sll_452_U182 ( .A(u4_sll_452_n65), .ZN(u4_sll_452_ML_int_6__2_) );
  NAND2_X1 u4_sll_452_U181 ( .A1(u4_sll_452_ML_int_5__30_), .A2(u4_sll_452_n43), .ZN(u4_sll_452_n64) );
  INV_X1 u4_sll_452_U180 ( .A(u4_sll_452_n64), .ZN(u4_sll_452_ML_int_6__30_)
         );
  NAND2_X1 u4_sll_452_U179 ( .A1(u4_sll_452_ML_int_5__31_), .A2(u4_sll_452_n43), .ZN(u4_sll_452_n63) );
  INV_X1 u4_sll_452_U178 ( .A(u4_sll_452_n63), .ZN(u4_sll_452_ML_int_6__31_)
         );
  NAND2_X1 u4_sll_452_U177 ( .A1(u4_sll_452_ML_int_5__3_), .A2(u4_sll_452_n43), 
        .ZN(u4_sll_452_n62) );
  INV_X1 u4_sll_452_U176 ( .A(u4_sll_452_n62), .ZN(u4_sll_452_ML_int_6__3_) );
  NAND2_X1 u4_sll_452_U175 ( .A1(u4_sll_452_ML_int_5__4_), .A2(u4_sll_452_n43), 
        .ZN(u4_sll_452_n61) );
  INV_X1 u4_sll_452_U174 ( .A(u4_sll_452_n61), .ZN(u4_sll_452_ML_int_6__4_) );
  NAND2_X1 u4_sll_452_U173 ( .A1(u4_sll_452_ML_int_5__5_), .A2(u4_sll_452_n43), 
        .ZN(u4_sll_452_n60) );
  INV_X1 u4_sll_452_U172 ( .A(u4_sll_452_n60), .ZN(u4_sll_452_ML_int_6__5_) );
  NAND2_X1 u4_sll_452_U171 ( .A1(u4_sll_452_ML_int_5__6_), .A2(u4_sll_452_n43), 
        .ZN(u4_sll_452_n58) );
  INV_X1 u4_sll_452_U170 ( .A(u4_sll_452_n58), .ZN(u4_sll_452_ML_int_6__6_) );
  NAND2_X1 u4_sll_452_U169 ( .A1(u4_sll_452_ML_int_5__7_), .A2(u4_sll_452_n43), 
        .ZN(u4_sll_452_n57) );
  INV_X1 u4_sll_452_U168 ( .A(u4_sll_452_n57), .ZN(u4_sll_452_ML_int_6__7_) );
  NAND2_X1 u4_sll_452_U167 ( .A1(u4_sll_452_ML_int_5__8_), .A2(u4_sll_452_n43), 
        .ZN(u4_sll_452_n56) );
  INV_X1 u4_sll_452_U166 ( .A(u4_sll_452_n56), .ZN(u4_sll_452_ML_int_6__8_) );
  NAND2_X1 u4_sll_452_U165 ( .A1(u4_sll_452_ML_int_5__9_), .A2(u4_sll_452_n43), 
        .ZN(u4_sll_452_n54) );
  INV_X1 u4_sll_452_U164 ( .A(u4_sll_452_n54), .ZN(u4_sll_452_ML_int_6__9_) );
  AOI21_X1 u4_sll_452_U163 ( .B1(u4_shift_left[6]), .B2(u4_sll_452_n88), .A(
        u4_sll_452_n89), .ZN(u4_sll_452_SHMAG_6_) );
  NOR2_X1 u4_sll_452_U162 ( .A1(u4_sll_452_n39), .A2(u4_shift_left[8]), .ZN(
        u4_sll_452_n59) );
  NOR2_X1 u4_sll_452_U161 ( .A1(u4_sll_452_n2), .A2(u4_sll_452_n87), .ZN(
        u4_N6008) );
  AND2_X1 u4_sll_452_U160 ( .A1(u4_sll_452_ML_int_7__100_), .A2(u4_sll_452_n1), 
        .ZN(u4_N6108) );
  AND2_X1 u4_sll_452_U159 ( .A1(u4_sll_452_ML_int_7__101_), .A2(u4_sll_452_n1), 
        .ZN(u4_N6109) );
  AND2_X1 u4_sll_452_U158 ( .A1(u4_sll_452_ML_int_7__102_), .A2(u4_sll_452_n1), 
        .ZN(u4_N6110) );
  AND2_X1 u4_sll_452_U157 ( .A1(u4_sll_452_ML_int_7__103_), .A2(u4_sll_452_n1), 
        .ZN(u4_N6111) );
  AND2_X1 u4_sll_452_U156 ( .A1(u4_sll_452_ML_int_7__104_), .A2(u4_sll_452_n1), 
        .ZN(u4_N6112) );
  AND2_X1 u4_sll_452_U155 ( .A1(u4_sll_452_ML_int_7__105_), .A2(u4_sll_452_n1), 
        .ZN(u4_N6113) );
  NOR2_X1 u4_sll_452_U154 ( .A1(u4_sll_452_n2), .A2(u4_sll_452_n86), .ZN(
        u4_N6018) );
  NOR2_X1 u4_sll_452_U153 ( .A1(u4_sll_452_n2), .A2(u4_sll_452_n85), .ZN(
        u4_N6019) );
  NOR2_X1 u4_sll_452_U152 ( .A1(u4_sll_452_n2), .A2(u4_sll_452_n84), .ZN(
        u4_N6020) );
  NOR2_X1 u4_sll_452_U151 ( .A1(u4_sll_452_n2), .A2(u4_sll_452_n83), .ZN(
        u4_N6021) );
  NOR2_X1 u4_sll_452_U150 ( .A1(u4_sll_452_n2), .A2(u4_sll_452_n82), .ZN(
        u4_N6022) );
  NOR2_X1 u4_sll_452_U149 ( .A1(u4_sll_452_n2), .A2(u4_sll_452_n81), .ZN(
        u4_N6023) );
  NOR2_X1 u4_sll_452_U148 ( .A1(u4_sll_452_n2), .A2(u4_sll_452_n80), .ZN(
        u4_N6024) );
  NOR2_X1 u4_sll_452_U147 ( .A1(u4_sll_452_n2), .A2(u4_sll_452_n79), .ZN(
        u4_N6025) );
  NOR2_X1 u4_sll_452_U146 ( .A1(u4_sll_452_n2), .A2(u4_sll_452_n78), .ZN(
        u4_N6026) );
  NOR2_X1 u4_sll_452_U145 ( .A1(u4_sll_452_n2), .A2(u4_sll_452_n77), .ZN(
        u4_N6027) );
  NOR2_X1 u4_sll_452_U144 ( .A1(u4_sll_452_n3), .A2(u4_sll_452_n76), .ZN(
        u4_N6009) );
  NOR2_X1 u4_sll_452_U143 ( .A1(u4_sll_452_n3), .A2(u4_sll_452_n75), .ZN(
        u4_N6028) );
  NOR2_X1 u4_sll_452_U142 ( .A1(u4_sll_452_n3), .A2(u4_sll_452_n74), .ZN(
        u4_N6029) );
  NOR2_X1 u4_sll_452_U141 ( .A1(u4_sll_452_n3), .A2(u4_sll_452_n73), .ZN(
        u4_N6030) );
  NOR2_X1 u4_sll_452_U140 ( .A1(u4_sll_452_n3), .A2(u4_sll_452_n72), .ZN(
        u4_N6031) );
  NOR2_X1 u4_sll_452_U139 ( .A1(u4_sll_452_n3), .A2(u4_sll_452_n71), .ZN(
        u4_N6032) );
  NOR2_X1 u4_sll_452_U138 ( .A1(u4_sll_452_n3), .A2(u4_sll_452_n70), .ZN(
        u4_N6033) );
  NOR2_X1 u4_sll_452_U137 ( .A1(u4_sll_452_n3), .A2(u4_sll_452_n69), .ZN(
        u4_N6034) );
  NOR2_X1 u4_sll_452_U136 ( .A1(u4_sll_452_n3), .A2(u4_sll_452_n68), .ZN(
        u4_N6035) );
  NOR2_X1 u4_sll_452_U135 ( .A1(u4_sll_452_n3), .A2(u4_sll_452_n67), .ZN(
        u4_N6036) );
  NOR2_X1 u4_sll_452_U134 ( .A1(u4_sll_452_n3), .A2(u4_sll_452_n66), .ZN(
        u4_N6037) );
  NOR2_X1 u4_sll_452_U133 ( .A1(u4_sll_452_n2), .A2(u4_sll_452_n65), .ZN(
        u4_N6010) );
  NOR2_X1 u4_sll_452_U132 ( .A1(u4_sll_452_n2), .A2(u4_sll_452_n64), .ZN(
        u4_N6038) );
  NOR2_X1 u4_sll_452_U131 ( .A1(u4_sll_452_n3), .A2(u4_sll_452_n63), .ZN(
        u4_N6039) );
  AND2_X1 u4_sll_452_U130 ( .A1(u4_sll_452_ML_int_6__32_), .A2(u4_sll_452_n59), 
        .ZN(u4_N6040) );
  AND2_X1 u4_sll_452_U129 ( .A1(u4_sll_452_ML_int_6__33_), .A2(u4_sll_452_n59), 
        .ZN(u4_N6041) );
  AND2_X1 u4_sll_452_U128 ( .A1(u4_sll_452_ML_int_6__34_), .A2(u4_sll_452_n59), 
        .ZN(u4_N6042) );
  AND2_X1 u4_sll_452_U127 ( .A1(u4_sll_452_ML_int_6__35_), .A2(u4_sll_452_n4), 
        .ZN(u4_N6043) );
  AND2_X1 u4_sll_452_U126 ( .A1(u4_sll_452_ML_int_6__36_), .A2(u4_sll_452_n4), 
        .ZN(u4_N6044) );
  AND2_X1 u4_sll_452_U125 ( .A1(u4_sll_452_ML_int_6__37_), .A2(u4_sll_452_n59), 
        .ZN(u4_N6045) );
  AND2_X1 u4_sll_452_U124 ( .A1(u4_sll_452_ML_int_6__38_), .A2(u4_sll_452_n59), 
        .ZN(u4_N6046) );
  AND2_X1 u4_sll_452_U123 ( .A1(u4_sll_452_ML_int_6__39_), .A2(u4_sll_452_n4), 
        .ZN(u4_N6047) );
  NOR2_X1 u4_sll_452_U122 ( .A1(u4_sll_452_n2), .A2(u4_sll_452_n62), .ZN(
        u4_N6011) );
  AND2_X1 u4_sll_452_U121 ( .A1(u4_sll_452_ML_int_6__40_), .A2(u4_sll_452_n59), 
        .ZN(u4_N6048) );
  AND2_X1 u4_sll_452_U120 ( .A1(u4_sll_452_ML_int_6__41_), .A2(u4_sll_452_n59), 
        .ZN(u4_N6049) );
  AND2_X1 u4_sll_452_U119 ( .A1(u4_sll_452_ML_int_6__42_), .A2(u4_sll_452_n59), 
        .ZN(u4_N6050) );
  AND2_X1 u4_sll_452_U118 ( .A1(u4_sll_452_ML_int_6__43_), .A2(u4_sll_452_n59), 
        .ZN(u4_N6051) );
  AND2_X1 u4_sll_452_U117 ( .A1(u4_sll_452_ML_int_6__44_), .A2(u4_sll_452_n59), 
        .ZN(u4_N6052) );
  AND2_X1 u4_sll_452_U116 ( .A1(u4_sll_452_ML_int_6__45_), .A2(u4_sll_452_n59), 
        .ZN(u4_N6053) );
  AND2_X1 u4_sll_452_U115 ( .A1(u4_sll_452_ML_int_6__46_), .A2(u4_sll_452_n59), 
        .ZN(u4_N6054) );
  AND2_X1 u4_sll_452_U114 ( .A1(u4_sll_452_ML_int_6__47_), .A2(u4_sll_452_n59), 
        .ZN(u4_N6055) );
  AND2_X1 u4_sll_452_U113 ( .A1(u4_sll_452_ML_int_6__48_), .A2(u4_sll_452_n59), 
        .ZN(u4_N6056) );
  AND2_X1 u4_sll_452_U112 ( .A1(u4_sll_452_ML_int_6__49_), .A2(u4_sll_452_n59), 
        .ZN(u4_N6057) );
  NOR2_X1 u4_sll_452_U111 ( .A1(u4_sll_452_n2), .A2(u4_sll_452_n61), .ZN(
        u4_N6012) );
  AND2_X1 u4_sll_452_U110 ( .A1(u4_sll_452_ML_int_6__50_), .A2(u4_sll_452_n59), 
        .ZN(u4_N6058) );
  AND2_X1 u4_sll_452_U109 ( .A1(u4_sll_452_ML_int_6__51_), .A2(u4_sll_452_n59), 
        .ZN(u4_N6059) );
  AND2_X1 u4_sll_452_U108 ( .A1(u4_sll_452_ML_int_6__52_), .A2(u4_sll_452_n59), 
        .ZN(u4_N6060) );
  AND2_X1 u4_sll_452_U107 ( .A1(u4_sll_452_ML_int_6__53_), .A2(u4_sll_452_n4), 
        .ZN(u4_N6061) );
  AND2_X1 u4_sll_452_U106 ( .A1(u4_sll_452_ML_int_6__54_), .A2(u4_sll_452_n59), 
        .ZN(u4_N6062) );
  AND2_X1 u4_sll_452_U105 ( .A1(u4_sll_452_ML_int_6__55_), .A2(u4_sll_452_n4), 
        .ZN(u4_N6063) );
  AND2_X1 u4_sll_452_U104 ( .A1(u4_sll_452_ML_int_6__56_), .A2(u4_sll_452_n4), 
        .ZN(u4_N6064) );
  AND2_X1 u4_sll_452_U103 ( .A1(u4_sll_452_ML_int_6__57_), .A2(u4_sll_452_n4), 
        .ZN(u4_N6065) );
  AND2_X1 u4_sll_452_U102 ( .A1(u4_sll_452_ML_int_6__58_), .A2(u4_sll_452_n4), 
        .ZN(u4_N6066) );
  AND2_X1 u4_sll_452_U101 ( .A1(u4_sll_452_ML_int_6__59_), .A2(u4_sll_452_n4), 
        .ZN(u4_N6067) );
  NOR2_X1 u4_sll_452_U100 ( .A1(u4_sll_452_n2), .A2(u4_sll_452_n60), .ZN(
        u4_N6013) );
  AND2_X1 u4_sll_452_U99 ( .A1(u4_sll_452_ML_int_6__60_), .A2(u4_sll_452_n4), 
        .ZN(u4_N6068) );
  AND2_X1 u4_sll_452_U98 ( .A1(u4_sll_452_ML_int_6__61_), .A2(u4_sll_452_n4), 
        .ZN(u4_N6069) );
  AND2_X1 u4_sll_452_U97 ( .A1(u4_sll_452_ML_int_6__62_), .A2(u4_sll_452_n4), 
        .ZN(u4_N6070) );
  AND2_X1 u4_sll_452_U96 ( .A1(u4_sll_452_ML_int_6__63_), .A2(u4_sll_452_n4), 
        .ZN(u4_N6071) );
  AND2_X1 u4_sll_452_U95 ( .A1(u4_sll_452_ML_int_7__64_), .A2(u4_sll_452_n1), 
        .ZN(u4_N6072) );
  AND2_X1 u4_sll_452_U94 ( .A1(u4_sll_452_ML_int_7__65_), .A2(u4_sll_452_n1), 
        .ZN(u4_N6073) );
  AND2_X1 u4_sll_452_U93 ( .A1(u4_sll_452_ML_int_7__66_), .A2(u4_sll_452_n1), 
        .ZN(u4_N6074) );
  AND2_X1 u4_sll_452_U92 ( .A1(u4_sll_452_ML_int_7__67_), .A2(u4_sll_452_n1), 
        .ZN(u4_N6075) );
  AND2_X1 u4_sll_452_U91 ( .A1(u4_sll_452_ML_int_7__68_), .A2(u4_sll_452_n55), 
        .ZN(u4_N6076) );
  AND2_X1 u4_sll_452_U90 ( .A1(u4_sll_452_ML_int_7__69_), .A2(u4_sll_452_n55), 
        .ZN(u4_N6077) );
  NOR2_X1 u4_sll_452_U89 ( .A1(u4_sll_452_n2), .A2(u4_sll_452_n58), .ZN(
        u4_N6014) );
  AND2_X1 u4_sll_452_U88 ( .A1(u4_sll_452_ML_int_7__70_), .A2(u4_sll_452_n55), 
        .ZN(u4_N6078) );
  AND2_X1 u4_sll_452_U87 ( .A1(u4_sll_452_ML_int_7__71_), .A2(u4_sll_452_n55), 
        .ZN(u4_N6079) );
  AND2_X1 u4_sll_452_U86 ( .A1(u4_sll_452_ML_int_7__72_), .A2(u4_sll_452_n55), 
        .ZN(u4_N6080) );
  AND2_X1 u4_sll_452_U85 ( .A1(u4_sll_452_ML_int_7__73_), .A2(u4_sll_452_n55), 
        .ZN(u4_N6081) );
  AND2_X1 u4_sll_452_U84 ( .A1(u4_sll_452_ML_int_7__74_), .A2(u4_sll_452_n55), 
        .ZN(u4_N6082) );
  AND2_X1 u4_sll_452_U83 ( .A1(u4_sll_452_ML_int_7__75_), .A2(u4_sll_452_n55), 
        .ZN(u4_N6083) );
  AND2_X1 u4_sll_452_U82 ( .A1(u4_sll_452_ML_int_7__76_), .A2(u4_sll_452_n55), 
        .ZN(u4_N6084) );
  AND2_X1 u4_sll_452_U81 ( .A1(u4_sll_452_ML_int_7__77_), .A2(u4_sll_452_n55), 
        .ZN(u4_N6085) );
  AND2_X1 u4_sll_452_U80 ( .A1(u4_sll_452_ML_int_7__78_), .A2(u4_sll_452_n55), 
        .ZN(u4_N6086) );
  AND2_X1 u4_sll_452_U79 ( .A1(u4_sll_452_ML_int_7__79_), .A2(u4_sll_452_n55), 
        .ZN(u4_N6087) );
  NOR2_X1 u4_sll_452_U78 ( .A1(u4_sll_452_n3), .A2(u4_sll_452_n57), .ZN(
        u4_N6015) );
  AND2_X1 u4_sll_452_U77 ( .A1(u4_sll_452_ML_int_7__80_), .A2(u4_sll_452_n55), 
        .ZN(u4_N6088) );
  AND2_X1 u4_sll_452_U76 ( .A1(u4_sll_452_ML_int_7__81_), .A2(u4_sll_452_n55), 
        .ZN(u4_N6089) );
  AND2_X1 u4_sll_452_U75 ( .A1(u4_sll_452_ML_int_7__82_), .A2(u4_sll_452_n55), 
        .ZN(u4_N6090) );
  AND2_X1 u4_sll_452_U74 ( .A1(u4_sll_452_ML_int_7__83_), .A2(u4_sll_452_n55), 
        .ZN(u4_N6091) );
  AND2_X1 u4_sll_452_U73 ( .A1(u4_sll_452_ML_int_7__84_), .A2(u4_sll_452_n55), 
        .ZN(u4_N6092) );
  AND2_X1 u4_sll_452_U72 ( .A1(u4_sll_452_ML_int_7__85_), .A2(u4_sll_452_n55), 
        .ZN(u4_N6093) );
  AND2_X1 u4_sll_452_U71 ( .A1(u4_sll_452_ML_int_7__86_), .A2(u4_sll_452_n55), 
        .ZN(u4_N6094) );
  AND2_X1 u4_sll_452_U70 ( .A1(u4_sll_452_ML_int_7__87_), .A2(u4_sll_452_n1), 
        .ZN(u4_N6095) );
  AND2_X1 u4_sll_452_U69 ( .A1(u4_sll_452_ML_int_7__88_), .A2(u4_sll_452_n1), 
        .ZN(u4_N6096) );
  AND2_X1 u4_sll_452_U68 ( .A1(u4_sll_452_ML_int_7__89_), .A2(u4_sll_452_n1), 
        .ZN(u4_N6097) );
  NOR2_X1 u4_sll_452_U67 ( .A1(u4_sll_452_n2), .A2(u4_sll_452_n56), .ZN(
        u4_N6016) );
  AND2_X1 u4_sll_452_U66 ( .A1(u4_sll_452_ML_int_7__90_), .A2(u4_sll_452_n1), 
        .ZN(u4_N6098) );
  AND2_X1 u4_sll_452_U65 ( .A1(u4_sll_452_ML_int_7__91_), .A2(u4_sll_452_n1), 
        .ZN(u4_N6099) );
  AND2_X1 u4_sll_452_U64 ( .A1(u4_sll_452_ML_int_7__92_), .A2(u4_sll_452_n1), 
        .ZN(u4_N6100) );
  AND2_X1 u4_sll_452_U63 ( .A1(u4_sll_452_ML_int_7__93_), .A2(u4_sll_452_n1), 
        .ZN(u4_N6101) );
  AND2_X1 u4_sll_452_U62 ( .A1(u4_sll_452_ML_int_7__94_), .A2(u4_sll_452_n1), 
        .ZN(u4_N6102) );
  AND2_X1 u4_sll_452_U61 ( .A1(u4_sll_452_ML_int_7__95_), .A2(u4_sll_452_n1), 
        .ZN(u4_N6103) );
  AND2_X1 u4_sll_452_U60 ( .A1(u4_sll_452_ML_int_7__96_), .A2(u4_sll_452_n1), 
        .ZN(u4_N6104) );
  AND2_X1 u4_sll_452_U59 ( .A1(u4_sll_452_ML_int_7__97_), .A2(u4_sll_452_n1), 
        .ZN(u4_N6105) );
  AND2_X1 u4_sll_452_U58 ( .A1(u4_sll_452_ML_int_7__98_), .A2(u4_sll_452_n1), 
        .ZN(u4_N6106) );
  AND2_X1 u4_sll_452_U57 ( .A1(u4_sll_452_ML_int_7__99_), .A2(u4_sll_452_n1), 
        .ZN(u4_N6107) );
  NOR2_X1 u4_sll_452_U56 ( .A1(u4_sll_452_n2), .A2(u4_sll_452_n54), .ZN(
        u4_N6017) );
  INV_X4 u4_sll_452_U55 ( .A(u4_sll_452_n4), .ZN(u4_sll_452_n3) );
  INV_X4 u4_sll_452_U54 ( .A(u4_sll_452_n4), .ZN(u4_sll_452_n2) );
  INV_X4 u4_sll_452_U53 ( .A(u4_sll_452_n41), .ZN(u4_sll_452_n45) );
  INV_X4 u4_sll_452_U52 ( .A(u4_sll_452_n52), .ZN(u4_sll_452_n50) );
  INV_X4 u4_sll_452_U51 ( .A(u4_sll_452_n37), .ZN(u4_sll_452_n30) );
  INV_X4 u4_sll_452_U50 ( .A(u4_sll_452_n26), .ZN(u4_sll_452_n24) );
  INV_X4 u4_sll_452_U49 ( .A(u4_sll_452_SHMAG_2_), .ZN(u4_sll_452_n15) );
  INV_X4 u4_sll_452_U48 ( .A(u4_sll_452_n5), .ZN(u4_sll_452_n4) );
  INV_X4 u4_sll_452_U47 ( .A(u4_sll_452_n59), .ZN(u4_sll_452_n5) );
  INV_X4 u4_sll_452_U46 ( .A(u4_sll_452_n41), .ZN(u4_sll_452_n44) );
  INV_X4 u4_sll_452_U45 ( .A(u4_sll_452_n30), .ZN(u4_sll_452_n27) );
  INV_X4 u4_sll_452_U44 ( .A(u4_sll_452_SHMAG_0_), .ZN(u4_sll_452_n7) );
  INV_X4 u4_sll_452_U43 ( .A(u4_sll_452_SHMAG_6_), .ZN(u4_sll_452_n40) );
  INV_X4 u4_sll_452_U42 ( .A(u4_sll_452_SHMAG_6_), .ZN(u4_sll_452_n39) );
  INV_X4 u4_sll_452_U41 ( .A(u4_sll_452_SHMAG_0_), .ZN(u4_sll_452_n6) );
  INV_X4 u4_sll_452_U40 ( .A(u4_sll_452_SHMAG_1_), .ZN(u4_sll_452_n10) );
  INV_X4 u4_sll_452_U39 ( .A(u4_sll_452_SHMAG_2_), .ZN(u4_sll_452_n14) );
  INV_X4 u4_sll_452_U38 ( .A(u4_shift_left[8]), .ZN(u4_sll_452_n1) );
  INV_X4 u4_sll_452_U37 ( .A(u4_sll_452_n38), .ZN(u4_sll_452_n37) );
  INV_X4 u4_sll_452_U36 ( .A(u4_sll_452_n45), .ZN(u4_sll_452_n42) );
  INV_X4 u4_sll_452_U35 ( .A(u4_sll_452_n51), .ZN(u4_sll_452_n46) );
  INV_X4 u4_sll_452_U34 ( .A(u4_sll_452_n19), .ZN(u4_sll_452_n18) );
  INV_X4 u4_sll_452_U33 ( .A(u4_sll_452_SHMAG_0_), .ZN(u4_sll_452_n9) );
  INV_X4 u4_sll_452_U32 ( .A(u4_sll_452_SHMAG_0_), .ZN(u4_sll_452_n8) );
  INV_X4 u4_sll_452_U31 ( .A(u4_sll_452_SHMAG_2_), .ZN(u4_sll_452_n16) );
  INV_X4 u4_sll_452_U30 ( .A(u4_sll_452_SHMAG_2_), .ZN(u4_sll_452_n17) );
  INV_X4 u4_sll_452_U29 ( .A(u4_sll_452_n52), .ZN(u4_sll_452_n51) );
  INV_X4 u4_sll_452_U28 ( .A(u4_sll_452_n38), .ZN(u4_sll_452_n36) );
  INV_X4 u4_sll_452_U27 ( .A(u4_sll_452_n26), .ZN(u4_sll_452_n25) );
  INV_X4 u4_sll_452_U26 ( .A(u4_sll_452_n29), .ZN(u4_sll_452_n28) );
  INV_X4 u4_sll_452_U25 ( .A(u4_sll_452_n37), .ZN(u4_sll_452_n29) );
  INV_X4 u4_sll_452_U24 ( .A(u4_sll_452_SHMAG_1_), .ZN(u4_sll_452_n11) );
  INV_X4 u4_sll_452_U23 ( .A(u4_sll_452_n25), .ZN(u4_sll_452_n19) );
  INV_X4 u4_sll_452_U22 ( .A(u4_sll_452_n24), .ZN(u4_sll_452_n20) );
  INV_X4 u4_sll_452_U21 ( .A(u4_sll_452_n46), .ZN(u4_sll_452_n41) );
  INV_X4 u4_sll_452_U20 ( .A(u4_sll_452_n53), .ZN(u4_sll_452_n52) );
  INV_X4 u4_sll_452_U19 ( .A(u4_sll_452_n38), .ZN(u4_sll_452_n35) );
  INV_X4 u4_sll_452_U18 ( .A(u4_sll_452_SHMAG_1_), .ZN(u4_sll_452_n13) );
  INV_X4 u4_sll_452_U17 ( .A(u4_sll_452_SHMAG_1_), .ZN(u4_sll_452_n12) );
  INV_X4 u4_sll_452_U16 ( .A(u4_sll_452_n44), .ZN(u4_sll_452_n43) );
  INV_X4 u4_sll_452_U15 ( .A(u4_sll_452_n23), .ZN(u4_sll_452_n21) );
  INV_X4 u4_sll_452_U14 ( .A(u4_sll_452_n23), .ZN(u4_sll_452_n22) );
  INV_X4 u4_sll_452_U13 ( .A(u4_sll_452_n26), .ZN(u4_sll_452_n23) );
  INV_X4 u4_sll_452_U12 ( .A(u4_sll_452_n50), .ZN(u4_sll_452_n49) );
  INV_X4 u4_sll_452_U11 ( .A(u4_sll_452_n36), .ZN(u4_sll_452_n31) );
  INV_X4 u4_sll_452_U10 ( .A(u4_sll_452_n50), .ZN(u4_sll_452_n48) );
  INV_X4 u4_sll_452_U9 ( .A(u4_sll_452_n51), .ZN(u4_sll_452_n47) );
  INV_X4 u4_sll_452_U8 ( .A(u4_sll_452_n36), .ZN(u4_sll_452_n32) );
  INV_X4 u4_sll_452_U7 ( .A(u4_sll_452_n35), .ZN(u4_sll_452_n33) );
  INV_X4 u4_sll_452_U6 ( .A(u4_sll_452_n35), .ZN(u4_sll_452_n34) );
  INV_X4 u4_sll_452_U5 ( .A(u4_sll_452_SHMAG_3_), .ZN(u4_sll_452_n26) );
  INV_X4 u4_sll_452_U4 ( .A(u4_sll_452_temp_int_SH_5_), .ZN(u4_sll_452_n53) );
  INV_X4 u4_sll_452_U3 ( .A(u4_sll_452_SHMAG_4_), .ZN(u4_sll_452_n38) );
  MUX2_X2 u4_sll_452_M1_0_1 ( .A(fract_denorm[1]), .B(fract_denorm[0]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__1_) );
  MUX2_X2 u4_sll_452_M1_0_2 ( .A(fract_denorm[2]), .B(fract_denorm[1]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__2_) );
  MUX2_X2 u4_sll_452_M1_0_3 ( .A(fract_denorm[3]), .B(fract_denorm[2]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__3_) );
  MUX2_X2 u4_sll_452_M1_0_4 ( .A(fract_denorm[4]), .B(fract_denorm[3]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__4_) );
  MUX2_X2 u4_sll_452_M1_0_5 ( .A(fract_denorm[5]), .B(fract_denorm[4]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__5_) );
  MUX2_X2 u4_sll_452_M1_0_6 ( .A(fract_denorm[6]), .B(fract_denorm[5]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__6_) );
  MUX2_X2 u4_sll_452_M1_0_7 ( .A(fract_denorm[7]), .B(fract_denorm[6]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__7_) );
  MUX2_X2 u4_sll_452_M1_0_8 ( .A(fract_denorm[8]), .B(fract_denorm[7]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__8_) );
  MUX2_X2 u4_sll_452_M1_0_9 ( .A(fract_denorm[9]), .B(fract_denorm[8]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__9_) );
  MUX2_X2 u4_sll_452_M1_0_10 ( .A(fract_denorm[10]), .B(fract_denorm[9]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__10_) );
  MUX2_X2 u4_sll_452_M1_0_11 ( .A(fract_denorm[11]), .B(fract_denorm[10]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__11_) );
  MUX2_X2 u4_sll_452_M1_0_12 ( .A(fract_denorm[12]), .B(fract_denorm[11]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__12_) );
  MUX2_X2 u4_sll_452_M1_0_13 ( .A(fract_denorm[13]), .B(fract_denorm[12]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__13_) );
  MUX2_X2 u4_sll_452_M1_0_14 ( .A(fract_denorm[14]), .B(fract_denorm[13]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__14_) );
  MUX2_X2 u4_sll_452_M1_0_15 ( .A(fract_denorm[15]), .B(fract_denorm[14]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__15_) );
  MUX2_X2 u4_sll_452_M1_0_16 ( .A(fract_denorm[16]), .B(fract_denorm[15]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__16_) );
  MUX2_X2 u4_sll_452_M1_0_17 ( .A(fract_denorm[17]), .B(fract_denorm[16]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__17_) );
  MUX2_X2 u4_sll_452_M1_0_18 ( .A(fract_denorm[18]), .B(fract_denorm[17]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__18_) );
  MUX2_X2 u4_sll_452_M1_0_19 ( .A(fract_denorm[19]), .B(fract_denorm[18]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__19_) );
  MUX2_X2 u4_sll_452_M1_0_20 ( .A(fract_denorm[20]), .B(fract_denorm[19]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__20_) );
  MUX2_X2 u4_sll_452_M1_0_21 ( .A(fract_denorm[21]), .B(fract_denorm[20]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__21_) );
  MUX2_X2 u4_sll_452_M1_0_22 ( .A(fract_denorm[22]), .B(fract_denorm[21]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__22_) );
  MUX2_X2 u4_sll_452_M1_0_23 ( .A(fract_denorm[23]), .B(fract_denorm[22]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__23_) );
  MUX2_X2 u4_sll_452_M1_0_24 ( .A(fract_denorm[24]), .B(fract_denorm[23]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__24_) );
  MUX2_X2 u4_sll_452_M1_0_25 ( .A(fract_denorm[25]), .B(fract_denorm[24]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__25_) );
  MUX2_X2 u4_sll_452_M1_0_26 ( .A(fract_denorm[26]), .B(fract_denorm[25]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__26_) );
  MUX2_X2 u4_sll_452_M1_0_27 ( .A(fract_denorm[27]), .B(fract_denorm[26]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__27_) );
  MUX2_X2 u4_sll_452_M1_0_28 ( .A(fract_denorm[28]), .B(fract_denorm[27]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__28_) );
  MUX2_X2 u4_sll_452_M1_0_29 ( .A(fract_denorm[29]), .B(fract_denorm[28]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__29_) );
  MUX2_X2 u4_sll_452_M1_0_30 ( .A(fract_denorm[30]), .B(fract_denorm[29]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__30_) );
  MUX2_X2 u4_sll_452_M1_0_31 ( .A(fract_denorm[31]), .B(fract_denorm[30]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__31_) );
  MUX2_X2 u4_sll_452_M1_0_32 ( .A(fract_denorm[32]), .B(fract_denorm[31]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__32_) );
  MUX2_X2 u4_sll_452_M1_0_33 ( .A(fract_denorm[33]), .B(fract_denorm[32]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__33_) );
  MUX2_X2 u4_sll_452_M1_0_34 ( .A(fract_denorm[34]), .B(fract_denorm[33]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__34_) );
  MUX2_X2 u4_sll_452_M1_0_35 ( .A(fract_denorm[35]), .B(fract_denorm[34]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__35_) );
  MUX2_X2 u4_sll_452_M1_0_36 ( .A(fract_denorm[36]), .B(fract_denorm[35]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__36_) );
  MUX2_X2 u4_sll_452_M1_0_37 ( .A(fract_denorm[37]), .B(fract_denorm[36]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__37_) );
  MUX2_X2 u4_sll_452_M1_0_38 ( .A(fract_denorm[38]), .B(fract_denorm[37]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__38_) );
  MUX2_X2 u4_sll_452_M1_0_39 ( .A(fract_denorm[39]), .B(fract_denorm[38]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__39_) );
  MUX2_X2 u4_sll_452_M1_0_40 ( .A(fract_denorm[40]), .B(fract_denorm[39]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__40_) );
  MUX2_X2 u4_sll_452_M1_0_41 ( .A(fract_denorm[41]), .B(fract_denorm[40]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__41_) );
  MUX2_X2 u4_sll_452_M1_0_42 ( .A(fract_denorm[42]), .B(fract_denorm[41]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__42_) );
  MUX2_X2 u4_sll_452_M1_0_43 ( .A(fract_denorm[43]), .B(fract_denorm[42]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__43_) );
  MUX2_X2 u4_sll_452_M1_0_44 ( .A(fract_denorm[44]), .B(fract_denorm[43]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__44_) );
  MUX2_X2 u4_sll_452_M1_0_45 ( .A(fract_denorm[45]), .B(fract_denorm[44]), .S(
        u4_sll_452_n6), .Z(u4_sll_452_ML_int_1__45_) );
  MUX2_X2 u4_sll_452_M1_0_46 ( .A(fract_denorm[46]), .B(fract_denorm[45]), .S(
        u4_sll_452_n6), .Z(u4_sll_452_ML_int_1__46_) );
  MUX2_X2 u4_sll_452_M1_0_47 ( .A(fract_denorm[47]), .B(fract_denorm[46]), .S(
        u4_sll_452_n6), .Z(u4_sll_452_ML_int_1__47_) );
  MUX2_X2 u4_sll_452_M1_0_48 ( .A(fract_denorm[48]), .B(fract_denorm[47]), .S(
        u4_sll_452_n6), .Z(u4_sll_452_ML_int_1__48_) );
  MUX2_X2 u4_sll_452_M1_0_49 ( .A(fract_denorm[49]), .B(fract_denorm[48]), .S(
        u4_sll_452_n6), .Z(u4_sll_452_ML_int_1__49_) );
  MUX2_X2 u4_sll_452_M1_0_50 ( .A(fract_denorm[50]), .B(fract_denorm[49]), .S(
        u4_sll_452_n6), .Z(u4_sll_452_ML_int_1__50_) );
  MUX2_X2 u4_sll_452_M1_0_51 ( .A(fract_denorm[51]), .B(fract_denorm[50]), .S(
        u4_sll_452_n6), .Z(u4_sll_452_ML_int_1__51_) );
  MUX2_X2 u4_sll_452_M1_0_52 ( .A(fract_denorm[52]), .B(fract_denorm[51]), .S(
        u4_sll_452_n6), .Z(u4_sll_452_ML_int_1__52_) );
  MUX2_X2 u4_sll_452_M1_0_53 ( .A(fract_denorm[53]), .B(fract_denorm[52]), .S(
        u4_sll_452_n6), .Z(u4_sll_452_ML_int_1__53_) );
  MUX2_X2 u4_sll_452_M1_0_54 ( .A(fract_denorm[54]), .B(fract_denorm[53]), .S(
        u4_sll_452_n6), .Z(u4_sll_452_ML_int_1__54_) );
  MUX2_X2 u4_sll_452_M1_0_55 ( .A(fract_denorm[55]), .B(fract_denorm[54]), .S(
        u4_sll_452_n6), .Z(u4_sll_452_ML_int_1__55_) );
  MUX2_X2 u4_sll_452_M1_0_56 ( .A(fract_denorm[56]), .B(fract_denorm[55]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__56_) );
  MUX2_X2 u4_sll_452_M1_0_57 ( .A(fract_denorm[57]), .B(fract_denorm[56]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__57_) );
  MUX2_X2 u4_sll_452_M1_0_58 ( .A(fract_denorm[58]), .B(fract_denorm[57]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__58_) );
  MUX2_X2 u4_sll_452_M1_0_59 ( .A(fract_denorm[59]), .B(fract_denorm[58]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__59_) );
  MUX2_X2 u4_sll_452_M1_0_60 ( .A(fract_denorm[60]), .B(fract_denorm[59]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__60_) );
  MUX2_X2 u4_sll_452_M1_0_61 ( .A(fract_denorm[61]), .B(fract_denorm[60]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__61_) );
  MUX2_X2 u4_sll_452_M1_0_62 ( .A(fract_denorm[62]), .B(fract_denorm[61]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__62_) );
  MUX2_X2 u4_sll_452_M1_0_63 ( .A(fract_denorm[63]), .B(fract_denorm[62]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__63_) );
  MUX2_X2 u4_sll_452_M1_0_64 ( .A(fract_denorm[64]), .B(fract_denorm[63]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__64_) );
  MUX2_X2 u4_sll_452_M1_0_65 ( .A(fract_denorm[65]), .B(fract_denorm[64]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__65_) );
  MUX2_X2 u4_sll_452_M1_0_66 ( .A(fract_denorm[66]), .B(fract_denorm[65]), .S(
        u4_sll_452_n6), .Z(u4_sll_452_ML_int_1__66_) );
  MUX2_X2 u4_sll_452_M1_0_67 ( .A(fract_denorm[67]), .B(fract_denorm[66]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__67_) );
  MUX2_X2 u4_sll_452_M1_0_68 ( .A(fract_denorm[68]), .B(fract_denorm[67]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__68_) );
  MUX2_X2 u4_sll_452_M1_0_69 ( .A(fract_denorm[69]), .B(fract_denorm[68]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__69_) );
  MUX2_X2 u4_sll_452_M1_0_70 ( .A(fract_denorm[70]), .B(fract_denorm[69]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__70_) );
  MUX2_X2 u4_sll_452_M1_0_71 ( .A(fract_denorm[71]), .B(fract_denorm[70]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__71_) );
  MUX2_X2 u4_sll_452_M1_0_72 ( .A(fract_denorm[72]), .B(fract_denorm[71]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__72_) );
  MUX2_X2 u4_sll_452_M1_0_73 ( .A(fract_denorm[73]), .B(fract_denorm[72]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__73_) );
  MUX2_X2 u4_sll_452_M1_0_74 ( .A(fract_denorm[74]), .B(fract_denorm[73]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__74_) );
  MUX2_X2 u4_sll_452_M1_0_75 ( .A(fract_denorm[75]), .B(fract_denorm[74]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__75_) );
  MUX2_X2 u4_sll_452_M1_0_76 ( .A(fract_denorm[76]), .B(fract_denorm[75]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__76_) );
  MUX2_X2 u4_sll_452_M1_0_77 ( .A(fract_denorm[77]), .B(fract_denorm[76]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__77_) );
  MUX2_X2 u4_sll_452_M1_0_78 ( .A(fract_denorm[78]), .B(fract_denorm[77]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__78_) );
  MUX2_X2 u4_sll_452_M1_0_79 ( .A(fract_denorm[79]), .B(fract_denorm[78]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__79_) );
  MUX2_X2 u4_sll_452_M1_0_80 ( .A(fract_denorm[80]), .B(fract_denorm[79]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__80_) );
  MUX2_X2 u4_sll_452_M1_0_81 ( .A(fract_denorm[81]), .B(fract_denorm[80]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__81_) );
  MUX2_X2 u4_sll_452_M1_0_82 ( .A(fract_denorm[82]), .B(fract_denorm[81]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__82_) );
  MUX2_X2 u4_sll_452_M1_0_83 ( .A(fract_denorm[83]), .B(fract_denorm[82]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__83_) );
  MUX2_X2 u4_sll_452_M1_0_84 ( .A(fract_denorm[84]), .B(fract_denorm[83]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__84_) );
  MUX2_X2 u4_sll_452_M1_0_85 ( .A(fract_denorm[85]), .B(fract_denorm[84]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__85_) );
  MUX2_X2 u4_sll_452_M1_0_86 ( .A(fract_denorm[86]), .B(fract_denorm[85]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__86_) );
  MUX2_X2 u4_sll_452_M1_0_87 ( .A(fract_denorm[87]), .B(fract_denorm[86]), .S(
        u4_sll_452_n9), .Z(u4_sll_452_ML_int_1__87_) );
  MUX2_X2 u4_sll_452_M1_0_88 ( .A(fract_denorm[88]), .B(fract_denorm[87]), .S(
        u4_sll_452_n8), .Z(u4_sll_452_ML_int_1__88_) );
  MUX2_X2 u4_sll_452_M1_0_89 ( .A(fract_denorm[89]), .B(fract_denorm[88]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__89_) );
  MUX2_X2 u4_sll_452_M1_0_90 ( .A(fract_denorm[90]), .B(fract_denorm[89]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__90_) );
  MUX2_X2 u4_sll_452_M1_0_91 ( .A(fract_denorm[91]), .B(fract_denorm[90]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__91_) );
  MUX2_X2 u4_sll_452_M1_0_92 ( .A(fract_denorm[92]), .B(fract_denorm[91]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__92_) );
  MUX2_X2 u4_sll_452_M1_0_93 ( .A(fract_denorm[93]), .B(fract_denorm[92]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__93_) );
  MUX2_X2 u4_sll_452_M1_0_94 ( .A(fract_denorm[94]), .B(fract_denorm[93]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__94_) );
  MUX2_X2 u4_sll_452_M1_0_95 ( .A(fract_denorm[95]), .B(fract_denorm[94]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__95_) );
  MUX2_X2 u4_sll_452_M1_0_96 ( .A(fract_denorm[96]), .B(fract_denorm[95]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__96_) );
  MUX2_X2 u4_sll_452_M1_0_97 ( .A(fract_denorm[97]), .B(fract_denorm[96]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__97_) );
  MUX2_X2 u4_sll_452_M1_0_98 ( .A(fract_denorm[98]), .B(fract_denorm[97]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__98_) );
  MUX2_X2 u4_sll_452_M1_0_99 ( .A(fract_denorm[99]), .B(fract_denorm[98]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__99_) );
  MUX2_X2 u4_sll_452_M1_0_100 ( .A(fract_denorm[100]), .B(fract_denorm[99]), 
        .S(u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__100_) );
  MUX2_X2 u4_sll_452_M1_0_101 ( .A(fract_denorm[101]), .B(fract_denorm[100]), 
        .S(u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__101_) );
  MUX2_X2 u4_sll_452_M1_0_102 ( .A(fract_denorm[102]), .B(fract_denorm[101]), 
        .S(u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__102_) );
  MUX2_X2 u4_sll_452_M1_0_103 ( .A(fract_denorm[103]), .B(fract_denorm[102]), 
        .S(u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__103_) );
  MUX2_X2 u4_sll_452_M1_0_104 ( .A(fract_denorm[104]), .B(fract_denorm[103]), 
        .S(u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__104_) );
  MUX2_X2 u4_sll_452_M1_0_105 ( .A(n4873), .B(fract_denorm[104]), .S(
        u4_sll_452_n7), .Z(u4_sll_452_ML_int_1__105_) );
  MUX2_X2 u4_sll_452_M1_1_2 ( .A(u4_sll_452_ML_int_1__2_), .B(
        u4_sll_452_ML_int_1__0_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__2_) );
  MUX2_X2 u4_sll_452_M1_1_3 ( .A(u4_sll_452_ML_int_1__3_), .B(
        u4_sll_452_ML_int_1__1_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__3_) );
  MUX2_X2 u4_sll_452_M1_1_4 ( .A(u4_sll_452_ML_int_1__4_), .B(
        u4_sll_452_ML_int_1__2_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__4_) );
  MUX2_X2 u4_sll_452_M1_1_5 ( .A(u4_sll_452_ML_int_1__5_), .B(
        u4_sll_452_ML_int_1__3_), .S(u4_sll_452_n13), .Z(
        u4_sll_452_ML_int_2__5_) );
  MUX2_X2 u4_sll_452_M1_1_6 ( .A(u4_sll_452_ML_int_1__6_), .B(
        u4_sll_452_ML_int_1__4_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__6_) );
  MUX2_X2 u4_sll_452_M1_1_7 ( .A(u4_sll_452_ML_int_1__7_), .B(
        u4_sll_452_ML_int_1__5_), .S(u4_sll_452_n13), .Z(
        u4_sll_452_ML_int_2__7_) );
  MUX2_X2 u4_sll_452_M1_1_8 ( .A(u4_sll_452_ML_int_1__8_), .B(
        u4_sll_452_ML_int_1__6_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__8_) );
  MUX2_X2 u4_sll_452_M1_1_9 ( .A(u4_sll_452_ML_int_1__9_), .B(
        u4_sll_452_ML_int_1__7_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__9_) );
  MUX2_X2 u4_sll_452_M1_1_10 ( .A(u4_sll_452_ML_int_1__10_), .B(
        u4_sll_452_ML_int_1__8_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__10_) );
  MUX2_X2 u4_sll_452_M1_1_11 ( .A(u4_sll_452_ML_int_1__11_), .B(
        u4_sll_452_ML_int_1__9_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__11_) );
  MUX2_X2 u4_sll_452_M1_1_12 ( .A(u4_sll_452_ML_int_1__12_), .B(
        u4_sll_452_ML_int_1__10_), .S(u4_sll_452_n13), .Z(
        u4_sll_452_ML_int_2__12_) );
  MUX2_X2 u4_sll_452_M1_1_13 ( .A(u4_sll_452_ML_int_1__13_), .B(
        u4_sll_452_ML_int_1__11_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__13_) );
  MUX2_X2 u4_sll_452_M1_1_14 ( .A(u4_sll_452_ML_int_1__14_), .B(
        u4_sll_452_ML_int_1__12_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__14_) );
  MUX2_X2 u4_sll_452_M1_1_15 ( .A(u4_sll_452_ML_int_1__15_), .B(
        u4_sll_452_ML_int_1__13_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__15_) );
  MUX2_X2 u4_sll_452_M1_1_16 ( .A(u4_sll_452_ML_int_1__16_), .B(
        u4_sll_452_ML_int_1__14_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__16_) );
  MUX2_X2 u4_sll_452_M1_1_17 ( .A(u4_sll_452_ML_int_1__17_), .B(
        u4_sll_452_ML_int_1__15_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__17_) );
  MUX2_X2 u4_sll_452_M1_1_18 ( .A(u4_sll_452_ML_int_1__18_), .B(
        u4_sll_452_ML_int_1__16_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__18_) );
  MUX2_X2 u4_sll_452_M1_1_19 ( .A(u4_sll_452_ML_int_1__19_), .B(
        u4_sll_452_ML_int_1__17_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__19_) );
  MUX2_X2 u4_sll_452_M1_1_20 ( .A(u4_sll_452_ML_int_1__20_), .B(
        u4_sll_452_ML_int_1__18_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__20_) );
  MUX2_X2 u4_sll_452_M1_1_21 ( .A(u4_sll_452_ML_int_1__21_), .B(
        u4_sll_452_ML_int_1__19_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__21_) );
  MUX2_X2 u4_sll_452_M1_1_22 ( .A(u4_sll_452_ML_int_1__22_), .B(
        u4_sll_452_ML_int_1__20_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__22_) );
  MUX2_X2 u4_sll_452_M1_1_23 ( .A(u4_sll_452_ML_int_1__23_), .B(
        u4_sll_452_ML_int_1__21_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__23_) );
  MUX2_X2 u4_sll_452_M1_1_24 ( .A(u4_sll_452_ML_int_1__24_), .B(
        u4_sll_452_ML_int_1__22_), .S(u4_sll_452_n13), .Z(
        u4_sll_452_ML_int_2__24_) );
  MUX2_X2 u4_sll_452_M1_1_25 ( .A(u4_sll_452_ML_int_1__25_), .B(
        u4_sll_452_ML_int_1__23_), .S(u4_sll_452_n13), .Z(
        u4_sll_452_ML_int_2__25_) );
  MUX2_X2 u4_sll_452_M1_1_26 ( .A(u4_sll_452_ML_int_1__26_), .B(
        u4_sll_452_ML_int_1__24_), .S(u4_sll_452_n13), .Z(
        u4_sll_452_ML_int_2__26_) );
  MUX2_X2 u4_sll_452_M1_1_27 ( .A(u4_sll_452_ML_int_1__27_), .B(
        u4_sll_452_ML_int_1__25_), .S(u4_sll_452_n13), .Z(
        u4_sll_452_ML_int_2__27_) );
  MUX2_X2 u4_sll_452_M1_1_28 ( .A(u4_sll_452_ML_int_1__28_), .B(
        u4_sll_452_ML_int_1__26_), .S(u4_sll_452_n13), .Z(
        u4_sll_452_ML_int_2__28_) );
  MUX2_X2 u4_sll_452_M1_1_29 ( .A(u4_sll_452_ML_int_1__29_), .B(
        u4_sll_452_ML_int_1__27_), .S(u4_sll_452_n13), .Z(
        u4_sll_452_ML_int_2__29_) );
  MUX2_X2 u4_sll_452_M1_1_30 ( .A(u4_sll_452_ML_int_1__30_), .B(
        u4_sll_452_ML_int_1__28_), .S(u4_sll_452_n13), .Z(
        u4_sll_452_ML_int_2__30_) );
  MUX2_X2 u4_sll_452_M1_1_31 ( .A(u4_sll_452_ML_int_1__31_), .B(
        u4_sll_452_ML_int_1__29_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__31_) );
  MUX2_X2 u4_sll_452_M1_1_32 ( .A(u4_sll_452_ML_int_1__32_), .B(
        u4_sll_452_ML_int_1__30_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__32_) );
  MUX2_X2 u4_sll_452_M1_1_33 ( .A(u4_sll_452_ML_int_1__33_), .B(
        u4_sll_452_ML_int_1__31_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__33_) );
  MUX2_X2 u4_sll_452_M1_1_34 ( .A(u4_sll_452_ML_int_1__34_), .B(
        u4_sll_452_ML_int_1__32_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__34_) );
  MUX2_X2 u4_sll_452_M1_1_35 ( .A(u4_sll_452_ML_int_1__35_), .B(
        u4_sll_452_ML_int_1__33_), .S(u4_sll_452_n13), .Z(
        u4_sll_452_ML_int_2__35_) );
  MUX2_X2 u4_sll_452_M1_1_36 ( .A(u4_sll_452_ML_int_1__36_), .B(
        u4_sll_452_ML_int_1__34_), .S(u4_sll_452_n13), .Z(
        u4_sll_452_ML_int_2__36_) );
  MUX2_X2 u4_sll_452_M1_1_37 ( .A(u4_sll_452_ML_int_1__37_), .B(
        u4_sll_452_ML_int_1__35_), .S(u4_sll_452_n13), .Z(
        u4_sll_452_ML_int_2__37_) );
  MUX2_X2 u4_sll_452_M1_1_38 ( .A(u4_sll_452_ML_int_1__38_), .B(
        u4_sll_452_ML_int_1__36_), .S(u4_sll_452_n13), .Z(
        u4_sll_452_ML_int_2__38_) );
  MUX2_X2 u4_sll_452_M1_1_39 ( .A(u4_sll_452_ML_int_1__39_), .B(
        u4_sll_452_ML_int_1__37_), .S(u4_sll_452_n13), .Z(
        u4_sll_452_ML_int_2__39_) );
  MUX2_X2 u4_sll_452_M1_1_40 ( .A(u4_sll_452_ML_int_1__40_), .B(
        u4_sll_452_ML_int_1__38_), .S(u4_sll_452_n13), .Z(
        u4_sll_452_ML_int_2__40_) );
  MUX2_X2 u4_sll_452_M1_1_41 ( .A(u4_sll_452_ML_int_1__41_), .B(
        u4_sll_452_ML_int_1__39_), .S(u4_sll_452_n13), .Z(
        u4_sll_452_ML_int_2__41_) );
  MUX2_X2 u4_sll_452_M1_1_42 ( .A(u4_sll_452_ML_int_1__42_), .B(
        u4_sll_452_ML_int_1__40_), .S(u4_sll_452_n13), .Z(
        u4_sll_452_ML_int_2__42_) );
  MUX2_X2 u4_sll_452_M1_1_43 ( .A(u4_sll_452_ML_int_1__43_), .B(
        u4_sll_452_ML_int_1__41_), .S(u4_sll_452_n13), .Z(
        u4_sll_452_ML_int_2__43_) );
  MUX2_X2 u4_sll_452_M1_1_44 ( .A(u4_sll_452_ML_int_1__44_), .B(
        u4_sll_452_ML_int_1__42_), .S(u4_sll_452_n13), .Z(
        u4_sll_452_ML_int_2__44_) );
  MUX2_X2 u4_sll_452_M1_1_45 ( .A(u4_sll_452_ML_int_1__45_), .B(
        u4_sll_452_ML_int_1__43_), .S(u4_sll_452_n13), .Z(
        u4_sll_452_ML_int_2__45_) );
  MUX2_X2 u4_sll_452_M1_1_46 ( .A(u4_sll_452_ML_int_1__46_), .B(
        u4_sll_452_ML_int_1__44_), .S(u4_sll_452_n10), .Z(
        u4_sll_452_ML_int_2__46_) );
  MUX2_X2 u4_sll_452_M1_1_47 ( .A(u4_sll_452_ML_int_1__47_), .B(
        u4_sll_452_ML_int_1__45_), .S(u4_sll_452_n10), .Z(
        u4_sll_452_ML_int_2__47_) );
  MUX2_X2 u4_sll_452_M1_1_48 ( .A(u4_sll_452_ML_int_1__48_), .B(
        u4_sll_452_ML_int_1__46_), .S(u4_sll_452_n10), .Z(
        u4_sll_452_ML_int_2__48_) );
  MUX2_X2 u4_sll_452_M1_1_49 ( .A(u4_sll_452_ML_int_1__49_), .B(
        u4_sll_452_ML_int_1__47_), .S(u4_sll_452_n10), .Z(
        u4_sll_452_ML_int_2__49_) );
  MUX2_X2 u4_sll_452_M1_1_50 ( .A(u4_sll_452_ML_int_1__50_), .B(
        u4_sll_452_ML_int_1__48_), .S(u4_sll_452_n10), .Z(
        u4_sll_452_ML_int_2__50_) );
  MUX2_X2 u4_sll_452_M1_1_51 ( .A(u4_sll_452_ML_int_1__51_), .B(
        u4_sll_452_ML_int_1__49_), .S(u4_sll_452_n10), .Z(
        u4_sll_452_ML_int_2__51_) );
  MUX2_X2 u4_sll_452_M1_1_52 ( .A(u4_sll_452_ML_int_1__52_), .B(
        u4_sll_452_ML_int_1__50_), .S(u4_sll_452_n10), .Z(
        u4_sll_452_ML_int_2__52_) );
  MUX2_X2 u4_sll_452_M1_1_53 ( .A(u4_sll_452_ML_int_1__53_), .B(
        u4_sll_452_ML_int_1__51_), .S(u4_sll_452_n10), .Z(
        u4_sll_452_ML_int_2__53_) );
  MUX2_X2 u4_sll_452_M1_1_54 ( .A(u4_sll_452_ML_int_1__54_), .B(
        u4_sll_452_ML_int_1__52_), .S(u4_sll_452_n10), .Z(
        u4_sll_452_ML_int_2__54_) );
  MUX2_X2 u4_sll_452_M1_1_55 ( .A(u4_sll_452_ML_int_1__55_), .B(
        u4_sll_452_ML_int_1__53_), .S(u4_sll_452_n10), .Z(
        u4_sll_452_ML_int_2__55_) );
  MUX2_X2 u4_sll_452_M1_1_56 ( .A(u4_sll_452_ML_int_1__56_), .B(
        u4_sll_452_ML_int_1__54_), .S(u4_sll_452_n10), .Z(
        u4_sll_452_ML_int_2__56_) );
  MUX2_X2 u4_sll_452_M1_1_57 ( .A(u4_sll_452_ML_int_1__57_), .B(
        u4_sll_452_ML_int_1__55_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__57_) );
  MUX2_X2 u4_sll_452_M1_1_58 ( .A(u4_sll_452_ML_int_1__58_), .B(
        u4_sll_452_ML_int_1__56_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__58_) );
  MUX2_X2 u4_sll_452_M1_1_59 ( .A(u4_sll_452_ML_int_1__59_), .B(
        u4_sll_452_ML_int_1__57_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__59_) );
  MUX2_X2 u4_sll_452_M1_1_60 ( .A(u4_sll_452_ML_int_1__60_), .B(
        u4_sll_452_ML_int_1__58_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__60_) );
  MUX2_X2 u4_sll_452_M1_1_61 ( .A(u4_sll_452_ML_int_1__61_), .B(
        u4_sll_452_ML_int_1__59_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__61_) );
  MUX2_X2 u4_sll_452_M1_1_62 ( .A(u4_sll_452_ML_int_1__62_), .B(
        u4_sll_452_ML_int_1__60_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__62_) );
  MUX2_X2 u4_sll_452_M1_1_63 ( .A(u4_sll_452_ML_int_1__63_), .B(
        u4_sll_452_ML_int_1__61_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__63_) );
  MUX2_X2 u4_sll_452_M1_1_64 ( .A(u4_sll_452_ML_int_1__64_), .B(
        u4_sll_452_ML_int_1__62_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__64_) );
  MUX2_X2 u4_sll_452_M1_1_65 ( .A(u4_sll_452_ML_int_1__65_), .B(
        u4_sll_452_ML_int_1__63_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__65_) );
  MUX2_X2 u4_sll_452_M1_1_66 ( .A(u4_sll_452_ML_int_1__66_), .B(
        u4_sll_452_ML_int_1__64_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__66_) );
  MUX2_X2 u4_sll_452_M1_1_67 ( .A(u4_sll_452_ML_int_1__67_), .B(
        u4_sll_452_ML_int_1__65_), .S(u4_sll_452_n10), .Z(
        u4_sll_452_ML_int_2__67_) );
  MUX2_X2 u4_sll_452_M1_1_68 ( .A(u4_sll_452_ML_int_1__68_), .B(
        u4_sll_452_ML_int_1__66_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__68_) );
  MUX2_X2 u4_sll_452_M1_1_69 ( .A(u4_sll_452_ML_int_1__69_), .B(
        u4_sll_452_ML_int_1__67_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__69_) );
  MUX2_X2 u4_sll_452_M1_1_70 ( .A(u4_sll_452_ML_int_1__70_), .B(
        u4_sll_452_ML_int_1__68_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__70_) );
  MUX2_X2 u4_sll_452_M1_1_71 ( .A(u4_sll_452_ML_int_1__71_), .B(
        u4_sll_452_ML_int_1__69_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__71_) );
  MUX2_X2 u4_sll_452_M1_1_72 ( .A(u4_sll_452_ML_int_1__72_), .B(
        u4_sll_452_ML_int_1__70_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__72_) );
  MUX2_X2 u4_sll_452_M1_1_73 ( .A(u4_sll_452_ML_int_1__73_), .B(
        u4_sll_452_ML_int_1__71_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__73_) );
  MUX2_X2 u4_sll_452_M1_1_74 ( .A(u4_sll_452_ML_int_1__74_), .B(
        u4_sll_452_ML_int_1__72_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__74_) );
  MUX2_X2 u4_sll_452_M1_1_75 ( .A(u4_sll_452_ML_int_1__75_), .B(
        u4_sll_452_ML_int_1__73_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__75_) );
  MUX2_X2 u4_sll_452_M1_1_76 ( .A(u4_sll_452_ML_int_1__76_), .B(
        u4_sll_452_ML_int_1__74_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__76_) );
  MUX2_X2 u4_sll_452_M1_1_77 ( .A(u4_sll_452_ML_int_1__77_), .B(
        u4_sll_452_ML_int_1__75_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__77_) );
  MUX2_X2 u4_sll_452_M1_1_78 ( .A(u4_sll_452_ML_int_1__78_), .B(
        u4_sll_452_ML_int_1__76_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__78_) );
  MUX2_X2 u4_sll_452_M1_1_79 ( .A(u4_sll_452_ML_int_1__79_), .B(
        u4_sll_452_ML_int_1__77_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__79_) );
  MUX2_X2 u4_sll_452_M1_1_80 ( .A(u4_sll_452_ML_int_1__80_), .B(
        u4_sll_452_ML_int_1__78_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__80_) );
  MUX2_X2 u4_sll_452_M1_1_81 ( .A(u4_sll_452_ML_int_1__81_), .B(
        u4_sll_452_ML_int_1__79_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__81_) );
  MUX2_X2 u4_sll_452_M1_1_82 ( .A(u4_sll_452_ML_int_1__82_), .B(
        u4_sll_452_ML_int_1__80_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__82_) );
  MUX2_X2 u4_sll_452_M1_1_83 ( .A(u4_sll_452_ML_int_1__83_), .B(
        u4_sll_452_ML_int_1__81_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__83_) );
  MUX2_X2 u4_sll_452_M1_1_84 ( .A(u4_sll_452_ML_int_1__84_), .B(
        u4_sll_452_ML_int_1__82_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__84_) );
  MUX2_X2 u4_sll_452_M1_1_85 ( .A(u4_sll_452_ML_int_1__85_), .B(
        u4_sll_452_ML_int_1__83_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__85_) );
  MUX2_X2 u4_sll_452_M1_1_86 ( .A(u4_sll_452_ML_int_1__86_), .B(
        u4_sll_452_ML_int_1__84_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__86_) );
  MUX2_X2 u4_sll_452_M1_1_87 ( .A(u4_sll_452_ML_int_1__87_), .B(
        u4_sll_452_ML_int_1__85_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__87_) );
  MUX2_X2 u4_sll_452_M1_1_88 ( .A(u4_sll_452_ML_int_1__88_), .B(
        u4_sll_452_ML_int_1__86_), .S(u4_sll_452_n13), .Z(
        u4_sll_452_ML_int_2__88_) );
  MUX2_X2 u4_sll_452_M1_1_89 ( .A(u4_sll_452_ML_int_1__89_), .B(
        u4_sll_452_ML_int_1__87_), .S(u4_sll_452_n12), .Z(
        u4_sll_452_ML_int_2__89_) );
  MUX2_X2 u4_sll_452_M1_1_90 ( .A(u4_sll_452_ML_int_1__90_), .B(
        u4_sll_452_ML_int_1__88_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__90_) );
  MUX2_X2 u4_sll_452_M1_1_91 ( .A(u4_sll_452_ML_int_1__91_), .B(
        u4_sll_452_ML_int_1__89_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__91_) );
  MUX2_X2 u4_sll_452_M1_1_92 ( .A(u4_sll_452_ML_int_1__92_), .B(
        u4_sll_452_ML_int_1__90_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__92_) );
  MUX2_X2 u4_sll_452_M1_1_93 ( .A(u4_sll_452_ML_int_1__93_), .B(
        u4_sll_452_ML_int_1__91_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__93_) );
  MUX2_X2 u4_sll_452_M1_1_94 ( .A(u4_sll_452_ML_int_1__94_), .B(
        u4_sll_452_ML_int_1__92_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__94_) );
  MUX2_X2 u4_sll_452_M1_1_95 ( .A(u4_sll_452_ML_int_1__95_), .B(
        u4_sll_452_ML_int_1__93_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__95_) );
  MUX2_X2 u4_sll_452_M1_1_96 ( .A(u4_sll_452_ML_int_1__96_), .B(
        u4_sll_452_ML_int_1__94_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__96_) );
  MUX2_X2 u4_sll_452_M1_1_97 ( .A(u4_sll_452_ML_int_1__97_), .B(
        u4_sll_452_ML_int_1__95_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__97_) );
  MUX2_X2 u4_sll_452_M1_1_98 ( .A(u4_sll_452_ML_int_1__98_), .B(
        u4_sll_452_ML_int_1__96_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__98_) );
  MUX2_X2 u4_sll_452_M1_1_99 ( .A(u4_sll_452_ML_int_1__99_), .B(
        u4_sll_452_ML_int_1__97_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__99_) );
  MUX2_X2 u4_sll_452_M1_1_100 ( .A(u4_sll_452_ML_int_1__100_), .B(
        u4_sll_452_ML_int_1__98_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__100_) );
  MUX2_X2 u4_sll_452_M1_1_101 ( .A(u4_sll_452_ML_int_1__101_), .B(
        u4_sll_452_ML_int_1__99_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__101_) );
  MUX2_X2 u4_sll_452_M1_1_102 ( .A(u4_sll_452_ML_int_1__102_), .B(
        u4_sll_452_ML_int_1__100_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__102_) );
  MUX2_X2 u4_sll_452_M1_1_103 ( .A(u4_sll_452_ML_int_1__103_), .B(
        u4_sll_452_ML_int_1__101_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__103_) );
  MUX2_X2 u4_sll_452_M1_1_104 ( .A(u4_sll_452_ML_int_1__104_), .B(
        u4_sll_452_ML_int_1__102_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__104_) );
  MUX2_X2 u4_sll_452_M1_1_105 ( .A(u4_sll_452_ML_int_1__105_), .B(
        u4_sll_452_ML_int_1__103_), .S(u4_sll_452_n11), .Z(
        u4_sll_452_ML_int_2__105_) );
  MUX2_X2 u4_sll_452_M1_2_4 ( .A(u4_sll_452_ML_int_2__4_), .B(
        u4_sll_452_ML_int_2__0_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__4_) );
  MUX2_X2 u4_sll_452_M1_2_5 ( .A(u4_sll_452_ML_int_2__5_), .B(
        u4_sll_452_ML_int_2__1_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__5_) );
  MUX2_X2 u4_sll_452_M1_2_6 ( .A(u4_sll_452_ML_int_2__6_), .B(
        u4_sll_452_ML_int_2__2_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__6_) );
  MUX2_X2 u4_sll_452_M1_2_7 ( .A(u4_sll_452_ML_int_2__7_), .B(
        u4_sll_452_ML_int_2__3_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__7_) );
  MUX2_X2 u4_sll_452_M1_2_8 ( .A(u4_sll_452_ML_int_2__8_), .B(
        u4_sll_452_ML_int_2__4_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__8_) );
  MUX2_X2 u4_sll_452_M1_2_9 ( .A(u4_sll_452_ML_int_2__9_), .B(
        u4_sll_452_ML_int_2__5_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__9_) );
  MUX2_X2 u4_sll_452_M1_2_10 ( .A(u4_sll_452_ML_int_2__10_), .B(
        u4_sll_452_ML_int_2__6_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__10_) );
  MUX2_X2 u4_sll_452_M1_2_11 ( .A(u4_sll_452_ML_int_2__11_), .B(
        u4_sll_452_ML_int_2__7_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__11_) );
  MUX2_X2 u4_sll_452_M1_2_12 ( .A(u4_sll_452_ML_int_2__12_), .B(
        u4_sll_452_ML_int_2__8_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__12_) );
  MUX2_X2 u4_sll_452_M1_2_13 ( .A(u4_sll_452_ML_int_2__13_), .B(
        u4_sll_452_ML_int_2__9_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__13_) );
  MUX2_X2 u4_sll_452_M1_2_14 ( .A(u4_sll_452_ML_int_2__14_), .B(
        u4_sll_452_ML_int_2__10_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__14_) );
  MUX2_X2 u4_sll_452_M1_2_15 ( .A(u4_sll_452_ML_int_2__15_), .B(
        u4_sll_452_ML_int_2__11_), .S(u4_sll_452_n14), .Z(
        u4_sll_452_ML_int_3__15_) );
  MUX2_X2 u4_sll_452_M1_2_16 ( .A(u4_sll_452_ML_int_2__16_), .B(
        u4_sll_452_ML_int_2__12_), .S(u4_sll_452_n14), .Z(
        u4_sll_452_ML_int_3__16_) );
  MUX2_X2 u4_sll_452_M1_2_17 ( .A(u4_sll_452_ML_int_2__17_), .B(
        u4_sll_452_ML_int_2__13_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__17_) );
  MUX2_X2 u4_sll_452_M1_2_18 ( .A(u4_sll_452_ML_int_2__18_), .B(
        u4_sll_452_ML_int_2__14_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__18_) );
  MUX2_X2 u4_sll_452_M1_2_19 ( .A(u4_sll_452_ML_int_2__19_), .B(
        u4_sll_452_ML_int_2__15_), .S(u4_sll_452_n16), .Z(
        u4_sll_452_ML_int_3__19_) );
  MUX2_X2 u4_sll_452_M1_2_20 ( .A(u4_sll_452_ML_int_2__20_), .B(
        u4_sll_452_ML_int_2__16_), .S(u4_sll_452_n16), .Z(
        u4_sll_452_ML_int_3__20_) );
  MUX2_X2 u4_sll_452_M1_2_21 ( .A(u4_sll_452_ML_int_2__21_), .B(
        u4_sll_452_ML_int_2__17_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__21_) );
  MUX2_X2 u4_sll_452_M1_2_22 ( .A(u4_sll_452_ML_int_2__22_), .B(
        u4_sll_452_ML_int_2__18_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__22_) );
  MUX2_X2 u4_sll_452_M1_2_23 ( .A(u4_sll_452_ML_int_2__23_), .B(
        u4_sll_452_ML_int_2__19_), .S(u4_sll_452_n14), .Z(
        u4_sll_452_ML_int_3__23_) );
  MUX2_X2 u4_sll_452_M1_2_24 ( .A(u4_sll_452_ML_int_2__24_), .B(
        u4_sll_452_ML_int_2__20_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__24_) );
  MUX2_X2 u4_sll_452_M1_2_25 ( .A(u4_sll_452_ML_int_2__25_), .B(
        u4_sll_452_ML_int_2__21_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__25_) );
  MUX2_X2 u4_sll_452_M1_2_26 ( .A(u4_sll_452_ML_int_2__26_), .B(
        u4_sll_452_ML_int_2__22_), .S(u4_sll_452_n16), .Z(
        u4_sll_452_ML_int_3__26_) );
  MUX2_X2 u4_sll_452_M1_2_27 ( .A(u4_sll_452_ML_int_2__27_), .B(
        u4_sll_452_ML_int_2__23_), .S(u4_sll_452_n16), .Z(
        u4_sll_452_ML_int_3__27_) );
  MUX2_X2 u4_sll_452_M1_2_28 ( .A(u4_sll_452_ML_int_2__28_), .B(
        u4_sll_452_ML_int_2__24_), .S(u4_sll_452_n16), .Z(
        u4_sll_452_ML_int_3__28_) );
  MUX2_X2 u4_sll_452_M1_2_29 ( .A(u4_sll_452_ML_int_2__29_), .B(
        u4_sll_452_ML_int_2__25_), .S(u4_sll_452_n16), .Z(
        u4_sll_452_ML_int_3__29_) );
  MUX2_X2 u4_sll_452_M1_2_30 ( .A(u4_sll_452_ML_int_2__30_), .B(
        u4_sll_452_ML_int_2__26_), .S(u4_sll_452_n16), .Z(
        u4_sll_452_ML_int_3__30_) );
  MUX2_X2 u4_sll_452_M1_2_31 ( .A(u4_sll_452_ML_int_2__31_), .B(
        u4_sll_452_ML_int_2__27_), .S(u4_sll_452_n16), .Z(
        u4_sll_452_ML_int_3__31_) );
  MUX2_X2 u4_sll_452_M1_2_32 ( .A(u4_sll_452_ML_int_2__32_), .B(
        u4_sll_452_ML_int_2__28_), .S(u4_sll_452_n16), .Z(
        u4_sll_452_ML_int_3__32_) );
  MUX2_X2 u4_sll_452_M1_2_33 ( .A(u4_sll_452_ML_int_2__33_), .B(
        u4_sll_452_ML_int_2__29_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__33_) );
  MUX2_X2 u4_sll_452_M1_2_34 ( .A(u4_sll_452_ML_int_2__34_), .B(
        u4_sll_452_ML_int_2__30_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__34_) );
  MUX2_X2 u4_sll_452_M1_2_35 ( .A(u4_sll_452_ML_int_2__35_), .B(
        u4_sll_452_ML_int_2__31_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__35_) );
  MUX2_X2 u4_sll_452_M1_2_36 ( .A(u4_sll_452_ML_int_2__36_), .B(
        u4_sll_452_ML_int_2__32_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__36_) );
  MUX2_X2 u4_sll_452_M1_2_37 ( .A(u4_sll_452_ML_int_2__37_), .B(
        u4_sll_452_ML_int_2__33_), .S(u4_sll_452_n16), .Z(
        u4_sll_452_ML_int_3__37_) );
  MUX2_X2 u4_sll_452_M1_2_38 ( .A(u4_sll_452_ML_int_2__38_), .B(
        u4_sll_452_ML_int_2__34_), .S(u4_sll_452_n16), .Z(
        u4_sll_452_ML_int_3__38_) );
  MUX2_X2 u4_sll_452_M1_2_39 ( .A(u4_sll_452_ML_int_2__39_), .B(
        u4_sll_452_ML_int_2__35_), .S(u4_sll_452_n16), .Z(
        u4_sll_452_ML_int_3__39_) );
  MUX2_X2 u4_sll_452_M1_2_40 ( .A(u4_sll_452_ML_int_2__40_), .B(
        u4_sll_452_ML_int_2__36_), .S(u4_sll_452_n16), .Z(
        u4_sll_452_ML_int_3__40_) );
  MUX2_X2 u4_sll_452_M1_2_41 ( .A(u4_sll_452_ML_int_2__41_), .B(
        u4_sll_452_ML_int_2__37_), .S(u4_sll_452_n16), .Z(
        u4_sll_452_ML_int_3__41_) );
  MUX2_X2 u4_sll_452_M1_2_42 ( .A(u4_sll_452_ML_int_2__42_), .B(
        u4_sll_452_ML_int_2__38_), .S(u4_sll_452_n16), .Z(
        u4_sll_452_ML_int_3__42_) );
  MUX2_X2 u4_sll_452_M1_2_43 ( .A(u4_sll_452_ML_int_2__43_), .B(
        u4_sll_452_ML_int_2__39_), .S(u4_sll_452_n16), .Z(
        u4_sll_452_ML_int_3__43_) );
  MUX2_X2 u4_sll_452_M1_2_44 ( .A(u4_sll_452_ML_int_2__44_), .B(
        u4_sll_452_ML_int_2__40_), .S(u4_sll_452_n16), .Z(
        u4_sll_452_ML_int_3__44_) );
  MUX2_X2 u4_sll_452_M1_2_45 ( .A(u4_sll_452_ML_int_2__45_), .B(
        u4_sll_452_ML_int_2__41_), .S(u4_sll_452_n16), .Z(
        u4_sll_452_ML_int_3__45_) );
  MUX2_X2 u4_sll_452_M1_2_46 ( .A(u4_sll_452_ML_int_2__46_), .B(
        u4_sll_452_ML_int_2__42_), .S(u4_sll_452_n16), .Z(
        u4_sll_452_ML_int_3__46_) );
  MUX2_X2 u4_sll_452_M1_2_47 ( .A(u4_sll_452_ML_int_2__47_), .B(
        u4_sll_452_ML_int_2__43_), .S(u4_sll_452_n16), .Z(
        u4_sll_452_ML_int_3__47_) );
  MUX2_X2 u4_sll_452_M1_2_48 ( .A(u4_sll_452_ML_int_2__48_), .B(
        u4_sll_452_ML_int_2__44_), .S(u4_sll_452_n14), .Z(
        u4_sll_452_ML_int_3__48_) );
  MUX2_X2 u4_sll_452_M1_2_49 ( .A(u4_sll_452_ML_int_2__49_), .B(
        u4_sll_452_ML_int_2__45_), .S(u4_sll_452_n14), .Z(
        u4_sll_452_ML_int_3__49_) );
  MUX2_X2 u4_sll_452_M1_2_50 ( .A(u4_sll_452_ML_int_2__50_), .B(
        u4_sll_452_ML_int_2__46_), .S(u4_sll_452_n14), .Z(
        u4_sll_452_ML_int_3__50_) );
  MUX2_X2 u4_sll_452_M1_2_51 ( .A(u4_sll_452_ML_int_2__51_), .B(
        u4_sll_452_ML_int_2__47_), .S(u4_sll_452_n14), .Z(
        u4_sll_452_ML_int_3__51_) );
  MUX2_X2 u4_sll_452_M1_2_52 ( .A(u4_sll_452_ML_int_2__52_), .B(
        u4_sll_452_ML_int_2__48_), .S(u4_sll_452_n14), .Z(
        u4_sll_452_ML_int_3__52_) );
  MUX2_X2 u4_sll_452_M1_2_53 ( .A(u4_sll_452_ML_int_2__53_), .B(
        u4_sll_452_ML_int_2__49_), .S(u4_sll_452_n14), .Z(
        u4_sll_452_ML_int_3__53_) );
  MUX2_X2 u4_sll_452_M1_2_54 ( .A(u4_sll_452_ML_int_2__54_), .B(
        u4_sll_452_ML_int_2__50_), .S(u4_sll_452_n14), .Z(
        u4_sll_452_ML_int_3__54_) );
  MUX2_X2 u4_sll_452_M1_2_55 ( .A(u4_sll_452_ML_int_2__55_), .B(
        u4_sll_452_ML_int_2__51_), .S(u4_sll_452_n14), .Z(
        u4_sll_452_ML_int_3__55_) );
  MUX2_X2 u4_sll_452_M1_2_56 ( .A(u4_sll_452_ML_int_2__56_), .B(
        u4_sll_452_ML_int_2__52_), .S(u4_sll_452_n14), .Z(
        u4_sll_452_ML_int_3__56_) );
  MUX2_X2 u4_sll_452_M1_2_57 ( .A(u4_sll_452_ML_int_2__57_), .B(
        u4_sll_452_ML_int_2__53_), .S(u4_sll_452_n14), .Z(
        u4_sll_452_ML_int_3__57_) );
  MUX2_X2 u4_sll_452_M1_2_58 ( .A(u4_sll_452_ML_int_2__58_), .B(
        u4_sll_452_ML_int_2__54_), .S(u4_sll_452_n14), .Z(
        u4_sll_452_ML_int_3__58_) );
  MUX2_X2 u4_sll_452_M1_2_59 ( .A(u4_sll_452_ML_int_2__59_), .B(
        u4_sll_452_ML_int_2__55_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__59_) );
  MUX2_X2 u4_sll_452_M1_2_60 ( .A(u4_sll_452_ML_int_2__60_), .B(
        u4_sll_452_ML_int_2__56_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__60_) );
  MUX2_X2 u4_sll_452_M1_2_61 ( .A(u4_sll_452_ML_int_2__61_), .B(
        u4_sll_452_ML_int_2__57_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__61_) );
  MUX2_X2 u4_sll_452_M1_2_62 ( .A(u4_sll_452_ML_int_2__62_), .B(
        u4_sll_452_ML_int_2__58_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__62_) );
  MUX2_X2 u4_sll_452_M1_2_63 ( .A(u4_sll_452_ML_int_2__63_), .B(
        u4_sll_452_ML_int_2__59_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__63_) );
  MUX2_X2 u4_sll_452_M1_2_64 ( .A(u4_sll_452_ML_int_2__64_), .B(
        u4_sll_452_ML_int_2__60_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__64_) );
  MUX2_X2 u4_sll_452_M1_2_65 ( .A(u4_sll_452_ML_int_2__65_), .B(
        u4_sll_452_ML_int_2__61_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__65_) );
  MUX2_X2 u4_sll_452_M1_2_66 ( .A(u4_sll_452_ML_int_2__66_), .B(
        u4_sll_452_ML_int_2__62_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__66_) );
  MUX2_X2 u4_sll_452_M1_2_67 ( .A(u4_sll_452_ML_int_2__67_), .B(
        u4_sll_452_ML_int_2__63_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__67_) );
  MUX2_X2 u4_sll_452_M1_2_68 ( .A(u4_sll_452_ML_int_2__68_), .B(
        u4_sll_452_ML_int_2__64_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__68_) );
  MUX2_X2 u4_sll_452_M1_2_69 ( .A(u4_sll_452_ML_int_2__69_), .B(
        u4_sll_452_ML_int_2__65_), .S(u4_sll_452_n14), .Z(
        u4_sll_452_ML_int_3__69_) );
  MUX2_X2 u4_sll_452_M1_2_70 ( .A(u4_sll_452_ML_int_2__70_), .B(
        u4_sll_452_ML_int_2__66_), .S(u4_sll_452_n16), .Z(
        u4_sll_452_ML_int_3__70_) );
  MUX2_X2 u4_sll_452_M1_2_71 ( .A(u4_sll_452_ML_int_2__71_), .B(
        u4_sll_452_ML_int_2__67_), .S(u4_sll_452_n14), .Z(
        u4_sll_452_ML_int_3__71_) );
  MUX2_X2 u4_sll_452_M1_2_72 ( .A(u4_sll_452_ML_int_2__72_), .B(
        u4_sll_452_ML_int_2__68_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__72_) );
  MUX2_X2 u4_sll_452_M1_2_73 ( .A(u4_sll_452_ML_int_2__73_), .B(
        u4_sll_452_ML_int_2__69_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__73_) );
  MUX2_X2 u4_sll_452_M1_2_74 ( .A(u4_sll_452_ML_int_2__74_), .B(
        u4_sll_452_ML_int_2__70_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__74_) );
  MUX2_X2 u4_sll_452_M1_2_75 ( .A(u4_sll_452_ML_int_2__75_), .B(
        u4_sll_452_ML_int_2__71_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__75_) );
  MUX2_X2 u4_sll_452_M1_2_76 ( .A(u4_sll_452_ML_int_2__76_), .B(
        u4_sll_452_ML_int_2__72_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__76_) );
  MUX2_X2 u4_sll_452_M1_2_77 ( .A(u4_sll_452_ML_int_2__77_), .B(
        u4_sll_452_ML_int_2__73_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__77_) );
  MUX2_X2 u4_sll_452_M1_2_78 ( .A(u4_sll_452_ML_int_2__78_), .B(
        u4_sll_452_ML_int_2__74_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__78_) );
  MUX2_X2 u4_sll_452_M1_2_79 ( .A(u4_sll_452_ML_int_2__79_), .B(
        u4_sll_452_ML_int_2__75_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__79_) );
  MUX2_X2 u4_sll_452_M1_2_80 ( .A(u4_sll_452_ML_int_2__80_), .B(
        u4_sll_452_ML_int_2__76_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__80_) );
  MUX2_X2 u4_sll_452_M1_2_81 ( .A(u4_sll_452_ML_int_2__81_), .B(
        u4_sll_452_ML_int_2__77_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__81_) );
  MUX2_X2 u4_sll_452_M1_2_82 ( .A(u4_sll_452_ML_int_2__82_), .B(
        u4_sll_452_ML_int_2__78_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__82_) );
  MUX2_X2 u4_sll_452_M1_2_83 ( .A(u4_sll_452_ML_int_2__83_), .B(
        u4_sll_452_ML_int_2__79_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__83_) );
  MUX2_X2 u4_sll_452_M1_2_84 ( .A(u4_sll_452_ML_int_2__84_), .B(
        u4_sll_452_ML_int_2__80_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__84_) );
  MUX2_X2 u4_sll_452_M1_2_85 ( .A(u4_sll_452_ML_int_2__85_), .B(
        u4_sll_452_ML_int_2__81_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__85_) );
  MUX2_X2 u4_sll_452_M1_2_86 ( .A(u4_sll_452_ML_int_2__86_), .B(
        u4_sll_452_ML_int_2__82_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__86_) );
  MUX2_X2 u4_sll_452_M1_2_87 ( .A(u4_sll_452_ML_int_2__87_), .B(
        u4_sll_452_ML_int_2__83_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__87_) );
  MUX2_X2 u4_sll_452_M1_2_88 ( .A(u4_sll_452_ML_int_2__88_), .B(
        u4_sll_452_ML_int_2__84_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__88_) );
  MUX2_X2 u4_sll_452_M1_2_89 ( .A(u4_sll_452_ML_int_2__89_), .B(
        u4_sll_452_ML_int_2__85_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__89_) );
  MUX2_X2 u4_sll_452_M1_2_90 ( .A(u4_sll_452_ML_int_2__90_), .B(
        u4_sll_452_ML_int_2__86_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__90_) );
  MUX2_X2 u4_sll_452_M1_2_91 ( .A(u4_sll_452_ML_int_2__91_), .B(
        u4_sll_452_ML_int_2__87_), .S(u4_sll_452_n17), .Z(
        u4_sll_452_ML_int_3__91_) );
  MUX2_X2 u4_sll_452_M1_2_92 ( .A(u4_sll_452_ML_int_2__92_), .B(
        u4_sll_452_ML_int_2__88_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__92_) );
  MUX2_X2 u4_sll_452_M1_2_93 ( .A(u4_sll_452_ML_int_2__93_), .B(
        u4_sll_452_ML_int_2__89_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__93_) );
  MUX2_X2 u4_sll_452_M1_2_94 ( .A(u4_sll_452_ML_int_2__94_), .B(
        u4_sll_452_ML_int_2__90_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__94_) );
  MUX2_X2 u4_sll_452_M1_2_95 ( .A(u4_sll_452_ML_int_2__95_), .B(
        u4_sll_452_ML_int_2__91_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__95_) );
  MUX2_X2 u4_sll_452_M1_2_96 ( .A(u4_sll_452_ML_int_2__96_), .B(
        u4_sll_452_ML_int_2__92_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__96_) );
  MUX2_X2 u4_sll_452_M1_2_97 ( .A(u4_sll_452_ML_int_2__97_), .B(
        u4_sll_452_ML_int_2__93_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__97_) );
  MUX2_X2 u4_sll_452_M1_2_98 ( .A(u4_sll_452_ML_int_2__98_), .B(
        u4_sll_452_ML_int_2__94_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__98_) );
  MUX2_X2 u4_sll_452_M1_2_99 ( .A(u4_sll_452_ML_int_2__99_), .B(
        u4_sll_452_ML_int_2__95_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__99_) );
  MUX2_X2 u4_sll_452_M1_2_100 ( .A(u4_sll_452_ML_int_2__100_), .B(
        u4_sll_452_ML_int_2__96_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__100_) );
  MUX2_X2 u4_sll_452_M1_2_101 ( .A(u4_sll_452_ML_int_2__101_), .B(
        u4_sll_452_ML_int_2__97_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__101_) );
  MUX2_X2 u4_sll_452_M1_2_102 ( .A(u4_sll_452_ML_int_2__102_), .B(
        u4_sll_452_ML_int_2__98_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__102_) );
  MUX2_X2 u4_sll_452_M1_2_103 ( .A(u4_sll_452_ML_int_2__103_), .B(
        u4_sll_452_ML_int_2__99_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__103_) );
  MUX2_X2 u4_sll_452_M1_2_104 ( .A(u4_sll_452_ML_int_2__104_), .B(
        u4_sll_452_ML_int_2__100_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__104_) );
  MUX2_X2 u4_sll_452_M1_2_105 ( .A(u4_sll_452_ML_int_2__105_), .B(
        u4_sll_452_ML_int_2__101_), .S(u4_sll_452_n15), .Z(
        u4_sll_452_ML_int_3__105_) );
  MUX2_X2 u4_sll_452_M1_3_8 ( .A(u4_sll_452_ML_int_3__8_), .B(
        u4_sll_452_ML_int_3__0_), .S(u4_sll_452_n22), .Z(
        u4_sll_452_ML_int_4__8_) );
  MUX2_X2 u4_sll_452_M1_3_9 ( .A(u4_sll_452_ML_int_3__9_), .B(
        u4_sll_452_ML_int_3__1_), .S(u4_sll_452_n22), .Z(
        u4_sll_452_ML_int_4__9_) );
  MUX2_X2 u4_sll_452_M1_3_10 ( .A(u4_sll_452_ML_int_3__10_), .B(
        u4_sll_452_ML_int_3__2_), .S(u4_sll_452_n22), .Z(
        u4_sll_452_ML_int_4__10_) );
  MUX2_X2 u4_sll_452_M1_3_11 ( .A(u4_sll_452_ML_int_3__11_), .B(
        u4_sll_452_ML_int_3__3_), .S(u4_sll_452_n22), .Z(
        u4_sll_452_ML_int_4__11_) );
  MUX2_X2 u4_sll_452_M1_3_12 ( .A(u4_sll_452_ML_int_3__12_), .B(
        u4_sll_452_ML_int_3__4_), .S(u4_sll_452_n22), .Z(
        u4_sll_452_ML_int_4__12_) );
  MUX2_X2 u4_sll_452_M1_3_13 ( .A(u4_sll_452_ML_int_3__13_), .B(
        u4_sll_452_ML_int_3__5_), .S(u4_sll_452_n22), .Z(
        u4_sll_452_ML_int_4__13_) );
  MUX2_X2 u4_sll_452_M1_3_14 ( .A(u4_sll_452_ML_int_3__14_), .B(
        u4_sll_452_ML_int_3__6_), .S(u4_sll_452_n22), .Z(
        u4_sll_452_ML_int_4__14_) );
  MUX2_X2 u4_sll_452_M1_3_15 ( .A(u4_sll_452_ML_int_3__15_), .B(
        u4_sll_452_ML_int_3__7_), .S(u4_sll_452_n22), .Z(
        u4_sll_452_ML_int_4__15_) );
  MUX2_X2 u4_sll_452_M1_3_16 ( .A(u4_sll_452_ML_int_3__16_), .B(
        u4_sll_452_ML_int_3__8_), .S(u4_sll_452_n22), .Z(
        u4_sll_452_ML_int_4__16_) );
  MUX2_X2 u4_sll_452_M1_3_17 ( .A(u4_sll_452_ML_int_3__17_), .B(
        u4_sll_452_ML_int_3__9_), .S(u4_sll_452_n22), .Z(
        u4_sll_452_ML_int_4__17_) );
  MUX2_X2 u4_sll_452_M1_3_18 ( .A(u4_sll_452_ML_int_3__18_), .B(
        u4_sll_452_ML_int_3__10_), .S(u4_sll_452_n21), .Z(
        u4_sll_452_ML_int_4__18_) );
  MUX2_X2 u4_sll_452_M1_3_19 ( .A(u4_sll_452_ML_int_3__19_), .B(
        u4_sll_452_ML_int_3__11_), .S(u4_sll_452_n19), .Z(
        u4_sll_452_ML_int_4__19_) );
  MUX2_X2 u4_sll_452_M1_3_20 ( .A(u4_sll_452_ML_int_3__20_), .B(
        u4_sll_452_ML_int_3__12_), .S(u4_sll_452_n21), .Z(
        u4_sll_452_ML_int_4__20_) );
  MUX2_X2 u4_sll_452_M1_3_21 ( .A(u4_sll_452_ML_int_3__21_), .B(
        u4_sll_452_ML_int_3__13_), .S(u4_sll_452_n21), .Z(
        u4_sll_452_ML_int_4__21_) );
  MUX2_X2 u4_sll_452_M1_3_22 ( .A(u4_sll_452_ML_int_3__22_), .B(
        u4_sll_452_ML_int_3__14_), .S(u4_sll_452_n22), .Z(
        u4_sll_452_ML_int_4__22_) );
  MUX2_X2 u4_sll_452_M1_3_23 ( .A(u4_sll_452_ML_int_3__23_), .B(
        u4_sll_452_ML_int_3__15_), .S(u4_sll_452_n22), .Z(
        u4_sll_452_ML_int_4__23_) );
  MUX2_X2 u4_sll_452_M1_3_24 ( .A(u4_sll_452_ML_int_3__24_), .B(
        u4_sll_452_ML_int_3__16_), .S(u4_sll_452_n22), .Z(
        u4_sll_452_ML_int_4__24_) );
  MUX2_X2 u4_sll_452_M1_3_25 ( .A(u4_sll_452_ML_int_3__25_), .B(
        u4_sll_452_ML_int_3__17_), .S(u4_sll_452_n22), .Z(
        u4_sll_452_ML_int_4__25_) );
  MUX2_X2 u4_sll_452_M1_3_26 ( .A(u4_sll_452_ML_int_3__26_), .B(
        u4_sll_452_ML_int_3__18_), .S(u4_sll_452_n22), .Z(
        u4_sll_452_ML_int_4__26_) );
  MUX2_X2 u4_sll_452_M1_3_27 ( .A(u4_sll_452_ML_int_3__27_), .B(
        u4_sll_452_ML_int_3__19_), .S(u4_sll_452_n22), .Z(
        u4_sll_452_ML_int_4__27_) );
  MUX2_X2 u4_sll_452_M1_3_28 ( .A(u4_sll_452_ML_int_3__28_), .B(
        u4_sll_452_ML_int_3__20_), .S(u4_sll_452_n22), .Z(
        u4_sll_452_ML_int_4__28_) );
  MUX2_X2 u4_sll_452_M1_3_29 ( .A(u4_sll_452_ML_int_3__29_), .B(
        u4_sll_452_ML_int_3__21_), .S(u4_sll_452_n22), .Z(
        u4_sll_452_ML_int_4__29_) );
  MUX2_X2 u4_sll_452_M1_3_30 ( .A(u4_sll_452_ML_int_3__30_), .B(
        u4_sll_452_ML_int_3__22_), .S(u4_sll_452_n19), .Z(
        u4_sll_452_ML_int_4__30_) );
  MUX2_X2 u4_sll_452_M1_3_31 ( .A(u4_sll_452_ML_int_3__31_), .B(
        u4_sll_452_ML_int_3__23_), .S(u4_sll_452_n19), .Z(
        u4_sll_452_ML_int_4__31_) );
  MUX2_X2 u4_sll_452_M1_3_32 ( .A(u4_sll_452_ML_int_3__32_), .B(
        u4_sll_452_ML_int_3__24_), .S(u4_sll_452_n19), .Z(
        u4_sll_452_ML_int_4__32_) );
  MUX2_X2 u4_sll_452_M1_3_33 ( .A(u4_sll_452_ML_int_3__33_), .B(
        u4_sll_452_ML_int_3__25_), .S(u4_sll_452_n19), .Z(
        u4_sll_452_ML_int_4__33_) );
  MUX2_X2 u4_sll_452_M1_3_34 ( .A(u4_sll_452_ML_int_3__34_), .B(
        u4_sll_452_ML_int_3__26_), .S(u4_sll_452_n19), .Z(
        u4_sll_452_ML_int_4__34_) );
  MUX2_X2 u4_sll_452_M1_3_35 ( .A(u4_sll_452_ML_int_3__35_), .B(
        u4_sll_452_ML_int_3__27_), .S(u4_sll_452_n19), .Z(
        u4_sll_452_ML_int_4__35_) );
  MUX2_X2 u4_sll_452_M1_3_36 ( .A(u4_sll_452_ML_int_3__36_), .B(
        u4_sll_452_ML_int_3__28_), .S(u4_sll_452_n21), .Z(
        u4_sll_452_ML_int_4__36_) );
  MUX2_X2 u4_sll_452_M1_3_37 ( .A(u4_sll_452_ML_int_3__37_), .B(
        u4_sll_452_ML_int_3__29_), .S(u4_sll_452_n21), .Z(
        u4_sll_452_ML_int_4__37_) );
  MUX2_X2 u4_sll_452_M1_3_38 ( .A(u4_sll_452_ML_int_3__38_), .B(
        u4_sll_452_ML_int_3__30_), .S(u4_sll_452_n22), .Z(
        u4_sll_452_ML_int_4__38_) );
  MUX2_X2 u4_sll_452_M1_3_39 ( .A(u4_sll_452_ML_int_3__39_), .B(
        u4_sll_452_ML_int_3__31_), .S(u4_sll_452_n19), .Z(
        u4_sll_452_ML_int_4__39_) );
  MUX2_X2 u4_sll_452_M1_3_40 ( .A(u4_sll_452_ML_int_3__40_), .B(
        u4_sll_452_ML_int_3__32_), .S(u4_sll_452_n19), .Z(
        u4_sll_452_ML_int_4__40_) );
  MUX2_X2 u4_sll_452_M1_3_41 ( .A(u4_sll_452_ML_int_3__41_), .B(
        u4_sll_452_ML_int_3__33_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__41_) );
  MUX2_X2 u4_sll_452_M1_3_42 ( .A(u4_sll_452_ML_int_3__42_), .B(
        u4_sll_452_ML_int_3__34_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__42_) );
  MUX2_X2 u4_sll_452_M1_3_43 ( .A(u4_sll_452_ML_int_3__43_), .B(
        u4_sll_452_ML_int_3__35_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__43_) );
  MUX2_X2 u4_sll_452_M1_3_44 ( .A(u4_sll_452_ML_int_3__44_), .B(
        u4_sll_452_ML_int_3__36_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__44_) );
  MUX2_X2 u4_sll_452_M1_3_45 ( .A(u4_sll_452_ML_int_3__45_), .B(
        u4_sll_452_ML_int_3__37_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__45_) );
  MUX2_X2 u4_sll_452_M1_3_46 ( .A(u4_sll_452_ML_int_3__46_), .B(
        u4_sll_452_ML_int_3__38_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__46_) );
  MUX2_X2 u4_sll_452_M1_3_47 ( .A(u4_sll_452_ML_int_3__47_), .B(
        u4_sll_452_ML_int_3__39_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__47_) );
  MUX2_X2 u4_sll_452_M1_3_48 ( .A(u4_sll_452_ML_int_3__48_), .B(
        u4_sll_452_ML_int_3__40_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__48_) );
  MUX2_X2 u4_sll_452_M1_3_49 ( .A(u4_sll_452_ML_int_3__49_), .B(
        u4_sll_452_ML_int_3__41_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__49_) );
  MUX2_X2 u4_sll_452_M1_3_50 ( .A(u4_sll_452_ML_int_3__50_), .B(
        u4_sll_452_ML_int_3__42_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__50_) );
  MUX2_X2 u4_sll_452_M1_3_51 ( .A(u4_sll_452_ML_int_3__51_), .B(
        u4_sll_452_ML_int_3__43_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__51_) );
  MUX2_X2 u4_sll_452_M1_3_52 ( .A(u4_sll_452_ML_int_3__52_), .B(
        u4_sll_452_ML_int_3__44_), .S(u4_sll_452_n21), .Z(
        u4_sll_452_ML_int_4__52_) );
  MUX2_X2 u4_sll_452_M1_3_53 ( .A(u4_sll_452_ML_int_3__53_), .B(
        u4_sll_452_ML_int_3__45_), .S(u4_sll_452_n21), .Z(
        u4_sll_452_ML_int_4__53_) );
  MUX2_X2 u4_sll_452_M1_3_54 ( .A(u4_sll_452_ML_int_3__54_), .B(
        u4_sll_452_ML_int_3__46_), .S(u4_sll_452_n21), .Z(
        u4_sll_452_ML_int_4__54_) );
  MUX2_X2 u4_sll_452_M1_3_55 ( .A(u4_sll_452_ML_int_3__55_), .B(
        u4_sll_452_ML_int_3__47_), .S(u4_sll_452_n21), .Z(
        u4_sll_452_ML_int_4__55_) );
  MUX2_X2 u4_sll_452_M1_3_56 ( .A(u4_sll_452_ML_int_3__56_), .B(
        u4_sll_452_ML_int_3__48_), .S(u4_sll_452_n21), .Z(
        u4_sll_452_ML_int_4__56_) );
  MUX2_X2 u4_sll_452_M1_3_57 ( .A(u4_sll_452_ML_int_3__57_), .B(
        u4_sll_452_ML_int_3__49_), .S(u4_sll_452_n21), .Z(
        u4_sll_452_ML_int_4__57_) );
  MUX2_X2 u4_sll_452_M1_3_58 ( .A(u4_sll_452_ML_int_3__58_), .B(
        u4_sll_452_ML_int_3__50_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__58_) );
  MUX2_X2 u4_sll_452_M1_3_59 ( .A(u4_sll_452_ML_int_3__59_), .B(
        u4_sll_452_ML_int_3__51_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__59_) );
  MUX2_X2 u4_sll_452_M1_3_60 ( .A(u4_sll_452_ML_int_3__60_), .B(
        u4_sll_452_ML_int_3__52_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__60_) );
  MUX2_X2 u4_sll_452_M1_3_61 ( .A(u4_sll_452_ML_int_3__61_), .B(
        u4_sll_452_ML_int_3__53_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__61_) );
  MUX2_X2 u4_sll_452_M1_3_62 ( .A(u4_sll_452_ML_int_3__62_), .B(
        u4_sll_452_ML_int_3__54_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__62_) );
  MUX2_X2 u4_sll_452_M1_3_63 ( .A(u4_sll_452_ML_int_3__63_), .B(
        u4_sll_452_ML_int_3__55_), .S(u4_sll_452_n21), .Z(
        u4_sll_452_ML_int_4__63_) );
  MUX2_X2 u4_sll_452_M1_3_64 ( .A(u4_sll_452_ML_int_3__64_), .B(
        u4_sll_452_ML_int_3__56_), .S(u4_sll_452_n21), .Z(
        u4_sll_452_ML_int_4__64_) );
  MUX2_X2 u4_sll_452_M1_3_65 ( .A(u4_sll_452_ML_int_3__65_), .B(
        u4_sll_452_ML_int_3__57_), .S(u4_sll_452_n21), .Z(
        u4_sll_452_ML_int_4__65_) );
  MUX2_X2 u4_sll_452_M1_3_66 ( .A(u4_sll_452_ML_int_3__66_), .B(
        u4_sll_452_ML_int_3__58_), .S(u4_sll_452_n21), .Z(
        u4_sll_452_ML_int_4__66_) );
  MUX2_X2 u4_sll_452_M1_3_67 ( .A(u4_sll_452_ML_int_3__67_), .B(
        u4_sll_452_ML_int_3__59_), .S(u4_sll_452_n21), .Z(
        u4_sll_452_ML_int_4__67_) );
  MUX2_X2 u4_sll_452_M1_3_68 ( .A(u4_sll_452_ML_int_3__68_), .B(
        u4_sll_452_ML_int_3__60_), .S(u4_sll_452_n21), .Z(
        u4_sll_452_ML_int_4__68_) );
  MUX2_X2 u4_sll_452_M1_3_69 ( .A(u4_sll_452_ML_int_3__69_), .B(
        u4_sll_452_ML_int_3__61_), .S(u4_sll_452_n21), .Z(
        u4_sll_452_ML_int_4__69_) );
  MUX2_X2 u4_sll_452_M1_3_70 ( .A(u4_sll_452_ML_int_3__70_), .B(
        u4_sll_452_ML_int_3__62_), .S(u4_sll_452_n21), .Z(
        u4_sll_452_ML_int_4__70_) );
  MUX2_X2 u4_sll_452_M1_3_71 ( .A(u4_sll_452_ML_int_3__71_), .B(
        u4_sll_452_ML_int_3__63_), .S(u4_sll_452_n21), .Z(
        u4_sll_452_ML_int_4__71_) );
  MUX2_X2 u4_sll_452_M1_3_72 ( .A(u4_sll_452_ML_int_3__72_), .B(
        u4_sll_452_ML_int_3__64_), .S(u4_sll_452_n21), .Z(
        u4_sll_452_ML_int_4__72_) );
  MUX2_X2 u4_sll_452_M1_3_73 ( .A(u4_sll_452_ML_int_3__73_), .B(
        u4_sll_452_ML_int_3__65_), .S(u4_sll_452_n21), .Z(
        u4_sll_452_ML_int_4__73_) );
  MUX2_X2 u4_sll_452_M1_3_74 ( .A(u4_sll_452_ML_int_3__74_), .B(
        u4_sll_452_ML_int_3__66_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__74_) );
  MUX2_X2 u4_sll_452_M1_3_75 ( .A(u4_sll_452_ML_int_3__75_), .B(
        u4_sll_452_ML_int_3__67_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__75_) );
  MUX2_X2 u4_sll_452_M1_3_76 ( .A(u4_sll_452_ML_int_3__76_), .B(
        u4_sll_452_ML_int_3__68_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__76_) );
  MUX2_X2 u4_sll_452_M1_3_77 ( .A(u4_sll_452_ML_int_3__77_), .B(
        u4_sll_452_ML_int_3__69_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__77_) );
  MUX2_X2 u4_sll_452_M1_3_78 ( .A(u4_sll_452_ML_int_3__78_), .B(
        u4_sll_452_ML_int_3__70_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__78_) );
  MUX2_X2 u4_sll_452_M1_3_79 ( .A(u4_sll_452_ML_int_3__79_), .B(
        u4_sll_452_ML_int_3__71_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__79_) );
  MUX2_X2 u4_sll_452_M1_3_80 ( .A(u4_sll_452_ML_int_3__80_), .B(
        u4_sll_452_ML_int_3__72_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__80_) );
  MUX2_X2 u4_sll_452_M1_3_81 ( .A(u4_sll_452_ML_int_3__81_), .B(
        u4_sll_452_ML_int_3__73_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__81_) );
  MUX2_X2 u4_sll_452_M1_3_82 ( .A(u4_sll_452_ML_int_3__82_), .B(
        u4_sll_452_ML_int_3__74_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__82_) );
  MUX2_X2 u4_sll_452_M1_3_83 ( .A(u4_sll_452_ML_int_3__83_), .B(
        u4_sll_452_ML_int_3__75_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__83_) );
  MUX2_X2 u4_sll_452_M1_3_84 ( .A(u4_sll_452_ML_int_3__84_), .B(
        u4_sll_452_ML_int_3__76_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__84_) );
  MUX2_X2 u4_sll_452_M1_3_85 ( .A(u4_sll_452_ML_int_3__85_), .B(
        u4_sll_452_ML_int_3__77_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__85_) );
  MUX2_X2 u4_sll_452_M1_3_86 ( .A(u4_sll_452_ML_int_3__86_), .B(
        u4_sll_452_ML_int_3__78_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__86_) );
  MUX2_X2 u4_sll_452_M1_3_87 ( .A(u4_sll_452_ML_int_3__87_), .B(
        u4_sll_452_ML_int_3__79_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__87_) );
  MUX2_X2 u4_sll_452_M1_3_88 ( .A(u4_sll_452_ML_int_3__88_), .B(
        u4_sll_452_ML_int_3__80_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__88_) );
  MUX2_X2 u4_sll_452_M1_3_89 ( .A(u4_sll_452_ML_int_3__89_), .B(
        u4_sll_452_ML_int_3__81_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__89_) );
  MUX2_X2 u4_sll_452_M1_3_90 ( .A(u4_sll_452_ML_int_3__90_), .B(
        u4_sll_452_ML_int_3__82_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__90_) );
  MUX2_X2 u4_sll_452_M1_3_91 ( .A(u4_sll_452_ML_int_3__91_), .B(
        u4_sll_452_ML_int_3__83_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__91_) );
  MUX2_X2 u4_sll_452_M1_3_92 ( .A(u4_sll_452_ML_int_3__92_), .B(
        u4_sll_452_ML_int_3__84_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__92_) );
  MUX2_X2 u4_sll_452_M1_3_93 ( .A(u4_sll_452_ML_int_3__93_), .B(
        u4_sll_452_ML_int_3__85_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__93_) );
  MUX2_X2 u4_sll_452_M1_3_94 ( .A(u4_sll_452_ML_int_3__94_), .B(
        u4_sll_452_ML_int_3__86_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__94_) );
  MUX2_X2 u4_sll_452_M1_3_95 ( .A(u4_sll_452_ML_int_3__95_), .B(
        u4_sll_452_ML_int_3__87_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__95_) );
  MUX2_X2 u4_sll_452_M1_3_96 ( .A(u4_sll_452_ML_int_3__96_), .B(
        u4_sll_452_ML_int_3__88_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__96_) );
  MUX2_X2 u4_sll_452_M1_3_97 ( .A(u4_sll_452_ML_int_3__97_), .B(
        u4_sll_452_ML_int_3__89_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__97_) );
  MUX2_X2 u4_sll_452_M1_3_98 ( .A(u4_sll_452_ML_int_3__98_), .B(
        u4_sll_452_ML_int_3__90_), .S(u4_sll_452_n19), .Z(
        u4_sll_452_ML_int_4__98_) );
  MUX2_X2 u4_sll_452_M1_3_99 ( .A(u4_sll_452_ML_int_3__99_), .B(
        u4_sll_452_ML_int_3__91_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__99_) );
  MUX2_X2 u4_sll_452_M1_3_100 ( .A(u4_sll_452_ML_int_3__100_), .B(
        u4_sll_452_ML_int_3__92_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__100_) );
  MUX2_X2 u4_sll_452_M1_3_101 ( .A(u4_sll_452_ML_int_3__101_), .B(
        u4_sll_452_ML_int_3__93_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__101_) );
  MUX2_X2 u4_sll_452_M1_3_102 ( .A(u4_sll_452_ML_int_3__102_), .B(
        u4_sll_452_ML_int_3__94_), .S(u4_sll_452_n19), .Z(
        u4_sll_452_ML_int_4__102_) );
  MUX2_X2 u4_sll_452_M1_3_103 ( .A(u4_sll_452_ML_int_3__103_), .B(
        u4_sll_452_ML_int_3__95_), .S(u4_sll_452_n19), .Z(
        u4_sll_452_ML_int_4__103_) );
  MUX2_X2 u4_sll_452_M1_3_104 ( .A(u4_sll_452_ML_int_3__104_), .B(
        u4_sll_452_ML_int_3__96_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__104_) );
  MUX2_X2 u4_sll_452_M1_3_105 ( .A(u4_sll_452_ML_int_3__105_), .B(
        u4_sll_452_ML_int_3__97_), .S(u4_sll_452_n20), .Z(
        u4_sll_452_ML_int_4__105_) );
  MUX2_X2 u4_sll_452_M1_4_16 ( .A(u4_sll_452_ML_int_4__16_), .B(
        u4_sll_452_ML_int_4__0_), .S(u4_sll_452_n34), .Z(
        u4_sll_452_ML_int_5__16_) );
  MUX2_X2 u4_sll_452_M1_4_17 ( .A(u4_sll_452_ML_int_4__17_), .B(
        u4_sll_452_ML_int_4__1_), .S(u4_sll_452_n34), .Z(
        u4_sll_452_ML_int_5__17_) );
  MUX2_X2 u4_sll_452_M1_4_18 ( .A(u4_sll_452_ML_int_4__18_), .B(
        u4_sll_452_ML_int_4__2_), .S(u4_sll_452_n33), .Z(
        u4_sll_452_ML_int_5__18_) );
  MUX2_X2 u4_sll_452_M1_4_19 ( .A(u4_sll_452_ML_int_4__19_), .B(
        u4_sll_452_ML_int_4__3_), .S(u4_sll_452_n33), .Z(
        u4_sll_452_ML_int_5__19_) );
  MUX2_X2 u4_sll_452_M1_4_20 ( .A(u4_sll_452_ML_int_4__20_), .B(
        u4_sll_452_ML_int_4__4_), .S(u4_sll_452_n33), .Z(
        u4_sll_452_ML_int_5__20_) );
  MUX2_X2 u4_sll_452_M1_4_21 ( .A(u4_sll_452_ML_int_4__21_), .B(
        u4_sll_452_ML_int_4__5_), .S(u4_sll_452_n33), .Z(
        u4_sll_452_ML_int_5__21_) );
  MUX2_X2 u4_sll_452_M1_4_22 ( .A(u4_sll_452_ML_int_4__22_), .B(
        u4_sll_452_ML_int_4__6_), .S(u4_sll_452_n33), .Z(
        u4_sll_452_ML_int_5__22_) );
  MUX2_X2 u4_sll_452_M1_4_23 ( .A(u4_sll_452_ML_int_4__23_), .B(
        u4_sll_452_ML_int_4__7_), .S(u4_sll_452_n33), .Z(
        u4_sll_452_ML_int_5__23_) );
  MUX2_X2 u4_sll_452_M1_4_24 ( .A(u4_sll_452_ML_int_4__24_), .B(
        u4_sll_452_ML_int_4__8_), .S(u4_sll_452_n33), .Z(
        u4_sll_452_ML_int_5__24_) );
  MUX2_X2 u4_sll_452_M1_4_25 ( .A(u4_sll_452_ML_int_4__25_), .B(
        u4_sll_452_ML_int_4__9_), .S(u4_sll_452_n33), .Z(
        u4_sll_452_ML_int_5__25_) );
  MUX2_X2 u4_sll_452_M1_4_26 ( .A(u4_sll_452_ML_int_4__26_), .B(
        u4_sll_452_ML_int_4__10_), .S(u4_sll_452_n33), .Z(
        u4_sll_452_ML_int_5__26_) );
  MUX2_X2 u4_sll_452_M1_4_27 ( .A(u4_sll_452_ML_int_4__27_), .B(
        u4_sll_452_ML_int_4__11_), .S(u4_sll_452_n34), .Z(
        u4_sll_452_ML_int_5__27_) );
  MUX2_X2 u4_sll_452_M1_4_28 ( .A(u4_sll_452_ML_int_4__28_), .B(
        u4_sll_452_ML_int_4__12_), .S(u4_sll_452_n34), .Z(
        u4_sll_452_ML_int_5__28_) );
  MUX2_X2 u4_sll_452_M1_4_29 ( .A(u4_sll_452_ML_int_4__29_), .B(
        u4_sll_452_ML_int_4__13_), .S(u4_sll_452_n34), .Z(
        u4_sll_452_ML_int_5__29_) );
  MUX2_X2 u4_sll_452_M1_4_30 ( .A(u4_sll_452_ML_int_4__30_), .B(
        u4_sll_452_ML_int_4__14_), .S(u4_sll_452_n34), .Z(
        u4_sll_452_ML_int_5__30_) );
  MUX2_X2 u4_sll_452_M1_4_31 ( .A(u4_sll_452_ML_int_4__31_), .B(
        u4_sll_452_ML_int_4__15_), .S(u4_sll_452_n34), .Z(
        u4_sll_452_ML_int_5__31_) );
  MUX2_X2 u4_sll_452_M1_4_32 ( .A(u4_sll_452_ML_int_4__32_), .B(
        u4_sll_452_ML_int_4__16_), .S(u4_sll_452_n34), .Z(
        u4_sll_452_ML_int_5__32_) );
  MUX2_X2 u4_sll_452_M1_4_33 ( .A(u4_sll_452_ML_int_4__33_), .B(
        u4_sll_452_ML_int_4__17_), .S(u4_sll_452_n34), .Z(
        u4_sll_452_ML_int_5__33_) );
  MUX2_X2 u4_sll_452_M1_4_34 ( .A(u4_sll_452_ML_int_4__34_), .B(
        u4_sll_452_ML_int_4__18_), .S(u4_sll_452_n34), .Z(
        u4_sll_452_ML_int_5__34_) );
  MUX2_X2 u4_sll_452_M1_4_35 ( .A(u4_sll_452_ML_int_4__35_), .B(
        u4_sll_452_ML_int_4__19_), .S(u4_sll_452_n34), .Z(
        u4_sll_452_ML_int_5__35_) );
  MUX2_X2 u4_sll_452_M1_4_36 ( .A(u4_sll_452_ML_int_4__36_), .B(
        u4_sll_452_ML_int_4__20_), .S(u4_sll_452_n34), .Z(
        u4_sll_452_ML_int_5__36_) );
  MUX2_X2 u4_sll_452_M1_4_37 ( .A(u4_sll_452_ML_int_4__37_), .B(
        u4_sll_452_ML_int_4__21_), .S(u4_sll_452_n34), .Z(
        u4_sll_452_ML_int_5__37_) );
  MUX2_X2 u4_sll_452_M1_4_38 ( .A(u4_sll_452_ML_int_4__38_), .B(
        u4_sll_452_ML_int_4__22_), .S(u4_sll_452_n30), .Z(
        u4_sll_452_ML_int_5__38_) );
  MUX2_X2 u4_sll_452_M1_4_39 ( .A(u4_sll_452_ML_int_4__39_), .B(
        u4_sll_452_ML_int_4__23_), .S(u4_sll_452_n30), .Z(
        u4_sll_452_ML_int_5__39_) );
  MUX2_X2 u4_sll_452_M1_4_40 ( .A(u4_sll_452_ML_int_4__40_), .B(
        u4_sll_452_ML_int_4__24_), .S(u4_sll_452_n30), .Z(
        u4_sll_452_ML_int_5__40_) );
  MUX2_X2 u4_sll_452_M1_4_41 ( .A(u4_sll_452_ML_int_4__41_), .B(
        u4_sll_452_ML_int_4__25_), .S(u4_sll_452_n30), .Z(
        u4_sll_452_ML_int_5__41_) );
  MUX2_X2 u4_sll_452_M1_4_42 ( .A(u4_sll_452_ML_int_4__42_), .B(
        u4_sll_452_ML_int_4__26_), .S(u4_sll_452_n30), .Z(
        u4_sll_452_ML_int_5__42_) );
  MUX2_X2 u4_sll_452_M1_4_43 ( .A(u4_sll_452_ML_int_4__43_), .B(
        u4_sll_452_ML_int_4__27_), .S(u4_sll_452_n30), .Z(
        u4_sll_452_ML_int_5__43_) );
  MUX2_X2 u4_sll_452_M1_4_44 ( .A(u4_sll_452_ML_int_4__44_), .B(
        u4_sll_452_ML_int_4__28_), .S(u4_sll_452_n34), .Z(
        u4_sll_452_ML_int_5__44_) );
  MUX2_X2 u4_sll_452_M1_4_45 ( .A(u4_sll_452_ML_int_4__45_), .B(
        u4_sll_452_ML_int_4__29_), .S(u4_sll_452_n34), .Z(
        u4_sll_452_ML_int_5__45_) );
  MUX2_X2 u4_sll_452_M1_4_46 ( .A(u4_sll_452_ML_int_4__46_), .B(
        u4_sll_452_ML_int_4__30_), .S(u4_sll_452_n34), .Z(
        u4_sll_452_ML_int_5__46_) );
  MUX2_X2 u4_sll_452_M1_4_47 ( .A(u4_sll_452_ML_int_4__47_), .B(
        u4_sll_452_ML_int_4__31_), .S(u4_sll_452_n34), .Z(
        u4_sll_452_ML_int_5__47_) );
  MUX2_X2 u4_sll_452_M1_4_48 ( .A(u4_sll_452_ML_int_4__48_), .B(
        u4_sll_452_ML_int_4__32_), .S(u4_sll_452_n34), .Z(
        u4_sll_452_ML_int_5__48_) );
  MUX2_X2 u4_sll_452_M1_4_49 ( .A(u4_sll_452_ML_int_4__49_), .B(
        u4_sll_452_ML_int_4__33_), .S(u4_sll_452_n32), .Z(
        u4_sll_452_ML_int_5__49_) );
  MUX2_X2 u4_sll_452_M1_4_50 ( .A(u4_sll_452_ML_int_4__50_), .B(
        u4_sll_452_ML_int_4__34_), .S(u4_sll_452_n32), .Z(
        u4_sll_452_ML_int_5__50_) );
  MUX2_X2 u4_sll_452_M1_4_51 ( .A(u4_sll_452_ML_int_4__51_), .B(
        u4_sll_452_ML_int_4__35_), .S(u4_sll_452_n32), .Z(
        u4_sll_452_ML_int_5__51_) );
  MUX2_X2 u4_sll_452_M1_4_52 ( .A(u4_sll_452_ML_int_4__52_), .B(
        u4_sll_452_ML_int_4__36_), .S(u4_sll_452_n32), .Z(
        u4_sll_452_ML_int_5__52_) );
  MUX2_X2 u4_sll_452_M1_4_53 ( .A(u4_sll_452_ML_int_4__53_), .B(
        u4_sll_452_ML_int_4__37_), .S(u4_sll_452_n32), .Z(
        u4_sll_452_ML_int_5__53_) );
  MUX2_X2 u4_sll_452_M1_4_54 ( .A(u4_sll_452_ML_int_4__54_), .B(
        u4_sll_452_ML_int_4__38_), .S(u4_sll_452_n31), .Z(
        u4_sll_452_ML_int_5__54_) );
  MUX2_X2 u4_sll_452_M1_4_55 ( .A(u4_sll_452_ML_int_4__55_), .B(
        u4_sll_452_ML_int_4__39_), .S(u4_sll_452_n31), .Z(
        u4_sll_452_ML_int_5__55_) );
  MUX2_X2 u4_sll_452_M1_4_56 ( .A(u4_sll_452_ML_int_4__56_), .B(
        u4_sll_452_ML_int_4__40_), .S(u4_sll_452_n31), .Z(
        u4_sll_452_ML_int_5__56_) );
  MUX2_X2 u4_sll_452_M1_4_57 ( .A(u4_sll_452_ML_int_4__57_), .B(
        u4_sll_452_ML_int_4__41_), .S(u4_sll_452_n31), .Z(
        u4_sll_452_ML_int_5__57_) );
  MUX2_X2 u4_sll_452_M1_4_58 ( .A(u4_sll_452_ML_int_4__58_), .B(
        u4_sll_452_ML_int_4__42_), .S(u4_sll_452_n31), .Z(
        u4_sll_452_ML_int_5__58_) );
  MUX2_X2 u4_sll_452_M1_4_59 ( .A(u4_sll_452_ML_int_4__59_), .B(
        u4_sll_452_ML_int_4__43_), .S(u4_sll_452_n31), .Z(
        u4_sll_452_ML_int_5__59_) );
  MUX2_X2 u4_sll_452_M1_4_60 ( .A(u4_sll_452_ML_int_4__60_), .B(
        u4_sll_452_ML_int_4__44_), .S(u4_sll_452_n32), .Z(
        u4_sll_452_ML_int_5__60_) );
  MUX2_X2 u4_sll_452_M1_4_61 ( .A(u4_sll_452_ML_int_4__61_), .B(
        u4_sll_452_ML_int_4__45_), .S(u4_sll_452_n32), .Z(
        u4_sll_452_ML_int_5__61_) );
  MUX2_X2 u4_sll_452_M1_4_62 ( .A(u4_sll_452_ML_int_4__62_), .B(
        u4_sll_452_ML_int_4__46_), .S(u4_sll_452_n32), .Z(
        u4_sll_452_ML_int_5__62_) );
  MUX2_X2 u4_sll_452_M1_4_63 ( .A(u4_sll_452_ML_int_4__63_), .B(
        u4_sll_452_ML_int_4__47_), .S(u4_sll_452_n32), .Z(
        u4_sll_452_ML_int_5__63_) );
  MUX2_X2 u4_sll_452_M1_4_64 ( .A(u4_sll_452_ML_int_4__64_), .B(
        u4_sll_452_ML_int_4__48_), .S(u4_sll_452_n32), .Z(
        u4_sll_452_ML_int_5__64_) );
  MUX2_X2 u4_sll_452_M1_4_65 ( .A(u4_sll_452_ML_int_4__65_), .B(
        u4_sll_452_ML_int_4__49_), .S(u4_sll_452_n32), .Z(
        u4_sll_452_ML_int_5__65_) );
  MUX2_X2 u4_sll_452_M1_4_66 ( .A(u4_sll_452_ML_int_4__66_), .B(
        u4_sll_452_ML_int_4__50_), .S(u4_sll_452_n32), .Z(
        u4_sll_452_ML_int_5__66_) );
  MUX2_X2 u4_sll_452_M1_4_67 ( .A(u4_sll_452_ML_int_4__67_), .B(
        u4_sll_452_ML_int_4__51_), .S(u4_sll_452_n32), .Z(
        u4_sll_452_ML_int_5__67_) );
  MUX2_X2 u4_sll_452_M1_4_68 ( .A(u4_sll_452_ML_int_4__68_), .B(
        u4_sll_452_ML_int_4__52_), .S(u4_sll_452_n32), .Z(
        u4_sll_452_ML_int_5__68_) );
  MUX2_X2 u4_sll_452_M1_4_69 ( .A(u4_sll_452_ML_int_4__69_), .B(
        u4_sll_452_ML_int_4__53_), .S(u4_sll_452_n32), .Z(
        u4_sll_452_ML_int_5__69_) );
  MUX2_X2 u4_sll_452_M1_4_70 ( .A(u4_sll_452_ML_int_4__70_), .B(
        u4_sll_452_ML_int_4__54_), .S(u4_sll_452_n32), .Z(
        u4_sll_452_ML_int_5__70_) );
  MUX2_X2 u4_sll_452_M1_4_71 ( .A(u4_sll_452_ML_int_4__71_), .B(
        u4_sll_452_ML_int_4__55_), .S(u4_sll_452_n33), .Z(
        u4_sll_452_ML_int_5__71_) );
  MUX2_X2 u4_sll_452_M1_4_72 ( .A(u4_sll_452_ML_int_4__72_), .B(
        u4_sll_452_ML_int_4__56_), .S(u4_sll_452_n33), .Z(
        u4_sll_452_ML_int_5__72_) );
  MUX2_X2 u4_sll_452_M1_4_73 ( .A(u4_sll_452_ML_int_4__73_), .B(
        u4_sll_452_ML_int_4__57_), .S(u4_sll_452_n33), .Z(
        u4_sll_452_ML_int_5__73_) );
  MUX2_X2 u4_sll_452_M1_4_74 ( .A(u4_sll_452_ML_int_4__74_), .B(
        u4_sll_452_ML_int_4__58_), .S(u4_sll_452_n33), .Z(
        u4_sll_452_ML_int_5__74_) );
  MUX2_X2 u4_sll_452_M1_4_75 ( .A(u4_sll_452_ML_int_4__75_), .B(
        u4_sll_452_ML_int_4__59_), .S(u4_sll_452_n33), .Z(
        u4_sll_452_ML_int_5__75_) );
  MUX2_X2 u4_sll_452_M1_4_76 ( .A(u4_sll_452_ML_int_4__76_), .B(
        u4_sll_452_ML_int_4__60_), .S(u4_sll_452_n33), .Z(
        u4_sll_452_ML_int_5__76_) );
  MUX2_X2 u4_sll_452_M1_4_77 ( .A(u4_sll_452_ML_int_4__77_), .B(
        u4_sll_452_ML_int_4__61_), .S(u4_sll_452_n33), .Z(
        u4_sll_452_ML_int_5__77_) );
  MUX2_X2 u4_sll_452_M1_4_78 ( .A(u4_sll_452_ML_int_4__78_), .B(
        u4_sll_452_ML_int_4__62_), .S(u4_sll_452_n33), .Z(
        u4_sll_452_ML_int_5__78_) );
  MUX2_X2 u4_sll_452_M1_4_79 ( .A(u4_sll_452_ML_int_4__79_), .B(
        u4_sll_452_ML_int_4__63_), .S(u4_sll_452_n33), .Z(
        u4_sll_452_ML_int_5__79_) );
  MUX2_X2 u4_sll_452_M1_4_80 ( .A(u4_sll_452_ML_int_4__80_), .B(
        u4_sll_452_ML_int_4__64_), .S(u4_sll_452_n32), .Z(
        u4_sll_452_ML_int_5__80_) );
  MUX2_X2 u4_sll_452_M1_4_81 ( .A(u4_sll_452_ML_int_4__81_), .B(
        u4_sll_452_ML_int_4__65_), .S(u4_sll_452_n32), .Z(
        u4_sll_452_ML_int_5__81_) );
  MUX2_X2 u4_sll_452_M1_4_82 ( .A(u4_sll_452_ML_int_4__82_), .B(
        u4_sll_452_ML_int_4__66_), .S(u4_sll_452_n30), .Z(
        u4_sll_452_ML_int_5__82_) );
  MUX2_X2 u4_sll_452_M1_4_83 ( .A(u4_sll_452_ML_int_4__83_), .B(
        u4_sll_452_ML_int_4__67_), .S(u4_sll_452_n30), .Z(
        u4_sll_452_ML_int_5__83_) );
  MUX2_X2 u4_sll_452_M1_4_84 ( .A(u4_sll_452_ML_int_4__84_), .B(
        u4_sll_452_ML_int_4__68_), .S(u4_sll_452_n30), .Z(
        u4_sll_452_ML_int_5__84_) );
  MUX2_X2 u4_sll_452_M1_4_85 ( .A(u4_sll_452_ML_int_4__85_), .B(
        u4_sll_452_ML_int_4__69_), .S(u4_sll_452_n30), .Z(
        u4_sll_452_ML_int_5__85_) );
  MUX2_X2 u4_sll_452_M1_4_86 ( .A(u4_sll_452_ML_int_4__86_), .B(
        u4_sll_452_ML_int_4__70_), .S(u4_sll_452_n30), .Z(
        u4_sll_452_ML_int_5__86_) );
  MUX2_X2 u4_sll_452_M1_4_87 ( .A(u4_sll_452_ML_int_4__87_), .B(
        u4_sll_452_ML_int_4__71_), .S(u4_sll_452_n30), .Z(
        u4_sll_452_ML_int_5__87_) );
  MUX2_X2 u4_sll_452_M1_4_88 ( .A(u4_sll_452_ML_int_4__88_), .B(
        u4_sll_452_ML_int_4__72_), .S(u4_sll_452_n30), .Z(
        u4_sll_452_ML_int_5__88_) );
  MUX2_X2 u4_sll_452_M1_4_89 ( .A(u4_sll_452_ML_int_4__89_), .B(
        u4_sll_452_ML_int_4__73_), .S(u4_sll_452_n30), .Z(
        u4_sll_452_ML_int_5__89_) );
  MUX2_X2 u4_sll_452_M1_4_90 ( .A(u4_sll_452_ML_int_4__90_), .B(
        u4_sll_452_ML_int_4__74_), .S(u4_sll_452_n30), .Z(
        u4_sll_452_ML_int_5__90_) );
  MUX2_X2 u4_sll_452_M1_4_91 ( .A(u4_sll_452_ML_int_4__91_), .B(
        u4_sll_452_ML_int_4__75_), .S(u4_sll_452_n30), .Z(
        u4_sll_452_ML_int_5__91_) );
  MUX2_X2 u4_sll_452_M1_4_92 ( .A(u4_sll_452_ML_int_4__92_), .B(
        u4_sll_452_ML_int_4__76_), .S(u4_sll_452_n30), .Z(
        u4_sll_452_ML_int_5__92_) );
  MUX2_X2 u4_sll_452_M1_4_93 ( .A(u4_sll_452_ML_int_4__93_), .B(
        u4_sll_452_ML_int_4__77_), .S(u4_sll_452_n31), .Z(
        u4_sll_452_ML_int_5__93_) );
  MUX2_X2 u4_sll_452_M1_4_94 ( .A(u4_sll_452_ML_int_4__94_), .B(
        u4_sll_452_ML_int_4__78_), .S(u4_sll_452_n31), .Z(
        u4_sll_452_ML_int_5__94_) );
  MUX2_X2 u4_sll_452_M1_4_95 ( .A(u4_sll_452_ML_int_4__95_), .B(
        u4_sll_452_ML_int_4__79_), .S(u4_sll_452_n31), .Z(
        u4_sll_452_ML_int_5__95_) );
  MUX2_X2 u4_sll_452_M1_4_96 ( .A(u4_sll_452_ML_int_4__96_), .B(
        u4_sll_452_ML_int_4__80_), .S(u4_sll_452_n31), .Z(
        u4_sll_452_ML_int_5__96_) );
  MUX2_X2 u4_sll_452_M1_4_97 ( .A(u4_sll_452_ML_int_4__97_), .B(
        u4_sll_452_ML_int_4__81_), .S(u4_sll_452_n31), .Z(
        u4_sll_452_ML_int_5__97_) );
  MUX2_X2 u4_sll_452_M1_4_98 ( .A(u4_sll_452_ML_int_4__98_), .B(
        u4_sll_452_ML_int_4__82_), .S(u4_sll_452_n31), .Z(
        u4_sll_452_ML_int_5__98_) );
  MUX2_X2 u4_sll_452_M1_4_99 ( .A(u4_sll_452_ML_int_4__99_), .B(
        u4_sll_452_ML_int_4__83_), .S(u4_sll_452_n31), .Z(
        u4_sll_452_ML_int_5__99_) );
  MUX2_X2 u4_sll_452_M1_4_100 ( .A(u4_sll_452_ML_int_4__100_), .B(
        u4_sll_452_ML_int_4__84_), .S(u4_sll_452_n31), .Z(
        u4_sll_452_ML_int_5__100_) );
  MUX2_X2 u4_sll_452_M1_4_101 ( .A(u4_sll_452_ML_int_4__101_), .B(
        u4_sll_452_ML_int_4__85_), .S(u4_sll_452_n31), .Z(
        u4_sll_452_ML_int_5__101_) );
  MUX2_X2 u4_sll_452_M1_4_102 ( .A(u4_sll_452_ML_int_4__102_), .B(
        u4_sll_452_ML_int_4__86_), .S(u4_sll_452_n31), .Z(
        u4_sll_452_ML_int_5__102_) );
  MUX2_X2 u4_sll_452_M1_4_103 ( .A(u4_sll_452_ML_int_4__103_), .B(
        u4_sll_452_ML_int_4__87_), .S(u4_sll_452_n30), .Z(
        u4_sll_452_ML_int_5__103_) );
  MUX2_X2 u4_sll_452_M1_4_104 ( .A(u4_sll_452_ML_int_4__104_), .B(
        u4_sll_452_ML_int_4__88_), .S(u4_sll_452_n31), .Z(
        u4_sll_452_ML_int_5__104_) );
  MUX2_X2 u4_sll_452_M1_4_105 ( .A(u4_sll_452_ML_int_4__105_), .B(
        u4_sll_452_ML_int_4__89_), .S(u4_sll_452_n31), .Z(
        u4_sll_452_ML_int_5__105_) );
  MUX2_X2 u4_sll_452_M1_5_32 ( .A(u4_sll_452_ML_int_5__32_), .B(
        u4_sll_452_ML_int_5__0_), .S(u4_sll_452_n46), .Z(
        u4_sll_452_ML_int_6__32_) );
  MUX2_X2 u4_sll_452_M1_5_33 ( .A(u4_sll_452_ML_int_5__33_), .B(
        u4_sll_452_ML_int_5__1_), .S(u4_sll_452_n46), .Z(
        u4_sll_452_ML_int_6__33_) );
  MUX2_X2 u4_sll_452_M1_5_34 ( .A(u4_sll_452_ML_int_5__34_), .B(
        u4_sll_452_ML_int_5__2_), .S(u4_sll_452_n46), .Z(
        u4_sll_452_ML_int_6__34_) );
  MUX2_X2 u4_sll_452_M1_5_35 ( .A(u4_sll_452_ML_int_5__35_), .B(
        u4_sll_452_ML_int_5__3_), .S(u4_sll_452_n46), .Z(
        u4_sll_452_ML_int_6__35_) );
  MUX2_X2 u4_sll_452_M1_5_36 ( .A(u4_sll_452_ML_int_5__36_), .B(
        u4_sll_452_ML_int_5__4_), .S(u4_sll_452_n46), .Z(
        u4_sll_452_ML_int_6__36_) );
  MUX2_X2 u4_sll_452_M1_5_37 ( .A(u4_sll_452_ML_int_5__37_), .B(
        u4_sll_452_ML_int_5__5_), .S(u4_sll_452_n46), .Z(
        u4_sll_452_ML_int_6__37_) );
  MUX2_X2 u4_sll_452_M1_5_38 ( .A(u4_sll_452_ML_int_5__38_), .B(
        u4_sll_452_ML_int_5__6_), .S(u4_sll_452_n47), .Z(
        u4_sll_452_ML_int_6__38_) );
  MUX2_X2 u4_sll_452_M1_5_39 ( .A(u4_sll_452_ML_int_5__39_), .B(
        u4_sll_452_ML_int_5__7_), .S(u4_sll_452_n47), .Z(
        u4_sll_452_ML_int_6__39_) );
  MUX2_X2 u4_sll_452_M1_5_40 ( .A(u4_sll_452_ML_int_5__40_), .B(
        u4_sll_452_ML_int_5__8_), .S(u4_sll_452_n47), .Z(
        u4_sll_452_ML_int_6__40_) );
  MUX2_X2 u4_sll_452_M1_5_41 ( .A(u4_sll_452_ML_int_5__41_), .B(
        u4_sll_452_ML_int_5__9_), .S(u4_sll_452_n47), .Z(
        u4_sll_452_ML_int_6__41_) );
  MUX2_X2 u4_sll_452_M1_5_42 ( .A(u4_sll_452_ML_int_5__42_), .B(
        u4_sll_452_ML_int_5__10_), .S(u4_sll_452_n47), .Z(
        u4_sll_452_ML_int_6__42_) );
  MUX2_X2 u4_sll_452_M1_5_43 ( .A(u4_sll_452_ML_int_5__43_), .B(
        u4_sll_452_ML_int_5__11_), .S(u4_sll_452_n47), .Z(
        u4_sll_452_ML_int_6__43_) );
  MUX2_X2 u4_sll_452_M1_5_44 ( .A(u4_sll_452_ML_int_5__44_), .B(
        u4_sll_452_ML_int_5__12_), .S(u4_sll_452_n47), .Z(
        u4_sll_452_ML_int_6__44_) );
  MUX2_X2 u4_sll_452_M1_5_45 ( .A(u4_sll_452_ML_int_5__45_), .B(
        u4_sll_452_ML_int_5__13_), .S(u4_sll_452_n47), .Z(
        u4_sll_452_ML_int_6__45_) );
  MUX2_X2 u4_sll_452_M1_5_46 ( .A(u4_sll_452_ML_int_5__46_), .B(
        u4_sll_452_ML_int_5__14_), .S(u4_sll_452_n47), .Z(
        u4_sll_452_ML_int_6__46_) );
  MUX2_X2 u4_sll_452_M1_5_47 ( .A(u4_sll_452_ML_int_5__47_), .B(
        u4_sll_452_ML_int_5__15_), .S(u4_sll_452_n47), .Z(
        u4_sll_452_ML_int_6__47_) );
  MUX2_X2 u4_sll_452_M1_5_48 ( .A(u4_sll_452_ML_int_5__48_), .B(
        u4_sll_452_ML_int_5__16_), .S(u4_sll_452_n47), .Z(
        u4_sll_452_ML_int_6__48_) );
  MUX2_X2 u4_sll_452_M1_5_49 ( .A(u4_sll_452_ML_int_5__49_), .B(
        u4_sll_452_ML_int_5__17_), .S(u4_sll_452_n47), .Z(
        u4_sll_452_ML_int_6__49_) );
  MUX2_X2 u4_sll_452_M1_5_50 ( .A(u4_sll_452_ML_int_5__50_), .B(
        u4_sll_452_ML_int_5__18_), .S(u4_sll_452_n47), .Z(
        u4_sll_452_ML_int_6__50_) );
  MUX2_X2 u4_sll_452_M1_5_51 ( .A(u4_sll_452_ML_int_5__51_), .B(
        u4_sll_452_ML_int_5__19_), .S(u4_sll_452_n47), .Z(
        u4_sll_452_ML_int_6__51_) );
  MUX2_X2 u4_sll_452_M1_5_52 ( .A(u4_sll_452_ML_int_5__52_), .B(
        u4_sll_452_ML_int_5__20_), .S(u4_sll_452_n47), .Z(
        u4_sll_452_ML_int_6__52_) );
  MUX2_X2 u4_sll_452_M1_5_53 ( .A(u4_sll_452_ML_int_5__53_), .B(
        u4_sll_452_ML_int_5__21_), .S(u4_sll_452_n47), .Z(
        u4_sll_452_ML_int_6__53_) );
  MUX2_X2 u4_sll_452_M1_5_54 ( .A(u4_sll_452_ML_int_5__54_), .B(
        u4_sll_452_ML_int_5__22_), .S(u4_sll_452_n47), .Z(
        u4_sll_452_ML_int_6__54_) );
  MUX2_X2 u4_sll_452_M1_5_55 ( .A(u4_sll_452_ML_int_5__55_), .B(
        u4_sll_452_ML_int_5__23_), .S(u4_sll_452_n47), .Z(
        u4_sll_452_ML_int_6__55_) );
  MUX2_X2 u4_sll_452_M1_5_56 ( .A(u4_sll_452_ML_int_5__56_), .B(
        u4_sll_452_ML_int_5__24_), .S(u4_sll_452_n48), .Z(
        u4_sll_452_ML_int_6__56_) );
  MUX2_X2 u4_sll_452_M1_5_57 ( .A(u4_sll_452_ML_int_5__57_), .B(
        u4_sll_452_ML_int_5__25_), .S(u4_sll_452_n48), .Z(
        u4_sll_452_ML_int_6__57_) );
  MUX2_X2 u4_sll_452_M1_5_58 ( .A(u4_sll_452_ML_int_5__58_), .B(
        u4_sll_452_ML_int_5__26_), .S(u4_sll_452_n48), .Z(
        u4_sll_452_ML_int_6__58_) );
  MUX2_X2 u4_sll_452_M1_5_59 ( .A(u4_sll_452_ML_int_5__59_), .B(
        u4_sll_452_ML_int_5__27_), .S(u4_sll_452_n48), .Z(
        u4_sll_452_ML_int_6__59_) );
  MUX2_X2 u4_sll_452_M1_5_60 ( .A(u4_sll_452_ML_int_5__60_), .B(
        u4_sll_452_ML_int_5__28_), .S(u4_sll_452_n48), .Z(
        u4_sll_452_ML_int_6__60_) );
  MUX2_X2 u4_sll_452_M1_5_61 ( .A(u4_sll_452_ML_int_5__61_), .B(
        u4_sll_452_ML_int_5__29_), .S(u4_sll_452_n48), .Z(
        u4_sll_452_ML_int_6__61_) );
  MUX2_X2 u4_sll_452_M1_5_62 ( .A(u4_sll_452_ML_int_5__62_), .B(
        u4_sll_452_ML_int_5__30_), .S(u4_sll_452_n48), .Z(
        u4_sll_452_ML_int_6__62_) );
  MUX2_X2 u4_sll_452_M1_5_63 ( .A(u4_sll_452_ML_int_5__63_), .B(
        u4_sll_452_ML_int_5__31_), .S(u4_sll_452_n48), .Z(
        u4_sll_452_ML_int_6__63_) );
  MUX2_X2 u4_sll_452_M1_5_64 ( .A(u4_sll_452_ML_int_5__64_), .B(
        u4_sll_452_ML_int_5__32_), .S(u4_sll_452_n48), .Z(
        u4_sll_452_ML_int_6__64_) );
  MUX2_X2 u4_sll_452_M1_5_65 ( .A(u4_sll_452_ML_int_5__65_), .B(
        u4_sll_452_ML_int_5__33_), .S(u4_sll_452_n48), .Z(
        u4_sll_452_ML_int_6__65_) );
  MUX2_X2 u4_sll_452_M1_5_66 ( .A(u4_sll_452_ML_int_5__66_), .B(
        u4_sll_452_ML_int_5__34_), .S(u4_sll_452_n48), .Z(
        u4_sll_452_ML_int_6__66_) );
  MUX2_X2 u4_sll_452_M1_5_67 ( .A(u4_sll_452_ML_int_5__67_), .B(
        u4_sll_452_ML_int_5__35_), .S(u4_sll_452_n48), .Z(
        u4_sll_452_ML_int_6__67_) );
  MUX2_X2 u4_sll_452_M1_5_68 ( .A(u4_sll_452_ML_int_5__68_), .B(
        u4_sll_452_ML_int_5__36_), .S(u4_sll_452_n48), .Z(
        u4_sll_452_ML_int_6__68_) );
  MUX2_X2 u4_sll_452_M1_5_69 ( .A(u4_sll_452_ML_int_5__69_), .B(
        u4_sll_452_ML_int_5__37_), .S(u4_sll_452_n48), .Z(
        u4_sll_452_ML_int_6__69_) );
  MUX2_X2 u4_sll_452_M1_5_70 ( .A(u4_sll_452_ML_int_5__70_), .B(
        u4_sll_452_ML_int_5__38_), .S(u4_sll_452_n48), .Z(
        u4_sll_452_ML_int_6__70_) );
  MUX2_X2 u4_sll_452_M1_5_71 ( .A(u4_sll_452_ML_int_5__71_), .B(
        u4_sll_452_ML_int_5__39_), .S(u4_sll_452_n48), .Z(
        u4_sll_452_ML_int_6__71_) );
  MUX2_X2 u4_sll_452_M1_5_72 ( .A(u4_sll_452_ML_int_5__72_), .B(
        u4_sll_452_ML_int_5__40_), .S(u4_sll_452_n48), .Z(
        u4_sll_452_ML_int_6__72_) );
  MUX2_X2 u4_sll_452_M1_5_73 ( .A(u4_sll_452_ML_int_5__73_), .B(
        u4_sll_452_ML_int_5__41_), .S(u4_sll_452_n48), .Z(
        u4_sll_452_ML_int_6__73_) );
  MUX2_X2 u4_sll_452_M1_5_74 ( .A(u4_sll_452_ML_int_5__74_), .B(
        u4_sll_452_ML_int_5__42_), .S(u4_sll_452_n49), .Z(
        u4_sll_452_ML_int_6__74_) );
  MUX2_X2 u4_sll_452_M1_5_75 ( .A(u4_sll_452_ML_int_5__75_), .B(
        u4_sll_452_ML_int_5__43_), .S(u4_sll_452_n49), .Z(
        u4_sll_452_ML_int_6__75_) );
  MUX2_X2 u4_sll_452_M1_5_76 ( .A(u4_sll_452_ML_int_5__76_), .B(
        u4_sll_452_ML_int_5__44_), .S(u4_sll_452_n49), .Z(
        u4_sll_452_ML_int_6__76_) );
  MUX2_X2 u4_sll_452_M1_5_77 ( .A(u4_sll_452_ML_int_5__77_), .B(
        u4_sll_452_ML_int_5__45_), .S(u4_sll_452_n49), .Z(
        u4_sll_452_ML_int_6__77_) );
  MUX2_X2 u4_sll_452_M1_5_78 ( .A(u4_sll_452_ML_int_5__78_), .B(
        u4_sll_452_ML_int_5__46_), .S(u4_sll_452_n49), .Z(
        u4_sll_452_ML_int_6__78_) );
  MUX2_X2 u4_sll_452_M1_5_79 ( .A(u4_sll_452_ML_int_5__79_), .B(
        u4_sll_452_ML_int_5__47_), .S(u4_sll_452_n49), .Z(
        u4_sll_452_ML_int_6__79_) );
  MUX2_X2 u4_sll_452_M1_5_80 ( .A(u4_sll_452_ML_int_5__80_), .B(
        u4_sll_452_ML_int_5__48_), .S(u4_sll_452_n49), .Z(
        u4_sll_452_ML_int_6__80_) );
  MUX2_X2 u4_sll_452_M1_5_81 ( .A(u4_sll_452_ML_int_5__81_), .B(
        u4_sll_452_ML_int_5__49_), .S(u4_sll_452_n49), .Z(
        u4_sll_452_ML_int_6__81_) );
  MUX2_X2 u4_sll_452_M1_5_82 ( .A(u4_sll_452_ML_int_5__82_), .B(
        u4_sll_452_ML_int_5__50_), .S(u4_sll_452_n49), .Z(
        u4_sll_452_ML_int_6__82_) );
  MUX2_X2 u4_sll_452_M1_5_83 ( .A(u4_sll_452_ML_int_5__83_), .B(
        u4_sll_452_ML_int_5__51_), .S(u4_sll_452_n49), .Z(
        u4_sll_452_ML_int_6__83_) );
  MUX2_X2 u4_sll_452_M1_5_84 ( .A(u4_sll_452_ML_int_5__84_), .B(
        u4_sll_452_ML_int_5__52_), .S(u4_sll_452_n49), .Z(
        u4_sll_452_ML_int_6__84_) );
  MUX2_X2 u4_sll_452_M1_5_85 ( .A(u4_sll_452_ML_int_5__85_), .B(
        u4_sll_452_ML_int_5__53_), .S(u4_sll_452_n49), .Z(
        u4_sll_452_ML_int_6__85_) );
  MUX2_X2 u4_sll_452_M1_5_86 ( .A(u4_sll_452_ML_int_5__86_), .B(
        u4_sll_452_ML_int_5__54_), .S(u4_sll_452_n49), .Z(
        u4_sll_452_ML_int_6__86_) );
  MUX2_X2 u4_sll_452_M1_5_87 ( .A(u4_sll_452_ML_int_5__87_), .B(
        u4_sll_452_ML_int_5__55_), .S(u4_sll_452_n49), .Z(
        u4_sll_452_ML_int_6__87_) );
  MUX2_X2 u4_sll_452_M1_5_88 ( .A(u4_sll_452_ML_int_5__88_), .B(
        u4_sll_452_ML_int_5__56_), .S(u4_sll_452_n49), .Z(
        u4_sll_452_ML_int_6__88_) );
  MUX2_X2 u4_sll_452_M1_5_89 ( .A(u4_sll_452_ML_int_5__89_), .B(
        u4_sll_452_ML_int_5__57_), .S(u4_sll_452_n49), .Z(
        u4_sll_452_ML_int_6__89_) );
  MUX2_X2 u4_sll_452_M1_5_90 ( .A(u4_sll_452_ML_int_5__90_), .B(
        u4_sll_452_ML_int_5__58_), .S(u4_sll_452_n49), .Z(
        u4_sll_452_ML_int_6__90_) );
  MUX2_X2 u4_sll_452_M1_5_91 ( .A(u4_sll_452_ML_int_5__91_), .B(
        u4_sll_452_ML_int_5__59_), .S(u4_sll_452_n49), .Z(
        u4_sll_452_ML_int_6__91_) );
  MUX2_X2 u4_sll_452_M1_5_92 ( .A(u4_sll_452_ML_int_5__92_), .B(
        u4_sll_452_ML_int_5__60_), .S(u4_sll_452_n45), .Z(
        u4_sll_452_ML_int_6__92_) );
  MUX2_X2 u4_sll_452_M1_5_93 ( .A(u4_sll_452_ML_int_5__93_), .B(
        u4_sll_452_ML_int_5__61_), .S(u4_sll_452_n45), .Z(
        u4_sll_452_ML_int_6__93_) );
  MUX2_X2 u4_sll_452_M1_5_94 ( .A(u4_sll_452_ML_int_5__94_), .B(
        u4_sll_452_ML_int_5__62_), .S(u4_sll_452_n45), .Z(
        u4_sll_452_ML_int_6__94_) );
  MUX2_X2 u4_sll_452_M1_5_95 ( .A(u4_sll_452_ML_int_5__95_), .B(
        u4_sll_452_ML_int_5__63_), .S(u4_sll_452_n45), .Z(
        u4_sll_452_ML_int_6__95_) );
  MUX2_X2 u4_sll_452_M1_5_96 ( .A(u4_sll_452_ML_int_5__96_), .B(
        u4_sll_452_ML_int_5__64_), .S(u4_sll_452_n45), .Z(
        u4_sll_452_ML_int_6__96_) );
  MUX2_X2 u4_sll_452_M1_5_97 ( .A(u4_sll_452_ML_int_5__97_), .B(
        u4_sll_452_ML_int_5__65_), .S(u4_sll_452_n45), .Z(
        u4_sll_452_ML_int_6__97_) );
  MUX2_X2 u4_sll_452_M1_5_98 ( .A(u4_sll_452_ML_int_5__98_), .B(
        u4_sll_452_ML_int_5__66_), .S(u4_sll_452_n45), .Z(
        u4_sll_452_ML_int_6__98_) );
  MUX2_X2 u4_sll_452_M1_5_99 ( .A(u4_sll_452_ML_int_5__99_), .B(
        u4_sll_452_ML_int_5__67_), .S(u4_sll_452_n45), .Z(
        u4_sll_452_ML_int_6__99_) );
  MUX2_X2 u4_sll_452_M1_5_100 ( .A(u4_sll_452_ML_int_5__100_), .B(
        u4_sll_452_ML_int_5__68_), .S(u4_sll_452_n45), .Z(
        u4_sll_452_ML_int_6__100_) );
  MUX2_X2 u4_sll_452_M1_5_101 ( .A(u4_sll_452_ML_int_5__101_), .B(
        u4_sll_452_ML_int_5__69_), .S(u4_sll_452_n45), .Z(
        u4_sll_452_ML_int_6__101_) );
  MUX2_X2 u4_sll_452_M1_5_102 ( .A(u4_sll_452_ML_int_5__102_), .B(
        u4_sll_452_ML_int_5__70_), .S(u4_sll_452_n45), .Z(
        u4_sll_452_ML_int_6__102_) );
  MUX2_X2 u4_sll_452_M1_5_103 ( .A(u4_sll_452_ML_int_5__103_), .B(
        u4_sll_452_ML_int_5__71_), .S(u4_sll_452_n45), .Z(
        u4_sll_452_ML_int_6__103_) );
  MUX2_X2 u4_sll_452_M1_5_104 ( .A(u4_sll_452_ML_int_5__104_), .B(
        u4_sll_452_ML_int_5__72_), .S(u4_sll_452_n45), .Z(
        u4_sll_452_ML_int_6__104_) );
  MUX2_X2 u4_sll_452_M1_5_105 ( .A(u4_sll_452_ML_int_5__105_), .B(
        u4_sll_452_ML_int_5__73_), .S(u4_sll_452_n45), .Z(
        u4_sll_452_ML_int_6__105_) );
  MUX2_X2 u4_sll_452_M1_6_64 ( .A(u4_sll_452_ML_int_6__64_), .B(
        u4_sll_452_ML_int_6__0_), .S(u4_sll_452_n39), .Z(
        u4_sll_452_ML_int_7__64_) );
  MUX2_X2 u4_sll_452_M1_6_65 ( .A(u4_sll_452_ML_int_6__65_), .B(
        u4_sll_452_ML_int_6__1_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__65_) );
  MUX2_X2 u4_sll_452_M1_6_66 ( .A(u4_sll_452_ML_int_6__66_), .B(
        u4_sll_452_ML_int_6__2_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__66_) );
  MUX2_X2 u4_sll_452_M1_6_67 ( .A(u4_sll_452_ML_int_6__67_), .B(
        u4_sll_452_ML_int_6__3_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__67_) );
  MUX2_X2 u4_sll_452_M1_6_68 ( .A(u4_sll_452_ML_int_6__68_), .B(
        u4_sll_452_ML_int_6__4_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__68_) );
  MUX2_X2 u4_sll_452_M1_6_69 ( .A(u4_sll_452_ML_int_6__69_), .B(
        u4_sll_452_ML_int_6__5_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__69_) );
  MUX2_X2 u4_sll_452_M1_6_70 ( .A(u4_sll_452_ML_int_6__70_), .B(
        u4_sll_452_ML_int_6__6_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__70_) );
  MUX2_X2 u4_sll_452_M1_6_71 ( .A(u4_sll_452_ML_int_6__71_), .B(
        u4_sll_452_ML_int_6__7_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__71_) );
  MUX2_X2 u4_sll_452_M1_6_72 ( .A(u4_sll_452_ML_int_6__72_), .B(
        u4_sll_452_ML_int_6__8_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__72_) );
  MUX2_X2 u4_sll_452_M1_6_73 ( .A(u4_sll_452_ML_int_6__73_), .B(
        u4_sll_452_ML_int_6__9_), .S(u4_sll_452_n39), .Z(
        u4_sll_452_ML_int_7__73_) );
  MUX2_X2 u4_sll_452_M1_6_74 ( .A(u4_sll_452_ML_int_6__74_), .B(
        u4_sll_452_ML_int_6__10_), .S(u4_sll_452_n39), .Z(
        u4_sll_452_ML_int_7__74_) );
  MUX2_X2 u4_sll_452_M1_6_75 ( .A(u4_sll_452_ML_int_6__75_), .B(
        u4_sll_452_ML_int_6__11_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__75_) );
  MUX2_X2 u4_sll_452_M1_6_76 ( .A(u4_sll_452_ML_int_6__76_), .B(
        u4_sll_452_ML_int_6__12_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__76_) );
  MUX2_X2 u4_sll_452_M1_6_77 ( .A(u4_sll_452_ML_int_6__77_), .B(
        u4_sll_452_ML_int_6__13_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__77_) );
  MUX2_X2 u4_sll_452_M1_6_78 ( .A(u4_sll_452_ML_int_6__78_), .B(
        u4_sll_452_ML_int_6__14_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__78_) );
  MUX2_X2 u4_sll_452_M1_6_79 ( .A(u4_sll_452_ML_int_6__79_), .B(
        u4_sll_452_ML_int_6__15_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__79_) );
  MUX2_X2 u4_sll_452_M1_6_80 ( .A(u4_sll_452_ML_int_6__80_), .B(
        u4_sll_452_ML_int_6__16_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__80_) );
  MUX2_X2 u4_sll_452_M1_6_81 ( .A(u4_sll_452_ML_int_6__81_), .B(
        u4_sll_452_ML_int_6__17_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__81_) );
  MUX2_X2 u4_sll_452_M1_6_82 ( .A(u4_sll_452_ML_int_6__82_), .B(
        u4_sll_452_ML_int_6__18_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__82_) );
  MUX2_X2 u4_sll_452_M1_6_83 ( .A(u4_sll_452_ML_int_6__83_), .B(
        u4_sll_452_ML_int_6__19_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__83_) );
  MUX2_X2 u4_sll_452_M1_6_84 ( .A(u4_sll_452_ML_int_6__84_), .B(
        u4_sll_452_ML_int_6__20_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__84_) );
  MUX2_X2 u4_sll_452_M1_6_85 ( .A(u4_sll_452_ML_int_6__85_), .B(
        u4_sll_452_ML_int_6__21_), .S(u4_sll_452_n39), .Z(
        u4_sll_452_ML_int_7__85_) );
  MUX2_X2 u4_sll_452_M1_6_86 ( .A(u4_sll_452_ML_int_6__86_), .B(
        u4_sll_452_ML_int_6__22_), .S(u4_sll_452_n39), .Z(
        u4_sll_452_ML_int_7__86_) );
  MUX2_X2 u4_sll_452_M1_6_87 ( .A(u4_sll_452_ML_int_6__87_), .B(
        u4_sll_452_ML_int_6__23_), .S(u4_sll_452_n39), .Z(
        u4_sll_452_ML_int_7__87_) );
  MUX2_X2 u4_sll_452_M1_6_88 ( .A(u4_sll_452_ML_int_6__88_), .B(
        u4_sll_452_ML_int_6__24_), .S(u4_sll_452_n39), .Z(
        u4_sll_452_ML_int_7__88_) );
  MUX2_X2 u4_sll_452_M1_6_89 ( .A(u4_sll_452_ML_int_6__89_), .B(
        u4_sll_452_ML_int_6__25_), .S(u4_sll_452_n39), .Z(
        u4_sll_452_ML_int_7__89_) );
  MUX2_X2 u4_sll_452_M1_6_90 ( .A(u4_sll_452_ML_int_6__90_), .B(
        u4_sll_452_ML_int_6__26_), .S(u4_sll_452_n39), .Z(
        u4_sll_452_ML_int_7__90_) );
  MUX2_X2 u4_sll_452_M1_6_91 ( .A(u4_sll_452_ML_int_6__91_), .B(
        u4_sll_452_ML_int_6__27_), .S(u4_sll_452_n39), .Z(
        u4_sll_452_ML_int_7__91_) );
  MUX2_X2 u4_sll_452_M1_6_92 ( .A(u4_sll_452_ML_int_6__92_), .B(
        u4_sll_452_ML_int_6__28_), .S(u4_sll_452_n39), .Z(
        u4_sll_452_ML_int_7__92_) );
  MUX2_X2 u4_sll_452_M1_6_93 ( .A(u4_sll_452_ML_int_6__93_), .B(
        u4_sll_452_ML_int_6__29_), .S(u4_sll_452_n39), .Z(
        u4_sll_452_ML_int_7__93_) );
  MUX2_X2 u4_sll_452_M1_6_94 ( .A(u4_sll_452_ML_int_6__94_), .B(
        u4_sll_452_ML_int_6__30_), .S(u4_sll_452_n39), .Z(
        u4_sll_452_ML_int_7__94_) );
  MUX2_X2 u4_sll_452_M1_6_95 ( .A(u4_sll_452_ML_int_6__95_), .B(
        u4_sll_452_ML_int_6__31_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__95_) );
  MUX2_X2 u4_sll_452_M1_6_96 ( .A(u4_sll_452_ML_int_6__96_), .B(
        u4_sll_452_ML_int_6__32_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__96_) );
  MUX2_X2 u4_sll_452_M1_6_97 ( .A(u4_sll_452_ML_int_6__97_), .B(
        u4_sll_452_ML_int_6__33_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__97_) );
  MUX2_X2 u4_sll_452_M1_6_98 ( .A(u4_sll_452_ML_int_6__98_), .B(
        u4_sll_452_ML_int_6__34_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__98_) );
  MUX2_X2 u4_sll_452_M1_6_99 ( .A(u4_sll_452_ML_int_6__99_), .B(
        u4_sll_452_ML_int_6__35_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__99_) );
  MUX2_X2 u4_sll_452_M1_6_100 ( .A(u4_sll_452_ML_int_6__100_), .B(
        u4_sll_452_ML_int_6__36_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__100_) );
  MUX2_X2 u4_sll_452_M1_6_101 ( .A(u4_sll_452_ML_int_6__101_), .B(
        u4_sll_452_ML_int_6__37_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__101_) );
  MUX2_X2 u4_sll_452_M1_6_102 ( .A(u4_sll_452_ML_int_6__102_), .B(
        u4_sll_452_ML_int_6__38_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__102_) );
  MUX2_X2 u4_sll_452_M1_6_103 ( .A(u4_sll_452_ML_int_6__103_), .B(
        u4_sll_452_ML_int_6__39_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__103_) );
  MUX2_X2 u4_sll_452_M1_6_104 ( .A(u4_sll_452_ML_int_6__104_), .B(
        u4_sll_452_ML_int_6__40_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__104_) );
  MUX2_X2 u4_sll_452_M1_6_105 ( .A(u4_sll_452_ML_int_6__105_), .B(
        u4_sll_452_ML_int_6__41_), .S(u4_sll_452_n40), .Z(
        u4_sll_452_ML_int_7__105_) );
  NOR2_X1 u4_srl_451_U991 ( .A1(u4_shift_right[1]), .A2(u4_shift_right[7]), 
        .ZN(u4_srl_451_n882) );
  INV_X1 u4_srl_451_U990 ( .A(u4_shift_right[0]), .ZN(u4_srl_451_n883) );
  NAND2_X1 u4_srl_451_U989 ( .A1(u4_srl_451_n882), .A2(u4_srl_451_n883), .ZN(
        u4_srl_451_n400) );
  AOI22_X1 u4_srl_451_U988 ( .A1(fract_denorm[71]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[70]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n881) );
  OAI221_X1 u4_srl_451_U987 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n131), .C1(
        u4_srl_451_n40), .C2(u4_srl_451_n130), .A(u4_srl_451_n881), .ZN(
        u4_srl_451_n508) );
  INV_X1 u4_srl_451_U986 ( .A(u4_srl_451_n508), .ZN(u4_srl_451_n603) );
  NOR2_X1 u4_srl_451_U985 ( .A1(u4_shift_right[3]), .A2(u4_shift_right[7]), 
        .ZN(u4_srl_451_n837) );
  INV_X1 u4_srl_451_U984 ( .A(u4_srl_451_n837), .ZN(u4_srl_451_n732) );
  INV_X1 u4_srl_451_U983 ( .A(u4_shift_right[2]), .ZN(u4_srl_451_n838) );
  NOR2_X1 u4_srl_451_U982 ( .A1(u4_srl_451_n732), .A2(u4_srl_451_n838), .ZN(
        u4_srl_451_n398) );
  AOI22_X1 u4_srl_451_U981 ( .A1(fract_denorm[67]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[66]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n880) );
  OAI221_X1 u4_srl_451_U980 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n127), .C1(
        u4_srl_451_n40), .C2(u4_srl_451_n126), .A(u4_srl_451_n880), .ZN(
        u4_srl_451_n509) );
  INV_X1 u4_srl_451_U979 ( .A(u4_srl_451_n509), .ZN(u4_srl_451_n750) );
  NOR2_X1 u4_srl_451_U978 ( .A1(u4_srl_451_n838), .A2(u4_srl_451_n837), .ZN(
        u4_srl_451_n399) );
  AOI22_X1 u4_srl_451_U977 ( .A1(fract_denorm[79]), .A2(u4_srl_451_n50), .B1(
        fract_denorm[78]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n879) );
  OAI221_X1 u4_srl_451_U976 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n139), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n138), .A(u4_srl_451_n879), .ZN(
        u4_srl_451_n605) );
  AOI22_X1 u4_srl_451_U975 ( .A1(fract_denorm[75]), .A2(u4_srl_451_n50), .B1(
        fract_denorm[74]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n878) );
  OAI221_X1 u4_srl_451_U974 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n135), .C1(
        u4_srl_451_n43), .C2(u4_srl_451_n134), .A(u4_srl_451_n878), .ZN(
        u4_srl_451_n606) );
  AOI22_X1 u4_srl_451_U973 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n605), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n606), .ZN(u4_srl_451_n877) );
  OAI221_X1 u4_srl_451_U972 ( .B1(u4_srl_451_n603), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n750), .C2(u4_srl_451_n64), .A(u4_srl_451_n877), .ZN(
        u4_srl_451_n427) );
  NOR2_X1 u4_srl_451_U971 ( .A1(u4_shift_right[5]), .A2(u4_shift_right[7]), 
        .ZN(u4_srl_451_n271) );
  INV_X1 u4_srl_451_U970 ( .A(u4_srl_451_n243), .ZN(u4_srl_451_n405) );
  AOI22_X1 u4_srl_451_U969 ( .A1(fract_denorm[103]), .A2(u4_srl_451_n50), .B1(
        fract_denorm[102]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n876) );
  OAI221_X1 u4_srl_451_U968 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n163), .C1(
        u4_srl_451_n41), .C2(u4_srl_451_n162), .A(u4_srl_451_n876), .ZN(
        u4_srl_451_n503) );
  AOI22_X1 u4_srl_451_U967 ( .A1(u4_srl_451_n45), .A2(fract_denorm[104]), .B1(
        u4_srl_451_n38), .B2(n4873), .ZN(u4_srl_451_n249) );
  INV_X1 u4_srl_451_U966 ( .A(u4_srl_451_n249), .ZN(u4_srl_451_n385) );
  AOI22_X1 u4_srl_451_U965 ( .A1(fract_denorm[99]), .A2(u4_srl_451_n50), .B1(
        fract_denorm[98]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n875) );
  OAI221_X1 u4_srl_451_U964 ( .B1(u4_srl_451_n32), .B2(u4_srl_451_n159), .C1(
        u4_srl_451_n44), .C2(u4_srl_451_n158), .A(u4_srl_451_n875), .ZN(
        u4_srl_451_n504) );
  AOI222_X1 u4_srl_451_U963 ( .A1(u4_srl_451_n503), .A2(u4_srl_451_n16), .B1(
        u4_srl_451_n385), .B2(u4_srl_451_n26), .C1(u4_srl_451_n504), .C2(
        u4_srl_451_n60), .ZN(u4_srl_451_n189) );
  INV_X1 u4_srl_451_U962 ( .A(u4_srl_451_n189), .ZN(u4_srl_451_n351) );
  NOR2_X1 u4_srl_451_U961 ( .A1(u4_shift_right[4]), .A2(u4_srl_451_n271), .ZN(
        u4_srl_451_n341) );
  AOI22_X1 u4_srl_451_U960 ( .A1(fract_denorm[87]), .A2(u4_srl_451_n50), .B1(
        fract_denorm[86]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n874) );
  OAI221_X1 u4_srl_451_U959 ( .B1(u4_srl_451_n36), .B2(u4_srl_451_n147), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n146), .A(u4_srl_451_n874), .ZN(
        u4_srl_451_n498) );
  INV_X1 u4_srl_451_U958 ( .A(u4_srl_451_n498), .ZN(u4_srl_451_n607) );
  AOI22_X1 u4_srl_451_U957 ( .A1(fract_denorm[83]), .A2(u4_srl_451_n50), .B1(
        fract_denorm[82]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n873) );
  OAI221_X1 u4_srl_451_U956 ( .B1(u4_srl_451_n36), .B2(u4_srl_451_n143), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n142), .A(u4_srl_451_n873), .ZN(
        u4_srl_451_n499) );
  INV_X1 u4_srl_451_U955 ( .A(u4_srl_451_n499), .ZN(u4_srl_451_n752) );
  AOI22_X1 u4_srl_451_U954 ( .A1(fract_denorm[95]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[94]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n872) );
  OAI221_X1 u4_srl_451_U953 ( .B1(u4_srl_451_n36), .B2(u4_srl_451_n155), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n154), .A(u4_srl_451_n872), .ZN(
        u4_srl_451_n609) );
  AOI22_X1 u4_srl_451_U952 ( .A1(fract_denorm[91]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[90]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n871) );
  OAI221_X1 u4_srl_451_U951 ( .B1(u4_srl_451_n36), .B2(u4_srl_451_n151), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n150), .A(u4_srl_451_n871), .ZN(
        u4_srl_451_n610) );
  AOI22_X1 u4_srl_451_U950 ( .A1(u4_srl_451_n24), .A2(u4_srl_451_n609), .B1(
        u4_srl_451_n30), .B2(u4_srl_451_n610), .ZN(u4_srl_451_n870) );
  OAI221_X1 u4_srl_451_U949 ( .B1(u4_srl_451_n607), .B2(u4_srl_451_n19), .C1(
        u4_srl_451_n752), .C2(u4_srl_451_n63), .A(u4_srl_451_n870), .ZN(
        u4_srl_451_n352) );
  INV_X1 u4_srl_451_U948 ( .A(u4_srl_451_n247), .ZN(u4_srl_451_n406) );
  AOI222_X1 u4_srl_451_U947 ( .A1(u4_srl_451_n427), .A2(u4_srl_451_n405), .B1(
        u4_srl_451_n351), .B2(u4_srl_451_n341), .C1(u4_srl_451_n352), .C2(
        u4_srl_451_n406), .ZN(u4_srl_451_n277) );
  NOR2_X1 u4_srl_451_U946 ( .A1(u4_shift_right[6]), .A2(u4_shift_right[7]), 
        .ZN(u4_srl_451_n863) );
  NOR2_X1 u4_srl_451_U945 ( .A1(u4_srl_451_n863), .A2(u4_shift_right[8]), .ZN(
        u4_srl_451_n381) );
  AOI22_X1 u4_srl_451_U944 ( .A1(fract_denorm[55]), .A2(u4_srl_451_n50), .B1(
        fract_denorm[54]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n869) );
  OAI221_X1 u4_srl_451_U943 ( .B1(u4_srl_451_n36), .B2(u4_srl_451_n115), .C1(
        u4_srl_451_n44), .C2(u4_srl_451_n114), .A(u4_srl_451_n869), .ZN(
        u4_srl_451_n521) );
  AOI22_X1 u4_srl_451_U942 ( .A1(fract_denorm[51]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[50]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n868) );
  OAI221_X1 u4_srl_451_U941 ( .B1(u4_srl_451_n36), .B2(u4_srl_451_n111), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n110), .A(u4_srl_451_n868), .ZN(
        u4_srl_451_n522) );
  AOI22_X1 u4_srl_451_U940 ( .A1(fract_denorm[63]), .A2(u4_srl_451_n50), .B1(
        fract_denorm[62]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n867) );
  OAI221_X1 u4_srl_451_U939 ( .B1(u4_srl_451_n36), .B2(u4_srl_451_n123), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n122), .A(u4_srl_451_n867), .ZN(
        u4_srl_451_n613) );
  AOI22_X1 u4_srl_451_U938 ( .A1(fract_denorm[59]), .A2(u4_srl_451_n50), .B1(
        fract_denorm[58]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n866) );
  OAI221_X1 u4_srl_451_U937 ( .B1(u4_srl_451_n36), .B2(u4_srl_451_n119), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n118), .A(u4_srl_451_n866), .ZN(
        u4_srl_451_n510) );
  AOI22_X1 u4_srl_451_U936 ( .A1(u4_srl_451_n24), .A2(u4_srl_451_n613), .B1(
        u4_srl_451_n30), .B2(u4_srl_451_n510), .ZN(u4_srl_451_n865) );
  INV_X1 u4_srl_451_U935 ( .A(u4_srl_451_n865), .ZN(u4_srl_451_n864) );
  AOI221_X1 u4_srl_451_U934 ( .B1(u4_srl_451_n521), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n522), .C2(u4_srl_451_n60), .A(u4_srl_451_n864), .ZN(
        u4_srl_451_n349) );
  NOR2_X1 u4_srl_451_U933 ( .A1(u4_srl_451_n179), .A2(u4_srl_451_n271), .ZN(
        u4_srl_451_n805) );
  INV_X1 u4_srl_451_U932 ( .A(u4_shift_right[8]), .ZN(u4_srl_451_n862) );
  NAND2_X1 u4_srl_451_U931 ( .A1(u4_srl_451_n805), .A2(u4_srl_451_n862), .ZN(
        u4_srl_451_n304) );
  NOR2_X1 u4_srl_451_U930 ( .A1(u4_srl_451_n304), .A2(u4_srl_451_n397), .ZN(
        u4_srl_451_n317) );
  AOI22_X1 u4_srl_451_U929 ( .A1(fract_denorm[39]), .A2(u4_srl_451_n50), .B1(
        fract_denorm[38]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n861) );
  OAI221_X1 u4_srl_451_U928 ( .B1(u4_srl_451_n36), .B2(u4_srl_451_n99), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n98), .A(u4_srl_451_n861), .ZN(
        u4_srl_451_n514) );
  AOI22_X1 u4_srl_451_U927 ( .A1(fract_denorm[35]), .A2(u4_srl_451_n50), .B1(
        fract_denorm[34]), .B2(u4_srl_451_n54), .ZN(u4_srl_451_n860) );
  OAI221_X1 u4_srl_451_U926 ( .B1(u4_srl_451_n36), .B2(u4_srl_451_n95), .C1(
        u4_srl_451_n44), .C2(u4_srl_451_n94), .A(u4_srl_451_n860), .ZN(
        u4_srl_451_n515) );
  AOI22_X1 u4_srl_451_U925 ( .A1(fract_denorm[47]), .A2(u4_srl_451_n50), .B1(
        fract_denorm[46]), .B2(u4_srl_451_n54), .ZN(u4_srl_451_n859) );
  OAI221_X1 u4_srl_451_U924 ( .B1(u4_srl_451_n36), .B2(u4_srl_451_n107), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n106), .A(u4_srl_451_n859), .ZN(
        u4_srl_451_n517) );
  AOI22_X1 u4_srl_451_U923 ( .A1(fract_denorm[43]), .A2(u4_srl_451_n50), .B1(
        fract_denorm[42]), .B2(u4_srl_451_n54), .ZN(u4_srl_451_n858) );
  OAI221_X1 u4_srl_451_U922 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n103), .C1(
        u4_srl_451_n44), .C2(u4_srl_451_n102), .A(u4_srl_451_n858), .ZN(
        u4_srl_451_n518) );
  AOI22_X1 u4_srl_451_U921 ( .A1(u4_srl_451_n24), .A2(u4_srl_451_n517), .B1(
        u4_srl_451_n30), .B2(u4_srl_451_n518), .ZN(u4_srl_451_n857) );
  INV_X1 u4_srl_451_U920 ( .A(u4_srl_451_n857), .ZN(u4_srl_451_n856) );
  AOI221_X1 u4_srl_451_U919 ( .B1(u4_srl_451_n514), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n515), .C2(u4_srl_451_n61), .A(u4_srl_451_n856), .ZN(
        u4_srl_451_n425) );
  INV_X1 u4_srl_451_U918 ( .A(u4_srl_451_n425), .ZN(u4_srl_451_n841) );
  NAND2_X1 u4_srl_451_U917 ( .A1(u4_srl_451_n215), .A2(u4_srl_451_n271), .ZN(
        u4_srl_451_n209) );
  INV_X1 u4_srl_451_U916 ( .A(u4_srl_451_n209), .ZN(u4_srl_451_n391) );
  OAI22_X1 u4_srl_451_U915 ( .A1(u4_srl_451_n58), .A2(u4_srl_451_n65), .B1(
        u4_srl_451_n1), .B2(u4_srl_451_n66), .ZN(u4_srl_451_n855) );
  AOI221_X1 u4_srl_451_U914 ( .B1(fract_denorm[1]), .B2(u4_srl_451_n38), .C1(
        fract_denorm[0]), .C2(u4_srl_451_n45), .A(u4_srl_451_n855), .ZN(
        u4_srl_451_n843) );
  NAND2_X1 u4_srl_451_U913 ( .A1(u4_srl_451_n61), .A2(u4_srl_451_n397), .ZN(
        u4_srl_451_n270) );
  OAI22_X1 u4_srl_451_U912 ( .A1(u4_srl_451_n85), .A2(u4_srl_451_n1), .B1(
        u4_srl_451_n84), .B2(u4_srl_451_n58), .ZN(u4_srl_451_n854) );
  AOI221_X1 u4_srl_451_U911 ( .B1(u4_srl_451_n38), .B2(fract_denorm[21]), .C1(
        u4_srl_451_n45), .C2(fract_denorm[20]), .A(u4_srl_451_n854), .ZN(
        u4_srl_451_n202) );
  AOI22_X1 u4_srl_451_U910 ( .A1(fract_denorm[19]), .A2(u4_srl_451_n50), .B1(
        fract_denorm[18]), .B2(u4_srl_451_n54), .ZN(u4_srl_451_n853) );
  OAI221_X1 u4_srl_451_U909 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n80), .C1(
        u4_srl_451_n44), .C2(u4_srl_451_n79), .A(u4_srl_451_n853), .ZN(
        u4_srl_451_n332) );
  INV_X1 u4_srl_451_U908 ( .A(u4_srl_451_n332), .ZN(u4_srl_451_n201) );
  AOI22_X1 u4_srl_451_U907 ( .A1(fract_denorm[31]), .A2(u4_srl_451_n50), .B1(
        fract_denorm[30]), .B2(u4_srl_451_n54), .ZN(u4_srl_451_n852) );
  OAI221_X1 u4_srl_451_U906 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n91), .C1(
        u4_srl_451_n44), .C2(u4_srl_451_n90), .A(u4_srl_451_n852), .ZN(
        u4_srl_451_n516) );
  AOI22_X1 u4_srl_451_U905 ( .A1(fract_denorm[27]), .A2(u4_srl_451_n50), .B1(
        fract_denorm[26]), .B2(u4_srl_451_n54), .ZN(u4_srl_451_n851) );
  OAI221_X1 u4_srl_451_U904 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n87), .C1(
        u4_srl_451_n86), .C2(u4_srl_451_n40), .A(u4_srl_451_n851), .ZN(
        u4_srl_451_n745) );
  AOI22_X1 u4_srl_451_U903 ( .A1(u4_srl_451_n24), .A2(u4_srl_451_n516), .B1(
        u4_srl_451_n30), .B2(u4_srl_451_n745), .ZN(u4_srl_451_n850) );
  OAI221_X1 u4_srl_451_U902 ( .B1(u4_srl_451_n202), .B2(u4_srl_451_n19), .C1(
        u4_srl_451_n201), .C2(u4_srl_451_n63), .A(u4_srl_451_n850), .ZN(
        u4_srl_451_n849) );
  INV_X1 u4_srl_451_U901 ( .A(u4_srl_451_n849), .ZN(u4_srl_451_n677) );
  AOI22_X1 u4_srl_451_U900 ( .A1(fract_denorm[7]), .A2(u4_srl_451_n50), .B1(
        fract_denorm[6]), .B2(u4_srl_451_n54), .ZN(u4_srl_451_n848) );
  OAI221_X1 u4_srl_451_U899 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n68), .C1(
        u4_srl_451_n44), .C2(u4_srl_451_n67), .A(u4_srl_451_n848), .ZN(
        u4_srl_451_n335) );
  AOI22_X1 u4_srl_451_U898 ( .A1(fract_denorm[15]), .A2(u4_srl_451_n50), .B1(
        fract_denorm[14]), .B2(u4_srl_451_n54), .ZN(u4_srl_451_n847) );
  OAI221_X1 u4_srl_451_U897 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n76), .C1(
        u4_srl_451_n44), .C2(u4_srl_451_n75), .A(u4_srl_451_n847), .ZN(
        u4_srl_451_n198) );
  AOI22_X1 u4_srl_451_U896 ( .A1(fract_denorm[11]), .A2(u4_srl_451_n50), .B1(
        fract_denorm[10]), .B2(u4_srl_451_n54), .ZN(u4_srl_451_n846) );
  OAI221_X1 u4_srl_451_U895 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n72), .C1(
        u4_srl_451_n44), .C2(u4_srl_451_n71), .A(u4_srl_451_n846), .ZN(
        u4_srl_451_n199) );
  AOI222_X1 u4_srl_451_U894 ( .A1(u4_srl_451_n16), .A2(u4_srl_451_n335), .B1(
        u4_srl_451_n21), .B2(u4_srl_451_n198), .C1(u4_srl_451_n26), .C2(
        u4_srl_451_n199), .ZN(u4_srl_451_n845) );
  MUX2_X1 u4_srl_451_U893 ( .A(u4_srl_451_n677), .B(u4_srl_451_n845), .S(
        u4_srl_451_n397), .Z(u4_srl_451_n844) );
  OAI21_X1 u4_srl_451_U892 ( .B1(u4_srl_451_n843), .B2(u4_srl_451_n270), .A(
        u4_srl_451_n844), .ZN(u4_srl_451_n842) );
  AOI22_X1 u4_srl_451_U891 ( .A1(u4_srl_451_n15), .A2(u4_srl_451_n841), .B1(
        u4_srl_451_n391), .B2(u4_srl_451_n842), .ZN(u4_srl_451_n840) );
  OAI221_X1 u4_srl_451_U890 ( .B1(u4_srl_451_n277), .B2(u4_srl_451_n388), .C1(
        u4_srl_451_n349), .C2(u4_srl_451_n12), .A(u4_srl_451_n840), .ZN(
        u4_N5900) );
  AOI22_X1 u4_srl_451_U889 ( .A1(u4_srl_451_n503), .A2(u4_srl_451_n61), .B1(
        u4_srl_451_n385), .B2(u4_srl_451_n17), .ZN(u4_srl_451_n339) );
  NAND2_X1 u4_srl_451_U888 ( .A1(u4_srl_451_n391), .A2(u4_srl_451_n397), .ZN(
        u4_srl_451_n186) );
  NOR2_X1 u4_srl_451_U887 ( .A1(u4_srl_451_n339), .A2(u4_srl_451_n9), .ZN(
        u4_N6000) );
  NAND2_X1 u4_srl_451_U886 ( .A1(n4873), .A2(u4_srl_451_n45), .ZN(
        u4_srl_451_n245) );
  INV_X1 u4_srl_451_U885 ( .A(u4_srl_451_n245), .ZN(u4_srl_451_n669) );
  AOI22_X1 u4_srl_451_U884 ( .A1(fract_denorm[104]), .A2(u4_srl_451_n50), .B1(
        fract_denorm[103]), .B2(u4_srl_451_n54), .ZN(u4_srl_451_n839) );
  OAI221_X1 u4_srl_451_U883 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n164), .C1(
        u4_srl_451_n44), .C2(u4_srl_451_n163), .A(u4_srl_451_n839), .ZN(
        u4_srl_451_n473) );
  MUX2_X1 u4_srl_451_U882 ( .A(u4_srl_451_n669), .B(u4_srl_451_n473), .S(
        u4_srl_451_n838), .Z(u4_srl_451_n733) );
  NAND2_X1 u4_srl_451_U881 ( .A1(u4_srl_451_n837), .A2(u4_srl_451_n733), .ZN(
        u4_srl_451_n297) );
  NOR2_X1 u4_srl_451_U880 ( .A1(u4_srl_451_n186), .A2(u4_srl_451_n297), .ZN(
        u4_N6001) );
  AOI22_X1 u4_srl_451_U879 ( .A1(n4873), .A2(u4_srl_451_n50), .B1(
        fract_denorm[104]), .B2(u4_srl_451_n54), .ZN(u4_srl_451_n836) );
  INV_X1 u4_srl_451_U878 ( .A(u4_srl_451_n836), .ZN(u4_srl_451_n835) );
  AOI221_X1 u4_srl_451_U877 ( .B1(u4_srl_451_n38), .B2(fract_denorm[103]), 
        .C1(u4_srl_451_n45), .C2(fract_denorm[102]), .A(u4_srl_451_n835), .ZN(
        u4_srl_451_n268) );
  OR2_X1 u4_srl_451_U876 ( .A1(u4_srl_451_n186), .A2(u4_srl_451_n64), .ZN(
        u4_srl_451_n834) );
  NOR2_X1 u4_srl_451_U875 ( .A1(u4_srl_451_n268), .A2(u4_srl_451_n834), .ZN(
        u4_N6002) );
  AOI222_X1 u4_srl_451_U874 ( .A1(u4_srl_451_n38), .A2(fract_denorm[104]), 
        .B1(u4_srl_451_n55), .B2(n4873), .C1(u4_srl_451_n45), .C2(
        fract_denorm[103]), .ZN(u4_srl_451_n252) );
  NOR2_X1 u4_srl_451_U873 ( .A1(u4_srl_451_n252), .A2(u4_srl_451_n834), .ZN(
        u4_N6003) );
  NOR2_X1 u4_srl_451_U872 ( .A1(u4_srl_451_n249), .A2(u4_srl_451_n834), .ZN(
        u4_N6004) );
  NOR3_X1 u4_srl_451_U871 ( .A1(u4_srl_451_n63), .A2(u4_srl_451_n243), .A3(
        u4_srl_451_n245), .ZN(u4_srl_451_n380) );
  AND2_X1 u4_srl_451_U870 ( .A1(u4_srl_451_n215), .A2(u4_srl_451_n380), .ZN(
        u4_N6005) );
  AOI22_X1 u4_srl_451_U869 ( .A1(fract_denorm[33]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[32]), .B2(u4_srl_451_n54), .ZN(u4_srl_451_n833) );
  OAI221_X1 u4_srl_451_U868 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n93), .C1(
        u4_srl_451_n44), .C2(u4_srl_451_n92), .A(u4_srl_451_n833), .ZN(
        u4_srl_451_n578) );
  AOI22_X1 u4_srl_451_U867 ( .A1(fract_denorm[29]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[28]), .B2(u4_srl_451_n53), .ZN(u4_srl_451_n832) );
  OAI221_X1 u4_srl_451_U866 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n89), .C1(
        u4_srl_451_n44), .C2(u4_srl_451_n88), .A(u4_srl_451_n832), .ZN(
        u4_srl_451_n659) );
  AOI22_X1 u4_srl_451_U865 ( .A1(fract_denorm[41]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[40]), .B2(u4_srl_451_n53), .ZN(u4_srl_451_n831) );
  OAI221_X1 u4_srl_451_U864 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n101), .C1(
        u4_srl_451_n44), .C2(u4_srl_451_n100), .A(u4_srl_451_n831), .ZN(
        u4_srl_451_n580) );
  AOI22_X1 u4_srl_451_U863 ( .A1(fract_denorm[37]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[36]), .B2(u4_srl_451_n53), .ZN(u4_srl_451_n830) );
  OAI221_X1 u4_srl_451_U862 ( .B1(u4_srl_451_n35), .B2(u4_srl_451_n97), .C1(
        u4_srl_451_n44), .C2(u4_srl_451_n96), .A(u4_srl_451_n830), .ZN(
        u4_srl_451_n577) );
  AOI22_X1 u4_srl_451_U861 ( .A1(u4_srl_451_n24), .A2(u4_srl_451_n580), .B1(
        u4_srl_451_n30), .B2(u4_srl_451_n577), .ZN(u4_srl_451_n829) );
  INV_X1 u4_srl_451_U860 ( .A(u4_srl_451_n829), .ZN(u4_srl_451_n828) );
  AOI221_X1 u4_srl_451_U859 ( .B1(u4_srl_451_n578), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n659), .C2(u4_srl_451_n61), .A(u4_srl_451_n828), .ZN(
        u4_srl_451_n456) );
  INV_X1 u4_srl_451_U858 ( .A(u4_srl_451_n456), .ZN(u4_srl_451_n803) );
  AOI22_X1 u4_srl_451_U857 ( .A1(fract_denorm[97]), .A2(u4_srl_451_n50), .B1(
        fract_denorm[96]), .B2(u4_srl_451_n53), .ZN(u4_srl_451_n827) );
  OAI221_X1 u4_srl_451_U856 ( .B1(u4_srl_451_n35), .B2(u4_srl_451_n157), .C1(
        u4_srl_451_n43), .C2(u4_srl_451_n156), .A(u4_srl_451_n827), .ZN(
        u4_srl_451_n567) );
  AOI22_X1 u4_srl_451_U855 ( .A1(fract_denorm[93]), .A2(u4_srl_451_n48), .B1(
        fract_denorm[92]), .B2(u4_srl_451_n53), .ZN(u4_srl_451_n826) );
  OAI221_X1 u4_srl_451_U854 ( .B1(u4_srl_451_n35), .B2(u4_srl_451_n153), .C1(
        u4_srl_451_n43), .C2(u4_srl_451_n152), .A(u4_srl_451_n826), .ZN(
        u4_srl_451_n562) );
  INV_X1 u4_srl_451_U853 ( .A(u4_srl_451_n268), .ZN(u4_srl_451_n411) );
  AOI22_X1 u4_srl_451_U852 ( .A1(fract_denorm[101]), .A2(u4_srl_451_n50), .B1(
        fract_denorm[100]), .B2(u4_srl_451_n53), .ZN(u4_srl_451_n825) );
  OAI221_X1 u4_srl_451_U851 ( .B1(u4_srl_451_n35), .B2(u4_srl_451_n161), .C1(
        u4_srl_451_n40), .C2(u4_srl_451_n160), .A(u4_srl_451_n825), .ZN(
        u4_srl_451_n566) );
  AOI22_X1 u4_srl_451_U850 ( .A1(u4_srl_451_n24), .A2(u4_srl_451_n411), .B1(
        u4_srl_451_n30), .B2(u4_srl_451_n566), .ZN(u4_srl_451_n824) );
  INV_X1 u4_srl_451_U849 ( .A(u4_srl_451_n824), .ZN(u4_srl_451_n823) );
  AOI221_X1 u4_srl_451_U848 ( .B1(u4_srl_451_n567), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n562), .C2(u4_srl_451_n61), .A(u4_srl_451_n823), .ZN(
        u4_srl_451_n195) );
  AOI22_X1 u4_srl_451_U847 ( .A1(fract_denorm[81]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[80]), .B2(u4_srl_451_n53), .ZN(u4_srl_451_n822) );
  OAI221_X1 u4_srl_451_U846 ( .B1(u4_srl_451_n35), .B2(u4_srl_451_n141), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n140), .A(u4_srl_451_n822), .ZN(
        u4_srl_451_n561) );
  INV_X1 u4_srl_451_U845 ( .A(u4_srl_451_n561), .ZN(u4_srl_451_n702) );
  AOI22_X1 u4_srl_451_U844 ( .A1(fract_denorm[77]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[76]), .B2(u4_srl_451_n53), .ZN(u4_srl_451_n821) );
  OAI221_X1 u4_srl_451_U843 ( .B1(u4_srl_451_n35), .B2(u4_srl_451_n137), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n136), .A(u4_srl_451_n821), .ZN(
        u4_srl_451_n649) );
  INV_X1 u4_srl_451_U842 ( .A(u4_srl_451_n649), .ZN(u4_srl_451_n557) );
  AOI22_X1 u4_srl_451_U841 ( .A1(fract_denorm[89]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[88]), .B2(u4_srl_451_n53), .ZN(u4_srl_451_n820) );
  OAI221_X1 u4_srl_451_U840 ( .B1(u4_srl_451_n35), .B2(u4_srl_451_n149), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n148), .A(u4_srl_451_n820), .ZN(
        u4_srl_451_n563) );
  AOI22_X1 u4_srl_451_U839 ( .A1(fract_denorm[85]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[84]), .B2(u4_srl_451_n53), .ZN(u4_srl_451_n819) );
  OAI221_X1 u4_srl_451_U838 ( .B1(u4_srl_451_n35), .B2(u4_srl_451_n145), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n144), .A(u4_srl_451_n819), .ZN(
        u4_srl_451_n560) );
  AOI22_X1 u4_srl_451_U837 ( .A1(u4_srl_451_n24), .A2(u4_srl_451_n563), .B1(
        u4_srl_451_n29), .B2(u4_srl_451_n560), .ZN(u4_srl_451_n818) );
  OAI221_X1 u4_srl_451_U836 ( .B1(u4_srl_451_n702), .B2(u4_srl_451_n19), .C1(
        u4_srl_451_n557), .C2(u4_srl_451_n64), .A(u4_srl_451_n818), .ZN(
        u4_srl_451_n376) );
  INV_X1 u4_srl_451_U835 ( .A(u4_srl_451_n376), .ZN(u4_srl_451_n302) );
  OAI22_X1 u4_srl_451_U834 ( .A1(u4_srl_451_n195), .A2(u4_srl_451_n247), .B1(
        u4_srl_451_n302), .B2(u4_srl_451_n243), .ZN(u4_srl_451_n241) );
  AOI22_X1 u4_srl_451_U833 ( .A1(fract_denorm[65]), .A2(u4_srl_451_n49), .B1(
        fract_denorm[64]), .B2(u4_srl_451_n53), .ZN(u4_srl_451_n817) );
  OAI221_X1 u4_srl_451_U832 ( .B1(u4_srl_451_n35), .B2(u4_srl_451_n125), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n124), .A(u4_srl_451_n817), .ZN(
        u4_srl_451_n573) );
  AOI22_X1 u4_srl_451_U831 ( .A1(fract_denorm[61]), .A2(u4_srl_451_n49), .B1(
        fract_denorm[60]), .B2(u4_srl_451_n53), .ZN(u4_srl_451_n816) );
  OAI221_X1 u4_srl_451_U830 ( .B1(u4_srl_451_n35), .B2(u4_srl_451_n121), .C1(
        u4_srl_451_n41), .C2(u4_srl_451_n120), .A(u4_srl_451_n816), .ZN(
        u4_srl_451_n568) );
  AOI22_X1 u4_srl_451_U829 ( .A1(fract_denorm[73]), .A2(u4_srl_451_n49), .B1(
        fract_denorm[72]), .B2(u4_srl_451_n52), .ZN(u4_srl_451_n815) );
  OAI221_X1 u4_srl_451_U828 ( .B1(u4_srl_451_n35), .B2(u4_srl_451_n133), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n132), .A(u4_srl_451_n815), .ZN(
        u4_srl_451_n650) );
  AOI22_X1 u4_srl_451_U827 ( .A1(fract_denorm[69]), .A2(u4_srl_451_n49), .B1(
        fract_denorm[68]), .B2(u4_srl_451_n52), .ZN(u4_srl_451_n814) );
  OAI221_X1 u4_srl_451_U826 ( .B1(u4_srl_451_n34), .B2(u4_srl_451_n129), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n128), .A(u4_srl_451_n814), .ZN(
        u4_srl_451_n572) );
  AOI22_X1 u4_srl_451_U825 ( .A1(u4_srl_451_n24), .A2(u4_srl_451_n650), .B1(
        u4_srl_451_n30), .B2(u4_srl_451_n572), .ZN(u4_srl_451_n813) );
  INV_X1 u4_srl_451_U824 ( .A(u4_srl_451_n813), .ZN(u4_srl_451_n812) );
  AOI221_X1 u4_srl_451_U823 ( .B1(u4_srl_451_n573), .B2(u4_srl_451_n18), .C1(
        u4_srl_451_n568), .C2(u4_srl_451_n62), .A(u4_srl_451_n812), .ZN(
        u4_srl_451_n303) );
  AOI22_X1 u4_srl_451_U822 ( .A1(fract_denorm[49]), .A2(u4_srl_451_n49), .B1(
        fract_denorm[48]), .B2(u4_srl_451_n52), .ZN(u4_srl_451_n811) );
  OAI221_X1 u4_srl_451_U821 ( .B1(u4_srl_451_n34), .B2(u4_srl_451_n109), .C1(
        u4_srl_451_n43), .C2(u4_srl_451_n108), .A(u4_srl_451_n811), .ZN(
        u4_srl_451_n584) );
  AOI22_X1 u4_srl_451_U820 ( .A1(fract_denorm[45]), .A2(u4_srl_451_n49), .B1(
        fract_denorm[44]), .B2(u4_srl_451_n52), .ZN(u4_srl_451_n810) );
  OAI221_X1 u4_srl_451_U819 ( .B1(u4_srl_451_n34), .B2(u4_srl_451_n105), .C1(
        u4_srl_451_n43), .C2(u4_srl_451_n104), .A(u4_srl_451_n810), .ZN(
        u4_srl_451_n579) );
  AOI22_X1 u4_srl_451_U818 ( .A1(fract_denorm[57]), .A2(u4_srl_451_n49), .B1(
        fract_denorm[56]), .B2(u4_srl_451_n52), .ZN(u4_srl_451_n809) );
  OAI221_X1 u4_srl_451_U817 ( .B1(u4_srl_451_n34), .B2(u4_srl_451_n117), .C1(
        u4_srl_451_n43), .C2(u4_srl_451_n116), .A(u4_srl_451_n809), .ZN(
        u4_srl_451_n569) );
  AOI22_X1 u4_srl_451_U816 ( .A1(fract_denorm[53]), .A2(u4_srl_451_n49), .B1(
        fract_denorm[52]), .B2(u4_srl_451_n52), .ZN(u4_srl_451_n808) );
  OAI221_X1 u4_srl_451_U815 ( .B1(u4_srl_451_n34), .B2(u4_srl_451_n113), .C1(
        u4_srl_451_n43), .C2(u4_srl_451_n112), .A(u4_srl_451_n808), .ZN(
        u4_srl_451_n583) );
  AOI22_X1 u4_srl_451_U814 ( .A1(u4_srl_451_n24), .A2(u4_srl_451_n569), .B1(
        u4_srl_451_n30), .B2(u4_srl_451_n583), .ZN(u4_srl_451_n807) );
  INV_X1 u4_srl_451_U813 ( .A(u4_srl_451_n807), .ZN(u4_srl_451_n806) );
  AOI221_X1 u4_srl_451_U812 ( .B1(u4_srl_451_n584), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n579), .C2(u4_srl_451_n62), .A(u4_srl_451_n806), .ZN(
        u4_srl_451_n378) );
  OAI22_X1 u4_srl_451_U811 ( .A1(u4_srl_451_n303), .A2(u4_srl_451_n182), .B1(
        u4_srl_451_n378), .B2(u4_srl_451_n184), .ZN(u4_srl_451_n804) );
  AOI221_X1 u4_srl_451_U810 ( .B1(u4_srl_451_n176), .B2(u4_srl_451_n803), .C1(
        u4_srl_451_n241), .C2(u4_srl_451_n179), .A(u4_srl_451_n804), .ZN(
        u4_srl_451_n795) );
  NOR2_X1 u4_srl_451_U809 ( .A1(u4_srl_451_n243), .A2(u4_srl_451_n179), .ZN(
        u4_srl_451_n798) );
  AOI22_X1 u4_srl_451_U808 ( .A1(fract_denorm[17]), .A2(u4_srl_451_n49), .B1(
        fract_denorm[16]), .B2(u4_srl_451_n52), .ZN(u4_srl_451_n802) );
  OAI221_X1 u4_srl_451_U807 ( .B1(u4_srl_451_n34), .B2(u4_srl_451_n78), .C1(
        u4_srl_451_n43), .C2(u4_srl_451_n77), .A(u4_srl_451_n802), .ZN(
        u4_srl_451_n258) );
  AOI22_X1 u4_srl_451_U806 ( .A1(fract_denorm[13]), .A2(u4_srl_451_n49), .B1(
        fract_denorm[12]), .B2(u4_srl_451_n52), .ZN(u4_srl_451_n801) );
  OAI221_X1 u4_srl_451_U805 ( .B1(u4_srl_451_n34), .B2(u4_srl_451_n74), .C1(
        u4_srl_451_n43), .C2(u4_srl_451_n73), .A(u4_srl_451_n801), .ZN(
        u4_srl_451_n262) );
  AOI22_X1 u4_srl_451_U804 ( .A1(fract_denorm[21]), .A2(u4_srl_451_n49), .B1(
        fract_denorm[20]), .B2(u4_srl_451_n52), .ZN(u4_srl_451_n800) );
  OAI221_X1 u4_srl_451_U803 ( .B1(u4_srl_451_n34), .B2(u4_srl_451_n82), .C1(
        u4_srl_451_n43), .C2(u4_srl_451_n81), .A(u4_srl_451_n800), .ZN(
        u4_srl_451_n257) );
  INV_X1 u4_srl_451_U802 ( .A(u4_srl_451_n257), .ZN(u4_srl_451_n657) );
  OAI22_X1 u4_srl_451_U801 ( .A1(u4_srl_451_n87), .A2(u4_srl_451_n1), .B1(
        u4_srl_451_n58), .B2(u4_srl_451_n86), .ZN(u4_srl_451_n799) );
  AOI221_X1 u4_srl_451_U800 ( .B1(fract_denorm[23]), .B2(u4_srl_451_n38), .C1(
        fract_denorm[22]), .C2(u4_srl_451_n45), .A(u4_srl_451_n799), .ZN(
        u4_srl_451_n575) );
  OAI22_X1 u4_srl_451_U799 ( .A1(u4_srl_451_n657), .A2(u4_srl_451_n173), .B1(
        u4_srl_451_n575), .B2(u4_srl_451_n175), .ZN(u4_srl_451_n797) );
  AOI221_X1 u4_srl_451_U798 ( .B1(u4_srl_451_n167), .B2(u4_srl_451_n258), .C1(
        u4_srl_451_n169), .C2(u4_srl_451_n262), .A(u4_srl_451_n797), .ZN(
        u4_srl_451_n796) );
  AOI21_X1 u4_srl_451_U797 ( .B1(u4_srl_451_n795), .B2(u4_srl_451_n796), .A(
        u4_shift_right[8]), .ZN(u4_N5910) );
  AOI22_X1 u4_srl_451_U796 ( .A1(fract_denorm[34]), .A2(u4_srl_451_n49), .B1(
        fract_denorm[33]), .B2(u4_srl_451_n52), .ZN(u4_srl_451_n794) );
  OAI221_X1 u4_srl_451_U795 ( .B1(u4_srl_451_n34), .B2(u4_srl_451_n94), .C1(
        u4_srl_451_n43), .C2(u4_srl_451_n93), .A(u4_srl_451_n794), .ZN(
        u4_srl_451_n547) );
  AOI22_X1 u4_srl_451_U794 ( .A1(fract_denorm[30]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[29]), .B2(u4_srl_451_n52), .ZN(u4_srl_451_n793) );
  OAI221_X1 u4_srl_451_U793 ( .B1(u4_srl_451_n34), .B2(u4_srl_451_n90), .C1(
        u4_srl_451_n43), .C2(u4_srl_451_n89), .A(u4_srl_451_n793), .ZN(
        u4_srl_451_n642) );
  AOI22_X1 u4_srl_451_U792 ( .A1(fract_denorm[42]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[41]), .B2(u4_srl_451_n51), .ZN(u4_srl_451_n792) );
  OAI221_X1 u4_srl_451_U791 ( .B1(u4_srl_451_n33), .B2(u4_srl_451_n102), .C1(
        u4_srl_451_n43), .C2(u4_srl_451_n101), .A(u4_srl_451_n792), .ZN(
        u4_srl_451_n549) );
  AOI22_X1 u4_srl_451_U790 ( .A1(fract_denorm[38]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[37]), .B2(u4_srl_451_n51), .ZN(u4_srl_451_n791) );
  OAI221_X1 u4_srl_451_U789 ( .B1(u4_srl_451_n33), .B2(u4_srl_451_n98), .C1(
        u4_srl_451_n43), .C2(u4_srl_451_n97), .A(u4_srl_451_n791), .ZN(
        u4_srl_451_n546) );
  AOI22_X1 u4_srl_451_U788 ( .A1(u4_srl_451_n23), .A2(u4_srl_451_n549), .B1(
        u4_srl_451_n29), .B2(u4_srl_451_n546), .ZN(u4_srl_451_n790) );
  INV_X1 u4_srl_451_U787 ( .A(u4_srl_451_n790), .ZN(u4_srl_451_n789) );
  AOI221_X1 u4_srl_451_U786 ( .B1(u4_srl_451_n547), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n642), .C2(u4_srl_451_n62), .A(u4_srl_451_n789), .ZN(
        u4_srl_451_n453) );
  INV_X1 u4_srl_451_U785 ( .A(u4_srl_451_n453), .ZN(u4_srl_451_n765) );
  AOI22_X1 u4_srl_451_U784 ( .A1(fract_denorm[98]), .A2(u4_srl_451_n49), .B1(
        fract_denorm[97]), .B2(u4_srl_451_n51), .ZN(u4_srl_451_n788) );
  OAI221_X1 u4_srl_451_U783 ( .B1(u4_srl_451_n33), .B2(u4_srl_451_n158), .C1(
        u4_srl_451_n41), .C2(u4_srl_451_n157), .A(u4_srl_451_n788), .ZN(
        u4_srl_451_n536) );
  AOI22_X1 u4_srl_451_U782 ( .A1(fract_denorm[94]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[93]), .B2(u4_srl_451_n51), .ZN(u4_srl_451_n787) );
  OAI221_X1 u4_srl_451_U781 ( .B1(u4_srl_451_n33), .B2(u4_srl_451_n154), .C1(
        u4_srl_451_n40), .C2(u4_srl_451_n153), .A(u4_srl_451_n787), .ZN(
        u4_srl_451_n531) );
  INV_X1 u4_srl_451_U780 ( .A(u4_srl_451_n252), .ZN(u4_srl_451_n408) );
  AOI22_X1 u4_srl_451_U779 ( .A1(fract_denorm[102]), .A2(u4_srl_451_n48), .B1(
        fract_denorm[101]), .B2(u4_srl_451_n51), .ZN(u4_srl_451_n786) );
  OAI221_X1 u4_srl_451_U778 ( .B1(u4_srl_451_n33), .B2(u4_srl_451_n162), .C1(
        u4_srl_451_n40), .C2(u4_srl_451_n161), .A(u4_srl_451_n786), .ZN(
        u4_srl_451_n535) );
  AOI22_X1 u4_srl_451_U777 ( .A1(u4_srl_451_n23), .A2(u4_srl_451_n408), .B1(
        u4_srl_451_n29), .B2(u4_srl_451_n535), .ZN(u4_srl_451_n785) );
  INV_X1 u4_srl_451_U776 ( .A(u4_srl_451_n785), .ZN(u4_srl_451_n784) );
  AOI221_X1 u4_srl_451_U775 ( .B1(u4_srl_451_n536), .B2(u4_srl_451_n18), .C1(
        u4_srl_451_n531), .C2(u4_srl_451_n62), .A(u4_srl_451_n784), .ZN(
        u4_srl_451_n194) );
  AOI22_X1 u4_srl_451_U774 ( .A1(fract_denorm[82]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[81]), .B2(u4_srl_451_n51), .ZN(u4_srl_451_n783) );
  OAI221_X1 u4_srl_451_U773 ( .B1(u4_srl_451_n33), .B2(u4_srl_451_n142), .C1(
        u4_srl_451_n40), .C2(u4_srl_451_n141), .A(u4_srl_451_n783), .ZN(
        u4_srl_451_n530) );
  INV_X1 u4_srl_451_U772 ( .A(u4_srl_451_n530), .ZN(u4_srl_451_n689) );
  AOI22_X1 u4_srl_451_U771 ( .A1(fract_denorm[78]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[77]), .B2(u4_srl_451_n51), .ZN(u4_srl_451_n782) );
  OAI221_X1 u4_srl_451_U770 ( .B1(u4_srl_451_n33), .B2(u4_srl_451_n138), .C1(
        u4_srl_451_n41), .C2(u4_srl_451_n137), .A(u4_srl_451_n782), .ZN(
        u4_srl_451_n632) );
  INV_X1 u4_srl_451_U769 ( .A(u4_srl_451_n632), .ZN(u4_srl_451_n526) );
  AOI22_X1 u4_srl_451_U768 ( .A1(fract_denorm[90]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[89]), .B2(u4_srl_451_n51), .ZN(u4_srl_451_n781) );
  OAI221_X1 u4_srl_451_U767 ( .B1(u4_srl_451_n33), .B2(u4_srl_451_n150), .C1(
        u4_srl_451_n40), .C2(u4_srl_451_n149), .A(u4_srl_451_n781), .ZN(
        u4_srl_451_n532) );
  AOI22_X1 u4_srl_451_U766 ( .A1(fract_denorm[86]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[85]), .B2(u4_srl_451_n51), .ZN(u4_srl_451_n780) );
  OAI221_X1 u4_srl_451_U765 ( .B1(u4_srl_451_n33), .B2(u4_srl_451_n146), .C1(
        u4_srl_451_n41), .C2(u4_srl_451_n145), .A(u4_srl_451_n780), .ZN(
        u4_srl_451_n529) );
  AOI22_X1 u4_srl_451_U764 ( .A1(u4_srl_451_n23), .A2(u4_srl_451_n532), .B1(
        u4_srl_451_n29), .B2(u4_srl_451_n529), .ZN(u4_srl_451_n779) );
  OAI221_X1 u4_srl_451_U763 ( .B1(u4_srl_451_n689), .B2(u4_srl_451_n19), .C1(
        u4_srl_451_n526), .C2(u4_srl_451_n64), .A(u4_srl_451_n779), .ZN(
        u4_srl_451_n371) );
  INV_X1 u4_srl_451_U762 ( .A(u4_srl_451_n371), .ZN(u4_srl_451_n300) );
  OAI22_X1 u4_srl_451_U761 ( .A1(u4_srl_451_n194), .A2(u4_srl_451_n247), .B1(
        u4_srl_451_n300), .B2(u4_srl_451_n243), .ZN(u4_srl_451_n240) );
  AOI22_X1 u4_srl_451_U760 ( .A1(fract_denorm[66]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[65]), .B2(u4_srl_451_n51), .ZN(u4_srl_451_n778) );
  OAI221_X1 u4_srl_451_U759 ( .B1(u4_srl_451_n33), .B2(u4_srl_451_n126), .C1(
        u4_srl_451_n41), .C2(u4_srl_451_n125), .A(u4_srl_451_n778), .ZN(
        u4_srl_451_n542) );
  AOI22_X1 u4_srl_451_U758 ( .A1(fract_denorm[62]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[61]), .B2(u4_srl_451_n51), .ZN(u4_srl_451_n777) );
  OAI221_X1 u4_srl_451_U757 ( .B1(u4_srl_451_n33), .B2(u4_srl_451_n122), .C1(
        u4_srl_451_n43), .C2(u4_srl_451_n121), .A(u4_srl_451_n777), .ZN(
        u4_srl_451_n537) );
  AOI22_X1 u4_srl_451_U756 ( .A1(fract_denorm[74]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[73]), .B2(u4_srl_451_n51), .ZN(u4_srl_451_n776) );
  OAI221_X1 u4_srl_451_U755 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n134), .C1(
        u4_srl_451_n43), .C2(u4_srl_451_n133), .A(u4_srl_451_n776), .ZN(
        u4_srl_451_n633) );
  AOI22_X1 u4_srl_451_U754 ( .A1(fract_denorm[70]), .A2(u4_srl_451_n48), .B1(
        fract_denorm[69]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n775) );
  OAI221_X1 u4_srl_451_U753 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n130), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n129), .A(u4_srl_451_n775), .ZN(
        u4_srl_451_n541) );
  AOI22_X1 u4_srl_451_U752 ( .A1(u4_srl_451_n23), .A2(u4_srl_451_n633), .B1(
        u4_srl_451_n29), .B2(u4_srl_451_n541), .ZN(u4_srl_451_n774) );
  INV_X1 u4_srl_451_U751 ( .A(u4_srl_451_n774), .ZN(u4_srl_451_n773) );
  AOI221_X1 u4_srl_451_U750 ( .B1(u4_srl_451_n542), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n537), .C2(u4_srl_451_n62), .A(u4_srl_451_n773), .ZN(
        u4_srl_451_n301) );
  AOI22_X1 u4_srl_451_U749 ( .A1(fract_denorm[50]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[49]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n772) );
  OAI221_X1 u4_srl_451_U748 ( .B1(u4_srl_451_n32), .B2(u4_srl_451_n110), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n109), .A(u4_srl_451_n772), .ZN(
        u4_srl_451_n553) );
  AOI22_X1 u4_srl_451_U747 ( .A1(fract_denorm[46]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[45]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n771) );
  OAI221_X1 u4_srl_451_U746 ( .B1(u4_srl_451_n32), .B2(u4_srl_451_n106), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n105), .A(u4_srl_451_n771), .ZN(
        u4_srl_451_n548) );
  AOI22_X1 u4_srl_451_U745 ( .A1(fract_denorm[58]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[57]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n770) );
  OAI221_X1 u4_srl_451_U744 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n118), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n117), .A(u4_srl_451_n770), .ZN(
        u4_srl_451_n538) );
  AOI22_X1 u4_srl_451_U743 ( .A1(fract_denorm[54]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[53]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n769) );
  OAI221_X1 u4_srl_451_U742 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n114), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n113), .A(u4_srl_451_n769), .ZN(
        u4_srl_451_n552) );
  AOI22_X1 u4_srl_451_U741 ( .A1(u4_srl_451_n23), .A2(u4_srl_451_n538), .B1(
        u4_srl_451_n29), .B2(u4_srl_451_n552), .ZN(u4_srl_451_n768) );
  INV_X1 u4_srl_451_U740 ( .A(u4_srl_451_n768), .ZN(u4_srl_451_n767) );
  AOI221_X1 u4_srl_451_U739 ( .B1(u4_srl_451_n553), .B2(u4_srl_451_n18), .C1(
        u4_srl_451_n548), .C2(u4_srl_451_n62), .A(u4_srl_451_n767), .ZN(
        u4_srl_451_n373) );
  OAI22_X1 u4_srl_451_U738 ( .A1(u4_srl_451_n301), .A2(u4_srl_451_n182), .B1(
        u4_srl_451_n373), .B2(u4_srl_451_n184), .ZN(u4_srl_451_n766) );
  AOI221_X1 u4_srl_451_U737 ( .B1(u4_srl_451_n176), .B2(u4_srl_451_n765), .C1(
        u4_srl_451_n240), .C2(u4_srl_451_n179), .A(u4_srl_451_n766), .ZN(
        u4_srl_451_n758) );
  AOI22_X1 u4_srl_451_U736 ( .A1(fract_denorm[18]), .A2(u4_srl_451_n48), .B1(
        fract_denorm[17]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n764) );
  OAI221_X1 u4_srl_451_U735 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n79), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n78), .A(u4_srl_451_n764), .ZN(
        u4_srl_451_n226) );
  AOI22_X1 u4_srl_451_U734 ( .A1(fract_denorm[14]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[13]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n763) );
  OAI221_X1 u4_srl_451_U733 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n75), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n74), .A(u4_srl_451_n763), .ZN(
        u4_srl_451_n230) );
  OAI22_X1 u4_srl_451_U732 ( .A1(u4_srl_451_n84), .A2(u4_srl_451_n1), .B1(
        u4_srl_451_n83), .B2(u4_srl_451_n58), .ZN(u4_srl_451_n762) );
  AOI221_X1 u4_srl_451_U731 ( .B1(u4_srl_451_n38), .B2(fract_denorm[20]), .C1(
        u4_srl_451_n45), .C2(fract_denorm[19]), .A(u4_srl_451_n762), .ZN(
        u4_srl_451_n640) );
  OAI22_X1 u4_srl_451_U730 ( .A1(u4_srl_451_n88), .A2(u4_srl_451_n1), .B1(
        u4_srl_451_n87), .B2(u4_srl_451_n58), .ZN(u4_srl_451_n761) );
  AOI221_X1 u4_srl_451_U729 ( .B1(fract_denorm[24]), .B2(u4_srl_451_n38), .C1(
        fract_denorm[23]), .C2(u4_srl_451_n45), .A(u4_srl_451_n761), .ZN(
        u4_srl_451_n544) );
  OAI22_X1 u4_srl_451_U728 ( .A1(u4_srl_451_n640), .A2(u4_srl_451_n173), .B1(
        u4_srl_451_n544), .B2(u4_srl_451_n175), .ZN(u4_srl_451_n760) );
  AOI221_X1 u4_srl_451_U727 ( .B1(u4_srl_451_n167), .B2(u4_srl_451_n226), .C1(
        u4_srl_451_n169), .C2(u4_srl_451_n230), .A(u4_srl_451_n760), .ZN(
        u4_srl_451_n759) );
  AOI21_X1 u4_srl_451_U726 ( .B1(u4_srl_451_n758), .B2(u4_srl_451_n759), .A(
        u4_shift_right[8]), .ZN(u4_N5911) );
  AOI22_X1 u4_srl_451_U725 ( .A1(u4_srl_451_n23), .A2(u4_srl_451_n518), .B1(
        u4_srl_451_n29), .B2(u4_srl_451_n514), .ZN(u4_srl_451_n757) );
  INV_X1 u4_srl_451_U724 ( .A(u4_srl_451_n757), .ZN(u4_srl_451_n756) );
  AOI221_X1 u4_srl_451_U723 ( .B1(u4_srl_451_n515), .B2(u4_srl_451_n18), .C1(
        u4_srl_451_n516), .C2(u4_srl_451_n62), .A(u4_srl_451_n756), .ZN(
        u4_srl_451_n450) );
  INV_X1 u4_srl_451_U722 ( .A(u4_srl_451_n450), .ZN(u4_srl_451_n746) );
  INV_X1 u4_srl_451_U721 ( .A(u4_srl_451_n504), .ZN(u4_srl_451_n754) );
  INV_X1 u4_srl_451_U720 ( .A(u4_srl_451_n609), .ZN(u4_srl_451_n500) );
  AOI22_X1 u4_srl_451_U719 ( .A1(u4_srl_451_n23), .A2(u4_srl_451_n385), .B1(
        u4_srl_451_n29), .B2(u4_srl_451_n503), .ZN(u4_srl_451_n755) );
  OAI221_X1 u4_srl_451_U718 ( .B1(u4_srl_451_n754), .B2(u4_srl_451_n19), .C1(
        u4_srl_451_n500), .C2(u4_srl_451_n64), .A(u4_srl_451_n755), .ZN(
        u4_srl_451_n365) );
  INV_X1 u4_srl_451_U717 ( .A(u4_srl_451_n365), .ZN(u4_srl_451_n193) );
  INV_X1 u4_srl_451_U716 ( .A(u4_srl_451_n605), .ZN(u4_srl_451_n495) );
  AOI22_X1 u4_srl_451_U715 ( .A1(u4_srl_451_n23), .A2(u4_srl_451_n610), .B1(
        u4_srl_451_n29), .B2(u4_srl_451_n498), .ZN(u4_srl_451_n753) );
  OAI221_X1 u4_srl_451_U714 ( .B1(u4_srl_451_n752), .B2(u4_srl_451_n19), .C1(
        u4_srl_451_n495), .C2(u4_srl_451_n64), .A(u4_srl_451_n753), .ZN(
        u4_srl_451_n366) );
  INV_X1 u4_srl_451_U713 ( .A(u4_srl_451_n366), .ZN(u4_srl_451_n284) );
  OAI22_X1 u4_srl_451_U712 ( .A1(u4_srl_451_n193), .A2(u4_srl_451_n247), .B1(
        u4_srl_451_n284), .B2(u4_srl_451_n243), .ZN(u4_srl_451_n239) );
  INV_X1 u4_srl_451_U711 ( .A(u4_srl_451_n613), .ZN(u4_srl_451_n505) );
  AOI22_X1 u4_srl_451_U710 ( .A1(u4_srl_451_n23), .A2(u4_srl_451_n606), .B1(
        u4_srl_451_n29), .B2(u4_srl_451_n508), .ZN(u4_srl_451_n751) );
  OAI221_X1 u4_srl_451_U709 ( .B1(u4_srl_451_n750), .B2(u4_srl_451_n19), .C1(
        u4_srl_451_n505), .C2(u4_srl_451_n64), .A(u4_srl_451_n751), .ZN(
        u4_srl_451_n452) );
  INV_X1 u4_srl_451_U708 ( .A(u4_srl_451_n452), .ZN(u4_srl_451_n285) );
  AOI22_X1 u4_srl_451_U707 ( .A1(u4_srl_451_n23), .A2(u4_srl_451_n510), .B1(
        u4_srl_451_n29), .B2(u4_srl_451_n521), .ZN(u4_srl_451_n749) );
  INV_X1 u4_srl_451_U706 ( .A(u4_srl_451_n749), .ZN(u4_srl_451_n748) );
  AOI221_X1 u4_srl_451_U705 ( .B1(u4_srl_451_n522), .B2(u4_srl_451_n18), .C1(
        u4_srl_451_n517), .C2(u4_srl_451_n62), .A(u4_srl_451_n748), .ZN(
        u4_srl_451_n368) );
  OAI22_X1 u4_srl_451_U704 ( .A1(u4_srl_451_n285), .A2(u4_srl_451_n182), .B1(
        u4_srl_451_n368), .B2(u4_srl_451_n184), .ZN(u4_srl_451_n747) );
  AOI221_X1 u4_srl_451_U703 ( .B1(u4_srl_451_n176), .B2(u4_srl_451_n746), .C1(
        u4_srl_451_n239), .C2(u4_srl_451_n179), .A(u4_srl_451_n747), .ZN(
        u4_srl_451_n742) );
  INV_X1 u4_srl_451_U702 ( .A(u4_srl_451_n745), .ZN(u4_srl_451_n512) );
  OAI22_X1 u4_srl_451_U701 ( .A1(u4_srl_451_n202), .A2(u4_srl_451_n173), .B1(
        u4_srl_451_n512), .B2(u4_srl_451_n175), .ZN(u4_srl_451_n744) );
  AOI221_X1 u4_srl_451_U700 ( .B1(u4_srl_451_n167), .B2(u4_srl_451_n332), .C1(
        u4_srl_451_n169), .C2(u4_srl_451_n198), .A(u4_srl_451_n744), .ZN(
        u4_srl_451_n743) );
  AOI21_X1 u4_srl_451_U699 ( .B1(u4_srl_451_n742), .B2(u4_srl_451_n743), .A(
        u4_shift_right[8]), .ZN(u4_N5912) );
  AOI22_X1 u4_srl_451_U698 ( .A1(fract_denorm[36]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[35]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n741) );
  OAI221_X1 u4_srl_451_U697 ( .B1(u4_srl_451_n32), .B2(u4_srl_451_n96), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n95), .A(u4_srl_451_n741), .ZN(
        u4_srl_451_n485) );
  AOI22_X1 u4_srl_451_U696 ( .A1(fract_denorm[32]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[31]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n740) );
  OAI221_X1 u4_srl_451_U695 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n92), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n91), .A(u4_srl_451_n740), .ZN(
        u4_srl_451_n486) );
  AOI22_X1 u4_srl_451_U694 ( .A1(fract_denorm[44]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[43]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n739) );
  OAI221_X1 u4_srl_451_U693 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n104), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n103), .A(u4_srl_451_n739), .ZN(
        u4_srl_451_n488) );
  AOI22_X1 u4_srl_451_U692 ( .A1(fract_denorm[40]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[39]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n738) );
  OAI221_X1 u4_srl_451_U691 ( .B1(u4_srl_451_n32), .B2(u4_srl_451_n100), .C1(
        u4_srl_451_n42), .C2(u4_srl_451_n99), .A(u4_srl_451_n738), .ZN(
        u4_srl_451_n484) );
  AOI22_X1 u4_srl_451_U690 ( .A1(u4_srl_451_n23), .A2(u4_srl_451_n488), .B1(
        u4_srl_451_n28), .B2(u4_srl_451_n484), .ZN(u4_srl_451_n737) );
  INV_X1 u4_srl_451_U689 ( .A(u4_srl_451_n737), .ZN(u4_srl_451_n736) );
  AOI221_X1 u4_srl_451_U688 ( .B1(u4_srl_451_n485), .B2(u4_srl_451_n18), .C1(
        u4_srl_451_n486), .C2(u4_srl_451_n62), .A(u4_srl_451_n736), .ZN(
        u4_srl_451_n447) );
  INV_X1 u4_srl_451_U687 ( .A(u4_srl_451_n447), .ZN(u4_srl_451_n713) );
  AOI22_X1 u4_srl_451_U686 ( .A1(fract_denorm[96]), .A2(u4_srl_451_n48), .B1(
        fract_denorm[95]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n735) );
  OAI221_X1 u4_srl_451_U685 ( .B1(u4_srl_451_n32), .B2(u4_srl_451_n156), .C1(
        u4_srl_451_n41), .C2(u4_srl_451_n155), .A(u4_srl_451_n735), .ZN(
        u4_srl_451_n469) );
  AOI22_X1 u4_srl_451_U684 ( .A1(fract_denorm[100]), .A2(u4_srl_451_n48), .B1(
        fract_denorm[99]), .B2(u4_srl_451_n52), .ZN(u4_srl_451_n734) );
  OAI221_X1 u4_srl_451_U683 ( .B1(u4_srl_451_n32), .B2(u4_srl_451_n160), .C1(
        u4_srl_451_n41), .C2(u4_srl_451_n159), .A(u4_srl_451_n734), .ZN(
        u4_srl_451_n474) );
  AOI222_X1 u4_srl_451_U682 ( .A1(u4_srl_451_n469), .A2(u4_srl_451_n60), .B1(
        u4_srl_451_n474), .B2(u4_srl_451_n17), .C1(u4_srl_451_n732), .C2(
        u4_srl_451_n733), .ZN(u4_srl_451_n192) );
  AOI22_X1 u4_srl_451_U681 ( .A1(fract_denorm[84]), .A2(u4_srl_451_n48), .B1(
        fract_denorm[83]), .B2(u4_srl_451_n52), .ZN(u4_srl_451_n731) );
  OAI221_X1 u4_srl_451_U680 ( .B1(u4_srl_451_n32), .B2(u4_srl_451_n144), .C1(
        u4_srl_451_n41), .C2(u4_srl_451_n143), .A(u4_srl_451_n731), .ZN(
        u4_srl_451_n467) );
  INV_X1 u4_srl_451_U679 ( .A(u4_srl_451_n467), .ZN(u4_srl_451_n667) );
  AOI22_X1 u4_srl_451_U678 ( .A1(fract_denorm[80]), .A2(u4_srl_451_n48), .B1(
        fract_denorm[79]), .B2(u4_srl_451_n52), .ZN(u4_srl_451_n730) );
  OAI221_X1 u4_srl_451_U677 ( .B1(u4_srl_451_n32), .B2(u4_srl_451_n140), .C1(
        u4_srl_451_n41), .C2(u4_srl_451_n139), .A(u4_srl_451_n730), .ZN(
        u4_srl_451_n591) );
  INV_X1 u4_srl_451_U676 ( .A(u4_srl_451_n591), .ZN(u4_srl_451_n463) );
  AOI22_X1 u4_srl_451_U675 ( .A1(fract_denorm[92]), .A2(u4_srl_451_n48), .B1(
        fract_denorm[91]), .B2(u4_srl_451_n52), .ZN(u4_srl_451_n729) );
  OAI221_X1 u4_srl_451_U674 ( .B1(u4_srl_451_n32), .B2(u4_srl_451_n152), .C1(
        u4_srl_451_n41), .C2(u4_srl_451_n151), .A(u4_srl_451_n729), .ZN(
        u4_srl_451_n470) );
  AOI22_X1 u4_srl_451_U673 ( .A1(fract_denorm[88]), .A2(u4_srl_451_n48), .B1(
        fract_denorm[87]), .B2(u4_srl_451_n52), .ZN(u4_srl_451_n728) );
  OAI221_X1 u4_srl_451_U672 ( .B1(u4_srl_451_n32), .B2(u4_srl_451_n148), .C1(
        u4_srl_451_n41), .C2(u4_srl_451_n147), .A(u4_srl_451_n728), .ZN(
        u4_srl_451_n466) );
  AOI22_X1 u4_srl_451_U671 ( .A1(u4_srl_451_n23), .A2(u4_srl_451_n470), .B1(
        u4_srl_451_n28), .B2(u4_srl_451_n466), .ZN(u4_srl_451_n727) );
  OAI221_X1 u4_srl_451_U670 ( .B1(u4_srl_451_n667), .B2(u4_srl_451_n19), .C1(
        u4_srl_451_n463), .C2(u4_srl_451_n64), .A(u4_srl_451_n727), .ZN(
        u4_srl_451_n361) );
  INV_X1 u4_srl_451_U669 ( .A(u4_srl_451_n361), .ZN(u4_srl_451_n282) );
  OAI22_X1 u4_srl_451_U668 ( .A1(u4_srl_451_n192), .A2(u4_srl_451_n247), .B1(
        u4_srl_451_n282), .B2(u4_srl_451_n243), .ZN(u4_srl_451_n238) );
  AOI22_X1 u4_srl_451_U667 ( .A1(fract_denorm[68]), .A2(u4_srl_451_n48), .B1(
        fract_denorm[67]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n726) );
  OAI221_X1 u4_srl_451_U666 ( .B1(u4_srl_451_n32), .B2(u4_srl_451_n128), .C1(
        u4_srl_451_n41), .C2(u4_srl_451_n127), .A(u4_srl_451_n726), .ZN(
        u4_srl_451_n480) );
  AOI22_X1 u4_srl_451_U665 ( .A1(fract_denorm[64]), .A2(u4_srl_451_n48), .B1(
        fract_denorm[63]), .B2(u4_srl_451_n52), .ZN(u4_srl_451_n725) );
  OAI221_X1 u4_srl_451_U664 ( .B1(u4_srl_451_n32), .B2(u4_srl_451_n124), .C1(
        u4_srl_451_n41), .C2(u4_srl_451_n123), .A(u4_srl_451_n725), .ZN(
        u4_srl_451_n475) );
  AOI22_X1 u4_srl_451_U663 ( .A1(fract_denorm[76]), .A2(u4_srl_451_n48), .B1(
        fract_denorm[75]), .B2(u4_srl_451_n52), .ZN(u4_srl_451_n724) );
  OAI221_X1 u4_srl_451_U662 ( .B1(u4_srl_451_n32), .B2(u4_srl_451_n136), .C1(
        u4_srl_451_n41), .C2(u4_srl_451_n135), .A(u4_srl_451_n724), .ZN(
        u4_srl_451_n592) );
  AOI22_X1 u4_srl_451_U661 ( .A1(fract_denorm[72]), .A2(u4_srl_451_n48), .B1(
        fract_denorm[71]), .B2(u4_srl_451_n52), .ZN(u4_srl_451_n723) );
  OAI221_X1 u4_srl_451_U660 ( .B1(u4_srl_451_n32), .B2(u4_srl_451_n132), .C1(
        u4_srl_451_n41), .C2(u4_srl_451_n131), .A(u4_srl_451_n723), .ZN(
        u4_srl_451_n479) );
  AOI22_X1 u4_srl_451_U659 ( .A1(u4_srl_451_n22), .A2(u4_srl_451_n592), .B1(
        u4_srl_451_n28), .B2(u4_srl_451_n479), .ZN(u4_srl_451_n722) );
  INV_X1 u4_srl_451_U658 ( .A(u4_srl_451_n722), .ZN(u4_srl_451_n721) );
  AOI221_X1 u4_srl_451_U657 ( .B1(u4_srl_451_n480), .B2(u4_srl_451_n18), .C1(
        u4_srl_451_n475), .C2(u4_srl_451_n62), .A(u4_srl_451_n721), .ZN(
        u4_srl_451_n283) );
  AOI22_X1 u4_srl_451_U656 ( .A1(fract_denorm[52]), .A2(u4_srl_451_n48), .B1(
        fract_denorm[51]), .B2(u4_srl_451_n52), .ZN(u4_srl_451_n720) );
  OAI221_X1 u4_srl_451_U655 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n112), .C1(
        u4_srl_451_n41), .C2(u4_srl_451_n111), .A(u4_srl_451_n720), .ZN(
        u4_srl_451_n492) );
  AOI22_X1 u4_srl_451_U654 ( .A1(fract_denorm[48]), .A2(u4_srl_451_n48), .B1(
        fract_denorm[47]), .B2(u4_srl_451_n52), .ZN(u4_srl_451_n719) );
  OAI221_X1 u4_srl_451_U653 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n108), .C1(
        u4_srl_451_n40), .C2(u4_srl_451_n107), .A(u4_srl_451_n719), .ZN(
        u4_srl_451_n487) );
  AOI22_X1 u4_srl_451_U652 ( .A1(fract_denorm[60]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[59]), .B2(u4_srl_451_n52), .ZN(u4_srl_451_n718) );
  OAI221_X1 u4_srl_451_U651 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n120), .C1(
        u4_srl_451_n40), .C2(u4_srl_451_n119), .A(u4_srl_451_n718), .ZN(
        u4_srl_451_n476) );
  AOI22_X1 u4_srl_451_U650 ( .A1(fract_denorm[56]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[55]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n717) );
  OAI221_X1 u4_srl_451_U649 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n116), .C1(
        u4_srl_451_n40), .C2(u4_srl_451_n115), .A(u4_srl_451_n717), .ZN(
        u4_srl_451_n491) );
  AOI22_X1 u4_srl_451_U648 ( .A1(u4_srl_451_n22), .A2(u4_srl_451_n476), .B1(
        u4_srl_451_n28), .B2(u4_srl_451_n491), .ZN(u4_srl_451_n716) );
  INV_X1 u4_srl_451_U647 ( .A(u4_srl_451_n716), .ZN(u4_srl_451_n715) );
  AOI221_X1 u4_srl_451_U646 ( .B1(u4_srl_451_n492), .B2(u4_srl_451_n18), .C1(
        u4_srl_451_n487), .C2(u4_srl_451_n62), .A(u4_srl_451_n715), .ZN(
        u4_srl_451_n363) );
  OAI22_X1 u4_srl_451_U645 ( .A1(u4_srl_451_n283), .A2(u4_srl_451_n182), .B1(
        u4_srl_451_n363), .B2(u4_srl_451_n184), .ZN(u4_srl_451_n714) );
  AOI221_X1 u4_srl_451_U644 ( .B1(u4_srl_451_n176), .B2(u4_srl_451_n713), .C1(
        u4_srl_451_n238), .C2(u4_srl_451_n179), .A(u4_srl_451_n714), .ZN(
        u4_srl_451_n706) );
  AOI22_X1 u4_srl_451_U643 ( .A1(fract_denorm[20]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[19]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n712) );
  OAI221_X1 u4_srl_451_U642 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n81), .C1(
        u4_srl_451_n40), .C2(u4_srl_451_n80), .A(u4_srl_451_n712), .ZN(
        u4_srl_451_n288) );
  AOI22_X1 u4_srl_451_U641 ( .A1(fract_denorm[16]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[15]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n711) );
  OAI221_X1 u4_srl_451_U640 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n77), .C1(
        u4_srl_451_n40), .C2(u4_srl_451_n76), .A(u4_srl_451_n711), .ZN(
        u4_srl_451_n168) );
  OAI22_X1 u4_srl_451_U639 ( .A1(u4_srl_451_n86), .A2(u4_srl_451_n1), .B1(
        u4_srl_451_n85), .B2(u4_srl_451_n58), .ZN(u4_srl_451_n710) );
  AOI221_X1 u4_srl_451_U638 ( .B1(u4_srl_451_n38), .B2(fract_denorm[22]), .C1(
        u4_srl_451_n45), .C2(fract_denorm[21]), .A(u4_srl_451_n710), .ZN(
        u4_srl_451_n174) );
  AOI22_X1 u4_srl_451_U637 ( .A1(fract_denorm[28]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[27]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n709) );
  OAI221_X1 u4_srl_451_U636 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n88), .C1(
        u4_srl_451_n40), .C2(u4_srl_451_n87), .A(u4_srl_451_n709), .ZN(
        u4_srl_451_n674) );
  INV_X1 u4_srl_451_U635 ( .A(u4_srl_451_n674), .ZN(u4_srl_451_n482) );
  OAI22_X1 u4_srl_451_U634 ( .A1(u4_srl_451_n174), .A2(u4_srl_451_n173), .B1(
        u4_srl_451_n482), .B2(u4_srl_451_n175), .ZN(u4_srl_451_n708) );
  AOI221_X1 u4_srl_451_U633 ( .B1(u4_srl_451_n167), .B2(u4_srl_451_n288), .C1(
        u4_srl_451_n169), .C2(u4_srl_451_n168), .A(u4_srl_451_n708), .ZN(
        u4_srl_451_n707) );
  AOI21_X1 u4_srl_451_U632 ( .B1(u4_srl_451_n706), .B2(u4_srl_451_n707), .A(
        u4_shift_right[8]), .ZN(u4_N5913) );
  AOI22_X1 u4_srl_451_U631 ( .A1(u4_srl_451_n22), .A2(u4_srl_451_n579), .B1(
        u4_srl_451_n28), .B2(u4_srl_451_n580), .ZN(u4_srl_451_n705) );
  INV_X1 u4_srl_451_U630 ( .A(u4_srl_451_n705), .ZN(u4_srl_451_n704) );
  AOI221_X1 u4_srl_451_U629 ( .B1(u4_srl_451_n577), .B2(u4_srl_451_n18), .C1(
        u4_srl_451_n578), .C2(u4_srl_451_n61), .A(u4_srl_451_n704), .ZN(
        u4_srl_451_n433) );
  INV_X1 u4_srl_451_U628 ( .A(u4_srl_451_n433), .ZN(u4_srl_451_n696) );
  AOI222_X1 u4_srl_451_U627 ( .A1(u4_srl_451_n566), .A2(u4_srl_451_n16), .B1(
        u4_srl_451_n411), .B2(u4_srl_451_n26), .C1(u4_srl_451_n567), .C2(
        u4_srl_451_n60), .ZN(u4_srl_451_n191) );
  INV_X1 u4_srl_451_U626 ( .A(u4_srl_451_n560), .ZN(u4_srl_451_n652) );
  AOI22_X1 u4_srl_451_U625 ( .A1(u4_srl_451_n22), .A2(u4_srl_451_n562), .B1(
        u4_srl_451_n28), .B2(u4_srl_451_n563), .ZN(u4_srl_451_n703) );
  OAI221_X1 u4_srl_451_U624 ( .B1(u4_srl_451_n652), .B2(u4_srl_451_n19), .C1(
        u4_srl_451_n702), .C2(u4_srl_451_n63), .A(u4_srl_451_n703), .ZN(
        u4_srl_451_n436) );
  INV_X1 u4_srl_451_U623 ( .A(u4_srl_451_n436), .ZN(u4_srl_451_n280) );
  OAI22_X1 u4_srl_451_U622 ( .A1(u4_srl_451_n191), .A2(u4_srl_451_n247), .B1(
        u4_srl_451_n280), .B2(u4_srl_451_n243), .ZN(u4_srl_451_n237) );
  AOI22_X1 u4_srl_451_U621 ( .A1(u4_srl_451_n22), .A2(u4_srl_451_n649), .B1(
        u4_srl_451_n28), .B2(u4_srl_451_n650), .ZN(u4_srl_451_n701) );
  INV_X1 u4_srl_451_U620 ( .A(u4_srl_451_n701), .ZN(u4_srl_451_n700) );
  AOI221_X1 u4_srl_451_U619 ( .B1(u4_srl_451_n572), .B2(u4_srl_451_n18), .C1(
        u4_srl_451_n573), .C2(u4_srl_451_n61), .A(u4_srl_451_n700), .ZN(
        u4_srl_451_n281) );
  AOI22_X1 u4_srl_451_U618 ( .A1(u4_srl_451_n22), .A2(u4_srl_451_n568), .B1(
        u4_srl_451_n28), .B2(u4_srl_451_n569), .ZN(u4_srl_451_n699) );
  INV_X1 u4_srl_451_U617 ( .A(u4_srl_451_n699), .ZN(u4_srl_451_n698) );
  AOI221_X1 u4_srl_451_U616 ( .B1(u4_srl_451_n583), .B2(u4_srl_451_n18), .C1(
        u4_srl_451_n584), .C2(u4_srl_451_n61), .A(u4_srl_451_n698), .ZN(
        u4_srl_451_n358) );
  OAI22_X1 u4_srl_451_U615 ( .A1(u4_srl_451_n281), .A2(u4_srl_451_n182), .B1(
        u4_srl_451_n358), .B2(u4_srl_451_n184), .ZN(u4_srl_451_n697) );
  AOI221_X1 u4_srl_451_U614 ( .B1(u4_srl_451_n176), .B2(u4_srl_451_n696), .C1(
        u4_srl_451_n237), .C2(u4_srl_451_n179), .A(u4_srl_451_n697), .ZN(
        u4_srl_451_n693) );
  INV_X1 u4_srl_451_U613 ( .A(u4_srl_451_n659), .ZN(u4_srl_451_n574) );
  OAI22_X1 u4_srl_451_U612 ( .A1(u4_srl_451_n575), .A2(u4_srl_451_n173), .B1(
        u4_srl_451_n574), .B2(u4_srl_451_n175), .ZN(u4_srl_451_n695) );
  AOI221_X1 u4_srl_451_U611 ( .B1(u4_srl_451_n167), .B2(u4_srl_451_n257), .C1(
        u4_srl_451_n169), .C2(u4_srl_451_n258), .A(u4_srl_451_n695), .ZN(
        u4_srl_451_n694) );
  AOI21_X1 u4_srl_451_U610 ( .B1(u4_srl_451_n693), .B2(u4_srl_451_n694), .A(
        u4_shift_right[8]), .ZN(u4_N5914) );
  AOI22_X1 u4_srl_451_U609 ( .A1(u4_srl_451_n22), .A2(u4_srl_451_n548), .B1(
        u4_srl_451_n28), .B2(u4_srl_451_n549), .ZN(u4_srl_451_n692) );
  INV_X1 u4_srl_451_U608 ( .A(u4_srl_451_n692), .ZN(u4_srl_451_n691) );
  AOI221_X1 u4_srl_451_U607 ( .B1(u4_srl_451_n546), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n547), .C2(u4_srl_451_n61), .A(u4_srl_451_n691), .ZN(
        u4_srl_451_n428) );
  INV_X1 u4_srl_451_U606 ( .A(u4_srl_451_n428), .ZN(u4_srl_451_n683) );
  AOI222_X1 u4_srl_451_U605 ( .A1(u4_srl_451_n535), .A2(u4_srl_451_n16), .B1(
        u4_srl_451_n408), .B2(u4_srl_451_n26), .C1(u4_srl_451_n536), .C2(
        u4_srl_451_n60), .ZN(u4_srl_451_n190) );
  INV_X1 u4_srl_451_U604 ( .A(u4_srl_451_n529), .ZN(u4_srl_451_n635) );
  AOI22_X1 u4_srl_451_U603 ( .A1(u4_srl_451_n22), .A2(u4_srl_451_n531), .B1(
        u4_srl_451_n28), .B2(u4_srl_451_n532), .ZN(u4_srl_451_n690) );
  OAI221_X1 u4_srl_451_U602 ( .B1(u4_srl_451_n635), .B2(u4_srl_451_n19), .C1(
        u4_srl_451_n689), .C2(u4_srl_451_n63), .A(u4_srl_451_n690), .ZN(
        u4_srl_451_n431) );
  INV_X1 u4_srl_451_U601 ( .A(u4_srl_451_n431), .ZN(u4_srl_451_n278) );
  OAI22_X1 u4_srl_451_U600 ( .A1(u4_srl_451_n190), .A2(u4_srl_451_n247), .B1(
        u4_srl_451_n278), .B2(u4_srl_451_n243), .ZN(u4_srl_451_n236) );
  INV_X1 u4_srl_451_U599 ( .A(u4_srl_451_n541), .ZN(u4_srl_451_n630) );
  INV_X1 u4_srl_451_U598 ( .A(u4_srl_451_n542), .ZN(u4_srl_451_n687) );
  AOI22_X1 u4_srl_451_U597 ( .A1(u4_srl_451_n22), .A2(u4_srl_451_n632), .B1(
        u4_srl_451_n28), .B2(u4_srl_451_n633), .ZN(u4_srl_451_n688) );
  OAI221_X1 u4_srl_451_U596 ( .B1(u4_srl_451_n630), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n687), .C2(u4_srl_451_n63), .A(u4_srl_451_n688), .ZN(
        u4_srl_451_n430) );
  INV_X1 u4_srl_451_U595 ( .A(u4_srl_451_n430), .ZN(u4_srl_451_n279) );
  AOI22_X1 u4_srl_451_U594 ( .A1(u4_srl_451_n22), .A2(u4_srl_451_n537), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n538), .ZN(u4_srl_451_n686) );
  INV_X1 u4_srl_451_U593 ( .A(u4_srl_451_n686), .ZN(u4_srl_451_n685) );
  AOI221_X1 u4_srl_451_U592 ( .B1(u4_srl_451_n552), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n553), .C2(u4_srl_451_n61), .A(u4_srl_451_n685), .ZN(
        u4_srl_451_n355) );
  OAI22_X1 u4_srl_451_U591 ( .A1(u4_srl_451_n279), .A2(u4_srl_451_n182), .B1(
        u4_srl_451_n355), .B2(u4_srl_451_n184), .ZN(u4_srl_451_n684) );
  AOI221_X1 u4_srl_451_U590 ( .B1(u4_srl_451_n176), .B2(u4_srl_451_n683), .C1(
        u4_srl_451_n236), .C2(u4_srl_451_n179), .A(u4_srl_451_n684), .ZN(
        u4_srl_451_n680) );
  INV_X1 u4_srl_451_U589 ( .A(u4_srl_451_n640), .ZN(u4_srl_451_n224) );
  INV_X1 u4_srl_451_U588 ( .A(u4_srl_451_n642), .ZN(u4_srl_451_n543) );
  OAI22_X1 u4_srl_451_U587 ( .A1(u4_srl_451_n544), .A2(u4_srl_451_n173), .B1(
        u4_srl_451_n543), .B2(u4_srl_451_n175), .ZN(u4_srl_451_n682) );
  AOI221_X1 u4_srl_451_U586 ( .B1(u4_srl_451_n167), .B2(u4_srl_451_n224), .C1(
        u4_srl_451_n169), .C2(u4_srl_451_n226), .A(u4_srl_451_n682), .ZN(
        u4_srl_451_n681) );
  AOI21_X1 u4_srl_451_U585 ( .B1(u4_srl_451_n680), .B2(u4_srl_451_n681), .A(
        u4_shift_right[8]), .ZN(u4_N5915) );
  AOI22_X1 u4_srl_451_U584 ( .A1(u4_srl_451_n351), .A2(u4_srl_451_n406), .B1(
        u4_srl_451_n352), .B2(u4_srl_451_n405), .ZN(u4_srl_451_n220) );
  INV_X1 u4_srl_451_U583 ( .A(u4_srl_451_n427), .ZN(u4_srl_451_n348) );
  OAI222_X1 u4_srl_451_U582 ( .A1(u4_srl_451_n3), .A2(u4_srl_451_n349), .B1(
        u4_srl_451_n388), .B2(u4_srl_451_n220), .C1(u4_srl_451_n12), .C2(
        u4_srl_451_n348), .ZN(u4_srl_451_n679) );
  INV_X1 u4_srl_451_U581 ( .A(u4_srl_451_n679), .ZN(u4_srl_451_n678) );
  OAI221_X1 u4_srl_451_U580 ( .B1(u4_srl_451_n425), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n677), .C2(u4_srl_451_n9), .A(u4_srl_451_n678), .ZN(
        u4_N5916) );
  AOI22_X1 u4_srl_451_U579 ( .A1(u4_srl_451_n22), .A2(u4_srl_451_n487), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n488), .ZN(u4_srl_451_n676) );
  INV_X1 u4_srl_451_U578 ( .A(u4_srl_451_n676), .ZN(u4_srl_451_n675) );
  AOI221_X1 u4_srl_451_U577 ( .B1(u4_srl_451_n484), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n485), .C2(u4_srl_451_n61), .A(u4_srl_451_n675), .ZN(
        u4_srl_451_n422) );
  INV_X1 u4_srl_451_U576 ( .A(u4_srl_451_n288), .ZN(u4_srl_451_n172) );
  AOI22_X1 u4_srl_451_U575 ( .A1(u4_srl_451_n22), .A2(u4_srl_451_n486), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n674), .ZN(u4_srl_451_n673) );
  OAI221_X1 u4_srl_451_U574 ( .B1(u4_srl_451_n174), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n172), .C2(u4_srl_451_n63), .A(u4_srl_451_n673), .ZN(
        u4_srl_451_n672) );
  INV_X1 u4_srl_451_U573 ( .A(u4_srl_451_n672), .ZN(u4_srl_451_n622) );
  AOI22_X1 u4_srl_451_U572 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n475), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n476), .ZN(u4_srl_451_n671) );
  INV_X1 u4_srl_451_U571 ( .A(u4_srl_451_n671), .ZN(u4_srl_451_n670) );
  AOI221_X1 u4_srl_451_U570 ( .B1(u4_srl_451_n491), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n492), .C2(u4_srl_451_n61), .A(u4_srl_451_n670), .ZN(
        u4_srl_451_n344) );
  AOI222_X1 u4_srl_451_U569 ( .A1(u4_srl_451_n473), .A2(u4_srl_451_n16), .B1(
        u4_srl_451_n26), .B2(u4_srl_451_n669), .C1(u4_srl_451_n474), .C2(
        u4_srl_451_n60), .ZN(u4_srl_451_n188) );
  INV_X1 u4_srl_451_U568 ( .A(u4_srl_451_n188), .ZN(u4_srl_451_n346) );
  INV_X1 u4_srl_451_U567 ( .A(u4_srl_451_n466), .ZN(u4_srl_451_n666) );
  AOI22_X1 u4_srl_451_U566 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n469), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n470), .ZN(u4_srl_451_n668) );
  OAI221_X1 u4_srl_451_U565 ( .B1(u4_srl_451_n666), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n667), .C2(u4_srl_451_n63), .A(u4_srl_451_n668), .ZN(
        u4_srl_451_n347) );
  AOI22_X1 u4_srl_451_U564 ( .A1(u4_srl_451_n346), .A2(u4_srl_451_n406), .B1(
        u4_srl_451_n347), .B2(u4_srl_451_n405), .ZN(u4_srl_451_n219) );
  AOI22_X1 u4_srl_451_U563 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n591), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n592), .ZN(u4_srl_451_n665) );
  INV_X1 u4_srl_451_U562 ( .A(u4_srl_451_n665), .ZN(u4_srl_451_n664) );
  AOI221_X1 u4_srl_451_U561 ( .B1(u4_srl_451_n479), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n480), .C2(u4_srl_451_n61), .A(u4_srl_451_n664), .ZN(
        u4_srl_451_n343) );
  OAI222_X1 u4_srl_451_U560 ( .A1(u4_srl_451_n3), .A2(u4_srl_451_n344), .B1(
        u4_srl_451_n388), .B2(u4_srl_451_n219), .C1(u4_srl_451_n12), .C2(
        u4_srl_451_n343), .ZN(u4_srl_451_n663) );
  INV_X1 u4_srl_451_U559 ( .A(u4_srl_451_n663), .ZN(u4_srl_451_n662) );
  OAI221_X1 u4_srl_451_U558 ( .B1(u4_srl_451_n422), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n622), .C2(u4_srl_451_n9), .A(u4_srl_451_n662), .ZN(
        u4_N5917) );
  AOI22_X1 u4_srl_451_U557 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n584), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n579), .ZN(u4_srl_451_n661) );
  INV_X1 u4_srl_451_U556 ( .A(u4_srl_451_n661), .ZN(u4_srl_451_n660) );
  AOI221_X1 u4_srl_451_U555 ( .B1(u4_srl_451_n580), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n577), .C2(u4_srl_451_n61), .A(u4_srl_451_n660), .ZN(
        u4_srl_451_n419) );
  AOI22_X1 u4_srl_451_U554 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n578), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n659), .ZN(u4_srl_451_n658) );
  OAI221_X1 u4_srl_451_U553 ( .B1(u4_srl_451_n575), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n657), .C2(u4_srl_451_n63), .A(u4_srl_451_n658), .ZN(
        u4_srl_451_n656) );
  INV_X1 u4_srl_451_U552 ( .A(u4_srl_451_n656), .ZN(u4_srl_451_n443) );
  AOI22_X1 u4_srl_451_U551 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n573), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n568), .ZN(u4_srl_451_n655) );
  INV_X1 u4_srl_451_U550 ( .A(u4_srl_451_n655), .ZN(u4_srl_451_n654) );
  AOI221_X1 u4_srl_451_U549 ( .B1(u4_srl_451_n569), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n583), .C2(u4_srl_451_n61), .A(u4_srl_451_n654), .ZN(
        u4_srl_451_n326) );
  AOI22_X1 u4_srl_451_U548 ( .A1(u4_srl_451_n566), .A2(u4_srl_451_n61), .B1(
        u4_srl_451_n411), .B2(u4_srl_451_n17), .ZN(u4_srl_451_n187) );
  INV_X1 u4_srl_451_U547 ( .A(u4_srl_451_n187), .ZN(u4_srl_451_n328) );
  INV_X1 u4_srl_451_U546 ( .A(u4_srl_451_n563), .ZN(u4_srl_451_n651) );
  AOI22_X1 u4_srl_451_U545 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n567), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n562), .ZN(u4_srl_451_n653) );
  OAI221_X1 u4_srl_451_U544 ( .B1(u4_srl_451_n651), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n652), .C2(u4_srl_451_n64), .A(u4_srl_451_n653), .ZN(
        u4_srl_451_n329) );
  AOI22_X1 u4_srl_451_U543 ( .A1(u4_srl_451_n328), .A2(u4_srl_451_n406), .B1(
        u4_srl_451_n329), .B2(u4_srl_451_n405), .ZN(u4_srl_451_n218) );
  INV_X1 u4_srl_451_U542 ( .A(u4_srl_451_n650), .ZN(u4_srl_451_n558) );
  INV_X1 u4_srl_451_U541 ( .A(u4_srl_451_n572), .ZN(u4_srl_451_n647) );
  AOI22_X1 u4_srl_451_U540 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n561), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n649), .ZN(u4_srl_451_n648) );
  OAI221_X1 u4_srl_451_U539 ( .B1(u4_srl_451_n558), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n647), .C2(u4_srl_451_n64), .A(u4_srl_451_n648), .ZN(
        u4_srl_451_n421) );
  INV_X1 u4_srl_451_U538 ( .A(u4_srl_451_n421), .ZN(u4_srl_451_n325) );
  OAI222_X1 u4_srl_451_U537 ( .A1(u4_srl_451_n3), .A2(u4_srl_451_n326), .B1(
        u4_srl_451_n388), .B2(u4_srl_451_n218), .C1(u4_srl_451_n12), .C2(
        u4_srl_451_n325), .ZN(u4_srl_451_n646) );
  INV_X1 u4_srl_451_U536 ( .A(u4_srl_451_n646), .ZN(u4_srl_451_n645) );
  OAI221_X1 u4_srl_451_U535 ( .B1(u4_srl_451_n419), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n443), .C2(u4_srl_451_n9), .A(u4_srl_451_n645), .ZN(
        u4_N5918) );
  AOI22_X1 u4_srl_451_U534 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n553), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n548), .ZN(u4_srl_451_n644) );
  INV_X1 u4_srl_451_U533 ( .A(u4_srl_451_n644), .ZN(u4_srl_451_n643) );
  AOI221_X1 u4_srl_451_U532 ( .B1(u4_srl_451_n549), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n546), .C2(u4_srl_451_n61), .A(u4_srl_451_n643), .ZN(
        u4_srl_451_n403) );
  AOI22_X1 u4_srl_451_U531 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n547), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n642), .ZN(u4_srl_451_n641) );
  OAI221_X1 u4_srl_451_U530 ( .B1(u4_srl_451_n544), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n640), .C2(u4_srl_451_n64), .A(u4_srl_451_n641), .ZN(
        u4_srl_451_n639) );
  INV_X1 u4_srl_451_U529 ( .A(u4_srl_451_n639), .ZN(u4_srl_451_n395) );
  AOI22_X1 u4_srl_451_U528 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n542), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n537), .ZN(u4_srl_451_n638) );
  INV_X1 u4_srl_451_U527 ( .A(u4_srl_451_n638), .ZN(u4_srl_451_n637) );
  AOI221_X1 u4_srl_451_U526 ( .B1(u4_srl_451_n538), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n552), .C2(u4_srl_451_n61), .A(u4_srl_451_n637), .ZN(
        u4_srl_451_n321) );
  AOI22_X1 u4_srl_451_U525 ( .A1(u4_srl_451_n535), .A2(u4_srl_451_n61), .B1(
        u4_srl_451_n408), .B2(u4_srl_451_n17), .ZN(u4_srl_451_n185) );
  INV_X1 u4_srl_451_U524 ( .A(u4_srl_451_n185), .ZN(u4_srl_451_n323) );
  INV_X1 u4_srl_451_U523 ( .A(u4_srl_451_n532), .ZN(u4_srl_451_n634) );
  AOI22_X1 u4_srl_451_U522 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n536), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n531), .ZN(u4_srl_451_n636) );
  OAI221_X1 u4_srl_451_U521 ( .B1(u4_srl_451_n634), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n635), .C2(u4_srl_451_n64), .A(u4_srl_451_n636), .ZN(
        u4_srl_451_n324) );
  AOI22_X1 u4_srl_451_U520 ( .A1(u4_srl_451_n323), .A2(u4_srl_451_n406), .B1(
        u4_srl_451_n324), .B2(u4_srl_451_n405), .ZN(u4_srl_451_n216) );
  INV_X1 u4_srl_451_U519 ( .A(u4_srl_451_n633), .ZN(u4_srl_451_n527) );
  AOI22_X1 u4_srl_451_U518 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n530), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n632), .ZN(u4_srl_451_n631) );
  OAI221_X1 u4_srl_451_U517 ( .B1(u4_srl_451_n527), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n630), .C2(u4_srl_451_n64), .A(u4_srl_451_n631), .ZN(
        u4_srl_451_n404) );
  INV_X1 u4_srl_451_U516 ( .A(u4_srl_451_n404), .ZN(u4_srl_451_n320) );
  OAI222_X1 u4_srl_451_U515 ( .A1(u4_srl_451_n3), .A2(u4_srl_451_n321), .B1(
        u4_srl_451_n388), .B2(u4_srl_451_n216), .C1(u4_srl_451_n12), .C2(
        u4_srl_451_n320), .ZN(u4_srl_451_n629) );
  INV_X1 u4_srl_451_U514 ( .A(u4_srl_451_n629), .ZN(u4_srl_451_n628) );
  OAI221_X1 u4_srl_451_U513 ( .B1(u4_srl_451_n403), .B2(u4_srl_451_n11), .C1(
        u4_srl_451_n395), .C2(u4_srl_451_n9), .A(u4_srl_451_n628), .ZN(
        u4_N5919) );
  INV_X1 u4_srl_451_U512 ( .A(u4_srl_451_n343), .ZN(u4_srl_451_n424) );
  AOI222_X1 u4_srl_451_U511 ( .A1(u4_srl_451_n424), .A2(u4_srl_451_n405), .B1(
        u4_srl_451_n346), .B2(u4_srl_451_n341), .C1(u4_srl_451_n347), .C2(
        u4_srl_451_n406), .ZN(u4_srl_451_n276) );
  INV_X1 u4_srl_451_U510 ( .A(u4_srl_451_n422), .ZN(u4_srl_451_n618) );
  AOI22_X1 u4_srl_451_U509 ( .A1(u4_srl_451_n45), .A2(fract_denorm[1]), .B1(
        u4_srl_451_n38), .B2(fract_denorm[2]), .ZN(u4_srl_451_n627) );
  INV_X1 u4_srl_451_U508 ( .A(u4_srl_451_n627), .ZN(u4_srl_451_n626) );
  AOI221_X1 u4_srl_451_U507 ( .B1(fract_denorm[4]), .B2(u4_srl_451_n47), .C1(
        fract_denorm[3]), .C2(u4_srl_451_n55), .A(u4_srl_451_n626), .ZN(
        u4_srl_451_n620) );
  AOI22_X1 u4_srl_451_U506 ( .A1(fract_denorm[8]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[7]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n625) );
  OAI221_X1 u4_srl_451_U505 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n69), .C1(
        u4_srl_451_n40), .C2(u4_srl_451_n68), .A(u4_srl_451_n625), .ZN(
        u4_srl_451_n291) );
  AOI22_X1 u4_srl_451_U504 ( .A1(fract_denorm[12]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[11]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n624) );
  OAI221_X1 u4_srl_451_U503 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n73), .C1(
        u4_srl_451_n40), .C2(u4_srl_451_n72), .A(u4_srl_451_n624), .ZN(
        u4_srl_451_n170) );
  AOI222_X1 u4_srl_451_U502 ( .A1(u4_srl_451_n16), .A2(u4_srl_451_n291), .B1(
        u4_srl_451_n21), .B2(u4_srl_451_n168), .C1(u4_srl_451_n26), .C2(
        u4_srl_451_n170), .ZN(u4_srl_451_n623) );
  MUX2_X1 u4_srl_451_U501 ( .A(u4_srl_451_n622), .B(u4_srl_451_n623), .S(
        u4_srl_451_n397), .Z(u4_srl_451_n621) );
  OAI21_X1 u4_srl_451_U500 ( .B1(u4_srl_451_n620), .B2(u4_srl_451_n270), .A(
        u4_srl_451_n621), .ZN(u4_srl_451_n619) );
  AOI22_X1 u4_srl_451_U499 ( .A1(u4_srl_451_n15), .A2(u4_srl_451_n618), .B1(
        u4_srl_451_n391), .B2(u4_srl_451_n619), .ZN(u4_srl_451_n617) );
  OAI221_X1 u4_srl_451_U498 ( .B1(u4_srl_451_n276), .B2(u4_srl_451_n388), .C1(
        u4_srl_451_n344), .C2(u4_srl_451_n12), .A(u4_srl_451_n617), .ZN(
        u4_N5901) );
  AOI22_X1 u4_srl_451_U497 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n522), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n517), .ZN(u4_srl_451_n616) );
  INV_X1 u4_srl_451_U496 ( .A(u4_srl_451_n616), .ZN(u4_srl_451_n615) );
  AOI221_X1 u4_srl_451_U495 ( .B1(u4_srl_451_n518), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n514), .C2(u4_srl_451_n61), .A(u4_srl_451_n615), .ZN(
        u4_srl_451_n338) );
  AOI22_X1 u4_srl_451_U494 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n515), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n516), .ZN(u4_srl_451_n614) );
  OAI221_X1 u4_srl_451_U493 ( .B1(u4_srl_451_n512), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n202), .C2(u4_srl_451_n64), .A(u4_srl_451_n614), .ZN(
        u4_srl_451_n336) );
  INV_X1 u4_srl_451_U492 ( .A(u4_srl_451_n336), .ZN(u4_srl_451_n600) );
  AOI22_X1 u4_srl_451_U491 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n509), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n613), .ZN(u4_srl_451_n612) );
  INV_X1 u4_srl_451_U490 ( .A(u4_srl_451_n612), .ZN(u4_srl_451_n611) );
  AOI221_X1 u4_srl_451_U489 ( .B1(u4_srl_451_n510), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n521), .C2(u4_srl_451_n61), .A(u4_srl_451_n611), .ZN(
        u4_srl_451_n315) );
  INV_X1 u4_srl_451_U488 ( .A(u4_srl_451_n315), .ZN(u4_srl_451_n602) );
  INV_X1 u4_srl_451_U487 ( .A(u4_srl_451_n610), .ZN(u4_srl_451_n501) );
  AOI22_X1 u4_srl_451_U486 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n504), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n609), .ZN(u4_srl_451_n608) );
  OAI221_X1 u4_srl_451_U485 ( .B1(u4_srl_451_n501), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n607), .C2(u4_srl_451_n64), .A(u4_srl_451_n608), .ZN(
        u4_srl_451_n319) );
  INV_X1 u4_srl_451_U484 ( .A(u4_srl_451_n319), .ZN(u4_srl_451_n340) );
  OAI22_X1 u4_srl_451_U483 ( .A1(u4_srl_451_n339), .A2(u4_srl_451_n247), .B1(
        u4_srl_451_n340), .B2(u4_srl_451_n243), .ZN(u4_srl_451_n214) );
  INV_X1 u4_srl_451_U482 ( .A(u4_srl_451_n606), .ZN(u4_srl_451_n496) );
  AOI22_X1 u4_srl_451_U481 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n499), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n605), .ZN(u4_srl_451_n604) );
  OAI221_X1 u4_srl_451_U480 ( .B1(u4_srl_451_n496), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n603), .C2(u4_srl_451_n64), .A(u4_srl_451_n604), .ZN(
        u4_srl_451_n342) );
  AOI222_X1 u4_srl_451_U479 ( .A1(u4_srl_451_n14), .A2(u4_srl_451_n602), .B1(
        u4_srl_451_n381), .B2(u4_srl_451_n214), .C1(u4_srl_451_n317), .C2(
        u4_srl_451_n342), .ZN(u4_srl_451_n601) );
  OAI221_X1 u4_srl_451_U478 ( .B1(u4_srl_451_n338), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n600), .C2(u4_srl_451_n9), .A(u4_srl_451_n601), .ZN(
        u4_N5920) );
  AOI22_X1 u4_srl_451_U477 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n492), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n487), .ZN(u4_srl_451_n599) );
  INV_X1 u4_srl_451_U476 ( .A(u4_srl_451_n599), .ZN(u4_srl_451_n598) );
  AOI221_X1 u4_srl_451_U475 ( .B1(u4_srl_451_n488), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n484), .C2(u4_srl_451_n61), .A(u4_srl_451_n598), .ZN(
        u4_srl_451_n295) );
  AOI22_X1 u4_srl_451_U474 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n485), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n486), .ZN(u4_srl_451_n597) );
  OAI221_X1 u4_srl_451_U473 ( .B1(u4_srl_451_n482), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n174), .C2(u4_srl_451_n64), .A(u4_srl_451_n597), .ZN(
        u4_srl_451_n292) );
  INV_X1 u4_srl_451_U472 ( .A(u4_srl_451_n292), .ZN(u4_srl_451_n585) );
  AOI22_X1 u4_srl_451_U471 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n480), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n475), .ZN(u4_srl_451_n596) );
  INV_X1 u4_srl_451_U470 ( .A(u4_srl_451_n596), .ZN(u4_srl_451_n595) );
  AOI221_X1 u4_srl_451_U469 ( .B1(u4_srl_451_n476), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n491), .C2(u4_srl_451_n61), .A(u4_srl_451_n595), .ZN(
        u4_srl_451_n294) );
  INV_X1 u4_srl_451_U468 ( .A(u4_srl_451_n294), .ZN(u4_srl_451_n587) );
  AND2_X1 u4_srl_451_U467 ( .A1(u4_srl_451_n381), .A2(u4_srl_451_n271), .ZN(
        u4_srl_451_n462) );
  AOI22_X1 u4_srl_451_U466 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n474), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n469), .ZN(u4_srl_451_n594) );
  INV_X1 u4_srl_451_U465 ( .A(u4_srl_451_n594), .ZN(u4_srl_451_n593) );
  AOI221_X1 u4_srl_451_U464 ( .B1(u4_srl_451_n470), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n466), .C2(u4_srl_451_n61), .A(u4_srl_451_n593), .ZN(
        u4_srl_451_n299) );
  MUX2_X1 u4_srl_451_U463 ( .A(u4_srl_451_n297), .B(u4_srl_451_n299), .S(
        u4_srl_451_n397), .Z(u4_srl_451_n213) );
  INV_X1 u4_srl_451_U462 ( .A(u4_srl_451_n213), .ZN(u4_srl_451_n588) );
  INV_X1 u4_srl_451_U461 ( .A(u4_srl_451_n592), .ZN(u4_srl_451_n464) );
  INV_X1 u4_srl_451_U460 ( .A(u4_srl_451_n479), .ZN(u4_srl_451_n589) );
  AOI22_X1 u4_srl_451_U459 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n467), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n591), .ZN(u4_srl_451_n590) );
  OAI221_X1 u4_srl_451_U458 ( .B1(u4_srl_451_n464), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n589), .C2(u4_srl_451_n64), .A(u4_srl_451_n590), .ZN(
        u4_srl_451_n313) );
  AOI222_X1 u4_srl_451_U457 ( .A1(u4_srl_451_n14), .A2(u4_srl_451_n587), .B1(
        u4_srl_451_n462), .B2(u4_srl_451_n588), .C1(u4_srl_451_n317), .C2(
        u4_srl_451_n313), .ZN(u4_srl_451_n586) );
  OAI221_X1 u4_srl_451_U456 ( .B1(u4_srl_451_n295), .B2(u4_srl_451_n11), .C1(
        u4_srl_451_n585), .C2(u4_srl_451_n9), .A(u4_srl_451_n586), .ZN(
        u4_N5921) );
  AOI22_X1 u4_srl_451_U455 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n583), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n584), .ZN(u4_srl_451_n582) );
  INV_X1 u4_srl_451_U454 ( .A(u4_srl_451_n582), .ZN(u4_srl_451_n581) );
  AOI221_X1 u4_srl_451_U453 ( .B1(u4_srl_451_n579), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n580), .C2(u4_srl_451_n61), .A(u4_srl_451_n581), .ZN(
        u4_srl_451_n266) );
  AOI22_X1 u4_srl_451_U452 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n577), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n578), .ZN(u4_srl_451_n576) );
  OAI221_X1 u4_srl_451_U451 ( .B1(u4_srl_451_n574), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n575), .C2(u4_srl_451_n63), .A(u4_srl_451_n576), .ZN(
        u4_srl_451_n263) );
  INV_X1 u4_srl_451_U450 ( .A(u4_srl_451_n263), .ZN(u4_srl_451_n554) );
  AOI22_X1 u4_srl_451_U449 ( .A1(u4_srl_451_n24), .A2(u4_srl_451_n572), .B1(
        u4_srl_451_n30), .B2(u4_srl_451_n573), .ZN(u4_srl_451_n571) );
  INV_X1 u4_srl_451_U448 ( .A(u4_srl_451_n571), .ZN(u4_srl_451_n570) );
  AOI221_X1 u4_srl_451_U447 ( .B1(u4_srl_451_n568), .B2(u4_srl_451_n18), .C1(
        u4_srl_451_n569), .C2(u4_srl_451_n62), .A(u4_srl_451_n570), .ZN(
        u4_srl_451_n265) );
  INV_X1 u4_srl_451_U446 ( .A(u4_srl_451_n265), .ZN(u4_srl_451_n556) );
  AOI22_X1 u4_srl_451_U445 ( .A1(u4_srl_451_n399), .A2(u4_srl_451_n566), .B1(
        u4_srl_451_n28), .B2(u4_srl_451_n567), .ZN(u4_srl_451_n565) );
  INV_X1 u4_srl_451_U444 ( .A(u4_srl_451_n565), .ZN(u4_srl_451_n564) );
  AOI221_X1 u4_srl_451_U443 ( .B1(u4_srl_451_n562), .B2(u4_srl_451_n16), .C1(
        u4_srl_451_n563), .C2(u4_srl_451_n5), .A(u4_srl_451_n564), .ZN(
        u4_srl_451_n269) );
  NAND2_X1 u4_srl_451_U442 ( .A1(u4_srl_451_n5), .A2(u4_shift_right[4]), .ZN(
        u4_srl_451_n468) );
  OAI22_X1 u4_srl_451_U441 ( .A1(u4_shift_right[4]), .A2(u4_srl_451_n269), 
        .B1(u4_srl_451_n268), .B2(u4_srl_451_n468), .ZN(u4_srl_451_n311) );
  AOI22_X1 u4_srl_451_U440 ( .A1(u4_srl_451_n22), .A2(u4_srl_451_n560), .B1(
        u4_srl_451_n29), .B2(u4_srl_451_n561), .ZN(u4_srl_451_n559) );
  OAI221_X1 u4_srl_451_U439 ( .B1(u4_srl_451_n557), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n558), .C2(u4_srl_451_n64), .A(u4_srl_451_n559), .ZN(
        u4_srl_451_n312) );
  AOI222_X1 u4_srl_451_U438 ( .A1(u4_srl_451_n14), .A2(u4_srl_451_n556), .B1(
        u4_srl_451_n462), .B2(u4_srl_451_n311), .C1(u4_srl_451_n317), .C2(
        u4_srl_451_n312), .ZN(u4_srl_451_n555) );
  OAI221_X1 u4_srl_451_U437 ( .B1(u4_srl_451_n266), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n554), .C2(u4_srl_451_n9), .A(u4_srl_451_n555), .ZN(
        u4_N5922) );
  AOI22_X1 u4_srl_451_U436 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n552), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n553), .ZN(u4_srl_451_n551) );
  INV_X1 u4_srl_451_U435 ( .A(u4_srl_451_n551), .ZN(u4_srl_451_n550) );
  AOI221_X1 u4_srl_451_U434 ( .B1(u4_srl_451_n548), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n549), .C2(u4_srl_451_n61), .A(u4_srl_451_n550), .ZN(
        u4_srl_451_n235) );
  AOI22_X1 u4_srl_451_U433 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n546), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n547), .ZN(u4_srl_451_n545) );
  OAI221_X1 u4_srl_451_U432 ( .B1(u4_srl_451_n543), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n544), .C2(u4_srl_451_n64), .A(u4_srl_451_n545), .ZN(
        u4_srl_451_n231) );
  INV_X1 u4_srl_451_U431 ( .A(u4_srl_451_n231), .ZN(u4_srl_451_n523) );
  AOI22_X1 u4_srl_451_U430 ( .A1(u4_srl_451_n23), .A2(u4_srl_451_n541), .B1(
        u4_srl_451_n29), .B2(u4_srl_451_n542), .ZN(u4_srl_451_n540) );
  INV_X1 u4_srl_451_U429 ( .A(u4_srl_451_n540), .ZN(u4_srl_451_n539) );
  AOI221_X1 u4_srl_451_U428 ( .B1(u4_srl_451_n537), .B2(u4_srl_451_n18), .C1(
        u4_srl_451_n538), .C2(u4_srl_451_n60), .A(u4_srl_451_n539), .ZN(
        u4_srl_451_n234) );
  INV_X1 u4_srl_451_U427 ( .A(u4_srl_451_n234), .ZN(u4_srl_451_n525) );
  AOI22_X1 u4_srl_451_U426 ( .A1(u4_srl_451_n399), .A2(u4_srl_451_n535), .B1(
        u4_srl_451_n26), .B2(u4_srl_451_n536), .ZN(u4_srl_451_n534) );
  INV_X1 u4_srl_451_U425 ( .A(u4_srl_451_n534), .ZN(u4_srl_451_n533) );
  AOI221_X1 u4_srl_451_U424 ( .B1(u4_srl_451_n531), .B2(u4_srl_451_n16), .C1(
        u4_srl_451_n532), .C2(u4_srl_451_n60), .A(u4_srl_451_n533), .ZN(
        u4_srl_451_n253) );
  OAI22_X1 u4_srl_451_U423 ( .A1(u4_shift_right[4]), .A2(u4_srl_451_n253), 
        .B1(u4_srl_451_n252), .B2(u4_srl_451_n468), .ZN(u4_srl_451_n309) );
  AOI22_X1 u4_srl_451_U422 ( .A1(u4_srl_451_n22), .A2(u4_srl_451_n529), .B1(
        u4_srl_451_n28), .B2(u4_srl_451_n530), .ZN(u4_srl_451_n528) );
  OAI221_X1 u4_srl_451_U421 ( .B1(u4_srl_451_n526), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n527), .C2(u4_srl_451_n64), .A(u4_srl_451_n528), .ZN(
        u4_srl_451_n310) );
  AOI222_X1 u4_srl_451_U420 ( .A1(u4_srl_451_n14), .A2(u4_srl_451_n525), .B1(
        u4_srl_451_n462), .B2(u4_srl_451_n309), .C1(u4_srl_451_n317), .C2(
        u4_srl_451_n310), .ZN(u4_srl_451_n524) );
  OAI221_X1 u4_srl_451_U419 ( .B1(u4_srl_451_n235), .B2(u4_srl_451_n11), .C1(
        u4_srl_451_n523), .C2(u4_srl_451_n9), .A(u4_srl_451_n524), .ZN(
        u4_N5923) );
  AOI22_X1 u4_srl_451_U418 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n521), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n522), .ZN(u4_srl_451_n520) );
  INV_X1 u4_srl_451_U417 ( .A(u4_srl_451_n520), .ZN(u4_srl_451_n519) );
  AOI221_X1 u4_srl_451_U416 ( .B1(u4_srl_451_n517), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n518), .C2(u4_srl_451_n60), .A(u4_srl_451_n519), .ZN(
        u4_srl_451_n207) );
  INV_X1 u4_srl_451_U415 ( .A(u4_srl_451_n516), .ZN(u4_srl_451_n511) );
  AOI22_X1 u4_srl_451_U414 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n514), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n515), .ZN(u4_srl_451_n513) );
  OAI221_X1 u4_srl_451_U413 ( .B1(u4_srl_451_n511), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n512), .C2(u4_srl_451_n64), .A(u4_srl_451_n513), .ZN(
        u4_srl_451_n203) );
  INV_X1 u4_srl_451_U412 ( .A(u4_srl_451_n203), .ZN(u4_srl_451_n493) );
  INV_X1 u4_srl_451_U411 ( .A(u4_srl_451_n510), .ZN(u4_srl_451_n506) );
  AOI22_X1 u4_srl_451_U410 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n508), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n509), .ZN(u4_srl_451_n507) );
  OAI221_X1 u4_srl_451_U409 ( .B1(u4_srl_451_n505), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n506), .C2(u4_srl_451_n64), .A(u4_srl_451_n507), .ZN(
        u4_srl_451_n387) );
  AOI22_X1 u4_srl_451_U408 ( .A1(u4_srl_451_n24), .A2(u4_srl_451_n503), .B1(
        u4_srl_451_n30), .B2(u4_srl_451_n504), .ZN(u4_srl_451_n502) );
  OAI221_X1 u4_srl_451_U407 ( .B1(u4_srl_451_n500), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n501), .C2(u4_srl_451_n64), .A(u4_srl_451_n502), .ZN(
        u4_srl_451_n386) );
  INV_X1 u4_srl_451_U406 ( .A(u4_srl_451_n386), .ZN(u4_srl_451_n250) );
  OAI22_X1 u4_srl_451_U405 ( .A1(u4_shift_right[4]), .A2(u4_srl_451_n250), 
        .B1(u4_srl_451_n249), .B2(u4_srl_451_n468), .ZN(u4_srl_451_n307) );
  AOI22_X1 u4_srl_451_U404 ( .A1(u4_srl_451_n22), .A2(u4_srl_451_n498), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n499), .ZN(u4_srl_451_n497) );
  OAI221_X1 u4_srl_451_U403 ( .B1(u4_srl_451_n495), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n496), .C2(u4_srl_451_n64), .A(u4_srl_451_n497), .ZN(
        u4_srl_451_n308) );
  AOI222_X1 u4_srl_451_U402 ( .A1(u4_srl_451_n14), .A2(u4_srl_451_n387), .B1(
        u4_srl_451_n462), .B2(u4_srl_451_n307), .C1(u4_srl_451_n317), .C2(
        u4_srl_451_n308), .ZN(u4_srl_451_n494) );
  OAI221_X1 u4_srl_451_U401 ( .B1(u4_srl_451_n207), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n493), .C2(u4_srl_451_n9), .A(u4_srl_451_n494), .ZN(
        u4_N5924) );
  AOI22_X1 u4_srl_451_U400 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n491), .B1(
        u4_srl_451_n27), .B2(u4_srl_451_n492), .ZN(u4_srl_451_n490) );
  INV_X1 u4_srl_451_U399 ( .A(u4_srl_451_n490), .ZN(u4_srl_451_n489) );
  AOI221_X1 u4_srl_451_U398 ( .B1(u4_srl_451_n487), .B2(u4_srl_451_n16), .C1(
        u4_srl_451_n488), .C2(u4_srl_451_n60), .A(u4_srl_451_n489), .ZN(
        u4_srl_451_n183) );
  INV_X1 u4_srl_451_U397 ( .A(u4_srl_451_n486), .ZN(u4_srl_451_n481) );
  AOI22_X1 u4_srl_451_U396 ( .A1(u4_srl_451_n21), .A2(u4_srl_451_n484), .B1(
        u4_srl_451_n26), .B2(u4_srl_451_n485), .ZN(u4_srl_451_n483) );
  OAI221_X1 u4_srl_451_U395 ( .B1(u4_srl_451_n481), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n482), .C2(u4_srl_451_n64), .A(u4_srl_451_n483), .ZN(
        u4_srl_451_n177) );
  INV_X1 u4_srl_451_U394 ( .A(u4_srl_451_n177), .ZN(u4_srl_451_n459) );
  AOI22_X1 u4_srl_451_U393 ( .A1(u4_srl_451_n23), .A2(u4_srl_451_n479), .B1(
        u4_srl_451_n26), .B2(u4_srl_451_n480), .ZN(u4_srl_451_n478) );
  INV_X1 u4_srl_451_U392 ( .A(u4_srl_451_n478), .ZN(u4_srl_451_n477) );
  AOI221_X1 u4_srl_451_U391 ( .B1(u4_srl_451_n475), .B2(u4_srl_451_n17), .C1(
        u4_srl_451_n476), .C2(u4_srl_451_n60), .A(u4_srl_451_n477), .ZN(
        u4_srl_451_n181) );
  INV_X1 u4_srl_451_U390 ( .A(u4_srl_451_n181), .ZN(u4_srl_451_n461) );
  AOI22_X1 u4_srl_451_U389 ( .A1(u4_srl_451_n24), .A2(u4_srl_451_n473), .B1(
        u4_srl_451_n30), .B2(u4_srl_451_n474), .ZN(u4_srl_451_n472) );
  INV_X1 u4_srl_451_U388 ( .A(u4_srl_451_n472), .ZN(u4_srl_451_n471) );
  AOI221_X1 u4_srl_451_U387 ( .B1(u4_srl_451_n469), .B2(u4_srl_451_n16), .C1(
        u4_srl_451_n470), .C2(u4_srl_451_n60), .A(u4_srl_451_n471), .ZN(
        u4_srl_451_n246) );
  OAI22_X1 u4_srl_451_U386 ( .A1(u4_srl_451_n246), .A2(u4_shift_right[4]), 
        .B1(u4_srl_451_n245), .B2(u4_srl_451_n468), .ZN(u4_srl_451_n305) );
  AOI22_X1 u4_srl_451_U385 ( .A1(u4_srl_451_n22), .A2(u4_srl_451_n466), .B1(
        u4_srl_451_n26), .B2(u4_srl_451_n467), .ZN(u4_srl_451_n465) );
  OAI221_X1 u4_srl_451_U384 ( .B1(u4_srl_451_n463), .B2(u4_srl_451_n20), .C1(
        u4_srl_451_n464), .C2(u4_srl_451_n64), .A(u4_srl_451_n465), .ZN(
        u4_srl_451_n306) );
  AOI222_X1 u4_srl_451_U383 ( .A1(u4_srl_451_n14), .A2(u4_srl_451_n461), .B1(
        u4_srl_451_n462), .B2(u4_srl_451_n305), .C1(u4_srl_451_n317), .C2(
        u4_srl_451_n306), .ZN(u4_srl_451_n460) );
  OAI221_X1 u4_srl_451_U382 ( .B1(u4_srl_451_n183), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n459), .C2(u4_srl_451_n9), .A(u4_srl_451_n460), .ZN(
        u4_N5925) );
  INV_X1 u4_srl_451_U381 ( .A(u4_srl_451_n303), .ZN(u4_srl_451_n458) );
  INV_X1 u4_srl_451_U380 ( .A(u4_srl_451_n195), .ZN(u4_srl_451_n375) );
  AOI222_X1 u4_srl_451_U379 ( .A1(u4_srl_451_n14), .A2(u4_srl_451_n458), .B1(
        u4_srl_451_n13), .B2(u4_srl_451_n376), .C1(u4_srl_451_n413), .C2(
        u4_srl_451_n375), .ZN(u4_srl_451_n457) );
  OAI221_X1 u4_srl_451_U378 ( .B1(u4_srl_451_n378), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n456), .C2(u4_srl_451_n9), .A(u4_srl_451_n457), .ZN(
        u4_N5926) );
  INV_X1 u4_srl_451_U377 ( .A(u4_srl_451_n301), .ZN(u4_srl_451_n455) );
  INV_X1 u4_srl_451_U376 ( .A(u4_srl_451_n194), .ZN(u4_srl_451_n370) );
  AOI222_X1 u4_srl_451_U375 ( .A1(u4_srl_451_n14), .A2(u4_srl_451_n455), .B1(
        u4_srl_451_n13), .B2(u4_srl_451_n371), .C1(u4_srl_451_n413), .C2(
        u4_srl_451_n370), .ZN(u4_srl_451_n454) );
  OAI221_X1 u4_srl_451_U374 ( .B1(u4_srl_451_n373), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n453), .C2(u4_srl_451_n9), .A(u4_srl_451_n454), .ZN(
        u4_N5927) );
  AOI222_X1 u4_srl_451_U373 ( .A1(u4_srl_451_n14), .A2(u4_srl_451_n452), .B1(
        u4_srl_451_n13), .B2(u4_srl_451_n366), .C1(u4_srl_451_n413), .C2(
        u4_srl_451_n365), .ZN(u4_srl_451_n451) );
  OAI221_X1 u4_srl_451_U372 ( .B1(u4_srl_451_n368), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n450), .C2(u4_srl_451_n9), .A(u4_srl_451_n451), .ZN(
        u4_N5928) );
  INV_X1 u4_srl_451_U371 ( .A(u4_srl_451_n283), .ZN(u4_srl_451_n449) );
  INV_X1 u4_srl_451_U370 ( .A(u4_srl_451_n192), .ZN(u4_srl_451_n360) );
  AOI222_X1 u4_srl_451_U369 ( .A1(u4_srl_451_n14), .A2(u4_srl_451_n449), .B1(
        u4_srl_451_n13), .B2(u4_srl_451_n361), .C1(u4_srl_451_n413), .C2(
        u4_srl_451_n360), .ZN(u4_srl_451_n448) );
  OAI221_X1 u4_srl_451_U368 ( .B1(u4_srl_451_n363), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n447), .C2(u4_srl_451_n9), .A(u4_srl_451_n448), .ZN(
        u4_N5929) );
  AOI222_X1 u4_srl_451_U367 ( .A1(u4_srl_451_n421), .A2(u4_srl_451_n405), .B1(
        u4_srl_451_n328), .B2(u4_srl_451_n341), .C1(u4_srl_451_n329), .C2(
        u4_srl_451_n406), .ZN(u4_srl_451_n275) );
  INV_X1 u4_srl_451_U366 ( .A(u4_srl_451_n419), .ZN(u4_srl_451_n439) );
  OAI22_X1 u4_srl_451_U365 ( .A1(u4_srl_451_n40), .A2(u4_srl_451_n65), .B1(
        u4_srl_451_n31), .B2(u4_srl_451_n66), .ZN(u4_srl_451_n446) );
  AOI221_X1 u4_srl_451_U364 ( .B1(fract_denorm[5]), .B2(u4_srl_451_n47), .C1(
        fract_denorm[4]), .C2(u4_srl_451_n55), .A(u4_srl_451_n446), .ZN(
        u4_srl_451_n441) );
  AOI22_X1 u4_srl_451_U363 ( .A1(fract_denorm[9]), .A2(u4_srl_451_n47), .B1(
        fract_denorm[8]), .B2(u4_srl_451_n55), .ZN(u4_srl_451_n445) );
  OAI221_X1 u4_srl_451_U362 ( .B1(u4_srl_451_n31), .B2(u4_srl_451_n70), .C1(
        u4_srl_451_n40), .C2(u4_srl_451_n69), .A(u4_srl_451_n445), .ZN(
        u4_srl_451_n261) );
  AOI222_X1 u4_srl_451_U361 ( .A1(u4_srl_451_n16), .A2(u4_srl_451_n261), .B1(
        u4_srl_451_n21), .B2(u4_srl_451_n258), .C1(u4_srl_451_n26), .C2(
        u4_srl_451_n262), .ZN(u4_srl_451_n444) );
  MUX2_X1 u4_srl_451_U360 ( .A(u4_srl_451_n443), .B(u4_srl_451_n444), .S(
        u4_srl_451_n397), .Z(u4_srl_451_n442) );
  OAI21_X1 u4_srl_451_U359 ( .B1(u4_srl_451_n441), .B2(u4_srl_451_n270), .A(
        u4_srl_451_n442), .ZN(u4_srl_451_n440) );
  AOI22_X1 u4_srl_451_U358 ( .A1(u4_srl_451_n15), .A2(u4_srl_451_n439), .B1(
        u4_srl_451_n391), .B2(u4_srl_451_n440), .ZN(u4_srl_451_n438) );
  OAI221_X1 u4_srl_451_U357 ( .B1(u4_srl_451_n275), .B2(u4_srl_451_n388), .C1(
        u4_srl_451_n326), .C2(u4_srl_451_n12), .A(u4_srl_451_n438), .ZN(
        u4_N5902) );
  INV_X1 u4_srl_451_U356 ( .A(u4_srl_451_n281), .ZN(u4_srl_451_n435) );
  INV_X1 u4_srl_451_U355 ( .A(u4_srl_451_n191), .ZN(u4_srl_451_n437) );
  AOI222_X1 u4_srl_451_U354 ( .A1(u4_srl_451_n14), .A2(u4_srl_451_n435), .B1(
        u4_srl_451_n13), .B2(u4_srl_451_n436), .C1(u4_srl_451_n413), .C2(
        u4_srl_451_n437), .ZN(u4_srl_451_n434) );
  OAI221_X1 u4_srl_451_U353 ( .B1(u4_srl_451_n358), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n433), .C2(u4_srl_451_n9), .A(u4_srl_451_n434), .ZN(
        u4_N5930) );
  INV_X1 u4_srl_451_U352 ( .A(u4_srl_451_n190), .ZN(u4_srl_451_n432) );
  AOI222_X1 u4_srl_451_U351 ( .A1(u4_srl_451_n15), .A2(u4_srl_451_n430), .B1(
        u4_srl_451_n13), .B2(u4_srl_451_n431), .C1(u4_srl_451_n413), .C2(
        u4_srl_451_n432), .ZN(u4_srl_451_n429) );
  OAI221_X1 u4_srl_451_U350 ( .B1(u4_srl_451_n355), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n428), .C2(u4_srl_451_n9), .A(u4_srl_451_n429), .ZN(
        u4_N5931) );
  AOI222_X1 u4_srl_451_U349 ( .A1(u4_srl_451_n14), .A2(u4_srl_451_n427), .B1(
        u4_srl_451_n13), .B2(u4_srl_451_n352), .C1(u4_srl_451_n413), .C2(
        u4_srl_451_n351), .ZN(u4_srl_451_n426) );
  OAI221_X1 u4_srl_451_U348 ( .B1(u4_srl_451_n349), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n425), .C2(u4_srl_451_n9), .A(u4_srl_451_n426), .ZN(
        u4_N5932) );
  AOI222_X1 u4_srl_451_U347 ( .A1(u4_srl_451_n15), .A2(u4_srl_451_n424), .B1(
        u4_srl_451_n13), .B2(u4_srl_451_n347), .C1(u4_srl_451_n413), .C2(
        u4_srl_451_n346), .ZN(u4_srl_451_n423) );
  OAI221_X1 u4_srl_451_U346 ( .B1(u4_srl_451_n344), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n422), .C2(u4_srl_451_n9), .A(u4_srl_451_n423), .ZN(
        u4_N5933) );
  AOI222_X1 u4_srl_451_U345 ( .A1(u4_srl_451_n15), .A2(u4_srl_451_n421), .B1(
        u4_srl_451_n13), .B2(u4_srl_451_n329), .C1(u4_srl_451_n413), .C2(
        u4_srl_451_n328), .ZN(u4_srl_451_n420) );
  OAI221_X1 u4_srl_451_U344 ( .B1(u4_srl_451_n326), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n419), .C2(u4_srl_451_n9), .A(u4_srl_451_n420), .ZN(
        u4_N5934) );
  AOI222_X1 u4_srl_451_U343 ( .A1(u4_srl_451_n14), .A2(u4_srl_451_n404), .B1(
        u4_srl_451_n13), .B2(u4_srl_451_n324), .C1(u4_srl_451_n413), .C2(
        u4_srl_451_n323), .ZN(u4_srl_451_n418) );
  OAI221_X1 u4_srl_451_U342 ( .B1(u4_srl_451_n321), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n403), .C2(u4_srl_451_n9), .A(u4_srl_451_n418), .ZN(
        u4_N5935) );
  INV_X1 u4_srl_451_U341 ( .A(u4_srl_451_n339), .ZN(u4_srl_451_n318) );
  AOI222_X1 u4_srl_451_U340 ( .A1(u4_srl_451_n14), .A2(u4_srl_451_n342), .B1(
        u4_srl_451_n13), .B2(u4_srl_451_n319), .C1(u4_srl_451_n413), .C2(
        u4_srl_451_n318), .ZN(u4_srl_451_n417) );
  OAI221_X1 u4_srl_451_U339 ( .B1(u4_srl_451_n315), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n338), .C2(u4_srl_451_n9), .A(u4_srl_451_n417), .ZN(
        u4_N5936) );
  INV_X1 u4_srl_451_U338 ( .A(u4_srl_451_n297), .ZN(u4_srl_451_n415) );
  INV_X1 u4_srl_451_U337 ( .A(u4_srl_451_n299), .ZN(u4_srl_451_n416) );
  AOI222_X1 u4_srl_451_U336 ( .A1(u4_srl_451_n15), .A2(u4_srl_451_n313), .B1(
        u4_srl_451_n413), .B2(u4_srl_451_n415), .C1(u4_srl_451_n13), .C2(
        u4_srl_451_n416), .ZN(u4_srl_451_n414) );
  OAI221_X1 u4_srl_451_U335 ( .B1(u4_srl_451_n294), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n295), .C2(u4_srl_451_n9), .A(u4_srl_451_n414), .ZN(
        u4_N5937) );
  AND2_X1 u4_srl_451_U334 ( .A1(u4_srl_451_n413), .A2(u4_srl_451_n61), .ZN(
        u4_srl_451_n384) );
  INV_X1 u4_srl_451_U333 ( .A(u4_srl_451_n269), .ZN(u4_srl_451_n412) );
  AOI222_X1 u4_srl_451_U332 ( .A1(u4_srl_451_n15), .A2(u4_srl_451_n312), .B1(
        u4_srl_451_n384), .B2(u4_srl_451_n411), .C1(u4_srl_451_n13), .C2(
        u4_srl_451_n412), .ZN(u4_srl_451_n410) );
  OAI221_X1 u4_srl_451_U331 ( .B1(u4_srl_451_n265), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n266), .C2(u4_srl_451_n9), .A(u4_srl_451_n410), .ZN(
        u4_N5938) );
  INV_X1 u4_srl_451_U330 ( .A(u4_srl_451_n253), .ZN(u4_srl_451_n409) );
  AOI222_X1 u4_srl_451_U329 ( .A1(u4_srl_451_n14), .A2(u4_srl_451_n310), .B1(
        u4_srl_451_n384), .B2(u4_srl_451_n408), .C1(u4_srl_451_n13), .C2(
        u4_srl_451_n409), .ZN(u4_srl_451_n407) );
  OAI221_X1 u4_srl_451_U328 ( .B1(u4_srl_451_n234), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n235), .C2(u4_srl_451_n9), .A(u4_srl_451_n407), .ZN(
        u4_N5939) );
  AOI222_X1 u4_srl_451_U327 ( .A1(u4_srl_451_n404), .A2(u4_srl_451_n405), .B1(
        u4_srl_451_n323), .B2(u4_srl_451_n341), .C1(u4_srl_451_n324), .C2(
        u4_srl_451_n406), .ZN(u4_srl_451_n274) );
  INV_X1 u4_srl_451_U326 ( .A(u4_srl_451_n403), .ZN(u4_srl_451_n390) );
  OAI22_X1 u4_srl_451_U325 ( .A1(u4_srl_451_n40), .A2(u4_srl_451_n66), .B1(
        u4_srl_451_n31), .B2(u4_srl_451_n67), .ZN(u4_srl_451_n402) );
  AOI221_X1 u4_srl_451_U324 ( .B1(fract_denorm[6]), .B2(u4_srl_451_n47), .C1(
        fract_denorm[5]), .C2(u4_srl_451_n55), .A(u4_srl_451_n402), .ZN(
        u4_srl_451_n393) );
  AOI22_X1 u4_srl_451_U323 ( .A1(fract_denorm[10]), .A2(u4_srl_451_n49), .B1(
        fract_denorm[9]), .B2(u4_srl_451_n52), .ZN(u4_srl_451_n401) );
  OAI221_X1 u4_srl_451_U322 ( .B1(u4_srl_451_n34), .B2(u4_srl_451_n71), .C1(
        u4_srl_451_n43), .C2(u4_srl_451_n70), .A(u4_srl_451_n401), .ZN(
        u4_srl_451_n229) );
  AOI222_X1 u4_srl_451_U321 ( .A1(u4_srl_451_n16), .A2(u4_srl_451_n229), .B1(
        u4_srl_451_n21), .B2(u4_srl_451_n226), .C1(u4_srl_451_n26), .C2(
        u4_srl_451_n230), .ZN(u4_srl_451_n396) );
  MUX2_X1 u4_srl_451_U320 ( .A(u4_srl_451_n395), .B(u4_srl_451_n396), .S(
        u4_srl_451_n397), .Z(u4_srl_451_n394) );
  OAI21_X1 u4_srl_451_U319 ( .B1(u4_srl_451_n393), .B2(u4_srl_451_n270), .A(
        u4_srl_451_n394), .ZN(u4_srl_451_n392) );
  AOI22_X1 u4_srl_451_U318 ( .A1(u4_srl_451_n15), .A2(u4_srl_451_n390), .B1(
        u4_srl_451_n391), .B2(u4_srl_451_n392), .ZN(u4_srl_451_n389) );
  OAI221_X1 u4_srl_451_U317 ( .B1(u4_srl_451_n274), .B2(u4_srl_451_n388), .C1(
        u4_srl_451_n321), .C2(u4_srl_451_n12), .A(u4_srl_451_n389), .ZN(
        u4_N5903) );
  INV_X1 u4_srl_451_U316 ( .A(u4_srl_451_n387), .ZN(u4_srl_451_n206) );
  AOI222_X1 u4_srl_451_U315 ( .A1(u4_srl_451_n15), .A2(u4_srl_451_n308), .B1(
        u4_srl_451_n384), .B2(u4_srl_451_n385), .C1(u4_srl_451_n13), .C2(
        u4_srl_451_n386), .ZN(u4_srl_451_n383) );
  OAI221_X1 u4_srl_451_U314 ( .B1(u4_srl_451_n206), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n207), .C2(u4_srl_451_n9), .A(u4_srl_451_n383), .ZN(
        u4_N5940) );
  INV_X1 u4_srl_451_U313 ( .A(u4_srl_451_n246), .ZN(u4_srl_451_n382) );
  AOI222_X1 u4_srl_451_U312 ( .A1(u4_srl_451_n14), .A2(u4_srl_451_n306), .B1(
        u4_srl_451_n380), .B2(u4_srl_451_n381), .C1(u4_srl_451_n317), .C2(
        u4_srl_451_n382), .ZN(u4_srl_451_n379) );
  OAI221_X1 u4_srl_451_U311 ( .B1(u4_srl_451_n181), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n183), .C2(u4_srl_451_n9), .A(u4_srl_451_n379), .ZN(
        u4_N5941) );
  OAI22_X1 u4_srl_451_U310 ( .A1(u4_srl_451_n11), .A2(u4_srl_451_n303), .B1(
        u4_srl_451_n9), .B2(u4_srl_451_n378), .ZN(u4_srl_451_n377) );
  AOI221_X1 u4_srl_451_U309 ( .B1(u4_srl_451_n375), .B2(u4_srl_451_n317), .C1(
        u4_srl_451_n376), .C2(u4_srl_451_n15), .A(u4_srl_451_n377), .ZN(
        u4_srl_451_n374) );
  INV_X1 u4_srl_451_U308 ( .A(u4_srl_451_n374), .ZN(u4_N5942) );
  OAI22_X1 u4_srl_451_U307 ( .A1(u4_srl_451_n10), .A2(u4_srl_451_n301), .B1(
        u4_srl_451_n9), .B2(u4_srl_451_n373), .ZN(u4_srl_451_n372) );
  AOI221_X1 u4_srl_451_U306 ( .B1(u4_srl_451_n370), .B2(u4_srl_451_n317), .C1(
        u4_srl_451_n371), .C2(u4_srl_451_n15), .A(u4_srl_451_n372), .ZN(
        u4_srl_451_n369) );
  INV_X1 u4_srl_451_U305 ( .A(u4_srl_451_n369), .ZN(u4_N5943) );
  OAI22_X1 u4_srl_451_U304 ( .A1(u4_srl_451_n11), .A2(u4_srl_451_n285), .B1(
        u4_srl_451_n9), .B2(u4_srl_451_n368), .ZN(u4_srl_451_n367) );
  AOI221_X1 u4_srl_451_U303 ( .B1(u4_srl_451_n365), .B2(u4_srl_451_n317), .C1(
        u4_srl_451_n366), .C2(u4_srl_451_n15), .A(u4_srl_451_n367), .ZN(
        u4_srl_451_n364) );
  INV_X1 u4_srl_451_U302 ( .A(u4_srl_451_n364), .ZN(u4_N5944) );
  OAI22_X1 u4_srl_451_U301 ( .A1(u4_srl_451_n10), .A2(u4_srl_451_n283), .B1(
        u4_srl_451_n9), .B2(u4_srl_451_n363), .ZN(u4_srl_451_n362) );
  AOI221_X1 u4_srl_451_U300 ( .B1(u4_srl_451_n360), .B2(u4_srl_451_n317), .C1(
        u4_srl_451_n361), .C2(u4_srl_451_n15), .A(u4_srl_451_n362), .ZN(
        u4_srl_451_n359) );
  INV_X1 u4_srl_451_U299 ( .A(u4_srl_451_n359), .ZN(u4_N5945) );
  OAI22_X1 u4_srl_451_U298 ( .A1(u4_srl_451_n10), .A2(u4_srl_451_n281), .B1(
        u4_srl_451_n9), .B2(u4_srl_451_n358), .ZN(u4_srl_451_n357) );
  INV_X1 u4_srl_451_U297 ( .A(u4_srl_451_n357), .ZN(u4_srl_451_n356) );
  OAI221_X1 u4_srl_451_U296 ( .B1(u4_srl_451_n191), .B2(u4_srl_451_n12), .C1(
        u4_srl_451_n280), .C2(u4_srl_451_n3), .A(u4_srl_451_n356), .ZN(
        u4_N5946) );
  OAI22_X1 u4_srl_451_U295 ( .A1(u4_srl_451_n10), .A2(u4_srl_451_n279), .B1(
        u4_srl_451_n9), .B2(u4_srl_451_n355), .ZN(u4_srl_451_n354) );
  INV_X1 u4_srl_451_U294 ( .A(u4_srl_451_n354), .ZN(u4_srl_451_n353) );
  OAI221_X1 u4_srl_451_U293 ( .B1(u4_srl_451_n190), .B2(u4_srl_451_n12), .C1(
        u4_srl_451_n278), .C2(u4_srl_451_n3), .A(u4_srl_451_n353), .ZN(
        u4_N5947) );
  AOI22_X1 u4_srl_451_U292 ( .A1(u4_srl_451_n13), .A2(u4_srl_451_n351), .B1(
        u4_srl_451_n15), .B2(u4_srl_451_n352), .ZN(u4_srl_451_n350) );
  OAI221_X1 u4_srl_451_U291 ( .B1(u4_srl_451_n348), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n349), .C2(u4_srl_451_n9), .A(u4_srl_451_n350), .ZN(
        u4_N5948) );
  AOI22_X1 u4_srl_451_U290 ( .A1(u4_srl_451_n13), .A2(u4_srl_451_n346), .B1(
        u4_srl_451_n15), .B2(u4_srl_451_n347), .ZN(u4_srl_451_n345) );
  OAI221_X1 u4_srl_451_U289 ( .B1(u4_srl_451_n343), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n344), .C2(u4_srl_451_n9), .A(u4_srl_451_n345), .ZN(
        u4_N5949) );
  INV_X1 u4_srl_451_U288 ( .A(u4_srl_451_n342), .ZN(u4_srl_451_n314) );
  INV_X1 u4_srl_451_U287 ( .A(u4_srl_451_n341), .ZN(u4_srl_451_n298) );
  OAI222_X1 u4_srl_451_U286 ( .A1(u4_srl_451_n314), .A2(u4_srl_451_n243), .B1(
        u4_srl_451_n339), .B2(u4_srl_451_n298), .C1(u4_srl_451_n340), .C2(
        u4_srl_451_n247), .ZN(u4_srl_451_n273) );
  OAI22_X1 u4_srl_451_U285 ( .A1(u4_srl_451_n315), .A2(u4_srl_451_n182), .B1(
        u4_srl_451_n338), .B2(u4_srl_451_n184), .ZN(u4_srl_451_n337) );
  AOI221_X1 u4_srl_451_U284 ( .B1(u4_srl_451_n176), .B2(u4_srl_451_n336), .C1(
        u4_srl_451_n273), .C2(u4_srl_451_n179), .A(u4_srl_451_n337), .ZN(
        u4_srl_451_n330) );
  INV_X1 u4_srl_451_U283 ( .A(u4_srl_451_n175), .ZN(u4_srl_451_n223) );
  INV_X1 u4_srl_451_U282 ( .A(u4_srl_451_n173), .ZN(u4_srl_451_n225) );
  AOI22_X1 u4_srl_451_U281 ( .A1(u4_srl_451_n335), .A2(u4_srl_451_n169), .B1(
        u4_srl_451_n199), .B2(u4_srl_451_n167), .ZN(u4_srl_451_n334) );
  INV_X1 u4_srl_451_U280 ( .A(u4_srl_451_n334), .ZN(u4_srl_451_n333) );
  AOI221_X1 u4_srl_451_U279 ( .B1(u4_srl_451_n223), .B2(u4_srl_451_n332), .C1(
        u4_srl_451_n225), .C2(u4_srl_451_n198), .A(u4_srl_451_n333), .ZN(
        u4_srl_451_n331) );
  AOI21_X1 u4_srl_451_U278 ( .B1(u4_srl_451_n330), .B2(u4_srl_451_n331), .A(
        u4_shift_right[8]), .ZN(u4_N5904) );
  AOI22_X1 u4_srl_451_U277 ( .A1(u4_srl_451_n13), .A2(u4_srl_451_n328), .B1(
        u4_srl_451_n15), .B2(u4_srl_451_n329), .ZN(u4_srl_451_n327) );
  OAI221_X1 u4_srl_451_U276 ( .B1(u4_srl_451_n325), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n326), .C2(u4_srl_451_n9), .A(u4_srl_451_n327), .ZN(
        u4_N5950) );
  AOI22_X1 u4_srl_451_U275 ( .A1(u4_srl_451_n13), .A2(u4_srl_451_n323), .B1(
        u4_srl_451_n15), .B2(u4_srl_451_n324), .ZN(u4_srl_451_n322) );
  OAI221_X1 u4_srl_451_U274 ( .B1(u4_srl_451_n320), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n321), .C2(u4_srl_451_n9), .A(u4_srl_451_n322), .ZN(
        u4_N5951) );
  AOI22_X1 u4_srl_451_U273 ( .A1(u4_srl_451_n13), .A2(u4_srl_451_n318), .B1(
        u4_srl_451_n15), .B2(u4_srl_451_n319), .ZN(u4_srl_451_n316) );
  OAI221_X1 u4_srl_451_U272 ( .B1(u4_srl_451_n314), .B2(u4_srl_451_n10), .C1(
        u4_srl_451_n315), .C2(u4_srl_451_n9), .A(u4_srl_451_n316), .ZN(
        u4_N5952) );
  INV_X1 u4_srl_451_U271 ( .A(u4_srl_451_n313), .ZN(u4_srl_451_n296) );
  OAI222_X1 u4_srl_451_U270 ( .A1(u4_srl_451_n294), .A2(u4_srl_451_n186), .B1(
        u4_srl_451_n296), .B2(u4_srl_451_n10), .C1(u4_srl_451_n213), .C2(
        u4_srl_451_n304), .ZN(u4_N5953) );
  INV_X1 u4_srl_451_U269 ( .A(u4_srl_451_n312), .ZN(u4_srl_451_n267) );
  INV_X1 u4_srl_451_U268 ( .A(u4_srl_451_n311), .ZN(u4_srl_451_n212) );
  OAI222_X1 u4_srl_451_U267 ( .A1(u4_srl_451_n265), .A2(u4_srl_451_n186), .B1(
        u4_srl_451_n267), .B2(u4_srl_451_n11), .C1(u4_srl_451_n212), .C2(
        u4_srl_451_n304), .ZN(u4_N5954) );
  INV_X1 u4_srl_451_U266 ( .A(u4_srl_451_n310), .ZN(u4_srl_451_n251) );
  INV_X1 u4_srl_451_U265 ( .A(u4_srl_451_n309), .ZN(u4_srl_451_n211) );
  OAI222_X1 u4_srl_451_U264 ( .A1(u4_srl_451_n234), .A2(u4_srl_451_n186), .B1(
        u4_srl_451_n251), .B2(u4_srl_451_n11), .C1(u4_srl_451_n211), .C2(
        u4_srl_451_n304), .ZN(u4_N5955) );
  INV_X1 u4_srl_451_U263 ( .A(u4_srl_451_n308), .ZN(u4_srl_451_n248) );
  INV_X1 u4_srl_451_U262 ( .A(u4_srl_451_n307), .ZN(u4_srl_451_n210) );
  OAI222_X1 u4_srl_451_U261 ( .A1(u4_srl_451_n206), .A2(u4_srl_451_n186), .B1(
        u4_srl_451_n248), .B2(u4_srl_451_n11), .C1(u4_srl_451_n210), .C2(
        u4_srl_451_n304), .ZN(u4_N5956) );
  INV_X1 u4_srl_451_U260 ( .A(u4_srl_451_n306), .ZN(u4_srl_451_n242) );
  INV_X1 u4_srl_451_U259 ( .A(u4_srl_451_n305), .ZN(u4_srl_451_n208) );
  OAI222_X1 u4_srl_451_U258 ( .A1(u4_srl_451_n181), .A2(u4_srl_451_n186), .B1(
        u4_srl_451_n242), .B2(u4_srl_451_n10), .C1(u4_srl_451_n208), .C2(
        u4_srl_451_n304), .ZN(u4_N5957) );
  OAI222_X1 u4_srl_451_U257 ( .A1(u4_srl_451_n302), .A2(u4_srl_451_n11), .B1(
        u4_srl_451_n195), .B2(u4_srl_451_n3), .C1(u4_srl_451_n303), .C2(
        u4_srl_451_n9), .ZN(u4_N5958) );
  OAI222_X1 u4_srl_451_U256 ( .A1(u4_srl_451_n300), .A2(u4_srl_451_n11), .B1(
        u4_srl_451_n194), .B2(u4_srl_451_n3), .C1(u4_srl_451_n301), .C2(
        u4_srl_451_n186), .ZN(u4_N5959) );
  OAI222_X1 u4_srl_451_U255 ( .A1(u4_srl_451_n296), .A2(u4_srl_451_n243), .B1(
        u4_srl_451_n297), .B2(u4_srl_451_n298), .C1(u4_srl_451_n299), .C2(
        u4_srl_451_n247), .ZN(u4_srl_451_n272) );
  OAI22_X1 u4_srl_451_U254 ( .A1(u4_srl_451_n294), .A2(u4_srl_451_n182), .B1(
        u4_srl_451_n295), .B2(u4_srl_451_n184), .ZN(u4_srl_451_n293) );
  AOI221_X1 u4_srl_451_U253 ( .B1(u4_srl_451_n176), .B2(u4_srl_451_n292), .C1(
        u4_srl_451_n272), .C2(u4_srl_451_n179), .A(u4_srl_451_n293), .ZN(
        u4_srl_451_n286) );
  AOI22_X1 u4_srl_451_U252 ( .A1(u4_srl_451_n291), .A2(u4_srl_451_n169), .B1(
        u4_srl_451_n170), .B2(u4_srl_451_n167), .ZN(u4_srl_451_n290) );
  INV_X1 u4_srl_451_U251 ( .A(u4_srl_451_n290), .ZN(u4_srl_451_n289) );
  AOI221_X1 u4_srl_451_U250 ( .B1(u4_srl_451_n223), .B2(u4_srl_451_n288), .C1(
        u4_srl_451_n225), .C2(u4_srl_451_n168), .A(u4_srl_451_n289), .ZN(
        u4_srl_451_n287) );
  AOI21_X1 u4_srl_451_U249 ( .B1(u4_srl_451_n286), .B2(u4_srl_451_n287), .A(
        u4_shift_right[8]), .ZN(u4_N5905) );
  OAI222_X1 u4_srl_451_U248 ( .A1(u4_srl_451_n284), .A2(u4_srl_451_n11), .B1(
        u4_srl_451_n193), .B2(u4_srl_451_n3), .C1(u4_srl_451_n285), .C2(
        u4_srl_451_n186), .ZN(u4_N5960) );
  OAI222_X1 u4_srl_451_U247 ( .A1(u4_srl_451_n282), .A2(u4_srl_451_n11), .B1(
        u4_srl_451_n192), .B2(u4_srl_451_n3), .C1(u4_srl_451_n283), .C2(
        u4_srl_451_n9), .ZN(u4_N5961) );
  OAI222_X1 u4_srl_451_U246 ( .A1(u4_srl_451_n280), .A2(u4_srl_451_n11), .B1(
        u4_srl_451_n191), .B2(u4_srl_451_n3), .C1(u4_srl_451_n281), .C2(
        u4_srl_451_n186), .ZN(u4_N5962) );
  OAI222_X1 u4_srl_451_U245 ( .A1(u4_srl_451_n278), .A2(u4_srl_451_n11), .B1(
        u4_srl_451_n190), .B2(u4_srl_451_n3), .C1(u4_srl_451_n279), .C2(
        u4_srl_451_n186), .ZN(u4_N5963) );
  INV_X1 u4_srl_451_U244 ( .A(u4_srl_451_n215), .ZN(u4_srl_451_n217) );
  NOR2_X1 u4_srl_451_U243 ( .A1(u4_srl_451_n277), .A2(u4_srl_451_n217), .ZN(
        u4_N5964) );
  NOR2_X1 u4_srl_451_U242 ( .A1(u4_srl_451_n276), .A2(u4_srl_451_n217), .ZN(
        u4_N5965) );
  NOR2_X1 u4_srl_451_U241 ( .A1(u4_srl_451_n275), .A2(u4_srl_451_n217), .ZN(
        u4_N5966) );
  NOR2_X1 u4_srl_451_U240 ( .A1(u4_srl_451_n274), .A2(u4_srl_451_n217), .ZN(
        u4_N5967) );
  AND2_X1 u4_srl_451_U239 ( .A1(u4_srl_451_n273), .A2(u4_srl_451_n215), .ZN(
        u4_N5968) );
  AND2_X1 u4_srl_451_U238 ( .A1(u4_srl_451_n272), .A2(u4_srl_451_n215), .ZN(
        u4_N5969) );
  OR2_X1 u4_srl_451_U237 ( .A1(u4_srl_451_n270), .A2(u4_srl_451_n271), .ZN(
        u4_srl_451_n244) );
  OAI222_X1 u4_srl_451_U236 ( .A1(u4_srl_451_n267), .A2(u4_srl_451_n243), .B1(
        u4_srl_451_n268), .B2(u4_srl_451_n244), .C1(u4_srl_451_n269), .C2(
        u4_srl_451_n247), .ZN(u4_srl_451_n254) );
  OAI22_X1 u4_srl_451_U235 ( .A1(u4_srl_451_n265), .A2(u4_srl_451_n182), .B1(
        u4_srl_451_n266), .B2(u4_srl_451_n184), .ZN(u4_srl_451_n264) );
  AOI221_X1 u4_srl_451_U234 ( .B1(u4_srl_451_n176), .B2(u4_srl_451_n263), .C1(
        u4_srl_451_n254), .C2(u4_srl_451_n179), .A(u4_srl_451_n264), .ZN(
        u4_srl_451_n255) );
  AOI22_X1 u4_srl_451_U233 ( .A1(u4_srl_451_n261), .A2(u4_srl_451_n169), .B1(
        u4_srl_451_n262), .B2(u4_srl_451_n167), .ZN(u4_srl_451_n260) );
  INV_X1 u4_srl_451_U232 ( .A(u4_srl_451_n260), .ZN(u4_srl_451_n259) );
  AOI221_X1 u4_srl_451_U231 ( .B1(u4_srl_451_n223), .B2(u4_srl_451_n257), .C1(
        u4_srl_451_n225), .C2(u4_srl_451_n258), .A(u4_srl_451_n259), .ZN(
        u4_srl_451_n256) );
  AOI21_X1 u4_srl_451_U230 ( .B1(u4_srl_451_n255), .B2(u4_srl_451_n256), .A(
        u4_shift_right[8]), .ZN(u4_N5906) );
  AND2_X1 u4_srl_451_U229 ( .A1(u4_srl_451_n254), .A2(u4_srl_451_n215), .ZN(
        u4_N5970) );
  OAI222_X1 u4_srl_451_U228 ( .A1(u4_srl_451_n251), .A2(u4_srl_451_n243), .B1(
        u4_srl_451_n252), .B2(u4_srl_451_n244), .C1(u4_srl_451_n253), .C2(
        u4_srl_451_n247), .ZN(u4_srl_451_n232) );
  AND2_X1 u4_srl_451_U227 ( .A1(u4_srl_451_n232), .A2(u4_srl_451_n215), .ZN(
        u4_N5971) );
  OAI222_X1 u4_srl_451_U226 ( .A1(u4_srl_451_n248), .A2(u4_srl_451_n243), .B1(
        u4_srl_451_n249), .B2(u4_srl_451_n244), .C1(u4_srl_451_n250), .C2(
        u4_srl_451_n247), .ZN(u4_srl_451_n204) );
  AND2_X1 u4_srl_451_U225 ( .A1(u4_srl_451_n204), .A2(u4_srl_451_n215), .ZN(
        u4_N5972) );
  OAI222_X1 u4_srl_451_U224 ( .A1(u4_srl_451_n242), .A2(u4_srl_451_n243), .B1(
        u4_srl_451_n244), .B2(u4_srl_451_n245), .C1(u4_srl_451_n246), .C2(
        u4_srl_451_n247), .ZN(u4_srl_451_n178) );
  AND2_X1 u4_srl_451_U223 ( .A1(u4_srl_451_n178), .A2(u4_srl_451_n215), .ZN(
        u4_N5973) );
  AND2_X1 u4_srl_451_U222 ( .A1(u4_srl_451_n241), .A2(u4_srl_451_n215), .ZN(
        u4_N5974) );
  AND2_X1 u4_srl_451_U221 ( .A1(u4_srl_451_n240), .A2(u4_srl_451_n215), .ZN(
        u4_N5975) );
  AND2_X1 u4_srl_451_U220 ( .A1(u4_srl_451_n239), .A2(u4_srl_451_n215), .ZN(
        u4_N5976) );
  AND2_X1 u4_srl_451_U219 ( .A1(u4_srl_451_n238), .A2(u4_srl_451_n215), .ZN(
        u4_N5977) );
  AND2_X1 u4_srl_451_U218 ( .A1(u4_srl_451_n237), .A2(u4_srl_451_n215), .ZN(
        u4_N5978) );
  AND2_X1 u4_srl_451_U217 ( .A1(u4_srl_451_n236), .A2(u4_srl_451_n215), .ZN(
        u4_N5979) );
  OAI22_X1 u4_srl_451_U216 ( .A1(u4_srl_451_n234), .A2(u4_srl_451_n182), .B1(
        u4_srl_451_n235), .B2(u4_srl_451_n184), .ZN(u4_srl_451_n233) );
  AOI221_X1 u4_srl_451_U215 ( .B1(u4_srl_451_n176), .B2(u4_srl_451_n231), .C1(
        u4_srl_451_n232), .C2(u4_srl_451_n179), .A(u4_srl_451_n233), .ZN(
        u4_srl_451_n221) );
  AOI22_X1 u4_srl_451_U214 ( .A1(u4_srl_451_n229), .A2(u4_srl_451_n169), .B1(
        u4_srl_451_n230), .B2(u4_srl_451_n167), .ZN(u4_srl_451_n228) );
  INV_X1 u4_srl_451_U213 ( .A(u4_srl_451_n228), .ZN(u4_srl_451_n227) );
  AOI221_X1 u4_srl_451_U212 ( .B1(u4_srl_451_n223), .B2(u4_srl_451_n224), .C1(
        u4_srl_451_n225), .C2(u4_srl_451_n226), .A(u4_srl_451_n227), .ZN(
        u4_srl_451_n222) );
  AOI21_X1 u4_srl_451_U211 ( .B1(u4_srl_451_n221), .B2(u4_srl_451_n222), .A(
        u4_shift_right[8]), .ZN(u4_N5907) );
  NOR2_X1 u4_srl_451_U210 ( .A1(u4_srl_451_n220), .A2(u4_srl_451_n217), .ZN(
        u4_N5980) );
  NOR2_X1 u4_srl_451_U209 ( .A1(u4_srl_451_n219), .A2(u4_srl_451_n217), .ZN(
        u4_N5981) );
  NOR2_X1 u4_srl_451_U208 ( .A1(u4_srl_451_n218), .A2(u4_srl_451_n217), .ZN(
        u4_N5982) );
  NOR2_X1 u4_srl_451_U207 ( .A1(u4_srl_451_n216), .A2(u4_srl_451_n217), .ZN(
        u4_N5983) );
  AND2_X1 u4_srl_451_U206 ( .A1(u4_srl_451_n214), .A2(u4_srl_451_n215), .ZN(
        u4_N5984) );
  NOR2_X1 u4_srl_451_U205 ( .A1(u4_srl_451_n213), .A2(u4_srl_451_n209), .ZN(
        u4_N5985) );
  NOR2_X1 u4_srl_451_U204 ( .A1(u4_srl_451_n212), .A2(u4_srl_451_n209), .ZN(
        u4_N5986) );
  NOR2_X1 u4_srl_451_U203 ( .A1(u4_srl_451_n211), .A2(u4_srl_451_n209), .ZN(
        u4_N5987) );
  NOR2_X1 u4_srl_451_U202 ( .A1(u4_srl_451_n210), .A2(u4_srl_451_n209), .ZN(
        u4_N5988) );
  NOR2_X1 u4_srl_451_U201 ( .A1(u4_srl_451_n208), .A2(u4_srl_451_n209), .ZN(
        u4_N5989) );
  OAI22_X1 u4_srl_451_U200 ( .A1(u4_srl_451_n206), .A2(u4_srl_451_n182), .B1(
        u4_srl_451_n207), .B2(u4_srl_451_n184), .ZN(u4_srl_451_n205) );
  AOI221_X1 u4_srl_451_U199 ( .B1(u4_srl_451_n176), .B2(u4_srl_451_n203), .C1(
        u4_srl_451_n204), .C2(u4_srl_451_n179), .A(u4_srl_451_n205), .ZN(
        u4_srl_451_n196) );
  OAI22_X1 u4_srl_451_U198 ( .A1(u4_srl_451_n201), .A2(u4_srl_451_n173), .B1(
        u4_srl_451_n202), .B2(u4_srl_451_n175), .ZN(u4_srl_451_n200) );
  AOI221_X1 u4_srl_451_U197 ( .B1(u4_srl_451_n167), .B2(u4_srl_451_n198), .C1(
        u4_srl_451_n169), .C2(u4_srl_451_n199), .A(u4_srl_451_n200), .ZN(
        u4_srl_451_n197) );
  AOI21_X1 u4_srl_451_U196 ( .B1(u4_srl_451_n196), .B2(u4_srl_451_n197), .A(
        u4_shift_right[8]), .ZN(u4_N5908) );
  NOR2_X1 u4_srl_451_U195 ( .A1(u4_srl_451_n195), .A2(u4_srl_451_n9), .ZN(
        u4_N5990) );
  NOR2_X1 u4_srl_451_U194 ( .A1(u4_srl_451_n194), .A2(u4_srl_451_n9), .ZN(
        u4_N5991) );
  NOR2_X1 u4_srl_451_U193 ( .A1(u4_srl_451_n193), .A2(u4_srl_451_n9), .ZN(
        u4_N5992) );
  NOR2_X1 u4_srl_451_U192 ( .A1(u4_srl_451_n192), .A2(u4_srl_451_n9), .ZN(
        u4_N5993) );
  NOR2_X1 u4_srl_451_U191 ( .A1(u4_srl_451_n191), .A2(u4_srl_451_n9), .ZN(
        u4_N5994) );
  NOR2_X1 u4_srl_451_U190 ( .A1(u4_srl_451_n190), .A2(u4_srl_451_n9), .ZN(
        u4_N5995) );
  NOR2_X1 u4_srl_451_U189 ( .A1(u4_srl_451_n189), .A2(u4_srl_451_n9), .ZN(
        u4_N5996) );
  NOR2_X1 u4_srl_451_U188 ( .A1(u4_srl_451_n188), .A2(u4_srl_451_n9), .ZN(
        u4_N5997) );
  NOR2_X1 u4_srl_451_U187 ( .A1(u4_srl_451_n187), .A2(u4_srl_451_n9), .ZN(
        u4_N5998) );
  NOR2_X1 u4_srl_451_U186 ( .A1(u4_srl_451_n185), .A2(u4_srl_451_n9), .ZN(
        u4_N5999) );
  OAI22_X1 u4_srl_451_U185 ( .A1(u4_srl_451_n181), .A2(u4_srl_451_n182), .B1(
        u4_srl_451_n183), .B2(u4_srl_451_n184), .ZN(u4_srl_451_n180) );
  AOI221_X1 u4_srl_451_U184 ( .B1(u4_srl_451_n176), .B2(u4_srl_451_n177), .C1(
        u4_srl_451_n178), .C2(u4_srl_451_n179), .A(u4_srl_451_n180), .ZN(
        u4_srl_451_n165) );
  OAI22_X1 u4_srl_451_U183 ( .A1(u4_srl_451_n172), .A2(u4_srl_451_n173), .B1(
        u4_srl_451_n174), .B2(u4_srl_451_n175), .ZN(u4_srl_451_n171) );
  AOI221_X1 u4_srl_451_U182 ( .B1(u4_srl_451_n167), .B2(u4_srl_451_n168), .C1(
        u4_srl_451_n169), .C2(u4_srl_451_n170), .A(u4_srl_451_n171), .ZN(
        u4_srl_451_n166) );
  AOI21_X1 u4_srl_451_U181 ( .B1(u4_srl_451_n165), .B2(u4_srl_451_n166), .A(
        u4_shift_right[8]), .ZN(u4_N5909) );
  INV_X4 u4_srl_451_U180 ( .A(fract_denorm[102]), .ZN(u4_srl_451_n164) );
  INV_X4 u4_srl_451_U179 ( .A(fract_denorm[101]), .ZN(u4_srl_451_n163) );
  INV_X4 u4_srl_451_U178 ( .A(fract_denorm[100]), .ZN(u4_srl_451_n162) );
  INV_X4 u4_srl_451_U177 ( .A(fract_denorm[99]), .ZN(u4_srl_451_n161) );
  INV_X4 u4_srl_451_U176 ( .A(fract_denorm[98]), .ZN(u4_srl_451_n160) );
  INV_X4 u4_srl_451_U175 ( .A(fract_denorm[97]), .ZN(u4_srl_451_n159) );
  INV_X4 u4_srl_451_U174 ( .A(fract_denorm[96]), .ZN(u4_srl_451_n158) );
  INV_X4 u4_srl_451_U173 ( .A(fract_denorm[95]), .ZN(u4_srl_451_n157) );
  INV_X4 u4_srl_451_U172 ( .A(fract_denorm[94]), .ZN(u4_srl_451_n156) );
  INV_X4 u4_srl_451_U171 ( .A(fract_denorm[93]), .ZN(u4_srl_451_n155) );
  INV_X4 u4_srl_451_U170 ( .A(fract_denorm[92]), .ZN(u4_srl_451_n154) );
  INV_X4 u4_srl_451_U169 ( .A(fract_denorm[91]), .ZN(u4_srl_451_n153) );
  INV_X4 u4_srl_451_U168 ( .A(fract_denorm[90]), .ZN(u4_srl_451_n152) );
  INV_X4 u4_srl_451_U167 ( .A(fract_denorm[89]), .ZN(u4_srl_451_n151) );
  INV_X4 u4_srl_451_U166 ( .A(fract_denorm[88]), .ZN(u4_srl_451_n150) );
  INV_X4 u4_srl_451_U165 ( .A(fract_denorm[87]), .ZN(u4_srl_451_n149) );
  INV_X4 u4_srl_451_U164 ( .A(fract_denorm[86]), .ZN(u4_srl_451_n148) );
  INV_X4 u4_srl_451_U163 ( .A(fract_denorm[85]), .ZN(u4_srl_451_n147) );
  INV_X4 u4_srl_451_U162 ( .A(fract_denorm[84]), .ZN(u4_srl_451_n146) );
  INV_X4 u4_srl_451_U161 ( .A(fract_denorm[83]), .ZN(u4_srl_451_n145) );
  INV_X4 u4_srl_451_U160 ( .A(fract_denorm[82]), .ZN(u4_srl_451_n144) );
  INV_X4 u4_srl_451_U159 ( .A(fract_denorm[81]), .ZN(u4_srl_451_n143) );
  INV_X4 u4_srl_451_U158 ( .A(fract_denorm[80]), .ZN(u4_srl_451_n142) );
  INV_X4 u4_srl_451_U157 ( .A(fract_denorm[79]), .ZN(u4_srl_451_n141) );
  INV_X4 u4_srl_451_U156 ( .A(fract_denorm[78]), .ZN(u4_srl_451_n140) );
  INV_X4 u4_srl_451_U155 ( .A(fract_denorm[77]), .ZN(u4_srl_451_n139) );
  INV_X4 u4_srl_451_U154 ( .A(fract_denorm[76]), .ZN(u4_srl_451_n138) );
  INV_X4 u4_srl_451_U153 ( .A(fract_denorm[75]), .ZN(u4_srl_451_n137) );
  INV_X4 u4_srl_451_U152 ( .A(fract_denorm[74]), .ZN(u4_srl_451_n136) );
  INV_X4 u4_srl_451_U151 ( .A(fract_denorm[73]), .ZN(u4_srl_451_n135) );
  INV_X4 u4_srl_451_U150 ( .A(fract_denorm[72]), .ZN(u4_srl_451_n134) );
  INV_X4 u4_srl_451_U149 ( .A(fract_denorm[71]), .ZN(u4_srl_451_n133) );
  INV_X4 u4_srl_451_U148 ( .A(fract_denorm[70]), .ZN(u4_srl_451_n132) );
  INV_X4 u4_srl_451_U147 ( .A(fract_denorm[69]), .ZN(u4_srl_451_n131) );
  INV_X4 u4_srl_451_U146 ( .A(fract_denorm[68]), .ZN(u4_srl_451_n130) );
  INV_X4 u4_srl_451_U145 ( .A(fract_denorm[67]), .ZN(u4_srl_451_n129) );
  INV_X4 u4_srl_451_U144 ( .A(fract_denorm[66]), .ZN(u4_srl_451_n128) );
  INV_X4 u4_srl_451_U143 ( .A(fract_denorm[65]), .ZN(u4_srl_451_n127) );
  INV_X4 u4_srl_451_U142 ( .A(fract_denorm[64]), .ZN(u4_srl_451_n126) );
  INV_X4 u4_srl_451_U141 ( .A(fract_denorm[63]), .ZN(u4_srl_451_n125) );
  INV_X4 u4_srl_451_U140 ( .A(fract_denorm[62]), .ZN(u4_srl_451_n124) );
  INV_X4 u4_srl_451_U139 ( .A(fract_denorm[61]), .ZN(u4_srl_451_n123) );
  INV_X4 u4_srl_451_U138 ( .A(fract_denorm[60]), .ZN(u4_srl_451_n122) );
  INV_X4 u4_srl_451_U137 ( .A(fract_denorm[59]), .ZN(u4_srl_451_n121) );
  INV_X4 u4_srl_451_U136 ( .A(fract_denorm[58]), .ZN(u4_srl_451_n120) );
  INV_X4 u4_srl_451_U135 ( .A(fract_denorm[57]), .ZN(u4_srl_451_n119) );
  INV_X4 u4_srl_451_U134 ( .A(fract_denorm[56]), .ZN(u4_srl_451_n118) );
  INV_X4 u4_srl_451_U133 ( .A(fract_denorm[55]), .ZN(u4_srl_451_n117) );
  INV_X4 u4_srl_451_U132 ( .A(fract_denorm[54]), .ZN(u4_srl_451_n116) );
  INV_X4 u4_srl_451_U131 ( .A(fract_denorm[53]), .ZN(u4_srl_451_n115) );
  INV_X4 u4_srl_451_U130 ( .A(fract_denorm[52]), .ZN(u4_srl_451_n114) );
  INV_X4 u4_srl_451_U129 ( .A(fract_denorm[51]), .ZN(u4_srl_451_n113) );
  INV_X4 u4_srl_451_U128 ( .A(fract_denorm[50]), .ZN(u4_srl_451_n112) );
  INV_X4 u4_srl_451_U127 ( .A(fract_denorm[49]), .ZN(u4_srl_451_n111) );
  INV_X4 u4_srl_451_U126 ( .A(fract_denorm[48]), .ZN(u4_srl_451_n110) );
  INV_X4 u4_srl_451_U125 ( .A(fract_denorm[47]), .ZN(u4_srl_451_n109) );
  INV_X4 u4_srl_451_U124 ( .A(fract_denorm[46]), .ZN(u4_srl_451_n108) );
  INV_X4 u4_srl_451_U123 ( .A(fract_denorm[45]), .ZN(u4_srl_451_n107) );
  INV_X4 u4_srl_451_U122 ( .A(fract_denorm[44]), .ZN(u4_srl_451_n106) );
  INV_X4 u4_srl_451_U121 ( .A(fract_denorm[43]), .ZN(u4_srl_451_n105) );
  INV_X4 u4_srl_451_U120 ( .A(fract_denorm[42]), .ZN(u4_srl_451_n104) );
  INV_X4 u4_srl_451_U119 ( .A(fract_denorm[41]), .ZN(u4_srl_451_n103) );
  INV_X4 u4_srl_451_U118 ( .A(fract_denorm[40]), .ZN(u4_srl_451_n102) );
  INV_X4 u4_srl_451_U117 ( .A(fract_denorm[39]), .ZN(u4_srl_451_n101) );
  INV_X4 u4_srl_451_U116 ( .A(fract_denorm[38]), .ZN(u4_srl_451_n100) );
  INV_X4 u4_srl_451_U115 ( .A(fract_denorm[37]), .ZN(u4_srl_451_n99) );
  INV_X4 u4_srl_451_U114 ( .A(fract_denorm[36]), .ZN(u4_srl_451_n98) );
  INV_X4 u4_srl_451_U113 ( .A(fract_denorm[35]), .ZN(u4_srl_451_n97) );
  INV_X4 u4_srl_451_U112 ( .A(fract_denorm[34]), .ZN(u4_srl_451_n96) );
  INV_X4 u4_srl_451_U111 ( .A(fract_denorm[33]), .ZN(u4_srl_451_n95) );
  INV_X4 u4_srl_451_U110 ( .A(fract_denorm[32]), .ZN(u4_srl_451_n94) );
  INV_X4 u4_srl_451_U109 ( .A(fract_denorm[31]), .ZN(u4_srl_451_n93) );
  INV_X4 u4_srl_451_U108 ( .A(fract_denorm[30]), .ZN(u4_srl_451_n92) );
  INV_X4 u4_srl_451_U107 ( .A(fract_denorm[29]), .ZN(u4_srl_451_n91) );
  INV_X4 u4_srl_451_U106 ( .A(fract_denorm[28]), .ZN(u4_srl_451_n90) );
  INV_X4 u4_srl_451_U105 ( .A(fract_denorm[27]), .ZN(u4_srl_451_n89) );
  INV_X4 u4_srl_451_U104 ( .A(fract_denorm[26]), .ZN(u4_srl_451_n88) );
  INV_X4 u4_srl_451_U103 ( .A(fract_denorm[25]), .ZN(u4_srl_451_n87) );
  INV_X4 u4_srl_451_U102 ( .A(fract_denorm[24]), .ZN(u4_srl_451_n86) );
  INV_X4 u4_srl_451_U101 ( .A(fract_denorm[23]), .ZN(u4_srl_451_n85) );
  INV_X4 u4_srl_451_U100 ( .A(fract_denorm[22]), .ZN(u4_srl_451_n84) );
  INV_X4 u4_srl_451_U99 ( .A(fract_denorm[21]), .ZN(u4_srl_451_n83) );
  INV_X4 u4_srl_451_U98 ( .A(fract_denorm[19]), .ZN(u4_srl_451_n82) );
  INV_X4 u4_srl_451_U97 ( .A(fract_denorm[18]), .ZN(u4_srl_451_n81) );
  INV_X4 u4_srl_451_U96 ( .A(fract_denorm[17]), .ZN(u4_srl_451_n80) );
  INV_X4 u4_srl_451_U95 ( .A(fract_denorm[16]), .ZN(u4_srl_451_n79) );
  INV_X4 u4_srl_451_U94 ( .A(fract_denorm[15]), .ZN(u4_srl_451_n78) );
  INV_X4 u4_srl_451_U93 ( .A(fract_denorm[14]), .ZN(u4_srl_451_n77) );
  INV_X4 u4_srl_451_U92 ( .A(fract_denorm[13]), .ZN(u4_srl_451_n76) );
  INV_X4 u4_srl_451_U91 ( .A(fract_denorm[12]), .ZN(u4_srl_451_n75) );
  INV_X4 u4_srl_451_U90 ( .A(fract_denorm[11]), .ZN(u4_srl_451_n74) );
  INV_X4 u4_srl_451_U89 ( .A(fract_denorm[10]), .ZN(u4_srl_451_n73) );
  INV_X4 u4_srl_451_U88 ( .A(fract_denorm[9]), .ZN(u4_srl_451_n72) );
  INV_X4 u4_srl_451_U87 ( .A(fract_denorm[8]), .ZN(u4_srl_451_n71) );
  INV_X4 u4_srl_451_U86 ( .A(fract_denorm[7]), .ZN(u4_srl_451_n70) );
  INV_X4 u4_srl_451_U85 ( .A(fract_denorm[6]), .ZN(u4_srl_451_n69) );
  INV_X4 u4_srl_451_U84 ( .A(fract_denorm[5]), .ZN(u4_srl_451_n68) );
  INV_X4 u4_srl_451_U83 ( .A(fract_denorm[4]), .ZN(u4_srl_451_n67) );
  INV_X4 u4_srl_451_U82 ( .A(fract_denorm[3]), .ZN(u4_srl_451_n66) );
  INV_X4 u4_srl_451_U81 ( .A(fract_denorm[2]), .ZN(u4_srl_451_n65) );
  INV_X4 u4_srl_451_U80 ( .A(u4_srl_451_n381), .ZN(u4_srl_451_n388) );
  INV_X4 u4_srl_451_U79 ( .A(u4_srl_451_n863), .ZN(u4_srl_451_n179) );
  AND2_X4 u4_srl_451_U78 ( .A1(u4_srl_451_n17), .A2(u4_srl_451_n798), .ZN(
        u4_srl_451_n167) );
  AND2_X4 u4_srl_451_U77 ( .A1(u4_srl_451_n61), .A2(u4_srl_451_n798), .ZN(
        u4_srl_451_n169) );
  INV_X4 u4_srl_451_U76 ( .A(u4_srl_451_n7), .ZN(u4_srl_451_n10) );
  INV_X4 u4_srl_451_U75 ( .A(u4_srl_451_n5), .ZN(u4_srl_451_n64) );
  INV_X4 u4_srl_451_U74 ( .A(u4_srl_451_n3), .ZN(u4_srl_451_n15) );
  INV_X4 u4_srl_451_U73 ( .A(u4_srl_451_n12), .ZN(u4_srl_451_n13) );
  INV_X4 u4_srl_451_U72 ( .A(u4_srl_451_n25), .ZN(u4_srl_451_n21) );
  INV_X4 u4_srl_451_U71 ( .A(u4_srl_451_n46), .ZN(u4_srl_451_n42) );
  INV_X4 u4_srl_451_U70 ( .A(u4_srl_451_n46), .ZN(u4_srl_451_n41) );
  INV_X4 u4_srl_451_U69 ( .A(u4_srl_451_n45), .ZN(u4_srl_451_n44) );
  INV_X4 u4_srl_451_U68 ( .A(u4_srl_451_n6), .ZN(u4_srl_451_n29) );
  INV_X4 u4_srl_451_U67 ( .A(u4_srl_451_n6), .ZN(u4_srl_451_n30) );
  INV_X4 u4_srl_451_U66 ( .A(u4_srl_451_n6), .ZN(u4_srl_451_n26) );
  INV_X4 u4_srl_451_U65 ( .A(u4_srl_451_n20), .ZN(u4_srl_451_n17) );
  INV_X4 u4_srl_451_U64 ( .A(u4_srl_451_n317), .ZN(u4_srl_451_n12) );
  INV_X4 u4_srl_451_U63 ( .A(u4_srl_451_n3), .ZN(u4_srl_451_n14) );
  INV_X4 u4_srl_451_U62 ( .A(u4_srl_451_n1), .ZN(u4_srl_451_n47) );
  INV_X4 u4_srl_451_U61 ( .A(u4_srl_451_n63), .ZN(u4_srl_451_n61) );
  INV_X4 u4_srl_451_U60 ( .A(u4_srl_451_n25), .ZN(u4_srl_451_n22) );
  INV_X4 u4_srl_451_U59 ( .A(u4_srl_451_n25), .ZN(u4_srl_451_n23) );
  INV_X4 u4_srl_451_U58 ( .A(u4_srl_451_n25), .ZN(u4_srl_451_n24) );
  INV_X4 u4_srl_451_U57 ( .A(u4_srl_451_n46), .ZN(u4_srl_451_n40) );
  INV_X4 u4_srl_451_U56 ( .A(u4_srl_451_n6), .ZN(u4_srl_451_n27) );
  INV_X4 u4_srl_451_U55 ( .A(u4_srl_451_n6), .ZN(u4_srl_451_n28) );
  INV_X4 u4_srl_451_U54 ( .A(u4_srl_451_n20), .ZN(u4_srl_451_n18) );
  INV_X4 u4_srl_451_U53 ( .A(u4_srl_451_n19), .ZN(u4_srl_451_n16) );
  INV_X4 u4_srl_451_U52 ( .A(u4_srl_451_n398), .ZN(u4_srl_451_n19) );
  INV_X4 u4_srl_451_U51 ( .A(u4_srl_451_n399), .ZN(u4_srl_451_n25) );
  INV_X4 u4_srl_451_U50 ( .A(u4_srl_451_n7), .ZN(u4_srl_451_n11) );
  INV_X4 u4_srl_451_U49 ( .A(u4_srl_451_n400), .ZN(u4_srl_451_n45) );
  INV_X4 u4_srl_451_U48 ( .A(u4_srl_451_n400), .ZN(u4_srl_451_n46) );
  INV_X4 u4_srl_451_U47 ( .A(u4_srl_451_n1), .ZN(u4_srl_451_n50) );
  INV_X4 u4_srl_451_U46 ( .A(u4_srl_451_n63), .ZN(u4_srl_451_n62) );
  INV_X4 u4_srl_451_U45 ( .A(u4_srl_451_n5), .ZN(u4_srl_451_n63) );
  INV_X4 u4_srl_451_U44 ( .A(u4_srl_451_n8), .ZN(u4_srl_451_n9) );
  INV_X4 u4_srl_451_U43 ( .A(u4_srl_451_n1), .ZN(u4_srl_451_n49) );
  INV_X4 u4_srl_451_U42 ( .A(u4_srl_451_n53), .ZN(u4_srl_451_n56) );
  INV_X4 u4_srl_451_U41 ( .A(u4_srl_451_n59), .ZN(u4_srl_451_n58) );
  INV_X4 u4_srl_451_U40 ( .A(u4_srl_451_n2), .ZN(u4_srl_451_n59) );
  INV_X4 u4_srl_451_U39 ( .A(u4_srl_451_n398), .ZN(u4_srl_451_n20) );
  INV_X4 u4_srl_451_U38 ( .A(u4_srl_451_n186), .ZN(u4_srl_451_n8) );
  INV_X4 u4_srl_451_U37 ( .A(u4_srl_451_n2), .ZN(u4_srl_451_n53) );
  INV_X4 u4_srl_451_U36 ( .A(u4_srl_451_n38), .ZN(u4_srl_451_n31) );
  INV_X4 u4_srl_451_U35 ( .A(u4_srl_451_n38), .ZN(u4_srl_451_n32) );
  INV_X4 u4_srl_451_U34 ( .A(u4_srl_451_n37), .ZN(u4_srl_451_n34) );
  INV_X4 u4_srl_451_U33 ( .A(u4_srl_451_n46), .ZN(u4_srl_451_n43) );
  INV_X4 u4_srl_451_U32 ( .A(u4_srl_451_n63), .ZN(u4_srl_451_n60) );
  AND2_X4 u4_srl_451_U31 ( .A1(u4_srl_451_n391), .A2(u4_shift_right[4]), .ZN(
        u4_srl_451_n7) );
  INV_X4 u4_srl_451_U30 ( .A(u4_srl_451_n1), .ZN(u4_srl_451_n48) );
  OR2_X4 u4_srl_451_U29 ( .A1(u4_shift_right[2]), .A2(u4_srl_451_n837), .ZN(
        u4_srl_451_n6) );
  NOR2_X2 u4_srl_451_U28 ( .A1(u4_srl_451_n732), .A2(u4_shift_right[2]), .ZN(
        u4_srl_451_n5) );
  AND2_X4 u4_srl_451_U27 ( .A1(u4_srl_451_n882), .A2(u4_shift_right[0]), .ZN(
        u4_srl_451_n4) );
  OR2_X4 u4_srl_451_U26 ( .A1(u4_srl_451_n304), .A2(u4_shift_right[4]), .ZN(
        u4_srl_451_n3) );
  OR2_X4 u4_srl_451_U25 ( .A1(u4_shift_right[0]), .A2(u4_srl_451_n882), .ZN(
        u4_srl_451_n2) );
  OR2_X4 u4_srl_451_U24 ( .A1(u4_srl_451_n883), .A2(u4_srl_451_n882), .ZN(
        u4_srl_451_n1) );
  NOR2_X2 u4_srl_451_U23 ( .A1(u4_srl_451_n179), .A2(u4_shift_right[8]), .ZN(
        u4_srl_451_n215) );
  NOR2_X2 u4_srl_451_U22 ( .A1(u4_srl_451_n247), .A2(u4_srl_451_n179), .ZN(
        u4_srl_451_n176) );
  NAND2_X2 u4_srl_451_U21 ( .A1(u4_srl_451_n30), .A2(u4_srl_451_n798), .ZN(
        u4_srl_451_n173) );
  NAND2_X2 u4_srl_451_U20 ( .A1(u4_srl_451_n798), .A2(u4_srl_451_n24), .ZN(
        u4_srl_451_n175) );
  NOR2_X2 u4_srl_451_U19 ( .A1(u4_srl_451_n388), .A2(u4_srl_451_n243), .ZN(
        u4_srl_451_n413) );
  INV_X4 u4_srl_451_U18 ( .A(u4_shift_right[4]), .ZN(u4_srl_451_n397) );
  INV_X4 u4_srl_451_U17 ( .A(u4_srl_451_n56), .ZN(u4_srl_451_n55) );
  INV_X4 u4_srl_451_U16 ( .A(u4_srl_451_n39), .ZN(u4_srl_451_n38) );
  INV_X4 u4_srl_451_U15 ( .A(u4_srl_451_n58), .ZN(u4_srl_451_n54) );
  NAND2_X2 u4_srl_451_U14 ( .A1(u4_srl_451_n271), .A2(u4_srl_451_n397), .ZN(
        u4_srl_451_n243) );
  NAND2_X2 u4_srl_451_U13 ( .A1(u4_srl_451_n271), .A2(u4_shift_right[4]), .ZN(
        u4_srl_451_n247) );
  NAND2_X2 u4_srl_451_U12 ( .A1(u4_srl_451_n805), .A2(u4_shift_right[4]), .ZN(
        u4_srl_451_n182) );
  NAND2_X2 u4_srl_451_U11 ( .A1(u4_srl_451_n805), .A2(u4_srl_451_n397), .ZN(
        u4_srl_451_n184) );
  INV_X4 u4_srl_451_U10 ( .A(u4_srl_451_n57), .ZN(u4_srl_451_n52) );
  INV_X4 u4_srl_451_U9 ( .A(u4_srl_451_n37), .ZN(u4_srl_451_n33) );
  INV_X4 u4_srl_451_U8 ( .A(u4_srl_451_n57), .ZN(u4_srl_451_n51) );
  INV_X4 u4_srl_451_U7 ( .A(u4_srl_451_n37), .ZN(u4_srl_451_n35) );
  INV_X4 u4_srl_451_U6 ( .A(u4_srl_451_n4), .ZN(u4_srl_451_n39) );
  INV_X4 u4_srl_451_U5 ( .A(u4_srl_451_n39), .ZN(u4_srl_451_n37) );
  INV_X4 u4_srl_451_U4 ( .A(u4_srl_451_n59), .ZN(u4_srl_451_n57) );
  INV_X4 u4_srl_451_U3 ( .A(u4_srl_451_n37), .ZN(u4_srl_451_n36) );
  OR3_X1 u4_sll_480_U89 ( .A1(u4_f2i_shft_8_), .A2(u4_f2i_shft_9_), .A3(
        u4_f2i_shft_7_), .ZN(u4_sll_480_n58) );
  NAND2_X1 u4_sll_480_U88 ( .A1(u4_sll_480_n58), .A2(u4_sll_480_n45), .ZN(
        u4_sll_480_n47) );
  NAND3_X1 u4_sll_480_U87 ( .A1(u4_f2i_shft_8_), .A2(u4_f2i_shft_7_), .A3(
        u4_f2i_shft_9_), .ZN(u4_sll_480_n57) );
  NAND2_X1 u4_sll_480_U86 ( .A1(u4_f2i_shft_10_), .A2(u4_sll_480_n57), .ZN(
        u4_sll_480_n46) );
  NAND2_X1 u4_sll_480_U85 ( .A1(n4400), .A2(u4_sll_480_n46), .ZN(
        u4_sll_480_n56) );
  NAND2_X1 u4_sll_480_U84 ( .A1(u4_sll_480_n47), .A2(u4_sll_480_n56), .ZN(
        u4_sll_480_temp_int_SH_0_) );
  AND2_X1 u4_sll_480_U83 ( .A1(fract_denorm[0]), .A2(u4_sll_480_n12), .ZN(
        u4_sll_480_ML_int_1__0_) );
  AND2_X1 u4_sll_480_U82 ( .A1(n4873), .A2(u4_sll_480_n6), .ZN(
        u4_sll_480_MR_int_1__113_) );
  NAND2_X1 u4_sll_480_U81 ( .A1(u4_f2i_shft_1_), .A2(u4_sll_480_n46), .ZN(
        u4_sll_480_n55) );
  NAND2_X1 u4_sll_480_U80 ( .A1(u4_sll_480_ML_int_1__0_), .A2(u4_sll_480_n1), 
        .ZN(u4_sll_480_n52) );
  NAND2_X1 u4_sll_480_U79 ( .A1(u4_sll_480_ML_int_1__1_), .A2(u4_sll_480_n1), 
        .ZN(u4_sll_480_n51) );
  NAND2_X1 u4_sll_480_U78 ( .A1(u4_f2i_shft_2_), .A2(u4_sll_480_n46), .ZN(
        u4_sll_480_n54) );
  NAND2_X1 u4_sll_480_U77 ( .A1(u4_sll_480_ML_int_2__3_), .A2(u4_sll_480_n2), 
        .ZN(u4_sll_480_n49) );
  NAND2_X1 u4_sll_480_U76 ( .A1(u4_f2i_shft_3_), .A2(u4_sll_480_n46), .ZN(
        u4_sll_480_n53) );
  NAND2_X1 u4_sll_480_U75 ( .A1(u4_sll_480_n47), .A2(u4_sll_480_n53), .ZN(
        u4_sll_480_temp_int_SH_3_) );
  NAND2_X1 u4_sll_480_U74 ( .A1(u4_sll_480_n2), .A2(u4_sll_480_n34), .ZN(
        u4_sll_480_n50) );
  NOR2_X1 u4_sll_480_U73 ( .A1(u4_sll_480_n50), .A2(u4_sll_480_n52), .ZN(
        u4_sll_480_ML_int_4__0_) );
  NOR2_X1 u4_sll_480_U72 ( .A1(u4_sll_480_n50), .A2(u4_sll_480_n51), .ZN(
        u4_sll_480_ML_int_4__1_) );
  NOR2_X1 u4_sll_480_U71 ( .A1(u4_sll_480_n39), .A2(u4_sll_480_n50), .ZN(
        u4_sll_480_ML_int_4__2_) );
  NOR2_X1 u4_sll_480_U70 ( .A1(u4_sll_480_n30), .A2(u4_sll_480_n49), .ZN(
        u4_sll_480_ML_int_4__3_) );
  AND2_X1 u4_sll_480_U69 ( .A1(u4_sll_480_ML_int_3__4_), .A2(u4_sll_480_n34), 
        .ZN(u4_sll_480_ML_int_4__4_) );
  AND2_X1 u4_sll_480_U68 ( .A1(u4_sll_480_ML_int_3__5_), .A2(u4_sll_480_n34), 
        .ZN(u4_sll_480_ML_int_4__5_) );
  NAND2_X1 u4_sll_480_U67 ( .A1(u4_f2i_shft_4_), .A2(u4_sll_480_n46), .ZN(
        u4_sll_480_n48) );
  NAND2_X1 u4_sll_480_U66 ( .A1(u4_sll_480_n47), .A2(u4_sll_480_n48), .ZN(
        u4_sll_480_temp_int_SH_4_) );
  AND2_X1 u4_sll_480_U65 ( .A1(u4_sll_480_ML_int_4__11_), .A2(u4_sll_480_n35), 
        .ZN(u4_sll_480_ML_int_5__11_) );
  AND2_X1 u4_sll_480_U64 ( .A1(u4_sll_480_ML_int_4__12_), .A2(u4_sll_480_n35), 
        .ZN(u4_sll_480_ML_int_5__12_) );
  AND2_X1 u4_sll_480_U63 ( .A1(u4_sll_480_ML_int_4__13_), .A2(u4_sll_480_n35), 
        .ZN(u4_sll_480_ML_int_5__13_) );
  AND2_X1 u4_sll_480_U62 ( .A1(u4_sll_480_ML_int_4__14_), .A2(u4_sll_480_n35), 
        .ZN(u4_sll_480_ML_int_5__14_) );
  AND2_X1 u4_sll_480_U61 ( .A1(u4_sll_480_ML_int_4__15_), .A2(u4_sll_480_n35), 
        .ZN(u4_sll_480_ML_int_5__15_) );
  AND2_X1 u4_sll_480_U60 ( .A1(u4_sll_480_ML_int_7__107_), .A2(u4_sll_480_n45), 
        .ZN(u4_exp_f2i_1[107]) );
  AND2_X1 u4_sll_480_U59 ( .A1(u4_sll_480_ML_int_7__108_), .A2(u4_sll_480_n45), 
        .ZN(u4_exp_f2i_1[108]) );
  AND2_X1 u4_sll_480_U58 ( .A1(u4_sll_480_ML_int_7__109_), .A2(u4_sll_480_n45), 
        .ZN(u4_exp_f2i_1[109]) );
  AND2_X1 u4_sll_480_U57 ( .A1(u4_sll_480_ML_int_7__110_), .A2(u4_sll_480_n45), 
        .ZN(u4_exp_f2i_1[110]) );
  AND2_X1 u4_sll_480_U56 ( .A1(u4_sll_480_ML_int_7__111_), .A2(u4_sll_480_n45), 
        .ZN(u4_exp_f2i_1[111]) );
  AND2_X1 u4_sll_480_U55 ( .A1(u4_sll_480_ML_int_7__112_), .A2(u4_sll_480_n45), 
        .ZN(u4_exp_f2i_1[112]) );
  AND2_X1 u4_sll_480_U54 ( .A1(u4_sll_480_ML_int_7__113_), .A2(u4_sll_480_n45), 
        .ZN(u4_exp_f2i_1[113]) );
  AND2_X1 u4_sll_480_U53 ( .A1(u4_sll_480_ML_int_7__114_), .A2(u4_sll_480_n45), 
        .ZN(u4_exp_f2i_1[114]) );
  AND2_X1 u4_sll_480_U52 ( .A1(u4_sll_480_ML_int_7__115_), .A2(u4_sll_480_n45), 
        .ZN(u4_exp_f2i_1[115]) );
  AND2_X1 u4_sll_480_U51 ( .A1(u4_sll_480_ML_int_7__116_), .A2(u4_sll_480_n45), 
        .ZN(u4_exp_f2i_1[116]) );
  AND2_X1 u4_sll_480_U50 ( .A1(u4_sll_480_ML_int_7__117_), .A2(u4_sll_480_n45), 
        .ZN(u4_exp_f2i_1[117]) );
  OAI21_X1 u4_sll_480_U49 ( .B1(u4_f2i_shft_5_), .B2(u4_sll_480_n44), .A(
        u4_sll_480_n46), .ZN(u4_sll_480_SHMAG[5]) );
  OAI21_X1 u4_sll_480_U48 ( .B1(u4_f2i_shft_6_), .B2(u4_sll_480_n44), .A(
        u4_sll_480_n46), .ZN(u4_sll_480_SHMAG[6]) );
  INV_X4 u4_sll_480_U47 ( .A(u4_f2i_shft_10_), .ZN(u4_sll_480_n45) );
  INV_X4 u4_sll_480_U46 ( .A(u4_sll_480_n47), .ZN(u4_sll_480_n44) );
  INV_X4 u4_sll_480_U45 ( .A(u4_sll_480_SHMAG[6]), .ZN(u4_sll_480_n43) );
  INV_X4 u4_sll_480_U44 ( .A(u4_sll_480_SHMAG[5]), .ZN(u4_sll_480_n42) );
  INV_X4 u4_sll_480_U43 ( .A(u4_sll_480_n49), .ZN(u4_sll_480_n41) );
  INV_X4 u4_sll_480_U42 ( .A(u4_sll_480_n51), .ZN(u4_sll_480_n40) );
  INV_X4 u4_sll_480_U41 ( .A(u4_sll_480_ML_int_2__2_), .ZN(u4_sll_480_n39) );
  INV_X4 u4_sll_480_U40 ( .A(u4_sll_480_n52), .ZN(u4_sll_480_n38) );
  AND2_X4 u4_sll_480_U39 ( .A1(u4_sll_480_n29), .A2(u4_sll_480_ML_int_2__113_), 
        .ZN(u4_sll_480_n5) );
  AND2_X4 u4_sll_480_U38 ( .A1(u4_sll_480_n20), .A2(u4_sll_480_MR_int_1__113_), 
        .ZN(u4_sll_480_n4) );
  INV_X4 u4_sll_480_U37 ( .A(u4_sll_480_n1), .ZN(u4_sll_480_n22) );
  INV_X4 u4_sll_480_U36 ( .A(u4_sll_480_n35), .ZN(u4_sll_480_n37) );
  INV_X4 u4_sll_480_U35 ( .A(u4_sll_480_n35), .ZN(u4_sll_480_n36) );
  INV_X4 u4_sll_480_U34 ( .A(u4_sll_480_n34), .ZN(u4_sll_480_n33) );
  INV_X4 u4_sll_480_U33 ( .A(u4_sll_480_n2), .ZN(u4_sll_480_n29) );
  INV_X4 u4_sll_480_U32 ( .A(u4_sll_480_n2), .ZN(u4_sll_480_n28) );
  INV_X4 u4_sll_480_U31 ( .A(u4_sll_480_n2), .ZN(u4_sll_480_n23) );
  INV_X4 u4_sll_480_U30 ( .A(u4_sll_480_temp_int_SH_4_), .ZN(u4_sll_480_n35)
         );
  INV_X4 u4_sll_480_U29 ( .A(u4_sll_480_n1), .ZN(u4_sll_480_n18) );
  INV_X4 u4_sll_480_U28 ( .A(u4_sll_480_n1), .ZN(u4_sll_480_n20) );
  INV_X4 u4_sll_480_U27 ( .A(u4_sll_480_n1), .ZN(u4_sll_480_n16) );
  AND2_X4 u4_sll_480_U26 ( .A1(u4_sll_480_n22), .A2(u4_sll_480_ML_int_1__113_), 
        .ZN(u4_sll_480_n3) );
  INV_X4 u4_sll_480_U25 ( .A(u4_sll_480_n34), .ZN(u4_sll_480_n30) );
  INV_X4 u4_sll_480_U24 ( .A(u4_sll_480_temp_int_SH_3_), .ZN(u4_sll_480_n34)
         );
  INV_X4 u4_sll_480_U23 ( .A(u4_sll_480_n34), .ZN(u4_sll_480_n32) );
  INV_X4 u4_sll_480_U22 ( .A(u4_sll_480_n1), .ZN(u4_sll_480_n17) );
  INV_X4 u4_sll_480_U21 ( .A(u4_sll_480_n1), .ZN(u4_sll_480_n19) );
  INV_X4 u4_sll_480_U20 ( .A(u4_sll_480_n12), .ZN(u4_sll_480_n6) );
  INV_X4 u4_sll_480_U19 ( .A(u4_sll_480_temp_int_SH_0_), .ZN(u4_sll_480_n15)
         );
  INV_X4 u4_sll_480_U18 ( .A(u4_sll_480_n12), .ZN(u4_sll_480_n7) );
  INV_X4 u4_sll_480_U17 ( .A(u4_sll_480_n34), .ZN(u4_sll_480_n31) );
  INV_X4 u4_sll_480_U16 ( .A(u4_sll_480_n11), .ZN(u4_sll_480_n9) );
  INV_X4 u4_sll_480_U15 ( .A(u4_sll_480_n15), .ZN(u4_sll_480_n13) );
  INV_X4 u4_sll_480_U14 ( .A(u4_sll_480_n2), .ZN(u4_sll_480_n26) );
  INV_X4 u4_sll_480_U13 ( .A(u4_sll_480_n2), .ZN(u4_sll_480_n27) );
  INV_X4 u4_sll_480_U12 ( .A(u4_sll_480_n11), .ZN(u4_sll_480_n8) );
  INV_X4 u4_sll_480_U11 ( .A(u4_sll_480_n11), .ZN(u4_sll_480_n10) );
  INV_X4 u4_sll_480_U10 ( .A(u4_sll_480_n14), .ZN(u4_sll_480_n11) );
  INV_X4 u4_sll_480_U9 ( .A(u4_sll_480_n15), .ZN(u4_sll_480_n14) );
  INV_X4 u4_sll_480_U8 ( .A(u4_sll_480_n2), .ZN(u4_sll_480_n25) );
  INV_X4 u4_sll_480_U7 ( .A(u4_sll_480_n13), .ZN(u4_sll_480_n12) );
  INV_X4 u4_sll_480_U6 ( .A(u4_sll_480_n2), .ZN(u4_sll_480_n24) );
  INV_X4 u4_sll_480_U5 ( .A(u4_sll_480_n1), .ZN(u4_sll_480_n21) );
  AND2_X4 u4_sll_480_U4 ( .A1(u4_sll_480_n47), .A2(u4_sll_480_n54), .ZN(
        u4_sll_480_n2) );
  AND2_X4 u4_sll_480_U3 ( .A1(u4_sll_480_n47), .A2(u4_sll_480_n55), .ZN(
        u4_sll_480_n1) );
  MUX2_X2 u4_sll_480_M1_0_1 ( .A(fract_denorm[1]), .B(fract_denorm[0]), .S(
        u4_sll_480_n6), .Z(u4_sll_480_ML_int_1__1_) );
  MUX2_X2 u4_sll_480_M1_0_2 ( .A(fract_denorm[2]), .B(fract_denorm[1]), .S(
        u4_sll_480_n6), .Z(u4_sll_480_ML_int_1__2_) );
  MUX2_X2 u4_sll_480_M1_0_3 ( .A(fract_denorm[3]), .B(fract_denorm[2]), .S(
        u4_sll_480_n6), .Z(u4_sll_480_ML_int_1__3_) );
  MUX2_X2 u4_sll_480_M1_0_4 ( .A(fract_denorm[4]), .B(fract_denorm[3]), .S(
        u4_sll_480_n10), .Z(u4_sll_480_ML_int_1__4_) );
  MUX2_X2 u4_sll_480_M1_0_5 ( .A(fract_denorm[5]), .B(fract_denorm[4]), .S(
        u4_sll_480_n10), .Z(u4_sll_480_ML_int_1__5_) );
  MUX2_X2 u4_sll_480_M1_0_6 ( .A(fract_denorm[6]), .B(fract_denorm[5]), .S(
        u4_sll_480_n10), .Z(u4_sll_480_ML_int_1__6_) );
  MUX2_X2 u4_sll_480_M1_0_7 ( .A(fract_denorm[7]), .B(fract_denorm[6]), .S(
        u4_sll_480_n10), .Z(u4_sll_480_ML_int_1__7_) );
  MUX2_X2 u4_sll_480_M1_0_8 ( .A(fract_denorm[8]), .B(fract_denorm[7]), .S(
        u4_sll_480_n10), .Z(u4_sll_480_ML_int_1__8_) );
  MUX2_X2 u4_sll_480_M1_0_9 ( .A(fract_denorm[9]), .B(fract_denorm[8]), .S(
        u4_sll_480_n10), .Z(u4_sll_480_ML_int_1__9_) );
  MUX2_X2 u4_sll_480_M1_0_10 ( .A(fract_denorm[10]), .B(fract_denorm[9]), .S(
        u4_sll_480_n10), .Z(u4_sll_480_ML_int_1__10_) );
  MUX2_X2 u4_sll_480_M1_0_11 ( .A(fract_denorm[11]), .B(fract_denorm[10]), .S(
        u4_sll_480_n10), .Z(u4_sll_480_ML_int_1__11_) );
  MUX2_X2 u4_sll_480_M1_0_12 ( .A(fract_denorm[12]), .B(fract_denorm[11]), .S(
        u4_sll_480_n10), .Z(u4_sll_480_ML_int_1__12_) );
  MUX2_X2 u4_sll_480_M1_0_13 ( .A(fract_denorm[13]), .B(fract_denorm[12]), .S(
        u4_sll_480_n10), .Z(u4_sll_480_ML_int_1__13_) );
  MUX2_X2 u4_sll_480_M1_0_14 ( .A(fract_denorm[14]), .B(fract_denorm[13]), .S(
        u4_sll_480_n10), .Z(u4_sll_480_ML_int_1__14_) );
  MUX2_X2 u4_sll_480_M1_0_15 ( .A(fract_denorm[15]), .B(fract_denorm[14]), .S(
        u4_sll_480_n9), .Z(u4_sll_480_ML_int_1__15_) );
  MUX2_X2 u4_sll_480_M1_0_16 ( .A(fract_denorm[16]), .B(fract_denorm[15]), .S(
        u4_sll_480_n9), .Z(u4_sll_480_ML_int_1__16_) );
  MUX2_X2 u4_sll_480_M1_0_17 ( .A(fract_denorm[17]), .B(fract_denorm[16]), .S(
        u4_sll_480_n9), .Z(u4_sll_480_ML_int_1__17_) );
  MUX2_X2 u4_sll_480_M1_0_18 ( .A(fract_denorm[18]), .B(fract_denorm[17]), .S(
        u4_sll_480_n9), .Z(u4_sll_480_ML_int_1__18_) );
  MUX2_X2 u4_sll_480_M1_0_19 ( .A(fract_denorm[19]), .B(fract_denorm[18]), .S(
        u4_sll_480_n9), .Z(u4_sll_480_ML_int_1__19_) );
  MUX2_X2 u4_sll_480_M1_0_20 ( .A(fract_denorm[20]), .B(fract_denorm[19]), .S(
        u4_sll_480_n9), .Z(u4_sll_480_ML_int_1__20_) );
  MUX2_X2 u4_sll_480_M1_0_21 ( .A(fract_denorm[21]), .B(fract_denorm[20]), .S(
        u4_sll_480_n9), .Z(u4_sll_480_ML_int_1__21_) );
  MUX2_X2 u4_sll_480_M1_0_22 ( .A(fract_denorm[22]), .B(fract_denorm[21]), .S(
        u4_sll_480_n9), .Z(u4_sll_480_ML_int_1__22_) );
  MUX2_X2 u4_sll_480_M1_0_23 ( .A(fract_denorm[23]), .B(fract_denorm[22]), .S(
        u4_sll_480_n9), .Z(u4_sll_480_ML_int_1__23_) );
  MUX2_X2 u4_sll_480_M1_0_24 ( .A(fract_denorm[24]), .B(fract_denorm[23]), .S(
        u4_sll_480_n9), .Z(u4_sll_480_ML_int_1__24_) );
  MUX2_X2 u4_sll_480_M1_0_25 ( .A(fract_denorm[25]), .B(fract_denorm[24]), .S(
        u4_sll_480_n9), .Z(u4_sll_480_ML_int_1__25_) );
  MUX2_X2 u4_sll_480_M1_0_26 ( .A(fract_denorm[26]), .B(fract_denorm[25]), .S(
        u4_sll_480_n14), .Z(u4_sll_480_ML_int_1__26_) );
  MUX2_X2 u4_sll_480_M1_0_27 ( .A(fract_denorm[27]), .B(fract_denorm[26]), .S(
        u4_sll_480_n13), .Z(u4_sll_480_ML_int_1__27_) );
  MUX2_X2 u4_sll_480_M1_0_28 ( .A(fract_denorm[28]), .B(fract_denorm[27]), .S(
        u4_sll_480_n9), .Z(u4_sll_480_ML_int_1__28_) );
  MUX2_X2 u4_sll_480_M1_0_29 ( .A(fract_denorm[29]), .B(fract_denorm[28]), .S(
        u4_sll_480_n14), .Z(u4_sll_480_ML_int_1__29_) );
  MUX2_X2 u4_sll_480_M1_0_30 ( .A(fract_denorm[30]), .B(fract_denorm[29]), .S(
        u4_sll_480_n9), .Z(u4_sll_480_ML_int_1__30_) );
  MUX2_X2 u4_sll_480_M1_0_31 ( .A(fract_denorm[31]), .B(fract_denorm[30]), .S(
        u4_sll_480_temp_int_SH_0_), .Z(u4_sll_480_ML_int_1__31_) );
  MUX2_X2 u4_sll_480_M1_0_32 ( .A(fract_denorm[32]), .B(fract_denorm[31]), .S(
        u4_sll_480_n14), .Z(u4_sll_480_ML_int_1__32_) );
  MUX2_X2 u4_sll_480_M1_0_33 ( .A(fract_denorm[33]), .B(fract_denorm[32]), .S(
        u4_sll_480_temp_int_SH_0_), .Z(u4_sll_480_ML_int_1__33_) );
  MUX2_X2 u4_sll_480_M1_0_34 ( .A(fract_denorm[34]), .B(fract_denorm[33]), .S(
        u4_sll_480_n14), .Z(u4_sll_480_ML_int_1__34_) );
  MUX2_X2 u4_sll_480_M1_0_35 ( .A(fract_denorm[35]), .B(fract_denorm[34]), .S(
        u4_sll_480_temp_int_SH_0_), .Z(u4_sll_480_ML_int_1__35_) );
  MUX2_X2 u4_sll_480_M1_0_36 ( .A(fract_denorm[36]), .B(fract_denorm[35]), .S(
        u4_sll_480_n9), .Z(u4_sll_480_ML_int_1__36_) );
  MUX2_X2 u4_sll_480_M1_0_37 ( .A(fract_denorm[37]), .B(fract_denorm[36]), .S(
        u4_sll_480_n8), .Z(u4_sll_480_ML_int_1__37_) );
  MUX2_X2 u4_sll_480_M1_0_38 ( .A(fract_denorm[38]), .B(fract_denorm[37]), .S(
        u4_sll_480_n8), .Z(u4_sll_480_ML_int_1__38_) );
  MUX2_X2 u4_sll_480_M1_0_39 ( .A(fract_denorm[39]), .B(fract_denorm[38]), .S(
        u4_sll_480_n8), .Z(u4_sll_480_ML_int_1__39_) );
  MUX2_X2 u4_sll_480_M1_0_40 ( .A(fract_denorm[40]), .B(fract_denorm[39]), .S(
        u4_sll_480_n8), .Z(u4_sll_480_ML_int_1__40_) );
  MUX2_X2 u4_sll_480_M1_0_41 ( .A(fract_denorm[41]), .B(fract_denorm[40]), .S(
        u4_sll_480_n8), .Z(u4_sll_480_ML_int_1__41_) );
  MUX2_X2 u4_sll_480_M1_0_42 ( .A(fract_denorm[42]), .B(fract_denorm[41]), .S(
        u4_sll_480_n8), .Z(u4_sll_480_ML_int_1__42_) );
  MUX2_X2 u4_sll_480_M1_0_43 ( .A(fract_denorm[43]), .B(fract_denorm[42]), .S(
        u4_sll_480_n8), .Z(u4_sll_480_ML_int_1__43_) );
  MUX2_X2 u4_sll_480_M1_0_44 ( .A(fract_denorm[44]), .B(fract_denorm[43]), .S(
        u4_sll_480_n8), .Z(u4_sll_480_ML_int_1__44_) );
  MUX2_X2 u4_sll_480_M1_0_45 ( .A(fract_denorm[45]), .B(fract_denorm[44]), .S(
        u4_sll_480_n8), .Z(u4_sll_480_ML_int_1__45_) );
  MUX2_X2 u4_sll_480_M1_0_46 ( .A(fract_denorm[46]), .B(fract_denorm[45]), .S(
        u4_sll_480_n8), .Z(u4_sll_480_ML_int_1__46_) );
  MUX2_X2 u4_sll_480_M1_0_47 ( .A(fract_denorm[47]), .B(fract_denorm[46]), .S(
        u4_sll_480_n8), .Z(u4_sll_480_ML_int_1__47_) );
  MUX2_X2 u4_sll_480_M1_0_48 ( .A(fract_denorm[48]), .B(fract_denorm[47]), .S(
        u4_sll_480_n8), .Z(u4_sll_480_ML_int_1__48_) );
  MUX2_X2 u4_sll_480_M1_0_49 ( .A(fract_denorm[49]), .B(fract_denorm[48]), .S(
        u4_sll_480_n10), .Z(u4_sll_480_ML_int_1__49_) );
  MUX2_X2 u4_sll_480_M1_0_50 ( .A(fract_denorm[50]), .B(fract_denorm[49]), .S(
        u4_sll_480_n10), .Z(u4_sll_480_ML_int_1__50_) );
  MUX2_X2 u4_sll_480_M1_0_51 ( .A(fract_denorm[51]), .B(fract_denorm[50]), .S(
        u4_sll_480_n10), .Z(u4_sll_480_ML_int_1__51_) );
  MUX2_X2 u4_sll_480_M1_0_52 ( .A(fract_denorm[52]), .B(fract_denorm[51]), .S(
        u4_sll_480_n10), .Z(u4_sll_480_ML_int_1__52_) );
  MUX2_X2 u4_sll_480_M1_0_53 ( .A(fract_denorm[53]), .B(fract_denorm[52]), .S(
        u4_sll_480_n6), .Z(u4_sll_480_ML_int_1__53_) );
  MUX2_X2 u4_sll_480_M1_0_54 ( .A(fract_denorm[54]), .B(fract_denorm[53]), .S(
        u4_sll_480_n8), .Z(u4_sll_480_ML_int_1__54_) );
  MUX2_X2 u4_sll_480_M1_0_55 ( .A(fract_denorm[55]), .B(fract_denorm[54]), .S(
        u4_sll_480_n8), .Z(u4_sll_480_ML_int_1__55_) );
  MUX2_X2 u4_sll_480_M1_0_56 ( .A(fract_denorm[56]), .B(fract_denorm[55]), .S(
        u4_sll_480_n10), .Z(u4_sll_480_ML_int_1__56_) );
  MUX2_X2 u4_sll_480_M1_0_57 ( .A(fract_denorm[57]), .B(fract_denorm[56]), .S(
        u4_sll_480_n10), .Z(u4_sll_480_ML_int_1__57_) );
  MUX2_X2 u4_sll_480_M1_0_58 ( .A(fract_denorm[58]), .B(fract_denorm[57]), .S(
        u4_sll_480_n8), .Z(u4_sll_480_ML_int_1__58_) );
  MUX2_X2 u4_sll_480_M1_0_59 ( .A(fract_denorm[59]), .B(fract_denorm[58]), .S(
        u4_sll_480_n7), .Z(u4_sll_480_ML_int_1__59_) );
  MUX2_X2 u4_sll_480_M1_0_60 ( .A(fract_denorm[60]), .B(fract_denorm[59]), .S(
        u4_sll_480_n7), .Z(u4_sll_480_ML_int_1__60_) );
  MUX2_X2 u4_sll_480_M1_0_61 ( .A(fract_denorm[61]), .B(fract_denorm[60]), .S(
        u4_sll_480_n7), .Z(u4_sll_480_ML_int_1__61_) );
  MUX2_X2 u4_sll_480_M1_0_62 ( .A(fract_denorm[62]), .B(fract_denorm[61]), .S(
        u4_sll_480_n7), .Z(u4_sll_480_ML_int_1__62_) );
  MUX2_X2 u4_sll_480_M1_0_63 ( .A(fract_denorm[63]), .B(fract_denorm[62]), .S(
        u4_sll_480_n7), .Z(u4_sll_480_ML_int_1__63_) );
  MUX2_X2 u4_sll_480_M1_0_64 ( .A(fract_denorm[64]), .B(fract_denorm[63]), .S(
        u4_sll_480_n7), .Z(u4_sll_480_ML_int_1__64_) );
  MUX2_X2 u4_sll_480_M1_0_65 ( .A(fract_denorm[65]), .B(fract_denorm[64]), .S(
        u4_sll_480_n7), .Z(u4_sll_480_ML_int_1__65_) );
  MUX2_X2 u4_sll_480_M1_0_66 ( .A(fract_denorm[66]), .B(fract_denorm[65]), .S(
        u4_sll_480_n7), .Z(u4_sll_480_ML_int_1__66_) );
  MUX2_X2 u4_sll_480_M1_0_67 ( .A(fract_denorm[67]), .B(fract_denorm[66]), .S(
        u4_sll_480_n7), .Z(u4_sll_480_ML_int_1__67_) );
  MUX2_X2 u4_sll_480_M1_0_68 ( .A(fract_denorm[68]), .B(fract_denorm[67]), .S(
        u4_sll_480_n7), .Z(u4_sll_480_ML_int_1__68_) );
  MUX2_X2 u4_sll_480_M1_0_69 ( .A(fract_denorm[69]), .B(fract_denorm[68]), .S(
        u4_sll_480_n7), .Z(u4_sll_480_ML_int_1__69_) );
  MUX2_X2 u4_sll_480_M1_0_70 ( .A(fract_denorm[70]), .B(fract_denorm[69]), .S(
        u4_sll_480_n13), .Z(u4_sll_480_ML_int_1__70_) );
  MUX2_X2 u4_sll_480_M1_0_71 ( .A(fract_denorm[71]), .B(fract_denorm[70]), .S(
        u4_sll_480_n13), .Z(u4_sll_480_ML_int_1__71_) );
  MUX2_X2 u4_sll_480_M1_0_72 ( .A(fract_denorm[72]), .B(fract_denorm[71]), .S(
        u4_sll_480_n13), .Z(u4_sll_480_ML_int_1__72_) );
  MUX2_X2 u4_sll_480_M1_0_73 ( .A(fract_denorm[73]), .B(fract_denorm[72]), .S(
        u4_sll_480_n13), .Z(u4_sll_480_ML_int_1__73_) );
  MUX2_X2 u4_sll_480_M1_0_74 ( .A(fract_denorm[74]), .B(fract_denorm[73]), .S(
        u4_sll_480_n6), .Z(u4_sll_480_ML_int_1__74_) );
  MUX2_X2 u4_sll_480_M1_0_75 ( .A(fract_denorm[75]), .B(fract_denorm[74]), .S(
        u4_sll_480_n13), .Z(u4_sll_480_ML_int_1__75_) );
  MUX2_X2 u4_sll_480_M1_0_76 ( .A(fract_denorm[76]), .B(fract_denorm[75]), .S(
        u4_sll_480_n13), .Z(u4_sll_480_ML_int_1__76_) );
  MUX2_X2 u4_sll_480_M1_0_77 ( .A(fract_denorm[77]), .B(fract_denorm[76]), .S(
        u4_sll_480_n6), .Z(u4_sll_480_ML_int_1__77_) );
  MUX2_X2 u4_sll_480_M1_0_78 ( .A(fract_denorm[78]), .B(fract_denorm[77]), .S(
        u4_sll_480_n13), .Z(u4_sll_480_ML_int_1__78_) );
  MUX2_X2 u4_sll_480_M1_0_79 ( .A(fract_denorm[79]), .B(fract_denorm[78]), .S(
        u4_sll_480_n13), .Z(u4_sll_480_ML_int_1__79_) );
  MUX2_X2 u4_sll_480_M1_0_80 ( .A(fract_denorm[80]), .B(fract_denorm[79]), .S(
        u4_sll_480_n13), .Z(u4_sll_480_ML_int_1__80_) );
  MUX2_X2 u4_sll_480_M1_0_81 ( .A(fract_denorm[81]), .B(fract_denorm[80]), .S(
        u4_sll_480_n8), .Z(u4_sll_480_ML_int_1__81_) );
  MUX2_X2 u4_sll_480_M1_0_82 ( .A(fract_denorm[82]), .B(fract_denorm[81]), .S(
        u4_sll_480_n9), .Z(u4_sll_480_ML_int_1__82_) );
  MUX2_X2 u4_sll_480_M1_0_83 ( .A(fract_denorm[83]), .B(fract_denorm[82]), .S(
        u4_sll_480_temp_int_SH_0_), .Z(u4_sll_480_ML_int_1__83_) );
  MUX2_X2 u4_sll_480_M1_0_84 ( .A(fract_denorm[84]), .B(fract_denorm[83]), .S(
        u4_sll_480_n9), .Z(u4_sll_480_ML_int_1__84_) );
  MUX2_X2 u4_sll_480_M1_0_85 ( .A(fract_denorm[85]), .B(fract_denorm[84]), .S(
        u4_sll_480_n13), .Z(u4_sll_480_ML_int_1__85_) );
  MUX2_X2 u4_sll_480_M1_0_86 ( .A(fract_denorm[86]), .B(fract_denorm[85]), .S(
        u4_sll_480_n8), .Z(u4_sll_480_ML_int_1__86_) );
  MUX2_X2 u4_sll_480_M1_0_87 ( .A(fract_denorm[87]), .B(fract_denorm[86]), .S(
        u4_sll_480_temp_int_SH_0_), .Z(u4_sll_480_ML_int_1__87_) );
  MUX2_X2 u4_sll_480_M1_0_88 ( .A(fract_denorm[88]), .B(fract_denorm[87]), .S(
        u4_sll_480_n7), .Z(u4_sll_480_ML_int_1__88_) );
  MUX2_X2 u4_sll_480_M1_0_89 ( .A(fract_denorm[89]), .B(fract_denorm[88]), .S(
        u4_sll_480_temp_int_SH_0_), .Z(u4_sll_480_ML_int_1__89_) );
  MUX2_X2 u4_sll_480_M1_0_90 ( .A(fract_denorm[90]), .B(fract_denorm[89]), .S(
        u4_sll_480_n14), .Z(u4_sll_480_ML_int_1__90_) );
  MUX2_X2 u4_sll_480_M1_0_91 ( .A(fract_denorm[91]), .B(fract_denorm[90]), .S(
        u4_sll_480_temp_int_SH_0_), .Z(u4_sll_480_ML_int_1__91_) );
  MUX2_X2 u4_sll_480_M1_0_92 ( .A(fract_denorm[92]), .B(fract_denorm[91]), .S(
        u4_sll_480_n14), .Z(u4_sll_480_ML_int_1__92_) );
  MUX2_X2 u4_sll_480_M1_0_93 ( .A(fract_denorm[93]), .B(fract_denorm[92]), .S(
        u4_sll_480_n13), .Z(u4_sll_480_ML_int_1__93_) );
  MUX2_X2 u4_sll_480_M1_0_94 ( .A(fract_denorm[94]), .B(fract_denorm[93]), .S(
        u4_sll_480_n9), .Z(u4_sll_480_ML_int_1__94_) );
  MUX2_X2 u4_sll_480_M1_0_95 ( .A(fract_denorm[95]), .B(fract_denorm[94]), .S(
        u4_sll_480_n7), .Z(u4_sll_480_ML_int_1__95_) );
  MUX2_X2 u4_sll_480_M1_0_96 ( .A(fract_denorm[96]), .B(fract_denorm[95]), .S(
        u4_sll_480_n6), .Z(u4_sll_480_ML_int_1__96_) );
  MUX2_X2 u4_sll_480_M1_0_97 ( .A(fract_denorm[97]), .B(fract_denorm[96]), .S(
        u4_sll_480_n13), .Z(u4_sll_480_ML_int_1__97_) );
  MUX2_X2 u4_sll_480_M1_0_98 ( .A(fract_denorm[98]), .B(fract_denorm[97]), .S(
        u4_sll_480_n13), .Z(u4_sll_480_ML_int_1__98_) );
  MUX2_X2 u4_sll_480_M1_0_99 ( .A(fract_denorm[99]), .B(fract_denorm[98]), .S(
        u4_sll_480_n9), .Z(u4_sll_480_ML_int_1__99_) );
  MUX2_X2 u4_sll_480_M1_0_100 ( .A(fract_denorm[100]), .B(fract_denorm[99]), 
        .S(u4_sll_480_n14), .Z(u4_sll_480_ML_int_1__100_) );
  MUX2_X2 u4_sll_480_M1_0_101 ( .A(fract_denorm[101]), .B(fract_denorm[100]), 
        .S(u4_sll_480_temp_int_SH_0_), .Z(u4_sll_480_ML_int_1__101_) );
  MUX2_X2 u4_sll_480_M1_0_102 ( .A(fract_denorm[102]), .B(fract_denorm[101]), 
        .S(u4_sll_480_n6), .Z(u4_sll_480_ML_int_1__102_) );
  MUX2_X2 u4_sll_480_M1_0_103 ( .A(fract_denorm[103]), .B(fract_denorm[102]), 
        .S(u4_sll_480_n6), .Z(u4_sll_480_ML_int_1__103_) );
  MUX2_X2 u4_sll_480_M1_0_104 ( .A(fract_denorm[104]), .B(fract_denorm[103]), 
        .S(u4_sll_480_n6), .Z(u4_sll_480_ML_int_1__104_) );
  MUX2_X2 u4_sll_480_M1_0_105 ( .A(n4873), .B(fract_denorm[104]), .S(
        u4_sll_480_n6), .Z(u4_sll_480_ML_int_1__105_) );
  MUX2_X2 u4_sll_480_M1_0_106 ( .A(n4873), .B(n4873), .S(u4_sll_480_n6), .Z(
        u4_sll_480_ML_int_1__106_) );
  MUX2_X2 u4_sll_480_M1_0_107 ( .A(n4873), .B(n4873), .S(u4_sll_480_n6), .Z(
        u4_sll_480_ML_int_1__107_) );
  MUX2_X2 u4_sll_480_M1_0_108 ( .A(n4873), .B(n4873), .S(u4_sll_480_n6), .Z(
        u4_sll_480_ML_int_1__108_) );
  MUX2_X2 u4_sll_480_M1_0_109 ( .A(n4873), .B(n4873), .S(u4_sll_480_n6), .Z(
        u4_sll_480_ML_int_1__109_) );
  MUX2_X2 u4_sll_480_M1_0_110 ( .A(n4873), .B(n4873), .S(u4_sll_480_n6), .Z(
        u4_sll_480_ML_int_1__110_) );
  MUX2_X2 u4_sll_480_M1_0_111 ( .A(n4873), .B(n4873), .S(u4_sll_480_n6), .Z(
        u4_sll_480_ML_int_1__111_) );
  MUX2_X2 u4_sll_480_M1_0_112 ( .A(n4873), .B(n4873), .S(u4_sll_480_n6), .Z(
        u4_sll_480_ML_int_1__112_) );
  MUX2_X2 u4_sll_480_M1_0_113 ( .A(n4873), .B(n4873), .S(u4_sll_480_n6), .Z(
        u4_sll_480_ML_int_1__113_) );
  MUX2_X2 u4_sll_480_M1_1_2 ( .A(u4_sll_480_ML_int_1__2_), .B(
        u4_sll_480_ML_int_1__0_), .S(u4_sll_480_n16), .Z(
        u4_sll_480_ML_int_2__2_) );
  MUX2_X2 u4_sll_480_M1_1_3 ( .A(u4_sll_480_ML_int_1__3_), .B(
        u4_sll_480_ML_int_1__1_), .S(u4_sll_480_n16), .Z(
        u4_sll_480_ML_int_2__3_) );
  MUX2_X2 u4_sll_480_M1_1_4 ( .A(u4_sll_480_ML_int_1__4_), .B(
        u4_sll_480_ML_int_1__2_), .S(u4_sll_480_n16), .Z(
        u4_sll_480_ML_int_2__4_) );
  MUX2_X2 u4_sll_480_M1_1_5 ( .A(u4_sll_480_ML_int_1__5_), .B(
        u4_sll_480_ML_int_1__3_), .S(u4_sll_480_n16), .Z(
        u4_sll_480_ML_int_2__5_) );
  MUX2_X2 u4_sll_480_M1_1_6 ( .A(u4_sll_480_ML_int_1__6_), .B(
        u4_sll_480_ML_int_1__4_), .S(u4_sll_480_n16), .Z(
        u4_sll_480_ML_int_2__6_) );
  MUX2_X2 u4_sll_480_M1_1_7 ( .A(u4_sll_480_ML_int_1__7_), .B(
        u4_sll_480_ML_int_1__5_), .S(u4_sll_480_n16), .Z(
        u4_sll_480_ML_int_2__7_) );
  MUX2_X2 u4_sll_480_M1_1_8 ( .A(u4_sll_480_ML_int_1__8_), .B(
        u4_sll_480_ML_int_1__6_), .S(u4_sll_480_n16), .Z(
        u4_sll_480_ML_int_2__8_) );
  MUX2_X2 u4_sll_480_M1_1_9 ( .A(u4_sll_480_ML_int_1__9_), .B(
        u4_sll_480_ML_int_1__7_), .S(u4_sll_480_n16), .Z(
        u4_sll_480_ML_int_2__9_) );
  MUX2_X2 u4_sll_480_M1_1_10 ( .A(u4_sll_480_ML_int_1__10_), .B(
        u4_sll_480_ML_int_1__8_), .S(u4_sll_480_n16), .Z(
        u4_sll_480_ML_int_2__10_) );
  MUX2_X2 u4_sll_480_M1_1_11 ( .A(u4_sll_480_ML_int_1__11_), .B(
        u4_sll_480_ML_int_1__9_), .S(u4_sll_480_n16), .Z(
        u4_sll_480_ML_int_2__11_) );
  MUX2_X2 u4_sll_480_M1_1_12 ( .A(u4_sll_480_ML_int_1__12_), .B(
        u4_sll_480_ML_int_1__10_), .S(u4_sll_480_n16), .Z(
        u4_sll_480_ML_int_2__12_) );
  MUX2_X2 u4_sll_480_M1_1_13 ( .A(u4_sll_480_ML_int_1__13_), .B(
        u4_sll_480_ML_int_1__11_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__13_) );
  MUX2_X2 u4_sll_480_M1_1_14 ( .A(u4_sll_480_ML_int_1__14_), .B(
        u4_sll_480_ML_int_1__12_), .S(u4_sll_480_n18), .Z(
        u4_sll_480_ML_int_2__14_) );
  MUX2_X2 u4_sll_480_M1_1_15 ( .A(u4_sll_480_ML_int_1__15_), .B(
        u4_sll_480_ML_int_1__13_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__15_) );
  MUX2_X2 u4_sll_480_M1_1_16 ( .A(u4_sll_480_ML_int_1__16_), .B(
        u4_sll_480_ML_int_1__14_), .S(u4_sll_480_n16), .Z(
        u4_sll_480_ML_int_2__16_) );
  MUX2_X2 u4_sll_480_M1_1_17 ( .A(u4_sll_480_ML_int_1__17_), .B(
        u4_sll_480_ML_int_1__15_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__17_) );
  MUX2_X2 u4_sll_480_M1_1_18 ( .A(u4_sll_480_ML_int_1__18_), .B(
        u4_sll_480_ML_int_1__16_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__18_) );
  MUX2_X2 u4_sll_480_M1_1_19 ( .A(u4_sll_480_ML_int_1__19_), .B(
        u4_sll_480_ML_int_1__17_), .S(u4_sll_480_n18), .Z(
        u4_sll_480_ML_int_2__19_) );
  MUX2_X2 u4_sll_480_M1_1_20 ( .A(u4_sll_480_ML_int_1__20_), .B(
        u4_sll_480_ML_int_1__18_), .S(u4_sll_480_n20), .Z(
        u4_sll_480_ML_int_2__20_) );
  MUX2_X2 u4_sll_480_M1_1_21 ( .A(u4_sll_480_ML_int_1__21_), .B(
        u4_sll_480_ML_int_1__19_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__21_) );
  MUX2_X2 u4_sll_480_M1_1_22 ( .A(u4_sll_480_ML_int_1__22_), .B(
        u4_sll_480_ML_int_1__20_), .S(u4_sll_480_n16), .Z(
        u4_sll_480_ML_int_2__22_) );
  MUX2_X2 u4_sll_480_M1_1_23 ( .A(u4_sll_480_ML_int_1__23_), .B(
        u4_sll_480_ML_int_1__21_), .S(u4_sll_480_n18), .Z(
        u4_sll_480_ML_int_2__23_) );
  MUX2_X2 u4_sll_480_M1_1_24 ( .A(u4_sll_480_ML_int_1__24_), .B(
        u4_sll_480_ML_int_1__22_), .S(u4_sll_480_n17), .Z(
        u4_sll_480_ML_int_2__24_) );
  MUX2_X2 u4_sll_480_M1_1_25 ( .A(u4_sll_480_ML_int_1__25_), .B(
        u4_sll_480_ML_int_1__23_), .S(u4_sll_480_n17), .Z(
        u4_sll_480_ML_int_2__25_) );
  MUX2_X2 u4_sll_480_M1_1_26 ( .A(u4_sll_480_ML_int_1__26_), .B(
        u4_sll_480_ML_int_1__24_), .S(u4_sll_480_n17), .Z(
        u4_sll_480_ML_int_2__26_) );
  MUX2_X2 u4_sll_480_M1_1_27 ( .A(u4_sll_480_ML_int_1__27_), .B(
        u4_sll_480_ML_int_1__25_), .S(u4_sll_480_n17), .Z(
        u4_sll_480_ML_int_2__27_) );
  MUX2_X2 u4_sll_480_M1_1_28 ( .A(u4_sll_480_ML_int_1__28_), .B(
        u4_sll_480_ML_int_1__26_), .S(u4_sll_480_n17), .Z(
        u4_sll_480_ML_int_2__28_) );
  MUX2_X2 u4_sll_480_M1_1_29 ( .A(u4_sll_480_ML_int_1__29_), .B(
        u4_sll_480_ML_int_1__27_), .S(u4_sll_480_n17), .Z(
        u4_sll_480_ML_int_2__29_) );
  MUX2_X2 u4_sll_480_M1_1_30 ( .A(u4_sll_480_ML_int_1__30_), .B(
        u4_sll_480_ML_int_1__28_), .S(u4_sll_480_n17), .Z(
        u4_sll_480_ML_int_2__30_) );
  MUX2_X2 u4_sll_480_M1_1_31 ( .A(u4_sll_480_ML_int_1__31_), .B(
        u4_sll_480_ML_int_1__29_), .S(u4_sll_480_n17), .Z(
        u4_sll_480_ML_int_2__31_) );
  MUX2_X2 u4_sll_480_M1_1_32 ( .A(u4_sll_480_ML_int_1__32_), .B(
        u4_sll_480_ML_int_1__30_), .S(u4_sll_480_n17), .Z(
        u4_sll_480_ML_int_2__32_) );
  MUX2_X2 u4_sll_480_M1_1_33 ( .A(u4_sll_480_ML_int_1__33_), .B(
        u4_sll_480_ML_int_1__31_), .S(u4_sll_480_n17), .Z(
        u4_sll_480_ML_int_2__33_) );
  MUX2_X2 u4_sll_480_M1_1_34 ( .A(u4_sll_480_ML_int_1__34_), .B(
        u4_sll_480_ML_int_1__32_), .S(u4_sll_480_n17), .Z(
        u4_sll_480_ML_int_2__34_) );
  MUX2_X2 u4_sll_480_M1_1_35 ( .A(u4_sll_480_ML_int_1__35_), .B(
        u4_sll_480_ML_int_1__33_), .S(u4_sll_480_n18), .Z(
        u4_sll_480_ML_int_2__35_) );
  MUX2_X2 u4_sll_480_M1_1_36 ( .A(u4_sll_480_ML_int_1__36_), .B(
        u4_sll_480_ML_int_1__34_), .S(u4_sll_480_n18), .Z(
        u4_sll_480_ML_int_2__36_) );
  MUX2_X2 u4_sll_480_M1_1_37 ( .A(u4_sll_480_ML_int_1__37_), .B(
        u4_sll_480_ML_int_1__35_), .S(u4_sll_480_n18), .Z(
        u4_sll_480_ML_int_2__37_) );
  MUX2_X2 u4_sll_480_M1_1_38 ( .A(u4_sll_480_ML_int_1__38_), .B(
        u4_sll_480_ML_int_1__36_), .S(u4_sll_480_n18), .Z(
        u4_sll_480_ML_int_2__38_) );
  MUX2_X2 u4_sll_480_M1_1_39 ( .A(u4_sll_480_ML_int_1__39_), .B(
        u4_sll_480_ML_int_1__37_), .S(u4_sll_480_n18), .Z(
        u4_sll_480_ML_int_2__39_) );
  MUX2_X2 u4_sll_480_M1_1_40 ( .A(u4_sll_480_ML_int_1__40_), .B(
        u4_sll_480_ML_int_1__38_), .S(u4_sll_480_n18), .Z(
        u4_sll_480_ML_int_2__40_) );
  MUX2_X2 u4_sll_480_M1_1_41 ( .A(u4_sll_480_ML_int_1__41_), .B(
        u4_sll_480_ML_int_1__39_), .S(u4_sll_480_n18), .Z(
        u4_sll_480_ML_int_2__41_) );
  MUX2_X2 u4_sll_480_M1_1_42 ( .A(u4_sll_480_ML_int_1__42_), .B(
        u4_sll_480_ML_int_1__40_), .S(u4_sll_480_n18), .Z(
        u4_sll_480_ML_int_2__42_) );
  MUX2_X2 u4_sll_480_M1_1_43 ( .A(u4_sll_480_ML_int_1__43_), .B(
        u4_sll_480_ML_int_1__41_), .S(u4_sll_480_n18), .Z(
        u4_sll_480_ML_int_2__43_) );
  MUX2_X2 u4_sll_480_M1_1_44 ( .A(u4_sll_480_ML_int_1__44_), .B(
        u4_sll_480_ML_int_1__42_), .S(u4_sll_480_n18), .Z(
        u4_sll_480_ML_int_2__44_) );
  MUX2_X2 u4_sll_480_M1_1_45 ( .A(u4_sll_480_ML_int_1__45_), .B(
        u4_sll_480_ML_int_1__43_), .S(u4_sll_480_n18), .Z(
        u4_sll_480_ML_int_2__45_) );
  MUX2_X2 u4_sll_480_M1_1_46 ( .A(u4_sll_480_ML_int_1__46_), .B(
        u4_sll_480_ML_int_1__44_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__46_) );
  MUX2_X2 u4_sll_480_M1_1_47 ( .A(u4_sll_480_ML_int_1__47_), .B(
        u4_sll_480_ML_int_1__45_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__47_) );
  MUX2_X2 u4_sll_480_M1_1_48 ( .A(u4_sll_480_ML_int_1__48_), .B(
        u4_sll_480_ML_int_1__46_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__48_) );
  MUX2_X2 u4_sll_480_M1_1_49 ( .A(u4_sll_480_ML_int_1__49_), .B(
        u4_sll_480_ML_int_1__47_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__49_) );
  MUX2_X2 u4_sll_480_M1_1_50 ( .A(u4_sll_480_ML_int_1__50_), .B(
        u4_sll_480_ML_int_1__48_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__50_) );
  MUX2_X2 u4_sll_480_M1_1_51 ( .A(u4_sll_480_ML_int_1__51_), .B(
        u4_sll_480_ML_int_1__49_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__51_) );
  MUX2_X2 u4_sll_480_M1_1_52 ( .A(u4_sll_480_ML_int_1__52_), .B(
        u4_sll_480_ML_int_1__50_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__52_) );
  MUX2_X2 u4_sll_480_M1_1_53 ( .A(u4_sll_480_ML_int_1__53_), .B(
        u4_sll_480_ML_int_1__51_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__53_) );
  MUX2_X2 u4_sll_480_M1_1_54 ( .A(u4_sll_480_ML_int_1__54_), .B(
        u4_sll_480_ML_int_1__52_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__54_) );
  MUX2_X2 u4_sll_480_M1_1_55 ( .A(u4_sll_480_ML_int_1__55_), .B(
        u4_sll_480_ML_int_1__53_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__55_) );
  MUX2_X2 u4_sll_480_M1_1_56 ( .A(u4_sll_480_ML_int_1__56_), .B(
        u4_sll_480_ML_int_1__54_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__56_) );
  MUX2_X2 u4_sll_480_M1_1_57 ( .A(u4_sll_480_ML_int_1__57_), .B(
        u4_sll_480_ML_int_1__55_), .S(u4_sll_480_n19), .Z(
        u4_sll_480_ML_int_2__57_) );
  MUX2_X2 u4_sll_480_M1_1_58 ( .A(u4_sll_480_ML_int_1__58_), .B(
        u4_sll_480_ML_int_1__56_), .S(u4_sll_480_n19), .Z(
        u4_sll_480_ML_int_2__58_) );
  MUX2_X2 u4_sll_480_M1_1_59 ( .A(u4_sll_480_ML_int_1__59_), .B(
        u4_sll_480_ML_int_1__57_), .S(u4_sll_480_n19), .Z(
        u4_sll_480_ML_int_2__59_) );
  MUX2_X2 u4_sll_480_M1_1_60 ( .A(u4_sll_480_ML_int_1__60_), .B(
        u4_sll_480_ML_int_1__58_), .S(u4_sll_480_n19), .Z(
        u4_sll_480_ML_int_2__60_) );
  MUX2_X2 u4_sll_480_M1_1_61 ( .A(u4_sll_480_ML_int_1__61_), .B(
        u4_sll_480_ML_int_1__59_), .S(u4_sll_480_n19), .Z(
        u4_sll_480_ML_int_2__61_) );
  MUX2_X2 u4_sll_480_M1_1_62 ( .A(u4_sll_480_ML_int_1__62_), .B(
        u4_sll_480_ML_int_1__60_), .S(u4_sll_480_n19), .Z(
        u4_sll_480_ML_int_2__62_) );
  MUX2_X2 u4_sll_480_M1_1_63 ( .A(u4_sll_480_ML_int_1__63_), .B(
        u4_sll_480_ML_int_1__61_), .S(u4_sll_480_n19), .Z(
        u4_sll_480_ML_int_2__63_) );
  MUX2_X2 u4_sll_480_M1_1_64 ( .A(u4_sll_480_ML_int_1__64_), .B(
        u4_sll_480_ML_int_1__62_), .S(u4_sll_480_n19), .Z(
        u4_sll_480_ML_int_2__64_) );
  MUX2_X2 u4_sll_480_M1_1_65 ( .A(u4_sll_480_ML_int_1__65_), .B(
        u4_sll_480_ML_int_1__63_), .S(u4_sll_480_n19), .Z(
        u4_sll_480_ML_int_2__65_) );
  MUX2_X2 u4_sll_480_M1_1_66 ( .A(u4_sll_480_ML_int_1__66_), .B(
        u4_sll_480_ML_int_1__64_), .S(u4_sll_480_n19), .Z(
        u4_sll_480_ML_int_2__66_) );
  MUX2_X2 u4_sll_480_M1_1_67 ( .A(u4_sll_480_ML_int_1__67_), .B(
        u4_sll_480_ML_int_1__65_), .S(u4_sll_480_n19), .Z(
        u4_sll_480_ML_int_2__67_) );
  MUX2_X2 u4_sll_480_M1_1_68 ( .A(u4_sll_480_ML_int_1__68_), .B(
        u4_sll_480_ML_int_1__66_), .S(u4_sll_480_n20), .Z(
        u4_sll_480_ML_int_2__68_) );
  MUX2_X2 u4_sll_480_M1_1_69 ( .A(u4_sll_480_ML_int_1__69_), .B(
        u4_sll_480_ML_int_1__67_), .S(u4_sll_480_n20), .Z(
        u4_sll_480_ML_int_2__69_) );
  MUX2_X2 u4_sll_480_M1_1_70 ( .A(u4_sll_480_ML_int_1__70_), .B(
        u4_sll_480_ML_int_1__68_), .S(u4_sll_480_n20), .Z(
        u4_sll_480_ML_int_2__70_) );
  MUX2_X2 u4_sll_480_M1_1_71 ( .A(u4_sll_480_ML_int_1__71_), .B(
        u4_sll_480_ML_int_1__69_), .S(u4_sll_480_n20), .Z(
        u4_sll_480_ML_int_2__71_) );
  MUX2_X2 u4_sll_480_M1_1_72 ( .A(u4_sll_480_ML_int_1__72_), .B(
        u4_sll_480_ML_int_1__70_), .S(u4_sll_480_n20), .Z(
        u4_sll_480_ML_int_2__72_) );
  MUX2_X2 u4_sll_480_M1_1_73 ( .A(u4_sll_480_ML_int_1__73_), .B(
        u4_sll_480_ML_int_1__71_), .S(u4_sll_480_n20), .Z(
        u4_sll_480_ML_int_2__73_) );
  MUX2_X2 u4_sll_480_M1_1_74 ( .A(u4_sll_480_ML_int_1__74_), .B(
        u4_sll_480_ML_int_1__72_), .S(u4_sll_480_n20), .Z(
        u4_sll_480_ML_int_2__74_) );
  MUX2_X2 u4_sll_480_M1_1_75 ( .A(u4_sll_480_ML_int_1__75_), .B(
        u4_sll_480_ML_int_1__73_), .S(u4_sll_480_n20), .Z(
        u4_sll_480_ML_int_2__75_) );
  MUX2_X2 u4_sll_480_M1_1_76 ( .A(u4_sll_480_ML_int_1__76_), .B(
        u4_sll_480_ML_int_1__74_), .S(u4_sll_480_n20), .Z(
        u4_sll_480_ML_int_2__76_) );
  MUX2_X2 u4_sll_480_M1_1_77 ( .A(u4_sll_480_ML_int_1__77_), .B(
        u4_sll_480_ML_int_1__75_), .S(u4_sll_480_n20), .Z(
        u4_sll_480_ML_int_2__77_) );
  MUX2_X2 u4_sll_480_M1_1_78 ( .A(u4_sll_480_ML_int_1__78_), .B(
        u4_sll_480_ML_int_1__76_), .S(u4_sll_480_n20), .Z(
        u4_sll_480_ML_int_2__78_) );
  MUX2_X2 u4_sll_480_M1_1_79 ( .A(u4_sll_480_ML_int_1__79_), .B(
        u4_sll_480_ML_int_1__77_), .S(u4_sll_480_n17), .Z(
        u4_sll_480_ML_int_2__79_) );
  MUX2_X2 u4_sll_480_M1_1_80 ( .A(u4_sll_480_ML_int_1__80_), .B(
        u4_sll_480_ML_int_1__78_), .S(u4_sll_480_n19), .Z(
        u4_sll_480_ML_int_2__80_) );
  MUX2_X2 u4_sll_480_M1_1_81 ( .A(u4_sll_480_ML_int_1__81_), .B(
        u4_sll_480_ML_int_1__79_), .S(u4_sll_480_n19), .Z(
        u4_sll_480_ML_int_2__81_) );
  MUX2_X2 u4_sll_480_M1_1_82 ( .A(u4_sll_480_ML_int_1__82_), .B(
        u4_sll_480_ML_int_1__80_), .S(u4_sll_480_n19), .Z(
        u4_sll_480_ML_int_2__82_) );
  MUX2_X2 u4_sll_480_M1_1_83 ( .A(u4_sll_480_ML_int_1__83_), .B(
        u4_sll_480_ML_int_1__81_), .S(u4_sll_480_n17), .Z(
        u4_sll_480_ML_int_2__83_) );
  MUX2_X2 u4_sll_480_M1_1_84 ( .A(u4_sll_480_ML_int_1__84_), .B(
        u4_sll_480_ML_int_1__82_), .S(u4_sll_480_n19), .Z(
        u4_sll_480_ML_int_2__84_) );
  MUX2_X2 u4_sll_480_M1_1_85 ( .A(u4_sll_480_ML_int_1__85_), .B(
        u4_sll_480_ML_int_1__83_), .S(u4_sll_480_n19), .Z(
        u4_sll_480_ML_int_2__85_) );
  MUX2_X2 u4_sll_480_M1_1_86 ( .A(u4_sll_480_ML_int_1__86_), .B(
        u4_sll_480_ML_int_1__84_), .S(u4_sll_480_n19), .Z(
        u4_sll_480_ML_int_2__86_) );
  MUX2_X2 u4_sll_480_M1_1_87 ( .A(u4_sll_480_ML_int_1__87_), .B(
        u4_sll_480_ML_int_1__85_), .S(u4_sll_480_n17), .Z(
        u4_sll_480_ML_int_2__87_) );
  MUX2_X2 u4_sll_480_M1_1_88 ( .A(u4_sll_480_ML_int_1__88_), .B(
        u4_sll_480_ML_int_1__86_), .S(u4_sll_480_n19), .Z(
        u4_sll_480_ML_int_2__88_) );
  MUX2_X2 u4_sll_480_M1_1_89 ( .A(u4_sll_480_ML_int_1__89_), .B(
        u4_sll_480_ML_int_1__87_), .S(u4_sll_480_n19), .Z(
        u4_sll_480_ML_int_2__89_) );
  MUX2_X2 u4_sll_480_M1_1_90 ( .A(u4_sll_480_ML_int_1__90_), .B(
        u4_sll_480_ML_int_1__88_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__90_) );
  MUX2_X2 u4_sll_480_M1_1_91 ( .A(u4_sll_480_ML_int_1__91_), .B(
        u4_sll_480_ML_int_1__89_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__91_) );
  MUX2_X2 u4_sll_480_M1_1_92 ( .A(u4_sll_480_ML_int_1__92_), .B(
        u4_sll_480_ML_int_1__90_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__92_) );
  MUX2_X2 u4_sll_480_M1_1_93 ( .A(u4_sll_480_ML_int_1__93_), .B(
        u4_sll_480_ML_int_1__91_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__93_) );
  MUX2_X2 u4_sll_480_M1_1_94 ( .A(u4_sll_480_ML_int_1__94_), .B(
        u4_sll_480_ML_int_1__92_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__94_) );
  MUX2_X2 u4_sll_480_M1_1_95 ( .A(u4_sll_480_ML_int_1__95_), .B(
        u4_sll_480_ML_int_1__93_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__95_) );
  MUX2_X2 u4_sll_480_M1_1_96 ( .A(u4_sll_480_ML_int_1__96_), .B(
        u4_sll_480_ML_int_1__94_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__96_) );
  MUX2_X2 u4_sll_480_M1_1_97 ( .A(u4_sll_480_ML_int_1__97_), .B(
        u4_sll_480_ML_int_1__95_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__97_) );
  MUX2_X2 u4_sll_480_M1_1_98 ( .A(u4_sll_480_ML_int_1__98_), .B(
        u4_sll_480_ML_int_1__96_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__98_) );
  MUX2_X2 u4_sll_480_M1_1_99 ( .A(u4_sll_480_ML_int_1__99_), .B(
        u4_sll_480_ML_int_1__97_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__99_) );
  MUX2_X2 u4_sll_480_M1_1_100 ( .A(u4_sll_480_ML_int_1__100_), .B(
        u4_sll_480_ML_int_1__98_), .S(u4_sll_480_n21), .Z(
        u4_sll_480_ML_int_2__100_) );
  MUX2_X2 u4_sll_480_M1_1_101 ( .A(u4_sll_480_ML_int_1__101_), .B(
        u4_sll_480_ML_int_1__99_), .S(u4_sll_480_n22), .Z(
        u4_sll_480_ML_int_2__101_) );
  MUX2_X2 u4_sll_480_M1_1_102 ( .A(u4_sll_480_ML_int_1__102_), .B(
        u4_sll_480_ML_int_1__100_), .S(u4_sll_480_n22), .Z(
        u4_sll_480_ML_int_2__102_) );
  MUX2_X2 u4_sll_480_M1_1_103 ( .A(u4_sll_480_ML_int_1__103_), .B(
        u4_sll_480_ML_int_1__101_), .S(u4_sll_480_n22), .Z(
        u4_sll_480_ML_int_2__103_) );
  MUX2_X2 u4_sll_480_M1_1_104 ( .A(u4_sll_480_ML_int_1__104_), .B(
        u4_sll_480_ML_int_1__102_), .S(u4_sll_480_n22), .Z(
        u4_sll_480_ML_int_2__104_) );
  MUX2_X2 u4_sll_480_M1_1_105 ( .A(u4_sll_480_ML_int_1__105_), .B(
        u4_sll_480_ML_int_1__103_), .S(u4_sll_480_n22), .Z(
        u4_sll_480_ML_int_2__105_) );
  MUX2_X2 u4_sll_480_M1_1_106 ( .A(u4_sll_480_ML_int_1__106_), .B(
        u4_sll_480_ML_int_1__104_), .S(u4_sll_480_n22), .Z(
        u4_sll_480_ML_int_2__106_) );
  MUX2_X2 u4_sll_480_M1_1_107 ( .A(u4_sll_480_ML_int_1__107_), .B(
        u4_sll_480_ML_int_1__105_), .S(u4_sll_480_n22), .Z(
        u4_sll_480_ML_int_2__107_) );
  MUX2_X2 u4_sll_480_M1_1_108 ( .A(u4_sll_480_ML_int_1__108_), .B(
        u4_sll_480_ML_int_1__106_), .S(u4_sll_480_n22), .Z(
        u4_sll_480_ML_int_2__108_) );
  MUX2_X2 u4_sll_480_M1_1_109 ( .A(u4_sll_480_ML_int_1__109_), .B(
        u4_sll_480_ML_int_1__107_), .S(u4_sll_480_n22), .Z(
        u4_sll_480_ML_int_2__109_) );
  MUX2_X2 u4_sll_480_M1_1_110 ( .A(u4_sll_480_ML_int_1__110_), .B(
        u4_sll_480_ML_int_1__108_), .S(u4_sll_480_n22), .Z(
        u4_sll_480_ML_int_2__110_) );
  MUX2_X2 u4_sll_480_M1_1_111 ( .A(u4_sll_480_ML_int_1__111_), .B(
        u4_sll_480_ML_int_1__109_), .S(u4_sll_480_n22), .Z(
        u4_sll_480_ML_int_2__111_) );
  MUX2_X2 u4_sll_480_M1_1_112 ( .A(u4_sll_480_ML_int_1__112_), .B(
        u4_sll_480_ML_int_1__110_), .S(u4_sll_480_n22), .Z(
        u4_sll_480_ML_int_2__112_) );
  MUX2_X2 u4_sll_480_M1_1_113 ( .A(u4_sll_480_ML_int_1__113_), .B(
        u4_sll_480_ML_int_1__111_), .S(u4_sll_480_n22), .Z(
        u4_sll_480_ML_int_2__113_) );
  MUX2_X2 u4_sll_480_M1_1_114 ( .A(u4_sll_480_MR_int_1__113_), .B(
        u4_sll_480_ML_int_1__112_), .S(u4_sll_480_n22), .Z(
        u4_sll_480_ML_int_2__114_) );
  MUX2_X2 u4_sll_480_M1_2_4 ( .A(u4_sll_480_ML_int_2__4_), .B(u4_sll_480_n38), 
        .S(u4_sll_480_n23), .Z(u4_sll_480_ML_int_3__4_) );
  MUX2_X2 u4_sll_480_M1_2_5 ( .A(u4_sll_480_ML_int_2__5_), .B(u4_sll_480_n40), 
        .S(u4_sll_480_n23), .Z(u4_sll_480_ML_int_3__5_) );
  MUX2_X2 u4_sll_480_M1_2_6 ( .A(u4_sll_480_ML_int_2__6_), .B(
        u4_sll_480_ML_int_2__2_), .S(u4_sll_480_n23), .Z(
        u4_sll_480_ML_int_3__6_) );
  MUX2_X2 u4_sll_480_M1_2_7 ( .A(u4_sll_480_ML_int_2__7_), .B(
        u4_sll_480_ML_int_2__3_), .S(u4_sll_480_n23), .Z(
        u4_sll_480_ML_int_3__7_) );
  MUX2_X2 u4_sll_480_M1_2_8 ( .A(u4_sll_480_ML_int_2__8_), .B(
        u4_sll_480_ML_int_2__4_), .S(u4_sll_480_n23), .Z(
        u4_sll_480_ML_int_3__8_) );
  MUX2_X2 u4_sll_480_M1_2_9 ( .A(u4_sll_480_ML_int_2__9_), .B(
        u4_sll_480_ML_int_2__5_), .S(u4_sll_480_n23), .Z(
        u4_sll_480_ML_int_3__9_) );
  MUX2_X2 u4_sll_480_M1_2_10 ( .A(u4_sll_480_ML_int_2__10_), .B(
        u4_sll_480_ML_int_2__6_), .S(u4_sll_480_n23), .Z(
        u4_sll_480_ML_int_3__10_) );
  MUX2_X2 u4_sll_480_M1_2_11 ( .A(u4_sll_480_ML_int_2__11_), .B(
        u4_sll_480_ML_int_2__7_), .S(u4_sll_480_n23), .Z(
        u4_sll_480_ML_int_3__11_) );
  MUX2_X2 u4_sll_480_M1_2_12 ( .A(u4_sll_480_ML_int_2__12_), .B(
        u4_sll_480_ML_int_2__8_), .S(u4_sll_480_n23), .Z(
        u4_sll_480_ML_int_3__12_) );
  MUX2_X2 u4_sll_480_M1_2_13 ( .A(u4_sll_480_ML_int_2__13_), .B(
        u4_sll_480_ML_int_2__9_), .S(u4_sll_480_n23), .Z(
        u4_sll_480_ML_int_3__13_) );
  MUX2_X2 u4_sll_480_M1_2_14 ( .A(u4_sll_480_ML_int_2__14_), .B(
        u4_sll_480_ML_int_2__10_), .S(u4_sll_480_n23), .Z(
        u4_sll_480_ML_int_3__14_) );
  MUX2_X2 u4_sll_480_M1_2_15 ( .A(u4_sll_480_ML_int_2__15_), .B(
        u4_sll_480_ML_int_2__11_), .S(u4_sll_480_n24), .Z(
        u4_sll_480_ML_int_3__15_) );
  MUX2_X2 u4_sll_480_M1_2_16 ( .A(u4_sll_480_ML_int_2__16_), .B(
        u4_sll_480_ML_int_2__12_), .S(u4_sll_480_n24), .Z(
        u4_sll_480_ML_int_3__16_) );
  MUX2_X2 u4_sll_480_M1_2_17 ( .A(u4_sll_480_ML_int_2__17_), .B(
        u4_sll_480_ML_int_2__13_), .S(u4_sll_480_n24), .Z(
        u4_sll_480_ML_int_3__17_) );
  MUX2_X2 u4_sll_480_M1_2_18 ( .A(u4_sll_480_ML_int_2__18_), .B(
        u4_sll_480_ML_int_2__14_), .S(u4_sll_480_n24), .Z(
        u4_sll_480_ML_int_3__18_) );
  MUX2_X2 u4_sll_480_M1_2_19 ( .A(u4_sll_480_ML_int_2__19_), .B(
        u4_sll_480_ML_int_2__15_), .S(u4_sll_480_n24), .Z(
        u4_sll_480_ML_int_3__19_) );
  MUX2_X2 u4_sll_480_M1_2_20 ( .A(u4_sll_480_ML_int_2__20_), .B(
        u4_sll_480_ML_int_2__16_), .S(u4_sll_480_n24), .Z(
        u4_sll_480_ML_int_3__20_) );
  MUX2_X2 u4_sll_480_M1_2_21 ( .A(u4_sll_480_ML_int_2__21_), .B(
        u4_sll_480_ML_int_2__17_), .S(u4_sll_480_n24), .Z(
        u4_sll_480_ML_int_3__21_) );
  MUX2_X2 u4_sll_480_M1_2_22 ( .A(u4_sll_480_ML_int_2__22_), .B(
        u4_sll_480_ML_int_2__18_), .S(u4_sll_480_n24), .Z(
        u4_sll_480_ML_int_3__22_) );
  MUX2_X2 u4_sll_480_M1_2_23 ( .A(u4_sll_480_ML_int_2__23_), .B(
        u4_sll_480_ML_int_2__19_), .S(u4_sll_480_n24), .Z(
        u4_sll_480_ML_int_3__23_) );
  MUX2_X2 u4_sll_480_M1_2_24 ( .A(u4_sll_480_ML_int_2__24_), .B(
        u4_sll_480_ML_int_2__20_), .S(u4_sll_480_n24), .Z(
        u4_sll_480_ML_int_3__24_) );
  MUX2_X2 u4_sll_480_M1_2_25 ( .A(u4_sll_480_ML_int_2__25_), .B(
        u4_sll_480_ML_int_2__21_), .S(u4_sll_480_n24), .Z(
        u4_sll_480_ML_int_3__25_) );
  MUX2_X2 u4_sll_480_M1_2_26 ( .A(u4_sll_480_ML_int_2__26_), .B(
        u4_sll_480_ML_int_2__22_), .S(u4_sll_480_n23), .Z(
        u4_sll_480_ML_int_3__26_) );
  MUX2_X2 u4_sll_480_M1_2_27 ( .A(u4_sll_480_ML_int_2__27_), .B(
        u4_sll_480_ML_int_2__23_), .S(u4_sll_480_n29), .Z(
        u4_sll_480_ML_int_3__27_) );
  MUX2_X2 u4_sll_480_M1_2_28 ( .A(u4_sll_480_ML_int_2__28_), .B(
        u4_sll_480_ML_int_2__24_), .S(u4_sll_480_n28), .Z(
        u4_sll_480_ML_int_3__28_) );
  MUX2_X2 u4_sll_480_M1_2_29 ( .A(u4_sll_480_ML_int_2__29_), .B(
        u4_sll_480_ML_int_2__25_), .S(u4_sll_480_n29), .Z(
        u4_sll_480_ML_int_3__29_) );
  MUX2_X2 u4_sll_480_M1_2_30 ( .A(u4_sll_480_ML_int_2__30_), .B(
        u4_sll_480_ML_int_2__26_), .S(u4_sll_480_n25), .Z(
        u4_sll_480_ML_int_3__30_) );
  MUX2_X2 u4_sll_480_M1_2_31 ( .A(u4_sll_480_ML_int_2__31_), .B(
        u4_sll_480_ML_int_2__27_), .S(u4_sll_480_n25), .Z(
        u4_sll_480_ML_int_3__31_) );
  MUX2_X2 u4_sll_480_M1_2_32 ( .A(u4_sll_480_ML_int_2__32_), .B(
        u4_sll_480_ML_int_2__28_), .S(u4_sll_480_n25), .Z(
        u4_sll_480_ML_int_3__32_) );
  MUX2_X2 u4_sll_480_M1_2_33 ( .A(u4_sll_480_ML_int_2__33_), .B(
        u4_sll_480_ML_int_2__29_), .S(u4_sll_480_n28), .Z(
        u4_sll_480_ML_int_3__33_) );
  MUX2_X2 u4_sll_480_M1_2_34 ( .A(u4_sll_480_ML_int_2__34_), .B(
        u4_sll_480_ML_int_2__30_), .S(u4_sll_480_n29), .Z(
        u4_sll_480_ML_int_3__34_) );
  MUX2_X2 u4_sll_480_M1_2_35 ( .A(u4_sll_480_ML_int_2__35_), .B(
        u4_sll_480_ML_int_2__31_), .S(u4_sll_480_n28), .Z(
        u4_sll_480_ML_int_3__35_) );
  MUX2_X2 u4_sll_480_M1_2_36 ( .A(u4_sll_480_ML_int_2__36_), .B(
        u4_sll_480_ML_int_2__32_), .S(u4_sll_480_n25), .Z(
        u4_sll_480_ML_int_3__36_) );
  MUX2_X2 u4_sll_480_M1_2_37 ( .A(u4_sll_480_ML_int_2__37_), .B(
        u4_sll_480_ML_int_2__33_), .S(u4_sll_480_n25), .Z(
        u4_sll_480_ML_int_3__37_) );
  MUX2_X2 u4_sll_480_M1_2_38 ( .A(u4_sll_480_ML_int_2__38_), .B(
        u4_sll_480_ML_int_2__34_), .S(u4_sll_480_n25), .Z(
        u4_sll_480_ML_int_3__38_) );
  MUX2_X2 u4_sll_480_M1_2_39 ( .A(u4_sll_480_ML_int_2__39_), .B(
        u4_sll_480_ML_int_2__35_), .S(u4_sll_480_n25), .Z(
        u4_sll_480_ML_int_3__39_) );
  MUX2_X2 u4_sll_480_M1_2_40 ( .A(u4_sll_480_ML_int_2__40_), .B(
        u4_sll_480_ML_int_2__36_), .S(u4_sll_480_n25), .Z(
        u4_sll_480_ML_int_3__40_) );
  MUX2_X2 u4_sll_480_M1_2_41 ( .A(u4_sll_480_ML_int_2__41_), .B(
        u4_sll_480_ML_int_2__37_), .S(u4_sll_480_n25), .Z(
        u4_sll_480_ML_int_3__41_) );
  MUX2_X2 u4_sll_480_M1_2_42 ( .A(u4_sll_480_ML_int_2__42_), .B(
        u4_sll_480_ML_int_2__38_), .S(u4_sll_480_n25), .Z(
        u4_sll_480_ML_int_3__42_) );
  MUX2_X2 u4_sll_480_M1_2_43 ( .A(u4_sll_480_ML_int_2__43_), .B(
        u4_sll_480_ML_int_2__39_), .S(u4_sll_480_n25), .Z(
        u4_sll_480_ML_int_3__43_) );
  MUX2_X2 u4_sll_480_M1_2_44 ( .A(u4_sll_480_ML_int_2__44_), .B(
        u4_sll_480_ML_int_2__40_), .S(u4_sll_480_n25), .Z(
        u4_sll_480_ML_int_3__44_) );
  MUX2_X2 u4_sll_480_M1_2_45 ( .A(u4_sll_480_ML_int_2__45_), .B(
        u4_sll_480_ML_int_2__41_), .S(u4_sll_480_n25), .Z(
        u4_sll_480_ML_int_3__45_) );
  MUX2_X2 u4_sll_480_M1_2_46 ( .A(u4_sll_480_ML_int_2__46_), .B(
        u4_sll_480_ML_int_2__42_), .S(u4_sll_480_n25), .Z(
        u4_sll_480_ML_int_3__46_) );
  MUX2_X2 u4_sll_480_M1_2_47 ( .A(u4_sll_480_ML_int_2__47_), .B(
        u4_sll_480_ML_int_2__43_), .S(u4_sll_480_n25), .Z(
        u4_sll_480_ML_int_3__47_) );
  MUX2_X2 u4_sll_480_M1_2_48 ( .A(u4_sll_480_ML_int_2__48_), .B(
        u4_sll_480_ML_int_2__44_), .S(u4_sll_480_n24), .Z(
        u4_sll_480_ML_int_3__48_) );
  MUX2_X2 u4_sll_480_M1_2_49 ( .A(u4_sll_480_ML_int_2__49_), .B(
        u4_sll_480_ML_int_2__45_), .S(u4_sll_480_n24), .Z(
        u4_sll_480_ML_int_3__49_) );
  MUX2_X2 u4_sll_480_M1_2_50 ( .A(u4_sll_480_ML_int_2__50_), .B(
        u4_sll_480_ML_int_2__46_), .S(u4_sll_480_n24), .Z(
        u4_sll_480_ML_int_3__50_) );
  MUX2_X2 u4_sll_480_M1_2_51 ( .A(u4_sll_480_ML_int_2__51_), .B(
        u4_sll_480_ML_int_2__47_), .S(u4_sll_480_n24), .Z(
        u4_sll_480_ML_int_3__51_) );
  MUX2_X2 u4_sll_480_M1_2_52 ( .A(u4_sll_480_ML_int_2__52_), .B(
        u4_sll_480_ML_int_2__48_), .S(u4_sll_480_n24), .Z(
        u4_sll_480_ML_int_3__52_) );
  MUX2_X2 u4_sll_480_M1_2_53 ( .A(u4_sll_480_ML_int_2__53_), .B(
        u4_sll_480_ML_int_2__49_), .S(u4_sll_480_n24), .Z(
        u4_sll_480_ML_int_3__53_) );
  MUX2_X2 u4_sll_480_M1_2_54 ( .A(u4_sll_480_ML_int_2__54_), .B(
        u4_sll_480_ML_int_2__50_), .S(u4_sll_480_n24), .Z(
        u4_sll_480_ML_int_3__54_) );
  MUX2_X2 u4_sll_480_M1_2_55 ( .A(u4_sll_480_ML_int_2__55_), .B(
        u4_sll_480_ML_int_2__51_), .S(u4_sll_480_n24), .Z(
        u4_sll_480_ML_int_3__55_) );
  MUX2_X2 u4_sll_480_M1_2_56 ( .A(u4_sll_480_ML_int_2__56_), .B(
        u4_sll_480_ML_int_2__52_), .S(u4_sll_480_n24), .Z(
        u4_sll_480_ML_int_3__56_) );
  MUX2_X2 u4_sll_480_M1_2_57 ( .A(u4_sll_480_ML_int_2__57_), .B(
        u4_sll_480_ML_int_2__53_), .S(u4_sll_480_n24), .Z(
        u4_sll_480_ML_int_3__57_) );
  MUX2_X2 u4_sll_480_M1_2_58 ( .A(u4_sll_480_ML_int_2__58_), .B(
        u4_sll_480_ML_int_2__54_), .S(u4_sll_480_n24), .Z(
        u4_sll_480_ML_int_3__58_) );
  MUX2_X2 u4_sll_480_M1_2_59 ( .A(u4_sll_480_ML_int_2__59_), .B(
        u4_sll_480_ML_int_2__55_), .S(u4_sll_480_n26), .Z(
        u4_sll_480_ML_int_3__59_) );
  MUX2_X2 u4_sll_480_M1_2_60 ( .A(u4_sll_480_ML_int_2__60_), .B(
        u4_sll_480_ML_int_2__56_), .S(u4_sll_480_n26), .Z(
        u4_sll_480_ML_int_3__60_) );
  MUX2_X2 u4_sll_480_M1_2_61 ( .A(u4_sll_480_ML_int_2__61_), .B(
        u4_sll_480_ML_int_2__57_), .S(u4_sll_480_n26), .Z(
        u4_sll_480_ML_int_3__61_) );
  MUX2_X2 u4_sll_480_M1_2_62 ( .A(u4_sll_480_ML_int_2__62_), .B(
        u4_sll_480_ML_int_2__58_), .S(u4_sll_480_n26), .Z(
        u4_sll_480_ML_int_3__62_) );
  MUX2_X2 u4_sll_480_M1_2_63 ( .A(u4_sll_480_ML_int_2__63_), .B(
        u4_sll_480_ML_int_2__59_), .S(u4_sll_480_n26), .Z(
        u4_sll_480_ML_int_3__63_) );
  MUX2_X2 u4_sll_480_M1_2_64 ( .A(u4_sll_480_ML_int_2__64_), .B(
        u4_sll_480_ML_int_2__60_), .S(u4_sll_480_n26), .Z(
        u4_sll_480_ML_int_3__64_) );
  MUX2_X2 u4_sll_480_M1_2_65 ( .A(u4_sll_480_ML_int_2__65_), .B(
        u4_sll_480_ML_int_2__61_), .S(u4_sll_480_n26), .Z(
        u4_sll_480_ML_int_3__65_) );
  MUX2_X2 u4_sll_480_M1_2_66 ( .A(u4_sll_480_ML_int_2__66_), .B(
        u4_sll_480_ML_int_2__62_), .S(u4_sll_480_n26), .Z(
        u4_sll_480_ML_int_3__66_) );
  MUX2_X2 u4_sll_480_M1_2_67 ( .A(u4_sll_480_ML_int_2__67_), .B(
        u4_sll_480_ML_int_2__63_), .S(u4_sll_480_n26), .Z(
        u4_sll_480_ML_int_3__67_) );
  MUX2_X2 u4_sll_480_M1_2_68 ( .A(u4_sll_480_ML_int_2__68_), .B(
        u4_sll_480_ML_int_2__64_), .S(u4_sll_480_n26), .Z(
        u4_sll_480_ML_int_3__68_) );
  MUX2_X2 u4_sll_480_M1_2_69 ( .A(u4_sll_480_ML_int_2__69_), .B(
        u4_sll_480_ML_int_2__65_), .S(u4_sll_480_n26), .Z(
        u4_sll_480_ML_int_3__69_) );
  MUX2_X2 u4_sll_480_M1_2_70 ( .A(u4_sll_480_ML_int_2__70_), .B(
        u4_sll_480_ML_int_2__66_), .S(u4_sll_480_n27), .Z(
        u4_sll_480_ML_int_3__70_) );
  MUX2_X2 u4_sll_480_M1_2_71 ( .A(u4_sll_480_ML_int_2__71_), .B(
        u4_sll_480_ML_int_2__67_), .S(u4_sll_480_n27), .Z(
        u4_sll_480_ML_int_3__71_) );
  MUX2_X2 u4_sll_480_M1_2_72 ( .A(u4_sll_480_ML_int_2__72_), .B(
        u4_sll_480_ML_int_2__68_), .S(u4_sll_480_n27), .Z(
        u4_sll_480_ML_int_3__72_) );
  MUX2_X2 u4_sll_480_M1_2_73 ( .A(u4_sll_480_ML_int_2__73_), .B(
        u4_sll_480_ML_int_2__69_), .S(u4_sll_480_n27), .Z(
        u4_sll_480_ML_int_3__73_) );
  MUX2_X2 u4_sll_480_M1_2_74 ( .A(u4_sll_480_ML_int_2__74_), .B(
        u4_sll_480_ML_int_2__70_), .S(u4_sll_480_n27), .Z(
        u4_sll_480_ML_int_3__74_) );
  MUX2_X2 u4_sll_480_M1_2_75 ( .A(u4_sll_480_ML_int_2__75_), .B(
        u4_sll_480_ML_int_2__71_), .S(u4_sll_480_n27), .Z(
        u4_sll_480_ML_int_3__75_) );
  MUX2_X2 u4_sll_480_M1_2_76 ( .A(u4_sll_480_ML_int_2__76_), .B(
        u4_sll_480_ML_int_2__72_), .S(u4_sll_480_n27), .Z(
        u4_sll_480_ML_int_3__76_) );
  MUX2_X2 u4_sll_480_M1_2_77 ( .A(u4_sll_480_ML_int_2__77_), .B(
        u4_sll_480_ML_int_2__73_), .S(u4_sll_480_n27), .Z(
        u4_sll_480_ML_int_3__77_) );
  MUX2_X2 u4_sll_480_M1_2_78 ( .A(u4_sll_480_ML_int_2__78_), .B(
        u4_sll_480_ML_int_2__74_), .S(u4_sll_480_n27), .Z(
        u4_sll_480_ML_int_3__78_) );
  MUX2_X2 u4_sll_480_M1_2_79 ( .A(u4_sll_480_ML_int_2__79_), .B(
        u4_sll_480_ML_int_2__75_), .S(u4_sll_480_n27), .Z(
        u4_sll_480_ML_int_3__79_) );
  MUX2_X2 u4_sll_480_M1_2_80 ( .A(u4_sll_480_ML_int_2__80_), .B(
        u4_sll_480_ML_int_2__76_), .S(u4_sll_480_n27), .Z(
        u4_sll_480_ML_int_3__80_) );
  MUX2_X2 u4_sll_480_M1_2_81 ( .A(u4_sll_480_ML_int_2__81_), .B(
        u4_sll_480_ML_int_2__77_), .S(u4_sll_480_n26), .Z(
        u4_sll_480_ML_int_3__81_) );
  MUX2_X2 u4_sll_480_M1_2_82 ( .A(u4_sll_480_ML_int_2__82_), .B(
        u4_sll_480_ML_int_2__78_), .S(u4_sll_480_n27), .Z(
        u4_sll_480_ML_int_3__82_) );
  MUX2_X2 u4_sll_480_M1_2_83 ( .A(u4_sll_480_ML_int_2__83_), .B(
        u4_sll_480_ML_int_2__79_), .S(u4_sll_480_n27), .Z(
        u4_sll_480_ML_int_3__83_) );
  MUX2_X2 u4_sll_480_M1_2_84 ( .A(u4_sll_480_ML_int_2__84_), .B(
        u4_sll_480_ML_int_2__80_), .S(u4_sll_480_n27), .Z(
        u4_sll_480_ML_int_3__84_) );
  MUX2_X2 u4_sll_480_M1_2_85 ( .A(u4_sll_480_ML_int_2__85_), .B(
        u4_sll_480_ML_int_2__81_), .S(u4_sll_480_n26), .Z(
        u4_sll_480_ML_int_3__85_) );
  MUX2_X2 u4_sll_480_M1_2_86 ( .A(u4_sll_480_ML_int_2__86_), .B(
        u4_sll_480_ML_int_2__82_), .S(u4_sll_480_n26), .Z(
        u4_sll_480_ML_int_3__86_) );
  MUX2_X2 u4_sll_480_M1_2_87 ( .A(u4_sll_480_ML_int_2__87_), .B(
        u4_sll_480_ML_int_2__83_), .S(u4_sll_480_n27), .Z(
        u4_sll_480_ML_int_3__87_) );
  MUX2_X2 u4_sll_480_M1_2_88 ( .A(u4_sll_480_ML_int_2__88_), .B(
        u4_sll_480_ML_int_2__84_), .S(u4_sll_480_n27), .Z(
        u4_sll_480_ML_int_3__88_) );
  MUX2_X2 u4_sll_480_M1_2_89 ( .A(u4_sll_480_ML_int_2__89_), .B(
        u4_sll_480_ML_int_2__85_), .S(u4_sll_480_n26), .Z(
        u4_sll_480_ML_int_3__89_) );
  MUX2_X2 u4_sll_480_M1_2_90 ( .A(u4_sll_480_ML_int_2__90_), .B(
        u4_sll_480_ML_int_2__86_), .S(u4_sll_480_n26), .Z(
        u4_sll_480_ML_int_3__90_) );
  MUX2_X2 u4_sll_480_M1_2_91 ( .A(u4_sll_480_ML_int_2__91_), .B(
        u4_sll_480_ML_int_2__87_), .S(u4_sll_480_n27), .Z(
        u4_sll_480_ML_int_3__91_) );
  MUX2_X2 u4_sll_480_M1_2_92 ( .A(u4_sll_480_ML_int_2__92_), .B(
        u4_sll_480_ML_int_2__88_), .S(u4_sll_480_n28), .Z(
        u4_sll_480_ML_int_3__92_) );
  MUX2_X2 u4_sll_480_M1_2_93 ( .A(u4_sll_480_ML_int_2__93_), .B(
        u4_sll_480_ML_int_2__89_), .S(u4_sll_480_n28), .Z(
        u4_sll_480_ML_int_3__93_) );
  MUX2_X2 u4_sll_480_M1_2_94 ( .A(u4_sll_480_ML_int_2__94_), .B(
        u4_sll_480_ML_int_2__90_), .S(u4_sll_480_n28), .Z(
        u4_sll_480_ML_int_3__94_) );
  MUX2_X2 u4_sll_480_M1_2_95 ( .A(u4_sll_480_ML_int_2__95_), .B(
        u4_sll_480_ML_int_2__91_), .S(u4_sll_480_n28), .Z(
        u4_sll_480_ML_int_3__95_) );
  MUX2_X2 u4_sll_480_M1_2_96 ( .A(u4_sll_480_ML_int_2__96_), .B(
        u4_sll_480_ML_int_2__92_), .S(u4_sll_480_n28), .Z(
        u4_sll_480_ML_int_3__96_) );
  MUX2_X2 u4_sll_480_M1_2_97 ( .A(u4_sll_480_ML_int_2__97_), .B(
        u4_sll_480_ML_int_2__93_), .S(u4_sll_480_n28), .Z(
        u4_sll_480_ML_int_3__97_) );
  MUX2_X2 u4_sll_480_M1_2_98 ( .A(u4_sll_480_ML_int_2__98_), .B(
        u4_sll_480_ML_int_2__94_), .S(u4_sll_480_n28), .Z(
        u4_sll_480_ML_int_3__98_) );
  MUX2_X2 u4_sll_480_M1_2_99 ( .A(u4_sll_480_ML_int_2__99_), .B(
        u4_sll_480_ML_int_2__95_), .S(u4_sll_480_n28), .Z(
        u4_sll_480_ML_int_3__99_) );
  MUX2_X2 u4_sll_480_M1_2_100 ( .A(u4_sll_480_ML_int_2__100_), .B(
        u4_sll_480_ML_int_2__96_), .S(u4_sll_480_n28), .Z(
        u4_sll_480_ML_int_3__100_) );
  MUX2_X2 u4_sll_480_M1_2_101 ( .A(u4_sll_480_ML_int_2__101_), .B(
        u4_sll_480_ML_int_2__97_), .S(u4_sll_480_n28), .Z(
        u4_sll_480_ML_int_3__101_) );
  MUX2_X2 u4_sll_480_M1_2_102 ( .A(u4_sll_480_ML_int_2__102_), .B(
        u4_sll_480_ML_int_2__98_), .S(u4_sll_480_n28), .Z(
        u4_sll_480_ML_int_3__102_) );
  MUX2_X2 u4_sll_480_M1_2_103 ( .A(u4_sll_480_ML_int_2__103_), .B(
        u4_sll_480_ML_int_2__99_), .S(u4_sll_480_n29), .Z(
        u4_sll_480_ML_int_3__103_) );
  MUX2_X2 u4_sll_480_M1_2_104 ( .A(u4_sll_480_ML_int_2__104_), .B(
        u4_sll_480_ML_int_2__100_), .S(u4_sll_480_n29), .Z(
        u4_sll_480_ML_int_3__104_) );
  MUX2_X2 u4_sll_480_M1_2_105 ( .A(u4_sll_480_ML_int_2__105_), .B(
        u4_sll_480_ML_int_2__101_), .S(u4_sll_480_n29), .Z(
        u4_sll_480_ML_int_3__105_) );
  MUX2_X2 u4_sll_480_M1_2_106 ( .A(u4_sll_480_ML_int_2__106_), .B(
        u4_sll_480_ML_int_2__102_), .S(u4_sll_480_n29), .Z(
        u4_sll_480_ML_int_3__106_) );
  MUX2_X2 u4_sll_480_M1_2_107 ( .A(u4_sll_480_ML_int_2__107_), .B(
        u4_sll_480_ML_int_2__103_), .S(u4_sll_480_n29), .Z(
        u4_sll_480_ML_int_3__107_) );
  MUX2_X2 u4_sll_480_M1_2_108 ( .A(u4_sll_480_ML_int_2__108_), .B(
        u4_sll_480_ML_int_2__104_), .S(u4_sll_480_n29), .Z(
        u4_sll_480_ML_int_3__108_) );
  MUX2_X2 u4_sll_480_M1_2_109 ( .A(u4_sll_480_ML_int_2__109_), .B(
        u4_sll_480_ML_int_2__105_), .S(u4_sll_480_n29), .Z(
        u4_sll_480_ML_int_3__109_) );
  MUX2_X2 u4_sll_480_M1_2_110 ( .A(u4_sll_480_ML_int_2__110_), .B(
        u4_sll_480_ML_int_2__106_), .S(u4_sll_480_n29), .Z(
        u4_sll_480_ML_int_3__110_) );
  MUX2_X2 u4_sll_480_M1_2_111 ( .A(u4_sll_480_ML_int_2__111_), .B(
        u4_sll_480_ML_int_2__107_), .S(u4_sll_480_n29), .Z(
        u4_sll_480_ML_int_3__111_) );
  MUX2_X2 u4_sll_480_M1_2_112 ( .A(u4_sll_480_ML_int_2__112_), .B(
        u4_sll_480_ML_int_2__108_), .S(u4_sll_480_n29), .Z(
        u4_sll_480_ML_int_3__112_) );
  MUX2_X2 u4_sll_480_M1_2_113 ( .A(u4_sll_480_ML_int_2__113_), .B(
        u4_sll_480_ML_int_2__109_), .S(u4_sll_480_n29), .Z(
        u4_sll_480_ML_int_3__113_) );
  MUX2_X2 u4_sll_480_M1_2_114 ( .A(u4_sll_480_ML_int_2__114_), .B(
        u4_sll_480_ML_int_2__110_), .S(u4_sll_480_n25), .Z(
        u4_sll_480_ML_int_3__114_) );
  MUX2_X2 u4_sll_480_M1_2_115 ( .A(u4_sll_480_n3), .B(
        u4_sll_480_ML_int_2__111_), .S(u4_sll_480_n25), .Z(
        u4_sll_480_ML_int_3__115_) );
  MUX2_X2 u4_sll_480_M1_2_116 ( .A(u4_sll_480_n4), .B(
        u4_sll_480_ML_int_2__112_), .S(u4_sll_480_n25), .Z(
        u4_sll_480_ML_int_3__116_) );
  MUX2_X2 u4_sll_480_M1_3_11 ( .A(u4_sll_480_ML_int_3__11_), .B(u4_sll_480_n41), .S(u4_sll_480_n33), .Z(u4_sll_480_ML_int_4__11_) );
  MUX2_X2 u4_sll_480_M1_3_12 ( .A(u4_sll_480_ML_int_3__12_), .B(
        u4_sll_480_ML_int_3__4_), .S(u4_sll_480_n32), .Z(
        u4_sll_480_ML_int_4__12_) );
  MUX2_X2 u4_sll_480_M1_3_13 ( .A(u4_sll_480_ML_int_3__13_), .B(
        u4_sll_480_ML_int_3__5_), .S(u4_sll_480_n32), .Z(
        u4_sll_480_ML_int_4__13_) );
  MUX2_X2 u4_sll_480_M1_3_14 ( .A(u4_sll_480_ML_int_3__14_), .B(
        u4_sll_480_ML_int_3__6_), .S(u4_sll_480_n32), .Z(
        u4_sll_480_ML_int_4__14_) );
  MUX2_X2 u4_sll_480_M1_3_15 ( .A(u4_sll_480_ML_int_3__15_), .B(
        u4_sll_480_ML_int_3__7_), .S(u4_sll_480_n32), .Z(
        u4_sll_480_ML_int_4__15_) );
  MUX2_X2 u4_sll_480_M1_3_16 ( .A(u4_sll_480_ML_int_3__16_), .B(
        u4_sll_480_ML_int_3__8_), .S(u4_sll_480_n32), .Z(
        u4_sll_480_ML_int_4__16_) );
  MUX2_X2 u4_sll_480_M1_3_17 ( .A(u4_sll_480_ML_int_3__17_), .B(
        u4_sll_480_ML_int_3__9_), .S(u4_sll_480_n32), .Z(
        u4_sll_480_ML_int_4__17_) );
  MUX2_X2 u4_sll_480_M1_3_18 ( .A(u4_sll_480_ML_int_3__18_), .B(
        u4_sll_480_ML_int_3__10_), .S(u4_sll_480_n32), .Z(
        u4_sll_480_ML_int_4__18_) );
  MUX2_X2 u4_sll_480_M1_3_19 ( .A(u4_sll_480_ML_int_3__19_), .B(
        u4_sll_480_ML_int_3__11_), .S(u4_sll_480_n32), .Z(
        u4_sll_480_ML_int_4__19_) );
  MUX2_X2 u4_sll_480_M1_3_20 ( .A(u4_sll_480_ML_int_3__20_), .B(
        u4_sll_480_ML_int_3__12_), .S(u4_sll_480_temp_int_SH_3_), .Z(
        u4_sll_480_ML_int_4__20_) );
  MUX2_X2 u4_sll_480_M1_3_21 ( .A(u4_sll_480_ML_int_3__21_), .B(
        u4_sll_480_ML_int_3__13_), .S(u4_sll_480_temp_int_SH_3_), .Z(
        u4_sll_480_ML_int_4__21_) );
  MUX2_X2 u4_sll_480_M1_3_27 ( .A(u4_sll_480_ML_int_3__27_), .B(
        u4_sll_480_ML_int_3__19_), .S(u4_sll_480_n31), .Z(
        u4_sll_480_ML_int_4__27_) );
  MUX2_X2 u4_sll_480_M1_3_28 ( .A(u4_sll_480_ML_int_3__28_), .B(
        u4_sll_480_ML_int_3__20_), .S(u4_sll_480_n31), .Z(
        u4_sll_480_ML_int_4__28_) );
  MUX2_X2 u4_sll_480_M1_3_29 ( .A(u4_sll_480_ML_int_3__29_), .B(
        u4_sll_480_ML_int_3__21_), .S(u4_sll_480_n31), .Z(
        u4_sll_480_ML_int_4__29_) );
  MUX2_X2 u4_sll_480_M1_3_30 ( .A(u4_sll_480_ML_int_3__30_), .B(
        u4_sll_480_ML_int_3__22_), .S(u4_sll_480_n31), .Z(
        u4_sll_480_ML_int_4__30_) );
  MUX2_X2 u4_sll_480_M1_3_31 ( .A(u4_sll_480_ML_int_3__31_), .B(
        u4_sll_480_ML_int_3__23_), .S(u4_sll_480_n31), .Z(
        u4_sll_480_ML_int_4__31_) );
  MUX2_X2 u4_sll_480_M1_3_32 ( .A(u4_sll_480_ML_int_3__32_), .B(
        u4_sll_480_ML_int_3__24_), .S(u4_sll_480_n31), .Z(
        u4_sll_480_ML_int_4__32_) );
  MUX2_X2 u4_sll_480_M1_3_33 ( .A(u4_sll_480_ML_int_3__33_), .B(
        u4_sll_480_ML_int_3__25_), .S(u4_sll_480_n31), .Z(
        u4_sll_480_ML_int_4__33_) );
  MUX2_X2 u4_sll_480_M1_3_34 ( .A(u4_sll_480_ML_int_3__34_), .B(
        u4_sll_480_ML_int_3__26_), .S(u4_sll_480_n31), .Z(
        u4_sll_480_ML_int_4__34_) );
  MUX2_X2 u4_sll_480_M1_3_35 ( .A(u4_sll_480_ML_int_3__35_), .B(
        u4_sll_480_ML_int_3__27_), .S(u4_sll_480_n31), .Z(
        u4_sll_480_ML_int_4__35_) );
  MUX2_X2 u4_sll_480_M1_3_36 ( .A(u4_sll_480_ML_int_3__36_), .B(
        u4_sll_480_ML_int_3__28_), .S(u4_sll_480_n31), .Z(
        u4_sll_480_ML_int_4__36_) );
  MUX2_X2 u4_sll_480_M1_3_37 ( .A(u4_sll_480_ML_int_3__37_), .B(
        u4_sll_480_ML_int_3__29_), .S(u4_sll_480_n31), .Z(
        u4_sll_480_ML_int_4__37_) );
  MUX2_X2 u4_sll_480_M1_3_43 ( .A(u4_sll_480_ML_int_3__43_), .B(
        u4_sll_480_ML_int_3__35_), .S(u4_sll_480_n32), .Z(
        u4_sll_480_ML_int_4__43_) );
  MUX2_X2 u4_sll_480_M1_3_44 ( .A(u4_sll_480_ML_int_3__44_), .B(
        u4_sll_480_ML_int_3__36_), .S(u4_sll_480_n32), .Z(
        u4_sll_480_ML_int_4__44_) );
  MUX2_X2 u4_sll_480_M1_3_45 ( .A(u4_sll_480_ML_int_3__45_), .B(
        u4_sll_480_ML_int_3__37_), .S(u4_sll_480_n32), .Z(
        u4_sll_480_ML_int_4__45_) );
  MUX2_X2 u4_sll_480_M1_3_46 ( .A(u4_sll_480_ML_int_3__46_), .B(
        u4_sll_480_ML_int_3__38_), .S(u4_sll_480_n30), .Z(
        u4_sll_480_ML_int_4__46_) );
  MUX2_X2 u4_sll_480_M1_3_47 ( .A(u4_sll_480_ML_int_3__47_), .B(
        u4_sll_480_ML_int_3__39_), .S(u4_sll_480_n33), .Z(
        u4_sll_480_ML_int_4__47_) );
  MUX2_X2 u4_sll_480_M1_3_48 ( .A(u4_sll_480_ML_int_3__48_), .B(
        u4_sll_480_ML_int_3__40_), .S(u4_sll_480_n32), .Z(
        u4_sll_480_ML_int_4__48_) );
  MUX2_X2 u4_sll_480_M1_3_49 ( .A(u4_sll_480_ML_int_3__49_), .B(
        u4_sll_480_ML_int_3__41_), .S(u4_sll_480_n30), .Z(
        u4_sll_480_ML_int_4__49_) );
  MUX2_X2 u4_sll_480_M1_3_50 ( .A(u4_sll_480_ML_int_3__50_), .B(
        u4_sll_480_ML_int_3__42_), .S(u4_sll_480_n31), .Z(
        u4_sll_480_ML_int_4__50_) );
  MUX2_X2 u4_sll_480_M1_3_51 ( .A(u4_sll_480_ML_int_3__51_), .B(
        u4_sll_480_ML_int_3__43_), .S(u4_sll_480_n32), .Z(
        u4_sll_480_ML_int_4__51_) );
  MUX2_X2 u4_sll_480_M1_3_52 ( .A(u4_sll_480_ML_int_3__52_), .B(
        u4_sll_480_ML_int_3__44_), .S(u4_sll_480_temp_int_SH_3_), .Z(
        u4_sll_480_ML_int_4__52_) );
  MUX2_X2 u4_sll_480_M1_3_53 ( .A(u4_sll_480_ML_int_3__53_), .B(
        u4_sll_480_ML_int_3__45_), .S(u4_sll_480_temp_int_SH_3_), .Z(
        u4_sll_480_ML_int_4__53_) );
  MUX2_X2 u4_sll_480_M1_3_59 ( .A(u4_sll_480_ML_int_3__59_), .B(
        u4_sll_480_ML_int_3__51_), .S(u4_sll_480_n33), .Z(
        u4_sll_480_ML_int_4__59_) );
  MUX2_X2 u4_sll_480_M1_3_60 ( .A(u4_sll_480_ML_int_3__60_), .B(
        u4_sll_480_ML_int_3__52_), .S(u4_sll_480_n31), .Z(
        u4_sll_480_ML_int_4__60_) );
  MUX2_X2 u4_sll_480_M1_3_61 ( .A(u4_sll_480_ML_int_3__61_), .B(
        u4_sll_480_ML_int_3__53_), .S(u4_sll_480_n32), .Z(
        u4_sll_480_ML_int_4__61_) );
  MUX2_X2 u4_sll_480_M1_3_62 ( .A(u4_sll_480_ML_int_3__62_), .B(
        u4_sll_480_ML_int_3__54_), .S(u4_sll_480_n32), .Z(
        u4_sll_480_ML_int_4__62_) );
  MUX2_X2 u4_sll_480_M1_3_63 ( .A(u4_sll_480_ML_int_3__63_), .B(
        u4_sll_480_ML_int_3__55_), .S(u4_sll_480_n32), .Z(
        u4_sll_480_ML_int_4__63_) );
  MUX2_X2 u4_sll_480_M1_3_64 ( .A(u4_sll_480_ML_int_3__64_), .B(
        u4_sll_480_ML_int_3__56_), .S(u4_sll_480_n32), .Z(
        u4_sll_480_ML_int_4__64_) );
  MUX2_X2 u4_sll_480_M1_3_65 ( .A(u4_sll_480_ML_int_3__65_), .B(
        u4_sll_480_ML_int_3__57_), .S(u4_sll_480_n32), .Z(
        u4_sll_480_ML_int_4__65_) );
  MUX2_X2 u4_sll_480_M1_3_66 ( .A(u4_sll_480_ML_int_3__66_), .B(
        u4_sll_480_ML_int_3__58_), .S(u4_sll_480_n32), .Z(
        u4_sll_480_ML_int_4__66_) );
  MUX2_X2 u4_sll_480_M1_3_67 ( .A(u4_sll_480_ML_int_3__67_), .B(
        u4_sll_480_ML_int_3__59_), .S(u4_sll_480_n32), .Z(
        u4_sll_480_ML_int_4__67_) );
  MUX2_X2 u4_sll_480_M1_3_68 ( .A(u4_sll_480_ML_int_3__68_), .B(
        u4_sll_480_ML_int_3__60_), .S(u4_sll_480_temp_int_SH_3_), .Z(
        u4_sll_480_ML_int_4__68_) );
  MUX2_X2 u4_sll_480_M1_3_69 ( .A(u4_sll_480_ML_int_3__69_), .B(
        u4_sll_480_ML_int_3__61_), .S(u4_sll_480_temp_int_SH_3_), .Z(
        u4_sll_480_ML_int_4__69_) );
  MUX2_X2 u4_sll_480_M1_3_75 ( .A(u4_sll_480_ML_int_3__75_), .B(
        u4_sll_480_ML_int_3__67_), .S(u4_sll_480_n30), .Z(
        u4_sll_480_ML_int_4__75_) );
  MUX2_X2 u4_sll_480_M1_3_76 ( .A(u4_sll_480_ML_int_3__76_), .B(
        u4_sll_480_ML_int_3__68_), .S(u4_sll_480_n32), .Z(
        u4_sll_480_ML_int_4__76_) );
  MUX2_X2 u4_sll_480_M1_3_77 ( .A(u4_sll_480_ML_int_3__77_), .B(
        u4_sll_480_ML_int_3__69_), .S(u4_sll_480_n31), .Z(
        u4_sll_480_ML_int_4__77_) );
  MUX2_X2 u4_sll_480_M1_3_78 ( .A(u4_sll_480_ML_int_3__78_), .B(
        u4_sll_480_ML_int_3__70_), .S(u4_sll_480_n30), .Z(
        u4_sll_480_ML_int_4__78_) );
  MUX2_X2 u4_sll_480_M1_3_79 ( .A(u4_sll_480_ML_int_3__79_), .B(
        u4_sll_480_ML_int_3__71_), .S(u4_sll_480_n31), .Z(
        u4_sll_480_ML_int_4__79_) );
  MUX2_X2 u4_sll_480_M1_3_80 ( .A(u4_sll_480_ML_int_3__80_), .B(
        u4_sll_480_ML_int_3__72_), .S(u4_sll_480_n30), .Z(
        u4_sll_480_ML_int_4__80_) );
  MUX2_X2 u4_sll_480_M1_3_81 ( .A(u4_sll_480_ML_int_3__81_), .B(
        u4_sll_480_ML_int_3__73_), .S(u4_sll_480_n32), .Z(
        u4_sll_480_ML_int_4__81_) );
  MUX2_X2 u4_sll_480_M1_3_82 ( .A(u4_sll_480_ML_int_3__82_), .B(
        u4_sll_480_ML_int_3__74_), .S(u4_sll_480_n33), .Z(
        u4_sll_480_ML_int_4__82_) );
  MUX2_X2 u4_sll_480_M1_3_83 ( .A(u4_sll_480_ML_int_3__83_), .B(
        u4_sll_480_ML_int_3__75_), .S(u4_sll_480_n31), .Z(
        u4_sll_480_ML_int_4__83_) );
  MUX2_X2 u4_sll_480_M1_3_84 ( .A(u4_sll_480_ML_int_3__84_), .B(
        u4_sll_480_ML_int_3__76_), .S(u4_sll_480_n31), .Z(
        u4_sll_480_ML_int_4__84_) );
  MUX2_X2 u4_sll_480_M1_3_85 ( .A(u4_sll_480_ML_int_3__85_), .B(
        u4_sll_480_ML_int_3__77_), .S(u4_sll_480_n30), .Z(
        u4_sll_480_ML_int_4__85_) );
  MUX2_X2 u4_sll_480_M1_3_91 ( .A(u4_sll_480_ML_int_3__91_), .B(
        u4_sll_480_ML_int_3__83_), .S(u4_sll_480_n33), .Z(
        u4_sll_480_ML_int_4__91_) );
  MUX2_X2 u4_sll_480_M1_3_92 ( .A(u4_sll_480_ML_int_3__92_), .B(
        u4_sll_480_ML_int_3__84_), .S(u4_sll_480_n33), .Z(
        u4_sll_480_ML_int_4__92_) );
  MUX2_X2 u4_sll_480_M1_3_93 ( .A(u4_sll_480_ML_int_3__93_), .B(
        u4_sll_480_ML_int_3__85_), .S(u4_sll_480_n33), .Z(
        u4_sll_480_ML_int_4__93_) );
  MUX2_X2 u4_sll_480_M1_3_94 ( .A(u4_sll_480_ML_int_3__94_), .B(
        u4_sll_480_ML_int_3__86_), .S(u4_sll_480_n33), .Z(
        u4_sll_480_ML_int_4__94_) );
  MUX2_X2 u4_sll_480_M1_3_95 ( .A(u4_sll_480_ML_int_3__95_), .B(
        u4_sll_480_ML_int_3__87_), .S(u4_sll_480_n33), .Z(
        u4_sll_480_ML_int_4__95_) );
  MUX2_X2 u4_sll_480_M1_3_96 ( .A(u4_sll_480_ML_int_3__96_), .B(
        u4_sll_480_ML_int_3__88_), .S(u4_sll_480_n33), .Z(
        u4_sll_480_ML_int_4__96_) );
  MUX2_X2 u4_sll_480_M1_3_97 ( .A(u4_sll_480_ML_int_3__97_), .B(
        u4_sll_480_ML_int_3__89_), .S(u4_sll_480_n33), .Z(
        u4_sll_480_ML_int_4__97_) );
  MUX2_X2 u4_sll_480_M1_3_98 ( .A(u4_sll_480_ML_int_3__98_), .B(
        u4_sll_480_ML_int_3__90_), .S(u4_sll_480_n33), .Z(
        u4_sll_480_ML_int_4__98_) );
  MUX2_X2 u4_sll_480_M1_3_99 ( .A(u4_sll_480_ML_int_3__99_), .B(
        u4_sll_480_ML_int_3__91_), .S(u4_sll_480_n33), .Z(
        u4_sll_480_ML_int_4__99_) );
  MUX2_X2 u4_sll_480_M1_3_100 ( .A(u4_sll_480_ML_int_3__100_), .B(
        u4_sll_480_ML_int_3__92_), .S(u4_sll_480_n33), .Z(
        u4_sll_480_ML_int_4__100_) );
  MUX2_X2 u4_sll_480_M1_3_101 ( .A(u4_sll_480_ML_int_3__101_), .B(
        u4_sll_480_ML_int_3__93_), .S(u4_sll_480_n33), .Z(
        u4_sll_480_ML_int_4__101_) );
  MUX2_X2 u4_sll_480_M1_3_107 ( .A(u4_sll_480_ML_int_3__107_), .B(
        u4_sll_480_ML_int_3__99_), .S(u4_sll_480_n30), .Z(
        u4_sll_480_ML_int_4__107_) );
  MUX2_X2 u4_sll_480_M1_3_108 ( .A(u4_sll_480_ML_int_3__108_), .B(
        u4_sll_480_ML_int_3__100_), .S(u4_sll_480_n30), .Z(
        u4_sll_480_ML_int_4__108_) );
  MUX2_X2 u4_sll_480_M1_3_109 ( .A(u4_sll_480_ML_int_3__109_), .B(
        u4_sll_480_ML_int_3__101_), .S(u4_sll_480_n30), .Z(
        u4_sll_480_ML_int_4__109_) );
  MUX2_X2 u4_sll_480_M1_3_110 ( .A(u4_sll_480_ML_int_3__110_), .B(
        u4_sll_480_ML_int_3__102_), .S(u4_sll_480_n30), .Z(
        u4_sll_480_ML_int_4__110_) );
  MUX2_X2 u4_sll_480_M1_3_111 ( .A(u4_sll_480_ML_int_3__111_), .B(
        u4_sll_480_ML_int_3__103_), .S(u4_sll_480_n30), .Z(
        u4_sll_480_ML_int_4__111_) );
  MUX2_X2 u4_sll_480_M1_3_112 ( .A(u4_sll_480_ML_int_3__112_), .B(
        u4_sll_480_ML_int_3__104_), .S(u4_sll_480_n30), .Z(
        u4_sll_480_ML_int_4__112_) );
  MUX2_X2 u4_sll_480_M1_3_113 ( .A(u4_sll_480_ML_int_3__113_), .B(
        u4_sll_480_ML_int_3__105_), .S(u4_sll_480_n30), .Z(
        u4_sll_480_ML_int_4__113_) );
  MUX2_X2 u4_sll_480_M1_3_114 ( .A(u4_sll_480_ML_int_3__114_), .B(
        u4_sll_480_ML_int_3__106_), .S(u4_sll_480_n30), .Z(
        u4_sll_480_ML_int_4__114_) );
  MUX2_X2 u4_sll_480_M1_3_115 ( .A(u4_sll_480_ML_int_3__115_), .B(
        u4_sll_480_ML_int_3__107_), .S(u4_sll_480_n30), .Z(
        u4_sll_480_ML_int_4__115_) );
  MUX2_X2 u4_sll_480_M1_3_116 ( .A(u4_sll_480_ML_int_3__116_), .B(
        u4_sll_480_ML_int_3__108_), .S(u4_sll_480_n30), .Z(
        u4_sll_480_ML_int_4__116_) );
  MUX2_X2 u4_sll_480_M1_3_117 ( .A(u4_sll_480_n5), .B(
        u4_sll_480_ML_int_3__109_), .S(u4_sll_480_n30), .Z(
        u4_sll_480_ML_int_4__117_) );
  MUX2_X2 u4_sll_480_M1_4_16 ( .A(u4_sll_480_ML_int_4__16_), .B(
        u4_sll_480_ML_int_4__0_), .S(u4_sll_480_temp_int_SH_4_), .Z(
        u4_sll_480_ML_int_5__16_) );
  MUX2_X2 u4_sll_480_M1_4_17 ( .A(u4_sll_480_ML_int_4__17_), .B(
        u4_sll_480_ML_int_4__1_), .S(u4_sll_480_temp_int_SH_4_), .Z(
        u4_sll_480_ML_int_5__17_) );
  MUX2_X2 u4_sll_480_M1_4_18 ( .A(u4_sll_480_ML_int_4__18_), .B(
        u4_sll_480_ML_int_4__2_), .S(u4_sll_480_n37), .Z(
        u4_sll_480_ML_int_5__18_) );
  MUX2_X2 u4_sll_480_M1_4_19 ( .A(u4_sll_480_ML_int_4__19_), .B(
        u4_sll_480_ML_int_4__3_), .S(u4_sll_480_n36), .Z(
        u4_sll_480_ML_int_5__19_) );
  MUX2_X2 u4_sll_480_M1_4_20 ( .A(u4_sll_480_ML_int_4__20_), .B(
        u4_sll_480_ML_int_4__4_), .S(u4_sll_480_temp_int_SH_4_), .Z(
        u4_sll_480_ML_int_5__20_) );
  MUX2_X2 u4_sll_480_M1_4_21 ( .A(u4_sll_480_ML_int_4__21_), .B(
        u4_sll_480_ML_int_4__5_), .S(u4_sll_480_temp_int_SH_4_), .Z(
        u4_sll_480_ML_int_5__21_) );
  MUX2_X2 u4_sll_480_M1_4_43 ( .A(u4_sll_480_ML_int_4__43_), .B(
        u4_sll_480_ML_int_4__27_), .S(u4_sll_480_temp_int_SH_4_), .Z(
        u4_sll_480_ML_int_5__43_) );
  MUX2_X2 u4_sll_480_M1_4_44 ( .A(u4_sll_480_ML_int_4__44_), .B(
        u4_sll_480_ML_int_4__28_), .S(u4_sll_480_n36), .Z(
        u4_sll_480_ML_int_5__44_) );
  MUX2_X2 u4_sll_480_M1_4_45 ( .A(u4_sll_480_ML_int_4__45_), .B(
        u4_sll_480_ML_int_4__29_), .S(u4_sll_480_temp_int_SH_4_), .Z(
        u4_sll_480_ML_int_5__45_) );
  MUX2_X2 u4_sll_480_M1_4_46 ( .A(u4_sll_480_ML_int_4__46_), .B(
        u4_sll_480_ML_int_4__30_), .S(u4_sll_480_n36), .Z(
        u4_sll_480_ML_int_5__46_) );
  MUX2_X2 u4_sll_480_M1_4_47 ( .A(u4_sll_480_ML_int_4__47_), .B(
        u4_sll_480_ML_int_4__31_), .S(u4_sll_480_temp_int_SH_4_), .Z(
        u4_sll_480_ML_int_5__47_) );
  MUX2_X2 u4_sll_480_M1_4_48 ( .A(u4_sll_480_ML_int_4__48_), .B(
        u4_sll_480_ML_int_4__32_), .S(u4_sll_480_n36), .Z(
        u4_sll_480_ML_int_5__48_) );
  MUX2_X2 u4_sll_480_M1_4_49 ( .A(u4_sll_480_ML_int_4__49_), .B(
        u4_sll_480_ML_int_4__33_), .S(u4_sll_480_n36), .Z(
        u4_sll_480_ML_int_5__49_) );
  MUX2_X2 u4_sll_480_M1_4_50 ( .A(u4_sll_480_ML_int_4__50_), .B(
        u4_sll_480_ML_int_4__34_), .S(u4_sll_480_n36), .Z(
        u4_sll_480_ML_int_5__50_) );
  MUX2_X2 u4_sll_480_M1_4_51 ( .A(u4_sll_480_ML_int_4__51_), .B(
        u4_sll_480_ML_int_4__35_), .S(u4_sll_480_n36), .Z(
        u4_sll_480_ML_int_5__51_) );
  MUX2_X2 u4_sll_480_M1_4_52 ( .A(u4_sll_480_ML_int_4__52_), .B(
        u4_sll_480_ML_int_4__36_), .S(u4_sll_480_n36), .Z(
        u4_sll_480_ML_int_5__52_) );
  MUX2_X2 u4_sll_480_M1_4_53 ( .A(u4_sll_480_ML_int_4__53_), .B(
        u4_sll_480_ML_int_4__37_), .S(u4_sll_480_n36), .Z(
        u4_sll_480_ML_int_5__53_) );
  MUX2_X2 u4_sll_480_M1_4_75 ( .A(u4_sll_480_ML_int_4__75_), .B(
        u4_sll_480_ML_int_4__59_), .S(u4_sll_480_n36), .Z(
        u4_sll_480_ML_int_5__75_) );
  MUX2_X2 u4_sll_480_M1_4_76 ( .A(u4_sll_480_ML_int_4__76_), .B(
        u4_sll_480_ML_int_4__60_), .S(u4_sll_480_n36), .Z(
        u4_sll_480_ML_int_5__76_) );
  MUX2_X2 u4_sll_480_M1_4_77 ( .A(u4_sll_480_ML_int_4__77_), .B(
        u4_sll_480_ML_int_4__61_), .S(u4_sll_480_n36), .Z(
        u4_sll_480_ML_int_5__77_) );
  MUX2_X2 u4_sll_480_M1_4_78 ( .A(u4_sll_480_ML_int_4__78_), .B(
        u4_sll_480_ML_int_4__62_), .S(u4_sll_480_n36), .Z(
        u4_sll_480_ML_int_5__78_) );
  MUX2_X2 u4_sll_480_M1_4_79 ( .A(u4_sll_480_ML_int_4__79_), .B(
        u4_sll_480_ML_int_4__63_), .S(u4_sll_480_n36), .Z(
        u4_sll_480_ML_int_5__79_) );
  MUX2_X2 u4_sll_480_M1_4_80 ( .A(u4_sll_480_ML_int_4__80_), .B(
        u4_sll_480_ML_int_4__64_), .S(u4_sll_480_n37), .Z(
        u4_sll_480_ML_int_5__80_) );
  MUX2_X2 u4_sll_480_M1_4_81 ( .A(u4_sll_480_ML_int_4__81_), .B(
        u4_sll_480_ML_int_4__65_), .S(u4_sll_480_n37), .Z(
        u4_sll_480_ML_int_5__81_) );
  MUX2_X2 u4_sll_480_M1_4_82 ( .A(u4_sll_480_ML_int_4__82_), .B(
        u4_sll_480_ML_int_4__66_), .S(u4_sll_480_n37), .Z(
        u4_sll_480_ML_int_5__82_) );
  MUX2_X2 u4_sll_480_M1_4_83 ( .A(u4_sll_480_ML_int_4__83_), .B(
        u4_sll_480_ML_int_4__67_), .S(u4_sll_480_n37), .Z(
        u4_sll_480_ML_int_5__83_) );
  MUX2_X2 u4_sll_480_M1_4_84 ( .A(u4_sll_480_ML_int_4__84_), .B(
        u4_sll_480_ML_int_4__68_), .S(u4_sll_480_n37), .Z(
        u4_sll_480_ML_int_5__84_) );
  MUX2_X2 u4_sll_480_M1_4_85 ( .A(u4_sll_480_ML_int_4__85_), .B(
        u4_sll_480_ML_int_4__69_), .S(u4_sll_480_n37), .Z(
        u4_sll_480_ML_int_5__85_) );
  MUX2_X2 u4_sll_480_M1_4_107 ( .A(u4_sll_480_ML_int_4__107_), .B(
        u4_sll_480_ML_int_4__91_), .S(u4_sll_480_n37), .Z(
        u4_sll_480_ML_int_5__107_) );
  MUX2_X2 u4_sll_480_M1_4_108 ( .A(u4_sll_480_ML_int_4__108_), .B(
        u4_sll_480_ML_int_4__92_), .S(u4_sll_480_n37), .Z(
        u4_sll_480_ML_int_5__108_) );
  MUX2_X2 u4_sll_480_M1_4_109 ( .A(u4_sll_480_ML_int_4__109_), .B(
        u4_sll_480_ML_int_4__93_), .S(u4_sll_480_n37), .Z(
        u4_sll_480_ML_int_5__109_) );
  MUX2_X2 u4_sll_480_M1_4_110 ( .A(u4_sll_480_ML_int_4__110_), .B(
        u4_sll_480_ML_int_4__94_), .S(u4_sll_480_n37), .Z(
        u4_sll_480_ML_int_5__110_) );
  MUX2_X2 u4_sll_480_M1_4_111 ( .A(u4_sll_480_ML_int_4__111_), .B(
        u4_sll_480_ML_int_4__95_), .S(u4_sll_480_n37), .Z(
        u4_sll_480_ML_int_5__111_) );
  MUX2_X2 u4_sll_480_M1_4_112 ( .A(u4_sll_480_ML_int_4__112_), .B(
        u4_sll_480_ML_int_4__96_), .S(u4_sll_480_n36), .Z(
        u4_sll_480_ML_int_5__112_) );
  MUX2_X2 u4_sll_480_M1_4_113 ( .A(u4_sll_480_ML_int_4__113_), .B(
        u4_sll_480_ML_int_4__97_), .S(u4_sll_480_n37), .Z(
        u4_sll_480_ML_int_5__113_) );
  MUX2_X2 u4_sll_480_M1_4_114 ( .A(u4_sll_480_ML_int_4__114_), .B(
        u4_sll_480_ML_int_4__98_), .S(u4_sll_480_n36), .Z(
        u4_sll_480_ML_int_5__114_) );
  MUX2_X2 u4_sll_480_M1_4_115 ( .A(u4_sll_480_ML_int_4__115_), .B(
        u4_sll_480_ML_int_4__99_), .S(u4_sll_480_n37), .Z(
        u4_sll_480_ML_int_5__115_) );
  MUX2_X2 u4_sll_480_M1_4_116 ( .A(u4_sll_480_ML_int_4__116_), .B(
        u4_sll_480_ML_int_4__100_), .S(u4_sll_480_n36), .Z(
        u4_sll_480_ML_int_5__116_) );
  MUX2_X2 u4_sll_480_M1_4_117 ( .A(u4_sll_480_ML_int_4__117_), .B(
        u4_sll_480_ML_int_4__101_), .S(u4_sll_480_n37), .Z(
        u4_sll_480_ML_int_5__117_) );
  MUX2_X2 u4_sll_480_M1_5_43 ( .A(u4_sll_480_ML_int_5__43_), .B(
        u4_sll_480_ML_int_5__11_), .S(u4_sll_480_n42), .Z(
        u4_sll_480_ML_int_6__43_) );
  MUX2_X2 u4_sll_480_M1_5_44 ( .A(u4_sll_480_ML_int_5__44_), .B(
        u4_sll_480_ML_int_5__12_), .S(u4_sll_480_n42), .Z(
        u4_sll_480_ML_int_6__44_) );
  MUX2_X2 u4_sll_480_M1_5_45 ( .A(u4_sll_480_ML_int_5__45_), .B(
        u4_sll_480_ML_int_5__13_), .S(u4_sll_480_n42), .Z(
        u4_sll_480_ML_int_6__45_) );
  MUX2_X2 u4_sll_480_M1_5_46 ( .A(u4_sll_480_ML_int_5__46_), .B(
        u4_sll_480_ML_int_5__14_), .S(u4_sll_480_n42), .Z(
        u4_sll_480_ML_int_6__46_) );
  MUX2_X2 u4_sll_480_M1_5_47 ( .A(u4_sll_480_ML_int_5__47_), .B(
        u4_sll_480_ML_int_5__15_), .S(u4_sll_480_n42), .Z(
        u4_sll_480_ML_int_6__47_) );
  MUX2_X2 u4_sll_480_M1_5_48 ( .A(u4_sll_480_ML_int_5__48_), .B(
        u4_sll_480_ML_int_5__16_), .S(u4_sll_480_n42), .Z(
        u4_sll_480_ML_int_6__48_) );
  MUX2_X2 u4_sll_480_M1_5_49 ( .A(u4_sll_480_ML_int_5__49_), .B(
        u4_sll_480_ML_int_5__17_), .S(u4_sll_480_n42), .Z(
        u4_sll_480_ML_int_6__49_) );
  MUX2_X2 u4_sll_480_M1_5_50 ( .A(u4_sll_480_ML_int_5__50_), .B(
        u4_sll_480_ML_int_5__18_), .S(u4_sll_480_n42), .Z(
        u4_sll_480_ML_int_6__50_) );
  MUX2_X2 u4_sll_480_M1_5_51 ( .A(u4_sll_480_ML_int_5__51_), .B(
        u4_sll_480_ML_int_5__19_), .S(u4_sll_480_n42), .Z(
        u4_sll_480_ML_int_6__51_) );
  MUX2_X2 u4_sll_480_M1_5_52 ( .A(u4_sll_480_ML_int_5__52_), .B(
        u4_sll_480_ML_int_5__20_), .S(u4_sll_480_n42), .Z(
        u4_sll_480_ML_int_6__52_) );
  MUX2_X2 u4_sll_480_M1_5_53 ( .A(u4_sll_480_ML_int_5__53_), .B(
        u4_sll_480_ML_int_5__21_), .S(u4_sll_480_n42), .Z(
        u4_sll_480_ML_int_6__53_) );
  MUX2_X2 u4_sll_480_M1_5_107 ( .A(u4_sll_480_ML_int_5__107_), .B(
        u4_sll_480_ML_int_5__75_), .S(u4_sll_480_n42), .Z(
        u4_sll_480_ML_int_6__107_) );
  MUX2_X2 u4_sll_480_M1_5_108 ( .A(u4_sll_480_ML_int_5__108_), .B(
        u4_sll_480_ML_int_5__76_), .S(u4_sll_480_n42), .Z(
        u4_sll_480_ML_int_6__108_) );
  MUX2_X2 u4_sll_480_M1_5_109 ( .A(u4_sll_480_ML_int_5__109_), .B(
        u4_sll_480_ML_int_5__77_), .S(u4_sll_480_n42), .Z(
        u4_sll_480_ML_int_6__109_) );
  MUX2_X2 u4_sll_480_M1_5_110 ( .A(u4_sll_480_ML_int_5__110_), .B(
        u4_sll_480_ML_int_5__78_), .S(u4_sll_480_n42), .Z(
        u4_sll_480_ML_int_6__110_) );
  MUX2_X2 u4_sll_480_M1_5_111 ( .A(u4_sll_480_ML_int_5__111_), .B(
        u4_sll_480_ML_int_5__79_), .S(u4_sll_480_n42), .Z(
        u4_sll_480_ML_int_6__111_) );
  MUX2_X2 u4_sll_480_M1_5_112 ( .A(u4_sll_480_ML_int_5__112_), .B(
        u4_sll_480_ML_int_5__80_), .S(u4_sll_480_n42), .Z(
        u4_sll_480_ML_int_6__112_) );
  MUX2_X2 u4_sll_480_M1_5_113 ( .A(u4_sll_480_ML_int_5__113_), .B(
        u4_sll_480_ML_int_5__81_), .S(u4_sll_480_n42), .Z(
        u4_sll_480_ML_int_6__113_) );
  MUX2_X2 u4_sll_480_M1_5_114 ( .A(u4_sll_480_ML_int_5__114_), .B(
        u4_sll_480_ML_int_5__82_), .S(u4_sll_480_n42), .Z(
        u4_sll_480_ML_int_6__114_) );
  MUX2_X2 u4_sll_480_M1_5_115 ( .A(u4_sll_480_ML_int_5__115_), .B(
        u4_sll_480_ML_int_5__83_), .S(u4_sll_480_n42), .Z(
        u4_sll_480_ML_int_6__115_) );
  MUX2_X2 u4_sll_480_M1_5_116 ( .A(u4_sll_480_ML_int_5__116_), .B(
        u4_sll_480_ML_int_5__84_), .S(u4_sll_480_n42), .Z(
        u4_sll_480_ML_int_6__116_) );
  MUX2_X2 u4_sll_480_M1_5_117 ( .A(u4_sll_480_ML_int_5__117_), .B(
        u4_sll_480_ML_int_5__85_), .S(u4_sll_480_n42), .Z(
        u4_sll_480_ML_int_6__117_) );
  MUX2_X2 u4_sll_480_M1_6_107 ( .A(u4_sll_480_ML_int_6__107_), .B(
        u4_sll_480_ML_int_6__43_), .S(u4_sll_480_n43), .Z(
        u4_sll_480_ML_int_7__107_) );
  MUX2_X2 u4_sll_480_M1_6_108 ( .A(u4_sll_480_ML_int_6__108_), .B(
        u4_sll_480_ML_int_6__44_), .S(u4_sll_480_n43), .Z(
        u4_sll_480_ML_int_7__108_) );
  MUX2_X2 u4_sll_480_M1_6_109 ( .A(u4_sll_480_ML_int_6__109_), .B(
        u4_sll_480_ML_int_6__45_), .S(u4_sll_480_n43), .Z(
        u4_sll_480_ML_int_7__109_) );
  MUX2_X2 u4_sll_480_M1_6_110 ( .A(u4_sll_480_ML_int_6__110_), .B(
        u4_sll_480_ML_int_6__46_), .S(u4_sll_480_n43), .Z(
        u4_sll_480_ML_int_7__110_) );
  MUX2_X2 u4_sll_480_M1_6_111 ( .A(u4_sll_480_ML_int_6__111_), .B(
        u4_sll_480_ML_int_6__47_), .S(u4_sll_480_n43), .Z(
        u4_sll_480_ML_int_7__111_) );
  MUX2_X2 u4_sll_480_M1_6_112 ( .A(u4_sll_480_ML_int_6__112_), .B(
        u4_sll_480_ML_int_6__48_), .S(u4_sll_480_n43), .Z(
        u4_sll_480_ML_int_7__112_) );
  MUX2_X2 u4_sll_480_M1_6_113 ( .A(u4_sll_480_ML_int_6__113_), .B(
        u4_sll_480_ML_int_6__49_), .S(u4_sll_480_n43), .Z(
        u4_sll_480_ML_int_7__113_) );
  MUX2_X2 u4_sll_480_M1_6_114 ( .A(u4_sll_480_ML_int_6__114_), .B(
        u4_sll_480_ML_int_6__50_), .S(u4_sll_480_n43), .Z(
        u4_sll_480_ML_int_7__114_) );
  MUX2_X2 u4_sll_480_M1_6_115 ( .A(u4_sll_480_ML_int_6__115_), .B(
        u4_sll_480_ML_int_6__51_), .S(u4_sll_480_n43), .Z(
        u4_sll_480_ML_int_7__115_) );
  MUX2_X2 u4_sll_480_M1_6_116 ( .A(u4_sll_480_ML_int_6__116_), .B(
        u4_sll_480_ML_int_6__52_), .S(u4_sll_480_n43), .Z(
        u4_sll_480_ML_int_7__116_) );
  MUX2_X2 u4_sll_480_M1_6_117 ( .A(u4_sll_480_ML_int_6__117_), .B(
        u4_sll_480_ML_int_6__53_), .S(u4_sll_480_n43), .Z(
        u4_sll_480_ML_int_7__117_) );
  INV_X4 u4_sub_468_U27 ( .A(u4_fi_ldz_mi1_0_), .ZN(u4_sub_468_n16) );
  INV_X4 u4_sub_468_U26 ( .A(u4_fi_ldz_mi1_6_), .ZN(u4_sub_468_n15) );
  INV_X4 u4_sub_468_U25 ( .A(u4_fi_ldz_mi1_5_), .ZN(u4_sub_468_n14) );
  INV_X4 u4_sub_468_U24 ( .A(u4_fi_ldz_mi1_4_), .ZN(u4_sub_468_n13) );
  INV_X4 u4_sub_468_U23 ( .A(u4_fi_ldz_mi1_3_), .ZN(u4_sub_468_n12) );
  INV_X4 u4_sub_468_U22 ( .A(u4_fi_ldz_mi1_2_), .ZN(u4_sub_468_n11) );
  INV_X4 u4_sub_468_U21 ( .A(u4_fi_ldz_mi1_1_), .ZN(u4_sub_468_n10) );
  INV_X4 u4_sub_468_U20 ( .A(u4_exp_in_pl1_0_), .ZN(u4_sub_468_n9) );
  XNOR2_X2 u4_sub_468_U19 ( .A(u4_sub_468_n16), .B(u4_exp_in_pl1_0_), .ZN(
        u4_exp_next_mi_0_) );
  NAND2_X2 u4_sub_468_U18 ( .A1(u4_fi_ldz_mi1_0_), .A2(u4_sub_468_n9), .ZN(
        u4_sub_468_carry_1_) );
  INV_X4 u4_sub_468_U17 ( .A(u4_sub_468_carry_9_), .ZN(u4_sub_468_n8) );
  INV_X4 u4_sub_468_U16 ( .A(u4_exp_in_pl1_9_), .ZN(u4_sub_468_n7) );
  XNOR2_X2 u4_sub_468_U15 ( .A(u4_exp_in_pl1_9_), .B(u4_sub_468_carry_9_), 
        .ZN(u4_exp_next_mi_9_) );
  NAND2_X2 u4_sub_468_U14 ( .A1(u4_sub_468_n7), .A2(u4_sub_468_n8), .ZN(
        u4_sub_468_carry_10_) );
  INV_X4 u4_sub_468_U13 ( .A(u4_sub_468_carry_8_), .ZN(u4_sub_468_n6) );
  INV_X4 u4_sub_468_U12 ( .A(u4_exp_in_pl1_8_), .ZN(u4_sub_468_n5) );
  XNOR2_X2 u4_sub_468_U11 ( .A(u4_exp_in_pl1_8_), .B(u4_sub_468_carry_8_), 
        .ZN(u4_exp_next_mi_8_) );
  NAND2_X2 u4_sub_468_U10 ( .A1(u4_sub_468_n5), .A2(u4_sub_468_n6), .ZN(
        u4_sub_468_carry_9_) );
  INV_X4 u4_sub_468_U9 ( .A(u4_sub_468_carry_7_), .ZN(u4_sub_468_n4) );
  INV_X4 u4_sub_468_U8 ( .A(u4_exp_in_pl1_7_), .ZN(u4_sub_468_n3) );
  XNOR2_X2 u4_sub_468_U7 ( .A(u4_exp_in_pl1_7_), .B(u4_sub_468_carry_7_), .ZN(
        u4_exp_next_mi_7_) );
  NAND2_X2 u4_sub_468_U6 ( .A1(u4_sub_468_n3), .A2(u4_sub_468_n4), .ZN(
        u4_sub_468_carry_8_) );
  XNOR2_X2 u4_sub_468_U5 ( .A(u4_exp_in_pl1_11_), .B(u4_sub_468_carry_11_), 
        .ZN(u4_exp_next_mi_11_) );
  INV_X4 u4_sub_468_U4 ( .A(u4_sub_468_carry_10_), .ZN(u4_sub_468_n2) );
  INV_X4 u4_sub_468_U3 ( .A(u4_exp_in_pl1_10_), .ZN(u4_sub_468_n1) );
  XNOR2_X2 u4_sub_468_U2 ( .A(u4_exp_in_pl1_10_), .B(u4_sub_468_carry_10_), 
        .ZN(u4_exp_next_mi_10_) );
  NAND2_X2 u4_sub_468_U1 ( .A1(u4_sub_468_n1), .A2(u4_sub_468_n2), .ZN(
        u4_sub_468_carry_11_) );
  FA_X1 u4_sub_468_U2_1 ( .A(u4_exp_in_pl1_1_), .B(u4_sub_468_n10), .CI(
        u4_sub_468_carry_1_), .CO(u4_sub_468_carry_2_), .S(u4_exp_next_mi_1_)
         );
  FA_X1 u4_sub_468_U2_2 ( .A(u4_exp_in_pl1_2_), .B(u4_sub_468_n11), .CI(
        u4_sub_468_carry_2_), .CO(u4_sub_468_carry_3_), .S(u4_exp_next_mi_2_)
         );
  FA_X1 u4_sub_468_U2_3 ( .A(u4_exp_in_pl1_3_), .B(u4_sub_468_n12), .CI(
        u4_sub_468_carry_3_), .CO(u4_sub_468_carry_4_), .S(u4_exp_next_mi_3_)
         );
  FA_X1 u4_sub_468_U2_4 ( .A(u4_exp_in_pl1_4_), .B(u4_sub_468_n13), .CI(
        u4_sub_468_carry_4_), .CO(u4_sub_468_carry_5_), .S(u4_exp_next_mi_4_)
         );
  FA_X1 u4_sub_468_U2_5 ( .A(u4_exp_in_pl1_5_), .B(u4_sub_468_n14), .CI(
        u4_sub_468_carry_5_), .CO(u4_sub_468_carry_6_), .S(u4_exp_next_mi_5_)
         );
  FA_X1 u4_sub_468_U2_6 ( .A(u4_exp_in_pl1_6_), .B(u4_sub_468_n15), .CI(
        u4_sub_468_carry_6_), .CO(u4_sub_468_carry_7_), .S(u4_exp_next_mi_6_)
         );
  INV_X4 u4_sub_494_U23 ( .A(u4_ldz_all_0_), .ZN(u4_sub_494_n14) );
  INV_X4 u4_sub_494_U22 ( .A(u4_ldz_all_1_), .ZN(u4_sub_494_n13) );
  INV_X4 u4_sub_494_U21 ( .A(u4_ldz_all_2_), .ZN(u4_sub_494_n12) );
  INV_X4 u4_sub_494_U20 ( .A(u4_ldz_all_3_), .ZN(u4_sub_494_n11) );
  INV_X4 u4_sub_494_U19 ( .A(u4_ldz_all_4_), .ZN(u4_sub_494_n10) );
  INV_X4 u4_sub_494_U18 ( .A(u4_ldz_all_5_), .ZN(u4_sub_494_n9) );
  INV_X4 u4_sub_494_U17 ( .A(u4_ldz_all_6_), .ZN(u4_sub_494_n8) );
  INV_X4 u4_sub_494_U16 ( .A(u4_exp_in_pl1_0_), .ZN(u4_sub_494_n7) );
  XNOR2_X2 u4_sub_494_U15 ( .A(u4_sub_494_n14), .B(u4_exp_in_pl1_0_), .ZN(
        u4_div_exp2_0_) );
  NAND2_X2 u4_sub_494_U14 ( .A1(u4_ldz_all_0_), .A2(u4_sub_494_n7), .ZN(
        u4_sub_494_carry_1_) );
  INV_X4 u4_sub_494_U13 ( .A(u4_sub_494_carry_9_), .ZN(u4_sub_494_n6) );
  INV_X4 u4_sub_494_U12 ( .A(u4_exp_in_pl1_9_), .ZN(u4_sub_494_n5) );
  XNOR2_X2 u4_sub_494_U11 ( .A(u4_exp_in_pl1_9_), .B(u4_sub_494_carry_9_), 
        .ZN(u4_div_exp2_9_) );
  NAND2_X2 u4_sub_494_U10 ( .A1(u4_sub_494_n5), .A2(u4_sub_494_n6), .ZN(
        u4_sub_494_carry_10_) );
  INV_X4 u4_sub_494_U9 ( .A(u4_sub_494_carry_8_), .ZN(u4_sub_494_n4) );
  INV_X4 u4_sub_494_U8 ( .A(u4_exp_in_pl1_8_), .ZN(u4_sub_494_n3) );
  XNOR2_X2 u4_sub_494_U7 ( .A(u4_exp_in_pl1_8_), .B(u4_sub_494_carry_8_), .ZN(
        u4_div_exp2_8_) );
  NAND2_X2 u4_sub_494_U6 ( .A1(u4_sub_494_n3), .A2(u4_sub_494_n4), .ZN(
        u4_sub_494_carry_9_) );
  INV_X4 u4_sub_494_U5 ( .A(u4_sub_494_carry_7_), .ZN(u4_sub_494_n2) );
  INV_X4 u4_sub_494_U4 ( .A(u4_exp_in_pl1_7_), .ZN(u4_sub_494_n1) );
  XNOR2_X2 u4_sub_494_U3 ( .A(u4_exp_in_pl1_7_), .B(u4_sub_494_carry_7_), .ZN(
        u4_div_exp2_7_) );
  NAND2_X2 u4_sub_494_U2 ( .A1(u4_sub_494_n1), .A2(u4_sub_494_n2), .ZN(
        u4_sub_494_carry_8_) );
  XNOR2_X2 u4_sub_494_U1 ( .A(u4_exp_in_pl1_10_), .B(u4_sub_494_carry_10_), 
        .ZN(u4_div_exp2_10_) );
  FA_X1 u4_sub_494_U2_1 ( .A(u4_exp_in_pl1_1_), .B(u4_sub_494_n13), .CI(
        u4_sub_494_carry_1_), .CO(u4_sub_494_carry_2_), .S(u4_div_exp2_1_) );
  FA_X1 u4_sub_494_U2_2 ( .A(u4_exp_in_pl1_2_), .B(u4_sub_494_n12), .CI(
        u4_sub_494_carry_2_), .CO(u4_sub_494_carry_3_), .S(u4_div_exp2_2_) );
  FA_X1 u4_sub_494_U2_3 ( .A(u4_exp_in_pl1_3_), .B(u4_sub_494_n11), .CI(
        u4_sub_494_carry_3_), .CO(u4_sub_494_carry_4_), .S(u4_div_exp2_3_) );
  FA_X1 u4_sub_494_U2_4 ( .A(u4_exp_in_pl1_4_), .B(u4_sub_494_n10), .CI(
        u4_sub_494_carry_4_), .CO(u4_sub_494_carry_5_), .S(u4_div_exp2_4_) );
  FA_X1 u4_sub_494_U2_5 ( .A(u4_exp_in_pl1_5_), .B(u4_sub_494_n9), .CI(
        u4_sub_494_carry_5_), .CO(u4_sub_494_carry_6_), .S(u4_div_exp2_5_) );
  FA_X1 u4_sub_494_U2_6 ( .A(u4_exp_in_pl1_6_), .B(u4_sub_494_n8), .CI(
        u4_sub_494_carry_6_), .CO(u4_sub_494_carry_7_), .S(u4_div_exp2_6_) );
  AND2_X4 u4_add_487_U5 ( .A1(u4_fi_ldz_5_), .A2(u4_add_487_carry_5_), .ZN(
        u4_add_487_n5) );
  AND2_X4 u4_add_487_U4 ( .A1(u4_fi_ldz_2a_0_), .A2(div_opa_ldz_r2[0]), .ZN(
        u4_add_487_n4) );
  XOR2_X2 u4_add_487_U3 ( .A(u4_fi_ldz_5_), .B(u4_add_487_carry_5_), .Z(
        u4_ldz_all_5_) );
  XOR2_X2 u4_add_487_U2 ( .A(u4_fi_ldz_6_), .B(u4_add_487_n5), .Z(
        u4_ldz_all_6_) );
  XOR2_X2 u4_add_487_U1 ( .A(u4_fi_ldz_2a_0_), .B(div_opa_ldz_r2[0]), .Z(
        u4_ldz_all_0_) );
  FA_X1 u4_add_487_U1_1 ( .A(div_opa_ldz_r2[1]), .B(u4_fi_ldz_1_), .CI(
        u4_add_487_n4), .CO(u4_add_487_carry_2_), .S(u4_ldz_all_1_) );
  FA_X1 u4_add_487_U1_2 ( .A(div_opa_ldz_r2[2]), .B(u4_fi_ldz_2_), .CI(
        u4_add_487_carry_2_), .CO(u4_add_487_carry_3_), .S(u4_ldz_all_2_) );
  FA_X1 u4_add_487_U1_3 ( .A(div_opa_ldz_r2[3]), .B(u4_fi_ldz_3_), .CI(
        u4_add_487_carry_3_), .CO(u4_add_487_carry_4_), .S(u4_ldz_all_3_) );
  FA_X1 u4_add_487_U1_4 ( .A(div_opa_ldz_r2[4]), .B(u4_fi_ldz_4_), .CI(
        u4_add_487_carry_4_), .CO(u4_add_487_carry_5_), .S(u4_ldz_all_4_) );
  INV_X4 u4_add_464_U1 ( .A(n4823), .ZN(u4_exp_in_pl1_0_) );
  HA_X1 u4_add_464_U1_1_1 ( .A(n4368), .B(n4823), .CO(u4_add_464_carry[2]), 
        .S(u4_exp_in_pl1_1_) );
  HA_X1 u4_add_464_U1_1_2 ( .A(exp_r[2]), .B(u4_add_464_carry[2]), .CO(
        u4_add_464_carry[3]), .S(u4_exp_in_pl1_2_) );
  HA_X1 u4_add_464_U1_1_3 ( .A(exp_r[3]), .B(u4_add_464_carry[3]), .CO(
        u4_add_464_carry[4]), .S(u4_exp_in_pl1_3_) );
  HA_X1 u4_add_464_U1_1_4 ( .A(n4399), .B(u4_add_464_carry[4]), .CO(
        u4_add_464_carry[5]), .S(u4_exp_in_pl1_4_) );
  HA_X1 u4_add_464_U1_1_5 ( .A(n4370), .B(u4_add_464_carry[5]), .CO(
        u4_add_464_carry[6]), .S(u4_exp_in_pl1_5_) );
  HA_X1 u4_add_464_U1_1_6 ( .A(n4382), .B(u4_add_464_carry[6]), .CO(
        u4_add_464_carry[7]), .S(u4_exp_in_pl1_6_) );
  HA_X1 u4_add_464_U1_1_7 ( .A(n4359), .B(u4_add_464_carry[7]), .CO(
        u4_add_464_carry[8]), .S(u4_exp_in_pl1_7_) );
  HA_X1 u4_add_464_U1_1_8 ( .A(n4369), .B(u4_add_464_carry[8]), .CO(
        u4_add_464_carry[9]), .S(u4_exp_in_pl1_8_) );
  HA_X1 u4_add_464_U1_1_9 ( .A(n4428), .B(u4_add_464_carry[9]), .CO(
        u4_add_464_carry[10]), .S(u4_exp_in_pl1_9_) );
  HA_X1 u4_add_464_U1_1_10 ( .A(n4875), .B(u4_add_464_carry[10]), .CO(
        u4_exp_in_pl1_11_), .S(u4_exp_in_pl1_10_) );
  XOR2_X2 u4_add_492_U7 ( .A(u4_exp_in_mi1_10_), .B(u4_add_492_n6), .Z(
        u4_div_exp1_10_) );
  AND2_X4 u4_add_492_U6 ( .A1(u4_exp_in_mi1_9_), .A2(u4_add_492_n4), .ZN(
        u4_add_492_n6) );
  XOR2_X2 u4_add_492_U5 ( .A(u4_exp_in_mi1_9_), .B(u4_add_492_n4), .Z(
        u4_div_exp1_9_) );
  AND2_X4 u4_add_492_U4 ( .A1(u4_exp_in_mi1_8_), .A2(u4_add_492_carry_8_), 
        .ZN(u4_add_492_n4) );
  AND2_X4 u4_add_492_U3 ( .A1(u4_fi_ldz_2a_0_), .A2(n4400), .ZN(u4_add_492_n3)
         );
  XOR2_X2 u4_add_492_U2 ( .A(u4_fi_ldz_2a_0_), .B(n4400), .Z(u4_div_exp1_0_)
         );
  XOR2_X2 u4_add_492_U1 ( .A(u4_exp_in_mi1_8_), .B(u4_add_492_carry_8_), .Z(
        u4_div_exp1_8_) );
  FA_X1 u4_add_492_U1_1 ( .A(u4_exp_in_mi1_1_), .B(u4_fi_ldz_2a_1_), .CI(
        u4_add_492_n3), .CO(u4_add_492_carry_2_), .S(u4_div_exp1_1_) );
  FA_X1 u4_add_492_U1_2 ( .A(u4_exp_in_mi1_2_), .B(u4_fi_ldz_2a_2_), .CI(
        u4_add_492_carry_2_), .CO(u4_add_492_carry_3_), .S(u4_div_exp1_2_) );
  FA_X1 u4_add_492_U1_3 ( .A(u4_exp_in_mi1_3_), .B(u4_fi_ldz_2a_3_), .CI(
        u4_add_492_carry_3_), .CO(u4_add_492_carry_4_), .S(u4_div_exp1_3_) );
  FA_X1 u4_add_492_U1_4 ( .A(u4_exp_in_mi1_4_), .B(u4_fi_ldz_2a_4_), .CI(
        u4_add_492_carry_4_), .CO(u4_add_492_carry_5_), .S(u4_div_exp1_4_) );
  FA_X1 u4_add_492_U1_5 ( .A(u4_exp_in_mi1_5_), .B(u4_fi_ldz_2a_5_), .CI(
        u4_add_492_carry_5_), .CO(u4_add_492_carry_6_), .S(u4_div_exp1_5_) );
  FA_X1 u4_add_492_U1_6 ( .A(u4_exp_in_mi1_6_), .B(u4_fi_ldz_2a_6_), .CI(
        u4_add_492_carry_6_), .CO(u4_add_492_carry_7_), .S(u4_div_exp1_6_) );
  FA_X1 u4_add_492_U1_7 ( .A(u4_exp_in_mi1_7_), .B(u4_fi_ldz_2a_6_), .CI(
        u4_add_492_carry_7_), .CO(u4_add_492_carry_8_), .S(u4_div_exp1_7_) );
  INV_X1 u4_add_394_U1 ( .A(u4_fract_out_0_), .ZN(u4_fract_out_pl1_0_) );
  HA_X1 u4_add_394_U1_1_1 ( .A(u4_fract_out_1_), .B(u4_fract_out_0_), .CO(
        u4_add_394_carry[2]), .S(u4_fract_out_pl1_1_) );
  HA_X1 u4_add_394_U1_1_2 ( .A(u4_fract_out_2_), .B(u4_add_394_carry[2]), .CO(
        u4_add_394_carry[3]), .S(u4_fract_out_pl1_2_) );
  HA_X1 u4_add_394_U1_1_3 ( .A(u4_fract_out_3_), .B(u4_add_394_carry[3]), .CO(
        u4_add_394_carry[4]), .S(u4_fract_out_pl1_3_) );
  HA_X1 u4_add_394_U1_1_4 ( .A(u4_fract_out_4_), .B(u4_add_394_carry[4]), .CO(
        u4_add_394_carry[5]), .S(u4_fract_out_pl1_4_) );
  HA_X1 u4_add_394_U1_1_5 ( .A(u4_fract_out_5_), .B(u4_add_394_carry[5]), .CO(
        u4_add_394_carry[6]), .S(u4_fract_out_pl1_5_) );
  HA_X1 u4_add_394_U1_1_6 ( .A(u4_fract_out_6_), .B(u4_add_394_carry[6]), .CO(
        u4_add_394_carry[7]), .S(u4_fract_out_pl1_6_) );
  HA_X1 u4_add_394_U1_1_7 ( .A(u4_fract_out_7_), .B(u4_add_394_carry[7]), .CO(
        u4_add_394_carry[8]), .S(u4_fract_out_pl1_7_) );
  HA_X1 u4_add_394_U1_1_8 ( .A(u4_fract_out_8_), .B(u4_add_394_carry[8]), .CO(
        u4_add_394_carry[9]), .S(u4_fract_out_pl1_8_) );
  HA_X1 u4_add_394_U1_1_9 ( .A(u4_fract_out_9_), .B(u4_add_394_carry[9]), .CO(
        u4_add_394_carry[10]), .S(u4_fract_out_pl1_9_) );
  HA_X1 u4_add_394_U1_1_10 ( .A(u4_fract_out_10_), .B(u4_add_394_carry[10]), 
        .CO(u4_add_394_carry[11]), .S(u4_fract_out_pl1_10_) );
  HA_X1 u4_add_394_U1_1_11 ( .A(u4_fract_out_11_), .B(u4_add_394_carry[11]), 
        .CO(u4_add_394_carry[12]), .S(u4_fract_out_pl1_11_) );
  HA_X1 u4_add_394_U1_1_12 ( .A(u4_fract_out_12_), .B(u4_add_394_carry[12]), 
        .CO(u4_add_394_carry[13]), .S(u4_fract_out_pl1_12_) );
  HA_X1 u4_add_394_U1_1_13 ( .A(u4_fract_out_13_), .B(u4_add_394_carry[13]), 
        .CO(u4_add_394_carry[14]), .S(u4_fract_out_pl1_13_) );
  HA_X1 u4_add_394_U1_1_14 ( .A(u4_fract_out_14_), .B(u4_add_394_carry[14]), 
        .CO(u4_add_394_carry[15]), .S(u4_fract_out_pl1_14_) );
  HA_X1 u4_add_394_U1_1_15 ( .A(u4_fract_out_15_), .B(u4_add_394_carry[15]), 
        .CO(u4_add_394_carry[16]), .S(u4_fract_out_pl1_15_) );
  HA_X1 u4_add_394_U1_1_16 ( .A(u4_fract_out_16_), .B(u4_add_394_carry[16]), 
        .CO(u4_add_394_carry[17]), .S(u4_fract_out_pl1_16_) );
  HA_X1 u4_add_394_U1_1_17 ( .A(u4_fract_out_17_), .B(u4_add_394_carry[17]), 
        .CO(u4_add_394_carry[18]), .S(u4_fract_out_pl1_17_) );
  HA_X1 u4_add_394_U1_1_18 ( .A(u4_fract_out_18_), .B(u4_add_394_carry[18]), 
        .CO(u4_add_394_carry[19]), .S(u4_fract_out_pl1_18_) );
  HA_X1 u4_add_394_U1_1_19 ( .A(u4_fract_out_19_), .B(u4_add_394_carry[19]), 
        .CO(u4_add_394_carry[20]), .S(u4_fract_out_pl1_19_) );
  HA_X1 u4_add_394_U1_1_20 ( .A(u4_fract_out_20_), .B(u4_add_394_carry[20]), 
        .CO(u4_add_394_carry[21]), .S(u4_fract_out_pl1_20_) );
  HA_X1 u4_add_394_U1_1_21 ( .A(u4_fract_out_21_), .B(u4_add_394_carry[21]), 
        .CO(u4_add_394_carry[22]), .S(u4_fract_out_pl1_21_) );
  HA_X1 u4_add_394_U1_1_22 ( .A(u4_fract_out_22_), .B(u4_add_394_carry[22]), 
        .CO(u4_add_394_carry[23]), .S(u4_fract_out_pl1_22_) );
  HA_X1 u4_add_394_U1_1_23 ( .A(u4_fract_out_23_), .B(u4_add_394_carry[23]), 
        .CO(u4_add_394_carry[24]), .S(u4_fract_out_pl1_23_) );
  HA_X1 u4_add_394_U1_1_24 ( .A(u4_fract_out_24_), .B(u4_add_394_carry[24]), 
        .CO(u4_add_394_carry[25]), .S(u4_fract_out_pl1_24_) );
  HA_X1 u4_add_394_U1_1_25 ( .A(u4_fract_out_25_), .B(u4_add_394_carry[25]), 
        .CO(u4_add_394_carry[26]), .S(u4_fract_out_pl1_25_) );
  HA_X1 u4_add_394_U1_1_26 ( .A(u4_fract_out_26_), .B(u4_add_394_carry[26]), 
        .CO(u4_add_394_carry[27]), .S(u4_fract_out_pl1_26_) );
  HA_X1 u4_add_394_U1_1_27 ( .A(u4_fract_out_27_), .B(u4_add_394_carry[27]), 
        .CO(u4_add_394_carry[28]), .S(u4_fract_out_pl1_27_) );
  HA_X1 u4_add_394_U1_1_28 ( .A(u4_fract_out_28_), .B(u4_add_394_carry[28]), 
        .CO(u4_add_394_carry[29]), .S(u4_fract_out_pl1_28_) );
  HA_X1 u4_add_394_U1_1_29 ( .A(u4_fract_out_29_), .B(u4_add_394_carry[29]), 
        .CO(u4_add_394_carry[30]), .S(u4_fract_out_pl1_29_) );
  HA_X1 u4_add_394_U1_1_30 ( .A(u4_fract_out_30_), .B(u4_add_394_carry[30]), 
        .CO(u4_add_394_carry[31]), .S(u4_fract_out_pl1_30_) );
  HA_X1 u4_add_394_U1_1_31 ( .A(u4_fract_out_31_), .B(u4_add_394_carry[31]), 
        .CO(u4_add_394_carry[32]), .S(u4_fract_out_pl1_31_) );
  HA_X1 u4_add_394_U1_1_32 ( .A(u4_fract_out_32_), .B(u4_add_394_carry[32]), 
        .CO(u4_add_394_carry[33]), .S(u4_fract_out_pl1_32_) );
  HA_X1 u4_add_394_U1_1_33 ( .A(u4_fract_out_33_), .B(u4_add_394_carry[33]), 
        .CO(u4_add_394_carry[34]), .S(u4_fract_out_pl1_33_) );
  HA_X1 u4_add_394_U1_1_34 ( .A(u4_fract_out_34_), .B(u4_add_394_carry[34]), 
        .CO(u4_add_394_carry[35]), .S(u4_fract_out_pl1_34_) );
  HA_X1 u4_add_394_U1_1_35 ( .A(u4_fract_out_35_), .B(u4_add_394_carry[35]), 
        .CO(u4_add_394_carry[36]), .S(u4_fract_out_pl1_35_) );
  HA_X1 u4_add_394_U1_1_36 ( .A(u4_fract_out_36_), .B(u4_add_394_carry[36]), 
        .CO(u4_add_394_carry[37]), .S(u4_fract_out_pl1_36_) );
  HA_X1 u4_add_394_U1_1_37 ( .A(u4_fract_out_37_), .B(u4_add_394_carry[37]), 
        .CO(u4_add_394_carry[38]), .S(u4_fract_out_pl1_37_) );
  HA_X1 u4_add_394_U1_1_38 ( .A(u4_fract_out_38_), .B(u4_add_394_carry[38]), 
        .CO(u4_add_394_carry[39]), .S(u4_fract_out_pl1_38_) );
  HA_X1 u4_add_394_U1_1_39 ( .A(u4_fract_out_39_), .B(u4_add_394_carry[39]), 
        .CO(u4_add_394_carry[40]), .S(u4_fract_out_pl1_39_) );
  HA_X1 u4_add_394_U1_1_40 ( .A(u4_fract_out_40_), .B(u4_add_394_carry[40]), 
        .CO(u4_add_394_carry[41]), .S(u4_fract_out_pl1_40_) );
  HA_X1 u4_add_394_U1_1_41 ( .A(u4_fract_out_41_), .B(u4_add_394_carry[41]), 
        .CO(u4_add_394_carry[42]), .S(u4_fract_out_pl1_41_) );
  HA_X1 u4_add_394_U1_1_42 ( .A(u4_fract_out_42_), .B(u4_add_394_carry[42]), 
        .CO(u4_add_394_carry[43]), .S(u4_fract_out_pl1_42_) );
  HA_X1 u4_add_394_U1_1_43 ( .A(u4_fract_out_43_), .B(u4_add_394_carry[43]), 
        .CO(u4_add_394_carry[44]), .S(u4_fract_out_pl1_43_) );
  HA_X1 u4_add_394_U1_1_44 ( .A(u4_fract_out_44_), .B(u4_add_394_carry[44]), 
        .CO(u4_add_394_carry[45]), .S(u4_fract_out_pl1_44_) );
  HA_X1 u4_add_394_U1_1_45 ( .A(u4_fract_out_45_), .B(u4_add_394_carry[45]), 
        .CO(u4_add_394_carry[46]), .S(u4_fract_out_pl1_45_) );
  HA_X1 u4_add_394_U1_1_46 ( .A(u4_fract_out_46_), .B(u4_add_394_carry[46]), 
        .CO(u4_add_394_carry[47]), .S(u4_fract_out_pl1_46_) );
  HA_X1 u4_add_394_U1_1_47 ( .A(u4_fract_out_47_), .B(u4_add_394_carry[47]), 
        .CO(u4_add_394_carry[48]), .S(u4_fract_out_pl1_47_) );
  HA_X1 u4_add_394_U1_1_48 ( .A(u4_fract_out_48_), .B(u4_add_394_carry[48]), 
        .CO(u4_add_394_carry[49]), .S(u4_fract_out_pl1_48_) );
  HA_X1 u4_add_394_U1_1_49 ( .A(u4_fract_out_49_), .B(u4_add_394_carry[49]), 
        .CO(u4_add_394_carry[50]), .S(u4_fract_out_pl1_49_) );
  HA_X1 u4_add_394_U1_1_50 ( .A(u4_fract_out_50_), .B(u4_add_394_carry[50]), 
        .CO(u4_add_394_carry[51]), .S(u4_fract_out_pl1_50_) );
  HA_X1 u4_add_394_U1_1_51 ( .A(u4_fract_out_51_), .B(u4_add_394_carry[51]), 
        .CO(u4_fract_out_pl1_52_), .S(u4_fract_out_pl1_51_) );
  INV_X4 u3_sub_61_U60 ( .A(fractb[0]), .ZN(u3_sub_61_n58) );
  INV_X4 u3_sub_61_U59 ( .A(fractb[10]), .ZN(u3_sub_61_n57) );
  INV_X4 u3_sub_61_U58 ( .A(fractb[11]), .ZN(u3_sub_61_n56) );
  INV_X4 u3_sub_61_U57 ( .A(fractb[12]), .ZN(u3_sub_61_n55) );
  INV_X4 u3_sub_61_U56 ( .A(fractb[13]), .ZN(u3_sub_61_n54) );
  INV_X4 u3_sub_61_U55 ( .A(fractb[14]), .ZN(u3_sub_61_n53) );
  INV_X4 u3_sub_61_U54 ( .A(fractb[15]), .ZN(u3_sub_61_n52) );
  INV_X4 u3_sub_61_U53 ( .A(fractb[16]), .ZN(u3_sub_61_n51) );
  INV_X4 u3_sub_61_U52 ( .A(fractb[17]), .ZN(u3_sub_61_n50) );
  INV_X4 u3_sub_61_U51 ( .A(fractb[18]), .ZN(u3_sub_61_n49) );
  INV_X4 u3_sub_61_U50 ( .A(fractb[19]), .ZN(u3_sub_61_n48) );
  INV_X4 u3_sub_61_U49 ( .A(fractb[1]), .ZN(u3_sub_61_n47) );
  INV_X4 u3_sub_61_U48 ( .A(fractb[20]), .ZN(u3_sub_61_n46) );
  INV_X4 u3_sub_61_U47 ( .A(fractb[21]), .ZN(u3_sub_61_n45) );
  INV_X4 u3_sub_61_U46 ( .A(fractb[22]), .ZN(u3_sub_61_n44) );
  INV_X4 u3_sub_61_U45 ( .A(fractb[23]), .ZN(u3_sub_61_n43) );
  INV_X4 u3_sub_61_U44 ( .A(fractb[24]), .ZN(u3_sub_61_n42) );
  INV_X4 u3_sub_61_U43 ( .A(fractb[25]), .ZN(u3_sub_61_n41) );
  INV_X4 u3_sub_61_U42 ( .A(fractb[26]), .ZN(u3_sub_61_n40) );
  INV_X4 u3_sub_61_U41 ( .A(fractb[27]), .ZN(u3_sub_61_n39) );
  INV_X4 u3_sub_61_U40 ( .A(fractb[28]), .ZN(u3_sub_61_n38) );
  INV_X4 u3_sub_61_U39 ( .A(fractb[29]), .ZN(u3_sub_61_n37) );
  INV_X4 u3_sub_61_U38 ( .A(fractb[2]), .ZN(u3_sub_61_n36) );
  INV_X4 u3_sub_61_U37 ( .A(fractb[30]), .ZN(u3_sub_61_n35) );
  INV_X4 u3_sub_61_U36 ( .A(fractb[31]), .ZN(u3_sub_61_n34) );
  INV_X4 u3_sub_61_U35 ( .A(fractb[32]), .ZN(u3_sub_61_n33) );
  INV_X4 u3_sub_61_U34 ( .A(fractb[33]), .ZN(u3_sub_61_n32) );
  INV_X4 u3_sub_61_U33 ( .A(fractb[34]), .ZN(u3_sub_61_n31) );
  INV_X4 u3_sub_61_U32 ( .A(fractb[35]), .ZN(u3_sub_61_n30) );
  INV_X4 u3_sub_61_U31 ( .A(fractb[36]), .ZN(u3_sub_61_n29) );
  INV_X4 u3_sub_61_U30 ( .A(fractb[37]), .ZN(u3_sub_61_n28) );
  INV_X4 u3_sub_61_U29 ( .A(fractb[38]), .ZN(u3_sub_61_n27) );
  INV_X4 u3_sub_61_U28 ( .A(fractb[39]), .ZN(u3_sub_61_n26) );
  INV_X4 u3_sub_61_U27 ( .A(fractb[3]), .ZN(u3_sub_61_n25) );
  INV_X4 u3_sub_61_U26 ( .A(fractb[40]), .ZN(u3_sub_61_n24) );
  INV_X4 u3_sub_61_U25 ( .A(fractb[41]), .ZN(u3_sub_61_n23) );
  INV_X4 u3_sub_61_U24 ( .A(fractb[42]), .ZN(u3_sub_61_n22) );
  INV_X4 u3_sub_61_U23 ( .A(fractb[43]), .ZN(u3_sub_61_n21) );
  INV_X4 u3_sub_61_U22 ( .A(fractb[44]), .ZN(u3_sub_61_n20) );
  INV_X4 u3_sub_61_U21 ( .A(fractb[45]), .ZN(u3_sub_61_n19) );
  INV_X4 u3_sub_61_U20 ( .A(fractb[46]), .ZN(u3_sub_61_n18) );
  INV_X4 u3_sub_61_U19 ( .A(fractb[47]), .ZN(u3_sub_61_n17) );
  INV_X4 u3_sub_61_U18 ( .A(fractb[48]), .ZN(u3_sub_61_n16) );
  INV_X4 u3_sub_61_U17 ( .A(fractb[49]), .ZN(u3_sub_61_n15) );
  INV_X4 u3_sub_61_U16 ( .A(fractb[4]), .ZN(u3_sub_61_n14) );
  INV_X4 u3_sub_61_U15 ( .A(fractb[50]), .ZN(u3_sub_61_n13) );
  INV_X4 u3_sub_61_U14 ( .A(fractb[51]), .ZN(u3_sub_61_n12) );
  INV_X4 u3_sub_61_U13 ( .A(fractb[52]), .ZN(u3_sub_61_n11) );
  INV_X4 u3_sub_61_U12 ( .A(fractb[53]), .ZN(u3_sub_61_n10) );
  INV_X4 u3_sub_61_U11 ( .A(fractb[54]), .ZN(u3_sub_61_n9) );
  INV_X4 u3_sub_61_U10 ( .A(fractb[55]), .ZN(u3_sub_61_n8) );
  INV_X4 u3_sub_61_U9 ( .A(fractb[5]), .ZN(u3_sub_61_n7) );
  INV_X4 u3_sub_61_U8 ( .A(fractb[6]), .ZN(u3_sub_61_n6) );
  INV_X4 u3_sub_61_U7 ( .A(fractb[7]), .ZN(u3_sub_61_n5) );
  INV_X4 u3_sub_61_U6 ( .A(fractb[8]), .ZN(u3_sub_61_n4) );
  INV_X4 u3_sub_61_U5 ( .A(fractb[9]), .ZN(u3_sub_61_n3) );
  INV_X4 u3_sub_61_U4 ( .A(u3_sub_61_carry[56]), .ZN(u3_N116) );
  INV_X4 u3_sub_61_U3 ( .A(fracta[0]), .ZN(u3_sub_61_n1) );
  XNOR2_X2 u3_sub_61_U2 ( .A(u3_sub_61_n58), .B(fracta[0]), .ZN(u3_N60) );
  NAND2_X2 u3_sub_61_U1 ( .A1(fractb[0]), .A2(u3_sub_61_n1), .ZN(
        u3_sub_61_carry[1]) );
  FA_X1 u3_sub_61_U2_1 ( .A(fracta[1]), .B(u3_sub_61_n47), .CI(
        u3_sub_61_carry[1]), .CO(u3_sub_61_carry[2]), .S(u3_N61) );
  FA_X1 u3_sub_61_U2_2 ( .A(fracta[2]), .B(u3_sub_61_n36), .CI(
        u3_sub_61_carry[2]), .CO(u3_sub_61_carry[3]), .S(u3_N62) );
  FA_X1 u3_sub_61_U2_3 ( .A(fracta[3]), .B(u3_sub_61_n25), .CI(
        u3_sub_61_carry[3]), .CO(u3_sub_61_carry[4]), .S(u3_N63) );
  FA_X1 u3_sub_61_U2_4 ( .A(fracta[4]), .B(u3_sub_61_n14), .CI(
        u3_sub_61_carry[4]), .CO(u3_sub_61_carry[5]), .S(u3_N64) );
  FA_X1 u3_sub_61_U2_5 ( .A(fracta[5]), .B(u3_sub_61_n7), .CI(
        u3_sub_61_carry[5]), .CO(u3_sub_61_carry[6]), .S(u3_N65) );
  FA_X1 u3_sub_61_U2_6 ( .A(fracta[6]), .B(u3_sub_61_n6), .CI(
        u3_sub_61_carry[6]), .CO(u3_sub_61_carry[7]), .S(u3_N66) );
  FA_X1 u3_sub_61_U2_7 ( .A(fracta[7]), .B(u3_sub_61_n5), .CI(
        u3_sub_61_carry[7]), .CO(u3_sub_61_carry[8]), .S(u3_N67) );
  FA_X1 u3_sub_61_U2_8 ( .A(fracta[8]), .B(u3_sub_61_n4), .CI(
        u3_sub_61_carry[8]), .CO(u3_sub_61_carry[9]), .S(u3_N68) );
  FA_X1 u3_sub_61_U2_9 ( .A(fracta[9]), .B(u3_sub_61_n3), .CI(
        u3_sub_61_carry[9]), .CO(u3_sub_61_carry[10]), .S(u3_N69) );
  FA_X1 u3_sub_61_U2_10 ( .A(fracta[10]), .B(u3_sub_61_n57), .CI(
        u3_sub_61_carry[10]), .CO(u3_sub_61_carry[11]), .S(u3_N70) );
  FA_X1 u3_sub_61_U2_11 ( .A(fracta[11]), .B(u3_sub_61_n56), .CI(
        u3_sub_61_carry[11]), .CO(u3_sub_61_carry[12]), .S(u3_N71) );
  FA_X1 u3_sub_61_U2_12 ( .A(fracta[12]), .B(u3_sub_61_n55), .CI(
        u3_sub_61_carry[12]), .CO(u3_sub_61_carry[13]), .S(u3_N72) );
  FA_X1 u3_sub_61_U2_13 ( .A(fracta[13]), .B(u3_sub_61_n54), .CI(
        u3_sub_61_carry[13]), .CO(u3_sub_61_carry[14]), .S(u3_N73) );
  FA_X1 u3_sub_61_U2_14 ( .A(fracta[14]), .B(u3_sub_61_n53), .CI(
        u3_sub_61_carry[14]), .CO(u3_sub_61_carry[15]), .S(u3_N74) );
  FA_X1 u3_sub_61_U2_15 ( .A(fracta[15]), .B(u3_sub_61_n52), .CI(
        u3_sub_61_carry[15]), .CO(u3_sub_61_carry[16]), .S(u3_N75) );
  FA_X1 u3_sub_61_U2_16 ( .A(fracta[16]), .B(u3_sub_61_n51), .CI(
        u3_sub_61_carry[16]), .CO(u3_sub_61_carry[17]), .S(u3_N76) );
  FA_X1 u3_sub_61_U2_17 ( .A(fracta[17]), .B(u3_sub_61_n50), .CI(
        u3_sub_61_carry[17]), .CO(u3_sub_61_carry[18]), .S(u3_N77) );
  FA_X1 u3_sub_61_U2_18 ( .A(fracta[18]), .B(u3_sub_61_n49), .CI(
        u3_sub_61_carry[18]), .CO(u3_sub_61_carry[19]), .S(u3_N78) );
  FA_X1 u3_sub_61_U2_19 ( .A(fracta[19]), .B(u3_sub_61_n48), .CI(
        u3_sub_61_carry[19]), .CO(u3_sub_61_carry[20]), .S(u3_N79) );
  FA_X1 u3_sub_61_U2_20 ( .A(fracta[20]), .B(u3_sub_61_n46), .CI(
        u3_sub_61_carry[20]), .CO(u3_sub_61_carry[21]), .S(u3_N80) );
  FA_X1 u3_sub_61_U2_21 ( .A(fracta[21]), .B(u3_sub_61_n45), .CI(
        u3_sub_61_carry[21]), .CO(u3_sub_61_carry[22]), .S(u3_N81) );
  FA_X1 u3_sub_61_U2_22 ( .A(fracta[22]), .B(u3_sub_61_n44), .CI(
        u3_sub_61_carry[22]), .CO(u3_sub_61_carry[23]), .S(u3_N82) );
  FA_X1 u3_sub_61_U2_23 ( .A(fracta[23]), .B(u3_sub_61_n43), .CI(
        u3_sub_61_carry[23]), .CO(u3_sub_61_carry[24]), .S(u3_N83) );
  FA_X1 u3_sub_61_U2_24 ( .A(fracta[24]), .B(u3_sub_61_n42), .CI(
        u3_sub_61_carry[24]), .CO(u3_sub_61_carry[25]), .S(u3_N84) );
  FA_X1 u3_sub_61_U2_25 ( .A(fracta[25]), .B(u3_sub_61_n41), .CI(
        u3_sub_61_carry[25]), .CO(u3_sub_61_carry[26]), .S(u3_N85) );
  FA_X1 u3_sub_61_U2_26 ( .A(fracta[26]), .B(u3_sub_61_n40), .CI(
        u3_sub_61_carry[26]), .CO(u3_sub_61_carry[27]), .S(u3_N86) );
  FA_X1 u3_sub_61_U2_27 ( .A(fracta[27]), .B(u3_sub_61_n39), .CI(
        u3_sub_61_carry[27]), .CO(u3_sub_61_carry[28]), .S(u3_N87) );
  FA_X1 u3_sub_61_U2_28 ( .A(fracta[28]), .B(u3_sub_61_n38), .CI(
        u3_sub_61_carry[28]), .CO(u3_sub_61_carry[29]), .S(u3_N88) );
  FA_X1 u3_sub_61_U2_29 ( .A(fracta[29]), .B(u3_sub_61_n37), .CI(
        u3_sub_61_carry[29]), .CO(u3_sub_61_carry[30]), .S(u3_N89) );
  FA_X1 u3_sub_61_U2_30 ( .A(fracta[30]), .B(u3_sub_61_n35), .CI(
        u3_sub_61_carry[30]), .CO(u3_sub_61_carry[31]), .S(u3_N90) );
  FA_X1 u3_sub_61_U2_31 ( .A(fracta[31]), .B(u3_sub_61_n34), .CI(
        u3_sub_61_carry[31]), .CO(u3_sub_61_carry[32]), .S(u3_N91) );
  FA_X1 u3_sub_61_U2_32 ( .A(fracta[32]), .B(u3_sub_61_n33), .CI(
        u3_sub_61_carry[32]), .CO(u3_sub_61_carry[33]), .S(u3_N92) );
  FA_X1 u3_sub_61_U2_33 ( .A(fracta[33]), .B(u3_sub_61_n32), .CI(
        u3_sub_61_carry[33]), .CO(u3_sub_61_carry[34]), .S(u3_N93) );
  FA_X1 u3_sub_61_U2_34 ( .A(fracta[34]), .B(u3_sub_61_n31), .CI(
        u3_sub_61_carry[34]), .CO(u3_sub_61_carry[35]), .S(u3_N94) );
  FA_X1 u3_sub_61_U2_35 ( .A(fracta[35]), .B(u3_sub_61_n30), .CI(
        u3_sub_61_carry[35]), .CO(u3_sub_61_carry[36]), .S(u3_N95) );
  FA_X1 u3_sub_61_U2_36 ( .A(fracta[36]), .B(u3_sub_61_n29), .CI(
        u3_sub_61_carry[36]), .CO(u3_sub_61_carry[37]), .S(u3_N96) );
  FA_X1 u3_sub_61_U2_37 ( .A(fracta[37]), .B(u3_sub_61_n28), .CI(
        u3_sub_61_carry[37]), .CO(u3_sub_61_carry[38]), .S(u3_N97) );
  FA_X1 u3_sub_61_U2_38 ( .A(fracta[38]), .B(u3_sub_61_n27), .CI(
        u3_sub_61_carry[38]), .CO(u3_sub_61_carry[39]), .S(u3_N98) );
  FA_X1 u3_sub_61_U2_39 ( .A(fracta[39]), .B(u3_sub_61_n26), .CI(
        u3_sub_61_carry[39]), .CO(u3_sub_61_carry[40]), .S(u3_N99) );
  FA_X1 u3_sub_61_U2_40 ( .A(fracta[40]), .B(u3_sub_61_n24), .CI(
        u3_sub_61_carry[40]), .CO(u3_sub_61_carry[41]), .S(u3_N100) );
  FA_X1 u3_sub_61_U2_41 ( .A(fracta[41]), .B(u3_sub_61_n23), .CI(
        u3_sub_61_carry[41]), .CO(u3_sub_61_carry[42]), .S(u3_N101) );
  FA_X1 u3_sub_61_U2_42 ( .A(fracta[42]), .B(u3_sub_61_n22), .CI(
        u3_sub_61_carry[42]), .CO(u3_sub_61_carry[43]), .S(u3_N102) );
  FA_X1 u3_sub_61_U2_43 ( .A(fracta[43]), .B(u3_sub_61_n21), .CI(
        u3_sub_61_carry[43]), .CO(u3_sub_61_carry[44]), .S(u3_N103) );
  FA_X1 u3_sub_61_U2_44 ( .A(fracta[44]), .B(u3_sub_61_n20), .CI(
        u3_sub_61_carry[44]), .CO(u3_sub_61_carry[45]), .S(u3_N104) );
  FA_X1 u3_sub_61_U2_45 ( .A(fracta[45]), .B(u3_sub_61_n19), .CI(
        u3_sub_61_carry[45]), .CO(u3_sub_61_carry[46]), .S(u3_N105) );
  FA_X1 u3_sub_61_U2_46 ( .A(fracta[46]), .B(u3_sub_61_n18), .CI(
        u3_sub_61_carry[46]), .CO(u3_sub_61_carry[47]), .S(u3_N106) );
  FA_X1 u3_sub_61_U2_47 ( .A(fracta[47]), .B(u3_sub_61_n17), .CI(
        u3_sub_61_carry[47]), .CO(u3_sub_61_carry[48]), .S(u3_N107) );
  FA_X1 u3_sub_61_U2_48 ( .A(fracta[48]), .B(u3_sub_61_n16), .CI(
        u3_sub_61_carry[48]), .CO(u3_sub_61_carry[49]), .S(u3_N108) );
  FA_X1 u3_sub_61_U2_49 ( .A(fracta[49]), .B(u3_sub_61_n15), .CI(
        u3_sub_61_carry[49]), .CO(u3_sub_61_carry[50]), .S(u3_N109) );
  FA_X1 u3_sub_61_U2_50 ( .A(fracta[50]), .B(u3_sub_61_n13), .CI(
        u3_sub_61_carry[50]), .CO(u3_sub_61_carry[51]), .S(u3_N110) );
  FA_X1 u3_sub_61_U2_51 ( .A(fracta[51]), .B(u3_sub_61_n12), .CI(
        u3_sub_61_carry[51]), .CO(u3_sub_61_carry[52]), .S(u3_N111) );
  FA_X1 u3_sub_61_U2_52 ( .A(fracta[52]), .B(u3_sub_61_n11), .CI(
        u3_sub_61_carry[52]), .CO(u3_sub_61_carry[53]), .S(u3_N112) );
  FA_X1 u3_sub_61_U2_53 ( .A(fracta[53]), .B(u3_sub_61_n10), .CI(
        u3_sub_61_carry[53]), .CO(u3_sub_61_carry[54]), .S(u3_N113) );
  FA_X1 u3_sub_61_U2_54 ( .A(fracta[54]), .B(u3_sub_61_n9), .CI(
        u3_sub_61_carry[54]), .CO(u3_sub_61_carry[55]), .S(u3_N114) );
  FA_X1 u3_sub_61_U2_55 ( .A(fracta[55]), .B(u3_sub_61_n8), .CI(
        u3_sub_61_carry[55]), .CO(u3_sub_61_carry[56]), .S(u3_N115) );
  XOR2_X2 u3_add_61_U2 ( .A(fractb[0]), .B(fracta[0]), .Z(u3_N3) );
  AND2_X4 u3_add_61_U1 ( .A1(fractb[0]), .A2(fracta[0]), .ZN(u3_add_61_n1) );
  FA_X1 u3_add_61_U1_1 ( .A(fracta[1]), .B(fractb[1]), .CI(u3_add_61_n1), .CO(
        u3_add_61_carry[2]), .S(u3_N4) );
  FA_X1 u3_add_61_U1_2 ( .A(fracta[2]), .B(fractb[2]), .CI(u3_add_61_carry[2]), 
        .CO(u3_add_61_carry[3]), .S(u3_N5) );
  FA_X1 u3_add_61_U1_3 ( .A(fracta[3]), .B(fractb[3]), .CI(u3_add_61_carry[3]), 
        .CO(u3_add_61_carry[4]), .S(u3_N6) );
  FA_X1 u3_add_61_U1_4 ( .A(fracta[4]), .B(fractb[4]), .CI(u3_add_61_carry[4]), 
        .CO(u3_add_61_carry[5]), .S(u3_N7) );
  FA_X1 u3_add_61_U1_5 ( .A(fracta[5]), .B(fractb[5]), .CI(u3_add_61_carry[5]), 
        .CO(u3_add_61_carry[6]), .S(u3_N8) );
  FA_X1 u3_add_61_U1_6 ( .A(fracta[6]), .B(fractb[6]), .CI(u3_add_61_carry[6]), 
        .CO(u3_add_61_carry[7]), .S(u3_N9) );
  FA_X1 u3_add_61_U1_7 ( .A(fracta[7]), .B(fractb[7]), .CI(u3_add_61_carry[7]), 
        .CO(u3_add_61_carry[8]), .S(u3_N10) );
  FA_X1 u3_add_61_U1_8 ( .A(fracta[8]), .B(fractb[8]), .CI(u3_add_61_carry[8]), 
        .CO(u3_add_61_carry[9]), .S(u3_N11) );
  FA_X1 u3_add_61_U1_9 ( .A(fracta[9]), .B(fractb[9]), .CI(u3_add_61_carry[9]), 
        .CO(u3_add_61_carry[10]), .S(u3_N12) );
  FA_X1 u3_add_61_U1_10 ( .A(fracta[10]), .B(fractb[10]), .CI(
        u3_add_61_carry[10]), .CO(u3_add_61_carry[11]), .S(u3_N13) );
  FA_X1 u3_add_61_U1_11 ( .A(fracta[11]), .B(fractb[11]), .CI(
        u3_add_61_carry[11]), .CO(u3_add_61_carry[12]), .S(u3_N14) );
  FA_X1 u3_add_61_U1_12 ( .A(fracta[12]), .B(fractb[12]), .CI(
        u3_add_61_carry[12]), .CO(u3_add_61_carry[13]), .S(u3_N15) );
  FA_X1 u3_add_61_U1_13 ( .A(fracta[13]), .B(fractb[13]), .CI(
        u3_add_61_carry[13]), .CO(u3_add_61_carry[14]), .S(u3_N16) );
  FA_X1 u3_add_61_U1_14 ( .A(fracta[14]), .B(fractb[14]), .CI(
        u3_add_61_carry[14]), .CO(u3_add_61_carry[15]), .S(u3_N17) );
  FA_X1 u3_add_61_U1_15 ( .A(fracta[15]), .B(fractb[15]), .CI(
        u3_add_61_carry[15]), .CO(u3_add_61_carry[16]), .S(u3_N18) );
  FA_X1 u3_add_61_U1_16 ( .A(fracta[16]), .B(fractb[16]), .CI(
        u3_add_61_carry[16]), .CO(u3_add_61_carry[17]), .S(u3_N19) );
  FA_X1 u3_add_61_U1_17 ( .A(fracta[17]), .B(fractb[17]), .CI(
        u3_add_61_carry[17]), .CO(u3_add_61_carry[18]), .S(u3_N20) );
  FA_X1 u3_add_61_U1_18 ( .A(fracta[18]), .B(fractb[18]), .CI(
        u3_add_61_carry[18]), .CO(u3_add_61_carry[19]), .S(u3_N21) );
  FA_X1 u3_add_61_U1_19 ( .A(fracta[19]), .B(fractb[19]), .CI(
        u3_add_61_carry[19]), .CO(u3_add_61_carry[20]), .S(u3_N22) );
  FA_X1 u3_add_61_U1_20 ( .A(fracta[20]), .B(fractb[20]), .CI(
        u3_add_61_carry[20]), .CO(u3_add_61_carry[21]), .S(u3_N23) );
  FA_X1 u3_add_61_U1_21 ( .A(fracta[21]), .B(fractb[21]), .CI(
        u3_add_61_carry[21]), .CO(u3_add_61_carry[22]), .S(u3_N24) );
  FA_X1 u3_add_61_U1_22 ( .A(fracta[22]), .B(fractb[22]), .CI(
        u3_add_61_carry[22]), .CO(u3_add_61_carry[23]), .S(u3_N25) );
  FA_X1 u3_add_61_U1_23 ( .A(fracta[23]), .B(fractb[23]), .CI(
        u3_add_61_carry[23]), .CO(u3_add_61_carry[24]), .S(u3_N26) );
  FA_X1 u3_add_61_U1_24 ( .A(fracta[24]), .B(fractb[24]), .CI(
        u3_add_61_carry[24]), .CO(u3_add_61_carry[25]), .S(u3_N27) );
  FA_X1 u3_add_61_U1_25 ( .A(fracta[25]), .B(fractb[25]), .CI(
        u3_add_61_carry[25]), .CO(u3_add_61_carry[26]), .S(u3_N28) );
  FA_X1 u3_add_61_U1_26 ( .A(fracta[26]), .B(fractb[26]), .CI(
        u3_add_61_carry[26]), .CO(u3_add_61_carry[27]), .S(u3_N29) );
  FA_X1 u3_add_61_U1_27 ( .A(fracta[27]), .B(fractb[27]), .CI(
        u3_add_61_carry[27]), .CO(u3_add_61_carry[28]), .S(u3_N30) );
  FA_X1 u3_add_61_U1_28 ( .A(fracta[28]), .B(fractb[28]), .CI(
        u3_add_61_carry[28]), .CO(u3_add_61_carry[29]), .S(u3_N31) );
  FA_X1 u3_add_61_U1_29 ( .A(fracta[29]), .B(fractb[29]), .CI(
        u3_add_61_carry[29]), .CO(u3_add_61_carry[30]), .S(u3_N32) );
  FA_X1 u3_add_61_U1_30 ( .A(fracta[30]), .B(fractb[30]), .CI(
        u3_add_61_carry[30]), .CO(u3_add_61_carry[31]), .S(u3_N33) );
  FA_X1 u3_add_61_U1_31 ( .A(fracta[31]), .B(fractb[31]), .CI(
        u3_add_61_carry[31]), .CO(u3_add_61_carry[32]), .S(u3_N34) );
  FA_X1 u3_add_61_U1_32 ( .A(fracta[32]), .B(fractb[32]), .CI(
        u3_add_61_carry[32]), .CO(u3_add_61_carry[33]), .S(u3_N35) );
  FA_X1 u3_add_61_U1_33 ( .A(fracta[33]), .B(fractb[33]), .CI(
        u3_add_61_carry[33]), .CO(u3_add_61_carry[34]), .S(u3_N36) );
  FA_X1 u3_add_61_U1_34 ( .A(fracta[34]), .B(fractb[34]), .CI(
        u3_add_61_carry[34]), .CO(u3_add_61_carry[35]), .S(u3_N37) );
  FA_X1 u3_add_61_U1_35 ( .A(fracta[35]), .B(fractb[35]), .CI(
        u3_add_61_carry[35]), .CO(u3_add_61_carry[36]), .S(u3_N38) );
  FA_X1 u3_add_61_U1_36 ( .A(fracta[36]), .B(fractb[36]), .CI(
        u3_add_61_carry[36]), .CO(u3_add_61_carry[37]), .S(u3_N39) );
  FA_X1 u3_add_61_U1_37 ( .A(fracta[37]), .B(fractb[37]), .CI(
        u3_add_61_carry[37]), .CO(u3_add_61_carry[38]), .S(u3_N40) );
  FA_X1 u3_add_61_U1_38 ( .A(fracta[38]), .B(fractb[38]), .CI(
        u3_add_61_carry[38]), .CO(u3_add_61_carry[39]), .S(u3_N41) );
  FA_X1 u3_add_61_U1_39 ( .A(fracta[39]), .B(fractb[39]), .CI(
        u3_add_61_carry[39]), .CO(u3_add_61_carry[40]), .S(u3_N42) );
  FA_X1 u3_add_61_U1_40 ( .A(fracta[40]), .B(fractb[40]), .CI(
        u3_add_61_carry[40]), .CO(u3_add_61_carry[41]), .S(u3_N43) );
  FA_X1 u3_add_61_U1_41 ( .A(fracta[41]), .B(fractb[41]), .CI(
        u3_add_61_carry[41]), .CO(u3_add_61_carry[42]), .S(u3_N44) );
  FA_X1 u3_add_61_U1_42 ( .A(fracta[42]), .B(fractb[42]), .CI(
        u3_add_61_carry[42]), .CO(u3_add_61_carry[43]), .S(u3_N45) );
  FA_X1 u3_add_61_U1_43 ( .A(fracta[43]), .B(fractb[43]), .CI(
        u3_add_61_carry[43]), .CO(u3_add_61_carry[44]), .S(u3_N46) );
  FA_X1 u3_add_61_U1_44 ( .A(fracta[44]), .B(fractb[44]), .CI(
        u3_add_61_carry[44]), .CO(u3_add_61_carry[45]), .S(u3_N47) );
  FA_X1 u3_add_61_U1_45 ( .A(fracta[45]), .B(fractb[45]), .CI(
        u3_add_61_carry[45]), .CO(u3_add_61_carry[46]), .S(u3_N48) );
  FA_X1 u3_add_61_U1_46 ( .A(fracta[46]), .B(fractb[46]), .CI(
        u3_add_61_carry[46]), .CO(u3_add_61_carry[47]), .S(u3_N49) );
  FA_X1 u3_add_61_U1_47 ( .A(fracta[47]), .B(fractb[47]), .CI(
        u3_add_61_carry[47]), .CO(u3_add_61_carry[48]), .S(u3_N50) );
  FA_X1 u3_add_61_U1_48 ( .A(fracta[48]), .B(fractb[48]), .CI(
        u3_add_61_carry[48]), .CO(u3_add_61_carry[49]), .S(u3_N51) );
  FA_X1 u3_add_61_U1_49 ( .A(fracta[49]), .B(fractb[49]), .CI(
        u3_add_61_carry[49]), .CO(u3_add_61_carry[50]), .S(u3_N52) );
  FA_X1 u3_add_61_U1_50 ( .A(fracta[50]), .B(fractb[50]), .CI(
        u3_add_61_carry[50]), .CO(u3_add_61_carry[51]), .S(u3_N53) );
  FA_X1 u3_add_61_U1_51 ( .A(fracta[51]), .B(fractb[51]), .CI(
        u3_add_61_carry[51]), .CO(u3_add_61_carry[52]), .S(u3_N54) );
  FA_X1 u3_add_61_U1_52 ( .A(fracta[52]), .B(fractb[52]), .CI(
        u3_add_61_carry[52]), .CO(u3_add_61_carry[53]), .S(u3_N55) );
  FA_X1 u3_add_61_U1_53 ( .A(fracta[53]), .B(fractb[53]), .CI(
        u3_add_61_carry[53]), .CO(u3_add_61_carry[54]), .S(u3_N56) );
  FA_X1 u3_add_61_U1_54 ( .A(fracta[54]), .B(fractb[54]), .CI(
        u3_add_61_carry[54]), .CO(u3_add_61_carry[55]), .S(u3_N57) );
  FA_X1 u3_add_61_U1_55 ( .A(fracta[55]), .B(fractb[55]), .CI(
        u3_add_61_carry[55]), .CO(u3_N59), .S(u3_N58) );
  XOR2_X1 u2_add_116_U2 ( .A(u2_add_116_carry[10]), .B(u2_exp_tmp4_10_), .Z(
        u2_N64) );
  INV_X4 u2_add_116_U1 ( .A(n1054), .ZN(u2_N54) );
  HA_X1 u2_add_116_U1_1_1 ( .A(u2_exp_tmp4_1_), .B(n1054), .CO(
        u2_add_116_carry[2]), .S(u2_N55) );
  HA_X1 u2_add_116_U1_1_2 ( .A(u2_exp_tmp4_2_), .B(u2_add_116_carry[2]), .CO(
        u2_add_116_carry[3]), .S(u2_N56) );
  HA_X1 u2_add_116_U1_1_3 ( .A(u2_exp_tmp4_3_), .B(u2_add_116_carry[3]), .CO(
        u2_add_116_carry[4]), .S(u2_N57) );
  HA_X1 u2_add_116_U1_1_4 ( .A(u2_exp_tmp4_4_), .B(u2_add_116_carry[4]), .CO(
        u2_add_116_carry[5]), .S(u2_N58) );
  HA_X1 u2_add_116_U1_1_5 ( .A(n1052), .B(u2_add_116_carry[5]), .CO(
        u2_add_116_carry[6]), .S(u2_N59) );
  HA_X1 u2_add_116_U1_1_6 ( .A(n1051), .B(u2_add_116_carry[6]), .CO(
        u2_add_116_carry[7]), .S(u2_N60) );
  HA_X1 u2_add_116_U1_1_7 ( .A(n1050), .B(u2_add_116_carry[7]), .CO(
        u2_add_116_carry[8]), .S(u2_N61) );
  HA_X1 u2_add_116_U1_1_8 ( .A(n1049), .B(u2_add_116_carry[8]), .CO(
        u2_add_116_carry[9]), .S(u2_N62) );
  HA_X1 u2_add_116_U1_1_9 ( .A(n1048), .B(u2_add_116_carry[9]), .CO(
        u2_add_116_carry[10]), .S(u2_N63) );
  XOR2_X1 u2_add_114_U2 ( .A(u2_add_114_carry[10]), .B(n6083), .Z(
        u2_exp_tmp3_10_) );
  INV_X4 u2_add_114_U1 ( .A(n6098), .ZN(u2_exp_tmp3_0_) );
  HA_X1 u2_add_114_U1_1_1 ( .A(n6096), .B(n6098), .CO(u2_add_114_carry[2]), 
        .S(u2_exp_tmp3_1_) );
  HA_X1 u2_add_114_U1_1_2 ( .A(n6094), .B(u2_add_114_carry[2]), .CO(
        u2_add_114_carry[3]), .S(u2_exp_tmp3_2_) );
  HA_X1 u2_add_114_U1_1_3 ( .A(n6092), .B(u2_add_114_carry[3]), .CO(
        u2_add_114_carry[4]), .S(u2_exp_tmp3_3_) );
  HA_X1 u2_add_114_U1_1_4 ( .A(n6090), .B(u2_add_114_carry[4]), .CO(
        u2_add_114_carry[5]), .S(u2_exp_tmp3_4_) );
  HA_X1 u2_add_114_U1_1_5 ( .A(n6089), .B(u2_add_114_carry[5]), .CO(
        u2_add_114_carry[6]), .S(u2_exp_tmp3_5_) );
  HA_X1 u2_add_114_U1_1_6 ( .A(n6088), .B(u2_add_114_carry[6]), .CO(
        u2_add_114_carry[7]), .S(u2_exp_tmp3_6_) );
  HA_X1 u2_add_114_U1_1_7 ( .A(n6087), .B(u2_add_114_carry[7]), .CO(
        u2_add_114_carry[8]), .S(u2_exp_tmp3_7_) );
  HA_X1 u2_add_114_U1_1_8 ( .A(n6086), .B(u2_add_114_carry[8]), .CO(
        u2_add_114_carry[9]), .S(u2_exp_tmp3_8_) );
  HA_X1 u2_add_114_U1_1_9 ( .A(n6085), .B(u2_add_114_carry[9]), .CO(
        u2_add_114_carry[10]), .S(u2_exp_tmp3_9_) );
  AND2_X4 u2_add_111_U2 ( .A1(opb_r[52]), .A2(opa_r[52]), .ZN(u2_add_111_n2)
         );
  XOR2_X2 u2_add_111_U1 ( .A(opb_r[52]), .B(opa_r[52]), .Z(u2_N18) );
  FA_X1 u2_add_111_U1_1 ( .A(opa_r[53]), .B(opb_r[53]), .CI(u2_add_111_n2), 
        .CO(u2_add_111_carry[2]), .S(u2_N19) );
  FA_X1 u2_add_111_U1_2 ( .A(opa_r[54]), .B(opb_r[54]), .CI(
        u2_add_111_carry[2]), .CO(u2_add_111_carry[3]), .S(u2_N20) );
  FA_X1 u2_add_111_U1_3 ( .A(opa_r[55]), .B(opb_r[55]), .CI(
        u2_add_111_carry[3]), .CO(u2_add_111_carry[4]), .S(u2_N21) );
  FA_X1 u2_add_111_U1_4 ( .A(opa_r[56]), .B(opb_r[56]), .CI(
        u2_add_111_carry[4]), .CO(u2_add_111_carry[5]), .S(u2_N22) );
  FA_X1 u2_add_111_U1_5 ( .A(opa_r[57]), .B(opb_r[57]), .CI(
        u2_add_111_carry[5]), .CO(u2_add_111_carry[6]), .S(u2_N23) );
  FA_X1 u2_add_111_U1_6 ( .A(opa_r[58]), .B(opb_r[58]), .CI(
        u2_add_111_carry[6]), .CO(u2_add_111_carry[7]), .S(u2_N24) );
  FA_X1 u2_add_111_U1_7 ( .A(opa_r[59]), .B(opb_r[59]), .CI(
        u2_add_111_carry[7]), .CO(u2_add_111_carry[8]), .S(u2_N25) );
  FA_X1 u2_add_111_U1_8 ( .A(opa_r[60]), .B(opb_r[60]), .CI(
        u2_add_111_carry[8]), .CO(u2_add_111_carry[9]), .S(u2_N26) );
  FA_X1 u2_add_111_U1_9 ( .A(opa_r[61]), .B(opb_r[61]), .CI(
        u2_add_111_carry[9]), .CO(u2_add_111_carry[10]), .S(u2_N27) );
  FA_X1 u2_add_111_U1_10 ( .A(opa_r[62]), .B(opb_r[62]), .CI(
        u2_add_111_carry[10]), .CO(u2_N29), .S(u2_N28) );
  INV_X4 u2_sub_111_U15 ( .A(opb_r[52]), .ZN(u2_sub_111_n13) );
  INV_X4 u2_sub_111_U14 ( .A(opb_r[53]), .ZN(u2_sub_111_n12) );
  INV_X4 u2_sub_111_U13 ( .A(opb_r[54]), .ZN(u2_sub_111_n11) );
  INV_X4 u2_sub_111_U12 ( .A(opb_r[55]), .ZN(u2_sub_111_n10) );
  INV_X4 u2_sub_111_U11 ( .A(opb_r[56]), .ZN(u2_sub_111_n9) );
  INV_X4 u2_sub_111_U10 ( .A(opb_r[57]), .ZN(u2_sub_111_n8) );
  INV_X4 u2_sub_111_U9 ( .A(opb_r[58]), .ZN(u2_sub_111_n7) );
  INV_X4 u2_sub_111_U8 ( .A(opb_r[59]), .ZN(u2_sub_111_n6) );
  INV_X4 u2_sub_111_U7 ( .A(opb_r[60]), .ZN(u2_sub_111_n5) );
  INV_X4 u2_sub_111_U6 ( .A(opb_r[61]), .ZN(u2_sub_111_n4) );
  INV_X4 u2_sub_111_U5 ( .A(opb_r[62]), .ZN(u2_sub_111_n3) );
  INV_X4 u2_sub_111_U4 ( .A(u2_sub_111_carry[11]), .ZN(u2_N17) );
  INV_X4 u2_sub_111_U3 ( .A(opa_r[52]), .ZN(u2_sub_111_n1) );
  XNOR2_X2 u2_sub_111_U2 ( .A(u2_sub_111_n13), .B(opa_r[52]), .ZN(u2_N6) );
  NAND2_X2 u2_sub_111_U1 ( .A1(opb_r[52]), .A2(u2_sub_111_n1), .ZN(
        u2_sub_111_carry[1]) );
  FA_X1 u2_sub_111_U2_1 ( .A(opa_r[53]), .B(u2_sub_111_n12), .CI(
        u2_sub_111_carry[1]), .CO(u2_sub_111_carry[2]), .S(u2_N7) );
  FA_X1 u2_sub_111_U2_2 ( .A(opa_r[54]), .B(u2_sub_111_n11), .CI(
        u2_sub_111_carry[2]), .CO(u2_sub_111_carry[3]), .S(u2_N8) );
  FA_X1 u2_sub_111_U2_3 ( .A(opa_r[55]), .B(u2_sub_111_n10), .CI(
        u2_sub_111_carry[3]), .CO(u2_sub_111_carry[4]), .S(u2_N9) );
  FA_X1 u2_sub_111_U2_4 ( .A(opa_r[56]), .B(u2_sub_111_n9), .CI(
        u2_sub_111_carry[4]), .CO(u2_sub_111_carry[5]), .S(u2_N10) );
  FA_X1 u2_sub_111_U2_5 ( .A(opa_r[57]), .B(u2_sub_111_n8), .CI(
        u2_sub_111_carry[5]), .CO(u2_sub_111_carry[6]), .S(u2_N11) );
  FA_X1 u2_sub_111_U2_6 ( .A(opa_r[58]), .B(u2_sub_111_n7), .CI(
        u2_sub_111_carry[6]), .CO(u2_sub_111_carry[7]), .S(u2_N12) );
  FA_X1 u2_sub_111_U2_7 ( .A(opa_r[59]), .B(u2_sub_111_n6), .CI(
        u2_sub_111_carry[7]), .CO(u2_sub_111_carry[8]), .S(u2_N13) );
  FA_X1 u2_sub_111_U2_8 ( .A(opa_r[60]), .B(u2_sub_111_n5), .CI(
        u2_sub_111_carry[8]), .CO(u2_sub_111_carry[9]), .S(u2_N14) );
  FA_X1 u2_sub_111_U2_9 ( .A(opa_r[61]), .B(u2_sub_111_n4), .CI(
        u2_sub_111_carry[9]), .CO(u2_sub_111_carry[10]), .S(u2_N15) );
  FA_X1 u2_sub_111_U2_10 ( .A(opa_r[62]), .B(u2_sub_111_n3), .CI(
        u2_sub_111_carry[10]), .CO(u2_sub_111_carry[11]), .S(u2_N16) );
  NOR2_X1 u1_gt_226_U168 ( .A1(n6227), .A2(u1_gt_226_n55), .ZN(u1_gt_226_n112)
         );
  NOR2_X1 u1_gt_226_U167 ( .A1(u1_gt_226_n2), .A2(n6172), .ZN(u1_gt_226_n167)
         );
  AOI21_X1 u1_gt_226_U166 ( .B1(u1_gt_226_n167), .B2(u1_gt_226_n90), .A(n6262), 
        .ZN(u1_gt_226_n166) );
  AOI221_X1 u1_gt_226_U165 ( .B1(n6211), .B2(u1_gt_226_n39), .C1(n6263), .C2(
        u1_gt_226_n1), .A(u1_gt_226_n166), .ZN(u1_gt_226_n165) );
  AOI221_X1 u1_gt_226_U164 ( .B1(n6238), .B2(u1_gt_226_n67), .C1(n6210), .C2(
        u1_gt_226_n40), .A(u1_gt_226_n165), .ZN(u1_gt_226_n164) );
  AOI221_X1 u1_gt_226_U163 ( .B1(n6183), .B2(u1_gt_226_n11), .C1(n6239), .C2(
        u1_gt_226_n66), .A(u1_gt_226_n164), .ZN(u1_gt_226_n163) );
  AOI221_X1 u1_gt_226_U162 ( .B1(n6268), .B2(u1_gt_226_n96), .C1(n6182), .C2(
        u1_gt_226_n12), .A(u1_gt_226_n163), .ZN(u1_gt_226_n162) );
  AOI221_X1 u1_gt_226_U161 ( .B1(n6215), .B2(u1_gt_226_n43), .C1(n6269), .C2(
        u1_gt_226_n95), .A(u1_gt_226_n162), .ZN(u1_gt_226_n161) );
  AOI221_X1 u1_gt_226_U160 ( .B1(n6242), .B2(u1_gt_226_n71), .C1(n6214), .C2(
        u1_gt_226_n44), .A(u1_gt_226_n161), .ZN(u1_gt_226_n160) );
  AOI221_X1 u1_gt_226_U159 ( .B1(n6187), .B2(u1_gt_226_n15), .C1(n6243), .C2(
        u1_gt_226_n70), .A(u1_gt_226_n160), .ZN(u1_gt_226_n159) );
  AOI221_X1 u1_gt_226_U158 ( .B1(n6272), .B2(u1_gt_226_n100), .C1(n6186), .C2(
        u1_gt_226_n16), .A(u1_gt_226_n159), .ZN(u1_gt_226_n158) );
  AOI221_X1 u1_gt_226_U157 ( .B1(n6273), .B2(u1_gt_226_n99), .C1(n6201), .C2(
        u1_gt_226_n29), .A(u1_gt_226_n158), .ZN(u1_gt_226_n157) );
  AOI221_X1 u1_gt_226_U156 ( .B1(n6228), .B2(u1_gt_226_n57), .C1(n6200), .C2(
        u1_gt_226_n30), .A(u1_gt_226_n157), .ZN(u1_gt_226_n156) );
  AOI221_X1 u1_gt_226_U155 ( .B1(n6177), .B2(u1_gt_226_n5), .C1(n6229), .C2(
        u1_gt_226_n56), .A(u1_gt_226_n156), .ZN(u1_gt_226_n155) );
  AOI221_X1 u1_gt_226_U154 ( .B1(n6256), .B2(u1_gt_226_n85), .C1(n6176), .C2(
        u1_gt_226_n6), .A(u1_gt_226_n155), .ZN(u1_gt_226_n154) );
  AOI221_X1 u1_gt_226_U153 ( .B1(n6205), .B2(u1_gt_226_n33), .C1(n6257), .C2(
        u1_gt_226_n84), .A(u1_gt_226_n154), .ZN(u1_gt_226_n153) );
  AOI221_X1 u1_gt_226_U152 ( .B1(n6232), .B2(u1_gt_226_n61), .C1(n6204), .C2(
        u1_gt_226_n34), .A(u1_gt_226_n153), .ZN(u1_gt_226_n152) );
  AOI221_X1 u1_gt_226_U151 ( .B1(n6175), .B2(u1_gt_226_n3), .C1(n6233), .C2(
        u1_gt_226_n60), .A(u1_gt_226_n152), .ZN(u1_gt_226_n151) );
  AOI221_X1 u1_gt_226_U150 ( .B1(n6260), .B2(u1_gt_226_n89), .C1(n6174), .C2(
        u1_gt_226_n4), .A(u1_gt_226_n151), .ZN(u1_gt_226_n150) );
  AOI221_X1 u1_gt_226_U149 ( .B1(n6209), .B2(u1_gt_226_n37), .C1(n6261), .C2(
        u1_gt_226_n88), .A(u1_gt_226_n150), .ZN(u1_gt_226_n149) );
  AOI221_X1 u1_gt_226_U148 ( .B1(n6236), .B2(u1_gt_226_n65), .C1(n6208), .C2(
        u1_gt_226_n38), .A(u1_gt_226_n149), .ZN(u1_gt_226_n148) );
  AOI221_X1 u1_gt_226_U147 ( .B1(n6181), .B2(u1_gt_226_n9), .C1(n6237), .C2(
        u1_gt_226_n64), .A(u1_gt_226_n148), .ZN(u1_gt_226_n147) );
  AOI221_X1 u1_gt_226_U146 ( .B1(n6266), .B2(u1_gt_226_n94), .C1(n6180), .C2(
        u1_gt_226_n10), .A(u1_gt_226_n147), .ZN(u1_gt_226_n146) );
  AOI221_X1 u1_gt_226_U145 ( .B1(n6213), .B2(u1_gt_226_n41), .C1(n6267), .C2(
        u1_gt_226_n93), .A(u1_gt_226_n146), .ZN(u1_gt_226_n145) );
  AOI221_X1 u1_gt_226_U144 ( .B1(n6240), .B2(u1_gt_226_n69), .C1(n6212), .C2(
        u1_gt_226_n42), .A(u1_gt_226_n145), .ZN(u1_gt_226_n144) );
  AOI221_X1 u1_gt_226_U143 ( .B1(n6185), .B2(u1_gt_226_n13), .C1(n6241), .C2(
        u1_gt_226_n68), .A(u1_gt_226_n144), .ZN(u1_gt_226_n143) );
  AOI221_X1 u1_gt_226_U142 ( .B1(n6270), .B2(u1_gt_226_n98), .C1(n6184), .C2(
        u1_gt_226_n14), .A(u1_gt_226_n143), .ZN(u1_gt_226_n142) );
  AOI221_X1 u1_gt_226_U141 ( .B1(n6203), .B2(u1_gt_226_n31), .C1(n6271), .C2(
        u1_gt_226_n97), .A(u1_gt_226_n142), .ZN(u1_gt_226_n141) );
  AOI221_X1 u1_gt_226_U140 ( .B1(n6230), .B2(u1_gt_226_n59), .C1(n6202), .C2(
        u1_gt_226_n32), .A(u1_gt_226_n141), .ZN(u1_gt_226_n140) );
  AOI221_X1 u1_gt_226_U139 ( .B1(n6179), .B2(u1_gt_226_n7), .C1(n6231), .C2(
        u1_gt_226_n58), .A(u1_gt_226_n140), .ZN(u1_gt_226_n139) );
  AOI221_X1 u1_gt_226_U138 ( .B1(n6258), .B2(u1_gt_226_n87), .C1(n6178), .C2(
        u1_gt_226_n8), .A(u1_gt_226_n139), .ZN(u1_gt_226_n138) );
  AOI221_X1 u1_gt_226_U137 ( .B1(n6207), .B2(u1_gt_226_n35), .C1(n6259), .C2(
        u1_gt_226_n86), .A(u1_gt_226_n138), .ZN(u1_gt_226_n137) );
  AOI221_X1 u1_gt_226_U136 ( .B1(n6234), .B2(u1_gt_226_n63), .C1(n6206), .C2(
        u1_gt_226_n36), .A(u1_gt_226_n137), .ZN(u1_gt_226_n136) );
  AOI221_X1 u1_gt_226_U135 ( .B1(n6189), .B2(u1_gt_226_n17), .C1(n6235), .C2(
        u1_gt_226_n62), .A(u1_gt_226_n136), .ZN(u1_gt_226_n135) );
  AOI221_X1 u1_gt_226_U134 ( .B1(n6264), .B2(u1_gt_226_n92), .C1(n6188), .C2(
        u1_gt_226_n18), .A(u1_gt_226_n135), .ZN(u1_gt_226_n134) );
  AOI221_X1 u1_gt_226_U133 ( .B1(n6217), .B2(u1_gt_226_n45), .C1(n6265), .C2(
        u1_gt_226_n91), .A(u1_gt_226_n134), .ZN(u1_gt_226_n133) );
  AOI221_X1 u1_gt_226_U132 ( .B1(n6244), .B2(u1_gt_226_n73), .C1(n6216), .C2(
        u1_gt_226_n46), .A(u1_gt_226_n133), .ZN(u1_gt_226_n132) );
  AOI221_X1 u1_gt_226_U131 ( .B1(n6191), .B2(u1_gt_226_n19), .C1(n6245), .C2(
        u1_gt_226_n72), .A(u1_gt_226_n132), .ZN(u1_gt_226_n131) );
  AOI221_X1 u1_gt_226_U130 ( .B1(n6274), .B2(u1_gt_226_n102), .C1(n6190), .C2(
        u1_gt_226_n20), .A(u1_gt_226_n131), .ZN(u1_gt_226_n130) );
  AOI221_X1 u1_gt_226_U129 ( .B1(n6219), .B2(u1_gt_226_n47), .C1(n6275), .C2(
        u1_gt_226_n101), .A(u1_gt_226_n130), .ZN(u1_gt_226_n129) );
  AOI221_X1 u1_gt_226_U128 ( .B1(n6246), .B2(u1_gt_226_n75), .C1(n6218), .C2(
        u1_gt_226_n48), .A(u1_gt_226_n129), .ZN(u1_gt_226_n128) );
  AOI221_X1 u1_gt_226_U127 ( .B1(n6195), .B2(u1_gt_226_n23), .C1(n6247), .C2(
        u1_gt_226_n74), .A(u1_gt_226_n128), .ZN(u1_gt_226_n127) );
  AOI221_X1 u1_gt_226_U126 ( .B1(n6276), .B2(u1_gt_226_n104), .C1(n6194), .C2(
        u1_gt_226_n24), .A(u1_gt_226_n127), .ZN(u1_gt_226_n126) );
  AOI221_X1 u1_gt_226_U125 ( .B1(n6221), .B2(u1_gt_226_n49), .C1(n6277), .C2(
        u1_gt_226_n103), .A(u1_gt_226_n126), .ZN(u1_gt_226_n125) );
  AOI221_X1 u1_gt_226_U124 ( .B1(n6248), .B2(u1_gt_226_n77), .C1(n6220), .C2(
        u1_gt_226_n50), .A(u1_gt_226_n125), .ZN(u1_gt_226_n124) );
  AOI221_X1 u1_gt_226_U123 ( .B1(n6193), .B2(u1_gt_226_n21), .C1(n6249), .C2(
        u1_gt_226_n76), .A(u1_gt_226_n124), .ZN(u1_gt_226_n123) );
  AOI221_X1 u1_gt_226_U122 ( .B1(n6278), .B2(u1_gt_226_n106), .C1(n6192), .C2(
        u1_gt_226_n22), .A(u1_gt_226_n123), .ZN(u1_gt_226_n122) );
  AOI221_X1 u1_gt_226_U121 ( .B1(n6223), .B2(u1_gt_226_n51), .C1(n6279), .C2(
        u1_gt_226_n105), .A(u1_gt_226_n122), .ZN(u1_gt_226_n121) );
  AOI221_X1 u1_gt_226_U120 ( .B1(n6250), .B2(u1_gt_226_n79), .C1(n6222), .C2(
        u1_gt_226_n52), .A(u1_gt_226_n121), .ZN(u1_gt_226_n120) );
  AOI221_X1 u1_gt_226_U119 ( .B1(n6197), .B2(u1_gt_226_n25), .C1(n6251), .C2(
        u1_gt_226_n78), .A(u1_gt_226_n120), .ZN(u1_gt_226_n119) );
  AOI221_X1 u1_gt_226_U118 ( .B1(n6280), .B2(u1_gt_226_n108), .C1(n6196), .C2(
        u1_gt_226_n26), .A(u1_gt_226_n119), .ZN(u1_gt_226_n118) );
  AOI221_X1 u1_gt_226_U117 ( .B1(n6225), .B2(u1_gt_226_n53), .C1(n6281), .C2(
        u1_gt_226_n107), .A(u1_gt_226_n118), .ZN(u1_gt_226_n117) );
  AOI221_X1 u1_gt_226_U116 ( .B1(n6252), .B2(u1_gt_226_n81), .C1(n6224), .C2(
        u1_gt_226_n54), .A(u1_gt_226_n117), .ZN(u1_gt_226_n116) );
  AOI221_X1 u1_gt_226_U115 ( .B1(n6199), .B2(u1_gt_226_n27), .C1(n6253), .C2(
        u1_gt_226_n80), .A(u1_gt_226_n116), .ZN(u1_gt_226_n115) );
  AOI221_X1 u1_gt_226_U114 ( .B1(n6282), .B2(u1_gt_226_n110), .C1(n6198), .C2(
        u1_gt_226_n28), .A(u1_gt_226_n115), .ZN(u1_gt_226_n114) );
  AOI221_X1 u1_gt_226_U113 ( .B1(n6227), .B2(u1_gt_226_n55), .C1(n6283), .C2(
        u1_gt_226_n109), .A(u1_gt_226_n114), .ZN(u1_gt_226_n113) );
  OAI22_X1 u1_gt_226_U112 ( .A1(u1_gt_226_n112), .A2(u1_gt_226_n113), .B1(
        n6254), .B2(u1_gt_226_n83), .ZN(u1_gt_226_n111) );
  OAI21_X1 u1_gt_226_U111 ( .B1(n6255), .B2(u1_gt_226_n82), .A(u1_gt_226_n111), 
        .ZN(u1_fractb_lt_fracta) );
  INV_X4 u1_gt_226_U110 ( .A(n6283), .ZN(u1_gt_226_n110) );
  INV_X4 u1_gt_226_U109 ( .A(n6282), .ZN(u1_gt_226_n109) );
  INV_X4 u1_gt_226_U108 ( .A(n6281), .ZN(u1_gt_226_n108) );
  INV_X4 u1_gt_226_U107 ( .A(n6280), .ZN(u1_gt_226_n107) );
  INV_X4 u1_gt_226_U106 ( .A(n6279), .ZN(u1_gt_226_n106) );
  INV_X4 u1_gt_226_U105 ( .A(n6278), .ZN(u1_gt_226_n105) );
  INV_X4 u1_gt_226_U104 ( .A(n6277), .ZN(u1_gt_226_n104) );
  INV_X4 u1_gt_226_U103 ( .A(n6276), .ZN(u1_gt_226_n103) );
  INV_X4 u1_gt_226_U102 ( .A(n6275), .ZN(u1_gt_226_n102) );
  INV_X4 u1_gt_226_U101 ( .A(n6274), .ZN(u1_gt_226_n101) );
  INV_X4 u1_gt_226_U100 ( .A(n6273), .ZN(u1_gt_226_n100) );
  INV_X4 u1_gt_226_U99 ( .A(n6272), .ZN(u1_gt_226_n99) );
  INV_X4 u1_gt_226_U98 ( .A(n6271), .ZN(u1_gt_226_n98) );
  INV_X4 u1_gt_226_U97 ( .A(n6270), .ZN(u1_gt_226_n97) );
  INV_X4 u1_gt_226_U96 ( .A(n6269), .ZN(u1_gt_226_n96) );
  INV_X4 u1_gt_226_U95 ( .A(n6268), .ZN(u1_gt_226_n95) );
  INV_X4 u1_gt_226_U94 ( .A(n6267), .ZN(u1_gt_226_n94) );
  INV_X4 u1_gt_226_U93 ( .A(n6266), .ZN(u1_gt_226_n93) );
  INV_X4 u1_gt_226_U92 ( .A(n6265), .ZN(u1_gt_226_n92) );
  INV_X4 u1_gt_226_U91 ( .A(n6264), .ZN(u1_gt_226_n91) );
  INV_X4 u1_gt_226_U90 ( .A(n6263), .ZN(u1_gt_226_n90) );
  INV_X4 u1_gt_226_U89 ( .A(n6261), .ZN(u1_gt_226_n89) );
  INV_X4 u1_gt_226_U88 ( .A(n6260), .ZN(u1_gt_226_n88) );
  INV_X4 u1_gt_226_U87 ( .A(n6259), .ZN(u1_gt_226_n87) );
  INV_X4 u1_gt_226_U86 ( .A(n6258), .ZN(u1_gt_226_n86) );
  INV_X4 u1_gt_226_U85 ( .A(n6257), .ZN(u1_gt_226_n85) );
  INV_X4 u1_gt_226_U84 ( .A(n6256), .ZN(u1_gt_226_n84) );
  INV_X4 u1_gt_226_U83 ( .A(n6255), .ZN(u1_gt_226_n83) );
  INV_X4 u1_gt_226_U82 ( .A(n6254), .ZN(u1_gt_226_n82) );
  INV_X4 u1_gt_226_U81 ( .A(n6253), .ZN(u1_gt_226_n81) );
  INV_X4 u1_gt_226_U80 ( .A(n6252), .ZN(u1_gt_226_n80) );
  INV_X4 u1_gt_226_U79 ( .A(n6251), .ZN(u1_gt_226_n79) );
  INV_X4 u1_gt_226_U78 ( .A(n6250), .ZN(u1_gt_226_n78) );
  INV_X4 u1_gt_226_U77 ( .A(n6249), .ZN(u1_gt_226_n77) );
  INV_X4 u1_gt_226_U76 ( .A(n6248), .ZN(u1_gt_226_n76) );
  INV_X4 u1_gt_226_U75 ( .A(n6247), .ZN(u1_gt_226_n75) );
  INV_X4 u1_gt_226_U74 ( .A(n6246), .ZN(u1_gt_226_n74) );
  INV_X4 u1_gt_226_U73 ( .A(n6245), .ZN(u1_gt_226_n73) );
  INV_X4 u1_gt_226_U72 ( .A(n6244), .ZN(u1_gt_226_n72) );
  INV_X4 u1_gt_226_U71 ( .A(n6243), .ZN(u1_gt_226_n71) );
  INV_X4 u1_gt_226_U70 ( .A(n6242), .ZN(u1_gt_226_n70) );
  INV_X4 u1_gt_226_U69 ( .A(n6241), .ZN(u1_gt_226_n69) );
  INV_X4 u1_gt_226_U68 ( .A(n6240), .ZN(u1_gt_226_n68) );
  INV_X4 u1_gt_226_U67 ( .A(n6239), .ZN(u1_gt_226_n67) );
  INV_X4 u1_gt_226_U66 ( .A(n6238), .ZN(u1_gt_226_n66) );
  INV_X4 u1_gt_226_U65 ( .A(n6237), .ZN(u1_gt_226_n65) );
  INV_X4 u1_gt_226_U64 ( .A(n6236), .ZN(u1_gt_226_n64) );
  INV_X4 u1_gt_226_U63 ( .A(n6235), .ZN(u1_gt_226_n63) );
  INV_X4 u1_gt_226_U62 ( .A(n6234), .ZN(u1_gt_226_n62) );
  INV_X4 u1_gt_226_U61 ( .A(n6233), .ZN(u1_gt_226_n61) );
  INV_X4 u1_gt_226_U60 ( .A(n6232), .ZN(u1_gt_226_n60) );
  INV_X4 u1_gt_226_U59 ( .A(n6231), .ZN(u1_gt_226_n59) );
  INV_X4 u1_gt_226_U58 ( .A(n6230), .ZN(u1_gt_226_n58) );
  INV_X4 u1_gt_226_U57 ( .A(n6229), .ZN(u1_gt_226_n57) );
  INV_X4 u1_gt_226_U56 ( .A(n6228), .ZN(u1_gt_226_n56) );
  INV_X4 u1_gt_226_U55 ( .A(n6226), .ZN(u1_gt_226_n55) );
  INV_X4 u1_gt_226_U54 ( .A(n6225), .ZN(u1_gt_226_n54) );
  INV_X4 u1_gt_226_U53 ( .A(n6224), .ZN(u1_gt_226_n53) );
  INV_X4 u1_gt_226_U52 ( .A(n6223), .ZN(u1_gt_226_n52) );
  INV_X4 u1_gt_226_U51 ( .A(n6222), .ZN(u1_gt_226_n51) );
  INV_X4 u1_gt_226_U50 ( .A(n6221), .ZN(u1_gt_226_n50) );
  INV_X4 u1_gt_226_U49 ( .A(n6220), .ZN(u1_gt_226_n49) );
  INV_X4 u1_gt_226_U48 ( .A(n6219), .ZN(u1_gt_226_n48) );
  INV_X4 u1_gt_226_U47 ( .A(n6218), .ZN(u1_gt_226_n47) );
  INV_X4 u1_gt_226_U46 ( .A(n6217), .ZN(u1_gt_226_n46) );
  INV_X4 u1_gt_226_U45 ( .A(n6216), .ZN(u1_gt_226_n45) );
  INV_X4 u1_gt_226_U44 ( .A(n6215), .ZN(u1_gt_226_n44) );
  INV_X4 u1_gt_226_U43 ( .A(n6214), .ZN(u1_gt_226_n43) );
  INV_X4 u1_gt_226_U42 ( .A(n6213), .ZN(u1_gt_226_n42) );
  INV_X4 u1_gt_226_U41 ( .A(n6212), .ZN(u1_gt_226_n41) );
  INV_X4 u1_gt_226_U40 ( .A(n6211), .ZN(u1_gt_226_n40) );
  INV_X4 u1_gt_226_U39 ( .A(n6210), .ZN(u1_gt_226_n39) );
  INV_X4 u1_gt_226_U38 ( .A(n6209), .ZN(u1_gt_226_n38) );
  INV_X4 u1_gt_226_U37 ( .A(n6208), .ZN(u1_gt_226_n37) );
  INV_X4 u1_gt_226_U36 ( .A(n6207), .ZN(u1_gt_226_n36) );
  INV_X4 u1_gt_226_U35 ( .A(n6206), .ZN(u1_gt_226_n35) );
  INV_X4 u1_gt_226_U34 ( .A(n6205), .ZN(u1_gt_226_n34) );
  INV_X4 u1_gt_226_U33 ( .A(n6204), .ZN(u1_gt_226_n33) );
  INV_X4 u1_gt_226_U32 ( .A(n6203), .ZN(u1_gt_226_n32) );
  INV_X4 u1_gt_226_U31 ( .A(n6202), .ZN(u1_gt_226_n31) );
  INV_X4 u1_gt_226_U30 ( .A(n6201), .ZN(u1_gt_226_n30) );
  INV_X4 u1_gt_226_U29 ( .A(n6200), .ZN(u1_gt_226_n29) );
  INV_X4 u1_gt_226_U28 ( .A(n6199), .ZN(u1_gt_226_n28) );
  INV_X4 u1_gt_226_U27 ( .A(n6198), .ZN(u1_gt_226_n27) );
  INV_X4 u1_gt_226_U26 ( .A(n6197), .ZN(u1_gt_226_n26) );
  INV_X4 u1_gt_226_U25 ( .A(n6196), .ZN(u1_gt_226_n25) );
  INV_X4 u1_gt_226_U24 ( .A(n6195), .ZN(u1_gt_226_n24) );
  INV_X4 u1_gt_226_U23 ( .A(n6194), .ZN(u1_gt_226_n23) );
  INV_X4 u1_gt_226_U22 ( .A(n6193), .ZN(u1_gt_226_n22) );
  INV_X4 u1_gt_226_U21 ( .A(n6192), .ZN(u1_gt_226_n21) );
  INV_X4 u1_gt_226_U20 ( .A(n6191), .ZN(u1_gt_226_n20) );
  INV_X4 u1_gt_226_U19 ( .A(n6190), .ZN(u1_gt_226_n19) );
  INV_X4 u1_gt_226_U18 ( .A(n6189), .ZN(u1_gt_226_n18) );
  INV_X4 u1_gt_226_U17 ( .A(n6188), .ZN(u1_gt_226_n17) );
  INV_X4 u1_gt_226_U16 ( .A(n6187), .ZN(u1_gt_226_n16) );
  INV_X4 u1_gt_226_U15 ( .A(n6186), .ZN(u1_gt_226_n15) );
  INV_X4 u1_gt_226_U14 ( .A(n6185), .ZN(u1_gt_226_n14) );
  INV_X4 u1_gt_226_U13 ( .A(n6184), .ZN(u1_gt_226_n13) );
  INV_X4 u1_gt_226_U12 ( .A(n6183), .ZN(u1_gt_226_n12) );
  INV_X4 u1_gt_226_U11 ( .A(n6182), .ZN(u1_gt_226_n11) );
  INV_X4 u1_gt_226_U10 ( .A(n6181), .ZN(u1_gt_226_n10) );
  INV_X4 u1_gt_226_U9 ( .A(n6180), .ZN(u1_gt_226_n9) );
  INV_X4 u1_gt_226_U8 ( .A(n6179), .ZN(u1_gt_226_n8) );
  INV_X4 u1_gt_226_U7 ( .A(n6178), .ZN(u1_gt_226_n7) );
  INV_X4 u1_gt_226_U6 ( .A(n6177), .ZN(u1_gt_226_n6) );
  INV_X4 u1_gt_226_U5 ( .A(n6176), .ZN(u1_gt_226_n5) );
  INV_X4 u1_gt_226_U4 ( .A(n6175), .ZN(u1_gt_226_n4) );
  INV_X4 u1_gt_226_U3 ( .A(n6174), .ZN(u1_gt_226_n3) );
  INV_X4 u1_gt_226_U2 ( .A(n6173), .ZN(u1_gt_226_n2) );
  INV_X4 u1_gt_226_U1 ( .A(u1_gt_226_n167), .ZN(u1_gt_226_n1) );
  NOR2_X1 u1_srl_148_U418 ( .A1(u1_srl_148_n97), .A2(n6302), .ZN(
        u1_srl_148_n162) );
  AND2_X1 u1_srl_148_U417 ( .A1(n6285), .A2(u1_exp_diff_sft_0_), .ZN(
        u1_srl_148_n197) );
  NOR2_X1 u1_srl_148_U416 ( .A1(u1_exp_diff_sft_0_), .A2(n6285), .ZN(
        u1_srl_148_n198) );
  AOI22_X1 u1_srl_148_U415 ( .A1(n4174), .A2(u1_srl_148_n14), .B1(n4177), .B2(
        u1_srl_148_n198), .ZN(u1_srl_148_n360) );
  OAI221_X1 u1_srl_148_U414 ( .B1(u1_srl_148_n5), .B2(u1_srl_148_n110), .C1(
        u1_srl_148_n2), .C2(u1_srl_148_n109), .A(u1_srl_148_n360), .ZN(
        u1_srl_148_n242) );
  AOI22_X1 u1_srl_148_U413 ( .A1(n6332), .A2(u1_srl_148_n197), .B1(
        u1_srl_148_n198), .B2(n4181), .ZN(u1_srl_148_n359) );
  OAI221_X1 u1_srl_148_U412 ( .B1(u1_srl_148_n5), .B2(u1_srl_148_n114), .C1(
        u1_srl_148_n2), .C2(u1_srl_148_n113), .A(u1_srl_148_n359), .ZN(
        u1_srl_148_n243) );
  AOI22_X1 u1_srl_148_U411 ( .A1(u1_srl_148_n14), .A2(n6333), .B1(n4185), .B2(
        u1_srl_148_n15), .ZN(u1_srl_148_n358) );
  OAI221_X1 u1_srl_148_U410 ( .B1(u1_srl_148_n6), .B2(u1_srl_148_n118), .C1(
        u1_srl_148_n117), .C2(u1_srl_148_n2), .A(u1_srl_148_n358), .ZN(
        u1_srl_148_n152) );
  NOR2_X1 u1_srl_148_U409 ( .A1(n6293), .A2(n6301), .ZN(u1_srl_148_n211) );
  AOI22_X1 u1_srl_148_U408 ( .A1(n4186), .A2(u1_srl_148_n14), .B1(n6338), .B2(
        u1_srl_148_n15), .ZN(u1_srl_148_n357) );
  OAI221_X1 u1_srl_148_U407 ( .B1(u1_srl_148_n6), .B2(u1_srl_148_n122), .C1(
        u1_srl_148_n2), .C2(u1_srl_148_n121), .A(u1_srl_148_n357), .ZN(
        u1_srl_148_n153) );
  AOI22_X1 u1_srl_148_U406 ( .A1(u1_srl_148_n9), .A2(u1_srl_148_n152), .B1(
        u1_srl_148_n211), .B2(u1_srl_148_n153), .ZN(u1_srl_148_n356) );
  AOI221_X1 u1_srl_148_U405 ( .B1(u1_srl_148_n242), .B2(u1_srl_148_n237), .C1(
        u1_srl_148_n243), .C2(u1_srl_148_n195), .A(u1_srl_148_n22), .ZN(
        u1_srl_148_n289) );
  AOI22_X1 u1_srl_148_U404 ( .A1(n6345), .A2(u1_srl_148_n197), .B1(n6347), 
        .B2(u1_srl_148_n15), .ZN(u1_srl_148_n355) );
  OAI221_X1 u1_srl_148_U403 ( .B1(u1_srl_148_n6), .B2(u1_srl_148_n104), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n133), .A(u1_srl_148_n355), .ZN(
        u1_srl_148_n183) );
  AOI22_X1 u1_srl_148_U402 ( .A1(u1_adj_op_36_), .A2(u1_srl_148_n14), .B1(
        n6330), .B2(u1_srl_148_n15), .ZN(u1_srl_148_n354) );
  OAI221_X1 u1_srl_148_U401 ( .B1(u1_srl_148_n6), .B2(u1_srl_148_n105), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n100), .A(u1_srl_148_n354), .ZN(
        u1_srl_148_n245) );
  AOI22_X1 u1_srl_148_U400 ( .A1(n4173), .A2(u1_srl_148_n14), .B1(
        u1_adj_op_29_), .B2(u1_srl_148_n15), .ZN(u1_srl_148_n353) );
  OAI221_X1 u1_srl_148_U399 ( .B1(u1_srl_148_n6), .B2(u1_srl_148_n102), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n101), .A(u1_srl_148_n353), .ZN(
        u1_srl_148_n246) );
  AOI22_X1 u1_srl_148_U398 ( .A1(n6324), .A2(u1_srl_148_n197), .B1(n6326), 
        .B2(u1_srl_148_n198), .ZN(u1_srl_148_n352) );
  AOI221_X1 u1_srl_148_U397 ( .B1(u1_srl_148_n224), .B2(n4166), .C1(
        u1_srl_148_n12), .C2(n6325), .A(u1_srl_148_n30), .ZN(u1_srl_148_n270)
         );
  AOI22_X1 u1_srl_148_U396 ( .A1(n6327), .A2(u1_srl_148_n197), .B1(n6304), 
        .B2(u1_srl_148_n198), .ZN(u1_srl_148_n351) );
  AOI221_X1 u1_srl_148_U395 ( .B1(u1_srl_148_n224), .B2(n4170), .C1(
        u1_srl_148_n12), .C2(n6328), .A(u1_srl_148_n32), .ZN(u1_srl_148_n312)
         );
  OAI22_X1 u1_srl_148_U394 ( .A1(u1_srl_148_n91), .A2(u1_srl_148_n270), .B1(
        u1_srl_148_n4), .B2(u1_srl_148_n312), .ZN(u1_srl_148_n350) );
  AOI221_X1 u1_srl_148_U393 ( .B1(u1_srl_148_n245), .B2(u1_srl_148_n10), .C1(
        u1_srl_148_n246), .C2(u1_srl_148_n211), .A(u1_srl_148_n350), .ZN(
        u1_srl_148_n215) );
  AOI222_X1 u1_srl_148_U392 ( .A1(u1_srl_148_n162), .A2(u1_srl_148_n19), .B1(
        u1_srl_148_n138), .B2(u1_srl_148_n183), .C1(u1_srl_148_n144), .C2(
        u1_srl_148_n23), .ZN(u1_srl_148_n342) );
  NAND2_X1 u1_srl_148_U391 ( .A1(n6303), .A2(n6302), .ZN(u1_srl_148_n223) );
  AOI22_X1 u1_srl_148_U390 ( .A1(n4160), .A2(u1_srl_148_n14), .B1(n6323), .B2(
        u1_srl_148_n198), .ZN(u1_srl_148_n349) );
  AOI221_X1 u1_srl_148_U389 ( .B1(u1_srl_148_n224), .B2(n6322), .C1(
        u1_srl_148_n12), .C2(n4161), .A(u1_srl_148_n35), .ZN(u1_srl_148_n241)
         );
  AOI22_X1 u1_srl_148_U388 ( .A1(n4348), .A2(u1_srl_148_n14), .B1(n4159), .B2(
        u1_srl_148_n15), .ZN(u1_srl_148_n348) );
  AOI221_X1 u1_srl_148_U387 ( .B1(u1_srl_148_n224), .B2(n4158), .C1(
        u1_srl_148_n12), .C2(n4157), .A(u1_srl_148_n37), .ZN(u1_srl_148_n178)
         );
  AOI22_X1 u1_srl_148_U386 ( .A1(u1_srl_148_n34), .A2(u1_srl_148_n17), .B1(
        u1_srl_148_n36), .B2(u1_srl_148_n10), .ZN(u1_srl_148_n186) );
  AOI22_X1 u1_srl_148_U385 ( .A1(n6341), .A2(u1_srl_148_n14), .B1(n6344), .B2(
        u1_srl_148_n15), .ZN(u1_srl_148_n347) );
  OAI221_X1 u1_srl_148_U384 ( .B1(u1_srl_148_n6), .B2(u1_srl_148_n130), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n129), .A(u1_srl_148_n347), .ZN(
        u1_srl_148_n154) );
  AOI22_X1 u1_srl_148_U383 ( .A1(n4190), .A2(u1_srl_148_n14), .B1(n4193), .B2(
        u1_srl_148_n198), .ZN(u1_srl_148_n346) );
  OAI221_X1 u1_srl_148_U382 ( .B1(u1_srl_148_n6), .B2(u1_srl_148_n126), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n125), .A(u1_srl_148_n346), .ZN(
        u1_srl_148_n151) );
  AOI22_X1 u1_srl_148_U381 ( .A1(u1_srl_148_n154), .A2(u1_srl_148_n142), .B1(
        u1_srl_148_n151), .B2(u1_srl_148_n140), .ZN(u1_srl_148_n344) );
  NAND3_X1 u1_srl_148_U380 ( .A1(n6348), .A2(u1_srl_148_n197), .A3(
        u1_srl_148_n145), .ZN(u1_srl_148_n345) );
  OAI211_X1 u1_srl_148_U379 ( .C1(u1_srl_148_n223), .C2(u1_srl_148_n186), .A(
        u1_srl_148_n344), .B(u1_srl_148_n345), .ZN(u1_srl_148_n343) );
  NAND2_X1 u1_srl_148_U378 ( .A1(u1_srl_148_n342), .A2(u1_srl_148_n33), .ZN(
        u1_adj_op_out_sft_0_) );
  AOI22_X1 u1_srl_148_U377 ( .A1(n6307), .A2(u1_srl_148_n14), .B1(n4175), .B2(
        u1_srl_148_n15), .ZN(u1_srl_148_n341) );
  OAI221_X1 u1_srl_148_U376 ( .B1(u1_srl_148_n6), .B2(u1_srl_148_n108), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n103), .A(u1_srl_148_n341), .ZN(
        u1_srl_148_n259) );
  AOI22_X1 u1_srl_148_U375 ( .A1(n6331), .A2(u1_srl_148_n14), .B1(n4179), .B2(
        u1_srl_148_n198), .ZN(u1_srl_148_n340) );
  OAI221_X1 u1_srl_148_U374 ( .B1(u1_srl_148_n6), .B2(u1_srl_148_n112), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n111), .A(u1_srl_148_n340), .ZN(
        u1_srl_148_n255) );
  AOI22_X1 u1_srl_148_U373 ( .A1(n4170), .A2(u1_srl_148_n14), .B1(n6305), .B2(
        u1_srl_148_n15), .ZN(u1_srl_148_n339) );
  OAI221_X1 u1_srl_148_U372 ( .B1(u1_srl_148_n6), .B2(u1_srl_148_n99), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n98), .A(u1_srl_148_n339), .ZN(
        u1_srl_148_n260) );
  AOI22_X1 u1_srl_148_U371 ( .A1(n6329), .A2(u1_srl_148_n14), .B1(n6306), .B2(
        u1_srl_148_n15), .ZN(u1_srl_148_n338) );
  OAI221_X1 u1_srl_148_U370 ( .B1(u1_srl_148_n6), .B2(u1_srl_148_n107), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n106), .A(u1_srl_148_n338), .ZN(
        u1_srl_148_n258) );
  AOI22_X1 u1_srl_148_U369 ( .A1(u1_srl_148_n237), .A2(u1_srl_148_n260), .B1(
        u1_srl_148_n195), .B2(u1_srl_148_n258), .ZN(u1_srl_148_n337) );
  AOI221_X1 u1_srl_148_U368 ( .B1(u1_srl_148_n259), .B2(u1_srl_148_n10), .C1(
        u1_srl_148_n255), .C2(u1_srl_148_n211), .A(u1_srl_148_n42), .ZN(
        u1_srl_148_n231) );
  AOI22_X1 u1_srl_148_U367 ( .A1(n6322), .A2(u1_srl_148_n14), .B1(n6325), .B2(
        u1_srl_148_n15), .ZN(u1_srl_148_n336) );
  AOI221_X1 u1_srl_148_U366 ( .B1(u1_srl_148_n224), .B2(n6324), .C1(
        u1_srl_148_n12), .C2(n6323), .A(u1_srl_148_n49), .ZN(u1_srl_148_n263)
         );
  AOI22_X1 u1_srl_148_U365 ( .A1(n4166), .A2(u1_srl_148_n14), .B1(n6328), .B2(
        u1_srl_148_n15), .ZN(u1_srl_148_n335) );
  AOI221_X1 u1_srl_148_U364 ( .B1(u1_srl_148_n224), .B2(n6327), .C1(
        u1_srl_148_n12), .C2(n6326), .A(u1_srl_148_n51), .ZN(u1_srl_148_n286)
         );
  AOI22_X1 u1_srl_148_U363 ( .A1(u1_srl_148_n15), .A2(n4157), .B1(
        u1_srl_148_n224), .B2(n4348), .ZN(u1_srl_148_n176) );
  AOI22_X1 u1_srl_148_U362 ( .A1(n4158), .A2(u1_srl_148_n14), .B1(n4161), .B2(
        u1_srl_148_n15), .ZN(u1_srl_148_n334) );
  AOI221_X1 u1_srl_148_U361 ( .B1(u1_srl_148_n224), .B2(n4160), .C1(
        u1_srl_148_n12), .C2(n4159), .A(u1_srl_148_n54), .ZN(u1_srl_148_n262)
         );
  OAI22_X1 u1_srl_148_U360 ( .A1(u1_srl_148_n91), .A2(u1_srl_148_n176), .B1(
        u1_srl_148_n4), .B2(u1_srl_148_n262), .ZN(u1_srl_148_n333) );
  AOI221_X1 u1_srl_148_U359 ( .B1(u1_srl_148_n48), .B2(u1_srl_148_n10), .C1(
        u1_srl_148_n50), .C2(u1_srl_148_n211), .A(u1_srl_148_n333), .ZN(
        u1_srl_148_n190) );
  AOI22_X1 u1_srl_148_U358 ( .A1(n6340), .A2(u1_srl_148_n14), .B1(n6342), .B2(
        u1_srl_148_n15), .ZN(u1_srl_148_n332) );
  OAI221_X1 u1_srl_148_U357 ( .B1(u1_srl_148_n6), .B2(u1_srl_148_n128), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n127), .A(u1_srl_148_n332), .ZN(
        u1_srl_148_n166) );
  AOI22_X1 u1_srl_148_U356 ( .A1(u1_srl_148_n144), .A2(u1_srl_148_n46), .B1(
        u1_srl_148_n145), .B2(u1_srl_148_n166), .ZN(u1_srl_148_n327) );
  AOI22_X1 u1_srl_148_U355 ( .A1(n6337), .A2(u1_srl_148_n14), .B1(n6339), .B2(
        u1_srl_148_n15), .ZN(u1_srl_148_n331) );
  OAI221_X1 u1_srl_148_U354 ( .B1(u1_srl_148_n5), .B2(u1_srl_148_n124), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n123), .A(u1_srl_148_n331), .ZN(
        u1_srl_148_n168) );
  AOI22_X1 u1_srl_148_U353 ( .A1(n4180), .A2(u1_srl_148_n14), .B1(
        u1_srl_148_n15), .B2(n6334), .ZN(u1_srl_148_n330) );
  OAI221_X1 u1_srl_148_U352 ( .B1(u1_srl_148_n5), .B2(u1_srl_148_n116), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n115), .A(u1_srl_148_n330), .ZN(
        u1_srl_148_n256) );
  AOI22_X1 u1_srl_148_U351 ( .A1(n6335), .A2(u1_srl_148_n14), .B1(n6336), .B2(
        u1_srl_148_n15), .ZN(u1_srl_148_n329) );
  OAI221_X1 u1_srl_148_U350 ( .B1(u1_srl_148_n5), .B2(u1_srl_148_n120), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n119), .A(u1_srl_148_n329), .ZN(
        u1_srl_148_n167) );
  AOI222_X1 u1_srl_148_U349 ( .A1(u1_srl_148_n138), .A2(u1_srl_148_n168), .B1(
        u1_srl_148_n140), .B2(u1_srl_148_n256), .C1(u1_srl_148_n142), .C2(
        u1_srl_148_n167), .ZN(u1_srl_148_n328) );
  OAI211_X1 u1_srl_148_U348 ( .C1(u1_srl_148_n231), .C2(u1_srl_148_n96), .A(
        u1_srl_148_n327), .B(u1_srl_148_n328), .ZN(u1_adj_op_out_sft_10_) );
  AOI22_X1 u1_srl_148_U347 ( .A1(n6306), .A2(u1_srl_148_n14), .B1(n4174), .B2(
        u1_srl_148_n15), .ZN(u1_srl_148_n326) );
  OAI221_X1 u1_srl_148_U346 ( .B1(u1_srl_148_n5), .B2(u1_srl_148_n103), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n102), .A(u1_srl_148_n326), .ZN(
        u1_srl_148_n279) );
  AOI22_X1 u1_srl_148_U345 ( .A1(n4175), .A2(u1_srl_148_n14), .B1(n6332), .B2(
        u1_srl_148_n15), .ZN(u1_srl_148_n325) );
  OAI221_X1 u1_srl_148_U344 ( .B1(u1_srl_148_n5), .B2(u1_srl_148_n111), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n110), .A(u1_srl_148_n325), .ZN(
        u1_srl_148_n248) );
  AOI22_X1 u1_srl_148_U343 ( .A1(n6328), .A2(u1_srl_148_n14), .B1(
        u1_adj_op_36_), .B2(u1_srl_148_n15), .ZN(u1_srl_148_n324) );
  AOI221_X1 u1_srl_148_U342 ( .B1(u1_srl_148_n224), .B2(n6304), .C1(
        u1_srl_148_n12), .C2(n4170), .A(u1_srl_148_n62), .ZN(u1_srl_148_n283)
         );
  AOI22_X1 u1_srl_148_U341 ( .A1(n6305), .A2(u1_srl_148_n14), .B1(n4173), .B2(
        u1_srl_148_n15), .ZN(u1_srl_148_n323) );
  OAI221_X1 u1_srl_148_U340 ( .B1(u1_srl_148_n5), .B2(u1_srl_148_n106), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n105), .A(u1_srl_148_n323), .ZN(
        u1_srl_148_n281) );
  OAI22_X1 u1_srl_148_U339 ( .A1(u1_srl_148_n91), .A2(u1_srl_148_n283), .B1(
        u1_srl_148_n4), .B2(u1_srl_148_n63), .ZN(u1_srl_148_n322) );
  AOI221_X1 u1_srl_148_U338 ( .B1(u1_srl_148_n279), .B2(u1_srl_148_n10), .C1(
        u1_srl_148_n248), .C2(u1_srl_148_n211), .A(u1_srl_148_n322), .ZN(
        u1_srl_148_n229) );
  AOI22_X1 u1_srl_148_U337 ( .A1(n6325), .A2(u1_srl_148_n14), .B1(n6327), .B2(
        u1_srl_148_n15), .ZN(u1_srl_148_n321) );
  AOI221_X1 u1_srl_148_U336 ( .B1(u1_srl_148_n224), .B2(n6326), .C1(
        u1_srl_148_n12), .C2(n4166), .A(u1_srl_148_n66), .ZN(u1_srl_148_n254)
         );
  AOI22_X1 u1_srl_148_U335 ( .A1(n4161), .A2(u1_srl_148_n14), .B1(n6324), .B2(
        u1_srl_148_n15), .ZN(u1_srl_148_n320) );
  AOI221_X1 u1_srl_148_U334 ( .B1(u1_srl_148_n224), .B2(n6323), .C1(
        u1_srl_148_n12), .C2(n6322), .A(u1_srl_148_n68), .ZN(u1_srl_148_n253)
         );
  NAND2_X1 u1_srl_148_U333 ( .A1(n4348), .A2(u1_srl_148_n15), .ZN(
        u1_srl_148_n175) );
  AOI22_X1 u1_srl_148_U332 ( .A1(n4157), .A2(u1_srl_148_n197), .B1(n4160), 
        .B2(u1_srl_148_n15), .ZN(u1_srl_148_n319) );
  AOI221_X1 u1_srl_148_U331 ( .B1(u1_srl_148_n224), .B2(n4159), .C1(
        u1_srl_148_n12), .C2(n4158), .A(u1_srl_148_n69), .ZN(u1_srl_148_n252)
         );
  MUX2_X1 u1_srl_148_U330 ( .A(u1_srl_148_n175), .B(u1_srl_148_n252), .S(
        u1_srl_148_n92), .Z(u1_srl_148_n280) );
  OAI222_X1 u1_srl_148_U329 ( .A1(u1_srl_148_n254), .A2(u1_srl_148_n18), .B1(
        u1_srl_148_n253), .B2(u1_srl_148_n1), .C1(u1_srl_148_n280), .C2(
        u1_srl_148_n93), .ZN(u1_srl_148_n230) );
  AOI22_X1 u1_srl_148_U328 ( .A1(n6339), .A2(u1_srl_148_n14), .B1(n6341), .B2(
        u1_srl_148_n15), .ZN(u1_srl_148_n318) );
  OAI221_X1 u1_srl_148_U327 ( .B1(u1_srl_148_n5), .B2(u1_srl_148_n127), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n126), .A(u1_srl_148_n318), .ZN(
        u1_srl_148_n158) );
  AOI22_X1 u1_srl_148_U326 ( .A1(u1_srl_148_n144), .A2(u1_srl_148_n230), .B1(
        u1_srl_148_n145), .B2(u1_srl_148_n158), .ZN(u1_srl_148_n313) );
  AOI22_X1 u1_srl_148_U325 ( .A1(n6336), .A2(u1_srl_148_n14), .B1(n4190), .B2(
        u1_srl_148_n15), .ZN(u1_srl_148_n317) );
  OAI221_X1 u1_srl_148_U324 ( .B1(u1_srl_148_n5), .B2(u1_srl_148_n123), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n122), .A(u1_srl_148_n317), .ZN(
        u1_srl_148_n160) );
  AOI22_X1 u1_srl_148_U323 ( .A1(n4179), .A2(u1_srl_148_n14), .B1(
        u1_srl_148_n198), .B2(n6333), .ZN(u1_srl_148_n316) );
  OAI221_X1 u1_srl_148_U322 ( .B1(u1_srl_148_n5), .B2(u1_srl_148_n115), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n114), .A(u1_srl_148_n316), .ZN(
        u1_srl_148_n249) );
  AOI22_X1 u1_srl_148_U321 ( .A1(u1_srl_148_n197), .A2(n6334), .B1(n4186), 
        .B2(u1_srl_148_n15), .ZN(u1_srl_148_n315) );
  OAI221_X1 u1_srl_148_U320 ( .B1(u1_srl_148_n5), .B2(u1_srl_148_n119), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n118), .A(u1_srl_148_n315), .ZN(
        u1_srl_148_n159) );
  AOI222_X1 u1_srl_148_U319 ( .A1(u1_srl_148_n138), .A2(u1_srl_148_n160), .B1(
        u1_srl_148_n140), .B2(u1_srl_148_n249), .C1(u1_srl_148_n142), .C2(
        u1_srl_148_n159), .ZN(u1_srl_148_n314) );
  OAI211_X1 u1_srl_148_U318 ( .C1(u1_srl_148_n229), .C2(u1_srl_148_n96), .A(
        u1_srl_148_n313), .B(u1_srl_148_n314), .ZN(u1_adj_op_out_sft_11_) );
  AOI22_X1 u1_srl_148_U317 ( .A1(u1_srl_148_n237), .A2(u1_srl_148_n31), .B1(
        u1_srl_148_n195), .B2(u1_srl_148_n245), .ZN(u1_srl_148_n311) );
  AOI221_X1 u1_srl_148_U316 ( .B1(u1_srl_148_n246), .B2(u1_srl_148_n10), .C1(
        u1_srl_148_n242), .C2(u1_srl_148_n211), .A(u1_srl_148_n24), .ZN(
        u1_srl_148_n228) );
  AOI222_X1 u1_srl_148_U315 ( .A1(u1_srl_148_n34), .A2(u1_srl_148_n9), .B1(
        u1_srl_148_n36), .B2(u1_srl_148_n195), .C1(u1_srl_148_n29), .C2(
        u1_srl_148_n211), .ZN(u1_srl_148_n189) );
  AOI22_X1 u1_srl_148_U314 ( .A1(u1_srl_148_n144), .A2(u1_srl_148_n27), .B1(
        u1_srl_148_n145), .B2(u1_srl_148_n151), .ZN(u1_srl_148_n309) );
  AOI222_X1 u1_srl_148_U313 ( .A1(u1_srl_148_n138), .A2(u1_srl_148_n153), .B1(
        u1_srl_148_n140), .B2(u1_srl_148_n243), .C1(u1_srl_148_n142), .C2(
        u1_srl_148_n152), .ZN(u1_srl_148_n310) );
  OAI211_X1 u1_srl_148_U312 ( .C1(u1_srl_148_n228), .C2(u1_srl_148_n96), .A(
        u1_srl_148_n309), .B(u1_srl_148_n310), .ZN(u1_adj_op_out_sft_12_) );
  AOI22_X1 u1_srl_148_U311 ( .A1(n6330), .A2(u1_srl_148_n197), .B1(n6307), 
        .B2(u1_srl_148_n15), .ZN(u1_srl_148_n308) );
  OAI221_X1 u1_srl_148_U310 ( .B1(u1_srl_148_n5), .B2(u1_srl_148_n101), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n107), .A(u1_srl_148_n308), .ZN(
        u1_srl_148_n239) );
  AOI22_X1 u1_srl_148_U309 ( .A1(u1_adj_op_29_), .A2(u1_srl_148_n14), .B1(
        n6331), .B2(u1_srl_148_n15), .ZN(u1_srl_148_n307) );
  OAI221_X1 u1_srl_148_U308 ( .B1(u1_srl_148_n5), .B2(u1_srl_148_n109), .C1(
        u1_srl_148_n2), .C2(u1_srl_148_n108), .A(u1_srl_148_n307), .ZN(
        u1_srl_148_n234) );
  AOI22_X1 u1_srl_148_U307 ( .A1(n6326), .A2(u1_srl_148_n14), .B1(n4170), .B2(
        u1_srl_148_n15), .ZN(u1_srl_148_n306) );
  AOI221_X1 u1_srl_148_U306 ( .B1(u1_srl_148_n224), .B2(n6328), .C1(
        u1_srl_148_n12), .C2(n6327), .A(u1_srl_148_n80), .ZN(u1_srl_148_n267)
         );
  AOI22_X1 u1_srl_148_U305 ( .A1(n6304), .A2(u1_srl_148_n197), .B1(n6329), 
        .B2(u1_srl_148_n15), .ZN(u1_srl_148_n305) );
  OAI221_X1 u1_srl_148_U304 ( .B1(u1_srl_148_n5), .B2(u1_srl_148_n100), .C1(
        u1_srl_148_n2), .C2(u1_srl_148_n99), .A(u1_srl_148_n305), .ZN(
        u1_srl_148_n238) );
  OAI22_X1 u1_srl_148_U303 ( .A1(u1_srl_148_n91), .A2(u1_srl_148_n267), .B1(
        u1_srl_148_n4), .B2(u1_srl_148_n81), .ZN(u1_srl_148_n304) );
  AOI221_X1 u1_srl_148_U302 ( .B1(u1_srl_148_n239), .B2(u1_srl_148_n10), .C1(
        u1_srl_148_n234), .C2(u1_srl_148_n211), .A(u1_srl_148_n304), .ZN(
        u1_srl_148_n227) );
  AOI22_X1 u1_srl_148_U301 ( .A1(n4159), .A2(u1_srl_148_n197), .B1(n6322), 
        .B2(u1_srl_148_n15), .ZN(u1_srl_148_n303) );
  AOI221_X1 u1_srl_148_U300 ( .B1(u1_srl_148_n224), .B2(n4161), .C1(
        u1_srl_148_n12), .C2(n4160), .A(u1_srl_148_n85), .ZN(u1_srl_148_n233)
         );
  AOI222_X1 u1_srl_148_U299 ( .A1(u1_srl_148_n12), .A2(n4348), .B1(
        u1_srl_148_n224), .B2(n4157), .C1(u1_srl_148_n198), .C2(n4158), .ZN(
        u1_srl_148_n177) );
  AOI22_X1 u1_srl_148_U298 ( .A1(n6323), .A2(u1_srl_148_n14), .B1(n4166), .B2(
        u1_srl_148_n15), .ZN(u1_srl_148_n302) );
  AOI221_X1 u1_srl_148_U297 ( .B1(u1_srl_148_n224), .B2(n6325), .C1(
        u1_srl_148_n12), .C2(n6324), .A(u1_srl_148_n88), .ZN(u1_srl_148_n266)
         );
  AOI222_X1 u1_srl_148_U296 ( .A1(u1_srl_148_n84), .A2(u1_srl_148_n9), .B1(
        u1_srl_148_n86), .B2(u1_srl_148_n195), .C1(u1_srl_148_n87), .C2(
        u1_srl_148_n211), .ZN(u1_srl_148_n188) );
  AOI22_X1 u1_srl_148_U295 ( .A1(n6338), .A2(u1_srl_148_n197), .B1(n6340), 
        .B2(u1_srl_148_n198), .ZN(u1_srl_148_n301) );
  OAI221_X1 u1_srl_148_U294 ( .B1(u1_srl_148_n5), .B2(u1_srl_148_n125), .C1(
        u1_srl_148_n2), .C2(u1_srl_148_n124), .A(u1_srl_148_n301), .ZN(
        u1_srl_148_n139) );
  AOI22_X1 u1_srl_148_U293 ( .A1(u1_srl_148_n144), .A2(u1_srl_148_n82), .B1(
        u1_srl_148_n145), .B2(u1_srl_148_n139), .ZN(u1_srl_148_n296) );
  AOI22_X1 u1_srl_148_U292 ( .A1(n4185), .A2(u1_srl_148_n197), .B1(n6337), 
        .B2(u1_srl_148_n15), .ZN(u1_srl_148_n300) );
  OAI221_X1 u1_srl_148_U291 ( .B1(u1_srl_148_n5), .B2(u1_srl_148_n121), .C1(
        u1_srl_148_n2), .C2(u1_srl_148_n120), .A(u1_srl_148_n300), .ZN(
        u1_srl_148_n143) );
  AOI22_X1 u1_srl_148_U290 ( .A1(n4177), .A2(u1_srl_148_n14), .B1(n4180), .B2(
        u1_srl_148_n198), .ZN(u1_srl_148_n299) );
  OAI221_X1 u1_srl_148_U289 ( .B1(u1_srl_148_n5), .B2(u1_srl_148_n113), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n112), .A(u1_srl_148_n299), .ZN(
        u1_srl_148_n235) );
  AOI22_X1 u1_srl_148_U288 ( .A1(n4181), .A2(u1_srl_148_n197), .B1(n6335), 
        .B2(u1_srl_148_n15), .ZN(u1_srl_148_n298) );
  OAI221_X1 u1_srl_148_U287 ( .B1(u1_srl_148_n5), .B2(u1_srl_148_n117), .C1(
        u1_srl_148_n2), .C2(u1_srl_148_n116), .A(u1_srl_148_n298), .ZN(
        u1_srl_148_n141) );
  AOI222_X1 u1_srl_148_U286 ( .A1(u1_srl_148_n138), .A2(u1_srl_148_n143), .B1(
        u1_srl_148_n140), .B2(u1_srl_148_n235), .C1(u1_srl_148_n142), .C2(
        u1_srl_148_n141), .ZN(u1_srl_148_n297) );
  OAI211_X1 u1_srl_148_U285 ( .C1(u1_srl_148_n227), .C2(u1_srl_148_n96), .A(
        u1_srl_148_n296), .B(u1_srl_148_n297), .ZN(u1_adj_op_out_sft_13_) );
  AOI22_X1 u1_srl_148_U284 ( .A1(u1_srl_148_n237), .A2(u1_srl_148_n50), .B1(
        u1_srl_148_n195), .B2(u1_srl_148_n260), .ZN(u1_srl_148_n295) );
  AOI221_X1 u1_srl_148_U283 ( .B1(u1_srl_148_n258), .B2(u1_srl_148_n9), .C1(
        u1_srl_148_n259), .C2(u1_srl_148_n17), .A(u1_srl_148_n43), .ZN(
        u1_srl_148_n218) );
  AOI222_X1 u1_srl_148_U282 ( .A1(u1_srl_148_n53), .A2(u1_srl_148_n9), .B1(
        u1_srl_148_n52), .B2(u1_srl_148_n195), .C1(u1_srl_148_n48), .C2(
        u1_srl_148_n211), .ZN(u1_srl_148_n187) );
  AOI22_X1 u1_srl_148_U281 ( .A1(u1_srl_148_n144), .A2(u1_srl_148_n47), .B1(
        u1_srl_148_n145), .B2(u1_srl_148_n168), .ZN(u1_srl_148_n293) );
  AOI222_X1 u1_srl_148_U280 ( .A1(u1_srl_148_n138), .A2(u1_srl_148_n167), .B1(
        u1_srl_148_n140), .B2(u1_srl_148_n255), .C1(u1_srl_148_n142), .C2(
        u1_srl_148_n256), .ZN(u1_srl_148_n294) );
  OAI211_X1 u1_srl_148_U279 ( .C1(u1_srl_148_n218), .C2(u1_srl_148_n96), .A(
        u1_srl_148_n293), .B(u1_srl_148_n294), .ZN(u1_adj_op_out_sft_14_) );
  OAI22_X1 u1_srl_148_U278 ( .A1(u1_srl_148_n91), .A2(u1_srl_148_n254), .B1(
        u1_srl_148_n4), .B2(u1_srl_148_n283), .ZN(u1_srl_148_n292) );
  AOI221_X1 u1_srl_148_U277 ( .B1(u1_srl_148_n281), .B2(u1_srl_148_n10), .C1(
        u1_srl_148_n279), .C2(u1_srl_148_n211), .A(u1_srl_148_n292), .ZN(
        u1_srl_148_n216) );
  OAI222_X1 u1_srl_148_U276 ( .A1(u1_srl_148_n252), .A2(u1_srl_148_n1), .B1(
        u1_srl_148_n4), .B2(u1_srl_148_n175), .C1(u1_srl_148_n253), .C2(
        u1_srl_148_n18), .ZN(u1_srl_148_n217) );
  AOI22_X1 u1_srl_148_U275 ( .A1(u1_srl_148_n144), .A2(u1_srl_148_n217), .B1(
        u1_srl_148_n145), .B2(u1_srl_148_n160), .ZN(u1_srl_148_n290) );
  AOI222_X1 u1_srl_148_U274 ( .A1(u1_srl_148_n138), .A2(u1_srl_148_n159), .B1(
        u1_srl_148_n140), .B2(u1_srl_148_n248), .C1(u1_srl_148_n142), .C2(
        u1_srl_148_n249), .ZN(u1_srl_148_n291) );
  OAI211_X1 u1_srl_148_U273 ( .C1(u1_srl_148_n216), .C2(u1_srl_148_n96), .A(
        u1_srl_148_n290), .B(u1_srl_148_n291), .ZN(u1_adj_op_out_sft_15_) );
  OAI222_X1 u1_srl_148_U272 ( .A1(u1_srl_148_n215), .A2(u1_srl_148_n96), .B1(
        u1_srl_148_n186), .B2(u1_srl_148_n94), .C1(u1_srl_148_n289), .C2(
        u1_srl_148_n8), .ZN(u1_adj_op_out_sft_16_) );
  OAI22_X1 u1_srl_148_U271 ( .A1(u1_srl_148_n91), .A2(u1_srl_148_n266), .B1(
        u1_srl_148_n4), .B2(u1_srl_148_n267), .ZN(u1_srl_148_n288) );
  AOI221_X1 u1_srl_148_U270 ( .B1(u1_srl_148_n238), .B2(u1_srl_148_n10), .C1(
        u1_srl_148_n239), .C2(u1_srl_148_n17), .A(u1_srl_148_n288), .ZN(
        u1_srl_148_n214) );
  AOI22_X1 u1_srl_148_U269 ( .A1(u1_srl_148_n84), .A2(u1_srl_148_n17), .B1(
        u1_srl_148_n86), .B2(u1_srl_148_n10), .ZN(u1_srl_148_n185) );
  AOI22_X1 u1_srl_148_U268 ( .A1(u1_srl_148_n237), .A2(u1_srl_148_n234), .B1(
        u1_srl_148_n195), .B2(u1_srl_148_n235), .ZN(u1_srl_148_n287) );
  AOI221_X1 u1_srl_148_U267 ( .B1(u1_srl_148_n141), .B2(u1_srl_148_n9), .C1(
        u1_srl_148_n143), .C2(u1_srl_148_n17), .A(u1_srl_148_n76), .ZN(
        u1_srl_148_n277) );
  OAI222_X1 u1_srl_148_U266 ( .A1(u1_srl_148_n214), .A2(u1_srl_148_n96), .B1(
        u1_srl_148_n185), .B2(u1_srl_148_n94), .C1(u1_srl_148_n277), .C2(
        u1_srl_148_n8), .ZN(u1_adj_op_out_sft_17_) );
  OAI22_X1 u1_srl_148_U265 ( .A1(u1_srl_148_n91), .A2(u1_srl_148_n263), .B1(
        u1_srl_148_n4), .B2(u1_srl_148_n286), .ZN(u1_srl_148_n285) );
  AOI221_X1 u1_srl_148_U264 ( .B1(u1_srl_148_n260), .B2(u1_srl_148_n9), .C1(
        u1_srl_148_n258), .C2(u1_srl_148_n17), .A(u1_srl_148_n285), .ZN(
        u1_srl_148_n213) );
  AOI22_X1 u1_srl_148_U263 ( .A1(u1_srl_148_n53), .A2(u1_srl_148_n17), .B1(
        u1_srl_148_n52), .B2(u1_srl_148_n10), .ZN(u1_srl_148_n180) );
  AOI22_X1 u1_srl_148_U262 ( .A1(u1_srl_148_n237), .A2(u1_srl_148_n259), .B1(
        u1_srl_148_n195), .B2(u1_srl_148_n255), .ZN(u1_srl_148_n284) );
  AOI221_X1 u1_srl_148_U261 ( .B1(u1_srl_148_n256), .B2(u1_srl_148_n9), .C1(
        u1_srl_148_n167), .C2(u1_srl_148_n17), .A(u1_srl_148_n39), .ZN(
        u1_srl_148_n226) );
  OAI222_X1 u1_srl_148_U260 ( .A1(u1_srl_148_n213), .A2(u1_srl_148_n96), .B1(
        u1_srl_148_n180), .B2(u1_srl_148_n94), .C1(u1_srl_148_n226), .C2(
        u1_srl_148_n8), .ZN(u1_adj_op_out_sft_18_) );
  OAI22_X1 u1_srl_148_U259 ( .A1(u1_srl_148_n91), .A2(u1_srl_148_n253), .B1(
        u1_srl_148_n4), .B2(u1_srl_148_n254), .ZN(u1_srl_148_n282) );
  AOI221_X1 u1_srl_148_U258 ( .B1(u1_srl_148_n61), .B2(u1_srl_148_n10), .C1(
        u1_srl_148_n281), .C2(u1_srl_148_n17), .A(u1_srl_148_n282), .ZN(
        u1_srl_148_n212) );
  OR2_X1 u1_srl_148_U257 ( .A1(u1_srl_148_n280), .A2(n6301), .ZN(
        u1_srl_148_n179) );
  OAI22_X1 u1_srl_148_U256 ( .A1(u1_srl_148_n91), .A2(u1_srl_148_n57), .B1(
        u1_srl_148_n4), .B2(u1_srl_148_n58), .ZN(u1_srl_148_n278) );
  AOI221_X1 u1_srl_148_U255 ( .B1(u1_srl_148_n249), .B2(u1_srl_148_n9), .C1(
        u1_srl_148_n159), .C2(u1_srl_148_n17), .A(u1_srl_148_n278), .ZN(
        u1_srl_148_n200) );
  OAI222_X1 u1_srl_148_U254 ( .A1(u1_srl_148_n212), .A2(u1_srl_148_n96), .B1(
        u1_srl_148_n94), .B2(u1_srl_148_n179), .C1(u1_srl_148_n200), .C2(
        u1_srl_148_n8), .ZN(u1_adj_op_out_sft_19_) );
  AOI22_X1 u1_srl_148_U253 ( .A1(n6344), .A2(u1_srl_148_n197), .B1(n6308), 
        .B2(u1_srl_148_n198), .ZN(u1_srl_148_n276) );
  OAI221_X1 u1_srl_148_U252 ( .B1(u1_srl_148_n5), .B2(u1_srl_148_n133), .C1(
        u1_srl_148_n2), .C2(u1_srl_148_n132), .A(u1_srl_148_n276), .ZN(
        u1_srl_148_n173) );
  AOI222_X1 u1_srl_148_U251 ( .A1(u1_srl_148_n162), .A2(u1_srl_148_n75), .B1(
        u1_srl_148_n138), .B2(u1_srl_148_n173), .C1(u1_srl_148_n144), .C2(
        u1_srl_148_n71), .ZN(u1_srl_148_n271) );
  AOI22_X1 u1_srl_148_U250 ( .A1(u1_srl_148_n197), .A2(n6347), .B1(
        u1_srl_148_n12), .B2(n6348), .ZN(u1_srl_148_n273) );
  AOI22_X1 u1_srl_148_U249 ( .A1(n4193), .A2(u1_srl_148_n197), .B1(n6343), 
        .B2(u1_srl_148_n198), .ZN(u1_srl_148_n275) );
  OAI221_X1 u1_srl_148_U248 ( .B1(u1_srl_148_n5), .B2(u1_srl_148_n129), .C1(
        u1_srl_148_n2), .C2(u1_srl_148_n128), .A(u1_srl_148_n275), .ZN(
        u1_srl_148_n146) );
  AOI22_X1 u1_srl_148_U247 ( .A1(u1_srl_148_n146), .A2(u1_srl_148_n142), .B1(
        u1_srl_148_n139), .B2(u1_srl_148_n140), .ZN(u1_srl_148_n274) );
  OAI221_X1 u1_srl_148_U246 ( .B1(u1_srl_148_n90), .B2(u1_srl_148_n273), .C1(
        u1_srl_148_n223), .C2(u1_srl_148_n185), .A(u1_srl_148_n274), .ZN(
        u1_srl_148_n272) );
  NAND2_X1 u1_srl_148_U245 ( .A1(u1_srl_148_n271), .A2(u1_srl_148_n83), .ZN(
        u1_adj_op_out_sft_1_) );
  OAI22_X1 u1_srl_148_U244 ( .A1(u1_srl_148_n91), .A2(u1_srl_148_n241), .B1(
        u1_srl_148_n4), .B2(u1_srl_148_n270), .ZN(u1_srl_148_n269) );
  AOI221_X1 u1_srl_148_U243 ( .B1(u1_srl_148_n31), .B2(u1_srl_148_n10), .C1(
        u1_srl_148_n245), .C2(u1_srl_148_n17), .A(u1_srl_148_n269), .ZN(
        u1_srl_148_n210) );
  NAND2_X1 u1_srl_148_U242 ( .A1(u1_srl_148_n144), .A2(u1_srl_148_n211), .ZN(
        u1_srl_148_n247) );
  AOI22_X1 u1_srl_148_U241 ( .A1(u1_srl_148_n237), .A2(u1_srl_148_n246), .B1(
        u1_srl_148_n195), .B2(u1_srl_148_n242), .ZN(u1_srl_148_n268) );
  AOI221_X1 u1_srl_148_U240 ( .B1(u1_srl_148_n243), .B2(u1_srl_148_n9), .C1(
        u1_srl_148_n152), .C2(u1_srl_148_n17), .A(u1_srl_148_n21), .ZN(
        u1_srl_148_n184) );
  OAI222_X1 u1_srl_148_U239 ( .A1(u1_srl_148_n210), .A2(u1_srl_148_n96), .B1(
        u1_srl_148_n178), .B2(u1_srl_148_n247), .C1(u1_srl_148_n184), .C2(
        u1_srl_148_n8), .ZN(u1_adj_op_out_sft_20_) );
  OAI22_X1 u1_srl_148_U238 ( .A1(u1_srl_148_n91), .A2(u1_srl_148_n233), .B1(
        u1_srl_148_n4), .B2(u1_srl_148_n266), .ZN(u1_srl_148_n265) );
  AOI221_X1 u1_srl_148_U237 ( .B1(u1_srl_148_n79), .B2(u1_srl_148_n10), .C1(
        u1_srl_148_n238), .C2(u1_srl_148_n17), .A(u1_srl_148_n265), .ZN(
        u1_srl_148_n208) );
  AOI22_X1 u1_srl_148_U236 ( .A1(u1_srl_148_n237), .A2(u1_srl_148_n239), .B1(
        u1_srl_148_n195), .B2(u1_srl_148_n234), .ZN(u1_srl_148_n264) );
  AOI221_X1 u1_srl_148_U235 ( .B1(u1_srl_148_n235), .B2(u1_srl_148_n9), .C1(
        u1_srl_148_n141), .C2(u1_srl_148_n17), .A(u1_srl_148_n73), .ZN(
        u1_srl_148_n174) );
  OAI222_X1 u1_srl_148_U234 ( .A1(u1_srl_148_n208), .A2(u1_srl_148_n96), .B1(
        u1_srl_148_n177), .B2(u1_srl_148_n247), .C1(u1_srl_148_n174), .C2(
        u1_srl_148_n8), .ZN(u1_adj_op_out_sft_21_) );
  OAI22_X1 u1_srl_148_U233 ( .A1(u1_srl_148_n91), .A2(u1_srl_148_n262), .B1(
        u1_srl_148_n4), .B2(u1_srl_148_n263), .ZN(u1_srl_148_n261) );
  AOI221_X1 u1_srl_148_U232 ( .B1(u1_srl_148_n50), .B2(u1_srl_148_n9), .C1(
        u1_srl_148_n260), .C2(u1_srl_148_n17), .A(u1_srl_148_n261), .ZN(
        u1_srl_148_n206) );
  AOI22_X1 u1_srl_148_U231 ( .A1(u1_srl_148_n237), .A2(u1_srl_148_n258), .B1(
        u1_srl_148_n195), .B2(u1_srl_148_n259), .ZN(u1_srl_148_n257) );
  AOI221_X1 u1_srl_148_U230 ( .B1(u1_srl_148_n255), .B2(u1_srl_148_n9), .C1(
        u1_srl_148_n256), .C2(u1_srl_148_n17), .A(u1_srl_148_n41), .ZN(
        u1_srl_148_n170) );
  OAI222_X1 u1_srl_148_U229 ( .A1(u1_srl_148_n206), .A2(u1_srl_148_n96), .B1(
        u1_srl_148_n176), .B2(u1_srl_148_n247), .C1(u1_srl_148_n170), .C2(
        u1_srl_148_n8), .ZN(u1_adj_op_out_sft_22_) );
  OAI22_X1 u1_srl_148_U228 ( .A1(u1_srl_148_n91), .A2(u1_srl_148_n252), .B1(
        u1_srl_148_n4), .B2(u1_srl_148_n253), .ZN(u1_srl_148_n251) );
  AOI221_X1 u1_srl_148_U227 ( .B1(u1_srl_148_n65), .B2(u1_srl_148_n9), .C1(
        u1_srl_148_n61), .C2(u1_srl_148_n211), .A(u1_srl_148_n251), .ZN(
        u1_srl_148_n203) );
  OAI22_X1 u1_srl_148_U226 ( .A1(u1_srl_148_n91), .A2(u1_srl_148_n63), .B1(
        u1_srl_148_n4), .B2(u1_srl_148_n57), .ZN(u1_srl_148_n250) );
  AOI221_X1 u1_srl_148_U225 ( .B1(u1_srl_148_n248), .B2(u1_srl_148_n9), .C1(
        u1_srl_148_n249), .C2(u1_srl_148_n17), .A(u1_srl_148_n250), .ZN(
        u1_srl_148_n163) );
  OAI222_X1 u1_srl_148_U224 ( .A1(u1_srl_148_n203), .A2(u1_srl_148_n96), .B1(
        u1_srl_148_n175), .B2(u1_srl_148_n247), .C1(u1_srl_148_n163), .C2(
        u1_srl_148_n8), .ZN(u1_adj_op_out_sft_23_) );
  AOI22_X1 u1_srl_148_U223 ( .A1(u1_srl_148_n237), .A2(u1_srl_148_n245), .B1(
        u1_srl_148_n195), .B2(u1_srl_148_n246), .ZN(u1_srl_148_n244) );
  AOI221_X1 u1_srl_148_U222 ( .B1(u1_srl_148_n242), .B2(u1_srl_148_n9), .C1(
        u1_srl_148_n243), .C2(u1_srl_148_n211), .A(u1_srl_148_n26), .ZN(
        u1_srl_148_n148) );
  OAI22_X1 u1_srl_148_U221 ( .A1(u1_srl_148_n91), .A2(u1_srl_148_n178), .B1(
        u1_srl_148_n4), .B2(u1_srl_148_n241), .ZN(u1_srl_148_n240) );
  AOI221_X1 u1_srl_148_U220 ( .B1(u1_srl_148_n29), .B2(u1_srl_148_n9), .C1(
        u1_srl_148_n31), .C2(u1_srl_148_n211), .A(u1_srl_148_n240), .ZN(
        u1_srl_148_n155) );
  OAI22_X1 u1_srl_148_U219 ( .A1(u1_srl_148_n148), .A2(u1_srl_148_n7), .B1(
        u1_srl_148_n155), .B2(u1_srl_148_n96), .ZN(u1_adj_op_out_sft_24_) );
  AOI22_X1 u1_srl_148_U218 ( .A1(u1_srl_148_n237), .A2(u1_srl_148_n238), .B1(
        u1_srl_148_n195), .B2(u1_srl_148_n239), .ZN(u1_srl_148_n236) );
  AOI221_X1 u1_srl_148_U217 ( .B1(u1_srl_148_n234), .B2(u1_srl_148_n9), .C1(
        u1_srl_148_n235), .C2(u1_srl_148_n211), .A(u1_srl_148_n74), .ZN(
        u1_srl_148_n135) );
  OAI22_X1 u1_srl_148_U216 ( .A1(u1_srl_148_n91), .A2(u1_srl_148_n177), .B1(
        u1_srl_148_n4), .B2(u1_srl_148_n233), .ZN(u1_srl_148_n232) );
  AOI221_X1 u1_srl_148_U215 ( .B1(u1_srl_148_n87), .B2(u1_srl_148_n9), .C1(
        u1_srl_148_n79), .C2(u1_srl_148_n211), .A(u1_srl_148_n232), .ZN(
        u1_srl_148_n147) );
  OAI22_X1 u1_srl_148_U214 ( .A1(u1_srl_148_n135), .A2(u1_srl_148_n7), .B1(
        u1_srl_148_n147), .B2(u1_srl_148_n96), .ZN(u1_adj_op_out_sft_25_) );
  OAI22_X1 u1_srl_148_U213 ( .A1(u1_srl_148_n231), .A2(u1_srl_148_n7), .B1(
        u1_srl_148_n190), .B2(u1_srl_148_n96), .ZN(u1_adj_op_out_sft_26_) );
  OAI22_X1 u1_srl_148_U212 ( .A1(u1_srl_148_n229), .A2(u1_srl_148_n7), .B1(
        u1_srl_148_n64), .B2(u1_srl_148_n96), .ZN(u1_adj_op_out_sft_27_) );
  OAI22_X1 u1_srl_148_U211 ( .A1(u1_srl_148_n228), .A2(u1_srl_148_n7), .B1(
        u1_srl_148_n189), .B2(u1_srl_148_n96), .ZN(u1_adj_op_out_sft_28_) );
  OAI22_X1 u1_srl_148_U210 ( .A1(u1_srl_148_n227), .A2(u1_srl_148_n7), .B1(
        u1_srl_148_n188), .B2(u1_srl_148_n96), .ZN(u1_adj_op_out_sft_29_) );
  AOI22_X1 u1_srl_148_U209 ( .A1(n6343), .A2(u1_srl_148_n197), .B1(n6346), 
        .B2(u1_srl_148_n198), .ZN(u1_srl_148_n225) );
  OAI221_X1 u1_srl_148_U208 ( .B1(u1_srl_148_n5), .B2(u1_srl_148_n132), .C1(
        u1_srl_148_n2), .C2(u1_srl_148_n131), .A(u1_srl_148_n225), .ZN(
        u1_srl_148_n169) );
  AOI222_X1 u1_srl_148_U207 ( .A1(u1_srl_148_n162), .A2(u1_srl_148_n38), .B1(
        u1_srl_148_n138), .B2(u1_srl_148_n169), .C1(u1_srl_148_n144), .C2(
        u1_srl_148_n44), .ZN(u1_srl_148_n219) );
  AOI222_X1 u1_srl_148_U206 ( .A1(n6308), .A2(u1_srl_148_n197), .B1(n6348), 
        .B2(u1_srl_148_n224), .C1(n6347), .C2(u1_srl_148_n12), .ZN(
        u1_srl_148_n222) );
  OAI22_X1 u1_srl_148_U205 ( .A1(u1_srl_148_n222), .A2(u1_srl_148_n90), .B1(
        u1_srl_148_n180), .B2(u1_srl_148_n223), .ZN(u1_srl_148_n221) );
  AOI221_X1 u1_srl_148_U204 ( .B1(u1_srl_148_n140), .B2(u1_srl_148_n168), .C1(
        u1_srl_148_n142), .C2(u1_srl_148_n166), .A(u1_srl_148_n221), .ZN(
        u1_srl_148_n220) );
  NAND2_X1 u1_srl_148_U203 ( .A1(u1_srl_148_n219), .A2(u1_srl_148_n220), .ZN(
        u1_adj_op_out_sft_2_) );
  OAI22_X1 u1_srl_148_U202 ( .A1(u1_srl_148_n218), .A2(u1_srl_148_n7), .B1(
        u1_srl_148_n187), .B2(u1_srl_148_n96), .ZN(u1_adj_op_out_sft_30_) );
  OAI22_X1 u1_srl_148_U201 ( .A1(u1_srl_148_n216), .A2(u1_srl_148_n8), .B1(
        u1_srl_148_n67), .B2(u1_srl_148_n96), .ZN(u1_adj_op_out_sft_31_) );
  OAI22_X1 u1_srl_148_U200 ( .A1(u1_srl_148_n215), .A2(u1_srl_148_n7), .B1(
        u1_srl_148_n186), .B2(u1_srl_148_n96), .ZN(u1_adj_op_out_sft_32_) );
  OAI22_X1 u1_srl_148_U199 ( .A1(u1_srl_148_n214), .A2(u1_srl_148_n8), .B1(
        u1_srl_148_n185), .B2(u1_srl_148_n96), .ZN(u1_adj_op_out_sft_33_) );
  OAI22_X1 u1_srl_148_U198 ( .A1(u1_srl_148_n213), .A2(u1_srl_148_n8), .B1(
        u1_srl_148_n180), .B2(u1_srl_148_n96), .ZN(u1_adj_op_out_sft_34_) );
  MUX2_X1 u1_srl_148_U197 ( .A(u1_srl_148_n179), .B(u1_srl_148_n212), .S(
        u1_srl_148_n97), .Z(u1_srl_148_n201) );
  NOR2_X1 u1_srl_148_U196 ( .A1(n6302), .A2(u1_srl_148_n201), .ZN(
        u1_adj_op_out_sft_35_) );
  NAND2_X1 u1_srl_148_U195 ( .A1(n6303), .A2(u1_srl_148_n17), .ZN(
        u1_srl_148_n204) );
  OAI22_X1 u1_srl_148_U194 ( .A1(n6303), .A2(u1_srl_148_n210), .B1(
        u1_srl_148_n178), .B2(u1_srl_148_n204), .ZN(u1_srl_148_n209) );
  NOR2_X1 u1_srl_148_U193 ( .A1(n6302), .A2(u1_srl_148_n25), .ZN(
        u1_adj_op_out_sft_36_) );
  OAI22_X1 u1_srl_148_U192 ( .A1(n6303), .A2(u1_srl_148_n208), .B1(
        u1_srl_148_n177), .B2(u1_srl_148_n204), .ZN(u1_srl_148_n207) );
  NOR2_X1 u1_srl_148_U191 ( .A1(n6302), .A2(u1_srl_148_n77), .ZN(
        u1_adj_op_out_sft_37_) );
  OAI22_X1 u1_srl_148_U190 ( .A1(n6303), .A2(u1_srl_148_n206), .B1(
        u1_srl_148_n176), .B2(u1_srl_148_n204), .ZN(u1_srl_148_n205) );
  NOR2_X1 u1_srl_148_U189 ( .A1(n6302), .A2(u1_srl_148_n45), .ZN(
        u1_adj_op_out_sft_38_) );
  OAI22_X1 u1_srl_148_U188 ( .A1(n6303), .A2(u1_srl_148_n203), .B1(
        u1_srl_148_n204), .B2(u1_srl_148_n175), .ZN(u1_srl_148_n202) );
  NOR2_X1 u1_srl_148_U187 ( .A1(n6302), .A2(u1_srl_148_n60), .ZN(
        u1_adj_op_out_sft_39_) );
  OAI22_X1 u1_srl_148_U186 ( .A1(u1_srl_148_n2), .A2(u1_srl_148_n104), .B1(
        u1_srl_148_n5), .B2(u1_srl_148_n134), .ZN(u1_srl_148_n199) );
  AOI221_X1 u1_srl_148_U185 ( .B1(n6346), .B2(u1_srl_148_n197), .C1(n6348), 
        .C2(u1_srl_148_n198), .A(u1_srl_148_n199), .ZN(u1_srl_148_n193) );
  AOI22_X1 u1_srl_148_U184 ( .A1(n6342), .A2(u1_srl_148_n14), .B1(n6345), .B2(
        u1_srl_148_n15), .ZN(u1_srl_148_n196) );
  OAI221_X1 u1_srl_148_U183 ( .B1(u1_srl_148_n5), .B2(u1_srl_148_n131), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n130), .A(u1_srl_148_n196), .ZN(
        u1_srl_148_n161) );
  AOI22_X1 u1_srl_148_U182 ( .A1(u1_srl_148_n195), .A2(u1_srl_148_n158), .B1(
        u1_srl_148_n10), .B2(u1_srl_148_n161), .ZN(u1_srl_148_n194) );
  OAI221_X1 u1_srl_148_U181 ( .B1(u1_srl_148_n193), .B2(u1_srl_148_n18), .C1(
        u1_srl_148_n70), .C2(u1_srl_148_n91), .A(u1_srl_148_n194), .ZN(
        u1_srl_148_n192) );
  MUX2_X1 u1_srl_148_U180 ( .A(u1_srl_148_n55), .B(u1_srl_148_n192), .S(
        u1_srl_148_n97), .Z(u1_srl_148_n191) );
  MUX2_X1 u1_srl_148_U179 ( .A(u1_srl_148_n59), .B(u1_srl_148_n191), .S(
        u1_srl_148_n95), .Z(u1_adj_op_out_sft_3_) );
  NOR2_X1 u1_srl_148_U178 ( .A1(u1_srl_148_n155), .A2(u1_srl_148_n7), .ZN(
        u1_adj_op_out_sft_40_) );
  NOR2_X1 u1_srl_148_U177 ( .A1(u1_srl_148_n147), .A2(u1_srl_148_n7), .ZN(
        u1_adj_op_out_sft_41_) );
  NOR2_X1 u1_srl_148_U176 ( .A1(u1_srl_148_n190), .A2(u1_srl_148_n7), .ZN(
        u1_adj_op_out_sft_42_) );
  NOR2_X1 u1_srl_148_U175 ( .A1(u1_srl_148_n64), .A2(u1_srl_148_n7), .ZN(
        u1_adj_op_out_sft_43_) );
  NOR2_X1 u1_srl_148_U174 ( .A1(u1_srl_148_n189), .A2(u1_srl_148_n7), .ZN(
        u1_adj_op_out_sft_44_) );
  NOR2_X1 u1_srl_148_U173 ( .A1(u1_srl_148_n188), .A2(u1_srl_148_n7), .ZN(
        u1_adj_op_out_sft_45_) );
  NOR2_X1 u1_srl_148_U172 ( .A1(u1_srl_148_n187), .A2(u1_srl_148_n7), .ZN(
        u1_adj_op_out_sft_46_) );
  NOR2_X1 u1_srl_148_U171 ( .A1(u1_srl_148_n67), .A2(u1_srl_148_n7), .ZN(
        u1_adj_op_out_sft_47_) );
  NOR2_X1 u1_srl_148_U170 ( .A1(u1_srl_148_n186), .A2(u1_srl_148_n7), .ZN(
        u1_adj_op_out_sft_48_) );
  NOR2_X1 u1_srl_148_U169 ( .A1(u1_srl_148_n185), .A2(u1_srl_148_n7), .ZN(
        u1_adj_op_out_sft_49_) );
  AOI22_X1 u1_srl_148_U168 ( .A1(u1_srl_148_n145), .A2(u1_srl_148_n183), .B1(
        u1_srl_148_n162), .B2(u1_srl_148_n20), .ZN(u1_srl_148_n181) );
  AOI222_X1 u1_srl_148_U167 ( .A1(u1_srl_148_n138), .A2(u1_srl_148_n154), .B1(
        u1_srl_148_n140), .B2(u1_srl_148_n153), .C1(u1_srl_148_n142), .C2(
        u1_srl_148_n151), .ZN(u1_srl_148_n182) );
  OAI211_X1 u1_srl_148_U166 ( .C1(u1_srl_148_n25), .C2(u1_srl_148_n95), .A(
        u1_srl_148_n181), .B(u1_srl_148_n182), .ZN(u1_adj_op_out_sft_4_) );
  NOR2_X1 u1_srl_148_U165 ( .A1(u1_srl_148_n180), .A2(u1_srl_148_n7), .ZN(
        u1_adj_op_out_sft_50_) );
  NOR2_X1 u1_srl_148_U164 ( .A1(u1_srl_148_n7), .A2(u1_srl_148_n179), .ZN(
        u1_adj_op_out_sft_51_) );
  NOR2_X1 u1_srl_148_U163 ( .A1(u1_srl_148_n178), .A2(u1_srl_148_n90), .ZN(
        u1_adj_op_out_sft_52_) );
  NOR2_X1 u1_srl_148_U162 ( .A1(u1_srl_148_n177), .A2(u1_srl_148_n90), .ZN(
        u1_adj_op_out_sft_53_) );
  NOR2_X1 u1_srl_148_U161 ( .A1(u1_srl_148_n176), .A2(u1_srl_148_n90), .ZN(
        u1_adj_op_out_sft_54_) );
  NOR2_X1 u1_srl_148_U160 ( .A1(u1_srl_148_n90), .A2(u1_srl_148_n175), .ZN(
        u1_adj_op_out_sft_55_) );
  AOI22_X1 u1_srl_148_U159 ( .A1(u1_srl_148_n145), .A2(u1_srl_148_n173), .B1(
        u1_srl_148_n162), .B2(u1_srl_148_n72), .ZN(u1_srl_148_n171) );
  AOI222_X1 u1_srl_148_U158 ( .A1(u1_srl_148_n138), .A2(u1_srl_148_n146), .B1(
        u1_srl_148_n140), .B2(u1_srl_148_n143), .C1(u1_srl_148_n142), .C2(
        u1_srl_148_n139), .ZN(u1_srl_148_n172) );
  OAI211_X1 u1_srl_148_U157 ( .C1(u1_srl_148_n77), .C2(u1_srl_148_n95), .A(
        u1_srl_148_n171), .B(u1_srl_148_n172), .ZN(u1_adj_op_out_sft_5_) );
  AOI22_X1 u1_srl_148_U156 ( .A1(u1_srl_148_n145), .A2(u1_srl_148_n169), .B1(
        u1_srl_148_n162), .B2(u1_srl_148_n40), .ZN(u1_srl_148_n164) );
  AOI222_X1 u1_srl_148_U155 ( .A1(u1_srl_148_n138), .A2(u1_srl_148_n166), .B1(
        u1_srl_148_n140), .B2(u1_srl_148_n167), .C1(u1_srl_148_n142), .C2(
        u1_srl_148_n168), .ZN(u1_srl_148_n165) );
  OAI211_X1 u1_srl_148_U154 ( .C1(u1_srl_148_n45), .C2(u1_srl_148_n95), .A(
        u1_srl_148_n164), .B(u1_srl_148_n165), .ZN(u1_adj_op_out_sft_6_) );
  AOI22_X1 u1_srl_148_U153 ( .A1(u1_srl_148_n145), .A2(u1_srl_148_n161), .B1(
        u1_srl_148_n162), .B2(u1_srl_148_n56), .ZN(u1_srl_148_n156) );
  AOI222_X1 u1_srl_148_U152 ( .A1(u1_srl_148_n138), .A2(u1_srl_148_n158), .B1(
        u1_srl_148_n140), .B2(u1_srl_148_n159), .C1(u1_srl_148_n142), .C2(
        u1_srl_148_n160), .ZN(u1_srl_148_n157) );
  OAI211_X1 u1_srl_148_U151 ( .C1(u1_srl_148_n60), .C2(u1_srl_148_n95), .A(
        u1_srl_148_n156), .B(u1_srl_148_n157), .ZN(u1_adj_op_out_sft_7_) );
  AOI22_X1 u1_srl_148_U150 ( .A1(u1_srl_148_n144), .A2(u1_srl_148_n28), .B1(
        u1_srl_148_n145), .B2(u1_srl_148_n154), .ZN(u1_srl_148_n149) );
  AOI222_X1 u1_srl_148_U149 ( .A1(u1_srl_148_n138), .A2(u1_srl_148_n151), .B1(
        u1_srl_148_n140), .B2(u1_srl_148_n152), .C1(u1_srl_148_n142), .C2(
        u1_srl_148_n153), .ZN(u1_srl_148_n150) );
  OAI211_X1 u1_srl_148_U148 ( .C1(u1_srl_148_n148), .C2(u1_srl_148_n96), .A(
        u1_srl_148_n149), .B(u1_srl_148_n150), .ZN(u1_adj_op_out_sft_8_) );
  AOI22_X1 u1_srl_148_U147 ( .A1(u1_srl_148_n144), .A2(u1_srl_148_n78), .B1(
        u1_srl_148_n145), .B2(u1_srl_148_n146), .ZN(u1_srl_148_n136) );
  AOI222_X1 u1_srl_148_U146 ( .A1(u1_srl_148_n138), .A2(u1_srl_148_n139), .B1(
        u1_srl_148_n140), .B2(u1_srl_148_n141), .C1(u1_srl_148_n142), .C2(
        u1_srl_148_n143), .ZN(u1_srl_148_n137) );
  OAI211_X1 u1_srl_148_U145 ( .C1(u1_srl_148_n135), .C2(u1_srl_148_n96), .A(
        u1_srl_148_n136), .B(u1_srl_148_n137), .ZN(u1_adj_op_out_sft_9_) );
  INV_X4 u1_srl_148_U144 ( .A(n6347), .ZN(u1_srl_148_n134) );
  INV_X4 u1_srl_148_U143 ( .A(n6346), .ZN(u1_srl_148_n133) );
  INV_X4 u1_srl_148_U142 ( .A(n6345), .ZN(u1_srl_148_n132) );
  INV_X4 u1_srl_148_U141 ( .A(n6344), .ZN(u1_srl_148_n131) );
  INV_X4 u1_srl_148_U140 ( .A(n6343), .ZN(u1_srl_148_n130) );
  INV_X4 u1_srl_148_U139 ( .A(n6342), .ZN(u1_srl_148_n129) );
  INV_X4 u1_srl_148_U138 ( .A(n6341), .ZN(u1_srl_148_n128) );
  INV_X4 u1_srl_148_U137 ( .A(n4193), .ZN(u1_srl_148_n127) );
  INV_X4 u1_srl_148_U136 ( .A(n6340), .ZN(u1_srl_148_n126) );
  INV_X4 u1_srl_148_U135 ( .A(n6339), .ZN(u1_srl_148_n125) );
  INV_X4 u1_srl_148_U134 ( .A(n4190), .ZN(u1_srl_148_n124) );
  INV_X4 u1_srl_148_U133 ( .A(n6338), .ZN(u1_srl_148_n123) );
  INV_X4 u1_srl_148_U132 ( .A(n6337), .ZN(u1_srl_148_n122) );
  INV_X4 u1_srl_148_U131 ( .A(n6336), .ZN(u1_srl_148_n121) );
  INV_X4 u1_srl_148_U130 ( .A(n4186), .ZN(u1_srl_148_n120) );
  INV_X4 u1_srl_148_U129 ( .A(n4185), .ZN(u1_srl_148_n119) );
  INV_X4 u1_srl_148_U128 ( .A(n6335), .ZN(u1_srl_148_n118) );
  INV_X4 u1_srl_148_U127 ( .A(n6334), .ZN(u1_srl_148_n117) );
  INV_X4 u1_srl_148_U126 ( .A(n6333), .ZN(u1_srl_148_n116) );
  INV_X4 u1_srl_148_U125 ( .A(n4181), .ZN(u1_srl_148_n115) );
  INV_X4 u1_srl_148_U124 ( .A(n4180), .ZN(u1_srl_148_n114) );
  INV_X4 u1_srl_148_U123 ( .A(n4179), .ZN(u1_srl_148_n113) );
  INV_X4 u1_srl_148_U122 ( .A(n6332), .ZN(u1_srl_148_n112) );
  INV_X4 u1_srl_148_U121 ( .A(n4177), .ZN(u1_srl_148_n111) );
  INV_X4 u1_srl_148_U120 ( .A(n6331), .ZN(u1_srl_148_n110) );
  INV_X4 u1_srl_148_U119 ( .A(n4175), .ZN(u1_srl_148_n109) );
  INV_X4 u1_srl_148_U118 ( .A(n4174), .ZN(u1_srl_148_n108) );
  INV_X4 u1_srl_148_U117 ( .A(n4173), .ZN(u1_srl_148_n107) );
  INV_X4 u1_srl_148_U116 ( .A(n6330), .ZN(u1_srl_148_n106) );
  INV_X4 u1_srl_148_U115 ( .A(n6329), .ZN(u1_srl_148_n105) );
  INV_X4 u1_srl_148_U114 ( .A(n6308), .ZN(u1_srl_148_n104) );
  INV_X4 u1_srl_148_U113 ( .A(u1_adj_op_29_), .ZN(u1_srl_148_n103) );
  INV_X4 u1_srl_148_U112 ( .A(n6307), .ZN(u1_srl_148_n102) );
  INV_X4 u1_srl_148_U111 ( .A(n6306), .ZN(u1_srl_148_n101) );
  INV_X4 u1_srl_148_U110 ( .A(n6305), .ZN(u1_srl_148_n100) );
  INV_X4 u1_srl_148_U109 ( .A(u1_adj_op_36_), .ZN(u1_srl_148_n99) );
  INV_X4 u1_srl_148_U108 ( .A(n6304), .ZN(u1_srl_148_n98) );
  INV_X4 u1_srl_148_U107 ( .A(n6303), .ZN(u1_srl_148_n97) );
  INV_X4 u1_srl_148_U106 ( .A(n6302), .ZN(u1_srl_148_n95) );
  INV_X4 u1_srl_148_U105 ( .A(u1_srl_148_n144), .ZN(u1_srl_148_n94) );
  INV_X4 u1_srl_148_U104 ( .A(n6301), .ZN(u1_srl_148_n93) );
  INV_X4 u1_srl_148_U103 ( .A(n6293), .ZN(u1_srl_148_n92) );
  INV_X4 u1_srl_148_U102 ( .A(u1_srl_148_n145), .ZN(u1_srl_148_n90) );
  INV_X4 u1_srl_148_U101 ( .A(u1_exp_diff_sft_0_), .ZN(u1_srl_148_n89) );
  INV_X4 u1_srl_148_U100 ( .A(u1_srl_148_n302), .ZN(u1_srl_148_n88) );
  INV_X4 u1_srl_148_U99 ( .A(u1_srl_148_n266), .ZN(u1_srl_148_n87) );
  INV_X4 u1_srl_148_U98 ( .A(u1_srl_148_n177), .ZN(u1_srl_148_n86) );
  INV_X4 u1_srl_148_U97 ( .A(u1_srl_148_n303), .ZN(u1_srl_148_n85) );
  INV_X4 u1_srl_148_U96 ( .A(u1_srl_148_n233), .ZN(u1_srl_148_n84) );
  INV_X4 u1_srl_148_U95 ( .A(u1_srl_148_n272), .ZN(u1_srl_148_n83) );
  INV_X4 u1_srl_148_U94 ( .A(u1_srl_148_n188), .ZN(u1_srl_148_n82) );
  INV_X4 u1_srl_148_U93 ( .A(u1_srl_148_n238), .ZN(u1_srl_148_n81) );
  INV_X4 u1_srl_148_U92 ( .A(u1_srl_148_n306), .ZN(u1_srl_148_n80) );
  INV_X4 u1_srl_148_U91 ( .A(u1_srl_148_n267), .ZN(u1_srl_148_n79) );
  INV_X4 u1_srl_148_U90 ( .A(u1_srl_148_n147), .ZN(u1_srl_148_n78) );
  INV_X4 u1_srl_148_U89 ( .A(u1_srl_148_n207), .ZN(u1_srl_148_n77) );
  INV_X4 u1_srl_148_U88 ( .A(u1_srl_148_n287), .ZN(u1_srl_148_n76) );
  INV_X4 u1_srl_148_U87 ( .A(u1_srl_148_n277), .ZN(u1_srl_148_n75) );
  INV_X4 u1_srl_148_U86 ( .A(u1_srl_148_n236), .ZN(u1_srl_148_n74) );
  INV_X4 u1_srl_148_U85 ( .A(u1_srl_148_n264), .ZN(u1_srl_148_n73) );
  INV_X4 u1_srl_148_U84 ( .A(u1_srl_148_n174), .ZN(u1_srl_148_n72) );
  INV_X4 u1_srl_148_U83 ( .A(u1_srl_148_n214), .ZN(u1_srl_148_n71) );
  INV_X4 u1_srl_148_U82 ( .A(u1_srl_148_n160), .ZN(u1_srl_148_n70) );
  INV_X4 u1_srl_148_U81 ( .A(u1_srl_148_n319), .ZN(u1_srl_148_n69) );
  INV_X4 u1_srl_148_U80 ( .A(u1_srl_148_n320), .ZN(u1_srl_148_n68) );
  INV_X4 u1_srl_148_U79 ( .A(u1_srl_148_n217), .ZN(u1_srl_148_n67) );
  INV_X4 u1_srl_148_U78 ( .A(u1_srl_148_n321), .ZN(u1_srl_148_n66) );
  INV_X4 u1_srl_148_U77 ( .A(u1_srl_148_n254), .ZN(u1_srl_148_n65) );
  INV_X4 u1_srl_148_U76 ( .A(u1_srl_148_n230), .ZN(u1_srl_148_n64) );
  INV_X4 u1_srl_148_U75 ( .A(u1_srl_148_n281), .ZN(u1_srl_148_n63) );
  INV_X4 u1_srl_148_U74 ( .A(u1_srl_148_n324), .ZN(u1_srl_148_n62) );
  INV_X4 u1_srl_148_U73 ( .A(u1_srl_148_n283), .ZN(u1_srl_148_n61) );
  INV_X4 u1_srl_148_U72 ( .A(u1_srl_148_n202), .ZN(u1_srl_148_n60) );
  INV_X4 u1_srl_148_U71 ( .A(u1_srl_148_n201), .ZN(u1_srl_148_n59) );
  INV_X4 u1_srl_148_U70 ( .A(u1_srl_148_n248), .ZN(u1_srl_148_n58) );
  INV_X4 u1_srl_148_U69 ( .A(u1_srl_148_n279), .ZN(u1_srl_148_n57) );
  INV_X4 u1_srl_148_U68 ( .A(u1_srl_148_n163), .ZN(u1_srl_148_n56) );
  INV_X4 u1_srl_148_U67 ( .A(u1_srl_148_n200), .ZN(u1_srl_148_n55) );
  INV_X4 u1_srl_148_U66 ( .A(u1_srl_148_n334), .ZN(u1_srl_148_n54) );
  INV_X4 u1_srl_148_U65 ( .A(u1_srl_148_n262), .ZN(u1_srl_148_n53) );
  INV_X4 u1_srl_148_U64 ( .A(u1_srl_148_n176), .ZN(u1_srl_148_n52) );
  INV_X4 u1_srl_148_U63 ( .A(u1_srl_148_n335), .ZN(u1_srl_148_n51) );
  INV_X4 u1_srl_148_U62 ( .A(u1_srl_148_n286), .ZN(u1_srl_148_n50) );
  INV_X4 u1_srl_148_U61 ( .A(u1_srl_148_n336), .ZN(u1_srl_148_n49) );
  INV_X4 u1_srl_148_U60 ( .A(u1_srl_148_n263), .ZN(u1_srl_148_n48) );
  INV_X4 u1_srl_148_U59 ( .A(u1_srl_148_n187), .ZN(u1_srl_148_n47) );
  INV_X4 u1_srl_148_U58 ( .A(u1_srl_148_n190), .ZN(u1_srl_148_n46) );
  INV_X4 u1_srl_148_U57 ( .A(u1_srl_148_n205), .ZN(u1_srl_148_n45) );
  INV_X4 u1_srl_148_U56 ( .A(u1_srl_148_n213), .ZN(u1_srl_148_n44) );
  INV_X4 u1_srl_148_U55 ( .A(u1_srl_148_n295), .ZN(u1_srl_148_n43) );
  INV_X4 u1_srl_148_U54 ( .A(u1_srl_148_n337), .ZN(u1_srl_148_n42) );
  INV_X4 u1_srl_148_U53 ( .A(u1_srl_148_n257), .ZN(u1_srl_148_n41) );
  INV_X4 u1_srl_148_U52 ( .A(u1_srl_148_n170), .ZN(u1_srl_148_n40) );
  INV_X4 u1_srl_148_U51 ( .A(u1_srl_148_n284), .ZN(u1_srl_148_n39) );
  INV_X4 u1_srl_148_U50 ( .A(u1_srl_148_n226), .ZN(u1_srl_148_n38) );
  INV_X4 u1_srl_148_U49 ( .A(u1_srl_148_n348), .ZN(u1_srl_148_n37) );
  INV_X4 u1_srl_148_U48 ( .A(u1_srl_148_n178), .ZN(u1_srl_148_n36) );
  INV_X4 u1_srl_148_U47 ( .A(u1_srl_148_n349), .ZN(u1_srl_148_n35) );
  INV_X4 u1_srl_148_U46 ( .A(u1_srl_148_n241), .ZN(u1_srl_148_n34) );
  INV_X4 u1_srl_148_U45 ( .A(u1_srl_148_n343), .ZN(u1_srl_148_n33) );
  INV_X4 u1_srl_148_U44 ( .A(u1_srl_148_n351), .ZN(u1_srl_148_n32) );
  INV_X4 u1_srl_148_U43 ( .A(u1_srl_148_n312), .ZN(u1_srl_148_n31) );
  INV_X4 u1_srl_148_U42 ( .A(u1_srl_148_n352), .ZN(u1_srl_148_n30) );
  INV_X4 u1_srl_148_U41 ( .A(u1_srl_148_n270), .ZN(u1_srl_148_n29) );
  INV_X4 u1_srl_148_U40 ( .A(u1_srl_148_n155), .ZN(u1_srl_148_n28) );
  INV_X4 u1_srl_148_U39 ( .A(u1_srl_148_n189), .ZN(u1_srl_148_n27) );
  INV_X4 u1_srl_148_U38 ( .A(u1_srl_148_n244), .ZN(u1_srl_148_n26) );
  INV_X4 u1_srl_148_U37 ( .A(u1_srl_148_n209), .ZN(u1_srl_148_n25) );
  INV_X4 u1_srl_148_U36 ( .A(u1_srl_148_n311), .ZN(u1_srl_148_n24) );
  INV_X4 u1_srl_148_U35 ( .A(u1_srl_148_n215), .ZN(u1_srl_148_n23) );
  INV_X4 u1_srl_148_U34 ( .A(u1_srl_148_n356), .ZN(u1_srl_148_n22) );
  INV_X4 u1_srl_148_U33 ( .A(u1_srl_148_n268), .ZN(u1_srl_148_n21) );
  INV_X4 u1_srl_148_U32 ( .A(u1_srl_148_n184), .ZN(u1_srl_148_n20) );
  INV_X4 u1_srl_148_U31 ( .A(u1_srl_148_n289), .ZN(u1_srl_148_n19) );
  INV_X4 u1_srl_148_U30 ( .A(u1_srl_148_n3), .ZN(u1_srl_148_n8) );
  INV_X4 u1_srl_148_U29 ( .A(u1_srl_148_n224), .ZN(u1_srl_148_n5) );
  INV_X4 u1_srl_148_U28 ( .A(u1_srl_148_n13), .ZN(u1_srl_148_n14) );
  INV_X4 u1_srl_148_U27 ( .A(u1_srl_148_n12), .ZN(u1_srl_148_n11) );
  INV_X4 u1_srl_148_U26 ( .A(u1_srl_148_n16), .ZN(u1_srl_148_n15) );
  NOR2_X2 u1_srl_148_U25 ( .A1(u1_srl_148_n1), .A2(u1_srl_148_n8), .ZN(
        u1_srl_148_n138) );
  INV_X4 u1_srl_148_U24 ( .A(u1_srl_148_n195), .ZN(u1_srl_148_n4) );
  INV_X4 u1_srl_148_U23 ( .A(u1_srl_148_n162), .ZN(u1_srl_148_n96) );
  INV_X4 u1_srl_148_U22 ( .A(u1_srl_148_n224), .ZN(u1_srl_148_n6) );
  INV_X4 u1_srl_148_U21 ( .A(u1_srl_148_n1), .ZN(u1_srl_148_n10) );
  INV_X4 u1_srl_148_U20 ( .A(u1_srl_148_n1), .ZN(u1_srl_148_n9) );
  INV_X4 u1_srl_148_U19 ( .A(u1_srl_148_n198), .ZN(u1_srl_148_n16) );
  INV_X4 u1_srl_148_U18 ( .A(u1_srl_148_n3), .ZN(u1_srl_148_n7) );
  INV_X4 u1_srl_148_U17 ( .A(u1_srl_148_n211), .ZN(u1_srl_148_n18) );
  NOR2_X2 u1_srl_148_U16 ( .A1(u1_srl_148_n93), .A2(n6293), .ZN(
        u1_srl_148_n195) );
  INV_X4 u1_srl_148_U15 ( .A(u1_srl_148_n197), .ZN(u1_srl_148_n13) );
  INV_X4 u1_srl_148_U14 ( .A(u1_srl_148_n18), .ZN(u1_srl_148_n17) );
  INV_X4 u1_srl_148_U13 ( .A(u1_srl_148_n2), .ZN(u1_srl_148_n12) );
  NOR2_X2 u1_srl_148_U12 ( .A1(u1_srl_148_n89), .A2(n6285), .ZN(
        u1_srl_148_n224) );
  AND2_X4 u1_srl_148_U11 ( .A1(u1_srl_148_n97), .A2(u1_srl_148_n95), .ZN(
        u1_srl_148_n3) );
  NAND2_X2 u1_srl_148_U10 ( .A1(n6285), .A2(u1_srl_148_n89), .ZN(u1_srl_148_n2) );
  OR2_X4 u1_srl_148_U9 ( .A1(u1_srl_148_n92), .A2(n6301), .ZN(u1_srl_148_n1)
         );
  NOR2_X2 u1_srl_148_U8 ( .A1(u1_srl_148_n95), .A2(n6303), .ZN(u1_srl_148_n144) );
  NOR2_X2 u1_srl_148_U7 ( .A1(u1_srl_148_n18), .A2(u1_srl_148_n7), .ZN(
        u1_srl_148_n145) );
  NOR2_X2 u1_srl_148_U6 ( .A1(u1_srl_148_n7), .A2(u1_srl_148_n91), .ZN(
        u1_srl_148_n140) );
  NOR2_X2 u1_srl_148_U5 ( .A1(u1_srl_148_n4), .A2(u1_srl_148_n7), .ZN(
        u1_srl_148_n142) );
  INV_X4 u1_srl_148_U4 ( .A(u1_srl_148_n237), .ZN(u1_srl_148_n91) );
  NOR2_X2 u1_srl_148_U3 ( .A1(u1_srl_148_n93), .A2(u1_srl_148_n92), .ZN(
        u1_srl_148_n237) );
  INV_X4 sub_1_root_u1_sub_130_aco_U12 ( .A(n4123), .ZN(
        sub_1_root_u1_sub_130_aco_n12) );
  INV_X4 sub_1_root_u1_sub_130_aco_U11 ( .A(n6311), .ZN(
        sub_1_root_u1_sub_130_aco_n11) );
  INV_X4 sub_1_root_u1_sub_130_aco_U10 ( .A(n6310), .ZN(
        sub_1_root_u1_sub_130_aco_n10) );
  INV_X4 sub_1_root_u1_sub_130_aco_U9 ( .A(u1_exp_small[0]), .ZN(
        sub_1_root_u1_sub_130_aco_n9) );
  INV_X4 sub_1_root_u1_sub_130_aco_U8 ( .A(u1_exp_small[10]), .ZN(
        sub_1_root_u1_sub_130_aco_n8) );
  INV_X4 sub_1_root_u1_sub_130_aco_U7 ( .A(u1_exp_small[1]), .ZN(
        sub_1_root_u1_sub_130_aco_n7) );
  INV_X4 sub_1_root_u1_sub_130_aco_U6 ( .A(u1_exp_small[2]), .ZN(
        sub_1_root_u1_sub_130_aco_n6) );
  INV_X4 sub_1_root_u1_sub_130_aco_U5 ( .A(u1_exp_small[3]), .ZN(
        sub_1_root_u1_sub_130_aco_n5) );
  INV_X4 sub_1_root_u1_sub_130_aco_U4 ( .A(u1_exp_small[4]), .ZN(
        sub_1_root_u1_sub_130_aco_n4) );
  INV_X4 sub_1_root_u1_sub_130_aco_U3 ( .A(u1_exp_small[5]), .ZN(
        sub_1_root_u1_sub_130_aco_n3) );
  INV_X4 sub_1_root_u1_sub_130_aco_U2 ( .A(u1_exp_small[6]), .ZN(
        sub_1_root_u1_sub_130_aco_n2) );
  INV_X4 sub_1_root_u1_sub_130_aco_U1 ( .A(u1_exp_small[7]), .ZN(
        sub_1_root_u1_sub_130_aco_n1) );
  FA_X1 sub_1_root_u1_sub_130_aco_U2_0 ( .A(n4156), .B(
        sub_1_root_u1_sub_130_aco_n9), .CI(sub_1_root_u1_sub_130_aco_n12), 
        .CO(sub_1_root_u1_sub_130_aco_carry[1]), .S(u1_exp_diff2[0]) );
  FA_X1 sub_1_root_u1_sub_130_aco_U2_1 ( .A(n4155), .B(
        sub_1_root_u1_sub_130_aco_n7), .CI(sub_1_root_u1_sub_130_aco_carry[1]), 
        .CO(sub_1_root_u1_sub_130_aco_carry[2]), .S(u1_exp_diff2[1]) );
  FA_X1 sub_1_root_u1_sub_130_aco_U2_2 ( .A(n4154), .B(
        sub_1_root_u1_sub_130_aco_n6), .CI(sub_1_root_u1_sub_130_aco_carry[2]), 
        .CO(sub_1_root_u1_sub_130_aco_carry[3]), .S(u1_exp_diff2[2]) );
  FA_X1 sub_1_root_u1_sub_130_aco_U2_3 ( .A(n4153), .B(
        sub_1_root_u1_sub_130_aco_n5), .CI(sub_1_root_u1_sub_130_aco_carry[3]), 
        .CO(sub_1_root_u1_sub_130_aco_carry[4]), .S(u1_exp_diff2[3]) );
  FA_X1 sub_1_root_u1_sub_130_aco_U2_4 ( .A(n4152), .B(
        sub_1_root_u1_sub_130_aco_n4), .CI(sub_1_root_u1_sub_130_aco_carry[4]), 
        .CO(sub_1_root_u1_sub_130_aco_carry[5]), .S(u1_exp_diff2[4]) );
  FA_X1 sub_1_root_u1_sub_130_aco_U2_5 ( .A(n4151), .B(
        sub_1_root_u1_sub_130_aco_n3), .CI(sub_1_root_u1_sub_130_aco_carry[5]), 
        .CO(sub_1_root_u1_sub_130_aco_carry[6]), .S(u1_exp_diff2[5]) );
  FA_X1 sub_1_root_u1_sub_130_aco_U2_6 ( .A(n4150), .B(
        sub_1_root_u1_sub_130_aco_n2), .CI(sub_1_root_u1_sub_130_aco_carry[6]), 
        .CO(sub_1_root_u1_sub_130_aco_carry[7]), .S(u1_exp_diff2[6]) );
  FA_X1 sub_1_root_u1_sub_130_aco_U2_7 ( .A(n4149), .B(
        sub_1_root_u1_sub_130_aco_n1), .CI(sub_1_root_u1_sub_130_aco_carry[7]), 
        .CO(sub_1_root_u1_sub_130_aco_carry[8]), .S(u1_exp_diff2[7]) );
  FA_X1 sub_1_root_u1_sub_130_aco_U2_8 ( .A(n6313), .B(
        sub_1_root_u1_sub_130_aco_n11), .CI(sub_1_root_u1_sub_130_aco_carry[8]), .CO(sub_1_root_u1_sub_130_aco_carry[9]), .S(u1_exp_diff2[8]) );
  FA_X1 sub_1_root_u1_sub_130_aco_U2_9 ( .A(n6312), .B(
        sub_1_root_u1_sub_130_aco_n10), .CI(sub_1_root_u1_sub_130_aco_carry[9]), .CO(sub_1_root_u1_sub_130_aco_carry[10]), .S(u1_exp_diff2[9]) );
  FA_X1 sub_1_root_u1_sub_130_aco_U2_10 ( .A(n4070), .B(
        sub_1_root_u1_sub_130_aco_n8), .CI(sub_1_root_u1_sub_130_aco_carry[10]), .S(u1_exp_diff2[10]) );
  INV_X4 sub_430_3_U171 ( .A(N347), .ZN(sub_430_3_n171) );
  INV_X4 sub_430_3_U170 ( .A(opa_r1[1]), .ZN(sub_430_3_n170) );
  INV_X4 sub_430_3_U169 ( .A(opa_r1[2]), .ZN(sub_430_3_n169) );
  INV_X4 sub_430_3_U168 ( .A(opa_r1[3]), .ZN(sub_430_3_n168) );
  INV_X4 sub_430_3_U167 ( .A(opa_r1[4]), .ZN(sub_430_3_n167) );
  INV_X4 sub_430_3_U166 ( .A(opa_r1[5]), .ZN(sub_430_3_n166) );
  INV_X4 sub_430_3_U165 ( .A(opa_r1[6]), .ZN(sub_430_3_n165) );
  INV_X4 sub_430_3_U164 ( .A(opa_r1[7]), .ZN(sub_430_3_n164) );
  INV_X4 sub_430_3_U163 ( .A(opa_r1[8]), .ZN(sub_430_3_n163) );
  INV_X4 sub_430_3_U162 ( .A(opa_r1[9]), .ZN(sub_430_3_n162) );
  INV_X4 sub_430_3_U161 ( .A(opa_r1[10]), .ZN(sub_430_3_n161) );
  INV_X4 sub_430_3_U160 ( .A(opa_r1[11]), .ZN(sub_430_3_n160) );
  INV_X4 sub_430_3_U159 ( .A(opa_r1[12]), .ZN(sub_430_3_n159) );
  INV_X4 sub_430_3_U158 ( .A(opa_r1[13]), .ZN(sub_430_3_n158) );
  INV_X4 sub_430_3_U157 ( .A(opa_r1[14]), .ZN(sub_430_3_n157) );
  INV_X4 sub_430_3_U156 ( .A(opa_r1[15]), .ZN(sub_430_3_n156) );
  INV_X4 sub_430_3_U155 ( .A(opa_r1[16]), .ZN(sub_430_3_n155) );
  INV_X4 sub_430_3_U154 ( .A(opa_r1[17]), .ZN(sub_430_3_n154) );
  INV_X4 sub_430_3_U153 ( .A(opa_r1[18]), .ZN(sub_430_3_n153) );
  INV_X4 sub_430_3_U152 ( .A(opa_r1[19]), .ZN(sub_430_3_n152) );
  INV_X4 sub_430_3_U151 ( .A(opa_r1[20]), .ZN(sub_430_3_n151) );
  INV_X4 sub_430_3_U150 ( .A(opa_r1[21]), .ZN(sub_430_3_n150) );
  INV_X4 sub_430_3_U149 ( .A(opa_r1[22]), .ZN(sub_430_3_n149) );
  INV_X4 sub_430_3_U148 ( .A(opa_r1[23]), .ZN(sub_430_3_n148) );
  INV_X4 sub_430_3_U147 ( .A(opa_r1[24]), .ZN(sub_430_3_n147) );
  INV_X4 sub_430_3_U146 ( .A(opa_r1[25]), .ZN(sub_430_3_n146) );
  INV_X4 sub_430_3_U145 ( .A(opa_r1[26]), .ZN(sub_430_3_n145) );
  INV_X4 sub_430_3_U144 ( .A(opa_r1[27]), .ZN(sub_430_3_n144) );
  INV_X4 sub_430_3_U143 ( .A(opa_r1[28]), .ZN(sub_430_3_n143) );
  INV_X4 sub_430_3_U142 ( .A(opa_r1[29]), .ZN(sub_430_3_n142) );
  INV_X4 sub_430_3_U141 ( .A(opa_r1[30]), .ZN(sub_430_3_n141) );
  INV_X4 sub_430_3_U140 ( .A(opa_r1[31]), .ZN(sub_430_3_n140) );
  INV_X4 sub_430_3_U139 ( .A(opa_r1[32]), .ZN(sub_430_3_n139) );
  INV_X4 sub_430_3_U138 ( .A(opa_r1[33]), .ZN(sub_430_3_n138) );
  INV_X4 sub_430_3_U137 ( .A(opa_r1[34]), .ZN(sub_430_3_n137) );
  INV_X4 sub_430_3_U136 ( .A(opa_r1[35]), .ZN(sub_430_3_n136) );
  INV_X4 sub_430_3_U135 ( .A(opa_r1[36]), .ZN(sub_430_3_n135) );
  INV_X4 sub_430_3_U134 ( .A(opa_r1[37]), .ZN(sub_430_3_n134) );
  INV_X4 sub_430_3_U133 ( .A(opa_r1[38]), .ZN(sub_430_3_n133) );
  INV_X4 sub_430_3_U132 ( .A(opa_r1[39]), .ZN(sub_430_3_n132) );
  INV_X4 sub_430_3_U131 ( .A(opa_r1[40]), .ZN(sub_430_3_n131) );
  INV_X4 sub_430_3_U130 ( .A(opa_r1[41]), .ZN(sub_430_3_n130) );
  INV_X4 sub_430_3_U129 ( .A(opa_r1[42]), .ZN(sub_430_3_n129) );
  INV_X4 sub_430_3_U128 ( .A(opa_r1[43]), .ZN(sub_430_3_n128) );
  INV_X4 sub_430_3_U127 ( .A(opa_r1[44]), .ZN(sub_430_3_n127) );
  INV_X4 sub_430_3_U126 ( .A(opa_r1[45]), .ZN(sub_430_3_n126) );
  INV_X4 sub_430_3_U125 ( .A(opa_r1[46]), .ZN(sub_430_3_n125) );
  INV_X4 sub_430_3_U124 ( .A(opa_r1[47]), .ZN(sub_430_3_n124) );
  INV_X4 sub_430_3_U123 ( .A(opa_r1[48]), .ZN(sub_430_3_n123) );
  INV_X4 sub_430_3_U122 ( .A(opa_r1[49]), .ZN(sub_430_3_n122) );
  INV_X4 sub_430_3_U121 ( .A(opa_r1[50]), .ZN(sub_430_3_n121) );
  INV_X4 sub_430_3_U120 ( .A(opa_r1[51]), .ZN(sub_430_3_n120) );
  INV_X4 sub_430_3_U119 ( .A(opa_r1[52]), .ZN(sub_430_3_n119) );
  INV_X4 sub_430_3_U118 ( .A(opa_r1[53]), .ZN(sub_430_3_n118) );
  INV_X4 sub_430_3_U117 ( .A(opa_r1[54]), .ZN(sub_430_3_n117) );
  INV_X4 sub_430_3_U116 ( .A(opa_r1[55]), .ZN(sub_430_3_n116) );
  INV_X4 sub_430_3_U115 ( .A(opa_r1[56]), .ZN(sub_430_3_n115) );
  INV_X4 sub_430_3_U114 ( .A(opa_r1[57]), .ZN(sub_430_3_n114) );
  XOR2_X2 sub_430_3_U113 ( .A(sub_430_3_n159), .B(sub_430_3_n40), .Z(N516) );
  XOR2_X2 sub_430_3_U112 ( .A(sub_430_3_n160), .B(sub_430_3_n35), .Z(N515) );
  XOR2_X2 sub_430_3_U111 ( .A(sub_430_3_n161), .B(sub_430_3_n13), .Z(N514) );
  XOR2_X2 sub_430_3_U110 ( .A(sub_430_3_n162), .B(sub_430_3_n36), .Z(N513) );
  XOR2_X2 sub_430_3_U109 ( .A(sub_430_3_n163), .B(sub_430_3_n14), .Z(N512) );
  XOR2_X2 sub_430_3_U108 ( .A(sub_430_3_n164), .B(sub_430_3_n37), .Z(N511) );
  XOR2_X2 sub_430_3_U107 ( .A(sub_430_3_n166), .B(sub_430_3_n38), .Z(N509) );
  XOR2_X2 sub_430_3_U106 ( .A(sub_430_3_n168), .B(sub_430_3_n39), .Z(N507) );
  XOR2_X2 sub_430_3_U105 ( .A(sub_430_3_n165), .B(sub_430_3_n15), .Z(N510) );
  XOR2_X2 sub_430_3_U104 ( .A(sub_430_3_n167), .B(sub_430_3_n16), .Z(N508) );
  XOR2_X2 sub_430_3_U103 ( .A(sub_430_3_n121), .B(sub_430_3_n41), .Z(N554) );
  AND2_X4 sub_430_3_U102 ( .A1(sub_430_3_n115), .A2(sub_430_3_n43), .ZN(
        sub_430_3_n102) );
  AND2_X4 sub_430_3_U101 ( .A1(sub_430_3_n119), .A2(sub_430_3_n12), .ZN(
        sub_430_3_n101) );
  AND2_X4 sub_430_3_U100 ( .A1(sub_430_3_n117), .A2(sub_430_3_n46), .ZN(
        sub_430_3_n100) );
  AND2_X4 sub_430_3_U99 ( .A1(sub_430_3_n170), .A2(sub_430_3_n171), .ZN(
        sub_430_3_n99) );
  AND2_X4 sub_430_3_U98 ( .A1(sub_430_3_n159), .A2(sub_430_3_n40), .ZN(
        sub_430_3_n98) );
  AND2_X4 sub_430_3_U97 ( .A1(sub_430_3_n157), .A2(sub_430_3_n17), .ZN(
        sub_430_3_n97) );
  AND2_X4 sub_430_3_U96 ( .A1(sub_430_3_n155), .A2(sub_430_3_n31), .ZN(
        sub_430_3_n96) );
  AND2_X4 sub_430_3_U95 ( .A1(sub_430_3_n153), .A2(sub_430_3_n30), .ZN(
        sub_430_3_n95) );
  AND2_X4 sub_430_3_U94 ( .A1(sub_430_3_n151), .A2(sub_430_3_n29), .ZN(
        sub_430_3_n94) );
  AND2_X4 sub_430_3_U93 ( .A1(sub_430_3_n149), .A2(sub_430_3_n28), .ZN(
        sub_430_3_n93) );
  AND2_X4 sub_430_3_U92 ( .A1(sub_430_3_n147), .A2(sub_430_3_n27), .ZN(
        sub_430_3_n92) );
  AND2_X4 sub_430_3_U91 ( .A1(sub_430_3_n145), .A2(sub_430_3_n26), .ZN(
        sub_430_3_n91) );
  AND2_X4 sub_430_3_U90 ( .A1(sub_430_3_n143), .A2(sub_430_3_n25), .ZN(
        sub_430_3_n90) );
  AND2_X4 sub_430_3_U89 ( .A1(sub_430_3_n141), .A2(sub_430_3_n24), .ZN(
        sub_430_3_n89) );
  AND2_X4 sub_430_3_U88 ( .A1(sub_430_3_n139), .A2(sub_430_3_n23), .ZN(
        sub_430_3_n88) );
  AND2_X4 sub_430_3_U87 ( .A1(sub_430_3_n137), .A2(sub_430_3_n22), .ZN(
        sub_430_3_n87) );
  AND2_X4 sub_430_3_U86 ( .A1(sub_430_3_n135), .A2(sub_430_3_n21), .ZN(
        sub_430_3_n86) );
  AND2_X4 sub_430_3_U85 ( .A1(sub_430_3_n133), .A2(sub_430_3_n20), .ZN(
        sub_430_3_n85) );
  AND2_X4 sub_430_3_U84 ( .A1(sub_430_3_n131), .A2(sub_430_3_n19), .ZN(
        sub_430_3_n84) );
  AND2_X4 sub_430_3_U83 ( .A1(sub_430_3_n129), .A2(sub_430_3_n18), .ZN(
        sub_430_3_n83) );
  AND2_X4 sub_430_3_U82 ( .A1(sub_430_3_n127), .A2(sub_430_3_n45), .ZN(
        sub_430_3_n82) );
  AND2_X4 sub_430_3_U81 ( .A1(sub_430_3_n125), .A2(sub_430_3_n44), .ZN(
        sub_430_3_n81) );
  AND2_X4 sub_430_3_U80 ( .A1(sub_430_3_n123), .A2(sub_430_3_n42), .ZN(
        sub_430_3_n80) );
  AND2_X4 sub_430_3_U79 ( .A1(sub_430_3_n121), .A2(sub_430_3_n41), .ZN(
        sub_430_3_n79) );
  XOR2_X2 sub_430_3_U78 ( .A(sub_430_3_n141), .B(sub_430_3_n24), .Z(N534) );
  XOR2_X2 sub_430_3_U77 ( .A(sub_430_3_n142), .B(sub_430_3_n90), .Z(N533) );
  XOR2_X2 sub_430_3_U76 ( .A(sub_430_3_n144), .B(sub_430_3_n91), .Z(N531) );
  XOR2_X2 sub_430_3_U75 ( .A(sub_430_3_n147), .B(sub_430_3_n27), .Z(N528) );
  XOR2_X2 sub_430_3_U74 ( .A(sub_430_3_n149), .B(sub_430_3_n28), .Z(N526) );
  XOR2_X2 sub_430_3_U73 ( .A(sub_430_3_n150), .B(sub_430_3_n94), .Z(N525) );
  XOR2_X2 sub_430_3_U72 ( .A(sub_430_3_n151), .B(sub_430_3_n29), .Z(N524) );
  XOR2_X2 sub_430_3_U71 ( .A(sub_430_3_n152), .B(sub_430_3_n95), .Z(N523) );
  XOR2_X2 sub_430_3_U70 ( .A(sub_430_3_n154), .B(sub_430_3_n96), .Z(N521) );
  XOR2_X2 sub_430_3_U69 ( .A(sub_430_3_n157), .B(sub_430_3_n17), .Z(N518) );
  XOR2_X2 sub_430_3_U68 ( .A(sub_430_3_n143), .B(sub_430_3_n25), .Z(N532) );
  XOR2_X2 sub_430_3_U67 ( .A(sub_430_3_n145), .B(sub_430_3_n26), .Z(N530) );
  XOR2_X2 sub_430_3_U66 ( .A(sub_430_3_n146), .B(sub_430_3_n92), .Z(N529) );
  XOR2_X2 sub_430_3_U65 ( .A(sub_430_3_n148), .B(sub_430_3_n93), .Z(N527) );
  XOR2_X2 sub_430_3_U64 ( .A(sub_430_3_n153), .B(sub_430_3_n30), .Z(N522) );
  XOR2_X2 sub_430_3_U63 ( .A(sub_430_3_n155), .B(sub_430_3_n31), .Z(N520) );
  XOR2_X2 sub_430_3_U62 ( .A(sub_430_3_n156), .B(sub_430_3_n97), .Z(N519) );
  XOR2_X2 sub_430_3_U61 ( .A(sub_430_3_n128), .B(sub_430_3_n83), .Z(N547) );
  XOR2_X2 sub_430_3_U60 ( .A(sub_430_3_n129), .B(sub_430_3_n18), .Z(N546) );
  XOR2_X2 sub_430_3_U59 ( .A(sub_430_3_n131), .B(sub_430_3_n19), .Z(N544) );
  XOR2_X2 sub_430_3_U58 ( .A(sub_430_3_n133), .B(sub_430_3_n20), .Z(N542) );
  XOR2_X2 sub_430_3_U57 ( .A(sub_430_3_n134), .B(sub_430_3_n86), .Z(N541) );
  XOR2_X2 sub_430_3_U56 ( .A(sub_430_3_n135), .B(sub_430_3_n21), .Z(N540) );
  XOR2_X2 sub_430_3_U55 ( .A(sub_430_3_n136), .B(sub_430_3_n87), .Z(N539) );
  XOR2_X2 sub_430_3_U54 ( .A(sub_430_3_n139), .B(sub_430_3_n23), .Z(N536) );
  XOR2_X2 sub_430_3_U53 ( .A(sub_430_3_n140), .B(sub_430_3_n89), .Z(N535) );
  XOR2_X2 sub_430_3_U52 ( .A(sub_430_3_n130), .B(sub_430_3_n84), .Z(N545) );
  XOR2_X2 sub_430_3_U51 ( .A(sub_430_3_n132), .B(sub_430_3_n85), .Z(N543) );
  XOR2_X2 sub_430_3_U50 ( .A(sub_430_3_n137), .B(sub_430_3_n22), .Z(N538) );
  XOR2_X2 sub_430_3_U49 ( .A(sub_430_3_n138), .B(sub_430_3_n88), .Z(N537) );
  XOR2_X2 sub_430_3_U48 ( .A(sub_430_3_n120), .B(sub_430_3_n79), .Z(N555) );
  XOR2_X2 sub_430_3_U47 ( .A(sub_430_3_n119), .B(sub_430_3_n12), .Z(N556) );
  AND2_X4 sub_430_3_U46 ( .A1(sub_430_3_n118), .A2(sub_430_3_n101), .ZN(
        sub_430_3_n46) );
  AND2_X4 sub_430_3_U45 ( .A1(sub_430_3_n128), .A2(sub_430_3_n83), .ZN(
        sub_430_3_n45) );
  AND2_X4 sub_430_3_U44 ( .A1(sub_430_3_n126), .A2(sub_430_3_n82), .ZN(
        sub_430_3_n44) );
  AND2_X4 sub_430_3_U43 ( .A1(sub_430_3_n116), .A2(sub_430_3_n100), .ZN(
        sub_430_3_n43) );
  AND2_X4 sub_430_3_U42 ( .A1(sub_430_3_n124), .A2(sub_430_3_n81), .ZN(
        sub_430_3_n42) );
  AND2_X4 sub_430_3_U41 ( .A1(sub_430_3_n122), .A2(sub_430_3_n80), .ZN(
        sub_430_3_n41) );
  AND2_X4 sub_430_3_U40 ( .A1(sub_430_3_n160), .A2(sub_430_3_n35), .ZN(
        sub_430_3_n40) );
  AND2_X4 sub_430_3_U39 ( .A1(sub_430_3_n169), .A2(sub_430_3_n99), .ZN(
        sub_430_3_n39) );
  AND2_X4 sub_430_3_U38 ( .A1(sub_430_3_n167), .A2(sub_430_3_n16), .ZN(
        sub_430_3_n38) );
  AND2_X4 sub_430_3_U37 ( .A1(sub_430_3_n165), .A2(sub_430_3_n15), .ZN(
        sub_430_3_n37) );
  AND2_X4 sub_430_3_U36 ( .A1(sub_430_3_n163), .A2(sub_430_3_n14), .ZN(
        sub_430_3_n36) );
  AND2_X4 sub_430_3_U35 ( .A1(sub_430_3_n161), .A2(sub_430_3_n13), .ZN(
        sub_430_3_n35) );
  XOR2_X2 sub_430_3_U34 ( .A(sub_430_3_n169), .B(sub_430_3_n99), .Z(N506) );
  XOR2_X2 sub_430_3_U33 ( .A(sub_430_3_n170), .B(sub_430_3_n171), .Z(N505) );
  XOR2_X2 sub_430_3_U32 ( .A(sub_430_3_n158), .B(sub_430_3_n98), .Z(N517) );
  AND2_X4 sub_430_3_U31 ( .A1(sub_430_3_n156), .A2(sub_430_3_n97), .ZN(
        sub_430_3_n31) );
  AND2_X4 sub_430_3_U30 ( .A1(sub_430_3_n154), .A2(sub_430_3_n96), .ZN(
        sub_430_3_n30) );
  AND2_X4 sub_430_3_U29 ( .A1(sub_430_3_n152), .A2(sub_430_3_n95), .ZN(
        sub_430_3_n29) );
  AND2_X4 sub_430_3_U28 ( .A1(sub_430_3_n150), .A2(sub_430_3_n94), .ZN(
        sub_430_3_n28) );
  AND2_X4 sub_430_3_U27 ( .A1(sub_430_3_n148), .A2(sub_430_3_n93), .ZN(
        sub_430_3_n27) );
  AND2_X4 sub_430_3_U26 ( .A1(sub_430_3_n146), .A2(sub_430_3_n92), .ZN(
        sub_430_3_n26) );
  AND2_X4 sub_430_3_U25 ( .A1(sub_430_3_n144), .A2(sub_430_3_n91), .ZN(
        sub_430_3_n25) );
  AND2_X4 sub_430_3_U24 ( .A1(sub_430_3_n142), .A2(sub_430_3_n90), .ZN(
        sub_430_3_n24) );
  AND2_X4 sub_430_3_U23 ( .A1(sub_430_3_n140), .A2(sub_430_3_n89), .ZN(
        sub_430_3_n23) );
  AND2_X4 sub_430_3_U22 ( .A1(sub_430_3_n138), .A2(sub_430_3_n88), .ZN(
        sub_430_3_n22) );
  AND2_X4 sub_430_3_U21 ( .A1(sub_430_3_n136), .A2(sub_430_3_n87), .ZN(
        sub_430_3_n21) );
  AND2_X4 sub_430_3_U20 ( .A1(sub_430_3_n134), .A2(sub_430_3_n86), .ZN(
        sub_430_3_n20) );
  AND2_X4 sub_430_3_U19 ( .A1(sub_430_3_n132), .A2(sub_430_3_n85), .ZN(
        sub_430_3_n19) );
  AND2_X4 sub_430_3_U18 ( .A1(sub_430_3_n130), .A2(sub_430_3_n84), .ZN(
        sub_430_3_n18) );
  AND2_X4 sub_430_3_U17 ( .A1(sub_430_3_n158), .A2(sub_430_3_n98), .ZN(
        sub_430_3_n17) );
  AND2_X4 sub_430_3_U16 ( .A1(sub_430_3_n168), .A2(sub_430_3_n39), .ZN(
        sub_430_3_n16) );
  AND2_X4 sub_430_3_U15 ( .A1(sub_430_3_n166), .A2(sub_430_3_n38), .ZN(
        sub_430_3_n15) );
  AND2_X4 sub_430_3_U14 ( .A1(sub_430_3_n164), .A2(sub_430_3_n37), .ZN(
        sub_430_3_n14) );
  AND2_X4 sub_430_3_U13 ( .A1(sub_430_3_n162), .A2(sub_430_3_n36), .ZN(
        sub_430_3_n13) );
  AND2_X4 sub_430_3_U12 ( .A1(sub_430_3_n120), .A2(sub_430_3_n79), .ZN(
        sub_430_3_n12) );
  XOR2_X2 sub_430_3_U11 ( .A(sub_430_3_n125), .B(sub_430_3_n44), .Z(N550) );
  XOR2_X2 sub_430_3_U10 ( .A(sub_430_3_n127), .B(sub_430_3_n45), .Z(N548) );
  XOR2_X2 sub_430_3_U9 ( .A(sub_430_3_n114), .B(sub_430_3_n102), .Z(N561) );
  XOR2_X2 sub_430_3_U8 ( .A(sub_430_3_n126), .B(sub_430_3_n82), .Z(N549) );
  XOR2_X2 sub_430_3_U7 ( .A(sub_430_3_n115), .B(sub_430_3_n43), .Z(N560) );
  XOR2_X2 sub_430_3_U6 ( .A(sub_430_3_n117), .B(sub_430_3_n46), .Z(N558) );
  XOR2_X2 sub_430_3_U5 ( .A(sub_430_3_n122), .B(sub_430_3_n80), .Z(N553) );
  XOR2_X2 sub_430_3_U4 ( .A(sub_430_3_n123), .B(sub_430_3_n42), .Z(N552) );
  XOR2_X2 sub_430_3_U3 ( .A(sub_430_3_n124), .B(sub_430_3_n81), .Z(N551) );
  XOR2_X2 sub_430_3_U2 ( .A(sub_430_3_n118), .B(sub_430_3_n101), .Z(N557) );
  XOR2_X2 sub_430_3_U1 ( .A(sub_430_3_n116), .B(sub_430_3_n100), .Z(N559) );
  INV_X4 sub_430_b0_U157 ( .A(N347), .ZN(sub_430_b0_n157) );
  INV_X4 sub_430_b0_U156 ( .A(opa_r1[1]), .ZN(sub_430_b0_n156) );
  INV_X4 sub_430_b0_U155 ( .A(opa_r1[2]), .ZN(sub_430_b0_n155) );
  INV_X4 sub_430_b0_U154 ( .A(opa_r1[3]), .ZN(sub_430_b0_n154) );
  INV_X4 sub_430_b0_U153 ( .A(opa_r1[4]), .ZN(sub_430_b0_n153) );
  INV_X4 sub_430_b0_U152 ( .A(opa_r1[5]), .ZN(sub_430_b0_n152) );
  INV_X4 sub_430_b0_U151 ( .A(opa_r1[6]), .ZN(sub_430_b0_n151) );
  INV_X4 sub_430_b0_U150 ( .A(opa_r1[7]), .ZN(sub_430_b0_n150) );
  INV_X4 sub_430_b0_U149 ( .A(opa_r1[8]), .ZN(sub_430_b0_n149) );
  INV_X4 sub_430_b0_U148 ( .A(opa_r1[9]), .ZN(sub_430_b0_n148) );
  INV_X4 sub_430_b0_U147 ( .A(opa_r1[10]), .ZN(sub_430_b0_n147) );
  INV_X4 sub_430_b0_U146 ( .A(opa_r1[11]), .ZN(sub_430_b0_n146) );
  INV_X4 sub_430_b0_U145 ( .A(opa_r1[12]), .ZN(sub_430_b0_n145) );
  INV_X4 sub_430_b0_U144 ( .A(opa_r1[13]), .ZN(sub_430_b0_n144) );
  INV_X4 sub_430_b0_U143 ( .A(opa_r1[14]), .ZN(sub_430_b0_n143) );
  INV_X4 sub_430_b0_U142 ( .A(opa_r1[15]), .ZN(sub_430_b0_n142) );
  INV_X4 sub_430_b0_U141 ( .A(opa_r1[16]), .ZN(sub_430_b0_n141) );
  INV_X4 sub_430_b0_U140 ( .A(opa_r1[17]), .ZN(sub_430_b0_n140) );
  INV_X4 sub_430_b0_U139 ( .A(opa_r1[18]), .ZN(sub_430_b0_n139) );
  INV_X4 sub_430_b0_U138 ( .A(opa_r1[19]), .ZN(sub_430_b0_n138) );
  INV_X4 sub_430_b0_U137 ( .A(opa_r1[20]), .ZN(sub_430_b0_n137) );
  INV_X4 sub_430_b0_U136 ( .A(opa_r1[21]), .ZN(sub_430_b0_n136) );
  INV_X4 sub_430_b0_U135 ( .A(opa_r1[22]), .ZN(sub_430_b0_n135) );
  INV_X4 sub_430_b0_U134 ( .A(opa_r1[23]), .ZN(sub_430_b0_n134) );
  INV_X4 sub_430_b0_U133 ( .A(opa_r1[24]), .ZN(sub_430_b0_n133) );
  INV_X4 sub_430_b0_U132 ( .A(opa_r1[25]), .ZN(sub_430_b0_n132) );
  INV_X4 sub_430_b0_U131 ( .A(opa_r1[26]), .ZN(sub_430_b0_n131) );
  INV_X4 sub_430_b0_U130 ( .A(opa_r1[27]), .ZN(sub_430_b0_n130) );
  INV_X4 sub_430_b0_U129 ( .A(opa_r1[28]), .ZN(sub_430_b0_n129) );
  INV_X4 sub_430_b0_U128 ( .A(opa_r1[29]), .ZN(sub_430_b0_n128) );
  INV_X4 sub_430_b0_U127 ( .A(opa_r1[30]), .ZN(sub_430_b0_n127) );
  INV_X4 sub_430_b0_U126 ( .A(opa_r1[31]), .ZN(sub_430_b0_n126) );
  INV_X4 sub_430_b0_U125 ( .A(opa_r1[32]), .ZN(sub_430_b0_n125) );
  INV_X4 sub_430_b0_U124 ( .A(opa_r1[33]), .ZN(sub_430_b0_n124) );
  INV_X4 sub_430_b0_U123 ( .A(opa_r1[34]), .ZN(sub_430_b0_n123) );
  INV_X4 sub_430_b0_U122 ( .A(opa_r1[35]), .ZN(sub_430_b0_n122) );
  INV_X4 sub_430_b0_U121 ( .A(opa_r1[36]), .ZN(sub_430_b0_n121) );
  INV_X4 sub_430_b0_U120 ( .A(opa_r1[37]), .ZN(sub_430_b0_n120) );
  INV_X4 sub_430_b0_U119 ( .A(opa_r1[38]), .ZN(sub_430_b0_n119) );
  INV_X4 sub_430_b0_U118 ( .A(opa_r1[39]), .ZN(sub_430_b0_n118) );
  INV_X4 sub_430_b0_U117 ( .A(opa_r1[40]), .ZN(sub_430_b0_n117) );
  INV_X4 sub_430_b0_U116 ( .A(opa_r1[41]), .ZN(sub_430_b0_n116) );
  INV_X4 sub_430_b0_U115 ( .A(opa_r1[42]), .ZN(sub_430_b0_n115) );
  INV_X4 sub_430_b0_U114 ( .A(opa_r1[43]), .ZN(sub_430_b0_n114) );
  INV_X4 sub_430_b0_U113 ( .A(opa_r1[44]), .ZN(sub_430_b0_n113) );
  INV_X4 sub_430_b0_U112 ( .A(opa_r1[45]), .ZN(sub_430_b0_n112) );
  INV_X4 sub_430_b0_U111 ( .A(opa_r1[46]), .ZN(sub_430_b0_n111) );
  INV_X4 sub_430_b0_U110 ( .A(opa_r1[47]), .ZN(sub_430_b0_n110) );
  INV_X4 sub_430_b0_U109 ( .A(opa_r1[48]), .ZN(sub_430_b0_n109) );
  INV_X4 sub_430_b0_U108 ( .A(opa_r1[49]), .ZN(sub_430_b0_n108) );
  INV_X4 sub_430_b0_U107 ( .A(opa_r1[50]), .ZN(sub_430_b0_n107) );
  INV_X4 sub_430_b0_U106 ( .A(opa_r1[51]), .ZN(sub_430_b0_n106) );
  INV_X4 sub_430_b0_U105 ( .A(N342), .ZN(sub_430_b0_n105) );
  NAND2_X2 sub_430_b0_U104 ( .A1(sub_430_b0_n105), .A2(sub_430_b0_n43), .ZN(
        N400) );
  XOR2_X2 sub_430_b0_U103 ( .A(sub_430_b0_n144), .B(sub_430_b0_n2), .Z(N360)
         );
  XOR2_X2 sub_430_b0_U102 ( .A(sub_430_b0_n145), .B(sub_430_b0_n63), .Z(N359)
         );
  XOR2_X2 sub_430_b0_U101 ( .A(sub_430_b0_n146), .B(sub_430_b0_n3), .Z(N358)
         );
  XOR2_X2 sub_430_b0_U100 ( .A(sub_430_b0_n147), .B(sub_430_b0_n64), .Z(N357)
         );
  XOR2_X2 sub_430_b0_U99 ( .A(sub_430_b0_n148), .B(sub_430_b0_n4), .Z(N356) );
  XOR2_X2 sub_430_b0_U98 ( .A(sub_430_b0_n122), .B(sub_430_b0_n9), .Z(N382) );
  XOR2_X2 sub_430_b0_U97 ( .A(sub_430_b0_n123), .B(sub_430_b0_n52), .Z(N381)
         );
  XOR2_X2 sub_430_b0_U96 ( .A(sub_430_b0_n124), .B(sub_430_b0_n10), .Z(N380)
         );
  XOR2_X2 sub_430_b0_U95 ( .A(sub_430_b0_n125), .B(sub_430_b0_n53), .Z(N379)
         );
  XOR2_X2 sub_430_b0_U94 ( .A(sub_430_b0_n126), .B(sub_430_b0_n11), .Z(N378)
         );
  XOR2_X2 sub_430_b0_U93 ( .A(sub_430_b0_n127), .B(sub_430_b0_n54), .Z(N377)
         );
  XOR2_X2 sub_430_b0_U92 ( .A(sub_430_b0_n128), .B(sub_430_b0_n12), .Z(N376)
         );
  XOR2_X2 sub_430_b0_U91 ( .A(sub_430_b0_n129), .B(sub_430_b0_n55), .Z(N375)
         );
  XOR2_X2 sub_430_b0_U90 ( .A(sub_430_b0_n130), .B(sub_430_b0_n13), .Z(N374)
         );
  XOR2_X2 sub_430_b0_U89 ( .A(sub_430_b0_n131), .B(sub_430_b0_n56), .Z(N373)
         );
  XOR2_X2 sub_430_b0_U88 ( .A(sub_430_b0_n132), .B(sub_430_b0_n14), .Z(N372)
         );
  XOR2_X2 sub_430_b0_U87 ( .A(sub_430_b0_n133), .B(sub_430_b0_n57), .Z(N371)
         );
  XOR2_X2 sub_430_b0_U86 ( .A(sub_430_b0_n134), .B(sub_430_b0_n15), .Z(N370)
         );
  XOR2_X2 sub_430_b0_U85 ( .A(sub_430_b0_n135), .B(sub_430_b0_n58), .Z(N369)
         );
  XOR2_X2 sub_430_b0_U84 ( .A(sub_430_b0_n136), .B(sub_430_b0_n16), .Z(N368)
         );
  XOR2_X2 sub_430_b0_U83 ( .A(sub_430_b0_n137), .B(sub_430_b0_n59), .Z(N367)
         );
  XOR2_X2 sub_430_b0_U82 ( .A(sub_430_b0_n138), .B(sub_430_b0_n17), .Z(N366)
         );
  XOR2_X2 sub_430_b0_U81 ( .A(sub_430_b0_n139), .B(sub_430_b0_n60), .Z(N365)
         );
  XOR2_X2 sub_430_b0_U80 ( .A(sub_430_b0_n140), .B(sub_430_b0_n18), .Z(N364)
         );
  XOR2_X2 sub_430_b0_U79 ( .A(sub_430_b0_n141), .B(sub_430_b0_n61), .Z(N363)
         );
  XOR2_X2 sub_430_b0_U78 ( .A(sub_430_b0_n142), .B(sub_430_b0_n1), .Z(N362) );
  XOR2_X2 sub_430_b0_U77 ( .A(sub_430_b0_n143), .B(sub_430_b0_n62), .Z(N361)
         );
  XOR2_X2 sub_430_b0_U76 ( .A(sub_430_b0_n114), .B(sub_430_b0_n5), .Z(N390) );
  XOR2_X2 sub_430_b0_U75 ( .A(sub_430_b0_n115), .B(sub_430_b0_n48), .Z(N389)
         );
  XOR2_X2 sub_430_b0_U74 ( .A(sub_430_b0_n116), .B(sub_430_b0_n6), .Z(N388) );
  XOR2_X2 sub_430_b0_U73 ( .A(sub_430_b0_n117), .B(sub_430_b0_n49), .Z(N387)
         );
  XOR2_X2 sub_430_b0_U72 ( .A(sub_430_b0_n118), .B(sub_430_b0_n7), .Z(N386) );
  XOR2_X2 sub_430_b0_U71 ( .A(sub_430_b0_n119), .B(sub_430_b0_n50), .Z(N385)
         );
  XOR2_X2 sub_430_b0_U70 ( .A(sub_430_b0_n120), .B(sub_430_b0_n8), .Z(N384) );
  XOR2_X2 sub_430_b0_U69 ( .A(sub_430_b0_n121), .B(sub_430_b0_n51), .Z(N383)
         );
  AND2_X4 sub_430_b0_U68 ( .A1(sub_430_b0_n156), .A2(sub_430_b0_n157), .ZN(
        sub_430_b0_n68) );
  AND2_X4 sub_430_b0_U67 ( .A1(sub_430_b0_n154), .A2(sub_430_b0_n24), .ZN(
        sub_430_b0_n67) );
  AND2_X4 sub_430_b0_U66 ( .A1(sub_430_b0_n152), .A2(sub_430_b0_n23), .ZN(
        sub_430_b0_n66) );
  AND2_X4 sub_430_b0_U65 ( .A1(sub_430_b0_n150), .A2(sub_430_b0_n22), .ZN(
        sub_430_b0_n65) );
  AND2_X4 sub_430_b0_U64 ( .A1(sub_430_b0_n148), .A2(sub_430_b0_n4), .ZN(
        sub_430_b0_n64) );
  AND2_X4 sub_430_b0_U63 ( .A1(sub_430_b0_n146), .A2(sub_430_b0_n3), .ZN(
        sub_430_b0_n63) );
  AND2_X4 sub_430_b0_U62 ( .A1(sub_430_b0_n144), .A2(sub_430_b0_n2), .ZN(
        sub_430_b0_n62) );
  AND2_X4 sub_430_b0_U61 ( .A1(sub_430_b0_n142), .A2(sub_430_b0_n1), .ZN(
        sub_430_b0_n61) );
  AND2_X4 sub_430_b0_U60 ( .A1(sub_430_b0_n140), .A2(sub_430_b0_n18), .ZN(
        sub_430_b0_n60) );
  AND2_X4 sub_430_b0_U59 ( .A1(sub_430_b0_n138), .A2(sub_430_b0_n17), .ZN(
        sub_430_b0_n59) );
  AND2_X4 sub_430_b0_U58 ( .A1(sub_430_b0_n136), .A2(sub_430_b0_n16), .ZN(
        sub_430_b0_n58) );
  AND2_X4 sub_430_b0_U57 ( .A1(sub_430_b0_n134), .A2(sub_430_b0_n15), .ZN(
        sub_430_b0_n57) );
  AND2_X4 sub_430_b0_U56 ( .A1(sub_430_b0_n132), .A2(sub_430_b0_n14), .ZN(
        sub_430_b0_n56) );
  AND2_X4 sub_430_b0_U55 ( .A1(sub_430_b0_n130), .A2(sub_430_b0_n13), .ZN(
        sub_430_b0_n55) );
  AND2_X4 sub_430_b0_U54 ( .A1(sub_430_b0_n128), .A2(sub_430_b0_n12), .ZN(
        sub_430_b0_n54) );
  AND2_X4 sub_430_b0_U53 ( .A1(sub_430_b0_n126), .A2(sub_430_b0_n11), .ZN(
        sub_430_b0_n53) );
  AND2_X4 sub_430_b0_U52 ( .A1(sub_430_b0_n124), .A2(sub_430_b0_n10), .ZN(
        sub_430_b0_n52) );
  AND2_X4 sub_430_b0_U51 ( .A1(sub_430_b0_n122), .A2(sub_430_b0_n9), .ZN(
        sub_430_b0_n51) );
  AND2_X4 sub_430_b0_U50 ( .A1(sub_430_b0_n120), .A2(sub_430_b0_n8), .ZN(
        sub_430_b0_n50) );
  AND2_X4 sub_430_b0_U49 ( .A1(sub_430_b0_n118), .A2(sub_430_b0_n7), .ZN(
        sub_430_b0_n49) );
  AND2_X4 sub_430_b0_U48 ( .A1(sub_430_b0_n116), .A2(sub_430_b0_n6), .ZN(
        sub_430_b0_n48) );
  AND2_X4 sub_430_b0_U47 ( .A1(sub_430_b0_n114), .A2(sub_430_b0_n5), .ZN(
        sub_430_b0_n47) );
  AND2_X4 sub_430_b0_U46 ( .A1(sub_430_b0_n112), .A2(sub_430_b0_n25), .ZN(
        sub_430_b0_n46) );
  AND2_X4 sub_430_b0_U45 ( .A1(sub_430_b0_n110), .A2(sub_430_b0_n21), .ZN(
        sub_430_b0_n45) );
  AND2_X4 sub_430_b0_U44 ( .A1(sub_430_b0_n108), .A2(sub_430_b0_n20), .ZN(
        sub_430_b0_n44) );
  AND2_X4 sub_430_b0_U43 ( .A1(sub_430_b0_n106), .A2(sub_430_b0_n19), .ZN(
        sub_430_b0_n43) );
  XOR2_X2 sub_430_b0_U42 ( .A(sub_430_b0_n149), .B(sub_430_b0_n65), .Z(N355)
         );
  XOR2_X2 sub_430_b0_U41 ( .A(sub_430_b0_n150), .B(sub_430_b0_n22), .Z(N354)
         );
  XOR2_X2 sub_430_b0_U40 ( .A(sub_430_b0_n151), .B(sub_430_b0_n66), .Z(N353)
         );
  XOR2_X2 sub_430_b0_U39 ( .A(sub_430_b0_n152), .B(sub_430_b0_n23), .Z(N352)
         );
  XOR2_X2 sub_430_b0_U38 ( .A(sub_430_b0_n153), .B(sub_430_b0_n67), .Z(N351)
         );
  XOR2_X2 sub_430_b0_U37 ( .A(sub_430_b0_n154), .B(sub_430_b0_n24), .Z(N350)
         );
  XOR2_X2 sub_430_b0_U36 ( .A(sub_430_b0_n155), .B(sub_430_b0_n68), .Z(N349)
         );
  XOR2_X2 sub_430_b0_U35 ( .A(sub_430_b0_n156), .B(sub_430_b0_n157), .Z(N348)
         );
  XOR2_X2 sub_430_b0_U34 ( .A(sub_430_b0_n109), .B(sub_430_b0_n45), .Z(N395)
         );
  XOR2_X2 sub_430_b0_U33 ( .A(sub_430_b0_n110), .B(sub_430_b0_n21), .Z(N394)
         );
  XOR2_X2 sub_430_b0_U32 ( .A(sub_430_b0_n111), .B(sub_430_b0_n46), .Z(N393)
         );
  XOR2_X2 sub_430_b0_U31 ( .A(sub_430_b0_n112), .B(sub_430_b0_n25), .Z(N392)
         );
  XOR2_X2 sub_430_b0_U30 ( .A(sub_430_b0_n113), .B(sub_430_b0_n47), .Z(N391)
         );
  XOR2_X2 sub_430_b0_U29 ( .A(sub_430_b0_n105), .B(sub_430_b0_n43), .Z(N399)
         );
  XOR2_X2 sub_430_b0_U28 ( .A(sub_430_b0_n106), .B(sub_430_b0_n19), .Z(N398)
         );
  XOR2_X2 sub_430_b0_U27 ( .A(sub_430_b0_n107), .B(sub_430_b0_n44), .Z(N397)
         );
  XOR2_X2 sub_430_b0_U26 ( .A(sub_430_b0_n108), .B(sub_430_b0_n20), .Z(N396)
         );
  AND2_X4 sub_430_b0_U25 ( .A1(sub_430_b0_n113), .A2(sub_430_b0_n47), .ZN(
        sub_430_b0_n25) );
  AND2_X4 sub_430_b0_U24 ( .A1(sub_430_b0_n155), .A2(sub_430_b0_n68), .ZN(
        sub_430_b0_n24) );
  AND2_X4 sub_430_b0_U23 ( .A1(sub_430_b0_n153), .A2(sub_430_b0_n67), .ZN(
        sub_430_b0_n23) );
  AND2_X4 sub_430_b0_U22 ( .A1(sub_430_b0_n151), .A2(sub_430_b0_n66), .ZN(
        sub_430_b0_n22) );
  AND2_X4 sub_430_b0_U21 ( .A1(sub_430_b0_n111), .A2(sub_430_b0_n46), .ZN(
        sub_430_b0_n21) );
  AND2_X4 sub_430_b0_U20 ( .A1(sub_430_b0_n109), .A2(sub_430_b0_n45), .ZN(
        sub_430_b0_n20) );
  AND2_X4 sub_430_b0_U19 ( .A1(sub_430_b0_n107), .A2(sub_430_b0_n44), .ZN(
        sub_430_b0_n19) );
  AND2_X4 sub_430_b0_U18 ( .A1(sub_430_b0_n141), .A2(sub_430_b0_n61), .ZN(
        sub_430_b0_n18) );
  AND2_X4 sub_430_b0_U17 ( .A1(sub_430_b0_n139), .A2(sub_430_b0_n60), .ZN(
        sub_430_b0_n17) );
  AND2_X4 sub_430_b0_U16 ( .A1(sub_430_b0_n137), .A2(sub_430_b0_n59), .ZN(
        sub_430_b0_n16) );
  AND2_X4 sub_430_b0_U15 ( .A1(sub_430_b0_n135), .A2(sub_430_b0_n58), .ZN(
        sub_430_b0_n15) );
  AND2_X4 sub_430_b0_U14 ( .A1(sub_430_b0_n133), .A2(sub_430_b0_n57), .ZN(
        sub_430_b0_n14) );
  AND2_X4 sub_430_b0_U13 ( .A1(sub_430_b0_n131), .A2(sub_430_b0_n56), .ZN(
        sub_430_b0_n13) );
  AND2_X4 sub_430_b0_U12 ( .A1(sub_430_b0_n129), .A2(sub_430_b0_n55), .ZN(
        sub_430_b0_n12) );
  AND2_X4 sub_430_b0_U11 ( .A1(sub_430_b0_n127), .A2(sub_430_b0_n54), .ZN(
        sub_430_b0_n11) );
  AND2_X4 sub_430_b0_U10 ( .A1(sub_430_b0_n125), .A2(sub_430_b0_n53), .ZN(
        sub_430_b0_n10) );
  AND2_X4 sub_430_b0_U9 ( .A1(sub_430_b0_n123), .A2(sub_430_b0_n52), .ZN(
        sub_430_b0_n9) );
  AND2_X4 sub_430_b0_U8 ( .A1(sub_430_b0_n121), .A2(sub_430_b0_n51), .ZN(
        sub_430_b0_n8) );
  AND2_X4 sub_430_b0_U7 ( .A1(sub_430_b0_n119), .A2(sub_430_b0_n50), .ZN(
        sub_430_b0_n7) );
  AND2_X4 sub_430_b0_U6 ( .A1(sub_430_b0_n117), .A2(sub_430_b0_n49), .ZN(
        sub_430_b0_n6) );
  AND2_X4 sub_430_b0_U5 ( .A1(sub_430_b0_n115), .A2(sub_430_b0_n48), .ZN(
        sub_430_b0_n5) );
  AND2_X4 sub_430_b0_U4 ( .A1(sub_430_b0_n149), .A2(sub_430_b0_n65), .ZN(
        sub_430_b0_n4) );
  AND2_X4 sub_430_b0_U3 ( .A1(sub_430_b0_n147), .A2(sub_430_b0_n64), .ZN(
        sub_430_b0_n3) );
  AND2_X4 sub_430_b0_U2 ( .A1(sub_430_b0_n145), .A2(sub_430_b0_n63), .ZN(
        sub_430_b0_n2) );
  AND2_X4 sub_430_b0_U1 ( .A1(sub_430_b0_n143), .A2(sub_430_b0_n62), .ZN(
        sub_430_b0_n1) );
  AND2_X1 sll_381_U55 ( .A1(fracta_mul[0]), .A2(sll_381_n2), .ZN(
        sll_381_ML_int_1__0_) );
  AND2_X1 sll_381_U54 ( .A1(sll_381_ML_int_1__0_), .A2(sll_381_n4), .ZN(
        sll_381_ML_int_2__0_) );
  AND2_X1 sll_381_U53 ( .A1(sll_381_ML_int_1__1_), .A2(sll_381_n4), .ZN(
        sll_381_ML_int_2__1_) );
  AND2_X1 sll_381_U52 ( .A1(sll_381_ML_int_2__0_), .A2(sll_381_n9), .ZN(
        sll_381_ML_int_3__0_) );
  AND2_X1 sll_381_U51 ( .A1(sll_381_ML_int_2__1_), .A2(sll_381_n9), .ZN(
        sll_381_ML_int_3__1_) );
  AND2_X1 sll_381_U50 ( .A1(sll_381_ML_int_2__2_), .A2(sll_381_n9), .ZN(
        sll_381_ML_int_3__2_) );
  AND2_X1 sll_381_U49 ( .A1(sll_381_ML_int_2__3_), .A2(sll_381_n9), .ZN(
        sll_381_ML_int_3__3_) );
  NAND2_X1 sll_381_U48 ( .A1(sll_381_ML_int_3__0_), .A2(sll_381_n11), .ZN(
        sll_381_n30) );
  NAND2_X1 sll_381_U47 ( .A1(sll_381_ML_int_3__1_), .A2(sll_381_n11), .ZN(
        sll_381_n29) );
  NAND2_X1 sll_381_U46 ( .A1(sll_381_ML_int_3__2_), .A2(sll_381_n11), .ZN(
        sll_381_n28) );
  NAND2_X1 sll_381_U45 ( .A1(sll_381_ML_int_3__3_), .A2(sll_381_n11), .ZN(
        sll_381_n27) );
  NAND2_X1 sll_381_U44 ( .A1(sll_381_ML_int_3__4_), .A2(sll_381_n11), .ZN(
        sll_381_n26) );
  NAND2_X1 sll_381_U43 ( .A1(sll_381_ML_int_3__5_), .A2(sll_381_n11), .ZN(
        sll_381_n25) );
  NAND2_X1 sll_381_U42 ( .A1(sll_381_ML_int_3__6_), .A2(sll_381_n11), .ZN(
        sll_381_n24) );
  NAND2_X1 sll_381_U41 ( .A1(sll_381_ML_int_3__7_), .A2(sll_381_n11), .ZN(
        sll_381_n23) );
  NOR2_X1 sll_381_U40 ( .A1(div_opa_ldz_d[4]), .A2(sll_381_n30), .ZN(N261) );
  AND2_X1 sll_381_U39 ( .A1(sll_381_ML_int_4__10_), .A2(sll_381_n13), .ZN(N271) );
  AND2_X1 sll_381_U38 ( .A1(sll_381_ML_int_4__11_), .A2(sll_381_n13), .ZN(N272) );
  AND2_X1 sll_381_U37 ( .A1(sll_381_ML_int_4__12_), .A2(sll_381_n13), .ZN(N273) );
  AND2_X1 sll_381_U36 ( .A1(sll_381_ML_int_4__13_), .A2(sll_381_n13), .ZN(N274) );
  AND2_X1 sll_381_U35 ( .A1(sll_381_ML_int_4__14_), .A2(sll_381_n13), .ZN(N275) );
  AND2_X1 sll_381_U34 ( .A1(sll_381_ML_int_4__15_), .A2(sll_381_n13), .ZN(N276) );
  NOR2_X1 sll_381_U33 ( .A1(sll_381_n14), .A2(sll_381_n29), .ZN(N262) );
  NOR2_X1 sll_381_U32 ( .A1(sll_381_n12), .A2(sll_381_n28), .ZN(N263) );
  NOR2_X1 sll_381_U31 ( .A1(sll_381_n12), .A2(sll_381_n27), .ZN(N264) );
  NOR2_X1 sll_381_U30 ( .A1(sll_381_n12), .A2(sll_381_n26), .ZN(N265) );
  NOR2_X1 sll_381_U29 ( .A1(div_opa_ldz_d[4]), .A2(sll_381_n25), .ZN(N266) );
  NOR2_X1 sll_381_U28 ( .A1(sll_381_n12), .A2(sll_381_n24), .ZN(N267) );
  NOR2_X1 sll_381_U27 ( .A1(sll_381_n12), .A2(sll_381_n23), .ZN(N268) );
  AND2_X1 sll_381_U26 ( .A1(sll_381_ML_int_4__8_), .A2(sll_381_n13), .ZN(N269)
         );
  AND2_X1 sll_381_U25 ( .A1(sll_381_ML_int_4__9_), .A2(sll_381_n13), .ZN(N270)
         );
  INV_X4 sll_381_U24 ( .A(sll_381_n23), .ZN(sll_381_n22) );
  INV_X4 sll_381_U23 ( .A(sll_381_n27), .ZN(sll_381_n21) );
  INV_X4 sll_381_U22 ( .A(sll_381_n24), .ZN(sll_381_n20) );
  INV_X4 sll_381_U21 ( .A(sll_381_n28), .ZN(sll_381_n19) );
  INV_X4 sll_381_U20 ( .A(sll_381_n26), .ZN(sll_381_n18) );
  INV_X4 sll_381_U19 ( .A(sll_381_n30), .ZN(sll_381_n17) );
  INV_X4 sll_381_U18 ( .A(sll_381_n25), .ZN(sll_381_n16) );
  INV_X4 sll_381_U17 ( .A(sll_381_n29), .ZN(sll_381_n15) );
  INV_X4 sll_381_U16 ( .A(sll_381_n11), .ZN(sll_381_n10) );
  INV_X4 sll_381_U15 ( .A(sll_381_n9), .ZN(sll_381_n8) );
  INV_X4 sll_381_U14 ( .A(sll_381_n4), .ZN(sll_381_n6) );
  INV_X4 sll_381_U13 ( .A(sll_381_n13), .ZN(sll_381_n14) );
  INV_X4 sll_381_U12 ( .A(sll_381_n13), .ZN(sll_381_n12) );
  INV_X4 sll_381_U11 ( .A(sll_381_n9), .ZN(sll_381_n7) );
  INV_X4 sll_381_U10 ( .A(div_opa_ldz_d[2]), .ZN(sll_381_n9) );
  INV_X4 sll_381_U9 ( .A(div_opa_ldz_d[3]), .ZN(sll_381_n11) );
  INV_X4 sll_381_U8 ( .A(div_opa_ldz_d[4]), .ZN(sll_381_n13) );
  INV_X4 sll_381_U7 ( .A(div_opa_ldz_d[0]), .ZN(sll_381_n2) );
  INV_X4 sll_381_U6 ( .A(sll_381_n2), .ZN(sll_381_n1) );
  INV_X4 sll_381_U5 ( .A(sll_381_n4), .ZN(sll_381_n5) );
  INV_X4 sll_381_U4 ( .A(sll_381_n2), .ZN(sll_381_n3) );
  INV_X4 sll_381_U3 ( .A(div_opa_ldz_d[1]), .ZN(sll_381_n4) );
  MUX2_X2 sll_381_M1_0_1 ( .A(fracta_mul[1]), .B(fracta_mul[0]), .S(sll_381_n3), .Z(sll_381_ML_int_1__1_) );
  MUX2_X2 sll_381_M1_0_2 ( .A(fracta_mul[2]), .B(fracta_mul[1]), .S(sll_381_n3), .Z(sll_381_ML_int_1__2_) );
  MUX2_X2 sll_381_M1_0_3 ( .A(fracta_mul[3]), .B(fracta_mul[2]), .S(sll_381_n3), .Z(sll_381_ML_int_1__3_) );
  MUX2_X2 sll_381_M1_0_4 ( .A(fracta_mul[4]), .B(fracta_mul[3]), .S(sll_381_n3), .Z(sll_381_ML_int_1__4_) );
  MUX2_X2 sll_381_M1_0_5 ( .A(fracta_mul[5]), .B(fracta_mul[4]), .S(sll_381_n3), .Z(sll_381_ML_int_1__5_) );
  MUX2_X2 sll_381_M1_0_6 ( .A(fracta_mul[6]), .B(fracta_mul[5]), .S(sll_381_n3), .Z(sll_381_ML_int_1__6_) );
  MUX2_X2 sll_381_M1_0_7 ( .A(fracta_mul[7]), .B(fracta_mul[6]), .S(sll_381_n3), .Z(sll_381_ML_int_1__7_) );
  MUX2_X2 sll_381_M1_0_8 ( .A(fracta_mul[8]), .B(fracta_mul[7]), .S(sll_381_n3), .Z(sll_381_ML_int_1__8_) );
  MUX2_X2 sll_381_M1_0_9 ( .A(fracta_mul[9]), .B(fracta_mul[8]), .S(sll_381_n3), .Z(sll_381_ML_int_1__9_) );
  MUX2_X2 sll_381_M1_0_10 ( .A(fracta_mul[10]), .B(fracta_mul[9]), .S(
        sll_381_n3), .Z(sll_381_ML_int_1__10_) );
  MUX2_X2 sll_381_M1_0_11 ( .A(fracta_mul[11]), .B(fracta_mul[10]), .S(
        sll_381_n3), .Z(sll_381_ML_int_1__11_) );
  MUX2_X2 sll_381_M1_0_12 ( .A(fracta_mul[12]), .B(fracta_mul[11]), .S(
        sll_381_n3), .Z(sll_381_ML_int_1__12_) );
  MUX2_X2 sll_381_M1_0_13 ( .A(fracta_mul[13]), .B(fracta_mul[12]), .S(
        sll_381_n3), .Z(sll_381_ML_int_1__13_) );
  MUX2_X2 sll_381_M1_0_14 ( .A(fracta_mul[14]), .B(fracta_mul[13]), .S(
        sll_381_n3), .Z(sll_381_ML_int_1__14_) );
  MUX2_X2 sll_381_M1_0_15 ( .A(fracta_mul[15]), .B(fracta_mul[14]), .S(
        sll_381_n3), .Z(sll_381_ML_int_1__15_) );
  MUX2_X2 sll_381_M1_0_16 ( .A(fracta_mul[16]), .B(fracta_mul[15]), .S(
        sll_381_n3), .Z(sll_381_ML_int_1__16_) );
  MUX2_X2 sll_381_M1_0_17 ( .A(fracta_mul[17]), .B(fracta_mul[16]), .S(
        sll_381_n3), .Z(sll_381_ML_int_1__17_) );
  MUX2_X2 sll_381_M1_0_18 ( .A(fracta_mul[18]), .B(fracta_mul[17]), .S(
        sll_381_n3), .Z(sll_381_ML_int_1__18_) );
  MUX2_X2 sll_381_M1_0_19 ( .A(fracta_mul[19]), .B(fracta_mul[18]), .S(
        sll_381_n3), .Z(sll_381_ML_int_1__19_) );
  MUX2_X2 sll_381_M1_0_20 ( .A(fracta_mul[20]), .B(fracta_mul[19]), .S(
        sll_381_n3), .Z(sll_381_ML_int_1__20_) );
  MUX2_X2 sll_381_M1_0_21 ( .A(fracta_mul[21]), .B(fracta_mul[20]), .S(
        sll_381_n3), .Z(sll_381_ML_int_1__21_) );
  MUX2_X2 sll_381_M1_0_22 ( .A(fracta_mul[22]), .B(fracta_mul[21]), .S(
        sll_381_n3), .Z(sll_381_ML_int_1__22_) );
  MUX2_X2 sll_381_M1_0_23 ( .A(fracta_mul[23]), .B(fracta_mul[22]), .S(
        sll_381_n1), .Z(sll_381_ML_int_1__23_) );
  MUX2_X2 sll_381_M1_0_24 ( .A(fracta_mul[24]), .B(fracta_mul[23]), .S(
        sll_381_n1), .Z(sll_381_ML_int_1__24_) );
  MUX2_X2 sll_381_M1_0_25 ( .A(fracta_mul[25]), .B(fracta_mul[24]), .S(
        div_opa_ldz_d[0]), .Z(sll_381_ML_int_1__25_) );
  MUX2_X2 sll_381_M1_0_26 ( .A(fracta_mul[26]), .B(fracta_mul[25]), .S(
        div_opa_ldz_d[0]), .Z(sll_381_ML_int_1__26_) );
  MUX2_X2 sll_381_M1_0_27 ( .A(fracta_mul[27]), .B(fracta_mul[26]), .S(
        div_opa_ldz_d[0]), .Z(sll_381_ML_int_1__27_) );
  MUX2_X2 sll_381_M1_0_28 ( .A(fracta_mul[28]), .B(fracta_mul[27]), .S(
        div_opa_ldz_d[0]), .Z(sll_381_ML_int_1__28_) );
  MUX2_X2 sll_381_M1_0_29 ( .A(fracta_mul[29]), .B(fracta_mul[28]), .S(
        div_opa_ldz_d[0]), .Z(sll_381_ML_int_1__29_) );
  MUX2_X2 sll_381_M1_0_30 ( .A(fracta_mul[30]), .B(fracta_mul[29]), .S(
        div_opa_ldz_d[0]), .Z(sll_381_ML_int_1__30_) );
  MUX2_X2 sll_381_M1_0_31 ( .A(fracta_mul[31]), .B(fracta_mul[30]), .S(
        div_opa_ldz_d[0]), .Z(sll_381_ML_int_1__31_) );
  MUX2_X2 sll_381_M1_0_32 ( .A(fracta_mul[32]), .B(fracta_mul[31]), .S(
        div_opa_ldz_d[0]), .Z(sll_381_ML_int_1__32_) );
  MUX2_X2 sll_381_M1_0_33 ( .A(fracta_mul[33]), .B(fracta_mul[32]), .S(
        div_opa_ldz_d[0]), .Z(sll_381_ML_int_1__33_) );
  MUX2_X2 sll_381_M1_0_34 ( .A(fracta_mul[34]), .B(fracta_mul[33]), .S(
        div_opa_ldz_d[0]), .Z(sll_381_ML_int_1__34_) );
  MUX2_X2 sll_381_M1_0_35 ( .A(fracta_mul[35]), .B(fracta_mul[34]), .S(
        div_opa_ldz_d[0]), .Z(sll_381_ML_int_1__35_) );
  MUX2_X2 sll_381_M1_0_36 ( .A(fracta_mul[36]), .B(fracta_mul[35]), .S(
        div_opa_ldz_d[0]), .Z(sll_381_ML_int_1__36_) );
  MUX2_X2 sll_381_M1_0_37 ( .A(fracta_mul[37]), .B(fracta_mul[36]), .S(
        div_opa_ldz_d[0]), .Z(sll_381_ML_int_1__37_) );
  MUX2_X2 sll_381_M1_0_38 ( .A(fracta_mul[38]), .B(fracta_mul[37]), .S(
        div_opa_ldz_d[0]), .Z(sll_381_ML_int_1__38_) );
  MUX2_X2 sll_381_M1_0_39 ( .A(fracta_mul[39]), .B(fracta_mul[38]), .S(
        div_opa_ldz_d[0]), .Z(sll_381_ML_int_1__39_) );
  MUX2_X2 sll_381_M1_0_40 ( .A(fracta_mul[40]), .B(fracta_mul[39]), .S(
        div_opa_ldz_d[0]), .Z(sll_381_ML_int_1__40_) );
  MUX2_X2 sll_381_M1_0_41 ( .A(fracta_mul[41]), .B(fracta_mul[40]), .S(
        div_opa_ldz_d[0]), .Z(sll_381_ML_int_1__41_) );
  MUX2_X2 sll_381_M1_0_42 ( .A(fracta_mul[42]), .B(fracta_mul[41]), .S(
        div_opa_ldz_d[0]), .Z(sll_381_ML_int_1__42_) );
  MUX2_X2 sll_381_M1_0_43 ( .A(fracta_mul[43]), .B(fracta_mul[42]), .S(
        div_opa_ldz_d[0]), .Z(sll_381_ML_int_1__43_) );
  MUX2_X2 sll_381_M1_0_44 ( .A(fracta_mul[44]), .B(fracta_mul[43]), .S(
        div_opa_ldz_d[0]), .Z(sll_381_ML_int_1__44_) );
  MUX2_X2 sll_381_M1_0_45 ( .A(fracta_mul[45]), .B(fracta_mul[44]), .S(
        div_opa_ldz_d[0]), .Z(sll_381_ML_int_1__45_) );
  MUX2_X2 sll_381_M1_0_46 ( .A(fracta_mul[46]), .B(fracta_mul[45]), .S(
        div_opa_ldz_d[0]), .Z(sll_381_ML_int_1__46_) );
  MUX2_X2 sll_381_M1_0_47 ( .A(fracta_mul[47]), .B(fracta_mul[46]), .S(
        div_opa_ldz_d[0]), .Z(sll_381_ML_int_1__47_) );
  MUX2_X2 sll_381_M1_0_48 ( .A(fracta_mul[48]), .B(fracta_mul[47]), .S(
        sll_381_n1), .Z(sll_381_ML_int_1__48_) );
  MUX2_X2 sll_381_M1_0_49 ( .A(fracta_mul[49]), .B(fracta_mul[48]), .S(
        sll_381_n1), .Z(sll_381_ML_int_1__49_) );
  MUX2_X2 sll_381_M1_0_50 ( .A(fracta_mul[50]), .B(fracta_mul[49]), .S(
        sll_381_n1), .Z(sll_381_ML_int_1__50_) );
  MUX2_X2 sll_381_M1_0_51 ( .A(fracta_mul[51]), .B(fracta_mul[50]), .S(
        sll_381_n1), .Z(sll_381_ML_int_1__51_) );
  MUX2_X2 sll_381_M1_0_52 ( .A(n4825), .B(fracta_mul[51]), .S(sll_381_n1), .Z(
        sll_381_ML_int_1__52_) );
  MUX2_X2 sll_381_M1_1_2 ( .A(sll_381_ML_int_1__2_), .B(sll_381_ML_int_1__0_), 
        .S(sll_381_n5), .Z(sll_381_ML_int_2__2_) );
  MUX2_X2 sll_381_M1_1_3 ( .A(sll_381_ML_int_1__3_), .B(sll_381_ML_int_1__1_), 
        .S(div_opa_ldz_d[1]), .Z(sll_381_ML_int_2__3_) );
  MUX2_X2 sll_381_M1_1_4 ( .A(sll_381_ML_int_1__4_), .B(sll_381_ML_int_1__2_), 
        .S(div_opa_ldz_d[1]), .Z(sll_381_ML_int_2__4_) );
  MUX2_X2 sll_381_M1_1_5 ( .A(sll_381_ML_int_1__5_), .B(sll_381_ML_int_1__3_), 
        .S(div_opa_ldz_d[1]), .Z(sll_381_ML_int_2__5_) );
  MUX2_X2 sll_381_M1_1_6 ( .A(sll_381_ML_int_1__6_), .B(sll_381_ML_int_1__4_), 
        .S(div_opa_ldz_d[1]), .Z(sll_381_ML_int_2__6_) );
  MUX2_X2 sll_381_M1_1_7 ( .A(sll_381_ML_int_1__7_), .B(sll_381_ML_int_1__5_), 
        .S(div_opa_ldz_d[1]), .Z(sll_381_ML_int_2__7_) );
  MUX2_X2 sll_381_M1_1_8 ( .A(sll_381_ML_int_1__8_), .B(sll_381_ML_int_1__6_), 
        .S(div_opa_ldz_d[1]), .Z(sll_381_ML_int_2__8_) );
  MUX2_X2 sll_381_M1_1_9 ( .A(sll_381_ML_int_1__9_), .B(sll_381_ML_int_1__7_), 
        .S(div_opa_ldz_d[1]), .Z(sll_381_ML_int_2__9_) );
  MUX2_X2 sll_381_M1_1_10 ( .A(sll_381_ML_int_1__10_), .B(sll_381_ML_int_1__8_), .S(div_opa_ldz_d[1]), .Z(sll_381_ML_int_2__10_) );
  MUX2_X2 sll_381_M1_1_11 ( .A(sll_381_ML_int_1__11_), .B(sll_381_ML_int_1__9_), .S(sll_381_n5), .Z(sll_381_ML_int_2__11_) );
  MUX2_X2 sll_381_M1_1_12 ( .A(sll_381_ML_int_1__12_), .B(
        sll_381_ML_int_1__10_), .S(div_opa_ldz_d[1]), .Z(sll_381_ML_int_2__12_) );
  MUX2_X2 sll_381_M1_1_13 ( .A(sll_381_ML_int_1__13_), .B(
        sll_381_ML_int_1__11_), .S(div_opa_ldz_d[1]), .Z(sll_381_ML_int_2__13_) );
  MUX2_X2 sll_381_M1_1_14 ( .A(sll_381_ML_int_1__14_), .B(
        sll_381_ML_int_1__12_), .S(div_opa_ldz_d[1]), .Z(sll_381_ML_int_2__14_) );
  MUX2_X2 sll_381_M1_1_15 ( .A(sll_381_ML_int_1__15_), .B(
        sll_381_ML_int_1__13_), .S(div_opa_ldz_d[1]), .Z(sll_381_ML_int_2__15_) );
  MUX2_X2 sll_381_M1_1_16 ( .A(sll_381_ML_int_1__16_), .B(
        sll_381_ML_int_1__14_), .S(sll_381_n5), .Z(sll_381_ML_int_2__16_) );
  MUX2_X2 sll_381_M1_1_17 ( .A(sll_381_ML_int_1__17_), .B(
        sll_381_ML_int_1__15_), .S(div_opa_ldz_d[1]), .Z(sll_381_ML_int_2__17_) );
  MUX2_X2 sll_381_M1_1_18 ( .A(sll_381_ML_int_1__18_), .B(
        sll_381_ML_int_1__16_), .S(div_opa_ldz_d[1]), .Z(sll_381_ML_int_2__18_) );
  MUX2_X2 sll_381_M1_1_19 ( .A(sll_381_ML_int_1__19_), .B(
        sll_381_ML_int_1__17_), .S(div_opa_ldz_d[1]), .Z(sll_381_ML_int_2__19_) );
  MUX2_X2 sll_381_M1_1_20 ( .A(sll_381_ML_int_1__20_), .B(
        sll_381_ML_int_1__18_), .S(div_opa_ldz_d[1]), .Z(sll_381_ML_int_2__20_) );
  MUX2_X2 sll_381_M1_1_21 ( .A(sll_381_ML_int_1__21_), .B(
        sll_381_ML_int_1__19_), .S(div_opa_ldz_d[1]), .Z(sll_381_ML_int_2__21_) );
  MUX2_X2 sll_381_M1_1_22 ( .A(sll_381_ML_int_1__22_), .B(
        sll_381_ML_int_1__20_), .S(div_opa_ldz_d[1]), .Z(sll_381_ML_int_2__22_) );
  MUX2_X2 sll_381_M1_1_23 ( .A(sll_381_ML_int_1__23_), .B(
        sll_381_ML_int_1__21_), .S(div_opa_ldz_d[1]), .Z(sll_381_ML_int_2__23_) );
  MUX2_X2 sll_381_M1_1_24 ( .A(sll_381_ML_int_1__24_), .B(
        sll_381_ML_int_1__22_), .S(sll_381_n5), .Z(sll_381_ML_int_2__24_) );
  MUX2_X2 sll_381_M1_1_25 ( .A(sll_381_ML_int_1__25_), .B(
        sll_381_ML_int_1__23_), .S(sll_381_n5), .Z(sll_381_ML_int_2__25_) );
  MUX2_X2 sll_381_M1_1_26 ( .A(sll_381_ML_int_1__26_), .B(
        sll_381_ML_int_1__24_), .S(sll_381_n5), .Z(sll_381_ML_int_2__26_) );
  MUX2_X2 sll_381_M1_1_27 ( .A(sll_381_ML_int_1__27_), .B(
        sll_381_ML_int_1__25_), .S(sll_381_n5), .Z(sll_381_ML_int_2__27_) );
  MUX2_X2 sll_381_M1_1_28 ( .A(sll_381_ML_int_1__28_), .B(
        sll_381_ML_int_1__26_), .S(sll_381_n5), .Z(sll_381_ML_int_2__28_) );
  MUX2_X2 sll_381_M1_1_29 ( .A(sll_381_ML_int_1__29_), .B(
        sll_381_ML_int_1__27_), .S(sll_381_n5), .Z(sll_381_ML_int_2__29_) );
  MUX2_X2 sll_381_M1_1_30 ( .A(sll_381_ML_int_1__30_), .B(
        sll_381_ML_int_1__28_), .S(sll_381_n5), .Z(sll_381_ML_int_2__30_) );
  MUX2_X2 sll_381_M1_1_31 ( .A(sll_381_ML_int_1__31_), .B(
        sll_381_ML_int_1__29_), .S(sll_381_n5), .Z(sll_381_ML_int_2__31_) );
  MUX2_X2 sll_381_M1_1_32 ( .A(sll_381_ML_int_1__32_), .B(
        sll_381_ML_int_1__30_), .S(sll_381_n5), .Z(sll_381_ML_int_2__32_) );
  MUX2_X2 sll_381_M1_1_33 ( .A(sll_381_ML_int_1__33_), .B(
        sll_381_ML_int_1__31_), .S(sll_381_n5), .Z(sll_381_ML_int_2__33_) );
  MUX2_X2 sll_381_M1_1_34 ( .A(sll_381_ML_int_1__34_), .B(
        sll_381_ML_int_1__32_), .S(sll_381_n5), .Z(sll_381_ML_int_2__34_) );
  MUX2_X2 sll_381_M1_1_35 ( .A(sll_381_ML_int_1__35_), .B(
        sll_381_ML_int_1__33_), .S(sll_381_n6), .Z(sll_381_ML_int_2__35_) );
  MUX2_X2 sll_381_M1_1_36 ( .A(sll_381_ML_int_1__36_), .B(
        sll_381_ML_int_1__34_), .S(sll_381_n6), .Z(sll_381_ML_int_2__36_) );
  MUX2_X2 sll_381_M1_1_37 ( .A(sll_381_ML_int_1__37_), .B(
        sll_381_ML_int_1__35_), .S(sll_381_n6), .Z(sll_381_ML_int_2__37_) );
  MUX2_X2 sll_381_M1_1_38 ( .A(sll_381_ML_int_1__38_), .B(
        sll_381_ML_int_1__36_), .S(sll_381_n6), .Z(sll_381_ML_int_2__38_) );
  MUX2_X2 sll_381_M1_1_39 ( .A(sll_381_ML_int_1__39_), .B(
        sll_381_ML_int_1__37_), .S(sll_381_n6), .Z(sll_381_ML_int_2__39_) );
  MUX2_X2 sll_381_M1_1_40 ( .A(sll_381_ML_int_1__40_), .B(
        sll_381_ML_int_1__38_), .S(sll_381_n6), .Z(sll_381_ML_int_2__40_) );
  MUX2_X2 sll_381_M1_1_41 ( .A(sll_381_ML_int_1__41_), .B(
        sll_381_ML_int_1__39_), .S(sll_381_n6), .Z(sll_381_ML_int_2__41_) );
  MUX2_X2 sll_381_M1_1_42 ( .A(sll_381_ML_int_1__42_), .B(
        sll_381_ML_int_1__40_), .S(sll_381_n6), .Z(sll_381_ML_int_2__42_) );
  MUX2_X2 sll_381_M1_1_43 ( .A(sll_381_ML_int_1__43_), .B(
        sll_381_ML_int_1__41_), .S(sll_381_n6), .Z(sll_381_ML_int_2__43_) );
  MUX2_X2 sll_381_M1_1_44 ( .A(sll_381_ML_int_1__44_), .B(
        sll_381_ML_int_1__42_), .S(sll_381_n6), .Z(sll_381_ML_int_2__44_) );
  MUX2_X2 sll_381_M1_1_45 ( .A(sll_381_ML_int_1__45_), .B(
        sll_381_ML_int_1__43_), .S(sll_381_n6), .Z(sll_381_ML_int_2__45_) );
  MUX2_X2 sll_381_M1_1_46 ( .A(sll_381_ML_int_1__46_), .B(
        sll_381_ML_int_1__44_), .S(sll_381_n6), .Z(sll_381_ML_int_2__46_) );
  MUX2_X2 sll_381_M1_1_47 ( .A(sll_381_ML_int_1__47_), .B(
        sll_381_ML_int_1__45_), .S(sll_381_n6), .Z(sll_381_ML_int_2__47_) );
  MUX2_X2 sll_381_M1_1_48 ( .A(sll_381_ML_int_1__48_), .B(
        sll_381_ML_int_1__46_), .S(sll_381_n6), .Z(sll_381_ML_int_2__48_) );
  MUX2_X2 sll_381_M1_1_49 ( .A(sll_381_ML_int_1__49_), .B(
        sll_381_ML_int_1__47_), .S(sll_381_n6), .Z(sll_381_ML_int_2__49_) );
  MUX2_X2 sll_381_M1_1_50 ( .A(sll_381_ML_int_1__50_), .B(
        sll_381_ML_int_1__48_), .S(sll_381_n6), .Z(sll_381_ML_int_2__50_) );
  MUX2_X2 sll_381_M1_1_51 ( .A(sll_381_ML_int_1__51_), .B(
        sll_381_ML_int_1__49_), .S(sll_381_n6), .Z(sll_381_ML_int_2__51_) );
  MUX2_X2 sll_381_M1_1_52 ( .A(sll_381_ML_int_1__52_), .B(
        sll_381_ML_int_1__50_), .S(sll_381_n6), .Z(sll_381_ML_int_2__52_) );
  MUX2_X2 sll_381_M1_2_4 ( .A(sll_381_ML_int_2__4_), .B(sll_381_ML_int_2__0_), 
        .S(sll_381_n7), .Z(sll_381_ML_int_3__4_) );
  MUX2_X2 sll_381_M1_2_5 ( .A(sll_381_ML_int_2__5_), .B(sll_381_ML_int_2__1_), 
        .S(sll_381_n7), .Z(sll_381_ML_int_3__5_) );
  MUX2_X2 sll_381_M1_2_6 ( .A(sll_381_ML_int_2__6_), .B(sll_381_ML_int_2__2_), 
        .S(sll_381_n7), .Z(sll_381_ML_int_3__6_) );
  MUX2_X2 sll_381_M1_2_7 ( .A(sll_381_ML_int_2__7_), .B(sll_381_ML_int_2__3_), 
        .S(sll_381_n7), .Z(sll_381_ML_int_3__7_) );
  MUX2_X2 sll_381_M1_2_8 ( .A(sll_381_ML_int_2__8_), .B(sll_381_ML_int_2__4_), 
        .S(sll_381_n7), .Z(sll_381_ML_int_3__8_) );
  MUX2_X2 sll_381_M1_2_9 ( .A(sll_381_ML_int_2__9_), .B(sll_381_ML_int_2__5_), 
        .S(sll_381_n7), .Z(sll_381_ML_int_3__9_) );
  MUX2_X2 sll_381_M1_2_10 ( .A(sll_381_ML_int_2__10_), .B(sll_381_ML_int_2__6_), .S(sll_381_n7), .Z(sll_381_ML_int_3__10_) );
  MUX2_X2 sll_381_M1_2_11 ( .A(sll_381_ML_int_2__11_), .B(sll_381_ML_int_2__7_), .S(sll_381_n7), .Z(sll_381_ML_int_3__11_) );
  MUX2_X2 sll_381_M1_2_12 ( .A(sll_381_ML_int_2__12_), .B(sll_381_ML_int_2__8_), .S(sll_381_n7), .Z(sll_381_ML_int_3__12_) );
  MUX2_X2 sll_381_M1_2_13 ( .A(sll_381_ML_int_2__13_), .B(sll_381_ML_int_2__9_), .S(sll_381_n7), .Z(sll_381_ML_int_3__13_) );
  MUX2_X2 sll_381_M1_2_14 ( .A(sll_381_ML_int_2__14_), .B(
        sll_381_ML_int_2__10_), .S(sll_381_n7), .Z(sll_381_ML_int_3__14_) );
  MUX2_X2 sll_381_M1_2_15 ( .A(sll_381_ML_int_2__15_), .B(
        sll_381_ML_int_2__11_), .S(sll_381_n8), .Z(sll_381_ML_int_3__15_) );
  MUX2_X2 sll_381_M1_2_16 ( .A(sll_381_ML_int_2__16_), .B(
        sll_381_ML_int_2__12_), .S(sll_381_n7), .Z(sll_381_ML_int_3__16_) );
  MUX2_X2 sll_381_M1_2_17 ( .A(sll_381_ML_int_2__17_), .B(
        sll_381_ML_int_2__13_), .S(sll_381_n7), .Z(sll_381_ML_int_3__17_) );
  MUX2_X2 sll_381_M1_2_18 ( .A(sll_381_ML_int_2__18_), .B(
        sll_381_ML_int_2__14_), .S(sll_381_n8), .Z(sll_381_ML_int_3__18_) );
  MUX2_X2 sll_381_M1_2_19 ( .A(sll_381_ML_int_2__19_), .B(
        sll_381_ML_int_2__15_), .S(sll_381_n7), .Z(sll_381_ML_int_3__19_) );
  MUX2_X2 sll_381_M1_2_20 ( .A(sll_381_ML_int_2__20_), .B(
        sll_381_ML_int_2__16_), .S(sll_381_n7), .Z(sll_381_ML_int_3__20_) );
  MUX2_X2 sll_381_M1_2_21 ( .A(sll_381_ML_int_2__21_), .B(
        sll_381_ML_int_2__17_), .S(sll_381_n8), .Z(sll_381_ML_int_3__21_) );
  MUX2_X2 sll_381_M1_2_22 ( .A(sll_381_ML_int_2__22_), .B(
        sll_381_ML_int_2__18_), .S(sll_381_n7), .Z(sll_381_ML_int_3__22_) );
  MUX2_X2 sll_381_M1_2_23 ( .A(sll_381_ML_int_2__23_), .B(
        sll_381_ML_int_2__19_), .S(sll_381_n7), .Z(sll_381_ML_int_3__23_) );
  MUX2_X2 sll_381_M1_2_24 ( .A(sll_381_ML_int_2__24_), .B(
        sll_381_ML_int_2__20_), .S(sll_381_n8), .Z(sll_381_ML_int_3__24_) );
  MUX2_X2 sll_381_M1_2_25 ( .A(sll_381_ML_int_2__25_), .B(
        sll_381_ML_int_2__21_), .S(sll_381_n7), .Z(sll_381_ML_int_3__25_) );
  MUX2_X2 sll_381_M1_2_26 ( .A(sll_381_ML_int_2__26_), .B(
        sll_381_ML_int_2__22_), .S(sll_381_n8), .Z(sll_381_ML_int_3__26_) );
  MUX2_X2 sll_381_M1_2_27 ( .A(sll_381_ML_int_2__27_), .B(
        sll_381_ML_int_2__23_), .S(sll_381_n8), .Z(sll_381_ML_int_3__27_) );
  MUX2_X2 sll_381_M1_2_28 ( .A(sll_381_ML_int_2__28_), .B(
        sll_381_ML_int_2__24_), .S(div_opa_ldz_d[2]), .Z(sll_381_ML_int_3__28_) );
  MUX2_X2 sll_381_M1_2_29 ( .A(sll_381_ML_int_2__29_), .B(
        sll_381_ML_int_2__25_), .S(div_opa_ldz_d[2]), .Z(sll_381_ML_int_3__29_) );
  MUX2_X2 sll_381_M1_2_30 ( .A(sll_381_ML_int_2__30_), .B(
        sll_381_ML_int_2__26_), .S(sll_381_n7), .Z(sll_381_ML_int_3__30_) );
  MUX2_X2 sll_381_M1_2_31 ( .A(sll_381_ML_int_2__31_), .B(
        sll_381_ML_int_2__27_), .S(div_opa_ldz_d[2]), .Z(sll_381_ML_int_3__31_) );
  MUX2_X2 sll_381_M1_2_32 ( .A(sll_381_ML_int_2__32_), .B(
        sll_381_ML_int_2__28_), .S(div_opa_ldz_d[2]), .Z(sll_381_ML_int_3__32_) );
  MUX2_X2 sll_381_M1_2_33 ( .A(sll_381_ML_int_2__33_), .B(
        sll_381_ML_int_2__29_), .S(div_opa_ldz_d[2]), .Z(sll_381_ML_int_3__33_) );
  MUX2_X2 sll_381_M1_2_34 ( .A(sll_381_ML_int_2__34_), .B(
        sll_381_ML_int_2__30_), .S(div_opa_ldz_d[2]), .Z(sll_381_ML_int_3__34_) );
  MUX2_X2 sll_381_M1_2_35 ( .A(sll_381_ML_int_2__35_), .B(
        sll_381_ML_int_2__31_), .S(div_opa_ldz_d[2]), .Z(sll_381_ML_int_3__35_) );
  MUX2_X2 sll_381_M1_2_36 ( .A(sll_381_ML_int_2__36_), .B(
        sll_381_ML_int_2__32_), .S(div_opa_ldz_d[2]), .Z(sll_381_ML_int_3__36_) );
  MUX2_X2 sll_381_M1_2_37 ( .A(sll_381_ML_int_2__37_), .B(
        sll_381_ML_int_2__33_), .S(sll_381_n8), .Z(sll_381_ML_int_3__37_) );
  MUX2_X2 sll_381_M1_2_38 ( .A(sll_381_ML_int_2__38_), .B(
        sll_381_ML_int_2__34_), .S(sll_381_n8), .Z(sll_381_ML_int_3__38_) );
  MUX2_X2 sll_381_M1_2_39 ( .A(sll_381_ML_int_2__39_), .B(
        sll_381_ML_int_2__35_), .S(sll_381_n8), .Z(sll_381_ML_int_3__39_) );
  MUX2_X2 sll_381_M1_2_40 ( .A(sll_381_ML_int_2__40_), .B(
        sll_381_ML_int_2__36_), .S(sll_381_n8), .Z(sll_381_ML_int_3__40_) );
  MUX2_X2 sll_381_M1_2_41 ( .A(sll_381_ML_int_2__41_), .B(
        sll_381_ML_int_2__37_), .S(sll_381_n8), .Z(sll_381_ML_int_3__41_) );
  MUX2_X2 sll_381_M1_2_42 ( .A(sll_381_ML_int_2__42_), .B(
        sll_381_ML_int_2__38_), .S(sll_381_n8), .Z(sll_381_ML_int_3__42_) );
  MUX2_X2 sll_381_M1_2_43 ( .A(sll_381_ML_int_2__43_), .B(
        sll_381_ML_int_2__39_), .S(sll_381_n8), .Z(sll_381_ML_int_3__43_) );
  MUX2_X2 sll_381_M1_2_44 ( .A(sll_381_ML_int_2__44_), .B(
        sll_381_ML_int_2__40_), .S(sll_381_n8), .Z(sll_381_ML_int_3__44_) );
  MUX2_X2 sll_381_M1_2_45 ( .A(sll_381_ML_int_2__45_), .B(
        sll_381_ML_int_2__41_), .S(sll_381_n8), .Z(sll_381_ML_int_3__45_) );
  MUX2_X2 sll_381_M1_2_46 ( .A(sll_381_ML_int_2__46_), .B(
        sll_381_ML_int_2__42_), .S(sll_381_n8), .Z(sll_381_ML_int_3__46_) );
  MUX2_X2 sll_381_M1_2_47 ( .A(sll_381_ML_int_2__47_), .B(
        sll_381_ML_int_2__43_), .S(sll_381_n8), .Z(sll_381_ML_int_3__47_) );
  MUX2_X2 sll_381_M1_2_48 ( .A(sll_381_ML_int_2__48_), .B(
        sll_381_ML_int_2__44_), .S(sll_381_n8), .Z(sll_381_ML_int_3__48_) );
  MUX2_X2 sll_381_M1_2_49 ( .A(sll_381_ML_int_2__49_), .B(
        sll_381_ML_int_2__45_), .S(sll_381_n8), .Z(sll_381_ML_int_3__49_) );
  MUX2_X2 sll_381_M1_2_50 ( .A(sll_381_ML_int_2__50_), .B(
        sll_381_ML_int_2__46_), .S(sll_381_n8), .Z(sll_381_ML_int_3__50_) );
  MUX2_X2 sll_381_M1_2_51 ( .A(sll_381_ML_int_2__51_), .B(
        sll_381_ML_int_2__47_), .S(sll_381_n8), .Z(sll_381_ML_int_3__51_) );
  MUX2_X2 sll_381_M1_2_52 ( .A(sll_381_ML_int_2__52_), .B(
        sll_381_ML_int_2__48_), .S(sll_381_n8), .Z(sll_381_ML_int_3__52_) );
  MUX2_X2 sll_381_M1_3_8 ( .A(sll_381_ML_int_3__8_), .B(sll_381_ML_int_3__0_), 
        .S(div_opa_ldz_d[3]), .Z(sll_381_ML_int_4__8_) );
  MUX2_X2 sll_381_M1_3_9 ( .A(sll_381_ML_int_3__9_), .B(sll_381_ML_int_3__1_), 
        .S(div_opa_ldz_d[3]), .Z(sll_381_ML_int_4__9_) );
  MUX2_X2 sll_381_M1_3_10 ( .A(sll_381_ML_int_3__10_), .B(sll_381_ML_int_3__2_), .S(div_opa_ldz_d[3]), .Z(sll_381_ML_int_4__10_) );
  MUX2_X2 sll_381_M1_3_11 ( .A(sll_381_ML_int_3__11_), .B(sll_381_ML_int_3__3_), .S(div_opa_ldz_d[3]), .Z(sll_381_ML_int_4__11_) );
  MUX2_X2 sll_381_M1_3_12 ( .A(sll_381_ML_int_3__12_), .B(sll_381_ML_int_3__4_), .S(div_opa_ldz_d[3]), .Z(sll_381_ML_int_4__12_) );
  MUX2_X2 sll_381_M1_3_13 ( .A(sll_381_ML_int_3__13_), .B(sll_381_ML_int_3__5_), .S(div_opa_ldz_d[3]), .Z(sll_381_ML_int_4__13_) );
  MUX2_X2 sll_381_M1_3_14 ( .A(sll_381_ML_int_3__14_), .B(sll_381_ML_int_3__6_), .S(div_opa_ldz_d[3]), .Z(sll_381_ML_int_4__14_) );
  MUX2_X2 sll_381_M1_3_15 ( .A(sll_381_ML_int_3__15_), .B(sll_381_ML_int_3__7_), .S(div_opa_ldz_d[3]), .Z(sll_381_ML_int_4__15_) );
  MUX2_X2 sll_381_M1_3_16 ( .A(sll_381_ML_int_3__16_), .B(sll_381_ML_int_3__8_), .S(div_opa_ldz_d[3]), .Z(sll_381_ML_int_4__16_) );
  MUX2_X2 sll_381_M1_3_17 ( .A(sll_381_ML_int_3__17_), .B(sll_381_ML_int_3__9_), .S(div_opa_ldz_d[3]), .Z(sll_381_ML_int_4__17_) );
  MUX2_X2 sll_381_M1_3_18 ( .A(sll_381_ML_int_3__18_), .B(
        sll_381_ML_int_3__10_), .S(div_opa_ldz_d[3]), .Z(sll_381_ML_int_4__18_) );
  MUX2_X2 sll_381_M1_3_19 ( .A(sll_381_ML_int_3__19_), .B(
        sll_381_ML_int_3__11_), .S(div_opa_ldz_d[3]), .Z(sll_381_ML_int_4__19_) );
  MUX2_X2 sll_381_M1_3_20 ( .A(sll_381_ML_int_3__20_), .B(
        sll_381_ML_int_3__12_), .S(div_opa_ldz_d[3]), .Z(sll_381_ML_int_4__20_) );
  MUX2_X2 sll_381_M1_3_21 ( .A(sll_381_ML_int_3__21_), .B(
        sll_381_ML_int_3__13_), .S(sll_381_n10), .Z(sll_381_ML_int_4__21_) );
  MUX2_X2 sll_381_M1_3_22 ( .A(sll_381_ML_int_3__22_), .B(
        sll_381_ML_int_3__14_), .S(div_opa_ldz_d[3]), .Z(sll_381_ML_int_4__22_) );
  MUX2_X2 sll_381_M1_3_23 ( .A(sll_381_ML_int_3__23_), .B(
        sll_381_ML_int_3__15_), .S(div_opa_ldz_d[3]), .Z(sll_381_ML_int_4__23_) );
  MUX2_X2 sll_381_M1_3_24 ( .A(sll_381_ML_int_3__24_), .B(
        sll_381_ML_int_3__16_), .S(div_opa_ldz_d[3]), .Z(sll_381_ML_int_4__24_) );
  MUX2_X2 sll_381_M1_3_25 ( .A(sll_381_ML_int_3__25_), .B(
        sll_381_ML_int_3__17_), .S(div_opa_ldz_d[3]), .Z(sll_381_ML_int_4__25_) );
  MUX2_X2 sll_381_M1_3_26 ( .A(sll_381_ML_int_3__26_), .B(
        sll_381_ML_int_3__18_), .S(div_opa_ldz_d[3]), .Z(sll_381_ML_int_4__26_) );
  MUX2_X2 sll_381_M1_3_27 ( .A(sll_381_ML_int_3__27_), .B(
        sll_381_ML_int_3__19_), .S(div_opa_ldz_d[3]), .Z(sll_381_ML_int_4__27_) );
  MUX2_X2 sll_381_M1_3_28 ( .A(sll_381_ML_int_3__28_), .B(
        sll_381_ML_int_3__20_), .S(div_opa_ldz_d[3]), .Z(sll_381_ML_int_4__28_) );
  MUX2_X2 sll_381_M1_3_29 ( .A(sll_381_ML_int_3__29_), .B(
        sll_381_ML_int_3__21_), .S(div_opa_ldz_d[3]), .Z(sll_381_ML_int_4__29_) );
  MUX2_X2 sll_381_M1_3_30 ( .A(sll_381_ML_int_3__30_), .B(
        sll_381_ML_int_3__22_), .S(sll_381_n10), .Z(sll_381_ML_int_4__30_) );
  MUX2_X2 sll_381_M1_3_31 ( .A(sll_381_ML_int_3__31_), .B(
        sll_381_ML_int_3__23_), .S(sll_381_n10), .Z(sll_381_ML_int_4__31_) );
  MUX2_X2 sll_381_M1_3_32 ( .A(sll_381_ML_int_3__32_), .B(
        sll_381_ML_int_3__24_), .S(sll_381_n10), .Z(sll_381_ML_int_4__32_) );
  MUX2_X2 sll_381_M1_3_33 ( .A(sll_381_ML_int_3__33_), .B(
        sll_381_ML_int_3__25_), .S(sll_381_n10), .Z(sll_381_ML_int_4__33_) );
  MUX2_X2 sll_381_M1_3_34 ( .A(sll_381_ML_int_3__34_), .B(
        sll_381_ML_int_3__26_), .S(sll_381_n10), .Z(sll_381_ML_int_4__34_) );
  MUX2_X2 sll_381_M1_3_35 ( .A(sll_381_ML_int_3__35_), .B(
        sll_381_ML_int_3__27_), .S(sll_381_n10), .Z(sll_381_ML_int_4__35_) );
  MUX2_X2 sll_381_M1_3_36 ( .A(sll_381_ML_int_3__36_), .B(
        sll_381_ML_int_3__28_), .S(sll_381_n10), .Z(sll_381_ML_int_4__36_) );
  MUX2_X2 sll_381_M1_3_37 ( .A(sll_381_ML_int_3__37_), .B(
        sll_381_ML_int_3__29_), .S(sll_381_n10), .Z(sll_381_ML_int_4__37_) );
  MUX2_X2 sll_381_M1_3_38 ( .A(sll_381_ML_int_3__38_), .B(
        sll_381_ML_int_3__30_), .S(sll_381_n10), .Z(sll_381_ML_int_4__38_) );
  MUX2_X2 sll_381_M1_3_39 ( .A(sll_381_ML_int_3__39_), .B(
        sll_381_ML_int_3__31_), .S(sll_381_n10), .Z(sll_381_ML_int_4__39_) );
  MUX2_X2 sll_381_M1_3_40 ( .A(sll_381_ML_int_3__40_), .B(
        sll_381_ML_int_3__32_), .S(sll_381_n10), .Z(sll_381_ML_int_4__40_) );
  MUX2_X2 sll_381_M1_3_41 ( .A(sll_381_ML_int_3__41_), .B(
        sll_381_ML_int_3__33_), .S(sll_381_n10), .Z(sll_381_ML_int_4__41_) );
  MUX2_X2 sll_381_M1_3_42 ( .A(sll_381_ML_int_3__42_), .B(
        sll_381_ML_int_3__34_), .S(sll_381_n10), .Z(sll_381_ML_int_4__42_) );
  MUX2_X2 sll_381_M1_3_43 ( .A(sll_381_ML_int_3__43_), .B(
        sll_381_ML_int_3__35_), .S(sll_381_n10), .Z(sll_381_ML_int_4__43_) );
  MUX2_X2 sll_381_M1_3_44 ( .A(sll_381_ML_int_3__44_), .B(
        sll_381_ML_int_3__36_), .S(sll_381_n10), .Z(sll_381_ML_int_4__44_) );
  MUX2_X2 sll_381_M1_3_45 ( .A(sll_381_ML_int_3__45_), .B(
        sll_381_ML_int_3__37_), .S(sll_381_n10), .Z(sll_381_ML_int_4__45_) );
  MUX2_X2 sll_381_M1_3_46 ( .A(sll_381_ML_int_3__46_), .B(
        sll_381_ML_int_3__38_), .S(sll_381_n10), .Z(sll_381_ML_int_4__46_) );
  MUX2_X2 sll_381_M1_3_47 ( .A(sll_381_ML_int_3__47_), .B(
        sll_381_ML_int_3__39_), .S(sll_381_n10), .Z(sll_381_ML_int_4__47_) );
  MUX2_X2 sll_381_M1_3_48 ( .A(sll_381_ML_int_3__48_), .B(
        sll_381_ML_int_3__40_), .S(sll_381_n10), .Z(sll_381_ML_int_4__48_) );
  MUX2_X2 sll_381_M1_3_49 ( .A(sll_381_ML_int_3__49_), .B(
        sll_381_ML_int_3__41_), .S(sll_381_n10), .Z(sll_381_ML_int_4__49_) );
  MUX2_X2 sll_381_M1_3_50 ( .A(sll_381_ML_int_3__50_), .B(
        sll_381_ML_int_3__42_), .S(sll_381_n10), .Z(sll_381_ML_int_4__50_) );
  MUX2_X2 sll_381_M1_3_51 ( .A(sll_381_ML_int_3__51_), .B(
        sll_381_ML_int_3__43_), .S(sll_381_n10), .Z(sll_381_ML_int_4__51_) );
  MUX2_X2 sll_381_M1_3_52 ( .A(sll_381_ML_int_3__52_), .B(
        sll_381_ML_int_3__44_), .S(sll_381_n10), .Z(sll_381_ML_int_4__52_) );
  MUX2_X2 sll_381_M1_4_16 ( .A(sll_381_ML_int_4__16_), .B(sll_381_n17), .S(
        sll_381_n12), .Z(N277) );
  MUX2_X2 sll_381_M1_4_17 ( .A(sll_381_ML_int_4__17_), .B(sll_381_n15), .S(
        sll_381_n12), .Z(N278) );
  MUX2_X2 sll_381_M1_4_18 ( .A(sll_381_ML_int_4__18_), .B(sll_381_n19), .S(
        sll_381_n14), .Z(N279) );
  MUX2_X2 sll_381_M1_4_19 ( .A(sll_381_ML_int_4__19_), .B(sll_381_n21), .S(
        sll_381_n12), .Z(N280) );
  MUX2_X2 sll_381_M1_4_20 ( .A(sll_381_ML_int_4__20_), .B(sll_381_n18), .S(
        sll_381_n12), .Z(N281) );
  MUX2_X2 sll_381_M1_4_21 ( .A(sll_381_ML_int_4__21_), .B(sll_381_n16), .S(
        sll_381_n14), .Z(N282) );
  MUX2_X2 sll_381_M1_4_22 ( .A(sll_381_ML_int_4__22_), .B(sll_381_n20), .S(
        sll_381_n12), .Z(N283) );
  MUX2_X2 sll_381_M1_4_23 ( .A(sll_381_ML_int_4__23_), .B(sll_381_n22), .S(
        div_opa_ldz_d[4]), .Z(N284) );
  MUX2_X2 sll_381_M1_4_24 ( .A(sll_381_ML_int_4__24_), .B(sll_381_ML_int_4__8_), .S(sll_381_n12), .Z(N285) );
  MUX2_X2 sll_381_M1_4_25 ( .A(sll_381_ML_int_4__25_), .B(sll_381_ML_int_4__9_), .S(div_opa_ldz_d[4]), .Z(N286) );
  MUX2_X2 sll_381_M1_4_26 ( .A(sll_381_ML_int_4__26_), .B(
        sll_381_ML_int_4__10_), .S(sll_381_n12), .Z(N287) );
  MUX2_X2 sll_381_M1_4_27 ( .A(sll_381_ML_int_4__27_), .B(
        sll_381_ML_int_4__11_), .S(div_opa_ldz_d[4]), .Z(N288) );
  MUX2_X2 sll_381_M1_4_28 ( .A(sll_381_ML_int_4__28_), .B(
        sll_381_ML_int_4__12_), .S(sll_381_n12), .Z(N289) );
  MUX2_X2 sll_381_M1_4_29 ( .A(sll_381_ML_int_4__29_), .B(
        sll_381_ML_int_4__13_), .S(div_opa_ldz_d[4]), .Z(N290) );
  MUX2_X2 sll_381_M1_4_30 ( .A(sll_381_ML_int_4__30_), .B(
        sll_381_ML_int_4__14_), .S(sll_381_n12), .Z(N291) );
  MUX2_X2 sll_381_M1_4_31 ( .A(sll_381_ML_int_4__31_), .B(
        sll_381_ML_int_4__15_), .S(sll_381_n14), .Z(N292) );
  MUX2_X2 sll_381_M1_4_32 ( .A(sll_381_ML_int_4__32_), .B(
        sll_381_ML_int_4__16_), .S(sll_381_n14), .Z(N293) );
  MUX2_X2 sll_381_M1_4_33 ( .A(sll_381_ML_int_4__33_), .B(
        sll_381_ML_int_4__17_), .S(sll_381_n14), .Z(N294) );
  MUX2_X2 sll_381_M1_4_34 ( .A(sll_381_ML_int_4__34_), .B(
        sll_381_ML_int_4__18_), .S(sll_381_n14), .Z(N295) );
  MUX2_X2 sll_381_M1_4_35 ( .A(sll_381_ML_int_4__35_), .B(
        sll_381_ML_int_4__19_), .S(sll_381_n14), .Z(N296) );
  MUX2_X2 sll_381_M1_4_36 ( .A(sll_381_ML_int_4__36_), .B(
        sll_381_ML_int_4__20_), .S(sll_381_n14), .Z(N297) );
  MUX2_X2 sll_381_M1_4_37 ( .A(sll_381_ML_int_4__37_), .B(
        sll_381_ML_int_4__21_), .S(sll_381_n14), .Z(N298) );
  MUX2_X2 sll_381_M1_4_38 ( .A(sll_381_ML_int_4__38_), .B(
        sll_381_ML_int_4__22_), .S(sll_381_n14), .Z(N299) );
  MUX2_X2 sll_381_M1_4_39 ( .A(sll_381_ML_int_4__39_), .B(
        sll_381_ML_int_4__23_), .S(sll_381_n14), .Z(N300) );
  MUX2_X2 sll_381_M1_4_40 ( .A(sll_381_ML_int_4__40_), .B(
        sll_381_ML_int_4__24_), .S(sll_381_n14), .Z(N301) );
  MUX2_X2 sll_381_M1_4_41 ( .A(sll_381_ML_int_4__41_), .B(
        sll_381_ML_int_4__25_), .S(sll_381_n14), .Z(N302) );
  MUX2_X2 sll_381_M1_4_42 ( .A(sll_381_ML_int_4__42_), .B(
        sll_381_ML_int_4__26_), .S(div_opa_ldz_d[4]), .Z(N303) );
  MUX2_X2 sll_381_M1_4_43 ( .A(sll_381_ML_int_4__43_), .B(
        sll_381_ML_int_4__27_), .S(sll_381_n12), .Z(N304) );
  MUX2_X2 sll_381_M1_4_44 ( .A(sll_381_ML_int_4__44_), .B(
        sll_381_ML_int_4__28_), .S(div_opa_ldz_d[4]), .Z(N305) );
  MUX2_X2 sll_381_M1_4_45 ( .A(sll_381_ML_int_4__45_), .B(
        sll_381_ML_int_4__29_), .S(div_opa_ldz_d[4]), .Z(N306) );
  MUX2_X2 sll_381_M1_4_46 ( .A(sll_381_ML_int_4__46_), .B(
        sll_381_ML_int_4__30_), .S(sll_381_n12), .Z(N307) );
  MUX2_X2 sll_381_M1_4_47 ( .A(sll_381_ML_int_4__47_), .B(
        sll_381_ML_int_4__31_), .S(div_opa_ldz_d[4]), .Z(N308) );
  MUX2_X2 sll_381_M1_4_48 ( .A(sll_381_ML_int_4__48_), .B(
        sll_381_ML_int_4__32_), .S(div_opa_ldz_d[4]), .Z(N309) );
  MUX2_X2 sll_381_M1_4_49 ( .A(sll_381_ML_int_4__49_), .B(
        sll_381_ML_int_4__33_), .S(div_opa_ldz_d[4]), .Z(N310) );
  MUX2_X2 sll_381_M1_4_50 ( .A(sll_381_ML_int_4__50_), .B(
        sll_381_ML_int_4__34_), .S(div_opa_ldz_d[4]), .Z(N311) );
  MUX2_X2 sll_381_M1_4_51 ( .A(sll_381_ML_int_4__51_), .B(
        sll_381_ML_int_4__35_), .S(div_opa_ldz_d[4]), .Z(N312) );
  MUX2_X2 sll_381_M1_4_52 ( .A(sll_381_ML_int_4__52_), .B(
        sll_381_ML_int_4__36_), .S(div_opa_ldz_d[4]), .Z(N313) );
  NAND2_X1 r466_U180 ( .A1(fracta_mul[49]), .A2(r466_n7), .ZN(r466_n168) );
  OR2_X1 r466_U179 ( .A1(r466_n1), .A2(u6_N50), .ZN(r466_n167) );
  AND2_X1 r466_U178 ( .A1(fracta_mul[0]), .A2(r466_n56), .ZN(r466_n178) );
  OAI22_X1 r466_U177 ( .A1(fracta_mul[1]), .A2(r466_n178), .B1(r466_n178), 
        .B2(r466_n55), .ZN(r466_n177) );
  AND3_X1 r466_U176 ( .A1(r466_n168), .A2(r466_n167), .A3(r466_n177), .ZN(
        r466_n176) );
  NAND2_X1 r466_U175 ( .A1(fracta_mul[48]), .A2(r466_n8), .ZN(r466_n93) );
  NAND2_X1 r466_U174 ( .A1(fracta_mul[46]), .A2(r466_n10), .ZN(r466_n97) );
  NAND2_X1 r466_U173 ( .A1(fracta_mul[47]), .A2(r466_n9), .ZN(r466_n94) );
  AND4_X1 r466_U172 ( .A1(r466_n176), .A2(r466_n93), .A3(r466_n97), .A4(
        r466_n94), .ZN(r466_n169) );
  NAND2_X1 r466_U171 ( .A1(fracta_mul[42]), .A2(r466_n14), .ZN(r466_n105) );
  NAND2_X1 r466_U170 ( .A1(fracta_mul[41]), .A2(r466_n15), .ZN(r466_n106) );
  NAND2_X1 r466_U169 ( .A1(fracta_mul[40]), .A2(r466_n16), .ZN(r466_n109) );
  NAND2_X1 r466_U168 ( .A1(fracta_mul[39]), .A2(r466_n17), .ZN(r466_n110) );
  AND4_X1 r466_U167 ( .A1(r466_n105), .A2(r466_n106), .A3(r466_n109), .A4(
        r466_n110), .ZN(r466_n175) );
  NAND2_X1 r466_U166 ( .A1(fracta_mul[45]), .A2(r466_n11), .ZN(r466_n98) );
  NAND2_X1 r466_U165 ( .A1(fracta_mul[43]), .A2(r466_n13), .ZN(r466_n102) );
  NAND2_X1 r466_U164 ( .A1(fracta_mul[44]), .A2(r466_n12), .ZN(r466_n101) );
  AND4_X1 r466_U163 ( .A1(r466_n175), .A2(r466_n98), .A3(r466_n102), .A4(
        r466_n101), .ZN(r466_n170) );
  NAND2_X1 r466_U162 ( .A1(fracta_mul[34]), .A2(r466_n22), .ZN(r466_n121) );
  NAND2_X1 r466_U161 ( .A1(fracta_mul[33]), .A2(r466_n23), .ZN(r466_n122) );
  NAND2_X1 r466_U160 ( .A1(fracta_mul[35]), .A2(r466_n21), .ZN(r466_n118) );
  AND3_X1 r466_U159 ( .A1(r466_n121), .A2(r466_n122), .A3(r466_n118), .ZN(
        r466_n174) );
  NAND2_X1 r466_U158 ( .A1(fracta_mul[38]), .A2(r466_n18), .ZN(r466_n113) );
  NAND2_X1 r466_U157 ( .A1(fracta_mul[36]), .A2(r466_n20), .ZN(r466_n117) );
  NAND2_X1 r466_U156 ( .A1(fracta_mul[37]), .A2(r466_n19), .ZN(r466_n114) );
  AND4_X1 r466_U155 ( .A1(r466_n174), .A2(r466_n113), .A3(r466_n117), .A4(
        r466_n114), .ZN(r466_n171) );
  NAND2_X1 r466_U154 ( .A1(fracta_mul[29]), .A2(r466_n27), .ZN(r466_n130) );
  NAND2_X1 r466_U153 ( .A1(fracta_mul[28]), .A2(r466_n28), .ZN(r466_n133) );
  NAND2_X1 r466_U152 ( .A1(fracta_mul[27]), .A2(r466_n29), .ZN(r466_n134) );
  NAND2_X1 r466_U151 ( .A1(fracta_mul[26]), .A2(r466_n30), .ZN(r466_n137) );
  AND4_X1 r466_U150 ( .A1(r466_n130), .A2(r466_n133), .A3(r466_n134), .A4(
        r466_n137), .ZN(r466_n173) );
  NAND2_X1 r466_U149 ( .A1(fracta_mul[32]), .A2(r466_n24), .ZN(r466_n125) );
  NAND2_X1 r466_U148 ( .A1(fracta_mul[30]), .A2(r466_n26), .ZN(r466_n129) );
  NAND2_X1 r466_U147 ( .A1(fracta_mul[31]), .A2(r466_n25), .ZN(r466_n126) );
  AND4_X1 r466_U146 ( .A1(r466_n173), .A2(r466_n125), .A3(r466_n129), .A4(
        r466_n126), .ZN(r466_n172) );
  NAND4_X1 r466_U145 ( .A1(r466_n169), .A2(r466_n170), .A3(r466_n171), .A4(
        r466_n172), .ZN(r466_n57) );
  NAND2_X1 r466_U144 ( .A1(fracta_mul[6]), .A2(r466_n50), .ZN(r466_n158) );
  NAND2_X1 r466_U143 ( .A1(fracta_mul[4]), .A2(r466_n52), .ZN(r466_n162) );
  NAND2_X1 r466_U142 ( .A1(fracta_mul[5]), .A2(r466_n51), .ZN(r466_n159) );
  AND3_X1 r466_U141 ( .A1(r466_n158), .A2(r466_n162), .A3(r466_n159), .ZN(
        r466_n76) );
  AND2_X1 r466_U140 ( .A1(fracta_mul[51]), .A2(r466_n6), .ZN(r466_n86) );
  AND2_X1 r466_U139 ( .A1(r466_n167), .A2(r466_n168), .ZN(r466_n90) );
  NAND2_X1 r466_U138 ( .A1(fracta_mul[25]), .A2(r466_n31), .ZN(r466_n63) );
  NAND2_X1 r466_U137 ( .A1(fracta_mul[24]), .A2(r466_n32), .ZN(r466_n61) );
  NAND2_X1 r466_U136 ( .A1(fracta_mul[23]), .A2(r466_n33), .ZN(r466_n62) );
  NAND2_X1 r466_U135 ( .A1(fracta_mul[22]), .A2(r466_n34), .ZN(r466_n65) );
  NAND2_X1 r466_U134 ( .A1(fracta_mul[21]), .A2(r466_n35), .ZN(r466_n67) );
  NAND2_X1 r466_U133 ( .A1(fracta_mul[20]), .A2(r466_n36), .ZN(r466_n66) );
  NAND2_X1 r466_U132 ( .A1(fracta_mul[19]), .A2(r466_n37), .ZN(r466_n70) );
  NAND2_X1 r466_U131 ( .A1(fracta_mul[18]), .A2(r466_n38), .ZN(r466_n68) );
  NAND2_X1 r466_U130 ( .A1(fracta_mul[17]), .A2(r466_n39), .ZN(r466_n69) );
  NAND2_X1 r466_U129 ( .A1(fracta_mul[16]), .A2(r466_n40), .ZN(r466_n75) );
  NAND2_X1 r466_U128 ( .A1(fracta_mul[15]), .A2(r466_n41), .ZN(r466_n74) );
  NAND2_X1 r466_U127 ( .A1(fracta_mul[14]), .A2(r466_n42), .ZN(r466_n73) );
  NAND2_X1 r466_U126 ( .A1(fracta_mul[13]), .A2(r466_n43), .ZN(r466_n72) );
  NAND2_X1 r466_U125 ( .A1(fracta_mul[12]), .A2(r466_n44), .ZN(r466_n80) );
  NAND2_X1 r466_U124 ( .A1(fracta_mul[11]), .A2(r466_n45), .ZN(r466_n82) );
  NAND2_X1 r466_U123 ( .A1(fracta_mul[10]), .A2(r466_n46), .ZN(r466_n81) );
  NAND2_X1 r466_U122 ( .A1(fracta_mul[9]), .A2(r466_n47), .ZN(r466_n85) );
  NAND2_X1 r466_U121 ( .A1(fracta_mul[8]), .A2(r466_n48), .ZN(r466_n83) );
  NAND2_X1 r466_U120 ( .A1(fracta_mul[7]), .A2(r466_n49), .ZN(r466_n84) );
  NAND2_X1 r466_U119 ( .A1(fracta_mul[3]), .A2(r466_n53), .ZN(r466_n87) );
  NOR2_X1 r466_U118 ( .A1(r466_n56), .A2(fracta_mul[0]), .ZN(r466_n165) );
  OAI21_X1 r466_U117 ( .B1(fracta_mul[1]), .B2(r466_n5), .A(r466_n55), .ZN(
        r466_n166) );
  NAND2_X1 r466_U116 ( .A1(fracta_mul[2]), .A2(r466_n54), .ZN(r466_n88) );
  OAI211_X1 r466_U115 ( .C1(r466_n165), .C2(r466_n4), .A(r466_n166), .B(
        r466_n88), .ZN(r466_n164) );
  OAI221_X1 r466_U114 ( .B1(fracta_mul[2]), .B2(r466_n54), .C1(fracta_mul[3]), 
        .C2(r466_n53), .A(r466_n164), .ZN(r466_n163) );
  NAND3_X1 r466_U113 ( .A1(r466_n162), .A2(r466_n87), .A3(r466_n163), .ZN(
        r466_n161) );
  OAI221_X1 r466_U112 ( .B1(fracta_mul[4]), .B2(r466_n52), .C1(fracta_mul[5]), 
        .C2(r466_n51), .A(r466_n161), .ZN(r466_n160) );
  NAND3_X1 r466_U111 ( .A1(r466_n158), .A2(r466_n159), .A3(r466_n160), .ZN(
        r466_n157) );
  OAI221_X1 r466_U110 ( .B1(fracta_mul[6]), .B2(r466_n50), .C1(fracta_mul[7]), 
        .C2(r466_n49), .A(r466_n157), .ZN(r466_n156) );
  NAND3_X1 r466_U109 ( .A1(r466_n83), .A2(r466_n84), .A3(r466_n156), .ZN(
        r466_n155) );
  OAI221_X1 r466_U108 ( .B1(fracta_mul[8]), .B2(r466_n48), .C1(fracta_mul[9]), 
        .C2(r466_n47), .A(r466_n155), .ZN(r466_n154) );
  NAND3_X1 r466_U107 ( .A1(r466_n81), .A2(r466_n85), .A3(r466_n154), .ZN(
        r466_n153) );
  OAI221_X1 r466_U106 ( .B1(fracta_mul[10]), .B2(r466_n46), .C1(fracta_mul[11]), .C2(r466_n45), .A(r466_n153), .ZN(r466_n152) );
  NAND3_X1 r466_U105 ( .A1(r466_n80), .A2(r466_n82), .A3(r466_n152), .ZN(
        r466_n151) );
  OAI221_X1 r466_U104 ( .B1(fracta_mul[12]), .B2(r466_n44), .C1(fracta_mul[13]), .C2(r466_n43), .A(r466_n151), .ZN(r466_n150) );
  NAND3_X1 r466_U103 ( .A1(r466_n73), .A2(r466_n72), .A3(r466_n150), .ZN(
        r466_n149) );
  OAI221_X1 r466_U102 ( .B1(fracta_mul[14]), .B2(r466_n42), .C1(fracta_mul[15]), .C2(r466_n41), .A(r466_n149), .ZN(r466_n148) );
  NAND3_X1 r466_U101 ( .A1(r466_n75), .A2(r466_n74), .A3(r466_n148), .ZN(
        r466_n147) );
  OAI221_X1 r466_U100 ( .B1(fracta_mul[16]), .B2(r466_n40), .C1(fracta_mul[17]), .C2(r466_n39), .A(r466_n147), .ZN(r466_n146) );
  NAND3_X1 r466_U99 ( .A1(r466_n68), .A2(r466_n69), .A3(r466_n146), .ZN(
        r466_n145) );
  OAI221_X1 r466_U98 ( .B1(fracta_mul[18]), .B2(r466_n38), .C1(fracta_mul[19]), 
        .C2(r466_n37), .A(r466_n145), .ZN(r466_n144) );
  NAND3_X1 r466_U97 ( .A1(r466_n66), .A2(r466_n70), .A3(r466_n144), .ZN(
        r466_n143) );
  OAI221_X1 r466_U96 ( .B1(fracta_mul[20]), .B2(r466_n36), .C1(fracta_mul[21]), 
        .C2(r466_n35), .A(r466_n143), .ZN(r466_n142) );
  NAND3_X1 r466_U95 ( .A1(r466_n65), .A2(r466_n67), .A3(r466_n142), .ZN(
        r466_n141) );
  OAI221_X1 r466_U94 ( .B1(fracta_mul[22]), .B2(r466_n34), .C1(fracta_mul[23]), 
        .C2(r466_n33), .A(r466_n141), .ZN(r466_n140) );
  NAND3_X1 r466_U93 ( .A1(r466_n61), .A2(r466_n62), .A3(r466_n140), .ZN(
        r466_n139) );
  OAI221_X1 r466_U92 ( .B1(fracta_mul[24]), .B2(r466_n32), .C1(fracta_mul[25]), 
        .C2(r466_n31), .A(r466_n139), .ZN(r466_n138) );
  NAND3_X1 r466_U91 ( .A1(r466_n137), .A2(r466_n63), .A3(r466_n138), .ZN(
        r466_n136) );
  OAI221_X1 r466_U90 ( .B1(fracta_mul[26]), .B2(r466_n30), .C1(fracta_mul[27]), 
        .C2(r466_n29), .A(r466_n136), .ZN(r466_n135) );
  NAND3_X1 r466_U89 ( .A1(r466_n133), .A2(r466_n134), .A3(r466_n135), .ZN(
        r466_n132) );
  OAI221_X1 r466_U88 ( .B1(fracta_mul[28]), .B2(r466_n28), .C1(fracta_mul[29]), 
        .C2(r466_n27), .A(r466_n132), .ZN(r466_n131) );
  NAND3_X1 r466_U87 ( .A1(r466_n129), .A2(r466_n130), .A3(r466_n131), .ZN(
        r466_n128) );
  OAI221_X1 r466_U86 ( .B1(fracta_mul[30]), .B2(r466_n26), .C1(fracta_mul[31]), 
        .C2(r466_n25), .A(r466_n128), .ZN(r466_n127) );
  NAND3_X1 r466_U85 ( .A1(r466_n125), .A2(r466_n126), .A3(r466_n127), .ZN(
        r466_n124) );
  OAI221_X1 r466_U84 ( .B1(fracta_mul[32]), .B2(r466_n24), .C1(fracta_mul[33]), 
        .C2(r466_n23), .A(r466_n124), .ZN(r466_n123) );
  NAND3_X1 r466_U83 ( .A1(r466_n121), .A2(r466_n122), .A3(r466_n123), .ZN(
        r466_n120) );
  OAI221_X1 r466_U82 ( .B1(fracta_mul[34]), .B2(r466_n22), .C1(fracta_mul[35]), 
        .C2(r466_n21), .A(r466_n120), .ZN(r466_n119) );
  NAND3_X1 r466_U81 ( .A1(r466_n117), .A2(r466_n118), .A3(r466_n119), .ZN(
        r466_n116) );
  OAI221_X1 r466_U80 ( .B1(fracta_mul[36]), .B2(r466_n20), .C1(fracta_mul[37]), 
        .C2(r466_n19), .A(r466_n116), .ZN(r466_n115) );
  NAND3_X1 r466_U79 ( .A1(r466_n113), .A2(r466_n114), .A3(r466_n115), .ZN(
        r466_n112) );
  OAI221_X1 r466_U78 ( .B1(fracta_mul[38]), .B2(r466_n18), .C1(fracta_mul[39]), 
        .C2(r466_n17), .A(r466_n112), .ZN(r466_n111) );
  NAND3_X1 r466_U77 ( .A1(r466_n109), .A2(r466_n110), .A3(r466_n111), .ZN(
        r466_n108) );
  OAI221_X1 r466_U76 ( .B1(fracta_mul[40]), .B2(r466_n16), .C1(fracta_mul[41]), 
        .C2(r466_n15), .A(r466_n108), .ZN(r466_n107) );
  NAND3_X1 r466_U75 ( .A1(r466_n105), .A2(r466_n106), .A3(r466_n107), .ZN(
        r466_n104) );
  OAI221_X1 r466_U74 ( .B1(fracta_mul[42]), .B2(r466_n14), .C1(fracta_mul[43]), 
        .C2(r466_n13), .A(r466_n104), .ZN(r466_n103) );
  NAND3_X1 r466_U73 ( .A1(r466_n101), .A2(r466_n102), .A3(r466_n103), .ZN(
        r466_n100) );
  OAI221_X1 r466_U72 ( .B1(fracta_mul[44]), .B2(r466_n12), .C1(fracta_mul[45]), 
        .C2(r466_n11), .A(r466_n100), .ZN(r466_n99) );
  NAND3_X1 r466_U71 ( .A1(r466_n97), .A2(r466_n98), .A3(r466_n99), .ZN(
        r466_n96) );
  OAI221_X1 r466_U70 ( .B1(fracta_mul[46]), .B2(r466_n10), .C1(fracta_mul[47]), 
        .C2(r466_n9), .A(r466_n96), .ZN(r466_n95) );
  NAND3_X1 r466_U69 ( .A1(r466_n93), .A2(r466_n94), .A3(r466_n95), .ZN(
        r466_n92) );
  OAI221_X1 r466_U68 ( .B1(fracta_mul[48]), .B2(r466_n8), .C1(fracta_mul[49]), 
        .C2(r466_n7), .A(r466_n92), .ZN(r466_n91) );
  AOI22_X1 r466_U67 ( .A1(u6_N50), .A2(r466_n1), .B1(r466_n90), .B2(r466_n91), 
        .ZN(r466_n89) );
  OAI22_X1 r466_U66 ( .A1(fracta_mul[51]), .A2(r466_n6), .B1(r466_n86), .B2(
        r466_n89), .ZN(u1_N324) );
  NOR4_X1 r466_U65 ( .A1(u1_N324), .A2(r466_n86), .A3(r466_n3), .A4(r466_n2), 
        .ZN(r466_n77) );
  AND3_X1 r466_U64 ( .A1(r466_n83), .A2(r466_n84), .A3(r466_n85), .ZN(r466_n79) );
  AND4_X1 r466_U63 ( .A1(r466_n79), .A2(r466_n80), .A3(r466_n81), .A4(r466_n82), .ZN(r466_n78) );
  NAND3_X1 r466_U62 ( .A1(r466_n76), .A2(r466_n77), .A3(r466_n78), .ZN(
        r466_n58) );
  AND4_X1 r466_U61 ( .A1(r466_n72), .A2(r466_n73), .A3(r466_n74), .A4(r466_n75), .ZN(r466_n71) );
  NAND4_X1 r466_U60 ( .A1(r466_n68), .A2(r466_n69), .A3(r466_n70), .A4(
        r466_n71), .ZN(r466_n59) );
  AND3_X1 r466_U59 ( .A1(r466_n65), .A2(r466_n66), .A3(r466_n67), .ZN(r466_n64) );
  NAND4_X1 r466_U58 ( .A1(r466_n61), .A2(r466_n62), .A3(r466_n63), .A4(
        r466_n64), .ZN(r466_n60) );
  NOR4_X1 r466_U57 ( .A1(r466_n57), .A2(r466_n58), .A3(r466_n59), .A4(r466_n60), .ZN(u1_N325) );
  INV_X4 r466_U56 ( .A(u6_N0), .ZN(r466_n56) );
  INV_X4 r466_U55 ( .A(u6_N1), .ZN(r466_n55) );
  INV_X4 r466_U54 ( .A(u6_N2), .ZN(r466_n54) );
  INV_X4 r466_U53 ( .A(u6_N3), .ZN(r466_n53) );
  INV_X4 r466_U52 ( .A(u6_N4), .ZN(r466_n52) );
  INV_X4 r466_U51 ( .A(u6_N5), .ZN(r466_n51) );
  INV_X4 r466_U50 ( .A(u6_N6), .ZN(r466_n50) );
  INV_X4 r466_U49 ( .A(u6_N7), .ZN(r466_n49) );
  INV_X4 r466_U48 ( .A(u6_N8), .ZN(r466_n48) );
  INV_X4 r466_U47 ( .A(u6_N9), .ZN(r466_n47) );
  INV_X4 r466_U46 ( .A(u6_N10), .ZN(r466_n46) );
  INV_X4 r466_U45 ( .A(u6_N11), .ZN(r466_n45) );
  INV_X4 r466_U44 ( .A(u6_N12), .ZN(r466_n44) );
  INV_X4 r466_U43 ( .A(u6_N13), .ZN(r466_n43) );
  INV_X4 r466_U42 ( .A(u6_N14), .ZN(r466_n42) );
  INV_X4 r466_U41 ( .A(u6_N15), .ZN(r466_n41) );
  INV_X4 r466_U40 ( .A(u6_N16), .ZN(r466_n40) );
  INV_X4 r466_U39 ( .A(u6_N17), .ZN(r466_n39) );
  INV_X4 r466_U38 ( .A(u6_N18), .ZN(r466_n38) );
  INV_X4 r466_U37 ( .A(u6_N19), .ZN(r466_n37) );
  INV_X4 r466_U36 ( .A(u6_N20), .ZN(r466_n36) );
  INV_X4 r466_U35 ( .A(u6_N21), .ZN(r466_n35) );
  INV_X4 r466_U34 ( .A(u6_N22), .ZN(r466_n34) );
  INV_X4 r466_U33 ( .A(u6_N23), .ZN(r466_n33) );
  INV_X4 r466_U32 ( .A(u6_N24), .ZN(r466_n32) );
  INV_X4 r466_U31 ( .A(u6_N25), .ZN(r466_n31) );
  INV_X4 r466_U30 ( .A(u6_N26), .ZN(r466_n30) );
  INV_X4 r466_U29 ( .A(u6_N27), .ZN(r466_n29) );
  INV_X4 r466_U28 ( .A(u6_N28), .ZN(r466_n28) );
  INV_X4 r466_U27 ( .A(u6_N29), .ZN(r466_n27) );
  INV_X4 r466_U26 ( .A(u6_N30), .ZN(r466_n26) );
  INV_X4 r466_U25 ( .A(u6_N31), .ZN(r466_n25) );
  INV_X4 r466_U24 ( .A(u6_N32), .ZN(r466_n24) );
  INV_X4 r466_U23 ( .A(u6_N33), .ZN(r466_n23) );
  INV_X4 r466_U22 ( .A(u6_N34), .ZN(r466_n22) );
  INV_X4 r466_U21 ( .A(u6_N35), .ZN(r466_n21) );
  INV_X4 r466_U20 ( .A(u6_N36), .ZN(r466_n20) );
  INV_X4 r466_U19 ( .A(u6_N37), .ZN(r466_n19) );
  INV_X4 r466_U18 ( .A(u6_N38), .ZN(r466_n18) );
  INV_X4 r466_U17 ( .A(u6_N39), .ZN(r466_n17) );
  INV_X4 r466_U16 ( .A(u6_N40), .ZN(r466_n16) );
  INV_X4 r466_U15 ( .A(u6_N41), .ZN(r466_n15) );
  INV_X4 r466_U14 ( .A(u6_N42), .ZN(r466_n14) );
  INV_X4 r466_U13 ( .A(u6_N43), .ZN(r466_n13) );
  INV_X4 r466_U12 ( .A(u6_N44), .ZN(r466_n12) );
  INV_X4 r466_U11 ( .A(u6_N45), .ZN(r466_n11) );
  INV_X4 r466_U10 ( .A(u6_N46), .ZN(r466_n10) );
  INV_X4 r466_U9 ( .A(u6_N47), .ZN(r466_n9) );
  INV_X4 r466_U8 ( .A(u6_N48), .ZN(r466_n8) );
  INV_X4 r466_U7 ( .A(u6_N49), .ZN(r466_n7) );
  INV_X4 r466_U6 ( .A(u6_N51), .ZN(r466_n6) );
  INV_X4 r466_U5 ( .A(r466_n165), .ZN(r466_n5) );
  INV_X4 r466_U4 ( .A(fracta_mul[1]), .ZN(r466_n4) );
  INV_X4 r466_U3 ( .A(r466_n88), .ZN(r466_n3) );
  INV_X4 r466_U2 ( .A(r466_n87), .ZN(r466_n2) );
  INV_X4 r466_U1 ( .A(fracta_mul[50]), .ZN(r466_n1) );
  XOR2_X2 add_0_root_sub_0_root_u4_add_495_U2 ( .A(u4_ldz_dif_0_), .B(n4823), 
        .Z(u4_div_exp3[0]) );
  AND2_X4 add_0_root_sub_0_root_u4_add_495_U1 ( .A1(u4_ldz_dif_0_), .A2(n4823), 
        .ZN(add_0_root_sub_0_root_u4_add_495_n1) );
  FA_X1 add_0_root_sub_0_root_u4_add_495_U1_1 ( .A(n4368), .B(u4_ldz_dif_1_), 
        .CI(add_0_root_sub_0_root_u4_add_495_n1), .CO(
        add_0_root_sub_0_root_u4_add_495_carry[2]), .S(u4_div_exp3[1]) );
  FA_X1 add_0_root_sub_0_root_u4_add_495_U1_2 ( .A(exp_r[2]), .B(u4_ldz_dif_2_), .CI(add_0_root_sub_0_root_u4_add_495_carry[2]), .CO(
        add_0_root_sub_0_root_u4_add_495_carry[3]), .S(u4_div_exp3[2]) );
  FA_X1 add_0_root_sub_0_root_u4_add_495_U1_3 ( .A(exp_r[3]), .B(u4_ldz_dif_3_), .CI(add_0_root_sub_0_root_u4_add_495_carry[3]), .CO(
        add_0_root_sub_0_root_u4_add_495_carry[4]), .S(u4_div_exp3[3]) );
  FA_X1 add_0_root_sub_0_root_u4_add_495_U1_4 ( .A(n4399), .B(u4_ldz_dif_4_), 
        .CI(add_0_root_sub_0_root_u4_add_495_carry[4]), .CO(
        add_0_root_sub_0_root_u4_add_495_carry[5]), .S(u4_div_exp3[4]) );
  FA_X1 add_0_root_sub_0_root_u4_add_495_U1_5 ( .A(n4370), .B(u4_ldz_dif_5_), 
        .CI(add_0_root_sub_0_root_u4_add_495_carry[5]), .CO(
        add_0_root_sub_0_root_u4_add_495_carry[6]), .S(u4_div_exp3[5]) );
  FA_X1 add_0_root_sub_0_root_u4_add_495_U1_6 ( .A(n4382), .B(u4_ldz_dif_6_), 
        .CI(add_0_root_sub_0_root_u4_add_495_carry[6]), .CO(
        add_0_root_sub_0_root_u4_add_495_carry[7]), .S(u4_div_exp3[6]) );
  FA_X1 add_0_root_sub_0_root_u4_add_495_U1_7 ( .A(n4359), .B(u4_ldz_dif_7_), 
        .CI(add_0_root_sub_0_root_u4_add_495_carry[7]), .CO(
        add_0_root_sub_0_root_u4_add_495_carry[8]), .S(u4_div_exp3[7]) );
  FA_X1 add_0_root_sub_0_root_u4_add_495_U1_8 ( .A(n4369), .B(n4480), .CI(
        add_0_root_sub_0_root_u4_add_495_carry[8]), .CO(
        add_0_root_sub_0_root_u4_add_495_carry[9]), .S(u4_div_exp3[8]) );
  FA_X1 add_0_root_sub_0_root_u4_add_495_U1_9 ( .A(n4428), .B(n4480), .CI(
        add_0_root_sub_0_root_u4_add_495_carry[9]), .CO(
        add_0_root_sub_0_root_u4_add_495_carry[10]), .S(u4_div_exp3[9]) );
  FA_X1 add_0_root_sub_0_root_u4_add_495_U1_10 ( .A(n4875), .B(n4480), .CI(
        add_0_root_sub_0_root_u4_add_495_carry[10]), .S(u4_div_exp3[10]) );
  NOR2_X1 u5_mult_87_U3292 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n339), .ZN(
        u5_N0) );
  NOR2_X1 u5_mult_87_U3291 ( .A1(u5_mult_87_n428), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__10_) );
  NOR2_X1 u5_mult_87_U3290 ( .A1(u5_mult_87_n425), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__11_) );
  NOR2_X1 u5_mult_87_U3289 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__12_) );
  NOR2_X1 u5_mult_87_U3288 ( .A1(u5_mult_87_n422), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__13_) );
  NOR2_X1 u5_mult_87_U3287 ( .A1(u5_mult_87_n418), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__14_) );
  NOR2_X1 u5_mult_87_U3286 ( .A1(u5_mult_87_n416), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__15_) );
  NOR2_X1 u5_mult_87_U3285 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__16_) );
  NOR2_X1 u5_mult_87_U3284 ( .A1(u5_mult_87_n413), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__17_) );
  NOR2_X1 u5_mult_87_U3283 ( .A1(u5_mult_87_n411), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__18_) );
  NOR2_X1 u5_mult_87_U3282 ( .A1(u5_mult_87_n409), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__19_) );
  NOR2_X1 u5_mult_87_U3281 ( .A1(u5_mult_87_n446), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__1_) );
  NOR2_X1 u5_mult_87_U3280 ( .A1(u5_mult_87_n407), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__20_) );
  NOR2_X1 u5_mult_87_U3279 ( .A1(u5_mult_87_n406), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__21_) );
  NOR2_X1 u5_mult_87_U3278 ( .A1(u5_mult_87_n404), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__22_) );
  NOR2_X1 u5_mult_87_U3277 ( .A1(u5_mult_87_n402), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__23_) );
  NOR2_X1 u5_mult_87_U3276 ( .A1(u5_mult_87_n399), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__24_) );
  NOR2_X1 u5_mult_87_U3275 ( .A1(u5_mult_87_n398), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__25_) );
  NOR2_X1 u5_mult_87_U3274 ( .A1(u5_mult_87_n395), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__26_) );
  NOR2_X1 u5_mult_87_U3273 ( .A1(u5_mult_87_n394), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__27_) );
  NOR2_X1 u5_mult_87_U3272 ( .A1(u5_mult_87_n392), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__28_) );
  NOR2_X1 u5_mult_87_U3271 ( .A1(u5_mult_87_n390), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__29_) );
  NOR2_X1 u5_mult_87_U3270 ( .A1(u5_mult_87_n444), .A2(u5_mult_87_n340), .ZN(
        u5_mult_87_ab_0__2_) );
  NOR2_X1 u5_mult_87_U3269 ( .A1(u5_mult_87_n387), .A2(u5_mult_87_n340), .ZN(
        u5_mult_87_ab_0__30_) );
  NOR2_X1 u5_mult_87_U3268 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n340), .ZN(
        u5_mult_87_ab_0__31_) );
  NOR2_X1 u5_mult_87_U3267 ( .A1(u5_mult_87_n383), .A2(u5_mult_87_n340), .ZN(
        u5_mult_87_ab_0__32_) );
  NOR2_X1 u5_mult_87_U3266 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n340), .ZN(
        u5_mult_87_ab_0__33_) );
  NOR2_X1 u5_mult_87_U3265 ( .A1(u5_mult_87_n379), .A2(u5_mult_87_n340), .ZN(
        u5_mult_87_ab_0__34_) );
  NOR2_X1 u5_mult_87_U3264 ( .A1(u5_mult_87_n377), .A2(u5_mult_87_n340), .ZN(
        u5_mult_87_ab_0__35_) );
  NOR2_X1 u5_mult_87_U3263 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n340), .ZN(
        u5_mult_87_ab_0__36_) );
  NOR2_X1 u5_mult_87_U3262 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n340), .ZN(
        u5_mult_87_ab_0__37_) );
  NOR2_X1 u5_mult_87_U3261 ( .A1(u5_mult_87_n372), .A2(u5_mult_87_n340), .ZN(
        u5_mult_87_ab_0__38_) );
  NOR2_X1 u5_mult_87_U3260 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n340), .ZN(
        u5_mult_87_ab_0__39_) );
  NOR2_X1 u5_mult_87_U3259 ( .A1(u5_mult_87_n442), .A2(u5_mult_87_n341), .ZN(
        u5_mult_87_ab_0__3_) );
  NOR2_X1 u5_mult_87_U3258 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n341), .ZN(
        u5_mult_87_ab_0__40_) );
  NOR2_X1 u5_mult_87_U3257 ( .A1(u5_mult_87_n365), .A2(u5_mult_87_n341), .ZN(
        u5_mult_87_ab_0__41_) );
  NOR2_X1 u5_mult_87_U3256 ( .A1(u5_mult_87_n363), .A2(u5_mult_87_n341), .ZN(
        u5_mult_87_ab_0__42_) );
  NOR2_X1 u5_mult_87_U3255 ( .A1(u5_mult_87_n360), .A2(u5_mult_87_n341), .ZN(
        u5_mult_87_ab_0__43_) );
  NOR2_X1 u5_mult_87_U3254 ( .A1(u5_mult_87_n358), .A2(u5_mult_87_n341), .ZN(
        u5_mult_87_ab_0__44_) );
  NOR2_X1 u5_mult_87_U3253 ( .A1(u5_mult_87_n356), .A2(u5_mult_87_n341), .ZN(
        u5_mult_87_ab_0__45_) );
  NOR2_X1 u5_mult_87_U3252 ( .A1(u5_mult_87_n354), .A2(u5_mult_87_n341), .ZN(
        u5_mult_87_ab_0__46_) );
  NOR2_X1 u5_mult_87_U3251 ( .A1(u5_mult_87_n353), .A2(u5_mult_87_n341), .ZN(
        u5_mult_87_ab_0__47_) );
  NOR2_X1 u5_mult_87_U3250 ( .A1(u5_mult_87_n350), .A2(u5_mult_87_n341), .ZN(
        u5_mult_87_ab_0__48_) );
  NOR2_X1 u5_mult_87_U3249 ( .A1(u5_mult_87_n348), .A2(u5_mult_87_n341), .ZN(
        u5_mult_87_ab_0__49_) );
  NOR2_X1 u5_mult_87_U3248 ( .A1(u5_mult_87_n440), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__4_) );
  NOR2_X1 u5_mult_87_U3247 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n340), .ZN(
        u5_mult_87_ab_0__50_) );
  NOR2_X1 u5_mult_87_U3246 ( .A1(u5_mult_87_n345), .A2(u5_mult_87_n341), .ZN(
        u5_mult_87_ab_0__51_) );
  NOR2_X1 u5_mult_87_U3245 ( .A1(u5_mult_87_n342), .A2(u5_mult_87_n341), .ZN(
        u5_mult_87_ab_0__52_) );
  NOR2_X1 u5_mult_87_U3244 ( .A1(u5_mult_87_n437), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__5_) );
  NOR2_X1 u5_mult_87_U3243 ( .A1(u5_mult_87_n436), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__6_) );
  NOR2_X1 u5_mult_87_U3242 ( .A1(u5_mult_87_n434), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__7_) );
  NOR2_X1 u5_mult_87_U3241 ( .A1(u5_mult_87_n432), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__8_) );
  NOR2_X1 u5_mult_87_U3240 ( .A1(u5_mult_87_n430), .A2(u5_mult_87_n339), .ZN(
        u5_mult_87_ab_0__9_) );
  NOR2_X1 u5_mult_87_U3239 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__0_) );
  NOR2_X1 u5_mult_87_U3238 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__10_) );
  NOR2_X1 u5_mult_87_U3237 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__11_) );
  NOR2_X1 u5_mult_87_U3236 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__12_) );
  NOR2_X1 u5_mult_87_U3235 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__13_) );
  NOR2_X1 u5_mult_87_U3234 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__14_) );
  NOR2_X1 u5_mult_87_U3233 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__15_) );
  NOR2_X1 u5_mult_87_U3232 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__16_) );
  NOR2_X1 u5_mult_87_U3231 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__17_) );
  NOR2_X1 u5_mult_87_U3230 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__18_) );
  NOR2_X1 u5_mult_87_U3229 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__19_) );
  NOR2_X1 u5_mult_87_U3228 ( .A1(u5_mult_87_n446), .A2(u5_mult_87_n311), .ZN(
        u5_mult_87_ab_10__1_) );
  NOR2_X1 u5_mult_87_U3227 ( .A1(u5_mult_87_n407), .A2(u5_mult_87_n311), .ZN(
        u5_mult_87_ab_10__20_) );
  NOR2_X1 u5_mult_87_U3226 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n311), .ZN(
        u5_mult_87_ab_10__21_) );
  NOR2_X1 u5_mult_87_U3225 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n311), .ZN(
        u5_mult_87_ab_10__22_) );
  NOR2_X1 u5_mult_87_U3224 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n311), .ZN(
        u5_mult_87_ab_10__23_) );
  NOR2_X1 u5_mult_87_U3223 ( .A1(u5_mult_87_n399), .A2(u5_mult_87_n311), .ZN(
        u5_mult_87_ab_10__24_) );
  NOR2_X1 u5_mult_87_U3222 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n311), .ZN(
        u5_mult_87_ab_10__25_) );
  NOR2_X1 u5_mult_87_U3221 ( .A1(u5_mult_87_n395), .A2(u5_mult_87_n311), .ZN(
        u5_mult_87_ab_10__26_) );
  NOR2_X1 u5_mult_87_U3220 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n311), .ZN(
        u5_mult_87_ab_10__27_) );
  NOR2_X1 u5_mult_87_U3219 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n311), .ZN(
        u5_mult_87_ab_10__28_) );
  NOR2_X1 u5_mult_87_U3218 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n311), .ZN(
        u5_mult_87_ab_10__29_) );
  NOR2_X1 u5_mult_87_U3217 ( .A1(u5_mult_87_n444), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__2_) );
  NOR2_X1 u5_mult_87_U3216 ( .A1(u5_mult_87_n387), .A2(u5_mult_87_n311), .ZN(
        u5_mult_87_ab_10__30_) );
  NOR2_X1 u5_mult_87_U3215 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n311), .ZN(
        u5_mult_87_ab_10__31_) );
  NOR2_X1 u5_mult_87_U3214 ( .A1(u5_mult_87_n383), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__32_) );
  NOR2_X1 u5_mult_87_U3213 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n311), .ZN(
        u5_mult_87_ab_10__33_) );
  NOR2_X1 u5_mult_87_U3212 ( .A1(u5_mult_87_n379), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__34_) );
  NOR2_X1 u5_mult_87_U3211 ( .A1(u5_mult_87_n377), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__35_) );
  NOR2_X1 u5_mult_87_U3210 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__36_) );
  NOR2_X1 u5_mult_87_U3209 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__37_) );
  NOR2_X1 u5_mult_87_U3208 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__38_) );
  NOR2_X1 u5_mult_87_U3207 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__39_) );
  NOR2_X1 u5_mult_87_U3206 ( .A1(u5_mult_87_n442), .A2(u5_mult_87_n475), .ZN(
        u5_mult_87_ab_10__3_) );
  NOR2_X1 u5_mult_87_U3205 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n475), .ZN(
        u5_mult_87_ab_10__40_) );
  NOR2_X1 u5_mult_87_U3204 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n475), .ZN(
        u5_mult_87_ab_10__41_) );
  NOR2_X1 u5_mult_87_U3203 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n475), .ZN(
        u5_mult_87_ab_10__42_) );
  NOR2_X1 u5_mult_87_U3202 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n311), .ZN(
        u5_mult_87_ab_10__43_) );
  NOR2_X1 u5_mult_87_U3201 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n475), .ZN(
        u5_mult_87_ab_10__44_) );
  NOR2_X1 u5_mult_87_U3200 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n475), .ZN(
        u5_mult_87_ab_10__45_) );
  NOR2_X1 u5_mult_87_U3199 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n475), .ZN(
        u5_mult_87_ab_10__46_) );
  NOR2_X1 u5_mult_87_U3198 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n475), .ZN(
        u5_mult_87_ab_10__47_) );
  NOR2_X1 u5_mult_87_U3197 ( .A1(u5_mult_87_n350), .A2(u5_mult_87_n475), .ZN(
        u5_mult_87_ab_10__48_) );
  NOR2_X1 u5_mult_87_U3196 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n475), .ZN(
        u5_mult_87_ab_10__49_) );
  NOR2_X1 u5_mult_87_U3195 ( .A1(u5_mult_87_n440), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__4_) );
  NOR2_X1 u5_mult_87_U3194 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n311), .ZN(
        u5_mult_87_ab_10__50_) );
  NOR2_X1 u5_mult_87_U3193 ( .A1(u5_mult_87_n345), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__51_) );
  NOR2_X1 u5_mult_87_U3192 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__52_) );
  NOR2_X1 u5_mult_87_U3191 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__5_) );
  NOR2_X1 u5_mult_87_U3190 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__6_) );
  NOR2_X1 u5_mult_87_U3189 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__7_) );
  NOR2_X1 u5_mult_87_U3188 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__8_) );
  NOR2_X1 u5_mult_87_U3187 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n310), .ZN(
        u5_mult_87_ab_10__9_) );
  NOR2_X1 u5_mult_87_U3186 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__0_) );
  NOR2_X1 u5_mult_87_U3185 ( .A1(u5_mult_87_n428), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__10_) );
  NOR2_X1 u5_mult_87_U3184 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__11_) );
  NOR2_X1 u5_mult_87_U3183 ( .A1(u5_mult_87_n481), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__12_) );
  NOR2_X1 u5_mult_87_U3182 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__13_) );
  NOR2_X1 u5_mult_87_U3181 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__14_) );
  NOR2_X1 u5_mult_87_U3180 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__15_) );
  NOR2_X1 u5_mult_87_U3179 ( .A1(u5_mult_87_n480), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__16_) );
  NOR2_X1 u5_mult_87_U3178 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__17_) );
  NOR2_X1 u5_mult_87_U3177 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__18_) );
  NOR2_X1 u5_mult_87_U3176 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__19_) );
  NOR2_X1 u5_mult_87_U3175 ( .A1(u5_mult_87_n446), .A2(u5_mult_87_n309), .ZN(
        u5_mult_87_ab_11__1_) );
  NOR2_X1 u5_mult_87_U3174 ( .A1(u5_mult_87_n407), .A2(u5_mult_87_n309), .ZN(
        u5_mult_87_ab_11__20_) );
  NOR2_X1 u5_mult_87_U3173 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n309), .ZN(
        u5_mult_87_ab_11__21_) );
  NOR2_X1 u5_mult_87_U3172 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n309), .ZN(
        u5_mult_87_ab_11__22_) );
  NOR2_X1 u5_mult_87_U3171 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n309), .ZN(
        u5_mult_87_ab_11__23_) );
  NOR2_X1 u5_mult_87_U3170 ( .A1(u5_mult_87_n399), .A2(u5_mult_87_n309), .ZN(
        u5_mult_87_ab_11__24_) );
  NOR2_X1 u5_mult_87_U3169 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n309), .ZN(
        u5_mult_87_ab_11__25_) );
  NOR2_X1 u5_mult_87_U3168 ( .A1(u5_mult_87_n395), .A2(u5_mult_87_n309), .ZN(
        u5_mult_87_ab_11__26_) );
  NOR2_X1 u5_mult_87_U3167 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n309), .ZN(
        u5_mult_87_ab_11__27_) );
  NOR2_X1 u5_mult_87_U3166 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n309), .ZN(
        u5_mult_87_ab_11__28_) );
  NOR2_X1 u5_mult_87_U3165 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n309), .ZN(
        u5_mult_87_ab_11__29_) );
  NOR2_X1 u5_mult_87_U3164 ( .A1(u5_mult_87_n444), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__2_) );
  NOR2_X1 u5_mult_87_U3163 ( .A1(u5_mult_87_n387), .A2(u5_mult_87_n309), .ZN(
        u5_mult_87_ab_11__30_) );
  NOR2_X1 u5_mult_87_U3162 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n309), .ZN(
        u5_mult_87_ab_11__31_) );
  NOR2_X1 u5_mult_87_U3161 ( .A1(u5_mult_87_n383), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__32_) );
  NOR2_X1 u5_mult_87_U3160 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__33_) );
  NOR2_X1 u5_mult_87_U3159 ( .A1(u5_mult_87_n379), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__34_) );
  NOR2_X1 u5_mult_87_U3158 ( .A1(u5_mult_87_n377), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__35_) );
  NOR2_X1 u5_mult_87_U3157 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__36_) );
  NOR2_X1 u5_mult_87_U3156 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__37_) );
  NOR2_X1 u5_mult_87_U3155 ( .A1(u5_mult_87_n372), .A2(u5_mult_87_n309), .ZN(
        u5_mult_87_ab_11__38_) );
  NOR2_X1 u5_mult_87_U3154 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n309), .ZN(
        u5_mult_87_ab_11__39_) );
  NOR2_X1 u5_mult_87_U3153 ( .A1(u5_mult_87_n442), .A2(u5_mult_87_n474), .ZN(
        u5_mult_87_ab_11__3_) );
  NOR2_X1 u5_mult_87_U3152 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n474), .ZN(
        u5_mult_87_ab_11__40_) );
  NOR2_X1 u5_mult_87_U3151 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n474), .ZN(
        u5_mult_87_ab_11__41_) );
  NOR2_X1 u5_mult_87_U3150 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n474), .ZN(
        u5_mult_87_ab_11__42_) );
  NOR2_X1 u5_mult_87_U3149 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n474), .ZN(
        u5_mult_87_ab_11__43_) );
  NOR2_X1 u5_mult_87_U3148 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n474), .ZN(
        u5_mult_87_ab_11__44_) );
  NOR2_X1 u5_mult_87_U3147 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n474), .ZN(
        u5_mult_87_ab_11__45_) );
  NOR2_X1 u5_mult_87_U3146 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n474), .ZN(
        u5_mult_87_ab_11__46_) );
  NOR2_X1 u5_mult_87_U3145 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n309), .ZN(
        u5_mult_87_ab_11__47_) );
  NOR2_X1 u5_mult_87_U3144 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n309), .ZN(
        u5_mult_87_ab_11__48_) );
  NOR2_X1 u5_mult_87_U3143 ( .A1(u5_mult_87_n348), .A2(u5_mult_87_n474), .ZN(
        u5_mult_87_ab_11__49_) );
  NOR2_X1 u5_mult_87_U3142 ( .A1(u5_mult_87_n440), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__4_) );
  NOR2_X1 u5_mult_87_U3141 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n309), .ZN(
        u5_mult_87_ab_11__50_) );
  NOR2_X1 u5_mult_87_U3140 ( .A1(u5_mult_87_n345), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__51_) );
  NOR2_X1 u5_mult_87_U3139 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__52_) );
  NOR2_X1 u5_mult_87_U3138 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__5_) );
  NOR2_X1 u5_mult_87_U3137 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__6_) );
  NOR2_X1 u5_mult_87_U3136 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__7_) );
  NOR2_X1 u5_mult_87_U3135 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__8_) );
  NOR2_X1 u5_mult_87_U3134 ( .A1(u5_mult_87_n430), .A2(u5_mult_87_n308), .ZN(
        u5_mult_87_ab_11__9_) );
  NOR2_X1 u5_mult_87_U3133 ( .A1(u5_mult_87_n450), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__0_) );
  NOR2_X1 u5_mult_87_U3132 ( .A1(u5_mult_87_n428), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__10_) );
  NOR2_X1 u5_mult_87_U3131 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__11_) );
  NOR2_X1 u5_mult_87_U3130 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__12_) );
  NOR2_X1 u5_mult_87_U3129 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__13_) );
  NOR2_X1 u5_mult_87_U3128 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__14_) );
  NOR2_X1 u5_mult_87_U3127 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__15_) );
  NOR2_X1 u5_mult_87_U3126 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__16_) );
  NOR2_X1 u5_mult_87_U3125 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__17_) );
  NOR2_X1 u5_mult_87_U3124 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__18_) );
  NOR2_X1 u5_mult_87_U3123 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__19_) );
  NOR2_X1 u5_mult_87_U3122 ( .A1(u5_mult_87_n446), .A2(u5_mult_87_n306), .ZN(
        u5_mult_87_ab_12__1_) );
  NOR2_X1 u5_mult_87_U3121 ( .A1(u5_mult_87_n407), .A2(u5_mult_87_n306), .ZN(
        u5_mult_87_ab_12__20_) );
  NOR2_X1 u5_mult_87_U3120 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n306), .ZN(
        u5_mult_87_ab_12__21_) );
  NOR2_X1 u5_mult_87_U3119 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n306), .ZN(
        u5_mult_87_ab_12__22_) );
  NOR2_X1 u5_mult_87_U3118 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n306), .ZN(
        u5_mult_87_ab_12__23_) );
  NOR2_X1 u5_mult_87_U3117 ( .A1(u5_mult_87_n399), .A2(u5_mult_87_n306), .ZN(
        u5_mult_87_ab_12__24_) );
  NOR2_X1 u5_mult_87_U3116 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n306), .ZN(
        u5_mult_87_ab_12__25_) );
  NOR2_X1 u5_mult_87_U3115 ( .A1(u5_mult_87_n395), .A2(u5_mult_87_n306), .ZN(
        u5_mult_87_ab_12__26_) );
  NOR2_X1 u5_mult_87_U3114 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n306), .ZN(
        u5_mult_87_ab_12__27_) );
  NOR2_X1 u5_mult_87_U3113 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n306), .ZN(
        u5_mult_87_ab_12__28_) );
  NOR2_X1 u5_mult_87_U3112 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n306), .ZN(
        u5_mult_87_ab_12__29_) );
  NOR2_X1 u5_mult_87_U3111 ( .A1(u5_mult_87_n444), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__2_) );
  NOR2_X1 u5_mult_87_U3110 ( .A1(u5_mult_87_n387), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__30_) );
  NOR2_X1 u5_mult_87_U3109 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__31_) );
  NOR2_X1 u5_mult_87_U3108 ( .A1(u5_mult_87_n383), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__32_) );
  NOR2_X1 u5_mult_87_U3107 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__33_) );
  NOR2_X1 u5_mult_87_U3106 ( .A1(u5_mult_87_n379), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__34_) );
  NOR2_X1 u5_mult_87_U3105 ( .A1(u5_mult_87_n377), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__35_) );
  NOR2_X1 u5_mult_87_U3104 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n306), .ZN(
        u5_mult_87_ab_12__36_) );
  NOR2_X1 u5_mult_87_U3103 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n306), .ZN(
        u5_mult_87_ab_12__37_) );
  NOR2_X1 u5_mult_87_U3102 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n306), .ZN(
        u5_mult_87_ab_12__38_) );
  NOR2_X1 u5_mult_87_U3101 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n306), .ZN(
        u5_mult_87_ab_12__39_) );
  NOR2_X1 u5_mult_87_U3100 ( .A1(u5_mult_87_n442), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__3_) );
  NOR2_X1 u5_mult_87_U3099 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n473), .ZN(
        u5_mult_87_ab_12__40_) );
  NOR2_X1 u5_mult_87_U3098 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n473), .ZN(
        u5_mult_87_ab_12__41_) );
  NOR2_X1 u5_mult_87_U3097 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n473), .ZN(
        u5_mult_87_ab_12__42_) );
  NOR2_X1 u5_mult_87_U3096 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n473), .ZN(
        u5_mult_87_ab_12__43_) );
  NOR2_X1 u5_mult_87_U3095 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n473), .ZN(
        u5_mult_87_ab_12__44_) );
  NOR2_X1 u5_mult_87_U3094 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n473), .ZN(
        u5_mult_87_ab_12__45_) );
  NOR2_X1 u5_mult_87_U3093 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n473), .ZN(
        u5_mult_87_ab_12__46_) );
  NOR2_X1 u5_mult_87_U3092 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n473), .ZN(
        u5_mult_87_ab_12__47_) );
  NOR2_X1 u5_mult_87_U3091 ( .A1(u5_mult_87_n350), .A2(u5_mult_87_n473), .ZN(
        u5_mult_87_ab_12__48_) );
  NOR2_X1 u5_mult_87_U3090 ( .A1(u5_mult_87_n348), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__49_) );
  NOR2_X1 u5_mult_87_U3089 ( .A1(u5_mult_87_n440), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__4_) );
  NOR2_X1 u5_mult_87_U3088 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__50_) );
  NOR2_X1 u5_mult_87_U3087 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__51_) );
  NOR2_X1 u5_mult_87_U3086 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__52_) );
  NOR2_X1 u5_mult_87_U3085 ( .A1(u5_mult_87_n439), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__5_) );
  NOR2_X1 u5_mult_87_U3084 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__6_) );
  NOR2_X1 u5_mult_87_U3083 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__7_) );
  NOR2_X1 u5_mult_87_U3082 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__8_) );
  NOR2_X1 u5_mult_87_U3081 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n307), .ZN(
        u5_mult_87_ab_12__9_) );
  NOR2_X1 u5_mult_87_U3080 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__0_) );
  NOR2_X1 u5_mult_87_U3079 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__10_) );
  NOR2_X1 u5_mult_87_U3078 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__11_) );
  NOR2_X1 u5_mult_87_U3077 ( .A1(u5_mult_87_n481), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__12_) );
  NOR2_X1 u5_mult_87_U3076 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__13_) );
  NOR2_X1 u5_mult_87_U3075 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__14_) );
  NOR2_X1 u5_mult_87_U3074 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__15_) );
  NOR2_X1 u5_mult_87_U3073 ( .A1(u5_mult_87_n480), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__16_) );
  NOR2_X1 u5_mult_87_U3072 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__17_) );
  NOR2_X1 u5_mult_87_U3071 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__18_) );
  NOR2_X1 u5_mult_87_U3070 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__19_) );
  NOR2_X1 u5_mult_87_U3069 ( .A1(u5_mult_87_n446), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__1_) );
  NOR2_X1 u5_mult_87_U3068 ( .A1(u5_mult_87_n407), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__20_) );
  NOR2_X1 u5_mult_87_U3067 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__21_) );
  NOR2_X1 u5_mult_87_U3066 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__22_) );
  NOR2_X1 u5_mult_87_U3065 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__23_) );
  NOR2_X1 u5_mult_87_U3064 ( .A1(u5_mult_87_n399), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__24_) );
  NOR2_X1 u5_mult_87_U3063 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__25_) );
  NOR2_X1 u5_mult_87_U3062 ( .A1(u5_mult_87_n395), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__26_) );
  NOR2_X1 u5_mult_87_U3061 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__27_) );
  NOR2_X1 u5_mult_87_U3060 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__28_) );
  NOR2_X1 u5_mult_87_U3059 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__29_) );
  NOR2_X1 u5_mult_87_U3058 ( .A1(u5_mult_87_n444), .A2(u5_mult_87_n305), .ZN(
        u5_mult_87_ab_13__2_) );
  NOR2_X1 u5_mult_87_U3057 ( .A1(u5_mult_87_n387), .A2(u5_mult_87_n305), .ZN(
        u5_mult_87_ab_13__30_) );
  NOR2_X1 u5_mult_87_U3056 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__31_) );
  NOR2_X1 u5_mult_87_U3055 ( .A1(u5_mult_87_n383), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__32_) );
  NOR2_X1 u5_mult_87_U3054 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__33_) );
  NOR2_X1 u5_mult_87_U3053 ( .A1(u5_mult_87_n379), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__34_) );
  NOR2_X1 u5_mult_87_U3052 ( .A1(u5_mult_87_n377), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__35_) );
  NOR2_X1 u5_mult_87_U3051 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n305), .ZN(
        u5_mult_87_ab_13__36_) );
  NOR2_X1 u5_mult_87_U3050 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n305), .ZN(
        u5_mult_87_ab_13__37_) );
  NOR2_X1 u5_mult_87_U3049 ( .A1(u5_mult_87_n372), .A2(u5_mult_87_n305), .ZN(
        u5_mult_87_ab_13__38_) );
  NOR2_X1 u5_mult_87_U3048 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n305), .ZN(
        u5_mult_87_ab_13__39_) );
  NOR2_X1 u5_mult_87_U3047 ( .A1(u5_mult_87_n442), .A2(u5_mult_87_n305), .ZN(
        u5_mult_87_ab_13__3_) );
  NOR2_X1 u5_mult_87_U3046 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n305), .ZN(
        u5_mult_87_ab_13__40_) );
  NOR2_X1 u5_mult_87_U3045 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n305), .ZN(
        u5_mult_87_ab_13__41_) );
  NOR2_X1 u5_mult_87_U3044 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n305), .ZN(
        u5_mult_87_ab_13__42_) );
  NOR2_X1 u5_mult_87_U3043 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n305), .ZN(
        u5_mult_87_ab_13__43_) );
  NOR2_X1 u5_mult_87_U3042 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n305), .ZN(
        u5_mult_87_ab_13__44_) );
  NOR2_X1 u5_mult_87_U3041 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n305), .ZN(
        u5_mult_87_ab_13__45_) );
  NOR2_X1 u5_mult_87_U3040 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n305), .ZN(
        u5_mult_87_ab_13__46_) );
  NOR2_X1 u5_mult_87_U3039 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n305), .ZN(
        u5_mult_87_ab_13__47_) );
  NOR2_X1 u5_mult_87_U3038 ( .A1(u5_mult_87_n350), .A2(u5_mult_87_n305), .ZN(
        u5_mult_87_ab_13__48_) );
  NOR2_X1 u5_mult_87_U3037 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n305), .ZN(
        u5_mult_87_ab_13__49_) );
  NOR2_X1 u5_mult_87_U3036 ( .A1(u5_mult_87_n440), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__4_) );
  NOR2_X1 u5_mult_87_U3035 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__50_) );
  NOR2_X1 u5_mult_87_U3034 ( .A1(u5_mult_87_n345), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__51_) );
  NOR2_X1 u5_mult_87_U3033 ( .A1(u5_mult_87_n342), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__52_) );
  NOR2_X1 u5_mult_87_U3032 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__5_) );
  NOR2_X1 u5_mult_87_U3031 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__6_) );
  NOR2_X1 u5_mult_87_U3030 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__7_) );
  NOR2_X1 u5_mult_87_U3029 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__8_) );
  NOR2_X1 u5_mult_87_U3028 ( .A1(u5_mult_87_n430), .A2(u5_mult_87_n304), .ZN(
        u5_mult_87_ab_13__9_) );
  NOR2_X1 u5_mult_87_U3027 ( .A1(u5_mult_87_n450), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__0_) );
  NOR2_X1 u5_mult_87_U3026 ( .A1(u5_mult_87_n428), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__10_) );
  NOR2_X1 u5_mult_87_U3025 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__11_) );
  NOR2_X1 u5_mult_87_U3024 ( .A1(u5_mult_87_n481), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__12_) );
  NOR2_X1 u5_mult_87_U3023 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__13_) );
  NOR2_X1 u5_mult_87_U3022 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__14_) );
  NOR2_X1 u5_mult_87_U3021 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__15_) );
  NOR2_X1 u5_mult_87_U3020 ( .A1(u5_mult_87_n480), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__16_) );
  NOR2_X1 u5_mult_87_U3019 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__17_) );
  NOR2_X1 u5_mult_87_U3018 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__18_) );
  NOR2_X1 u5_mult_87_U3017 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__19_) );
  NOR2_X1 u5_mult_87_U3016 ( .A1(u5_mult_87_n446), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__1_) );
  NOR2_X1 u5_mult_87_U3015 ( .A1(u5_mult_87_n407), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__20_) );
  NOR2_X1 u5_mult_87_U3014 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__21_) );
  NOR2_X1 u5_mult_87_U3013 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__22_) );
  NOR2_X1 u5_mult_87_U3012 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__23_) );
  NOR2_X1 u5_mult_87_U3011 ( .A1(u5_mult_87_n399), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__24_) );
  NOR2_X1 u5_mult_87_U3010 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__25_) );
  NOR2_X1 u5_mult_87_U3009 ( .A1(u5_mult_87_n395), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__26_) );
  NOR2_X1 u5_mult_87_U3008 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__27_) );
  NOR2_X1 u5_mult_87_U3007 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__28_) );
  NOR2_X1 u5_mult_87_U3006 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__29_) );
  NOR2_X1 u5_mult_87_U3005 ( .A1(u5_mult_87_n444), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__2_) );
  NOR2_X1 u5_mult_87_U3004 ( .A1(u5_mult_87_n387), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__30_) );
  NOR2_X1 u5_mult_87_U3003 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__31_) );
  NOR2_X1 u5_mult_87_U3002 ( .A1(u5_mult_87_n383), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__32_) );
  NOR2_X1 u5_mult_87_U3001 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__33_) );
  NOR2_X1 u5_mult_87_U3000 ( .A1(u5_mult_87_n379), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__34_) );
  NOR2_X1 u5_mult_87_U2999 ( .A1(u5_mult_87_n377), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__35_) );
  NOR2_X1 u5_mult_87_U2998 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__36_) );
  NOR2_X1 u5_mult_87_U2997 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__37_) );
  NOR2_X1 u5_mult_87_U2996 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__38_) );
  NOR2_X1 u5_mult_87_U2995 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__39_) );
  NOR2_X1 u5_mult_87_U2994 ( .A1(u5_mult_87_n442), .A2(u5_mult_87_n472), .ZN(
        u5_mult_87_ab_14__3_) );
  NOR2_X1 u5_mult_87_U2993 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n472), .ZN(
        u5_mult_87_ab_14__40_) );
  NOR2_X1 u5_mult_87_U2992 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__41_) );
  NOR2_X1 u5_mult_87_U2991 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n472), .ZN(
        u5_mult_87_ab_14__42_) );
  NOR2_X1 u5_mult_87_U2990 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n472), .ZN(
        u5_mult_87_ab_14__43_) );
  NOR2_X1 u5_mult_87_U2989 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n472), .ZN(
        u5_mult_87_ab_14__44_) );
  NOR2_X1 u5_mult_87_U2988 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n472), .ZN(
        u5_mult_87_ab_14__45_) );
  NOR2_X1 u5_mult_87_U2987 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n472), .ZN(
        u5_mult_87_ab_14__46_) );
  NOR2_X1 u5_mult_87_U2986 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n472), .ZN(
        u5_mult_87_ab_14__47_) );
  NOR2_X1 u5_mult_87_U2985 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n472), .ZN(
        u5_mult_87_ab_14__48_) );
  NOR2_X1 u5_mult_87_U2984 ( .A1(u5_mult_87_n348), .A2(u5_mult_87_n472), .ZN(
        u5_mult_87_ab_14__49_) );
  NOR2_X1 u5_mult_87_U2983 ( .A1(u5_mult_87_n440), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__4_) );
  NOR2_X1 u5_mult_87_U2982 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__50_) );
  NOR2_X1 u5_mult_87_U2981 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__51_) );
  NOR2_X1 u5_mult_87_U2980 ( .A1(u5_mult_87_n342), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__52_) );
  NOR2_X1 u5_mult_87_U2979 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__5_) );
  NOR2_X1 u5_mult_87_U2978 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__6_) );
  NOR2_X1 u5_mult_87_U2977 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__7_) );
  NOR2_X1 u5_mult_87_U2976 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__8_) );
  NOR2_X1 u5_mult_87_U2975 ( .A1(u5_mult_87_n430), .A2(u5_mult_87_n303), .ZN(
        u5_mult_87_ab_14__9_) );
  NOR2_X1 u5_mult_87_U2974 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__0_) );
  NOR2_X1 u5_mult_87_U2973 ( .A1(u5_mult_87_n428), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__10_) );
  NOR2_X1 u5_mult_87_U2972 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__11_) );
  NOR2_X1 u5_mult_87_U2971 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__12_) );
  NOR2_X1 u5_mult_87_U2970 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__13_) );
  NOR2_X1 u5_mult_87_U2969 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__14_) );
  NOR2_X1 u5_mult_87_U2968 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__15_) );
  NOR2_X1 u5_mult_87_U2967 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__16_) );
  NOR2_X1 u5_mult_87_U2966 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__17_) );
  NOR2_X1 u5_mult_87_U2965 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__18_) );
  NOR2_X1 u5_mult_87_U2964 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__19_) );
  NOR2_X1 u5_mult_87_U2963 ( .A1(u5_mult_87_n446), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__1_) );
  NOR2_X1 u5_mult_87_U2962 ( .A1(u5_mult_87_n407), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__20_) );
  NOR2_X1 u5_mult_87_U2961 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__21_) );
  NOR2_X1 u5_mult_87_U2960 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__22_) );
  NOR2_X1 u5_mult_87_U2959 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__23_) );
  NOR2_X1 u5_mult_87_U2958 ( .A1(u5_mult_87_n399), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__24_) );
  NOR2_X1 u5_mult_87_U2957 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__25_) );
  NOR2_X1 u5_mult_87_U2956 ( .A1(u5_mult_87_n395), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__26_) );
  NOR2_X1 u5_mult_87_U2955 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__27_) );
  NOR2_X1 u5_mult_87_U2954 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__28_) );
  NOR2_X1 u5_mult_87_U2953 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__29_) );
  NOR2_X1 u5_mult_87_U2952 ( .A1(u5_mult_87_n444), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__2_) );
  NOR2_X1 u5_mult_87_U2951 ( .A1(u5_mult_87_n387), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__30_) );
  NOR2_X1 u5_mult_87_U2950 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__31_) );
  NOR2_X1 u5_mult_87_U2949 ( .A1(u5_mult_87_n383), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__32_) );
  NOR2_X1 u5_mult_87_U2948 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__33_) );
  NOR2_X1 u5_mult_87_U2947 ( .A1(u5_mult_87_n379), .A2(u5_mult_87_n302), .ZN(
        u5_mult_87_ab_15__34_) );
  NOR2_X1 u5_mult_87_U2946 ( .A1(u5_mult_87_n377), .A2(u5_mult_87_n302), .ZN(
        u5_mult_87_ab_15__35_) );
  NOR2_X1 u5_mult_87_U2945 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n302), .ZN(
        u5_mult_87_ab_15__36_) );
  NOR2_X1 u5_mult_87_U2944 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n302), .ZN(
        u5_mult_87_ab_15__37_) );
  NOR2_X1 u5_mult_87_U2943 ( .A1(u5_mult_87_n372), .A2(u5_mult_87_n302), .ZN(
        u5_mult_87_ab_15__38_) );
  NOR2_X1 u5_mult_87_U2942 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n302), .ZN(
        u5_mult_87_ab_15__39_) );
  NOR2_X1 u5_mult_87_U2941 ( .A1(u5_mult_87_n442), .A2(u5_mult_87_n302), .ZN(
        u5_mult_87_ab_15__3_) );
  NOR2_X1 u5_mult_87_U2940 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n302), .ZN(
        u5_mult_87_ab_15__40_) );
  NOR2_X1 u5_mult_87_U2939 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n302), .ZN(
        u5_mult_87_ab_15__41_) );
  NOR2_X1 u5_mult_87_U2938 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n302), .ZN(
        u5_mult_87_ab_15__42_) );
  NOR2_X1 u5_mult_87_U2937 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n302), .ZN(
        u5_mult_87_ab_15__43_) );
  NOR2_X1 u5_mult_87_U2936 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n302), .ZN(
        u5_mult_87_ab_15__44_) );
  NOR2_X1 u5_mult_87_U2935 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n302), .ZN(
        u5_mult_87_ab_15__45_) );
  NOR2_X1 u5_mult_87_U2934 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n302), .ZN(
        u5_mult_87_ab_15__46_) );
  NOR2_X1 u5_mult_87_U2933 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n302), .ZN(
        u5_mult_87_ab_15__47_) );
  NOR2_X1 u5_mult_87_U2932 ( .A1(u5_mult_87_n350), .A2(u5_mult_87_n302), .ZN(
        u5_mult_87_ab_15__48_) );
  NOR2_X1 u5_mult_87_U2931 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n302), .ZN(
        u5_mult_87_ab_15__49_) );
  NOR2_X1 u5_mult_87_U2930 ( .A1(u5_mult_87_n440), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__4_) );
  NOR2_X1 u5_mult_87_U2929 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__50_) );
  NOR2_X1 u5_mult_87_U2928 ( .A1(u5_mult_87_n345), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__51_) );
  NOR2_X1 u5_mult_87_U2927 ( .A1(u5_mult_87_n342), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__52_) );
  NOR2_X1 u5_mult_87_U2926 ( .A1(u5_mult_87_n439), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__5_) );
  NOR2_X1 u5_mult_87_U2925 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__6_) );
  NOR2_X1 u5_mult_87_U2924 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__7_) );
  NOR2_X1 u5_mult_87_U2923 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__8_) );
  NOR2_X1 u5_mult_87_U2922 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n301), .ZN(
        u5_mult_87_ab_15__9_) );
  NOR2_X1 u5_mult_87_U2921 ( .A1(u5_mult_87_n450), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__0_) );
  NOR2_X1 u5_mult_87_U2920 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__10_) );
  NOR2_X1 u5_mult_87_U2919 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__11_) );
  NOR2_X1 u5_mult_87_U2918 ( .A1(u5_mult_87_n481), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__12_) );
  NOR2_X1 u5_mult_87_U2917 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__13_) );
  NOR2_X1 u5_mult_87_U2916 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__14_) );
  NOR2_X1 u5_mult_87_U2915 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__15_) );
  NOR2_X1 u5_mult_87_U2914 ( .A1(u5_mult_87_n480), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__16_) );
  NOR2_X1 u5_mult_87_U2913 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__17_) );
  NOR2_X1 u5_mult_87_U2912 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__18_) );
  NOR2_X1 u5_mult_87_U2911 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__19_) );
  NOR2_X1 u5_mult_87_U2910 ( .A1(u5_mult_87_n446), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__1_) );
  NOR2_X1 u5_mult_87_U2909 ( .A1(u5_mult_87_n407), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__20_) );
  NOR2_X1 u5_mult_87_U2908 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__21_) );
  NOR2_X1 u5_mult_87_U2907 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__22_) );
  NOR2_X1 u5_mult_87_U2906 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__23_) );
  NOR2_X1 u5_mult_87_U2905 ( .A1(u5_mult_87_n399), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__24_) );
  NOR2_X1 u5_mult_87_U2904 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__25_) );
  NOR2_X1 u5_mult_87_U2903 ( .A1(u5_mult_87_n395), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__26_) );
  NOR2_X1 u5_mult_87_U2902 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__27_) );
  NOR2_X1 u5_mult_87_U2901 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__28_) );
  NOR2_X1 u5_mult_87_U2900 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__29_) );
  NOR2_X1 u5_mult_87_U2899 ( .A1(u5_mult_87_n444), .A2(u5_mult_87_n471), .ZN(
        u5_mult_87_ab_16__2_) );
  NOR2_X1 u5_mult_87_U2898 ( .A1(u5_mult_87_n387), .A2(u5_mult_87_n471), .ZN(
        u5_mult_87_ab_16__30_) );
  NOR2_X1 u5_mult_87_U2897 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n471), .ZN(
        u5_mult_87_ab_16__31_) );
  NOR2_X1 u5_mult_87_U2896 ( .A1(u5_mult_87_n383), .A2(u5_mult_87_n471), .ZN(
        u5_mult_87_ab_16__32_) );
  NOR2_X1 u5_mult_87_U2895 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n471), .ZN(
        u5_mult_87_ab_16__33_) );
  NOR2_X1 u5_mult_87_U2894 ( .A1(u5_mult_87_n379), .A2(u5_mult_87_n471), .ZN(
        u5_mult_87_ab_16__34_) );
  NOR2_X1 u5_mult_87_U2893 ( .A1(u5_mult_87_n377), .A2(u5_mult_87_n300), .ZN(
        u5_mult_87_ab_16__35_) );
  NOR2_X1 u5_mult_87_U2892 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n471), .ZN(
        u5_mult_87_ab_16__36_) );
  NOR2_X1 u5_mult_87_U2891 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n300), .ZN(
        u5_mult_87_ab_16__37_) );
  NOR2_X1 u5_mult_87_U2890 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n471), .ZN(
        u5_mult_87_ab_16__38_) );
  NOR2_X1 u5_mult_87_U2889 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n471), .ZN(
        u5_mult_87_ab_16__39_) );
  NOR2_X1 u5_mult_87_U2888 ( .A1(u5_mult_87_n442), .A2(u5_mult_87_n300), .ZN(
        u5_mult_87_ab_16__3_) );
  NOR2_X1 u5_mult_87_U2887 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n300), .ZN(
        u5_mult_87_ab_16__40_) );
  NOR2_X1 u5_mult_87_U2886 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n300), .ZN(
        u5_mult_87_ab_16__41_) );
  NOR2_X1 u5_mult_87_U2885 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n300), .ZN(
        u5_mult_87_ab_16__42_) );
  NOR2_X1 u5_mult_87_U2884 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n300), .ZN(
        u5_mult_87_ab_16__43_) );
  NOR2_X1 u5_mult_87_U2883 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n300), .ZN(
        u5_mult_87_ab_16__44_) );
  NOR2_X1 u5_mult_87_U2882 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n300), .ZN(
        u5_mult_87_ab_16__45_) );
  NOR2_X1 u5_mult_87_U2881 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n300), .ZN(
        u5_mult_87_ab_16__46_) );
  NOR2_X1 u5_mult_87_U2880 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n300), .ZN(
        u5_mult_87_ab_16__47_) );
  NOR2_X1 u5_mult_87_U2879 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n300), .ZN(
        u5_mult_87_ab_16__48_) );
  NOR2_X1 u5_mult_87_U2878 ( .A1(u5_mult_87_n348), .A2(u5_mult_87_n300), .ZN(
        u5_mult_87_ab_16__49_) );
  NOR2_X1 u5_mult_87_U2877 ( .A1(u5_mult_87_n440), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__4_) );
  NOR2_X1 u5_mult_87_U2876 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__50_) );
  NOR2_X1 u5_mult_87_U2875 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__51_) );
  NOR2_X1 u5_mult_87_U2874 ( .A1(u5_mult_87_n342), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__52_) );
  NOR2_X1 u5_mult_87_U2873 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__5_) );
  NOR2_X1 u5_mult_87_U2872 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__6_) );
  NOR2_X1 u5_mult_87_U2871 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__7_) );
  NOR2_X1 u5_mult_87_U2870 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__8_) );
  NOR2_X1 u5_mult_87_U2869 ( .A1(u5_mult_87_n430), .A2(u5_mult_87_n299), .ZN(
        u5_mult_87_ab_16__9_) );
  NOR2_X1 u5_mult_87_U2868 ( .A1(u5_mult_87_n450), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__0_) );
  NOR2_X1 u5_mult_87_U2867 ( .A1(u5_mult_87_n428), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__10_) );
  NOR2_X1 u5_mult_87_U2866 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__11_) );
  NOR2_X1 u5_mult_87_U2865 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__12_) );
  NOR2_X1 u5_mult_87_U2864 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__13_) );
  NOR2_X1 u5_mult_87_U2863 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__14_) );
  NOR2_X1 u5_mult_87_U2862 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__15_) );
  NOR2_X1 u5_mult_87_U2861 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__16_) );
  NOR2_X1 u5_mult_87_U2860 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__17_) );
  NOR2_X1 u5_mult_87_U2859 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__18_) );
  NOR2_X1 u5_mult_87_U2858 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__19_) );
  NOR2_X1 u5_mult_87_U2857 ( .A1(u5_mult_87_n446), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__1_) );
  NOR2_X1 u5_mult_87_U2856 ( .A1(u5_mult_87_n407), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__20_) );
  NOR2_X1 u5_mult_87_U2855 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__21_) );
  NOR2_X1 u5_mult_87_U2854 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__22_) );
  NOR2_X1 u5_mult_87_U2853 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__23_) );
  NOR2_X1 u5_mult_87_U2852 ( .A1(u5_mult_87_n399), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__24_) );
  NOR2_X1 u5_mult_87_U2851 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__25_) );
  NOR2_X1 u5_mult_87_U2850 ( .A1(u5_mult_87_n395), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__26_) );
  NOR2_X1 u5_mult_87_U2849 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__27_) );
  NOR2_X1 u5_mult_87_U2848 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__28_) );
  NOR2_X1 u5_mult_87_U2847 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__29_) );
  NOR2_X1 u5_mult_87_U2846 ( .A1(u5_mult_87_n444), .A2(u5_mult_87_n470), .ZN(
        u5_mult_87_ab_17__2_) );
  NOR2_X1 u5_mult_87_U2845 ( .A1(u5_mult_87_n387), .A2(u5_mult_87_n470), .ZN(
        u5_mult_87_ab_17__30_) );
  NOR2_X1 u5_mult_87_U2844 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n470), .ZN(
        u5_mult_87_ab_17__31_) );
  NOR2_X1 u5_mult_87_U2843 ( .A1(u5_mult_87_n383), .A2(u5_mult_87_n470), .ZN(
        u5_mult_87_ab_17__32_) );
  NOR2_X1 u5_mult_87_U2842 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n470), .ZN(
        u5_mult_87_ab_17__33_) );
  NOR2_X1 u5_mult_87_U2841 ( .A1(u5_mult_87_n379), .A2(u5_mult_87_n470), .ZN(
        u5_mult_87_ab_17__34_) );
  NOR2_X1 u5_mult_87_U2840 ( .A1(u5_mult_87_n377), .A2(u5_mult_87_n298), .ZN(
        u5_mult_87_ab_17__35_) );
  NOR2_X1 u5_mult_87_U2839 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n470), .ZN(
        u5_mult_87_ab_17__36_) );
  NOR2_X1 u5_mult_87_U2838 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n298), .ZN(
        u5_mult_87_ab_17__37_) );
  NOR2_X1 u5_mult_87_U2837 ( .A1(u5_mult_87_n372), .A2(u5_mult_87_n470), .ZN(
        u5_mult_87_ab_17__38_) );
  NOR2_X1 u5_mult_87_U2836 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n470), .ZN(
        u5_mult_87_ab_17__39_) );
  NOR2_X1 u5_mult_87_U2835 ( .A1(u5_mult_87_n442), .A2(u5_mult_87_n298), .ZN(
        u5_mult_87_ab_17__3_) );
  NOR2_X1 u5_mult_87_U2834 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n298), .ZN(
        u5_mult_87_ab_17__40_) );
  NOR2_X1 u5_mult_87_U2833 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n298), .ZN(
        u5_mult_87_ab_17__41_) );
  NOR2_X1 u5_mult_87_U2832 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n298), .ZN(
        u5_mult_87_ab_17__42_) );
  NOR2_X1 u5_mult_87_U2831 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n298), .ZN(
        u5_mult_87_ab_17__43_) );
  NOR2_X1 u5_mult_87_U2830 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n298), .ZN(
        u5_mult_87_ab_17__44_) );
  NOR2_X1 u5_mult_87_U2829 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n298), .ZN(
        u5_mult_87_ab_17__45_) );
  NOR2_X1 u5_mult_87_U2828 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n298), .ZN(
        u5_mult_87_ab_17__46_) );
  NOR2_X1 u5_mult_87_U2827 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n298), .ZN(
        u5_mult_87_ab_17__47_) );
  NOR2_X1 u5_mult_87_U2826 ( .A1(u5_mult_87_n350), .A2(u5_mult_87_n298), .ZN(
        u5_mult_87_ab_17__48_) );
  NOR2_X1 u5_mult_87_U2825 ( .A1(u5_mult_87_n348), .A2(u5_mult_87_n298), .ZN(
        u5_mult_87_ab_17__49_) );
  NOR2_X1 u5_mult_87_U2824 ( .A1(u5_mult_87_n440), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__4_) );
  NOR2_X1 u5_mult_87_U2823 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__50_) );
  NOR2_X1 u5_mult_87_U2822 ( .A1(u5_mult_87_n345), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__51_) );
  NOR2_X1 u5_mult_87_U2821 ( .A1(u5_mult_87_n342), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__52_) );
  NOR2_X1 u5_mult_87_U2820 ( .A1(u5_mult_87_n439), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__5_) );
  NOR2_X1 u5_mult_87_U2819 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__6_) );
  NOR2_X1 u5_mult_87_U2818 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__7_) );
  NOR2_X1 u5_mult_87_U2817 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__8_) );
  NOR2_X1 u5_mult_87_U2816 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n297), .ZN(
        u5_mult_87_ab_17__9_) );
  NOR2_X1 u5_mult_87_U2815 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__0_) );
  NOR2_X1 u5_mult_87_U2814 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__10_) );
  NOR2_X1 u5_mult_87_U2813 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__11_) );
  NOR2_X1 u5_mult_87_U2812 ( .A1(u5_mult_87_n481), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__12_) );
  NOR2_X1 u5_mult_87_U2811 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__13_) );
  NOR2_X1 u5_mult_87_U2810 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__14_) );
  NOR2_X1 u5_mult_87_U2809 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__15_) );
  NOR2_X1 u5_mult_87_U2808 ( .A1(u5_mult_87_n480), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__16_) );
  NOR2_X1 u5_mult_87_U2807 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__17_) );
  NOR2_X1 u5_mult_87_U2806 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__18_) );
  NOR2_X1 u5_mult_87_U2805 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__19_) );
  NOR2_X1 u5_mult_87_U2804 ( .A1(u5_mult_87_n446), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__1_) );
  NOR2_X1 u5_mult_87_U2803 ( .A1(u5_mult_87_n407), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__20_) );
  NOR2_X1 u5_mult_87_U2802 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__21_) );
  NOR2_X1 u5_mult_87_U2801 ( .A1(u5_mult_87_n404), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__22_) );
  NOR2_X1 u5_mult_87_U2800 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__23_) );
  NOR2_X1 u5_mult_87_U2799 ( .A1(u5_mult_87_n399), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__24_) );
  NOR2_X1 u5_mult_87_U2798 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__25_) );
  NOR2_X1 u5_mult_87_U2797 ( .A1(u5_mult_87_n395), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__26_) );
  NOR2_X1 u5_mult_87_U2796 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__27_) );
  NOR2_X1 u5_mult_87_U2795 ( .A1(u5_mult_87_n392), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__28_) );
  NOR2_X1 u5_mult_87_U2794 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__29_) );
  NOR2_X1 u5_mult_87_U2793 ( .A1(u5_mult_87_n444), .A2(u5_mult_87_n469), .ZN(
        u5_mult_87_ab_18__2_) );
  NOR2_X1 u5_mult_87_U2792 ( .A1(u5_mult_87_n387), .A2(u5_mult_87_n469), .ZN(
        u5_mult_87_ab_18__30_) );
  NOR2_X1 u5_mult_87_U2791 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n469), .ZN(
        u5_mult_87_ab_18__31_) );
  NOR2_X1 u5_mult_87_U2790 ( .A1(u5_mult_87_n383), .A2(u5_mult_87_n469), .ZN(
        u5_mult_87_ab_18__32_) );
  NOR2_X1 u5_mult_87_U2789 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n296), .ZN(
        u5_mult_87_ab_18__33_) );
  NOR2_X1 u5_mult_87_U2788 ( .A1(u5_mult_87_n379), .A2(u5_mult_87_n296), .ZN(
        u5_mult_87_ab_18__34_) );
  NOR2_X1 u5_mult_87_U2787 ( .A1(u5_mult_87_n377), .A2(u5_mult_87_n296), .ZN(
        u5_mult_87_ab_18__35_) );
  NOR2_X1 u5_mult_87_U2786 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n296), .ZN(
        u5_mult_87_ab_18__36_) );
  NOR2_X1 u5_mult_87_U2785 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n296), .ZN(
        u5_mult_87_ab_18__37_) );
  NOR2_X1 u5_mult_87_U2784 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n296), .ZN(
        u5_mult_87_ab_18__38_) );
  NOR2_X1 u5_mult_87_U2783 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n469), .ZN(
        u5_mult_87_ab_18__39_) );
  NOR2_X1 u5_mult_87_U2782 ( .A1(u5_mult_87_n442), .A2(u5_mult_87_n296), .ZN(
        u5_mult_87_ab_18__3_) );
  NOR2_X1 u5_mult_87_U2781 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n296), .ZN(
        u5_mult_87_ab_18__40_) );
  NOR2_X1 u5_mult_87_U2780 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n296), .ZN(
        u5_mult_87_ab_18__41_) );
  NOR2_X1 u5_mult_87_U2779 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n296), .ZN(
        u5_mult_87_ab_18__42_) );
  NOR2_X1 u5_mult_87_U2778 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n296), .ZN(
        u5_mult_87_ab_18__43_) );
  NOR2_X1 u5_mult_87_U2777 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n296), .ZN(
        u5_mult_87_ab_18__44_) );
  NOR2_X1 u5_mult_87_U2776 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n296), .ZN(
        u5_mult_87_ab_18__45_) );
  NOR2_X1 u5_mult_87_U2775 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n296), .ZN(
        u5_mult_87_ab_18__46_) );
  NOR2_X1 u5_mult_87_U2774 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n296), .ZN(
        u5_mult_87_ab_18__47_) );
  NOR2_X1 u5_mult_87_U2773 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n296), .ZN(
        u5_mult_87_ab_18__48_) );
  NOR2_X1 u5_mult_87_U2772 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n296), .ZN(
        u5_mult_87_ab_18__49_) );
  NOR2_X1 u5_mult_87_U2771 ( .A1(u5_mult_87_n440), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__4_) );
  NOR2_X1 u5_mult_87_U2770 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__50_) );
  NOR2_X1 u5_mult_87_U2769 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__51_) );
  NOR2_X1 u5_mult_87_U2768 ( .A1(u5_mult_87_n342), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__52_) );
  NOR2_X1 u5_mult_87_U2767 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__5_) );
  NOR2_X1 u5_mult_87_U2766 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__6_) );
  NOR2_X1 u5_mult_87_U2765 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__7_) );
  NOR2_X1 u5_mult_87_U2764 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__8_) );
  NOR2_X1 u5_mult_87_U2763 ( .A1(u5_mult_87_n430), .A2(u5_mult_87_n295), .ZN(
        u5_mult_87_ab_18__9_) );
  NOR2_X1 u5_mult_87_U2762 ( .A1(u5_mult_87_n450), .A2(u5_mult_87_n293), .ZN(
        u5_mult_87_ab_19__0_) );
  NOR2_X1 u5_mult_87_U2761 ( .A1(u5_mult_87_n428), .A2(u5_mult_87_n293), .ZN(
        u5_mult_87_ab_19__10_) );
  NOR2_X1 u5_mult_87_U2760 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n293), .ZN(
        u5_mult_87_ab_19__11_) );
  NOR2_X1 u5_mult_87_U2759 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n293), .ZN(
        u5_mult_87_ab_19__12_) );
  NOR2_X1 u5_mult_87_U2758 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n293), .ZN(
        u5_mult_87_ab_19__13_) );
  NOR2_X1 u5_mult_87_U2757 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n293), .ZN(
        u5_mult_87_ab_19__14_) );
  NOR2_X1 u5_mult_87_U2756 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n293), .ZN(
        u5_mult_87_ab_19__15_) );
  NOR2_X1 u5_mult_87_U2755 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n293), .ZN(
        u5_mult_87_ab_19__16_) );
  NOR2_X1 u5_mult_87_U2754 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n293), .ZN(
        u5_mult_87_ab_19__17_) );
  NOR2_X1 u5_mult_87_U2753 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n293), .ZN(
        u5_mult_87_ab_19__18_) );
  NOR2_X1 u5_mult_87_U2752 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n293), .ZN(
        u5_mult_87_ab_19__19_) );
  NOR2_X1 u5_mult_87_U2751 ( .A1(u5_mult_87_n446), .A2(u5_mult_87_n292), .ZN(
        u5_mult_87_ab_19__1_) );
  NOR2_X1 u5_mult_87_U2750 ( .A1(u5_mult_87_n407), .A2(u5_mult_87_n292), .ZN(
        u5_mult_87_ab_19__20_) );
  NOR2_X1 u5_mult_87_U2749 ( .A1(u5_mult_87_n406), .A2(u5_mult_87_n292), .ZN(
        u5_mult_87_ab_19__21_) );
  NOR2_X1 u5_mult_87_U2748 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n292), .ZN(
        u5_mult_87_ab_19__22_) );
  NOR2_X1 u5_mult_87_U2747 ( .A1(u5_mult_87_n402), .A2(u5_mult_87_n292), .ZN(
        u5_mult_87_ab_19__23_) );
  NOR2_X1 u5_mult_87_U2746 ( .A1(u5_mult_87_n399), .A2(u5_mult_87_n292), .ZN(
        u5_mult_87_ab_19__24_) );
  NOR2_X1 u5_mult_87_U2745 ( .A1(u5_mult_87_n398), .A2(u5_mult_87_n292), .ZN(
        u5_mult_87_ab_19__25_) );
  NOR2_X1 u5_mult_87_U2744 ( .A1(u5_mult_87_n395), .A2(u5_mult_87_n292), .ZN(
        u5_mult_87_ab_19__26_) );
  NOR2_X1 u5_mult_87_U2743 ( .A1(u5_mult_87_n394), .A2(u5_mult_87_n292), .ZN(
        u5_mult_87_ab_19__27_) );
  NOR2_X1 u5_mult_87_U2742 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n292), .ZN(
        u5_mult_87_ab_19__28_) );
  NOR2_X1 u5_mult_87_U2741 ( .A1(u5_mult_87_n390), .A2(u5_mult_87_n292), .ZN(
        u5_mult_87_ab_19__29_) );
  NOR2_X1 u5_mult_87_U2740 ( .A1(u5_mult_87_n444), .A2(u5_mult_87_n293), .ZN(
        u5_mult_87_ab_19__2_) );
  NOR2_X1 u5_mult_87_U2739 ( .A1(u5_mult_87_n387), .A2(u5_mult_87_n293), .ZN(
        u5_mult_87_ab_19__30_) );
  NOR2_X1 u5_mult_87_U2738 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n292), .ZN(
        u5_mult_87_ab_19__31_) );
  NOR2_X1 u5_mult_87_U2737 ( .A1(u5_mult_87_n383), .A2(u5_mult_87_n292), .ZN(
        u5_mult_87_ab_19__32_) );
  NOR2_X1 u5_mult_87_U2736 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n292), .ZN(
        u5_mult_87_ab_19__33_) );
  NOR2_X1 u5_mult_87_U2735 ( .A1(u5_mult_87_n379), .A2(u5_mult_87_n292), .ZN(
        u5_mult_87_ab_19__34_) );
  NOR2_X1 u5_mult_87_U2734 ( .A1(u5_mult_87_n377), .A2(u5_mult_87_n294), .ZN(
        u5_mult_87_ab_19__35_) );
  NOR2_X1 u5_mult_87_U2733 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n294), .ZN(
        u5_mult_87_ab_19__36_) );
  NOR2_X1 u5_mult_87_U2732 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n292), .ZN(
        u5_mult_87_ab_19__37_) );
  NOR2_X1 u5_mult_87_U2731 ( .A1(u5_mult_87_n372), .A2(u5_mult_87_n292), .ZN(
        u5_mult_87_ab_19__38_) );
  NOR2_X1 u5_mult_87_U2730 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n292), .ZN(
        u5_mult_87_ab_19__39_) );
  NOR2_X1 u5_mult_87_U2729 ( .A1(u5_mult_87_n442), .A2(u5_mult_87_n294), .ZN(
        u5_mult_87_ab_19__3_) );
  NOR2_X1 u5_mult_87_U2728 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n294), .ZN(
        u5_mult_87_ab_19__40_) );
  NOR2_X1 u5_mult_87_U2727 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n292), .ZN(
        u5_mult_87_ab_19__41_) );
  NOR2_X1 u5_mult_87_U2726 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n294), .ZN(
        u5_mult_87_ab_19__42_) );
  NOR2_X1 u5_mult_87_U2725 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n294), .ZN(
        u5_mult_87_ab_19__43_) );
  NOR2_X1 u5_mult_87_U2724 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n294), .ZN(
        u5_mult_87_ab_19__44_) );
  NOR2_X1 u5_mult_87_U2723 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n292), .ZN(
        u5_mult_87_ab_19__45_) );
  NOR2_X1 u5_mult_87_U2722 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n292), .ZN(
        u5_mult_87_ab_19__46_) );
  NOR2_X1 u5_mult_87_U2721 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n294), .ZN(
        u5_mult_87_ab_19__47_) );
  NOR2_X1 u5_mult_87_U2720 ( .A1(u5_mult_87_n350), .A2(u5_mult_87_n292), .ZN(
        u5_mult_87_ab_19__48_) );
  NOR2_X1 u5_mult_87_U2719 ( .A1(u5_mult_87_n348), .A2(u5_mult_87_n294), .ZN(
        u5_mult_87_ab_19__49_) );
  NOR2_X1 u5_mult_87_U2718 ( .A1(u5_mult_87_n440), .A2(u5_mult_87_n293), .ZN(
        u5_mult_87_ab_19__4_) );
  NOR2_X1 u5_mult_87_U2717 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n293), .ZN(
        u5_mult_87_ab_19__50_) );
  NOR2_X1 u5_mult_87_U2716 ( .A1(u5_mult_87_n345), .A2(u5_mult_87_n293), .ZN(
        u5_mult_87_ab_19__51_) );
  NOR2_X1 u5_mult_87_U2715 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n293), .ZN(
        u5_mult_87_ab_19__52_) );
  NOR2_X1 u5_mult_87_U2714 ( .A1(u5_mult_87_n439), .A2(u5_mult_87_n293), .ZN(
        u5_mult_87_ab_19__5_) );
  NOR2_X1 u5_mult_87_U2713 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n293), .ZN(
        u5_mult_87_ab_19__6_) );
  NOR2_X1 u5_mult_87_U2712 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n293), .ZN(
        u5_mult_87_ab_19__7_) );
  NOR2_X1 u5_mult_87_U2711 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n293), .ZN(
        u5_mult_87_ab_19__8_) );
  NOR2_X1 u5_mult_87_U2710 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n293), .ZN(
        u5_mult_87_ab_19__9_) );
  NOR2_X1 u5_mult_87_U2709 ( .A1(u5_mult_87_n450), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__0_) );
  NOR2_X1 u5_mult_87_U2708 ( .A1(u5_mult_87_n428), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__10_) );
  NOR2_X1 u5_mult_87_U2707 ( .A1(u5_mult_87_n425), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__11_) );
  NOR2_X1 u5_mult_87_U2706 ( .A1(u5_mult_87_n481), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__12_) );
  NOR2_X1 u5_mult_87_U2705 ( .A1(u5_mult_87_n422), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__13_) );
  NOR2_X1 u5_mult_87_U2704 ( .A1(u5_mult_87_n421), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__14_) );
  NOR2_X1 u5_mult_87_U2703 ( .A1(u5_mult_87_n416), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__15_) );
  NOR2_X1 u5_mult_87_U2702 ( .A1(u5_mult_87_n480), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__16_) );
  NOR2_X1 u5_mult_87_U2701 ( .A1(u5_mult_87_n413), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__17_) );
  NOR2_X1 u5_mult_87_U2700 ( .A1(u5_mult_87_n411), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__18_) );
  NOR2_X1 u5_mult_87_U2699 ( .A1(u5_mult_87_n409), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__19_) );
  NOR2_X1 u5_mult_87_U2698 ( .A1(u5_mult_87_n482), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__1_) );
  NOR2_X1 u5_mult_87_U2697 ( .A1(u5_mult_87_n407), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__20_) );
  NOR2_X1 u5_mult_87_U2696 ( .A1(u5_mult_87_n406), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__21_) );
  NOR2_X1 u5_mult_87_U2695 ( .A1(u5_mult_87_n404), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__22_) );
  NOR2_X1 u5_mult_87_U2694 ( .A1(u5_mult_87_n402), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__23_) );
  NOR2_X1 u5_mult_87_U2693 ( .A1(u5_mult_87_n399), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__24_) );
  NOR2_X1 u5_mult_87_U2692 ( .A1(u5_mult_87_n398), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__25_) );
  NOR2_X1 u5_mult_87_U2691 ( .A1(u5_mult_87_n395), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__26_) );
  NOR2_X1 u5_mult_87_U2690 ( .A1(u5_mult_87_n394), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__27_) );
  NOR2_X1 u5_mult_87_U2689 ( .A1(u5_mult_87_n392), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__28_) );
  NOR2_X1 u5_mult_87_U2688 ( .A1(u5_mult_87_n390), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__29_) );
  NOR2_X1 u5_mult_87_U2687 ( .A1(u5_mult_87_n444), .A2(u5_mult_87_n337), .ZN(
        u5_mult_87_ab_1__2_) );
  NOR2_X1 u5_mult_87_U2686 ( .A1(u5_mult_87_n387), .A2(u5_mult_87_n337), .ZN(
        u5_mult_87_ab_1__30_) );
  NOR2_X1 u5_mult_87_U2685 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n337), .ZN(
        u5_mult_87_ab_1__31_) );
  NOR2_X1 u5_mult_87_U2684 ( .A1(u5_mult_87_n383), .A2(u5_mult_87_n337), .ZN(
        u5_mult_87_ab_1__32_) );
  NOR2_X1 u5_mult_87_U2683 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n337), .ZN(
        u5_mult_87_ab_1__33_) );
  NOR2_X1 u5_mult_87_U2682 ( .A1(u5_mult_87_n379), .A2(u5_mult_87_n337), .ZN(
        u5_mult_87_ab_1__34_) );
  NOR2_X1 u5_mult_87_U2681 ( .A1(u5_mult_87_n377), .A2(u5_mult_87_n337), .ZN(
        u5_mult_87_ab_1__35_) );
  NOR2_X1 u5_mult_87_U2680 ( .A1(u5_mult_87_n376), .A2(u5_mult_87_n337), .ZN(
        u5_mult_87_ab_1__36_) );
  NOR2_X1 u5_mult_87_U2679 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n337), .ZN(
        u5_mult_87_ab_1__37_) );
  NOR2_X1 u5_mult_87_U2678 ( .A1(u5_mult_87_n372), .A2(u5_mult_87_n337), .ZN(
        u5_mult_87_ab_1__38_) );
  NOR2_X1 u5_mult_87_U2677 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n337), .ZN(
        u5_mult_87_ab_1__39_) );
  NOR2_X1 u5_mult_87_U2676 ( .A1(u5_mult_87_n442), .A2(u5_mult_87_n338), .ZN(
        u5_mult_87_ab_1__3_) );
  NOR2_X1 u5_mult_87_U2675 ( .A1(u5_mult_87_n367), .A2(u5_mult_87_n338), .ZN(
        u5_mult_87_ab_1__40_) );
  NOR2_X1 u5_mult_87_U2674 ( .A1(u5_mult_87_n365), .A2(u5_mult_87_n338), .ZN(
        u5_mult_87_ab_1__41_) );
  NOR2_X1 u5_mult_87_U2673 ( .A1(u5_mult_87_n363), .A2(u5_mult_87_n338), .ZN(
        u5_mult_87_ab_1__42_) );
  NOR2_X1 u5_mult_87_U2672 ( .A1(u5_mult_87_n360), .A2(u5_mult_87_n338), .ZN(
        u5_mult_87_ab_1__43_) );
  NOR2_X1 u5_mult_87_U2671 ( .A1(u5_mult_87_n358), .A2(u5_mult_87_n338), .ZN(
        u5_mult_87_ab_1__44_) );
  NOR2_X1 u5_mult_87_U2670 ( .A1(u5_mult_87_n356), .A2(u5_mult_87_n338), .ZN(
        u5_mult_87_ab_1__45_) );
  NOR2_X1 u5_mult_87_U2669 ( .A1(u5_mult_87_n354), .A2(u5_mult_87_n338), .ZN(
        u5_mult_87_ab_1__46_) );
  NOR2_X1 u5_mult_87_U2668 ( .A1(u5_mult_87_n351), .A2(u5_mult_87_n338), .ZN(
        u5_mult_87_ab_1__47_) );
  NOR2_X1 u5_mult_87_U2667 ( .A1(u5_mult_87_n350), .A2(u5_mult_87_n338), .ZN(
        u5_mult_87_ab_1__48_) );
  NOR2_X1 u5_mult_87_U2666 ( .A1(u5_mult_87_n348), .A2(u5_mult_87_n338), .ZN(
        u5_mult_87_ab_1__49_) );
  NOR2_X1 u5_mult_87_U2665 ( .A1(u5_mult_87_n440), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__4_) );
  NOR2_X1 u5_mult_87_U2664 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n338), .ZN(
        u5_mult_87_ab_1__50_) );
  NOR2_X1 u5_mult_87_U2663 ( .A1(u5_mult_87_n345), .A2(u5_mult_87_n337), .ZN(
        u5_mult_87_ab_1__51_) );
  NOR2_X1 u5_mult_87_U2662 ( .A1(u5_mult_87_n342), .A2(u5_mult_87_n337), .ZN(
        u5_mult_87_ab_1__52_) );
  NOR2_X1 u5_mult_87_U2661 ( .A1(u5_mult_87_n437), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__5_) );
  NOR2_X1 u5_mult_87_U2660 ( .A1(u5_mult_87_n436), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__6_) );
  NOR2_X1 u5_mult_87_U2659 ( .A1(u5_mult_87_n434), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__7_) );
  NOR2_X1 u5_mult_87_U2658 ( .A1(u5_mult_87_n432), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__8_) );
  NOR2_X1 u5_mult_87_U2657 ( .A1(u5_mult_87_n430), .A2(u5_mult_87_n336), .ZN(
        u5_mult_87_ab_1__9_) );
  NOR2_X1 u5_mult_87_U2656 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__0_) );
  NOR2_X1 u5_mult_87_U2655 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__10_) );
  NOR2_X1 u5_mult_87_U2654 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__11_) );
  NOR2_X1 u5_mult_87_U2653 ( .A1(u5_mult_87_n481), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__12_) );
  NOR2_X1 u5_mult_87_U2652 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__13_) );
  NOR2_X1 u5_mult_87_U2651 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__14_) );
  NOR2_X1 u5_mult_87_U2650 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__15_) );
  NOR2_X1 u5_mult_87_U2649 ( .A1(u5_mult_87_n480), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__16_) );
  NOR2_X1 u5_mult_87_U2648 ( .A1(u5_mult_87_n413), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__17_) );
  NOR2_X1 u5_mult_87_U2647 ( .A1(u5_mult_87_n411), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__18_) );
  NOR2_X1 u5_mult_87_U2646 ( .A1(u5_mult_87_n409), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__19_) );
  NOR2_X1 u5_mult_87_U2645 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n291), .ZN(
        u5_mult_87_ab_20__1_) );
  NOR2_X1 u5_mult_87_U2644 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n291), .ZN(
        u5_mult_87_ab_20__20_) );
  NOR2_X1 u5_mult_87_U2643 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__21_) );
  NOR2_X1 u5_mult_87_U2642 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__22_) );
  NOR2_X1 u5_mult_87_U2641 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__23_) );
  NOR2_X1 u5_mult_87_U2640 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__24_) );
  NOR2_X1 u5_mult_87_U2639 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__25_) );
  NOR2_X1 u5_mult_87_U2638 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__26_) );
  NOR2_X1 u5_mult_87_U2637 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__27_) );
  NOR2_X1 u5_mult_87_U2636 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__28_) );
  NOR2_X1 u5_mult_87_U2635 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n291), .ZN(
        u5_mult_87_ab_20__29_) );
  NOR2_X1 u5_mult_87_U2634 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n468), .ZN(
        u5_mult_87_ab_20__2_) );
  NOR2_X1 u5_mult_87_U2633 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n468), .ZN(
        u5_mult_87_ab_20__30_) );
  NOR2_X1 u5_mult_87_U2632 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n291), .ZN(
        u5_mult_87_ab_20__31_) );
  NOR2_X1 u5_mult_87_U2631 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n468), .ZN(
        u5_mult_87_ab_20__32_) );
  NOR2_X1 u5_mult_87_U2630 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n291), .ZN(
        u5_mult_87_ab_20__33_) );
  NOR2_X1 u5_mult_87_U2629 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n468), .ZN(
        u5_mult_87_ab_20__34_) );
  NOR2_X1 u5_mult_87_U2628 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n468), .ZN(
        u5_mult_87_ab_20__35_) );
  NOR2_X1 u5_mult_87_U2627 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n291), .ZN(
        u5_mult_87_ab_20__36_) );
  NOR2_X1 u5_mult_87_U2626 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n291), .ZN(
        u5_mult_87_ab_20__37_) );
  NOR2_X1 u5_mult_87_U2625 ( .A1(u5_mult_87_n372), .A2(u5_mult_87_n468), .ZN(
        u5_mult_87_ab_20__38_) );
  NOR2_X1 u5_mult_87_U2624 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n468), .ZN(
        u5_mult_87_ab_20__39_) );
  NOR2_X1 u5_mult_87_U2623 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n291), .ZN(
        u5_mult_87_ab_20__3_) );
  NOR2_X1 u5_mult_87_U2622 ( .A1(u5_mult_87_n367), .A2(u5_mult_87_n291), .ZN(
        u5_mult_87_ab_20__40_) );
  NOR2_X1 u5_mult_87_U2621 ( .A1(u5_mult_87_n365), .A2(u5_mult_87_n291), .ZN(
        u5_mult_87_ab_20__41_) );
  NOR2_X1 u5_mult_87_U2620 ( .A1(u5_mult_87_n363), .A2(u5_mult_87_n291), .ZN(
        u5_mult_87_ab_20__42_) );
  NOR2_X1 u5_mult_87_U2619 ( .A1(u5_mult_87_n360), .A2(u5_mult_87_n291), .ZN(
        u5_mult_87_ab_20__43_) );
  NOR2_X1 u5_mult_87_U2618 ( .A1(u5_mult_87_n358), .A2(u5_mult_87_n291), .ZN(
        u5_mult_87_ab_20__44_) );
  NOR2_X1 u5_mult_87_U2617 ( .A1(u5_mult_87_n356), .A2(u5_mult_87_n291), .ZN(
        u5_mult_87_ab_20__45_) );
  NOR2_X1 u5_mult_87_U2616 ( .A1(u5_mult_87_n354), .A2(u5_mult_87_n291), .ZN(
        u5_mult_87_ab_20__46_) );
  NOR2_X1 u5_mult_87_U2615 ( .A1(u5_mult_87_n351), .A2(u5_mult_87_n291), .ZN(
        u5_mult_87_ab_20__47_) );
  NOR2_X1 u5_mult_87_U2614 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n291), .ZN(
        u5_mult_87_ab_20__48_) );
  NOR2_X1 u5_mult_87_U2613 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n291), .ZN(
        u5_mult_87_ab_20__49_) );
  NOR2_X1 u5_mult_87_U2612 ( .A1(u5_mult_87_n440), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__4_) );
  NOR2_X1 u5_mult_87_U2611 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__50_) );
  NOR2_X1 u5_mult_87_U2610 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__51_) );
  NOR2_X1 u5_mult_87_U2609 ( .A1(u5_mult_87_n342), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__52_) );
  NOR2_X1 u5_mult_87_U2608 ( .A1(u5_mult_87_n437), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__5_) );
  NOR2_X1 u5_mult_87_U2607 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__6_) );
  NOR2_X1 u5_mult_87_U2606 ( .A1(u5_mult_87_n434), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__7_) );
  NOR2_X1 u5_mult_87_U2605 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__8_) );
  NOR2_X1 u5_mult_87_U2604 ( .A1(u5_mult_87_n430), .A2(u5_mult_87_n290), .ZN(
        u5_mult_87_ab_20__9_) );
  NOR2_X1 u5_mult_87_U2603 ( .A1(u5_mult_87_n450), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__0_) );
  NOR2_X1 u5_mult_87_U2602 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__10_) );
  NOR2_X1 u5_mult_87_U2601 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__11_) );
  NOR2_X1 u5_mult_87_U2600 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__12_) );
  NOR2_X1 u5_mult_87_U2599 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__13_) );
  NOR2_X1 u5_mult_87_U2598 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__14_) );
  NOR2_X1 u5_mult_87_U2597 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__15_) );
  NOR2_X1 u5_mult_87_U2596 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__16_) );
  NOR2_X1 u5_mult_87_U2595 ( .A1(u5_mult_87_n413), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__17_) );
  NOR2_X1 u5_mult_87_U2594 ( .A1(u5_mult_87_n411), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__18_) );
  NOR2_X1 u5_mult_87_U2593 ( .A1(u5_mult_87_n409), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__19_) );
  NOR2_X1 u5_mult_87_U2592 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n289), .ZN(
        u5_mult_87_ab_21__1_) );
  NOR2_X1 u5_mult_87_U2591 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__20_) );
  NOR2_X1 u5_mult_87_U2590 ( .A1(u5_mult_87_n406), .A2(u5_mult_87_n289), .ZN(
        u5_mult_87_ab_21__21_) );
  NOR2_X1 u5_mult_87_U2589 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n289), .ZN(
        u5_mult_87_ab_21__22_) );
  NOR2_X1 u5_mult_87_U2588 ( .A1(u5_mult_87_n402), .A2(u5_mult_87_n289), .ZN(
        u5_mult_87_ab_21__23_) );
  NOR2_X1 u5_mult_87_U2587 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n289), .ZN(
        u5_mult_87_ab_21__24_) );
  NOR2_X1 u5_mult_87_U2586 ( .A1(u5_mult_87_n398), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__25_) );
  NOR2_X1 u5_mult_87_U2585 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__26_) );
  NOR2_X1 u5_mult_87_U2584 ( .A1(u5_mult_87_n394), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__27_) );
  NOR2_X1 u5_mult_87_U2583 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__28_) );
  NOR2_X1 u5_mult_87_U2582 ( .A1(u5_mult_87_n390), .A2(u5_mult_87_n289), .ZN(
        u5_mult_87_ab_21__29_) );
  NOR2_X1 u5_mult_87_U2581 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n467), .ZN(
        u5_mult_87_ab_21__2_) );
  NOR2_X1 u5_mult_87_U2580 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n467), .ZN(
        u5_mult_87_ab_21__30_) );
  NOR2_X1 u5_mult_87_U2579 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n289), .ZN(
        u5_mult_87_ab_21__31_) );
  NOR2_X1 u5_mult_87_U2578 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n467), .ZN(
        u5_mult_87_ab_21__32_) );
  NOR2_X1 u5_mult_87_U2577 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n467), .ZN(
        u5_mult_87_ab_21__33_) );
  NOR2_X1 u5_mult_87_U2576 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n467), .ZN(
        u5_mult_87_ab_21__34_) );
  NOR2_X1 u5_mult_87_U2575 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n289), .ZN(
        u5_mult_87_ab_21__35_) );
  NOR2_X1 u5_mult_87_U2574 ( .A1(u5_mult_87_n376), .A2(u5_mult_87_n289), .ZN(
        u5_mult_87_ab_21__36_) );
  NOR2_X1 u5_mult_87_U2573 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n289), .ZN(
        u5_mult_87_ab_21__37_) );
  NOR2_X1 u5_mult_87_U2572 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n289), .ZN(
        u5_mult_87_ab_21__38_) );
  NOR2_X1 u5_mult_87_U2571 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n289), .ZN(
        u5_mult_87_ab_21__39_) );
  NOR2_X1 u5_mult_87_U2570 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n289), .ZN(
        u5_mult_87_ab_21__3_) );
  NOR2_X1 u5_mult_87_U2569 ( .A1(u5_mult_87_n367), .A2(u5_mult_87_n289), .ZN(
        u5_mult_87_ab_21__40_) );
  NOR2_X1 u5_mult_87_U2568 ( .A1(u5_mult_87_n365), .A2(u5_mult_87_n289), .ZN(
        u5_mult_87_ab_21__41_) );
  NOR2_X1 u5_mult_87_U2567 ( .A1(u5_mult_87_n363), .A2(u5_mult_87_n289), .ZN(
        u5_mult_87_ab_21__42_) );
  NOR2_X1 u5_mult_87_U2566 ( .A1(u5_mult_87_n360), .A2(u5_mult_87_n289), .ZN(
        u5_mult_87_ab_21__43_) );
  NOR2_X1 u5_mult_87_U2565 ( .A1(u5_mult_87_n358), .A2(u5_mult_87_n289), .ZN(
        u5_mult_87_ab_21__44_) );
  NOR2_X1 u5_mult_87_U2564 ( .A1(u5_mult_87_n356), .A2(u5_mult_87_n289), .ZN(
        u5_mult_87_ab_21__45_) );
  NOR2_X1 u5_mult_87_U2563 ( .A1(u5_mult_87_n354), .A2(u5_mult_87_n289), .ZN(
        u5_mult_87_ab_21__46_) );
  NOR2_X1 u5_mult_87_U2562 ( .A1(u5_mult_87_n351), .A2(u5_mult_87_n289), .ZN(
        u5_mult_87_ab_21__47_) );
  NOR2_X1 u5_mult_87_U2561 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n289), .ZN(
        u5_mult_87_ab_21__48_) );
  NOR2_X1 u5_mult_87_U2560 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n289), .ZN(
        u5_mult_87_ab_21__49_) );
  NOR2_X1 u5_mult_87_U2559 ( .A1(u5_mult_87_n440), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__4_) );
  NOR2_X1 u5_mult_87_U2558 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__50_) );
  NOR2_X1 u5_mult_87_U2557 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__51_) );
  NOR2_X1 u5_mult_87_U2556 ( .A1(u5_mult_87_n342), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__52_) );
  NOR2_X1 u5_mult_87_U2555 ( .A1(u5_mult_87_n437), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__5_) );
  NOR2_X1 u5_mult_87_U2554 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__6_) );
  NOR2_X1 u5_mult_87_U2553 ( .A1(u5_mult_87_n434), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__7_) );
  NOR2_X1 u5_mult_87_U2552 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__8_) );
  NOR2_X1 u5_mult_87_U2551 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n288), .ZN(
        u5_mult_87_ab_21__9_) );
  NOR2_X1 u5_mult_87_U2550 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__0_) );
  NOR2_X1 u5_mult_87_U2549 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__10_) );
  NOR2_X1 u5_mult_87_U2548 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__11_) );
  NOR2_X1 u5_mult_87_U2547 ( .A1(u5_mult_87_n481), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__12_) );
  NOR2_X1 u5_mult_87_U2546 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__13_) );
  NOR2_X1 u5_mult_87_U2545 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__14_) );
  NOR2_X1 u5_mult_87_U2544 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__15_) );
  NOR2_X1 u5_mult_87_U2543 ( .A1(u5_mult_87_n480), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__16_) );
  NOR2_X1 u5_mult_87_U2542 ( .A1(u5_mult_87_n413), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__17_) );
  NOR2_X1 u5_mult_87_U2541 ( .A1(u5_mult_87_n411), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__18_) );
  NOR2_X1 u5_mult_87_U2540 ( .A1(u5_mult_87_n409), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__19_) );
  NOR2_X1 u5_mult_87_U2539 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n287), .ZN(
        u5_mult_87_ab_22__1_) );
  NOR2_X1 u5_mult_87_U2538 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__20_) );
  NOR2_X1 u5_mult_87_U2537 ( .A1(u5_mult_87_n406), .A2(u5_mult_87_n287), .ZN(
        u5_mult_87_ab_22__21_) );
  NOR2_X1 u5_mult_87_U2536 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n287), .ZN(
        u5_mult_87_ab_22__22_) );
  NOR2_X1 u5_mult_87_U2535 ( .A1(u5_mult_87_n402), .A2(u5_mult_87_n287), .ZN(
        u5_mult_87_ab_22__23_) );
  NOR2_X1 u5_mult_87_U2534 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n287), .ZN(
        u5_mult_87_ab_22__24_) );
  NOR2_X1 u5_mult_87_U2533 ( .A1(u5_mult_87_n398), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__25_) );
  NOR2_X1 u5_mult_87_U2532 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__26_) );
  NOR2_X1 u5_mult_87_U2531 ( .A1(u5_mult_87_n394), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__27_) );
  NOR2_X1 u5_mult_87_U2530 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__28_) );
  NOR2_X1 u5_mult_87_U2529 ( .A1(u5_mult_87_n390), .A2(u5_mult_87_n287), .ZN(
        u5_mult_87_ab_22__29_) );
  NOR2_X1 u5_mult_87_U2528 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n466), .ZN(
        u5_mult_87_ab_22__2_) );
  NOR2_X1 u5_mult_87_U2527 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n287), .ZN(
        u5_mult_87_ab_22__30_) );
  NOR2_X1 u5_mult_87_U2526 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n287), .ZN(
        u5_mult_87_ab_22__31_) );
  NOR2_X1 u5_mult_87_U2525 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n466), .ZN(
        u5_mult_87_ab_22__32_) );
  NOR2_X1 u5_mult_87_U2524 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n466), .ZN(
        u5_mult_87_ab_22__33_) );
  NOR2_X1 u5_mult_87_U2523 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n287), .ZN(
        u5_mult_87_ab_22__34_) );
  NOR2_X1 u5_mult_87_U2522 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n287), .ZN(
        u5_mult_87_ab_22__35_) );
  NOR2_X1 u5_mult_87_U2521 ( .A1(u5_mult_87_n376), .A2(u5_mult_87_n466), .ZN(
        u5_mult_87_ab_22__36_) );
  NOR2_X1 u5_mult_87_U2520 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n466), .ZN(
        u5_mult_87_ab_22__37_) );
  NOR2_X1 u5_mult_87_U2519 ( .A1(u5_mult_87_n372), .A2(u5_mult_87_n466), .ZN(
        u5_mult_87_ab_22__38_) );
  NOR2_X1 u5_mult_87_U2518 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n466), .ZN(
        u5_mult_87_ab_22__39_) );
  NOR2_X1 u5_mult_87_U2517 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n287), .ZN(
        u5_mult_87_ab_22__3_) );
  NOR2_X1 u5_mult_87_U2516 ( .A1(u5_mult_87_n367), .A2(u5_mult_87_n287), .ZN(
        u5_mult_87_ab_22__40_) );
  NOR2_X1 u5_mult_87_U2515 ( .A1(u5_mult_87_n365), .A2(u5_mult_87_n287), .ZN(
        u5_mult_87_ab_22__41_) );
  NOR2_X1 u5_mult_87_U2514 ( .A1(u5_mult_87_n364), .A2(u5_mult_87_n287), .ZN(
        u5_mult_87_ab_22__42_) );
  NOR2_X1 u5_mult_87_U2513 ( .A1(u5_mult_87_n360), .A2(u5_mult_87_n287), .ZN(
        u5_mult_87_ab_22__43_) );
  NOR2_X1 u5_mult_87_U2512 ( .A1(u5_mult_87_n358), .A2(u5_mult_87_n287), .ZN(
        u5_mult_87_ab_22__44_) );
  NOR2_X1 u5_mult_87_U2511 ( .A1(u5_mult_87_n356), .A2(u5_mult_87_n287), .ZN(
        u5_mult_87_ab_22__45_) );
  NOR2_X1 u5_mult_87_U2510 ( .A1(u5_mult_87_n354), .A2(u5_mult_87_n287), .ZN(
        u5_mult_87_ab_22__46_) );
  NOR2_X1 u5_mult_87_U2509 ( .A1(u5_mult_87_n351), .A2(u5_mult_87_n287), .ZN(
        u5_mult_87_ab_22__47_) );
  NOR2_X1 u5_mult_87_U2508 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n287), .ZN(
        u5_mult_87_ab_22__48_) );
  NOR2_X1 u5_mult_87_U2507 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n287), .ZN(
        u5_mult_87_ab_22__49_) );
  NOR2_X1 u5_mult_87_U2506 ( .A1(u5_mult_87_n440), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__4_) );
  NOR2_X1 u5_mult_87_U2505 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__50_) );
  NOR2_X1 u5_mult_87_U2504 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__51_) );
  NOR2_X1 u5_mult_87_U2503 ( .A1(u5_mult_87_n342), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__52_) );
  NOR2_X1 u5_mult_87_U2502 ( .A1(u5_mult_87_n437), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__5_) );
  NOR2_X1 u5_mult_87_U2501 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__6_) );
  NOR2_X1 u5_mult_87_U2500 ( .A1(u5_mult_87_n434), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__7_) );
  NOR2_X1 u5_mult_87_U2499 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__8_) );
  NOR2_X1 u5_mult_87_U2498 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n286), .ZN(
        u5_mult_87_ab_22__9_) );
  NOR2_X1 u5_mult_87_U2497 ( .A1(u5_mult_87_n450), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__0_) );
  NOR2_X1 u5_mult_87_U2496 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__10_) );
  NOR2_X1 u5_mult_87_U2495 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__11_) );
  NOR2_X1 u5_mult_87_U2494 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__12_) );
  NOR2_X1 u5_mult_87_U2493 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__13_) );
  NOR2_X1 u5_mult_87_U2492 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__14_) );
  NOR2_X1 u5_mult_87_U2491 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__15_) );
  NOR2_X1 u5_mult_87_U2490 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__16_) );
  NOR2_X1 u5_mult_87_U2489 ( .A1(u5_mult_87_n413), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__17_) );
  NOR2_X1 u5_mult_87_U2488 ( .A1(u5_mult_87_n411), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__18_) );
  NOR2_X1 u5_mult_87_U2487 ( .A1(u5_mult_87_n409), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__19_) );
  NOR2_X1 u5_mult_87_U2486 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n285), .ZN(
        u5_mult_87_ab_23__1_) );
  NOR2_X1 u5_mult_87_U2485 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__20_) );
  NOR2_X1 u5_mult_87_U2484 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n285), .ZN(
        u5_mult_87_ab_23__21_) );
  NOR2_X1 u5_mult_87_U2483 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n285), .ZN(
        u5_mult_87_ab_23__22_) );
  NOR2_X1 u5_mult_87_U2482 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n285), .ZN(
        u5_mult_87_ab_23__23_) );
  NOR2_X1 u5_mult_87_U2481 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n285), .ZN(
        u5_mult_87_ab_23__24_) );
  NOR2_X1 u5_mult_87_U2480 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__25_) );
  NOR2_X1 u5_mult_87_U2479 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__26_) );
  NOR2_X1 u5_mult_87_U2478 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__27_) );
  NOR2_X1 u5_mult_87_U2477 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__28_) );
  NOR2_X1 u5_mult_87_U2476 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n285), .ZN(
        u5_mult_87_ab_23__29_) );
  NOR2_X1 u5_mult_87_U2475 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n465), .ZN(
        u5_mult_87_ab_23__2_) );
  NOR2_X1 u5_mult_87_U2474 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n285), .ZN(
        u5_mult_87_ab_23__30_) );
  NOR2_X1 u5_mult_87_U2473 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n285), .ZN(
        u5_mult_87_ab_23__31_) );
  NOR2_X1 u5_mult_87_U2472 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n285), .ZN(
        u5_mult_87_ab_23__32_) );
  NOR2_X1 u5_mult_87_U2471 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n285), .ZN(
        u5_mult_87_ab_23__33_) );
  NOR2_X1 u5_mult_87_U2470 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n465), .ZN(
        u5_mult_87_ab_23__34_) );
  NOR2_X1 u5_mult_87_U2469 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n285), .ZN(
        u5_mult_87_ab_23__35_) );
  NOR2_X1 u5_mult_87_U2468 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n465), .ZN(
        u5_mult_87_ab_23__36_) );
  NOR2_X1 u5_mult_87_U2467 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n465), .ZN(
        u5_mult_87_ab_23__37_) );
  NOR2_X1 u5_mult_87_U2466 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n465), .ZN(
        u5_mult_87_ab_23__38_) );
  NOR2_X1 u5_mult_87_U2465 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n465), .ZN(
        u5_mult_87_ab_23__39_) );
  NOR2_X1 u5_mult_87_U2464 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n285), .ZN(
        u5_mult_87_ab_23__3_) );
  NOR2_X1 u5_mult_87_U2463 ( .A1(u5_mult_87_n367), .A2(u5_mult_87_n285), .ZN(
        u5_mult_87_ab_23__40_) );
  NOR2_X1 u5_mult_87_U2462 ( .A1(u5_mult_87_n365), .A2(u5_mult_87_n285), .ZN(
        u5_mult_87_ab_23__41_) );
  NOR2_X1 u5_mult_87_U2461 ( .A1(u5_mult_87_n364), .A2(u5_mult_87_n285), .ZN(
        u5_mult_87_ab_23__42_) );
  NOR2_X1 u5_mult_87_U2460 ( .A1(u5_mult_87_n360), .A2(u5_mult_87_n285), .ZN(
        u5_mult_87_ab_23__43_) );
  NOR2_X1 u5_mult_87_U2459 ( .A1(u5_mult_87_n358), .A2(u5_mult_87_n285), .ZN(
        u5_mult_87_ab_23__44_) );
  NOR2_X1 u5_mult_87_U2458 ( .A1(u5_mult_87_n356), .A2(u5_mult_87_n285), .ZN(
        u5_mult_87_ab_23__45_) );
  NOR2_X1 u5_mult_87_U2457 ( .A1(u5_mult_87_n354), .A2(u5_mult_87_n285), .ZN(
        u5_mult_87_ab_23__46_) );
  NOR2_X1 u5_mult_87_U2456 ( .A1(u5_mult_87_n351), .A2(u5_mult_87_n285), .ZN(
        u5_mult_87_ab_23__47_) );
  NOR2_X1 u5_mult_87_U2455 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n285), .ZN(
        u5_mult_87_ab_23__48_) );
  NOR2_X1 u5_mult_87_U2454 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n285), .ZN(
        u5_mult_87_ab_23__49_) );
  NOR2_X1 u5_mult_87_U2453 ( .A1(u5_mult_87_n440), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__4_) );
  NOR2_X1 u5_mult_87_U2452 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__50_) );
  NOR2_X1 u5_mult_87_U2451 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__51_) );
  NOR2_X1 u5_mult_87_U2450 ( .A1(u5_mult_87_n342), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__52_) );
  NOR2_X1 u5_mult_87_U2449 ( .A1(u5_mult_87_n437), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__5_) );
  NOR2_X1 u5_mult_87_U2448 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__6_) );
  NOR2_X1 u5_mult_87_U2447 ( .A1(u5_mult_87_n434), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__7_) );
  NOR2_X1 u5_mult_87_U2446 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__8_) );
  NOR2_X1 u5_mult_87_U2445 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n284), .ZN(
        u5_mult_87_ab_23__9_) );
  NOR2_X1 u5_mult_87_U2444 ( .A1(u5_mult_87_n450), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__0_) );
  NOR2_X1 u5_mult_87_U2443 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__10_) );
  NOR2_X1 u5_mult_87_U2442 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__11_) );
  NOR2_X1 u5_mult_87_U2441 ( .A1(u5_mult_87_n481), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__12_) );
  NOR2_X1 u5_mult_87_U2440 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__13_) );
  NOR2_X1 u5_mult_87_U2439 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__14_) );
  NOR2_X1 u5_mult_87_U2438 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__15_) );
  NOR2_X1 u5_mult_87_U2437 ( .A1(u5_mult_87_n480), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__16_) );
  NOR2_X1 u5_mult_87_U2436 ( .A1(u5_mult_87_n413), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__17_) );
  NOR2_X1 u5_mult_87_U2435 ( .A1(u5_mult_87_n411), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__18_) );
  NOR2_X1 u5_mult_87_U2434 ( .A1(u5_mult_87_n409), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__19_) );
  NOR2_X1 u5_mult_87_U2433 ( .A1(u5_mult_87_n446), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__1_) );
  NOR2_X1 u5_mult_87_U2432 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__20_) );
  NOR2_X1 u5_mult_87_U2431 ( .A1(u5_mult_87_n406), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__21_) );
  NOR2_X1 u5_mult_87_U2430 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__22_) );
  NOR2_X1 u5_mult_87_U2429 ( .A1(u5_mult_87_n402), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__23_) );
  NOR2_X1 u5_mult_87_U2428 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__24_) );
  NOR2_X1 u5_mult_87_U2427 ( .A1(u5_mult_87_n398), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__25_) );
  NOR2_X1 u5_mult_87_U2426 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__26_) );
  NOR2_X1 u5_mult_87_U2425 ( .A1(u5_mult_87_n394), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__27_) );
  NOR2_X1 u5_mult_87_U2424 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__28_) );
  NOR2_X1 u5_mult_87_U2423 ( .A1(u5_mult_87_n390), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__29_) );
  NOR2_X1 u5_mult_87_U2422 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__2_) );
  NOR2_X1 u5_mult_87_U2421 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__30_) );
  NOR2_X1 u5_mult_87_U2420 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__31_) );
  NOR2_X1 u5_mult_87_U2419 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__32_) );
  NOR2_X1 u5_mult_87_U2418 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__33_) );
  NOR2_X1 u5_mult_87_U2417 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__34_) );
  NOR2_X1 u5_mult_87_U2416 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__35_) );
  NOR2_X1 u5_mult_87_U2415 ( .A1(u5_mult_87_n376), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__36_) );
  NOR2_X1 u5_mult_87_U2414 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__37_) );
  NOR2_X1 u5_mult_87_U2413 ( .A1(u5_mult_87_n372), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__38_) );
  NOR2_X1 u5_mult_87_U2412 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__39_) );
  NOR2_X1 u5_mult_87_U2411 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__3_) );
  NOR2_X1 u5_mult_87_U2410 ( .A1(u5_mult_87_n367), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__40_) );
  NOR2_X1 u5_mult_87_U2409 ( .A1(u5_mult_87_n365), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__41_) );
  NOR2_X1 u5_mult_87_U2408 ( .A1(u5_mult_87_n364), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__42_) );
  NOR2_X1 u5_mult_87_U2407 ( .A1(u5_mult_87_n360), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__43_) );
  NOR2_X1 u5_mult_87_U2406 ( .A1(u5_mult_87_n358), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__44_) );
  NOR2_X1 u5_mult_87_U2405 ( .A1(u5_mult_87_n356), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__45_) );
  NOR2_X1 u5_mult_87_U2404 ( .A1(u5_mult_87_n354), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__46_) );
  NOR2_X1 u5_mult_87_U2403 ( .A1(u5_mult_87_n351), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__47_) );
  NOR2_X1 u5_mult_87_U2402 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__48_) );
  NOR2_X1 u5_mult_87_U2401 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n283), .ZN(
        u5_mult_87_ab_24__49_) );
  NOR2_X1 u5_mult_87_U2400 ( .A1(u5_mult_87_n440), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__4_) );
  NOR2_X1 u5_mult_87_U2399 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__50_) );
  NOR2_X1 u5_mult_87_U2398 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__51_) );
  NOR2_X1 u5_mult_87_U2397 ( .A1(u5_mult_87_n342), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__52_) );
  NOR2_X1 u5_mult_87_U2396 ( .A1(u5_mult_87_n437), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__5_) );
  NOR2_X1 u5_mult_87_U2395 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__6_) );
  NOR2_X1 u5_mult_87_U2394 ( .A1(u5_mult_87_n434), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__7_) );
  NOR2_X1 u5_mult_87_U2393 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__8_) );
  NOR2_X1 u5_mult_87_U2392 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n282), .ZN(
        u5_mult_87_ab_24__9_) );
  NOR2_X1 u5_mult_87_U2391 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__0_) );
  NOR2_X1 u5_mult_87_U2390 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__10_) );
  NOR2_X1 u5_mult_87_U2389 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__11_) );
  NOR2_X1 u5_mult_87_U2388 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__12_) );
  NOR2_X1 u5_mult_87_U2387 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__13_) );
  NOR2_X1 u5_mult_87_U2386 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__14_) );
  NOR2_X1 u5_mult_87_U2385 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__15_) );
  NOR2_X1 u5_mult_87_U2384 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__16_) );
  NOR2_X1 u5_mult_87_U2383 ( .A1(u5_mult_87_n413), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__17_) );
  NOR2_X1 u5_mult_87_U2382 ( .A1(u5_mult_87_n411), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__18_) );
  NOR2_X1 u5_mult_87_U2381 ( .A1(u5_mult_87_n409), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__19_) );
  NOR2_X1 u5_mult_87_U2380 ( .A1(u5_mult_87_n446), .A2(u5_mult_87_n464), .ZN(
        u5_mult_87_ab_25__1_) );
  NOR2_X1 u5_mult_87_U2379 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__20_) );
  NOR2_X1 u5_mult_87_U2378 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__21_) );
  NOR2_X1 u5_mult_87_U2377 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__22_) );
  NOR2_X1 u5_mult_87_U2376 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__23_) );
  NOR2_X1 u5_mult_87_U2375 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n464), .ZN(
        u5_mult_87_ab_25__24_) );
  NOR2_X1 u5_mult_87_U2374 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n464), .ZN(
        u5_mult_87_ab_25__25_) );
  NOR2_X1 u5_mult_87_U2373 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n464), .ZN(
        u5_mult_87_ab_25__26_) );
  NOR2_X1 u5_mult_87_U2372 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n464), .ZN(
        u5_mult_87_ab_25__27_) );
  NOR2_X1 u5_mult_87_U2371 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n464), .ZN(
        u5_mult_87_ab_25__28_) );
  NOR2_X1 u5_mult_87_U2370 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n464), .ZN(
        u5_mult_87_ab_25__29_) );
  NOR2_X1 u5_mult_87_U2369 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n464), .ZN(
        u5_mult_87_ab_25__2_) );
  NOR2_X1 u5_mult_87_U2368 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n464), .ZN(
        u5_mult_87_ab_25__30_) );
  NOR2_X1 u5_mult_87_U2367 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n464), .ZN(
        u5_mult_87_ab_25__31_) );
  NOR2_X1 u5_mult_87_U2366 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n464), .ZN(
        u5_mult_87_ab_25__32_) );
  NOR2_X1 u5_mult_87_U2365 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n464), .ZN(
        u5_mult_87_ab_25__33_) );
  NOR2_X1 u5_mult_87_U2364 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n464), .ZN(
        u5_mult_87_ab_25__34_) );
  NOR2_X1 u5_mult_87_U2363 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n464), .ZN(
        u5_mult_87_ab_25__35_) );
  NOR2_X1 u5_mult_87_U2362 ( .A1(u5_mult_87_n376), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__36_) );
  NOR2_X1 u5_mult_87_U2361 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__37_) );
  NOR2_X1 u5_mult_87_U2360 ( .A1(u5_mult_87_n372), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__38_) );
  NOR2_X1 u5_mult_87_U2359 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__39_) );
  NOR2_X1 u5_mult_87_U2358 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__3_) );
  NOR2_X1 u5_mult_87_U2357 ( .A1(u5_mult_87_n367), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__40_) );
  NOR2_X1 u5_mult_87_U2356 ( .A1(u5_mult_87_n365), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__41_) );
  NOR2_X1 u5_mult_87_U2355 ( .A1(u5_mult_87_n364), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__42_) );
  NOR2_X1 u5_mult_87_U2354 ( .A1(u5_mult_87_n360), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__43_) );
  NOR2_X1 u5_mult_87_U2353 ( .A1(u5_mult_87_n358), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__44_) );
  NOR2_X1 u5_mult_87_U2352 ( .A1(u5_mult_87_n356), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__45_) );
  NOR2_X1 u5_mult_87_U2351 ( .A1(u5_mult_87_n354), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__46_) );
  NOR2_X1 u5_mult_87_U2350 ( .A1(u5_mult_87_n351), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__47_) );
  NOR2_X1 u5_mult_87_U2349 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__48_) );
  NOR2_X1 u5_mult_87_U2348 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__49_) );
  NOR2_X1 u5_mult_87_U2347 ( .A1(u5_mult_87_n440), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__4_) );
  NOR2_X1 u5_mult_87_U2346 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__50_) );
  NOR2_X1 u5_mult_87_U2345 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__51_) );
  NOR2_X1 u5_mult_87_U2344 ( .A1(u5_mult_87_n342), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__52_) );
  NOR2_X1 u5_mult_87_U2343 ( .A1(u5_mult_87_n437), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__5_) );
  NOR2_X1 u5_mult_87_U2342 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__6_) );
  NOR2_X1 u5_mult_87_U2341 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__7_) );
  NOR2_X1 u5_mult_87_U2340 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__8_) );
  NOR2_X1 u5_mult_87_U2339 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n281), .ZN(
        u5_mult_87_ab_25__9_) );
  NOR2_X1 u5_mult_87_U2338 ( .A1(u5_mult_87_n450), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__0_) );
  NOR2_X1 u5_mult_87_U2337 ( .A1(u5_mult_87_n428), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__10_) );
  NOR2_X1 u5_mult_87_U2336 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__11_) );
  NOR2_X1 u5_mult_87_U2335 ( .A1(u5_mult_87_n481), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__12_) );
  NOR2_X1 u5_mult_87_U2334 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__13_) );
  NOR2_X1 u5_mult_87_U2333 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__14_) );
  NOR2_X1 u5_mult_87_U2332 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__15_) );
  NOR2_X1 u5_mult_87_U2331 ( .A1(u5_mult_87_n480), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__16_) );
  NOR2_X1 u5_mult_87_U2330 ( .A1(u5_mult_87_n413), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__17_) );
  NOR2_X1 u5_mult_87_U2329 ( .A1(u5_mult_87_n411), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__18_) );
  NOR2_X1 u5_mult_87_U2328 ( .A1(u5_mult_87_n409), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__19_) );
  NOR2_X1 u5_mult_87_U2327 ( .A1(u5_mult_87_n446), .A2(u5_mult_87_n280), .ZN(
        u5_mult_87_ab_26__1_) );
  NOR2_X1 u5_mult_87_U2326 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n280), .ZN(
        u5_mult_87_ab_26__20_) );
  NOR2_X1 u5_mult_87_U2325 ( .A1(u5_mult_87_n406), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__21_) );
  NOR2_X1 u5_mult_87_U2324 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__22_) );
  NOR2_X1 u5_mult_87_U2323 ( .A1(u5_mult_87_n402), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__23_) );
  NOR2_X1 u5_mult_87_U2322 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n280), .ZN(
        u5_mult_87_ab_26__24_) );
  NOR2_X1 u5_mult_87_U2321 ( .A1(u5_mult_87_n398), .A2(u5_mult_87_n280), .ZN(
        u5_mult_87_ab_26__25_) );
  NOR2_X1 u5_mult_87_U2320 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n280), .ZN(
        u5_mult_87_ab_26__26_) );
  NOR2_X1 u5_mult_87_U2319 ( .A1(u5_mult_87_n394), .A2(u5_mult_87_n280), .ZN(
        u5_mult_87_ab_26__27_) );
  NOR2_X1 u5_mult_87_U2318 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n280), .ZN(
        u5_mult_87_ab_26__28_) );
  NOR2_X1 u5_mult_87_U2317 ( .A1(u5_mult_87_n390), .A2(u5_mult_87_n280), .ZN(
        u5_mult_87_ab_26__29_) );
  NOR2_X1 u5_mult_87_U2316 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__2_) );
  NOR2_X1 u5_mult_87_U2315 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n280), .ZN(
        u5_mult_87_ab_26__30_) );
  NOR2_X1 u5_mult_87_U2314 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n280), .ZN(
        u5_mult_87_ab_26__31_) );
  NOR2_X1 u5_mult_87_U2313 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n280), .ZN(
        u5_mult_87_ab_26__32_) );
  NOR2_X1 u5_mult_87_U2312 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n280), .ZN(
        u5_mult_87_ab_26__33_) );
  NOR2_X1 u5_mult_87_U2311 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n280), .ZN(
        u5_mult_87_ab_26__34_) );
  NOR2_X1 u5_mult_87_U2310 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__35_) );
  NOR2_X1 u5_mult_87_U2309 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n280), .ZN(
        u5_mult_87_ab_26__36_) );
  NOR2_X1 u5_mult_87_U2308 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n280), .ZN(
        u5_mult_87_ab_26__37_) );
  NOR2_X1 u5_mult_87_U2307 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__38_) );
  NOR2_X1 u5_mult_87_U2306 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__39_) );
  NOR2_X1 u5_mult_87_U2305 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__3_) );
  NOR2_X1 u5_mult_87_U2304 ( .A1(u5_mult_87_n367), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__40_) );
  NOR2_X1 u5_mult_87_U2303 ( .A1(u5_mult_87_n365), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__41_) );
  NOR2_X1 u5_mult_87_U2302 ( .A1(u5_mult_87_n364), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__42_) );
  NOR2_X1 u5_mult_87_U2301 ( .A1(u5_mult_87_n360), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__43_) );
  NOR2_X1 u5_mult_87_U2300 ( .A1(u5_mult_87_n358), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__44_) );
  NOR2_X1 u5_mult_87_U2299 ( .A1(u5_mult_87_n356), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__45_) );
  NOR2_X1 u5_mult_87_U2298 ( .A1(u5_mult_87_n354), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__46_) );
  NOR2_X1 u5_mult_87_U2297 ( .A1(u5_mult_87_n351), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__47_) );
  NOR2_X1 u5_mult_87_U2296 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__48_) );
  NOR2_X1 u5_mult_87_U2295 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__49_) );
  NOR2_X1 u5_mult_87_U2294 ( .A1(u5_mult_87_n440), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__4_) );
  NOR2_X1 u5_mult_87_U2293 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__50_) );
  NOR2_X1 u5_mult_87_U2292 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__51_) );
  NOR2_X1 u5_mult_87_U2291 ( .A1(u5_mult_87_n342), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__52_) );
  NOR2_X1 u5_mult_87_U2290 ( .A1(u5_mult_87_n437), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__5_) );
  NOR2_X1 u5_mult_87_U2289 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__6_) );
  NOR2_X1 u5_mult_87_U2288 ( .A1(u5_mult_87_n434), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__7_) );
  NOR2_X1 u5_mult_87_U2287 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__8_) );
  NOR2_X1 u5_mult_87_U2286 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n279), .ZN(
        u5_mult_87_ab_26__9_) );
  NOR2_X1 u5_mult_87_U2285 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n278), .ZN(
        u5_mult_87_ab_27__0_) );
  NOR2_X1 u5_mult_87_U2284 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n278), .ZN(
        u5_mult_87_ab_27__10_) );
  NOR2_X1 u5_mult_87_U2283 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n463), .ZN(
        u5_mult_87_ab_27__11_) );
  NOR2_X1 u5_mult_87_U2282 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n278), .ZN(
        u5_mult_87_ab_27__12_) );
  NOR2_X1 u5_mult_87_U2281 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n278), .ZN(
        u5_mult_87_ab_27__13_) );
  NOR2_X1 u5_mult_87_U2280 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n463), .ZN(
        u5_mult_87_ab_27__14_) );
  NOR2_X1 u5_mult_87_U2279 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n278), .ZN(
        u5_mult_87_ab_27__15_) );
  NOR2_X1 u5_mult_87_U2278 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n277), .ZN(
        u5_mult_87_ab_27__16_) );
  NOR2_X1 u5_mult_87_U2277 ( .A1(u5_mult_87_n413), .A2(u5_mult_87_n278), .ZN(
        u5_mult_87_ab_27__17_) );
  NOR2_X1 u5_mult_87_U2276 ( .A1(u5_mult_87_n411), .A2(u5_mult_87_n278), .ZN(
        u5_mult_87_ab_27__18_) );
  NOR2_X1 u5_mult_87_U2275 ( .A1(u5_mult_87_n409), .A2(u5_mult_87_n278), .ZN(
        u5_mult_87_ab_27__19_) );
  NOR2_X1 u5_mult_87_U2274 ( .A1(u5_mult_87_n446), .A2(u5_mult_87_n277), .ZN(
        u5_mult_87_ab_27__1_) );
  NOR2_X1 u5_mult_87_U2273 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n277), .ZN(
        u5_mult_87_ab_27__20_) );
  NOR2_X1 u5_mult_87_U2272 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n277), .ZN(
        u5_mult_87_ab_27__21_) );
  NOR2_X1 u5_mult_87_U2271 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n277), .ZN(
        u5_mult_87_ab_27__22_) );
  NOR2_X1 u5_mult_87_U2270 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n277), .ZN(
        u5_mult_87_ab_27__23_) );
  NOR2_X1 u5_mult_87_U2269 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n277), .ZN(
        u5_mult_87_ab_27__24_) );
  NOR2_X1 u5_mult_87_U2268 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n277), .ZN(
        u5_mult_87_ab_27__25_) );
  NOR2_X1 u5_mult_87_U2267 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n277), .ZN(
        u5_mult_87_ab_27__26_) );
  NOR2_X1 u5_mult_87_U2266 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n277), .ZN(
        u5_mult_87_ab_27__27_) );
  NOR2_X1 u5_mult_87_U2265 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n277), .ZN(
        u5_mult_87_ab_27__28_) );
  NOR2_X1 u5_mult_87_U2264 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n277), .ZN(
        u5_mult_87_ab_27__29_) );
  NOR2_X1 u5_mult_87_U2263 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n278), .ZN(
        u5_mult_87_ab_27__2_) );
  NOR2_X1 u5_mult_87_U2262 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n278), .ZN(
        u5_mult_87_ab_27__30_) );
  NOR2_X1 u5_mult_87_U2261 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n278), .ZN(
        u5_mult_87_ab_27__31_) );
  NOR2_X1 u5_mult_87_U2260 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n278), .ZN(
        u5_mult_87_ab_27__32_) );
  NOR2_X1 u5_mult_87_U2259 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n278), .ZN(
        u5_mult_87_ab_27__33_) );
  NOR2_X1 u5_mult_87_U2258 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n278), .ZN(
        u5_mult_87_ab_27__34_) );
  NOR2_X1 u5_mult_87_U2257 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n278), .ZN(
        u5_mult_87_ab_27__35_) );
  NOR2_X1 u5_mult_87_U2256 ( .A1(u5_mult_87_n376), .A2(u5_mult_87_n278), .ZN(
        u5_mult_87_ab_27__36_) );
  NOR2_X1 u5_mult_87_U2255 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n278), .ZN(
        u5_mult_87_ab_27__37_) );
  NOR2_X1 u5_mult_87_U2254 ( .A1(u5_mult_87_n372), .A2(u5_mult_87_n278), .ZN(
        u5_mult_87_ab_27__38_) );
  NOR2_X1 u5_mult_87_U2253 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n278), .ZN(
        u5_mult_87_ab_27__39_) );
  NOR2_X1 u5_mult_87_U2252 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n463), .ZN(
        u5_mult_87_ab_27__3_) );
  NOR2_X1 u5_mult_87_U2251 ( .A1(u5_mult_87_n367), .A2(u5_mult_87_n277), .ZN(
        u5_mult_87_ab_27__40_) );
  NOR2_X1 u5_mult_87_U2250 ( .A1(u5_mult_87_n365), .A2(u5_mult_87_n277), .ZN(
        u5_mult_87_ab_27__41_) );
  NOR2_X1 u5_mult_87_U2249 ( .A1(u5_mult_87_n364), .A2(u5_mult_87_n277), .ZN(
        u5_mult_87_ab_27__42_) );
  NOR2_X1 u5_mult_87_U2248 ( .A1(u5_mult_87_n360), .A2(u5_mult_87_n277), .ZN(
        u5_mult_87_ab_27__43_) );
  NOR2_X1 u5_mult_87_U2247 ( .A1(u5_mult_87_n358), .A2(u5_mult_87_n278), .ZN(
        u5_mult_87_ab_27__44_) );
  NOR2_X1 u5_mult_87_U2246 ( .A1(u5_mult_87_n356), .A2(u5_mult_87_n463), .ZN(
        u5_mult_87_ab_27__45_) );
  NOR2_X1 u5_mult_87_U2245 ( .A1(u5_mult_87_n354), .A2(u5_mult_87_n463), .ZN(
        u5_mult_87_ab_27__46_) );
  NOR2_X1 u5_mult_87_U2244 ( .A1(u5_mult_87_n351), .A2(u5_mult_87_n463), .ZN(
        u5_mult_87_ab_27__47_) );
  NOR2_X1 u5_mult_87_U2243 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n463), .ZN(
        u5_mult_87_ab_27__48_) );
  NOR2_X1 u5_mult_87_U2242 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n463), .ZN(
        u5_mult_87_ab_27__49_) );
  NOR2_X1 u5_mult_87_U2241 ( .A1(u5_mult_87_n440), .A2(u5_mult_87_n463), .ZN(
        u5_mult_87_ab_27__4_) );
  NOR2_X1 u5_mult_87_U2240 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n463), .ZN(
        u5_mult_87_ab_27__50_) );
  NOR2_X1 u5_mult_87_U2239 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n463), .ZN(
        u5_mult_87_ab_27__51_) );
  NOR2_X1 u5_mult_87_U2238 ( .A1(u5_mult_87_n342), .A2(u5_mult_87_n463), .ZN(
        u5_mult_87_ab_27__52_) );
  NOR2_X1 u5_mult_87_U2237 ( .A1(u5_mult_87_n437), .A2(u5_mult_87_n463), .ZN(
        u5_mult_87_ab_27__5_) );
  NOR2_X1 u5_mult_87_U2236 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n463), .ZN(
        u5_mult_87_ab_27__6_) );
  NOR2_X1 u5_mult_87_U2235 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n463), .ZN(
        u5_mult_87_ab_27__7_) );
  NOR2_X1 u5_mult_87_U2234 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n463), .ZN(
        u5_mult_87_ab_27__8_) );
  NOR2_X1 u5_mult_87_U2233 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n463), .ZN(
        u5_mult_87_ab_27__9_) );
  NOR2_X1 u5_mult_87_U2232 ( .A1(u5_mult_87_n450), .A2(u5_mult_87_n275), .ZN(
        u5_mult_87_ab_28__0_) );
  NOR2_X1 u5_mult_87_U2231 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n275), .ZN(
        u5_mult_87_ab_28__10_) );
  NOR2_X1 u5_mult_87_U2230 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n275), .ZN(
        u5_mult_87_ab_28__11_) );
  NOR2_X1 u5_mult_87_U2229 ( .A1(u5_mult_87_n481), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__12_) );
  NOR2_X1 u5_mult_87_U2228 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__13_) );
  NOR2_X1 u5_mult_87_U2227 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__14_) );
  NOR2_X1 u5_mult_87_U2226 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__15_) );
  NOR2_X1 u5_mult_87_U2225 ( .A1(u5_mult_87_n480), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__16_) );
  NOR2_X1 u5_mult_87_U2224 ( .A1(u5_mult_87_n413), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__17_) );
  NOR2_X1 u5_mult_87_U2223 ( .A1(u5_mult_87_n411), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__18_) );
  NOR2_X1 u5_mult_87_U2222 ( .A1(u5_mult_87_n409), .A2(u5_mult_87_n275), .ZN(
        u5_mult_87_ab_28__19_) );
  NOR2_X1 u5_mult_87_U2221 ( .A1(u5_mult_87_n446), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__1_) );
  NOR2_X1 u5_mult_87_U2220 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__20_) );
  NOR2_X1 u5_mult_87_U2219 ( .A1(u5_mult_87_n406), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__21_) );
  NOR2_X1 u5_mult_87_U2218 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n462), .ZN(
        u5_mult_87_ab_28__22_) );
  NOR2_X1 u5_mult_87_U2217 ( .A1(u5_mult_87_n402), .A2(u5_mult_87_n462), .ZN(
        u5_mult_87_ab_28__23_) );
  NOR2_X1 u5_mult_87_U2216 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n462), .ZN(
        u5_mult_87_ab_28__24_) );
  NOR2_X1 u5_mult_87_U2215 ( .A1(u5_mult_87_n398), .A2(u5_mult_87_n462), .ZN(
        u5_mult_87_ab_28__25_) );
  NOR2_X1 u5_mult_87_U2214 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n462), .ZN(
        u5_mult_87_ab_28__26_) );
  NOR2_X1 u5_mult_87_U2213 ( .A1(u5_mult_87_n394), .A2(u5_mult_87_n462), .ZN(
        u5_mult_87_ab_28__27_) );
  NOR2_X1 u5_mult_87_U2212 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n462), .ZN(
        u5_mult_87_ab_28__28_) );
  NOR2_X1 u5_mult_87_U2211 ( .A1(u5_mult_87_n390), .A2(u5_mult_87_n462), .ZN(
        u5_mult_87_ab_28__29_) );
  NOR2_X1 u5_mult_87_U2210 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n275), .ZN(
        u5_mult_87_ab_28__2_) );
  NOR2_X1 u5_mult_87_U2209 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n275), .ZN(
        u5_mult_87_ab_28__30_) );
  NOR2_X1 u5_mult_87_U2208 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n275), .ZN(
        u5_mult_87_ab_28__31_) );
  NOR2_X1 u5_mult_87_U2207 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n275), .ZN(
        u5_mult_87_ab_28__32_) );
  NOR2_X1 u5_mult_87_U2206 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n275), .ZN(
        u5_mult_87_ab_28__33_) );
  NOR2_X1 u5_mult_87_U2205 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n275), .ZN(
        u5_mult_87_ab_28__34_) );
  NOR2_X1 u5_mult_87_U2204 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n275), .ZN(
        u5_mult_87_ab_28__35_) );
  NOR2_X1 u5_mult_87_U2203 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n275), .ZN(
        u5_mult_87_ab_28__36_) );
  NOR2_X1 u5_mult_87_U2202 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n275), .ZN(
        u5_mult_87_ab_28__37_) );
  NOR2_X1 u5_mult_87_U2201 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n275), .ZN(
        u5_mult_87_ab_28__38_) );
  NOR2_X1 u5_mult_87_U2200 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n275), .ZN(
        u5_mult_87_ab_28__39_) );
  NOR2_X1 u5_mult_87_U2199 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__3_) );
  NOR2_X1 u5_mult_87_U2198 ( .A1(u5_mult_87_n367), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__40_) );
  NOR2_X1 u5_mult_87_U2197 ( .A1(u5_mult_87_n365), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__41_) );
  NOR2_X1 u5_mult_87_U2196 ( .A1(u5_mult_87_n364), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__42_) );
  NOR2_X1 u5_mult_87_U2195 ( .A1(u5_mult_87_n360), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__43_) );
  NOR2_X1 u5_mult_87_U2194 ( .A1(u5_mult_87_n358), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__44_) );
  NOR2_X1 u5_mult_87_U2193 ( .A1(u5_mult_87_n356), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__45_) );
  NOR2_X1 u5_mult_87_U2192 ( .A1(u5_mult_87_n354), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__46_) );
  NOR2_X1 u5_mult_87_U2191 ( .A1(u5_mult_87_n351), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__47_) );
  NOR2_X1 u5_mult_87_U2190 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__48_) );
  NOR2_X1 u5_mult_87_U2189 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__49_) );
  NOR2_X1 u5_mult_87_U2188 ( .A1(u5_mult_87_n440), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__4_) );
  NOR2_X1 u5_mult_87_U2187 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__50_) );
  NOR2_X1 u5_mult_87_U2186 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__51_) );
  NOR2_X1 u5_mult_87_U2185 ( .A1(u5_mult_87_n342), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__52_) );
  NOR2_X1 u5_mult_87_U2184 ( .A1(u5_mult_87_n437), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__5_) );
  NOR2_X1 u5_mult_87_U2183 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__6_) );
  NOR2_X1 u5_mult_87_U2182 ( .A1(u5_mult_87_n434), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__7_) );
  NOR2_X1 u5_mult_87_U2181 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__8_) );
  NOR2_X1 u5_mult_87_U2180 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n276), .ZN(
        u5_mult_87_ab_28__9_) );
  NOR2_X1 u5_mult_87_U2179 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n273), .ZN(
        u5_mult_87_ab_29__0_) );
  NOR2_X1 u5_mult_87_U2178 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n273), .ZN(
        u5_mult_87_ab_29__10_) );
  NOR2_X1 u5_mult_87_U2177 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__11_) );
  NOR2_X1 u5_mult_87_U2176 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n273), .ZN(
        u5_mult_87_ab_29__12_) );
  NOR2_X1 u5_mult_87_U2175 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n273), .ZN(
        u5_mult_87_ab_29__13_) );
  NOR2_X1 u5_mult_87_U2174 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__14_) );
  NOR2_X1 u5_mult_87_U2173 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__15_) );
  NOR2_X1 u5_mult_87_U2172 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__16_) );
  NOR2_X1 u5_mult_87_U2171 ( .A1(u5_mult_87_n413), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__17_) );
  NOR2_X1 u5_mult_87_U2170 ( .A1(u5_mult_87_n411), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__18_) );
  NOR2_X1 u5_mult_87_U2169 ( .A1(u5_mult_87_n409), .A2(u5_mult_87_n273), .ZN(
        u5_mult_87_ab_29__19_) );
  NOR2_X1 u5_mult_87_U2168 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n461), .ZN(
        u5_mult_87_ab_29__1_) );
  NOR2_X1 u5_mult_87_U2167 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n461), .ZN(
        u5_mult_87_ab_29__20_) );
  NOR2_X1 u5_mult_87_U2166 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n461), .ZN(
        u5_mult_87_ab_29__21_) );
  NOR2_X1 u5_mult_87_U2165 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n461), .ZN(
        u5_mult_87_ab_29__22_) );
  NOR2_X1 u5_mult_87_U2164 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n461), .ZN(
        u5_mult_87_ab_29__23_) );
  NOR2_X1 u5_mult_87_U2163 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n461), .ZN(
        u5_mult_87_ab_29__24_) );
  NOR2_X1 u5_mult_87_U2162 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n461), .ZN(
        u5_mult_87_ab_29__25_) );
  NOR2_X1 u5_mult_87_U2161 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n461), .ZN(
        u5_mult_87_ab_29__26_) );
  NOR2_X1 u5_mult_87_U2160 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n461), .ZN(
        u5_mult_87_ab_29__27_) );
  NOR2_X1 u5_mult_87_U2159 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n461), .ZN(
        u5_mult_87_ab_29__28_) );
  NOR2_X1 u5_mult_87_U2158 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n461), .ZN(
        u5_mult_87_ab_29__29_) );
  NOR2_X1 u5_mult_87_U2157 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n273), .ZN(
        u5_mult_87_ab_29__2_) );
  NOR2_X1 u5_mult_87_U2156 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n273), .ZN(
        u5_mult_87_ab_29__30_) );
  NOR2_X1 u5_mult_87_U2155 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n273), .ZN(
        u5_mult_87_ab_29__31_) );
  NOR2_X1 u5_mult_87_U2154 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n273), .ZN(
        u5_mult_87_ab_29__32_) );
  NOR2_X1 u5_mult_87_U2153 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n273), .ZN(
        u5_mult_87_ab_29__33_) );
  NOR2_X1 u5_mult_87_U2152 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n273), .ZN(
        u5_mult_87_ab_29__34_) );
  NOR2_X1 u5_mult_87_U2151 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n273), .ZN(
        u5_mult_87_ab_29__35_) );
  NOR2_X1 u5_mult_87_U2150 ( .A1(u5_mult_87_n376), .A2(u5_mult_87_n273), .ZN(
        u5_mult_87_ab_29__36_) );
  NOR2_X1 u5_mult_87_U2149 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n273), .ZN(
        u5_mult_87_ab_29__37_) );
  NOR2_X1 u5_mult_87_U2148 ( .A1(u5_mult_87_n372), .A2(u5_mult_87_n273), .ZN(
        u5_mult_87_ab_29__38_) );
  NOR2_X1 u5_mult_87_U2147 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n273), .ZN(
        u5_mult_87_ab_29__39_) );
  NOR2_X1 u5_mult_87_U2146 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__3_) );
  NOR2_X1 u5_mult_87_U2145 ( .A1(u5_mult_87_n367), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__40_) );
  NOR2_X1 u5_mult_87_U2144 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__41_) );
  NOR2_X1 u5_mult_87_U2143 ( .A1(u5_mult_87_n364), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__42_) );
  NOR2_X1 u5_mult_87_U2142 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__43_) );
  NOR2_X1 u5_mult_87_U2141 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__44_) );
  NOR2_X1 u5_mult_87_U2140 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__45_) );
  NOR2_X1 u5_mult_87_U2139 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__46_) );
  NOR2_X1 u5_mult_87_U2138 ( .A1(u5_mult_87_n351), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__47_) );
  NOR2_X1 u5_mult_87_U2137 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__48_) );
  NOR2_X1 u5_mult_87_U2136 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__49_) );
  NOR2_X1 u5_mult_87_U2135 ( .A1(u5_mult_87_n440), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__4_) );
  NOR2_X1 u5_mult_87_U2134 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__50_) );
  NOR2_X1 u5_mult_87_U2133 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__51_) );
  NOR2_X1 u5_mult_87_U2132 ( .A1(u5_mult_87_n342), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__52_) );
  NOR2_X1 u5_mult_87_U2131 ( .A1(u5_mult_87_n437), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__5_) );
  NOR2_X1 u5_mult_87_U2130 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__6_) );
  NOR2_X1 u5_mult_87_U2129 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__7_) );
  NOR2_X1 u5_mult_87_U2128 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__8_) );
  NOR2_X1 u5_mult_87_U2127 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n274), .ZN(
        u5_mult_87_ab_29__9_) );
  NOR2_X1 u5_mult_87_U2126 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__0_) );
  NOR2_X1 u5_mult_87_U2125 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__10_) );
  NOR2_X1 u5_mult_87_U2124 ( .A1(u5_mult_87_n425), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__11_) );
  NOR2_X1 u5_mult_87_U2123 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__12_) );
  NOR2_X1 u5_mult_87_U2122 ( .A1(u5_mult_87_n422), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__13_) );
  NOR2_X1 u5_mult_87_U2121 ( .A1(u5_mult_87_n418), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__14_) );
  NOR2_X1 u5_mult_87_U2120 ( .A1(u5_mult_87_n416), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__15_) );
  NOR2_X1 u5_mult_87_U2119 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__16_) );
  NOR2_X1 u5_mult_87_U2118 ( .A1(u5_mult_87_n413), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__17_) );
  NOR2_X1 u5_mult_87_U2117 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__18_) );
  NOR2_X1 u5_mult_87_U2116 ( .A1(u5_mult_87_n409), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__19_) );
  NOR2_X1 u5_mult_87_U2115 ( .A1(u5_mult_87_n447), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__1_) );
  NOR2_X1 u5_mult_87_U2114 ( .A1(u5_mult_87_n407), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__20_) );
  NOR2_X1 u5_mult_87_U2113 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__21_) );
  NOR2_X1 u5_mult_87_U2112 ( .A1(u5_mult_87_n404), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__22_) );
  NOR2_X1 u5_mult_87_U2111 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__23_) );
  NOR2_X1 u5_mult_87_U2110 ( .A1(u5_mult_87_n399), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__24_) );
  NOR2_X1 u5_mult_87_U2109 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__25_) );
  NOR2_X1 u5_mult_87_U2108 ( .A1(u5_mult_87_n395), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__26_) );
  NOR2_X1 u5_mult_87_U2107 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__27_) );
  NOR2_X1 u5_mult_87_U2106 ( .A1(u5_mult_87_n392), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__28_) );
  NOR2_X1 u5_mult_87_U2105 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__29_) );
  NOR2_X1 u5_mult_87_U2104 ( .A1(u5_mult_87_n444), .A2(u5_mult_87_n333), .ZN(
        u5_mult_87_ab_2__2_) );
  NOR2_X1 u5_mult_87_U2103 ( .A1(u5_mult_87_n387), .A2(u5_mult_87_n333), .ZN(
        u5_mult_87_ab_2__30_) );
  NOR2_X1 u5_mult_87_U2102 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n333), .ZN(
        u5_mult_87_ab_2__31_) );
  NOR2_X1 u5_mult_87_U2101 ( .A1(u5_mult_87_n383), .A2(u5_mult_87_n333), .ZN(
        u5_mult_87_ab_2__32_) );
  NOR2_X1 u5_mult_87_U2100 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n333), .ZN(
        u5_mult_87_ab_2__33_) );
  NOR2_X1 u5_mult_87_U2099 ( .A1(u5_mult_87_n379), .A2(u5_mult_87_n333), .ZN(
        u5_mult_87_ab_2__34_) );
  NOR2_X1 u5_mult_87_U2098 ( .A1(u5_mult_87_n377), .A2(u5_mult_87_n333), .ZN(
        u5_mult_87_ab_2__35_) );
  NOR2_X1 u5_mult_87_U2097 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n333), .ZN(
        u5_mult_87_ab_2__36_) );
  NOR2_X1 u5_mult_87_U2096 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n333), .ZN(
        u5_mult_87_ab_2__37_) );
  NOR2_X1 u5_mult_87_U2095 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n333), .ZN(
        u5_mult_87_ab_2__38_) );
  NOR2_X1 u5_mult_87_U2094 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n333), .ZN(
        u5_mult_87_ab_2__39_) );
  NOR2_X1 u5_mult_87_U2093 ( .A1(u5_mult_87_n442), .A2(u5_mult_87_n334), .ZN(
        u5_mult_87_ab_2__3_) );
  NOR2_X1 u5_mult_87_U2092 ( .A1(u5_mult_87_n367), .A2(u5_mult_87_n334), .ZN(
        u5_mult_87_ab_2__40_) );
  NOR2_X1 u5_mult_87_U2091 ( .A1(u5_mult_87_n365), .A2(u5_mult_87_n334), .ZN(
        u5_mult_87_ab_2__41_) );
  NOR2_X1 u5_mult_87_U2090 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n334), .ZN(
        u5_mult_87_ab_2__42_) );
  NOR2_X1 u5_mult_87_U2089 ( .A1(u5_mult_87_n360), .A2(u5_mult_87_n334), .ZN(
        u5_mult_87_ab_2__43_) );
  NOR2_X1 u5_mult_87_U2088 ( .A1(u5_mult_87_n358), .A2(u5_mult_87_n334), .ZN(
        u5_mult_87_ab_2__44_) );
  NOR2_X1 u5_mult_87_U2087 ( .A1(u5_mult_87_n356), .A2(u5_mult_87_n334), .ZN(
        u5_mult_87_ab_2__45_) );
  NOR2_X1 u5_mult_87_U2086 ( .A1(u5_mult_87_n354), .A2(u5_mult_87_n334), .ZN(
        u5_mult_87_ab_2__46_) );
  NOR2_X1 u5_mult_87_U2085 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n334), .ZN(
        u5_mult_87_ab_2__47_) );
  NOR2_X1 u5_mult_87_U2084 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n334), .ZN(
        u5_mult_87_ab_2__48_) );
  NOR2_X1 u5_mult_87_U2083 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n334), .ZN(
        u5_mult_87_ab_2__49_) );
  NOR2_X1 u5_mult_87_U2082 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__4_) );
  NOR2_X1 u5_mult_87_U2081 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n334), .ZN(
        u5_mult_87_ab_2__50_) );
  NOR2_X1 u5_mult_87_U2080 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n335), .ZN(
        u5_mult_87_ab_2__51_) );
  NOR2_X1 u5_mult_87_U2079 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n333), .ZN(
        u5_mult_87_ab_2__52_) );
  NOR2_X1 u5_mult_87_U2078 ( .A1(u5_mult_87_n439), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__5_) );
  NOR2_X1 u5_mult_87_U2077 ( .A1(u5_mult_87_n436), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__6_) );
  NOR2_X1 u5_mult_87_U2076 ( .A1(u5_mult_87_n434), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__7_) );
  NOR2_X1 u5_mult_87_U2075 ( .A1(u5_mult_87_n432), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__8_) );
  NOR2_X1 u5_mult_87_U2074 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n332), .ZN(
        u5_mult_87_ab_2__9_) );
  NOR2_X1 u5_mult_87_U2073 ( .A1(u5_mult_87_n450), .A2(u5_mult_87_n270), .ZN(
        u5_mult_87_ab_30__0_) );
  NOR2_X1 u5_mult_87_U2072 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n270), .ZN(
        u5_mult_87_ab_30__10_) );
  NOR2_X1 u5_mult_87_U2071 ( .A1(u5_mult_87_n425), .A2(u5_mult_87_n270), .ZN(
        u5_mult_87_ab_30__11_) );
  NOR2_X1 u5_mult_87_U2070 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n270), .ZN(
        u5_mult_87_ab_30__12_) );
  NOR2_X1 u5_mult_87_U2069 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__13_) );
  NOR2_X1 u5_mult_87_U2068 ( .A1(u5_mult_87_n418), .A2(u5_mult_87_n270), .ZN(
        u5_mult_87_ab_30__14_) );
  NOR2_X1 u5_mult_87_U2067 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n270), .ZN(
        u5_mult_87_ab_30__15_) );
  NOR2_X1 u5_mult_87_U2066 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n270), .ZN(
        u5_mult_87_ab_30__16_) );
  NOR2_X1 u5_mult_87_U2065 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__17_) );
  NOR2_X1 u5_mult_87_U2064 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n270), .ZN(
        u5_mult_87_ab_30__18_) );
  NOR2_X1 u5_mult_87_U2063 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n270), .ZN(
        u5_mult_87_ab_30__19_) );
  NOR2_X1 u5_mult_87_U2062 ( .A1(u5_mult_87_n447), .A2(u5_mult_87_n272), .ZN(
        u5_mult_87_ab_30__1_) );
  NOR2_X1 u5_mult_87_U2061 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n272), .ZN(
        u5_mult_87_ab_30__20_) );
  NOR2_X1 u5_mult_87_U2060 ( .A1(u5_mult_87_n406), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__21_) );
  NOR2_X1 u5_mult_87_U2059 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n272), .ZN(
        u5_mult_87_ab_30__22_) );
  NOR2_X1 u5_mult_87_U2058 ( .A1(u5_mult_87_n402), .A2(u5_mult_87_n272), .ZN(
        u5_mult_87_ab_30__23_) );
  NOR2_X1 u5_mult_87_U2057 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n272), .ZN(
        u5_mult_87_ab_30__24_) );
  NOR2_X1 u5_mult_87_U2056 ( .A1(u5_mult_87_n398), .A2(u5_mult_87_n272), .ZN(
        u5_mult_87_ab_30__25_) );
  NOR2_X1 u5_mult_87_U2055 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n272), .ZN(
        u5_mult_87_ab_30__26_) );
  NOR2_X1 u5_mult_87_U2054 ( .A1(u5_mult_87_n394), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__27_) );
  NOR2_X1 u5_mult_87_U2053 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n272), .ZN(
        u5_mult_87_ab_30__28_) );
  NOR2_X1 u5_mult_87_U2052 ( .A1(u5_mult_87_n390), .A2(u5_mult_87_n272), .ZN(
        u5_mult_87_ab_30__29_) );
  NOR2_X1 u5_mult_87_U2051 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n270), .ZN(
        u5_mult_87_ab_30__2_) );
  NOR2_X1 u5_mult_87_U2050 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n270), .ZN(
        u5_mult_87_ab_30__30_) );
  NOR2_X1 u5_mult_87_U2049 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n270), .ZN(
        u5_mult_87_ab_30__31_) );
  NOR2_X1 u5_mult_87_U2048 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n270), .ZN(
        u5_mult_87_ab_30__32_) );
  NOR2_X1 u5_mult_87_U2047 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n270), .ZN(
        u5_mult_87_ab_30__33_) );
  NOR2_X1 u5_mult_87_U2046 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n270), .ZN(
        u5_mult_87_ab_30__34_) );
  NOR2_X1 u5_mult_87_U2045 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n270), .ZN(
        u5_mult_87_ab_30__35_) );
  NOR2_X1 u5_mult_87_U2044 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n270), .ZN(
        u5_mult_87_ab_30__36_) );
  NOR2_X1 u5_mult_87_U2043 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n270), .ZN(
        u5_mult_87_ab_30__37_) );
  NOR2_X1 u5_mult_87_U2042 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n270), .ZN(
        u5_mult_87_ab_30__38_) );
  NOR2_X1 u5_mult_87_U2041 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n270), .ZN(
        u5_mult_87_ab_30__39_) );
  NOR2_X1 u5_mult_87_U2040 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__3_) );
  NOR2_X1 u5_mult_87_U2039 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__40_) );
  NOR2_X1 u5_mult_87_U2038 ( .A1(u5_mult_87_n365), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__41_) );
  NOR2_X1 u5_mult_87_U2037 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__42_) );
  NOR2_X1 u5_mult_87_U2036 ( .A1(u5_mult_87_n360), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__43_) );
  NOR2_X1 u5_mult_87_U2035 ( .A1(u5_mult_87_n358), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__44_) );
  NOR2_X1 u5_mult_87_U2034 ( .A1(u5_mult_87_n356), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__45_) );
  NOR2_X1 u5_mult_87_U2033 ( .A1(u5_mult_87_n354), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__46_) );
  NOR2_X1 u5_mult_87_U2032 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__47_) );
  NOR2_X1 u5_mult_87_U2031 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__48_) );
  NOR2_X1 u5_mult_87_U2030 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__49_) );
  NOR2_X1 u5_mult_87_U2029 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__4_) );
  NOR2_X1 u5_mult_87_U2028 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__50_) );
  NOR2_X1 u5_mult_87_U2027 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__51_) );
  NOR2_X1 u5_mult_87_U2026 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__52_) );
  NOR2_X1 u5_mult_87_U2025 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__5_) );
  NOR2_X1 u5_mult_87_U2024 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__6_) );
  NOR2_X1 u5_mult_87_U2023 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__7_) );
  NOR2_X1 u5_mult_87_U2022 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__8_) );
  NOR2_X1 u5_mult_87_U2021 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n271), .ZN(
        u5_mult_87_ab_30__9_) );
  NOR2_X1 u5_mult_87_U2020 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n268), .ZN(
        u5_mult_87_ab_31__0_) );
  NOR2_X1 u5_mult_87_U2019 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n268), .ZN(
        u5_mult_87_ab_31__10_) );
  NOR2_X1 u5_mult_87_U2018 ( .A1(u5_mult_87_n425), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__11_) );
  NOR2_X1 u5_mult_87_U2017 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n268), .ZN(
        u5_mult_87_ab_31__12_) );
  NOR2_X1 u5_mult_87_U2016 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n268), .ZN(
        u5_mult_87_ab_31__13_) );
  NOR2_X1 u5_mult_87_U2015 ( .A1(u5_mult_87_n418), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__14_) );
  NOR2_X1 u5_mult_87_U2014 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__15_) );
  NOR2_X1 u5_mult_87_U2013 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__16_) );
  NOR2_X1 u5_mult_87_U2012 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n268), .ZN(
        u5_mult_87_ab_31__17_) );
  NOR2_X1 u5_mult_87_U2011 ( .A1(u5_mult_87_n411), .A2(u5_mult_87_n268), .ZN(
        u5_mult_87_ab_31__18_) );
  NOR2_X1 u5_mult_87_U2010 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n268), .ZN(
        u5_mult_87_ab_31__19_) );
  NOR2_X1 u5_mult_87_U2009 ( .A1(u5_mult_87_n447), .A2(u5_mult_87_n460), .ZN(
        u5_mult_87_ab_31__1_) );
  NOR2_X1 u5_mult_87_U2008 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n460), .ZN(
        u5_mult_87_ab_31__20_) );
  NOR2_X1 u5_mult_87_U2007 ( .A1(u5_mult_87_n406), .A2(u5_mult_87_n460), .ZN(
        u5_mult_87_ab_31__21_) );
  NOR2_X1 u5_mult_87_U2006 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n460), .ZN(
        u5_mult_87_ab_31__22_) );
  NOR2_X1 u5_mult_87_U2005 ( .A1(u5_mult_87_n402), .A2(u5_mult_87_n460), .ZN(
        u5_mult_87_ab_31__23_) );
  NOR2_X1 u5_mult_87_U2004 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n460), .ZN(
        u5_mult_87_ab_31__24_) );
  NOR2_X1 u5_mult_87_U2003 ( .A1(u5_mult_87_n398), .A2(u5_mult_87_n460), .ZN(
        u5_mult_87_ab_31__25_) );
  NOR2_X1 u5_mult_87_U2002 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n460), .ZN(
        u5_mult_87_ab_31__26_) );
  NOR2_X1 u5_mult_87_U2001 ( .A1(u5_mult_87_n394), .A2(u5_mult_87_n460), .ZN(
        u5_mult_87_ab_31__27_) );
  NOR2_X1 u5_mult_87_U2000 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n460), .ZN(
        u5_mult_87_ab_31__28_) );
  NOR2_X1 u5_mult_87_U1999 ( .A1(u5_mult_87_n390), .A2(u5_mult_87_n460), .ZN(
        u5_mult_87_ab_31__29_) );
  NOR2_X1 u5_mult_87_U1998 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n268), .ZN(
        u5_mult_87_ab_31__2_) );
  NOR2_X1 u5_mult_87_U1997 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n268), .ZN(
        u5_mult_87_ab_31__30_) );
  NOR2_X1 u5_mult_87_U1996 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n268), .ZN(
        u5_mult_87_ab_31__31_) );
  NOR2_X1 u5_mult_87_U1995 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n268), .ZN(
        u5_mult_87_ab_31__32_) );
  NOR2_X1 u5_mult_87_U1994 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n268), .ZN(
        u5_mult_87_ab_31__33_) );
  NOR2_X1 u5_mult_87_U1993 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n268), .ZN(
        u5_mult_87_ab_31__34_) );
  NOR2_X1 u5_mult_87_U1992 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n268), .ZN(
        u5_mult_87_ab_31__35_) );
  NOR2_X1 u5_mult_87_U1991 ( .A1(u5_mult_87_n376), .A2(u5_mult_87_n268), .ZN(
        u5_mult_87_ab_31__36_) );
  NOR2_X1 u5_mult_87_U1990 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n268), .ZN(
        u5_mult_87_ab_31__37_) );
  NOR2_X1 u5_mult_87_U1989 ( .A1(u5_mult_87_n372), .A2(u5_mult_87_n268), .ZN(
        u5_mult_87_ab_31__38_) );
  NOR2_X1 u5_mult_87_U1988 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n268), .ZN(
        u5_mult_87_ab_31__39_) );
  NOR2_X1 u5_mult_87_U1987 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__3_) );
  NOR2_X1 u5_mult_87_U1986 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__40_) );
  NOR2_X1 u5_mult_87_U1985 ( .A1(u5_mult_87_n365), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__41_) );
  NOR2_X1 u5_mult_87_U1984 ( .A1(u5_mult_87_n363), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__42_) );
  NOR2_X1 u5_mult_87_U1983 ( .A1(u5_mult_87_n360), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__43_) );
  NOR2_X1 u5_mult_87_U1982 ( .A1(u5_mult_87_n358), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__44_) );
  NOR2_X1 u5_mult_87_U1981 ( .A1(u5_mult_87_n356), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__45_) );
  NOR2_X1 u5_mult_87_U1980 ( .A1(u5_mult_87_n354), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__46_) );
  NOR2_X1 u5_mult_87_U1979 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__47_) );
  NOR2_X1 u5_mult_87_U1978 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__48_) );
  NOR2_X1 u5_mult_87_U1977 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__49_) );
  NOR2_X1 u5_mult_87_U1976 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__4_) );
  NOR2_X1 u5_mult_87_U1975 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__50_) );
  NOR2_X1 u5_mult_87_U1974 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__51_) );
  NOR2_X1 u5_mult_87_U1973 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__52_) );
  NOR2_X1 u5_mult_87_U1972 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__5_) );
  NOR2_X1 u5_mult_87_U1971 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__6_) );
  NOR2_X1 u5_mult_87_U1970 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__7_) );
  NOR2_X1 u5_mult_87_U1969 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__8_) );
  NOR2_X1 u5_mult_87_U1968 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n269), .ZN(
        u5_mult_87_ab_31__9_) );
  NOR2_X1 u5_mult_87_U1967 ( .A1(u5_mult_87_n450), .A2(u5_mult_87_n265), .ZN(
        u5_mult_87_ab_32__0_) );
  NOR2_X1 u5_mult_87_U1966 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n265), .ZN(
        u5_mult_87_ab_32__10_) );
  NOR2_X1 u5_mult_87_U1965 ( .A1(u5_mult_87_n425), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__11_) );
  NOR2_X1 u5_mult_87_U1964 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n265), .ZN(
        u5_mult_87_ab_32__12_) );
  NOR2_X1 u5_mult_87_U1963 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n265), .ZN(
        u5_mult_87_ab_32__13_) );
  NOR2_X1 u5_mult_87_U1962 ( .A1(u5_mult_87_n418), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__14_) );
  NOR2_X1 u5_mult_87_U1961 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__15_) );
  NOR2_X1 u5_mult_87_U1960 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__16_) );
  NOR2_X1 u5_mult_87_U1959 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n265), .ZN(
        u5_mult_87_ab_32__17_) );
  NOR2_X1 u5_mult_87_U1958 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n265), .ZN(
        u5_mult_87_ab_32__18_) );
  NOR2_X1 u5_mult_87_U1957 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n265), .ZN(
        u5_mult_87_ab_32__19_) );
  NOR2_X1 u5_mult_87_U1956 ( .A1(u5_mult_87_n447), .A2(u5_mult_87_n267), .ZN(
        u5_mult_87_ab_32__1_) );
  NOR2_X1 u5_mult_87_U1955 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n267), .ZN(
        u5_mult_87_ab_32__20_) );
  NOR2_X1 u5_mult_87_U1954 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n267), .ZN(
        u5_mult_87_ab_32__21_) );
  NOR2_X1 u5_mult_87_U1953 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n267), .ZN(
        u5_mult_87_ab_32__22_) );
  NOR2_X1 u5_mult_87_U1952 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n267), .ZN(
        u5_mult_87_ab_32__23_) );
  NOR2_X1 u5_mult_87_U1951 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n267), .ZN(
        u5_mult_87_ab_32__24_) );
  NOR2_X1 u5_mult_87_U1950 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__25_) );
  NOR2_X1 u5_mult_87_U1949 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n267), .ZN(
        u5_mult_87_ab_32__26_) );
  NOR2_X1 u5_mult_87_U1948 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n267), .ZN(
        u5_mult_87_ab_32__27_) );
  NOR2_X1 u5_mult_87_U1947 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n267), .ZN(
        u5_mult_87_ab_32__28_) );
  NOR2_X1 u5_mult_87_U1946 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n267), .ZN(
        u5_mult_87_ab_32__29_) );
  NOR2_X1 u5_mult_87_U1945 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n265), .ZN(
        u5_mult_87_ab_32__2_) );
  NOR2_X1 u5_mult_87_U1944 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n265), .ZN(
        u5_mult_87_ab_32__30_) );
  NOR2_X1 u5_mult_87_U1943 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n265), .ZN(
        u5_mult_87_ab_32__31_) );
  NOR2_X1 u5_mult_87_U1942 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n265), .ZN(
        u5_mult_87_ab_32__32_) );
  NOR2_X1 u5_mult_87_U1941 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n265), .ZN(
        u5_mult_87_ab_32__33_) );
  NOR2_X1 u5_mult_87_U1940 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n265), .ZN(
        u5_mult_87_ab_32__34_) );
  NOR2_X1 u5_mult_87_U1939 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n265), .ZN(
        u5_mult_87_ab_32__35_) );
  NOR2_X1 u5_mult_87_U1938 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n265), .ZN(
        u5_mult_87_ab_32__36_) );
  NOR2_X1 u5_mult_87_U1937 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n265), .ZN(
        u5_mult_87_ab_32__37_) );
  NOR2_X1 u5_mult_87_U1936 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n265), .ZN(
        u5_mult_87_ab_32__38_) );
  NOR2_X1 u5_mult_87_U1935 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n265), .ZN(
        u5_mult_87_ab_32__39_) );
  NOR2_X1 u5_mult_87_U1934 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__3_) );
  NOR2_X1 u5_mult_87_U1933 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__40_) );
  NOR2_X1 u5_mult_87_U1932 ( .A1(u5_mult_87_n365), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__41_) );
  NOR2_X1 u5_mult_87_U1931 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__42_) );
  NOR2_X1 u5_mult_87_U1930 ( .A1(u5_mult_87_n360), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__43_) );
  NOR2_X1 u5_mult_87_U1929 ( .A1(u5_mult_87_n358), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__44_) );
  NOR2_X1 u5_mult_87_U1928 ( .A1(u5_mult_87_n356), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__45_) );
  NOR2_X1 u5_mult_87_U1927 ( .A1(u5_mult_87_n354), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__46_) );
  NOR2_X1 u5_mult_87_U1926 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__47_) );
  NOR2_X1 u5_mult_87_U1925 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__48_) );
  NOR2_X1 u5_mult_87_U1924 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__49_) );
  NOR2_X1 u5_mult_87_U1923 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__4_) );
  NOR2_X1 u5_mult_87_U1922 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__50_) );
  NOR2_X1 u5_mult_87_U1921 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__51_) );
  NOR2_X1 u5_mult_87_U1920 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__52_) );
  NOR2_X1 u5_mult_87_U1919 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__5_) );
  NOR2_X1 u5_mult_87_U1918 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__6_) );
  NOR2_X1 u5_mult_87_U1917 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__7_) );
  NOR2_X1 u5_mult_87_U1916 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__8_) );
  NOR2_X1 u5_mult_87_U1915 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n266), .ZN(
        u5_mult_87_ab_32__9_) );
  NOR2_X1 u5_mult_87_U1914 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n264), .ZN(
        u5_mult_87_ab_33__0_) );
  NOR2_X1 u5_mult_87_U1913 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n264), .ZN(
        u5_mult_87_ab_33__10_) );
  NOR2_X1 u5_mult_87_U1912 ( .A1(u5_mult_87_n425), .A2(u5_mult_87_n264), .ZN(
        u5_mult_87_ab_33__11_) );
  NOR2_X1 u5_mult_87_U1911 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n264), .ZN(
        u5_mult_87_ab_33__12_) );
  NOR2_X1 u5_mult_87_U1910 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__13_) );
  NOR2_X1 u5_mult_87_U1909 ( .A1(u5_mult_87_n418), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__14_) );
  NOR2_X1 u5_mult_87_U1908 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__15_) );
  NOR2_X1 u5_mult_87_U1907 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n264), .ZN(
        u5_mult_87_ab_33__16_) );
  NOR2_X1 u5_mult_87_U1906 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n264), .ZN(
        u5_mult_87_ab_33__17_) );
  NOR2_X1 u5_mult_87_U1905 ( .A1(u5_mult_87_n411), .A2(u5_mult_87_n264), .ZN(
        u5_mult_87_ab_33__18_) );
  NOR2_X1 u5_mult_87_U1904 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n264), .ZN(
        u5_mult_87_ab_33__19_) );
  NOR2_X1 u5_mult_87_U1903 ( .A1(u5_mult_87_n447), .A2(u5_mult_87_n459), .ZN(
        u5_mult_87_ab_33__1_) );
  NOR2_X1 u5_mult_87_U1902 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n264), .ZN(
        u5_mult_87_ab_33__20_) );
  NOR2_X1 u5_mult_87_U1901 ( .A1(u5_mult_87_n406), .A2(u5_mult_87_n264), .ZN(
        u5_mult_87_ab_33__21_) );
  NOR2_X1 u5_mult_87_U1900 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n264), .ZN(
        u5_mult_87_ab_33__22_) );
  NOR2_X1 u5_mult_87_U1899 ( .A1(u5_mult_87_n402), .A2(u5_mult_87_n459), .ZN(
        u5_mult_87_ab_33__23_) );
  NOR2_X1 u5_mult_87_U1898 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n459), .ZN(
        u5_mult_87_ab_33__24_) );
  NOR2_X1 u5_mult_87_U1897 ( .A1(u5_mult_87_n398), .A2(u5_mult_87_n459), .ZN(
        u5_mult_87_ab_33__25_) );
  NOR2_X1 u5_mult_87_U1896 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n459), .ZN(
        u5_mult_87_ab_33__26_) );
  NOR2_X1 u5_mult_87_U1895 ( .A1(u5_mult_87_n394), .A2(u5_mult_87_n459), .ZN(
        u5_mult_87_ab_33__27_) );
  NOR2_X1 u5_mult_87_U1894 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n459), .ZN(
        u5_mult_87_ab_33__28_) );
  NOR2_X1 u5_mult_87_U1893 ( .A1(u5_mult_87_n390), .A2(u5_mult_87_n459), .ZN(
        u5_mult_87_ab_33__29_) );
  NOR2_X1 u5_mult_87_U1892 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__2_) );
  NOR2_X1 u5_mult_87_U1891 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__30_) );
  NOR2_X1 u5_mult_87_U1890 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__31_) );
  NOR2_X1 u5_mult_87_U1889 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__32_) );
  NOR2_X1 u5_mult_87_U1888 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__33_) );
  NOR2_X1 u5_mult_87_U1887 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__34_) );
  NOR2_X1 u5_mult_87_U1886 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__35_) );
  NOR2_X1 u5_mult_87_U1885 ( .A1(u5_mult_87_n376), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__36_) );
  NOR2_X1 u5_mult_87_U1884 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__37_) );
  NOR2_X1 u5_mult_87_U1883 ( .A1(u5_mult_87_n372), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__38_) );
  NOR2_X1 u5_mult_87_U1882 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__39_) );
  NOR2_X1 u5_mult_87_U1881 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__3_) );
  NOR2_X1 u5_mult_87_U1880 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__40_) );
  NOR2_X1 u5_mult_87_U1879 ( .A1(u5_mult_87_n365), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__41_) );
  NOR2_X1 u5_mult_87_U1878 ( .A1(u5_mult_87_n363), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__42_) );
  NOR2_X1 u5_mult_87_U1877 ( .A1(u5_mult_87_n360), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__43_) );
  NOR2_X1 u5_mult_87_U1876 ( .A1(u5_mult_87_n358), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__44_) );
  NOR2_X1 u5_mult_87_U1875 ( .A1(u5_mult_87_n356), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__45_) );
  NOR2_X1 u5_mult_87_U1874 ( .A1(u5_mult_87_n354), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__46_) );
  NOR2_X1 u5_mult_87_U1873 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__47_) );
  NOR2_X1 u5_mult_87_U1872 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__48_) );
  NOR2_X1 u5_mult_87_U1871 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__49_) );
  NOR2_X1 u5_mult_87_U1870 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__4_) );
  NOR2_X1 u5_mult_87_U1869 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__50_) );
  NOR2_X1 u5_mult_87_U1868 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__51_) );
  NOR2_X1 u5_mult_87_U1867 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__52_) );
  NOR2_X1 u5_mult_87_U1866 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__5_) );
  NOR2_X1 u5_mult_87_U1865 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__6_) );
  NOR2_X1 u5_mult_87_U1864 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__7_) );
  NOR2_X1 u5_mult_87_U1863 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__8_) );
  NOR2_X1 u5_mult_87_U1862 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n263), .ZN(
        u5_mult_87_ab_33__9_) );
  NOR2_X1 u5_mult_87_U1861 ( .A1(u5_mult_87_n450), .A2(u5_mult_87_n261), .ZN(
        u5_mult_87_ab_34__0_) );
  NOR2_X1 u5_mult_87_U1860 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n261), .ZN(
        u5_mult_87_ab_34__10_) );
  NOR2_X1 u5_mult_87_U1859 ( .A1(u5_mult_87_n425), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__11_) );
  NOR2_X1 u5_mult_87_U1858 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n261), .ZN(
        u5_mult_87_ab_34__12_) );
  NOR2_X1 u5_mult_87_U1857 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__13_) );
  NOR2_X1 u5_mult_87_U1856 ( .A1(u5_mult_87_n418), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__14_) );
  NOR2_X1 u5_mult_87_U1855 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__15_) );
  NOR2_X1 u5_mult_87_U1854 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n261), .ZN(
        u5_mult_87_ab_34__16_) );
  NOR2_X1 u5_mult_87_U1853 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n261), .ZN(
        u5_mult_87_ab_34__17_) );
  NOR2_X1 u5_mult_87_U1852 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n261), .ZN(
        u5_mult_87_ab_34__18_) );
  NOR2_X1 u5_mult_87_U1851 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n261), .ZN(
        u5_mult_87_ab_34__19_) );
  NOR2_X1 u5_mult_87_U1850 ( .A1(u5_mult_87_n447), .A2(u5_mult_87_n458), .ZN(
        u5_mult_87_ab_34__1_) );
  NOR2_X1 u5_mult_87_U1849 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n458), .ZN(
        u5_mult_87_ab_34__20_) );
  NOR2_X1 u5_mult_87_U1848 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n458), .ZN(
        u5_mult_87_ab_34__21_) );
  NOR2_X1 u5_mult_87_U1847 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__22_) );
  NOR2_X1 u5_mult_87_U1846 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__23_) );
  NOR2_X1 u5_mult_87_U1845 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__24_) );
  NOR2_X1 u5_mult_87_U1844 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n458), .ZN(
        u5_mult_87_ab_34__25_) );
  NOR2_X1 u5_mult_87_U1843 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n458), .ZN(
        u5_mult_87_ab_34__26_) );
  NOR2_X1 u5_mult_87_U1842 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n458), .ZN(
        u5_mult_87_ab_34__27_) );
  NOR2_X1 u5_mult_87_U1841 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n458), .ZN(
        u5_mult_87_ab_34__28_) );
  NOR2_X1 u5_mult_87_U1840 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n458), .ZN(
        u5_mult_87_ab_34__29_) );
  NOR2_X1 u5_mult_87_U1839 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n261), .ZN(
        u5_mult_87_ab_34__2_) );
  NOR2_X1 u5_mult_87_U1838 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n261), .ZN(
        u5_mult_87_ab_34__30_) );
  NOR2_X1 u5_mult_87_U1837 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n261), .ZN(
        u5_mult_87_ab_34__31_) );
  NOR2_X1 u5_mult_87_U1836 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n261), .ZN(
        u5_mult_87_ab_34__32_) );
  NOR2_X1 u5_mult_87_U1835 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n261), .ZN(
        u5_mult_87_ab_34__33_) );
  NOR2_X1 u5_mult_87_U1834 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n261), .ZN(
        u5_mult_87_ab_34__34_) );
  NOR2_X1 u5_mult_87_U1833 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n261), .ZN(
        u5_mult_87_ab_34__35_) );
  NOR2_X1 u5_mult_87_U1832 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n261), .ZN(
        u5_mult_87_ab_34__36_) );
  NOR2_X1 u5_mult_87_U1831 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n261), .ZN(
        u5_mult_87_ab_34__37_) );
  NOR2_X1 u5_mult_87_U1830 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n261), .ZN(
        u5_mult_87_ab_34__38_) );
  NOR2_X1 u5_mult_87_U1829 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n261), .ZN(
        u5_mult_87_ab_34__39_) );
  NOR2_X1 u5_mult_87_U1828 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__3_) );
  NOR2_X1 u5_mult_87_U1827 ( .A1(u5_mult_87_n367), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__40_) );
  NOR2_X1 u5_mult_87_U1826 ( .A1(u5_mult_87_n365), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__41_) );
  NOR2_X1 u5_mult_87_U1825 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__42_) );
  NOR2_X1 u5_mult_87_U1824 ( .A1(u5_mult_87_n360), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__43_) );
  NOR2_X1 u5_mult_87_U1823 ( .A1(u5_mult_87_n358), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__44_) );
  NOR2_X1 u5_mult_87_U1822 ( .A1(u5_mult_87_n356), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__45_) );
  NOR2_X1 u5_mult_87_U1821 ( .A1(u5_mult_87_n354), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__46_) );
  NOR2_X1 u5_mult_87_U1820 ( .A1(u5_mult_87_n351), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__47_) );
  NOR2_X1 u5_mult_87_U1819 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__48_) );
  NOR2_X1 u5_mult_87_U1818 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__49_) );
  NOR2_X1 u5_mult_87_U1817 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__4_) );
  NOR2_X1 u5_mult_87_U1816 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__50_) );
  NOR2_X1 u5_mult_87_U1815 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__51_) );
  NOR2_X1 u5_mult_87_U1814 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__52_) );
  NOR2_X1 u5_mult_87_U1813 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__5_) );
  NOR2_X1 u5_mult_87_U1812 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__6_) );
  NOR2_X1 u5_mult_87_U1811 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__7_) );
  NOR2_X1 u5_mult_87_U1810 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__8_) );
  NOR2_X1 u5_mult_87_U1809 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n262), .ZN(
        u5_mult_87_ab_34__9_) );
  NOR2_X1 u5_mult_87_U1808 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n457), .ZN(
        u5_mult_87_ab_35__0_) );
  NOR2_X1 u5_mult_87_U1807 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n259), .ZN(
        u5_mult_87_ab_35__10_) );
  NOR2_X1 u5_mult_87_U1806 ( .A1(u5_mult_87_n425), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__11_) );
  NOR2_X1 u5_mult_87_U1805 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__12_) );
  NOR2_X1 u5_mult_87_U1804 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__13_) );
  NOR2_X1 u5_mult_87_U1803 ( .A1(u5_mult_87_n418), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__14_) );
  NOR2_X1 u5_mult_87_U1802 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__15_) );
  NOR2_X1 u5_mult_87_U1801 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n259), .ZN(
        u5_mult_87_ab_35__16_) );
  NOR2_X1 u5_mult_87_U1800 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n259), .ZN(
        u5_mult_87_ab_35__17_) );
  NOR2_X1 u5_mult_87_U1799 ( .A1(u5_mult_87_n411), .A2(u5_mult_87_n457), .ZN(
        u5_mult_87_ab_35__18_) );
  NOR2_X1 u5_mult_87_U1798 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n457), .ZN(
        u5_mult_87_ab_35__19_) );
  NOR2_X1 u5_mult_87_U1797 ( .A1(u5_mult_87_n447), .A2(u5_mult_87_n457), .ZN(
        u5_mult_87_ab_35__1_) );
  NOR2_X1 u5_mult_87_U1796 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n457), .ZN(
        u5_mult_87_ab_35__20_) );
  NOR2_X1 u5_mult_87_U1795 ( .A1(u5_mult_87_n406), .A2(u5_mult_87_n259), .ZN(
        u5_mult_87_ab_35__21_) );
  NOR2_X1 u5_mult_87_U1794 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n457), .ZN(
        u5_mult_87_ab_35__22_) );
  NOR2_X1 u5_mult_87_U1793 ( .A1(u5_mult_87_n402), .A2(u5_mult_87_n259), .ZN(
        u5_mult_87_ab_35__23_) );
  NOR2_X1 u5_mult_87_U1792 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n259), .ZN(
        u5_mult_87_ab_35__24_) );
  NOR2_X1 u5_mult_87_U1791 ( .A1(u5_mult_87_n398), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__25_) );
  NOR2_X1 u5_mult_87_U1790 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n457), .ZN(
        u5_mult_87_ab_35__26_) );
  NOR2_X1 u5_mult_87_U1789 ( .A1(u5_mult_87_n394), .A2(u5_mult_87_n457), .ZN(
        u5_mult_87_ab_35__27_) );
  NOR2_X1 u5_mult_87_U1788 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n457), .ZN(
        u5_mult_87_ab_35__28_) );
  NOR2_X1 u5_mult_87_U1787 ( .A1(u5_mult_87_n390), .A2(u5_mult_87_n457), .ZN(
        u5_mult_87_ab_35__29_) );
  NOR2_X1 u5_mult_87_U1786 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n259), .ZN(
        u5_mult_87_ab_35__2_) );
  NOR2_X1 u5_mult_87_U1785 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n259), .ZN(
        u5_mult_87_ab_35__30_) );
  NOR2_X1 u5_mult_87_U1784 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n259), .ZN(
        u5_mult_87_ab_35__31_) );
  NOR2_X1 u5_mult_87_U1783 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n259), .ZN(
        u5_mult_87_ab_35__32_) );
  NOR2_X1 u5_mult_87_U1782 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n259), .ZN(
        u5_mult_87_ab_35__33_) );
  NOR2_X1 u5_mult_87_U1781 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n259), .ZN(
        u5_mult_87_ab_35__34_) );
  NOR2_X1 u5_mult_87_U1780 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n259), .ZN(
        u5_mult_87_ab_35__35_) );
  NOR2_X1 u5_mult_87_U1779 ( .A1(u5_mult_87_n376), .A2(u5_mult_87_n259), .ZN(
        u5_mult_87_ab_35__36_) );
  NOR2_X1 u5_mult_87_U1778 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n259), .ZN(
        u5_mult_87_ab_35__37_) );
  NOR2_X1 u5_mult_87_U1777 ( .A1(u5_mult_87_n372), .A2(u5_mult_87_n259), .ZN(
        u5_mult_87_ab_35__38_) );
  NOR2_X1 u5_mult_87_U1776 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n259), .ZN(
        u5_mult_87_ab_35__39_) );
  NOR2_X1 u5_mult_87_U1775 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__3_) );
  NOR2_X1 u5_mult_87_U1774 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__40_) );
  NOR2_X1 u5_mult_87_U1773 ( .A1(u5_mult_87_n365), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__41_) );
  NOR2_X1 u5_mult_87_U1772 ( .A1(u5_mult_87_n363), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__42_) );
  NOR2_X1 u5_mult_87_U1771 ( .A1(u5_mult_87_n360), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__43_) );
  NOR2_X1 u5_mult_87_U1770 ( .A1(u5_mult_87_n358), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__44_) );
  NOR2_X1 u5_mult_87_U1769 ( .A1(u5_mult_87_n356), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__45_) );
  NOR2_X1 u5_mult_87_U1768 ( .A1(u5_mult_87_n354), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__46_) );
  NOR2_X1 u5_mult_87_U1767 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__47_) );
  NOR2_X1 u5_mult_87_U1766 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__48_) );
  NOR2_X1 u5_mult_87_U1765 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__49_) );
  NOR2_X1 u5_mult_87_U1764 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__4_) );
  NOR2_X1 u5_mult_87_U1763 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__50_) );
  NOR2_X1 u5_mult_87_U1762 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__51_) );
  NOR2_X1 u5_mult_87_U1761 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__52_) );
  NOR2_X1 u5_mult_87_U1760 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__5_) );
  NOR2_X1 u5_mult_87_U1759 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__6_) );
  NOR2_X1 u5_mult_87_U1758 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__7_) );
  NOR2_X1 u5_mult_87_U1757 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n260), .ZN(
        u5_mult_87_ab_35__8_) );
  NOR2_X1 u5_mult_87_U1756 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n259), .ZN(
        u5_mult_87_ab_35__9_) );
  NOR2_X1 u5_mult_87_U1755 ( .A1(u5_mult_87_n450), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__0_) );
  NOR2_X1 u5_mult_87_U1754 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__10_) );
  NOR2_X1 u5_mult_87_U1753 ( .A1(u5_mult_87_n425), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__11_) );
  NOR2_X1 u5_mult_87_U1752 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__12_) );
  NOR2_X1 u5_mult_87_U1751 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__13_) );
  NOR2_X1 u5_mult_87_U1750 ( .A1(u5_mult_87_n418), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__14_) );
  NOR2_X1 u5_mult_87_U1749 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n256), .ZN(
        u5_mult_87_ab_36__15_) );
  NOR2_X1 u5_mult_87_U1748 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n256), .ZN(
        u5_mult_87_ab_36__16_) );
  NOR2_X1 u5_mult_87_U1747 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n258), .ZN(
        u5_mult_87_ab_36__17_) );
  NOR2_X1 u5_mult_87_U1746 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n258), .ZN(
        u5_mult_87_ab_36__18_) );
  NOR2_X1 u5_mult_87_U1745 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n258), .ZN(
        u5_mult_87_ab_36__19_) );
  NOR2_X1 u5_mult_87_U1744 ( .A1(u5_mult_87_n447), .A2(u5_mult_87_n256), .ZN(
        u5_mult_87_ab_36__1_) );
  NOR2_X1 u5_mult_87_U1743 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n256), .ZN(
        u5_mult_87_ab_36__20_) );
  NOR2_X1 u5_mult_87_U1742 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n256), .ZN(
        u5_mult_87_ab_36__21_) );
  NOR2_X1 u5_mult_87_U1741 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n256), .ZN(
        u5_mult_87_ab_36__22_) );
  NOR2_X1 u5_mult_87_U1740 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n256), .ZN(
        u5_mult_87_ab_36__23_) );
  NOR2_X1 u5_mult_87_U1739 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n256), .ZN(
        u5_mult_87_ab_36__24_) );
  NOR2_X1 u5_mult_87_U1738 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n256), .ZN(
        u5_mult_87_ab_36__25_) );
  NOR2_X1 u5_mult_87_U1737 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n256), .ZN(
        u5_mult_87_ab_36__26_) );
  NOR2_X1 u5_mult_87_U1736 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n256), .ZN(
        u5_mult_87_ab_36__27_) );
  NOR2_X1 u5_mult_87_U1735 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n256), .ZN(
        u5_mult_87_ab_36__28_) );
  NOR2_X1 u5_mult_87_U1734 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n256), .ZN(
        u5_mult_87_ab_36__29_) );
  NOR2_X1 u5_mult_87_U1733 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__2_) );
  NOR2_X1 u5_mult_87_U1732 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__30_) );
  NOR2_X1 u5_mult_87_U1731 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__31_) );
  NOR2_X1 u5_mult_87_U1730 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__32_) );
  NOR2_X1 u5_mult_87_U1729 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__33_) );
  NOR2_X1 u5_mult_87_U1728 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__34_) );
  NOR2_X1 u5_mult_87_U1727 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__35_) );
  NOR2_X1 u5_mult_87_U1726 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__36_) );
  NOR2_X1 u5_mult_87_U1725 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__37_) );
  NOR2_X1 u5_mult_87_U1724 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__38_) );
  NOR2_X1 u5_mult_87_U1723 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__39_) );
  NOR2_X1 u5_mult_87_U1722 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__3_) );
  NOR2_X1 u5_mult_87_U1721 ( .A1(u5_mult_87_n367), .A2(u5_mult_87_n258), .ZN(
        u5_mult_87_ab_36__40_) );
  NOR2_X1 u5_mult_87_U1720 ( .A1(u5_mult_87_n365), .A2(u5_mult_87_n258), .ZN(
        u5_mult_87_ab_36__41_) );
  NOR2_X1 u5_mult_87_U1719 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__42_) );
  NOR2_X1 u5_mult_87_U1718 ( .A1(u5_mult_87_n360), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__43_) );
  NOR2_X1 u5_mult_87_U1717 ( .A1(u5_mult_87_n358), .A2(u5_mult_87_n256), .ZN(
        u5_mult_87_ab_36__44_) );
  NOR2_X1 u5_mult_87_U1716 ( .A1(u5_mult_87_n356), .A2(u5_mult_87_n256), .ZN(
        u5_mult_87_ab_36__45_) );
  NOR2_X1 u5_mult_87_U1715 ( .A1(u5_mult_87_n354), .A2(u5_mult_87_n256), .ZN(
        u5_mult_87_ab_36__46_) );
  NOR2_X1 u5_mult_87_U1714 ( .A1(u5_mult_87_n351), .A2(u5_mult_87_n258), .ZN(
        u5_mult_87_ab_36__47_) );
  NOR2_X1 u5_mult_87_U1713 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n258), .ZN(
        u5_mult_87_ab_36__48_) );
  NOR2_X1 u5_mult_87_U1712 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__49_) );
  NOR2_X1 u5_mult_87_U1711 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n258), .ZN(
        u5_mult_87_ab_36__4_) );
  NOR2_X1 u5_mult_87_U1710 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n258), .ZN(
        u5_mult_87_ab_36__50_) );
  NOR2_X1 u5_mult_87_U1709 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n258), .ZN(
        u5_mult_87_ab_36__51_) );
  NOR2_X1 u5_mult_87_U1708 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__52_) );
  NOR2_X1 u5_mult_87_U1707 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n258), .ZN(
        u5_mult_87_ab_36__5_) );
  NOR2_X1 u5_mult_87_U1706 ( .A1(u5_mult_87_n436), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__6_) );
  NOR2_X1 u5_mult_87_U1705 ( .A1(u5_mult_87_n434), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__7_) );
  NOR2_X1 u5_mult_87_U1704 ( .A1(u5_mult_87_n432), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__8_) );
  NOR2_X1 u5_mult_87_U1703 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n257), .ZN(
        u5_mult_87_ab_36__9_) );
  NOR2_X1 u5_mult_87_U1702 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__0_) );
  NOR2_X1 u5_mult_87_U1701 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__10_) );
  NOR2_X1 u5_mult_87_U1700 ( .A1(u5_mult_87_n425), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__11_) );
  NOR2_X1 u5_mult_87_U1699 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__12_) );
  NOR2_X1 u5_mult_87_U1698 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n254), .ZN(
        u5_mult_87_ab_37__13_) );
  NOR2_X1 u5_mult_87_U1697 ( .A1(u5_mult_87_n418), .A2(u5_mult_87_n254), .ZN(
        u5_mult_87_ab_37__14_) );
  NOR2_X1 u5_mult_87_U1696 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n254), .ZN(
        u5_mult_87_ab_37__15_) );
  NOR2_X1 u5_mult_87_U1695 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n456), .ZN(
        u5_mult_87_ab_37__16_) );
  NOR2_X1 u5_mult_87_U1694 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n456), .ZN(
        u5_mult_87_ab_37__17_) );
  NOR2_X1 u5_mult_87_U1693 ( .A1(u5_mult_87_n411), .A2(u5_mult_87_n456), .ZN(
        u5_mult_87_ab_37__18_) );
  NOR2_X1 u5_mult_87_U1692 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n254), .ZN(
        u5_mult_87_ab_37__19_) );
  NOR2_X1 u5_mult_87_U1691 ( .A1(u5_mult_87_n447), .A2(u5_mult_87_n456), .ZN(
        u5_mult_87_ab_37__1_) );
  NOR2_X1 u5_mult_87_U1690 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n456), .ZN(
        u5_mult_87_ab_37__20_) );
  NOR2_X1 u5_mult_87_U1689 ( .A1(u5_mult_87_n406), .A2(u5_mult_87_n254), .ZN(
        u5_mult_87_ab_37__21_) );
  NOR2_X1 u5_mult_87_U1688 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__22_) );
  NOR2_X1 u5_mult_87_U1687 ( .A1(u5_mult_87_n402), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__23_) );
  NOR2_X1 u5_mult_87_U1686 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n456), .ZN(
        u5_mult_87_ab_37__24_) );
  NOR2_X1 u5_mult_87_U1685 ( .A1(u5_mult_87_n398), .A2(u5_mult_87_n456), .ZN(
        u5_mult_87_ab_37__25_) );
  NOR2_X1 u5_mult_87_U1684 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n456), .ZN(
        u5_mult_87_ab_37__26_) );
  NOR2_X1 u5_mult_87_U1683 ( .A1(u5_mult_87_n394), .A2(u5_mult_87_n456), .ZN(
        u5_mult_87_ab_37__27_) );
  NOR2_X1 u5_mult_87_U1682 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n456), .ZN(
        u5_mult_87_ab_37__28_) );
  NOR2_X1 u5_mult_87_U1681 ( .A1(u5_mult_87_n390), .A2(u5_mult_87_n456), .ZN(
        u5_mult_87_ab_37__29_) );
  NOR2_X1 u5_mult_87_U1680 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n254), .ZN(
        u5_mult_87_ab_37__2_) );
  NOR2_X1 u5_mult_87_U1679 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n254), .ZN(
        u5_mult_87_ab_37__30_) );
  NOR2_X1 u5_mult_87_U1678 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n254), .ZN(
        u5_mult_87_ab_37__31_) );
  NOR2_X1 u5_mult_87_U1677 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n254), .ZN(
        u5_mult_87_ab_37__32_) );
  NOR2_X1 u5_mult_87_U1676 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n254), .ZN(
        u5_mult_87_ab_37__33_) );
  NOR2_X1 u5_mult_87_U1675 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n254), .ZN(
        u5_mult_87_ab_37__34_) );
  NOR2_X1 u5_mult_87_U1674 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n254), .ZN(
        u5_mult_87_ab_37__35_) );
  NOR2_X1 u5_mult_87_U1673 ( .A1(u5_mult_87_n376), .A2(u5_mult_87_n254), .ZN(
        u5_mult_87_ab_37__36_) );
  NOR2_X1 u5_mult_87_U1672 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n254), .ZN(
        u5_mult_87_ab_37__37_) );
  NOR2_X1 u5_mult_87_U1671 ( .A1(u5_mult_87_n372), .A2(u5_mult_87_n254), .ZN(
        u5_mult_87_ab_37__38_) );
  NOR2_X1 u5_mult_87_U1670 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n254), .ZN(
        u5_mult_87_ab_37__39_) );
  NOR2_X1 u5_mult_87_U1669 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__3_) );
  NOR2_X1 u5_mult_87_U1668 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__40_) );
  NOR2_X1 u5_mult_87_U1667 ( .A1(u5_mult_87_n365), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__41_) );
  NOR2_X1 u5_mult_87_U1666 ( .A1(u5_mult_87_n363), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__42_) );
  NOR2_X1 u5_mult_87_U1665 ( .A1(u5_mult_87_n360), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__43_) );
  NOR2_X1 u5_mult_87_U1664 ( .A1(u5_mult_87_n358), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__44_) );
  NOR2_X1 u5_mult_87_U1663 ( .A1(u5_mult_87_n356), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__45_) );
  NOR2_X1 u5_mult_87_U1662 ( .A1(u5_mult_87_n354), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__46_) );
  NOR2_X1 u5_mult_87_U1661 ( .A1(u5_mult_87_n351), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__47_) );
  NOR2_X1 u5_mult_87_U1660 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__48_) );
  NOR2_X1 u5_mult_87_U1659 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__49_) );
  NOR2_X1 u5_mult_87_U1658 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__4_) );
  NOR2_X1 u5_mult_87_U1657 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__50_) );
  NOR2_X1 u5_mult_87_U1656 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__51_) );
  NOR2_X1 u5_mult_87_U1655 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__52_) );
  NOR2_X1 u5_mult_87_U1654 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__5_) );
  NOR2_X1 u5_mult_87_U1653 ( .A1(u5_mult_87_n436), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__6_) );
  NOR2_X1 u5_mult_87_U1652 ( .A1(u5_mult_87_n434), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__7_) );
  NOR2_X1 u5_mult_87_U1651 ( .A1(u5_mult_87_n432), .A2(u5_mult_87_n255), .ZN(
        u5_mult_87_ab_37__8_) );
  NOR2_X1 u5_mult_87_U1650 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n254), .ZN(
        u5_mult_87_ab_37__9_) );
  NOR2_X1 u5_mult_87_U1649 ( .A1(u5_mult_87_n450), .A2(u5_mult_87_n252), .ZN(
        u5_mult_87_ab_38__0_) );
  NOR2_X1 u5_mult_87_U1648 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n252), .ZN(
        u5_mult_87_ab_38__10_) );
  NOR2_X1 u5_mult_87_U1647 ( .A1(u5_mult_87_n425), .A2(u5_mult_87_n251), .ZN(
        u5_mult_87_ab_38__11_) );
  NOR2_X1 u5_mult_87_U1646 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n251), .ZN(
        u5_mult_87_ab_38__12_) );
  NOR2_X1 u5_mult_87_U1645 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n253), .ZN(
        u5_mult_87_ab_38__13_) );
  NOR2_X1 u5_mult_87_U1644 ( .A1(u5_mult_87_n418), .A2(u5_mult_87_n253), .ZN(
        u5_mult_87_ab_38__14_) );
  NOR2_X1 u5_mult_87_U1643 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n253), .ZN(
        u5_mult_87_ab_38__15_) );
  NOR2_X1 u5_mult_87_U1642 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n253), .ZN(
        u5_mult_87_ab_38__16_) );
  NOR2_X1 u5_mult_87_U1641 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n253), .ZN(
        u5_mult_87_ab_38__17_) );
  NOR2_X1 u5_mult_87_U1640 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n251), .ZN(
        u5_mult_87_ab_38__18_) );
  NOR2_X1 u5_mult_87_U1639 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n253), .ZN(
        u5_mult_87_ab_38__19_) );
  NOR2_X1 u5_mult_87_U1638 ( .A1(u5_mult_87_n447), .A2(u5_mult_87_n253), .ZN(
        u5_mult_87_ab_38__1_) );
  NOR2_X1 u5_mult_87_U1637 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n253), .ZN(
        u5_mult_87_ab_38__20_) );
  NOR2_X1 u5_mult_87_U1636 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n253), .ZN(
        u5_mult_87_ab_38__21_) );
  NOR2_X1 u5_mult_87_U1635 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n253), .ZN(
        u5_mult_87_ab_38__22_) );
  NOR2_X1 u5_mult_87_U1634 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n253), .ZN(
        u5_mult_87_ab_38__23_) );
  NOR2_X1 u5_mult_87_U1633 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n253), .ZN(
        u5_mult_87_ab_38__24_) );
  NOR2_X1 u5_mult_87_U1632 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n253), .ZN(
        u5_mult_87_ab_38__25_) );
  NOR2_X1 u5_mult_87_U1631 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n253), .ZN(
        u5_mult_87_ab_38__26_) );
  NOR2_X1 u5_mult_87_U1630 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n253), .ZN(
        u5_mult_87_ab_38__27_) );
  NOR2_X1 u5_mult_87_U1629 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n253), .ZN(
        u5_mult_87_ab_38__28_) );
  NOR2_X1 u5_mult_87_U1628 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n253), .ZN(
        u5_mult_87_ab_38__29_) );
  NOR2_X1 u5_mult_87_U1627 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n251), .ZN(
        u5_mult_87_ab_38__2_) );
  NOR2_X1 u5_mult_87_U1626 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n251), .ZN(
        u5_mult_87_ab_38__30_) );
  NOR2_X1 u5_mult_87_U1625 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n251), .ZN(
        u5_mult_87_ab_38__31_) );
  NOR2_X1 u5_mult_87_U1624 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n251), .ZN(
        u5_mult_87_ab_38__32_) );
  NOR2_X1 u5_mult_87_U1623 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n251), .ZN(
        u5_mult_87_ab_38__33_) );
  NOR2_X1 u5_mult_87_U1622 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n251), .ZN(
        u5_mult_87_ab_38__34_) );
  NOR2_X1 u5_mult_87_U1621 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n251), .ZN(
        u5_mult_87_ab_38__35_) );
  NOR2_X1 u5_mult_87_U1620 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n251), .ZN(
        u5_mult_87_ab_38__36_) );
  NOR2_X1 u5_mult_87_U1619 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n251), .ZN(
        u5_mult_87_ab_38__37_) );
  NOR2_X1 u5_mult_87_U1618 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n251), .ZN(
        u5_mult_87_ab_38__38_) );
  NOR2_X1 u5_mult_87_U1617 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n251), .ZN(
        u5_mult_87_ab_38__39_) );
  NOR2_X1 u5_mult_87_U1616 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n252), .ZN(
        u5_mult_87_ab_38__3_) );
  NOR2_X1 u5_mult_87_U1615 ( .A1(u5_mult_87_n367), .A2(u5_mult_87_n252), .ZN(
        u5_mult_87_ab_38__40_) );
  NOR2_X1 u5_mult_87_U1614 ( .A1(u5_mult_87_n365), .A2(u5_mult_87_n252), .ZN(
        u5_mult_87_ab_38__41_) );
  NOR2_X1 u5_mult_87_U1613 ( .A1(u5_mult_87_n364), .A2(u5_mult_87_n252), .ZN(
        u5_mult_87_ab_38__42_) );
  NOR2_X1 u5_mult_87_U1612 ( .A1(u5_mult_87_n360), .A2(u5_mult_87_n252), .ZN(
        u5_mult_87_ab_38__43_) );
  NOR2_X1 u5_mult_87_U1611 ( .A1(u5_mult_87_n358), .A2(u5_mult_87_n252), .ZN(
        u5_mult_87_ab_38__44_) );
  NOR2_X1 u5_mult_87_U1610 ( .A1(u5_mult_87_n356), .A2(u5_mult_87_n252), .ZN(
        u5_mult_87_ab_38__45_) );
  NOR2_X1 u5_mult_87_U1609 ( .A1(u5_mult_87_n354), .A2(u5_mult_87_n252), .ZN(
        u5_mult_87_ab_38__46_) );
  NOR2_X1 u5_mult_87_U1608 ( .A1(u5_mult_87_n351), .A2(u5_mult_87_n252), .ZN(
        u5_mult_87_ab_38__47_) );
  NOR2_X1 u5_mult_87_U1607 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n252), .ZN(
        u5_mult_87_ab_38__48_) );
  NOR2_X1 u5_mult_87_U1606 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n252), .ZN(
        u5_mult_87_ab_38__49_) );
  NOR2_X1 u5_mult_87_U1605 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n252), .ZN(
        u5_mult_87_ab_38__4_) );
  NOR2_X1 u5_mult_87_U1604 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n252), .ZN(
        u5_mult_87_ab_38__50_) );
  NOR2_X1 u5_mult_87_U1603 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n252), .ZN(
        u5_mult_87_ab_38__51_) );
  NOR2_X1 u5_mult_87_U1602 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n252), .ZN(
        u5_mult_87_ab_38__52_) );
  NOR2_X1 u5_mult_87_U1601 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n252), .ZN(
        u5_mult_87_ab_38__5_) );
  NOR2_X1 u5_mult_87_U1600 ( .A1(u5_mult_87_n436), .A2(u5_mult_87_n252), .ZN(
        u5_mult_87_ab_38__6_) );
  NOR2_X1 u5_mult_87_U1599 ( .A1(u5_mult_87_n434), .A2(u5_mult_87_n252), .ZN(
        u5_mult_87_ab_38__7_) );
  NOR2_X1 u5_mult_87_U1598 ( .A1(u5_mult_87_n432), .A2(u5_mult_87_n252), .ZN(
        u5_mult_87_ab_38__8_) );
  NOR2_X1 u5_mult_87_U1597 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n251), .ZN(
        u5_mult_87_ab_38__9_) );
  NOR2_X1 u5_mult_87_U1596 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n249), .ZN(
        u5_mult_87_ab_39__0_) );
  NOR2_X1 u5_mult_87_U1595 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n250), .ZN(
        u5_mult_87_ab_39__10_) );
  NOR2_X1 u5_mult_87_U1594 ( .A1(u5_mult_87_n425), .A2(u5_mult_87_n250), .ZN(
        u5_mult_87_ab_39__11_) );
  NOR2_X1 u5_mult_87_U1593 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n248), .ZN(
        u5_mult_87_ab_39__12_) );
  NOR2_X1 u5_mult_87_U1592 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n248), .ZN(
        u5_mult_87_ab_39__13_) );
  NOR2_X1 u5_mult_87_U1591 ( .A1(u5_mult_87_n418), .A2(u5_mult_87_n248), .ZN(
        u5_mult_87_ab_39__14_) );
  NOR2_X1 u5_mult_87_U1590 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n250), .ZN(
        u5_mult_87_ab_39__15_) );
  NOR2_X1 u5_mult_87_U1589 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n250), .ZN(
        u5_mult_87_ab_39__16_) );
  NOR2_X1 u5_mult_87_U1588 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n248), .ZN(
        u5_mult_87_ab_39__17_) );
  NOR2_X1 u5_mult_87_U1587 ( .A1(u5_mult_87_n411), .A2(u5_mult_87_n248), .ZN(
        u5_mult_87_ab_39__18_) );
  NOR2_X1 u5_mult_87_U1586 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n248), .ZN(
        u5_mult_87_ab_39__19_) );
  NOR2_X1 u5_mult_87_U1585 ( .A1(u5_mult_87_n447), .A2(u5_mult_87_n248), .ZN(
        u5_mult_87_ab_39__1_) );
  NOR2_X1 u5_mult_87_U1584 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n248), .ZN(
        u5_mult_87_ab_39__20_) );
  NOR2_X1 u5_mult_87_U1583 ( .A1(u5_mult_87_n406), .A2(u5_mult_87_n248), .ZN(
        u5_mult_87_ab_39__21_) );
  NOR2_X1 u5_mult_87_U1582 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n248), .ZN(
        u5_mult_87_ab_39__22_) );
  NOR2_X1 u5_mult_87_U1581 ( .A1(u5_mult_87_n402), .A2(u5_mult_87_n248), .ZN(
        u5_mult_87_ab_39__23_) );
  NOR2_X1 u5_mult_87_U1580 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n248), .ZN(
        u5_mult_87_ab_39__24_) );
  NOR2_X1 u5_mult_87_U1579 ( .A1(u5_mult_87_n398), .A2(u5_mult_87_n248), .ZN(
        u5_mult_87_ab_39__25_) );
  NOR2_X1 u5_mult_87_U1578 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n248), .ZN(
        u5_mult_87_ab_39__26_) );
  NOR2_X1 u5_mult_87_U1577 ( .A1(u5_mult_87_n394), .A2(u5_mult_87_n248), .ZN(
        u5_mult_87_ab_39__27_) );
  NOR2_X1 u5_mult_87_U1576 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n248), .ZN(
        u5_mult_87_ab_39__28_) );
  NOR2_X1 u5_mult_87_U1575 ( .A1(u5_mult_87_n390), .A2(u5_mult_87_n248), .ZN(
        u5_mult_87_ab_39__29_) );
  NOR2_X1 u5_mult_87_U1574 ( .A1(u5_mult_87_n444), .A2(u5_mult_87_n249), .ZN(
        u5_mult_87_ab_39__2_) );
  NOR2_X1 u5_mult_87_U1573 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n249), .ZN(
        u5_mult_87_ab_39__30_) );
  NOR2_X1 u5_mult_87_U1572 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n249), .ZN(
        u5_mult_87_ab_39__31_) );
  NOR2_X1 u5_mult_87_U1571 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n249), .ZN(
        u5_mult_87_ab_39__32_) );
  NOR2_X1 u5_mult_87_U1570 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n249), .ZN(
        u5_mult_87_ab_39__33_) );
  NOR2_X1 u5_mult_87_U1569 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n249), .ZN(
        u5_mult_87_ab_39__34_) );
  NOR2_X1 u5_mult_87_U1568 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n249), .ZN(
        u5_mult_87_ab_39__35_) );
  NOR2_X1 u5_mult_87_U1567 ( .A1(u5_mult_87_n376), .A2(u5_mult_87_n249), .ZN(
        u5_mult_87_ab_39__36_) );
  NOR2_X1 u5_mult_87_U1566 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n249), .ZN(
        u5_mult_87_ab_39__37_) );
  NOR2_X1 u5_mult_87_U1565 ( .A1(u5_mult_87_n372), .A2(u5_mult_87_n249), .ZN(
        u5_mult_87_ab_39__38_) );
  NOR2_X1 u5_mult_87_U1564 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n249), .ZN(
        u5_mult_87_ab_39__39_) );
  NOR2_X1 u5_mult_87_U1563 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n249), .ZN(
        u5_mult_87_ab_39__3_) );
  NOR2_X1 u5_mult_87_U1562 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n249), .ZN(
        u5_mult_87_ab_39__40_) );
  NOR2_X1 u5_mult_87_U1561 ( .A1(u5_mult_87_n365), .A2(u5_mult_87_n249), .ZN(
        u5_mult_87_ab_39__41_) );
  NOR2_X1 u5_mult_87_U1560 ( .A1(u5_mult_87_n364), .A2(u5_mult_87_n249), .ZN(
        u5_mult_87_ab_39__42_) );
  NOR2_X1 u5_mult_87_U1559 ( .A1(u5_mult_87_n360), .A2(u5_mult_87_n249), .ZN(
        u5_mult_87_ab_39__43_) );
  NOR2_X1 u5_mult_87_U1558 ( .A1(u5_mult_87_n358), .A2(u5_mult_87_n249), .ZN(
        u5_mult_87_ab_39__44_) );
  NOR2_X1 u5_mult_87_U1557 ( .A1(u5_mult_87_n356), .A2(u5_mult_87_n249), .ZN(
        u5_mult_87_ab_39__45_) );
  NOR2_X1 u5_mult_87_U1556 ( .A1(u5_mult_87_n354), .A2(u5_mult_87_n249), .ZN(
        u5_mult_87_ab_39__46_) );
  NOR2_X1 u5_mult_87_U1555 ( .A1(u5_mult_87_n351), .A2(u5_mult_87_n249), .ZN(
        u5_mult_87_ab_39__47_) );
  NOR2_X1 u5_mult_87_U1554 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n249), .ZN(
        u5_mult_87_ab_39__48_) );
  NOR2_X1 u5_mult_87_U1553 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n249), .ZN(
        u5_mult_87_ab_39__49_) );
  NOR2_X1 u5_mult_87_U1552 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n250), .ZN(
        u5_mult_87_ab_39__4_) );
  NOR2_X1 u5_mult_87_U1551 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n250), .ZN(
        u5_mult_87_ab_39__50_) );
  NOR2_X1 u5_mult_87_U1550 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n250), .ZN(
        u5_mult_87_ab_39__51_) );
  NOR2_X1 u5_mult_87_U1549 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n250), .ZN(
        u5_mult_87_ab_39__52_) );
  NOR2_X1 u5_mult_87_U1548 ( .A1(u5_mult_87_n439), .A2(u5_mult_87_n250), .ZN(
        u5_mult_87_ab_39__5_) );
  NOR2_X1 u5_mult_87_U1547 ( .A1(u5_mult_87_n436), .A2(u5_mult_87_n250), .ZN(
        u5_mult_87_ab_39__6_) );
  NOR2_X1 u5_mult_87_U1546 ( .A1(u5_mult_87_n434), .A2(u5_mult_87_n250), .ZN(
        u5_mult_87_ab_39__7_) );
  NOR2_X1 u5_mult_87_U1545 ( .A1(u5_mult_87_n432), .A2(u5_mult_87_n250), .ZN(
        u5_mult_87_ab_39__8_) );
  NOR2_X1 u5_mult_87_U1544 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n250), .ZN(
        u5_mult_87_ab_39__9_) );
  NOR2_X1 u5_mult_87_U1543 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__0_) );
  NOR2_X1 u5_mult_87_U1542 ( .A1(u5_mult_87_n428), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__10_) );
  NOR2_X1 u5_mult_87_U1541 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__11_) );
  NOR2_X1 u5_mult_87_U1540 ( .A1(u5_mult_87_n481), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__12_) );
  NOR2_X1 u5_mult_87_U1539 ( .A1(u5_mult_87_n422), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__13_) );
  NOR2_X1 u5_mult_87_U1538 ( .A1(u5_mult_87_n419), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__14_) );
  NOR2_X1 u5_mult_87_U1537 ( .A1(u5_mult_87_n416), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__15_) );
  NOR2_X1 u5_mult_87_U1536 ( .A1(u5_mult_87_n480), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__16_) );
  NOR2_X1 u5_mult_87_U1535 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__17_) );
  NOR2_X1 u5_mult_87_U1534 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__18_) );
  NOR2_X1 u5_mult_87_U1533 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__19_) );
  NOR2_X1 u5_mult_87_U1532 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__1_) );
  NOR2_X1 u5_mult_87_U1531 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__20_) );
  NOR2_X1 u5_mult_87_U1530 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__21_) );
  NOR2_X1 u5_mult_87_U1529 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__22_) );
  NOR2_X1 u5_mult_87_U1528 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__23_) );
  NOR2_X1 u5_mult_87_U1527 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__24_) );
  NOR2_X1 u5_mult_87_U1526 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__25_) );
  NOR2_X1 u5_mult_87_U1525 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__26_) );
  NOR2_X1 u5_mult_87_U1524 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__27_) );
  NOR2_X1 u5_mult_87_U1523 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__28_) );
  NOR2_X1 u5_mult_87_U1522 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__29_) );
  NOR2_X1 u5_mult_87_U1521 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n330), .ZN(
        u5_mult_87_ab_3__2_) );
  NOR2_X1 u5_mult_87_U1520 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n330), .ZN(
        u5_mult_87_ab_3__30_) );
  NOR2_X1 u5_mult_87_U1519 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n330), .ZN(
        u5_mult_87_ab_3__31_) );
  NOR2_X1 u5_mult_87_U1518 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n330), .ZN(
        u5_mult_87_ab_3__32_) );
  NOR2_X1 u5_mult_87_U1517 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n330), .ZN(
        u5_mult_87_ab_3__33_) );
  NOR2_X1 u5_mult_87_U1516 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n330), .ZN(
        u5_mult_87_ab_3__34_) );
  NOR2_X1 u5_mult_87_U1515 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n330), .ZN(
        u5_mult_87_ab_3__35_) );
  NOR2_X1 u5_mult_87_U1514 ( .A1(u5_mult_87_n376), .A2(u5_mult_87_n330), .ZN(
        u5_mult_87_ab_3__36_) );
  NOR2_X1 u5_mult_87_U1513 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n330), .ZN(
        u5_mult_87_ab_3__37_) );
  NOR2_X1 u5_mult_87_U1512 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n330), .ZN(
        u5_mult_87_ab_3__38_) );
  NOR2_X1 u5_mult_87_U1511 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n330), .ZN(
        u5_mult_87_ab_3__39_) );
  NOR2_X1 u5_mult_87_U1510 ( .A1(u5_mult_87_n442), .A2(u5_mult_87_n331), .ZN(
        u5_mult_87_ab_3__3_) );
  NOR2_X1 u5_mult_87_U1509 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n331), .ZN(
        u5_mult_87_ab_3__40_) );
  NOR2_X1 u5_mult_87_U1508 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n331), .ZN(
        u5_mult_87_ab_3__41_) );
  NOR2_X1 u5_mult_87_U1507 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n331), .ZN(
        u5_mult_87_ab_3__42_) );
  NOR2_X1 u5_mult_87_U1506 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n331), .ZN(
        u5_mult_87_ab_3__43_) );
  NOR2_X1 u5_mult_87_U1505 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n331), .ZN(
        u5_mult_87_ab_3__44_) );
  NOR2_X1 u5_mult_87_U1504 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n331), .ZN(
        u5_mult_87_ab_3__45_) );
  NOR2_X1 u5_mult_87_U1503 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n331), .ZN(
        u5_mult_87_ab_3__46_) );
  NOR2_X1 u5_mult_87_U1502 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n331), .ZN(
        u5_mult_87_ab_3__47_) );
  NOR2_X1 u5_mult_87_U1501 ( .A1(u5_mult_87_n350), .A2(u5_mult_87_n331), .ZN(
        u5_mult_87_ab_3__48_) );
  NOR2_X1 u5_mult_87_U1500 ( .A1(u5_mult_87_n348), .A2(u5_mult_87_n331), .ZN(
        u5_mult_87_ab_3__49_) );
  NOR2_X1 u5_mult_87_U1499 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__4_) );
  NOR2_X1 u5_mult_87_U1498 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n331), .ZN(
        u5_mult_87_ab_3__50_) );
  NOR2_X1 u5_mult_87_U1497 ( .A1(u5_mult_87_n345), .A2(u5_mult_87_n478), .ZN(
        u5_mult_87_ab_3__51_) );
  NOR2_X1 u5_mult_87_U1496 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n330), .ZN(
        u5_mult_87_ab_3__52_) );
  NOR2_X1 u5_mult_87_U1495 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__5_) );
  NOR2_X1 u5_mult_87_U1494 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__6_) );
  NOR2_X1 u5_mult_87_U1493 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__7_) );
  NOR2_X1 u5_mult_87_U1492 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__8_) );
  NOR2_X1 u5_mult_87_U1491 ( .A1(u5_mult_87_n430), .A2(u5_mult_87_n329), .ZN(
        u5_mult_87_ab_3__9_) );
  NOR2_X1 u5_mult_87_U1490 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n246), .ZN(
        u5_mult_87_ab_40__0_) );
  NOR2_X1 u5_mult_87_U1489 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n455), .ZN(
        u5_mult_87_ab_40__10_) );
  NOR2_X1 u5_mult_87_U1488 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n455), .ZN(
        u5_mult_87_ab_40__11_) );
  NOR2_X1 u5_mult_87_U1487 ( .A1(u5_mult_87_n481), .A2(u5_mult_87_n455), .ZN(
        u5_mult_87_ab_40__12_) );
  NOR2_X1 u5_mult_87_U1486 ( .A1(u5_mult_87_n422), .A2(u5_mult_87_n455), .ZN(
        u5_mult_87_ab_40__13_) );
  NOR2_X1 u5_mult_87_U1485 ( .A1(u5_mult_87_n419), .A2(u5_mult_87_n455), .ZN(
        u5_mult_87_ab_40__14_) );
  NOR2_X1 u5_mult_87_U1484 ( .A1(u5_mult_87_n416), .A2(u5_mult_87_n455), .ZN(
        u5_mult_87_ab_40__15_) );
  NOR2_X1 u5_mult_87_U1483 ( .A1(u5_mult_87_n480), .A2(u5_mult_87_n455), .ZN(
        u5_mult_87_ab_40__16_) );
  NOR2_X1 u5_mult_87_U1482 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n245), .ZN(
        u5_mult_87_ab_40__17_) );
  NOR2_X1 u5_mult_87_U1481 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n455), .ZN(
        u5_mult_87_ab_40__18_) );
  NOR2_X1 u5_mult_87_U1480 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n455), .ZN(
        u5_mult_87_ab_40__19_) );
  NOR2_X1 u5_mult_87_U1479 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n244), .ZN(
        u5_mult_87_ab_40__1_) );
  NOR2_X1 u5_mult_87_U1478 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n244), .ZN(
        u5_mult_87_ab_40__20_) );
  NOR2_X1 u5_mult_87_U1477 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n244), .ZN(
        u5_mult_87_ab_40__21_) );
  NOR2_X1 u5_mult_87_U1476 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n244), .ZN(
        u5_mult_87_ab_40__22_) );
  NOR2_X1 u5_mult_87_U1475 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n244), .ZN(
        u5_mult_87_ab_40__23_) );
  NOR2_X1 u5_mult_87_U1474 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n244), .ZN(
        u5_mult_87_ab_40__24_) );
  NOR2_X1 u5_mult_87_U1473 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n244), .ZN(
        u5_mult_87_ab_40__25_) );
  NOR2_X1 u5_mult_87_U1472 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n244), .ZN(
        u5_mult_87_ab_40__26_) );
  NOR2_X1 u5_mult_87_U1471 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n244), .ZN(
        u5_mult_87_ab_40__27_) );
  NOR2_X1 u5_mult_87_U1470 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n244), .ZN(
        u5_mult_87_ab_40__28_) );
  NOR2_X1 u5_mult_87_U1469 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n244), .ZN(
        u5_mult_87_ab_40__29_) );
  NOR2_X1 u5_mult_87_U1468 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n245), .ZN(
        u5_mult_87_ab_40__2_) );
  NOR2_X1 u5_mult_87_U1467 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n245), .ZN(
        u5_mult_87_ab_40__30_) );
  NOR2_X1 u5_mult_87_U1466 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n245), .ZN(
        u5_mult_87_ab_40__31_) );
  NOR2_X1 u5_mult_87_U1465 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n245), .ZN(
        u5_mult_87_ab_40__32_) );
  NOR2_X1 u5_mult_87_U1464 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n245), .ZN(
        u5_mult_87_ab_40__33_) );
  NOR2_X1 u5_mult_87_U1463 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n245), .ZN(
        u5_mult_87_ab_40__34_) );
  NOR2_X1 u5_mult_87_U1462 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n245), .ZN(
        u5_mult_87_ab_40__35_) );
  NOR2_X1 u5_mult_87_U1461 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n245), .ZN(
        u5_mult_87_ab_40__36_) );
  NOR2_X1 u5_mult_87_U1460 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n245), .ZN(
        u5_mult_87_ab_40__37_) );
  NOR2_X1 u5_mult_87_U1459 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n245), .ZN(
        u5_mult_87_ab_40__38_) );
  NOR2_X1 u5_mult_87_U1458 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n245), .ZN(
        u5_mult_87_ab_40__39_) );
  NOR2_X1 u5_mult_87_U1457 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n246), .ZN(
        u5_mult_87_ab_40__3_) );
  NOR2_X1 u5_mult_87_U1456 ( .A1(u5_mult_87_n367), .A2(u5_mult_87_n246), .ZN(
        u5_mult_87_ab_40__40_) );
  NOR2_X1 u5_mult_87_U1455 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n246), .ZN(
        u5_mult_87_ab_40__41_) );
  NOR2_X1 u5_mult_87_U1454 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n246), .ZN(
        u5_mult_87_ab_40__42_) );
  NOR2_X1 u5_mult_87_U1453 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n246), .ZN(
        u5_mult_87_ab_40__43_) );
  NOR2_X1 u5_mult_87_U1452 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n246), .ZN(
        u5_mult_87_ab_40__44_) );
  NOR2_X1 u5_mult_87_U1451 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n246), .ZN(
        u5_mult_87_ab_40__45_) );
  NOR2_X1 u5_mult_87_U1450 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n246), .ZN(
        u5_mult_87_ab_40__46_) );
  NOR2_X1 u5_mult_87_U1449 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n246), .ZN(
        u5_mult_87_ab_40__47_) );
  NOR2_X1 u5_mult_87_U1448 ( .A1(u5_mult_87_n350), .A2(u5_mult_87_n246), .ZN(
        u5_mult_87_ab_40__48_) );
  NOR2_X1 u5_mult_87_U1447 ( .A1(u5_mult_87_n348), .A2(u5_mult_87_n246), .ZN(
        u5_mult_87_ab_40__49_) );
  NOR2_X1 u5_mult_87_U1446 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n245), .ZN(
        u5_mult_87_ab_40__4_) );
  NOR2_X1 u5_mult_87_U1445 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n246), .ZN(
        u5_mult_87_ab_40__50_) );
  NOR2_X1 u5_mult_87_U1444 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n245), .ZN(
        u5_mult_87_ab_40__51_) );
  NOR2_X1 u5_mult_87_U1443 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n246), .ZN(
        u5_mult_87_ab_40__52_) );
  NOR2_X1 u5_mult_87_U1442 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n246), .ZN(
        u5_mult_87_ab_40__5_) );
  NOR2_X1 u5_mult_87_U1441 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n246), .ZN(
        u5_mult_87_ab_40__6_) );
  NOR2_X1 u5_mult_87_U1440 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n246), .ZN(
        u5_mult_87_ab_40__7_) );
  NOR2_X1 u5_mult_87_U1439 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n245), .ZN(
        u5_mult_87_ab_40__8_) );
  NOR2_X1 u5_mult_87_U1438 ( .A1(u5_mult_87_n430), .A2(u5_mult_87_n244), .ZN(
        u5_mult_87_ab_40__9_) );
  NOR2_X1 u5_mult_87_U1437 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n241), .ZN(
        u5_mult_87_ab_41__0_) );
  NOR2_X1 u5_mult_87_U1436 ( .A1(u5_mult_87_n428), .A2(u5_mult_87_n243), .ZN(
        u5_mult_87_ab_41__10_) );
  NOR2_X1 u5_mult_87_U1435 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n240), .ZN(
        u5_mult_87_ab_41__11_) );
  NOR2_X1 u5_mult_87_U1434 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n243), .ZN(
        u5_mult_87_ab_41__12_) );
  NOR2_X1 u5_mult_87_U1433 ( .A1(u5_mult_87_n422), .A2(u5_mult_87_n243), .ZN(
        u5_mult_87_ab_41__13_) );
  NOR2_X1 u5_mult_87_U1432 ( .A1(u5_mult_87_n419), .A2(u5_mult_87_n243), .ZN(
        u5_mult_87_ab_41__14_) );
  NOR2_X1 u5_mult_87_U1431 ( .A1(u5_mult_87_n416), .A2(u5_mult_87_n243), .ZN(
        u5_mult_87_ab_41__15_) );
  NOR2_X1 u5_mult_87_U1430 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n243), .ZN(
        u5_mult_87_ab_41__16_) );
  NOR2_X1 u5_mult_87_U1429 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n243), .ZN(
        u5_mult_87_ab_41__17_) );
  NOR2_X1 u5_mult_87_U1428 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n243), .ZN(
        u5_mult_87_ab_41__18_) );
  NOR2_X1 u5_mult_87_U1427 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n241), .ZN(
        u5_mult_87_ab_41__19_) );
  NOR2_X1 u5_mult_87_U1426 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n240), .ZN(
        u5_mult_87_ab_41__1_) );
  NOR2_X1 u5_mult_87_U1425 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n240), .ZN(
        u5_mult_87_ab_41__20_) );
  NOR2_X1 u5_mult_87_U1424 ( .A1(u5_mult_87_n406), .A2(u5_mult_87_n240), .ZN(
        u5_mult_87_ab_41__21_) );
  NOR2_X1 u5_mult_87_U1423 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n240), .ZN(
        u5_mult_87_ab_41__22_) );
  NOR2_X1 u5_mult_87_U1422 ( .A1(u5_mult_87_n402), .A2(u5_mult_87_n240), .ZN(
        u5_mult_87_ab_41__23_) );
  NOR2_X1 u5_mult_87_U1421 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n240), .ZN(
        u5_mult_87_ab_41__24_) );
  NOR2_X1 u5_mult_87_U1420 ( .A1(u5_mult_87_n398), .A2(u5_mult_87_n240), .ZN(
        u5_mult_87_ab_41__25_) );
  NOR2_X1 u5_mult_87_U1419 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n240), .ZN(
        u5_mult_87_ab_41__26_) );
  NOR2_X1 u5_mult_87_U1418 ( .A1(u5_mult_87_n394), .A2(u5_mult_87_n240), .ZN(
        u5_mult_87_ab_41__27_) );
  NOR2_X1 u5_mult_87_U1417 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n240), .ZN(
        u5_mult_87_ab_41__28_) );
  NOR2_X1 u5_mult_87_U1416 ( .A1(u5_mult_87_n390), .A2(u5_mult_87_n240), .ZN(
        u5_mult_87_ab_41__29_) );
  NOR2_X1 u5_mult_87_U1415 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n241), .ZN(
        u5_mult_87_ab_41__2_) );
  NOR2_X1 u5_mult_87_U1414 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n241), .ZN(
        u5_mult_87_ab_41__30_) );
  NOR2_X1 u5_mult_87_U1413 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n241), .ZN(
        u5_mult_87_ab_41__31_) );
  NOR2_X1 u5_mult_87_U1412 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n241), .ZN(
        u5_mult_87_ab_41__32_) );
  NOR2_X1 u5_mult_87_U1411 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n241), .ZN(
        u5_mult_87_ab_41__33_) );
  NOR2_X1 u5_mult_87_U1410 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n241), .ZN(
        u5_mult_87_ab_41__34_) );
  NOR2_X1 u5_mult_87_U1409 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n241), .ZN(
        u5_mult_87_ab_41__35_) );
  NOR2_X1 u5_mult_87_U1408 ( .A1(u5_mult_87_n376), .A2(u5_mult_87_n241), .ZN(
        u5_mult_87_ab_41__36_) );
  NOR2_X1 u5_mult_87_U1407 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n241), .ZN(
        u5_mult_87_ab_41__37_) );
  NOR2_X1 u5_mult_87_U1406 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n241), .ZN(
        u5_mult_87_ab_41__38_) );
  NOR2_X1 u5_mult_87_U1405 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n241), .ZN(
        u5_mult_87_ab_41__39_) );
  NOR2_X1 u5_mult_87_U1404 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n242), .ZN(
        u5_mult_87_ab_41__3_) );
  NOR2_X1 u5_mult_87_U1403 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n242), .ZN(
        u5_mult_87_ab_41__40_) );
  NOR2_X1 u5_mult_87_U1402 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n242), .ZN(
        u5_mult_87_ab_41__41_) );
  NOR2_X1 u5_mult_87_U1401 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n242), .ZN(
        u5_mult_87_ab_41__42_) );
  NOR2_X1 u5_mult_87_U1400 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n242), .ZN(
        u5_mult_87_ab_41__43_) );
  NOR2_X1 u5_mult_87_U1399 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n242), .ZN(
        u5_mult_87_ab_41__44_) );
  NOR2_X1 u5_mult_87_U1398 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n242), .ZN(
        u5_mult_87_ab_41__45_) );
  NOR2_X1 u5_mult_87_U1397 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n242), .ZN(
        u5_mult_87_ab_41__46_) );
  NOR2_X1 u5_mult_87_U1396 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n242), .ZN(
        u5_mult_87_ab_41__47_) );
  NOR2_X1 u5_mult_87_U1395 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n242), .ZN(
        u5_mult_87_ab_41__48_) );
  NOR2_X1 u5_mult_87_U1394 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n242), .ZN(
        u5_mult_87_ab_41__49_) );
  NOR2_X1 u5_mult_87_U1393 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n241), .ZN(
        u5_mult_87_ab_41__4_) );
  NOR2_X1 u5_mult_87_U1392 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n242), .ZN(
        u5_mult_87_ab_41__50_) );
  NOR2_X1 u5_mult_87_U1391 ( .A1(u5_mult_87_n345), .A2(u5_mult_87_n241), .ZN(
        u5_mult_87_ab_41__51_) );
  NOR2_X1 u5_mult_87_U1390 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n242), .ZN(
        u5_mult_87_ab_41__52_) );
  NOR2_X1 u5_mult_87_U1389 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n242), .ZN(
        u5_mult_87_ab_41__5_) );
  NOR2_X1 u5_mult_87_U1388 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n241), .ZN(
        u5_mult_87_ab_41__6_) );
  NOR2_X1 u5_mult_87_U1387 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n241), .ZN(
        u5_mult_87_ab_41__7_) );
  NOR2_X1 u5_mult_87_U1386 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n242), .ZN(
        u5_mult_87_ab_41__8_) );
  NOR2_X1 u5_mult_87_U1385 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n240), .ZN(
        u5_mult_87_ab_41__9_) );
  NOR2_X1 u5_mult_87_U1384 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n239), .ZN(
        u5_mult_87_ab_42__0_) );
  NOR2_X1 u5_mult_87_U1383 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n236), .ZN(
        u5_mult_87_ab_42__10_) );
  NOR2_X1 u5_mult_87_U1382 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n239), .ZN(
        u5_mult_87_ab_42__11_) );
  NOR2_X1 u5_mult_87_U1381 ( .A1(u5_mult_87_n481), .A2(u5_mult_87_n239), .ZN(
        u5_mult_87_ab_42__12_) );
  NOR2_X1 u5_mult_87_U1380 ( .A1(u5_mult_87_n422), .A2(u5_mult_87_n239), .ZN(
        u5_mult_87_ab_42__13_) );
  NOR2_X1 u5_mult_87_U1379 ( .A1(u5_mult_87_n419), .A2(u5_mult_87_n239), .ZN(
        u5_mult_87_ab_42__14_) );
  NOR2_X1 u5_mult_87_U1378 ( .A1(u5_mult_87_n416), .A2(u5_mult_87_n236), .ZN(
        u5_mult_87_ab_42__15_) );
  NOR2_X1 u5_mult_87_U1377 ( .A1(u5_mult_87_n480), .A2(u5_mult_87_n237), .ZN(
        u5_mult_87_ab_42__16_) );
  NOR2_X1 u5_mult_87_U1376 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n237), .ZN(
        u5_mult_87_ab_42__17_) );
  NOR2_X1 u5_mult_87_U1375 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n237), .ZN(
        u5_mult_87_ab_42__18_) );
  NOR2_X1 u5_mult_87_U1374 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n239), .ZN(
        u5_mult_87_ab_42__19_) );
  NOR2_X1 u5_mult_87_U1373 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n236), .ZN(
        u5_mult_87_ab_42__1_) );
  NOR2_X1 u5_mult_87_U1372 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n236), .ZN(
        u5_mult_87_ab_42__20_) );
  NOR2_X1 u5_mult_87_U1371 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n236), .ZN(
        u5_mult_87_ab_42__21_) );
  NOR2_X1 u5_mult_87_U1370 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n236), .ZN(
        u5_mult_87_ab_42__22_) );
  NOR2_X1 u5_mult_87_U1369 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n236), .ZN(
        u5_mult_87_ab_42__23_) );
  NOR2_X1 u5_mult_87_U1368 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n236), .ZN(
        u5_mult_87_ab_42__24_) );
  NOR2_X1 u5_mult_87_U1367 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n236), .ZN(
        u5_mult_87_ab_42__25_) );
  NOR2_X1 u5_mult_87_U1366 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n236), .ZN(
        u5_mult_87_ab_42__26_) );
  NOR2_X1 u5_mult_87_U1365 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n236), .ZN(
        u5_mult_87_ab_42__27_) );
  NOR2_X1 u5_mult_87_U1364 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n236), .ZN(
        u5_mult_87_ab_42__28_) );
  NOR2_X1 u5_mult_87_U1363 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n236), .ZN(
        u5_mult_87_ab_42__29_) );
  NOR2_X1 u5_mult_87_U1362 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n237), .ZN(
        u5_mult_87_ab_42__2_) );
  NOR2_X1 u5_mult_87_U1361 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n237), .ZN(
        u5_mult_87_ab_42__30_) );
  NOR2_X1 u5_mult_87_U1360 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n237), .ZN(
        u5_mult_87_ab_42__31_) );
  NOR2_X1 u5_mult_87_U1359 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n237), .ZN(
        u5_mult_87_ab_42__32_) );
  NOR2_X1 u5_mult_87_U1358 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n237), .ZN(
        u5_mult_87_ab_42__33_) );
  NOR2_X1 u5_mult_87_U1357 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n237), .ZN(
        u5_mult_87_ab_42__34_) );
  NOR2_X1 u5_mult_87_U1356 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n237), .ZN(
        u5_mult_87_ab_42__35_) );
  NOR2_X1 u5_mult_87_U1355 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n237), .ZN(
        u5_mult_87_ab_42__36_) );
  NOR2_X1 u5_mult_87_U1354 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n237), .ZN(
        u5_mult_87_ab_42__37_) );
  NOR2_X1 u5_mult_87_U1353 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n237), .ZN(
        u5_mult_87_ab_42__38_) );
  NOR2_X1 u5_mult_87_U1352 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n237), .ZN(
        u5_mult_87_ab_42__39_) );
  NOR2_X1 u5_mult_87_U1351 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n238), .ZN(
        u5_mult_87_ab_42__3_) );
  NOR2_X1 u5_mult_87_U1350 ( .A1(u5_mult_87_n367), .A2(u5_mult_87_n238), .ZN(
        u5_mult_87_ab_42__40_) );
  NOR2_X1 u5_mult_87_U1349 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n238), .ZN(
        u5_mult_87_ab_42__41_) );
  NOR2_X1 u5_mult_87_U1348 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n238), .ZN(
        u5_mult_87_ab_42__42_) );
  NOR2_X1 u5_mult_87_U1347 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n238), .ZN(
        u5_mult_87_ab_42__43_) );
  NOR2_X1 u5_mult_87_U1346 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n238), .ZN(
        u5_mult_87_ab_42__44_) );
  NOR2_X1 u5_mult_87_U1345 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n238), .ZN(
        u5_mult_87_ab_42__45_) );
  NOR2_X1 u5_mult_87_U1344 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n238), .ZN(
        u5_mult_87_ab_42__46_) );
  NOR2_X1 u5_mult_87_U1343 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n238), .ZN(
        u5_mult_87_ab_42__47_) );
  NOR2_X1 u5_mult_87_U1342 ( .A1(u5_mult_87_n350), .A2(u5_mult_87_n238), .ZN(
        u5_mult_87_ab_42__48_) );
  NOR2_X1 u5_mult_87_U1341 ( .A1(u5_mult_87_n348), .A2(u5_mult_87_n238), .ZN(
        u5_mult_87_ab_42__49_) );
  NOR2_X1 u5_mult_87_U1340 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n236), .ZN(
        u5_mult_87_ab_42__4_) );
  NOR2_X1 u5_mult_87_U1339 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n237), .ZN(
        u5_mult_87_ab_42__50_) );
  NOR2_X1 u5_mult_87_U1338 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n236), .ZN(
        u5_mult_87_ab_42__51_) );
  NOR2_X1 u5_mult_87_U1337 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n237), .ZN(
        u5_mult_87_ab_42__52_) );
  NOR2_X1 u5_mult_87_U1336 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n237), .ZN(
        u5_mult_87_ab_42__5_) );
  NOR2_X1 u5_mult_87_U1335 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n237), .ZN(
        u5_mult_87_ab_42__6_) );
  NOR2_X1 u5_mult_87_U1334 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n237), .ZN(
        u5_mult_87_ab_42__7_) );
  NOR2_X1 u5_mult_87_U1333 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n236), .ZN(
        u5_mult_87_ab_42__8_) );
  NOR2_X1 u5_mult_87_U1332 ( .A1(u5_mult_87_n430), .A2(u5_mult_87_n238), .ZN(
        u5_mult_87_ab_42__9_) );
  NOR2_X1 u5_mult_87_U1331 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n234), .ZN(
        u5_mult_87_ab_43__0_) );
  NOR2_X1 u5_mult_87_U1330 ( .A1(u5_mult_87_n428), .A2(u5_mult_87_n234), .ZN(
        u5_mult_87_ab_43__10_) );
  NOR2_X1 u5_mult_87_U1329 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n235), .ZN(
        u5_mult_87_ab_43__11_) );
  NOR2_X1 u5_mult_87_U1328 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n235), .ZN(
        u5_mult_87_ab_43__12_) );
  NOR2_X1 u5_mult_87_U1327 ( .A1(u5_mult_87_n422), .A2(u5_mult_87_n234), .ZN(
        u5_mult_87_ab_43__13_) );
  NOR2_X1 u5_mult_87_U1326 ( .A1(u5_mult_87_n419), .A2(u5_mult_87_n234), .ZN(
        u5_mult_87_ab_43__14_) );
  NOR2_X1 u5_mult_87_U1325 ( .A1(u5_mult_87_n416), .A2(u5_mult_87_n233), .ZN(
        u5_mult_87_ab_43__15_) );
  NOR2_X1 u5_mult_87_U1324 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n234), .ZN(
        u5_mult_87_ab_43__16_) );
  NOR2_X1 u5_mult_87_U1323 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n233), .ZN(
        u5_mult_87_ab_43__17_) );
  NOR2_X1 u5_mult_87_U1322 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n234), .ZN(
        u5_mult_87_ab_43__18_) );
  NOR2_X1 u5_mult_87_U1321 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n233), .ZN(
        u5_mult_87_ab_43__19_) );
  NOR2_X1 u5_mult_87_U1320 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n233), .ZN(
        u5_mult_87_ab_43__1_) );
  NOR2_X1 u5_mult_87_U1319 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n233), .ZN(
        u5_mult_87_ab_43__20_) );
  NOR2_X1 u5_mult_87_U1318 ( .A1(u5_mult_87_n406), .A2(u5_mult_87_n233), .ZN(
        u5_mult_87_ab_43__21_) );
  NOR2_X1 u5_mult_87_U1317 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n233), .ZN(
        u5_mult_87_ab_43__22_) );
  NOR2_X1 u5_mult_87_U1316 ( .A1(u5_mult_87_n402), .A2(u5_mult_87_n233), .ZN(
        u5_mult_87_ab_43__23_) );
  NOR2_X1 u5_mult_87_U1315 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n233), .ZN(
        u5_mult_87_ab_43__24_) );
  NOR2_X1 u5_mult_87_U1314 ( .A1(u5_mult_87_n398), .A2(u5_mult_87_n233), .ZN(
        u5_mult_87_ab_43__25_) );
  NOR2_X1 u5_mult_87_U1313 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n233), .ZN(
        u5_mult_87_ab_43__26_) );
  NOR2_X1 u5_mult_87_U1312 ( .A1(u5_mult_87_n394), .A2(u5_mult_87_n233), .ZN(
        u5_mult_87_ab_43__27_) );
  NOR2_X1 u5_mult_87_U1311 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n233), .ZN(
        u5_mult_87_ab_43__28_) );
  NOR2_X1 u5_mult_87_U1310 ( .A1(u5_mult_87_n390), .A2(u5_mult_87_n233), .ZN(
        u5_mult_87_ab_43__29_) );
  NOR2_X1 u5_mult_87_U1309 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n234), .ZN(
        u5_mult_87_ab_43__2_) );
  NOR2_X1 u5_mult_87_U1308 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n234), .ZN(
        u5_mult_87_ab_43__30_) );
  NOR2_X1 u5_mult_87_U1307 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n234), .ZN(
        u5_mult_87_ab_43__31_) );
  NOR2_X1 u5_mult_87_U1306 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n234), .ZN(
        u5_mult_87_ab_43__32_) );
  NOR2_X1 u5_mult_87_U1305 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n234), .ZN(
        u5_mult_87_ab_43__33_) );
  NOR2_X1 u5_mult_87_U1304 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n234), .ZN(
        u5_mult_87_ab_43__34_) );
  NOR2_X1 u5_mult_87_U1303 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n234), .ZN(
        u5_mult_87_ab_43__35_) );
  NOR2_X1 u5_mult_87_U1302 ( .A1(u5_mult_87_n376), .A2(u5_mult_87_n234), .ZN(
        u5_mult_87_ab_43__36_) );
  NOR2_X1 u5_mult_87_U1301 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n234), .ZN(
        u5_mult_87_ab_43__37_) );
  NOR2_X1 u5_mult_87_U1300 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n234), .ZN(
        u5_mult_87_ab_43__38_) );
  NOR2_X1 u5_mult_87_U1299 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n234), .ZN(
        u5_mult_87_ab_43__39_) );
  NOR2_X1 u5_mult_87_U1298 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n235), .ZN(
        u5_mult_87_ab_43__3_) );
  NOR2_X1 u5_mult_87_U1297 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n235), .ZN(
        u5_mult_87_ab_43__40_) );
  NOR2_X1 u5_mult_87_U1296 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n235), .ZN(
        u5_mult_87_ab_43__41_) );
  NOR2_X1 u5_mult_87_U1295 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n235), .ZN(
        u5_mult_87_ab_43__42_) );
  NOR2_X1 u5_mult_87_U1294 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n235), .ZN(
        u5_mult_87_ab_43__43_) );
  NOR2_X1 u5_mult_87_U1293 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n235), .ZN(
        u5_mult_87_ab_43__44_) );
  NOR2_X1 u5_mult_87_U1292 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n235), .ZN(
        u5_mult_87_ab_43__45_) );
  NOR2_X1 u5_mult_87_U1291 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n235), .ZN(
        u5_mult_87_ab_43__46_) );
  NOR2_X1 u5_mult_87_U1290 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n235), .ZN(
        u5_mult_87_ab_43__47_) );
  NOR2_X1 u5_mult_87_U1289 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n235), .ZN(
        u5_mult_87_ab_43__48_) );
  NOR2_X1 u5_mult_87_U1288 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n235), .ZN(
        u5_mult_87_ab_43__49_) );
  NOR2_X1 u5_mult_87_U1287 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n234), .ZN(
        u5_mult_87_ab_43__4_) );
  NOR2_X1 u5_mult_87_U1286 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n233), .ZN(
        u5_mult_87_ab_43__50_) );
  NOR2_X1 u5_mult_87_U1285 ( .A1(u5_mult_87_n345), .A2(u5_mult_87_n234), .ZN(
        u5_mult_87_ab_43__51_) );
  NOR2_X1 u5_mult_87_U1284 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n233), .ZN(
        u5_mult_87_ab_43__52_) );
  NOR2_X1 u5_mult_87_U1283 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n233), .ZN(
        u5_mult_87_ab_43__5_) );
  NOR2_X1 u5_mult_87_U1282 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n233), .ZN(
        u5_mult_87_ab_43__6_) );
  NOR2_X1 u5_mult_87_U1281 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n233), .ZN(
        u5_mult_87_ab_43__7_) );
  NOR2_X1 u5_mult_87_U1280 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n234), .ZN(
        u5_mult_87_ab_43__8_) );
  NOR2_X1 u5_mult_87_U1279 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n235), .ZN(
        u5_mult_87_ab_43__9_) );
  NOR2_X1 u5_mult_87_U1278 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__0_) );
  NOR2_X1 u5_mult_87_U1277 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n232), .ZN(
        u5_mult_87_ab_44__10_) );
  NOR2_X1 u5_mult_87_U1276 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n232), .ZN(
        u5_mult_87_ab_44__11_) );
  NOR2_X1 u5_mult_87_U1275 ( .A1(u5_mult_87_n481), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__12_) );
  NOR2_X1 u5_mult_87_U1274 ( .A1(u5_mult_87_n422), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__13_) );
  NOR2_X1 u5_mult_87_U1273 ( .A1(u5_mult_87_n419), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__14_) );
  NOR2_X1 u5_mult_87_U1272 ( .A1(u5_mult_87_n416), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__15_) );
  NOR2_X1 u5_mult_87_U1271 ( .A1(u5_mult_87_n480), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__16_) );
  NOR2_X1 u5_mult_87_U1270 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__17_) );
  NOR2_X1 u5_mult_87_U1269 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__18_) );
  NOR2_X1 u5_mult_87_U1268 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__19_) );
  NOR2_X1 u5_mult_87_U1267 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__1_) );
  NOR2_X1 u5_mult_87_U1266 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__20_) );
  NOR2_X1 u5_mult_87_U1265 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__21_) );
  NOR2_X1 u5_mult_87_U1264 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__22_) );
  NOR2_X1 u5_mult_87_U1263 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__23_) );
  NOR2_X1 u5_mult_87_U1262 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__24_) );
  NOR2_X1 u5_mult_87_U1261 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__25_) );
  NOR2_X1 u5_mult_87_U1260 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__26_) );
  NOR2_X1 u5_mult_87_U1259 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__27_) );
  NOR2_X1 u5_mult_87_U1258 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__28_) );
  NOR2_X1 u5_mult_87_U1257 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__29_) );
  NOR2_X1 u5_mult_87_U1256 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n231), .ZN(
        u5_mult_87_ab_44__2_) );
  NOR2_X1 u5_mult_87_U1255 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n231), .ZN(
        u5_mult_87_ab_44__30_) );
  NOR2_X1 u5_mult_87_U1254 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n231), .ZN(
        u5_mult_87_ab_44__31_) );
  NOR2_X1 u5_mult_87_U1253 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n231), .ZN(
        u5_mult_87_ab_44__32_) );
  NOR2_X1 u5_mult_87_U1252 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n231), .ZN(
        u5_mult_87_ab_44__33_) );
  NOR2_X1 u5_mult_87_U1251 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n231), .ZN(
        u5_mult_87_ab_44__34_) );
  NOR2_X1 u5_mult_87_U1250 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n231), .ZN(
        u5_mult_87_ab_44__35_) );
  NOR2_X1 u5_mult_87_U1249 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n231), .ZN(
        u5_mult_87_ab_44__36_) );
  NOR2_X1 u5_mult_87_U1248 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n231), .ZN(
        u5_mult_87_ab_44__37_) );
  NOR2_X1 u5_mult_87_U1247 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n231), .ZN(
        u5_mult_87_ab_44__38_) );
  NOR2_X1 u5_mult_87_U1246 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n231), .ZN(
        u5_mult_87_ab_44__39_) );
  NOR2_X1 u5_mult_87_U1245 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n232), .ZN(
        u5_mult_87_ab_44__3_) );
  NOR2_X1 u5_mult_87_U1244 ( .A1(u5_mult_87_n367), .A2(u5_mult_87_n232), .ZN(
        u5_mult_87_ab_44__40_) );
  NOR2_X1 u5_mult_87_U1243 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n232), .ZN(
        u5_mult_87_ab_44__41_) );
  NOR2_X1 u5_mult_87_U1242 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n232), .ZN(
        u5_mult_87_ab_44__42_) );
  NOR2_X1 u5_mult_87_U1241 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n232), .ZN(
        u5_mult_87_ab_44__43_) );
  NOR2_X1 u5_mult_87_U1240 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n232), .ZN(
        u5_mult_87_ab_44__44_) );
  NOR2_X1 u5_mult_87_U1239 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n232), .ZN(
        u5_mult_87_ab_44__45_) );
  NOR2_X1 u5_mult_87_U1238 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n232), .ZN(
        u5_mult_87_ab_44__46_) );
  NOR2_X1 u5_mult_87_U1237 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n232), .ZN(
        u5_mult_87_ab_44__47_) );
  NOR2_X1 u5_mult_87_U1236 ( .A1(u5_mult_87_n350), .A2(u5_mult_87_n232), .ZN(
        u5_mult_87_ab_44__48_) );
  NOR2_X1 u5_mult_87_U1235 ( .A1(u5_mult_87_n348), .A2(u5_mult_87_n232), .ZN(
        u5_mult_87_ab_44__49_) );
  NOR2_X1 u5_mult_87_U1234 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__4_) );
  NOR2_X1 u5_mult_87_U1233 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n231), .ZN(
        u5_mult_87_ab_44__50_) );
  NOR2_X1 u5_mult_87_U1232 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__51_) );
  NOR2_X1 u5_mult_87_U1231 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n231), .ZN(
        u5_mult_87_ab_44__52_) );
  NOR2_X1 u5_mult_87_U1230 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n231), .ZN(
        u5_mult_87_ab_44__5_) );
  NOR2_X1 u5_mult_87_U1229 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__6_) );
  NOR2_X1 u5_mult_87_U1228 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n230), .ZN(
        u5_mult_87_ab_44__7_) );
  NOR2_X1 u5_mult_87_U1227 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n231), .ZN(
        u5_mult_87_ab_44__8_) );
  NOR2_X1 u5_mult_87_U1226 ( .A1(u5_mult_87_n430), .A2(u5_mult_87_n232), .ZN(
        u5_mult_87_ab_44__9_) );
  NOR2_X1 u5_mult_87_U1225 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__0_) );
  NOR2_X1 u5_mult_87_U1224 ( .A1(u5_mult_87_n428), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__10_) );
  NOR2_X1 u5_mult_87_U1223 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__11_) );
  NOR2_X1 u5_mult_87_U1222 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__12_) );
  NOR2_X1 u5_mult_87_U1221 ( .A1(u5_mult_87_n422), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__13_) );
  NOR2_X1 u5_mult_87_U1220 ( .A1(u5_mult_87_n419), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__14_) );
  NOR2_X1 u5_mult_87_U1219 ( .A1(u5_mult_87_n416), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__15_) );
  NOR2_X1 u5_mult_87_U1218 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__16_) );
  NOR2_X1 u5_mult_87_U1217 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__17_) );
  NOR2_X1 u5_mult_87_U1216 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n228), .ZN(
        u5_mult_87_ab_45__18_) );
  NOR2_X1 u5_mult_87_U1215 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__19_) );
  NOR2_X1 u5_mult_87_U1214 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__1_) );
  NOR2_X1 u5_mult_87_U1213 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__20_) );
  NOR2_X1 u5_mult_87_U1212 ( .A1(u5_mult_87_n406), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__21_) );
  NOR2_X1 u5_mult_87_U1211 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__22_) );
  NOR2_X1 u5_mult_87_U1210 ( .A1(u5_mult_87_n402), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__23_) );
  NOR2_X1 u5_mult_87_U1209 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__24_) );
  NOR2_X1 u5_mult_87_U1208 ( .A1(u5_mult_87_n398), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__25_) );
  NOR2_X1 u5_mult_87_U1207 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__26_) );
  NOR2_X1 u5_mult_87_U1206 ( .A1(u5_mult_87_n394), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__27_) );
  NOR2_X1 u5_mult_87_U1205 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__28_) );
  NOR2_X1 u5_mult_87_U1204 ( .A1(u5_mult_87_n390), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__29_) );
  NOR2_X1 u5_mult_87_U1203 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n228), .ZN(
        u5_mult_87_ab_45__2_) );
  NOR2_X1 u5_mult_87_U1202 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n228), .ZN(
        u5_mult_87_ab_45__30_) );
  NOR2_X1 u5_mult_87_U1201 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n228), .ZN(
        u5_mult_87_ab_45__31_) );
  NOR2_X1 u5_mult_87_U1200 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n228), .ZN(
        u5_mult_87_ab_45__32_) );
  NOR2_X1 u5_mult_87_U1199 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n228), .ZN(
        u5_mult_87_ab_45__33_) );
  NOR2_X1 u5_mult_87_U1198 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n228), .ZN(
        u5_mult_87_ab_45__34_) );
  NOR2_X1 u5_mult_87_U1197 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n228), .ZN(
        u5_mult_87_ab_45__35_) );
  NOR2_X1 u5_mult_87_U1196 ( .A1(u5_mult_87_n376), .A2(u5_mult_87_n228), .ZN(
        u5_mult_87_ab_45__36_) );
  NOR2_X1 u5_mult_87_U1195 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n228), .ZN(
        u5_mult_87_ab_45__37_) );
  NOR2_X1 u5_mult_87_U1194 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n228), .ZN(
        u5_mult_87_ab_45__38_) );
  NOR2_X1 u5_mult_87_U1193 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n228), .ZN(
        u5_mult_87_ab_45__39_) );
  NOR2_X1 u5_mult_87_U1192 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n229), .ZN(
        u5_mult_87_ab_45__3_) );
  NOR2_X1 u5_mult_87_U1191 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n229), .ZN(
        u5_mult_87_ab_45__40_) );
  NOR2_X1 u5_mult_87_U1190 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n229), .ZN(
        u5_mult_87_ab_45__41_) );
  NOR2_X1 u5_mult_87_U1189 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n229), .ZN(
        u5_mult_87_ab_45__42_) );
  NOR2_X1 u5_mult_87_U1188 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n229), .ZN(
        u5_mult_87_ab_45__43_) );
  NOR2_X1 u5_mult_87_U1187 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n229), .ZN(
        u5_mult_87_ab_45__44_) );
  NOR2_X1 u5_mult_87_U1186 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n229), .ZN(
        u5_mult_87_ab_45__45_) );
  NOR2_X1 u5_mult_87_U1185 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n229), .ZN(
        u5_mult_87_ab_45__46_) );
  NOR2_X1 u5_mult_87_U1184 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n229), .ZN(
        u5_mult_87_ab_45__47_) );
  NOR2_X1 u5_mult_87_U1183 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n229), .ZN(
        u5_mult_87_ab_45__48_) );
  NOR2_X1 u5_mult_87_U1182 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n229), .ZN(
        u5_mult_87_ab_45__49_) );
  NOR2_X1 u5_mult_87_U1181 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__4_) );
  NOR2_X1 u5_mult_87_U1180 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__50_) );
  NOR2_X1 u5_mult_87_U1179 ( .A1(u5_mult_87_n345), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__51_) );
  NOR2_X1 u5_mult_87_U1178 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__52_) );
  NOR2_X1 u5_mult_87_U1177 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__5_) );
  NOR2_X1 u5_mult_87_U1176 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n227), .ZN(
        u5_mult_87_ab_45__6_) );
  NOR2_X1 u5_mult_87_U1175 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n228), .ZN(
        u5_mult_87_ab_45__7_) );
  NOR2_X1 u5_mult_87_U1174 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n229), .ZN(
        u5_mult_87_ab_45__8_) );
  NOR2_X1 u5_mult_87_U1173 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n228), .ZN(
        u5_mult_87_ab_45__9_) );
  NOR2_X1 u5_mult_87_U1172 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n454), .ZN(
        u5_mult_87_ab_46__0_) );
  NOR2_X1 u5_mult_87_U1171 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__10_) );
  NOR2_X1 u5_mult_87_U1170 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__11_) );
  NOR2_X1 u5_mult_87_U1169 ( .A1(u5_mult_87_n481), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__12_) );
  NOR2_X1 u5_mult_87_U1168 ( .A1(u5_mult_87_n422), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__13_) );
  NOR2_X1 u5_mult_87_U1167 ( .A1(u5_mult_87_n419), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__14_) );
  NOR2_X1 u5_mult_87_U1166 ( .A1(u5_mult_87_n416), .A2(u5_mult_87_n454), .ZN(
        u5_mult_87_ab_46__15_) );
  NOR2_X1 u5_mult_87_U1165 ( .A1(u5_mult_87_n480), .A2(u5_mult_87_n454), .ZN(
        u5_mult_87_ab_46__16_) );
  NOR2_X1 u5_mult_87_U1164 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n454), .ZN(
        u5_mult_87_ab_46__17_) );
  NOR2_X1 u5_mult_87_U1163 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n454), .ZN(
        u5_mult_87_ab_46__18_) );
  NOR2_X1 u5_mult_87_U1162 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n454), .ZN(
        u5_mult_87_ab_46__19_) );
  NOR2_X1 u5_mult_87_U1161 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__1_) );
  NOR2_X1 u5_mult_87_U1160 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__20_) );
  NOR2_X1 u5_mult_87_U1159 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__21_) );
  NOR2_X1 u5_mult_87_U1158 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__22_) );
  NOR2_X1 u5_mult_87_U1157 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__23_) );
  NOR2_X1 u5_mult_87_U1156 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__24_) );
  NOR2_X1 u5_mult_87_U1155 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__25_) );
  NOR2_X1 u5_mult_87_U1154 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__26_) );
  NOR2_X1 u5_mult_87_U1153 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__27_) );
  NOR2_X1 u5_mult_87_U1152 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__28_) );
  NOR2_X1 u5_mult_87_U1151 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__29_) );
  NOR2_X1 u5_mult_87_U1150 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__2_) );
  NOR2_X1 u5_mult_87_U1149 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__30_) );
  NOR2_X1 u5_mult_87_U1148 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__31_) );
  NOR2_X1 u5_mult_87_U1147 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__32_) );
  NOR2_X1 u5_mult_87_U1146 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__33_) );
  NOR2_X1 u5_mult_87_U1145 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__34_) );
  NOR2_X1 u5_mult_87_U1144 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__35_) );
  NOR2_X1 u5_mult_87_U1143 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__36_) );
  NOR2_X1 u5_mult_87_U1142 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__37_) );
  NOR2_X1 u5_mult_87_U1141 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__38_) );
  NOR2_X1 u5_mult_87_U1140 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n225), .ZN(
        u5_mult_87_ab_46__39_) );
  NOR2_X1 u5_mult_87_U1139 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n226), .ZN(
        u5_mult_87_ab_46__3_) );
  NOR2_X1 u5_mult_87_U1138 ( .A1(u5_mult_87_n367), .A2(u5_mult_87_n226), .ZN(
        u5_mult_87_ab_46__40_) );
  NOR2_X1 u5_mult_87_U1137 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n226), .ZN(
        u5_mult_87_ab_46__41_) );
  NOR2_X1 u5_mult_87_U1136 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n226), .ZN(
        u5_mult_87_ab_46__42_) );
  NOR2_X1 u5_mult_87_U1135 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n226), .ZN(
        u5_mult_87_ab_46__43_) );
  NOR2_X1 u5_mult_87_U1134 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n226), .ZN(
        u5_mult_87_ab_46__44_) );
  NOR2_X1 u5_mult_87_U1133 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n226), .ZN(
        u5_mult_87_ab_46__45_) );
  NOR2_X1 u5_mult_87_U1132 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n226), .ZN(
        u5_mult_87_ab_46__46_) );
  NOR2_X1 u5_mult_87_U1131 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n226), .ZN(
        u5_mult_87_ab_46__47_) );
  NOR2_X1 u5_mult_87_U1130 ( .A1(u5_mult_87_n350), .A2(u5_mult_87_n226), .ZN(
        u5_mult_87_ab_46__48_) );
  NOR2_X1 u5_mult_87_U1129 ( .A1(u5_mult_87_n348), .A2(u5_mult_87_n226), .ZN(
        u5_mult_87_ab_46__49_) );
  NOR2_X1 u5_mult_87_U1128 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n226), .ZN(
        u5_mult_87_ab_46__4_) );
  NOR2_X1 u5_mult_87_U1127 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n226), .ZN(
        u5_mult_87_ab_46__50_) );
  NOR2_X1 u5_mult_87_U1126 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n226), .ZN(
        u5_mult_87_ab_46__51_) );
  NOR2_X1 u5_mult_87_U1125 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n226), .ZN(
        u5_mult_87_ab_46__52_) );
  NOR2_X1 u5_mult_87_U1124 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n226), .ZN(
        u5_mult_87_ab_46__5_) );
  NOR2_X1 u5_mult_87_U1123 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n226), .ZN(
        u5_mult_87_ab_46__6_) );
  NOR2_X1 u5_mult_87_U1122 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n454), .ZN(
        u5_mult_87_ab_46__7_) );
  NOR2_X1 u5_mult_87_U1121 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n454), .ZN(
        u5_mult_87_ab_46__8_) );
  NOR2_X1 u5_mult_87_U1120 ( .A1(u5_mult_87_n430), .A2(u5_mult_87_n454), .ZN(
        u5_mult_87_ab_46__9_) );
  NOR2_X1 u5_mult_87_U1119 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n222), .ZN(
        u5_mult_87_ab_47__0_) );
  NOR2_X1 u5_mult_87_U1118 ( .A1(u5_mult_87_n428), .A2(u5_mult_87_n222), .ZN(
        u5_mult_87_ab_47__10_) );
  NOR2_X1 u5_mult_87_U1117 ( .A1(u5_mult_87_n425), .A2(u5_mult_87_n222), .ZN(
        u5_mult_87_ab_47__11_) );
  NOR2_X1 u5_mult_87_U1116 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n222), .ZN(
        u5_mult_87_ab_47__12_) );
  NOR2_X1 u5_mult_87_U1115 ( .A1(u5_mult_87_n422), .A2(u5_mult_87_n222), .ZN(
        u5_mult_87_ab_47__13_) );
  NOR2_X1 u5_mult_87_U1114 ( .A1(u5_mult_87_n419), .A2(u5_mult_87_n222), .ZN(
        u5_mult_87_ab_47__14_) );
  NOR2_X1 u5_mult_87_U1113 ( .A1(u5_mult_87_n416), .A2(u5_mult_87_n222), .ZN(
        u5_mult_87_ab_47__15_) );
  NOR2_X1 u5_mult_87_U1112 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n222), .ZN(
        u5_mult_87_ab_47__16_) );
  NOR2_X1 u5_mult_87_U1111 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n222), .ZN(
        u5_mult_87_ab_47__17_) );
  NOR2_X1 u5_mult_87_U1110 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n222), .ZN(
        u5_mult_87_ab_47__18_) );
  NOR2_X1 u5_mult_87_U1109 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n222), .ZN(
        u5_mult_87_ab_47__19_) );
  NOR2_X1 u5_mult_87_U1108 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__1_) );
  NOR2_X1 u5_mult_87_U1107 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__20_) );
  NOR2_X1 u5_mult_87_U1106 ( .A1(u5_mult_87_n406), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__21_) );
  NOR2_X1 u5_mult_87_U1105 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__22_) );
  NOR2_X1 u5_mult_87_U1104 ( .A1(u5_mult_87_n402), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__23_) );
  NOR2_X1 u5_mult_87_U1103 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__24_) );
  NOR2_X1 u5_mult_87_U1102 ( .A1(u5_mult_87_n398), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__25_) );
  NOR2_X1 u5_mult_87_U1101 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__26_) );
  NOR2_X1 u5_mult_87_U1100 ( .A1(u5_mult_87_n394), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__27_) );
  NOR2_X1 u5_mult_87_U1099 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__28_) );
  NOR2_X1 u5_mult_87_U1098 ( .A1(u5_mult_87_n390), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__29_) );
  NOR2_X1 u5_mult_87_U1097 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n224), .ZN(
        u5_mult_87_ab_47__2_) );
  NOR2_X1 u5_mult_87_U1096 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n224), .ZN(
        u5_mult_87_ab_47__30_) );
  NOR2_X1 u5_mult_87_U1095 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n224), .ZN(
        u5_mult_87_ab_47__31_) );
  NOR2_X1 u5_mult_87_U1094 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n224), .ZN(
        u5_mult_87_ab_47__32_) );
  NOR2_X1 u5_mult_87_U1093 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n224), .ZN(
        u5_mult_87_ab_47__33_) );
  NOR2_X1 u5_mult_87_U1092 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n224), .ZN(
        u5_mult_87_ab_47__34_) );
  NOR2_X1 u5_mult_87_U1091 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n224), .ZN(
        u5_mult_87_ab_47__35_) );
  NOR2_X1 u5_mult_87_U1090 ( .A1(u5_mult_87_n376), .A2(u5_mult_87_n224), .ZN(
        u5_mult_87_ab_47__36_) );
  NOR2_X1 u5_mult_87_U1089 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n224), .ZN(
        u5_mult_87_ab_47__37_) );
  NOR2_X1 u5_mult_87_U1088 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n224), .ZN(
        u5_mult_87_ab_47__38_) );
  NOR2_X1 u5_mult_87_U1087 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n224), .ZN(
        u5_mult_87_ab_47__39_) );
  NOR2_X1 u5_mult_87_U1086 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__3_) );
  NOR2_X1 u5_mult_87_U1085 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__40_) );
  NOR2_X1 u5_mult_87_U1084 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__41_) );
  NOR2_X1 u5_mult_87_U1083 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__42_) );
  NOR2_X1 u5_mult_87_U1082 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__43_) );
  NOR2_X1 u5_mult_87_U1081 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__44_) );
  NOR2_X1 u5_mult_87_U1080 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__45_) );
  NOR2_X1 u5_mult_87_U1079 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__46_) );
  NOR2_X1 u5_mult_87_U1078 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__47_) );
  NOR2_X1 u5_mult_87_U1077 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__48_) );
  NOR2_X1 u5_mult_87_U1076 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__49_) );
  NOR2_X1 u5_mult_87_U1075 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__4_) );
  NOR2_X1 u5_mult_87_U1074 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__50_) );
  NOR2_X1 u5_mult_87_U1073 ( .A1(u5_mult_87_n345), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__51_) );
  NOR2_X1 u5_mult_87_U1072 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__52_) );
  NOR2_X1 u5_mult_87_U1071 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n224), .ZN(
        u5_mult_87_ab_47__5_) );
  NOR2_X1 u5_mult_87_U1070 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n222), .ZN(
        u5_mult_87_ab_47__6_) );
  NOR2_X1 u5_mult_87_U1069 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n224), .ZN(
        u5_mult_87_ab_47__7_) );
  NOR2_X1 u5_mult_87_U1068 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n224), .ZN(
        u5_mult_87_ab_47__8_) );
  NOR2_X1 u5_mult_87_U1067 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n223), .ZN(
        u5_mult_87_ab_47__9_) );
  NOR2_X1 u5_mult_87_U1066 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n220), .ZN(
        u5_mult_87_ab_48__0_) );
  NOR2_X1 u5_mult_87_U1065 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n221), .ZN(
        u5_mult_87_ab_48__10_) );
  NOR2_X1 u5_mult_87_U1064 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n220), .ZN(
        u5_mult_87_ab_48__11_) );
  NOR2_X1 u5_mult_87_U1063 ( .A1(u5_mult_87_n481), .A2(u5_mult_87_n221), .ZN(
        u5_mult_87_ab_48__12_) );
  NOR2_X1 u5_mult_87_U1062 ( .A1(u5_mult_87_n422), .A2(u5_mult_87_n220), .ZN(
        u5_mult_87_ab_48__13_) );
  NOR2_X1 u5_mult_87_U1061 ( .A1(u5_mult_87_n419), .A2(u5_mult_87_n221), .ZN(
        u5_mult_87_ab_48__14_) );
  NOR2_X1 u5_mult_87_U1060 ( .A1(u5_mult_87_n416), .A2(u5_mult_87_n220), .ZN(
        u5_mult_87_ab_48__15_) );
  NOR2_X1 u5_mult_87_U1059 ( .A1(u5_mult_87_n480), .A2(u5_mult_87_n221), .ZN(
        u5_mult_87_ab_48__16_) );
  NOR2_X1 u5_mult_87_U1058 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n221), .ZN(
        u5_mult_87_ab_48__17_) );
  NOR2_X1 u5_mult_87_U1057 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n221), .ZN(
        u5_mult_87_ab_48__18_) );
  NOR2_X1 u5_mult_87_U1056 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n221), .ZN(
        u5_mult_87_ab_48__19_) );
  NOR2_X1 u5_mult_87_U1055 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__1_) );
  NOR2_X1 u5_mult_87_U1054 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__20_) );
  NOR2_X1 u5_mult_87_U1053 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__21_) );
  NOR2_X1 u5_mult_87_U1052 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__22_) );
  NOR2_X1 u5_mult_87_U1051 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__23_) );
  NOR2_X1 u5_mult_87_U1050 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__24_) );
  NOR2_X1 u5_mult_87_U1049 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__25_) );
  NOR2_X1 u5_mult_87_U1048 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__26_) );
  NOR2_X1 u5_mult_87_U1047 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__27_) );
  NOR2_X1 u5_mult_87_U1046 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__28_) );
  NOR2_X1 u5_mult_87_U1045 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__29_) );
  NOR2_X1 u5_mult_87_U1044 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__2_) );
  NOR2_X1 u5_mult_87_U1043 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__30_) );
  NOR2_X1 u5_mult_87_U1042 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__31_) );
  NOR2_X1 u5_mult_87_U1041 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__32_) );
  NOR2_X1 u5_mult_87_U1040 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__33_) );
  NOR2_X1 u5_mult_87_U1039 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__34_) );
  NOR2_X1 u5_mult_87_U1038 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__35_) );
  NOR2_X1 u5_mult_87_U1037 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__36_) );
  NOR2_X1 u5_mult_87_U1036 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__37_) );
  NOR2_X1 u5_mult_87_U1035 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__38_) );
  NOR2_X1 u5_mult_87_U1034 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__39_) );
  NOR2_X1 u5_mult_87_U1033 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n220), .ZN(
        u5_mult_87_ab_48__3_) );
  NOR2_X1 u5_mult_87_U1032 ( .A1(u5_mult_87_n367), .A2(u5_mult_87_n220), .ZN(
        u5_mult_87_ab_48__40_) );
  NOR2_X1 u5_mult_87_U1031 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n220), .ZN(
        u5_mult_87_ab_48__41_) );
  NOR2_X1 u5_mult_87_U1030 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n220), .ZN(
        u5_mult_87_ab_48__42_) );
  NOR2_X1 u5_mult_87_U1029 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n220), .ZN(
        u5_mult_87_ab_48__43_) );
  NOR2_X1 u5_mult_87_U1028 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n220), .ZN(
        u5_mult_87_ab_48__44_) );
  NOR2_X1 u5_mult_87_U1027 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n220), .ZN(
        u5_mult_87_ab_48__45_) );
  NOR2_X1 u5_mult_87_U1026 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n220), .ZN(
        u5_mult_87_ab_48__46_) );
  NOR2_X1 u5_mult_87_U1025 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n220), .ZN(
        u5_mult_87_ab_48__47_) );
  NOR2_X1 u5_mult_87_U1024 ( .A1(u5_mult_87_n350), .A2(u5_mult_87_n220), .ZN(
        u5_mult_87_ab_48__48_) );
  NOR2_X1 u5_mult_87_U1023 ( .A1(u5_mult_87_n348), .A2(u5_mult_87_n220), .ZN(
        u5_mult_87_ab_48__49_) );
  NOR2_X1 u5_mult_87_U1022 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n220), .ZN(
        u5_mult_87_ab_48__4_) );
  NOR2_X1 u5_mult_87_U1021 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__50_) );
  NOR2_X1 u5_mult_87_U1020 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__51_) );
  NOR2_X1 u5_mult_87_U1019 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__52_) );
  NOR2_X1 u5_mult_87_U1018 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n221), .ZN(
        u5_mult_87_ab_48__5_) );
  NOR2_X1 u5_mult_87_U1017 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n221), .ZN(
        u5_mult_87_ab_48__6_) );
  NOR2_X1 u5_mult_87_U1016 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n221), .ZN(
        u5_mult_87_ab_48__7_) );
  NOR2_X1 u5_mult_87_U1015 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n221), .ZN(
        u5_mult_87_ab_48__8_) );
  NOR2_X1 u5_mult_87_U1014 ( .A1(u5_mult_87_n430), .A2(u5_mult_87_n219), .ZN(
        u5_mult_87_ab_48__9_) );
  NOR2_X1 u5_mult_87_U1013 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n218), .ZN(
        u5_mult_87_ab_49__0_) );
  NOR2_X1 u5_mult_87_U1012 ( .A1(u5_mult_87_n428), .A2(u5_mult_87_n218), .ZN(
        u5_mult_87_ab_49__10_) );
  NOR2_X1 u5_mult_87_U1011 ( .A1(u5_mult_87_n425), .A2(u5_mult_87_n218), .ZN(
        u5_mult_87_ab_49__11_) );
  NOR2_X1 u5_mult_87_U1010 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n218), .ZN(
        u5_mult_87_ab_49__12_) );
  NOR2_X1 u5_mult_87_U1009 ( .A1(u5_mult_87_n422), .A2(u5_mult_87_n218), .ZN(
        u5_mult_87_ab_49__13_) );
  NOR2_X1 u5_mult_87_U1008 ( .A1(u5_mult_87_n419), .A2(u5_mult_87_n218), .ZN(
        u5_mult_87_ab_49__14_) );
  NOR2_X1 u5_mult_87_U1007 ( .A1(u5_mult_87_n416), .A2(u5_mult_87_n217), .ZN(
        u5_mult_87_ab_49__15_) );
  NOR2_X1 u5_mult_87_U1006 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n218), .ZN(
        u5_mult_87_ab_49__16_) );
  NOR2_X1 u5_mult_87_U1005 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n218), .ZN(
        u5_mult_87_ab_49__17_) );
  NOR2_X1 u5_mult_87_U1004 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n218), .ZN(
        u5_mult_87_ab_49__18_) );
  NOR2_X1 u5_mult_87_U1003 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n218), .ZN(
        u5_mult_87_ab_49__19_) );
  NOR2_X1 u5_mult_87_U1002 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__1_) );
  NOR2_X1 u5_mult_87_U1001 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__20_) );
  NOR2_X1 u5_mult_87_U1000 ( .A1(u5_mult_87_n406), .A2(u5_mult_87_n218), .ZN(
        u5_mult_87_ab_49__21_) );
  NOR2_X1 u5_mult_87_U999 ( .A1(u5_mult_87_n403), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__22_) );
  NOR2_X1 u5_mult_87_U998 ( .A1(u5_mult_87_n402), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__23_) );
  NOR2_X1 u5_mult_87_U997 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__24_) );
  NOR2_X1 u5_mult_87_U996 ( .A1(u5_mult_87_n398), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__25_) );
  NOR2_X1 u5_mult_87_U995 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__26_) );
  NOR2_X1 u5_mult_87_U994 ( .A1(u5_mult_87_n394), .A2(u5_mult_87_n217), .ZN(
        u5_mult_87_ab_49__27_) );
  NOR2_X1 u5_mult_87_U993 ( .A1(u5_mult_87_n391), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__28_) );
  NOR2_X1 u5_mult_87_U992 ( .A1(u5_mult_87_n390), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__29_) );
  NOR2_X1 u5_mult_87_U991 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__2_) );
  NOR2_X1 u5_mult_87_U990 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__30_) );
  NOR2_X1 u5_mult_87_U989 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__31_) );
  NOR2_X1 u5_mult_87_U988 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__32_) );
  NOR2_X1 u5_mult_87_U987 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__33_) );
  NOR2_X1 u5_mult_87_U986 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__34_) );
  NOR2_X1 u5_mult_87_U985 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__35_) );
  NOR2_X1 u5_mult_87_U984 ( .A1(u5_mult_87_n376), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__36_) );
  NOR2_X1 u5_mult_87_U983 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__37_) );
  NOR2_X1 u5_mult_87_U982 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__38_) );
  NOR2_X1 u5_mult_87_U981 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__39_) );
  NOR2_X1 u5_mult_87_U980 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n217), .ZN(
        u5_mult_87_ab_49__3_) );
  NOR2_X1 u5_mult_87_U979 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n217), .ZN(
        u5_mult_87_ab_49__40_) );
  NOR2_X1 u5_mult_87_U978 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n217), .ZN(
        u5_mult_87_ab_49__41_) );
  NOR2_X1 u5_mult_87_U977 ( .A1(u5_mult_87_n362), .A2(u5_mult_87_n217), .ZN(
        u5_mult_87_ab_49__42_) );
  NOR2_X1 u5_mult_87_U976 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n217), .ZN(
        u5_mult_87_ab_49__43_) );
  NOR2_X1 u5_mult_87_U975 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n217), .ZN(
        u5_mult_87_ab_49__44_) );
  NOR2_X1 u5_mult_87_U974 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n217), .ZN(
        u5_mult_87_ab_49__45_) );
  NOR2_X1 u5_mult_87_U973 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n217), .ZN(
        u5_mult_87_ab_49__46_) );
  NOR2_X1 u5_mult_87_U972 ( .A1(u5_mult_87_n352), .A2(u5_mult_87_n217), .ZN(
        u5_mult_87_ab_49__47_) );
  NOR2_X1 u5_mult_87_U971 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n217), .ZN(
        u5_mult_87_ab_49__48_) );
  NOR2_X1 u5_mult_87_U970 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n217), .ZN(
        u5_mult_87_ab_49__49_) );
  NOR2_X1 u5_mult_87_U969 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n217), .ZN(
        u5_mult_87_ab_49__4_) );
  NOR2_X1 u5_mult_87_U968 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__50_) );
  NOR2_X1 u5_mult_87_U967 ( .A1(u5_mult_87_n345), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__51_) );
  NOR2_X1 u5_mult_87_U966 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__52_) );
  NOR2_X1 u5_mult_87_U965 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n218), .ZN(
        u5_mult_87_ab_49__5_) );
  NOR2_X1 u5_mult_87_U964 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n218), .ZN(
        u5_mult_87_ab_49__6_) );
  NOR2_X1 u5_mult_87_U963 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n218), .ZN(
        u5_mult_87_ab_49__7_) );
  NOR2_X1 u5_mult_87_U962 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n218), .ZN(
        u5_mult_87_ab_49__8_) );
  NOR2_X1 u5_mult_87_U961 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n216), .ZN(
        u5_mult_87_ab_49__9_) );
  NOR2_X1 u5_mult_87_U960 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__0_) );
  NOR2_X1 u5_mult_87_U959 ( .A1(u5_mult_87_n428), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__10_) );
  NOR2_X1 u5_mult_87_U958 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__11_) );
  NOR2_X1 u5_mult_87_U957 ( .A1(u5_mult_87_n481), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__12_) );
  NOR2_X1 u5_mult_87_U956 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__13_) );
  NOR2_X1 u5_mult_87_U955 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__14_) );
  NOR2_X1 u5_mult_87_U954 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__15_) );
  NOR2_X1 u5_mult_87_U953 ( .A1(u5_mult_87_n480), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__16_) );
  NOR2_X1 u5_mult_87_U952 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__17_) );
  NOR2_X1 u5_mult_87_U951 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__18_) );
  NOR2_X1 u5_mult_87_U950 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__19_) );
  NOR2_X1 u5_mult_87_U949 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n327), .ZN(
        u5_mult_87_ab_4__1_) );
  NOR2_X1 u5_mult_87_U948 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n327), .ZN(
        u5_mult_87_ab_4__20_) );
  NOR2_X1 u5_mult_87_U947 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n327), .ZN(
        u5_mult_87_ab_4__21_) );
  NOR2_X1 u5_mult_87_U946 ( .A1(u5_mult_87_n404), .A2(u5_mult_87_n327), .ZN(
        u5_mult_87_ab_4__22_) );
  NOR2_X1 u5_mult_87_U945 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n327), .ZN(
        u5_mult_87_ab_4__23_) );
  NOR2_X1 u5_mult_87_U944 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n327), .ZN(
        u5_mult_87_ab_4__24_) );
  NOR2_X1 u5_mult_87_U943 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n327), .ZN(
        u5_mult_87_ab_4__25_) );
  NOR2_X1 u5_mult_87_U942 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n327), .ZN(
        u5_mult_87_ab_4__26_) );
  NOR2_X1 u5_mult_87_U941 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n327), .ZN(
        u5_mult_87_ab_4__27_) );
  NOR2_X1 u5_mult_87_U940 ( .A1(u5_mult_87_n392), .A2(u5_mult_87_n327), .ZN(
        u5_mult_87_ab_4__28_) );
  NOR2_X1 u5_mult_87_U939 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n327), .ZN(
        u5_mult_87_ab_4__29_) );
  NOR2_X1 u5_mult_87_U938 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n328), .ZN(
        u5_mult_87_ab_4__2_) );
  NOR2_X1 u5_mult_87_U937 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n328), .ZN(
        u5_mult_87_ab_4__30_) );
  NOR2_X1 u5_mult_87_U936 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n328), .ZN(
        u5_mult_87_ab_4__31_) );
  NOR2_X1 u5_mult_87_U935 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n328), .ZN(
        u5_mult_87_ab_4__32_) );
  NOR2_X1 u5_mult_87_U934 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n328), .ZN(
        u5_mult_87_ab_4__33_) );
  NOR2_X1 u5_mult_87_U933 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n328), .ZN(
        u5_mult_87_ab_4__34_) );
  NOR2_X1 u5_mult_87_U932 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n328), .ZN(
        u5_mult_87_ab_4__35_) );
  NOR2_X1 u5_mult_87_U931 ( .A1(u5_mult_87_n376), .A2(u5_mult_87_n328), .ZN(
        u5_mult_87_ab_4__36_) );
  NOR2_X1 u5_mult_87_U930 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n328), .ZN(
        u5_mult_87_ab_4__37_) );
  NOR2_X1 u5_mult_87_U929 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n328), .ZN(
        u5_mult_87_ab_4__38_) );
  NOR2_X1 u5_mult_87_U928 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n328), .ZN(
        u5_mult_87_ab_4__39_) );
  NOR2_X1 u5_mult_87_U927 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__3_) );
  NOR2_X1 u5_mult_87_U926 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__40_) );
  NOR2_X1 u5_mult_87_U925 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__41_) );
  NOR2_X1 u5_mult_87_U924 ( .A1(u5_mult_87_n363), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__42_) );
  NOR2_X1 u5_mult_87_U923 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__43_) );
  NOR2_X1 u5_mult_87_U922 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__44_) );
  NOR2_X1 u5_mult_87_U921 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n327), .ZN(
        u5_mult_87_ab_4__45_) );
  NOR2_X1 u5_mult_87_U920 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__46_) );
  NOR2_X1 u5_mult_87_U919 ( .A1(u5_mult_87_n353), .A2(u5_mult_87_n327), .ZN(
        u5_mult_87_ab_4__47_) );
  NOR2_X1 u5_mult_87_U918 ( .A1(u5_mult_87_n350), .A2(u5_mult_87_n327), .ZN(
        u5_mult_87_ab_4__48_) );
  NOR2_X1 u5_mult_87_U917 ( .A1(u5_mult_87_n348), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__49_) );
  NOR2_X1 u5_mult_87_U916 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__4_) );
  NOR2_X1 u5_mult_87_U915 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n328), .ZN(
        u5_mult_87_ab_4__50_) );
  NOR2_X1 u5_mult_87_U914 ( .A1(u5_mult_87_n345), .A2(u5_mult_87_n327), .ZN(
        u5_mult_87_ab_4__51_) );
  NOR2_X1 u5_mult_87_U913 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n327), .ZN(
        u5_mult_87_ab_4__52_) );
  NOR2_X1 u5_mult_87_U912 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__5_) );
  NOR2_X1 u5_mult_87_U911 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__6_) );
  NOR2_X1 u5_mult_87_U910 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__7_) );
  NOR2_X1 u5_mult_87_U909 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__8_) );
  NOR2_X1 u5_mult_87_U908 ( .A1(u5_mult_87_n430), .A2(u5_mult_87_n326), .ZN(
        u5_mult_87_ab_4__9_) );
  NOR2_X1 u5_mult_87_U907 ( .A1(u5_mult_87_n450), .A2(u5_mult_87_n215), .ZN(
        u5_mult_87_ab_50__0_) );
  NOR2_X1 u5_mult_87_U906 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n215), .ZN(
        u5_mult_87_ab_50__10_) );
  NOR2_X1 u5_mult_87_U905 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n215), .ZN(
        u5_mult_87_ab_50__11_) );
  NOR2_X1 u5_mult_87_U904 ( .A1(u5_mult_87_n481), .A2(u5_mult_87_n215), .ZN(
        u5_mult_87_ab_50__12_) );
  NOR2_X1 u5_mult_87_U903 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n215), .ZN(
        u5_mult_87_ab_50__13_) );
  NOR2_X1 u5_mult_87_U902 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n215), .ZN(
        u5_mult_87_ab_50__14_) );
  NOR2_X1 u5_mult_87_U901 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n215), .ZN(
        u5_mult_87_ab_50__15_) );
  NOR2_X1 u5_mult_87_U900 ( .A1(u5_mult_87_n480), .A2(u5_mult_87_n215), .ZN(
        u5_mult_87_ab_50__16_) );
  NOR2_X1 u5_mult_87_U899 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n215), .ZN(
        u5_mult_87_ab_50__17_) );
  NOR2_X1 u5_mult_87_U898 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n215), .ZN(
        u5_mult_87_ab_50__18_) );
  NOR2_X1 u5_mult_87_U897 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n215), .ZN(
        u5_mult_87_ab_50__19_) );
  NOR2_X1 u5_mult_87_U896 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__1_) );
  NOR2_X1 u5_mult_87_U895 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__20_) );
  NOR2_X1 u5_mult_87_U894 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__21_) );
  NOR2_X1 u5_mult_87_U893 ( .A1(u5_mult_87_n404), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__22_) );
  NOR2_X1 u5_mult_87_U892 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__23_) );
  NOR2_X1 u5_mult_87_U891 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__24_) );
  NOR2_X1 u5_mult_87_U890 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__25_) );
  NOR2_X1 u5_mult_87_U889 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__26_) );
  NOR2_X1 u5_mult_87_U888 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__27_) );
  NOR2_X1 u5_mult_87_U887 ( .A1(u5_mult_87_n392), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__28_) );
  NOR2_X1 u5_mult_87_U886 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__29_) );
  NOR2_X1 u5_mult_87_U885 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n214), .ZN(
        u5_mult_87_ab_50__2_) );
  NOR2_X1 u5_mult_87_U884 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n214), .ZN(
        u5_mult_87_ab_50__30_) );
  NOR2_X1 u5_mult_87_U883 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n214), .ZN(
        u5_mult_87_ab_50__31_) );
  NOR2_X1 u5_mult_87_U882 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n214), .ZN(
        u5_mult_87_ab_50__32_) );
  NOR2_X1 u5_mult_87_U881 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n214), .ZN(
        u5_mult_87_ab_50__33_) );
  NOR2_X1 u5_mult_87_U880 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n214), .ZN(
        u5_mult_87_ab_50__34_) );
  NOR2_X1 u5_mult_87_U879 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n214), .ZN(
        u5_mult_87_ab_50__35_) );
  NOR2_X1 u5_mult_87_U878 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n214), .ZN(
        u5_mult_87_ab_50__36_) );
  NOR2_X1 u5_mult_87_U877 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n214), .ZN(
        u5_mult_87_ab_50__37_) );
  NOR2_X1 u5_mult_87_U876 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n214), .ZN(
        u5_mult_87_ab_50__38_) );
  NOR2_X1 u5_mult_87_U875 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n214), .ZN(
        u5_mult_87_ab_50__39_) );
  NOR2_X1 u5_mult_87_U874 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__3_) );
  NOR2_X1 u5_mult_87_U873 ( .A1(u5_mult_87_n367), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__40_) );
  NOR2_X1 u5_mult_87_U872 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__41_) );
  NOR2_X1 u5_mult_87_U871 ( .A1(u5_mult_87_n363), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__42_) );
  NOR2_X1 u5_mult_87_U870 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__43_) );
  NOR2_X1 u5_mult_87_U869 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__44_) );
  NOR2_X1 u5_mult_87_U868 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__45_) );
  NOR2_X1 u5_mult_87_U867 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__46_) );
  NOR2_X1 u5_mult_87_U866 ( .A1(u5_mult_87_n353), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__47_) );
  NOR2_X1 u5_mult_87_U865 ( .A1(u5_mult_87_n350), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__48_) );
  NOR2_X1 u5_mult_87_U864 ( .A1(u5_mult_87_n348), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__49_) );
  NOR2_X1 u5_mult_87_U863 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n214), .ZN(
        u5_mult_87_ab_50__4_) );
  NOR2_X1 u5_mult_87_U862 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__50_) );
  NOR2_X1 u5_mult_87_U861 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__51_) );
  NOR2_X1 u5_mult_87_U860 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__52_) );
  NOR2_X1 u5_mult_87_U859 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n215), .ZN(
        u5_mult_87_ab_50__5_) );
  NOR2_X1 u5_mult_87_U858 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n215), .ZN(
        u5_mult_87_ab_50__6_) );
  NOR2_X1 u5_mult_87_U857 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__7_) );
  NOR2_X1 u5_mult_87_U856 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__8_) );
  NOR2_X1 u5_mult_87_U855 ( .A1(u5_mult_87_n430), .A2(u5_mult_87_n213), .ZN(
        u5_mult_87_ab_50__9_) );
  NOR2_X1 u5_mult_87_U854 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n210), .ZN(
        u5_mult_87_ab_51__0_) );
  NOR2_X1 u5_mult_87_U853 ( .A1(u5_mult_87_n428), .A2(u5_mult_87_n210), .ZN(
        u5_mult_87_ab_51__10_) );
  NOR2_X1 u5_mult_87_U852 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n210), .ZN(
        u5_mult_87_ab_51__11_) );
  NOR2_X1 u5_mult_87_U851 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n210), .ZN(
        u5_mult_87_ab_51__12_) );
  NOR2_X1 u5_mult_87_U850 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n210), .ZN(
        u5_mult_87_ab_51__13_) );
  NOR2_X1 u5_mult_87_U849 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n210), .ZN(
        u5_mult_87_ab_51__14_) );
  NOR2_X1 u5_mult_87_U848 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n210), .ZN(
        u5_mult_87_ab_51__15_) );
  NOR2_X1 u5_mult_87_U847 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n210), .ZN(
        u5_mult_87_ab_51__16_) );
  NOR2_X1 u5_mult_87_U846 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n210), .ZN(
        u5_mult_87_ab_51__17_) );
  NOR2_X1 u5_mult_87_U845 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n210), .ZN(
        u5_mult_87_ab_51__18_) );
  NOR2_X1 u5_mult_87_U844 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n210), .ZN(
        u5_mult_87_ab_51__19_) );
  NOR2_X1 u5_mult_87_U843 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n211), .ZN(
        u5_mult_87_ab_51__1_) );
  NOR2_X1 u5_mult_87_U842 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n211), .ZN(
        u5_mult_87_ab_51__20_) );
  NOR2_X1 u5_mult_87_U841 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n211), .ZN(
        u5_mult_87_ab_51__21_) );
  NOR2_X1 u5_mult_87_U840 ( .A1(u5_mult_87_n404), .A2(u5_mult_87_n211), .ZN(
        u5_mult_87_ab_51__22_) );
  NOR2_X1 u5_mult_87_U839 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n211), .ZN(
        u5_mult_87_ab_51__23_) );
  NOR2_X1 u5_mult_87_U838 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n211), .ZN(
        u5_mult_87_ab_51__24_) );
  NOR2_X1 u5_mult_87_U837 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n211), .ZN(
        u5_mult_87_ab_51__25_) );
  NOR2_X1 u5_mult_87_U836 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n211), .ZN(
        u5_mult_87_ab_51__26_) );
  NOR2_X1 u5_mult_87_U835 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n211), .ZN(
        u5_mult_87_ab_51__27_) );
  NOR2_X1 u5_mult_87_U834 ( .A1(u5_mult_87_n392), .A2(u5_mult_87_n211), .ZN(
        u5_mult_87_ab_51__28_) );
  NOR2_X1 u5_mult_87_U833 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n211), .ZN(
        u5_mult_87_ab_51__29_) );
  NOR2_X1 u5_mult_87_U832 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n212), .ZN(
        u5_mult_87_ab_51__2_) );
  NOR2_X1 u5_mult_87_U831 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n212), .ZN(
        u5_mult_87_ab_51__30_) );
  NOR2_X1 u5_mult_87_U830 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n212), .ZN(
        u5_mult_87_ab_51__31_) );
  NOR2_X1 u5_mult_87_U829 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n212), .ZN(
        u5_mult_87_ab_51__32_) );
  NOR2_X1 u5_mult_87_U828 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n212), .ZN(
        u5_mult_87_ab_51__33_) );
  NOR2_X1 u5_mult_87_U827 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n212), .ZN(
        u5_mult_87_ab_51__34_) );
  NOR2_X1 u5_mult_87_U826 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n212), .ZN(
        u5_mult_87_ab_51__35_) );
  NOR2_X1 u5_mult_87_U825 ( .A1(u5_mult_87_n376), .A2(u5_mult_87_n212), .ZN(
        u5_mult_87_ab_51__36_) );
  NOR2_X1 u5_mult_87_U824 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n212), .ZN(
        u5_mult_87_ab_51__37_) );
  NOR2_X1 u5_mult_87_U823 ( .A1(u5_mult_87_n372), .A2(u5_mult_87_n212), .ZN(
        u5_mult_87_ab_51__38_) );
  NOR2_X1 u5_mult_87_U822 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n212), .ZN(
        u5_mult_87_ab_51__39_) );
  NOR2_X1 u5_mult_87_U821 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n211), .ZN(
        u5_mult_87_ab_51__3_) );
  NOR2_X1 u5_mult_87_U820 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n210), .ZN(
        u5_mult_87_ab_51__40_) );
  NOR2_X1 u5_mult_87_U819 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n210), .ZN(
        u5_mult_87_ab_51__41_) );
  NOR2_X1 u5_mult_87_U818 ( .A1(u5_mult_87_n363), .A2(u5_mult_87_n211), .ZN(
        u5_mult_87_ab_51__42_) );
  NOR2_X1 u5_mult_87_U817 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n211), .ZN(
        u5_mult_87_ab_51__43_) );
  NOR2_X1 u5_mult_87_U816 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n210), .ZN(
        u5_mult_87_ab_51__44_) );
  NOR2_X1 u5_mult_87_U815 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n210), .ZN(
        u5_mult_87_ab_51__45_) );
  NOR2_X1 u5_mult_87_U814 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n211), .ZN(
        u5_mult_87_ab_51__46_) );
  NOR2_X1 u5_mult_87_U813 ( .A1(u5_mult_87_n353), .A2(u5_mult_87_n212), .ZN(
        u5_mult_87_ab_51__47_) );
  NOR2_X1 u5_mult_87_U812 ( .A1(u5_mult_87_n349), .A2(u5_mult_87_n210), .ZN(
        u5_mult_87_ab_51__48_) );
  NOR2_X1 u5_mult_87_U811 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n212), .ZN(
        u5_mult_87_ab_51__49_) );
  NOR2_X1 u5_mult_87_U810 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n212), .ZN(
        u5_mult_87_ab_51__4_) );
  NOR2_X1 u5_mult_87_U809 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n210), .ZN(
        u5_mult_87_ab_51__50_) );
  NOR2_X1 u5_mult_87_U808 ( .A1(u5_mult_87_n345), .A2(u5_mult_87_n210), .ZN(
        u5_mult_87_ab_51__51_) );
  NOR2_X1 u5_mult_87_U807 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n211), .ZN(
        u5_mult_87_ab_51__52_) );
  NOR2_X1 u5_mult_87_U806 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n210), .ZN(
        u5_mult_87_ab_51__5_) );
  NOR2_X1 u5_mult_87_U805 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n210), .ZN(
        u5_mult_87_ab_51__6_) );
  NOR2_X1 u5_mult_87_U804 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n210), .ZN(
        u5_mult_87_ab_51__7_) );
  NOR2_X1 u5_mult_87_U803 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n210), .ZN(
        u5_mult_87_ab_51__8_) );
  NOR2_X1 u5_mult_87_U802 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n210), .ZN(
        u5_mult_87_ab_51__9_) );
  NOR2_X1 u5_mult_87_U801 ( .A1(u5_mult_87_n450), .A2(u5_mult_87_n453), .ZN(
        u5_mult_87_ab_52__0_) );
  NOR2_X1 u5_mult_87_U800 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n453), .ZN(
        u5_mult_87_ab_52__10_) );
  NOR2_X1 u5_mult_87_U799 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n453), .ZN(
        u5_mult_87_ab_52__11_) );
  NOR2_X1 u5_mult_87_U798 ( .A1(u5_mult_87_n481), .A2(u5_mult_87_n453), .ZN(
        u5_mult_87_ab_52__12_) );
  NOR2_X1 u5_mult_87_U797 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n453), .ZN(
        u5_mult_87_ab_52__13_) );
  NOR2_X1 u5_mult_87_U796 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n453), .ZN(
        u5_mult_87_ab_52__14_) );
  NOR2_X1 u5_mult_87_U795 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n453), .ZN(
        u5_mult_87_ab_52__15_) );
  NOR2_X1 u5_mult_87_U794 ( .A1(u5_mult_87_n480), .A2(u5_mult_87_n453), .ZN(
        u5_mult_87_ab_52__16_) );
  NOR2_X1 u5_mult_87_U793 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n451), .ZN(
        u5_mult_87_ab_52__17_) );
  NOR2_X1 u5_mult_87_U792 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n453), .ZN(
        u5_mult_87_ab_52__18_) );
  NOR2_X1 u5_mult_87_U791 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n453), .ZN(
        u5_mult_87_ab_52__19_) );
  NOR2_X1 u5_mult_87_U790 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n453), .ZN(
        u5_mult_87_ab_52__1_) );
  NOR2_X1 u5_mult_87_U789 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n453), .ZN(
        u5_mult_87_ab_52__20_) );
  NOR2_X1 u5_mult_87_U788 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n453), .ZN(
        u5_mult_87_ab_52__21_) );
  NOR2_X1 u5_mult_87_U787 ( .A1(u5_mult_87_n404), .A2(u5_mult_87_n453), .ZN(
        u5_mult_87_ab_52__22_) );
  NOR2_X1 u5_mult_87_U786 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n453), .ZN(
        u5_mult_87_ab_52__23_) );
  NOR2_X1 u5_mult_87_U785 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n453), .ZN(
        u5_mult_87_ab_52__24_) );
  NOR2_X1 u5_mult_87_U784 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n453), .ZN(
        u5_mult_87_ab_52__25_) );
  NOR2_X1 u5_mult_87_U783 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n453), .ZN(
        u5_mult_87_ab_52__26_) );
  NOR2_X1 u5_mult_87_U782 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n453), .ZN(
        u5_mult_87_ab_52__27_) );
  NOR2_X1 u5_mult_87_U781 ( .A1(u5_mult_87_n392), .A2(u5_mult_87_n452), .ZN(
        u5_mult_87_ab_52__28_) );
  NOR2_X1 u5_mult_87_U780 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n452), .ZN(
        u5_mult_87_ab_52__29_) );
  NOR2_X1 u5_mult_87_U779 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n452), .ZN(
        u5_mult_87_ab_52__2_) );
  NOR2_X1 u5_mult_87_U778 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n452), .ZN(
        u5_mult_87_ab_52__30_) );
  NOR2_X1 u5_mult_87_U777 ( .A1(u5_mult_87_n385), .A2(u5_mult_87_n452), .ZN(
        u5_mult_87_ab_52__31_) );
  NOR2_X1 u5_mult_87_U776 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n452), .ZN(
        u5_mult_87_ab_52__32_) );
  NOR2_X1 u5_mult_87_U775 ( .A1(u5_mult_87_n381), .A2(u5_mult_87_n452), .ZN(
        u5_mult_87_ab_52__33_) );
  NOR2_X1 u5_mult_87_U774 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n452), .ZN(
        u5_mult_87_ab_52__34_) );
  NOR2_X1 u5_mult_87_U773 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n452), .ZN(
        u5_mult_87_ab_52__35_) );
  NOR2_X1 u5_mult_87_U772 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n452), .ZN(
        u5_mult_87_ab_52__36_) );
  NOR2_X1 u5_mult_87_U771 ( .A1(u5_mult_87_n373), .A2(u5_mult_87_n452), .ZN(
        u5_mult_87_ab_52__37_) );
  NOR2_X1 u5_mult_87_U770 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n451), .ZN(
        u5_mult_87_ab_52__38_) );
  NOR2_X1 u5_mult_87_U769 ( .A1(u5_mult_87_n369), .A2(u5_mult_87_n451), .ZN(
        u5_mult_87_ab_52__39_) );
  NOR2_X1 u5_mult_87_U768 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n451), .ZN(
        u5_mult_87_ab_52__3_) );
  NOR2_X1 u5_mult_87_U767 ( .A1(u5_mult_87_n367), .A2(u5_mult_87_n451), .ZN(
        u5_mult_87_ab_52__40_) );
  NOR2_X1 u5_mult_87_U766 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n451), .ZN(
        u5_mult_87_ab_52__41_) );
  NOR2_X1 u5_mult_87_U765 ( .A1(u5_mult_87_n363), .A2(u5_mult_87_n451), .ZN(
        u5_mult_87_ab_52__42_) );
  NOR2_X1 u5_mult_87_U764 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n451), .ZN(
        u5_mult_87_ab_52__43_) );
  NOR2_X1 u5_mult_87_U763 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n452), .ZN(
        u5_mult_87_ab_52__44_) );
  NOR2_X1 u5_mult_87_U762 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n452), .ZN(
        u5_mult_87_ab_52__45_) );
  NOR2_X1 u5_mult_87_U761 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n452), .ZN(
        u5_mult_87_ab_52__46_) );
  NOR2_X1 u5_mult_87_U760 ( .A1(u5_mult_87_n353), .A2(u5_mult_87_n452), .ZN(
        u5_mult_87_ab_52__47_) );
  NOR2_X1 u5_mult_87_U759 ( .A1(u5_mult_87_n350), .A2(u5_mult_87_n451), .ZN(
        u5_mult_87_ab_52__48_) );
  NOR2_X1 u5_mult_87_U758 ( .A1(u5_mult_87_n348), .A2(u5_mult_87_n451), .ZN(
        u5_mult_87_ab_52__49_) );
  NOR2_X1 u5_mult_87_U757 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n451), .ZN(
        u5_mult_87_ab_52__4_) );
  NOR2_X1 u5_mult_87_U756 ( .A1(u5_mult_87_n346), .A2(u5_mult_87_n451), .ZN(
        u5_mult_87_ab_52__50_) );
  NOR2_X1 u5_mult_87_U755 ( .A1(u5_mult_87_n344), .A2(u5_mult_87_n451), .ZN(
        u5_mult_87_ab_52__51_) );
  NOR2_X1 u5_mult_87_U754 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n451), .ZN(
        u5_mult_87_ab_52__52_) );
  NOR2_X1 u5_mult_87_U753 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n451), .ZN(
        u5_mult_87_ab_52__5_) );
  NOR2_X1 u5_mult_87_U752 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n451), .ZN(
        u5_mult_87_ab_52__6_) );
  NOR2_X1 u5_mult_87_U751 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n451), .ZN(
        u5_mult_87_ab_52__7_) );
  NOR2_X1 u5_mult_87_U750 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n451), .ZN(
        u5_mult_87_ab_52__8_) );
  NOR2_X1 u5_mult_87_U749 ( .A1(u5_mult_87_n430), .A2(u5_mult_87_n451), .ZN(
        u5_mult_87_ab_52__9_) );
  NOR2_X1 u5_mult_87_U748 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__0_) );
  NOR2_X1 u5_mult_87_U747 ( .A1(u5_mult_87_n428), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__10_) );
  NOR2_X1 u5_mult_87_U746 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__11_) );
  NOR2_X1 u5_mult_87_U745 ( .A1(u5_mult_87_n481), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__12_) );
  NOR2_X1 u5_mult_87_U744 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__13_) );
  NOR2_X1 u5_mult_87_U743 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__14_) );
  NOR2_X1 u5_mult_87_U742 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__15_) );
  NOR2_X1 u5_mult_87_U741 ( .A1(u5_mult_87_n480), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__16_) );
  NOR2_X1 u5_mult_87_U740 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__17_) );
  NOR2_X1 u5_mult_87_U739 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__18_) );
  NOR2_X1 u5_mult_87_U738 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__19_) );
  NOR2_X1 u5_mult_87_U737 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n324), .ZN(
        u5_mult_87_ab_5__1_) );
  NOR2_X1 u5_mult_87_U736 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n324), .ZN(
        u5_mult_87_ab_5__20_) );
  NOR2_X1 u5_mult_87_U735 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n324), .ZN(
        u5_mult_87_ab_5__21_) );
  NOR2_X1 u5_mult_87_U734 ( .A1(u5_mult_87_n404), .A2(u5_mult_87_n324), .ZN(
        u5_mult_87_ab_5__22_) );
  NOR2_X1 u5_mult_87_U733 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n324), .ZN(
        u5_mult_87_ab_5__23_) );
  NOR2_X1 u5_mult_87_U732 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n324), .ZN(
        u5_mult_87_ab_5__24_) );
  NOR2_X1 u5_mult_87_U731 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n324), .ZN(
        u5_mult_87_ab_5__25_) );
  NOR2_X1 u5_mult_87_U730 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n324), .ZN(
        u5_mult_87_ab_5__26_) );
  NOR2_X1 u5_mult_87_U729 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n324), .ZN(
        u5_mult_87_ab_5__27_) );
  NOR2_X1 u5_mult_87_U728 ( .A1(u5_mult_87_n392), .A2(u5_mult_87_n324), .ZN(
        u5_mult_87_ab_5__28_) );
  NOR2_X1 u5_mult_87_U727 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n324), .ZN(
        u5_mult_87_ab_5__29_) );
  NOR2_X1 u5_mult_87_U726 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n325), .ZN(
        u5_mult_87_ab_5__2_) );
  NOR2_X1 u5_mult_87_U725 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n325), .ZN(
        u5_mult_87_ab_5__30_) );
  NOR2_X1 u5_mult_87_U724 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n325), .ZN(
        u5_mult_87_ab_5__31_) );
  NOR2_X1 u5_mult_87_U723 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n325), .ZN(
        u5_mult_87_ab_5__32_) );
  NOR2_X1 u5_mult_87_U722 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n325), .ZN(
        u5_mult_87_ab_5__33_) );
  NOR2_X1 u5_mult_87_U721 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n325), .ZN(
        u5_mult_87_ab_5__34_) );
  NOR2_X1 u5_mult_87_U720 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n325), .ZN(
        u5_mult_87_ab_5__35_) );
  NOR2_X1 u5_mult_87_U719 ( .A1(u5_mult_87_n376), .A2(u5_mult_87_n325), .ZN(
        u5_mult_87_ab_5__36_) );
  NOR2_X1 u5_mult_87_U718 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n325), .ZN(
        u5_mult_87_ab_5__37_) );
  NOR2_X1 u5_mult_87_U717 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n325), .ZN(
        u5_mult_87_ab_5__38_) );
  NOR2_X1 u5_mult_87_U716 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n325), .ZN(
        u5_mult_87_ab_5__39_) );
  NOR2_X1 u5_mult_87_U715 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n325), .ZN(
        u5_mult_87_ab_5__3_) );
  NOR2_X1 u5_mult_87_U714 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n325), .ZN(
        u5_mult_87_ab_5__40_) );
  NOR2_X1 u5_mult_87_U713 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__41_) );
  NOR2_X1 u5_mult_87_U712 ( .A1(u5_mult_87_n363), .A2(u5_mult_87_n325), .ZN(
        u5_mult_87_ab_5__42_) );
  NOR2_X1 u5_mult_87_U711 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__43_) );
  NOR2_X1 u5_mult_87_U710 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__44_) );
  NOR2_X1 u5_mult_87_U709 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__45_) );
  NOR2_X1 u5_mult_87_U708 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__46_) );
  NOR2_X1 u5_mult_87_U707 ( .A1(u5_mult_87_n353), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__47_) );
  NOR2_X1 u5_mult_87_U706 ( .A1(u5_mult_87_n350), .A2(u5_mult_87_n324), .ZN(
        u5_mult_87_ab_5__48_) );
  NOR2_X1 u5_mult_87_U705 ( .A1(u5_mult_87_n348), .A2(u5_mult_87_n324), .ZN(
        u5_mult_87_ab_5__49_) );
  NOR2_X1 u5_mult_87_U704 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__4_) );
  NOR2_X1 u5_mult_87_U703 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n325), .ZN(
        u5_mult_87_ab_5__50_) );
  NOR2_X1 u5_mult_87_U702 ( .A1(u5_mult_87_n345), .A2(u5_mult_87_n324), .ZN(
        u5_mult_87_ab_5__51_) );
  NOR2_X1 u5_mult_87_U701 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__52_) );
  NOR2_X1 u5_mult_87_U700 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__5_) );
  NOR2_X1 u5_mult_87_U699 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__6_) );
  NOR2_X1 u5_mult_87_U698 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__7_) );
  NOR2_X1 u5_mult_87_U697 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__8_) );
  NOR2_X1 u5_mult_87_U696 ( .A1(u5_mult_87_n430), .A2(u5_mult_87_n323), .ZN(
        u5_mult_87_ab_5__9_) );
  NOR2_X1 u5_mult_87_U695 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__0_) );
  NOR2_X1 u5_mult_87_U694 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__10_) );
  NOR2_X1 u5_mult_87_U693 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__11_) );
  NOR2_X1 u5_mult_87_U692 ( .A1(u5_mult_87_n481), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__12_) );
  NOR2_X1 u5_mult_87_U691 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__13_) );
  NOR2_X1 u5_mult_87_U690 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__14_) );
  NOR2_X1 u5_mult_87_U689 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__15_) );
  NOR2_X1 u5_mult_87_U688 ( .A1(u5_mult_87_n480), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__16_) );
  NOR2_X1 u5_mult_87_U687 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__17_) );
  NOR2_X1 u5_mult_87_U686 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__18_) );
  NOR2_X1 u5_mult_87_U685 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__19_) );
  NOR2_X1 u5_mult_87_U684 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__1_) );
  NOR2_X1 u5_mult_87_U683 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__20_) );
  NOR2_X1 u5_mult_87_U682 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__21_) );
  NOR2_X1 u5_mult_87_U681 ( .A1(u5_mult_87_n404), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__22_) );
  NOR2_X1 u5_mult_87_U680 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__23_) );
  NOR2_X1 u5_mult_87_U679 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__24_) );
  NOR2_X1 u5_mult_87_U678 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__25_) );
  NOR2_X1 u5_mult_87_U677 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__26_) );
  NOR2_X1 u5_mult_87_U676 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__27_) );
  NOR2_X1 u5_mult_87_U675 ( .A1(u5_mult_87_n392), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__28_) );
  NOR2_X1 u5_mult_87_U674 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__29_) );
  NOR2_X1 u5_mult_87_U673 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__2_) );
  NOR2_X1 u5_mult_87_U672 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__30_) );
  NOR2_X1 u5_mult_87_U671 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__31_) );
  NOR2_X1 u5_mult_87_U670 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__32_) );
  NOR2_X1 u5_mult_87_U669 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__33_) );
  NOR2_X1 u5_mult_87_U668 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__34_) );
  NOR2_X1 u5_mult_87_U667 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__35_) );
  NOR2_X1 u5_mult_87_U666 ( .A1(u5_mult_87_n376), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__36_) );
  NOR2_X1 u5_mult_87_U665 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__37_) );
  NOR2_X1 u5_mult_87_U664 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__38_) );
  NOR2_X1 u5_mult_87_U663 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__39_) );
  NOR2_X1 u5_mult_87_U662 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n322), .ZN(
        u5_mult_87_ab_6__3_) );
  NOR2_X1 u5_mult_87_U661 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n322), .ZN(
        u5_mult_87_ab_6__40_) );
  NOR2_X1 u5_mult_87_U660 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n322), .ZN(
        u5_mult_87_ab_6__41_) );
  NOR2_X1 u5_mult_87_U659 ( .A1(u5_mult_87_n363), .A2(u5_mult_87_n322), .ZN(
        u5_mult_87_ab_6__42_) );
  NOR2_X1 u5_mult_87_U658 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n322), .ZN(
        u5_mult_87_ab_6__43_) );
  NOR2_X1 u5_mult_87_U657 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n322), .ZN(
        u5_mult_87_ab_6__44_) );
  NOR2_X1 u5_mult_87_U656 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n322), .ZN(
        u5_mult_87_ab_6__45_) );
  NOR2_X1 u5_mult_87_U655 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n322), .ZN(
        u5_mult_87_ab_6__46_) );
  NOR2_X1 u5_mult_87_U654 ( .A1(u5_mult_87_n353), .A2(u5_mult_87_n322), .ZN(
        u5_mult_87_ab_6__47_) );
  NOR2_X1 u5_mult_87_U653 ( .A1(u5_mult_87_n350), .A2(u5_mult_87_n322), .ZN(
        u5_mult_87_ab_6__48_) );
  NOR2_X1 u5_mult_87_U652 ( .A1(u5_mult_87_n348), .A2(u5_mult_87_n322), .ZN(
        u5_mult_87_ab_6__49_) );
  NOR2_X1 u5_mult_87_U651 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__4_) );
  NOR2_X1 u5_mult_87_U650 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n322), .ZN(
        u5_mult_87_ab_6__50_) );
  NOR2_X1 u5_mult_87_U649 ( .A1(u5_mult_87_n345), .A2(u5_mult_87_n322), .ZN(
        u5_mult_87_ab_6__51_) );
  NOR2_X1 u5_mult_87_U648 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__52_) );
  NOR2_X1 u5_mult_87_U647 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__5_) );
  NOR2_X1 u5_mult_87_U646 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__6_) );
  NOR2_X1 u5_mult_87_U645 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__7_) );
  NOR2_X1 u5_mult_87_U644 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__8_) );
  NOR2_X1 u5_mult_87_U643 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n321), .ZN(
        u5_mult_87_ab_6__9_) );
  NOR2_X1 u5_mult_87_U642 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__0_) );
  NOR2_X1 u5_mult_87_U641 ( .A1(u5_mult_87_n428), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__10_) );
  NOR2_X1 u5_mult_87_U640 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__11_) );
  NOR2_X1 u5_mult_87_U639 ( .A1(u5_mult_87_n481), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__12_) );
  NOR2_X1 u5_mult_87_U638 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__13_) );
  NOR2_X1 u5_mult_87_U637 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__14_) );
  NOR2_X1 u5_mult_87_U636 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__15_) );
  NOR2_X1 u5_mult_87_U635 ( .A1(u5_mult_87_n480), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__16_) );
  NOR2_X1 u5_mult_87_U634 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__17_) );
  NOR2_X1 u5_mult_87_U633 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__18_) );
  NOR2_X1 u5_mult_87_U632 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__19_) );
  NOR2_X1 u5_mult_87_U631 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__1_) );
  NOR2_X1 u5_mult_87_U630 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__20_) );
  NOR2_X1 u5_mult_87_U629 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__21_) );
  NOR2_X1 u5_mult_87_U628 ( .A1(u5_mult_87_n404), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__22_) );
  NOR2_X1 u5_mult_87_U627 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__23_) );
  NOR2_X1 u5_mult_87_U626 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__24_) );
  NOR2_X1 u5_mult_87_U625 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__25_) );
  NOR2_X1 u5_mult_87_U624 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__26_) );
  NOR2_X1 u5_mult_87_U623 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__27_) );
  NOR2_X1 u5_mult_87_U622 ( .A1(u5_mult_87_n392), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__28_) );
  NOR2_X1 u5_mult_87_U621 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__29_) );
  NOR2_X1 u5_mult_87_U620 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__2_) );
  NOR2_X1 u5_mult_87_U619 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__30_) );
  NOR2_X1 u5_mult_87_U618 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__31_) );
  NOR2_X1 u5_mult_87_U617 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__32_) );
  NOR2_X1 u5_mult_87_U616 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__33_) );
  NOR2_X1 u5_mult_87_U615 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__34_) );
  NOR2_X1 u5_mult_87_U614 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__35_) );
  NOR2_X1 u5_mult_87_U613 ( .A1(u5_mult_87_n376), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__36_) );
  NOR2_X1 u5_mult_87_U612 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__37_) );
  NOR2_X1 u5_mult_87_U611 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__38_) );
  NOR2_X1 u5_mult_87_U610 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__39_) );
  NOR2_X1 u5_mult_87_U609 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n320), .ZN(
        u5_mult_87_ab_7__3_) );
  NOR2_X1 u5_mult_87_U608 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__40_) );
  NOR2_X1 u5_mult_87_U607 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__41_) );
  NOR2_X1 u5_mult_87_U606 ( .A1(u5_mult_87_n363), .A2(u5_mult_87_n320), .ZN(
        u5_mult_87_ab_7__42_) );
  NOR2_X1 u5_mult_87_U605 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n320), .ZN(
        u5_mult_87_ab_7__43_) );
  NOR2_X1 u5_mult_87_U604 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n320), .ZN(
        u5_mult_87_ab_7__44_) );
  NOR2_X1 u5_mult_87_U603 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n320), .ZN(
        u5_mult_87_ab_7__45_) );
  NOR2_X1 u5_mult_87_U602 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n320), .ZN(
        u5_mult_87_ab_7__46_) );
  NOR2_X1 u5_mult_87_U601 ( .A1(u5_mult_87_n353), .A2(u5_mult_87_n320), .ZN(
        u5_mult_87_ab_7__47_) );
  NOR2_X1 u5_mult_87_U600 ( .A1(u5_mult_87_n350), .A2(u5_mult_87_n320), .ZN(
        u5_mult_87_ab_7__48_) );
  NOR2_X1 u5_mult_87_U599 ( .A1(u5_mult_87_n348), .A2(u5_mult_87_n320), .ZN(
        u5_mult_87_ab_7__49_) );
  NOR2_X1 u5_mult_87_U598 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__4_) );
  NOR2_X1 u5_mult_87_U597 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n320), .ZN(
        u5_mult_87_ab_7__50_) );
  NOR2_X1 u5_mult_87_U596 ( .A1(u5_mult_87_n345), .A2(u5_mult_87_n320), .ZN(
        u5_mult_87_ab_7__51_) );
  NOR2_X1 u5_mult_87_U595 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n320), .ZN(
        u5_mult_87_ab_7__52_) );
  NOR2_X1 u5_mult_87_U594 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__5_) );
  NOR2_X1 u5_mult_87_U593 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n320), .ZN(
        u5_mult_87_ab_7__6_) );
  NOR2_X1 u5_mult_87_U592 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__7_) );
  NOR2_X1 u5_mult_87_U591 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n320), .ZN(
        u5_mult_87_ab_7__8_) );
  NOR2_X1 u5_mult_87_U590 ( .A1(u5_mult_87_n430), .A2(u5_mult_87_n319), .ZN(
        u5_mult_87_ab_7__9_) );
  NOR2_X1 u5_mult_87_U589 ( .A1(u5_mult_87_n449), .A2(u5_mult_87_n315), .ZN(
        u5_mult_87_ab_8__0_) );
  NOR2_X1 u5_mult_87_U588 ( .A1(u5_mult_87_n427), .A2(u5_mult_87_n315), .ZN(
        u5_mult_87_ab_8__10_) );
  NOR2_X1 u5_mult_87_U587 ( .A1(u5_mult_87_n426), .A2(u5_mult_87_n315), .ZN(
        u5_mult_87_ab_8__11_) );
  NOR2_X1 u5_mult_87_U586 ( .A1(u5_mult_87_n424), .A2(u5_mult_87_n315), .ZN(
        u5_mult_87_ab_8__12_) );
  NOR2_X1 u5_mult_87_U585 ( .A1(u5_mult_87_n423), .A2(u5_mult_87_n315), .ZN(
        u5_mult_87_ab_8__13_) );
  NOR2_X1 u5_mult_87_U584 ( .A1(u5_mult_87_n420), .A2(u5_mult_87_n315), .ZN(
        u5_mult_87_ab_8__14_) );
  NOR2_X1 u5_mult_87_U583 ( .A1(u5_mult_87_n417), .A2(u5_mult_87_n315), .ZN(
        u5_mult_87_ab_8__15_) );
  NOR2_X1 u5_mult_87_U582 ( .A1(u5_mult_87_n415), .A2(u5_mult_87_n315), .ZN(
        u5_mult_87_ab_8__16_) );
  NOR2_X1 u5_mult_87_U581 ( .A1(u5_mult_87_n414), .A2(u5_mult_87_n315), .ZN(
        u5_mult_87_ab_8__17_) );
  NOR2_X1 u5_mult_87_U580 ( .A1(u5_mult_87_n412), .A2(u5_mult_87_n315), .ZN(
        u5_mult_87_ab_8__18_) );
  NOR2_X1 u5_mult_87_U579 ( .A1(u5_mult_87_n410), .A2(u5_mult_87_n315), .ZN(
        u5_mult_87_ab_8__19_) );
  NOR2_X1 u5_mult_87_U578 ( .A1(u5_mult_87_n448), .A2(u5_mult_87_n316), .ZN(
        u5_mult_87_ab_8__1_) );
  NOR2_X1 u5_mult_87_U577 ( .A1(u5_mult_87_n408), .A2(u5_mult_87_n316), .ZN(
        u5_mult_87_ab_8__20_) );
  NOR2_X1 u5_mult_87_U576 ( .A1(u5_mult_87_n405), .A2(u5_mult_87_n316), .ZN(
        u5_mult_87_ab_8__21_) );
  NOR2_X1 u5_mult_87_U575 ( .A1(u5_mult_87_n404), .A2(u5_mult_87_n316), .ZN(
        u5_mult_87_ab_8__22_) );
  NOR2_X1 u5_mult_87_U574 ( .A1(u5_mult_87_n401), .A2(u5_mult_87_n316), .ZN(
        u5_mult_87_ab_8__23_) );
  NOR2_X1 u5_mult_87_U573 ( .A1(u5_mult_87_n400), .A2(u5_mult_87_n316), .ZN(
        u5_mult_87_ab_8__24_) );
  NOR2_X1 u5_mult_87_U572 ( .A1(u5_mult_87_n397), .A2(u5_mult_87_n316), .ZN(
        u5_mult_87_ab_8__25_) );
  NOR2_X1 u5_mult_87_U571 ( .A1(u5_mult_87_n396), .A2(u5_mult_87_n316), .ZN(
        u5_mult_87_ab_8__26_) );
  NOR2_X1 u5_mult_87_U570 ( .A1(u5_mult_87_n393), .A2(u5_mult_87_n316), .ZN(
        u5_mult_87_ab_8__27_) );
  NOR2_X1 u5_mult_87_U569 ( .A1(u5_mult_87_n392), .A2(u5_mult_87_n316), .ZN(
        u5_mult_87_ab_8__28_) );
  NOR2_X1 u5_mult_87_U568 ( .A1(u5_mult_87_n389), .A2(u5_mult_87_n316), .ZN(
        u5_mult_87_ab_8__29_) );
  NOR2_X1 u5_mult_87_U567 ( .A1(u5_mult_87_n445), .A2(u5_mult_87_n317), .ZN(
        u5_mult_87_ab_8__2_) );
  NOR2_X1 u5_mult_87_U566 ( .A1(u5_mult_87_n388), .A2(u5_mult_87_n317), .ZN(
        u5_mult_87_ab_8__30_) );
  NOR2_X1 u5_mult_87_U565 ( .A1(u5_mult_87_n386), .A2(u5_mult_87_n317), .ZN(
        u5_mult_87_ab_8__31_) );
  NOR2_X1 u5_mult_87_U564 ( .A1(u5_mult_87_n384), .A2(u5_mult_87_n317), .ZN(
        u5_mult_87_ab_8__32_) );
  NOR2_X1 u5_mult_87_U563 ( .A1(u5_mult_87_n382), .A2(u5_mult_87_n317), .ZN(
        u5_mult_87_ab_8__33_) );
  NOR2_X1 u5_mult_87_U562 ( .A1(u5_mult_87_n380), .A2(u5_mult_87_n317), .ZN(
        u5_mult_87_ab_8__34_) );
  NOR2_X1 u5_mult_87_U561 ( .A1(u5_mult_87_n378), .A2(u5_mult_87_n317), .ZN(
        u5_mult_87_ab_8__35_) );
  NOR2_X1 u5_mult_87_U560 ( .A1(u5_mult_87_n375), .A2(u5_mult_87_n317), .ZN(
        u5_mult_87_ab_8__36_) );
  NOR2_X1 u5_mult_87_U559 ( .A1(u5_mult_87_n374), .A2(u5_mult_87_n317), .ZN(
        u5_mult_87_ab_8__37_) );
  NOR2_X1 u5_mult_87_U558 ( .A1(u5_mult_87_n371), .A2(u5_mult_87_n317), .ZN(
        u5_mult_87_ab_8__38_) );
  NOR2_X1 u5_mult_87_U557 ( .A1(u5_mult_87_n370), .A2(u5_mult_87_n317), .ZN(
        u5_mult_87_ab_8__39_) );
  NOR2_X1 u5_mult_87_U556 ( .A1(u5_mult_87_n443), .A2(u5_mult_87_n477), .ZN(
        u5_mult_87_ab_8__3_) );
  NOR2_X1 u5_mult_87_U555 ( .A1(u5_mult_87_n368), .A2(u5_mult_87_n477), .ZN(
        u5_mult_87_ab_8__40_) );
  NOR2_X1 u5_mult_87_U554 ( .A1(u5_mult_87_n366), .A2(u5_mult_87_n477), .ZN(
        u5_mult_87_ab_8__41_) );
  NOR2_X1 u5_mult_87_U553 ( .A1(u5_mult_87_n363), .A2(u5_mult_87_n477), .ZN(
        u5_mult_87_ab_8__42_) );
  NOR2_X1 u5_mult_87_U552 ( .A1(u5_mult_87_n361), .A2(u5_mult_87_n315), .ZN(
        u5_mult_87_ab_8__43_) );
  NOR2_X1 u5_mult_87_U551 ( .A1(u5_mult_87_n359), .A2(u5_mult_87_n477), .ZN(
        u5_mult_87_ab_8__44_) );
  NOR2_X1 u5_mult_87_U550 ( .A1(u5_mult_87_n357), .A2(u5_mult_87_n477), .ZN(
        u5_mult_87_ab_8__45_) );
  NOR2_X1 u5_mult_87_U549 ( .A1(u5_mult_87_n355), .A2(u5_mult_87_n477), .ZN(
        u5_mult_87_ab_8__46_) );
  NOR2_X1 u5_mult_87_U548 ( .A1(u5_mult_87_n353), .A2(u5_mult_87_n477), .ZN(
        u5_mult_87_ab_8__47_) );
  NOR2_X1 u5_mult_87_U547 ( .A1(u5_mult_87_n350), .A2(u5_mult_87_n317), .ZN(
        u5_mult_87_ab_8__48_) );
  NOR2_X1 u5_mult_87_U546 ( .A1(u5_mult_87_n347), .A2(u5_mult_87_n477), .ZN(
        u5_mult_87_ab_8__49_) );
  NOR2_X1 u5_mult_87_U545 ( .A1(u5_mult_87_n441), .A2(u5_mult_87_n315), .ZN(
        u5_mult_87_ab_8__4_) );
  NOR2_X1 u5_mult_87_U544 ( .A1(u5_mult_87_n479), .A2(u5_mult_87_n317), .ZN(
        u5_mult_87_ab_8__50_) );
  NOR2_X1 u5_mult_87_U543 ( .A1(u5_mult_87_n345), .A2(u5_mult_87_n316), .ZN(
        u5_mult_87_ab_8__51_) );
  NOR2_X1 u5_mult_87_U542 ( .A1(u5_mult_87_n343), .A2(u5_mult_87_n315), .ZN(
        u5_mult_87_ab_8__52_) );
  NOR2_X1 u5_mult_87_U541 ( .A1(u5_mult_87_n438), .A2(u5_mult_87_n315), .ZN(
        u5_mult_87_ab_8__5_) );
  NOR2_X1 u5_mult_87_U540 ( .A1(u5_mult_87_n435), .A2(u5_mult_87_n315), .ZN(
        u5_mult_87_ab_8__6_) );
  NOR2_X1 u5_mult_87_U539 ( .A1(u5_mult_87_n433), .A2(u5_mult_87_n315), .ZN(
        u5_mult_87_ab_8__7_) );
  NOR2_X1 u5_mult_87_U538 ( .A1(u5_mult_87_n431), .A2(u5_mult_87_n315), .ZN(
        u5_mult_87_ab_8__8_) );
  NOR2_X1 u5_mult_87_U537 ( .A1(u5_mult_87_n429), .A2(u5_mult_87_n315), .ZN(
        u5_mult_87_ab_8__9_) );
  NOR2_X1 u5_mult_87_U536 ( .A1(u5_mult_87_n312), .A2(u5_mult_87_n450), .ZN(
        u5_mult_87_ab_9__0_) );
  NOR2_X1 u5_mult_87_U535 ( .A1(u5_mult_87_n312), .A2(u5_mult_87_n428), .ZN(
        u5_mult_87_ab_9__10_) );
  NOR2_X1 u5_mult_87_U534 ( .A1(u5_mult_87_n312), .A2(u5_mult_87_n426), .ZN(
        u5_mult_87_ab_9__11_) );
  NOR2_X1 u5_mult_87_U533 ( .A1(u5_mult_87_n312), .A2(u5_mult_87_n481), .ZN(
        u5_mult_87_ab_9__12_) );
  NOR2_X1 u5_mult_87_U532 ( .A1(u5_mult_87_n312), .A2(u5_mult_87_n423), .ZN(
        u5_mult_87_ab_9__13_) );
  NOR2_X1 u5_mult_87_U531 ( .A1(u5_mult_87_n312), .A2(u5_mult_87_n420), .ZN(
        u5_mult_87_ab_9__14_) );
  NOR2_X1 u5_mult_87_U530 ( .A1(u5_mult_87_n312), .A2(u5_mult_87_n417), .ZN(
        u5_mult_87_ab_9__15_) );
  NOR2_X1 u5_mult_87_U529 ( .A1(u5_mult_87_n312), .A2(u5_mult_87_n480), .ZN(
        u5_mult_87_ab_9__16_) );
  NOR2_X1 u5_mult_87_U528 ( .A1(u5_mult_87_n312), .A2(u5_mult_87_n414), .ZN(
        u5_mult_87_ab_9__17_) );
  NOR2_X1 u5_mult_87_U527 ( .A1(u5_mult_87_n312), .A2(u5_mult_87_n412), .ZN(
        u5_mult_87_ab_9__18_) );
  NOR2_X1 u5_mult_87_U526 ( .A1(u5_mult_87_n312), .A2(u5_mult_87_n410), .ZN(
        u5_mult_87_ab_9__19_) );
  NOR2_X1 u5_mult_87_U525 ( .A1(u5_mult_87_n313), .A2(u5_mult_87_n448), .ZN(
        u5_mult_87_ab_9__1_) );
  NOR2_X1 u5_mult_87_U524 ( .A1(u5_mult_87_n313), .A2(u5_mult_87_n408), .ZN(
        u5_mult_87_ab_9__20_) );
  NOR2_X1 u5_mult_87_U523 ( .A1(u5_mult_87_n313), .A2(u5_mult_87_n405), .ZN(
        u5_mult_87_ab_9__21_) );
  NOR2_X1 u5_mult_87_U522 ( .A1(u5_mult_87_n313), .A2(u5_mult_87_n404), .ZN(
        u5_mult_87_ab_9__22_) );
  NOR2_X1 u5_mult_87_U521 ( .A1(u5_mult_87_n313), .A2(u5_mult_87_n401), .ZN(
        u5_mult_87_ab_9__23_) );
  NOR2_X1 u5_mult_87_U520 ( .A1(u5_mult_87_n313), .A2(u5_mult_87_n400), .ZN(
        u5_mult_87_ab_9__24_) );
  NOR2_X1 u5_mult_87_U519 ( .A1(u5_mult_87_n313), .A2(u5_mult_87_n397), .ZN(
        u5_mult_87_ab_9__25_) );
  NOR2_X1 u5_mult_87_U518 ( .A1(u5_mult_87_n313), .A2(u5_mult_87_n396), .ZN(
        u5_mult_87_ab_9__26_) );
  NOR2_X1 u5_mult_87_U517 ( .A1(u5_mult_87_n313), .A2(u5_mult_87_n393), .ZN(
        u5_mult_87_ab_9__27_) );
  NOR2_X1 u5_mult_87_U516 ( .A1(u5_mult_87_n313), .A2(u5_mult_87_n392), .ZN(
        u5_mult_87_ab_9__28_) );
  NOR2_X1 u5_mult_87_U515 ( .A1(u5_mult_87_n313), .A2(u5_mult_87_n389), .ZN(
        u5_mult_87_ab_9__29_) );
  NOR2_X1 u5_mult_87_U514 ( .A1(u5_mult_87_n314), .A2(u5_mult_87_n445), .ZN(
        u5_mult_87_ab_9__2_) );
  NOR2_X1 u5_mult_87_U513 ( .A1(u5_mult_87_n314), .A2(u5_mult_87_n388), .ZN(
        u5_mult_87_ab_9__30_) );
  NOR2_X1 u5_mult_87_U512 ( .A1(u5_mult_87_n314), .A2(u5_mult_87_n386), .ZN(
        u5_mult_87_ab_9__31_) );
  NOR2_X1 u5_mult_87_U511 ( .A1(u5_mult_87_n314), .A2(u5_mult_87_n384), .ZN(
        u5_mult_87_ab_9__32_) );
  NOR2_X1 u5_mult_87_U510 ( .A1(u5_mult_87_n314), .A2(u5_mult_87_n382), .ZN(
        u5_mult_87_ab_9__33_) );
  NOR2_X1 u5_mult_87_U509 ( .A1(u5_mult_87_n314), .A2(u5_mult_87_n380), .ZN(
        u5_mult_87_ab_9__34_) );
  NOR2_X1 u5_mult_87_U508 ( .A1(u5_mult_87_n314), .A2(u5_mult_87_n378), .ZN(
        u5_mult_87_ab_9__35_) );
  NOR2_X1 u5_mult_87_U507 ( .A1(u5_mult_87_n314), .A2(u5_mult_87_n376), .ZN(
        u5_mult_87_ab_9__36_) );
  NOR2_X1 u5_mult_87_U506 ( .A1(u5_mult_87_n314), .A2(u5_mult_87_n374), .ZN(
        u5_mult_87_ab_9__37_) );
  NOR2_X1 u5_mult_87_U505 ( .A1(u5_mult_87_n314), .A2(u5_mult_87_n371), .ZN(
        u5_mult_87_ab_9__38_) );
  NOR2_X1 u5_mult_87_U504 ( .A1(u5_mult_87_n314), .A2(u5_mult_87_n370), .ZN(
        u5_mult_87_ab_9__39_) );
  NOR2_X1 u5_mult_87_U503 ( .A1(u5_mult_87_n312), .A2(u5_mult_87_n443), .ZN(
        u5_mult_87_ab_9__3_) );
  NOR2_X1 u5_mult_87_U502 ( .A1(u5_mult_87_n313), .A2(u5_mult_87_n368), .ZN(
        u5_mult_87_ab_9__40_) );
  NOR2_X1 u5_mult_87_U501 ( .A1(u5_mult_87_n313), .A2(u5_mult_87_n366), .ZN(
        u5_mult_87_ab_9__41_) );
  NOR2_X1 u5_mult_87_U500 ( .A1(u5_mult_87_n476), .A2(u5_mult_87_n363), .ZN(
        u5_mult_87_ab_9__42_) );
  NOR2_X1 u5_mult_87_U499 ( .A1(u5_mult_87_n476), .A2(u5_mult_87_n361), .ZN(
        u5_mult_87_ab_9__43_) );
  NOR2_X1 u5_mult_87_U498 ( .A1(u5_mult_87_n476), .A2(u5_mult_87_n359), .ZN(
        u5_mult_87_ab_9__44_) );
  NOR2_X1 u5_mult_87_U497 ( .A1(u5_mult_87_n476), .A2(u5_mult_87_n357), .ZN(
        u5_mult_87_ab_9__45_) );
  NOR2_X1 u5_mult_87_U496 ( .A1(u5_mult_87_n476), .A2(u5_mult_87_n355), .ZN(
        u5_mult_87_ab_9__46_) );
  NOR2_X1 u5_mult_87_U495 ( .A1(u5_mult_87_n476), .A2(u5_mult_87_n353), .ZN(
        u5_mult_87_ab_9__47_) );
  NOR2_X1 u5_mult_87_U494 ( .A1(u5_mult_87_n476), .A2(u5_mult_87_n349), .ZN(
        u5_mult_87_ab_9__48_) );
  NOR2_X1 u5_mult_87_U493 ( .A1(u5_mult_87_n476), .A2(u5_mult_87_n348), .ZN(
        u5_mult_87_ab_9__49_) );
  NOR2_X1 u5_mult_87_U492 ( .A1(u5_mult_87_n312), .A2(u5_mult_87_n441), .ZN(
        u5_mult_87_ab_9__4_) );
  NOR2_X1 u5_mult_87_U491 ( .A1(u5_mult_87_n314), .A2(u5_mult_87_n346), .ZN(
        u5_mult_87_ab_9__50_) );
  NOR2_X1 u5_mult_87_U490 ( .A1(u5_mult_87_n313), .A2(u5_mult_87_n344), .ZN(
        u5_mult_87_ab_9__51_) );
  NOR2_X1 u5_mult_87_U489 ( .A1(u5_mult_87_n312), .A2(u5_mult_87_n343), .ZN(
        u5_mult_87_ab_9__52_) );
  NOR2_X1 u5_mult_87_U488 ( .A1(u5_mult_87_n312), .A2(u5_mult_87_n438), .ZN(
        u5_mult_87_ab_9__5_) );
  NOR2_X1 u5_mult_87_U487 ( .A1(u5_mult_87_n312), .A2(u5_mult_87_n435), .ZN(
        u5_mult_87_ab_9__6_) );
  NOR2_X1 u5_mult_87_U486 ( .A1(u5_mult_87_n312), .A2(u5_mult_87_n433), .ZN(
        u5_mult_87_ab_9__7_) );
  NOR2_X1 u5_mult_87_U485 ( .A1(u5_mult_87_n312), .A2(u5_mult_87_n431), .ZN(
        u5_mult_87_ab_9__8_) );
  NOR2_X1 u5_mult_87_U484 ( .A1(u5_mult_87_n312), .A2(u5_mult_87_n430), .ZN(
        u5_mult_87_ab_9__9_) );
  INV_X4 u5_mult_87_U482 ( .A(u6_N1), .ZN(u5_mult_87_n482) );
  INV_X4 u5_mult_87_U481 ( .A(u6_N12), .ZN(u5_mult_87_n481) );
  INV_X4 u5_mult_87_U480 ( .A(u6_N16), .ZN(u5_mult_87_n480) );
  INV_X4 u5_mult_87_U479 ( .A(u6_N50), .ZN(u5_mult_87_n479) );
  INV_X4 u5_mult_87_U478 ( .A(fracta_mul[3]), .ZN(u5_mult_87_n478) );
  INV_X4 u5_mult_87_U477 ( .A(fracta_mul[8]), .ZN(u5_mult_87_n477) );
  INV_X4 u5_mult_87_U476 ( .A(fracta_mul[9]), .ZN(u5_mult_87_n476) );
  INV_X4 u5_mult_87_U475 ( .A(fracta_mul[10]), .ZN(u5_mult_87_n475) );
  INV_X4 u5_mult_87_U474 ( .A(fracta_mul[11]), .ZN(u5_mult_87_n474) );
  INV_X4 u5_mult_87_U473 ( .A(fracta_mul[12]), .ZN(u5_mult_87_n473) );
  INV_X4 u5_mult_87_U472 ( .A(fracta_mul[14]), .ZN(u5_mult_87_n472) );
  INV_X4 u5_mult_87_U471 ( .A(fracta_mul[16]), .ZN(u5_mult_87_n471) );
  INV_X4 u5_mult_87_U470 ( .A(fracta_mul[17]), .ZN(u5_mult_87_n470) );
  INV_X4 u5_mult_87_U469 ( .A(fracta_mul[18]), .ZN(u5_mult_87_n469) );
  INV_X4 u5_mult_87_U468 ( .A(fracta_mul[20]), .ZN(u5_mult_87_n468) );
  INV_X4 u5_mult_87_U467 ( .A(fracta_mul[21]), .ZN(u5_mult_87_n467) );
  INV_X4 u5_mult_87_U466 ( .A(fracta_mul[22]), .ZN(u5_mult_87_n466) );
  INV_X4 u5_mult_87_U465 ( .A(fracta_mul[23]), .ZN(u5_mult_87_n465) );
  INV_X4 u5_mult_87_U464 ( .A(fracta_mul[25]), .ZN(u5_mult_87_n464) );
  INV_X4 u5_mult_87_U463 ( .A(fracta_mul[27]), .ZN(u5_mult_87_n463) );
  INV_X4 u5_mult_87_U462 ( .A(fracta_mul[28]), .ZN(u5_mult_87_n462) );
  INV_X4 u5_mult_87_U461 ( .A(fracta_mul[29]), .ZN(u5_mult_87_n461) );
  INV_X4 u5_mult_87_U460 ( .A(fracta_mul[31]), .ZN(u5_mult_87_n460) );
  INV_X4 u5_mult_87_U459 ( .A(fracta_mul[33]), .ZN(u5_mult_87_n459) );
  INV_X4 u5_mult_87_U458 ( .A(fracta_mul[34]), .ZN(u5_mult_87_n458) );
  INV_X4 u5_mult_87_U457 ( .A(fracta_mul[35]), .ZN(u5_mult_87_n457) );
  INV_X4 u5_mult_87_U456 ( .A(fracta_mul[37]), .ZN(u5_mult_87_n456) );
  INV_X4 u5_mult_87_U455 ( .A(fracta_mul[40]), .ZN(u5_mult_87_n455) );
  INV_X4 u5_mult_87_U454 ( .A(fracta_mul[46]), .ZN(u5_mult_87_n454) );
  XOR2_X2 u5_mult_87_U453 ( .A(u5_mult_87_ab_1__0_), .B(u5_mult_87_ab_0__1_), 
        .Z(u5_N1) );
  INV_X4 u5_mult_87_U452 ( .A(fracta_mul[50]), .ZN(u5_mult_87_n214) );
  INV_X4 u5_mult_87_U451 ( .A(fracta_mul[50]), .ZN(u5_mult_87_n215) );
  INV_X4 u5_mult_87_U450 ( .A(fracta_mul[47]), .ZN(u5_mult_87_n222) );
  INV_X4 u5_mult_87_U449 ( .A(fracta_mul[47]), .ZN(u5_mult_87_n224) );
  INV_X4 u5_mult_87_U448 ( .A(fracta_mul[48]), .ZN(u5_mult_87_n220) );
  INV_X4 u5_mult_87_U447 ( .A(fracta_mul[48]), .ZN(u5_mult_87_n221) );
  INV_X4 u5_mult_87_U446 ( .A(fracta_mul[49]), .ZN(u5_mult_87_n217) );
  INV_X4 u5_mult_87_U445 ( .A(fracta_mul[49]), .ZN(u5_mult_87_n218) );
  INV_X4 u5_mult_87_U444 ( .A(fracta_mul[51]), .ZN(u5_mult_87_n211) );
  INV_X4 u5_mult_87_U443 ( .A(fracta_mul[51]), .ZN(u5_mult_87_n210) );
  INV_X4 u5_mult_87_U442 ( .A(fracta_mul[51]), .ZN(u5_mult_87_n212) );
  INV_X4 u5_mult_87_U441 ( .A(n4825), .ZN(u5_mult_87_n451) );
  INV_X4 u5_mult_87_U440 ( .A(n4825), .ZN(u5_mult_87_n453) );
  INV_X4 u5_mult_87_U439 ( .A(fracta_mul[46]), .ZN(u5_mult_87_n225) );
  INV_X4 u5_mult_87_U438 ( .A(fracta_mul[42]), .ZN(u5_mult_87_n237) );
  INV_X4 u5_mult_87_U437 ( .A(fracta_mul[42]), .ZN(u5_mult_87_n236) );
  INV_X4 u5_mult_87_U436 ( .A(fracta_mul[42]), .ZN(u5_mult_87_n238) );
  INV_X4 u5_mult_87_U435 ( .A(fracta_mul[45]), .ZN(u5_mult_87_n228) );
  INV_X4 u5_mult_87_U434 ( .A(fracta_mul[45]), .ZN(u5_mult_87_n229) );
  INV_X4 u5_mult_87_U433 ( .A(u5_mult_87_n247), .ZN(u5_mult_87_n246) );
  INV_X4 u5_mult_87_U432 ( .A(u5_mult_87_n247), .ZN(u5_mult_87_n245) );
  INV_X4 u5_mult_87_U431 ( .A(u5_mult_87_n247), .ZN(u5_mult_87_n244) );
  INV_X4 u5_mult_87_U430 ( .A(fracta_mul[43]), .ZN(u5_mult_87_n233) );
  INV_X4 u5_mult_87_U429 ( .A(fracta_mul[43]), .ZN(u5_mult_87_n234) );
  INV_X4 u5_mult_87_U428 ( .A(fracta_mul[43]), .ZN(u5_mult_87_n235) );
  INV_X4 u5_mult_87_U427 ( .A(fracta_mul[36]), .ZN(u5_mult_87_n257) );
  INV_X4 u5_mult_87_U426 ( .A(fracta_mul[38]), .ZN(u5_mult_87_n252) );
  INV_X4 u5_mult_87_U425 ( .A(fracta_mul[38]), .ZN(u5_mult_87_n251) );
  INV_X4 u5_mult_87_U424 ( .A(fracta_mul[33]), .ZN(u5_mult_87_n263) );
  INV_X4 u5_mult_87_U423 ( .A(fracta_mul[37]), .ZN(u5_mult_87_n255) );
  INV_X4 u5_mult_87_U422 ( .A(fracta_mul[37]), .ZN(u5_mult_87_n254) );
  INV_X4 u5_mult_87_U421 ( .A(fracta_mul[32]), .ZN(u5_mult_87_n266) );
  INV_X4 u5_mult_87_U420 ( .A(fracta_mul[28]), .ZN(u5_mult_87_n276) );
  INV_X4 u5_mult_87_U419 ( .A(fracta_mul[29]), .ZN(u5_mult_87_n274) );
  INV_X4 u5_mult_87_U418 ( .A(fracta_mul[31]), .ZN(u5_mult_87_n269) );
  INV_X4 u5_mult_87_U417 ( .A(fracta_mul[22]), .ZN(u5_mult_87_n286) );
  INV_X4 u5_mult_87_U416 ( .A(fracta_mul[23]), .ZN(u5_mult_87_n284) );
  INV_X4 u5_mult_87_U415 ( .A(fracta_mul[21]), .ZN(u5_mult_87_n288) );
  INV_X4 u5_mult_87_U414 ( .A(fracta_mul[25]), .ZN(u5_mult_87_n281) );
  INV_X4 u5_mult_87_U413 ( .A(fracta_mul[24]), .ZN(u5_mult_87_n282) );
  INV_X4 u5_mult_87_U412 ( .A(fracta_mul[20]), .ZN(u5_mult_87_n290) );
  INV_X4 u5_mult_87_U411 ( .A(fracta_mul[19]), .ZN(u5_mult_87_n293) );
  INV_X4 u5_mult_87_U410 ( .A(fracta_mul[16]), .ZN(u5_mult_87_n299) );
  INV_X4 u5_mult_87_U409 ( .A(fracta_mul[17]), .ZN(u5_mult_87_n297) );
  INV_X4 u5_mult_87_U408 ( .A(fracta_mul[13]), .ZN(u5_mult_87_n304) );
  INV_X4 u5_mult_87_U407 ( .A(fracta_mul[15]), .ZN(u5_mult_87_n301) );
  INV_X4 u5_mult_87_U406 ( .A(fracta_mul[12]), .ZN(u5_mult_87_n307) );
  AND2_X4 u5_mult_87_U405 ( .A1(u5_mult_87_ab_52__52_), .A2(
        u5_mult_87_CARRYB_52__51_), .ZN(u5_mult_87_n208) );
  INV_X4 u5_mult_87_U404 ( .A(fracta_mul[11]), .ZN(u5_mult_87_n308) );
  INV_X4 u5_mult_87_U403 ( .A(fracta_mul[11]), .ZN(u5_mult_87_n309) );
  INV_X4 u5_mult_87_U402 ( .A(fracta_mul[10]), .ZN(u5_mult_87_n310) );
  INV_X4 u5_mult_87_U401 ( .A(fracta_mul[10]), .ZN(u5_mult_87_n311) );
  INV_X4 u5_mult_87_U400 ( .A(u5_mult_87_n318), .ZN(u5_mult_87_n315) );
  INV_X4 u5_mult_87_U399 ( .A(u5_mult_87_n318), .ZN(u5_mult_87_n316) );
  INV_X4 u5_mult_87_U398 ( .A(u5_mult_87_n318), .ZN(u5_mult_87_n317) );
  INV_X4 u5_mult_87_U397 ( .A(u6_N18), .ZN(u5_mult_87_n412) );
  INV_X4 u5_mult_87_U396 ( .A(u6_N1), .ZN(u5_mult_87_n448) );
  INV_X4 u5_mult_87_U395 ( .A(u6_N2), .ZN(u5_mult_87_n445) );
  INV_X4 u5_mult_87_U394 ( .A(fracta_mul[9]), .ZN(u5_mult_87_n312) );
  INV_X4 u5_mult_87_U393 ( .A(fracta_mul[9]), .ZN(u5_mult_87_n313) );
  INV_X4 u5_mult_87_U392 ( .A(fracta_mul[9]), .ZN(u5_mult_87_n314) );
  INV_X4 u5_mult_87_U391 ( .A(u6_N0), .ZN(u5_mult_87_n450) );
  XOR2_X2 u5_mult_87_U390 ( .A(u5_mult_87_CARRYB_52__0_), .B(
        u5_mult_87_SUMB_52__1_), .Z(u5_N53) );
  AND2_X4 u5_mult_87_U389 ( .A1(u5_mult_87_SUMB_52__48_), .A2(
        u5_mult_87_CARRYB_52__47_), .ZN(u5_mult_87_n206) );
  AND2_X4 u5_mult_87_U388 ( .A1(u5_mult_87_SUMB_52__47_), .A2(
        u5_mult_87_CARRYB_52__46_), .ZN(u5_mult_87_n205) );
  AND2_X4 u5_mult_87_U387 ( .A1(u5_mult_87_SUMB_52__46_), .A2(
        u5_mult_87_CARRYB_52__45_), .ZN(u5_mult_87_n204) );
  AND2_X4 u5_mult_87_U386 ( .A1(u5_mult_87_SUMB_52__36_), .A2(
        u5_mult_87_CARRYB_52__35_), .ZN(u5_mult_87_n203) );
  AND2_X4 u5_mult_87_U385 ( .A1(u5_mult_87_SUMB_52__37_), .A2(
        u5_mult_87_CARRYB_52__36_), .ZN(u5_mult_87_n202) );
  AND2_X4 u5_mult_87_U384 ( .A1(u5_mult_87_SUMB_52__40_), .A2(
        u5_mult_87_CARRYB_52__39_), .ZN(u5_mult_87_n201) );
  AND2_X4 u5_mult_87_U383 ( .A1(u5_mult_87_SUMB_52__39_), .A2(
        u5_mult_87_CARRYB_52__38_), .ZN(u5_mult_87_n200) );
  AND2_X4 u5_mult_87_U382 ( .A1(u5_mult_87_SUMB_52__38_), .A2(
        u5_mult_87_CARRYB_52__37_), .ZN(u5_mult_87_n199) );
  AND2_X4 u5_mult_87_U381 ( .A1(u5_mult_87_SUMB_52__41_), .A2(
        u5_mult_87_CARRYB_52__40_), .ZN(u5_mult_87_n198) );
  AND2_X4 u5_mult_87_U380 ( .A1(u5_mult_87_SUMB_52__44_), .A2(
        u5_mult_87_CARRYB_52__43_), .ZN(u5_mult_87_n197) );
  AND2_X4 u5_mult_87_U379 ( .A1(u5_mult_87_SUMB_52__42_), .A2(
        u5_mult_87_CARRYB_52__41_), .ZN(u5_mult_87_n196) );
  AND2_X4 u5_mult_87_U378 ( .A1(u5_mult_87_SUMB_52__32_), .A2(
        u5_mult_87_CARRYB_52__31_), .ZN(u5_mult_87_n195) );
  AND2_X4 u5_mult_87_U377 ( .A1(u5_mult_87_SUMB_52__50_), .A2(
        u5_mult_87_CARRYB_52__49_), .ZN(u5_mult_87_n194) );
  AND2_X4 u5_mult_87_U376 ( .A1(u5_mult_87_SUMB_52__35_), .A2(
        u5_mult_87_CARRYB_52__34_), .ZN(u5_mult_87_n193) );
  AND2_X4 u5_mult_87_U375 ( .A1(u5_mult_87_SUMB_52__43_), .A2(
        u5_mult_87_CARRYB_52__42_), .ZN(u5_mult_87_n192) );
  AND2_X4 u5_mult_87_U374 ( .A1(u5_mult_87_SUMB_52__49_), .A2(
        u5_mult_87_CARRYB_52__48_), .ZN(u5_mult_87_n191) );
  AND2_X4 u5_mult_87_U373 ( .A1(u5_mult_87_SUMB_52__51_), .A2(
        u5_mult_87_CARRYB_52__50_), .ZN(u5_mult_87_n190) );
  AND2_X4 u5_mult_87_U372 ( .A1(u5_mult_87_SUMB_52__45_), .A2(
        u5_mult_87_CARRYB_52__44_), .ZN(u5_mult_87_n189) );
  INV_X4 u5_mult_87_U371 ( .A(fracta_mul[7]), .ZN(u5_mult_87_n320) );
  XOR2_X2 u5_mult_87_U370 ( .A(u5_mult_87_ab_1__1_), .B(u5_mult_87_ab_0__2_), 
        .Z(u5_mult_87_n188) );
  INV_X4 u5_mult_87_U369 ( .A(fracta_mul[0]), .ZN(u5_mult_87_n340) );
  INV_X4 u5_mult_87_U368 ( .A(fracta_mul[0]), .ZN(u5_mult_87_n341) );
  INV_X4 u5_mult_87_U367 ( .A(fracta_mul[3]), .ZN(u5_mult_87_n330) );
  INV_X4 u5_mult_87_U366 ( .A(fracta_mul[3]), .ZN(u5_mult_87_n331) );
  INV_X4 u5_mult_87_U365 ( .A(fracta_mul[4]), .ZN(u5_mult_87_n327) );
  INV_X4 u5_mult_87_U364 ( .A(fracta_mul[4]), .ZN(u5_mult_87_n328) );
  INV_X4 u5_mult_87_U363 ( .A(fracta_mul[5]), .ZN(u5_mult_87_n323) );
  INV_X4 u5_mult_87_U362 ( .A(fracta_mul[5]), .ZN(u5_mult_87_n324) );
  INV_X4 u5_mult_87_U361 ( .A(fracta_mul[5]), .ZN(u5_mult_87_n325) );
  INV_X4 u5_mult_87_U360 ( .A(fracta_mul[2]), .ZN(u5_mult_87_n333) );
  INV_X4 u5_mult_87_U359 ( .A(fracta_mul[2]), .ZN(u5_mult_87_n334) );
  INV_X4 u5_mult_87_U358 ( .A(fracta_mul[2]), .ZN(u5_mult_87_n335) );
  INV_X4 u5_mult_87_U357 ( .A(fracta_mul[1]), .ZN(u5_mult_87_n337) );
  INV_X4 u5_mult_87_U356 ( .A(fracta_mul[1]), .ZN(u5_mult_87_n338) );
  INV_X4 u5_mult_87_U355 ( .A(u6_N19), .ZN(u5_mult_87_n410) );
  INV_X4 u5_mult_87_U354 ( .A(u6_N20), .ZN(u5_mult_87_n408) );
  INV_X4 u5_mult_87_U353 ( .A(u6_N24), .ZN(u5_mult_87_n400) );
  INV_X4 u5_mult_87_U352 ( .A(u6_N26), .ZN(u5_mult_87_n396) );
  INV_X4 u5_mult_87_U351 ( .A(u6_N30), .ZN(u5_mult_87_n388) );
  INV_X4 u5_mult_87_U350 ( .A(u6_N34), .ZN(u5_mult_87_n380) );
  INV_X4 u5_mult_87_U349 ( .A(u6_N41), .ZN(u5_mult_87_n366) );
  INV_X4 u5_mult_87_U348 ( .A(u6_N43), .ZN(u5_mult_87_n361) );
  INV_X4 u5_mult_87_U347 ( .A(u6_N44), .ZN(u5_mult_87_n359) );
  INV_X4 u5_mult_87_U346 ( .A(u6_N45), .ZN(u5_mult_87_n357) );
  INV_X4 u5_mult_87_U345 ( .A(u6_N46), .ZN(u5_mult_87_n355) );
  INV_X4 u5_mult_87_U344 ( .A(u6_N35), .ZN(u5_mult_87_n378) );
  INV_X4 u5_mult_87_U343 ( .A(u6_N11), .ZN(u5_mult_87_n426) );
  INV_X4 u5_mult_87_U342 ( .A(u6_N13), .ZN(u5_mult_87_n423) );
  INV_X4 u5_mult_87_U341 ( .A(u6_N14), .ZN(u5_mult_87_n420) );
  INV_X4 u5_mult_87_U340 ( .A(u6_N14), .ZN(u5_mult_87_n421) );
  INV_X4 u5_mult_87_U339 ( .A(u6_N15), .ZN(u5_mult_87_n417) );
  AND2_X4 u5_mult_87_U338 ( .A1(u5_mult_87_SUMB_52__33_), .A2(
        u5_mult_87_CARRYB_52__32_), .ZN(u5_mult_87_n187) );
  AND2_X4 u5_mult_87_U337 ( .A1(u5_mult_87_SUMB_52__34_), .A2(
        u5_mult_87_CARRYB_52__33_), .ZN(u5_mult_87_n186) );
  AND2_X4 u5_mult_87_U336 ( .A1(u5_mult_87_SUMB_52__30_), .A2(
        u5_mult_87_CARRYB_52__29_), .ZN(u5_mult_87_n185) );
  AND2_X4 u5_mult_87_U335 ( .A1(u5_mult_87_SUMB_52__17_), .A2(
        u5_mult_87_CARRYB_52__16_), .ZN(u5_mult_87_n184) );
  AND2_X4 u5_mult_87_U334 ( .A1(u5_mult_87_SUMB_52__20_), .A2(
        u5_mult_87_CARRYB_52__19_), .ZN(u5_mult_87_n183) );
  AND2_X4 u5_mult_87_U333 ( .A1(u5_mult_87_SUMB_52__18_), .A2(
        u5_mult_87_CARRYB_52__17_), .ZN(u5_mult_87_n182) );
  AND2_X4 u5_mult_87_U332 ( .A1(u5_mult_87_SUMB_52__21_), .A2(
        u5_mult_87_CARRYB_52__20_), .ZN(u5_mult_87_n181) );
  AND2_X4 u5_mult_87_U331 ( .A1(u5_mult_87_SUMB_52__24_), .A2(
        u5_mult_87_CARRYB_52__23_), .ZN(u5_mult_87_n180) );
  AND2_X4 u5_mult_87_U330 ( .A1(u5_mult_87_SUMB_52__23_), .A2(
        u5_mult_87_CARRYB_52__22_), .ZN(u5_mult_87_n179) );
  AND2_X4 u5_mult_87_U329 ( .A1(u5_mult_87_SUMB_52__22_), .A2(
        u5_mult_87_CARRYB_52__21_), .ZN(u5_mult_87_n178) );
  AND2_X4 u5_mult_87_U328 ( .A1(u5_mult_87_SUMB_52__25_), .A2(
        u5_mult_87_CARRYB_52__24_), .ZN(u5_mult_87_n177) );
  AND2_X4 u5_mult_87_U327 ( .A1(u5_mult_87_SUMB_52__28_), .A2(
        u5_mult_87_CARRYB_52__27_), .ZN(u5_mult_87_n176) );
  AND2_X4 u5_mult_87_U326 ( .A1(u5_mult_87_SUMB_52__26_), .A2(
        u5_mult_87_CARRYB_52__25_), .ZN(u5_mult_87_n175) );
  AND2_X4 u5_mult_87_U325 ( .A1(u5_mult_87_SUMB_52__14_), .A2(
        u5_mult_87_CARRYB_52__13_), .ZN(u5_mult_87_n174) );
  AND2_X4 u5_mult_87_U324 ( .A1(u5_mult_87_SUMB_52__10_), .A2(
        u5_mult_87_CARRYB_52__9_), .ZN(u5_mult_87_n173) );
  AND2_X4 u5_mult_87_U323 ( .A1(u5_mult_87_SUMB_52__9_), .A2(
        u5_mult_87_CARRYB_52__8_), .ZN(u5_mult_87_n172) );
  AND2_X4 u5_mult_87_U322 ( .A1(u5_mult_87_SUMB_52__12_), .A2(
        u5_mult_87_CARRYB_52__11_), .ZN(u5_mult_87_n171) );
  AND2_X4 u5_mult_87_U321 ( .A1(u5_mult_87_SUMB_52__6_), .A2(
        u5_mult_87_CARRYB_52__5_), .ZN(u5_mult_87_n170) );
  AND2_X4 u5_mult_87_U320 ( .A1(u5_mult_87_SUMB_52__5_), .A2(
        u5_mult_87_CARRYB_52__4_), .ZN(u5_mult_87_n169) );
  AND2_X4 u5_mult_87_U319 ( .A1(u5_mult_87_SUMB_52__8_), .A2(
        u5_mult_87_CARRYB_52__7_), .ZN(u5_mult_87_n168) );
  AND2_X4 u5_mult_87_U318 ( .A1(u5_mult_87_SUMB_52__4_), .A2(
        u5_mult_87_CARRYB_52__3_), .ZN(u5_mult_87_n167) );
  AND2_X4 u5_mult_87_U317 ( .A1(u5_mult_87_SUMB_52__15_), .A2(
        u5_mult_87_CARRYB_52__14_), .ZN(u5_mult_87_n166) );
  AND2_X4 u5_mult_87_U316 ( .A1(u5_mult_87_SUMB_52__16_), .A2(
        u5_mult_87_CARRYB_52__15_), .ZN(u5_mult_87_n165) );
  AND2_X4 u5_mult_87_U315 ( .A1(u5_mult_87_SUMB_52__13_), .A2(
        u5_mult_87_CARRYB_52__12_), .ZN(u5_mult_87_n164) );
  AND2_X4 u5_mult_87_U314 ( .A1(u5_mult_87_SUMB_52__29_), .A2(
        u5_mult_87_CARRYB_52__28_), .ZN(u5_mult_87_n163) );
  AND2_X4 u5_mult_87_U313 ( .A1(u5_mult_87_SUMB_52__19_), .A2(
        u5_mult_87_CARRYB_52__18_), .ZN(u5_mult_87_n162) );
  AND2_X4 u5_mult_87_U312 ( .A1(u5_mult_87_SUMB_52__27_), .A2(
        u5_mult_87_CARRYB_52__26_), .ZN(u5_mult_87_n161) );
  AND2_X4 u5_mult_87_U311 ( .A1(u5_mult_87_SUMB_52__7_), .A2(
        u5_mult_87_CARRYB_52__6_), .ZN(u5_mult_87_n160) );
  AND2_X4 u5_mult_87_U310 ( .A1(u5_mult_87_SUMB_52__31_), .A2(
        u5_mult_87_CARRYB_52__30_), .ZN(u5_mult_87_n159) );
  AND2_X4 u5_mult_87_U309 ( .A1(u5_mult_87_SUMB_52__11_), .A2(
        u5_mult_87_CARRYB_52__10_), .ZN(u5_mult_87_n158) );
  INV_X4 u5_mult_87_U308 ( .A(u6_N5), .ZN(u5_mult_87_n439) );
  INV_X4 u5_mult_87_U307 ( .A(u6_N6), .ZN(u5_mult_87_n436) );
  INV_X4 u5_mult_87_U306 ( .A(u6_N7), .ZN(u5_mult_87_n434) );
  INV_X4 u5_mult_87_U305 ( .A(u6_N8), .ZN(u5_mult_87_n432) );
  XOR2_X2 u5_mult_87_U304 ( .A(u5_mult_87_ab_1__2_), .B(u5_mult_87_ab_0__3_), 
        .Z(u5_mult_87_n157) );
  XOR2_X2 u5_mult_87_U303 ( .A(u5_mult_87_ab_1__3_), .B(u5_mult_87_ab_0__4_), 
        .Z(u5_mult_87_n156) );
  XOR2_X2 u5_mult_87_U302 ( .A(u5_mult_87_ab_1__4_), .B(u5_mult_87_ab_0__5_), 
        .Z(u5_mult_87_n155) );
  XOR2_X2 u5_mult_87_U301 ( .A(u5_mult_87_ab_1__5_), .B(u5_mult_87_ab_0__6_), 
        .Z(u5_mult_87_n154) );
  XOR2_X2 u5_mult_87_U300 ( .A(u5_mult_87_ab_1__6_), .B(u5_mult_87_ab_0__7_), 
        .Z(u5_mult_87_n153) );
  XOR2_X2 u5_mult_87_U299 ( .A(u5_mult_87_ab_1__7_), .B(u5_mult_87_ab_0__8_), 
        .Z(u5_mult_87_n152) );
  XOR2_X2 u5_mult_87_U298 ( .A(u5_mult_87_ab_1__8_), .B(u5_mult_87_ab_0__9_), 
        .Z(u5_mult_87_n151) );
  XOR2_X2 u5_mult_87_U297 ( .A(u5_mult_87_ab_1__9_), .B(u5_mult_87_ab_0__10_), 
        .Z(u5_mult_87_n150) );
  XOR2_X2 u5_mult_87_U296 ( .A(u5_mult_87_ab_1__10_), .B(u5_mult_87_ab_0__11_), 
        .Z(u5_mult_87_n149) );
  XOR2_X2 u5_mult_87_U295 ( .A(u5_mult_87_ab_1__11_), .B(u5_mult_87_ab_0__12_), 
        .Z(u5_mult_87_n148) );
  XOR2_X2 u5_mult_87_U294 ( .A(u5_mult_87_ab_1__12_), .B(u5_mult_87_ab_0__13_), 
        .Z(u5_mult_87_n147) );
  XOR2_X2 u5_mult_87_U293 ( .A(u5_mult_87_ab_1__13_), .B(u5_mult_87_ab_0__14_), 
        .Z(u5_mult_87_n146) );
  XOR2_X2 u5_mult_87_U292 ( .A(u5_mult_87_ab_1__14_), .B(u5_mult_87_ab_0__15_), 
        .Z(u5_mult_87_n145) );
  XOR2_X2 u5_mult_87_U291 ( .A(u5_mult_87_ab_1__15_), .B(u5_mult_87_ab_0__16_), 
        .Z(u5_mult_87_n144) );
  XOR2_X2 u5_mult_87_U290 ( .A(u5_mult_87_ab_1__16_), .B(u5_mult_87_ab_0__17_), 
        .Z(u5_mult_87_n143) );
  XOR2_X2 u5_mult_87_U289 ( .A(u5_mult_87_ab_1__17_), .B(u5_mult_87_ab_0__18_), 
        .Z(u5_mult_87_n142) );
  XOR2_X2 u5_mult_87_U288 ( .A(u5_mult_87_ab_1__18_), .B(u5_mult_87_ab_0__19_), 
        .Z(u5_mult_87_n141) );
  XOR2_X2 u5_mult_87_U287 ( .A(u5_mult_87_ab_1__19_), .B(u5_mult_87_ab_0__20_), 
        .Z(u5_mult_87_n140) );
  XOR2_X2 u5_mult_87_U286 ( .A(u5_mult_87_ab_1__20_), .B(u5_mult_87_ab_0__21_), 
        .Z(u5_mult_87_n139) );
  XOR2_X2 u5_mult_87_U285 ( .A(u5_mult_87_ab_1__21_), .B(u5_mult_87_ab_0__22_), 
        .Z(u5_mult_87_n138) );
  XOR2_X2 u5_mult_87_U284 ( .A(u5_mult_87_ab_1__22_), .B(u5_mult_87_ab_0__23_), 
        .Z(u5_mult_87_n137) );
  XOR2_X2 u5_mult_87_U283 ( .A(u5_mult_87_ab_1__23_), .B(u5_mult_87_ab_0__24_), 
        .Z(u5_mult_87_n136) );
  XOR2_X2 u5_mult_87_U282 ( .A(u5_mult_87_ab_1__24_), .B(u5_mult_87_ab_0__25_), 
        .Z(u5_mult_87_n135) );
  XOR2_X2 u5_mult_87_U281 ( .A(u5_mult_87_ab_1__25_), .B(u5_mult_87_ab_0__26_), 
        .Z(u5_mult_87_n134) );
  XOR2_X2 u5_mult_87_U280 ( .A(u5_mult_87_ab_1__26_), .B(u5_mult_87_ab_0__27_), 
        .Z(u5_mult_87_n133) );
  XOR2_X2 u5_mult_87_U279 ( .A(u5_mult_87_ab_1__27_), .B(u5_mult_87_ab_0__28_), 
        .Z(u5_mult_87_n132) );
  XOR2_X2 u5_mult_87_U278 ( .A(u5_mult_87_ab_1__28_), .B(u5_mult_87_ab_0__29_), 
        .Z(u5_mult_87_n131) );
  XOR2_X2 u5_mult_87_U277 ( .A(u5_mult_87_ab_1__29_), .B(u5_mult_87_ab_0__30_), 
        .Z(u5_mult_87_n130) );
  XOR2_X2 u5_mult_87_U276 ( .A(u5_mult_87_ab_1__30_), .B(u5_mult_87_ab_0__31_), 
        .Z(u5_mult_87_n129) );
  XOR2_X2 u5_mult_87_U275 ( .A(u5_mult_87_ab_1__31_), .B(u5_mult_87_ab_0__32_), 
        .Z(u5_mult_87_n128) );
  XOR2_X2 u5_mult_87_U274 ( .A(u5_mult_87_ab_1__32_), .B(u5_mult_87_ab_0__33_), 
        .Z(u5_mult_87_n127) );
  XOR2_X2 u5_mult_87_U273 ( .A(u5_mult_87_ab_1__33_), .B(u5_mult_87_ab_0__34_), 
        .Z(u5_mult_87_n126) );
  XOR2_X2 u5_mult_87_U272 ( .A(u5_mult_87_ab_1__34_), .B(u5_mult_87_ab_0__35_), 
        .Z(u5_mult_87_n125) );
  XOR2_X2 u5_mult_87_U271 ( .A(u5_mult_87_ab_1__35_), .B(u5_mult_87_ab_0__36_), 
        .Z(u5_mult_87_n124) );
  XOR2_X2 u5_mult_87_U270 ( .A(u5_mult_87_ab_1__36_), .B(u5_mult_87_ab_0__37_), 
        .Z(u5_mult_87_n123) );
  XOR2_X2 u5_mult_87_U269 ( .A(u5_mult_87_ab_1__37_), .B(u5_mult_87_ab_0__38_), 
        .Z(u5_mult_87_n122) );
  XOR2_X2 u5_mult_87_U268 ( .A(u5_mult_87_ab_1__38_), .B(u5_mult_87_ab_0__39_), 
        .Z(u5_mult_87_n121) );
  XOR2_X2 u5_mult_87_U267 ( .A(u5_mult_87_ab_1__39_), .B(u5_mult_87_ab_0__40_), 
        .Z(u5_mult_87_n120) );
  XOR2_X2 u5_mult_87_U266 ( .A(u5_mult_87_ab_1__40_), .B(u5_mult_87_ab_0__41_), 
        .Z(u5_mult_87_n119) );
  XOR2_X2 u5_mult_87_U265 ( .A(u5_mult_87_ab_1__41_), .B(u5_mult_87_ab_0__42_), 
        .Z(u5_mult_87_n118) );
  XOR2_X2 u5_mult_87_U264 ( .A(u5_mult_87_ab_1__42_), .B(u5_mult_87_ab_0__43_), 
        .Z(u5_mult_87_n117) );
  XOR2_X2 u5_mult_87_U263 ( .A(u5_mult_87_ab_1__43_), .B(u5_mult_87_ab_0__44_), 
        .Z(u5_mult_87_n116) );
  XOR2_X2 u5_mult_87_U262 ( .A(u5_mult_87_ab_1__44_), .B(u5_mult_87_ab_0__45_), 
        .Z(u5_mult_87_n115) );
  XOR2_X2 u5_mult_87_U261 ( .A(u5_mult_87_ab_1__45_), .B(u5_mult_87_ab_0__46_), 
        .Z(u5_mult_87_n114) );
  XOR2_X2 u5_mult_87_U260 ( .A(u5_mult_87_ab_1__46_), .B(u5_mult_87_ab_0__47_), 
        .Z(u5_mult_87_n113) );
  XOR2_X2 u5_mult_87_U259 ( .A(u5_mult_87_ab_1__47_), .B(u5_mult_87_ab_0__48_), 
        .Z(u5_mult_87_n112) );
  XOR2_X2 u5_mult_87_U258 ( .A(u5_mult_87_ab_1__48_), .B(u5_mult_87_ab_0__49_), 
        .Z(u5_mult_87_n111) );
  XOR2_X2 u5_mult_87_U257 ( .A(u5_mult_87_ab_1__49_), .B(u5_mult_87_ab_0__50_), 
        .Z(u5_mult_87_n110) );
  XOR2_X2 u5_mult_87_U256 ( .A(u5_mult_87_ab_1__50_), .B(u5_mult_87_ab_0__51_), 
        .Z(u5_mult_87_n109) );
  AND2_X4 u5_mult_87_U255 ( .A1(u5_mult_87_ab_0__51_), .A2(
        u5_mult_87_ab_1__50_), .ZN(u5_mult_87_n108) );
  AND2_X4 u5_mult_87_U254 ( .A1(u5_mult_87_SUMB_52__3_), .A2(
        u5_mult_87_CARRYB_52__2_), .ZN(u5_mult_87_n107) );
  AND2_X4 u5_mult_87_U253 ( .A1(u5_mult_87_SUMB_52__2_), .A2(
        u5_mult_87_CARRYB_52__1_), .ZN(u5_mult_87_n106) );
  AND2_X4 u5_mult_87_U252 ( .A1(u5_mult_87_SUMB_52__1_), .A2(
        u5_mult_87_CARRYB_52__0_), .ZN(u5_mult_87_n105) );
  AND2_X4 u5_mult_87_U251 ( .A1(u5_mult_87_ab_0__52_), .A2(
        u5_mult_87_ab_1__51_), .ZN(u5_mult_87_n104) );
  INV_X4 u5_mult_87_U250 ( .A(n4825), .ZN(u5_mult_87_n452) );
  INV_X4 u5_mult_87_U249 ( .A(fracta_mul[46]), .ZN(u5_mult_87_n226) );
  INV_X4 u5_mult_87_U248 ( .A(fracta_mul[42]), .ZN(u5_mult_87_n239) );
  INV_X4 u5_mult_87_U247 ( .A(fracta_mul[44]), .ZN(u5_mult_87_n230) );
  INV_X4 u5_mult_87_U246 ( .A(fracta_mul[44]), .ZN(u5_mult_87_n231) );
  INV_X4 u5_mult_87_U245 ( .A(fracta_mul[44]), .ZN(u5_mult_87_n232) );
  INV_X4 u5_mult_87_U244 ( .A(fracta_mul[41]), .ZN(u5_mult_87_n241) );
  INV_X4 u5_mult_87_U243 ( .A(fracta_mul[41]), .ZN(u5_mult_87_n242) );
  INV_X4 u5_mult_87_U242 ( .A(fracta_mul[41]), .ZN(u5_mult_87_n240) );
  INV_X4 u5_mult_87_U241 ( .A(fracta_mul[39]), .ZN(u5_mult_87_n249) );
  INV_X4 u5_mult_87_U240 ( .A(u5_mult_87_n455), .ZN(u5_mult_87_n247) );
  INV_X4 u5_mult_87_U239 ( .A(fracta_mul[34]), .ZN(u5_mult_87_n262) );
  INV_X4 u5_mult_87_U238 ( .A(fracta_mul[35]), .ZN(u5_mult_87_n260) );
  INV_X4 u5_mult_87_U237 ( .A(fracta_mul[35]), .ZN(u5_mult_87_n259) );
  INV_X4 u5_mult_87_U236 ( .A(fracta_mul[36]), .ZN(u5_mult_87_n256) );
  INV_X4 u5_mult_87_U235 ( .A(fracta_mul[36]), .ZN(u5_mult_87_n258) );
  INV_X4 u5_mult_87_U234 ( .A(fracta_mul[38]), .ZN(u5_mult_87_n253) );
  INV_X4 u5_mult_87_U233 ( .A(fracta_mul[30]), .ZN(u5_mult_87_n271) );
  INV_X4 u5_mult_87_U232 ( .A(fracta_mul[26]), .ZN(u5_mult_87_n279) );
  INV_X4 u5_mult_87_U231 ( .A(fracta_mul[32]), .ZN(u5_mult_87_n265) );
  INV_X4 u5_mult_87_U230 ( .A(fracta_mul[28]), .ZN(u5_mult_87_n275) );
  INV_X4 u5_mult_87_U229 ( .A(fracta_mul[29]), .ZN(u5_mult_87_n273) );
  INV_X4 u5_mult_87_U228 ( .A(fracta_mul[27]), .ZN(u5_mult_87_n278) );
  INV_X4 u5_mult_87_U227 ( .A(fracta_mul[31]), .ZN(u5_mult_87_n268) );
  INV_X4 u5_mult_87_U226 ( .A(fracta_mul[22]), .ZN(u5_mult_87_n287) );
  INV_X4 u5_mult_87_U225 ( .A(fracta_mul[23]), .ZN(u5_mult_87_n285) );
  INV_X4 u5_mult_87_U224 ( .A(fracta_mul[21]), .ZN(u5_mult_87_n289) );
  INV_X4 u5_mult_87_U223 ( .A(fracta_mul[24]), .ZN(u5_mult_87_n283) );
  INV_X4 u5_mult_87_U222 ( .A(fracta_mul[20]), .ZN(u5_mult_87_n291) );
  INV_X4 u5_mult_87_U221 ( .A(fracta_mul[18]), .ZN(u5_mult_87_n295) );
  INV_X4 u5_mult_87_U220 ( .A(fracta_mul[19]), .ZN(u5_mult_87_n292) );
  INV_X4 u5_mult_87_U219 ( .A(fracta_mul[19]), .ZN(u5_mult_87_n294) );
  INV_X4 u5_mult_87_U218 ( .A(u5_mult_87_n477), .ZN(u5_mult_87_n318) );
  INV_X4 u5_mult_87_U217 ( .A(u6_N17), .ZN(u5_mult_87_n414) );
  INV_X4 u5_mult_87_U216 ( .A(u6_N6), .ZN(u5_mult_87_n435) );
  INV_X4 u5_mult_87_U215 ( .A(u6_N7), .ZN(u5_mult_87_n433) );
  INV_X4 u5_mult_87_U214 ( .A(u6_N8), .ZN(u5_mult_87_n431) );
  INV_X4 u5_mult_87_U213 ( .A(u6_N3), .ZN(u5_mult_87_n442) );
  XOR2_X2 u5_mult_87_U212 ( .A(u5_mult_87_CARRYB_52__47_), .B(
        u5_mult_87_SUMB_52__48_), .Z(u5_mult_87_n103) );
  XOR2_X2 u5_mult_87_U211 ( .A(u5_mult_87_CARRYB_52__46_), .B(
        u5_mult_87_SUMB_52__47_), .Z(u5_mult_87_n102) );
  XOR2_X2 u5_mult_87_U210 ( .A(u5_mult_87_CARRYB_52__40_), .B(
        u5_mult_87_SUMB_52__41_), .Z(u5_mult_87_n101) );
  XOR2_X2 u5_mult_87_U209 ( .A(u5_mult_87_CARRYB_52__41_), .B(
        u5_mult_87_SUMB_52__42_), .Z(u5_mult_87_n100) );
  XOR2_X2 u5_mult_87_U208 ( .A(u5_mult_87_CARRYB_52__44_), .B(
        u5_mult_87_SUMB_52__45_), .Z(u5_mult_87_n99) );
  XOR2_X2 u5_mult_87_U207 ( .A(u5_mult_87_CARRYB_52__42_), .B(
        u5_mult_87_SUMB_52__43_), .Z(u5_mult_87_n98) );
  XOR2_X2 u5_mult_87_U206 ( .A(u5_mult_87_CARRYB_52__50_), .B(
        u5_mult_87_SUMB_52__51_), .Z(u5_mult_87_n97) );
  XOR2_X2 u5_mult_87_U205 ( .A(u5_mult_87_CARRYB_52__45_), .B(
        u5_mult_87_SUMB_52__46_), .Z(u5_mult_87_n96) );
  XOR2_X2 u5_mult_87_U204 ( .A(u5_mult_87_CARRYB_52__48_), .B(
        u5_mult_87_SUMB_52__49_), .Z(u5_mult_87_n95) );
  XOR2_X2 u5_mult_87_U203 ( .A(u5_mult_87_CARRYB_52__43_), .B(
        u5_mult_87_SUMB_52__44_), .Z(u5_mult_87_n94) );
  XOR2_X2 u5_mult_87_U202 ( .A(u5_mult_87_CARRYB_52__49_), .B(
        u5_mult_87_SUMB_52__50_), .Z(u5_mult_87_n93) );
  XOR2_X2 u5_mult_87_U201 ( .A(u5_mult_87_CARRYB_52__51_), .B(
        u5_mult_87_ab_52__52_), .Z(u5_mult_87_n92) );
  AND2_X4 u5_mult_87_U200 ( .A1(u5_mult_87_ab_0__1_), .A2(u5_mult_87_ab_1__0_), 
        .ZN(u5_mult_87_n91) );
  INV_X4 u5_mult_87_U199 ( .A(u6_N32), .ZN(u5_mult_87_n384) );
  INV_X4 u5_mult_87_U198 ( .A(u6_N10), .ZN(u5_mult_87_n428) );
  INV_X4 u5_mult_87_U197 ( .A(u6_N48), .ZN(u5_mult_87_n350) );
  INV_X4 u5_mult_87_U196 ( .A(u6_N40), .ZN(u5_mult_87_n368) );
  INV_X4 u5_mult_87_U195 ( .A(u6_N31), .ZN(u5_mult_87_n386) );
  INV_X4 u5_mult_87_U194 ( .A(u6_N33), .ZN(u5_mult_87_n382) );
  INV_X4 u5_mult_87_U193 ( .A(u6_N37), .ZN(u5_mult_87_n374) );
  INV_X4 u5_mult_87_U192 ( .A(u6_N39), .ZN(u5_mult_87_n370) );
  INV_X4 u5_mult_87_U191 ( .A(u6_N42), .ZN(u5_mult_87_n362) );
  INV_X4 u5_mult_87_U190 ( .A(u6_N42), .ZN(u5_mult_87_n363) );
  INV_X4 u5_mult_87_U189 ( .A(u6_N47), .ZN(u5_mult_87_n352) );
  INV_X4 u5_mult_87_U188 ( .A(u6_N47), .ZN(u5_mult_87_n353) );
  INV_X4 u5_mult_87_U187 ( .A(u6_N38), .ZN(u5_mult_87_n372) );
  INV_X4 u5_mult_87_U186 ( .A(u6_N21), .ZN(u5_mult_87_n405) );
  INV_X4 u5_mult_87_U185 ( .A(u6_N22), .ZN(u5_mult_87_n403) );
  INV_X4 u5_mult_87_U184 ( .A(u6_N22), .ZN(u5_mult_87_n404) );
  INV_X4 u5_mult_87_U183 ( .A(u6_N23), .ZN(u5_mult_87_n401) );
  INV_X4 u5_mult_87_U182 ( .A(u6_N25), .ZN(u5_mult_87_n397) );
  INV_X4 u5_mult_87_U181 ( .A(u6_N27), .ZN(u5_mult_87_n393) );
  INV_X4 u5_mult_87_U180 ( .A(u6_N28), .ZN(u5_mult_87_n391) );
  INV_X4 u5_mult_87_U179 ( .A(u6_N28), .ZN(u5_mult_87_n392) );
  INV_X4 u5_mult_87_U178 ( .A(u6_N29), .ZN(u5_mult_87_n389) );
  INV_X4 u5_mult_87_U177 ( .A(fracta_mul[0]), .ZN(u5_mult_87_n339) );
  INV_X4 u5_mult_87_U176 ( .A(u6_N52), .ZN(u5_mult_87_n343) );
  INV_X4 u5_mult_87_U175 ( .A(u6_N20), .ZN(u5_mult_87_n407) );
  INV_X4 u5_mult_87_U174 ( .A(u6_N24), .ZN(u5_mult_87_n399) );
  INV_X4 u5_mult_87_U173 ( .A(u6_N26), .ZN(u5_mult_87_n395) );
  INV_X4 u5_mult_87_U172 ( .A(fracta_mul[4]), .ZN(u5_mult_87_n326) );
  XOR2_X2 u5_mult_87_U171 ( .A(u5_mult_87_CARRYB_52__33_), .B(
        u5_mult_87_SUMB_52__34_), .Z(u5_mult_87_n90) );
  XOR2_X2 u5_mult_87_U170 ( .A(u5_mult_87_CARRYB_52__36_), .B(
        u5_mult_87_SUMB_52__37_), .Z(u5_mult_87_n89) );
  XOR2_X2 u5_mult_87_U169 ( .A(u5_mult_87_CARRYB_52__34_), .B(
        u5_mult_87_SUMB_52__35_), .Z(u5_mult_87_n88) );
  XOR2_X2 u5_mult_87_U168 ( .A(u5_mult_87_CARRYB_52__37_), .B(
        u5_mult_87_SUMB_52__38_), .Z(u5_mult_87_n87) );
  XOR2_X2 u5_mult_87_U167 ( .A(u5_mult_87_CARRYB_52__39_), .B(
        u5_mult_87_SUMB_52__40_), .Z(u5_mult_87_n86) );
  XOR2_X2 u5_mult_87_U166 ( .A(u5_mult_87_CARRYB_52__38_), .B(
        u5_mult_87_SUMB_52__39_), .Z(u5_mult_87_n85) );
  XOR2_X2 u5_mult_87_U165 ( .A(u5_mult_87_CARRYB_52__30_), .B(
        u5_mult_87_SUMB_52__31_), .Z(u5_mult_87_n84) );
  XOR2_X2 u5_mult_87_U164 ( .A(u5_mult_87_CARRYB_52__17_), .B(
        u5_mult_87_SUMB_52__18_), .Z(u5_mult_87_n83) );
  XOR2_X2 u5_mult_87_U163 ( .A(u5_mult_87_CARRYB_52__20_), .B(
        u5_mult_87_SUMB_52__21_), .Z(u5_mult_87_n82) );
  XOR2_X2 u5_mult_87_U162 ( .A(u5_mult_87_CARRYB_52__18_), .B(
        u5_mult_87_SUMB_52__19_), .Z(u5_mult_87_n81) );
  XOR2_X2 u5_mult_87_U161 ( .A(u5_mult_87_CARRYB_52__21_), .B(
        u5_mult_87_SUMB_52__22_), .Z(u5_mult_87_n80) );
  XOR2_X2 u5_mult_87_U160 ( .A(u5_mult_87_CARRYB_52__24_), .B(
        u5_mult_87_SUMB_52__25_), .Z(u5_mult_87_n79) );
  XOR2_X2 u5_mult_87_U159 ( .A(u5_mult_87_CARRYB_52__23_), .B(
        u5_mult_87_SUMB_52__24_), .Z(u5_mult_87_n78) );
  XOR2_X2 u5_mult_87_U158 ( .A(u5_mult_87_CARRYB_52__22_), .B(
        u5_mult_87_SUMB_52__23_), .Z(u5_mult_87_n77) );
  XOR2_X2 u5_mult_87_U157 ( .A(u5_mult_87_CARRYB_52__25_), .B(
        u5_mult_87_SUMB_52__26_), .Z(u5_mult_87_n76) );
  XOR2_X2 u5_mult_87_U156 ( .A(u5_mult_87_CARRYB_52__28_), .B(
        u5_mult_87_SUMB_52__29_), .Z(u5_mult_87_n75) );
  XOR2_X2 u5_mult_87_U155 ( .A(u5_mult_87_CARRYB_52__26_), .B(
        u5_mult_87_SUMB_52__27_), .Z(u5_mult_87_n74) );
  XOR2_X2 u5_mult_87_U154 ( .A(u5_mult_87_CARRYB_52__14_), .B(
        u5_mult_87_SUMB_52__15_), .Z(u5_mult_87_n73) );
  XOR2_X2 u5_mult_87_U153 ( .A(u5_mult_87_CARRYB_52__10_), .B(
        u5_mult_87_SUMB_52__11_), .Z(u5_mult_87_n72) );
  XOR2_X2 u5_mult_87_U152 ( .A(u5_mult_87_CARRYB_52__9_), .B(
        u5_mult_87_SUMB_52__10_), .Z(u5_mult_87_n71) );
  XOR2_X2 u5_mult_87_U151 ( .A(u5_mult_87_CARRYB_52__12_), .B(
        u5_mult_87_SUMB_52__13_), .Z(u5_mult_87_n70) );
  XOR2_X2 u5_mult_87_U150 ( .A(u5_mult_87_CARRYB_52__8_), .B(
        u5_mult_87_SUMB_52__9_), .Z(u5_mult_87_n69) );
  XOR2_X2 u5_mult_87_U149 ( .A(u5_mult_87_CARRYB_52__15_), .B(
        u5_mult_87_SUMB_52__16_), .Z(u5_mult_87_n68) );
  XOR2_X2 u5_mult_87_U148 ( .A(u5_mult_87_CARRYB_52__16_), .B(
        u5_mult_87_SUMB_52__17_), .Z(u5_mult_87_n67) );
  XOR2_X2 u5_mult_87_U147 ( .A(u5_mult_87_CARRYB_52__13_), .B(
        u5_mult_87_SUMB_52__14_), .Z(u5_mult_87_n66) );
  XOR2_X2 u5_mult_87_U146 ( .A(u5_mult_87_CARRYB_52__32_), .B(
        u5_mult_87_SUMB_52__33_), .Z(u5_mult_87_n65) );
  XOR2_X2 u5_mult_87_U145 ( .A(u5_mult_87_CARRYB_52__29_), .B(
        u5_mult_87_SUMB_52__30_), .Z(u5_mult_87_n64) );
  XOR2_X2 u5_mult_87_U144 ( .A(u5_mult_87_CARRYB_52__11_), .B(
        u5_mult_87_SUMB_52__12_), .Z(u5_mult_87_n63) );
  XOR2_X2 u5_mult_87_U143 ( .A(u5_mult_87_CARRYB_52__35_), .B(
        u5_mult_87_SUMB_52__36_), .Z(u5_mult_87_n62) );
  XOR2_X2 u5_mult_87_U142 ( .A(u5_mult_87_CARRYB_52__19_), .B(
        u5_mult_87_SUMB_52__20_), .Z(u5_mult_87_n61) );
  XOR2_X2 u5_mult_87_U141 ( .A(u5_mult_87_CARRYB_52__27_), .B(
        u5_mult_87_SUMB_52__28_), .Z(u5_mult_87_n60) );
  XOR2_X2 u5_mult_87_U140 ( .A(u5_mult_87_CARRYB_52__31_), .B(
        u5_mult_87_SUMB_52__32_), .Z(u5_mult_87_n59) );
  AND2_X4 u5_mult_87_U139 ( .A1(u5_mult_87_ab_0__5_), .A2(u5_mult_87_ab_1__4_), 
        .ZN(u5_mult_87_n58) );
  AND2_X4 u5_mult_87_U138 ( .A1(u5_mult_87_ab_0__6_), .A2(u5_mult_87_ab_1__5_), 
        .ZN(u5_mult_87_n57) );
  AND2_X4 u5_mult_87_U137 ( .A1(u5_mult_87_ab_0__7_), .A2(u5_mult_87_ab_1__6_), 
        .ZN(u5_mult_87_n56) );
  AND2_X4 u5_mult_87_U136 ( .A1(u5_mult_87_ab_0__8_), .A2(u5_mult_87_ab_1__7_), 
        .ZN(u5_mult_87_n55) );
  AND2_X4 u5_mult_87_U135 ( .A1(u5_mult_87_ab_0__9_), .A2(u5_mult_87_ab_1__8_), 
        .ZN(u5_mult_87_n54) );
  AND2_X4 u5_mult_87_U134 ( .A1(u5_mult_87_ab_0__10_), .A2(u5_mult_87_ab_1__9_), .ZN(u5_mult_87_n53) );
  AND2_X4 u5_mult_87_U133 ( .A1(u5_mult_87_ab_0__11_), .A2(
        u5_mult_87_ab_1__10_), .ZN(u5_mult_87_n52) );
  AND2_X4 u5_mult_87_U132 ( .A1(u5_mult_87_ab_0__12_), .A2(
        u5_mult_87_ab_1__11_), .ZN(u5_mult_87_n51) );
  AND2_X4 u5_mult_87_U131 ( .A1(u5_mult_87_ab_0__13_), .A2(
        u5_mult_87_ab_1__12_), .ZN(u5_mult_87_n50) );
  AND2_X4 u5_mult_87_U130 ( .A1(u5_mult_87_ab_0__14_), .A2(
        u5_mult_87_ab_1__13_), .ZN(u5_mult_87_n49) );
  AND2_X4 u5_mult_87_U129 ( .A1(u5_mult_87_ab_0__15_), .A2(
        u5_mult_87_ab_1__14_), .ZN(u5_mult_87_n48) );
  AND2_X4 u5_mult_87_U128 ( .A1(u5_mult_87_ab_0__16_), .A2(
        u5_mult_87_ab_1__15_), .ZN(u5_mult_87_n47) );
  AND2_X4 u5_mult_87_U127 ( .A1(u5_mult_87_ab_0__17_), .A2(
        u5_mult_87_ab_1__16_), .ZN(u5_mult_87_n46) );
  AND2_X4 u5_mult_87_U126 ( .A1(u5_mult_87_ab_0__18_), .A2(
        u5_mult_87_ab_1__17_), .ZN(u5_mult_87_n45) );
  AND2_X4 u5_mult_87_U125 ( .A1(u5_mult_87_ab_0__19_), .A2(
        u5_mult_87_ab_1__18_), .ZN(u5_mult_87_n44) );
  AND2_X4 u5_mult_87_U124 ( .A1(u5_mult_87_ab_0__20_), .A2(
        u5_mult_87_ab_1__19_), .ZN(u5_mult_87_n43) );
  AND2_X4 u5_mult_87_U123 ( .A1(u5_mult_87_ab_0__21_), .A2(
        u5_mult_87_ab_1__20_), .ZN(u5_mult_87_n42) );
  AND2_X4 u5_mult_87_U122 ( .A1(u5_mult_87_ab_0__22_), .A2(
        u5_mult_87_ab_1__21_), .ZN(u5_mult_87_n41) );
  AND2_X4 u5_mult_87_U121 ( .A1(u5_mult_87_ab_0__23_), .A2(
        u5_mult_87_ab_1__22_), .ZN(u5_mult_87_n40) );
  AND2_X4 u5_mult_87_U120 ( .A1(u5_mult_87_ab_0__24_), .A2(
        u5_mult_87_ab_1__23_), .ZN(u5_mult_87_n39) );
  AND2_X4 u5_mult_87_U119 ( .A1(u5_mult_87_ab_0__25_), .A2(
        u5_mult_87_ab_1__24_), .ZN(u5_mult_87_n38) );
  AND2_X4 u5_mult_87_U118 ( .A1(u5_mult_87_ab_0__26_), .A2(
        u5_mult_87_ab_1__25_), .ZN(u5_mult_87_n37) );
  AND2_X4 u5_mult_87_U117 ( .A1(u5_mult_87_ab_0__27_), .A2(
        u5_mult_87_ab_1__26_), .ZN(u5_mult_87_n36) );
  AND2_X4 u5_mult_87_U116 ( .A1(u5_mult_87_ab_0__28_), .A2(
        u5_mult_87_ab_1__27_), .ZN(u5_mult_87_n35) );
  AND2_X4 u5_mult_87_U115 ( .A1(u5_mult_87_ab_0__29_), .A2(
        u5_mult_87_ab_1__28_), .ZN(u5_mult_87_n34) );
  AND2_X4 u5_mult_87_U114 ( .A1(u5_mult_87_ab_0__4_), .A2(u5_mult_87_ab_1__3_), 
        .ZN(u5_mult_87_n33) );
  AND2_X4 u5_mult_87_U113 ( .A1(u5_mult_87_ab_0__2_), .A2(u5_mult_87_ab_1__1_), 
        .ZN(u5_mult_87_n32) );
  AND2_X4 u5_mult_87_U112 ( .A1(u5_mult_87_ab_0__3_), .A2(u5_mult_87_ab_1__2_), 
        .ZN(u5_mult_87_n31) );
  AND2_X4 u5_mult_87_U111 ( .A1(u5_mult_87_ab_0__30_), .A2(
        u5_mult_87_ab_1__29_), .ZN(u5_mult_87_n30) );
  AND2_X4 u5_mult_87_U110 ( .A1(u5_mult_87_ab_0__31_), .A2(
        u5_mult_87_ab_1__30_), .ZN(u5_mult_87_n29) );
  AND2_X4 u5_mult_87_U109 ( .A1(u5_mult_87_ab_0__32_), .A2(
        u5_mult_87_ab_1__31_), .ZN(u5_mult_87_n28) );
  AND2_X4 u5_mult_87_U108 ( .A1(u5_mult_87_ab_0__33_), .A2(
        u5_mult_87_ab_1__32_), .ZN(u5_mult_87_n27) );
  AND2_X4 u5_mult_87_U107 ( .A1(u5_mult_87_ab_0__34_), .A2(
        u5_mult_87_ab_1__33_), .ZN(u5_mult_87_n26) );
  AND2_X4 u5_mult_87_U106 ( .A1(u5_mult_87_ab_0__35_), .A2(
        u5_mult_87_ab_1__34_), .ZN(u5_mult_87_n25) );
  AND2_X4 u5_mult_87_U105 ( .A1(u5_mult_87_ab_0__36_), .A2(
        u5_mult_87_ab_1__35_), .ZN(u5_mult_87_n24) );
  AND2_X4 u5_mult_87_U104 ( .A1(u5_mult_87_ab_0__37_), .A2(
        u5_mult_87_ab_1__36_), .ZN(u5_mult_87_n23) );
  AND2_X4 u5_mult_87_U103 ( .A1(u5_mult_87_ab_0__38_), .A2(
        u5_mult_87_ab_1__37_), .ZN(u5_mult_87_n22) );
  AND2_X4 u5_mult_87_U102 ( .A1(u5_mult_87_ab_0__39_), .A2(
        u5_mult_87_ab_1__38_), .ZN(u5_mult_87_n21) );
  AND2_X4 u5_mult_87_U101 ( .A1(u5_mult_87_ab_0__40_), .A2(
        u5_mult_87_ab_1__39_), .ZN(u5_mult_87_n20) );
  AND2_X4 u5_mult_87_U100 ( .A1(u5_mult_87_ab_0__41_), .A2(
        u5_mult_87_ab_1__40_), .ZN(u5_mult_87_n19) );
  AND2_X4 u5_mult_87_U99 ( .A1(u5_mult_87_ab_0__42_), .A2(u5_mult_87_ab_1__41_), .ZN(u5_mult_87_n18) );
  AND2_X4 u5_mult_87_U98 ( .A1(u5_mult_87_ab_0__43_), .A2(u5_mult_87_ab_1__42_), .ZN(u5_mult_87_n17) );
  AND2_X4 u5_mult_87_U97 ( .A1(u5_mult_87_ab_0__44_), .A2(u5_mult_87_ab_1__43_), .ZN(u5_mult_87_n16) );
  AND2_X4 u5_mult_87_U96 ( .A1(u5_mult_87_ab_0__45_), .A2(u5_mult_87_ab_1__44_), .ZN(u5_mult_87_n15) );
  AND2_X4 u5_mult_87_U95 ( .A1(u5_mult_87_ab_0__46_), .A2(u5_mult_87_ab_1__45_), .ZN(u5_mult_87_n14) );
  AND2_X4 u5_mult_87_U94 ( .A1(u5_mult_87_ab_0__47_), .A2(u5_mult_87_ab_1__46_), .ZN(u5_mult_87_n13) );
  AND2_X4 u5_mult_87_U93 ( .A1(u5_mult_87_ab_0__48_), .A2(u5_mult_87_ab_1__47_), .ZN(u5_mult_87_n12) );
  AND2_X4 u5_mult_87_U92 ( .A1(u5_mult_87_ab_0__49_), .A2(u5_mult_87_ab_1__48_), .ZN(u5_mult_87_n11) );
  XOR2_X2 u5_mult_87_U91 ( .A(u5_mult_87_CARRYB_52__6_), .B(
        u5_mult_87_SUMB_52__7_), .Z(u5_mult_87_n10) );
  XOR2_X2 u5_mult_87_U90 ( .A(u5_mult_87_CARRYB_52__5_), .B(
        u5_mult_87_SUMB_52__6_), .Z(u5_mult_87_n9) );
  XOR2_X2 u5_mult_87_U89 ( .A(u5_mult_87_CARRYB_52__3_), .B(
        u5_mult_87_SUMB_52__4_), .Z(u5_mult_87_n8) );
  XOR2_X2 u5_mult_87_U88 ( .A(u5_mult_87_CARRYB_52__2_), .B(
        u5_mult_87_SUMB_52__3_), .Z(u5_mult_87_n7) );
  XOR2_X2 u5_mult_87_U87 ( .A(u5_mult_87_CARRYB_52__4_), .B(
        u5_mult_87_SUMB_52__5_), .Z(u5_mult_87_n6) );
  XOR2_X2 u5_mult_87_U86 ( .A(u5_mult_87_CARRYB_52__1_), .B(
        u5_mult_87_SUMB_52__2_), .Z(u5_mult_87_n5) );
  XOR2_X2 u5_mult_87_U85 ( .A(u5_mult_87_CARRYB_52__7_), .B(
        u5_mult_87_SUMB_52__8_), .Z(u5_mult_87_n4) );
  XOR2_X2 u5_mult_87_U84 ( .A(u5_mult_87_ab_1__51_), .B(u5_mult_87_ab_0__52_), 
        .Z(u5_mult_87_n3) );
  AND2_X4 u5_mult_87_U83 ( .A1(u5_mult_87_ab_0__50_), .A2(u5_mult_87_ab_1__49_), .ZN(u5_mult_87_n2) );
  INV_X4 u5_mult_87_U82 ( .A(fracta_mul[48]), .ZN(u5_mult_87_n219) );
  INV_X4 u5_mult_87_U81 ( .A(fracta_mul[47]), .ZN(u5_mult_87_n223) );
  INV_X4 u5_mult_87_U80 ( .A(fracta_mul[49]), .ZN(u5_mult_87_n216) );
  INV_X4 u5_mult_87_U79 ( .A(fracta_mul[50]), .ZN(u5_mult_87_n213) );
  INV_X4 u5_mult_87_U78 ( .A(fracta_mul[41]), .ZN(u5_mult_87_n243) );
  INV_X4 u5_mult_87_U77 ( .A(fracta_mul[45]), .ZN(u5_mult_87_n227) );
  INV_X4 u5_mult_87_U76 ( .A(fracta_mul[34]), .ZN(u5_mult_87_n261) );
  INV_X4 u5_mult_87_U75 ( .A(fracta_mul[39]), .ZN(u5_mult_87_n250) );
  INV_X4 u5_mult_87_U74 ( .A(fracta_mul[39]), .ZN(u5_mult_87_n248) );
  INV_X4 u5_mult_87_U73 ( .A(fracta_mul[30]), .ZN(u5_mult_87_n270) );
  INV_X4 u5_mult_87_U72 ( .A(fracta_mul[33]), .ZN(u5_mult_87_n264) );
  INV_X4 u5_mult_87_U71 ( .A(fracta_mul[32]), .ZN(u5_mult_87_n267) );
  INV_X4 u5_mult_87_U70 ( .A(fracta_mul[12]), .ZN(u5_mult_87_n306) );
  INV_X4 u5_mult_87_U69 ( .A(u6_N3), .ZN(u5_mult_87_n443) );
  INV_X4 u5_mult_87_U68 ( .A(u6_N1), .ZN(u5_mult_87_n446) );
  INV_X4 u5_mult_87_U67 ( .A(u6_N5), .ZN(u5_mult_87_n438) );
  INV_X4 u5_mult_87_U66 ( .A(u6_N2), .ZN(u5_mult_87_n444) );
  INV_X4 u5_mult_87_U65 ( .A(fracta_mul[6]), .ZN(u5_mult_87_n321) );
  INV_X4 u5_mult_87_U64 ( .A(fracta_mul[7]), .ZN(u5_mult_87_n319) );
  INV_X4 u5_mult_87_U63 ( .A(u6_N47), .ZN(u5_mult_87_n351) );
  INV_X4 u5_mult_87_U62 ( .A(u6_N42), .ZN(u5_mult_87_n364) );
  INV_X4 u5_mult_87_U61 ( .A(u6_N49), .ZN(u5_mult_87_n348) );
  INV_X4 u5_mult_87_U60 ( .A(u6_N12), .ZN(u5_mult_87_n424) );
  INV_X4 u5_mult_87_U59 ( .A(u6_N16), .ZN(u5_mult_87_n415) );
  INV_X4 u5_mult_87_U58 ( .A(u6_N50), .ZN(u5_mult_87_n346) );
  INV_X4 u5_mult_87_U57 ( .A(u6_N9), .ZN(u5_mult_87_n430) );
  INV_X4 u5_mult_87_U56 ( .A(u6_N21), .ZN(u5_mult_87_n406) );
  INV_X4 u5_mult_87_U55 ( .A(u6_N23), .ZN(u5_mult_87_n402) );
  INV_X4 u5_mult_87_U54 ( .A(u6_N25), .ZN(u5_mult_87_n398) );
  INV_X4 u5_mult_87_U53 ( .A(u6_N27), .ZN(u5_mult_87_n394) );
  INV_X4 u5_mult_87_U52 ( .A(u6_N29), .ZN(u5_mult_87_n390) );
  INV_X4 u5_mult_87_U51 ( .A(u6_N36), .ZN(u5_mult_87_n376) );
  INV_X4 u5_mult_87_U50 ( .A(u6_N51), .ZN(u5_mult_87_n345) );
  INV_X4 u5_mult_87_U49 ( .A(fracta_mul[3]), .ZN(u5_mult_87_n329) );
  INV_X4 u5_mult_87_U48 ( .A(fracta_mul[2]), .ZN(u5_mult_87_n332) );
  INV_X4 u5_mult_87_U47 ( .A(u6_N41), .ZN(u5_mult_87_n365) );
  INV_X4 u5_mult_87_U46 ( .A(u6_N43), .ZN(u5_mult_87_n360) );
  INV_X4 u5_mult_87_U45 ( .A(u6_N44), .ZN(u5_mult_87_n358) );
  INV_X4 u5_mult_87_U44 ( .A(u6_N45), .ZN(u5_mult_87_n356) );
  INV_X4 u5_mult_87_U43 ( .A(u6_N46), .ZN(u5_mult_87_n354) );
  INV_X4 u5_mult_87_U42 ( .A(u6_N30), .ZN(u5_mult_87_n387) );
  INV_X4 u5_mult_87_U41 ( .A(u6_N34), .ZN(u5_mult_87_n379) );
  INV_X4 u5_mult_87_U40 ( .A(u6_N35), .ZN(u5_mult_87_n377) );
  INV_X4 u5_mult_87_U39 ( .A(u6_N14), .ZN(u5_mult_87_n418) );
  INV_X4 u5_mult_87_U38 ( .A(fracta_mul[30]), .ZN(u5_mult_87_n272) );
  INV_X4 u5_mult_87_U37 ( .A(fracta_mul[27]), .ZN(u5_mult_87_n277) );
  INV_X4 u5_mult_87_U36 ( .A(fracta_mul[26]), .ZN(u5_mult_87_n280) );
  INV_X4 u5_mult_87_U35 ( .A(u6_N11), .ZN(u5_mult_87_n425) );
  INV_X4 u5_mult_87_U34 ( .A(u6_N4), .ZN(u5_mult_87_n441) );
  INV_X4 u5_mult_87_U33 ( .A(u6_N38), .ZN(u5_mult_87_n371) );
  INV_X4 u5_mult_87_U32 ( .A(u6_N10), .ZN(u5_mult_87_n427) );
  INV_X4 u5_mult_87_U31 ( .A(u6_N37), .ZN(u5_mult_87_n373) );
  INV_X4 u5_mult_87_U30 ( .A(u6_N17), .ZN(u5_mult_87_n413) );
  INV_X4 u5_mult_87_U29 ( .A(u6_N31), .ZN(u5_mult_87_n385) );
  INV_X4 u5_mult_87_U28 ( .A(u6_N32), .ZN(u5_mult_87_n383) );
  INV_X4 u5_mult_87_U27 ( .A(u6_N40), .ZN(u5_mult_87_n367) );
  INV_X4 u5_mult_87_U26 ( .A(u6_N33), .ZN(u5_mult_87_n381) );
  INV_X4 u5_mult_87_U25 ( .A(u6_N39), .ZN(u5_mult_87_n369) );
  INV_X4 u5_mult_87_U24 ( .A(u6_N18), .ZN(u5_mult_87_n411) );
  INV_X4 u5_mult_87_U23 ( .A(u6_N19), .ZN(u5_mult_87_n409) );
  INV_X4 u5_mult_87_U22 ( .A(u6_N15), .ZN(u5_mult_87_n416) );
  INV_X4 u5_mult_87_U21 ( .A(fracta_mul[14]), .ZN(u5_mult_87_n303) );
  INV_X4 u5_mult_87_U20 ( .A(fracta_mul[13]), .ZN(u5_mult_87_n305) );
  INV_X4 u5_mult_87_U19 ( .A(u6_N0), .ZN(u5_mult_87_n449) );
  INV_X4 u5_mult_87_U18 ( .A(u6_N48), .ZN(u5_mult_87_n349) );
  INV_X4 u5_mult_87_U17 ( .A(u6_N49), .ZN(u5_mult_87_n347) );
  INV_X4 u5_mult_87_U16 ( .A(u6_N9), .ZN(u5_mult_87_n429) );
  INV_X4 u5_mult_87_U15 ( .A(u6_N51), .ZN(u5_mult_87_n344) );
  INV_X4 u5_mult_87_U14 ( .A(u6_N36), .ZN(u5_mult_87_n375) );
  INV_X4 u5_mult_87_U13 ( .A(fracta_mul[6]), .ZN(u5_mult_87_n322) );
  INV_X4 u5_mult_87_U12 ( .A(u6_N13), .ZN(u5_mult_87_n422) );
  INV_X4 u5_mult_87_U11 ( .A(u6_N4), .ZN(u5_mult_87_n440) );
  INV_X4 u5_mult_87_U10 ( .A(fracta_mul[1]), .ZN(u5_mult_87_n336) );
  INV_X4 u5_mult_87_U9 ( .A(u6_N52), .ZN(u5_mult_87_n342) );
  INV_X4 u5_mult_87_U8 ( .A(fracta_mul[15]), .ZN(u5_mult_87_n302) );
  INV_X4 u5_mult_87_U7 ( .A(fracta_mul[17]), .ZN(u5_mult_87_n298) );
  INV_X4 u5_mult_87_U6 ( .A(fracta_mul[18]), .ZN(u5_mult_87_n296) );
  INV_X4 u5_mult_87_U5 ( .A(fracta_mul[16]), .ZN(u5_mult_87_n300) );
  INV_X4 u5_mult_87_U4 ( .A(u6_N5), .ZN(u5_mult_87_n437) );
  INV_X4 u5_mult_87_U3 ( .A(u6_N1), .ZN(u5_mult_87_n447) );
  INV_X4 u5_mult_87_U2 ( .A(u6_N14), .ZN(u5_mult_87_n419) );
  FA_X1 u5_mult_87_S3_2_51 ( .A(u5_mult_87_ab_2__51_), .B(u5_mult_87_n104), 
        .CI(u5_mult_87_ab_1__52_), .CO(u5_mult_87_CARRYB_2__51_), .S(
        u5_mult_87_SUMB_2__51_) );
  FA_X1 u5_mult_87_S2_2_50 ( .A(u5_mult_87_ab_2__50_), .B(u5_mult_87_n108), 
        .CI(u5_mult_87_n3), .CO(u5_mult_87_CARRYB_2__50_), .S(
        u5_mult_87_SUMB_2__50_) );
  FA_X1 u5_mult_87_S2_2_49 ( .A(u5_mult_87_ab_2__49_), .B(u5_mult_87_n2), .CI(
        u5_mult_87_n109), .CO(u5_mult_87_CARRYB_2__49_), .S(
        u5_mult_87_SUMB_2__49_) );
  FA_X1 u5_mult_87_S2_2_48 ( .A(u5_mult_87_ab_2__48_), .B(u5_mult_87_n11), 
        .CI(u5_mult_87_n110), .CO(u5_mult_87_CARRYB_2__48_), .S(
        u5_mult_87_SUMB_2__48_) );
  FA_X1 u5_mult_87_S2_2_47 ( .A(u5_mult_87_ab_2__47_), .B(u5_mult_87_n12), 
        .CI(u5_mult_87_n111), .CO(u5_mult_87_CARRYB_2__47_), .S(
        u5_mult_87_SUMB_2__47_) );
  FA_X1 u5_mult_87_S2_2_46 ( .A(u5_mult_87_ab_2__46_), .B(u5_mult_87_n13), 
        .CI(u5_mult_87_n112), .CO(u5_mult_87_CARRYB_2__46_), .S(
        u5_mult_87_SUMB_2__46_) );
  FA_X1 u5_mult_87_S2_2_45 ( .A(u5_mult_87_ab_2__45_), .B(u5_mult_87_n14), 
        .CI(u5_mult_87_n113), .CO(u5_mult_87_CARRYB_2__45_), .S(
        u5_mult_87_SUMB_2__45_) );
  FA_X1 u5_mult_87_S2_2_44 ( .A(u5_mult_87_ab_2__44_), .B(u5_mult_87_n15), 
        .CI(u5_mult_87_n114), .CO(u5_mult_87_CARRYB_2__44_), .S(
        u5_mult_87_SUMB_2__44_) );
  FA_X1 u5_mult_87_S2_2_43 ( .A(u5_mult_87_ab_2__43_), .B(u5_mult_87_n16), 
        .CI(u5_mult_87_n115), .CO(u5_mult_87_CARRYB_2__43_), .S(
        u5_mult_87_SUMB_2__43_) );
  FA_X1 u5_mult_87_S2_2_42 ( .A(u5_mult_87_ab_2__42_), .B(u5_mult_87_n17), 
        .CI(u5_mult_87_n116), .CO(u5_mult_87_CARRYB_2__42_), .S(
        u5_mult_87_SUMB_2__42_) );
  FA_X1 u5_mult_87_S2_2_41 ( .A(u5_mult_87_ab_2__41_), .B(u5_mult_87_n18), 
        .CI(u5_mult_87_n117), .CO(u5_mult_87_CARRYB_2__41_), .S(
        u5_mult_87_SUMB_2__41_) );
  FA_X1 u5_mult_87_S2_2_40 ( .A(u5_mult_87_ab_2__40_), .B(u5_mult_87_n19), 
        .CI(u5_mult_87_n118), .CO(u5_mult_87_CARRYB_2__40_), .S(
        u5_mult_87_SUMB_2__40_) );
  FA_X1 u5_mult_87_S2_2_39 ( .A(u5_mult_87_ab_2__39_), .B(u5_mult_87_n20), 
        .CI(u5_mult_87_n119), .CO(u5_mult_87_CARRYB_2__39_), .S(
        u5_mult_87_SUMB_2__39_) );
  FA_X1 u5_mult_87_S2_2_38 ( .A(u5_mult_87_ab_2__38_), .B(u5_mult_87_n21), 
        .CI(u5_mult_87_n120), .CO(u5_mult_87_CARRYB_2__38_), .S(
        u5_mult_87_SUMB_2__38_) );
  FA_X1 u5_mult_87_S2_2_37 ( .A(u5_mult_87_ab_2__37_), .B(u5_mult_87_n22), 
        .CI(u5_mult_87_n121), .CO(u5_mult_87_CARRYB_2__37_), .S(
        u5_mult_87_SUMB_2__37_) );
  FA_X1 u5_mult_87_S2_2_36 ( .A(u5_mult_87_ab_2__36_), .B(u5_mult_87_n23), 
        .CI(u5_mult_87_n122), .CO(u5_mult_87_CARRYB_2__36_), .S(
        u5_mult_87_SUMB_2__36_) );
  FA_X1 u5_mult_87_S2_2_35 ( .A(u5_mult_87_ab_2__35_), .B(u5_mult_87_n24), 
        .CI(u5_mult_87_n123), .CO(u5_mult_87_CARRYB_2__35_), .S(
        u5_mult_87_SUMB_2__35_) );
  FA_X1 u5_mult_87_S2_2_34 ( .A(u5_mult_87_ab_2__34_), .B(u5_mult_87_n25), 
        .CI(u5_mult_87_n124), .CO(u5_mult_87_CARRYB_2__34_), .S(
        u5_mult_87_SUMB_2__34_) );
  FA_X1 u5_mult_87_S2_2_33 ( .A(u5_mult_87_ab_2__33_), .B(u5_mult_87_n26), 
        .CI(u5_mult_87_n125), .CO(u5_mult_87_CARRYB_2__33_), .S(
        u5_mult_87_SUMB_2__33_) );
  FA_X1 u5_mult_87_S2_2_32 ( .A(u5_mult_87_ab_2__32_), .B(u5_mult_87_n27), 
        .CI(u5_mult_87_n126), .CO(u5_mult_87_CARRYB_2__32_), .S(
        u5_mult_87_SUMB_2__32_) );
  FA_X1 u5_mult_87_S2_2_31 ( .A(u5_mult_87_ab_2__31_), .B(u5_mult_87_n28), 
        .CI(u5_mult_87_n127), .CO(u5_mult_87_CARRYB_2__31_), .S(
        u5_mult_87_SUMB_2__31_) );
  FA_X1 u5_mult_87_S2_2_30 ( .A(u5_mult_87_ab_2__30_), .B(u5_mult_87_n29), 
        .CI(u5_mult_87_n128), .CO(u5_mult_87_CARRYB_2__30_), .S(
        u5_mult_87_SUMB_2__30_) );
  FA_X1 u5_mult_87_S2_2_29 ( .A(u5_mult_87_ab_2__29_), .B(u5_mult_87_n30), 
        .CI(u5_mult_87_n129), .CO(u5_mult_87_CARRYB_2__29_), .S(
        u5_mult_87_SUMB_2__29_) );
  FA_X1 u5_mult_87_S2_2_28 ( .A(u5_mult_87_ab_2__28_), .B(u5_mult_87_n34), 
        .CI(u5_mult_87_n130), .CO(u5_mult_87_CARRYB_2__28_), .S(
        u5_mult_87_SUMB_2__28_) );
  FA_X1 u5_mult_87_S2_2_27 ( .A(u5_mult_87_ab_2__27_), .B(u5_mult_87_n35), 
        .CI(u5_mult_87_n131), .CO(u5_mult_87_CARRYB_2__27_), .S(
        u5_mult_87_SUMB_2__27_) );
  FA_X1 u5_mult_87_S2_2_26 ( .A(u5_mult_87_ab_2__26_), .B(u5_mult_87_n36), 
        .CI(u5_mult_87_n132), .CO(u5_mult_87_CARRYB_2__26_), .S(
        u5_mult_87_SUMB_2__26_) );
  FA_X1 u5_mult_87_S2_2_25 ( .A(u5_mult_87_ab_2__25_), .B(u5_mult_87_n37), 
        .CI(u5_mult_87_n133), .CO(u5_mult_87_CARRYB_2__25_), .S(
        u5_mult_87_SUMB_2__25_) );
  FA_X1 u5_mult_87_S2_2_24 ( .A(u5_mult_87_ab_2__24_), .B(u5_mult_87_n38), 
        .CI(u5_mult_87_n134), .CO(u5_mult_87_CARRYB_2__24_), .S(
        u5_mult_87_SUMB_2__24_) );
  FA_X1 u5_mult_87_S2_2_23 ( .A(u5_mult_87_ab_2__23_), .B(u5_mult_87_n39), 
        .CI(u5_mult_87_n135), .CO(u5_mult_87_CARRYB_2__23_), .S(
        u5_mult_87_SUMB_2__23_) );
  FA_X1 u5_mult_87_S2_2_22 ( .A(u5_mult_87_ab_2__22_), .B(u5_mult_87_n40), 
        .CI(u5_mult_87_n136), .CO(u5_mult_87_CARRYB_2__22_), .S(
        u5_mult_87_SUMB_2__22_) );
  FA_X1 u5_mult_87_S2_2_21 ( .A(u5_mult_87_ab_2__21_), .B(u5_mult_87_n41), 
        .CI(u5_mult_87_n137), .CO(u5_mult_87_CARRYB_2__21_), .S(
        u5_mult_87_SUMB_2__21_) );
  FA_X1 u5_mult_87_S2_2_20 ( .A(u5_mult_87_ab_2__20_), .B(u5_mult_87_n42), 
        .CI(u5_mult_87_n138), .CO(u5_mult_87_CARRYB_2__20_), .S(
        u5_mult_87_SUMB_2__20_) );
  FA_X1 u5_mult_87_S2_2_19 ( .A(u5_mult_87_ab_2__19_), .B(u5_mult_87_n43), 
        .CI(u5_mult_87_n139), .CO(u5_mult_87_CARRYB_2__19_), .S(
        u5_mult_87_SUMB_2__19_) );
  FA_X1 u5_mult_87_S2_2_18 ( .A(u5_mult_87_ab_2__18_), .B(u5_mult_87_n44), 
        .CI(u5_mult_87_n140), .CO(u5_mult_87_CARRYB_2__18_), .S(
        u5_mult_87_SUMB_2__18_) );
  FA_X1 u5_mult_87_S2_2_17 ( .A(u5_mult_87_ab_2__17_), .B(u5_mult_87_n45), 
        .CI(u5_mult_87_n141), .CO(u5_mult_87_CARRYB_2__17_), .S(
        u5_mult_87_SUMB_2__17_) );
  FA_X1 u5_mult_87_S2_2_16 ( .A(u5_mult_87_ab_2__16_), .B(u5_mult_87_n46), 
        .CI(u5_mult_87_n142), .CO(u5_mult_87_CARRYB_2__16_), .S(
        u5_mult_87_SUMB_2__16_) );
  FA_X1 u5_mult_87_S2_2_15 ( .A(u5_mult_87_ab_2__15_), .B(u5_mult_87_n47), 
        .CI(u5_mult_87_n143), .CO(u5_mult_87_CARRYB_2__15_), .S(
        u5_mult_87_SUMB_2__15_) );
  FA_X1 u5_mult_87_S2_2_14 ( .A(u5_mult_87_ab_2__14_), .B(u5_mult_87_n48), 
        .CI(u5_mult_87_n144), .CO(u5_mult_87_CARRYB_2__14_), .S(
        u5_mult_87_SUMB_2__14_) );
  FA_X1 u5_mult_87_S2_2_13 ( .A(u5_mult_87_ab_2__13_), .B(u5_mult_87_n49), 
        .CI(u5_mult_87_n145), .CO(u5_mult_87_CARRYB_2__13_), .S(
        u5_mult_87_SUMB_2__13_) );
  FA_X1 u5_mult_87_S2_2_12 ( .A(u5_mult_87_ab_2__12_), .B(u5_mult_87_n50), 
        .CI(u5_mult_87_n146), .CO(u5_mult_87_CARRYB_2__12_), .S(
        u5_mult_87_SUMB_2__12_) );
  FA_X1 u5_mult_87_S2_2_11 ( .A(u5_mult_87_ab_2__11_), .B(u5_mult_87_n51), 
        .CI(u5_mult_87_n147), .CO(u5_mult_87_CARRYB_2__11_), .S(
        u5_mult_87_SUMB_2__11_) );
  FA_X1 u5_mult_87_S2_2_10 ( .A(u5_mult_87_ab_2__10_), .B(u5_mult_87_n52), 
        .CI(u5_mult_87_n148), .CO(u5_mult_87_CARRYB_2__10_), .S(
        u5_mult_87_SUMB_2__10_) );
  FA_X1 u5_mult_87_S2_2_9 ( .A(u5_mult_87_ab_2__9_), .B(u5_mult_87_n53), .CI(
        u5_mult_87_n149), .CO(u5_mult_87_CARRYB_2__9_), .S(
        u5_mult_87_SUMB_2__9_) );
  FA_X1 u5_mult_87_S2_2_8 ( .A(u5_mult_87_ab_2__8_), .B(u5_mult_87_n54), .CI(
        u5_mult_87_n150), .CO(u5_mult_87_CARRYB_2__8_), .S(
        u5_mult_87_SUMB_2__8_) );
  FA_X1 u5_mult_87_S2_2_7 ( .A(u5_mult_87_ab_2__7_), .B(u5_mult_87_n55), .CI(
        u5_mult_87_n151), .CO(u5_mult_87_CARRYB_2__7_), .S(
        u5_mult_87_SUMB_2__7_) );
  FA_X1 u5_mult_87_S2_2_6 ( .A(u5_mult_87_ab_2__6_), .B(u5_mult_87_n56), .CI(
        u5_mult_87_n152), .CO(u5_mult_87_CARRYB_2__6_), .S(
        u5_mult_87_SUMB_2__6_) );
  FA_X1 u5_mult_87_S2_2_5 ( .A(u5_mult_87_ab_2__5_), .B(u5_mult_87_n57), .CI(
        u5_mult_87_n153), .CO(u5_mult_87_CARRYB_2__5_), .S(
        u5_mult_87_SUMB_2__5_) );
  FA_X1 u5_mult_87_S2_2_4 ( .A(u5_mult_87_ab_2__4_), .B(u5_mult_87_n58), .CI(
        u5_mult_87_n154), .CO(u5_mult_87_CARRYB_2__4_), .S(
        u5_mult_87_SUMB_2__4_) );
  FA_X1 u5_mult_87_S2_2_3 ( .A(u5_mult_87_ab_2__3_), .B(u5_mult_87_n33), .CI(
        u5_mult_87_n155), .CO(u5_mult_87_CARRYB_2__3_), .S(
        u5_mult_87_SUMB_2__3_) );
  FA_X1 u5_mult_87_S2_2_2 ( .A(u5_mult_87_ab_2__2_), .B(u5_mult_87_n31), .CI(
        u5_mult_87_n156), .CO(u5_mult_87_CARRYB_2__2_), .S(
        u5_mult_87_SUMB_2__2_) );
  FA_X1 u5_mult_87_S2_2_1 ( .A(u5_mult_87_ab_2__1_), .B(u5_mult_87_n32), .CI(
        u5_mult_87_n157), .CO(u5_mult_87_CARRYB_2__1_), .S(
        u5_mult_87_SUMB_2__1_) );
  FA_X1 u5_mult_87_S1_2_0 ( .A(u5_mult_87_ab_2__0_), .B(u5_mult_87_n91), .CI(
        u5_mult_87_n188), .CO(u5_mult_87_CARRYB_2__0_), .S(u5_N2) );
  FA_X1 u5_mult_87_S3_3_51 ( .A(u5_mult_87_ab_3__51_), .B(
        u5_mult_87_CARRYB_2__51_), .CI(u5_mult_87_ab_2__52_), .CO(
        u5_mult_87_CARRYB_3__51_), .S(u5_mult_87_SUMB_3__51_) );
  FA_X1 u5_mult_87_S2_3_50 ( .A(u5_mult_87_ab_3__50_), .B(
        u5_mult_87_CARRYB_2__50_), .CI(u5_mult_87_SUMB_2__51_), .CO(
        u5_mult_87_CARRYB_3__50_), .S(u5_mult_87_SUMB_3__50_) );
  FA_X1 u5_mult_87_S2_3_49 ( .A(u5_mult_87_ab_3__49_), .B(
        u5_mult_87_CARRYB_2__49_), .CI(u5_mult_87_SUMB_2__50_), .CO(
        u5_mult_87_CARRYB_3__49_), .S(u5_mult_87_SUMB_3__49_) );
  FA_X1 u5_mult_87_S2_3_48 ( .A(u5_mult_87_ab_3__48_), .B(
        u5_mult_87_CARRYB_2__48_), .CI(u5_mult_87_SUMB_2__49_), .CO(
        u5_mult_87_CARRYB_3__48_), .S(u5_mult_87_SUMB_3__48_) );
  FA_X1 u5_mult_87_S2_3_47 ( .A(u5_mult_87_ab_3__47_), .B(
        u5_mult_87_CARRYB_2__47_), .CI(u5_mult_87_SUMB_2__48_), .CO(
        u5_mult_87_CARRYB_3__47_), .S(u5_mult_87_SUMB_3__47_) );
  FA_X1 u5_mult_87_S2_3_46 ( .A(u5_mult_87_ab_3__46_), .B(
        u5_mult_87_CARRYB_2__46_), .CI(u5_mult_87_SUMB_2__47_), .CO(
        u5_mult_87_CARRYB_3__46_), .S(u5_mult_87_SUMB_3__46_) );
  FA_X1 u5_mult_87_S2_3_45 ( .A(u5_mult_87_ab_3__45_), .B(
        u5_mult_87_CARRYB_2__45_), .CI(u5_mult_87_SUMB_2__46_), .CO(
        u5_mult_87_CARRYB_3__45_), .S(u5_mult_87_SUMB_3__45_) );
  FA_X1 u5_mult_87_S2_3_44 ( .A(u5_mult_87_ab_3__44_), .B(
        u5_mult_87_CARRYB_2__44_), .CI(u5_mult_87_SUMB_2__45_), .CO(
        u5_mult_87_CARRYB_3__44_), .S(u5_mult_87_SUMB_3__44_) );
  FA_X1 u5_mult_87_S2_3_43 ( .A(u5_mult_87_ab_3__43_), .B(
        u5_mult_87_CARRYB_2__43_), .CI(u5_mult_87_SUMB_2__44_), .CO(
        u5_mult_87_CARRYB_3__43_), .S(u5_mult_87_SUMB_3__43_) );
  FA_X1 u5_mult_87_S2_3_42 ( .A(u5_mult_87_ab_3__42_), .B(
        u5_mult_87_CARRYB_2__42_), .CI(u5_mult_87_SUMB_2__43_), .CO(
        u5_mult_87_CARRYB_3__42_), .S(u5_mult_87_SUMB_3__42_) );
  FA_X1 u5_mult_87_S2_3_41 ( .A(u5_mult_87_ab_3__41_), .B(
        u5_mult_87_CARRYB_2__41_), .CI(u5_mult_87_SUMB_2__42_), .CO(
        u5_mult_87_CARRYB_3__41_), .S(u5_mult_87_SUMB_3__41_) );
  FA_X1 u5_mult_87_S2_3_40 ( .A(u5_mult_87_ab_3__40_), .B(
        u5_mult_87_CARRYB_2__40_), .CI(u5_mult_87_SUMB_2__41_), .CO(
        u5_mult_87_CARRYB_3__40_), .S(u5_mult_87_SUMB_3__40_) );
  FA_X1 u5_mult_87_S2_3_39 ( .A(u5_mult_87_ab_3__39_), .B(
        u5_mult_87_CARRYB_2__39_), .CI(u5_mult_87_SUMB_2__40_), .CO(
        u5_mult_87_CARRYB_3__39_), .S(u5_mult_87_SUMB_3__39_) );
  FA_X1 u5_mult_87_S2_3_38 ( .A(u5_mult_87_ab_3__38_), .B(
        u5_mult_87_CARRYB_2__38_), .CI(u5_mult_87_SUMB_2__39_), .CO(
        u5_mult_87_CARRYB_3__38_), .S(u5_mult_87_SUMB_3__38_) );
  FA_X1 u5_mult_87_S2_3_37 ( .A(u5_mult_87_ab_3__37_), .B(
        u5_mult_87_CARRYB_2__37_), .CI(u5_mult_87_SUMB_2__38_), .CO(
        u5_mult_87_CARRYB_3__37_), .S(u5_mult_87_SUMB_3__37_) );
  FA_X1 u5_mult_87_S2_3_36 ( .A(u5_mult_87_ab_3__36_), .B(
        u5_mult_87_CARRYB_2__36_), .CI(u5_mult_87_SUMB_2__37_), .CO(
        u5_mult_87_CARRYB_3__36_), .S(u5_mult_87_SUMB_3__36_) );
  FA_X1 u5_mult_87_S2_3_35 ( .A(u5_mult_87_ab_3__35_), .B(
        u5_mult_87_CARRYB_2__35_), .CI(u5_mult_87_SUMB_2__36_), .CO(
        u5_mult_87_CARRYB_3__35_), .S(u5_mult_87_SUMB_3__35_) );
  FA_X1 u5_mult_87_S2_3_34 ( .A(u5_mult_87_ab_3__34_), .B(
        u5_mult_87_CARRYB_2__34_), .CI(u5_mult_87_SUMB_2__35_), .CO(
        u5_mult_87_CARRYB_3__34_), .S(u5_mult_87_SUMB_3__34_) );
  FA_X1 u5_mult_87_S2_3_33 ( .A(u5_mult_87_ab_3__33_), .B(
        u5_mult_87_CARRYB_2__33_), .CI(u5_mult_87_SUMB_2__34_), .CO(
        u5_mult_87_CARRYB_3__33_), .S(u5_mult_87_SUMB_3__33_) );
  FA_X1 u5_mult_87_S2_3_32 ( .A(u5_mult_87_ab_3__32_), .B(
        u5_mult_87_CARRYB_2__32_), .CI(u5_mult_87_SUMB_2__33_), .CO(
        u5_mult_87_CARRYB_3__32_), .S(u5_mult_87_SUMB_3__32_) );
  FA_X1 u5_mult_87_S2_3_31 ( .A(u5_mult_87_ab_3__31_), .B(
        u5_mult_87_CARRYB_2__31_), .CI(u5_mult_87_SUMB_2__32_), .CO(
        u5_mult_87_CARRYB_3__31_), .S(u5_mult_87_SUMB_3__31_) );
  FA_X1 u5_mult_87_S2_3_30 ( .A(u5_mult_87_ab_3__30_), .B(
        u5_mult_87_CARRYB_2__30_), .CI(u5_mult_87_SUMB_2__31_), .CO(
        u5_mult_87_CARRYB_3__30_), .S(u5_mult_87_SUMB_3__30_) );
  FA_X1 u5_mult_87_S2_3_29 ( .A(u5_mult_87_ab_3__29_), .B(
        u5_mult_87_CARRYB_2__29_), .CI(u5_mult_87_SUMB_2__30_), .CO(
        u5_mult_87_CARRYB_3__29_), .S(u5_mult_87_SUMB_3__29_) );
  FA_X1 u5_mult_87_S2_3_28 ( .A(u5_mult_87_ab_3__28_), .B(
        u5_mult_87_CARRYB_2__28_), .CI(u5_mult_87_SUMB_2__29_), .CO(
        u5_mult_87_CARRYB_3__28_), .S(u5_mult_87_SUMB_3__28_) );
  FA_X1 u5_mult_87_S2_3_27 ( .A(u5_mult_87_ab_3__27_), .B(
        u5_mult_87_CARRYB_2__27_), .CI(u5_mult_87_SUMB_2__28_), .CO(
        u5_mult_87_CARRYB_3__27_), .S(u5_mult_87_SUMB_3__27_) );
  FA_X1 u5_mult_87_S2_3_26 ( .A(u5_mult_87_ab_3__26_), .B(
        u5_mult_87_CARRYB_2__26_), .CI(u5_mult_87_SUMB_2__27_), .CO(
        u5_mult_87_CARRYB_3__26_), .S(u5_mult_87_SUMB_3__26_) );
  FA_X1 u5_mult_87_S2_3_25 ( .A(u5_mult_87_ab_3__25_), .B(
        u5_mult_87_CARRYB_2__25_), .CI(u5_mult_87_SUMB_2__26_), .CO(
        u5_mult_87_CARRYB_3__25_), .S(u5_mult_87_SUMB_3__25_) );
  FA_X1 u5_mult_87_S2_3_24 ( .A(u5_mult_87_ab_3__24_), .B(
        u5_mult_87_CARRYB_2__24_), .CI(u5_mult_87_SUMB_2__25_), .CO(
        u5_mult_87_CARRYB_3__24_), .S(u5_mult_87_SUMB_3__24_) );
  FA_X1 u5_mult_87_S2_3_23 ( .A(u5_mult_87_ab_3__23_), .B(
        u5_mult_87_CARRYB_2__23_), .CI(u5_mult_87_SUMB_2__24_), .CO(
        u5_mult_87_CARRYB_3__23_), .S(u5_mult_87_SUMB_3__23_) );
  FA_X1 u5_mult_87_S2_3_22 ( .A(u5_mult_87_ab_3__22_), .B(
        u5_mult_87_CARRYB_2__22_), .CI(u5_mult_87_SUMB_2__23_), .CO(
        u5_mult_87_CARRYB_3__22_), .S(u5_mult_87_SUMB_3__22_) );
  FA_X1 u5_mult_87_S2_3_21 ( .A(u5_mult_87_ab_3__21_), .B(
        u5_mult_87_CARRYB_2__21_), .CI(u5_mult_87_SUMB_2__22_), .CO(
        u5_mult_87_CARRYB_3__21_), .S(u5_mult_87_SUMB_3__21_) );
  FA_X1 u5_mult_87_S2_3_20 ( .A(u5_mult_87_ab_3__20_), .B(
        u5_mult_87_CARRYB_2__20_), .CI(u5_mult_87_SUMB_2__21_), .CO(
        u5_mult_87_CARRYB_3__20_), .S(u5_mult_87_SUMB_3__20_) );
  FA_X1 u5_mult_87_S2_3_19 ( .A(u5_mult_87_ab_3__19_), .B(
        u5_mult_87_CARRYB_2__19_), .CI(u5_mult_87_SUMB_2__20_), .CO(
        u5_mult_87_CARRYB_3__19_), .S(u5_mult_87_SUMB_3__19_) );
  FA_X1 u5_mult_87_S2_3_18 ( .A(u5_mult_87_ab_3__18_), .B(
        u5_mult_87_CARRYB_2__18_), .CI(u5_mult_87_SUMB_2__19_), .CO(
        u5_mult_87_CARRYB_3__18_), .S(u5_mult_87_SUMB_3__18_) );
  FA_X1 u5_mult_87_S2_3_17 ( .A(u5_mult_87_ab_3__17_), .B(
        u5_mult_87_CARRYB_2__17_), .CI(u5_mult_87_SUMB_2__18_), .CO(
        u5_mult_87_CARRYB_3__17_), .S(u5_mult_87_SUMB_3__17_) );
  FA_X1 u5_mult_87_S2_3_16 ( .A(u5_mult_87_ab_3__16_), .B(
        u5_mult_87_CARRYB_2__16_), .CI(u5_mult_87_SUMB_2__17_), .CO(
        u5_mult_87_CARRYB_3__16_), .S(u5_mult_87_SUMB_3__16_) );
  FA_X1 u5_mult_87_S2_3_15 ( .A(u5_mult_87_ab_3__15_), .B(
        u5_mult_87_CARRYB_2__15_), .CI(u5_mult_87_SUMB_2__16_), .CO(
        u5_mult_87_CARRYB_3__15_), .S(u5_mult_87_SUMB_3__15_) );
  FA_X1 u5_mult_87_S2_3_14 ( .A(u5_mult_87_ab_3__14_), .B(
        u5_mult_87_CARRYB_2__14_), .CI(u5_mult_87_SUMB_2__15_), .CO(
        u5_mult_87_CARRYB_3__14_), .S(u5_mult_87_SUMB_3__14_) );
  FA_X1 u5_mult_87_S2_3_13 ( .A(u5_mult_87_ab_3__13_), .B(
        u5_mult_87_CARRYB_2__13_), .CI(u5_mult_87_SUMB_2__14_), .CO(
        u5_mult_87_CARRYB_3__13_), .S(u5_mult_87_SUMB_3__13_) );
  FA_X1 u5_mult_87_S2_3_12 ( .A(u5_mult_87_ab_3__12_), .B(
        u5_mult_87_CARRYB_2__12_), .CI(u5_mult_87_SUMB_2__13_), .CO(
        u5_mult_87_CARRYB_3__12_), .S(u5_mult_87_SUMB_3__12_) );
  FA_X1 u5_mult_87_S2_3_11 ( .A(u5_mult_87_ab_3__11_), .B(
        u5_mult_87_CARRYB_2__11_), .CI(u5_mult_87_SUMB_2__12_), .CO(
        u5_mult_87_CARRYB_3__11_), .S(u5_mult_87_SUMB_3__11_) );
  FA_X1 u5_mult_87_S2_3_10 ( .A(u5_mult_87_ab_3__10_), .B(
        u5_mult_87_CARRYB_2__10_), .CI(u5_mult_87_SUMB_2__11_), .CO(
        u5_mult_87_CARRYB_3__10_), .S(u5_mult_87_SUMB_3__10_) );
  FA_X1 u5_mult_87_S2_3_9 ( .A(u5_mult_87_ab_3__9_), .B(
        u5_mult_87_CARRYB_2__9_), .CI(u5_mult_87_SUMB_2__10_), .CO(
        u5_mult_87_CARRYB_3__9_), .S(u5_mult_87_SUMB_3__9_) );
  FA_X1 u5_mult_87_S2_3_8 ( .A(u5_mult_87_ab_3__8_), .B(
        u5_mult_87_CARRYB_2__8_), .CI(u5_mult_87_SUMB_2__9_), .CO(
        u5_mult_87_CARRYB_3__8_), .S(u5_mult_87_SUMB_3__8_) );
  FA_X1 u5_mult_87_S2_3_7 ( .A(u5_mult_87_ab_3__7_), .B(
        u5_mult_87_CARRYB_2__7_), .CI(u5_mult_87_SUMB_2__8_), .CO(
        u5_mult_87_CARRYB_3__7_), .S(u5_mult_87_SUMB_3__7_) );
  FA_X1 u5_mult_87_S2_3_6 ( .A(u5_mult_87_ab_3__6_), .B(
        u5_mult_87_CARRYB_2__6_), .CI(u5_mult_87_SUMB_2__7_), .CO(
        u5_mult_87_CARRYB_3__6_), .S(u5_mult_87_SUMB_3__6_) );
  FA_X1 u5_mult_87_S2_3_5 ( .A(u5_mult_87_ab_3__5_), .B(
        u5_mult_87_CARRYB_2__5_), .CI(u5_mult_87_SUMB_2__6_), .CO(
        u5_mult_87_CARRYB_3__5_), .S(u5_mult_87_SUMB_3__5_) );
  FA_X1 u5_mult_87_S2_3_4 ( .A(u5_mult_87_ab_3__4_), .B(
        u5_mult_87_CARRYB_2__4_), .CI(u5_mult_87_SUMB_2__5_), .CO(
        u5_mult_87_CARRYB_3__4_), .S(u5_mult_87_SUMB_3__4_) );
  FA_X1 u5_mult_87_S2_3_3 ( .A(u5_mult_87_ab_3__3_), .B(
        u5_mult_87_CARRYB_2__3_), .CI(u5_mult_87_SUMB_2__4_), .CO(
        u5_mult_87_CARRYB_3__3_), .S(u5_mult_87_SUMB_3__3_) );
  FA_X1 u5_mult_87_S2_3_2 ( .A(u5_mult_87_ab_3__2_), .B(
        u5_mult_87_CARRYB_2__2_), .CI(u5_mult_87_SUMB_2__3_), .CO(
        u5_mult_87_CARRYB_3__2_), .S(u5_mult_87_SUMB_3__2_) );
  FA_X1 u5_mult_87_S2_3_1 ( .A(u5_mult_87_ab_3__1_), .B(
        u5_mult_87_CARRYB_2__1_), .CI(u5_mult_87_SUMB_2__2_), .CO(
        u5_mult_87_CARRYB_3__1_), .S(u5_mult_87_SUMB_3__1_) );
  FA_X1 u5_mult_87_S1_3_0 ( .A(u5_mult_87_ab_3__0_), .B(
        u5_mult_87_CARRYB_2__0_), .CI(u5_mult_87_SUMB_2__1_), .CO(
        u5_mult_87_CARRYB_3__0_), .S(u5_N3) );
  FA_X1 u5_mult_87_S3_4_51 ( .A(u5_mult_87_ab_4__51_), .B(
        u5_mult_87_CARRYB_3__51_), .CI(u5_mult_87_ab_3__52_), .CO(
        u5_mult_87_CARRYB_4__51_), .S(u5_mult_87_SUMB_4__51_) );
  FA_X1 u5_mult_87_S2_4_50 ( .A(u5_mult_87_ab_4__50_), .B(
        u5_mult_87_CARRYB_3__50_), .CI(u5_mult_87_SUMB_3__51_), .CO(
        u5_mult_87_CARRYB_4__50_), .S(u5_mult_87_SUMB_4__50_) );
  FA_X1 u5_mult_87_S2_4_49 ( .A(u5_mult_87_ab_4__49_), .B(
        u5_mult_87_CARRYB_3__49_), .CI(u5_mult_87_SUMB_3__50_), .CO(
        u5_mult_87_CARRYB_4__49_), .S(u5_mult_87_SUMB_4__49_) );
  FA_X1 u5_mult_87_S2_4_48 ( .A(u5_mult_87_ab_4__48_), .B(
        u5_mult_87_CARRYB_3__48_), .CI(u5_mult_87_SUMB_3__49_), .CO(
        u5_mult_87_CARRYB_4__48_), .S(u5_mult_87_SUMB_4__48_) );
  FA_X1 u5_mult_87_S2_4_47 ( .A(u5_mult_87_ab_4__47_), .B(
        u5_mult_87_CARRYB_3__47_), .CI(u5_mult_87_SUMB_3__48_), .CO(
        u5_mult_87_CARRYB_4__47_), .S(u5_mult_87_SUMB_4__47_) );
  FA_X1 u5_mult_87_S2_4_46 ( .A(u5_mult_87_ab_4__46_), .B(
        u5_mult_87_CARRYB_3__46_), .CI(u5_mult_87_SUMB_3__47_), .CO(
        u5_mult_87_CARRYB_4__46_), .S(u5_mult_87_SUMB_4__46_) );
  FA_X1 u5_mult_87_S2_4_45 ( .A(u5_mult_87_ab_4__45_), .B(
        u5_mult_87_CARRYB_3__45_), .CI(u5_mult_87_SUMB_3__46_), .CO(
        u5_mult_87_CARRYB_4__45_), .S(u5_mult_87_SUMB_4__45_) );
  FA_X1 u5_mult_87_S2_4_44 ( .A(u5_mult_87_ab_4__44_), .B(
        u5_mult_87_CARRYB_3__44_), .CI(u5_mult_87_SUMB_3__45_), .CO(
        u5_mult_87_CARRYB_4__44_), .S(u5_mult_87_SUMB_4__44_) );
  FA_X1 u5_mult_87_S2_4_43 ( .A(u5_mult_87_ab_4__43_), .B(
        u5_mult_87_CARRYB_3__43_), .CI(u5_mult_87_SUMB_3__44_), .CO(
        u5_mult_87_CARRYB_4__43_), .S(u5_mult_87_SUMB_4__43_) );
  FA_X1 u5_mult_87_S2_4_42 ( .A(u5_mult_87_ab_4__42_), .B(
        u5_mult_87_CARRYB_3__42_), .CI(u5_mult_87_SUMB_3__43_), .CO(
        u5_mult_87_CARRYB_4__42_), .S(u5_mult_87_SUMB_4__42_) );
  FA_X1 u5_mult_87_S2_4_41 ( .A(u5_mult_87_ab_4__41_), .B(
        u5_mult_87_CARRYB_3__41_), .CI(u5_mult_87_SUMB_3__42_), .CO(
        u5_mult_87_CARRYB_4__41_), .S(u5_mult_87_SUMB_4__41_) );
  FA_X1 u5_mult_87_S2_4_40 ( .A(u5_mult_87_ab_4__40_), .B(
        u5_mult_87_CARRYB_3__40_), .CI(u5_mult_87_SUMB_3__41_), .CO(
        u5_mult_87_CARRYB_4__40_), .S(u5_mult_87_SUMB_4__40_) );
  FA_X1 u5_mult_87_S2_4_39 ( .A(u5_mult_87_ab_4__39_), .B(
        u5_mult_87_CARRYB_3__39_), .CI(u5_mult_87_SUMB_3__40_), .CO(
        u5_mult_87_CARRYB_4__39_), .S(u5_mult_87_SUMB_4__39_) );
  FA_X1 u5_mult_87_S2_4_38 ( .A(u5_mult_87_ab_4__38_), .B(
        u5_mult_87_CARRYB_3__38_), .CI(u5_mult_87_SUMB_3__39_), .CO(
        u5_mult_87_CARRYB_4__38_), .S(u5_mult_87_SUMB_4__38_) );
  FA_X1 u5_mult_87_S2_4_37 ( .A(u5_mult_87_ab_4__37_), .B(
        u5_mult_87_CARRYB_3__37_), .CI(u5_mult_87_SUMB_3__38_), .CO(
        u5_mult_87_CARRYB_4__37_), .S(u5_mult_87_SUMB_4__37_) );
  FA_X1 u5_mult_87_S2_4_36 ( .A(u5_mult_87_ab_4__36_), .B(
        u5_mult_87_CARRYB_3__36_), .CI(u5_mult_87_SUMB_3__37_), .CO(
        u5_mult_87_CARRYB_4__36_), .S(u5_mult_87_SUMB_4__36_) );
  FA_X1 u5_mult_87_S2_4_35 ( .A(u5_mult_87_ab_4__35_), .B(
        u5_mult_87_CARRYB_3__35_), .CI(u5_mult_87_SUMB_3__36_), .CO(
        u5_mult_87_CARRYB_4__35_), .S(u5_mult_87_SUMB_4__35_) );
  FA_X1 u5_mult_87_S2_4_34 ( .A(u5_mult_87_ab_4__34_), .B(
        u5_mult_87_CARRYB_3__34_), .CI(u5_mult_87_SUMB_3__35_), .CO(
        u5_mult_87_CARRYB_4__34_), .S(u5_mult_87_SUMB_4__34_) );
  FA_X1 u5_mult_87_S2_4_33 ( .A(u5_mult_87_ab_4__33_), .B(
        u5_mult_87_CARRYB_3__33_), .CI(u5_mult_87_SUMB_3__34_), .CO(
        u5_mult_87_CARRYB_4__33_), .S(u5_mult_87_SUMB_4__33_) );
  FA_X1 u5_mult_87_S2_4_32 ( .A(u5_mult_87_ab_4__32_), .B(
        u5_mult_87_CARRYB_3__32_), .CI(u5_mult_87_SUMB_3__33_), .CO(
        u5_mult_87_CARRYB_4__32_), .S(u5_mult_87_SUMB_4__32_) );
  FA_X1 u5_mult_87_S2_4_31 ( .A(u5_mult_87_ab_4__31_), .B(
        u5_mult_87_CARRYB_3__31_), .CI(u5_mult_87_SUMB_3__32_), .CO(
        u5_mult_87_CARRYB_4__31_), .S(u5_mult_87_SUMB_4__31_) );
  FA_X1 u5_mult_87_S2_4_30 ( .A(u5_mult_87_ab_4__30_), .B(
        u5_mult_87_CARRYB_3__30_), .CI(u5_mult_87_SUMB_3__31_), .CO(
        u5_mult_87_CARRYB_4__30_), .S(u5_mult_87_SUMB_4__30_) );
  FA_X1 u5_mult_87_S2_4_29 ( .A(u5_mult_87_ab_4__29_), .B(
        u5_mult_87_CARRYB_3__29_), .CI(u5_mult_87_SUMB_3__30_), .CO(
        u5_mult_87_CARRYB_4__29_), .S(u5_mult_87_SUMB_4__29_) );
  FA_X1 u5_mult_87_S2_4_28 ( .A(u5_mult_87_ab_4__28_), .B(
        u5_mult_87_CARRYB_3__28_), .CI(u5_mult_87_SUMB_3__29_), .CO(
        u5_mult_87_CARRYB_4__28_), .S(u5_mult_87_SUMB_4__28_) );
  FA_X1 u5_mult_87_S2_4_27 ( .A(u5_mult_87_ab_4__27_), .B(
        u5_mult_87_CARRYB_3__27_), .CI(u5_mult_87_SUMB_3__28_), .CO(
        u5_mult_87_CARRYB_4__27_), .S(u5_mult_87_SUMB_4__27_) );
  FA_X1 u5_mult_87_S2_4_26 ( .A(u5_mult_87_ab_4__26_), .B(
        u5_mult_87_CARRYB_3__26_), .CI(u5_mult_87_SUMB_3__27_), .CO(
        u5_mult_87_CARRYB_4__26_), .S(u5_mult_87_SUMB_4__26_) );
  FA_X1 u5_mult_87_S2_4_25 ( .A(u5_mult_87_ab_4__25_), .B(
        u5_mult_87_CARRYB_3__25_), .CI(u5_mult_87_SUMB_3__26_), .CO(
        u5_mult_87_CARRYB_4__25_), .S(u5_mult_87_SUMB_4__25_) );
  FA_X1 u5_mult_87_S2_4_24 ( .A(u5_mult_87_ab_4__24_), .B(
        u5_mult_87_CARRYB_3__24_), .CI(u5_mult_87_SUMB_3__25_), .CO(
        u5_mult_87_CARRYB_4__24_), .S(u5_mult_87_SUMB_4__24_) );
  FA_X1 u5_mult_87_S2_4_23 ( .A(u5_mult_87_ab_4__23_), .B(
        u5_mult_87_CARRYB_3__23_), .CI(u5_mult_87_SUMB_3__24_), .CO(
        u5_mult_87_CARRYB_4__23_), .S(u5_mult_87_SUMB_4__23_) );
  FA_X1 u5_mult_87_S2_4_22 ( .A(u5_mult_87_ab_4__22_), .B(
        u5_mult_87_CARRYB_3__22_), .CI(u5_mult_87_SUMB_3__23_), .CO(
        u5_mult_87_CARRYB_4__22_), .S(u5_mult_87_SUMB_4__22_) );
  FA_X1 u5_mult_87_S2_4_21 ( .A(u5_mult_87_ab_4__21_), .B(
        u5_mult_87_CARRYB_3__21_), .CI(u5_mult_87_SUMB_3__22_), .CO(
        u5_mult_87_CARRYB_4__21_), .S(u5_mult_87_SUMB_4__21_) );
  FA_X1 u5_mult_87_S2_4_20 ( .A(u5_mult_87_ab_4__20_), .B(
        u5_mult_87_CARRYB_3__20_), .CI(u5_mult_87_SUMB_3__21_), .CO(
        u5_mult_87_CARRYB_4__20_), .S(u5_mult_87_SUMB_4__20_) );
  FA_X1 u5_mult_87_S2_4_19 ( .A(u5_mult_87_ab_4__19_), .B(
        u5_mult_87_CARRYB_3__19_), .CI(u5_mult_87_SUMB_3__20_), .CO(
        u5_mult_87_CARRYB_4__19_), .S(u5_mult_87_SUMB_4__19_) );
  FA_X1 u5_mult_87_S2_4_18 ( .A(u5_mult_87_ab_4__18_), .B(
        u5_mult_87_CARRYB_3__18_), .CI(u5_mult_87_SUMB_3__19_), .CO(
        u5_mult_87_CARRYB_4__18_), .S(u5_mult_87_SUMB_4__18_) );
  FA_X1 u5_mult_87_S2_4_17 ( .A(u5_mult_87_ab_4__17_), .B(
        u5_mult_87_CARRYB_3__17_), .CI(u5_mult_87_SUMB_3__18_), .CO(
        u5_mult_87_CARRYB_4__17_), .S(u5_mult_87_SUMB_4__17_) );
  FA_X1 u5_mult_87_S2_4_16 ( .A(u5_mult_87_ab_4__16_), .B(
        u5_mult_87_CARRYB_3__16_), .CI(u5_mult_87_SUMB_3__17_), .CO(
        u5_mult_87_CARRYB_4__16_), .S(u5_mult_87_SUMB_4__16_) );
  FA_X1 u5_mult_87_S2_4_15 ( .A(u5_mult_87_ab_4__15_), .B(
        u5_mult_87_CARRYB_3__15_), .CI(u5_mult_87_SUMB_3__16_), .CO(
        u5_mult_87_CARRYB_4__15_), .S(u5_mult_87_SUMB_4__15_) );
  FA_X1 u5_mult_87_S2_4_14 ( .A(u5_mult_87_ab_4__14_), .B(
        u5_mult_87_CARRYB_3__14_), .CI(u5_mult_87_SUMB_3__15_), .CO(
        u5_mult_87_CARRYB_4__14_), .S(u5_mult_87_SUMB_4__14_) );
  FA_X1 u5_mult_87_S2_4_13 ( .A(u5_mult_87_ab_4__13_), .B(
        u5_mult_87_CARRYB_3__13_), .CI(u5_mult_87_SUMB_3__14_), .CO(
        u5_mult_87_CARRYB_4__13_), .S(u5_mult_87_SUMB_4__13_) );
  FA_X1 u5_mult_87_S2_4_12 ( .A(u5_mult_87_ab_4__12_), .B(
        u5_mult_87_CARRYB_3__12_), .CI(u5_mult_87_SUMB_3__13_), .CO(
        u5_mult_87_CARRYB_4__12_), .S(u5_mult_87_SUMB_4__12_) );
  FA_X1 u5_mult_87_S2_4_11 ( .A(u5_mult_87_ab_4__11_), .B(
        u5_mult_87_CARRYB_3__11_), .CI(u5_mult_87_SUMB_3__12_), .CO(
        u5_mult_87_CARRYB_4__11_), .S(u5_mult_87_SUMB_4__11_) );
  FA_X1 u5_mult_87_S2_4_10 ( .A(u5_mult_87_ab_4__10_), .B(
        u5_mult_87_CARRYB_3__10_), .CI(u5_mult_87_SUMB_3__11_), .CO(
        u5_mult_87_CARRYB_4__10_), .S(u5_mult_87_SUMB_4__10_) );
  FA_X1 u5_mult_87_S2_4_9 ( .A(u5_mult_87_ab_4__9_), .B(
        u5_mult_87_CARRYB_3__9_), .CI(u5_mult_87_SUMB_3__10_), .CO(
        u5_mult_87_CARRYB_4__9_), .S(u5_mult_87_SUMB_4__9_) );
  FA_X1 u5_mult_87_S2_4_8 ( .A(u5_mult_87_ab_4__8_), .B(
        u5_mult_87_CARRYB_3__8_), .CI(u5_mult_87_SUMB_3__9_), .CO(
        u5_mult_87_CARRYB_4__8_), .S(u5_mult_87_SUMB_4__8_) );
  FA_X1 u5_mult_87_S2_4_7 ( .A(u5_mult_87_ab_4__7_), .B(
        u5_mult_87_CARRYB_3__7_), .CI(u5_mult_87_SUMB_3__8_), .CO(
        u5_mult_87_CARRYB_4__7_), .S(u5_mult_87_SUMB_4__7_) );
  FA_X1 u5_mult_87_S2_4_6 ( .A(u5_mult_87_ab_4__6_), .B(
        u5_mult_87_CARRYB_3__6_), .CI(u5_mult_87_SUMB_3__7_), .CO(
        u5_mult_87_CARRYB_4__6_), .S(u5_mult_87_SUMB_4__6_) );
  FA_X1 u5_mult_87_S2_4_5 ( .A(u5_mult_87_ab_4__5_), .B(
        u5_mult_87_CARRYB_3__5_), .CI(u5_mult_87_SUMB_3__6_), .CO(
        u5_mult_87_CARRYB_4__5_), .S(u5_mult_87_SUMB_4__5_) );
  FA_X1 u5_mult_87_S2_4_4 ( .A(u5_mult_87_ab_4__4_), .B(
        u5_mult_87_CARRYB_3__4_), .CI(u5_mult_87_SUMB_3__5_), .CO(
        u5_mult_87_CARRYB_4__4_), .S(u5_mult_87_SUMB_4__4_) );
  FA_X1 u5_mult_87_S2_4_3 ( .A(u5_mult_87_ab_4__3_), .B(
        u5_mult_87_CARRYB_3__3_), .CI(u5_mult_87_SUMB_3__4_), .CO(
        u5_mult_87_CARRYB_4__3_), .S(u5_mult_87_SUMB_4__3_) );
  FA_X1 u5_mult_87_S2_4_2 ( .A(u5_mult_87_ab_4__2_), .B(
        u5_mult_87_CARRYB_3__2_), .CI(u5_mult_87_SUMB_3__3_), .CO(
        u5_mult_87_CARRYB_4__2_), .S(u5_mult_87_SUMB_4__2_) );
  FA_X1 u5_mult_87_S2_4_1 ( .A(u5_mult_87_ab_4__1_), .B(
        u5_mult_87_CARRYB_3__1_), .CI(u5_mult_87_SUMB_3__2_), .CO(
        u5_mult_87_CARRYB_4__1_), .S(u5_mult_87_SUMB_4__1_) );
  FA_X1 u5_mult_87_S1_4_0 ( .A(u5_mult_87_ab_4__0_), .B(
        u5_mult_87_CARRYB_3__0_), .CI(u5_mult_87_SUMB_3__1_), .CO(
        u5_mult_87_CARRYB_4__0_), .S(u5_N4) );
  FA_X1 u5_mult_87_S3_5_51 ( .A(u5_mult_87_ab_5__51_), .B(
        u5_mult_87_CARRYB_4__51_), .CI(u5_mult_87_ab_4__52_), .CO(
        u5_mult_87_CARRYB_5__51_), .S(u5_mult_87_SUMB_5__51_) );
  FA_X1 u5_mult_87_S2_5_50 ( .A(u5_mult_87_ab_5__50_), .B(
        u5_mult_87_CARRYB_4__50_), .CI(u5_mult_87_SUMB_4__51_), .CO(
        u5_mult_87_CARRYB_5__50_), .S(u5_mult_87_SUMB_5__50_) );
  FA_X1 u5_mult_87_S2_5_49 ( .A(u5_mult_87_ab_5__49_), .B(
        u5_mult_87_CARRYB_4__49_), .CI(u5_mult_87_SUMB_4__50_), .CO(
        u5_mult_87_CARRYB_5__49_), .S(u5_mult_87_SUMB_5__49_) );
  FA_X1 u5_mult_87_S2_5_48 ( .A(u5_mult_87_ab_5__48_), .B(
        u5_mult_87_CARRYB_4__48_), .CI(u5_mult_87_SUMB_4__49_), .CO(
        u5_mult_87_CARRYB_5__48_), .S(u5_mult_87_SUMB_5__48_) );
  FA_X1 u5_mult_87_S2_5_47 ( .A(u5_mult_87_ab_5__47_), .B(
        u5_mult_87_CARRYB_4__47_), .CI(u5_mult_87_SUMB_4__48_), .CO(
        u5_mult_87_CARRYB_5__47_), .S(u5_mult_87_SUMB_5__47_) );
  FA_X1 u5_mult_87_S2_5_46 ( .A(u5_mult_87_ab_5__46_), .B(
        u5_mult_87_CARRYB_4__46_), .CI(u5_mult_87_SUMB_4__47_), .CO(
        u5_mult_87_CARRYB_5__46_), .S(u5_mult_87_SUMB_5__46_) );
  FA_X1 u5_mult_87_S2_5_45 ( .A(u5_mult_87_ab_5__45_), .B(
        u5_mult_87_CARRYB_4__45_), .CI(u5_mult_87_SUMB_4__46_), .CO(
        u5_mult_87_CARRYB_5__45_), .S(u5_mult_87_SUMB_5__45_) );
  FA_X1 u5_mult_87_S2_5_44 ( .A(u5_mult_87_ab_5__44_), .B(
        u5_mult_87_CARRYB_4__44_), .CI(u5_mult_87_SUMB_4__45_), .CO(
        u5_mult_87_CARRYB_5__44_), .S(u5_mult_87_SUMB_5__44_) );
  FA_X1 u5_mult_87_S2_5_43 ( .A(u5_mult_87_ab_5__43_), .B(
        u5_mult_87_CARRYB_4__43_), .CI(u5_mult_87_SUMB_4__44_), .CO(
        u5_mult_87_CARRYB_5__43_), .S(u5_mult_87_SUMB_5__43_) );
  FA_X1 u5_mult_87_S2_5_42 ( .A(u5_mult_87_ab_5__42_), .B(
        u5_mult_87_CARRYB_4__42_), .CI(u5_mult_87_SUMB_4__43_), .CO(
        u5_mult_87_CARRYB_5__42_), .S(u5_mult_87_SUMB_5__42_) );
  FA_X1 u5_mult_87_S2_5_41 ( .A(u5_mult_87_ab_5__41_), .B(
        u5_mult_87_CARRYB_4__41_), .CI(u5_mult_87_SUMB_4__42_), .CO(
        u5_mult_87_CARRYB_5__41_), .S(u5_mult_87_SUMB_5__41_) );
  FA_X1 u5_mult_87_S2_5_40 ( .A(u5_mult_87_ab_5__40_), .B(
        u5_mult_87_CARRYB_4__40_), .CI(u5_mult_87_SUMB_4__41_), .CO(
        u5_mult_87_CARRYB_5__40_), .S(u5_mult_87_SUMB_5__40_) );
  FA_X1 u5_mult_87_S2_5_39 ( .A(u5_mult_87_ab_5__39_), .B(
        u5_mult_87_CARRYB_4__39_), .CI(u5_mult_87_SUMB_4__40_), .CO(
        u5_mult_87_CARRYB_5__39_), .S(u5_mult_87_SUMB_5__39_) );
  FA_X1 u5_mult_87_S2_5_38 ( .A(u5_mult_87_ab_5__38_), .B(
        u5_mult_87_CARRYB_4__38_), .CI(u5_mult_87_SUMB_4__39_), .CO(
        u5_mult_87_CARRYB_5__38_), .S(u5_mult_87_SUMB_5__38_) );
  FA_X1 u5_mult_87_S2_5_37 ( .A(u5_mult_87_ab_5__37_), .B(
        u5_mult_87_CARRYB_4__37_), .CI(u5_mult_87_SUMB_4__38_), .CO(
        u5_mult_87_CARRYB_5__37_), .S(u5_mult_87_SUMB_5__37_) );
  FA_X1 u5_mult_87_S2_5_36 ( .A(u5_mult_87_ab_5__36_), .B(
        u5_mult_87_CARRYB_4__36_), .CI(u5_mult_87_SUMB_4__37_), .CO(
        u5_mult_87_CARRYB_5__36_), .S(u5_mult_87_SUMB_5__36_) );
  FA_X1 u5_mult_87_S2_5_35 ( .A(u5_mult_87_ab_5__35_), .B(
        u5_mult_87_CARRYB_4__35_), .CI(u5_mult_87_SUMB_4__36_), .CO(
        u5_mult_87_CARRYB_5__35_), .S(u5_mult_87_SUMB_5__35_) );
  FA_X1 u5_mult_87_S2_5_34 ( .A(u5_mult_87_ab_5__34_), .B(
        u5_mult_87_CARRYB_4__34_), .CI(u5_mult_87_SUMB_4__35_), .CO(
        u5_mult_87_CARRYB_5__34_), .S(u5_mult_87_SUMB_5__34_) );
  FA_X1 u5_mult_87_S2_5_33 ( .A(u5_mult_87_ab_5__33_), .B(
        u5_mult_87_CARRYB_4__33_), .CI(u5_mult_87_SUMB_4__34_), .CO(
        u5_mult_87_CARRYB_5__33_), .S(u5_mult_87_SUMB_5__33_) );
  FA_X1 u5_mult_87_S2_5_32 ( .A(u5_mult_87_ab_5__32_), .B(
        u5_mult_87_CARRYB_4__32_), .CI(u5_mult_87_SUMB_4__33_), .CO(
        u5_mult_87_CARRYB_5__32_), .S(u5_mult_87_SUMB_5__32_) );
  FA_X1 u5_mult_87_S2_5_31 ( .A(u5_mult_87_ab_5__31_), .B(
        u5_mult_87_CARRYB_4__31_), .CI(u5_mult_87_SUMB_4__32_), .CO(
        u5_mult_87_CARRYB_5__31_), .S(u5_mult_87_SUMB_5__31_) );
  FA_X1 u5_mult_87_S2_5_30 ( .A(u5_mult_87_ab_5__30_), .B(
        u5_mult_87_CARRYB_4__30_), .CI(u5_mult_87_SUMB_4__31_), .CO(
        u5_mult_87_CARRYB_5__30_), .S(u5_mult_87_SUMB_5__30_) );
  FA_X1 u5_mult_87_S2_5_29 ( .A(u5_mult_87_ab_5__29_), .B(
        u5_mult_87_CARRYB_4__29_), .CI(u5_mult_87_SUMB_4__30_), .CO(
        u5_mult_87_CARRYB_5__29_), .S(u5_mult_87_SUMB_5__29_) );
  FA_X1 u5_mult_87_S2_5_28 ( .A(u5_mult_87_ab_5__28_), .B(
        u5_mult_87_CARRYB_4__28_), .CI(u5_mult_87_SUMB_4__29_), .CO(
        u5_mult_87_CARRYB_5__28_), .S(u5_mult_87_SUMB_5__28_) );
  FA_X1 u5_mult_87_S2_5_27 ( .A(u5_mult_87_ab_5__27_), .B(
        u5_mult_87_CARRYB_4__27_), .CI(u5_mult_87_SUMB_4__28_), .CO(
        u5_mult_87_CARRYB_5__27_), .S(u5_mult_87_SUMB_5__27_) );
  FA_X1 u5_mult_87_S2_5_26 ( .A(u5_mult_87_ab_5__26_), .B(
        u5_mult_87_CARRYB_4__26_), .CI(u5_mult_87_SUMB_4__27_), .CO(
        u5_mult_87_CARRYB_5__26_), .S(u5_mult_87_SUMB_5__26_) );
  FA_X1 u5_mult_87_S2_5_25 ( .A(u5_mult_87_ab_5__25_), .B(
        u5_mult_87_CARRYB_4__25_), .CI(u5_mult_87_SUMB_4__26_), .CO(
        u5_mult_87_CARRYB_5__25_), .S(u5_mult_87_SUMB_5__25_) );
  FA_X1 u5_mult_87_S2_5_24 ( .A(u5_mult_87_ab_5__24_), .B(
        u5_mult_87_CARRYB_4__24_), .CI(u5_mult_87_SUMB_4__25_), .CO(
        u5_mult_87_CARRYB_5__24_), .S(u5_mult_87_SUMB_5__24_) );
  FA_X1 u5_mult_87_S2_5_23 ( .A(u5_mult_87_ab_5__23_), .B(
        u5_mult_87_CARRYB_4__23_), .CI(u5_mult_87_SUMB_4__24_), .CO(
        u5_mult_87_CARRYB_5__23_), .S(u5_mult_87_SUMB_5__23_) );
  FA_X1 u5_mult_87_S2_5_22 ( .A(u5_mult_87_ab_5__22_), .B(
        u5_mult_87_CARRYB_4__22_), .CI(u5_mult_87_SUMB_4__23_), .CO(
        u5_mult_87_CARRYB_5__22_), .S(u5_mult_87_SUMB_5__22_) );
  FA_X1 u5_mult_87_S2_5_21 ( .A(u5_mult_87_ab_5__21_), .B(
        u5_mult_87_CARRYB_4__21_), .CI(u5_mult_87_SUMB_4__22_), .CO(
        u5_mult_87_CARRYB_5__21_), .S(u5_mult_87_SUMB_5__21_) );
  FA_X1 u5_mult_87_S2_5_20 ( .A(u5_mult_87_ab_5__20_), .B(
        u5_mult_87_CARRYB_4__20_), .CI(u5_mult_87_SUMB_4__21_), .CO(
        u5_mult_87_CARRYB_5__20_), .S(u5_mult_87_SUMB_5__20_) );
  FA_X1 u5_mult_87_S2_5_19 ( .A(u5_mult_87_ab_5__19_), .B(
        u5_mult_87_CARRYB_4__19_), .CI(u5_mult_87_SUMB_4__20_), .CO(
        u5_mult_87_CARRYB_5__19_), .S(u5_mult_87_SUMB_5__19_) );
  FA_X1 u5_mult_87_S2_5_18 ( .A(u5_mult_87_ab_5__18_), .B(
        u5_mult_87_CARRYB_4__18_), .CI(u5_mult_87_SUMB_4__19_), .CO(
        u5_mult_87_CARRYB_5__18_), .S(u5_mult_87_SUMB_5__18_) );
  FA_X1 u5_mult_87_S2_5_17 ( .A(u5_mult_87_ab_5__17_), .B(
        u5_mult_87_CARRYB_4__17_), .CI(u5_mult_87_SUMB_4__18_), .CO(
        u5_mult_87_CARRYB_5__17_), .S(u5_mult_87_SUMB_5__17_) );
  FA_X1 u5_mult_87_S2_5_16 ( .A(u5_mult_87_ab_5__16_), .B(
        u5_mult_87_CARRYB_4__16_), .CI(u5_mult_87_SUMB_4__17_), .CO(
        u5_mult_87_CARRYB_5__16_), .S(u5_mult_87_SUMB_5__16_) );
  FA_X1 u5_mult_87_S2_5_15 ( .A(u5_mult_87_ab_5__15_), .B(
        u5_mult_87_CARRYB_4__15_), .CI(u5_mult_87_SUMB_4__16_), .CO(
        u5_mult_87_CARRYB_5__15_), .S(u5_mult_87_SUMB_5__15_) );
  FA_X1 u5_mult_87_S2_5_14 ( .A(u5_mult_87_ab_5__14_), .B(
        u5_mult_87_CARRYB_4__14_), .CI(u5_mult_87_SUMB_4__15_), .CO(
        u5_mult_87_CARRYB_5__14_), .S(u5_mult_87_SUMB_5__14_) );
  FA_X1 u5_mult_87_S2_5_13 ( .A(u5_mult_87_ab_5__13_), .B(
        u5_mult_87_CARRYB_4__13_), .CI(u5_mult_87_SUMB_4__14_), .CO(
        u5_mult_87_CARRYB_5__13_), .S(u5_mult_87_SUMB_5__13_) );
  FA_X1 u5_mult_87_S2_5_12 ( .A(u5_mult_87_ab_5__12_), .B(
        u5_mult_87_CARRYB_4__12_), .CI(u5_mult_87_SUMB_4__13_), .CO(
        u5_mult_87_CARRYB_5__12_), .S(u5_mult_87_SUMB_5__12_) );
  FA_X1 u5_mult_87_S2_5_11 ( .A(u5_mult_87_ab_5__11_), .B(
        u5_mult_87_CARRYB_4__11_), .CI(u5_mult_87_SUMB_4__12_), .CO(
        u5_mult_87_CARRYB_5__11_), .S(u5_mult_87_SUMB_5__11_) );
  FA_X1 u5_mult_87_S2_5_10 ( .A(u5_mult_87_ab_5__10_), .B(
        u5_mult_87_CARRYB_4__10_), .CI(u5_mult_87_SUMB_4__11_), .CO(
        u5_mult_87_CARRYB_5__10_), .S(u5_mult_87_SUMB_5__10_) );
  FA_X1 u5_mult_87_S2_5_9 ( .A(u5_mult_87_ab_5__9_), .B(
        u5_mult_87_CARRYB_4__9_), .CI(u5_mult_87_SUMB_4__10_), .CO(
        u5_mult_87_CARRYB_5__9_), .S(u5_mult_87_SUMB_5__9_) );
  FA_X1 u5_mult_87_S2_5_8 ( .A(u5_mult_87_ab_5__8_), .B(
        u5_mult_87_CARRYB_4__8_), .CI(u5_mult_87_SUMB_4__9_), .CO(
        u5_mult_87_CARRYB_5__8_), .S(u5_mult_87_SUMB_5__8_) );
  FA_X1 u5_mult_87_S2_5_7 ( .A(u5_mult_87_ab_5__7_), .B(
        u5_mult_87_CARRYB_4__7_), .CI(u5_mult_87_SUMB_4__8_), .CO(
        u5_mult_87_CARRYB_5__7_), .S(u5_mult_87_SUMB_5__7_) );
  FA_X1 u5_mult_87_S2_5_6 ( .A(u5_mult_87_ab_5__6_), .B(
        u5_mult_87_CARRYB_4__6_), .CI(u5_mult_87_SUMB_4__7_), .CO(
        u5_mult_87_CARRYB_5__6_), .S(u5_mult_87_SUMB_5__6_) );
  FA_X1 u5_mult_87_S2_5_5 ( .A(u5_mult_87_ab_5__5_), .B(
        u5_mult_87_CARRYB_4__5_), .CI(u5_mult_87_SUMB_4__6_), .CO(
        u5_mult_87_CARRYB_5__5_), .S(u5_mult_87_SUMB_5__5_) );
  FA_X1 u5_mult_87_S2_5_4 ( .A(u5_mult_87_ab_5__4_), .B(
        u5_mult_87_CARRYB_4__4_), .CI(u5_mult_87_SUMB_4__5_), .CO(
        u5_mult_87_CARRYB_5__4_), .S(u5_mult_87_SUMB_5__4_) );
  FA_X1 u5_mult_87_S2_5_3 ( .A(u5_mult_87_ab_5__3_), .B(
        u5_mult_87_CARRYB_4__3_), .CI(u5_mult_87_SUMB_4__4_), .CO(
        u5_mult_87_CARRYB_5__3_), .S(u5_mult_87_SUMB_5__3_) );
  FA_X1 u5_mult_87_S2_5_2 ( .A(u5_mult_87_ab_5__2_), .B(
        u5_mult_87_CARRYB_4__2_), .CI(u5_mult_87_SUMB_4__3_), .CO(
        u5_mult_87_CARRYB_5__2_), .S(u5_mult_87_SUMB_5__2_) );
  FA_X1 u5_mult_87_S2_5_1 ( .A(u5_mult_87_ab_5__1_), .B(
        u5_mult_87_CARRYB_4__1_), .CI(u5_mult_87_SUMB_4__2_), .CO(
        u5_mult_87_CARRYB_5__1_), .S(u5_mult_87_SUMB_5__1_) );
  FA_X1 u5_mult_87_S1_5_0 ( .A(u5_mult_87_ab_5__0_), .B(
        u5_mult_87_CARRYB_4__0_), .CI(u5_mult_87_SUMB_4__1_), .CO(
        u5_mult_87_CARRYB_5__0_), .S(u5_N5) );
  FA_X1 u5_mult_87_S3_6_51 ( .A(u5_mult_87_ab_6__51_), .B(
        u5_mult_87_CARRYB_5__51_), .CI(u5_mult_87_ab_5__52_), .CO(
        u5_mult_87_CARRYB_6__51_), .S(u5_mult_87_SUMB_6__51_) );
  FA_X1 u5_mult_87_S2_6_50 ( .A(u5_mult_87_ab_6__50_), .B(
        u5_mult_87_CARRYB_5__50_), .CI(u5_mult_87_SUMB_5__51_), .CO(
        u5_mult_87_CARRYB_6__50_), .S(u5_mult_87_SUMB_6__50_) );
  FA_X1 u5_mult_87_S2_6_49 ( .A(u5_mult_87_ab_6__49_), .B(
        u5_mult_87_CARRYB_5__49_), .CI(u5_mult_87_SUMB_5__50_), .CO(
        u5_mult_87_CARRYB_6__49_), .S(u5_mult_87_SUMB_6__49_) );
  FA_X1 u5_mult_87_S2_6_48 ( .A(u5_mult_87_ab_6__48_), .B(
        u5_mult_87_CARRYB_5__48_), .CI(u5_mult_87_SUMB_5__49_), .CO(
        u5_mult_87_CARRYB_6__48_), .S(u5_mult_87_SUMB_6__48_) );
  FA_X1 u5_mult_87_S2_6_47 ( .A(u5_mult_87_ab_6__47_), .B(
        u5_mult_87_CARRYB_5__47_), .CI(u5_mult_87_SUMB_5__48_), .CO(
        u5_mult_87_CARRYB_6__47_), .S(u5_mult_87_SUMB_6__47_) );
  FA_X1 u5_mult_87_S2_6_46 ( .A(u5_mult_87_ab_6__46_), .B(
        u5_mult_87_CARRYB_5__46_), .CI(u5_mult_87_SUMB_5__47_), .CO(
        u5_mult_87_CARRYB_6__46_), .S(u5_mult_87_SUMB_6__46_) );
  FA_X1 u5_mult_87_S2_6_45 ( .A(u5_mult_87_ab_6__45_), .B(
        u5_mult_87_CARRYB_5__45_), .CI(u5_mult_87_SUMB_5__46_), .CO(
        u5_mult_87_CARRYB_6__45_), .S(u5_mult_87_SUMB_6__45_) );
  FA_X1 u5_mult_87_S2_6_44 ( .A(u5_mult_87_ab_6__44_), .B(
        u5_mult_87_CARRYB_5__44_), .CI(u5_mult_87_SUMB_5__45_), .CO(
        u5_mult_87_CARRYB_6__44_), .S(u5_mult_87_SUMB_6__44_) );
  FA_X1 u5_mult_87_S2_6_43 ( .A(u5_mult_87_ab_6__43_), .B(
        u5_mult_87_CARRYB_5__43_), .CI(u5_mult_87_SUMB_5__44_), .CO(
        u5_mult_87_CARRYB_6__43_), .S(u5_mult_87_SUMB_6__43_) );
  FA_X1 u5_mult_87_S2_6_42 ( .A(u5_mult_87_ab_6__42_), .B(
        u5_mult_87_CARRYB_5__42_), .CI(u5_mult_87_SUMB_5__43_), .CO(
        u5_mult_87_CARRYB_6__42_), .S(u5_mult_87_SUMB_6__42_) );
  FA_X1 u5_mult_87_S2_6_41 ( .A(u5_mult_87_ab_6__41_), .B(
        u5_mult_87_CARRYB_5__41_), .CI(u5_mult_87_SUMB_5__42_), .CO(
        u5_mult_87_CARRYB_6__41_), .S(u5_mult_87_SUMB_6__41_) );
  FA_X1 u5_mult_87_S2_6_40 ( .A(u5_mult_87_ab_6__40_), .B(
        u5_mult_87_CARRYB_5__40_), .CI(u5_mult_87_SUMB_5__41_), .CO(
        u5_mult_87_CARRYB_6__40_), .S(u5_mult_87_SUMB_6__40_) );
  FA_X1 u5_mult_87_S2_6_39 ( .A(u5_mult_87_ab_6__39_), .B(
        u5_mult_87_CARRYB_5__39_), .CI(u5_mult_87_SUMB_5__40_), .CO(
        u5_mult_87_CARRYB_6__39_), .S(u5_mult_87_SUMB_6__39_) );
  FA_X1 u5_mult_87_S2_6_38 ( .A(u5_mult_87_ab_6__38_), .B(
        u5_mult_87_CARRYB_5__38_), .CI(u5_mult_87_SUMB_5__39_), .CO(
        u5_mult_87_CARRYB_6__38_), .S(u5_mult_87_SUMB_6__38_) );
  FA_X1 u5_mult_87_S2_6_37 ( .A(u5_mult_87_ab_6__37_), .B(
        u5_mult_87_CARRYB_5__37_), .CI(u5_mult_87_SUMB_5__38_), .CO(
        u5_mult_87_CARRYB_6__37_), .S(u5_mult_87_SUMB_6__37_) );
  FA_X1 u5_mult_87_S2_6_36 ( .A(u5_mult_87_ab_6__36_), .B(
        u5_mult_87_CARRYB_5__36_), .CI(u5_mult_87_SUMB_5__37_), .CO(
        u5_mult_87_CARRYB_6__36_), .S(u5_mult_87_SUMB_6__36_) );
  FA_X1 u5_mult_87_S2_6_35 ( .A(u5_mult_87_ab_6__35_), .B(
        u5_mult_87_CARRYB_5__35_), .CI(u5_mult_87_SUMB_5__36_), .CO(
        u5_mult_87_CARRYB_6__35_), .S(u5_mult_87_SUMB_6__35_) );
  FA_X1 u5_mult_87_S2_6_34 ( .A(u5_mult_87_ab_6__34_), .B(
        u5_mult_87_CARRYB_5__34_), .CI(u5_mult_87_SUMB_5__35_), .CO(
        u5_mult_87_CARRYB_6__34_), .S(u5_mult_87_SUMB_6__34_) );
  FA_X1 u5_mult_87_S2_6_33 ( .A(u5_mult_87_ab_6__33_), .B(
        u5_mult_87_CARRYB_5__33_), .CI(u5_mult_87_SUMB_5__34_), .CO(
        u5_mult_87_CARRYB_6__33_), .S(u5_mult_87_SUMB_6__33_) );
  FA_X1 u5_mult_87_S2_6_32 ( .A(u5_mult_87_ab_6__32_), .B(
        u5_mult_87_CARRYB_5__32_), .CI(u5_mult_87_SUMB_5__33_), .CO(
        u5_mult_87_CARRYB_6__32_), .S(u5_mult_87_SUMB_6__32_) );
  FA_X1 u5_mult_87_S2_6_31 ( .A(u5_mult_87_ab_6__31_), .B(
        u5_mult_87_CARRYB_5__31_), .CI(u5_mult_87_SUMB_5__32_), .CO(
        u5_mult_87_CARRYB_6__31_), .S(u5_mult_87_SUMB_6__31_) );
  FA_X1 u5_mult_87_S2_6_30 ( .A(u5_mult_87_ab_6__30_), .B(
        u5_mult_87_CARRYB_5__30_), .CI(u5_mult_87_SUMB_5__31_), .CO(
        u5_mult_87_CARRYB_6__30_), .S(u5_mult_87_SUMB_6__30_) );
  FA_X1 u5_mult_87_S2_6_29 ( .A(u5_mult_87_ab_6__29_), .B(
        u5_mult_87_CARRYB_5__29_), .CI(u5_mult_87_SUMB_5__30_), .CO(
        u5_mult_87_CARRYB_6__29_), .S(u5_mult_87_SUMB_6__29_) );
  FA_X1 u5_mult_87_S2_6_28 ( .A(u5_mult_87_ab_6__28_), .B(
        u5_mult_87_CARRYB_5__28_), .CI(u5_mult_87_SUMB_5__29_), .CO(
        u5_mult_87_CARRYB_6__28_), .S(u5_mult_87_SUMB_6__28_) );
  FA_X1 u5_mult_87_S2_6_27 ( .A(u5_mult_87_ab_6__27_), .B(
        u5_mult_87_CARRYB_5__27_), .CI(u5_mult_87_SUMB_5__28_), .CO(
        u5_mult_87_CARRYB_6__27_), .S(u5_mult_87_SUMB_6__27_) );
  FA_X1 u5_mult_87_S2_6_26 ( .A(u5_mult_87_ab_6__26_), .B(
        u5_mult_87_CARRYB_5__26_), .CI(u5_mult_87_SUMB_5__27_), .CO(
        u5_mult_87_CARRYB_6__26_), .S(u5_mult_87_SUMB_6__26_) );
  FA_X1 u5_mult_87_S2_6_25 ( .A(u5_mult_87_ab_6__25_), .B(
        u5_mult_87_CARRYB_5__25_), .CI(u5_mult_87_SUMB_5__26_), .CO(
        u5_mult_87_CARRYB_6__25_), .S(u5_mult_87_SUMB_6__25_) );
  FA_X1 u5_mult_87_S2_6_24 ( .A(u5_mult_87_ab_6__24_), .B(
        u5_mult_87_CARRYB_5__24_), .CI(u5_mult_87_SUMB_5__25_), .CO(
        u5_mult_87_CARRYB_6__24_), .S(u5_mult_87_SUMB_6__24_) );
  FA_X1 u5_mult_87_S2_6_23 ( .A(u5_mult_87_ab_6__23_), .B(
        u5_mult_87_CARRYB_5__23_), .CI(u5_mult_87_SUMB_5__24_), .CO(
        u5_mult_87_CARRYB_6__23_), .S(u5_mult_87_SUMB_6__23_) );
  FA_X1 u5_mult_87_S2_6_22 ( .A(u5_mult_87_ab_6__22_), .B(
        u5_mult_87_CARRYB_5__22_), .CI(u5_mult_87_SUMB_5__23_), .CO(
        u5_mult_87_CARRYB_6__22_), .S(u5_mult_87_SUMB_6__22_) );
  FA_X1 u5_mult_87_S2_6_21 ( .A(u5_mult_87_ab_6__21_), .B(
        u5_mult_87_CARRYB_5__21_), .CI(u5_mult_87_SUMB_5__22_), .CO(
        u5_mult_87_CARRYB_6__21_), .S(u5_mult_87_SUMB_6__21_) );
  FA_X1 u5_mult_87_S2_6_20 ( .A(u5_mult_87_ab_6__20_), .B(
        u5_mult_87_CARRYB_5__20_), .CI(u5_mult_87_SUMB_5__21_), .CO(
        u5_mult_87_CARRYB_6__20_), .S(u5_mult_87_SUMB_6__20_) );
  FA_X1 u5_mult_87_S2_6_19 ( .A(u5_mult_87_ab_6__19_), .B(
        u5_mult_87_CARRYB_5__19_), .CI(u5_mult_87_SUMB_5__20_), .CO(
        u5_mult_87_CARRYB_6__19_), .S(u5_mult_87_SUMB_6__19_) );
  FA_X1 u5_mult_87_S2_6_18 ( .A(u5_mult_87_ab_6__18_), .B(
        u5_mult_87_CARRYB_5__18_), .CI(u5_mult_87_SUMB_5__19_), .CO(
        u5_mult_87_CARRYB_6__18_), .S(u5_mult_87_SUMB_6__18_) );
  FA_X1 u5_mult_87_S2_6_17 ( .A(u5_mult_87_ab_6__17_), .B(
        u5_mult_87_CARRYB_5__17_), .CI(u5_mult_87_SUMB_5__18_), .CO(
        u5_mult_87_CARRYB_6__17_), .S(u5_mult_87_SUMB_6__17_) );
  FA_X1 u5_mult_87_S2_6_16 ( .A(u5_mult_87_ab_6__16_), .B(
        u5_mult_87_CARRYB_5__16_), .CI(u5_mult_87_SUMB_5__17_), .CO(
        u5_mult_87_CARRYB_6__16_), .S(u5_mult_87_SUMB_6__16_) );
  FA_X1 u5_mult_87_S2_6_15 ( .A(u5_mult_87_ab_6__15_), .B(
        u5_mult_87_CARRYB_5__15_), .CI(u5_mult_87_SUMB_5__16_), .CO(
        u5_mult_87_CARRYB_6__15_), .S(u5_mult_87_SUMB_6__15_) );
  FA_X1 u5_mult_87_S2_6_14 ( .A(u5_mult_87_ab_6__14_), .B(
        u5_mult_87_CARRYB_5__14_), .CI(u5_mult_87_SUMB_5__15_), .CO(
        u5_mult_87_CARRYB_6__14_), .S(u5_mult_87_SUMB_6__14_) );
  FA_X1 u5_mult_87_S2_6_13 ( .A(u5_mult_87_ab_6__13_), .B(
        u5_mult_87_CARRYB_5__13_), .CI(u5_mult_87_SUMB_5__14_), .CO(
        u5_mult_87_CARRYB_6__13_), .S(u5_mult_87_SUMB_6__13_) );
  FA_X1 u5_mult_87_S2_6_12 ( .A(u5_mult_87_ab_6__12_), .B(
        u5_mult_87_CARRYB_5__12_), .CI(u5_mult_87_SUMB_5__13_), .CO(
        u5_mult_87_CARRYB_6__12_), .S(u5_mult_87_SUMB_6__12_) );
  FA_X1 u5_mult_87_S2_6_11 ( .A(u5_mult_87_ab_6__11_), .B(
        u5_mult_87_CARRYB_5__11_), .CI(u5_mult_87_SUMB_5__12_), .CO(
        u5_mult_87_CARRYB_6__11_), .S(u5_mult_87_SUMB_6__11_) );
  FA_X1 u5_mult_87_S2_6_10 ( .A(u5_mult_87_ab_6__10_), .B(
        u5_mult_87_CARRYB_5__10_), .CI(u5_mult_87_SUMB_5__11_), .CO(
        u5_mult_87_CARRYB_6__10_), .S(u5_mult_87_SUMB_6__10_) );
  FA_X1 u5_mult_87_S2_6_9 ( .A(u5_mult_87_ab_6__9_), .B(
        u5_mult_87_CARRYB_5__9_), .CI(u5_mult_87_SUMB_5__10_), .CO(
        u5_mult_87_CARRYB_6__9_), .S(u5_mult_87_SUMB_6__9_) );
  FA_X1 u5_mult_87_S2_6_8 ( .A(u5_mult_87_ab_6__8_), .B(
        u5_mult_87_CARRYB_5__8_), .CI(u5_mult_87_SUMB_5__9_), .CO(
        u5_mult_87_CARRYB_6__8_), .S(u5_mult_87_SUMB_6__8_) );
  FA_X1 u5_mult_87_S2_6_7 ( .A(u5_mult_87_ab_6__7_), .B(
        u5_mult_87_CARRYB_5__7_), .CI(u5_mult_87_SUMB_5__8_), .CO(
        u5_mult_87_CARRYB_6__7_), .S(u5_mult_87_SUMB_6__7_) );
  FA_X1 u5_mult_87_S2_6_6 ( .A(u5_mult_87_ab_6__6_), .B(
        u5_mult_87_CARRYB_5__6_), .CI(u5_mult_87_SUMB_5__7_), .CO(
        u5_mult_87_CARRYB_6__6_), .S(u5_mult_87_SUMB_6__6_) );
  FA_X1 u5_mult_87_S2_6_5 ( .A(u5_mult_87_ab_6__5_), .B(
        u5_mult_87_CARRYB_5__5_), .CI(u5_mult_87_SUMB_5__6_), .CO(
        u5_mult_87_CARRYB_6__5_), .S(u5_mult_87_SUMB_6__5_) );
  FA_X1 u5_mult_87_S2_6_4 ( .A(u5_mult_87_ab_6__4_), .B(
        u5_mult_87_CARRYB_5__4_), .CI(u5_mult_87_SUMB_5__5_), .CO(
        u5_mult_87_CARRYB_6__4_), .S(u5_mult_87_SUMB_6__4_) );
  FA_X1 u5_mult_87_S2_6_3 ( .A(u5_mult_87_ab_6__3_), .B(
        u5_mult_87_CARRYB_5__3_), .CI(u5_mult_87_SUMB_5__4_), .CO(
        u5_mult_87_CARRYB_6__3_), .S(u5_mult_87_SUMB_6__3_) );
  FA_X1 u5_mult_87_S2_6_2 ( .A(u5_mult_87_ab_6__2_), .B(
        u5_mult_87_CARRYB_5__2_), .CI(u5_mult_87_SUMB_5__3_), .CO(
        u5_mult_87_CARRYB_6__2_), .S(u5_mult_87_SUMB_6__2_) );
  FA_X1 u5_mult_87_S2_6_1 ( .A(u5_mult_87_ab_6__1_), .B(
        u5_mult_87_CARRYB_5__1_), .CI(u5_mult_87_SUMB_5__2_), .CO(
        u5_mult_87_CARRYB_6__1_), .S(u5_mult_87_SUMB_6__1_) );
  FA_X1 u5_mult_87_S1_6_0 ( .A(u5_mult_87_ab_6__0_), .B(
        u5_mult_87_CARRYB_5__0_), .CI(u5_mult_87_SUMB_5__1_), .CO(
        u5_mult_87_CARRYB_6__0_), .S(u5_N6) );
  FA_X1 u5_mult_87_S3_7_51 ( .A(u5_mult_87_ab_7__51_), .B(
        u5_mult_87_CARRYB_6__51_), .CI(u5_mult_87_ab_6__52_), .CO(
        u5_mult_87_CARRYB_7__51_), .S(u5_mult_87_SUMB_7__51_) );
  FA_X1 u5_mult_87_S2_7_50 ( .A(u5_mult_87_ab_7__50_), .B(
        u5_mult_87_CARRYB_6__50_), .CI(u5_mult_87_SUMB_6__51_), .CO(
        u5_mult_87_CARRYB_7__50_), .S(u5_mult_87_SUMB_7__50_) );
  FA_X1 u5_mult_87_S2_7_49 ( .A(u5_mult_87_ab_7__49_), .B(
        u5_mult_87_CARRYB_6__49_), .CI(u5_mult_87_SUMB_6__50_), .CO(
        u5_mult_87_CARRYB_7__49_), .S(u5_mult_87_SUMB_7__49_) );
  FA_X1 u5_mult_87_S2_7_48 ( .A(u5_mult_87_ab_7__48_), .B(
        u5_mult_87_CARRYB_6__48_), .CI(u5_mult_87_SUMB_6__49_), .CO(
        u5_mult_87_CARRYB_7__48_), .S(u5_mult_87_SUMB_7__48_) );
  FA_X1 u5_mult_87_S2_7_47 ( .A(u5_mult_87_ab_7__47_), .B(
        u5_mult_87_CARRYB_6__47_), .CI(u5_mult_87_SUMB_6__48_), .CO(
        u5_mult_87_CARRYB_7__47_), .S(u5_mult_87_SUMB_7__47_) );
  FA_X1 u5_mult_87_S2_7_46 ( .A(u5_mult_87_ab_7__46_), .B(
        u5_mult_87_CARRYB_6__46_), .CI(u5_mult_87_SUMB_6__47_), .CO(
        u5_mult_87_CARRYB_7__46_), .S(u5_mult_87_SUMB_7__46_) );
  FA_X1 u5_mult_87_S2_7_45 ( .A(u5_mult_87_ab_7__45_), .B(
        u5_mult_87_CARRYB_6__45_), .CI(u5_mult_87_SUMB_6__46_), .CO(
        u5_mult_87_CARRYB_7__45_), .S(u5_mult_87_SUMB_7__45_) );
  FA_X1 u5_mult_87_S2_7_44 ( .A(u5_mult_87_ab_7__44_), .B(
        u5_mult_87_CARRYB_6__44_), .CI(u5_mult_87_SUMB_6__45_), .CO(
        u5_mult_87_CARRYB_7__44_), .S(u5_mult_87_SUMB_7__44_) );
  FA_X1 u5_mult_87_S2_7_43 ( .A(u5_mult_87_ab_7__43_), .B(
        u5_mult_87_CARRYB_6__43_), .CI(u5_mult_87_SUMB_6__44_), .CO(
        u5_mult_87_CARRYB_7__43_), .S(u5_mult_87_SUMB_7__43_) );
  FA_X1 u5_mult_87_S2_7_42 ( .A(u5_mult_87_ab_7__42_), .B(
        u5_mult_87_CARRYB_6__42_), .CI(u5_mult_87_SUMB_6__43_), .CO(
        u5_mult_87_CARRYB_7__42_), .S(u5_mult_87_SUMB_7__42_) );
  FA_X1 u5_mult_87_S2_7_41 ( .A(u5_mult_87_ab_7__41_), .B(
        u5_mult_87_CARRYB_6__41_), .CI(u5_mult_87_SUMB_6__42_), .CO(
        u5_mult_87_CARRYB_7__41_), .S(u5_mult_87_SUMB_7__41_) );
  FA_X1 u5_mult_87_S2_7_40 ( .A(u5_mult_87_ab_7__40_), .B(
        u5_mult_87_CARRYB_6__40_), .CI(u5_mult_87_SUMB_6__41_), .CO(
        u5_mult_87_CARRYB_7__40_), .S(u5_mult_87_SUMB_7__40_) );
  FA_X1 u5_mult_87_S2_7_39 ( .A(u5_mult_87_ab_7__39_), .B(
        u5_mult_87_CARRYB_6__39_), .CI(u5_mult_87_SUMB_6__40_), .CO(
        u5_mult_87_CARRYB_7__39_), .S(u5_mult_87_SUMB_7__39_) );
  FA_X1 u5_mult_87_S2_7_38 ( .A(u5_mult_87_ab_7__38_), .B(
        u5_mult_87_CARRYB_6__38_), .CI(u5_mult_87_SUMB_6__39_), .CO(
        u5_mult_87_CARRYB_7__38_), .S(u5_mult_87_SUMB_7__38_) );
  FA_X1 u5_mult_87_S2_7_37 ( .A(u5_mult_87_ab_7__37_), .B(
        u5_mult_87_CARRYB_6__37_), .CI(u5_mult_87_SUMB_6__38_), .CO(
        u5_mult_87_CARRYB_7__37_), .S(u5_mult_87_SUMB_7__37_) );
  FA_X1 u5_mult_87_S2_7_36 ( .A(u5_mult_87_ab_7__36_), .B(
        u5_mult_87_CARRYB_6__36_), .CI(u5_mult_87_SUMB_6__37_), .CO(
        u5_mult_87_CARRYB_7__36_), .S(u5_mult_87_SUMB_7__36_) );
  FA_X1 u5_mult_87_S2_7_35 ( .A(u5_mult_87_ab_7__35_), .B(
        u5_mult_87_CARRYB_6__35_), .CI(u5_mult_87_SUMB_6__36_), .CO(
        u5_mult_87_CARRYB_7__35_), .S(u5_mult_87_SUMB_7__35_) );
  FA_X1 u5_mult_87_S2_7_34 ( .A(u5_mult_87_ab_7__34_), .B(
        u5_mult_87_CARRYB_6__34_), .CI(u5_mult_87_SUMB_6__35_), .CO(
        u5_mult_87_CARRYB_7__34_), .S(u5_mult_87_SUMB_7__34_) );
  FA_X1 u5_mult_87_S2_7_33 ( .A(u5_mult_87_ab_7__33_), .B(
        u5_mult_87_CARRYB_6__33_), .CI(u5_mult_87_SUMB_6__34_), .CO(
        u5_mult_87_CARRYB_7__33_), .S(u5_mult_87_SUMB_7__33_) );
  FA_X1 u5_mult_87_S2_7_32 ( .A(u5_mult_87_ab_7__32_), .B(
        u5_mult_87_CARRYB_6__32_), .CI(u5_mult_87_SUMB_6__33_), .CO(
        u5_mult_87_CARRYB_7__32_), .S(u5_mult_87_SUMB_7__32_) );
  FA_X1 u5_mult_87_S2_7_31 ( .A(u5_mult_87_ab_7__31_), .B(
        u5_mult_87_CARRYB_6__31_), .CI(u5_mult_87_SUMB_6__32_), .CO(
        u5_mult_87_CARRYB_7__31_), .S(u5_mult_87_SUMB_7__31_) );
  FA_X1 u5_mult_87_S2_7_30 ( .A(u5_mult_87_ab_7__30_), .B(
        u5_mult_87_CARRYB_6__30_), .CI(u5_mult_87_SUMB_6__31_), .CO(
        u5_mult_87_CARRYB_7__30_), .S(u5_mult_87_SUMB_7__30_) );
  FA_X1 u5_mult_87_S2_7_29 ( .A(u5_mult_87_ab_7__29_), .B(
        u5_mult_87_CARRYB_6__29_), .CI(u5_mult_87_SUMB_6__30_), .CO(
        u5_mult_87_CARRYB_7__29_), .S(u5_mult_87_SUMB_7__29_) );
  FA_X1 u5_mult_87_S2_7_28 ( .A(u5_mult_87_ab_7__28_), .B(
        u5_mult_87_CARRYB_6__28_), .CI(u5_mult_87_SUMB_6__29_), .CO(
        u5_mult_87_CARRYB_7__28_), .S(u5_mult_87_SUMB_7__28_) );
  FA_X1 u5_mult_87_S2_7_27 ( .A(u5_mult_87_ab_7__27_), .B(
        u5_mult_87_CARRYB_6__27_), .CI(u5_mult_87_SUMB_6__28_), .CO(
        u5_mult_87_CARRYB_7__27_), .S(u5_mult_87_SUMB_7__27_) );
  FA_X1 u5_mult_87_S2_7_26 ( .A(u5_mult_87_ab_7__26_), .B(
        u5_mult_87_CARRYB_6__26_), .CI(u5_mult_87_SUMB_6__27_), .CO(
        u5_mult_87_CARRYB_7__26_), .S(u5_mult_87_SUMB_7__26_) );
  FA_X1 u5_mult_87_S2_7_25 ( .A(u5_mult_87_ab_7__25_), .B(
        u5_mult_87_CARRYB_6__25_), .CI(u5_mult_87_SUMB_6__26_), .CO(
        u5_mult_87_CARRYB_7__25_), .S(u5_mult_87_SUMB_7__25_) );
  FA_X1 u5_mult_87_S2_7_24 ( .A(u5_mult_87_ab_7__24_), .B(
        u5_mult_87_CARRYB_6__24_), .CI(u5_mult_87_SUMB_6__25_), .CO(
        u5_mult_87_CARRYB_7__24_), .S(u5_mult_87_SUMB_7__24_) );
  FA_X1 u5_mult_87_S2_7_23 ( .A(u5_mult_87_ab_7__23_), .B(
        u5_mult_87_CARRYB_6__23_), .CI(u5_mult_87_SUMB_6__24_), .CO(
        u5_mult_87_CARRYB_7__23_), .S(u5_mult_87_SUMB_7__23_) );
  FA_X1 u5_mult_87_S2_7_22 ( .A(u5_mult_87_ab_7__22_), .B(
        u5_mult_87_CARRYB_6__22_), .CI(u5_mult_87_SUMB_6__23_), .CO(
        u5_mult_87_CARRYB_7__22_), .S(u5_mult_87_SUMB_7__22_) );
  FA_X1 u5_mult_87_S2_7_21 ( .A(u5_mult_87_ab_7__21_), .B(
        u5_mult_87_CARRYB_6__21_), .CI(u5_mult_87_SUMB_6__22_), .CO(
        u5_mult_87_CARRYB_7__21_), .S(u5_mult_87_SUMB_7__21_) );
  FA_X1 u5_mult_87_S2_7_20 ( .A(u5_mult_87_ab_7__20_), .B(
        u5_mult_87_CARRYB_6__20_), .CI(u5_mult_87_SUMB_6__21_), .CO(
        u5_mult_87_CARRYB_7__20_), .S(u5_mult_87_SUMB_7__20_) );
  FA_X1 u5_mult_87_S2_7_19 ( .A(u5_mult_87_ab_7__19_), .B(
        u5_mult_87_CARRYB_6__19_), .CI(u5_mult_87_SUMB_6__20_), .CO(
        u5_mult_87_CARRYB_7__19_), .S(u5_mult_87_SUMB_7__19_) );
  FA_X1 u5_mult_87_S2_7_18 ( .A(u5_mult_87_ab_7__18_), .B(
        u5_mult_87_CARRYB_6__18_), .CI(u5_mult_87_SUMB_6__19_), .CO(
        u5_mult_87_CARRYB_7__18_), .S(u5_mult_87_SUMB_7__18_) );
  FA_X1 u5_mult_87_S2_7_17 ( .A(u5_mult_87_ab_7__17_), .B(
        u5_mult_87_CARRYB_6__17_), .CI(u5_mult_87_SUMB_6__18_), .CO(
        u5_mult_87_CARRYB_7__17_), .S(u5_mult_87_SUMB_7__17_) );
  FA_X1 u5_mult_87_S2_7_16 ( .A(u5_mult_87_ab_7__16_), .B(
        u5_mult_87_CARRYB_6__16_), .CI(u5_mult_87_SUMB_6__17_), .CO(
        u5_mult_87_CARRYB_7__16_), .S(u5_mult_87_SUMB_7__16_) );
  FA_X1 u5_mult_87_S2_7_15 ( .A(u5_mult_87_ab_7__15_), .B(
        u5_mult_87_CARRYB_6__15_), .CI(u5_mult_87_SUMB_6__16_), .CO(
        u5_mult_87_CARRYB_7__15_), .S(u5_mult_87_SUMB_7__15_) );
  FA_X1 u5_mult_87_S2_7_14 ( .A(u5_mult_87_ab_7__14_), .B(
        u5_mult_87_CARRYB_6__14_), .CI(u5_mult_87_SUMB_6__15_), .CO(
        u5_mult_87_CARRYB_7__14_), .S(u5_mult_87_SUMB_7__14_) );
  FA_X1 u5_mult_87_S2_7_13 ( .A(u5_mult_87_ab_7__13_), .B(
        u5_mult_87_CARRYB_6__13_), .CI(u5_mult_87_SUMB_6__14_), .CO(
        u5_mult_87_CARRYB_7__13_), .S(u5_mult_87_SUMB_7__13_) );
  FA_X1 u5_mult_87_S2_7_12 ( .A(u5_mult_87_ab_7__12_), .B(
        u5_mult_87_CARRYB_6__12_), .CI(u5_mult_87_SUMB_6__13_), .CO(
        u5_mult_87_CARRYB_7__12_), .S(u5_mult_87_SUMB_7__12_) );
  FA_X1 u5_mult_87_S2_7_11 ( .A(u5_mult_87_ab_7__11_), .B(
        u5_mult_87_CARRYB_6__11_), .CI(u5_mult_87_SUMB_6__12_), .CO(
        u5_mult_87_CARRYB_7__11_), .S(u5_mult_87_SUMB_7__11_) );
  FA_X1 u5_mult_87_S2_7_10 ( .A(u5_mult_87_ab_7__10_), .B(
        u5_mult_87_CARRYB_6__10_), .CI(u5_mult_87_SUMB_6__11_), .CO(
        u5_mult_87_CARRYB_7__10_), .S(u5_mult_87_SUMB_7__10_) );
  FA_X1 u5_mult_87_S2_7_9 ( .A(u5_mult_87_ab_7__9_), .B(
        u5_mult_87_CARRYB_6__9_), .CI(u5_mult_87_SUMB_6__10_), .CO(
        u5_mult_87_CARRYB_7__9_), .S(u5_mult_87_SUMB_7__9_) );
  FA_X1 u5_mult_87_S2_7_8 ( .A(u5_mult_87_ab_7__8_), .B(
        u5_mult_87_CARRYB_6__8_), .CI(u5_mult_87_SUMB_6__9_), .CO(
        u5_mult_87_CARRYB_7__8_), .S(u5_mult_87_SUMB_7__8_) );
  FA_X1 u5_mult_87_S2_7_7 ( .A(u5_mult_87_ab_7__7_), .B(
        u5_mult_87_CARRYB_6__7_), .CI(u5_mult_87_SUMB_6__8_), .CO(
        u5_mult_87_CARRYB_7__7_), .S(u5_mult_87_SUMB_7__7_) );
  FA_X1 u5_mult_87_S2_7_6 ( .A(u5_mult_87_ab_7__6_), .B(
        u5_mult_87_CARRYB_6__6_), .CI(u5_mult_87_SUMB_6__7_), .CO(
        u5_mult_87_CARRYB_7__6_), .S(u5_mult_87_SUMB_7__6_) );
  FA_X1 u5_mult_87_S2_7_5 ( .A(u5_mult_87_ab_7__5_), .B(
        u5_mult_87_CARRYB_6__5_), .CI(u5_mult_87_SUMB_6__6_), .CO(
        u5_mult_87_CARRYB_7__5_), .S(u5_mult_87_SUMB_7__5_) );
  FA_X1 u5_mult_87_S2_7_4 ( .A(u5_mult_87_ab_7__4_), .B(
        u5_mult_87_CARRYB_6__4_), .CI(u5_mult_87_SUMB_6__5_), .CO(
        u5_mult_87_CARRYB_7__4_), .S(u5_mult_87_SUMB_7__4_) );
  FA_X1 u5_mult_87_S2_7_3 ( .A(u5_mult_87_ab_7__3_), .B(
        u5_mult_87_CARRYB_6__3_), .CI(u5_mult_87_SUMB_6__4_), .CO(
        u5_mult_87_CARRYB_7__3_), .S(u5_mult_87_SUMB_7__3_) );
  FA_X1 u5_mult_87_S2_7_2 ( .A(u5_mult_87_ab_7__2_), .B(
        u5_mult_87_CARRYB_6__2_), .CI(u5_mult_87_SUMB_6__3_), .CO(
        u5_mult_87_CARRYB_7__2_), .S(u5_mult_87_SUMB_7__2_) );
  FA_X1 u5_mult_87_S2_7_1 ( .A(u5_mult_87_ab_7__1_), .B(
        u5_mult_87_CARRYB_6__1_), .CI(u5_mult_87_SUMB_6__2_), .CO(
        u5_mult_87_CARRYB_7__1_), .S(u5_mult_87_SUMB_7__1_) );
  FA_X1 u5_mult_87_S1_7_0 ( .A(u5_mult_87_ab_7__0_), .B(
        u5_mult_87_CARRYB_6__0_), .CI(u5_mult_87_SUMB_6__1_), .CO(
        u5_mult_87_CARRYB_7__0_), .S(u5_N7) );
  FA_X1 u5_mult_87_S3_8_51 ( .A(u5_mult_87_ab_8__51_), .B(
        u5_mult_87_CARRYB_7__51_), .CI(u5_mult_87_ab_7__52_), .CO(
        u5_mult_87_CARRYB_8__51_), .S(u5_mult_87_SUMB_8__51_) );
  FA_X1 u5_mult_87_S2_8_50 ( .A(u5_mult_87_ab_8__50_), .B(
        u5_mult_87_CARRYB_7__50_), .CI(u5_mult_87_SUMB_7__51_), .CO(
        u5_mult_87_CARRYB_8__50_), .S(u5_mult_87_SUMB_8__50_) );
  FA_X1 u5_mult_87_S2_8_49 ( .A(u5_mult_87_ab_8__49_), .B(
        u5_mult_87_CARRYB_7__49_), .CI(u5_mult_87_SUMB_7__50_), .CO(
        u5_mult_87_CARRYB_8__49_), .S(u5_mult_87_SUMB_8__49_) );
  FA_X1 u5_mult_87_S2_8_48 ( .A(u5_mult_87_ab_8__48_), .B(
        u5_mult_87_CARRYB_7__48_), .CI(u5_mult_87_SUMB_7__49_), .CO(
        u5_mult_87_CARRYB_8__48_), .S(u5_mult_87_SUMB_8__48_) );
  FA_X1 u5_mult_87_S2_8_47 ( .A(u5_mult_87_ab_8__47_), .B(
        u5_mult_87_CARRYB_7__47_), .CI(u5_mult_87_SUMB_7__48_), .CO(
        u5_mult_87_CARRYB_8__47_), .S(u5_mult_87_SUMB_8__47_) );
  FA_X1 u5_mult_87_S2_8_46 ( .A(u5_mult_87_ab_8__46_), .B(
        u5_mult_87_CARRYB_7__46_), .CI(u5_mult_87_SUMB_7__47_), .CO(
        u5_mult_87_CARRYB_8__46_), .S(u5_mult_87_SUMB_8__46_) );
  FA_X1 u5_mult_87_S2_8_45 ( .A(u5_mult_87_ab_8__45_), .B(
        u5_mult_87_CARRYB_7__45_), .CI(u5_mult_87_SUMB_7__46_), .CO(
        u5_mult_87_CARRYB_8__45_), .S(u5_mult_87_SUMB_8__45_) );
  FA_X1 u5_mult_87_S2_8_44 ( .A(u5_mult_87_ab_8__44_), .B(
        u5_mult_87_CARRYB_7__44_), .CI(u5_mult_87_SUMB_7__45_), .CO(
        u5_mult_87_CARRYB_8__44_), .S(u5_mult_87_SUMB_8__44_) );
  FA_X1 u5_mult_87_S2_8_43 ( .A(u5_mult_87_ab_8__43_), .B(
        u5_mult_87_CARRYB_7__43_), .CI(u5_mult_87_SUMB_7__44_), .CO(
        u5_mult_87_CARRYB_8__43_), .S(u5_mult_87_SUMB_8__43_) );
  FA_X1 u5_mult_87_S2_8_42 ( .A(u5_mult_87_ab_8__42_), .B(
        u5_mult_87_CARRYB_7__42_), .CI(u5_mult_87_SUMB_7__43_), .CO(
        u5_mult_87_CARRYB_8__42_), .S(u5_mult_87_SUMB_8__42_) );
  FA_X1 u5_mult_87_S2_8_41 ( .A(u5_mult_87_ab_8__41_), .B(
        u5_mult_87_CARRYB_7__41_), .CI(u5_mult_87_SUMB_7__42_), .CO(
        u5_mult_87_CARRYB_8__41_), .S(u5_mult_87_SUMB_8__41_) );
  FA_X1 u5_mult_87_S2_8_40 ( .A(u5_mult_87_ab_8__40_), .B(
        u5_mult_87_CARRYB_7__40_), .CI(u5_mult_87_SUMB_7__41_), .CO(
        u5_mult_87_CARRYB_8__40_), .S(u5_mult_87_SUMB_8__40_) );
  FA_X1 u5_mult_87_S2_8_39 ( .A(u5_mult_87_ab_8__39_), .B(
        u5_mult_87_CARRYB_7__39_), .CI(u5_mult_87_SUMB_7__40_), .CO(
        u5_mult_87_CARRYB_8__39_), .S(u5_mult_87_SUMB_8__39_) );
  FA_X1 u5_mult_87_S2_8_38 ( .A(u5_mult_87_ab_8__38_), .B(
        u5_mult_87_CARRYB_7__38_), .CI(u5_mult_87_SUMB_7__39_), .CO(
        u5_mult_87_CARRYB_8__38_), .S(u5_mult_87_SUMB_8__38_) );
  FA_X1 u5_mult_87_S2_8_37 ( .A(u5_mult_87_ab_8__37_), .B(
        u5_mult_87_CARRYB_7__37_), .CI(u5_mult_87_SUMB_7__38_), .CO(
        u5_mult_87_CARRYB_8__37_), .S(u5_mult_87_SUMB_8__37_) );
  FA_X1 u5_mult_87_S2_8_36 ( .A(u5_mult_87_ab_8__36_), .B(
        u5_mult_87_CARRYB_7__36_), .CI(u5_mult_87_SUMB_7__37_), .CO(
        u5_mult_87_CARRYB_8__36_), .S(u5_mult_87_SUMB_8__36_) );
  FA_X1 u5_mult_87_S2_8_35 ( .A(u5_mult_87_ab_8__35_), .B(
        u5_mult_87_CARRYB_7__35_), .CI(u5_mult_87_SUMB_7__36_), .CO(
        u5_mult_87_CARRYB_8__35_), .S(u5_mult_87_SUMB_8__35_) );
  FA_X1 u5_mult_87_S2_8_34 ( .A(u5_mult_87_ab_8__34_), .B(
        u5_mult_87_CARRYB_7__34_), .CI(u5_mult_87_SUMB_7__35_), .CO(
        u5_mult_87_CARRYB_8__34_), .S(u5_mult_87_SUMB_8__34_) );
  FA_X1 u5_mult_87_S2_8_33 ( .A(u5_mult_87_ab_8__33_), .B(
        u5_mult_87_CARRYB_7__33_), .CI(u5_mult_87_SUMB_7__34_), .CO(
        u5_mult_87_CARRYB_8__33_), .S(u5_mult_87_SUMB_8__33_) );
  FA_X1 u5_mult_87_S2_8_32 ( .A(u5_mult_87_ab_8__32_), .B(
        u5_mult_87_CARRYB_7__32_), .CI(u5_mult_87_SUMB_7__33_), .CO(
        u5_mult_87_CARRYB_8__32_), .S(u5_mult_87_SUMB_8__32_) );
  FA_X1 u5_mult_87_S2_8_31 ( .A(u5_mult_87_ab_8__31_), .B(
        u5_mult_87_CARRYB_7__31_), .CI(u5_mult_87_SUMB_7__32_), .CO(
        u5_mult_87_CARRYB_8__31_), .S(u5_mult_87_SUMB_8__31_) );
  FA_X1 u5_mult_87_S2_8_30 ( .A(u5_mult_87_ab_8__30_), .B(
        u5_mult_87_CARRYB_7__30_), .CI(u5_mult_87_SUMB_7__31_), .CO(
        u5_mult_87_CARRYB_8__30_), .S(u5_mult_87_SUMB_8__30_) );
  FA_X1 u5_mult_87_S2_8_29 ( .A(u5_mult_87_ab_8__29_), .B(
        u5_mult_87_CARRYB_7__29_), .CI(u5_mult_87_SUMB_7__30_), .CO(
        u5_mult_87_CARRYB_8__29_), .S(u5_mult_87_SUMB_8__29_) );
  FA_X1 u5_mult_87_S2_8_28 ( .A(u5_mult_87_ab_8__28_), .B(
        u5_mult_87_CARRYB_7__28_), .CI(u5_mult_87_SUMB_7__29_), .CO(
        u5_mult_87_CARRYB_8__28_), .S(u5_mult_87_SUMB_8__28_) );
  FA_X1 u5_mult_87_S2_8_27 ( .A(u5_mult_87_ab_8__27_), .B(
        u5_mult_87_CARRYB_7__27_), .CI(u5_mult_87_SUMB_7__28_), .CO(
        u5_mult_87_CARRYB_8__27_), .S(u5_mult_87_SUMB_8__27_) );
  FA_X1 u5_mult_87_S2_8_26 ( .A(u5_mult_87_ab_8__26_), .B(
        u5_mult_87_CARRYB_7__26_), .CI(u5_mult_87_SUMB_7__27_), .CO(
        u5_mult_87_CARRYB_8__26_), .S(u5_mult_87_SUMB_8__26_) );
  FA_X1 u5_mult_87_S2_8_25 ( .A(u5_mult_87_ab_8__25_), .B(
        u5_mult_87_CARRYB_7__25_), .CI(u5_mult_87_SUMB_7__26_), .CO(
        u5_mult_87_CARRYB_8__25_), .S(u5_mult_87_SUMB_8__25_) );
  FA_X1 u5_mult_87_S2_8_24 ( .A(u5_mult_87_ab_8__24_), .B(
        u5_mult_87_CARRYB_7__24_), .CI(u5_mult_87_SUMB_7__25_), .CO(
        u5_mult_87_CARRYB_8__24_), .S(u5_mult_87_SUMB_8__24_) );
  FA_X1 u5_mult_87_S2_8_23 ( .A(u5_mult_87_ab_8__23_), .B(
        u5_mult_87_CARRYB_7__23_), .CI(u5_mult_87_SUMB_7__24_), .CO(
        u5_mult_87_CARRYB_8__23_), .S(u5_mult_87_SUMB_8__23_) );
  FA_X1 u5_mult_87_S2_8_22 ( .A(u5_mult_87_ab_8__22_), .B(
        u5_mult_87_CARRYB_7__22_), .CI(u5_mult_87_SUMB_7__23_), .CO(
        u5_mult_87_CARRYB_8__22_), .S(u5_mult_87_SUMB_8__22_) );
  FA_X1 u5_mult_87_S2_8_21 ( .A(u5_mult_87_ab_8__21_), .B(
        u5_mult_87_CARRYB_7__21_), .CI(u5_mult_87_SUMB_7__22_), .CO(
        u5_mult_87_CARRYB_8__21_), .S(u5_mult_87_SUMB_8__21_) );
  FA_X1 u5_mult_87_S2_8_20 ( .A(u5_mult_87_ab_8__20_), .B(
        u5_mult_87_CARRYB_7__20_), .CI(u5_mult_87_SUMB_7__21_), .CO(
        u5_mult_87_CARRYB_8__20_), .S(u5_mult_87_SUMB_8__20_) );
  FA_X1 u5_mult_87_S2_8_19 ( .A(u5_mult_87_ab_8__19_), .B(
        u5_mult_87_CARRYB_7__19_), .CI(u5_mult_87_SUMB_7__20_), .CO(
        u5_mult_87_CARRYB_8__19_), .S(u5_mult_87_SUMB_8__19_) );
  FA_X1 u5_mult_87_S2_8_18 ( .A(u5_mult_87_ab_8__18_), .B(
        u5_mult_87_CARRYB_7__18_), .CI(u5_mult_87_SUMB_7__19_), .CO(
        u5_mult_87_CARRYB_8__18_), .S(u5_mult_87_SUMB_8__18_) );
  FA_X1 u5_mult_87_S2_8_17 ( .A(u5_mult_87_ab_8__17_), .B(
        u5_mult_87_CARRYB_7__17_), .CI(u5_mult_87_SUMB_7__18_), .CO(
        u5_mult_87_CARRYB_8__17_), .S(u5_mult_87_SUMB_8__17_) );
  FA_X1 u5_mult_87_S2_8_16 ( .A(u5_mult_87_ab_8__16_), .B(
        u5_mult_87_CARRYB_7__16_), .CI(u5_mult_87_SUMB_7__17_), .CO(
        u5_mult_87_CARRYB_8__16_), .S(u5_mult_87_SUMB_8__16_) );
  FA_X1 u5_mult_87_S2_8_15 ( .A(u5_mult_87_ab_8__15_), .B(
        u5_mult_87_CARRYB_7__15_), .CI(u5_mult_87_SUMB_7__16_), .CO(
        u5_mult_87_CARRYB_8__15_), .S(u5_mult_87_SUMB_8__15_) );
  FA_X1 u5_mult_87_S2_8_14 ( .A(u5_mult_87_ab_8__14_), .B(
        u5_mult_87_CARRYB_7__14_), .CI(u5_mult_87_SUMB_7__15_), .CO(
        u5_mult_87_CARRYB_8__14_), .S(u5_mult_87_SUMB_8__14_) );
  FA_X1 u5_mult_87_S2_8_13 ( .A(u5_mult_87_ab_8__13_), .B(
        u5_mult_87_CARRYB_7__13_), .CI(u5_mult_87_SUMB_7__14_), .CO(
        u5_mult_87_CARRYB_8__13_), .S(u5_mult_87_SUMB_8__13_) );
  FA_X1 u5_mult_87_S2_8_12 ( .A(u5_mult_87_ab_8__12_), .B(
        u5_mult_87_CARRYB_7__12_), .CI(u5_mult_87_SUMB_7__13_), .CO(
        u5_mult_87_CARRYB_8__12_), .S(u5_mult_87_SUMB_8__12_) );
  FA_X1 u5_mult_87_S2_8_11 ( .A(u5_mult_87_ab_8__11_), .B(
        u5_mult_87_CARRYB_7__11_), .CI(u5_mult_87_SUMB_7__12_), .CO(
        u5_mult_87_CARRYB_8__11_), .S(u5_mult_87_SUMB_8__11_) );
  FA_X1 u5_mult_87_S2_8_10 ( .A(u5_mult_87_ab_8__10_), .B(
        u5_mult_87_CARRYB_7__10_), .CI(u5_mult_87_SUMB_7__11_), .CO(
        u5_mult_87_CARRYB_8__10_), .S(u5_mult_87_SUMB_8__10_) );
  FA_X1 u5_mult_87_S2_8_9 ( .A(u5_mult_87_ab_8__9_), .B(
        u5_mult_87_CARRYB_7__9_), .CI(u5_mult_87_SUMB_7__10_), .CO(
        u5_mult_87_CARRYB_8__9_), .S(u5_mult_87_SUMB_8__9_) );
  FA_X1 u5_mult_87_S2_8_8 ( .A(u5_mult_87_ab_8__8_), .B(
        u5_mult_87_CARRYB_7__8_), .CI(u5_mult_87_SUMB_7__9_), .CO(
        u5_mult_87_CARRYB_8__8_), .S(u5_mult_87_SUMB_8__8_) );
  FA_X1 u5_mult_87_S2_8_7 ( .A(u5_mult_87_ab_8__7_), .B(
        u5_mult_87_CARRYB_7__7_), .CI(u5_mult_87_SUMB_7__8_), .CO(
        u5_mult_87_CARRYB_8__7_), .S(u5_mult_87_SUMB_8__7_) );
  FA_X1 u5_mult_87_S2_8_6 ( .A(u5_mult_87_ab_8__6_), .B(
        u5_mult_87_CARRYB_7__6_), .CI(u5_mult_87_SUMB_7__7_), .CO(
        u5_mult_87_CARRYB_8__6_), .S(u5_mult_87_SUMB_8__6_) );
  FA_X1 u5_mult_87_S2_8_5 ( .A(u5_mult_87_ab_8__5_), .B(
        u5_mult_87_CARRYB_7__5_), .CI(u5_mult_87_SUMB_7__6_), .CO(
        u5_mult_87_CARRYB_8__5_), .S(u5_mult_87_SUMB_8__5_) );
  FA_X1 u5_mult_87_S2_8_4 ( .A(u5_mult_87_ab_8__4_), .B(
        u5_mult_87_CARRYB_7__4_), .CI(u5_mult_87_SUMB_7__5_), .CO(
        u5_mult_87_CARRYB_8__4_), .S(u5_mult_87_SUMB_8__4_) );
  FA_X1 u5_mult_87_S2_8_3 ( .A(u5_mult_87_ab_8__3_), .B(
        u5_mult_87_CARRYB_7__3_), .CI(u5_mult_87_SUMB_7__4_), .CO(
        u5_mult_87_CARRYB_8__3_), .S(u5_mult_87_SUMB_8__3_) );
  FA_X1 u5_mult_87_S2_8_2 ( .A(u5_mult_87_ab_8__2_), .B(
        u5_mult_87_CARRYB_7__2_), .CI(u5_mult_87_SUMB_7__3_), .CO(
        u5_mult_87_CARRYB_8__2_), .S(u5_mult_87_SUMB_8__2_) );
  FA_X1 u5_mult_87_S2_8_1 ( .A(u5_mult_87_ab_8__1_), .B(
        u5_mult_87_CARRYB_7__1_), .CI(u5_mult_87_SUMB_7__2_), .CO(
        u5_mult_87_CARRYB_8__1_), .S(u5_mult_87_SUMB_8__1_) );
  FA_X1 u5_mult_87_S1_8_0 ( .A(u5_mult_87_ab_8__0_), .B(
        u5_mult_87_CARRYB_7__0_), .CI(u5_mult_87_SUMB_7__1_), .CO(
        u5_mult_87_CARRYB_8__0_), .S(u5_N8) );
  FA_X1 u5_mult_87_S3_9_51 ( .A(u5_mult_87_ab_9__51_), .B(
        u5_mult_87_CARRYB_8__51_), .CI(u5_mult_87_ab_8__52_), .CO(
        u5_mult_87_CARRYB_9__51_), .S(u5_mult_87_SUMB_9__51_) );
  FA_X1 u5_mult_87_S2_9_50 ( .A(u5_mult_87_ab_9__50_), .B(
        u5_mult_87_CARRYB_8__50_), .CI(u5_mult_87_SUMB_8__51_), .CO(
        u5_mult_87_CARRYB_9__50_), .S(u5_mult_87_SUMB_9__50_) );
  FA_X1 u5_mult_87_S2_9_49 ( .A(u5_mult_87_ab_9__49_), .B(
        u5_mult_87_CARRYB_8__49_), .CI(u5_mult_87_SUMB_8__50_), .CO(
        u5_mult_87_CARRYB_9__49_), .S(u5_mult_87_SUMB_9__49_) );
  FA_X1 u5_mult_87_S2_9_48 ( .A(u5_mult_87_ab_9__48_), .B(
        u5_mult_87_CARRYB_8__48_), .CI(u5_mult_87_SUMB_8__49_), .CO(
        u5_mult_87_CARRYB_9__48_), .S(u5_mult_87_SUMB_9__48_) );
  FA_X1 u5_mult_87_S2_9_47 ( .A(u5_mult_87_ab_9__47_), .B(
        u5_mult_87_CARRYB_8__47_), .CI(u5_mult_87_SUMB_8__48_), .CO(
        u5_mult_87_CARRYB_9__47_), .S(u5_mult_87_SUMB_9__47_) );
  FA_X1 u5_mult_87_S2_9_46 ( .A(u5_mult_87_ab_9__46_), .B(
        u5_mult_87_CARRYB_8__46_), .CI(u5_mult_87_SUMB_8__47_), .CO(
        u5_mult_87_CARRYB_9__46_), .S(u5_mult_87_SUMB_9__46_) );
  FA_X1 u5_mult_87_S2_9_45 ( .A(u5_mult_87_ab_9__45_), .B(
        u5_mult_87_CARRYB_8__45_), .CI(u5_mult_87_SUMB_8__46_), .CO(
        u5_mult_87_CARRYB_9__45_), .S(u5_mult_87_SUMB_9__45_) );
  FA_X1 u5_mult_87_S2_9_44 ( .A(u5_mult_87_ab_9__44_), .B(
        u5_mult_87_CARRYB_8__44_), .CI(u5_mult_87_SUMB_8__45_), .CO(
        u5_mult_87_CARRYB_9__44_), .S(u5_mult_87_SUMB_9__44_) );
  FA_X1 u5_mult_87_S2_9_43 ( .A(u5_mult_87_ab_9__43_), .B(
        u5_mult_87_CARRYB_8__43_), .CI(u5_mult_87_SUMB_8__44_), .CO(
        u5_mult_87_CARRYB_9__43_), .S(u5_mult_87_SUMB_9__43_) );
  FA_X1 u5_mult_87_S2_9_42 ( .A(u5_mult_87_ab_9__42_), .B(
        u5_mult_87_CARRYB_8__42_), .CI(u5_mult_87_SUMB_8__43_), .CO(
        u5_mult_87_CARRYB_9__42_), .S(u5_mult_87_SUMB_9__42_) );
  FA_X1 u5_mult_87_S2_9_41 ( .A(u5_mult_87_ab_9__41_), .B(
        u5_mult_87_CARRYB_8__41_), .CI(u5_mult_87_SUMB_8__42_), .CO(
        u5_mult_87_CARRYB_9__41_), .S(u5_mult_87_SUMB_9__41_) );
  FA_X1 u5_mult_87_S2_9_40 ( .A(u5_mult_87_ab_9__40_), .B(
        u5_mult_87_CARRYB_8__40_), .CI(u5_mult_87_SUMB_8__41_), .CO(
        u5_mult_87_CARRYB_9__40_), .S(u5_mult_87_SUMB_9__40_) );
  FA_X1 u5_mult_87_S2_9_39 ( .A(u5_mult_87_ab_9__39_), .B(
        u5_mult_87_CARRYB_8__39_), .CI(u5_mult_87_SUMB_8__40_), .CO(
        u5_mult_87_CARRYB_9__39_), .S(u5_mult_87_SUMB_9__39_) );
  FA_X1 u5_mult_87_S2_9_38 ( .A(u5_mult_87_ab_9__38_), .B(
        u5_mult_87_CARRYB_8__38_), .CI(u5_mult_87_SUMB_8__39_), .CO(
        u5_mult_87_CARRYB_9__38_), .S(u5_mult_87_SUMB_9__38_) );
  FA_X1 u5_mult_87_S2_9_37 ( .A(u5_mult_87_ab_9__37_), .B(
        u5_mult_87_CARRYB_8__37_), .CI(u5_mult_87_SUMB_8__38_), .CO(
        u5_mult_87_CARRYB_9__37_), .S(u5_mult_87_SUMB_9__37_) );
  FA_X1 u5_mult_87_S2_9_36 ( .A(u5_mult_87_ab_9__36_), .B(
        u5_mult_87_CARRYB_8__36_), .CI(u5_mult_87_SUMB_8__37_), .CO(
        u5_mult_87_CARRYB_9__36_), .S(u5_mult_87_SUMB_9__36_) );
  FA_X1 u5_mult_87_S2_9_35 ( .A(u5_mult_87_ab_9__35_), .B(
        u5_mult_87_CARRYB_8__35_), .CI(u5_mult_87_SUMB_8__36_), .CO(
        u5_mult_87_CARRYB_9__35_), .S(u5_mult_87_SUMB_9__35_) );
  FA_X1 u5_mult_87_S2_9_34 ( .A(u5_mult_87_ab_9__34_), .B(
        u5_mult_87_CARRYB_8__34_), .CI(u5_mult_87_SUMB_8__35_), .CO(
        u5_mult_87_CARRYB_9__34_), .S(u5_mult_87_SUMB_9__34_) );
  FA_X1 u5_mult_87_S2_9_33 ( .A(u5_mult_87_ab_9__33_), .B(
        u5_mult_87_CARRYB_8__33_), .CI(u5_mult_87_SUMB_8__34_), .CO(
        u5_mult_87_CARRYB_9__33_), .S(u5_mult_87_SUMB_9__33_) );
  FA_X1 u5_mult_87_S2_9_32 ( .A(u5_mult_87_ab_9__32_), .B(
        u5_mult_87_CARRYB_8__32_), .CI(u5_mult_87_SUMB_8__33_), .CO(
        u5_mult_87_CARRYB_9__32_), .S(u5_mult_87_SUMB_9__32_) );
  FA_X1 u5_mult_87_S2_9_31 ( .A(u5_mult_87_ab_9__31_), .B(
        u5_mult_87_CARRYB_8__31_), .CI(u5_mult_87_SUMB_8__32_), .CO(
        u5_mult_87_CARRYB_9__31_), .S(u5_mult_87_SUMB_9__31_) );
  FA_X1 u5_mult_87_S2_9_30 ( .A(u5_mult_87_ab_9__30_), .B(
        u5_mult_87_CARRYB_8__30_), .CI(u5_mult_87_SUMB_8__31_), .CO(
        u5_mult_87_CARRYB_9__30_), .S(u5_mult_87_SUMB_9__30_) );
  FA_X1 u5_mult_87_S2_9_29 ( .A(u5_mult_87_ab_9__29_), .B(
        u5_mult_87_CARRYB_8__29_), .CI(u5_mult_87_SUMB_8__30_), .CO(
        u5_mult_87_CARRYB_9__29_), .S(u5_mult_87_SUMB_9__29_) );
  FA_X1 u5_mult_87_S2_9_28 ( .A(u5_mult_87_ab_9__28_), .B(
        u5_mult_87_CARRYB_8__28_), .CI(u5_mult_87_SUMB_8__29_), .CO(
        u5_mult_87_CARRYB_9__28_), .S(u5_mult_87_SUMB_9__28_) );
  FA_X1 u5_mult_87_S2_9_27 ( .A(u5_mult_87_ab_9__27_), .B(
        u5_mult_87_CARRYB_8__27_), .CI(u5_mult_87_SUMB_8__28_), .CO(
        u5_mult_87_CARRYB_9__27_), .S(u5_mult_87_SUMB_9__27_) );
  FA_X1 u5_mult_87_S2_9_26 ( .A(u5_mult_87_ab_9__26_), .B(
        u5_mult_87_CARRYB_8__26_), .CI(u5_mult_87_SUMB_8__27_), .CO(
        u5_mult_87_CARRYB_9__26_), .S(u5_mult_87_SUMB_9__26_) );
  FA_X1 u5_mult_87_S2_9_25 ( .A(u5_mult_87_ab_9__25_), .B(
        u5_mult_87_CARRYB_8__25_), .CI(u5_mult_87_SUMB_8__26_), .CO(
        u5_mult_87_CARRYB_9__25_), .S(u5_mult_87_SUMB_9__25_) );
  FA_X1 u5_mult_87_S2_9_24 ( .A(u5_mult_87_ab_9__24_), .B(
        u5_mult_87_CARRYB_8__24_), .CI(u5_mult_87_SUMB_8__25_), .CO(
        u5_mult_87_CARRYB_9__24_), .S(u5_mult_87_SUMB_9__24_) );
  FA_X1 u5_mult_87_S2_9_23 ( .A(u5_mult_87_ab_9__23_), .B(
        u5_mult_87_CARRYB_8__23_), .CI(u5_mult_87_SUMB_8__24_), .CO(
        u5_mult_87_CARRYB_9__23_), .S(u5_mult_87_SUMB_9__23_) );
  FA_X1 u5_mult_87_S2_9_22 ( .A(u5_mult_87_ab_9__22_), .B(
        u5_mult_87_CARRYB_8__22_), .CI(u5_mult_87_SUMB_8__23_), .CO(
        u5_mult_87_CARRYB_9__22_), .S(u5_mult_87_SUMB_9__22_) );
  FA_X1 u5_mult_87_S2_9_21 ( .A(u5_mult_87_ab_9__21_), .B(
        u5_mult_87_CARRYB_8__21_), .CI(u5_mult_87_SUMB_8__22_), .CO(
        u5_mult_87_CARRYB_9__21_), .S(u5_mult_87_SUMB_9__21_) );
  FA_X1 u5_mult_87_S2_9_20 ( .A(u5_mult_87_ab_9__20_), .B(
        u5_mult_87_CARRYB_8__20_), .CI(u5_mult_87_SUMB_8__21_), .CO(
        u5_mult_87_CARRYB_9__20_), .S(u5_mult_87_SUMB_9__20_) );
  FA_X1 u5_mult_87_S2_9_19 ( .A(u5_mult_87_ab_9__19_), .B(
        u5_mult_87_CARRYB_8__19_), .CI(u5_mult_87_SUMB_8__20_), .CO(
        u5_mult_87_CARRYB_9__19_), .S(u5_mult_87_SUMB_9__19_) );
  FA_X1 u5_mult_87_S2_9_18 ( .A(u5_mult_87_ab_9__18_), .B(
        u5_mult_87_CARRYB_8__18_), .CI(u5_mult_87_SUMB_8__19_), .CO(
        u5_mult_87_CARRYB_9__18_), .S(u5_mult_87_SUMB_9__18_) );
  FA_X1 u5_mult_87_S2_9_17 ( .A(u5_mult_87_ab_9__17_), .B(
        u5_mult_87_CARRYB_8__17_), .CI(u5_mult_87_SUMB_8__18_), .CO(
        u5_mult_87_CARRYB_9__17_), .S(u5_mult_87_SUMB_9__17_) );
  FA_X1 u5_mult_87_S2_9_16 ( .A(u5_mult_87_ab_9__16_), .B(
        u5_mult_87_CARRYB_8__16_), .CI(u5_mult_87_SUMB_8__17_), .CO(
        u5_mult_87_CARRYB_9__16_), .S(u5_mult_87_SUMB_9__16_) );
  FA_X1 u5_mult_87_S2_9_15 ( .A(u5_mult_87_ab_9__15_), .B(
        u5_mult_87_CARRYB_8__15_), .CI(u5_mult_87_SUMB_8__16_), .CO(
        u5_mult_87_CARRYB_9__15_), .S(u5_mult_87_SUMB_9__15_) );
  FA_X1 u5_mult_87_S2_9_14 ( .A(u5_mult_87_ab_9__14_), .B(
        u5_mult_87_CARRYB_8__14_), .CI(u5_mult_87_SUMB_8__15_), .CO(
        u5_mult_87_CARRYB_9__14_), .S(u5_mult_87_SUMB_9__14_) );
  FA_X1 u5_mult_87_S2_9_13 ( .A(u5_mult_87_ab_9__13_), .B(
        u5_mult_87_CARRYB_8__13_), .CI(u5_mult_87_SUMB_8__14_), .CO(
        u5_mult_87_CARRYB_9__13_), .S(u5_mult_87_SUMB_9__13_) );
  FA_X1 u5_mult_87_S2_9_12 ( .A(u5_mult_87_ab_9__12_), .B(
        u5_mult_87_CARRYB_8__12_), .CI(u5_mult_87_SUMB_8__13_), .CO(
        u5_mult_87_CARRYB_9__12_), .S(u5_mult_87_SUMB_9__12_) );
  FA_X1 u5_mult_87_S2_9_11 ( .A(u5_mult_87_ab_9__11_), .B(
        u5_mult_87_CARRYB_8__11_), .CI(u5_mult_87_SUMB_8__12_), .CO(
        u5_mult_87_CARRYB_9__11_), .S(u5_mult_87_SUMB_9__11_) );
  FA_X1 u5_mult_87_S2_9_10 ( .A(u5_mult_87_ab_9__10_), .B(
        u5_mult_87_CARRYB_8__10_), .CI(u5_mult_87_SUMB_8__11_), .CO(
        u5_mult_87_CARRYB_9__10_), .S(u5_mult_87_SUMB_9__10_) );
  FA_X1 u5_mult_87_S2_9_9 ( .A(u5_mult_87_ab_9__9_), .B(
        u5_mult_87_CARRYB_8__9_), .CI(u5_mult_87_SUMB_8__10_), .CO(
        u5_mult_87_CARRYB_9__9_), .S(u5_mult_87_SUMB_9__9_) );
  FA_X1 u5_mult_87_S2_9_8 ( .A(u5_mult_87_ab_9__8_), .B(
        u5_mult_87_CARRYB_8__8_), .CI(u5_mult_87_SUMB_8__9_), .CO(
        u5_mult_87_CARRYB_9__8_), .S(u5_mult_87_SUMB_9__8_) );
  FA_X1 u5_mult_87_S2_9_7 ( .A(u5_mult_87_ab_9__7_), .B(
        u5_mult_87_CARRYB_8__7_), .CI(u5_mult_87_SUMB_8__8_), .CO(
        u5_mult_87_CARRYB_9__7_), .S(u5_mult_87_SUMB_9__7_) );
  FA_X1 u5_mult_87_S2_9_6 ( .A(u5_mult_87_ab_9__6_), .B(
        u5_mult_87_CARRYB_8__6_), .CI(u5_mult_87_SUMB_8__7_), .CO(
        u5_mult_87_CARRYB_9__6_), .S(u5_mult_87_SUMB_9__6_) );
  FA_X1 u5_mult_87_S2_9_5 ( .A(u5_mult_87_ab_9__5_), .B(
        u5_mult_87_CARRYB_8__5_), .CI(u5_mult_87_SUMB_8__6_), .CO(
        u5_mult_87_CARRYB_9__5_), .S(u5_mult_87_SUMB_9__5_) );
  FA_X1 u5_mult_87_S2_9_4 ( .A(u5_mult_87_ab_9__4_), .B(
        u5_mult_87_CARRYB_8__4_), .CI(u5_mult_87_SUMB_8__5_), .CO(
        u5_mult_87_CARRYB_9__4_), .S(u5_mult_87_SUMB_9__4_) );
  FA_X1 u5_mult_87_S2_9_3 ( .A(u5_mult_87_ab_9__3_), .B(
        u5_mult_87_CARRYB_8__3_), .CI(u5_mult_87_SUMB_8__4_), .CO(
        u5_mult_87_CARRYB_9__3_), .S(u5_mult_87_SUMB_9__3_) );
  FA_X1 u5_mult_87_S2_9_2 ( .A(u5_mult_87_ab_9__2_), .B(
        u5_mult_87_CARRYB_8__2_), .CI(u5_mult_87_SUMB_8__3_), .CO(
        u5_mult_87_CARRYB_9__2_), .S(u5_mult_87_SUMB_9__2_) );
  FA_X1 u5_mult_87_S2_9_1 ( .A(u5_mult_87_ab_9__1_), .B(
        u5_mult_87_CARRYB_8__1_), .CI(u5_mult_87_SUMB_8__2_), .CO(
        u5_mult_87_CARRYB_9__1_), .S(u5_mult_87_SUMB_9__1_) );
  FA_X1 u5_mult_87_S1_9_0 ( .A(u5_mult_87_ab_9__0_), .B(
        u5_mult_87_CARRYB_8__0_), .CI(u5_mult_87_SUMB_8__1_), .CO(
        u5_mult_87_CARRYB_9__0_), .S(u5_N9) );
  FA_X1 u5_mult_87_S3_10_51 ( .A(u5_mult_87_ab_10__51_), .B(
        u5_mult_87_CARRYB_9__51_), .CI(u5_mult_87_ab_9__52_), .CO(
        u5_mult_87_CARRYB_10__51_), .S(u5_mult_87_SUMB_10__51_) );
  FA_X1 u5_mult_87_S2_10_50 ( .A(u5_mult_87_ab_10__50_), .B(
        u5_mult_87_CARRYB_9__50_), .CI(u5_mult_87_SUMB_9__51_), .CO(
        u5_mult_87_CARRYB_10__50_), .S(u5_mult_87_SUMB_10__50_) );
  FA_X1 u5_mult_87_S2_10_49 ( .A(u5_mult_87_ab_10__49_), .B(
        u5_mult_87_CARRYB_9__49_), .CI(u5_mult_87_SUMB_9__50_), .CO(
        u5_mult_87_CARRYB_10__49_), .S(u5_mult_87_SUMB_10__49_) );
  FA_X1 u5_mult_87_S2_10_48 ( .A(u5_mult_87_ab_10__48_), .B(
        u5_mult_87_CARRYB_9__48_), .CI(u5_mult_87_SUMB_9__49_), .CO(
        u5_mult_87_CARRYB_10__48_), .S(u5_mult_87_SUMB_10__48_) );
  FA_X1 u5_mult_87_S2_10_47 ( .A(u5_mult_87_ab_10__47_), .B(
        u5_mult_87_CARRYB_9__47_), .CI(u5_mult_87_SUMB_9__48_), .CO(
        u5_mult_87_CARRYB_10__47_), .S(u5_mult_87_SUMB_10__47_) );
  FA_X1 u5_mult_87_S2_10_46 ( .A(u5_mult_87_ab_10__46_), .B(
        u5_mult_87_CARRYB_9__46_), .CI(u5_mult_87_SUMB_9__47_), .CO(
        u5_mult_87_CARRYB_10__46_), .S(u5_mult_87_SUMB_10__46_) );
  FA_X1 u5_mult_87_S2_10_45 ( .A(u5_mult_87_ab_10__45_), .B(
        u5_mult_87_CARRYB_9__45_), .CI(u5_mult_87_SUMB_9__46_), .CO(
        u5_mult_87_CARRYB_10__45_), .S(u5_mult_87_SUMB_10__45_) );
  FA_X1 u5_mult_87_S2_10_44 ( .A(u5_mult_87_ab_10__44_), .B(
        u5_mult_87_CARRYB_9__44_), .CI(u5_mult_87_SUMB_9__45_), .CO(
        u5_mult_87_CARRYB_10__44_), .S(u5_mult_87_SUMB_10__44_) );
  FA_X1 u5_mult_87_S2_10_43 ( .A(u5_mult_87_ab_10__43_), .B(
        u5_mult_87_CARRYB_9__43_), .CI(u5_mult_87_SUMB_9__44_), .CO(
        u5_mult_87_CARRYB_10__43_), .S(u5_mult_87_SUMB_10__43_) );
  FA_X1 u5_mult_87_S2_10_42 ( .A(u5_mult_87_ab_10__42_), .B(
        u5_mult_87_CARRYB_9__42_), .CI(u5_mult_87_SUMB_9__43_), .CO(
        u5_mult_87_CARRYB_10__42_), .S(u5_mult_87_SUMB_10__42_) );
  FA_X1 u5_mult_87_S2_10_41 ( .A(u5_mult_87_ab_10__41_), .B(
        u5_mult_87_CARRYB_9__41_), .CI(u5_mult_87_SUMB_9__42_), .CO(
        u5_mult_87_CARRYB_10__41_), .S(u5_mult_87_SUMB_10__41_) );
  FA_X1 u5_mult_87_S2_10_40 ( .A(u5_mult_87_ab_10__40_), .B(
        u5_mult_87_CARRYB_9__40_), .CI(u5_mult_87_SUMB_9__41_), .CO(
        u5_mult_87_CARRYB_10__40_), .S(u5_mult_87_SUMB_10__40_) );
  FA_X1 u5_mult_87_S2_10_39 ( .A(u5_mult_87_ab_10__39_), .B(
        u5_mult_87_CARRYB_9__39_), .CI(u5_mult_87_SUMB_9__40_), .CO(
        u5_mult_87_CARRYB_10__39_), .S(u5_mult_87_SUMB_10__39_) );
  FA_X1 u5_mult_87_S2_10_38 ( .A(u5_mult_87_ab_10__38_), .B(
        u5_mult_87_CARRYB_9__38_), .CI(u5_mult_87_SUMB_9__39_), .CO(
        u5_mult_87_CARRYB_10__38_), .S(u5_mult_87_SUMB_10__38_) );
  FA_X1 u5_mult_87_S2_10_37 ( .A(u5_mult_87_ab_10__37_), .B(
        u5_mult_87_CARRYB_9__37_), .CI(u5_mult_87_SUMB_9__38_), .CO(
        u5_mult_87_CARRYB_10__37_), .S(u5_mult_87_SUMB_10__37_) );
  FA_X1 u5_mult_87_S2_10_36 ( .A(u5_mult_87_ab_10__36_), .B(
        u5_mult_87_CARRYB_9__36_), .CI(u5_mult_87_SUMB_9__37_), .CO(
        u5_mult_87_CARRYB_10__36_), .S(u5_mult_87_SUMB_10__36_) );
  FA_X1 u5_mult_87_S2_10_35 ( .A(u5_mult_87_ab_10__35_), .B(
        u5_mult_87_CARRYB_9__35_), .CI(u5_mult_87_SUMB_9__36_), .CO(
        u5_mult_87_CARRYB_10__35_), .S(u5_mult_87_SUMB_10__35_) );
  FA_X1 u5_mult_87_S2_10_34 ( .A(u5_mult_87_ab_10__34_), .B(
        u5_mult_87_CARRYB_9__34_), .CI(u5_mult_87_SUMB_9__35_), .CO(
        u5_mult_87_CARRYB_10__34_), .S(u5_mult_87_SUMB_10__34_) );
  FA_X1 u5_mult_87_S2_10_33 ( .A(u5_mult_87_ab_10__33_), .B(
        u5_mult_87_CARRYB_9__33_), .CI(u5_mult_87_SUMB_9__34_), .CO(
        u5_mult_87_CARRYB_10__33_), .S(u5_mult_87_SUMB_10__33_) );
  FA_X1 u5_mult_87_S2_10_32 ( .A(u5_mult_87_ab_10__32_), .B(
        u5_mult_87_CARRYB_9__32_), .CI(u5_mult_87_SUMB_9__33_), .CO(
        u5_mult_87_CARRYB_10__32_), .S(u5_mult_87_SUMB_10__32_) );
  FA_X1 u5_mult_87_S2_10_31 ( .A(u5_mult_87_ab_10__31_), .B(
        u5_mult_87_CARRYB_9__31_), .CI(u5_mult_87_SUMB_9__32_), .CO(
        u5_mult_87_CARRYB_10__31_), .S(u5_mult_87_SUMB_10__31_) );
  FA_X1 u5_mult_87_S2_10_30 ( .A(u5_mult_87_ab_10__30_), .B(
        u5_mult_87_CARRYB_9__30_), .CI(u5_mult_87_SUMB_9__31_), .CO(
        u5_mult_87_CARRYB_10__30_), .S(u5_mult_87_SUMB_10__30_) );
  FA_X1 u5_mult_87_S2_10_29 ( .A(u5_mult_87_ab_10__29_), .B(
        u5_mult_87_CARRYB_9__29_), .CI(u5_mult_87_SUMB_9__30_), .CO(
        u5_mult_87_CARRYB_10__29_), .S(u5_mult_87_SUMB_10__29_) );
  FA_X1 u5_mult_87_S2_10_28 ( .A(u5_mult_87_ab_10__28_), .B(
        u5_mult_87_CARRYB_9__28_), .CI(u5_mult_87_SUMB_9__29_), .CO(
        u5_mult_87_CARRYB_10__28_), .S(u5_mult_87_SUMB_10__28_) );
  FA_X1 u5_mult_87_S2_10_27 ( .A(u5_mult_87_ab_10__27_), .B(
        u5_mult_87_CARRYB_9__27_), .CI(u5_mult_87_SUMB_9__28_), .CO(
        u5_mult_87_CARRYB_10__27_), .S(u5_mult_87_SUMB_10__27_) );
  FA_X1 u5_mult_87_S2_10_26 ( .A(u5_mult_87_ab_10__26_), .B(
        u5_mult_87_CARRYB_9__26_), .CI(u5_mult_87_SUMB_9__27_), .CO(
        u5_mult_87_CARRYB_10__26_), .S(u5_mult_87_SUMB_10__26_) );
  FA_X1 u5_mult_87_S2_10_25 ( .A(u5_mult_87_ab_10__25_), .B(
        u5_mult_87_CARRYB_9__25_), .CI(u5_mult_87_SUMB_9__26_), .CO(
        u5_mult_87_CARRYB_10__25_), .S(u5_mult_87_SUMB_10__25_) );
  FA_X1 u5_mult_87_S2_10_24 ( .A(u5_mult_87_ab_10__24_), .B(
        u5_mult_87_CARRYB_9__24_), .CI(u5_mult_87_SUMB_9__25_), .CO(
        u5_mult_87_CARRYB_10__24_), .S(u5_mult_87_SUMB_10__24_) );
  FA_X1 u5_mult_87_S2_10_23 ( .A(u5_mult_87_ab_10__23_), .B(
        u5_mult_87_CARRYB_9__23_), .CI(u5_mult_87_SUMB_9__24_), .CO(
        u5_mult_87_CARRYB_10__23_), .S(u5_mult_87_SUMB_10__23_) );
  FA_X1 u5_mult_87_S2_10_22 ( .A(u5_mult_87_ab_10__22_), .B(
        u5_mult_87_CARRYB_9__22_), .CI(u5_mult_87_SUMB_9__23_), .CO(
        u5_mult_87_CARRYB_10__22_), .S(u5_mult_87_SUMB_10__22_) );
  FA_X1 u5_mult_87_S2_10_21 ( .A(u5_mult_87_ab_10__21_), .B(
        u5_mult_87_CARRYB_9__21_), .CI(u5_mult_87_SUMB_9__22_), .CO(
        u5_mult_87_CARRYB_10__21_), .S(u5_mult_87_SUMB_10__21_) );
  FA_X1 u5_mult_87_S2_10_20 ( .A(u5_mult_87_ab_10__20_), .B(
        u5_mult_87_CARRYB_9__20_), .CI(u5_mult_87_SUMB_9__21_), .CO(
        u5_mult_87_CARRYB_10__20_), .S(u5_mult_87_SUMB_10__20_) );
  FA_X1 u5_mult_87_S2_10_19 ( .A(u5_mult_87_ab_10__19_), .B(
        u5_mult_87_CARRYB_9__19_), .CI(u5_mult_87_SUMB_9__20_), .CO(
        u5_mult_87_CARRYB_10__19_), .S(u5_mult_87_SUMB_10__19_) );
  FA_X1 u5_mult_87_S2_10_18 ( .A(u5_mult_87_ab_10__18_), .B(
        u5_mult_87_CARRYB_9__18_), .CI(u5_mult_87_SUMB_9__19_), .CO(
        u5_mult_87_CARRYB_10__18_), .S(u5_mult_87_SUMB_10__18_) );
  FA_X1 u5_mult_87_S2_10_17 ( .A(u5_mult_87_ab_10__17_), .B(
        u5_mult_87_CARRYB_9__17_), .CI(u5_mult_87_SUMB_9__18_), .CO(
        u5_mult_87_CARRYB_10__17_), .S(u5_mult_87_SUMB_10__17_) );
  FA_X1 u5_mult_87_S2_10_16 ( .A(u5_mult_87_ab_10__16_), .B(
        u5_mult_87_CARRYB_9__16_), .CI(u5_mult_87_SUMB_9__17_), .CO(
        u5_mult_87_CARRYB_10__16_), .S(u5_mult_87_SUMB_10__16_) );
  FA_X1 u5_mult_87_S2_10_15 ( .A(u5_mult_87_ab_10__15_), .B(
        u5_mult_87_CARRYB_9__15_), .CI(u5_mult_87_SUMB_9__16_), .CO(
        u5_mult_87_CARRYB_10__15_), .S(u5_mult_87_SUMB_10__15_) );
  FA_X1 u5_mult_87_S2_10_14 ( .A(u5_mult_87_ab_10__14_), .B(
        u5_mult_87_CARRYB_9__14_), .CI(u5_mult_87_SUMB_9__15_), .CO(
        u5_mult_87_CARRYB_10__14_), .S(u5_mult_87_SUMB_10__14_) );
  FA_X1 u5_mult_87_S2_10_13 ( .A(u5_mult_87_ab_10__13_), .B(
        u5_mult_87_CARRYB_9__13_), .CI(u5_mult_87_SUMB_9__14_), .CO(
        u5_mult_87_CARRYB_10__13_), .S(u5_mult_87_SUMB_10__13_) );
  FA_X1 u5_mult_87_S2_10_12 ( .A(u5_mult_87_ab_10__12_), .B(
        u5_mult_87_CARRYB_9__12_), .CI(u5_mult_87_SUMB_9__13_), .CO(
        u5_mult_87_CARRYB_10__12_), .S(u5_mult_87_SUMB_10__12_) );
  FA_X1 u5_mult_87_S2_10_11 ( .A(u5_mult_87_ab_10__11_), .B(
        u5_mult_87_CARRYB_9__11_), .CI(u5_mult_87_SUMB_9__12_), .CO(
        u5_mult_87_CARRYB_10__11_), .S(u5_mult_87_SUMB_10__11_) );
  FA_X1 u5_mult_87_S2_10_10 ( .A(u5_mult_87_ab_10__10_), .B(
        u5_mult_87_CARRYB_9__10_), .CI(u5_mult_87_SUMB_9__11_), .CO(
        u5_mult_87_CARRYB_10__10_), .S(u5_mult_87_SUMB_10__10_) );
  FA_X1 u5_mult_87_S2_10_9 ( .A(u5_mult_87_ab_10__9_), .B(
        u5_mult_87_CARRYB_9__9_), .CI(u5_mult_87_SUMB_9__10_), .CO(
        u5_mult_87_CARRYB_10__9_), .S(u5_mult_87_SUMB_10__9_) );
  FA_X1 u5_mult_87_S2_10_8 ( .A(u5_mult_87_ab_10__8_), .B(
        u5_mult_87_CARRYB_9__8_), .CI(u5_mult_87_SUMB_9__9_), .CO(
        u5_mult_87_CARRYB_10__8_), .S(u5_mult_87_SUMB_10__8_) );
  FA_X1 u5_mult_87_S2_10_7 ( .A(u5_mult_87_ab_10__7_), .B(
        u5_mult_87_CARRYB_9__7_), .CI(u5_mult_87_SUMB_9__8_), .CO(
        u5_mult_87_CARRYB_10__7_), .S(u5_mult_87_SUMB_10__7_) );
  FA_X1 u5_mult_87_S2_10_6 ( .A(u5_mult_87_ab_10__6_), .B(
        u5_mult_87_CARRYB_9__6_), .CI(u5_mult_87_SUMB_9__7_), .CO(
        u5_mult_87_CARRYB_10__6_), .S(u5_mult_87_SUMB_10__6_) );
  FA_X1 u5_mult_87_S2_10_5 ( .A(u5_mult_87_ab_10__5_), .B(
        u5_mult_87_CARRYB_9__5_), .CI(u5_mult_87_SUMB_9__6_), .CO(
        u5_mult_87_CARRYB_10__5_), .S(u5_mult_87_SUMB_10__5_) );
  FA_X1 u5_mult_87_S2_10_4 ( .A(u5_mult_87_ab_10__4_), .B(
        u5_mult_87_CARRYB_9__4_), .CI(u5_mult_87_SUMB_9__5_), .CO(
        u5_mult_87_CARRYB_10__4_), .S(u5_mult_87_SUMB_10__4_) );
  FA_X1 u5_mult_87_S2_10_3 ( .A(u5_mult_87_ab_10__3_), .B(
        u5_mult_87_CARRYB_9__3_), .CI(u5_mult_87_SUMB_9__4_), .CO(
        u5_mult_87_CARRYB_10__3_), .S(u5_mult_87_SUMB_10__3_) );
  FA_X1 u5_mult_87_S2_10_2 ( .A(u5_mult_87_ab_10__2_), .B(
        u5_mult_87_CARRYB_9__2_), .CI(u5_mult_87_SUMB_9__3_), .CO(
        u5_mult_87_CARRYB_10__2_), .S(u5_mult_87_SUMB_10__2_) );
  FA_X1 u5_mult_87_S2_10_1 ( .A(u5_mult_87_ab_10__1_), .B(
        u5_mult_87_CARRYB_9__1_), .CI(u5_mult_87_SUMB_9__2_), .CO(
        u5_mult_87_CARRYB_10__1_), .S(u5_mult_87_SUMB_10__1_) );
  FA_X1 u5_mult_87_S1_10_0 ( .A(u5_mult_87_ab_10__0_), .B(
        u5_mult_87_CARRYB_9__0_), .CI(u5_mult_87_SUMB_9__1_), .CO(
        u5_mult_87_CARRYB_10__0_), .S(u5_N10) );
  FA_X1 u5_mult_87_S3_11_51 ( .A(u5_mult_87_ab_11__51_), .B(
        u5_mult_87_CARRYB_10__51_), .CI(u5_mult_87_ab_10__52_), .CO(
        u5_mult_87_CARRYB_11__51_), .S(u5_mult_87_SUMB_11__51_) );
  FA_X1 u5_mult_87_S2_11_50 ( .A(u5_mult_87_ab_11__50_), .B(
        u5_mult_87_CARRYB_10__50_), .CI(u5_mult_87_SUMB_10__51_), .CO(
        u5_mult_87_CARRYB_11__50_), .S(u5_mult_87_SUMB_11__50_) );
  FA_X1 u5_mult_87_S2_11_49 ( .A(u5_mult_87_ab_11__49_), .B(
        u5_mult_87_CARRYB_10__49_), .CI(u5_mult_87_SUMB_10__50_), .CO(
        u5_mult_87_CARRYB_11__49_), .S(u5_mult_87_SUMB_11__49_) );
  FA_X1 u5_mult_87_S2_11_48 ( .A(u5_mult_87_ab_11__48_), .B(
        u5_mult_87_CARRYB_10__48_), .CI(u5_mult_87_SUMB_10__49_), .CO(
        u5_mult_87_CARRYB_11__48_), .S(u5_mult_87_SUMB_11__48_) );
  FA_X1 u5_mult_87_S2_11_47 ( .A(u5_mult_87_ab_11__47_), .B(
        u5_mult_87_CARRYB_10__47_), .CI(u5_mult_87_SUMB_10__48_), .CO(
        u5_mult_87_CARRYB_11__47_), .S(u5_mult_87_SUMB_11__47_) );
  FA_X1 u5_mult_87_S2_11_46 ( .A(u5_mult_87_ab_11__46_), .B(
        u5_mult_87_CARRYB_10__46_), .CI(u5_mult_87_SUMB_10__47_), .CO(
        u5_mult_87_CARRYB_11__46_), .S(u5_mult_87_SUMB_11__46_) );
  FA_X1 u5_mult_87_S2_11_45 ( .A(u5_mult_87_ab_11__45_), .B(
        u5_mult_87_CARRYB_10__45_), .CI(u5_mult_87_SUMB_10__46_), .CO(
        u5_mult_87_CARRYB_11__45_), .S(u5_mult_87_SUMB_11__45_) );
  FA_X1 u5_mult_87_S2_11_44 ( .A(u5_mult_87_ab_11__44_), .B(
        u5_mult_87_CARRYB_10__44_), .CI(u5_mult_87_SUMB_10__45_), .CO(
        u5_mult_87_CARRYB_11__44_), .S(u5_mult_87_SUMB_11__44_) );
  FA_X1 u5_mult_87_S2_11_43 ( .A(u5_mult_87_ab_11__43_), .B(
        u5_mult_87_CARRYB_10__43_), .CI(u5_mult_87_SUMB_10__44_), .CO(
        u5_mult_87_CARRYB_11__43_), .S(u5_mult_87_SUMB_11__43_) );
  FA_X1 u5_mult_87_S2_11_42 ( .A(u5_mult_87_ab_11__42_), .B(
        u5_mult_87_CARRYB_10__42_), .CI(u5_mult_87_SUMB_10__43_), .CO(
        u5_mult_87_CARRYB_11__42_), .S(u5_mult_87_SUMB_11__42_) );
  FA_X1 u5_mult_87_S2_11_41 ( .A(u5_mult_87_ab_11__41_), .B(
        u5_mult_87_CARRYB_10__41_), .CI(u5_mult_87_SUMB_10__42_), .CO(
        u5_mult_87_CARRYB_11__41_), .S(u5_mult_87_SUMB_11__41_) );
  FA_X1 u5_mult_87_S2_11_40 ( .A(u5_mult_87_ab_11__40_), .B(
        u5_mult_87_CARRYB_10__40_), .CI(u5_mult_87_SUMB_10__41_), .CO(
        u5_mult_87_CARRYB_11__40_), .S(u5_mult_87_SUMB_11__40_) );
  FA_X1 u5_mult_87_S2_11_39 ( .A(u5_mult_87_ab_11__39_), .B(
        u5_mult_87_CARRYB_10__39_), .CI(u5_mult_87_SUMB_10__40_), .CO(
        u5_mult_87_CARRYB_11__39_), .S(u5_mult_87_SUMB_11__39_) );
  FA_X1 u5_mult_87_S2_11_38 ( .A(u5_mult_87_ab_11__38_), .B(
        u5_mult_87_CARRYB_10__38_), .CI(u5_mult_87_SUMB_10__39_), .CO(
        u5_mult_87_CARRYB_11__38_), .S(u5_mult_87_SUMB_11__38_) );
  FA_X1 u5_mult_87_S2_11_37 ( .A(u5_mult_87_ab_11__37_), .B(
        u5_mult_87_CARRYB_10__37_), .CI(u5_mult_87_SUMB_10__38_), .CO(
        u5_mult_87_CARRYB_11__37_), .S(u5_mult_87_SUMB_11__37_) );
  FA_X1 u5_mult_87_S2_11_36 ( .A(u5_mult_87_ab_11__36_), .B(
        u5_mult_87_CARRYB_10__36_), .CI(u5_mult_87_SUMB_10__37_), .CO(
        u5_mult_87_CARRYB_11__36_), .S(u5_mult_87_SUMB_11__36_) );
  FA_X1 u5_mult_87_S2_11_35 ( .A(u5_mult_87_ab_11__35_), .B(
        u5_mult_87_CARRYB_10__35_), .CI(u5_mult_87_SUMB_10__36_), .CO(
        u5_mult_87_CARRYB_11__35_), .S(u5_mult_87_SUMB_11__35_) );
  FA_X1 u5_mult_87_S2_11_34 ( .A(u5_mult_87_ab_11__34_), .B(
        u5_mult_87_CARRYB_10__34_), .CI(u5_mult_87_SUMB_10__35_), .CO(
        u5_mult_87_CARRYB_11__34_), .S(u5_mult_87_SUMB_11__34_) );
  FA_X1 u5_mult_87_S2_11_33 ( .A(u5_mult_87_ab_11__33_), .B(
        u5_mult_87_CARRYB_10__33_), .CI(u5_mult_87_SUMB_10__34_), .CO(
        u5_mult_87_CARRYB_11__33_), .S(u5_mult_87_SUMB_11__33_) );
  FA_X1 u5_mult_87_S2_11_32 ( .A(u5_mult_87_ab_11__32_), .B(
        u5_mult_87_CARRYB_10__32_), .CI(u5_mult_87_SUMB_10__33_), .CO(
        u5_mult_87_CARRYB_11__32_), .S(u5_mult_87_SUMB_11__32_) );
  FA_X1 u5_mult_87_S2_11_31 ( .A(u5_mult_87_ab_11__31_), .B(
        u5_mult_87_CARRYB_10__31_), .CI(u5_mult_87_SUMB_10__32_), .CO(
        u5_mult_87_CARRYB_11__31_), .S(u5_mult_87_SUMB_11__31_) );
  FA_X1 u5_mult_87_S2_11_30 ( .A(u5_mult_87_ab_11__30_), .B(
        u5_mult_87_CARRYB_10__30_), .CI(u5_mult_87_SUMB_10__31_), .CO(
        u5_mult_87_CARRYB_11__30_), .S(u5_mult_87_SUMB_11__30_) );
  FA_X1 u5_mult_87_S2_11_29 ( .A(u5_mult_87_ab_11__29_), .B(
        u5_mult_87_CARRYB_10__29_), .CI(u5_mult_87_SUMB_10__30_), .CO(
        u5_mult_87_CARRYB_11__29_), .S(u5_mult_87_SUMB_11__29_) );
  FA_X1 u5_mult_87_S2_11_28 ( .A(u5_mult_87_ab_11__28_), .B(
        u5_mult_87_CARRYB_10__28_), .CI(u5_mult_87_SUMB_10__29_), .CO(
        u5_mult_87_CARRYB_11__28_), .S(u5_mult_87_SUMB_11__28_) );
  FA_X1 u5_mult_87_S2_11_27 ( .A(u5_mult_87_ab_11__27_), .B(
        u5_mult_87_CARRYB_10__27_), .CI(u5_mult_87_SUMB_10__28_), .CO(
        u5_mult_87_CARRYB_11__27_), .S(u5_mult_87_SUMB_11__27_) );
  FA_X1 u5_mult_87_S2_11_26 ( .A(u5_mult_87_ab_11__26_), .B(
        u5_mult_87_CARRYB_10__26_), .CI(u5_mult_87_SUMB_10__27_), .CO(
        u5_mult_87_CARRYB_11__26_), .S(u5_mult_87_SUMB_11__26_) );
  FA_X1 u5_mult_87_S2_11_25 ( .A(u5_mult_87_ab_11__25_), .B(
        u5_mult_87_CARRYB_10__25_), .CI(u5_mult_87_SUMB_10__26_), .CO(
        u5_mult_87_CARRYB_11__25_), .S(u5_mult_87_SUMB_11__25_) );
  FA_X1 u5_mult_87_S2_11_24 ( .A(u5_mult_87_ab_11__24_), .B(
        u5_mult_87_CARRYB_10__24_), .CI(u5_mult_87_SUMB_10__25_), .CO(
        u5_mult_87_CARRYB_11__24_), .S(u5_mult_87_SUMB_11__24_) );
  FA_X1 u5_mult_87_S2_11_23 ( .A(u5_mult_87_ab_11__23_), .B(
        u5_mult_87_CARRYB_10__23_), .CI(u5_mult_87_SUMB_10__24_), .CO(
        u5_mult_87_CARRYB_11__23_), .S(u5_mult_87_SUMB_11__23_) );
  FA_X1 u5_mult_87_S2_11_22 ( .A(u5_mult_87_ab_11__22_), .B(
        u5_mult_87_CARRYB_10__22_), .CI(u5_mult_87_SUMB_10__23_), .CO(
        u5_mult_87_CARRYB_11__22_), .S(u5_mult_87_SUMB_11__22_) );
  FA_X1 u5_mult_87_S2_11_21 ( .A(u5_mult_87_ab_11__21_), .B(
        u5_mult_87_CARRYB_10__21_), .CI(u5_mult_87_SUMB_10__22_), .CO(
        u5_mult_87_CARRYB_11__21_), .S(u5_mult_87_SUMB_11__21_) );
  FA_X1 u5_mult_87_S2_11_20 ( .A(u5_mult_87_ab_11__20_), .B(
        u5_mult_87_CARRYB_10__20_), .CI(u5_mult_87_SUMB_10__21_), .CO(
        u5_mult_87_CARRYB_11__20_), .S(u5_mult_87_SUMB_11__20_) );
  FA_X1 u5_mult_87_S2_11_19 ( .A(u5_mult_87_ab_11__19_), .B(
        u5_mult_87_CARRYB_10__19_), .CI(u5_mult_87_SUMB_10__20_), .CO(
        u5_mult_87_CARRYB_11__19_), .S(u5_mult_87_SUMB_11__19_) );
  FA_X1 u5_mult_87_S2_11_18 ( .A(u5_mult_87_ab_11__18_), .B(
        u5_mult_87_CARRYB_10__18_), .CI(u5_mult_87_SUMB_10__19_), .CO(
        u5_mult_87_CARRYB_11__18_), .S(u5_mult_87_SUMB_11__18_) );
  FA_X1 u5_mult_87_S2_11_17 ( .A(u5_mult_87_ab_11__17_), .B(
        u5_mult_87_CARRYB_10__17_), .CI(u5_mult_87_SUMB_10__18_), .CO(
        u5_mult_87_CARRYB_11__17_), .S(u5_mult_87_SUMB_11__17_) );
  FA_X1 u5_mult_87_S2_11_16 ( .A(u5_mult_87_ab_11__16_), .B(
        u5_mult_87_CARRYB_10__16_), .CI(u5_mult_87_SUMB_10__17_), .CO(
        u5_mult_87_CARRYB_11__16_), .S(u5_mult_87_SUMB_11__16_) );
  FA_X1 u5_mult_87_S2_11_15 ( .A(u5_mult_87_ab_11__15_), .B(
        u5_mult_87_CARRYB_10__15_), .CI(u5_mult_87_SUMB_10__16_), .CO(
        u5_mult_87_CARRYB_11__15_), .S(u5_mult_87_SUMB_11__15_) );
  FA_X1 u5_mult_87_S2_11_14 ( .A(u5_mult_87_ab_11__14_), .B(
        u5_mult_87_CARRYB_10__14_), .CI(u5_mult_87_SUMB_10__15_), .CO(
        u5_mult_87_CARRYB_11__14_), .S(u5_mult_87_SUMB_11__14_) );
  FA_X1 u5_mult_87_S2_11_13 ( .A(u5_mult_87_ab_11__13_), .B(
        u5_mult_87_CARRYB_10__13_), .CI(u5_mult_87_SUMB_10__14_), .CO(
        u5_mult_87_CARRYB_11__13_), .S(u5_mult_87_SUMB_11__13_) );
  FA_X1 u5_mult_87_S2_11_12 ( .A(u5_mult_87_ab_11__12_), .B(
        u5_mult_87_CARRYB_10__12_), .CI(u5_mult_87_SUMB_10__13_), .CO(
        u5_mult_87_CARRYB_11__12_), .S(u5_mult_87_SUMB_11__12_) );
  FA_X1 u5_mult_87_S2_11_11 ( .A(u5_mult_87_ab_11__11_), .B(
        u5_mult_87_CARRYB_10__11_), .CI(u5_mult_87_SUMB_10__12_), .CO(
        u5_mult_87_CARRYB_11__11_), .S(u5_mult_87_SUMB_11__11_) );
  FA_X1 u5_mult_87_S2_11_10 ( .A(u5_mult_87_ab_11__10_), .B(
        u5_mult_87_CARRYB_10__10_), .CI(u5_mult_87_SUMB_10__11_), .CO(
        u5_mult_87_CARRYB_11__10_), .S(u5_mult_87_SUMB_11__10_) );
  FA_X1 u5_mult_87_S2_11_9 ( .A(u5_mult_87_ab_11__9_), .B(
        u5_mult_87_CARRYB_10__9_), .CI(u5_mult_87_SUMB_10__10_), .CO(
        u5_mult_87_CARRYB_11__9_), .S(u5_mult_87_SUMB_11__9_) );
  FA_X1 u5_mult_87_S2_11_8 ( .A(u5_mult_87_ab_11__8_), .B(
        u5_mult_87_CARRYB_10__8_), .CI(u5_mult_87_SUMB_10__9_), .CO(
        u5_mult_87_CARRYB_11__8_), .S(u5_mult_87_SUMB_11__8_) );
  FA_X1 u5_mult_87_S2_11_7 ( .A(u5_mult_87_ab_11__7_), .B(
        u5_mult_87_CARRYB_10__7_), .CI(u5_mult_87_SUMB_10__8_), .CO(
        u5_mult_87_CARRYB_11__7_), .S(u5_mult_87_SUMB_11__7_) );
  FA_X1 u5_mult_87_S2_11_6 ( .A(u5_mult_87_ab_11__6_), .B(
        u5_mult_87_CARRYB_10__6_), .CI(u5_mult_87_SUMB_10__7_), .CO(
        u5_mult_87_CARRYB_11__6_), .S(u5_mult_87_SUMB_11__6_) );
  FA_X1 u5_mult_87_S2_11_5 ( .A(u5_mult_87_ab_11__5_), .B(
        u5_mult_87_CARRYB_10__5_), .CI(u5_mult_87_SUMB_10__6_), .CO(
        u5_mult_87_CARRYB_11__5_), .S(u5_mult_87_SUMB_11__5_) );
  FA_X1 u5_mult_87_S2_11_4 ( .A(u5_mult_87_ab_11__4_), .B(
        u5_mult_87_CARRYB_10__4_), .CI(u5_mult_87_SUMB_10__5_), .CO(
        u5_mult_87_CARRYB_11__4_), .S(u5_mult_87_SUMB_11__4_) );
  FA_X1 u5_mult_87_S2_11_3 ( .A(u5_mult_87_ab_11__3_), .B(
        u5_mult_87_CARRYB_10__3_), .CI(u5_mult_87_SUMB_10__4_), .CO(
        u5_mult_87_CARRYB_11__3_), .S(u5_mult_87_SUMB_11__3_) );
  FA_X1 u5_mult_87_S2_11_2 ( .A(u5_mult_87_ab_11__2_), .B(
        u5_mult_87_CARRYB_10__2_), .CI(u5_mult_87_SUMB_10__3_), .CO(
        u5_mult_87_CARRYB_11__2_), .S(u5_mult_87_SUMB_11__2_) );
  FA_X1 u5_mult_87_S2_11_1 ( .A(u5_mult_87_ab_11__1_), .B(
        u5_mult_87_CARRYB_10__1_), .CI(u5_mult_87_SUMB_10__2_), .CO(
        u5_mult_87_CARRYB_11__1_), .S(u5_mult_87_SUMB_11__1_) );
  FA_X1 u5_mult_87_S1_11_0 ( .A(u5_mult_87_ab_11__0_), .B(
        u5_mult_87_CARRYB_10__0_), .CI(u5_mult_87_SUMB_10__1_), .CO(
        u5_mult_87_CARRYB_11__0_), .S(u5_N11) );
  FA_X1 u5_mult_87_S3_12_51 ( .A(u5_mult_87_ab_12__51_), .B(
        u5_mult_87_CARRYB_11__51_), .CI(u5_mult_87_ab_11__52_), .CO(
        u5_mult_87_CARRYB_12__51_), .S(u5_mult_87_SUMB_12__51_) );
  FA_X1 u5_mult_87_S2_12_50 ( .A(u5_mult_87_ab_12__50_), .B(
        u5_mult_87_CARRYB_11__50_), .CI(u5_mult_87_SUMB_11__51_), .CO(
        u5_mult_87_CARRYB_12__50_), .S(u5_mult_87_SUMB_12__50_) );
  FA_X1 u5_mult_87_S2_12_49 ( .A(u5_mult_87_ab_12__49_), .B(
        u5_mult_87_CARRYB_11__49_), .CI(u5_mult_87_SUMB_11__50_), .CO(
        u5_mult_87_CARRYB_12__49_), .S(u5_mult_87_SUMB_12__49_) );
  FA_X1 u5_mult_87_S2_12_48 ( .A(u5_mult_87_ab_12__48_), .B(
        u5_mult_87_CARRYB_11__48_), .CI(u5_mult_87_SUMB_11__49_), .CO(
        u5_mult_87_CARRYB_12__48_), .S(u5_mult_87_SUMB_12__48_) );
  FA_X1 u5_mult_87_S2_12_47 ( .A(u5_mult_87_ab_12__47_), .B(
        u5_mult_87_CARRYB_11__47_), .CI(u5_mult_87_SUMB_11__48_), .CO(
        u5_mult_87_CARRYB_12__47_), .S(u5_mult_87_SUMB_12__47_) );
  FA_X1 u5_mult_87_S2_12_46 ( .A(u5_mult_87_ab_12__46_), .B(
        u5_mult_87_CARRYB_11__46_), .CI(u5_mult_87_SUMB_11__47_), .CO(
        u5_mult_87_CARRYB_12__46_), .S(u5_mult_87_SUMB_12__46_) );
  FA_X1 u5_mult_87_S2_12_45 ( .A(u5_mult_87_ab_12__45_), .B(
        u5_mult_87_CARRYB_11__45_), .CI(u5_mult_87_SUMB_11__46_), .CO(
        u5_mult_87_CARRYB_12__45_), .S(u5_mult_87_SUMB_12__45_) );
  FA_X1 u5_mult_87_S2_12_44 ( .A(u5_mult_87_ab_12__44_), .B(
        u5_mult_87_CARRYB_11__44_), .CI(u5_mult_87_SUMB_11__45_), .CO(
        u5_mult_87_CARRYB_12__44_), .S(u5_mult_87_SUMB_12__44_) );
  FA_X1 u5_mult_87_S2_12_43 ( .A(u5_mult_87_ab_12__43_), .B(
        u5_mult_87_CARRYB_11__43_), .CI(u5_mult_87_SUMB_11__44_), .CO(
        u5_mult_87_CARRYB_12__43_), .S(u5_mult_87_SUMB_12__43_) );
  FA_X1 u5_mult_87_S2_12_42 ( .A(u5_mult_87_ab_12__42_), .B(
        u5_mult_87_CARRYB_11__42_), .CI(u5_mult_87_SUMB_11__43_), .CO(
        u5_mult_87_CARRYB_12__42_), .S(u5_mult_87_SUMB_12__42_) );
  FA_X1 u5_mult_87_S2_12_41 ( .A(u5_mult_87_ab_12__41_), .B(
        u5_mult_87_CARRYB_11__41_), .CI(u5_mult_87_SUMB_11__42_), .CO(
        u5_mult_87_CARRYB_12__41_), .S(u5_mult_87_SUMB_12__41_) );
  FA_X1 u5_mult_87_S2_12_40 ( .A(u5_mult_87_ab_12__40_), .B(
        u5_mult_87_CARRYB_11__40_), .CI(u5_mult_87_SUMB_11__41_), .CO(
        u5_mult_87_CARRYB_12__40_), .S(u5_mult_87_SUMB_12__40_) );
  FA_X1 u5_mult_87_S2_12_39 ( .A(u5_mult_87_ab_12__39_), .B(
        u5_mult_87_CARRYB_11__39_), .CI(u5_mult_87_SUMB_11__40_), .CO(
        u5_mult_87_CARRYB_12__39_), .S(u5_mult_87_SUMB_12__39_) );
  FA_X1 u5_mult_87_S2_12_38 ( .A(u5_mult_87_ab_12__38_), .B(
        u5_mult_87_CARRYB_11__38_), .CI(u5_mult_87_SUMB_11__39_), .CO(
        u5_mult_87_CARRYB_12__38_), .S(u5_mult_87_SUMB_12__38_) );
  FA_X1 u5_mult_87_S2_12_37 ( .A(u5_mult_87_ab_12__37_), .B(
        u5_mult_87_CARRYB_11__37_), .CI(u5_mult_87_SUMB_11__38_), .CO(
        u5_mult_87_CARRYB_12__37_), .S(u5_mult_87_SUMB_12__37_) );
  FA_X1 u5_mult_87_S2_12_36 ( .A(u5_mult_87_ab_12__36_), .B(
        u5_mult_87_CARRYB_11__36_), .CI(u5_mult_87_SUMB_11__37_), .CO(
        u5_mult_87_CARRYB_12__36_), .S(u5_mult_87_SUMB_12__36_) );
  FA_X1 u5_mult_87_S2_12_35 ( .A(u5_mult_87_ab_12__35_), .B(
        u5_mult_87_CARRYB_11__35_), .CI(u5_mult_87_SUMB_11__36_), .CO(
        u5_mult_87_CARRYB_12__35_), .S(u5_mult_87_SUMB_12__35_) );
  FA_X1 u5_mult_87_S2_12_34 ( .A(u5_mult_87_ab_12__34_), .B(
        u5_mult_87_CARRYB_11__34_), .CI(u5_mult_87_SUMB_11__35_), .CO(
        u5_mult_87_CARRYB_12__34_), .S(u5_mult_87_SUMB_12__34_) );
  FA_X1 u5_mult_87_S2_12_33 ( .A(u5_mult_87_ab_12__33_), .B(
        u5_mult_87_CARRYB_11__33_), .CI(u5_mult_87_SUMB_11__34_), .CO(
        u5_mult_87_CARRYB_12__33_), .S(u5_mult_87_SUMB_12__33_) );
  FA_X1 u5_mult_87_S2_12_32 ( .A(u5_mult_87_ab_12__32_), .B(
        u5_mult_87_CARRYB_11__32_), .CI(u5_mult_87_SUMB_11__33_), .CO(
        u5_mult_87_CARRYB_12__32_), .S(u5_mult_87_SUMB_12__32_) );
  FA_X1 u5_mult_87_S2_12_31 ( .A(u5_mult_87_ab_12__31_), .B(
        u5_mult_87_CARRYB_11__31_), .CI(u5_mult_87_SUMB_11__32_), .CO(
        u5_mult_87_CARRYB_12__31_), .S(u5_mult_87_SUMB_12__31_) );
  FA_X1 u5_mult_87_S2_12_30 ( .A(u5_mult_87_ab_12__30_), .B(
        u5_mult_87_CARRYB_11__30_), .CI(u5_mult_87_SUMB_11__31_), .CO(
        u5_mult_87_CARRYB_12__30_), .S(u5_mult_87_SUMB_12__30_) );
  FA_X1 u5_mult_87_S2_12_29 ( .A(u5_mult_87_ab_12__29_), .B(
        u5_mult_87_CARRYB_11__29_), .CI(u5_mult_87_SUMB_11__30_), .CO(
        u5_mult_87_CARRYB_12__29_), .S(u5_mult_87_SUMB_12__29_) );
  FA_X1 u5_mult_87_S2_12_28 ( .A(u5_mult_87_ab_12__28_), .B(
        u5_mult_87_CARRYB_11__28_), .CI(u5_mult_87_SUMB_11__29_), .CO(
        u5_mult_87_CARRYB_12__28_), .S(u5_mult_87_SUMB_12__28_) );
  FA_X1 u5_mult_87_S2_12_27 ( .A(u5_mult_87_ab_12__27_), .B(
        u5_mult_87_CARRYB_11__27_), .CI(u5_mult_87_SUMB_11__28_), .CO(
        u5_mult_87_CARRYB_12__27_), .S(u5_mult_87_SUMB_12__27_) );
  FA_X1 u5_mult_87_S2_12_26 ( .A(u5_mult_87_ab_12__26_), .B(
        u5_mult_87_CARRYB_11__26_), .CI(u5_mult_87_SUMB_11__27_), .CO(
        u5_mult_87_CARRYB_12__26_), .S(u5_mult_87_SUMB_12__26_) );
  FA_X1 u5_mult_87_S2_12_25 ( .A(u5_mult_87_ab_12__25_), .B(
        u5_mult_87_CARRYB_11__25_), .CI(u5_mult_87_SUMB_11__26_), .CO(
        u5_mult_87_CARRYB_12__25_), .S(u5_mult_87_SUMB_12__25_) );
  FA_X1 u5_mult_87_S2_12_24 ( .A(u5_mult_87_ab_12__24_), .B(
        u5_mult_87_CARRYB_11__24_), .CI(u5_mult_87_SUMB_11__25_), .CO(
        u5_mult_87_CARRYB_12__24_), .S(u5_mult_87_SUMB_12__24_) );
  FA_X1 u5_mult_87_S2_12_23 ( .A(u5_mult_87_ab_12__23_), .B(
        u5_mult_87_CARRYB_11__23_), .CI(u5_mult_87_SUMB_11__24_), .CO(
        u5_mult_87_CARRYB_12__23_), .S(u5_mult_87_SUMB_12__23_) );
  FA_X1 u5_mult_87_S2_12_22 ( .A(u5_mult_87_ab_12__22_), .B(
        u5_mult_87_CARRYB_11__22_), .CI(u5_mult_87_SUMB_11__23_), .CO(
        u5_mult_87_CARRYB_12__22_), .S(u5_mult_87_SUMB_12__22_) );
  FA_X1 u5_mult_87_S2_12_21 ( .A(u5_mult_87_ab_12__21_), .B(
        u5_mult_87_CARRYB_11__21_), .CI(u5_mult_87_SUMB_11__22_), .CO(
        u5_mult_87_CARRYB_12__21_), .S(u5_mult_87_SUMB_12__21_) );
  FA_X1 u5_mult_87_S2_12_20 ( .A(u5_mult_87_ab_12__20_), .B(
        u5_mult_87_CARRYB_11__20_), .CI(u5_mult_87_SUMB_11__21_), .CO(
        u5_mult_87_CARRYB_12__20_), .S(u5_mult_87_SUMB_12__20_) );
  FA_X1 u5_mult_87_S2_12_19 ( .A(u5_mult_87_ab_12__19_), .B(
        u5_mult_87_CARRYB_11__19_), .CI(u5_mult_87_SUMB_11__20_), .CO(
        u5_mult_87_CARRYB_12__19_), .S(u5_mult_87_SUMB_12__19_) );
  FA_X1 u5_mult_87_S2_12_18 ( .A(u5_mult_87_ab_12__18_), .B(
        u5_mult_87_CARRYB_11__18_), .CI(u5_mult_87_SUMB_11__19_), .CO(
        u5_mult_87_CARRYB_12__18_), .S(u5_mult_87_SUMB_12__18_) );
  FA_X1 u5_mult_87_S2_12_17 ( .A(u5_mult_87_ab_12__17_), .B(
        u5_mult_87_CARRYB_11__17_), .CI(u5_mult_87_SUMB_11__18_), .CO(
        u5_mult_87_CARRYB_12__17_), .S(u5_mult_87_SUMB_12__17_) );
  FA_X1 u5_mult_87_S2_12_16 ( .A(u5_mult_87_ab_12__16_), .B(
        u5_mult_87_CARRYB_11__16_), .CI(u5_mult_87_SUMB_11__17_), .CO(
        u5_mult_87_CARRYB_12__16_), .S(u5_mult_87_SUMB_12__16_) );
  FA_X1 u5_mult_87_S2_12_15 ( .A(u5_mult_87_ab_12__15_), .B(
        u5_mult_87_CARRYB_11__15_), .CI(u5_mult_87_SUMB_11__16_), .CO(
        u5_mult_87_CARRYB_12__15_), .S(u5_mult_87_SUMB_12__15_) );
  FA_X1 u5_mult_87_S2_12_14 ( .A(u5_mult_87_ab_12__14_), .B(
        u5_mult_87_CARRYB_11__14_), .CI(u5_mult_87_SUMB_11__15_), .CO(
        u5_mult_87_CARRYB_12__14_), .S(u5_mult_87_SUMB_12__14_) );
  FA_X1 u5_mult_87_S2_12_13 ( .A(u5_mult_87_ab_12__13_), .B(
        u5_mult_87_CARRYB_11__13_), .CI(u5_mult_87_SUMB_11__14_), .CO(
        u5_mult_87_CARRYB_12__13_), .S(u5_mult_87_SUMB_12__13_) );
  FA_X1 u5_mult_87_S2_12_12 ( .A(u5_mult_87_ab_12__12_), .B(
        u5_mult_87_CARRYB_11__12_), .CI(u5_mult_87_SUMB_11__13_), .CO(
        u5_mult_87_CARRYB_12__12_), .S(u5_mult_87_SUMB_12__12_) );
  FA_X1 u5_mult_87_S2_12_11 ( .A(u5_mult_87_ab_12__11_), .B(
        u5_mult_87_CARRYB_11__11_), .CI(u5_mult_87_SUMB_11__12_), .CO(
        u5_mult_87_CARRYB_12__11_), .S(u5_mult_87_SUMB_12__11_) );
  FA_X1 u5_mult_87_S2_12_10 ( .A(u5_mult_87_ab_12__10_), .B(
        u5_mult_87_CARRYB_11__10_), .CI(u5_mult_87_SUMB_11__11_), .CO(
        u5_mult_87_CARRYB_12__10_), .S(u5_mult_87_SUMB_12__10_) );
  FA_X1 u5_mult_87_S2_12_9 ( .A(u5_mult_87_ab_12__9_), .B(
        u5_mult_87_CARRYB_11__9_), .CI(u5_mult_87_SUMB_11__10_), .CO(
        u5_mult_87_CARRYB_12__9_), .S(u5_mult_87_SUMB_12__9_) );
  FA_X1 u5_mult_87_S2_12_8 ( .A(u5_mult_87_ab_12__8_), .B(
        u5_mult_87_CARRYB_11__8_), .CI(u5_mult_87_SUMB_11__9_), .CO(
        u5_mult_87_CARRYB_12__8_), .S(u5_mult_87_SUMB_12__8_) );
  FA_X1 u5_mult_87_S2_12_7 ( .A(u5_mult_87_ab_12__7_), .B(
        u5_mult_87_CARRYB_11__7_), .CI(u5_mult_87_SUMB_11__8_), .CO(
        u5_mult_87_CARRYB_12__7_), .S(u5_mult_87_SUMB_12__7_) );
  FA_X1 u5_mult_87_S2_12_6 ( .A(u5_mult_87_ab_12__6_), .B(
        u5_mult_87_CARRYB_11__6_), .CI(u5_mult_87_SUMB_11__7_), .CO(
        u5_mult_87_CARRYB_12__6_), .S(u5_mult_87_SUMB_12__6_) );
  FA_X1 u5_mult_87_S2_12_5 ( .A(u5_mult_87_ab_12__5_), .B(
        u5_mult_87_CARRYB_11__5_), .CI(u5_mult_87_SUMB_11__6_), .CO(
        u5_mult_87_CARRYB_12__5_), .S(u5_mult_87_SUMB_12__5_) );
  FA_X1 u5_mult_87_S2_12_4 ( .A(u5_mult_87_ab_12__4_), .B(
        u5_mult_87_CARRYB_11__4_), .CI(u5_mult_87_SUMB_11__5_), .CO(
        u5_mult_87_CARRYB_12__4_), .S(u5_mult_87_SUMB_12__4_) );
  FA_X1 u5_mult_87_S2_12_3 ( .A(u5_mult_87_ab_12__3_), .B(
        u5_mult_87_CARRYB_11__3_), .CI(u5_mult_87_SUMB_11__4_), .CO(
        u5_mult_87_CARRYB_12__3_), .S(u5_mult_87_SUMB_12__3_) );
  FA_X1 u5_mult_87_S2_12_2 ( .A(u5_mult_87_ab_12__2_), .B(
        u5_mult_87_CARRYB_11__2_), .CI(u5_mult_87_SUMB_11__3_), .CO(
        u5_mult_87_CARRYB_12__2_), .S(u5_mult_87_SUMB_12__2_) );
  FA_X1 u5_mult_87_S2_12_1 ( .A(u5_mult_87_ab_12__1_), .B(
        u5_mult_87_CARRYB_11__1_), .CI(u5_mult_87_SUMB_11__2_), .CO(
        u5_mult_87_CARRYB_12__1_), .S(u5_mult_87_SUMB_12__1_) );
  FA_X1 u5_mult_87_S1_12_0 ( .A(u5_mult_87_ab_12__0_), .B(
        u5_mult_87_CARRYB_11__0_), .CI(u5_mult_87_SUMB_11__1_), .CO(
        u5_mult_87_CARRYB_12__0_), .S(u5_N12) );
  FA_X1 u5_mult_87_S3_13_51 ( .A(u5_mult_87_ab_13__51_), .B(
        u5_mult_87_CARRYB_12__51_), .CI(u5_mult_87_ab_12__52_), .CO(
        u5_mult_87_CARRYB_13__51_), .S(u5_mult_87_SUMB_13__51_) );
  FA_X1 u5_mult_87_S2_13_50 ( .A(u5_mult_87_ab_13__50_), .B(
        u5_mult_87_CARRYB_12__50_), .CI(u5_mult_87_SUMB_12__51_), .CO(
        u5_mult_87_CARRYB_13__50_), .S(u5_mult_87_SUMB_13__50_) );
  FA_X1 u5_mult_87_S2_13_49 ( .A(u5_mult_87_ab_13__49_), .B(
        u5_mult_87_CARRYB_12__49_), .CI(u5_mult_87_SUMB_12__50_), .CO(
        u5_mult_87_CARRYB_13__49_), .S(u5_mult_87_SUMB_13__49_) );
  FA_X1 u5_mult_87_S2_13_48 ( .A(u5_mult_87_ab_13__48_), .B(
        u5_mult_87_CARRYB_12__48_), .CI(u5_mult_87_SUMB_12__49_), .CO(
        u5_mult_87_CARRYB_13__48_), .S(u5_mult_87_SUMB_13__48_) );
  FA_X1 u5_mult_87_S2_13_47 ( .A(u5_mult_87_ab_13__47_), .B(
        u5_mult_87_CARRYB_12__47_), .CI(u5_mult_87_SUMB_12__48_), .CO(
        u5_mult_87_CARRYB_13__47_), .S(u5_mult_87_SUMB_13__47_) );
  FA_X1 u5_mult_87_S2_13_46 ( .A(u5_mult_87_ab_13__46_), .B(
        u5_mult_87_CARRYB_12__46_), .CI(u5_mult_87_SUMB_12__47_), .CO(
        u5_mult_87_CARRYB_13__46_), .S(u5_mult_87_SUMB_13__46_) );
  FA_X1 u5_mult_87_S2_13_45 ( .A(u5_mult_87_ab_13__45_), .B(
        u5_mult_87_CARRYB_12__45_), .CI(u5_mult_87_SUMB_12__46_), .CO(
        u5_mult_87_CARRYB_13__45_), .S(u5_mult_87_SUMB_13__45_) );
  FA_X1 u5_mult_87_S2_13_44 ( .A(u5_mult_87_ab_13__44_), .B(
        u5_mult_87_CARRYB_12__44_), .CI(u5_mult_87_SUMB_12__45_), .CO(
        u5_mult_87_CARRYB_13__44_), .S(u5_mult_87_SUMB_13__44_) );
  FA_X1 u5_mult_87_S2_13_43 ( .A(u5_mult_87_ab_13__43_), .B(
        u5_mult_87_CARRYB_12__43_), .CI(u5_mult_87_SUMB_12__44_), .CO(
        u5_mult_87_CARRYB_13__43_), .S(u5_mult_87_SUMB_13__43_) );
  FA_X1 u5_mult_87_S2_13_42 ( .A(u5_mult_87_ab_13__42_), .B(
        u5_mult_87_CARRYB_12__42_), .CI(u5_mult_87_SUMB_12__43_), .CO(
        u5_mult_87_CARRYB_13__42_), .S(u5_mult_87_SUMB_13__42_) );
  FA_X1 u5_mult_87_S2_13_41 ( .A(u5_mult_87_ab_13__41_), .B(
        u5_mult_87_CARRYB_12__41_), .CI(u5_mult_87_SUMB_12__42_), .CO(
        u5_mult_87_CARRYB_13__41_), .S(u5_mult_87_SUMB_13__41_) );
  FA_X1 u5_mult_87_S2_13_40 ( .A(u5_mult_87_ab_13__40_), .B(
        u5_mult_87_CARRYB_12__40_), .CI(u5_mult_87_SUMB_12__41_), .CO(
        u5_mult_87_CARRYB_13__40_), .S(u5_mult_87_SUMB_13__40_) );
  FA_X1 u5_mult_87_S2_13_39 ( .A(u5_mult_87_ab_13__39_), .B(
        u5_mult_87_CARRYB_12__39_), .CI(u5_mult_87_SUMB_12__40_), .CO(
        u5_mult_87_CARRYB_13__39_), .S(u5_mult_87_SUMB_13__39_) );
  FA_X1 u5_mult_87_S2_13_38 ( .A(u5_mult_87_ab_13__38_), .B(
        u5_mult_87_CARRYB_12__38_), .CI(u5_mult_87_SUMB_12__39_), .CO(
        u5_mult_87_CARRYB_13__38_), .S(u5_mult_87_SUMB_13__38_) );
  FA_X1 u5_mult_87_S2_13_37 ( .A(u5_mult_87_ab_13__37_), .B(
        u5_mult_87_CARRYB_12__37_), .CI(u5_mult_87_SUMB_12__38_), .CO(
        u5_mult_87_CARRYB_13__37_), .S(u5_mult_87_SUMB_13__37_) );
  FA_X1 u5_mult_87_S2_13_36 ( .A(u5_mult_87_ab_13__36_), .B(
        u5_mult_87_CARRYB_12__36_), .CI(u5_mult_87_SUMB_12__37_), .CO(
        u5_mult_87_CARRYB_13__36_), .S(u5_mult_87_SUMB_13__36_) );
  FA_X1 u5_mult_87_S2_13_35 ( .A(u5_mult_87_ab_13__35_), .B(
        u5_mult_87_CARRYB_12__35_), .CI(u5_mult_87_SUMB_12__36_), .CO(
        u5_mult_87_CARRYB_13__35_), .S(u5_mult_87_SUMB_13__35_) );
  FA_X1 u5_mult_87_S2_13_34 ( .A(u5_mult_87_ab_13__34_), .B(
        u5_mult_87_CARRYB_12__34_), .CI(u5_mult_87_SUMB_12__35_), .CO(
        u5_mult_87_CARRYB_13__34_), .S(u5_mult_87_SUMB_13__34_) );
  FA_X1 u5_mult_87_S2_13_33 ( .A(u5_mult_87_ab_13__33_), .B(
        u5_mult_87_CARRYB_12__33_), .CI(u5_mult_87_SUMB_12__34_), .CO(
        u5_mult_87_CARRYB_13__33_), .S(u5_mult_87_SUMB_13__33_) );
  FA_X1 u5_mult_87_S2_13_32 ( .A(u5_mult_87_ab_13__32_), .B(
        u5_mult_87_CARRYB_12__32_), .CI(u5_mult_87_SUMB_12__33_), .CO(
        u5_mult_87_CARRYB_13__32_), .S(u5_mult_87_SUMB_13__32_) );
  FA_X1 u5_mult_87_S2_13_31 ( .A(u5_mult_87_ab_13__31_), .B(
        u5_mult_87_CARRYB_12__31_), .CI(u5_mult_87_SUMB_12__32_), .CO(
        u5_mult_87_CARRYB_13__31_), .S(u5_mult_87_SUMB_13__31_) );
  FA_X1 u5_mult_87_S2_13_30 ( .A(u5_mult_87_ab_13__30_), .B(
        u5_mult_87_CARRYB_12__30_), .CI(u5_mult_87_SUMB_12__31_), .CO(
        u5_mult_87_CARRYB_13__30_), .S(u5_mult_87_SUMB_13__30_) );
  FA_X1 u5_mult_87_S2_13_29 ( .A(u5_mult_87_ab_13__29_), .B(
        u5_mult_87_CARRYB_12__29_), .CI(u5_mult_87_SUMB_12__30_), .CO(
        u5_mult_87_CARRYB_13__29_), .S(u5_mult_87_SUMB_13__29_) );
  FA_X1 u5_mult_87_S2_13_28 ( .A(u5_mult_87_ab_13__28_), .B(
        u5_mult_87_CARRYB_12__28_), .CI(u5_mult_87_SUMB_12__29_), .CO(
        u5_mult_87_CARRYB_13__28_), .S(u5_mult_87_SUMB_13__28_) );
  FA_X1 u5_mult_87_S2_13_27 ( .A(u5_mult_87_ab_13__27_), .B(
        u5_mult_87_CARRYB_12__27_), .CI(u5_mult_87_SUMB_12__28_), .CO(
        u5_mult_87_CARRYB_13__27_), .S(u5_mult_87_SUMB_13__27_) );
  FA_X1 u5_mult_87_S2_13_26 ( .A(u5_mult_87_ab_13__26_), .B(
        u5_mult_87_CARRYB_12__26_), .CI(u5_mult_87_SUMB_12__27_), .CO(
        u5_mult_87_CARRYB_13__26_), .S(u5_mult_87_SUMB_13__26_) );
  FA_X1 u5_mult_87_S2_13_25 ( .A(u5_mult_87_ab_13__25_), .B(
        u5_mult_87_CARRYB_12__25_), .CI(u5_mult_87_SUMB_12__26_), .CO(
        u5_mult_87_CARRYB_13__25_), .S(u5_mult_87_SUMB_13__25_) );
  FA_X1 u5_mult_87_S2_13_24 ( .A(u5_mult_87_ab_13__24_), .B(
        u5_mult_87_CARRYB_12__24_), .CI(u5_mult_87_SUMB_12__25_), .CO(
        u5_mult_87_CARRYB_13__24_), .S(u5_mult_87_SUMB_13__24_) );
  FA_X1 u5_mult_87_S2_13_23 ( .A(u5_mult_87_ab_13__23_), .B(
        u5_mult_87_CARRYB_12__23_), .CI(u5_mult_87_SUMB_12__24_), .CO(
        u5_mult_87_CARRYB_13__23_), .S(u5_mult_87_SUMB_13__23_) );
  FA_X1 u5_mult_87_S2_13_22 ( .A(u5_mult_87_ab_13__22_), .B(
        u5_mult_87_CARRYB_12__22_), .CI(u5_mult_87_SUMB_12__23_), .CO(
        u5_mult_87_CARRYB_13__22_), .S(u5_mult_87_SUMB_13__22_) );
  FA_X1 u5_mult_87_S2_13_21 ( .A(u5_mult_87_ab_13__21_), .B(
        u5_mult_87_CARRYB_12__21_), .CI(u5_mult_87_SUMB_12__22_), .CO(
        u5_mult_87_CARRYB_13__21_), .S(u5_mult_87_SUMB_13__21_) );
  FA_X1 u5_mult_87_S2_13_20 ( .A(u5_mult_87_ab_13__20_), .B(
        u5_mult_87_CARRYB_12__20_), .CI(u5_mult_87_SUMB_12__21_), .CO(
        u5_mult_87_CARRYB_13__20_), .S(u5_mult_87_SUMB_13__20_) );
  FA_X1 u5_mult_87_S2_13_19 ( .A(u5_mult_87_ab_13__19_), .B(
        u5_mult_87_CARRYB_12__19_), .CI(u5_mult_87_SUMB_12__20_), .CO(
        u5_mult_87_CARRYB_13__19_), .S(u5_mult_87_SUMB_13__19_) );
  FA_X1 u5_mult_87_S2_13_18 ( .A(u5_mult_87_ab_13__18_), .B(
        u5_mult_87_CARRYB_12__18_), .CI(u5_mult_87_SUMB_12__19_), .CO(
        u5_mult_87_CARRYB_13__18_), .S(u5_mult_87_SUMB_13__18_) );
  FA_X1 u5_mult_87_S2_13_17 ( .A(u5_mult_87_ab_13__17_), .B(
        u5_mult_87_CARRYB_12__17_), .CI(u5_mult_87_SUMB_12__18_), .CO(
        u5_mult_87_CARRYB_13__17_), .S(u5_mult_87_SUMB_13__17_) );
  FA_X1 u5_mult_87_S2_13_16 ( .A(u5_mult_87_ab_13__16_), .B(
        u5_mult_87_CARRYB_12__16_), .CI(u5_mult_87_SUMB_12__17_), .CO(
        u5_mult_87_CARRYB_13__16_), .S(u5_mult_87_SUMB_13__16_) );
  FA_X1 u5_mult_87_S2_13_15 ( .A(u5_mult_87_ab_13__15_), .B(
        u5_mult_87_CARRYB_12__15_), .CI(u5_mult_87_SUMB_12__16_), .CO(
        u5_mult_87_CARRYB_13__15_), .S(u5_mult_87_SUMB_13__15_) );
  FA_X1 u5_mult_87_S2_13_14 ( .A(u5_mult_87_ab_13__14_), .B(
        u5_mult_87_CARRYB_12__14_), .CI(u5_mult_87_SUMB_12__15_), .CO(
        u5_mult_87_CARRYB_13__14_), .S(u5_mult_87_SUMB_13__14_) );
  FA_X1 u5_mult_87_S2_13_13 ( .A(u5_mult_87_ab_13__13_), .B(
        u5_mult_87_CARRYB_12__13_), .CI(u5_mult_87_SUMB_12__14_), .CO(
        u5_mult_87_CARRYB_13__13_), .S(u5_mult_87_SUMB_13__13_) );
  FA_X1 u5_mult_87_S2_13_12 ( .A(u5_mult_87_ab_13__12_), .B(
        u5_mult_87_CARRYB_12__12_), .CI(u5_mult_87_SUMB_12__13_), .CO(
        u5_mult_87_CARRYB_13__12_), .S(u5_mult_87_SUMB_13__12_) );
  FA_X1 u5_mult_87_S2_13_11 ( .A(u5_mult_87_ab_13__11_), .B(
        u5_mult_87_CARRYB_12__11_), .CI(u5_mult_87_SUMB_12__12_), .CO(
        u5_mult_87_CARRYB_13__11_), .S(u5_mult_87_SUMB_13__11_) );
  FA_X1 u5_mult_87_S2_13_10 ( .A(u5_mult_87_ab_13__10_), .B(
        u5_mult_87_CARRYB_12__10_), .CI(u5_mult_87_SUMB_12__11_), .CO(
        u5_mult_87_CARRYB_13__10_), .S(u5_mult_87_SUMB_13__10_) );
  FA_X1 u5_mult_87_S2_13_9 ( .A(u5_mult_87_ab_13__9_), .B(
        u5_mult_87_CARRYB_12__9_), .CI(u5_mult_87_SUMB_12__10_), .CO(
        u5_mult_87_CARRYB_13__9_), .S(u5_mult_87_SUMB_13__9_) );
  FA_X1 u5_mult_87_S2_13_8 ( .A(u5_mult_87_ab_13__8_), .B(
        u5_mult_87_CARRYB_12__8_), .CI(u5_mult_87_SUMB_12__9_), .CO(
        u5_mult_87_CARRYB_13__8_), .S(u5_mult_87_SUMB_13__8_) );
  FA_X1 u5_mult_87_S2_13_7 ( .A(u5_mult_87_ab_13__7_), .B(
        u5_mult_87_CARRYB_12__7_), .CI(u5_mult_87_SUMB_12__8_), .CO(
        u5_mult_87_CARRYB_13__7_), .S(u5_mult_87_SUMB_13__7_) );
  FA_X1 u5_mult_87_S2_13_6 ( .A(u5_mult_87_ab_13__6_), .B(
        u5_mult_87_CARRYB_12__6_), .CI(u5_mult_87_SUMB_12__7_), .CO(
        u5_mult_87_CARRYB_13__6_), .S(u5_mult_87_SUMB_13__6_) );
  FA_X1 u5_mult_87_S2_13_5 ( .A(u5_mult_87_ab_13__5_), .B(
        u5_mult_87_CARRYB_12__5_), .CI(u5_mult_87_SUMB_12__6_), .CO(
        u5_mult_87_CARRYB_13__5_), .S(u5_mult_87_SUMB_13__5_) );
  FA_X1 u5_mult_87_S2_13_4 ( .A(u5_mult_87_ab_13__4_), .B(
        u5_mult_87_CARRYB_12__4_), .CI(u5_mult_87_SUMB_12__5_), .CO(
        u5_mult_87_CARRYB_13__4_), .S(u5_mult_87_SUMB_13__4_) );
  FA_X1 u5_mult_87_S2_13_3 ( .A(u5_mult_87_ab_13__3_), .B(
        u5_mult_87_CARRYB_12__3_), .CI(u5_mult_87_SUMB_12__4_), .CO(
        u5_mult_87_CARRYB_13__3_), .S(u5_mult_87_SUMB_13__3_) );
  FA_X1 u5_mult_87_S2_13_2 ( .A(u5_mult_87_ab_13__2_), .B(
        u5_mult_87_CARRYB_12__2_), .CI(u5_mult_87_SUMB_12__3_), .CO(
        u5_mult_87_CARRYB_13__2_), .S(u5_mult_87_SUMB_13__2_) );
  FA_X1 u5_mult_87_S2_13_1 ( .A(u5_mult_87_ab_13__1_), .B(
        u5_mult_87_CARRYB_12__1_), .CI(u5_mult_87_SUMB_12__2_), .CO(
        u5_mult_87_CARRYB_13__1_), .S(u5_mult_87_SUMB_13__1_) );
  FA_X1 u5_mult_87_S1_13_0 ( .A(u5_mult_87_ab_13__0_), .B(
        u5_mult_87_CARRYB_12__0_), .CI(u5_mult_87_SUMB_12__1_), .CO(
        u5_mult_87_CARRYB_13__0_), .S(u5_N13) );
  FA_X1 u5_mult_87_S3_14_51 ( .A(u5_mult_87_ab_14__51_), .B(
        u5_mult_87_CARRYB_13__51_), .CI(u5_mult_87_ab_13__52_), .CO(
        u5_mult_87_CARRYB_14__51_), .S(u5_mult_87_SUMB_14__51_) );
  FA_X1 u5_mult_87_S2_14_50 ( .A(u5_mult_87_ab_14__50_), .B(
        u5_mult_87_CARRYB_13__50_), .CI(u5_mult_87_SUMB_13__51_), .CO(
        u5_mult_87_CARRYB_14__50_), .S(u5_mult_87_SUMB_14__50_) );
  FA_X1 u5_mult_87_S2_14_49 ( .A(u5_mult_87_ab_14__49_), .B(
        u5_mult_87_CARRYB_13__49_), .CI(u5_mult_87_SUMB_13__50_), .CO(
        u5_mult_87_CARRYB_14__49_), .S(u5_mult_87_SUMB_14__49_) );
  FA_X1 u5_mult_87_S2_14_48 ( .A(u5_mult_87_ab_14__48_), .B(
        u5_mult_87_CARRYB_13__48_), .CI(u5_mult_87_SUMB_13__49_), .CO(
        u5_mult_87_CARRYB_14__48_), .S(u5_mult_87_SUMB_14__48_) );
  FA_X1 u5_mult_87_S2_14_47 ( .A(u5_mult_87_ab_14__47_), .B(
        u5_mult_87_CARRYB_13__47_), .CI(u5_mult_87_SUMB_13__48_), .CO(
        u5_mult_87_CARRYB_14__47_), .S(u5_mult_87_SUMB_14__47_) );
  FA_X1 u5_mult_87_S2_14_46 ( .A(u5_mult_87_ab_14__46_), .B(
        u5_mult_87_CARRYB_13__46_), .CI(u5_mult_87_SUMB_13__47_), .CO(
        u5_mult_87_CARRYB_14__46_), .S(u5_mult_87_SUMB_14__46_) );
  FA_X1 u5_mult_87_S2_14_45 ( .A(u5_mult_87_ab_14__45_), .B(
        u5_mult_87_CARRYB_13__45_), .CI(u5_mult_87_SUMB_13__46_), .CO(
        u5_mult_87_CARRYB_14__45_), .S(u5_mult_87_SUMB_14__45_) );
  FA_X1 u5_mult_87_S2_14_44 ( .A(u5_mult_87_ab_14__44_), .B(
        u5_mult_87_CARRYB_13__44_), .CI(u5_mult_87_SUMB_13__45_), .CO(
        u5_mult_87_CARRYB_14__44_), .S(u5_mult_87_SUMB_14__44_) );
  FA_X1 u5_mult_87_S2_14_43 ( .A(u5_mult_87_ab_14__43_), .B(
        u5_mult_87_CARRYB_13__43_), .CI(u5_mult_87_SUMB_13__44_), .CO(
        u5_mult_87_CARRYB_14__43_), .S(u5_mult_87_SUMB_14__43_) );
  FA_X1 u5_mult_87_S2_14_42 ( .A(u5_mult_87_ab_14__42_), .B(
        u5_mult_87_CARRYB_13__42_), .CI(u5_mult_87_SUMB_13__43_), .CO(
        u5_mult_87_CARRYB_14__42_), .S(u5_mult_87_SUMB_14__42_) );
  FA_X1 u5_mult_87_S2_14_41 ( .A(u5_mult_87_ab_14__41_), .B(
        u5_mult_87_CARRYB_13__41_), .CI(u5_mult_87_SUMB_13__42_), .CO(
        u5_mult_87_CARRYB_14__41_), .S(u5_mult_87_SUMB_14__41_) );
  FA_X1 u5_mult_87_S2_14_40 ( .A(u5_mult_87_ab_14__40_), .B(
        u5_mult_87_CARRYB_13__40_), .CI(u5_mult_87_SUMB_13__41_), .CO(
        u5_mult_87_CARRYB_14__40_), .S(u5_mult_87_SUMB_14__40_) );
  FA_X1 u5_mult_87_S2_14_39 ( .A(u5_mult_87_ab_14__39_), .B(
        u5_mult_87_CARRYB_13__39_), .CI(u5_mult_87_SUMB_13__40_), .CO(
        u5_mult_87_CARRYB_14__39_), .S(u5_mult_87_SUMB_14__39_) );
  FA_X1 u5_mult_87_S2_14_38 ( .A(u5_mult_87_ab_14__38_), .B(
        u5_mult_87_CARRYB_13__38_), .CI(u5_mult_87_SUMB_13__39_), .CO(
        u5_mult_87_CARRYB_14__38_), .S(u5_mult_87_SUMB_14__38_) );
  FA_X1 u5_mult_87_S2_14_37 ( .A(u5_mult_87_ab_14__37_), .B(
        u5_mult_87_CARRYB_13__37_), .CI(u5_mult_87_SUMB_13__38_), .CO(
        u5_mult_87_CARRYB_14__37_), .S(u5_mult_87_SUMB_14__37_) );
  FA_X1 u5_mult_87_S2_14_36 ( .A(u5_mult_87_ab_14__36_), .B(
        u5_mult_87_CARRYB_13__36_), .CI(u5_mult_87_SUMB_13__37_), .CO(
        u5_mult_87_CARRYB_14__36_), .S(u5_mult_87_SUMB_14__36_) );
  FA_X1 u5_mult_87_S2_14_35 ( .A(u5_mult_87_ab_14__35_), .B(
        u5_mult_87_CARRYB_13__35_), .CI(u5_mult_87_SUMB_13__36_), .CO(
        u5_mult_87_CARRYB_14__35_), .S(u5_mult_87_SUMB_14__35_) );
  FA_X1 u5_mult_87_S2_14_34 ( .A(u5_mult_87_ab_14__34_), .B(
        u5_mult_87_CARRYB_13__34_), .CI(u5_mult_87_SUMB_13__35_), .CO(
        u5_mult_87_CARRYB_14__34_), .S(u5_mult_87_SUMB_14__34_) );
  FA_X1 u5_mult_87_S2_14_33 ( .A(u5_mult_87_ab_14__33_), .B(
        u5_mult_87_CARRYB_13__33_), .CI(u5_mult_87_SUMB_13__34_), .CO(
        u5_mult_87_CARRYB_14__33_), .S(u5_mult_87_SUMB_14__33_) );
  FA_X1 u5_mult_87_S2_14_32 ( .A(u5_mult_87_ab_14__32_), .B(
        u5_mult_87_CARRYB_13__32_), .CI(u5_mult_87_SUMB_13__33_), .CO(
        u5_mult_87_CARRYB_14__32_), .S(u5_mult_87_SUMB_14__32_) );
  FA_X1 u5_mult_87_S2_14_31 ( .A(u5_mult_87_ab_14__31_), .B(
        u5_mult_87_CARRYB_13__31_), .CI(u5_mult_87_SUMB_13__32_), .CO(
        u5_mult_87_CARRYB_14__31_), .S(u5_mult_87_SUMB_14__31_) );
  FA_X1 u5_mult_87_S2_14_30 ( .A(u5_mult_87_ab_14__30_), .B(
        u5_mult_87_CARRYB_13__30_), .CI(u5_mult_87_SUMB_13__31_), .CO(
        u5_mult_87_CARRYB_14__30_), .S(u5_mult_87_SUMB_14__30_) );
  FA_X1 u5_mult_87_S2_14_29 ( .A(u5_mult_87_ab_14__29_), .B(
        u5_mult_87_CARRYB_13__29_), .CI(u5_mult_87_SUMB_13__30_), .CO(
        u5_mult_87_CARRYB_14__29_), .S(u5_mult_87_SUMB_14__29_) );
  FA_X1 u5_mult_87_S2_14_28 ( .A(u5_mult_87_ab_14__28_), .B(
        u5_mult_87_CARRYB_13__28_), .CI(u5_mult_87_SUMB_13__29_), .CO(
        u5_mult_87_CARRYB_14__28_), .S(u5_mult_87_SUMB_14__28_) );
  FA_X1 u5_mult_87_S2_14_27 ( .A(u5_mult_87_ab_14__27_), .B(
        u5_mult_87_CARRYB_13__27_), .CI(u5_mult_87_SUMB_13__28_), .CO(
        u5_mult_87_CARRYB_14__27_), .S(u5_mult_87_SUMB_14__27_) );
  FA_X1 u5_mult_87_S2_14_26 ( .A(u5_mult_87_ab_14__26_), .B(
        u5_mult_87_CARRYB_13__26_), .CI(u5_mult_87_SUMB_13__27_), .CO(
        u5_mult_87_CARRYB_14__26_), .S(u5_mult_87_SUMB_14__26_) );
  FA_X1 u5_mult_87_S2_14_25 ( .A(u5_mult_87_ab_14__25_), .B(
        u5_mult_87_CARRYB_13__25_), .CI(u5_mult_87_SUMB_13__26_), .CO(
        u5_mult_87_CARRYB_14__25_), .S(u5_mult_87_SUMB_14__25_) );
  FA_X1 u5_mult_87_S2_14_24 ( .A(u5_mult_87_ab_14__24_), .B(
        u5_mult_87_CARRYB_13__24_), .CI(u5_mult_87_SUMB_13__25_), .CO(
        u5_mult_87_CARRYB_14__24_), .S(u5_mult_87_SUMB_14__24_) );
  FA_X1 u5_mult_87_S2_14_23 ( .A(u5_mult_87_ab_14__23_), .B(
        u5_mult_87_CARRYB_13__23_), .CI(u5_mult_87_SUMB_13__24_), .CO(
        u5_mult_87_CARRYB_14__23_), .S(u5_mult_87_SUMB_14__23_) );
  FA_X1 u5_mult_87_S2_14_22 ( .A(u5_mult_87_ab_14__22_), .B(
        u5_mult_87_CARRYB_13__22_), .CI(u5_mult_87_SUMB_13__23_), .CO(
        u5_mult_87_CARRYB_14__22_), .S(u5_mult_87_SUMB_14__22_) );
  FA_X1 u5_mult_87_S2_14_21 ( .A(u5_mult_87_ab_14__21_), .B(
        u5_mult_87_CARRYB_13__21_), .CI(u5_mult_87_SUMB_13__22_), .CO(
        u5_mult_87_CARRYB_14__21_), .S(u5_mult_87_SUMB_14__21_) );
  FA_X1 u5_mult_87_S2_14_20 ( .A(u5_mult_87_ab_14__20_), .B(
        u5_mult_87_CARRYB_13__20_), .CI(u5_mult_87_SUMB_13__21_), .CO(
        u5_mult_87_CARRYB_14__20_), .S(u5_mult_87_SUMB_14__20_) );
  FA_X1 u5_mult_87_S2_14_19 ( .A(u5_mult_87_ab_14__19_), .B(
        u5_mult_87_CARRYB_13__19_), .CI(u5_mult_87_SUMB_13__20_), .CO(
        u5_mult_87_CARRYB_14__19_), .S(u5_mult_87_SUMB_14__19_) );
  FA_X1 u5_mult_87_S2_14_18 ( .A(u5_mult_87_ab_14__18_), .B(
        u5_mult_87_CARRYB_13__18_), .CI(u5_mult_87_SUMB_13__19_), .CO(
        u5_mult_87_CARRYB_14__18_), .S(u5_mult_87_SUMB_14__18_) );
  FA_X1 u5_mult_87_S2_14_17 ( .A(u5_mult_87_ab_14__17_), .B(
        u5_mult_87_CARRYB_13__17_), .CI(u5_mult_87_SUMB_13__18_), .CO(
        u5_mult_87_CARRYB_14__17_), .S(u5_mult_87_SUMB_14__17_) );
  FA_X1 u5_mult_87_S2_14_16 ( .A(u5_mult_87_ab_14__16_), .B(
        u5_mult_87_CARRYB_13__16_), .CI(u5_mult_87_SUMB_13__17_), .CO(
        u5_mult_87_CARRYB_14__16_), .S(u5_mult_87_SUMB_14__16_) );
  FA_X1 u5_mult_87_S2_14_15 ( .A(u5_mult_87_ab_14__15_), .B(
        u5_mult_87_CARRYB_13__15_), .CI(u5_mult_87_SUMB_13__16_), .CO(
        u5_mult_87_CARRYB_14__15_), .S(u5_mult_87_SUMB_14__15_) );
  FA_X1 u5_mult_87_S2_14_14 ( .A(u5_mult_87_ab_14__14_), .B(
        u5_mult_87_CARRYB_13__14_), .CI(u5_mult_87_SUMB_13__15_), .CO(
        u5_mult_87_CARRYB_14__14_), .S(u5_mult_87_SUMB_14__14_) );
  FA_X1 u5_mult_87_S2_14_13 ( .A(u5_mult_87_ab_14__13_), .B(
        u5_mult_87_CARRYB_13__13_), .CI(u5_mult_87_SUMB_13__14_), .CO(
        u5_mult_87_CARRYB_14__13_), .S(u5_mult_87_SUMB_14__13_) );
  FA_X1 u5_mult_87_S2_14_12 ( .A(u5_mult_87_ab_14__12_), .B(
        u5_mult_87_CARRYB_13__12_), .CI(u5_mult_87_SUMB_13__13_), .CO(
        u5_mult_87_CARRYB_14__12_), .S(u5_mult_87_SUMB_14__12_) );
  FA_X1 u5_mult_87_S2_14_11 ( .A(u5_mult_87_ab_14__11_), .B(
        u5_mult_87_CARRYB_13__11_), .CI(u5_mult_87_SUMB_13__12_), .CO(
        u5_mult_87_CARRYB_14__11_), .S(u5_mult_87_SUMB_14__11_) );
  FA_X1 u5_mult_87_S2_14_10 ( .A(u5_mult_87_ab_14__10_), .B(
        u5_mult_87_CARRYB_13__10_), .CI(u5_mult_87_SUMB_13__11_), .CO(
        u5_mult_87_CARRYB_14__10_), .S(u5_mult_87_SUMB_14__10_) );
  FA_X1 u5_mult_87_S2_14_9 ( .A(u5_mult_87_ab_14__9_), .B(
        u5_mult_87_CARRYB_13__9_), .CI(u5_mult_87_SUMB_13__10_), .CO(
        u5_mult_87_CARRYB_14__9_), .S(u5_mult_87_SUMB_14__9_) );
  FA_X1 u5_mult_87_S2_14_8 ( .A(u5_mult_87_ab_14__8_), .B(
        u5_mult_87_CARRYB_13__8_), .CI(u5_mult_87_SUMB_13__9_), .CO(
        u5_mult_87_CARRYB_14__8_), .S(u5_mult_87_SUMB_14__8_) );
  FA_X1 u5_mult_87_S2_14_7 ( .A(u5_mult_87_ab_14__7_), .B(
        u5_mult_87_CARRYB_13__7_), .CI(u5_mult_87_SUMB_13__8_), .CO(
        u5_mult_87_CARRYB_14__7_), .S(u5_mult_87_SUMB_14__7_) );
  FA_X1 u5_mult_87_S2_14_6 ( .A(u5_mult_87_ab_14__6_), .B(
        u5_mult_87_CARRYB_13__6_), .CI(u5_mult_87_SUMB_13__7_), .CO(
        u5_mult_87_CARRYB_14__6_), .S(u5_mult_87_SUMB_14__6_) );
  FA_X1 u5_mult_87_S2_14_5 ( .A(u5_mult_87_ab_14__5_), .B(
        u5_mult_87_CARRYB_13__5_), .CI(u5_mult_87_SUMB_13__6_), .CO(
        u5_mult_87_CARRYB_14__5_), .S(u5_mult_87_SUMB_14__5_) );
  FA_X1 u5_mult_87_S2_14_4 ( .A(u5_mult_87_ab_14__4_), .B(
        u5_mult_87_CARRYB_13__4_), .CI(u5_mult_87_SUMB_13__5_), .CO(
        u5_mult_87_CARRYB_14__4_), .S(u5_mult_87_SUMB_14__4_) );
  FA_X1 u5_mult_87_S2_14_3 ( .A(u5_mult_87_ab_14__3_), .B(
        u5_mult_87_CARRYB_13__3_), .CI(u5_mult_87_SUMB_13__4_), .CO(
        u5_mult_87_CARRYB_14__3_), .S(u5_mult_87_SUMB_14__3_) );
  FA_X1 u5_mult_87_S2_14_2 ( .A(u5_mult_87_ab_14__2_), .B(
        u5_mult_87_CARRYB_13__2_), .CI(u5_mult_87_SUMB_13__3_), .CO(
        u5_mult_87_CARRYB_14__2_), .S(u5_mult_87_SUMB_14__2_) );
  FA_X1 u5_mult_87_S2_14_1 ( .A(u5_mult_87_ab_14__1_), .B(
        u5_mult_87_CARRYB_13__1_), .CI(u5_mult_87_SUMB_13__2_), .CO(
        u5_mult_87_CARRYB_14__1_), .S(u5_mult_87_SUMB_14__1_) );
  FA_X1 u5_mult_87_S1_14_0 ( .A(u5_mult_87_ab_14__0_), .B(
        u5_mult_87_CARRYB_13__0_), .CI(u5_mult_87_SUMB_13__1_), .CO(
        u5_mult_87_CARRYB_14__0_), .S(u5_N14) );
  FA_X1 u5_mult_87_S3_15_51 ( .A(u5_mult_87_ab_15__51_), .B(
        u5_mult_87_CARRYB_14__51_), .CI(u5_mult_87_ab_14__52_), .CO(
        u5_mult_87_CARRYB_15__51_), .S(u5_mult_87_SUMB_15__51_) );
  FA_X1 u5_mult_87_S2_15_50 ( .A(u5_mult_87_ab_15__50_), .B(
        u5_mult_87_CARRYB_14__50_), .CI(u5_mult_87_SUMB_14__51_), .CO(
        u5_mult_87_CARRYB_15__50_), .S(u5_mult_87_SUMB_15__50_) );
  FA_X1 u5_mult_87_S2_15_49 ( .A(u5_mult_87_ab_15__49_), .B(
        u5_mult_87_CARRYB_14__49_), .CI(u5_mult_87_SUMB_14__50_), .CO(
        u5_mult_87_CARRYB_15__49_), .S(u5_mult_87_SUMB_15__49_) );
  FA_X1 u5_mult_87_S2_15_48 ( .A(u5_mult_87_ab_15__48_), .B(
        u5_mult_87_CARRYB_14__48_), .CI(u5_mult_87_SUMB_14__49_), .CO(
        u5_mult_87_CARRYB_15__48_), .S(u5_mult_87_SUMB_15__48_) );
  FA_X1 u5_mult_87_S2_15_47 ( .A(u5_mult_87_ab_15__47_), .B(
        u5_mult_87_CARRYB_14__47_), .CI(u5_mult_87_SUMB_14__48_), .CO(
        u5_mult_87_CARRYB_15__47_), .S(u5_mult_87_SUMB_15__47_) );
  FA_X1 u5_mult_87_S2_15_46 ( .A(u5_mult_87_ab_15__46_), .B(
        u5_mult_87_CARRYB_14__46_), .CI(u5_mult_87_SUMB_14__47_), .CO(
        u5_mult_87_CARRYB_15__46_), .S(u5_mult_87_SUMB_15__46_) );
  FA_X1 u5_mult_87_S2_15_45 ( .A(u5_mult_87_ab_15__45_), .B(
        u5_mult_87_CARRYB_14__45_), .CI(u5_mult_87_SUMB_14__46_), .CO(
        u5_mult_87_CARRYB_15__45_), .S(u5_mult_87_SUMB_15__45_) );
  FA_X1 u5_mult_87_S2_15_44 ( .A(u5_mult_87_ab_15__44_), .B(
        u5_mult_87_CARRYB_14__44_), .CI(u5_mult_87_SUMB_14__45_), .CO(
        u5_mult_87_CARRYB_15__44_), .S(u5_mult_87_SUMB_15__44_) );
  FA_X1 u5_mult_87_S2_15_43 ( .A(u5_mult_87_ab_15__43_), .B(
        u5_mult_87_CARRYB_14__43_), .CI(u5_mult_87_SUMB_14__44_), .CO(
        u5_mult_87_CARRYB_15__43_), .S(u5_mult_87_SUMB_15__43_) );
  FA_X1 u5_mult_87_S2_15_42 ( .A(u5_mult_87_ab_15__42_), .B(
        u5_mult_87_CARRYB_14__42_), .CI(u5_mult_87_SUMB_14__43_), .CO(
        u5_mult_87_CARRYB_15__42_), .S(u5_mult_87_SUMB_15__42_) );
  FA_X1 u5_mult_87_S2_15_41 ( .A(u5_mult_87_ab_15__41_), .B(
        u5_mult_87_CARRYB_14__41_), .CI(u5_mult_87_SUMB_14__42_), .CO(
        u5_mult_87_CARRYB_15__41_), .S(u5_mult_87_SUMB_15__41_) );
  FA_X1 u5_mult_87_S2_15_40 ( .A(u5_mult_87_ab_15__40_), .B(
        u5_mult_87_CARRYB_14__40_), .CI(u5_mult_87_SUMB_14__41_), .CO(
        u5_mult_87_CARRYB_15__40_), .S(u5_mult_87_SUMB_15__40_) );
  FA_X1 u5_mult_87_S2_15_39 ( .A(u5_mult_87_ab_15__39_), .B(
        u5_mult_87_CARRYB_14__39_), .CI(u5_mult_87_SUMB_14__40_), .CO(
        u5_mult_87_CARRYB_15__39_), .S(u5_mult_87_SUMB_15__39_) );
  FA_X1 u5_mult_87_S2_15_38 ( .A(u5_mult_87_ab_15__38_), .B(
        u5_mult_87_CARRYB_14__38_), .CI(u5_mult_87_SUMB_14__39_), .CO(
        u5_mult_87_CARRYB_15__38_), .S(u5_mult_87_SUMB_15__38_) );
  FA_X1 u5_mult_87_S2_15_37 ( .A(u5_mult_87_ab_15__37_), .B(
        u5_mult_87_CARRYB_14__37_), .CI(u5_mult_87_SUMB_14__38_), .CO(
        u5_mult_87_CARRYB_15__37_), .S(u5_mult_87_SUMB_15__37_) );
  FA_X1 u5_mult_87_S2_15_36 ( .A(u5_mult_87_ab_15__36_), .B(
        u5_mult_87_CARRYB_14__36_), .CI(u5_mult_87_SUMB_14__37_), .CO(
        u5_mult_87_CARRYB_15__36_), .S(u5_mult_87_SUMB_15__36_) );
  FA_X1 u5_mult_87_S2_15_35 ( .A(u5_mult_87_ab_15__35_), .B(
        u5_mult_87_CARRYB_14__35_), .CI(u5_mult_87_SUMB_14__36_), .CO(
        u5_mult_87_CARRYB_15__35_), .S(u5_mult_87_SUMB_15__35_) );
  FA_X1 u5_mult_87_S2_15_34 ( .A(u5_mult_87_ab_15__34_), .B(
        u5_mult_87_CARRYB_14__34_), .CI(u5_mult_87_SUMB_14__35_), .CO(
        u5_mult_87_CARRYB_15__34_), .S(u5_mult_87_SUMB_15__34_) );
  FA_X1 u5_mult_87_S2_15_33 ( .A(u5_mult_87_ab_15__33_), .B(
        u5_mult_87_CARRYB_14__33_), .CI(u5_mult_87_SUMB_14__34_), .CO(
        u5_mult_87_CARRYB_15__33_), .S(u5_mult_87_SUMB_15__33_) );
  FA_X1 u5_mult_87_S2_15_32 ( .A(u5_mult_87_ab_15__32_), .B(
        u5_mult_87_CARRYB_14__32_), .CI(u5_mult_87_SUMB_14__33_), .CO(
        u5_mult_87_CARRYB_15__32_), .S(u5_mult_87_SUMB_15__32_) );
  FA_X1 u5_mult_87_S2_15_31 ( .A(u5_mult_87_ab_15__31_), .B(
        u5_mult_87_CARRYB_14__31_), .CI(u5_mult_87_SUMB_14__32_), .CO(
        u5_mult_87_CARRYB_15__31_), .S(u5_mult_87_SUMB_15__31_) );
  FA_X1 u5_mult_87_S2_15_30 ( .A(u5_mult_87_ab_15__30_), .B(
        u5_mult_87_CARRYB_14__30_), .CI(u5_mult_87_SUMB_14__31_), .CO(
        u5_mult_87_CARRYB_15__30_), .S(u5_mult_87_SUMB_15__30_) );
  FA_X1 u5_mult_87_S2_15_29 ( .A(u5_mult_87_ab_15__29_), .B(
        u5_mult_87_CARRYB_14__29_), .CI(u5_mult_87_SUMB_14__30_), .CO(
        u5_mult_87_CARRYB_15__29_), .S(u5_mult_87_SUMB_15__29_) );
  FA_X1 u5_mult_87_S2_15_28 ( .A(u5_mult_87_ab_15__28_), .B(
        u5_mult_87_CARRYB_14__28_), .CI(u5_mult_87_SUMB_14__29_), .CO(
        u5_mult_87_CARRYB_15__28_), .S(u5_mult_87_SUMB_15__28_) );
  FA_X1 u5_mult_87_S2_15_27 ( .A(u5_mult_87_ab_15__27_), .B(
        u5_mult_87_CARRYB_14__27_), .CI(u5_mult_87_SUMB_14__28_), .CO(
        u5_mult_87_CARRYB_15__27_), .S(u5_mult_87_SUMB_15__27_) );
  FA_X1 u5_mult_87_S2_15_26 ( .A(u5_mult_87_ab_15__26_), .B(
        u5_mult_87_CARRYB_14__26_), .CI(u5_mult_87_SUMB_14__27_), .CO(
        u5_mult_87_CARRYB_15__26_), .S(u5_mult_87_SUMB_15__26_) );
  FA_X1 u5_mult_87_S2_15_25 ( .A(u5_mult_87_ab_15__25_), .B(
        u5_mult_87_CARRYB_14__25_), .CI(u5_mult_87_SUMB_14__26_), .CO(
        u5_mult_87_CARRYB_15__25_), .S(u5_mult_87_SUMB_15__25_) );
  FA_X1 u5_mult_87_S2_15_24 ( .A(u5_mult_87_ab_15__24_), .B(
        u5_mult_87_CARRYB_14__24_), .CI(u5_mult_87_SUMB_14__25_), .CO(
        u5_mult_87_CARRYB_15__24_), .S(u5_mult_87_SUMB_15__24_) );
  FA_X1 u5_mult_87_S2_15_23 ( .A(u5_mult_87_ab_15__23_), .B(
        u5_mult_87_CARRYB_14__23_), .CI(u5_mult_87_SUMB_14__24_), .CO(
        u5_mult_87_CARRYB_15__23_), .S(u5_mult_87_SUMB_15__23_) );
  FA_X1 u5_mult_87_S2_15_22 ( .A(u5_mult_87_ab_15__22_), .B(
        u5_mult_87_CARRYB_14__22_), .CI(u5_mult_87_SUMB_14__23_), .CO(
        u5_mult_87_CARRYB_15__22_), .S(u5_mult_87_SUMB_15__22_) );
  FA_X1 u5_mult_87_S2_15_21 ( .A(u5_mult_87_ab_15__21_), .B(
        u5_mult_87_CARRYB_14__21_), .CI(u5_mult_87_SUMB_14__22_), .CO(
        u5_mult_87_CARRYB_15__21_), .S(u5_mult_87_SUMB_15__21_) );
  FA_X1 u5_mult_87_S2_15_20 ( .A(u5_mult_87_ab_15__20_), .B(
        u5_mult_87_CARRYB_14__20_), .CI(u5_mult_87_SUMB_14__21_), .CO(
        u5_mult_87_CARRYB_15__20_), .S(u5_mult_87_SUMB_15__20_) );
  FA_X1 u5_mult_87_S2_15_19 ( .A(u5_mult_87_ab_15__19_), .B(
        u5_mult_87_CARRYB_14__19_), .CI(u5_mult_87_SUMB_14__20_), .CO(
        u5_mult_87_CARRYB_15__19_), .S(u5_mult_87_SUMB_15__19_) );
  FA_X1 u5_mult_87_S2_15_18 ( .A(u5_mult_87_ab_15__18_), .B(
        u5_mult_87_CARRYB_14__18_), .CI(u5_mult_87_SUMB_14__19_), .CO(
        u5_mult_87_CARRYB_15__18_), .S(u5_mult_87_SUMB_15__18_) );
  FA_X1 u5_mult_87_S2_15_17 ( .A(u5_mult_87_ab_15__17_), .B(
        u5_mult_87_CARRYB_14__17_), .CI(u5_mult_87_SUMB_14__18_), .CO(
        u5_mult_87_CARRYB_15__17_), .S(u5_mult_87_SUMB_15__17_) );
  FA_X1 u5_mult_87_S2_15_16 ( .A(u5_mult_87_ab_15__16_), .B(
        u5_mult_87_CARRYB_14__16_), .CI(u5_mult_87_SUMB_14__17_), .CO(
        u5_mult_87_CARRYB_15__16_), .S(u5_mult_87_SUMB_15__16_) );
  FA_X1 u5_mult_87_S2_15_15 ( .A(u5_mult_87_ab_15__15_), .B(
        u5_mult_87_CARRYB_14__15_), .CI(u5_mult_87_SUMB_14__16_), .CO(
        u5_mult_87_CARRYB_15__15_), .S(u5_mult_87_SUMB_15__15_) );
  FA_X1 u5_mult_87_S2_15_14 ( .A(u5_mult_87_ab_15__14_), .B(
        u5_mult_87_CARRYB_14__14_), .CI(u5_mult_87_SUMB_14__15_), .CO(
        u5_mult_87_CARRYB_15__14_), .S(u5_mult_87_SUMB_15__14_) );
  FA_X1 u5_mult_87_S2_15_13 ( .A(u5_mult_87_ab_15__13_), .B(
        u5_mult_87_CARRYB_14__13_), .CI(u5_mult_87_SUMB_14__14_), .CO(
        u5_mult_87_CARRYB_15__13_), .S(u5_mult_87_SUMB_15__13_) );
  FA_X1 u5_mult_87_S2_15_12 ( .A(u5_mult_87_ab_15__12_), .B(
        u5_mult_87_CARRYB_14__12_), .CI(u5_mult_87_SUMB_14__13_), .CO(
        u5_mult_87_CARRYB_15__12_), .S(u5_mult_87_SUMB_15__12_) );
  FA_X1 u5_mult_87_S2_15_11 ( .A(u5_mult_87_ab_15__11_), .B(
        u5_mult_87_CARRYB_14__11_), .CI(u5_mult_87_SUMB_14__12_), .CO(
        u5_mult_87_CARRYB_15__11_), .S(u5_mult_87_SUMB_15__11_) );
  FA_X1 u5_mult_87_S2_15_10 ( .A(u5_mult_87_ab_15__10_), .B(
        u5_mult_87_CARRYB_14__10_), .CI(u5_mult_87_SUMB_14__11_), .CO(
        u5_mult_87_CARRYB_15__10_), .S(u5_mult_87_SUMB_15__10_) );
  FA_X1 u5_mult_87_S2_15_9 ( .A(u5_mult_87_ab_15__9_), .B(
        u5_mult_87_CARRYB_14__9_), .CI(u5_mult_87_SUMB_14__10_), .CO(
        u5_mult_87_CARRYB_15__9_), .S(u5_mult_87_SUMB_15__9_) );
  FA_X1 u5_mult_87_S2_15_8 ( .A(u5_mult_87_ab_15__8_), .B(
        u5_mult_87_CARRYB_14__8_), .CI(u5_mult_87_SUMB_14__9_), .CO(
        u5_mult_87_CARRYB_15__8_), .S(u5_mult_87_SUMB_15__8_) );
  FA_X1 u5_mult_87_S2_15_7 ( .A(u5_mult_87_ab_15__7_), .B(
        u5_mult_87_CARRYB_14__7_), .CI(u5_mult_87_SUMB_14__8_), .CO(
        u5_mult_87_CARRYB_15__7_), .S(u5_mult_87_SUMB_15__7_) );
  FA_X1 u5_mult_87_S2_15_6 ( .A(u5_mult_87_ab_15__6_), .B(
        u5_mult_87_CARRYB_14__6_), .CI(u5_mult_87_SUMB_14__7_), .CO(
        u5_mult_87_CARRYB_15__6_), .S(u5_mult_87_SUMB_15__6_) );
  FA_X1 u5_mult_87_S2_15_5 ( .A(u5_mult_87_ab_15__5_), .B(
        u5_mult_87_CARRYB_14__5_), .CI(u5_mult_87_SUMB_14__6_), .CO(
        u5_mult_87_CARRYB_15__5_), .S(u5_mult_87_SUMB_15__5_) );
  FA_X1 u5_mult_87_S2_15_4 ( .A(u5_mult_87_ab_15__4_), .B(
        u5_mult_87_CARRYB_14__4_), .CI(u5_mult_87_SUMB_14__5_), .CO(
        u5_mult_87_CARRYB_15__4_), .S(u5_mult_87_SUMB_15__4_) );
  FA_X1 u5_mult_87_S2_15_3 ( .A(u5_mult_87_ab_15__3_), .B(
        u5_mult_87_CARRYB_14__3_), .CI(u5_mult_87_SUMB_14__4_), .CO(
        u5_mult_87_CARRYB_15__3_), .S(u5_mult_87_SUMB_15__3_) );
  FA_X1 u5_mult_87_S2_15_2 ( .A(u5_mult_87_ab_15__2_), .B(
        u5_mult_87_CARRYB_14__2_), .CI(u5_mult_87_SUMB_14__3_), .CO(
        u5_mult_87_CARRYB_15__2_), .S(u5_mult_87_SUMB_15__2_) );
  FA_X1 u5_mult_87_S2_15_1 ( .A(u5_mult_87_ab_15__1_), .B(
        u5_mult_87_CARRYB_14__1_), .CI(u5_mult_87_SUMB_14__2_), .CO(
        u5_mult_87_CARRYB_15__1_), .S(u5_mult_87_SUMB_15__1_) );
  FA_X1 u5_mult_87_S1_15_0 ( .A(u5_mult_87_ab_15__0_), .B(
        u5_mult_87_CARRYB_14__0_), .CI(u5_mult_87_SUMB_14__1_), .CO(
        u5_mult_87_CARRYB_15__0_), .S(u5_N15) );
  FA_X1 u5_mult_87_S3_16_51 ( .A(u5_mult_87_ab_16__51_), .B(
        u5_mult_87_CARRYB_15__51_), .CI(u5_mult_87_ab_15__52_), .CO(
        u5_mult_87_CARRYB_16__51_), .S(u5_mult_87_SUMB_16__51_) );
  FA_X1 u5_mult_87_S2_16_50 ( .A(u5_mult_87_ab_16__50_), .B(
        u5_mult_87_CARRYB_15__50_), .CI(u5_mult_87_SUMB_15__51_), .CO(
        u5_mult_87_CARRYB_16__50_), .S(u5_mult_87_SUMB_16__50_) );
  FA_X1 u5_mult_87_S2_16_49 ( .A(u5_mult_87_ab_16__49_), .B(
        u5_mult_87_CARRYB_15__49_), .CI(u5_mult_87_SUMB_15__50_), .CO(
        u5_mult_87_CARRYB_16__49_), .S(u5_mult_87_SUMB_16__49_) );
  FA_X1 u5_mult_87_S2_16_48 ( .A(u5_mult_87_ab_16__48_), .B(
        u5_mult_87_CARRYB_15__48_), .CI(u5_mult_87_SUMB_15__49_), .CO(
        u5_mult_87_CARRYB_16__48_), .S(u5_mult_87_SUMB_16__48_) );
  FA_X1 u5_mult_87_S2_16_47 ( .A(u5_mult_87_ab_16__47_), .B(
        u5_mult_87_CARRYB_15__47_), .CI(u5_mult_87_SUMB_15__48_), .CO(
        u5_mult_87_CARRYB_16__47_), .S(u5_mult_87_SUMB_16__47_) );
  FA_X1 u5_mult_87_S2_16_46 ( .A(u5_mult_87_ab_16__46_), .B(
        u5_mult_87_CARRYB_15__46_), .CI(u5_mult_87_SUMB_15__47_), .CO(
        u5_mult_87_CARRYB_16__46_), .S(u5_mult_87_SUMB_16__46_) );
  FA_X1 u5_mult_87_S2_16_45 ( .A(u5_mult_87_ab_16__45_), .B(
        u5_mult_87_CARRYB_15__45_), .CI(u5_mult_87_SUMB_15__46_), .CO(
        u5_mult_87_CARRYB_16__45_), .S(u5_mult_87_SUMB_16__45_) );
  FA_X1 u5_mult_87_S2_16_44 ( .A(u5_mult_87_ab_16__44_), .B(
        u5_mult_87_CARRYB_15__44_), .CI(u5_mult_87_SUMB_15__45_), .CO(
        u5_mult_87_CARRYB_16__44_), .S(u5_mult_87_SUMB_16__44_) );
  FA_X1 u5_mult_87_S2_16_43 ( .A(u5_mult_87_ab_16__43_), .B(
        u5_mult_87_CARRYB_15__43_), .CI(u5_mult_87_SUMB_15__44_), .CO(
        u5_mult_87_CARRYB_16__43_), .S(u5_mult_87_SUMB_16__43_) );
  FA_X1 u5_mult_87_S2_16_42 ( .A(u5_mult_87_ab_16__42_), .B(
        u5_mult_87_CARRYB_15__42_), .CI(u5_mult_87_SUMB_15__43_), .CO(
        u5_mult_87_CARRYB_16__42_), .S(u5_mult_87_SUMB_16__42_) );
  FA_X1 u5_mult_87_S2_16_41 ( .A(u5_mult_87_ab_16__41_), .B(
        u5_mult_87_CARRYB_15__41_), .CI(u5_mult_87_SUMB_15__42_), .CO(
        u5_mult_87_CARRYB_16__41_), .S(u5_mult_87_SUMB_16__41_) );
  FA_X1 u5_mult_87_S2_16_40 ( .A(u5_mult_87_ab_16__40_), .B(
        u5_mult_87_CARRYB_15__40_), .CI(u5_mult_87_SUMB_15__41_), .CO(
        u5_mult_87_CARRYB_16__40_), .S(u5_mult_87_SUMB_16__40_) );
  FA_X1 u5_mult_87_S2_16_39 ( .A(u5_mult_87_ab_16__39_), .B(
        u5_mult_87_CARRYB_15__39_), .CI(u5_mult_87_SUMB_15__40_), .CO(
        u5_mult_87_CARRYB_16__39_), .S(u5_mult_87_SUMB_16__39_) );
  FA_X1 u5_mult_87_S2_16_38 ( .A(u5_mult_87_ab_16__38_), .B(
        u5_mult_87_CARRYB_15__38_), .CI(u5_mult_87_SUMB_15__39_), .CO(
        u5_mult_87_CARRYB_16__38_), .S(u5_mult_87_SUMB_16__38_) );
  FA_X1 u5_mult_87_S2_16_37 ( .A(u5_mult_87_ab_16__37_), .B(
        u5_mult_87_CARRYB_15__37_), .CI(u5_mult_87_SUMB_15__38_), .CO(
        u5_mult_87_CARRYB_16__37_), .S(u5_mult_87_SUMB_16__37_) );
  FA_X1 u5_mult_87_S2_16_36 ( .A(u5_mult_87_ab_16__36_), .B(
        u5_mult_87_CARRYB_15__36_), .CI(u5_mult_87_SUMB_15__37_), .CO(
        u5_mult_87_CARRYB_16__36_), .S(u5_mult_87_SUMB_16__36_) );
  FA_X1 u5_mult_87_S2_16_35 ( .A(u5_mult_87_ab_16__35_), .B(
        u5_mult_87_CARRYB_15__35_), .CI(u5_mult_87_SUMB_15__36_), .CO(
        u5_mult_87_CARRYB_16__35_), .S(u5_mult_87_SUMB_16__35_) );
  FA_X1 u5_mult_87_S2_16_34 ( .A(u5_mult_87_ab_16__34_), .B(
        u5_mult_87_CARRYB_15__34_), .CI(u5_mult_87_SUMB_15__35_), .CO(
        u5_mult_87_CARRYB_16__34_), .S(u5_mult_87_SUMB_16__34_) );
  FA_X1 u5_mult_87_S2_16_33 ( .A(u5_mult_87_ab_16__33_), .B(
        u5_mult_87_CARRYB_15__33_), .CI(u5_mult_87_SUMB_15__34_), .CO(
        u5_mult_87_CARRYB_16__33_), .S(u5_mult_87_SUMB_16__33_) );
  FA_X1 u5_mult_87_S2_16_32 ( .A(u5_mult_87_ab_16__32_), .B(
        u5_mult_87_CARRYB_15__32_), .CI(u5_mult_87_SUMB_15__33_), .CO(
        u5_mult_87_CARRYB_16__32_), .S(u5_mult_87_SUMB_16__32_) );
  FA_X1 u5_mult_87_S2_16_31 ( .A(u5_mult_87_ab_16__31_), .B(
        u5_mult_87_CARRYB_15__31_), .CI(u5_mult_87_SUMB_15__32_), .CO(
        u5_mult_87_CARRYB_16__31_), .S(u5_mult_87_SUMB_16__31_) );
  FA_X1 u5_mult_87_S2_16_30 ( .A(u5_mult_87_ab_16__30_), .B(
        u5_mult_87_CARRYB_15__30_), .CI(u5_mult_87_SUMB_15__31_), .CO(
        u5_mult_87_CARRYB_16__30_), .S(u5_mult_87_SUMB_16__30_) );
  FA_X1 u5_mult_87_S2_16_29 ( .A(u5_mult_87_ab_16__29_), .B(
        u5_mult_87_CARRYB_15__29_), .CI(u5_mult_87_SUMB_15__30_), .CO(
        u5_mult_87_CARRYB_16__29_), .S(u5_mult_87_SUMB_16__29_) );
  FA_X1 u5_mult_87_S2_16_28 ( .A(u5_mult_87_ab_16__28_), .B(
        u5_mult_87_CARRYB_15__28_), .CI(u5_mult_87_SUMB_15__29_), .CO(
        u5_mult_87_CARRYB_16__28_), .S(u5_mult_87_SUMB_16__28_) );
  FA_X1 u5_mult_87_S2_16_27 ( .A(u5_mult_87_ab_16__27_), .B(
        u5_mult_87_CARRYB_15__27_), .CI(u5_mult_87_SUMB_15__28_), .CO(
        u5_mult_87_CARRYB_16__27_), .S(u5_mult_87_SUMB_16__27_) );
  FA_X1 u5_mult_87_S2_16_26 ( .A(u5_mult_87_ab_16__26_), .B(
        u5_mult_87_CARRYB_15__26_), .CI(u5_mult_87_SUMB_15__27_), .CO(
        u5_mult_87_CARRYB_16__26_), .S(u5_mult_87_SUMB_16__26_) );
  FA_X1 u5_mult_87_S2_16_25 ( .A(u5_mult_87_ab_16__25_), .B(
        u5_mult_87_CARRYB_15__25_), .CI(u5_mult_87_SUMB_15__26_), .CO(
        u5_mult_87_CARRYB_16__25_), .S(u5_mult_87_SUMB_16__25_) );
  FA_X1 u5_mult_87_S2_16_24 ( .A(u5_mult_87_ab_16__24_), .B(
        u5_mult_87_CARRYB_15__24_), .CI(u5_mult_87_SUMB_15__25_), .CO(
        u5_mult_87_CARRYB_16__24_), .S(u5_mult_87_SUMB_16__24_) );
  FA_X1 u5_mult_87_S2_16_23 ( .A(u5_mult_87_ab_16__23_), .B(
        u5_mult_87_CARRYB_15__23_), .CI(u5_mult_87_SUMB_15__24_), .CO(
        u5_mult_87_CARRYB_16__23_), .S(u5_mult_87_SUMB_16__23_) );
  FA_X1 u5_mult_87_S2_16_22 ( .A(u5_mult_87_ab_16__22_), .B(
        u5_mult_87_CARRYB_15__22_), .CI(u5_mult_87_SUMB_15__23_), .CO(
        u5_mult_87_CARRYB_16__22_), .S(u5_mult_87_SUMB_16__22_) );
  FA_X1 u5_mult_87_S2_16_21 ( .A(u5_mult_87_ab_16__21_), .B(
        u5_mult_87_CARRYB_15__21_), .CI(u5_mult_87_SUMB_15__22_), .CO(
        u5_mult_87_CARRYB_16__21_), .S(u5_mult_87_SUMB_16__21_) );
  FA_X1 u5_mult_87_S2_16_20 ( .A(u5_mult_87_ab_16__20_), .B(
        u5_mult_87_CARRYB_15__20_), .CI(u5_mult_87_SUMB_15__21_), .CO(
        u5_mult_87_CARRYB_16__20_), .S(u5_mult_87_SUMB_16__20_) );
  FA_X1 u5_mult_87_S2_16_19 ( .A(u5_mult_87_ab_16__19_), .B(
        u5_mult_87_CARRYB_15__19_), .CI(u5_mult_87_SUMB_15__20_), .CO(
        u5_mult_87_CARRYB_16__19_), .S(u5_mult_87_SUMB_16__19_) );
  FA_X1 u5_mult_87_S2_16_18 ( .A(u5_mult_87_ab_16__18_), .B(
        u5_mult_87_CARRYB_15__18_), .CI(u5_mult_87_SUMB_15__19_), .CO(
        u5_mult_87_CARRYB_16__18_), .S(u5_mult_87_SUMB_16__18_) );
  FA_X1 u5_mult_87_S2_16_17 ( .A(u5_mult_87_ab_16__17_), .B(
        u5_mult_87_CARRYB_15__17_), .CI(u5_mult_87_SUMB_15__18_), .CO(
        u5_mult_87_CARRYB_16__17_), .S(u5_mult_87_SUMB_16__17_) );
  FA_X1 u5_mult_87_S2_16_16 ( .A(u5_mult_87_ab_16__16_), .B(
        u5_mult_87_CARRYB_15__16_), .CI(u5_mult_87_SUMB_15__17_), .CO(
        u5_mult_87_CARRYB_16__16_), .S(u5_mult_87_SUMB_16__16_) );
  FA_X1 u5_mult_87_S2_16_15 ( .A(u5_mult_87_ab_16__15_), .B(
        u5_mult_87_CARRYB_15__15_), .CI(u5_mult_87_SUMB_15__16_), .CO(
        u5_mult_87_CARRYB_16__15_), .S(u5_mult_87_SUMB_16__15_) );
  FA_X1 u5_mult_87_S2_16_14 ( .A(u5_mult_87_ab_16__14_), .B(
        u5_mult_87_CARRYB_15__14_), .CI(u5_mult_87_SUMB_15__15_), .CO(
        u5_mult_87_CARRYB_16__14_), .S(u5_mult_87_SUMB_16__14_) );
  FA_X1 u5_mult_87_S2_16_13 ( .A(u5_mult_87_ab_16__13_), .B(
        u5_mult_87_CARRYB_15__13_), .CI(u5_mult_87_SUMB_15__14_), .CO(
        u5_mult_87_CARRYB_16__13_), .S(u5_mult_87_SUMB_16__13_) );
  FA_X1 u5_mult_87_S2_16_12 ( .A(u5_mult_87_ab_16__12_), .B(
        u5_mult_87_CARRYB_15__12_), .CI(u5_mult_87_SUMB_15__13_), .CO(
        u5_mult_87_CARRYB_16__12_), .S(u5_mult_87_SUMB_16__12_) );
  FA_X1 u5_mult_87_S2_16_11 ( .A(u5_mult_87_ab_16__11_), .B(
        u5_mult_87_CARRYB_15__11_), .CI(u5_mult_87_SUMB_15__12_), .CO(
        u5_mult_87_CARRYB_16__11_), .S(u5_mult_87_SUMB_16__11_) );
  FA_X1 u5_mult_87_S2_16_10 ( .A(u5_mult_87_ab_16__10_), .B(
        u5_mult_87_CARRYB_15__10_), .CI(u5_mult_87_SUMB_15__11_), .CO(
        u5_mult_87_CARRYB_16__10_), .S(u5_mult_87_SUMB_16__10_) );
  FA_X1 u5_mult_87_S2_16_9 ( .A(u5_mult_87_ab_16__9_), .B(
        u5_mult_87_CARRYB_15__9_), .CI(u5_mult_87_SUMB_15__10_), .CO(
        u5_mult_87_CARRYB_16__9_), .S(u5_mult_87_SUMB_16__9_) );
  FA_X1 u5_mult_87_S2_16_8 ( .A(u5_mult_87_ab_16__8_), .B(
        u5_mult_87_CARRYB_15__8_), .CI(u5_mult_87_SUMB_15__9_), .CO(
        u5_mult_87_CARRYB_16__8_), .S(u5_mult_87_SUMB_16__8_) );
  FA_X1 u5_mult_87_S2_16_7 ( .A(u5_mult_87_ab_16__7_), .B(
        u5_mult_87_CARRYB_15__7_), .CI(u5_mult_87_SUMB_15__8_), .CO(
        u5_mult_87_CARRYB_16__7_), .S(u5_mult_87_SUMB_16__7_) );
  FA_X1 u5_mult_87_S2_16_6 ( .A(u5_mult_87_ab_16__6_), .B(
        u5_mult_87_CARRYB_15__6_), .CI(u5_mult_87_SUMB_15__7_), .CO(
        u5_mult_87_CARRYB_16__6_), .S(u5_mult_87_SUMB_16__6_) );
  FA_X1 u5_mult_87_S2_16_5 ( .A(u5_mult_87_ab_16__5_), .B(
        u5_mult_87_CARRYB_15__5_), .CI(u5_mult_87_SUMB_15__6_), .CO(
        u5_mult_87_CARRYB_16__5_), .S(u5_mult_87_SUMB_16__5_) );
  FA_X1 u5_mult_87_S2_16_4 ( .A(u5_mult_87_ab_16__4_), .B(
        u5_mult_87_CARRYB_15__4_), .CI(u5_mult_87_SUMB_15__5_), .CO(
        u5_mult_87_CARRYB_16__4_), .S(u5_mult_87_SUMB_16__4_) );
  FA_X1 u5_mult_87_S2_16_3 ( .A(u5_mult_87_ab_16__3_), .B(
        u5_mult_87_CARRYB_15__3_), .CI(u5_mult_87_SUMB_15__4_), .CO(
        u5_mult_87_CARRYB_16__3_), .S(u5_mult_87_SUMB_16__3_) );
  FA_X1 u5_mult_87_S2_16_2 ( .A(u5_mult_87_ab_16__2_), .B(
        u5_mult_87_CARRYB_15__2_), .CI(u5_mult_87_SUMB_15__3_), .CO(
        u5_mult_87_CARRYB_16__2_), .S(u5_mult_87_SUMB_16__2_) );
  FA_X1 u5_mult_87_S2_16_1 ( .A(u5_mult_87_ab_16__1_), .B(
        u5_mult_87_CARRYB_15__1_), .CI(u5_mult_87_SUMB_15__2_), .CO(
        u5_mult_87_CARRYB_16__1_), .S(u5_mult_87_SUMB_16__1_) );
  FA_X1 u5_mult_87_S1_16_0 ( .A(u5_mult_87_ab_16__0_), .B(
        u5_mult_87_CARRYB_15__0_), .CI(u5_mult_87_SUMB_15__1_), .CO(
        u5_mult_87_CARRYB_16__0_), .S(u5_N16) );
  FA_X1 u5_mult_87_S3_17_51 ( .A(u5_mult_87_ab_17__51_), .B(
        u5_mult_87_CARRYB_16__51_), .CI(u5_mult_87_ab_16__52_), .CO(
        u5_mult_87_CARRYB_17__51_), .S(u5_mult_87_SUMB_17__51_) );
  FA_X1 u5_mult_87_S2_17_50 ( .A(u5_mult_87_ab_17__50_), .B(
        u5_mult_87_CARRYB_16__50_), .CI(u5_mult_87_SUMB_16__51_), .CO(
        u5_mult_87_CARRYB_17__50_), .S(u5_mult_87_SUMB_17__50_) );
  FA_X1 u5_mult_87_S2_17_49 ( .A(u5_mult_87_ab_17__49_), .B(
        u5_mult_87_CARRYB_16__49_), .CI(u5_mult_87_SUMB_16__50_), .CO(
        u5_mult_87_CARRYB_17__49_), .S(u5_mult_87_SUMB_17__49_) );
  FA_X1 u5_mult_87_S2_17_48 ( .A(u5_mult_87_ab_17__48_), .B(
        u5_mult_87_CARRYB_16__48_), .CI(u5_mult_87_SUMB_16__49_), .CO(
        u5_mult_87_CARRYB_17__48_), .S(u5_mult_87_SUMB_17__48_) );
  FA_X1 u5_mult_87_S2_17_47 ( .A(u5_mult_87_ab_17__47_), .B(
        u5_mult_87_CARRYB_16__47_), .CI(u5_mult_87_SUMB_16__48_), .CO(
        u5_mult_87_CARRYB_17__47_), .S(u5_mult_87_SUMB_17__47_) );
  FA_X1 u5_mult_87_S2_17_46 ( .A(u5_mult_87_ab_17__46_), .B(
        u5_mult_87_CARRYB_16__46_), .CI(u5_mult_87_SUMB_16__47_), .CO(
        u5_mult_87_CARRYB_17__46_), .S(u5_mult_87_SUMB_17__46_) );
  FA_X1 u5_mult_87_S2_17_45 ( .A(u5_mult_87_ab_17__45_), .B(
        u5_mult_87_CARRYB_16__45_), .CI(u5_mult_87_SUMB_16__46_), .CO(
        u5_mult_87_CARRYB_17__45_), .S(u5_mult_87_SUMB_17__45_) );
  FA_X1 u5_mult_87_S2_17_44 ( .A(u5_mult_87_ab_17__44_), .B(
        u5_mult_87_CARRYB_16__44_), .CI(u5_mult_87_SUMB_16__45_), .CO(
        u5_mult_87_CARRYB_17__44_), .S(u5_mult_87_SUMB_17__44_) );
  FA_X1 u5_mult_87_S2_17_43 ( .A(u5_mult_87_ab_17__43_), .B(
        u5_mult_87_CARRYB_16__43_), .CI(u5_mult_87_SUMB_16__44_), .CO(
        u5_mult_87_CARRYB_17__43_), .S(u5_mult_87_SUMB_17__43_) );
  FA_X1 u5_mult_87_S2_17_42 ( .A(u5_mult_87_ab_17__42_), .B(
        u5_mult_87_CARRYB_16__42_), .CI(u5_mult_87_SUMB_16__43_), .CO(
        u5_mult_87_CARRYB_17__42_), .S(u5_mult_87_SUMB_17__42_) );
  FA_X1 u5_mult_87_S2_17_41 ( .A(u5_mult_87_ab_17__41_), .B(
        u5_mult_87_CARRYB_16__41_), .CI(u5_mult_87_SUMB_16__42_), .CO(
        u5_mult_87_CARRYB_17__41_), .S(u5_mult_87_SUMB_17__41_) );
  FA_X1 u5_mult_87_S2_17_40 ( .A(u5_mult_87_ab_17__40_), .B(
        u5_mult_87_CARRYB_16__40_), .CI(u5_mult_87_SUMB_16__41_), .CO(
        u5_mult_87_CARRYB_17__40_), .S(u5_mult_87_SUMB_17__40_) );
  FA_X1 u5_mult_87_S2_17_39 ( .A(u5_mult_87_ab_17__39_), .B(
        u5_mult_87_CARRYB_16__39_), .CI(u5_mult_87_SUMB_16__40_), .CO(
        u5_mult_87_CARRYB_17__39_), .S(u5_mult_87_SUMB_17__39_) );
  FA_X1 u5_mult_87_S2_17_38 ( .A(u5_mult_87_ab_17__38_), .B(
        u5_mult_87_CARRYB_16__38_), .CI(u5_mult_87_SUMB_16__39_), .CO(
        u5_mult_87_CARRYB_17__38_), .S(u5_mult_87_SUMB_17__38_) );
  FA_X1 u5_mult_87_S2_17_37 ( .A(u5_mult_87_ab_17__37_), .B(
        u5_mult_87_CARRYB_16__37_), .CI(u5_mult_87_SUMB_16__38_), .CO(
        u5_mult_87_CARRYB_17__37_), .S(u5_mult_87_SUMB_17__37_) );
  FA_X1 u5_mult_87_S2_17_36 ( .A(u5_mult_87_ab_17__36_), .B(
        u5_mult_87_CARRYB_16__36_), .CI(u5_mult_87_SUMB_16__37_), .CO(
        u5_mult_87_CARRYB_17__36_), .S(u5_mult_87_SUMB_17__36_) );
  FA_X1 u5_mult_87_S2_17_35 ( .A(u5_mult_87_ab_17__35_), .B(
        u5_mult_87_CARRYB_16__35_), .CI(u5_mult_87_SUMB_16__36_), .CO(
        u5_mult_87_CARRYB_17__35_), .S(u5_mult_87_SUMB_17__35_) );
  FA_X1 u5_mult_87_S2_17_34 ( .A(u5_mult_87_ab_17__34_), .B(
        u5_mult_87_CARRYB_16__34_), .CI(u5_mult_87_SUMB_16__35_), .CO(
        u5_mult_87_CARRYB_17__34_), .S(u5_mult_87_SUMB_17__34_) );
  FA_X1 u5_mult_87_S2_17_33 ( .A(u5_mult_87_ab_17__33_), .B(
        u5_mult_87_CARRYB_16__33_), .CI(u5_mult_87_SUMB_16__34_), .CO(
        u5_mult_87_CARRYB_17__33_), .S(u5_mult_87_SUMB_17__33_) );
  FA_X1 u5_mult_87_S2_17_32 ( .A(u5_mult_87_ab_17__32_), .B(
        u5_mult_87_CARRYB_16__32_), .CI(u5_mult_87_SUMB_16__33_), .CO(
        u5_mult_87_CARRYB_17__32_), .S(u5_mult_87_SUMB_17__32_) );
  FA_X1 u5_mult_87_S2_17_31 ( .A(u5_mult_87_ab_17__31_), .B(
        u5_mult_87_CARRYB_16__31_), .CI(u5_mult_87_SUMB_16__32_), .CO(
        u5_mult_87_CARRYB_17__31_), .S(u5_mult_87_SUMB_17__31_) );
  FA_X1 u5_mult_87_S2_17_30 ( .A(u5_mult_87_ab_17__30_), .B(
        u5_mult_87_CARRYB_16__30_), .CI(u5_mult_87_SUMB_16__31_), .CO(
        u5_mult_87_CARRYB_17__30_), .S(u5_mult_87_SUMB_17__30_) );
  FA_X1 u5_mult_87_S2_17_29 ( .A(u5_mult_87_ab_17__29_), .B(
        u5_mult_87_CARRYB_16__29_), .CI(u5_mult_87_SUMB_16__30_), .CO(
        u5_mult_87_CARRYB_17__29_), .S(u5_mult_87_SUMB_17__29_) );
  FA_X1 u5_mult_87_S2_17_28 ( .A(u5_mult_87_ab_17__28_), .B(
        u5_mult_87_CARRYB_16__28_), .CI(u5_mult_87_SUMB_16__29_), .CO(
        u5_mult_87_CARRYB_17__28_), .S(u5_mult_87_SUMB_17__28_) );
  FA_X1 u5_mult_87_S2_17_27 ( .A(u5_mult_87_ab_17__27_), .B(
        u5_mult_87_CARRYB_16__27_), .CI(u5_mult_87_SUMB_16__28_), .CO(
        u5_mult_87_CARRYB_17__27_), .S(u5_mult_87_SUMB_17__27_) );
  FA_X1 u5_mult_87_S2_17_26 ( .A(u5_mult_87_ab_17__26_), .B(
        u5_mult_87_CARRYB_16__26_), .CI(u5_mult_87_SUMB_16__27_), .CO(
        u5_mult_87_CARRYB_17__26_), .S(u5_mult_87_SUMB_17__26_) );
  FA_X1 u5_mult_87_S2_17_25 ( .A(u5_mult_87_ab_17__25_), .B(
        u5_mult_87_CARRYB_16__25_), .CI(u5_mult_87_SUMB_16__26_), .CO(
        u5_mult_87_CARRYB_17__25_), .S(u5_mult_87_SUMB_17__25_) );
  FA_X1 u5_mult_87_S2_17_24 ( .A(u5_mult_87_ab_17__24_), .B(
        u5_mult_87_CARRYB_16__24_), .CI(u5_mult_87_SUMB_16__25_), .CO(
        u5_mult_87_CARRYB_17__24_), .S(u5_mult_87_SUMB_17__24_) );
  FA_X1 u5_mult_87_S2_17_23 ( .A(u5_mult_87_ab_17__23_), .B(
        u5_mult_87_CARRYB_16__23_), .CI(u5_mult_87_SUMB_16__24_), .CO(
        u5_mult_87_CARRYB_17__23_), .S(u5_mult_87_SUMB_17__23_) );
  FA_X1 u5_mult_87_S2_17_22 ( .A(u5_mult_87_ab_17__22_), .B(
        u5_mult_87_CARRYB_16__22_), .CI(u5_mult_87_SUMB_16__23_), .CO(
        u5_mult_87_CARRYB_17__22_), .S(u5_mult_87_SUMB_17__22_) );
  FA_X1 u5_mult_87_S2_17_21 ( .A(u5_mult_87_ab_17__21_), .B(
        u5_mult_87_CARRYB_16__21_), .CI(u5_mult_87_SUMB_16__22_), .CO(
        u5_mult_87_CARRYB_17__21_), .S(u5_mult_87_SUMB_17__21_) );
  FA_X1 u5_mult_87_S2_17_20 ( .A(u5_mult_87_ab_17__20_), .B(
        u5_mult_87_CARRYB_16__20_), .CI(u5_mult_87_SUMB_16__21_), .CO(
        u5_mult_87_CARRYB_17__20_), .S(u5_mult_87_SUMB_17__20_) );
  FA_X1 u5_mult_87_S2_17_19 ( .A(u5_mult_87_ab_17__19_), .B(
        u5_mult_87_CARRYB_16__19_), .CI(u5_mult_87_SUMB_16__20_), .CO(
        u5_mult_87_CARRYB_17__19_), .S(u5_mult_87_SUMB_17__19_) );
  FA_X1 u5_mult_87_S2_17_18 ( .A(u5_mult_87_ab_17__18_), .B(
        u5_mult_87_CARRYB_16__18_), .CI(u5_mult_87_SUMB_16__19_), .CO(
        u5_mult_87_CARRYB_17__18_), .S(u5_mult_87_SUMB_17__18_) );
  FA_X1 u5_mult_87_S2_17_17 ( .A(u5_mult_87_ab_17__17_), .B(
        u5_mult_87_CARRYB_16__17_), .CI(u5_mult_87_SUMB_16__18_), .CO(
        u5_mult_87_CARRYB_17__17_), .S(u5_mult_87_SUMB_17__17_) );
  FA_X1 u5_mult_87_S2_17_16 ( .A(u5_mult_87_ab_17__16_), .B(
        u5_mult_87_CARRYB_16__16_), .CI(u5_mult_87_SUMB_16__17_), .CO(
        u5_mult_87_CARRYB_17__16_), .S(u5_mult_87_SUMB_17__16_) );
  FA_X1 u5_mult_87_S2_17_15 ( .A(u5_mult_87_ab_17__15_), .B(
        u5_mult_87_CARRYB_16__15_), .CI(u5_mult_87_SUMB_16__16_), .CO(
        u5_mult_87_CARRYB_17__15_), .S(u5_mult_87_SUMB_17__15_) );
  FA_X1 u5_mult_87_S2_17_14 ( .A(u5_mult_87_ab_17__14_), .B(
        u5_mult_87_CARRYB_16__14_), .CI(u5_mult_87_SUMB_16__15_), .CO(
        u5_mult_87_CARRYB_17__14_), .S(u5_mult_87_SUMB_17__14_) );
  FA_X1 u5_mult_87_S2_17_13 ( .A(u5_mult_87_ab_17__13_), .B(
        u5_mult_87_CARRYB_16__13_), .CI(u5_mult_87_SUMB_16__14_), .CO(
        u5_mult_87_CARRYB_17__13_), .S(u5_mult_87_SUMB_17__13_) );
  FA_X1 u5_mult_87_S2_17_12 ( .A(u5_mult_87_ab_17__12_), .B(
        u5_mult_87_CARRYB_16__12_), .CI(u5_mult_87_SUMB_16__13_), .CO(
        u5_mult_87_CARRYB_17__12_), .S(u5_mult_87_SUMB_17__12_) );
  FA_X1 u5_mult_87_S2_17_11 ( .A(u5_mult_87_ab_17__11_), .B(
        u5_mult_87_CARRYB_16__11_), .CI(u5_mult_87_SUMB_16__12_), .CO(
        u5_mult_87_CARRYB_17__11_), .S(u5_mult_87_SUMB_17__11_) );
  FA_X1 u5_mult_87_S2_17_10 ( .A(u5_mult_87_ab_17__10_), .B(
        u5_mult_87_CARRYB_16__10_), .CI(u5_mult_87_SUMB_16__11_), .CO(
        u5_mult_87_CARRYB_17__10_), .S(u5_mult_87_SUMB_17__10_) );
  FA_X1 u5_mult_87_S2_17_9 ( .A(u5_mult_87_ab_17__9_), .B(
        u5_mult_87_CARRYB_16__9_), .CI(u5_mult_87_SUMB_16__10_), .CO(
        u5_mult_87_CARRYB_17__9_), .S(u5_mult_87_SUMB_17__9_) );
  FA_X1 u5_mult_87_S2_17_8 ( .A(u5_mult_87_ab_17__8_), .B(
        u5_mult_87_CARRYB_16__8_), .CI(u5_mult_87_SUMB_16__9_), .CO(
        u5_mult_87_CARRYB_17__8_), .S(u5_mult_87_SUMB_17__8_) );
  FA_X1 u5_mult_87_S2_17_7 ( .A(u5_mult_87_ab_17__7_), .B(
        u5_mult_87_CARRYB_16__7_), .CI(u5_mult_87_SUMB_16__8_), .CO(
        u5_mult_87_CARRYB_17__7_), .S(u5_mult_87_SUMB_17__7_) );
  FA_X1 u5_mult_87_S2_17_6 ( .A(u5_mult_87_ab_17__6_), .B(
        u5_mult_87_CARRYB_16__6_), .CI(u5_mult_87_SUMB_16__7_), .CO(
        u5_mult_87_CARRYB_17__6_), .S(u5_mult_87_SUMB_17__6_) );
  FA_X1 u5_mult_87_S2_17_5 ( .A(u5_mult_87_ab_17__5_), .B(
        u5_mult_87_CARRYB_16__5_), .CI(u5_mult_87_SUMB_16__6_), .CO(
        u5_mult_87_CARRYB_17__5_), .S(u5_mult_87_SUMB_17__5_) );
  FA_X1 u5_mult_87_S2_17_4 ( .A(u5_mult_87_ab_17__4_), .B(
        u5_mult_87_CARRYB_16__4_), .CI(u5_mult_87_SUMB_16__5_), .CO(
        u5_mult_87_CARRYB_17__4_), .S(u5_mult_87_SUMB_17__4_) );
  FA_X1 u5_mult_87_S2_17_3 ( .A(u5_mult_87_ab_17__3_), .B(
        u5_mult_87_CARRYB_16__3_), .CI(u5_mult_87_SUMB_16__4_), .CO(
        u5_mult_87_CARRYB_17__3_), .S(u5_mult_87_SUMB_17__3_) );
  FA_X1 u5_mult_87_S2_17_2 ( .A(u5_mult_87_ab_17__2_), .B(
        u5_mult_87_CARRYB_16__2_), .CI(u5_mult_87_SUMB_16__3_), .CO(
        u5_mult_87_CARRYB_17__2_), .S(u5_mult_87_SUMB_17__2_) );
  FA_X1 u5_mult_87_S2_17_1 ( .A(u5_mult_87_ab_17__1_), .B(
        u5_mult_87_CARRYB_16__1_), .CI(u5_mult_87_SUMB_16__2_), .CO(
        u5_mult_87_CARRYB_17__1_), .S(u5_mult_87_SUMB_17__1_) );
  FA_X1 u5_mult_87_S1_17_0 ( .A(u5_mult_87_ab_17__0_), .B(
        u5_mult_87_CARRYB_16__0_), .CI(u5_mult_87_SUMB_16__1_), .CO(
        u5_mult_87_CARRYB_17__0_), .S(u5_N17) );
  FA_X1 u5_mult_87_S3_18_51 ( .A(u5_mult_87_ab_18__51_), .B(
        u5_mult_87_CARRYB_17__51_), .CI(u5_mult_87_ab_17__52_), .CO(
        u5_mult_87_CARRYB_18__51_), .S(u5_mult_87_SUMB_18__51_) );
  FA_X1 u5_mult_87_S2_18_50 ( .A(u5_mult_87_ab_18__50_), .B(
        u5_mult_87_CARRYB_17__50_), .CI(u5_mult_87_SUMB_17__51_), .CO(
        u5_mult_87_CARRYB_18__50_), .S(u5_mult_87_SUMB_18__50_) );
  FA_X1 u5_mult_87_S2_18_49 ( .A(u5_mult_87_ab_18__49_), .B(
        u5_mult_87_CARRYB_17__49_), .CI(u5_mult_87_SUMB_17__50_), .CO(
        u5_mult_87_CARRYB_18__49_), .S(u5_mult_87_SUMB_18__49_) );
  FA_X1 u5_mult_87_S2_18_48 ( .A(u5_mult_87_ab_18__48_), .B(
        u5_mult_87_CARRYB_17__48_), .CI(u5_mult_87_SUMB_17__49_), .CO(
        u5_mult_87_CARRYB_18__48_), .S(u5_mult_87_SUMB_18__48_) );
  FA_X1 u5_mult_87_S2_18_47 ( .A(u5_mult_87_ab_18__47_), .B(
        u5_mult_87_CARRYB_17__47_), .CI(u5_mult_87_SUMB_17__48_), .CO(
        u5_mult_87_CARRYB_18__47_), .S(u5_mult_87_SUMB_18__47_) );
  FA_X1 u5_mult_87_S2_18_46 ( .A(u5_mult_87_ab_18__46_), .B(
        u5_mult_87_CARRYB_17__46_), .CI(u5_mult_87_SUMB_17__47_), .CO(
        u5_mult_87_CARRYB_18__46_), .S(u5_mult_87_SUMB_18__46_) );
  FA_X1 u5_mult_87_S2_18_45 ( .A(u5_mult_87_ab_18__45_), .B(
        u5_mult_87_CARRYB_17__45_), .CI(u5_mult_87_SUMB_17__46_), .CO(
        u5_mult_87_CARRYB_18__45_), .S(u5_mult_87_SUMB_18__45_) );
  FA_X1 u5_mult_87_S2_18_44 ( .A(u5_mult_87_ab_18__44_), .B(
        u5_mult_87_CARRYB_17__44_), .CI(u5_mult_87_SUMB_17__45_), .CO(
        u5_mult_87_CARRYB_18__44_), .S(u5_mult_87_SUMB_18__44_) );
  FA_X1 u5_mult_87_S2_18_43 ( .A(u5_mult_87_ab_18__43_), .B(
        u5_mult_87_CARRYB_17__43_), .CI(u5_mult_87_SUMB_17__44_), .CO(
        u5_mult_87_CARRYB_18__43_), .S(u5_mult_87_SUMB_18__43_) );
  FA_X1 u5_mult_87_S2_18_42 ( .A(u5_mult_87_ab_18__42_), .B(
        u5_mult_87_CARRYB_17__42_), .CI(u5_mult_87_SUMB_17__43_), .CO(
        u5_mult_87_CARRYB_18__42_), .S(u5_mult_87_SUMB_18__42_) );
  FA_X1 u5_mult_87_S2_18_41 ( .A(u5_mult_87_ab_18__41_), .B(
        u5_mult_87_CARRYB_17__41_), .CI(u5_mult_87_SUMB_17__42_), .CO(
        u5_mult_87_CARRYB_18__41_), .S(u5_mult_87_SUMB_18__41_) );
  FA_X1 u5_mult_87_S2_18_40 ( .A(u5_mult_87_ab_18__40_), .B(
        u5_mult_87_CARRYB_17__40_), .CI(u5_mult_87_SUMB_17__41_), .CO(
        u5_mult_87_CARRYB_18__40_), .S(u5_mult_87_SUMB_18__40_) );
  FA_X1 u5_mult_87_S2_18_39 ( .A(u5_mult_87_ab_18__39_), .B(
        u5_mult_87_CARRYB_17__39_), .CI(u5_mult_87_SUMB_17__40_), .CO(
        u5_mult_87_CARRYB_18__39_), .S(u5_mult_87_SUMB_18__39_) );
  FA_X1 u5_mult_87_S2_18_38 ( .A(u5_mult_87_ab_18__38_), .B(
        u5_mult_87_CARRYB_17__38_), .CI(u5_mult_87_SUMB_17__39_), .CO(
        u5_mult_87_CARRYB_18__38_), .S(u5_mult_87_SUMB_18__38_) );
  FA_X1 u5_mult_87_S2_18_37 ( .A(u5_mult_87_ab_18__37_), .B(
        u5_mult_87_CARRYB_17__37_), .CI(u5_mult_87_SUMB_17__38_), .CO(
        u5_mult_87_CARRYB_18__37_), .S(u5_mult_87_SUMB_18__37_) );
  FA_X1 u5_mult_87_S2_18_36 ( .A(u5_mult_87_ab_18__36_), .B(
        u5_mult_87_CARRYB_17__36_), .CI(u5_mult_87_SUMB_17__37_), .CO(
        u5_mult_87_CARRYB_18__36_), .S(u5_mult_87_SUMB_18__36_) );
  FA_X1 u5_mult_87_S2_18_35 ( .A(u5_mult_87_ab_18__35_), .B(
        u5_mult_87_CARRYB_17__35_), .CI(u5_mult_87_SUMB_17__36_), .CO(
        u5_mult_87_CARRYB_18__35_), .S(u5_mult_87_SUMB_18__35_) );
  FA_X1 u5_mult_87_S2_18_34 ( .A(u5_mult_87_ab_18__34_), .B(
        u5_mult_87_CARRYB_17__34_), .CI(u5_mult_87_SUMB_17__35_), .CO(
        u5_mult_87_CARRYB_18__34_), .S(u5_mult_87_SUMB_18__34_) );
  FA_X1 u5_mult_87_S2_18_33 ( .A(u5_mult_87_ab_18__33_), .B(
        u5_mult_87_CARRYB_17__33_), .CI(u5_mult_87_SUMB_17__34_), .CO(
        u5_mult_87_CARRYB_18__33_), .S(u5_mult_87_SUMB_18__33_) );
  FA_X1 u5_mult_87_S2_18_32 ( .A(u5_mult_87_ab_18__32_), .B(
        u5_mult_87_CARRYB_17__32_), .CI(u5_mult_87_SUMB_17__33_), .CO(
        u5_mult_87_CARRYB_18__32_), .S(u5_mult_87_SUMB_18__32_) );
  FA_X1 u5_mult_87_S2_18_31 ( .A(u5_mult_87_ab_18__31_), .B(
        u5_mult_87_CARRYB_17__31_), .CI(u5_mult_87_SUMB_17__32_), .CO(
        u5_mult_87_CARRYB_18__31_), .S(u5_mult_87_SUMB_18__31_) );
  FA_X1 u5_mult_87_S2_18_30 ( .A(u5_mult_87_ab_18__30_), .B(
        u5_mult_87_CARRYB_17__30_), .CI(u5_mult_87_SUMB_17__31_), .CO(
        u5_mult_87_CARRYB_18__30_), .S(u5_mult_87_SUMB_18__30_) );
  FA_X1 u5_mult_87_S2_18_29 ( .A(u5_mult_87_ab_18__29_), .B(
        u5_mult_87_CARRYB_17__29_), .CI(u5_mult_87_SUMB_17__30_), .CO(
        u5_mult_87_CARRYB_18__29_), .S(u5_mult_87_SUMB_18__29_) );
  FA_X1 u5_mult_87_S2_18_28 ( .A(u5_mult_87_ab_18__28_), .B(
        u5_mult_87_CARRYB_17__28_), .CI(u5_mult_87_SUMB_17__29_), .CO(
        u5_mult_87_CARRYB_18__28_), .S(u5_mult_87_SUMB_18__28_) );
  FA_X1 u5_mult_87_S2_18_27 ( .A(u5_mult_87_ab_18__27_), .B(
        u5_mult_87_CARRYB_17__27_), .CI(u5_mult_87_SUMB_17__28_), .CO(
        u5_mult_87_CARRYB_18__27_), .S(u5_mult_87_SUMB_18__27_) );
  FA_X1 u5_mult_87_S2_18_26 ( .A(u5_mult_87_ab_18__26_), .B(
        u5_mult_87_CARRYB_17__26_), .CI(u5_mult_87_SUMB_17__27_), .CO(
        u5_mult_87_CARRYB_18__26_), .S(u5_mult_87_SUMB_18__26_) );
  FA_X1 u5_mult_87_S2_18_25 ( .A(u5_mult_87_ab_18__25_), .B(
        u5_mult_87_CARRYB_17__25_), .CI(u5_mult_87_SUMB_17__26_), .CO(
        u5_mult_87_CARRYB_18__25_), .S(u5_mult_87_SUMB_18__25_) );
  FA_X1 u5_mult_87_S2_18_24 ( .A(u5_mult_87_ab_18__24_), .B(
        u5_mult_87_CARRYB_17__24_), .CI(u5_mult_87_SUMB_17__25_), .CO(
        u5_mult_87_CARRYB_18__24_), .S(u5_mult_87_SUMB_18__24_) );
  FA_X1 u5_mult_87_S2_18_23 ( .A(u5_mult_87_ab_18__23_), .B(
        u5_mult_87_CARRYB_17__23_), .CI(u5_mult_87_SUMB_17__24_), .CO(
        u5_mult_87_CARRYB_18__23_), .S(u5_mult_87_SUMB_18__23_) );
  FA_X1 u5_mult_87_S2_18_22 ( .A(u5_mult_87_ab_18__22_), .B(
        u5_mult_87_CARRYB_17__22_), .CI(u5_mult_87_SUMB_17__23_), .CO(
        u5_mult_87_CARRYB_18__22_), .S(u5_mult_87_SUMB_18__22_) );
  FA_X1 u5_mult_87_S2_18_21 ( .A(u5_mult_87_ab_18__21_), .B(
        u5_mult_87_CARRYB_17__21_), .CI(u5_mult_87_SUMB_17__22_), .CO(
        u5_mult_87_CARRYB_18__21_), .S(u5_mult_87_SUMB_18__21_) );
  FA_X1 u5_mult_87_S2_18_20 ( .A(u5_mult_87_ab_18__20_), .B(
        u5_mult_87_CARRYB_17__20_), .CI(u5_mult_87_SUMB_17__21_), .CO(
        u5_mult_87_CARRYB_18__20_), .S(u5_mult_87_SUMB_18__20_) );
  FA_X1 u5_mult_87_S2_18_19 ( .A(u5_mult_87_ab_18__19_), .B(
        u5_mult_87_CARRYB_17__19_), .CI(u5_mult_87_SUMB_17__20_), .CO(
        u5_mult_87_CARRYB_18__19_), .S(u5_mult_87_SUMB_18__19_) );
  FA_X1 u5_mult_87_S2_18_18 ( .A(u5_mult_87_ab_18__18_), .B(
        u5_mult_87_CARRYB_17__18_), .CI(u5_mult_87_SUMB_17__19_), .CO(
        u5_mult_87_CARRYB_18__18_), .S(u5_mult_87_SUMB_18__18_) );
  FA_X1 u5_mult_87_S2_18_17 ( .A(u5_mult_87_ab_18__17_), .B(
        u5_mult_87_CARRYB_17__17_), .CI(u5_mult_87_SUMB_17__18_), .CO(
        u5_mult_87_CARRYB_18__17_), .S(u5_mult_87_SUMB_18__17_) );
  FA_X1 u5_mult_87_S2_18_16 ( .A(u5_mult_87_ab_18__16_), .B(
        u5_mult_87_CARRYB_17__16_), .CI(u5_mult_87_SUMB_17__17_), .CO(
        u5_mult_87_CARRYB_18__16_), .S(u5_mult_87_SUMB_18__16_) );
  FA_X1 u5_mult_87_S2_18_15 ( .A(u5_mult_87_ab_18__15_), .B(
        u5_mult_87_CARRYB_17__15_), .CI(u5_mult_87_SUMB_17__16_), .CO(
        u5_mult_87_CARRYB_18__15_), .S(u5_mult_87_SUMB_18__15_) );
  FA_X1 u5_mult_87_S2_18_14 ( .A(u5_mult_87_ab_18__14_), .B(
        u5_mult_87_CARRYB_17__14_), .CI(u5_mult_87_SUMB_17__15_), .CO(
        u5_mult_87_CARRYB_18__14_), .S(u5_mult_87_SUMB_18__14_) );
  FA_X1 u5_mult_87_S2_18_13 ( .A(u5_mult_87_ab_18__13_), .B(
        u5_mult_87_CARRYB_17__13_), .CI(u5_mult_87_SUMB_17__14_), .CO(
        u5_mult_87_CARRYB_18__13_), .S(u5_mult_87_SUMB_18__13_) );
  FA_X1 u5_mult_87_S2_18_12 ( .A(u5_mult_87_ab_18__12_), .B(
        u5_mult_87_CARRYB_17__12_), .CI(u5_mult_87_SUMB_17__13_), .CO(
        u5_mult_87_CARRYB_18__12_), .S(u5_mult_87_SUMB_18__12_) );
  FA_X1 u5_mult_87_S2_18_11 ( .A(u5_mult_87_ab_18__11_), .B(
        u5_mult_87_CARRYB_17__11_), .CI(u5_mult_87_SUMB_17__12_), .CO(
        u5_mult_87_CARRYB_18__11_), .S(u5_mult_87_SUMB_18__11_) );
  FA_X1 u5_mult_87_S2_18_10 ( .A(u5_mult_87_ab_18__10_), .B(
        u5_mult_87_CARRYB_17__10_), .CI(u5_mult_87_SUMB_17__11_), .CO(
        u5_mult_87_CARRYB_18__10_), .S(u5_mult_87_SUMB_18__10_) );
  FA_X1 u5_mult_87_S2_18_9 ( .A(u5_mult_87_ab_18__9_), .B(
        u5_mult_87_CARRYB_17__9_), .CI(u5_mult_87_SUMB_17__10_), .CO(
        u5_mult_87_CARRYB_18__9_), .S(u5_mult_87_SUMB_18__9_) );
  FA_X1 u5_mult_87_S2_18_8 ( .A(u5_mult_87_ab_18__8_), .B(
        u5_mult_87_CARRYB_17__8_), .CI(u5_mult_87_SUMB_17__9_), .CO(
        u5_mult_87_CARRYB_18__8_), .S(u5_mult_87_SUMB_18__8_) );
  FA_X1 u5_mult_87_S2_18_7 ( .A(u5_mult_87_ab_18__7_), .B(
        u5_mult_87_CARRYB_17__7_), .CI(u5_mult_87_SUMB_17__8_), .CO(
        u5_mult_87_CARRYB_18__7_), .S(u5_mult_87_SUMB_18__7_) );
  FA_X1 u5_mult_87_S2_18_6 ( .A(u5_mult_87_ab_18__6_), .B(
        u5_mult_87_CARRYB_17__6_), .CI(u5_mult_87_SUMB_17__7_), .CO(
        u5_mult_87_CARRYB_18__6_), .S(u5_mult_87_SUMB_18__6_) );
  FA_X1 u5_mult_87_S2_18_5 ( .A(u5_mult_87_ab_18__5_), .B(
        u5_mult_87_CARRYB_17__5_), .CI(u5_mult_87_SUMB_17__6_), .CO(
        u5_mult_87_CARRYB_18__5_), .S(u5_mult_87_SUMB_18__5_) );
  FA_X1 u5_mult_87_S2_18_4 ( .A(u5_mult_87_ab_18__4_), .B(
        u5_mult_87_CARRYB_17__4_), .CI(u5_mult_87_SUMB_17__5_), .CO(
        u5_mult_87_CARRYB_18__4_), .S(u5_mult_87_SUMB_18__4_) );
  FA_X1 u5_mult_87_S2_18_3 ( .A(u5_mult_87_ab_18__3_), .B(
        u5_mult_87_CARRYB_17__3_), .CI(u5_mult_87_SUMB_17__4_), .CO(
        u5_mult_87_CARRYB_18__3_), .S(u5_mult_87_SUMB_18__3_) );
  FA_X1 u5_mult_87_S2_18_2 ( .A(u5_mult_87_ab_18__2_), .B(
        u5_mult_87_CARRYB_17__2_), .CI(u5_mult_87_SUMB_17__3_), .CO(
        u5_mult_87_CARRYB_18__2_), .S(u5_mult_87_SUMB_18__2_) );
  FA_X1 u5_mult_87_S2_18_1 ( .A(u5_mult_87_ab_18__1_), .B(
        u5_mult_87_CARRYB_17__1_), .CI(u5_mult_87_SUMB_17__2_), .CO(
        u5_mult_87_CARRYB_18__1_), .S(u5_mult_87_SUMB_18__1_) );
  FA_X1 u5_mult_87_S1_18_0 ( .A(u5_mult_87_ab_18__0_), .B(
        u5_mult_87_CARRYB_17__0_), .CI(u5_mult_87_SUMB_17__1_), .CO(
        u5_mult_87_CARRYB_18__0_), .S(u5_N18) );
  FA_X1 u5_mult_87_S3_19_51 ( .A(u5_mult_87_ab_19__51_), .B(
        u5_mult_87_CARRYB_18__51_), .CI(u5_mult_87_ab_18__52_), .CO(
        u5_mult_87_CARRYB_19__51_), .S(u5_mult_87_SUMB_19__51_) );
  FA_X1 u5_mult_87_S2_19_50 ( .A(u5_mult_87_ab_19__50_), .B(
        u5_mult_87_CARRYB_18__50_), .CI(u5_mult_87_SUMB_18__51_), .CO(
        u5_mult_87_CARRYB_19__50_), .S(u5_mult_87_SUMB_19__50_) );
  FA_X1 u5_mult_87_S2_19_49 ( .A(u5_mult_87_ab_19__49_), .B(
        u5_mult_87_CARRYB_18__49_), .CI(u5_mult_87_SUMB_18__50_), .CO(
        u5_mult_87_CARRYB_19__49_), .S(u5_mult_87_SUMB_19__49_) );
  FA_X1 u5_mult_87_S2_19_48 ( .A(u5_mult_87_ab_19__48_), .B(
        u5_mult_87_CARRYB_18__48_), .CI(u5_mult_87_SUMB_18__49_), .CO(
        u5_mult_87_CARRYB_19__48_), .S(u5_mult_87_SUMB_19__48_) );
  FA_X1 u5_mult_87_S2_19_47 ( .A(u5_mult_87_ab_19__47_), .B(
        u5_mult_87_CARRYB_18__47_), .CI(u5_mult_87_SUMB_18__48_), .CO(
        u5_mult_87_CARRYB_19__47_), .S(u5_mult_87_SUMB_19__47_) );
  FA_X1 u5_mult_87_S2_19_46 ( .A(u5_mult_87_ab_19__46_), .B(
        u5_mult_87_CARRYB_18__46_), .CI(u5_mult_87_SUMB_18__47_), .CO(
        u5_mult_87_CARRYB_19__46_), .S(u5_mult_87_SUMB_19__46_) );
  FA_X1 u5_mult_87_S2_19_45 ( .A(u5_mult_87_ab_19__45_), .B(
        u5_mult_87_CARRYB_18__45_), .CI(u5_mult_87_SUMB_18__46_), .CO(
        u5_mult_87_CARRYB_19__45_), .S(u5_mult_87_SUMB_19__45_) );
  FA_X1 u5_mult_87_S2_19_44 ( .A(u5_mult_87_ab_19__44_), .B(
        u5_mult_87_CARRYB_18__44_), .CI(u5_mult_87_SUMB_18__45_), .CO(
        u5_mult_87_CARRYB_19__44_), .S(u5_mult_87_SUMB_19__44_) );
  FA_X1 u5_mult_87_S2_19_43 ( .A(u5_mult_87_ab_19__43_), .B(
        u5_mult_87_CARRYB_18__43_), .CI(u5_mult_87_SUMB_18__44_), .CO(
        u5_mult_87_CARRYB_19__43_), .S(u5_mult_87_SUMB_19__43_) );
  FA_X1 u5_mult_87_S2_19_42 ( .A(u5_mult_87_ab_19__42_), .B(
        u5_mult_87_CARRYB_18__42_), .CI(u5_mult_87_SUMB_18__43_), .CO(
        u5_mult_87_CARRYB_19__42_), .S(u5_mult_87_SUMB_19__42_) );
  FA_X1 u5_mult_87_S2_19_41 ( .A(u5_mult_87_ab_19__41_), .B(
        u5_mult_87_CARRYB_18__41_), .CI(u5_mult_87_SUMB_18__42_), .CO(
        u5_mult_87_CARRYB_19__41_), .S(u5_mult_87_SUMB_19__41_) );
  FA_X1 u5_mult_87_S2_19_40 ( .A(u5_mult_87_ab_19__40_), .B(
        u5_mult_87_CARRYB_18__40_), .CI(u5_mult_87_SUMB_18__41_), .CO(
        u5_mult_87_CARRYB_19__40_), .S(u5_mult_87_SUMB_19__40_) );
  FA_X1 u5_mult_87_S2_19_39 ( .A(u5_mult_87_ab_19__39_), .B(
        u5_mult_87_CARRYB_18__39_), .CI(u5_mult_87_SUMB_18__40_), .CO(
        u5_mult_87_CARRYB_19__39_), .S(u5_mult_87_SUMB_19__39_) );
  FA_X1 u5_mult_87_S2_19_38 ( .A(u5_mult_87_ab_19__38_), .B(
        u5_mult_87_CARRYB_18__38_), .CI(u5_mult_87_SUMB_18__39_), .CO(
        u5_mult_87_CARRYB_19__38_), .S(u5_mult_87_SUMB_19__38_) );
  FA_X1 u5_mult_87_S2_19_37 ( .A(u5_mult_87_ab_19__37_), .B(
        u5_mult_87_CARRYB_18__37_), .CI(u5_mult_87_SUMB_18__38_), .CO(
        u5_mult_87_CARRYB_19__37_), .S(u5_mult_87_SUMB_19__37_) );
  FA_X1 u5_mult_87_S2_19_36 ( .A(u5_mult_87_ab_19__36_), .B(
        u5_mult_87_CARRYB_18__36_), .CI(u5_mult_87_SUMB_18__37_), .CO(
        u5_mult_87_CARRYB_19__36_), .S(u5_mult_87_SUMB_19__36_) );
  FA_X1 u5_mult_87_S2_19_35 ( .A(u5_mult_87_ab_19__35_), .B(
        u5_mult_87_CARRYB_18__35_), .CI(u5_mult_87_SUMB_18__36_), .CO(
        u5_mult_87_CARRYB_19__35_), .S(u5_mult_87_SUMB_19__35_) );
  FA_X1 u5_mult_87_S2_19_34 ( .A(u5_mult_87_ab_19__34_), .B(
        u5_mult_87_CARRYB_18__34_), .CI(u5_mult_87_SUMB_18__35_), .CO(
        u5_mult_87_CARRYB_19__34_), .S(u5_mult_87_SUMB_19__34_) );
  FA_X1 u5_mult_87_S2_19_33 ( .A(u5_mult_87_ab_19__33_), .B(
        u5_mult_87_CARRYB_18__33_), .CI(u5_mult_87_SUMB_18__34_), .CO(
        u5_mult_87_CARRYB_19__33_), .S(u5_mult_87_SUMB_19__33_) );
  FA_X1 u5_mult_87_S2_19_32 ( .A(u5_mult_87_ab_19__32_), .B(
        u5_mult_87_CARRYB_18__32_), .CI(u5_mult_87_SUMB_18__33_), .CO(
        u5_mult_87_CARRYB_19__32_), .S(u5_mult_87_SUMB_19__32_) );
  FA_X1 u5_mult_87_S2_19_31 ( .A(u5_mult_87_ab_19__31_), .B(
        u5_mult_87_CARRYB_18__31_), .CI(u5_mult_87_SUMB_18__32_), .CO(
        u5_mult_87_CARRYB_19__31_), .S(u5_mult_87_SUMB_19__31_) );
  FA_X1 u5_mult_87_S2_19_30 ( .A(u5_mult_87_ab_19__30_), .B(
        u5_mult_87_CARRYB_18__30_), .CI(u5_mult_87_SUMB_18__31_), .CO(
        u5_mult_87_CARRYB_19__30_), .S(u5_mult_87_SUMB_19__30_) );
  FA_X1 u5_mult_87_S2_19_29 ( .A(u5_mult_87_ab_19__29_), .B(
        u5_mult_87_CARRYB_18__29_), .CI(u5_mult_87_SUMB_18__30_), .CO(
        u5_mult_87_CARRYB_19__29_), .S(u5_mult_87_SUMB_19__29_) );
  FA_X1 u5_mult_87_S2_19_28 ( .A(u5_mult_87_ab_19__28_), .B(
        u5_mult_87_CARRYB_18__28_), .CI(u5_mult_87_SUMB_18__29_), .CO(
        u5_mult_87_CARRYB_19__28_), .S(u5_mult_87_SUMB_19__28_) );
  FA_X1 u5_mult_87_S2_19_27 ( .A(u5_mult_87_ab_19__27_), .B(
        u5_mult_87_CARRYB_18__27_), .CI(u5_mult_87_SUMB_18__28_), .CO(
        u5_mult_87_CARRYB_19__27_), .S(u5_mult_87_SUMB_19__27_) );
  FA_X1 u5_mult_87_S2_19_26 ( .A(u5_mult_87_ab_19__26_), .B(
        u5_mult_87_CARRYB_18__26_), .CI(u5_mult_87_SUMB_18__27_), .CO(
        u5_mult_87_CARRYB_19__26_), .S(u5_mult_87_SUMB_19__26_) );
  FA_X1 u5_mult_87_S2_19_25 ( .A(u5_mult_87_ab_19__25_), .B(
        u5_mult_87_CARRYB_18__25_), .CI(u5_mult_87_SUMB_18__26_), .CO(
        u5_mult_87_CARRYB_19__25_), .S(u5_mult_87_SUMB_19__25_) );
  FA_X1 u5_mult_87_S2_19_24 ( .A(u5_mult_87_ab_19__24_), .B(
        u5_mult_87_CARRYB_18__24_), .CI(u5_mult_87_SUMB_18__25_), .CO(
        u5_mult_87_CARRYB_19__24_), .S(u5_mult_87_SUMB_19__24_) );
  FA_X1 u5_mult_87_S2_19_23 ( .A(u5_mult_87_ab_19__23_), .B(
        u5_mult_87_CARRYB_18__23_), .CI(u5_mult_87_SUMB_18__24_), .CO(
        u5_mult_87_CARRYB_19__23_), .S(u5_mult_87_SUMB_19__23_) );
  FA_X1 u5_mult_87_S2_19_22 ( .A(u5_mult_87_ab_19__22_), .B(
        u5_mult_87_CARRYB_18__22_), .CI(u5_mult_87_SUMB_18__23_), .CO(
        u5_mult_87_CARRYB_19__22_), .S(u5_mult_87_SUMB_19__22_) );
  FA_X1 u5_mult_87_S2_19_21 ( .A(u5_mult_87_ab_19__21_), .B(
        u5_mult_87_CARRYB_18__21_), .CI(u5_mult_87_SUMB_18__22_), .CO(
        u5_mult_87_CARRYB_19__21_), .S(u5_mult_87_SUMB_19__21_) );
  FA_X1 u5_mult_87_S2_19_20 ( .A(u5_mult_87_ab_19__20_), .B(
        u5_mult_87_CARRYB_18__20_), .CI(u5_mult_87_SUMB_18__21_), .CO(
        u5_mult_87_CARRYB_19__20_), .S(u5_mult_87_SUMB_19__20_) );
  FA_X1 u5_mult_87_S2_19_19 ( .A(u5_mult_87_ab_19__19_), .B(
        u5_mult_87_CARRYB_18__19_), .CI(u5_mult_87_SUMB_18__20_), .CO(
        u5_mult_87_CARRYB_19__19_), .S(u5_mult_87_SUMB_19__19_) );
  FA_X1 u5_mult_87_S2_19_18 ( .A(u5_mult_87_ab_19__18_), .B(
        u5_mult_87_CARRYB_18__18_), .CI(u5_mult_87_SUMB_18__19_), .CO(
        u5_mult_87_CARRYB_19__18_), .S(u5_mult_87_SUMB_19__18_) );
  FA_X1 u5_mult_87_S2_19_17 ( .A(u5_mult_87_ab_19__17_), .B(
        u5_mult_87_CARRYB_18__17_), .CI(u5_mult_87_SUMB_18__18_), .CO(
        u5_mult_87_CARRYB_19__17_), .S(u5_mult_87_SUMB_19__17_) );
  FA_X1 u5_mult_87_S2_19_16 ( .A(u5_mult_87_ab_19__16_), .B(
        u5_mult_87_CARRYB_18__16_), .CI(u5_mult_87_SUMB_18__17_), .CO(
        u5_mult_87_CARRYB_19__16_), .S(u5_mult_87_SUMB_19__16_) );
  FA_X1 u5_mult_87_S2_19_15 ( .A(u5_mult_87_ab_19__15_), .B(
        u5_mult_87_CARRYB_18__15_), .CI(u5_mult_87_SUMB_18__16_), .CO(
        u5_mult_87_CARRYB_19__15_), .S(u5_mult_87_SUMB_19__15_) );
  FA_X1 u5_mult_87_S2_19_14 ( .A(u5_mult_87_ab_19__14_), .B(
        u5_mult_87_CARRYB_18__14_), .CI(u5_mult_87_SUMB_18__15_), .CO(
        u5_mult_87_CARRYB_19__14_), .S(u5_mult_87_SUMB_19__14_) );
  FA_X1 u5_mult_87_S2_19_13 ( .A(u5_mult_87_ab_19__13_), .B(
        u5_mult_87_CARRYB_18__13_), .CI(u5_mult_87_SUMB_18__14_), .CO(
        u5_mult_87_CARRYB_19__13_), .S(u5_mult_87_SUMB_19__13_) );
  FA_X1 u5_mult_87_S2_19_12 ( .A(u5_mult_87_ab_19__12_), .B(
        u5_mult_87_CARRYB_18__12_), .CI(u5_mult_87_SUMB_18__13_), .CO(
        u5_mult_87_CARRYB_19__12_), .S(u5_mult_87_SUMB_19__12_) );
  FA_X1 u5_mult_87_S2_19_11 ( .A(u5_mult_87_ab_19__11_), .B(
        u5_mult_87_CARRYB_18__11_), .CI(u5_mult_87_SUMB_18__12_), .CO(
        u5_mult_87_CARRYB_19__11_), .S(u5_mult_87_SUMB_19__11_) );
  FA_X1 u5_mult_87_S2_19_10 ( .A(u5_mult_87_ab_19__10_), .B(
        u5_mult_87_CARRYB_18__10_), .CI(u5_mult_87_SUMB_18__11_), .CO(
        u5_mult_87_CARRYB_19__10_), .S(u5_mult_87_SUMB_19__10_) );
  FA_X1 u5_mult_87_S2_19_9 ( .A(u5_mult_87_ab_19__9_), .B(
        u5_mult_87_CARRYB_18__9_), .CI(u5_mult_87_SUMB_18__10_), .CO(
        u5_mult_87_CARRYB_19__9_), .S(u5_mult_87_SUMB_19__9_) );
  FA_X1 u5_mult_87_S2_19_8 ( .A(u5_mult_87_ab_19__8_), .B(
        u5_mult_87_CARRYB_18__8_), .CI(u5_mult_87_SUMB_18__9_), .CO(
        u5_mult_87_CARRYB_19__8_), .S(u5_mult_87_SUMB_19__8_) );
  FA_X1 u5_mult_87_S2_19_7 ( .A(u5_mult_87_ab_19__7_), .B(
        u5_mult_87_CARRYB_18__7_), .CI(u5_mult_87_SUMB_18__8_), .CO(
        u5_mult_87_CARRYB_19__7_), .S(u5_mult_87_SUMB_19__7_) );
  FA_X1 u5_mult_87_S2_19_6 ( .A(u5_mult_87_ab_19__6_), .B(
        u5_mult_87_CARRYB_18__6_), .CI(u5_mult_87_SUMB_18__7_), .CO(
        u5_mult_87_CARRYB_19__6_), .S(u5_mult_87_SUMB_19__6_) );
  FA_X1 u5_mult_87_S2_19_5 ( .A(u5_mult_87_ab_19__5_), .B(
        u5_mult_87_CARRYB_18__5_), .CI(u5_mult_87_SUMB_18__6_), .CO(
        u5_mult_87_CARRYB_19__5_), .S(u5_mult_87_SUMB_19__5_) );
  FA_X1 u5_mult_87_S2_19_4 ( .A(u5_mult_87_ab_19__4_), .B(
        u5_mult_87_CARRYB_18__4_), .CI(u5_mult_87_SUMB_18__5_), .CO(
        u5_mult_87_CARRYB_19__4_), .S(u5_mult_87_SUMB_19__4_) );
  FA_X1 u5_mult_87_S2_19_3 ( .A(u5_mult_87_ab_19__3_), .B(
        u5_mult_87_CARRYB_18__3_), .CI(u5_mult_87_SUMB_18__4_), .CO(
        u5_mult_87_CARRYB_19__3_), .S(u5_mult_87_SUMB_19__3_) );
  FA_X1 u5_mult_87_S2_19_2 ( .A(u5_mult_87_ab_19__2_), .B(
        u5_mult_87_CARRYB_18__2_), .CI(u5_mult_87_SUMB_18__3_), .CO(
        u5_mult_87_CARRYB_19__2_), .S(u5_mult_87_SUMB_19__2_) );
  FA_X1 u5_mult_87_S2_19_1 ( .A(u5_mult_87_ab_19__1_), .B(
        u5_mult_87_CARRYB_18__1_), .CI(u5_mult_87_SUMB_18__2_), .CO(
        u5_mult_87_CARRYB_19__1_), .S(u5_mult_87_SUMB_19__1_) );
  FA_X1 u5_mult_87_S1_19_0 ( .A(u5_mult_87_ab_19__0_), .B(
        u5_mult_87_CARRYB_18__0_), .CI(u5_mult_87_SUMB_18__1_), .CO(
        u5_mult_87_CARRYB_19__0_), .S(u5_N19) );
  FA_X1 u5_mult_87_S3_20_51 ( .A(u5_mult_87_ab_20__51_), .B(
        u5_mult_87_CARRYB_19__51_), .CI(u5_mult_87_ab_19__52_), .CO(
        u5_mult_87_CARRYB_20__51_), .S(u5_mult_87_SUMB_20__51_) );
  FA_X1 u5_mult_87_S2_20_50 ( .A(u5_mult_87_ab_20__50_), .B(
        u5_mult_87_CARRYB_19__50_), .CI(u5_mult_87_SUMB_19__51_), .CO(
        u5_mult_87_CARRYB_20__50_), .S(u5_mult_87_SUMB_20__50_) );
  FA_X1 u5_mult_87_S2_20_49 ( .A(u5_mult_87_ab_20__49_), .B(
        u5_mult_87_CARRYB_19__49_), .CI(u5_mult_87_SUMB_19__50_), .CO(
        u5_mult_87_CARRYB_20__49_), .S(u5_mult_87_SUMB_20__49_) );
  FA_X1 u5_mult_87_S2_20_48 ( .A(u5_mult_87_ab_20__48_), .B(
        u5_mult_87_CARRYB_19__48_), .CI(u5_mult_87_SUMB_19__49_), .CO(
        u5_mult_87_CARRYB_20__48_), .S(u5_mult_87_SUMB_20__48_) );
  FA_X1 u5_mult_87_S2_20_47 ( .A(u5_mult_87_ab_20__47_), .B(
        u5_mult_87_CARRYB_19__47_), .CI(u5_mult_87_SUMB_19__48_), .CO(
        u5_mult_87_CARRYB_20__47_), .S(u5_mult_87_SUMB_20__47_) );
  FA_X1 u5_mult_87_S2_20_46 ( .A(u5_mult_87_ab_20__46_), .B(
        u5_mult_87_CARRYB_19__46_), .CI(u5_mult_87_SUMB_19__47_), .CO(
        u5_mult_87_CARRYB_20__46_), .S(u5_mult_87_SUMB_20__46_) );
  FA_X1 u5_mult_87_S2_20_45 ( .A(u5_mult_87_ab_20__45_), .B(
        u5_mult_87_CARRYB_19__45_), .CI(u5_mult_87_SUMB_19__46_), .CO(
        u5_mult_87_CARRYB_20__45_), .S(u5_mult_87_SUMB_20__45_) );
  FA_X1 u5_mult_87_S2_20_44 ( .A(u5_mult_87_ab_20__44_), .B(
        u5_mult_87_CARRYB_19__44_), .CI(u5_mult_87_SUMB_19__45_), .CO(
        u5_mult_87_CARRYB_20__44_), .S(u5_mult_87_SUMB_20__44_) );
  FA_X1 u5_mult_87_S2_20_43 ( .A(u5_mult_87_ab_20__43_), .B(
        u5_mult_87_CARRYB_19__43_), .CI(u5_mult_87_SUMB_19__44_), .CO(
        u5_mult_87_CARRYB_20__43_), .S(u5_mult_87_SUMB_20__43_) );
  FA_X1 u5_mult_87_S2_20_42 ( .A(u5_mult_87_ab_20__42_), .B(
        u5_mult_87_CARRYB_19__42_), .CI(u5_mult_87_SUMB_19__43_), .CO(
        u5_mult_87_CARRYB_20__42_), .S(u5_mult_87_SUMB_20__42_) );
  FA_X1 u5_mult_87_S2_20_41 ( .A(u5_mult_87_ab_20__41_), .B(
        u5_mult_87_CARRYB_19__41_), .CI(u5_mult_87_SUMB_19__42_), .CO(
        u5_mult_87_CARRYB_20__41_), .S(u5_mult_87_SUMB_20__41_) );
  FA_X1 u5_mult_87_S2_20_40 ( .A(u5_mult_87_ab_20__40_), .B(
        u5_mult_87_CARRYB_19__40_), .CI(u5_mult_87_SUMB_19__41_), .CO(
        u5_mult_87_CARRYB_20__40_), .S(u5_mult_87_SUMB_20__40_) );
  FA_X1 u5_mult_87_S2_20_39 ( .A(u5_mult_87_ab_20__39_), .B(
        u5_mult_87_CARRYB_19__39_), .CI(u5_mult_87_SUMB_19__40_), .CO(
        u5_mult_87_CARRYB_20__39_), .S(u5_mult_87_SUMB_20__39_) );
  FA_X1 u5_mult_87_S2_20_38 ( .A(u5_mult_87_ab_20__38_), .B(
        u5_mult_87_CARRYB_19__38_), .CI(u5_mult_87_SUMB_19__39_), .CO(
        u5_mult_87_CARRYB_20__38_), .S(u5_mult_87_SUMB_20__38_) );
  FA_X1 u5_mult_87_S2_20_37 ( .A(u5_mult_87_ab_20__37_), .B(
        u5_mult_87_CARRYB_19__37_), .CI(u5_mult_87_SUMB_19__38_), .CO(
        u5_mult_87_CARRYB_20__37_), .S(u5_mult_87_SUMB_20__37_) );
  FA_X1 u5_mult_87_S2_20_36 ( .A(u5_mult_87_ab_20__36_), .B(
        u5_mult_87_CARRYB_19__36_), .CI(u5_mult_87_SUMB_19__37_), .CO(
        u5_mult_87_CARRYB_20__36_), .S(u5_mult_87_SUMB_20__36_) );
  FA_X1 u5_mult_87_S2_20_35 ( .A(u5_mult_87_ab_20__35_), .B(
        u5_mult_87_CARRYB_19__35_), .CI(u5_mult_87_SUMB_19__36_), .CO(
        u5_mult_87_CARRYB_20__35_), .S(u5_mult_87_SUMB_20__35_) );
  FA_X1 u5_mult_87_S2_20_34 ( .A(u5_mult_87_ab_20__34_), .B(
        u5_mult_87_CARRYB_19__34_), .CI(u5_mult_87_SUMB_19__35_), .CO(
        u5_mult_87_CARRYB_20__34_), .S(u5_mult_87_SUMB_20__34_) );
  FA_X1 u5_mult_87_S2_20_33 ( .A(u5_mult_87_ab_20__33_), .B(
        u5_mult_87_CARRYB_19__33_), .CI(u5_mult_87_SUMB_19__34_), .CO(
        u5_mult_87_CARRYB_20__33_), .S(u5_mult_87_SUMB_20__33_) );
  FA_X1 u5_mult_87_S2_20_32 ( .A(u5_mult_87_ab_20__32_), .B(
        u5_mult_87_CARRYB_19__32_), .CI(u5_mult_87_SUMB_19__33_), .CO(
        u5_mult_87_CARRYB_20__32_), .S(u5_mult_87_SUMB_20__32_) );
  FA_X1 u5_mult_87_S2_20_31 ( .A(u5_mult_87_ab_20__31_), .B(
        u5_mult_87_CARRYB_19__31_), .CI(u5_mult_87_SUMB_19__32_), .CO(
        u5_mult_87_CARRYB_20__31_), .S(u5_mult_87_SUMB_20__31_) );
  FA_X1 u5_mult_87_S2_20_30 ( .A(u5_mult_87_ab_20__30_), .B(
        u5_mult_87_CARRYB_19__30_), .CI(u5_mult_87_SUMB_19__31_), .CO(
        u5_mult_87_CARRYB_20__30_), .S(u5_mult_87_SUMB_20__30_) );
  FA_X1 u5_mult_87_S2_20_29 ( .A(u5_mult_87_ab_20__29_), .B(
        u5_mult_87_CARRYB_19__29_), .CI(u5_mult_87_SUMB_19__30_), .CO(
        u5_mult_87_CARRYB_20__29_), .S(u5_mult_87_SUMB_20__29_) );
  FA_X1 u5_mult_87_S2_20_28 ( .A(u5_mult_87_ab_20__28_), .B(
        u5_mult_87_CARRYB_19__28_), .CI(u5_mult_87_SUMB_19__29_), .CO(
        u5_mult_87_CARRYB_20__28_), .S(u5_mult_87_SUMB_20__28_) );
  FA_X1 u5_mult_87_S2_20_27 ( .A(u5_mult_87_ab_20__27_), .B(
        u5_mult_87_CARRYB_19__27_), .CI(u5_mult_87_SUMB_19__28_), .CO(
        u5_mult_87_CARRYB_20__27_), .S(u5_mult_87_SUMB_20__27_) );
  FA_X1 u5_mult_87_S2_20_26 ( .A(u5_mult_87_ab_20__26_), .B(
        u5_mult_87_CARRYB_19__26_), .CI(u5_mult_87_SUMB_19__27_), .CO(
        u5_mult_87_CARRYB_20__26_), .S(u5_mult_87_SUMB_20__26_) );
  FA_X1 u5_mult_87_S2_20_25 ( .A(u5_mult_87_ab_20__25_), .B(
        u5_mult_87_CARRYB_19__25_), .CI(u5_mult_87_SUMB_19__26_), .CO(
        u5_mult_87_CARRYB_20__25_), .S(u5_mult_87_SUMB_20__25_) );
  FA_X1 u5_mult_87_S2_20_24 ( .A(u5_mult_87_ab_20__24_), .B(
        u5_mult_87_CARRYB_19__24_), .CI(u5_mult_87_SUMB_19__25_), .CO(
        u5_mult_87_CARRYB_20__24_), .S(u5_mult_87_SUMB_20__24_) );
  FA_X1 u5_mult_87_S2_20_23 ( .A(u5_mult_87_ab_20__23_), .B(
        u5_mult_87_CARRYB_19__23_), .CI(u5_mult_87_SUMB_19__24_), .CO(
        u5_mult_87_CARRYB_20__23_), .S(u5_mult_87_SUMB_20__23_) );
  FA_X1 u5_mult_87_S2_20_22 ( .A(u5_mult_87_ab_20__22_), .B(
        u5_mult_87_CARRYB_19__22_), .CI(u5_mult_87_SUMB_19__23_), .CO(
        u5_mult_87_CARRYB_20__22_), .S(u5_mult_87_SUMB_20__22_) );
  FA_X1 u5_mult_87_S2_20_21 ( .A(u5_mult_87_ab_20__21_), .B(
        u5_mult_87_CARRYB_19__21_), .CI(u5_mult_87_SUMB_19__22_), .CO(
        u5_mult_87_CARRYB_20__21_), .S(u5_mult_87_SUMB_20__21_) );
  FA_X1 u5_mult_87_S2_20_20 ( .A(u5_mult_87_ab_20__20_), .B(
        u5_mult_87_CARRYB_19__20_), .CI(u5_mult_87_SUMB_19__21_), .CO(
        u5_mult_87_CARRYB_20__20_), .S(u5_mult_87_SUMB_20__20_) );
  FA_X1 u5_mult_87_S2_20_19 ( .A(u5_mult_87_ab_20__19_), .B(
        u5_mult_87_CARRYB_19__19_), .CI(u5_mult_87_SUMB_19__20_), .CO(
        u5_mult_87_CARRYB_20__19_), .S(u5_mult_87_SUMB_20__19_) );
  FA_X1 u5_mult_87_S2_20_18 ( .A(u5_mult_87_ab_20__18_), .B(
        u5_mult_87_CARRYB_19__18_), .CI(u5_mult_87_SUMB_19__19_), .CO(
        u5_mult_87_CARRYB_20__18_), .S(u5_mult_87_SUMB_20__18_) );
  FA_X1 u5_mult_87_S2_20_17 ( .A(u5_mult_87_ab_20__17_), .B(
        u5_mult_87_CARRYB_19__17_), .CI(u5_mult_87_SUMB_19__18_), .CO(
        u5_mult_87_CARRYB_20__17_), .S(u5_mult_87_SUMB_20__17_) );
  FA_X1 u5_mult_87_S2_20_16 ( .A(u5_mult_87_ab_20__16_), .B(
        u5_mult_87_CARRYB_19__16_), .CI(u5_mult_87_SUMB_19__17_), .CO(
        u5_mult_87_CARRYB_20__16_), .S(u5_mult_87_SUMB_20__16_) );
  FA_X1 u5_mult_87_S2_20_15 ( .A(u5_mult_87_ab_20__15_), .B(
        u5_mult_87_CARRYB_19__15_), .CI(u5_mult_87_SUMB_19__16_), .CO(
        u5_mult_87_CARRYB_20__15_), .S(u5_mult_87_SUMB_20__15_) );
  FA_X1 u5_mult_87_S2_20_14 ( .A(u5_mult_87_ab_20__14_), .B(
        u5_mult_87_CARRYB_19__14_), .CI(u5_mult_87_SUMB_19__15_), .CO(
        u5_mult_87_CARRYB_20__14_), .S(u5_mult_87_SUMB_20__14_) );
  FA_X1 u5_mult_87_S2_20_13 ( .A(u5_mult_87_ab_20__13_), .B(
        u5_mult_87_CARRYB_19__13_), .CI(u5_mult_87_SUMB_19__14_), .CO(
        u5_mult_87_CARRYB_20__13_), .S(u5_mult_87_SUMB_20__13_) );
  FA_X1 u5_mult_87_S2_20_12 ( .A(u5_mult_87_ab_20__12_), .B(
        u5_mult_87_CARRYB_19__12_), .CI(u5_mult_87_SUMB_19__13_), .CO(
        u5_mult_87_CARRYB_20__12_), .S(u5_mult_87_SUMB_20__12_) );
  FA_X1 u5_mult_87_S2_20_11 ( .A(u5_mult_87_ab_20__11_), .B(
        u5_mult_87_CARRYB_19__11_), .CI(u5_mult_87_SUMB_19__12_), .CO(
        u5_mult_87_CARRYB_20__11_), .S(u5_mult_87_SUMB_20__11_) );
  FA_X1 u5_mult_87_S2_20_10 ( .A(u5_mult_87_ab_20__10_), .B(
        u5_mult_87_CARRYB_19__10_), .CI(u5_mult_87_SUMB_19__11_), .CO(
        u5_mult_87_CARRYB_20__10_), .S(u5_mult_87_SUMB_20__10_) );
  FA_X1 u5_mult_87_S2_20_9 ( .A(u5_mult_87_ab_20__9_), .B(
        u5_mult_87_CARRYB_19__9_), .CI(u5_mult_87_SUMB_19__10_), .CO(
        u5_mult_87_CARRYB_20__9_), .S(u5_mult_87_SUMB_20__9_) );
  FA_X1 u5_mult_87_S2_20_8 ( .A(u5_mult_87_ab_20__8_), .B(
        u5_mult_87_CARRYB_19__8_), .CI(u5_mult_87_SUMB_19__9_), .CO(
        u5_mult_87_CARRYB_20__8_), .S(u5_mult_87_SUMB_20__8_) );
  FA_X1 u5_mult_87_S2_20_7 ( .A(u5_mult_87_ab_20__7_), .B(
        u5_mult_87_CARRYB_19__7_), .CI(u5_mult_87_SUMB_19__8_), .CO(
        u5_mult_87_CARRYB_20__7_), .S(u5_mult_87_SUMB_20__7_) );
  FA_X1 u5_mult_87_S2_20_6 ( .A(u5_mult_87_ab_20__6_), .B(
        u5_mult_87_CARRYB_19__6_), .CI(u5_mult_87_SUMB_19__7_), .CO(
        u5_mult_87_CARRYB_20__6_), .S(u5_mult_87_SUMB_20__6_) );
  FA_X1 u5_mult_87_S2_20_5 ( .A(u5_mult_87_ab_20__5_), .B(
        u5_mult_87_CARRYB_19__5_), .CI(u5_mult_87_SUMB_19__6_), .CO(
        u5_mult_87_CARRYB_20__5_), .S(u5_mult_87_SUMB_20__5_) );
  FA_X1 u5_mult_87_S2_20_4 ( .A(u5_mult_87_ab_20__4_), .B(
        u5_mult_87_CARRYB_19__4_), .CI(u5_mult_87_SUMB_19__5_), .CO(
        u5_mult_87_CARRYB_20__4_), .S(u5_mult_87_SUMB_20__4_) );
  FA_X1 u5_mult_87_S2_20_3 ( .A(u5_mult_87_ab_20__3_), .B(
        u5_mult_87_CARRYB_19__3_), .CI(u5_mult_87_SUMB_19__4_), .CO(
        u5_mult_87_CARRYB_20__3_), .S(u5_mult_87_SUMB_20__3_) );
  FA_X1 u5_mult_87_S2_20_2 ( .A(u5_mult_87_ab_20__2_), .B(
        u5_mult_87_CARRYB_19__2_), .CI(u5_mult_87_SUMB_19__3_), .CO(
        u5_mult_87_CARRYB_20__2_), .S(u5_mult_87_SUMB_20__2_) );
  FA_X1 u5_mult_87_S2_20_1 ( .A(u5_mult_87_ab_20__1_), .B(
        u5_mult_87_CARRYB_19__1_), .CI(u5_mult_87_SUMB_19__2_), .CO(
        u5_mult_87_CARRYB_20__1_), .S(u5_mult_87_SUMB_20__1_) );
  FA_X1 u5_mult_87_S1_20_0 ( .A(u5_mult_87_ab_20__0_), .B(
        u5_mult_87_CARRYB_19__0_), .CI(u5_mult_87_SUMB_19__1_), .CO(
        u5_mult_87_CARRYB_20__0_), .S(u5_N20) );
  FA_X1 u5_mult_87_S3_21_51 ( .A(u5_mult_87_ab_21__51_), .B(
        u5_mult_87_CARRYB_20__51_), .CI(u5_mult_87_ab_20__52_), .CO(
        u5_mult_87_CARRYB_21__51_), .S(u5_mult_87_SUMB_21__51_) );
  FA_X1 u5_mult_87_S2_21_50 ( .A(u5_mult_87_ab_21__50_), .B(
        u5_mult_87_CARRYB_20__50_), .CI(u5_mult_87_SUMB_20__51_), .CO(
        u5_mult_87_CARRYB_21__50_), .S(u5_mult_87_SUMB_21__50_) );
  FA_X1 u5_mult_87_S2_21_49 ( .A(u5_mult_87_ab_21__49_), .B(
        u5_mult_87_CARRYB_20__49_), .CI(u5_mult_87_SUMB_20__50_), .CO(
        u5_mult_87_CARRYB_21__49_), .S(u5_mult_87_SUMB_21__49_) );
  FA_X1 u5_mult_87_S2_21_48 ( .A(u5_mult_87_ab_21__48_), .B(
        u5_mult_87_CARRYB_20__48_), .CI(u5_mult_87_SUMB_20__49_), .CO(
        u5_mult_87_CARRYB_21__48_), .S(u5_mult_87_SUMB_21__48_) );
  FA_X1 u5_mult_87_S2_21_47 ( .A(u5_mult_87_ab_21__47_), .B(
        u5_mult_87_CARRYB_20__47_), .CI(u5_mult_87_SUMB_20__48_), .CO(
        u5_mult_87_CARRYB_21__47_), .S(u5_mult_87_SUMB_21__47_) );
  FA_X1 u5_mult_87_S2_21_46 ( .A(u5_mult_87_ab_21__46_), .B(
        u5_mult_87_CARRYB_20__46_), .CI(u5_mult_87_SUMB_20__47_), .CO(
        u5_mult_87_CARRYB_21__46_), .S(u5_mult_87_SUMB_21__46_) );
  FA_X1 u5_mult_87_S2_21_45 ( .A(u5_mult_87_ab_21__45_), .B(
        u5_mult_87_CARRYB_20__45_), .CI(u5_mult_87_SUMB_20__46_), .CO(
        u5_mult_87_CARRYB_21__45_), .S(u5_mult_87_SUMB_21__45_) );
  FA_X1 u5_mult_87_S2_21_44 ( .A(u5_mult_87_ab_21__44_), .B(
        u5_mult_87_CARRYB_20__44_), .CI(u5_mult_87_SUMB_20__45_), .CO(
        u5_mult_87_CARRYB_21__44_), .S(u5_mult_87_SUMB_21__44_) );
  FA_X1 u5_mult_87_S2_21_43 ( .A(u5_mult_87_ab_21__43_), .B(
        u5_mult_87_CARRYB_20__43_), .CI(u5_mult_87_SUMB_20__44_), .CO(
        u5_mult_87_CARRYB_21__43_), .S(u5_mult_87_SUMB_21__43_) );
  FA_X1 u5_mult_87_S2_21_42 ( .A(u5_mult_87_ab_21__42_), .B(
        u5_mult_87_CARRYB_20__42_), .CI(u5_mult_87_SUMB_20__43_), .CO(
        u5_mult_87_CARRYB_21__42_), .S(u5_mult_87_SUMB_21__42_) );
  FA_X1 u5_mult_87_S2_21_41 ( .A(u5_mult_87_ab_21__41_), .B(
        u5_mult_87_CARRYB_20__41_), .CI(u5_mult_87_SUMB_20__42_), .CO(
        u5_mult_87_CARRYB_21__41_), .S(u5_mult_87_SUMB_21__41_) );
  FA_X1 u5_mult_87_S2_21_40 ( .A(u5_mult_87_ab_21__40_), .B(
        u5_mult_87_CARRYB_20__40_), .CI(u5_mult_87_SUMB_20__41_), .CO(
        u5_mult_87_CARRYB_21__40_), .S(u5_mult_87_SUMB_21__40_) );
  FA_X1 u5_mult_87_S2_21_39 ( .A(u5_mult_87_ab_21__39_), .B(
        u5_mult_87_CARRYB_20__39_), .CI(u5_mult_87_SUMB_20__40_), .CO(
        u5_mult_87_CARRYB_21__39_), .S(u5_mult_87_SUMB_21__39_) );
  FA_X1 u5_mult_87_S2_21_38 ( .A(u5_mult_87_ab_21__38_), .B(
        u5_mult_87_CARRYB_20__38_), .CI(u5_mult_87_SUMB_20__39_), .CO(
        u5_mult_87_CARRYB_21__38_), .S(u5_mult_87_SUMB_21__38_) );
  FA_X1 u5_mult_87_S2_21_37 ( .A(u5_mult_87_ab_21__37_), .B(
        u5_mult_87_CARRYB_20__37_), .CI(u5_mult_87_SUMB_20__38_), .CO(
        u5_mult_87_CARRYB_21__37_), .S(u5_mult_87_SUMB_21__37_) );
  FA_X1 u5_mult_87_S2_21_36 ( .A(u5_mult_87_ab_21__36_), .B(
        u5_mult_87_CARRYB_20__36_), .CI(u5_mult_87_SUMB_20__37_), .CO(
        u5_mult_87_CARRYB_21__36_), .S(u5_mult_87_SUMB_21__36_) );
  FA_X1 u5_mult_87_S2_21_35 ( .A(u5_mult_87_ab_21__35_), .B(
        u5_mult_87_CARRYB_20__35_), .CI(u5_mult_87_SUMB_20__36_), .CO(
        u5_mult_87_CARRYB_21__35_), .S(u5_mult_87_SUMB_21__35_) );
  FA_X1 u5_mult_87_S2_21_34 ( .A(u5_mult_87_ab_21__34_), .B(
        u5_mult_87_CARRYB_20__34_), .CI(u5_mult_87_SUMB_20__35_), .CO(
        u5_mult_87_CARRYB_21__34_), .S(u5_mult_87_SUMB_21__34_) );
  FA_X1 u5_mult_87_S2_21_33 ( .A(u5_mult_87_ab_21__33_), .B(
        u5_mult_87_CARRYB_20__33_), .CI(u5_mult_87_SUMB_20__34_), .CO(
        u5_mult_87_CARRYB_21__33_), .S(u5_mult_87_SUMB_21__33_) );
  FA_X1 u5_mult_87_S2_21_32 ( .A(u5_mult_87_ab_21__32_), .B(
        u5_mult_87_CARRYB_20__32_), .CI(u5_mult_87_SUMB_20__33_), .CO(
        u5_mult_87_CARRYB_21__32_), .S(u5_mult_87_SUMB_21__32_) );
  FA_X1 u5_mult_87_S2_21_31 ( .A(u5_mult_87_ab_21__31_), .B(
        u5_mult_87_CARRYB_20__31_), .CI(u5_mult_87_SUMB_20__32_), .CO(
        u5_mult_87_CARRYB_21__31_), .S(u5_mult_87_SUMB_21__31_) );
  FA_X1 u5_mult_87_S2_21_30 ( .A(u5_mult_87_ab_21__30_), .B(
        u5_mult_87_CARRYB_20__30_), .CI(u5_mult_87_SUMB_20__31_), .CO(
        u5_mult_87_CARRYB_21__30_), .S(u5_mult_87_SUMB_21__30_) );
  FA_X1 u5_mult_87_S2_21_29 ( .A(u5_mult_87_ab_21__29_), .B(
        u5_mult_87_CARRYB_20__29_), .CI(u5_mult_87_SUMB_20__30_), .CO(
        u5_mult_87_CARRYB_21__29_), .S(u5_mult_87_SUMB_21__29_) );
  FA_X1 u5_mult_87_S2_21_28 ( .A(u5_mult_87_ab_21__28_), .B(
        u5_mult_87_CARRYB_20__28_), .CI(u5_mult_87_SUMB_20__29_), .CO(
        u5_mult_87_CARRYB_21__28_), .S(u5_mult_87_SUMB_21__28_) );
  FA_X1 u5_mult_87_S2_21_27 ( .A(u5_mult_87_ab_21__27_), .B(
        u5_mult_87_CARRYB_20__27_), .CI(u5_mult_87_SUMB_20__28_), .CO(
        u5_mult_87_CARRYB_21__27_), .S(u5_mult_87_SUMB_21__27_) );
  FA_X1 u5_mult_87_S2_21_26 ( .A(u5_mult_87_ab_21__26_), .B(
        u5_mult_87_CARRYB_20__26_), .CI(u5_mult_87_SUMB_20__27_), .CO(
        u5_mult_87_CARRYB_21__26_), .S(u5_mult_87_SUMB_21__26_) );
  FA_X1 u5_mult_87_S2_21_25 ( .A(u5_mult_87_ab_21__25_), .B(
        u5_mult_87_CARRYB_20__25_), .CI(u5_mult_87_SUMB_20__26_), .CO(
        u5_mult_87_CARRYB_21__25_), .S(u5_mult_87_SUMB_21__25_) );
  FA_X1 u5_mult_87_S2_21_24 ( .A(u5_mult_87_ab_21__24_), .B(
        u5_mult_87_CARRYB_20__24_), .CI(u5_mult_87_SUMB_20__25_), .CO(
        u5_mult_87_CARRYB_21__24_), .S(u5_mult_87_SUMB_21__24_) );
  FA_X1 u5_mult_87_S2_21_23 ( .A(u5_mult_87_ab_21__23_), .B(
        u5_mult_87_CARRYB_20__23_), .CI(u5_mult_87_SUMB_20__24_), .CO(
        u5_mult_87_CARRYB_21__23_), .S(u5_mult_87_SUMB_21__23_) );
  FA_X1 u5_mult_87_S2_21_22 ( .A(u5_mult_87_ab_21__22_), .B(
        u5_mult_87_CARRYB_20__22_), .CI(u5_mult_87_SUMB_20__23_), .CO(
        u5_mult_87_CARRYB_21__22_), .S(u5_mult_87_SUMB_21__22_) );
  FA_X1 u5_mult_87_S2_21_21 ( .A(u5_mult_87_ab_21__21_), .B(
        u5_mult_87_CARRYB_20__21_), .CI(u5_mult_87_SUMB_20__22_), .CO(
        u5_mult_87_CARRYB_21__21_), .S(u5_mult_87_SUMB_21__21_) );
  FA_X1 u5_mult_87_S2_21_20 ( .A(u5_mult_87_ab_21__20_), .B(
        u5_mult_87_CARRYB_20__20_), .CI(u5_mult_87_SUMB_20__21_), .CO(
        u5_mult_87_CARRYB_21__20_), .S(u5_mult_87_SUMB_21__20_) );
  FA_X1 u5_mult_87_S2_21_19 ( .A(u5_mult_87_ab_21__19_), .B(
        u5_mult_87_CARRYB_20__19_), .CI(u5_mult_87_SUMB_20__20_), .CO(
        u5_mult_87_CARRYB_21__19_), .S(u5_mult_87_SUMB_21__19_) );
  FA_X1 u5_mult_87_S2_21_18 ( .A(u5_mult_87_ab_21__18_), .B(
        u5_mult_87_CARRYB_20__18_), .CI(u5_mult_87_SUMB_20__19_), .CO(
        u5_mult_87_CARRYB_21__18_), .S(u5_mult_87_SUMB_21__18_) );
  FA_X1 u5_mult_87_S2_21_17 ( .A(u5_mult_87_ab_21__17_), .B(
        u5_mult_87_CARRYB_20__17_), .CI(u5_mult_87_SUMB_20__18_), .CO(
        u5_mult_87_CARRYB_21__17_), .S(u5_mult_87_SUMB_21__17_) );
  FA_X1 u5_mult_87_S2_21_16 ( .A(u5_mult_87_ab_21__16_), .B(
        u5_mult_87_CARRYB_20__16_), .CI(u5_mult_87_SUMB_20__17_), .CO(
        u5_mult_87_CARRYB_21__16_), .S(u5_mult_87_SUMB_21__16_) );
  FA_X1 u5_mult_87_S2_21_15 ( .A(u5_mult_87_ab_21__15_), .B(
        u5_mult_87_CARRYB_20__15_), .CI(u5_mult_87_SUMB_20__16_), .CO(
        u5_mult_87_CARRYB_21__15_), .S(u5_mult_87_SUMB_21__15_) );
  FA_X1 u5_mult_87_S2_21_14 ( .A(u5_mult_87_ab_21__14_), .B(
        u5_mult_87_CARRYB_20__14_), .CI(u5_mult_87_SUMB_20__15_), .CO(
        u5_mult_87_CARRYB_21__14_), .S(u5_mult_87_SUMB_21__14_) );
  FA_X1 u5_mult_87_S2_21_13 ( .A(u5_mult_87_ab_21__13_), .B(
        u5_mult_87_CARRYB_20__13_), .CI(u5_mult_87_SUMB_20__14_), .CO(
        u5_mult_87_CARRYB_21__13_), .S(u5_mult_87_SUMB_21__13_) );
  FA_X1 u5_mult_87_S2_21_12 ( .A(u5_mult_87_ab_21__12_), .B(
        u5_mult_87_CARRYB_20__12_), .CI(u5_mult_87_SUMB_20__13_), .CO(
        u5_mult_87_CARRYB_21__12_), .S(u5_mult_87_SUMB_21__12_) );
  FA_X1 u5_mult_87_S2_21_11 ( .A(u5_mult_87_ab_21__11_), .B(
        u5_mult_87_CARRYB_20__11_), .CI(u5_mult_87_SUMB_20__12_), .CO(
        u5_mult_87_CARRYB_21__11_), .S(u5_mult_87_SUMB_21__11_) );
  FA_X1 u5_mult_87_S2_21_10 ( .A(u5_mult_87_ab_21__10_), .B(
        u5_mult_87_CARRYB_20__10_), .CI(u5_mult_87_SUMB_20__11_), .CO(
        u5_mult_87_CARRYB_21__10_), .S(u5_mult_87_SUMB_21__10_) );
  FA_X1 u5_mult_87_S2_21_9 ( .A(u5_mult_87_ab_21__9_), .B(
        u5_mult_87_CARRYB_20__9_), .CI(u5_mult_87_SUMB_20__10_), .CO(
        u5_mult_87_CARRYB_21__9_), .S(u5_mult_87_SUMB_21__9_) );
  FA_X1 u5_mult_87_S2_21_8 ( .A(u5_mult_87_ab_21__8_), .B(
        u5_mult_87_CARRYB_20__8_), .CI(u5_mult_87_SUMB_20__9_), .CO(
        u5_mult_87_CARRYB_21__8_), .S(u5_mult_87_SUMB_21__8_) );
  FA_X1 u5_mult_87_S2_21_7 ( .A(u5_mult_87_ab_21__7_), .B(
        u5_mult_87_CARRYB_20__7_), .CI(u5_mult_87_SUMB_20__8_), .CO(
        u5_mult_87_CARRYB_21__7_), .S(u5_mult_87_SUMB_21__7_) );
  FA_X1 u5_mult_87_S2_21_6 ( .A(u5_mult_87_ab_21__6_), .B(
        u5_mult_87_CARRYB_20__6_), .CI(u5_mult_87_SUMB_20__7_), .CO(
        u5_mult_87_CARRYB_21__6_), .S(u5_mult_87_SUMB_21__6_) );
  FA_X1 u5_mult_87_S2_21_5 ( .A(u5_mult_87_ab_21__5_), .B(
        u5_mult_87_CARRYB_20__5_), .CI(u5_mult_87_SUMB_20__6_), .CO(
        u5_mult_87_CARRYB_21__5_), .S(u5_mult_87_SUMB_21__5_) );
  FA_X1 u5_mult_87_S2_21_4 ( .A(u5_mult_87_ab_21__4_), .B(
        u5_mult_87_CARRYB_20__4_), .CI(u5_mult_87_SUMB_20__5_), .CO(
        u5_mult_87_CARRYB_21__4_), .S(u5_mult_87_SUMB_21__4_) );
  FA_X1 u5_mult_87_S2_21_3 ( .A(u5_mult_87_ab_21__3_), .B(
        u5_mult_87_CARRYB_20__3_), .CI(u5_mult_87_SUMB_20__4_), .CO(
        u5_mult_87_CARRYB_21__3_), .S(u5_mult_87_SUMB_21__3_) );
  FA_X1 u5_mult_87_S2_21_2 ( .A(u5_mult_87_ab_21__2_), .B(
        u5_mult_87_CARRYB_20__2_), .CI(u5_mult_87_SUMB_20__3_), .CO(
        u5_mult_87_CARRYB_21__2_), .S(u5_mult_87_SUMB_21__2_) );
  FA_X1 u5_mult_87_S2_21_1 ( .A(u5_mult_87_ab_21__1_), .B(
        u5_mult_87_CARRYB_20__1_), .CI(u5_mult_87_SUMB_20__2_), .CO(
        u5_mult_87_CARRYB_21__1_), .S(u5_mult_87_SUMB_21__1_) );
  FA_X1 u5_mult_87_S1_21_0 ( .A(u5_mult_87_ab_21__0_), .B(
        u5_mult_87_CARRYB_20__0_), .CI(u5_mult_87_SUMB_20__1_), .CO(
        u5_mult_87_CARRYB_21__0_), .S(u5_N21) );
  FA_X1 u5_mult_87_S3_22_51 ( .A(u5_mult_87_ab_22__51_), .B(
        u5_mult_87_CARRYB_21__51_), .CI(u5_mult_87_ab_21__52_), .CO(
        u5_mult_87_CARRYB_22__51_), .S(u5_mult_87_SUMB_22__51_) );
  FA_X1 u5_mult_87_S2_22_50 ( .A(u5_mult_87_ab_22__50_), .B(
        u5_mult_87_CARRYB_21__50_), .CI(u5_mult_87_SUMB_21__51_), .CO(
        u5_mult_87_CARRYB_22__50_), .S(u5_mult_87_SUMB_22__50_) );
  FA_X1 u5_mult_87_S2_22_49 ( .A(u5_mult_87_ab_22__49_), .B(
        u5_mult_87_CARRYB_21__49_), .CI(u5_mult_87_SUMB_21__50_), .CO(
        u5_mult_87_CARRYB_22__49_), .S(u5_mult_87_SUMB_22__49_) );
  FA_X1 u5_mult_87_S2_22_48 ( .A(u5_mult_87_ab_22__48_), .B(
        u5_mult_87_CARRYB_21__48_), .CI(u5_mult_87_SUMB_21__49_), .CO(
        u5_mult_87_CARRYB_22__48_), .S(u5_mult_87_SUMB_22__48_) );
  FA_X1 u5_mult_87_S2_22_47 ( .A(u5_mult_87_ab_22__47_), .B(
        u5_mult_87_CARRYB_21__47_), .CI(u5_mult_87_SUMB_21__48_), .CO(
        u5_mult_87_CARRYB_22__47_), .S(u5_mult_87_SUMB_22__47_) );
  FA_X1 u5_mult_87_S2_22_46 ( .A(u5_mult_87_ab_22__46_), .B(
        u5_mult_87_CARRYB_21__46_), .CI(u5_mult_87_SUMB_21__47_), .CO(
        u5_mult_87_CARRYB_22__46_), .S(u5_mult_87_SUMB_22__46_) );
  FA_X1 u5_mult_87_S2_22_45 ( .A(u5_mult_87_ab_22__45_), .B(
        u5_mult_87_CARRYB_21__45_), .CI(u5_mult_87_SUMB_21__46_), .CO(
        u5_mult_87_CARRYB_22__45_), .S(u5_mult_87_SUMB_22__45_) );
  FA_X1 u5_mult_87_S2_22_44 ( .A(u5_mult_87_ab_22__44_), .B(
        u5_mult_87_CARRYB_21__44_), .CI(u5_mult_87_SUMB_21__45_), .CO(
        u5_mult_87_CARRYB_22__44_), .S(u5_mult_87_SUMB_22__44_) );
  FA_X1 u5_mult_87_S2_22_43 ( .A(u5_mult_87_ab_22__43_), .B(
        u5_mult_87_CARRYB_21__43_), .CI(u5_mult_87_SUMB_21__44_), .CO(
        u5_mult_87_CARRYB_22__43_), .S(u5_mult_87_SUMB_22__43_) );
  FA_X1 u5_mult_87_S2_22_42 ( .A(u5_mult_87_ab_22__42_), .B(
        u5_mult_87_CARRYB_21__42_), .CI(u5_mult_87_SUMB_21__43_), .CO(
        u5_mult_87_CARRYB_22__42_), .S(u5_mult_87_SUMB_22__42_) );
  FA_X1 u5_mult_87_S2_22_41 ( .A(u5_mult_87_ab_22__41_), .B(
        u5_mult_87_CARRYB_21__41_), .CI(u5_mult_87_SUMB_21__42_), .CO(
        u5_mult_87_CARRYB_22__41_), .S(u5_mult_87_SUMB_22__41_) );
  FA_X1 u5_mult_87_S2_22_40 ( .A(u5_mult_87_ab_22__40_), .B(
        u5_mult_87_CARRYB_21__40_), .CI(u5_mult_87_SUMB_21__41_), .CO(
        u5_mult_87_CARRYB_22__40_), .S(u5_mult_87_SUMB_22__40_) );
  FA_X1 u5_mult_87_S2_22_39 ( .A(u5_mult_87_ab_22__39_), .B(
        u5_mult_87_CARRYB_21__39_), .CI(u5_mult_87_SUMB_21__40_), .CO(
        u5_mult_87_CARRYB_22__39_), .S(u5_mult_87_SUMB_22__39_) );
  FA_X1 u5_mult_87_S2_22_38 ( .A(u5_mult_87_ab_22__38_), .B(
        u5_mult_87_CARRYB_21__38_), .CI(u5_mult_87_SUMB_21__39_), .CO(
        u5_mult_87_CARRYB_22__38_), .S(u5_mult_87_SUMB_22__38_) );
  FA_X1 u5_mult_87_S2_22_37 ( .A(u5_mult_87_ab_22__37_), .B(
        u5_mult_87_CARRYB_21__37_), .CI(u5_mult_87_SUMB_21__38_), .CO(
        u5_mult_87_CARRYB_22__37_), .S(u5_mult_87_SUMB_22__37_) );
  FA_X1 u5_mult_87_S2_22_36 ( .A(u5_mult_87_ab_22__36_), .B(
        u5_mult_87_CARRYB_21__36_), .CI(u5_mult_87_SUMB_21__37_), .CO(
        u5_mult_87_CARRYB_22__36_), .S(u5_mult_87_SUMB_22__36_) );
  FA_X1 u5_mult_87_S2_22_35 ( .A(u5_mult_87_ab_22__35_), .B(
        u5_mult_87_CARRYB_21__35_), .CI(u5_mult_87_SUMB_21__36_), .CO(
        u5_mult_87_CARRYB_22__35_), .S(u5_mult_87_SUMB_22__35_) );
  FA_X1 u5_mult_87_S2_22_34 ( .A(u5_mult_87_ab_22__34_), .B(
        u5_mult_87_CARRYB_21__34_), .CI(u5_mult_87_SUMB_21__35_), .CO(
        u5_mult_87_CARRYB_22__34_), .S(u5_mult_87_SUMB_22__34_) );
  FA_X1 u5_mult_87_S2_22_33 ( .A(u5_mult_87_ab_22__33_), .B(
        u5_mult_87_CARRYB_21__33_), .CI(u5_mult_87_SUMB_21__34_), .CO(
        u5_mult_87_CARRYB_22__33_), .S(u5_mult_87_SUMB_22__33_) );
  FA_X1 u5_mult_87_S2_22_32 ( .A(u5_mult_87_ab_22__32_), .B(
        u5_mult_87_CARRYB_21__32_), .CI(u5_mult_87_SUMB_21__33_), .CO(
        u5_mult_87_CARRYB_22__32_), .S(u5_mult_87_SUMB_22__32_) );
  FA_X1 u5_mult_87_S2_22_31 ( .A(u5_mult_87_ab_22__31_), .B(
        u5_mult_87_CARRYB_21__31_), .CI(u5_mult_87_SUMB_21__32_), .CO(
        u5_mult_87_CARRYB_22__31_), .S(u5_mult_87_SUMB_22__31_) );
  FA_X1 u5_mult_87_S2_22_30 ( .A(u5_mult_87_ab_22__30_), .B(
        u5_mult_87_CARRYB_21__30_), .CI(u5_mult_87_SUMB_21__31_), .CO(
        u5_mult_87_CARRYB_22__30_), .S(u5_mult_87_SUMB_22__30_) );
  FA_X1 u5_mult_87_S2_22_29 ( .A(u5_mult_87_ab_22__29_), .B(
        u5_mult_87_CARRYB_21__29_), .CI(u5_mult_87_SUMB_21__30_), .CO(
        u5_mult_87_CARRYB_22__29_), .S(u5_mult_87_SUMB_22__29_) );
  FA_X1 u5_mult_87_S2_22_28 ( .A(u5_mult_87_ab_22__28_), .B(
        u5_mult_87_CARRYB_21__28_), .CI(u5_mult_87_SUMB_21__29_), .CO(
        u5_mult_87_CARRYB_22__28_), .S(u5_mult_87_SUMB_22__28_) );
  FA_X1 u5_mult_87_S2_22_27 ( .A(u5_mult_87_ab_22__27_), .B(
        u5_mult_87_CARRYB_21__27_), .CI(u5_mult_87_SUMB_21__28_), .CO(
        u5_mult_87_CARRYB_22__27_), .S(u5_mult_87_SUMB_22__27_) );
  FA_X1 u5_mult_87_S2_22_26 ( .A(u5_mult_87_ab_22__26_), .B(
        u5_mult_87_CARRYB_21__26_), .CI(u5_mult_87_SUMB_21__27_), .CO(
        u5_mult_87_CARRYB_22__26_), .S(u5_mult_87_SUMB_22__26_) );
  FA_X1 u5_mult_87_S2_22_25 ( .A(u5_mult_87_ab_22__25_), .B(
        u5_mult_87_CARRYB_21__25_), .CI(u5_mult_87_SUMB_21__26_), .CO(
        u5_mult_87_CARRYB_22__25_), .S(u5_mult_87_SUMB_22__25_) );
  FA_X1 u5_mult_87_S2_22_24 ( .A(u5_mult_87_ab_22__24_), .B(
        u5_mult_87_CARRYB_21__24_), .CI(u5_mult_87_SUMB_21__25_), .CO(
        u5_mult_87_CARRYB_22__24_), .S(u5_mult_87_SUMB_22__24_) );
  FA_X1 u5_mult_87_S2_22_23 ( .A(u5_mult_87_ab_22__23_), .B(
        u5_mult_87_CARRYB_21__23_), .CI(u5_mult_87_SUMB_21__24_), .CO(
        u5_mult_87_CARRYB_22__23_), .S(u5_mult_87_SUMB_22__23_) );
  FA_X1 u5_mult_87_S2_22_22 ( .A(u5_mult_87_ab_22__22_), .B(
        u5_mult_87_CARRYB_21__22_), .CI(u5_mult_87_SUMB_21__23_), .CO(
        u5_mult_87_CARRYB_22__22_), .S(u5_mult_87_SUMB_22__22_) );
  FA_X1 u5_mult_87_S2_22_21 ( .A(u5_mult_87_ab_22__21_), .B(
        u5_mult_87_CARRYB_21__21_), .CI(u5_mult_87_SUMB_21__22_), .CO(
        u5_mult_87_CARRYB_22__21_), .S(u5_mult_87_SUMB_22__21_) );
  FA_X1 u5_mult_87_S2_22_20 ( .A(u5_mult_87_ab_22__20_), .B(
        u5_mult_87_CARRYB_21__20_), .CI(u5_mult_87_SUMB_21__21_), .CO(
        u5_mult_87_CARRYB_22__20_), .S(u5_mult_87_SUMB_22__20_) );
  FA_X1 u5_mult_87_S2_22_19 ( .A(u5_mult_87_ab_22__19_), .B(
        u5_mult_87_CARRYB_21__19_), .CI(u5_mult_87_SUMB_21__20_), .CO(
        u5_mult_87_CARRYB_22__19_), .S(u5_mult_87_SUMB_22__19_) );
  FA_X1 u5_mult_87_S2_22_18 ( .A(u5_mult_87_ab_22__18_), .B(
        u5_mult_87_CARRYB_21__18_), .CI(u5_mult_87_SUMB_21__19_), .CO(
        u5_mult_87_CARRYB_22__18_), .S(u5_mult_87_SUMB_22__18_) );
  FA_X1 u5_mult_87_S2_22_17 ( .A(u5_mult_87_ab_22__17_), .B(
        u5_mult_87_CARRYB_21__17_), .CI(u5_mult_87_SUMB_21__18_), .CO(
        u5_mult_87_CARRYB_22__17_), .S(u5_mult_87_SUMB_22__17_) );
  FA_X1 u5_mult_87_S2_22_16 ( .A(u5_mult_87_ab_22__16_), .B(
        u5_mult_87_CARRYB_21__16_), .CI(u5_mult_87_SUMB_21__17_), .CO(
        u5_mult_87_CARRYB_22__16_), .S(u5_mult_87_SUMB_22__16_) );
  FA_X1 u5_mult_87_S2_22_15 ( .A(u5_mult_87_ab_22__15_), .B(
        u5_mult_87_CARRYB_21__15_), .CI(u5_mult_87_SUMB_21__16_), .CO(
        u5_mult_87_CARRYB_22__15_), .S(u5_mult_87_SUMB_22__15_) );
  FA_X1 u5_mult_87_S2_22_14 ( .A(u5_mult_87_ab_22__14_), .B(
        u5_mult_87_CARRYB_21__14_), .CI(u5_mult_87_SUMB_21__15_), .CO(
        u5_mult_87_CARRYB_22__14_), .S(u5_mult_87_SUMB_22__14_) );
  FA_X1 u5_mult_87_S2_22_13 ( .A(u5_mult_87_ab_22__13_), .B(
        u5_mult_87_CARRYB_21__13_), .CI(u5_mult_87_SUMB_21__14_), .CO(
        u5_mult_87_CARRYB_22__13_), .S(u5_mult_87_SUMB_22__13_) );
  FA_X1 u5_mult_87_S2_22_12 ( .A(u5_mult_87_ab_22__12_), .B(
        u5_mult_87_CARRYB_21__12_), .CI(u5_mult_87_SUMB_21__13_), .CO(
        u5_mult_87_CARRYB_22__12_), .S(u5_mult_87_SUMB_22__12_) );
  FA_X1 u5_mult_87_S2_22_11 ( .A(u5_mult_87_ab_22__11_), .B(
        u5_mult_87_CARRYB_21__11_), .CI(u5_mult_87_SUMB_21__12_), .CO(
        u5_mult_87_CARRYB_22__11_), .S(u5_mult_87_SUMB_22__11_) );
  FA_X1 u5_mult_87_S2_22_10 ( .A(u5_mult_87_ab_22__10_), .B(
        u5_mult_87_CARRYB_21__10_), .CI(u5_mult_87_SUMB_21__11_), .CO(
        u5_mult_87_CARRYB_22__10_), .S(u5_mult_87_SUMB_22__10_) );
  FA_X1 u5_mult_87_S2_22_9 ( .A(u5_mult_87_ab_22__9_), .B(
        u5_mult_87_CARRYB_21__9_), .CI(u5_mult_87_SUMB_21__10_), .CO(
        u5_mult_87_CARRYB_22__9_), .S(u5_mult_87_SUMB_22__9_) );
  FA_X1 u5_mult_87_S2_22_8 ( .A(u5_mult_87_ab_22__8_), .B(
        u5_mult_87_CARRYB_21__8_), .CI(u5_mult_87_SUMB_21__9_), .CO(
        u5_mult_87_CARRYB_22__8_), .S(u5_mult_87_SUMB_22__8_) );
  FA_X1 u5_mult_87_S2_22_7 ( .A(u5_mult_87_ab_22__7_), .B(
        u5_mult_87_CARRYB_21__7_), .CI(u5_mult_87_SUMB_21__8_), .CO(
        u5_mult_87_CARRYB_22__7_), .S(u5_mult_87_SUMB_22__7_) );
  FA_X1 u5_mult_87_S2_22_6 ( .A(u5_mult_87_ab_22__6_), .B(
        u5_mult_87_CARRYB_21__6_), .CI(u5_mult_87_SUMB_21__7_), .CO(
        u5_mult_87_CARRYB_22__6_), .S(u5_mult_87_SUMB_22__6_) );
  FA_X1 u5_mult_87_S2_22_5 ( .A(u5_mult_87_ab_22__5_), .B(
        u5_mult_87_CARRYB_21__5_), .CI(u5_mult_87_SUMB_21__6_), .CO(
        u5_mult_87_CARRYB_22__5_), .S(u5_mult_87_SUMB_22__5_) );
  FA_X1 u5_mult_87_S2_22_4 ( .A(u5_mult_87_ab_22__4_), .B(
        u5_mult_87_CARRYB_21__4_), .CI(u5_mult_87_SUMB_21__5_), .CO(
        u5_mult_87_CARRYB_22__4_), .S(u5_mult_87_SUMB_22__4_) );
  FA_X1 u5_mult_87_S2_22_3 ( .A(u5_mult_87_ab_22__3_), .B(
        u5_mult_87_CARRYB_21__3_), .CI(u5_mult_87_SUMB_21__4_), .CO(
        u5_mult_87_CARRYB_22__3_), .S(u5_mult_87_SUMB_22__3_) );
  FA_X1 u5_mult_87_S2_22_2 ( .A(u5_mult_87_ab_22__2_), .B(
        u5_mult_87_CARRYB_21__2_), .CI(u5_mult_87_SUMB_21__3_), .CO(
        u5_mult_87_CARRYB_22__2_), .S(u5_mult_87_SUMB_22__2_) );
  FA_X1 u5_mult_87_S2_22_1 ( .A(u5_mult_87_ab_22__1_), .B(
        u5_mult_87_CARRYB_21__1_), .CI(u5_mult_87_SUMB_21__2_), .CO(
        u5_mult_87_CARRYB_22__1_), .S(u5_mult_87_SUMB_22__1_) );
  FA_X1 u5_mult_87_S1_22_0 ( .A(u5_mult_87_ab_22__0_), .B(
        u5_mult_87_CARRYB_21__0_), .CI(u5_mult_87_SUMB_21__1_), .CO(
        u5_mult_87_CARRYB_22__0_), .S(u5_N22) );
  FA_X1 u5_mult_87_S3_23_51 ( .A(u5_mult_87_ab_23__51_), .B(
        u5_mult_87_CARRYB_22__51_), .CI(u5_mult_87_ab_22__52_), .CO(
        u5_mult_87_CARRYB_23__51_), .S(u5_mult_87_SUMB_23__51_) );
  FA_X1 u5_mult_87_S2_23_50 ( .A(u5_mult_87_ab_23__50_), .B(
        u5_mult_87_CARRYB_22__50_), .CI(u5_mult_87_SUMB_22__51_), .CO(
        u5_mult_87_CARRYB_23__50_), .S(u5_mult_87_SUMB_23__50_) );
  FA_X1 u5_mult_87_S2_23_49 ( .A(u5_mult_87_ab_23__49_), .B(
        u5_mult_87_CARRYB_22__49_), .CI(u5_mult_87_SUMB_22__50_), .CO(
        u5_mult_87_CARRYB_23__49_), .S(u5_mult_87_SUMB_23__49_) );
  FA_X1 u5_mult_87_S2_23_48 ( .A(u5_mult_87_ab_23__48_), .B(
        u5_mult_87_CARRYB_22__48_), .CI(u5_mult_87_SUMB_22__49_), .CO(
        u5_mult_87_CARRYB_23__48_), .S(u5_mult_87_SUMB_23__48_) );
  FA_X1 u5_mult_87_S2_23_47 ( .A(u5_mult_87_ab_23__47_), .B(
        u5_mult_87_CARRYB_22__47_), .CI(u5_mult_87_SUMB_22__48_), .CO(
        u5_mult_87_CARRYB_23__47_), .S(u5_mult_87_SUMB_23__47_) );
  FA_X1 u5_mult_87_S2_23_46 ( .A(u5_mult_87_ab_23__46_), .B(
        u5_mult_87_CARRYB_22__46_), .CI(u5_mult_87_SUMB_22__47_), .CO(
        u5_mult_87_CARRYB_23__46_), .S(u5_mult_87_SUMB_23__46_) );
  FA_X1 u5_mult_87_S2_23_45 ( .A(u5_mult_87_ab_23__45_), .B(
        u5_mult_87_CARRYB_22__45_), .CI(u5_mult_87_SUMB_22__46_), .CO(
        u5_mult_87_CARRYB_23__45_), .S(u5_mult_87_SUMB_23__45_) );
  FA_X1 u5_mult_87_S2_23_44 ( .A(u5_mult_87_ab_23__44_), .B(
        u5_mult_87_CARRYB_22__44_), .CI(u5_mult_87_SUMB_22__45_), .CO(
        u5_mult_87_CARRYB_23__44_), .S(u5_mult_87_SUMB_23__44_) );
  FA_X1 u5_mult_87_S2_23_43 ( .A(u5_mult_87_ab_23__43_), .B(
        u5_mult_87_CARRYB_22__43_), .CI(u5_mult_87_SUMB_22__44_), .CO(
        u5_mult_87_CARRYB_23__43_), .S(u5_mult_87_SUMB_23__43_) );
  FA_X1 u5_mult_87_S2_23_42 ( .A(u5_mult_87_ab_23__42_), .B(
        u5_mult_87_CARRYB_22__42_), .CI(u5_mult_87_SUMB_22__43_), .CO(
        u5_mult_87_CARRYB_23__42_), .S(u5_mult_87_SUMB_23__42_) );
  FA_X1 u5_mult_87_S2_23_41 ( .A(u5_mult_87_ab_23__41_), .B(
        u5_mult_87_CARRYB_22__41_), .CI(u5_mult_87_SUMB_22__42_), .CO(
        u5_mult_87_CARRYB_23__41_), .S(u5_mult_87_SUMB_23__41_) );
  FA_X1 u5_mult_87_S2_23_40 ( .A(u5_mult_87_ab_23__40_), .B(
        u5_mult_87_CARRYB_22__40_), .CI(u5_mult_87_SUMB_22__41_), .CO(
        u5_mult_87_CARRYB_23__40_), .S(u5_mult_87_SUMB_23__40_) );
  FA_X1 u5_mult_87_S2_23_39 ( .A(u5_mult_87_ab_23__39_), .B(
        u5_mult_87_CARRYB_22__39_), .CI(u5_mult_87_SUMB_22__40_), .CO(
        u5_mult_87_CARRYB_23__39_), .S(u5_mult_87_SUMB_23__39_) );
  FA_X1 u5_mult_87_S2_23_38 ( .A(u5_mult_87_ab_23__38_), .B(
        u5_mult_87_CARRYB_22__38_), .CI(u5_mult_87_SUMB_22__39_), .CO(
        u5_mult_87_CARRYB_23__38_), .S(u5_mult_87_SUMB_23__38_) );
  FA_X1 u5_mult_87_S2_23_37 ( .A(u5_mult_87_ab_23__37_), .B(
        u5_mult_87_CARRYB_22__37_), .CI(u5_mult_87_SUMB_22__38_), .CO(
        u5_mult_87_CARRYB_23__37_), .S(u5_mult_87_SUMB_23__37_) );
  FA_X1 u5_mult_87_S2_23_36 ( .A(u5_mult_87_ab_23__36_), .B(
        u5_mult_87_CARRYB_22__36_), .CI(u5_mult_87_SUMB_22__37_), .CO(
        u5_mult_87_CARRYB_23__36_), .S(u5_mult_87_SUMB_23__36_) );
  FA_X1 u5_mult_87_S2_23_35 ( .A(u5_mult_87_ab_23__35_), .B(
        u5_mult_87_CARRYB_22__35_), .CI(u5_mult_87_SUMB_22__36_), .CO(
        u5_mult_87_CARRYB_23__35_), .S(u5_mult_87_SUMB_23__35_) );
  FA_X1 u5_mult_87_S2_23_34 ( .A(u5_mult_87_ab_23__34_), .B(
        u5_mult_87_CARRYB_22__34_), .CI(u5_mult_87_SUMB_22__35_), .CO(
        u5_mult_87_CARRYB_23__34_), .S(u5_mult_87_SUMB_23__34_) );
  FA_X1 u5_mult_87_S2_23_33 ( .A(u5_mult_87_ab_23__33_), .B(
        u5_mult_87_CARRYB_22__33_), .CI(u5_mult_87_SUMB_22__34_), .CO(
        u5_mult_87_CARRYB_23__33_), .S(u5_mult_87_SUMB_23__33_) );
  FA_X1 u5_mult_87_S2_23_32 ( .A(u5_mult_87_ab_23__32_), .B(
        u5_mult_87_CARRYB_22__32_), .CI(u5_mult_87_SUMB_22__33_), .CO(
        u5_mult_87_CARRYB_23__32_), .S(u5_mult_87_SUMB_23__32_) );
  FA_X1 u5_mult_87_S2_23_31 ( .A(u5_mult_87_ab_23__31_), .B(
        u5_mult_87_CARRYB_22__31_), .CI(u5_mult_87_SUMB_22__32_), .CO(
        u5_mult_87_CARRYB_23__31_), .S(u5_mult_87_SUMB_23__31_) );
  FA_X1 u5_mult_87_S2_23_30 ( .A(u5_mult_87_ab_23__30_), .B(
        u5_mult_87_CARRYB_22__30_), .CI(u5_mult_87_SUMB_22__31_), .CO(
        u5_mult_87_CARRYB_23__30_), .S(u5_mult_87_SUMB_23__30_) );
  FA_X1 u5_mult_87_S2_23_29 ( .A(u5_mult_87_ab_23__29_), .B(
        u5_mult_87_CARRYB_22__29_), .CI(u5_mult_87_SUMB_22__30_), .CO(
        u5_mult_87_CARRYB_23__29_), .S(u5_mult_87_SUMB_23__29_) );
  FA_X1 u5_mult_87_S2_23_28 ( .A(u5_mult_87_ab_23__28_), .B(
        u5_mult_87_CARRYB_22__28_), .CI(u5_mult_87_SUMB_22__29_), .CO(
        u5_mult_87_CARRYB_23__28_), .S(u5_mult_87_SUMB_23__28_) );
  FA_X1 u5_mult_87_S2_23_27 ( .A(u5_mult_87_ab_23__27_), .B(
        u5_mult_87_CARRYB_22__27_), .CI(u5_mult_87_SUMB_22__28_), .CO(
        u5_mult_87_CARRYB_23__27_), .S(u5_mult_87_SUMB_23__27_) );
  FA_X1 u5_mult_87_S2_23_26 ( .A(u5_mult_87_ab_23__26_), .B(
        u5_mult_87_CARRYB_22__26_), .CI(u5_mult_87_SUMB_22__27_), .CO(
        u5_mult_87_CARRYB_23__26_), .S(u5_mult_87_SUMB_23__26_) );
  FA_X1 u5_mult_87_S2_23_25 ( .A(u5_mult_87_ab_23__25_), .B(
        u5_mult_87_CARRYB_22__25_), .CI(u5_mult_87_SUMB_22__26_), .CO(
        u5_mult_87_CARRYB_23__25_), .S(u5_mult_87_SUMB_23__25_) );
  FA_X1 u5_mult_87_S2_23_24 ( .A(u5_mult_87_ab_23__24_), .B(
        u5_mult_87_CARRYB_22__24_), .CI(u5_mult_87_SUMB_22__25_), .CO(
        u5_mult_87_CARRYB_23__24_), .S(u5_mult_87_SUMB_23__24_) );
  FA_X1 u5_mult_87_S2_23_23 ( .A(u5_mult_87_ab_23__23_), .B(
        u5_mult_87_CARRYB_22__23_), .CI(u5_mult_87_SUMB_22__24_), .CO(
        u5_mult_87_CARRYB_23__23_), .S(u5_mult_87_SUMB_23__23_) );
  FA_X1 u5_mult_87_S2_23_22 ( .A(u5_mult_87_ab_23__22_), .B(
        u5_mult_87_CARRYB_22__22_), .CI(u5_mult_87_SUMB_22__23_), .CO(
        u5_mult_87_CARRYB_23__22_), .S(u5_mult_87_SUMB_23__22_) );
  FA_X1 u5_mult_87_S2_23_21 ( .A(u5_mult_87_ab_23__21_), .B(
        u5_mult_87_CARRYB_22__21_), .CI(u5_mult_87_SUMB_22__22_), .CO(
        u5_mult_87_CARRYB_23__21_), .S(u5_mult_87_SUMB_23__21_) );
  FA_X1 u5_mult_87_S2_23_20 ( .A(u5_mult_87_ab_23__20_), .B(
        u5_mult_87_CARRYB_22__20_), .CI(u5_mult_87_SUMB_22__21_), .CO(
        u5_mult_87_CARRYB_23__20_), .S(u5_mult_87_SUMB_23__20_) );
  FA_X1 u5_mult_87_S2_23_19 ( .A(u5_mult_87_ab_23__19_), .B(
        u5_mult_87_CARRYB_22__19_), .CI(u5_mult_87_SUMB_22__20_), .CO(
        u5_mult_87_CARRYB_23__19_), .S(u5_mult_87_SUMB_23__19_) );
  FA_X1 u5_mult_87_S2_23_18 ( .A(u5_mult_87_ab_23__18_), .B(
        u5_mult_87_CARRYB_22__18_), .CI(u5_mult_87_SUMB_22__19_), .CO(
        u5_mult_87_CARRYB_23__18_), .S(u5_mult_87_SUMB_23__18_) );
  FA_X1 u5_mult_87_S2_23_17 ( .A(u5_mult_87_ab_23__17_), .B(
        u5_mult_87_CARRYB_22__17_), .CI(u5_mult_87_SUMB_22__18_), .CO(
        u5_mult_87_CARRYB_23__17_), .S(u5_mult_87_SUMB_23__17_) );
  FA_X1 u5_mult_87_S2_23_16 ( .A(u5_mult_87_ab_23__16_), .B(
        u5_mult_87_CARRYB_22__16_), .CI(u5_mult_87_SUMB_22__17_), .CO(
        u5_mult_87_CARRYB_23__16_), .S(u5_mult_87_SUMB_23__16_) );
  FA_X1 u5_mult_87_S2_23_15 ( .A(u5_mult_87_ab_23__15_), .B(
        u5_mult_87_CARRYB_22__15_), .CI(u5_mult_87_SUMB_22__16_), .CO(
        u5_mult_87_CARRYB_23__15_), .S(u5_mult_87_SUMB_23__15_) );
  FA_X1 u5_mult_87_S2_23_14 ( .A(u5_mult_87_ab_23__14_), .B(
        u5_mult_87_CARRYB_22__14_), .CI(u5_mult_87_SUMB_22__15_), .CO(
        u5_mult_87_CARRYB_23__14_), .S(u5_mult_87_SUMB_23__14_) );
  FA_X1 u5_mult_87_S2_23_13 ( .A(u5_mult_87_ab_23__13_), .B(
        u5_mult_87_CARRYB_22__13_), .CI(u5_mult_87_SUMB_22__14_), .CO(
        u5_mult_87_CARRYB_23__13_), .S(u5_mult_87_SUMB_23__13_) );
  FA_X1 u5_mult_87_S2_23_12 ( .A(u5_mult_87_ab_23__12_), .B(
        u5_mult_87_CARRYB_22__12_), .CI(u5_mult_87_SUMB_22__13_), .CO(
        u5_mult_87_CARRYB_23__12_), .S(u5_mult_87_SUMB_23__12_) );
  FA_X1 u5_mult_87_S2_23_11 ( .A(u5_mult_87_ab_23__11_), .B(
        u5_mult_87_CARRYB_22__11_), .CI(u5_mult_87_SUMB_22__12_), .CO(
        u5_mult_87_CARRYB_23__11_), .S(u5_mult_87_SUMB_23__11_) );
  FA_X1 u5_mult_87_S2_23_10 ( .A(u5_mult_87_ab_23__10_), .B(
        u5_mult_87_CARRYB_22__10_), .CI(u5_mult_87_SUMB_22__11_), .CO(
        u5_mult_87_CARRYB_23__10_), .S(u5_mult_87_SUMB_23__10_) );
  FA_X1 u5_mult_87_S2_23_9 ( .A(u5_mult_87_ab_23__9_), .B(
        u5_mult_87_CARRYB_22__9_), .CI(u5_mult_87_SUMB_22__10_), .CO(
        u5_mult_87_CARRYB_23__9_), .S(u5_mult_87_SUMB_23__9_) );
  FA_X1 u5_mult_87_S2_23_8 ( .A(u5_mult_87_ab_23__8_), .B(
        u5_mult_87_CARRYB_22__8_), .CI(u5_mult_87_SUMB_22__9_), .CO(
        u5_mult_87_CARRYB_23__8_), .S(u5_mult_87_SUMB_23__8_) );
  FA_X1 u5_mult_87_S2_23_7 ( .A(u5_mult_87_ab_23__7_), .B(
        u5_mult_87_CARRYB_22__7_), .CI(u5_mult_87_SUMB_22__8_), .CO(
        u5_mult_87_CARRYB_23__7_), .S(u5_mult_87_SUMB_23__7_) );
  FA_X1 u5_mult_87_S2_23_6 ( .A(u5_mult_87_ab_23__6_), .B(
        u5_mult_87_CARRYB_22__6_), .CI(u5_mult_87_SUMB_22__7_), .CO(
        u5_mult_87_CARRYB_23__6_), .S(u5_mult_87_SUMB_23__6_) );
  FA_X1 u5_mult_87_S2_23_5 ( .A(u5_mult_87_ab_23__5_), .B(
        u5_mult_87_CARRYB_22__5_), .CI(u5_mult_87_SUMB_22__6_), .CO(
        u5_mult_87_CARRYB_23__5_), .S(u5_mult_87_SUMB_23__5_) );
  FA_X1 u5_mult_87_S2_23_4 ( .A(u5_mult_87_ab_23__4_), .B(
        u5_mult_87_CARRYB_22__4_), .CI(u5_mult_87_SUMB_22__5_), .CO(
        u5_mult_87_CARRYB_23__4_), .S(u5_mult_87_SUMB_23__4_) );
  FA_X1 u5_mult_87_S2_23_3 ( .A(u5_mult_87_ab_23__3_), .B(
        u5_mult_87_CARRYB_22__3_), .CI(u5_mult_87_SUMB_22__4_), .CO(
        u5_mult_87_CARRYB_23__3_), .S(u5_mult_87_SUMB_23__3_) );
  FA_X1 u5_mult_87_S2_23_2 ( .A(u5_mult_87_ab_23__2_), .B(
        u5_mult_87_CARRYB_22__2_), .CI(u5_mult_87_SUMB_22__3_), .CO(
        u5_mult_87_CARRYB_23__2_), .S(u5_mult_87_SUMB_23__2_) );
  FA_X1 u5_mult_87_S2_23_1 ( .A(u5_mult_87_ab_23__1_), .B(
        u5_mult_87_CARRYB_22__1_), .CI(u5_mult_87_SUMB_22__2_), .CO(
        u5_mult_87_CARRYB_23__1_), .S(u5_mult_87_SUMB_23__1_) );
  FA_X1 u5_mult_87_S1_23_0 ( .A(u5_mult_87_ab_23__0_), .B(
        u5_mult_87_CARRYB_22__0_), .CI(u5_mult_87_SUMB_22__1_), .CO(
        u5_mult_87_CARRYB_23__0_), .S(u5_N23) );
  FA_X1 u5_mult_87_S3_24_51 ( .A(u5_mult_87_ab_24__51_), .B(
        u5_mult_87_CARRYB_23__51_), .CI(u5_mult_87_ab_23__52_), .CO(
        u5_mult_87_CARRYB_24__51_), .S(u5_mult_87_SUMB_24__51_) );
  FA_X1 u5_mult_87_S2_24_50 ( .A(u5_mult_87_ab_24__50_), .B(
        u5_mult_87_CARRYB_23__50_), .CI(u5_mult_87_SUMB_23__51_), .CO(
        u5_mult_87_CARRYB_24__50_), .S(u5_mult_87_SUMB_24__50_) );
  FA_X1 u5_mult_87_S2_24_49 ( .A(u5_mult_87_ab_24__49_), .B(
        u5_mult_87_CARRYB_23__49_), .CI(u5_mult_87_SUMB_23__50_), .CO(
        u5_mult_87_CARRYB_24__49_), .S(u5_mult_87_SUMB_24__49_) );
  FA_X1 u5_mult_87_S2_24_48 ( .A(u5_mult_87_ab_24__48_), .B(
        u5_mult_87_CARRYB_23__48_), .CI(u5_mult_87_SUMB_23__49_), .CO(
        u5_mult_87_CARRYB_24__48_), .S(u5_mult_87_SUMB_24__48_) );
  FA_X1 u5_mult_87_S2_24_47 ( .A(u5_mult_87_ab_24__47_), .B(
        u5_mult_87_CARRYB_23__47_), .CI(u5_mult_87_SUMB_23__48_), .CO(
        u5_mult_87_CARRYB_24__47_), .S(u5_mult_87_SUMB_24__47_) );
  FA_X1 u5_mult_87_S2_24_46 ( .A(u5_mult_87_ab_24__46_), .B(
        u5_mult_87_CARRYB_23__46_), .CI(u5_mult_87_SUMB_23__47_), .CO(
        u5_mult_87_CARRYB_24__46_), .S(u5_mult_87_SUMB_24__46_) );
  FA_X1 u5_mult_87_S2_24_45 ( .A(u5_mult_87_ab_24__45_), .B(
        u5_mult_87_CARRYB_23__45_), .CI(u5_mult_87_SUMB_23__46_), .CO(
        u5_mult_87_CARRYB_24__45_), .S(u5_mult_87_SUMB_24__45_) );
  FA_X1 u5_mult_87_S2_24_44 ( .A(u5_mult_87_ab_24__44_), .B(
        u5_mult_87_CARRYB_23__44_), .CI(u5_mult_87_SUMB_23__45_), .CO(
        u5_mult_87_CARRYB_24__44_), .S(u5_mult_87_SUMB_24__44_) );
  FA_X1 u5_mult_87_S2_24_43 ( .A(u5_mult_87_ab_24__43_), .B(
        u5_mult_87_CARRYB_23__43_), .CI(u5_mult_87_SUMB_23__44_), .CO(
        u5_mult_87_CARRYB_24__43_), .S(u5_mult_87_SUMB_24__43_) );
  FA_X1 u5_mult_87_S2_24_42 ( .A(u5_mult_87_ab_24__42_), .B(
        u5_mult_87_CARRYB_23__42_), .CI(u5_mult_87_SUMB_23__43_), .CO(
        u5_mult_87_CARRYB_24__42_), .S(u5_mult_87_SUMB_24__42_) );
  FA_X1 u5_mult_87_S2_24_41 ( .A(u5_mult_87_ab_24__41_), .B(
        u5_mult_87_CARRYB_23__41_), .CI(u5_mult_87_SUMB_23__42_), .CO(
        u5_mult_87_CARRYB_24__41_), .S(u5_mult_87_SUMB_24__41_) );
  FA_X1 u5_mult_87_S2_24_40 ( .A(u5_mult_87_ab_24__40_), .B(
        u5_mult_87_CARRYB_23__40_), .CI(u5_mult_87_SUMB_23__41_), .CO(
        u5_mult_87_CARRYB_24__40_), .S(u5_mult_87_SUMB_24__40_) );
  FA_X1 u5_mult_87_S2_24_39 ( .A(u5_mult_87_ab_24__39_), .B(
        u5_mult_87_CARRYB_23__39_), .CI(u5_mult_87_SUMB_23__40_), .CO(
        u5_mult_87_CARRYB_24__39_), .S(u5_mult_87_SUMB_24__39_) );
  FA_X1 u5_mult_87_S2_24_38 ( .A(u5_mult_87_ab_24__38_), .B(
        u5_mult_87_CARRYB_23__38_), .CI(u5_mult_87_SUMB_23__39_), .CO(
        u5_mult_87_CARRYB_24__38_), .S(u5_mult_87_SUMB_24__38_) );
  FA_X1 u5_mult_87_S2_24_37 ( .A(u5_mult_87_ab_24__37_), .B(
        u5_mult_87_CARRYB_23__37_), .CI(u5_mult_87_SUMB_23__38_), .CO(
        u5_mult_87_CARRYB_24__37_), .S(u5_mult_87_SUMB_24__37_) );
  FA_X1 u5_mult_87_S2_24_36 ( .A(u5_mult_87_ab_24__36_), .B(
        u5_mult_87_CARRYB_23__36_), .CI(u5_mult_87_SUMB_23__37_), .CO(
        u5_mult_87_CARRYB_24__36_), .S(u5_mult_87_SUMB_24__36_) );
  FA_X1 u5_mult_87_S2_24_35 ( .A(u5_mult_87_ab_24__35_), .B(
        u5_mult_87_CARRYB_23__35_), .CI(u5_mult_87_SUMB_23__36_), .CO(
        u5_mult_87_CARRYB_24__35_), .S(u5_mult_87_SUMB_24__35_) );
  FA_X1 u5_mult_87_S2_24_34 ( .A(u5_mult_87_ab_24__34_), .B(
        u5_mult_87_CARRYB_23__34_), .CI(u5_mult_87_SUMB_23__35_), .CO(
        u5_mult_87_CARRYB_24__34_), .S(u5_mult_87_SUMB_24__34_) );
  FA_X1 u5_mult_87_S2_24_33 ( .A(u5_mult_87_ab_24__33_), .B(
        u5_mult_87_CARRYB_23__33_), .CI(u5_mult_87_SUMB_23__34_), .CO(
        u5_mult_87_CARRYB_24__33_), .S(u5_mult_87_SUMB_24__33_) );
  FA_X1 u5_mult_87_S2_24_32 ( .A(u5_mult_87_ab_24__32_), .B(
        u5_mult_87_CARRYB_23__32_), .CI(u5_mult_87_SUMB_23__33_), .CO(
        u5_mult_87_CARRYB_24__32_), .S(u5_mult_87_SUMB_24__32_) );
  FA_X1 u5_mult_87_S2_24_31 ( .A(u5_mult_87_ab_24__31_), .B(
        u5_mult_87_CARRYB_23__31_), .CI(u5_mult_87_SUMB_23__32_), .CO(
        u5_mult_87_CARRYB_24__31_), .S(u5_mult_87_SUMB_24__31_) );
  FA_X1 u5_mult_87_S2_24_30 ( .A(u5_mult_87_ab_24__30_), .B(
        u5_mult_87_CARRYB_23__30_), .CI(u5_mult_87_SUMB_23__31_), .CO(
        u5_mult_87_CARRYB_24__30_), .S(u5_mult_87_SUMB_24__30_) );
  FA_X1 u5_mult_87_S2_24_29 ( .A(u5_mult_87_ab_24__29_), .B(
        u5_mult_87_CARRYB_23__29_), .CI(u5_mult_87_SUMB_23__30_), .CO(
        u5_mult_87_CARRYB_24__29_), .S(u5_mult_87_SUMB_24__29_) );
  FA_X1 u5_mult_87_S2_24_28 ( .A(u5_mult_87_ab_24__28_), .B(
        u5_mult_87_CARRYB_23__28_), .CI(u5_mult_87_SUMB_23__29_), .CO(
        u5_mult_87_CARRYB_24__28_), .S(u5_mult_87_SUMB_24__28_) );
  FA_X1 u5_mult_87_S2_24_27 ( .A(u5_mult_87_ab_24__27_), .B(
        u5_mult_87_CARRYB_23__27_), .CI(u5_mult_87_SUMB_23__28_), .CO(
        u5_mult_87_CARRYB_24__27_), .S(u5_mult_87_SUMB_24__27_) );
  FA_X1 u5_mult_87_S2_24_26 ( .A(u5_mult_87_ab_24__26_), .B(
        u5_mult_87_CARRYB_23__26_), .CI(u5_mult_87_SUMB_23__27_), .CO(
        u5_mult_87_CARRYB_24__26_), .S(u5_mult_87_SUMB_24__26_) );
  FA_X1 u5_mult_87_S2_24_25 ( .A(u5_mult_87_ab_24__25_), .B(
        u5_mult_87_CARRYB_23__25_), .CI(u5_mult_87_SUMB_23__26_), .CO(
        u5_mult_87_CARRYB_24__25_), .S(u5_mult_87_SUMB_24__25_) );
  FA_X1 u5_mult_87_S2_24_24 ( .A(u5_mult_87_ab_24__24_), .B(
        u5_mult_87_CARRYB_23__24_), .CI(u5_mult_87_SUMB_23__25_), .CO(
        u5_mult_87_CARRYB_24__24_), .S(u5_mult_87_SUMB_24__24_) );
  FA_X1 u5_mult_87_S2_24_23 ( .A(u5_mult_87_ab_24__23_), .B(
        u5_mult_87_CARRYB_23__23_), .CI(u5_mult_87_SUMB_23__24_), .CO(
        u5_mult_87_CARRYB_24__23_), .S(u5_mult_87_SUMB_24__23_) );
  FA_X1 u5_mult_87_S2_24_22 ( .A(u5_mult_87_ab_24__22_), .B(
        u5_mult_87_CARRYB_23__22_), .CI(u5_mult_87_SUMB_23__23_), .CO(
        u5_mult_87_CARRYB_24__22_), .S(u5_mult_87_SUMB_24__22_) );
  FA_X1 u5_mult_87_S2_24_21 ( .A(u5_mult_87_ab_24__21_), .B(
        u5_mult_87_CARRYB_23__21_), .CI(u5_mult_87_SUMB_23__22_), .CO(
        u5_mult_87_CARRYB_24__21_), .S(u5_mult_87_SUMB_24__21_) );
  FA_X1 u5_mult_87_S2_24_20 ( .A(u5_mult_87_ab_24__20_), .B(
        u5_mult_87_CARRYB_23__20_), .CI(u5_mult_87_SUMB_23__21_), .CO(
        u5_mult_87_CARRYB_24__20_), .S(u5_mult_87_SUMB_24__20_) );
  FA_X1 u5_mult_87_S2_24_19 ( .A(u5_mult_87_ab_24__19_), .B(
        u5_mult_87_CARRYB_23__19_), .CI(u5_mult_87_SUMB_23__20_), .CO(
        u5_mult_87_CARRYB_24__19_), .S(u5_mult_87_SUMB_24__19_) );
  FA_X1 u5_mult_87_S2_24_18 ( .A(u5_mult_87_ab_24__18_), .B(
        u5_mult_87_CARRYB_23__18_), .CI(u5_mult_87_SUMB_23__19_), .CO(
        u5_mult_87_CARRYB_24__18_), .S(u5_mult_87_SUMB_24__18_) );
  FA_X1 u5_mult_87_S2_24_17 ( .A(u5_mult_87_ab_24__17_), .B(
        u5_mult_87_CARRYB_23__17_), .CI(u5_mult_87_SUMB_23__18_), .CO(
        u5_mult_87_CARRYB_24__17_), .S(u5_mult_87_SUMB_24__17_) );
  FA_X1 u5_mult_87_S2_24_16 ( .A(u5_mult_87_ab_24__16_), .B(
        u5_mult_87_CARRYB_23__16_), .CI(u5_mult_87_SUMB_23__17_), .CO(
        u5_mult_87_CARRYB_24__16_), .S(u5_mult_87_SUMB_24__16_) );
  FA_X1 u5_mult_87_S2_24_15 ( .A(u5_mult_87_ab_24__15_), .B(
        u5_mult_87_CARRYB_23__15_), .CI(u5_mult_87_SUMB_23__16_), .CO(
        u5_mult_87_CARRYB_24__15_), .S(u5_mult_87_SUMB_24__15_) );
  FA_X1 u5_mult_87_S2_24_14 ( .A(u5_mult_87_ab_24__14_), .B(
        u5_mult_87_CARRYB_23__14_), .CI(u5_mult_87_SUMB_23__15_), .CO(
        u5_mult_87_CARRYB_24__14_), .S(u5_mult_87_SUMB_24__14_) );
  FA_X1 u5_mult_87_S2_24_13 ( .A(u5_mult_87_ab_24__13_), .B(
        u5_mult_87_CARRYB_23__13_), .CI(u5_mult_87_SUMB_23__14_), .CO(
        u5_mult_87_CARRYB_24__13_), .S(u5_mult_87_SUMB_24__13_) );
  FA_X1 u5_mult_87_S2_24_12 ( .A(u5_mult_87_ab_24__12_), .B(
        u5_mult_87_CARRYB_23__12_), .CI(u5_mult_87_SUMB_23__13_), .CO(
        u5_mult_87_CARRYB_24__12_), .S(u5_mult_87_SUMB_24__12_) );
  FA_X1 u5_mult_87_S2_24_11 ( .A(u5_mult_87_ab_24__11_), .B(
        u5_mult_87_CARRYB_23__11_), .CI(u5_mult_87_SUMB_23__12_), .CO(
        u5_mult_87_CARRYB_24__11_), .S(u5_mult_87_SUMB_24__11_) );
  FA_X1 u5_mult_87_S2_24_10 ( .A(u5_mult_87_ab_24__10_), .B(
        u5_mult_87_CARRYB_23__10_), .CI(u5_mult_87_SUMB_23__11_), .CO(
        u5_mult_87_CARRYB_24__10_), .S(u5_mult_87_SUMB_24__10_) );
  FA_X1 u5_mult_87_S2_24_9 ( .A(u5_mult_87_ab_24__9_), .B(
        u5_mult_87_CARRYB_23__9_), .CI(u5_mult_87_SUMB_23__10_), .CO(
        u5_mult_87_CARRYB_24__9_), .S(u5_mult_87_SUMB_24__9_) );
  FA_X1 u5_mult_87_S2_24_8 ( .A(u5_mult_87_ab_24__8_), .B(
        u5_mult_87_CARRYB_23__8_), .CI(u5_mult_87_SUMB_23__9_), .CO(
        u5_mult_87_CARRYB_24__8_), .S(u5_mult_87_SUMB_24__8_) );
  FA_X1 u5_mult_87_S2_24_7 ( .A(u5_mult_87_ab_24__7_), .B(
        u5_mult_87_CARRYB_23__7_), .CI(u5_mult_87_SUMB_23__8_), .CO(
        u5_mult_87_CARRYB_24__7_), .S(u5_mult_87_SUMB_24__7_) );
  FA_X1 u5_mult_87_S2_24_6 ( .A(u5_mult_87_ab_24__6_), .B(
        u5_mult_87_CARRYB_23__6_), .CI(u5_mult_87_SUMB_23__7_), .CO(
        u5_mult_87_CARRYB_24__6_), .S(u5_mult_87_SUMB_24__6_) );
  FA_X1 u5_mult_87_S2_24_5 ( .A(u5_mult_87_ab_24__5_), .B(
        u5_mult_87_CARRYB_23__5_), .CI(u5_mult_87_SUMB_23__6_), .CO(
        u5_mult_87_CARRYB_24__5_), .S(u5_mult_87_SUMB_24__5_) );
  FA_X1 u5_mult_87_S2_24_4 ( .A(u5_mult_87_ab_24__4_), .B(
        u5_mult_87_CARRYB_23__4_), .CI(u5_mult_87_SUMB_23__5_), .CO(
        u5_mult_87_CARRYB_24__4_), .S(u5_mult_87_SUMB_24__4_) );
  FA_X1 u5_mult_87_S2_24_3 ( .A(u5_mult_87_ab_24__3_), .B(
        u5_mult_87_CARRYB_23__3_), .CI(u5_mult_87_SUMB_23__4_), .CO(
        u5_mult_87_CARRYB_24__3_), .S(u5_mult_87_SUMB_24__3_) );
  FA_X1 u5_mult_87_S2_24_2 ( .A(u5_mult_87_ab_24__2_), .B(
        u5_mult_87_CARRYB_23__2_), .CI(u5_mult_87_SUMB_23__3_), .CO(
        u5_mult_87_CARRYB_24__2_), .S(u5_mult_87_SUMB_24__2_) );
  FA_X1 u5_mult_87_S2_24_1 ( .A(u5_mult_87_ab_24__1_), .B(
        u5_mult_87_CARRYB_23__1_), .CI(u5_mult_87_SUMB_23__2_), .CO(
        u5_mult_87_CARRYB_24__1_), .S(u5_mult_87_SUMB_24__1_) );
  FA_X1 u5_mult_87_S1_24_0 ( .A(u5_mult_87_ab_24__0_), .B(
        u5_mult_87_CARRYB_23__0_), .CI(u5_mult_87_SUMB_23__1_), .CO(
        u5_mult_87_CARRYB_24__0_), .S(u5_N24) );
  FA_X1 u5_mult_87_S3_25_51 ( .A(u5_mult_87_ab_25__51_), .B(
        u5_mult_87_CARRYB_24__51_), .CI(u5_mult_87_ab_24__52_), .CO(
        u5_mult_87_CARRYB_25__51_), .S(u5_mult_87_SUMB_25__51_) );
  FA_X1 u5_mult_87_S2_25_50 ( .A(u5_mult_87_ab_25__50_), .B(
        u5_mult_87_CARRYB_24__50_), .CI(u5_mult_87_SUMB_24__51_), .CO(
        u5_mult_87_CARRYB_25__50_), .S(u5_mult_87_SUMB_25__50_) );
  FA_X1 u5_mult_87_S2_25_49 ( .A(u5_mult_87_ab_25__49_), .B(
        u5_mult_87_CARRYB_24__49_), .CI(u5_mult_87_SUMB_24__50_), .CO(
        u5_mult_87_CARRYB_25__49_), .S(u5_mult_87_SUMB_25__49_) );
  FA_X1 u5_mult_87_S2_25_48 ( .A(u5_mult_87_ab_25__48_), .B(
        u5_mult_87_CARRYB_24__48_), .CI(u5_mult_87_SUMB_24__49_), .CO(
        u5_mult_87_CARRYB_25__48_), .S(u5_mult_87_SUMB_25__48_) );
  FA_X1 u5_mult_87_S2_25_47 ( .A(u5_mult_87_ab_25__47_), .B(
        u5_mult_87_CARRYB_24__47_), .CI(u5_mult_87_SUMB_24__48_), .CO(
        u5_mult_87_CARRYB_25__47_), .S(u5_mult_87_SUMB_25__47_) );
  FA_X1 u5_mult_87_S2_25_46 ( .A(u5_mult_87_ab_25__46_), .B(
        u5_mult_87_CARRYB_24__46_), .CI(u5_mult_87_SUMB_24__47_), .CO(
        u5_mult_87_CARRYB_25__46_), .S(u5_mult_87_SUMB_25__46_) );
  FA_X1 u5_mult_87_S2_25_45 ( .A(u5_mult_87_ab_25__45_), .B(
        u5_mult_87_CARRYB_24__45_), .CI(u5_mult_87_SUMB_24__46_), .CO(
        u5_mult_87_CARRYB_25__45_), .S(u5_mult_87_SUMB_25__45_) );
  FA_X1 u5_mult_87_S2_25_44 ( .A(u5_mult_87_ab_25__44_), .B(
        u5_mult_87_CARRYB_24__44_), .CI(u5_mult_87_SUMB_24__45_), .CO(
        u5_mult_87_CARRYB_25__44_), .S(u5_mult_87_SUMB_25__44_) );
  FA_X1 u5_mult_87_S2_25_43 ( .A(u5_mult_87_ab_25__43_), .B(
        u5_mult_87_CARRYB_24__43_), .CI(u5_mult_87_SUMB_24__44_), .CO(
        u5_mult_87_CARRYB_25__43_), .S(u5_mult_87_SUMB_25__43_) );
  FA_X1 u5_mult_87_S2_25_42 ( .A(u5_mult_87_ab_25__42_), .B(
        u5_mult_87_CARRYB_24__42_), .CI(u5_mult_87_SUMB_24__43_), .CO(
        u5_mult_87_CARRYB_25__42_), .S(u5_mult_87_SUMB_25__42_) );
  FA_X1 u5_mult_87_S2_25_41 ( .A(u5_mult_87_ab_25__41_), .B(
        u5_mult_87_CARRYB_24__41_), .CI(u5_mult_87_SUMB_24__42_), .CO(
        u5_mult_87_CARRYB_25__41_), .S(u5_mult_87_SUMB_25__41_) );
  FA_X1 u5_mult_87_S2_25_40 ( .A(u5_mult_87_ab_25__40_), .B(
        u5_mult_87_CARRYB_24__40_), .CI(u5_mult_87_SUMB_24__41_), .CO(
        u5_mult_87_CARRYB_25__40_), .S(u5_mult_87_SUMB_25__40_) );
  FA_X1 u5_mult_87_S2_25_39 ( .A(u5_mult_87_ab_25__39_), .B(
        u5_mult_87_CARRYB_24__39_), .CI(u5_mult_87_SUMB_24__40_), .CO(
        u5_mult_87_CARRYB_25__39_), .S(u5_mult_87_SUMB_25__39_) );
  FA_X1 u5_mult_87_S2_25_38 ( .A(u5_mult_87_ab_25__38_), .B(
        u5_mult_87_CARRYB_24__38_), .CI(u5_mult_87_SUMB_24__39_), .CO(
        u5_mult_87_CARRYB_25__38_), .S(u5_mult_87_SUMB_25__38_) );
  FA_X1 u5_mult_87_S2_25_37 ( .A(u5_mult_87_ab_25__37_), .B(
        u5_mult_87_CARRYB_24__37_), .CI(u5_mult_87_SUMB_24__38_), .CO(
        u5_mult_87_CARRYB_25__37_), .S(u5_mult_87_SUMB_25__37_) );
  FA_X1 u5_mult_87_S2_25_36 ( .A(u5_mult_87_ab_25__36_), .B(
        u5_mult_87_CARRYB_24__36_), .CI(u5_mult_87_SUMB_24__37_), .CO(
        u5_mult_87_CARRYB_25__36_), .S(u5_mult_87_SUMB_25__36_) );
  FA_X1 u5_mult_87_S2_25_35 ( .A(u5_mult_87_ab_25__35_), .B(
        u5_mult_87_CARRYB_24__35_), .CI(u5_mult_87_SUMB_24__36_), .CO(
        u5_mult_87_CARRYB_25__35_), .S(u5_mult_87_SUMB_25__35_) );
  FA_X1 u5_mult_87_S2_25_34 ( .A(u5_mult_87_ab_25__34_), .B(
        u5_mult_87_CARRYB_24__34_), .CI(u5_mult_87_SUMB_24__35_), .CO(
        u5_mult_87_CARRYB_25__34_), .S(u5_mult_87_SUMB_25__34_) );
  FA_X1 u5_mult_87_S2_25_33 ( .A(u5_mult_87_ab_25__33_), .B(
        u5_mult_87_CARRYB_24__33_), .CI(u5_mult_87_SUMB_24__34_), .CO(
        u5_mult_87_CARRYB_25__33_), .S(u5_mult_87_SUMB_25__33_) );
  FA_X1 u5_mult_87_S2_25_32 ( .A(u5_mult_87_ab_25__32_), .B(
        u5_mult_87_CARRYB_24__32_), .CI(u5_mult_87_SUMB_24__33_), .CO(
        u5_mult_87_CARRYB_25__32_), .S(u5_mult_87_SUMB_25__32_) );
  FA_X1 u5_mult_87_S2_25_31 ( .A(u5_mult_87_ab_25__31_), .B(
        u5_mult_87_CARRYB_24__31_), .CI(u5_mult_87_SUMB_24__32_), .CO(
        u5_mult_87_CARRYB_25__31_), .S(u5_mult_87_SUMB_25__31_) );
  FA_X1 u5_mult_87_S2_25_30 ( .A(u5_mult_87_ab_25__30_), .B(
        u5_mult_87_CARRYB_24__30_), .CI(u5_mult_87_SUMB_24__31_), .CO(
        u5_mult_87_CARRYB_25__30_), .S(u5_mult_87_SUMB_25__30_) );
  FA_X1 u5_mult_87_S2_25_29 ( .A(u5_mult_87_ab_25__29_), .B(
        u5_mult_87_CARRYB_24__29_), .CI(u5_mult_87_SUMB_24__30_), .CO(
        u5_mult_87_CARRYB_25__29_), .S(u5_mult_87_SUMB_25__29_) );
  FA_X1 u5_mult_87_S2_25_28 ( .A(u5_mult_87_ab_25__28_), .B(
        u5_mult_87_CARRYB_24__28_), .CI(u5_mult_87_SUMB_24__29_), .CO(
        u5_mult_87_CARRYB_25__28_), .S(u5_mult_87_SUMB_25__28_) );
  FA_X1 u5_mult_87_S2_25_27 ( .A(u5_mult_87_ab_25__27_), .B(
        u5_mult_87_CARRYB_24__27_), .CI(u5_mult_87_SUMB_24__28_), .CO(
        u5_mult_87_CARRYB_25__27_), .S(u5_mult_87_SUMB_25__27_) );
  FA_X1 u5_mult_87_S2_25_26 ( .A(u5_mult_87_ab_25__26_), .B(
        u5_mult_87_CARRYB_24__26_), .CI(u5_mult_87_SUMB_24__27_), .CO(
        u5_mult_87_CARRYB_25__26_), .S(u5_mult_87_SUMB_25__26_) );
  FA_X1 u5_mult_87_S2_25_25 ( .A(u5_mult_87_ab_25__25_), .B(
        u5_mult_87_CARRYB_24__25_), .CI(u5_mult_87_SUMB_24__26_), .CO(
        u5_mult_87_CARRYB_25__25_), .S(u5_mult_87_SUMB_25__25_) );
  FA_X1 u5_mult_87_S2_25_24 ( .A(u5_mult_87_ab_25__24_), .B(
        u5_mult_87_CARRYB_24__24_), .CI(u5_mult_87_SUMB_24__25_), .CO(
        u5_mult_87_CARRYB_25__24_), .S(u5_mult_87_SUMB_25__24_) );
  FA_X1 u5_mult_87_S2_25_23 ( .A(u5_mult_87_ab_25__23_), .B(
        u5_mult_87_CARRYB_24__23_), .CI(u5_mult_87_SUMB_24__24_), .CO(
        u5_mult_87_CARRYB_25__23_), .S(u5_mult_87_SUMB_25__23_) );
  FA_X1 u5_mult_87_S2_25_22 ( .A(u5_mult_87_ab_25__22_), .B(
        u5_mult_87_CARRYB_24__22_), .CI(u5_mult_87_SUMB_24__23_), .CO(
        u5_mult_87_CARRYB_25__22_), .S(u5_mult_87_SUMB_25__22_) );
  FA_X1 u5_mult_87_S2_25_21 ( .A(u5_mult_87_ab_25__21_), .B(
        u5_mult_87_CARRYB_24__21_), .CI(u5_mult_87_SUMB_24__22_), .CO(
        u5_mult_87_CARRYB_25__21_), .S(u5_mult_87_SUMB_25__21_) );
  FA_X1 u5_mult_87_S2_25_20 ( .A(u5_mult_87_ab_25__20_), .B(
        u5_mult_87_CARRYB_24__20_), .CI(u5_mult_87_SUMB_24__21_), .CO(
        u5_mult_87_CARRYB_25__20_), .S(u5_mult_87_SUMB_25__20_) );
  FA_X1 u5_mult_87_S2_25_19 ( .A(u5_mult_87_ab_25__19_), .B(
        u5_mult_87_CARRYB_24__19_), .CI(u5_mult_87_SUMB_24__20_), .CO(
        u5_mult_87_CARRYB_25__19_), .S(u5_mult_87_SUMB_25__19_) );
  FA_X1 u5_mult_87_S2_25_18 ( .A(u5_mult_87_ab_25__18_), .B(
        u5_mult_87_CARRYB_24__18_), .CI(u5_mult_87_SUMB_24__19_), .CO(
        u5_mult_87_CARRYB_25__18_), .S(u5_mult_87_SUMB_25__18_) );
  FA_X1 u5_mult_87_S2_25_17 ( .A(u5_mult_87_ab_25__17_), .B(
        u5_mult_87_CARRYB_24__17_), .CI(u5_mult_87_SUMB_24__18_), .CO(
        u5_mult_87_CARRYB_25__17_), .S(u5_mult_87_SUMB_25__17_) );
  FA_X1 u5_mult_87_S2_25_16 ( .A(u5_mult_87_ab_25__16_), .B(
        u5_mult_87_CARRYB_24__16_), .CI(u5_mult_87_SUMB_24__17_), .CO(
        u5_mult_87_CARRYB_25__16_), .S(u5_mult_87_SUMB_25__16_) );
  FA_X1 u5_mult_87_S2_25_15 ( .A(u5_mult_87_ab_25__15_), .B(
        u5_mult_87_CARRYB_24__15_), .CI(u5_mult_87_SUMB_24__16_), .CO(
        u5_mult_87_CARRYB_25__15_), .S(u5_mult_87_SUMB_25__15_) );
  FA_X1 u5_mult_87_S2_25_14 ( .A(u5_mult_87_ab_25__14_), .B(
        u5_mult_87_CARRYB_24__14_), .CI(u5_mult_87_SUMB_24__15_), .CO(
        u5_mult_87_CARRYB_25__14_), .S(u5_mult_87_SUMB_25__14_) );
  FA_X1 u5_mult_87_S2_25_13 ( .A(u5_mult_87_ab_25__13_), .B(
        u5_mult_87_CARRYB_24__13_), .CI(u5_mult_87_SUMB_24__14_), .CO(
        u5_mult_87_CARRYB_25__13_), .S(u5_mult_87_SUMB_25__13_) );
  FA_X1 u5_mult_87_S2_25_12 ( .A(u5_mult_87_ab_25__12_), .B(
        u5_mult_87_CARRYB_24__12_), .CI(u5_mult_87_SUMB_24__13_), .CO(
        u5_mult_87_CARRYB_25__12_), .S(u5_mult_87_SUMB_25__12_) );
  FA_X1 u5_mult_87_S2_25_11 ( .A(u5_mult_87_ab_25__11_), .B(
        u5_mult_87_CARRYB_24__11_), .CI(u5_mult_87_SUMB_24__12_), .CO(
        u5_mult_87_CARRYB_25__11_), .S(u5_mult_87_SUMB_25__11_) );
  FA_X1 u5_mult_87_S2_25_10 ( .A(u5_mult_87_ab_25__10_), .B(
        u5_mult_87_CARRYB_24__10_), .CI(u5_mult_87_SUMB_24__11_), .CO(
        u5_mult_87_CARRYB_25__10_), .S(u5_mult_87_SUMB_25__10_) );
  FA_X1 u5_mult_87_S2_25_9 ( .A(u5_mult_87_ab_25__9_), .B(
        u5_mult_87_CARRYB_24__9_), .CI(u5_mult_87_SUMB_24__10_), .CO(
        u5_mult_87_CARRYB_25__9_), .S(u5_mult_87_SUMB_25__9_) );
  FA_X1 u5_mult_87_S2_25_8 ( .A(u5_mult_87_ab_25__8_), .B(
        u5_mult_87_CARRYB_24__8_), .CI(u5_mult_87_SUMB_24__9_), .CO(
        u5_mult_87_CARRYB_25__8_), .S(u5_mult_87_SUMB_25__8_) );
  FA_X1 u5_mult_87_S2_25_7 ( .A(u5_mult_87_ab_25__7_), .B(
        u5_mult_87_CARRYB_24__7_), .CI(u5_mult_87_SUMB_24__8_), .CO(
        u5_mult_87_CARRYB_25__7_), .S(u5_mult_87_SUMB_25__7_) );
  FA_X1 u5_mult_87_S2_25_6 ( .A(u5_mult_87_ab_25__6_), .B(
        u5_mult_87_CARRYB_24__6_), .CI(u5_mult_87_SUMB_24__7_), .CO(
        u5_mult_87_CARRYB_25__6_), .S(u5_mult_87_SUMB_25__6_) );
  FA_X1 u5_mult_87_S2_25_5 ( .A(u5_mult_87_ab_25__5_), .B(
        u5_mult_87_CARRYB_24__5_), .CI(u5_mult_87_SUMB_24__6_), .CO(
        u5_mult_87_CARRYB_25__5_), .S(u5_mult_87_SUMB_25__5_) );
  FA_X1 u5_mult_87_S2_25_4 ( .A(u5_mult_87_ab_25__4_), .B(
        u5_mult_87_CARRYB_24__4_), .CI(u5_mult_87_SUMB_24__5_), .CO(
        u5_mult_87_CARRYB_25__4_), .S(u5_mult_87_SUMB_25__4_) );
  FA_X1 u5_mult_87_S2_25_3 ( .A(u5_mult_87_ab_25__3_), .B(
        u5_mult_87_CARRYB_24__3_), .CI(u5_mult_87_SUMB_24__4_), .CO(
        u5_mult_87_CARRYB_25__3_), .S(u5_mult_87_SUMB_25__3_) );
  FA_X1 u5_mult_87_S2_25_2 ( .A(u5_mult_87_ab_25__2_), .B(
        u5_mult_87_CARRYB_24__2_), .CI(u5_mult_87_SUMB_24__3_), .CO(
        u5_mult_87_CARRYB_25__2_), .S(u5_mult_87_SUMB_25__2_) );
  FA_X1 u5_mult_87_S2_25_1 ( .A(u5_mult_87_ab_25__1_), .B(
        u5_mult_87_CARRYB_24__1_), .CI(u5_mult_87_SUMB_24__2_), .CO(
        u5_mult_87_CARRYB_25__1_), .S(u5_mult_87_SUMB_25__1_) );
  FA_X1 u5_mult_87_S1_25_0 ( .A(u5_mult_87_ab_25__0_), .B(
        u5_mult_87_CARRYB_24__0_), .CI(u5_mult_87_SUMB_24__1_), .CO(
        u5_mult_87_CARRYB_25__0_), .S(u5_N25) );
  FA_X1 u5_mult_87_S3_26_51 ( .A(u5_mult_87_ab_26__51_), .B(
        u5_mult_87_CARRYB_25__51_), .CI(u5_mult_87_ab_25__52_), .CO(
        u5_mult_87_CARRYB_26__51_), .S(u5_mult_87_SUMB_26__51_) );
  FA_X1 u5_mult_87_S2_26_50 ( .A(u5_mult_87_ab_26__50_), .B(
        u5_mult_87_CARRYB_25__50_), .CI(u5_mult_87_SUMB_25__51_), .CO(
        u5_mult_87_CARRYB_26__50_), .S(u5_mult_87_SUMB_26__50_) );
  FA_X1 u5_mult_87_S2_26_49 ( .A(u5_mult_87_ab_26__49_), .B(
        u5_mult_87_CARRYB_25__49_), .CI(u5_mult_87_SUMB_25__50_), .CO(
        u5_mult_87_CARRYB_26__49_), .S(u5_mult_87_SUMB_26__49_) );
  FA_X1 u5_mult_87_S2_26_48 ( .A(u5_mult_87_ab_26__48_), .B(
        u5_mult_87_CARRYB_25__48_), .CI(u5_mult_87_SUMB_25__49_), .CO(
        u5_mult_87_CARRYB_26__48_), .S(u5_mult_87_SUMB_26__48_) );
  FA_X1 u5_mult_87_S2_26_47 ( .A(u5_mult_87_ab_26__47_), .B(
        u5_mult_87_CARRYB_25__47_), .CI(u5_mult_87_SUMB_25__48_), .CO(
        u5_mult_87_CARRYB_26__47_), .S(u5_mult_87_SUMB_26__47_) );
  FA_X1 u5_mult_87_S2_26_46 ( .A(u5_mult_87_ab_26__46_), .B(
        u5_mult_87_CARRYB_25__46_), .CI(u5_mult_87_SUMB_25__47_), .CO(
        u5_mult_87_CARRYB_26__46_), .S(u5_mult_87_SUMB_26__46_) );
  FA_X1 u5_mult_87_S2_26_45 ( .A(u5_mult_87_ab_26__45_), .B(
        u5_mult_87_CARRYB_25__45_), .CI(u5_mult_87_SUMB_25__46_), .CO(
        u5_mult_87_CARRYB_26__45_), .S(u5_mult_87_SUMB_26__45_) );
  FA_X1 u5_mult_87_S2_26_44 ( .A(u5_mult_87_ab_26__44_), .B(
        u5_mult_87_CARRYB_25__44_), .CI(u5_mult_87_SUMB_25__45_), .CO(
        u5_mult_87_CARRYB_26__44_), .S(u5_mult_87_SUMB_26__44_) );
  FA_X1 u5_mult_87_S2_26_43 ( .A(u5_mult_87_ab_26__43_), .B(
        u5_mult_87_CARRYB_25__43_), .CI(u5_mult_87_SUMB_25__44_), .CO(
        u5_mult_87_CARRYB_26__43_), .S(u5_mult_87_SUMB_26__43_) );
  FA_X1 u5_mult_87_S2_26_42 ( .A(u5_mult_87_ab_26__42_), .B(
        u5_mult_87_CARRYB_25__42_), .CI(u5_mult_87_SUMB_25__43_), .CO(
        u5_mult_87_CARRYB_26__42_), .S(u5_mult_87_SUMB_26__42_) );
  FA_X1 u5_mult_87_S2_26_41 ( .A(u5_mult_87_ab_26__41_), .B(
        u5_mult_87_CARRYB_25__41_), .CI(u5_mult_87_SUMB_25__42_), .CO(
        u5_mult_87_CARRYB_26__41_), .S(u5_mult_87_SUMB_26__41_) );
  FA_X1 u5_mult_87_S2_26_40 ( .A(u5_mult_87_ab_26__40_), .B(
        u5_mult_87_CARRYB_25__40_), .CI(u5_mult_87_SUMB_25__41_), .CO(
        u5_mult_87_CARRYB_26__40_), .S(u5_mult_87_SUMB_26__40_) );
  FA_X1 u5_mult_87_S2_26_39 ( .A(u5_mult_87_ab_26__39_), .B(
        u5_mult_87_CARRYB_25__39_), .CI(u5_mult_87_SUMB_25__40_), .CO(
        u5_mult_87_CARRYB_26__39_), .S(u5_mult_87_SUMB_26__39_) );
  FA_X1 u5_mult_87_S2_26_38 ( .A(u5_mult_87_ab_26__38_), .B(
        u5_mult_87_CARRYB_25__38_), .CI(u5_mult_87_SUMB_25__39_), .CO(
        u5_mult_87_CARRYB_26__38_), .S(u5_mult_87_SUMB_26__38_) );
  FA_X1 u5_mult_87_S2_26_37 ( .A(u5_mult_87_ab_26__37_), .B(
        u5_mult_87_CARRYB_25__37_), .CI(u5_mult_87_SUMB_25__38_), .CO(
        u5_mult_87_CARRYB_26__37_), .S(u5_mult_87_SUMB_26__37_) );
  FA_X1 u5_mult_87_S2_26_36 ( .A(u5_mult_87_ab_26__36_), .B(
        u5_mult_87_CARRYB_25__36_), .CI(u5_mult_87_SUMB_25__37_), .CO(
        u5_mult_87_CARRYB_26__36_), .S(u5_mult_87_SUMB_26__36_) );
  FA_X1 u5_mult_87_S2_26_35 ( .A(u5_mult_87_ab_26__35_), .B(
        u5_mult_87_CARRYB_25__35_), .CI(u5_mult_87_SUMB_25__36_), .CO(
        u5_mult_87_CARRYB_26__35_), .S(u5_mult_87_SUMB_26__35_) );
  FA_X1 u5_mult_87_S2_26_34 ( .A(u5_mult_87_ab_26__34_), .B(
        u5_mult_87_CARRYB_25__34_), .CI(u5_mult_87_SUMB_25__35_), .CO(
        u5_mult_87_CARRYB_26__34_), .S(u5_mult_87_SUMB_26__34_) );
  FA_X1 u5_mult_87_S2_26_33 ( .A(u5_mult_87_ab_26__33_), .B(
        u5_mult_87_CARRYB_25__33_), .CI(u5_mult_87_SUMB_25__34_), .CO(
        u5_mult_87_CARRYB_26__33_), .S(u5_mult_87_SUMB_26__33_) );
  FA_X1 u5_mult_87_S2_26_32 ( .A(u5_mult_87_ab_26__32_), .B(
        u5_mult_87_CARRYB_25__32_), .CI(u5_mult_87_SUMB_25__33_), .CO(
        u5_mult_87_CARRYB_26__32_), .S(u5_mult_87_SUMB_26__32_) );
  FA_X1 u5_mult_87_S2_26_31 ( .A(u5_mult_87_ab_26__31_), .B(
        u5_mult_87_CARRYB_25__31_), .CI(u5_mult_87_SUMB_25__32_), .CO(
        u5_mult_87_CARRYB_26__31_), .S(u5_mult_87_SUMB_26__31_) );
  FA_X1 u5_mult_87_S2_26_30 ( .A(u5_mult_87_ab_26__30_), .B(
        u5_mult_87_CARRYB_25__30_), .CI(u5_mult_87_SUMB_25__31_), .CO(
        u5_mult_87_CARRYB_26__30_), .S(u5_mult_87_SUMB_26__30_) );
  FA_X1 u5_mult_87_S2_26_29 ( .A(u5_mult_87_ab_26__29_), .B(
        u5_mult_87_CARRYB_25__29_), .CI(u5_mult_87_SUMB_25__30_), .CO(
        u5_mult_87_CARRYB_26__29_), .S(u5_mult_87_SUMB_26__29_) );
  FA_X1 u5_mult_87_S2_26_28 ( .A(u5_mult_87_ab_26__28_), .B(
        u5_mult_87_CARRYB_25__28_), .CI(u5_mult_87_SUMB_25__29_), .CO(
        u5_mult_87_CARRYB_26__28_), .S(u5_mult_87_SUMB_26__28_) );
  FA_X1 u5_mult_87_S2_26_27 ( .A(u5_mult_87_ab_26__27_), .B(
        u5_mult_87_CARRYB_25__27_), .CI(u5_mult_87_SUMB_25__28_), .CO(
        u5_mult_87_CARRYB_26__27_), .S(u5_mult_87_SUMB_26__27_) );
  FA_X1 u5_mult_87_S2_26_26 ( .A(u5_mult_87_ab_26__26_), .B(
        u5_mult_87_CARRYB_25__26_), .CI(u5_mult_87_SUMB_25__27_), .CO(
        u5_mult_87_CARRYB_26__26_), .S(u5_mult_87_SUMB_26__26_) );
  FA_X1 u5_mult_87_S2_26_25 ( .A(u5_mult_87_ab_26__25_), .B(
        u5_mult_87_CARRYB_25__25_), .CI(u5_mult_87_SUMB_25__26_), .CO(
        u5_mult_87_CARRYB_26__25_), .S(u5_mult_87_SUMB_26__25_) );
  FA_X1 u5_mult_87_S2_26_24 ( .A(u5_mult_87_ab_26__24_), .B(
        u5_mult_87_CARRYB_25__24_), .CI(u5_mult_87_SUMB_25__25_), .CO(
        u5_mult_87_CARRYB_26__24_), .S(u5_mult_87_SUMB_26__24_) );
  FA_X1 u5_mult_87_S2_26_23 ( .A(u5_mult_87_ab_26__23_), .B(
        u5_mult_87_CARRYB_25__23_), .CI(u5_mult_87_SUMB_25__24_), .CO(
        u5_mult_87_CARRYB_26__23_), .S(u5_mult_87_SUMB_26__23_) );
  FA_X1 u5_mult_87_S2_26_22 ( .A(u5_mult_87_ab_26__22_), .B(
        u5_mult_87_CARRYB_25__22_), .CI(u5_mult_87_SUMB_25__23_), .CO(
        u5_mult_87_CARRYB_26__22_), .S(u5_mult_87_SUMB_26__22_) );
  FA_X1 u5_mult_87_S2_26_21 ( .A(u5_mult_87_ab_26__21_), .B(
        u5_mult_87_CARRYB_25__21_), .CI(u5_mult_87_SUMB_25__22_), .CO(
        u5_mult_87_CARRYB_26__21_), .S(u5_mult_87_SUMB_26__21_) );
  FA_X1 u5_mult_87_S2_26_20 ( .A(u5_mult_87_ab_26__20_), .B(
        u5_mult_87_CARRYB_25__20_), .CI(u5_mult_87_SUMB_25__21_), .CO(
        u5_mult_87_CARRYB_26__20_), .S(u5_mult_87_SUMB_26__20_) );
  FA_X1 u5_mult_87_S2_26_19 ( .A(u5_mult_87_ab_26__19_), .B(
        u5_mult_87_CARRYB_25__19_), .CI(u5_mult_87_SUMB_25__20_), .CO(
        u5_mult_87_CARRYB_26__19_), .S(u5_mult_87_SUMB_26__19_) );
  FA_X1 u5_mult_87_S2_26_18 ( .A(u5_mult_87_ab_26__18_), .B(
        u5_mult_87_CARRYB_25__18_), .CI(u5_mult_87_SUMB_25__19_), .CO(
        u5_mult_87_CARRYB_26__18_), .S(u5_mult_87_SUMB_26__18_) );
  FA_X1 u5_mult_87_S2_26_17 ( .A(u5_mult_87_ab_26__17_), .B(
        u5_mult_87_CARRYB_25__17_), .CI(u5_mult_87_SUMB_25__18_), .CO(
        u5_mult_87_CARRYB_26__17_), .S(u5_mult_87_SUMB_26__17_) );
  FA_X1 u5_mult_87_S2_26_16 ( .A(u5_mult_87_ab_26__16_), .B(
        u5_mult_87_CARRYB_25__16_), .CI(u5_mult_87_SUMB_25__17_), .CO(
        u5_mult_87_CARRYB_26__16_), .S(u5_mult_87_SUMB_26__16_) );
  FA_X1 u5_mult_87_S2_26_15 ( .A(u5_mult_87_ab_26__15_), .B(
        u5_mult_87_CARRYB_25__15_), .CI(u5_mult_87_SUMB_25__16_), .CO(
        u5_mult_87_CARRYB_26__15_), .S(u5_mult_87_SUMB_26__15_) );
  FA_X1 u5_mult_87_S2_26_14 ( .A(u5_mult_87_ab_26__14_), .B(
        u5_mult_87_CARRYB_25__14_), .CI(u5_mult_87_SUMB_25__15_), .CO(
        u5_mult_87_CARRYB_26__14_), .S(u5_mult_87_SUMB_26__14_) );
  FA_X1 u5_mult_87_S2_26_13 ( .A(u5_mult_87_ab_26__13_), .B(
        u5_mult_87_CARRYB_25__13_), .CI(u5_mult_87_SUMB_25__14_), .CO(
        u5_mult_87_CARRYB_26__13_), .S(u5_mult_87_SUMB_26__13_) );
  FA_X1 u5_mult_87_S2_26_12 ( .A(u5_mult_87_ab_26__12_), .B(
        u5_mult_87_CARRYB_25__12_), .CI(u5_mult_87_SUMB_25__13_), .CO(
        u5_mult_87_CARRYB_26__12_), .S(u5_mult_87_SUMB_26__12_) );
  FA_X1 u5_mult_87_S2_26_11 ( .A(u5_mult_87_ab_26__11_), .B(
        u5_mult_87_CARRYB_25__11_), .CI(u5_mult_87_SUMB_25__12_), .CO(
        u5_mult_87_CARRYB_26__11_), .S(u5_mult_87_SUMB_26__11_) );
  FA_X1 u5_mult_87_S2_26_10 ( .A(u5_mult_87_ab_26__10_), .B(
        u5_mult_87_CARRYB_25__10_), .CI(u5_mult_87_SUMB_25__11_), .CO(
        u5_mult_87_CARRYB_26__10_), .S(u5_mult_87_SUMB_26__10_) );
  FA_X1 u5_mult_87_S2_26_9 ( .A(u5_mult_87_ab_26__9_), .B(
        u5_mult_87_CARRYB_25__9_), .CI(u5_mult_87_SUMB_25__10_), .CO(
        u5_mult_87_CARRYB_26__9_), .S(u5_mult_87_SUMB_26__9_) );
  FA_X1 u5_mult_87_S2_26_8 ( .A(u5_mult_87_ab_26__8_), .B(
        u5_mult_87_CARRYB_25__8_), .CI(u5_mult_87_SUMB_25__9_), .CO(
        u5_mult_87_CARRYB_26__8_), .S(u5_mult_87_SUMB_26__8_) );
  FA_X1 u5_mult_87_S2_26_7 ( .A(u5_mult_87_ab_26__7_), .B(
        u5_mult_87_CARRYB_25__7_), .CI(u5_mult_87_SUMB_25__8_), .CO(
        u5_mult_87_CARRYB_26__7_), .S(u5_mult_87_SUMB_26__7_) );
  FA_X1 u5_mult_87_S2_26_6 ( .A(u5_mult_87_ab_26__6_), .B(
        u5_mult_87_CARRYB_25__6_), .CI(u5_mult_87_SUMB_25__7_), .CO(
        u5_mult_87_CARRYB_26__6_), .S(u5_mult_87_SUMB_26__6_) );
  FA_X1 u5_mult_87_S2_26_5 ( .A(u5_mult_87_ab_26__5_), .B(
        u5_mult_87_CARRYB_25__5_), .CI(u5_mult_87_SUMB_25__6_), .CO(
        u5_mult_87_CARRYB_26__5_), .S(u5_mult_87_SUMB_26__5_) );
  FA_X1 u5_mult_87_S2_26_4 ( .A(u5_mult_87_ab_26__4_), .B(
        u5_mult_87_CARRYB_25__4_), .CI(u5_mult_87_SUMB_25__5_), .CO(
        u5_mult_87_CARRYB_26__4_), .S(u5_mult_87_SUMB_26__4_) );
  FA_X1 u5_mult_87_S2_26_3 ( .A(u5_mult_87_ab_26__3_), .B(
        u5_mult_87_CARRYB_25__3_), .CI(u5_mult_87_SUMB_25__4_), .CO(
        u5_mult_87_CARRYB_26__3_), .S(u5_mult_87_SUMB_26__3_) );
  FA_X1 u5_mult_87_S2_26_2 ( .A(u5_mult_87_ab_26__2_), .B(
        u5_mult_87_CARRYB_25__2_), .CI(u5_mult_87_SUMB_25__3_), .CO(
        u5_mult_87_CARRYB_26__2_), .S(u5_mult_87_SUMB_26__2_) );
  FA_X1 u5_mult_87_S2_26_1 ( .A(u5_mult_87_ab_26__1_), .B(
        u5_mult_87_CARRYB_25__1_), .CI(u5_mult_87_SUMB_25__2_), .CO(
        u5_mult_87_CARRYB_26__1_), .S(u5_mult_87_SUMB_26__1_) );
  FA_X1 u5_mult_87_S1_26_0 ( .A(u5_mult_87_ab_26__0_), .B(
        u5_mult_87_CARRYB_25__0_), .CI(u5_mult_87_SUMB_25__1_), .CO(
        u5_mult_87_CARRYB_26__0_), .S(u5_N26) );
  FA_X1 u5_mult_87_S3_27_51 ( .A(u5_mult_87_ab_27__51_), .B(
        u5_mult_87_CARRYB_26__51_), .CI(u5_mult_87_ab_26__52_), .CO(
        u5_mult_87_CARRYB_27__51_), .S(u5_mult_87_SUMB_27__51_) );
  FA_X1 u5_mult_87_S2_27_50 ( .A(u5_mult_87_ab_27__50_), .B(
        u5_mult_87_CARRYB_26__50_), .CI(u5_mult_87_SUMB_26__51_), .CO(
        u5_mult_87_CARRYB_27__50_), .S(u5_mult_87_SUMB_27__50_) );
  FA_X1 u5_mult_87_S2_27_49 ( .A(u5_mult_87_ab_27__49_), .B(
        u5_mult_87_CARRYB_26__49_), .CI(u5_mult_87_SUMB_26__50_), .CO(
        u5_mult_87_CARRYB_27__49_), .S(u5_mult_87_SUMB_27__49_) );
  FA_X1 u5_mult_87_S2_27_48 ( .A(u5_mult_87_ab_27__48_), .B(
        u5_mult_87_CARRYB_26__48_), .CI(u5_mult_87_SUMB_26__49_), .CO(
        u5_mult_87_CARRYB_27__48_), .S(u5_mult_87_SUMB_27__48_) );
  FA_X1 u5_mult_87_S2_27_47 ( .A(u5_mult_87_ab_27__47_), .B(
        u5_mult_87_CARRYB_26__47_), .CI(u5_mult_87_SUMB_26__48_), .CO(
        u5_mult_87_CARRYB_27__47_), .S(u5_mult_87_SUMB_27__47_) );
  FA_X1 u5_mult_87_S2_27_46 ( .A(u5_mult_87_ab_27__46_), .B(
        u5_mult_87_CARRYB_26__46_), .CI(u5_mult_87_SUMB_26__47_), .CO(
        u5_mult_87_CARRYB_27__46_), .S(u5_mult_87_SUMB_27__46_) );
  FA_X1 u5_mult_87_S2_27_45 ( .A(u5_mult_87_ab_27__45_), .B(
        u5_mult_87_CARRYB_26__45_), .CI(u5_mult_87_SUMB_26__46_), .CO(
        u5_mult_87_CARRYB_27__45_), .S(u5_mult_87_SUMB_27__45_) );
  FA_X1 u5_mult_87_S2_27_44 ( .A(u5_mult_87_ab_27__44_), .B(
        u5_mult_87_CARRYB_26__44_), .CI(u5_mult_87_SUMB_26__45_), .CO(
        u5_mult_87_CARRYB_27__44_), .S(u5_mult_87_SUMB_27__44_) );
  FA_X1 u5_mult_87_S2_27_43 ( .A(u5_mult_87_ab_27__43_), .B(
        u5_mult_87_CARRYB_26__43_), .CI(u5_mult_87_SUMB_26__44_), .CO(
        u5_mult_87_CARRYB_27__43_), .S(u5_mult_87_SUMB_27__43_) );
  FA_X1 u5_mult_87_S2_27_42 ( .A(u5_mult_87_ab_27__42_), .B(
        u5_mult_87_CARRYB_26__42_), .CI(u5_mult_87_SUMB_26__43_), .CO(
        u5_mult_87_CARRYB_27__42_), .S(u5_mult_87_SUMB_27__42_) );
  FA_X1 u5_mult_87_S2_27_41 ( .A(u5_mult_87_ab_27__41_), .B(
        u5_mult_87_CARRYB_26__41_), .CI(u5_mult_87_SUMB_26__42_), .CO(
        u5_mult_87_CARRYB_27__41_), .S(u5_mult_87_SUMB_27__41_) );
  FA_X1 u5_mult_87_S2_27_40 ( .A(u5_mult_87_ab_27__40_), .B(
        u5_mult_87_CARRYB_26__40_), .CI(u5_mult_87_SUMB_26__41_), .CO(
        u5_mult_87_CARRYB_27__40_), .S(u5_mult_87_SUMB_27__40_) );
  FA_X1 u5_mult_87_S2_27_39 ( .A(u5_mult_87_ab_27__39_), .B(
        u5_mult_87_CARRYB_26__39_), .CI(u5_mult_87_SUMB_26__40_), .CO(
        u5_mult_87_CARRYB_27__39_), .S(u5_mult_87_SUMB_27__39_) );
  FA_X1 u5_mult_87_S2_27_38 ( .A(u5_mult_87_ab_27__38_), .B(
        u5_mult_87_CARRYB_26__38_), .CI(u5_mult_87_SUMB_26__39_), .CO(
        u5_mult_87_CARRYB_27__38_), .S(u5_mult_87_SUMB_27__38_) );
  FA_X1 u5_mult_87_S2_27_37 ( .A(u5_mult_87_ab_27__37_), .B(
        u5_mult_87_CARRYB_26__37_), .CI(u5_mult_87_SUMB_26__38_), .CO(
        u5_mult_87_CARRYB_27__37_), .S(u5_mult_87_SUMB_27__37_) );
  FA_X1 u5_mult_87_S2_27_36 ( .A(u5_mult_87_ab_27__36_), .B(
        u5_mult_87_CARRYB_26__36_), .CI(u5_mult_87_SUMB_26__37_), .CO(
        u5_mult_87_CARRYB_27__36_), .S(u5_mult_87_SUMB_27__36_) );
  FA_X1 u5_mult_87_S2_27_35 ( .A(u5_mult_87_ab_27__35_), .B(
        u5_mult_87_CARRYB_26__35_), .CI(u5_mult_87_SUMB_26__36_), .CO(
        u5_mult_87_CARRYB_27__35_), .S(u5_mult_87_SUMB_27__35_) );
  FA_X1 u5_mult_87_S2_27_34 ( .A(u5_mult_87_ab_27__34_), .B(
        u5_mult_87_CARRYB_26__34_), .CI(u5_mult_87_SUMB_26__35_), .CO(
        u5_mult_87_CARRYB_27__34_), .S(u5_mult_87_SUMB_27__34_) );
  FA_X1 u5_mult_87_S2_27_33 ( .A(u5_mult_87_ab_27__33_), .B(
        u5_mult_87_CARRYB_26__33_), .CI(u5_mult_87_SUMB_26__34_), .CO(
        u5_mult_87_CARRYB_27__33_), .S(u5_mult_87_SUMB_27__33_) );
  FA_X1 u5_mult_87_S2_27_32 ( .A(u5_mult_87_ab_27__32_), .B(
        u5_mult_87_CARRYB_26__32_), .CI(u5_mult_87_SUMB_26__33_), .CO(
        u5_mult_87_CARRYB_27__32_), .S(u5_mult_87_SUMB_27__32_) );
  FA_X1 u5_mult_87_S2_27_31 ( .A(u5_mult_87_ab_27__31_), .B(
        u5_mult_87_CARRYB_26__31_), .CI(u5_mult_87_SUMB_26__32_), .CO(
        u5_mult_87_CARRYB_27__31_), .S(u5_mult_87_SUMB_27__31_) );
  FA_X1 u5_mult_87_S2_27_30 ( .A(u5_mult_87_ab_27__30_), .B(
        u5_mult_87_CARRYB_26__30_), .CI(u5_mult_87_SUMB_26__31_), .CO(
        u5_mult_87_CARRYB_27__30_), .S(u5_mult_87_SUMB_27__30_) );
  FA_X1 u5_mult_87_S2_27_29 ( .A(u5_mult_87_ab_27__29_), .B(
        u5_mult_87_CARRYB_26__29_), .CI(u5_mult_87_SUMB_26__30_), .CO(
        u5_mult_87_CARRYB_27__29_), .S(u5_mult_87_SUMB_27__29_) );
  FA_X1 u5_mult_87_S2_27_28 ( .A(u5_mult_87_ab_27__28_), .B(
        u5_mult_87_CARRYB_26__28_), .CI(u5_mult_87_SUMB_26__29_), .CO(
        u5_mult_87_CARRYB_27__28_), .S(u5_mult_87_SUMB_27__28_) );
  FA_X1 u5_mult_87_S2_27_27 ( .A(u5_mult_87_ab_27__27_), .B(
        u5_mult_87_CARRYB_26__27_), .CI(u5_mult_87_SUMB_26__28_), .CO(
        u5_mult_87_CARRYB_27__27_), .S(u5_mult_87_SUMB_27__27_) );
  FA_X1 u5_mult_87_S2_27_26 ( .A(u5_mult_87_ab_27__26_), .B(
        u5_mult_87_CARRYB_26__26_), .CI(u5_mult_87_SUMB_26__27_), .CO(
        u5_mult_87_CARRYB_27__26_), .S(u5_mult_87_SUMB_27__26_) );
  FA_X1 u5_mult_87_S2_27_25 ( .A(u5_mult_87_ab_27__25_), .B(
        u5_mult_87_CARRYB_26__25_), .CI(u5_mult_87_SUMB_26__26_), .CO(
        u5_mult_87_CARRYB_27__25_), .S(u5_mult_87_SUMB_27__25_) );
  FA_X1 u5_mult_87_S2_27_24 ( .A(u5_mult_87_ab_27__24_), .B(
        u5_mult_87_CARRYB_26__24_), .CI(u5_mult_87_SUMB_26__25_), .CO(
        u5_mult_87_CARRYB_27__24_), .S(u5_mult_87_SUMB_27__24_) );
  FA_X1 u5_mult_87_S2_27_23 ( .A(u5_mult_87_ab_27__23_), .B(
        u5_mult_87_CARRYB_26__23_), .CI(u5_mult_87_SUMB_26__24_), .CO(
        u5_mult_87_CARRYB_27__23_), .S(u5_mult_87_SUMB_27__23_) );
  FA_X1 u5_mult_87_S2_27_22 ( .A(u5_mult_87_ab_27__22_), .B(
        u5_mult_87_CARRYB_26__22_), .CI(u5_mult_87_SUMB_26__23_), .CO(
        u5_mult_87_CARRYB_27__22_), .S(u5_mult_87_SUMB_27__22_) );
  FA_X1 u5_mult_87_S2_27_21 ( .A(u5_mult_87_ab_27__21_), .B(
        u5_mult_87_CARRYB_26__21_), .CI(u5_mult_87_SUMB_26__22_), .CO(
        u5_mult_87_CARRYB_27__21_), .S(u5_mult_87_SUMB_27__21_) );
  FA_X1 u5_mult_87_S2_27_20 ( .A(u5_mult_87_ab_27__20_), .B(
        u5_mult_87_CARRYB_26__20_), .CI(u5_mult_87_SUMB_26__21_), .CO(
        u5_mult_87_CARRYB_27__20_), .S(u5_mult_87_SUMB_27__20_) );
  FA_X1 u5_mult_87_S2_27_19 ( .A(u5_mult_87_ab_27__19_), .B(
        u5_mult_87_CARRYB_26__19_), .CI(u5_mult_87_SUMB_26__20_), .CO(
        u5_mult_87_CARRYB_27__19_), .S(u5_mult_87_SUMB_27__19_) );
  FA_X1 u5_mult_87_S2_27_18 ( .A(u5_mult_87_ab_27__18_), .B(
        u5_mult_87_CARRYB_26__18_), .CI(u5_mult_87_SUMB_26__19_), .CO(
        u5_mult_87_CARRYB_27__18_), .S(u5_mult_87_SUMB_27__18_) );
  FA_X1 u5_mult_87_S2_27_17 ( .A(u5_mult_87_ab_27__17_), .B(
        u5_mult_87_CARRYB_26__17_), .CI(u5_mult_87_SUMB_26__18_), .CO(
        u5_mult_87_CARRYB_27__17_), .S(u5_mult_87_SUMB_27__17_) );
  FA_X1 u5_mult_87_S2_27_16 ( .A(u5_mult_87_ab_27__16_), .B(
        u5_mult_87_CARRYB_26__16_), .CI(u5_mult_87_SUMB_26__17_), .CO(
        u5_mult_87_CARRYB_27__16_), .S(u5_mult_87_SUMB_27__16_) );
  FA_X1 u5_mult_87_S2_27_15 ( .A(u5_mult_87_ab_27__15_), .B(
        u5_mult_87_CARRYB_26__15_), .CI(u5_mult_87_SUMB_26__16_), .CO(
        u5_mult_87_CARRYB_27__15_), .S(u5_mult_87_SUMB_27__15_) );
  FA_X1 u5_mult_87_S2_27_14 ( .A(u5_mult_87_ab_27__14_), .B(
        u5_mult_87_CARRYB_26__14_), .CI(u5_mult_87_SUMB_26__15_), .CO(
        u5_mult_87_CARRYB_27__14_), .S(u5_mult_87_SUMB_27__14_) );
  FA_X1 u5_mult_87_S2_27_13 ( .A(u5_mult_87_ab_27__13_), .B(
        u5_mult_87_CARRYB_26__13_), .CI(u5_mult_87_SUMB_26__14_), .CO(
        u5_mult_87_CARRYB_27__13_), .S(u5_mult_87_SUMB_27__13_) );
  FA_X1 u5_mult_87_S2_27_12 ( .A(u5_mult_87_ab_27__12_), .B(
        u5_mult_87_CARRYB_26__12_), .CI(u5_mult_87_SUMB_26__13_), .CO(
        u5_mult_87_CARRYB_27__12_), .S(u5_mult_87_SUMB_27__12_) );
  FA_X1 u5_mult_87_S2_27_11 ( .A(u5_mult_87_ab_27__11_), .B(
        u5_mult_87_CARRYB_26__11_), .CI(u5_mult_87_SUMB_26__12_), .CO(
        u5_mult_87_CARRYB_27__11_), .S(u5_mult_87_SUMB_27__11_) );
  FA_X1 u5_mult_87_S2_27_10 ( .A(u5_mult_87_ab_27__10_), .B(
        u5_mult_87_CARRYB_26__10_), .CI(u5_mult_87_SUMB_26__11_), .CO(
        u5_mult_87_CARRYB_27__10_), .S(u5_mult_87_SUMB_27__10_) );
  FA_X1 u5_mult_87_S2_27_9 ( .A(u5_mult_87_ab_27__9_), .B(
        u5_mult_87_CARRYB_26__9_), .CI(u5_mult_87_SUMB_26__10_), .CO(
        u5_mult_87_CARRYB_27__9_), .S(u5_mult_87_SUMB_27__9_) );
  FA_X1 u5_mult_87_S2_27_8 ( .A(u5_mult_87_ab_27__8_), .B(
        u5_mult_87_CARRYB_26__8_), .CI(u5_mult_87_SUMB_26__9_), .CO(
        u5_mult_87_CARRYB_27__8_), .S(u5_mult_87_SUMB_27__8_) );
  FA_X1 u5_mult_87_S2_27_7 ( .A(u5_mult_87_ab_27__7_), .B(
        u5_mult_87_CARRYB_26__7_), .CI(u5_mult_87_SUMB_26__8_), .CO(
        u5_mult_87_CARRYB_27__7_), .S(u5_mult_87_SUMB_27__7_) );
  FA_X1 u5_mult_87_S2_27_6 ( .A(u5_mult_87_ab_27__6_), .B(
        u5_mult_87_CARRYB_26__6_), .CI(u5_mult_87_SUMB_26__7_), .CO(
        u5_mult_87_CARRYB_27__6_), .S(u5_mult_87_SUMB_27__6_) );
  FA_X1 u5_mult_87_S2_27_5 ( .A(u5_mult_87_ab_27__5_), .B(
        u5_mult_87_CARRYB_26__5_), .CI(u5_mult_87_SUMB_26__6_), .CO(
        u5_mult_87_CARRYB_27__5_), .S(u5_mult_87_SUMB_27__5_) );
  FA_X1 u5_mult_87_S2_27_4 ( .A(u5_mult_87_ab_27__4_), .B(
        u5_mult_87_CARRYB_26__4_), .CI(u5_mult_87_SUMB_26__5_), .CO(
        u5_mult_87_CARRYB_27__4_), .S(u5_mult_87_SUMB_27__4_) );
  FA_X1 u5_mult_87_S2_27_3 ( .A(u5_mult_87_ab_27__3_), .B(
        u5_mult_87_CARRYB_26__3_), .CI(u5_mult_87_SUMB_26__4_), .CO(
        u5_mult_87_CARRYB_27__3_), .S(u5_mult_87_SUMB_27__3_) );
  FA_X1 u5_mult_87_S2_27_2 ( .A(u5_mult_87_ab_27__2_), .B(
        u5_mult_87_CARRYB_26__2_), .CI(u5_mult_87_SUMB_26__3_), .CO(
        u5_mult_87_CARRYB_27__2_), .S(u5_mult_87_SUMB_27__2_) );
  FA_X1 u5_mult_87_S2_27_1 ( .A(u5_mult_87_ab_27__1_), .B(
        u5_mult_87_CARRYB_26__1_), .CI(u5_mult_87_SUMB_26__2_), .CO(
        u5_mult_87_CARRYB_27__1_), .S(u5_mult_87_SUMB_27__1_) );
  FA_X1 u5_mult_87_S1_27_0 ( .A(u5_mult_87_ab_27__0_), .B(
        u5_mult_87_CARRYB_26__0_), .CI(u5_mult_87_SUMB_26__1_), .CO(
        u5_mult_87_CARRYB_27__0_), .S(u5_N27) );
  FA_X1 u5_mult_87_S3_28_51 ( .A(u5_mult_87_ab_28__51_), .B(
        u5_mult_87_CARRYB_27__51_), .CI(u5_mult_87_ab_27__52_), .CO(
        u5_mult_87_CARRYB_28__51_), .S(u5_mult_87_SUMB_28__51_) );
  FA_X1 u5_mult_87_S2_28_50 ( .A(u5_mult_87_ab_28__50_), .B(
        u5_mult_87_CARRYB_27__50_), .CI(u5_mult_87_SUMB_27__51_), .CO(
        u5_mult_87_CARRYB_28__50_), .S(u5_mult_87_SUMB_28__50_) );
  FA_X1 u5_mult_87_S2_28_49 ( .A(u5_mult_87_ab_28__49_), .B(
        u5_mult_87_CARRYB_27__49_), .CI(u5_mult_87_SUMB_27__50_), .CO(
        u5_mult_87_CARRYB_28__49_), .S(u5_mult_87_SUMB_28__49_) );
  FA_X1 u5_mult_87_S2_28_48 ( .A(u5_mult_87_ab_28__48_), .B(
        u5_mult_87_CARRYB_27__48_), .CI(u5_mult_87_SUMB_27__49_), .CO(
        u5_mult_87_CARRYB_28__48_), .S(u5_mult_87_SUMB_28__48_) );
  FA_X1 u5_mult_87_S2_28_47 ( .A(u5_mult_87_ab_28__47_), .B(
        u5_mult_87_CARRYB_27__47_), .CI(u5_mult_87_SUMB_27__48_), .CO(
        u5_mult_87_CARRYB_28__47_), .S(u5_mult_87_SUMB_28__47_) );
  FA_X1 u5_mult_87_S2_28_46 ( .A(u5_mult_87_ab_28__46_), .B(
        u5_mult_87_CARRYB_27__46_), .CI(u5_mult_87_SUMB_27__47_), .CO(
        u5_mult_87_CARRYB_28__46_), .S(u5_mult_87_SUMB_28__46_) );
  FA_X1 u5_mult_87_S2_28_45 ( .A(u5_mult_87_ab_28__45_), .B(
        u5_mult_87_CARRYB_27__45_), .CI(u5_mult_87_SUMB_27__46_), .CO(
        u5_mult_87_CARRYB_28__45_), .S(u5_mult_87_SUMB_28__45_) );
  FA_X1 u5_mult_87_S2_28_44 ( .A(u5_mult_87_ab_28__44_), .B(
        u5_mult_87_CARRYB_27__44_), .CI(u5_mult_87_SUMB_27__45_), .CO(
        u5_mult_87_CARRYB_28__44_), .S(u5_mult_87_SUMB_28__44_) );
  FA_X1 u5_mult_87_S2_28_43 ( .A(u5_mult_87_ab_28__43_), .B(
        u5_mult_87_CARRYB_27__43_), .CI(u5_mult_87_SUMB_27__44_), .CO(
        u5_mult_87_CARRYB_28__43_), .S(u5_mult_87_SUMB_28__43_) );
  FA_X1 u5_mult_87_S2_28_42 ( .A(u5_mult_87_ab_28__42_), .B(
        u5_mult_87_CARRYB_27__42_), .CI(u5_mult_87_SUMB_27__43_), .CO(
        u5_mult_87_CARRYB_28__42_), .S(u5_mult_87_SUMB_28__42_) );
  FA_X1 u5_mult_87_S2_28_41 ( .A(u5_mult_87_ab_28__41_), .B(
        u5_mult_87_CARRYB_27__41_), .CI(u5_mult_87_SUMB_27__42_), .CO(
        u5_mult_87_CARRYB_28__41_), .S(u5_mult_87_SUMB_28__41_) );
  FA_X1 u5_mult_87_S2_28_40 ( .A(u5_mult_87_ab_28__40_), .B(
        u5_mult_87_CARRYB_27__40_), .CI(u5_mult_87_SUMB_27__41_), .CO(
        u5_mult_87_CARRYB_28__40_), .S(u5_mult_87_SUMB_28__40_) );
  FA_X1 u5_mult_87_S2_28_39 ( .A(u5_mult_87_ab_28__39_), .B(
        u5_mult_87_CARRYB_27__39_), .CI(u5_mult_87_SUMB_27__40_), .CO(
        u5_mult_87_CARRYB_28__39_), .S(u5_mult_87_SUMB_28__39_) );
  FA_X1 u5_mult_87_S2_28_38 ( .A(u5_mult_87_ab_28__38_), .B(
        u5_mult_87_CARRYB_27__38_), .CI(u5_mult_87_SUMB_27__39_), .CO(
        u5_mult_87_CARRYB_28__38_), .S(u5_mult_87_SUMB_28__38_) );
  FA_X1 u5_mult_87_S2_28_37 ( .A(u5_mult_87_ab_28__37_), .B(
        u5_mult_87_CARRYB_27__37_), .CI(u5_mult_87_SUMB_27__38_), .CO(
        u5_mult_87_CARRYB_28__37_), .S(u5_mult_87_SUMB_28__37_) );
  FA_X1 u5_mult_87_S2_28_36 ( .A(u5_mult_87_ab_28__36_), .B(
        u5_mult_87_CARRYB_27__36_), .CI(u5_mult_87_SUMB_27__37_), .CO(
        u5_mult_87_CARRYB_28__36_), .S(u5_mult_87_SUMB_28__36_) );
  FA_X1 u5_mult_87_S2_28_35 ( .A(u5_mult_87_ab_28__35_), .B(
        u5_mult_87_CARRYB_27__35_), .CI(u5_mult_87_SUMB_27__36_), .CO(
        u5_mult_87_CARRYB_28__35_), .S(u5_mult_87_SUMB_28__35_) );
  FA_X1 u5_mult_87_S2_28_34 ( .A(u5_mult_87_ab_28__34_), .B(
        u5_mult_87_CARRYB_27__34_), .CI(u5_mult_87_SUMB_27__35_), .CO(
        u5_mult_87_CARRYB_28__34_), .S(u5_mult_87_SUMB_28__34_) );
  FA_X1 u5_mult_87_S2_28_33 ( .A(u5_mult_87_ab_28__33_), .B(
        u5_mult_87_CARRYB_27__33_), .CI(u5_mult_87_SUMB_27__34_), .CO(
        u5_mult_87_CARRYB_28__33_), .S(u5_mult_87_SUMB_28__33_) );
  FA_X1 u5_mult_87_S2_28_32 ( .A(u5_mult_87_ab_28__32_), .B(
        u5_mult_87_CARRYB_27__32_), .CI(u5_mult_87_SUMB_27__33_), .CO(
        u5_mult_87_CARRYB_28__32_), .S(u5_mult_87_SUMB_28__32_) );
  FA_X1 u5_mult_87_S2_28_31 ( .A(u5_mult_87_ab_28__31_), .B(
        u5_mult_87_CARRYB_27__31_), .CI(u5_mult_87_SUMB_27__32_), .CO(
        u5_mult_87_CARRYB_28__31_), .S(u5_mult_87_SUMB_28__31_) );
  FA_X1 u5_mult_87_S2_28_30 ( .A(u5_mult_87_ab_28__30_), .B(
        u5_mult_87_CARRYB_27__30_), .CI(u5_mult_87_SUMB_27__31_), .CO(
        u5_mult_87_CARRYB_28__30_), .S(u5_mult_87_SUMB_28__30_) );
  FA_X1 u5_mult_87_S2_28_29 ( .A(u5_mult_87_ab_28__29_), .B(
        u5_mult_87_CARRYB_27__29_), .CI(u5_mult_87_SUMB_27__30_), .CO(
        u5_mult_87_CARRYB_28__29_), .S(u5_mult_87_SUMB_28__29_) );
  FA_X1 u5_mult_87_S2_28_28 ( .A(u5_mult_87_ab_28__28_), .B(
        u5_mult_87_CARRYB_27__28_), .CI(u5_mult_87_SUMB_27__29_), .CO(
        u5_mult_87_CARRYB_28__28_), .S(u5_mult_87_SUMB_28__28_) );
  FA_X1 u5_mult_87_S2_28_27 ( .A(u5_mult_87_ab_28__27_), .B(
        u5_mult_87_CARRYB_27__27_), .CI(u5_mult_87_SUMB_27__28_), .CO(
        u5_mult_87_CARRYB_28__27_), .S(u5_mult_87_SUMB_28__27_) );
  FA_X1 u5_mult_87_S2_28_26 ( .A(u5_mult_87_ab_28__26_), .B(
        u5_mult_87_CARRYB_27__26_), .CI(u5_mult_87_SUMB_27__27_), .CO(
        u5_mult_87_CARRYB_28__26_), .S(u5_mult_87_SUMB_28__26_) );
  FA_X1 u5_mult_87_S2_28_25 ( .A(u5_mult_87_ab_28__25_), .B(
        u5_mult_87_CARRYB_27__25_), .CI(u5_mult_87_SUMB_27__26_), .CO(
        u5_mult_87_CARRYB_28__25_), .S(u5_mult_87_SUMB_28__25_) );
  FA_X1 u5_mult_87_S2_28_24 ( .A(u5_mult_87_ab_28__24_), .B(
        u5_mult_87_CARRYB_27__24_), .CI(u5_mult_87_SUMB_27__25_), .CO(
        u5_mult_87_CARRYB_28__24_), .S(u5_mult_87_SUMB_28__24_) );
  FA_X1 u5_mult_87_S2_28_23 ( .A(u5_mult_87_ab_28__23_), .B(
        u5_mult_87_CARRYB_27__23_), .CI(u5_mult_87_SUMB_27__24_), .CO(
        u5_mult_87_CARRYB_28__23_), .S(u5_mult_87_SUMB_28__23_) );
  FA_X1 u5_mult_87_S2_28_22 ( .A(u5_mult_87_ab_28__22_), .B(
        u5_mult_87_CARRYB_27__22_), .CI(u5_mult_87_SUMB_27__23_), .CO(
        u5_mult_87_CARRYB_28__22_), .S(u5_mult_87_SUMB_28__22_) );
  FA_X1 u5_mult_87_S2_28_21 ( .A(u5_mult_87_ab_28__21_), .B(
        u5_mult_87_CARRYB_27__21_), .CI(u5_mult_87_SUMB_27__22_), .CO(
        u5_mult_87_CARRYB_28__21_), .S(u5_mult_87_SUMB_28__21_) );
  FA_X1 u5_mult_87_S2_28_20 ( .A(u5_mult_87_ab_28__20_), .B(
        u5_mult_87_CARRYB_27__20_), .CI(u5_mult_87_SUMB_27__21_), .CO(
        u5_mult_87_CARRYB_28__20_), .S(u5_mult_87_SUMB_28__20_) );
  FA_X1 u5_mult_87_S2_28_19 ( .A(u5_mult_87_ab_28__19_), .B(
        u5_mult_87_CARRYB_27__19_), .CI(u5_mult_87_SUMB_27__20_), .CO(
        u5_mult_87_CARRYB_28__19_), .S(u5_mult_87_SUMB_28__19_) );
  FA_X1 u5_mult_87_S2_28_18 ( .A(u5_mult_87_ab_28__18_), .B(
        u5_mult_87_CARRYB_27__18_), .CI(u5_mult_87_SUMB_27__19_), .CO(
        u5_mult_87_CARRYB_28__18_), .S(u5_mult_87_SUMB_28__18_) );
  FA_X1 u5_mult_87_S2_28_17 ( .A(u5_mult_87_ab_28__17_), .B(
        u5_mult_87_CARRYB_27__17_), .CI(u5_mult_87_SUMB_27__18_), .CO(
        u5_mult_87_CARRYB_28__17_), .S(u5_mult_87_SUMB_28__17_) );
  FA_X1 u5_mult_87_S2_28_16 ( .A(u5_mult_87_ab_28__16_), .B(
        u5_mult_87_CARRYB_27__16_), .CI(u5_mult_87_SUMB_27__17_), .CO(
        u5_mult_87_CARRYB_28__16_), .S(u5_mult_87_SUMB_28__16_) );
  FA_X1 u5_mult_87_S2_28_15 ( .A(u5_mult_87_ab_28__15_), .B(
        u5_mult_87_CARRYB_27__15_), .CI(u5_mult_87_SUMB_27__16_), .CO(
        u5_mult_87_CARRYB_28__15_), .S(u5_mult_87_SUMB_28__15_) );
  FA_X1 u5_mult_87_S2_28_14 ( .A(u5_mult_87_ab_28__14_), .B(
        u5_mult_87_CARRYB_27__14_), .CI(u5_mult_87_SUMB_27__15_), .CO(
        u5_mult_87_CARRYB_28__14_), .S(u5_mult_87_SUMB_28__14_) );
  FA_X1 u5_mult_87_S2_28_13 ( .A(u5_mult_87_ab_28__13_), .B(
        u5_mult_87_CARRYB_27__13_), .CI(u5_mult_87_SUMB_27__14_), .CO(
        u5_mult_87_CARRYB_28__13_), .S(u5_mult_87_SUMB_28__13_) );
  FA_X1 u5_mult_87_S2_28_12 ( .A(u5_mult_87_ab_28__12_), .B(
        u5_mult_87_CARRYB_27__12_), .CI(u5_mult_87_SUMB_27__13_), .CO(
        u5_mult_87_CARRYB_28__12_), .S(u5_mult_87_SUMB_28__12_) );
  FA_X1 u5_mult_87_S2_28_11 ( .A(u5_mult_87_ab_28__11_), .B(
        u5_mult_87_CARRYB_27__11_), .CI(u5_mult_87_SUMB_27__12_), .CO(
        u5_mult_87_CARRYB_28__11_), .S(u5_mult_87_SUMB_28__11_) );
  FA_X1 u5_mult_87_S2_28_10 ( .A(u5_mult_87_ab_28__10_), .B(
        u5_mult_87_CARRYB_27__10_), .CI(u5_mult_87_SUMB_27__11_), .CO(
        u5_mult_87_CARRYB_28__10_), .S(u5_mult_87_SUMB_28__10_) );
  FA_X1 u5_mult_87_S2_28_9 ( .A(u5_mult_87_ab_28__9_), .B(
        u5_mult_87_CARRYB_27__9_), .CI(u5_mult_87_SUMB_27__10_), .CO(
        u5_mult_87_CARRYB_28__9_), .S(u5_mult_87_SUMB_28__9_) );
  FA_X1 u5_mult_87_S2_28_8 ( .A(u5_mult_87_ab_28__8_), .B(
        u5_mult_87_CARRYB_27__8_), .CI(u5_mult_87_SUMB_27__9_), .CO(
        u5_mult_87_CARRYB_28__8_), .S(u5_mult_87_SUMB_28__8_) );
  FA_X1 u5_mult_87_S2_28_7 ( .A(u5_mult_87_ab_28__7_), .B(
        u5_mult_87_CARRYB_27__7_), .CI(u5_mult_87_SUMB_27__8_), .CO(
        u5_mult_87_CARRYB_28__7_), .S(u5_mult_87_SUMB_28__7_) );
  FA_X1 u5_mult_87_S2_28_6 ( .A(u5_mult_87_ab_28__6_), .B(
        u5_mult_87_CARRYB_27__6_), .CI(u5_mult_87_SUMB_27__7_), .CO(
        u5_mult_87_CARRYB_28__6_), .S(u5_mult_87_SUMB_28__6_) );
  FA_X1 u5_mult_87_S2_28_5 ( .A(u5_mult_87_ab_28__5_), .B(
        u5_mult_87_CARRYB_27__5_), .CI(u5_mult_87_SUMB_27__6_), .CO(
        u5_mult_87_CARRYB_28__5_), .S(u5_mult_87_SUMB_28__5_) );
  FA_X1 u5_mult_87_S2_28_4 ( .A(u5_mult_87_ab_28__4_), .B(
        u5_mult_87_CARRYB_27__4_), .CI(u5_mult_87_SUMB_27__5_), .CO(
        u5_mult_87_CARRYB_28__4_), .S(u5_mult_87_SUMB_28__4_) );
  FA_X1 u5_mult_87_S2_28_3 ( .A(u5_mult_87_ab_28__3_), .B(
        u5_mult_87_CARRYB_27__3_), .CI(u5_mult_87_SUMB_27__4_), .CO(
        u5_mult_87_CARRYB_28__3_), .S(u5_mult_87_SUMB_28__3_) );
  FA_X1 u5_mult_87_S2_28_2 ( .A(u5_mult_87_ab_28__2_), .B(
        u5_mult_87_CARRYB_27__2_), .CI(u5_mult_87_SUMB_27__3_), .CO(
        u5_mult_87_CARRYB_28__2_), .S(u5_mult_87_SUMB_28__2_) );
  FA_X1 u5_mult_87_S2_28_1 ( .A(u5_mult_87_ab_28__1_), .B(
        u5_mult_87_CARRYB_27__1_), .CI(u5_mult_87_SUMB_27__2_), .CO(
        u5_mult_87_CARRYB_28__1_), .S(u5_mult_87_SUMB_28__1_) );
  FA_X1 u5_mult_87_S1_28_0 ( .A(u5_mult_87_ab_28__0_), .B(
        u5_mult_87_CARRYB_27__0_), .CI(u5_mult_87_SUMB_27__1_), .CO(
        u5_mult_87_CARRYB_28__0_), .S(u5_N28) );
  FA_X1 u5_mult_87_S3_29_51 ( .A(u5_mult_87_ab_29__51_), .B(
        u5_mult_87_CARRYB_28__51_), .CI(u5_mult_87_ab_28__52_), .CO(
        u5_mult_87_CARRYB_29__51_), .S(u5_mult_87_SUMB_29__51_) );
  FA_X1 u5_mult_87_S2_29_50 ( .A(u5_mult_87_ab_29__50_), .B(
        u5_mult_87_CARRYB_28__50_), .CI(u5_mult_87_SUMB_28__51_), .CO(
        u5_mult_87_CARRYB_29__50_), .S(u5_mult_87_SUMB_29__50_) );
  FA_X1 u5_mult_87_S2_29_49 ( .A(u5_mult_87_ab_29__49_), .B(
        u5_mult_87_CARRYB_28__49_), .CI(u5_mult_87_SUMB_28__50_), .CO(
        u5_mult_87_CARRYB_29__49_), .S(u5_mult_87_SUMB_29__49_) );
  FA_X1 u5_mult_87_S2_29_48 ( .A(u5_mult_87_ab_29__48_), .B(
        u5_mult_87_CARRYB_28__48_), .CI(u5_mult_87_SUMB_28__49_), .CO(
        u5_mult_87_CARRYB_29__48_), .S(u5_mult_87_SUMB_29__48_) );
  FA_X1 u5_mult_87_S2_29_47 ( .A(u5_mult_87_ab_29__47_), .B(
        u5_mult_87_CARRYB_28__47_), .CI(u5_mult_87_SUMB_28__48_), .CO(
        u5_mult_87_CARRYB_29__47_), .S(u5_mult_87_SUMB_29__47_) );
  FA_X1 u5_mult_87_S2_29_46 ( .A(u5_mult_87_ab_29__46_), .B(
        u5_mult_87_CARRYB_28__46_), .CI(u5_mult_87_SUMB_28__47_), .CO(
        u5_mult_87_CARRYB_29__46_), .S(u5_mult_87_SUMB_29__46_) );
  FA_X1 u5_mult_87_S2_29_45 ( .A(u5_mult_87_ab_29__45_), .B(
        u5_mult_87_CARRYB_28__45_), .CI(u5_mult_87_SUMB_28__46_), .CO(
        u5_mult_87_CARRYB_29__45_), .S(u5_mult_87_SUMB_29__45_) );
  FA_X1 u5_mult_87_S2_29_44 ( .A(u5_mult_87_ab_29__44_), .B(
        u5_mult_87_CARRYB_28__44_), .CI(u5_mult_87_SUMB_28__45_), .CO(
        u5_mult_87_CARRYB_29__44_), .S(u5_mult_87_SUMB_29__44_) );
  FA_X1 u5_mult_87_S2_29_43 ( .A(u5_mult_87_ab_29__43_), .B(
        u5_mult_87_CARRYB_28__43_), .CI(u5_mult_87_SUMB_28__44_), .CO(
        u5_mult_87_CARRYB_29__43_), .S(u5_mult_87_SUMB_29__43_) );
  FA_X1 u5_mult_87_S2_29_42 ( .A(u5_mult_87_ab_29__42_), .B(
        u5_mult_87_CARRYB_28__42_), .CI(u5_mult_87_SUMB_28__43_), .CO(
        u5_mult_87_CARRYB_29__42_), .S(u5_mult_87_SUMB_29__42_) );
  FA_X1 u5_mult_87_S2_29_41 ( .A(u5_mult_87_ab_29__41_), .B(
        u5_mult_87_CARRYB_28__41_), .CI(u5_mult_87_SUMB_28__42_), .CO(
        u5_mult_87_CARRYB_29__41_), .S(u5_mult_87_SUMB_29__41_) );
  FA_X1 u5_mult_87_S2_29_40 ( .A(u5_mult_87_ab_29__40_), .B(
        u5_mult_87_CARRYB_28__40_), .CI(u5_mult_87_SUMB_28__41_), .CO(
        u5_mult_87_CARRYB_29__40_), .S(u5_mult_87_SUMB_29__40_) );
  FA_X1 u5_mult_87_S2_29_39 ( .A(u5_mult_87_ab_29__39_), .B(
        u5_mult_87_CARRYB_28__39_), .CI(u5_mult_87_SUMB_28__40_), .CO(
        u5_mult_87_CARRYB_29__39_), .S(u5_mult_87_SUMB_29__39_) );
  FA_X1 u5_mult_87_S2_29_38 ( .A(u5_mult_87_ab_29__38_), .B(
        u5_mult_87_CARRYB_28__38_), .CI(u5_mult_87_SUMB_28__39_), .CO(
        u5_mult_87_CARRYB_29__38_), .S(u5_mult_87_SUMB_29__38_) );
  FA_X1 u5_mult_87_S2_29_37 ( .A(u5_mult_87_ab_29__37_), .B(
        u5_mult_87_CARRYB_28__37_), .CI(u5_mult_87_SUMB_28__38_), .CO(
        u5_mult_87_CARRYB_29__37_), .S(u5_mult_87_SUMB_29__37_) );
  FA_X1 u5_mult_87_S2_29_36 ( .A(u5_mult_87_ab_29__36_), .B(
        u5_mult_87_CARRYB_28__36_), .CI(u5_mult_87_SUMB_28__37_), .CO(
        u5_mult_87_CARRYB_29__36_), .S(u5_mult_87_SUMB_29__36_) );
  FA_X1 u5_mult_87_S2_29_35 ( .A(u5_mult_87_ab_29__35_), .B(
        u5_mult_87_CARRYB_28__35_), .CI(u5_mult_87_SUMB_28__36_), .CO(
        u5_mult_87_CARRYB_29__35_), .S(u5_mult_87_SUMB_29__35_) );
  FA_X1 u5_mult_87_S2_29_34 ( .A(u5_mult_87_ab_29__34_), .B(
        u5_mult_87_CARRYB_28__34_), .CI(u5_mult_87_SUMB_28__35_), .CO(
        u5_mult_87_CARRYB_29__34_), .S(u5_mult_87_SUMB_29__34_) );
  FA_X1 u5_mult_87_S2_29_33 ( .A(u5_mult_87_ab_29__33_), .B(
        u5_mult_87_CARRYB_28__33_), .CI(u5_mult_87_SUMB_28__34_), .CO(
        u5_mult_87_CARRYB_29__33_), .S(u5_mult_87_SUMB_29__33_) );
  FA_X1 u5_mult_87_S2_29_32 ( .A(u5_mult_87_ab_29__32_), .B(
        u5_mult_87_CARRYB_28__32_), .CI(u5_mult_87_SUMB_28__33_), .CO(
        u5_mult_87_CARRYB_29__32_), .S(u5_mult_87_SUMB_29__32_) );
  FA_X1 u5_mult_87_S2_29_31 ( .A(u5_mult_87_ab_29__31_), .B(
        u5_mult_87_CARRYB_28__31_), .CI(u5_mult_87_SUMB_28__32_), .CO(
        u5_mult_87_CARRYB_29__31_), .S(u5_mult_87_SUMB_29__31_) );
  FA_X1 u5_mult_87_S2_29_30 ( .A(u5_mult_87_ab_29__30_), .B(
        u5_mult_87_CARRYB_28__30_), .CI(u5_mult_87_SUMB_28__31_), .CO(
        u5_mult_87_CARRYB_29__30_), .S(u5_mult_87_SUMB_29__30_) );
  FA_X1 u5_mult_87_S2_29_29 ( .A(u5_mult_87_ab_29__29_), .B(
        u5_mult_87_CARRYB_28__29_), .CI(u5_mult_87_SUMB_28__30_), .CO(
        u5_mult_87_CARRYB_29__29_), .S(u5_mult_87_SUMB_29__29_) );
  FA_X1 u5_mult_87_S2_29_28 ( .A(u5_mult_87_ab_29__28_), .B(
        u5_mult_87_CARRYB_28__28_), .CI(u5_mult_87_SUMB_28__29_), .CO(
        u5_mult_87_CARRYB_29__28_), .S(u5_mult_87_SUMB_29__28_) );
  FA_X1 u5_mult_87_S2_29_27 ( .A(u5_mult_87_ab_29__27_), .B(
        u5_mult_87_CARRYB_28__27_), .CI(u5_mult_87_SUMB_28__28_), .CO(
        u5_mult_87_CARRYB_29__27_), .S(u5_mult_87_SUMB_29__27_) );
  FA_X1 u5_mult_87_S2_29_26 ( .A(u5_mult_87_ab_29__26_), .B(
        u5_mult_87_CARRYB_28__26_), .CI(u5_mult_87_SUMB_28__27_), .CO(
        u5_mult_87_CARRYB_29__26_), .S(u5_mult_87_SUMB_29__26_) );
  FA_X1 u5_mult_87_S2_29_25 ( .A(u5_mult_87_ab_29__25_), .B(
        u5_mult_87_CARRYB_28__25_), .CI(u5_mult_87_SUMB_28__26_), .CO(
        u5_mult_87_CARRYB_29__25_), .S(u5_mult_87_SUMB_29__25_) );
  FA_X1 u5_mult_87_S2_29_24 ( .A(u5_mult_87_ab_29__24_), .B(
        u5_mult_87_CARRYB_28__24_), .CI(u5_mult_87_SUMB_28__25_), .CO(
        u5_mult_87_CARRYB_29__24_), .S(u5_mult_87_SUMB_29__24_) );
  FA_X1 u5_mult_87_S2_29_23 ( .A(u5_mult_87_ab_29__23_), .B(
        u5_mult_87_CARRYB_28__23_), .CI(u5_mult_87_SUMB_28__24_), .CO(
        u5_mult_87_CARRYB_29__23_), .S(u5_mult_87_SUMB_29__23_) );
  FA_X1 u5_mult_87_S2_29_22 ( .A(u5_mult_87_ab_29__22_), .B(
        u5_mult_87_CARRYB_28__22_), .CI(u5_mult_87_SUMB_28__23_), .CO(
        u5_mult_87_CARRYB_29__22_), .S(u5_mult_87_SUMB_29__22_) );
  FA_X1 u5_mult_87_S2_29_21 ( .A(u5_mult_87_ab_29__21_), .B(
        u5_mult_87_CARRYB_28__21_), .CI(u5_mult_87_SUMB_28__22_), .CO(
        u5_mult_87_CARRYB_29__21_), .S(u5_mult_87_SUMB_29__21_) );
  FA_X1 u5_mult_87_S2_29_20 ( .A(u5_mult_87_ab_29__20_), .B(
        u5_mult_87_CARRYB_28__20_), .CI(u5_mult_87_SUMB_28__21_), .CO(
        u5_mult_87_CARRYB_29__20_), .S(u5_mult_87_SUMB_29__20_) );
  FA_X1 u5_mult_87_S2_29_19 ( .A(u5_mult_87_ab_29__19_), .B(
        u5_mult_87_CARRYB_28__19_), .CI(u5_mult_87_SUMB_28__20_), .CO(
        u5_mult_87_CARRYB_29__19_), .S(u5_mult_87_SUMB_29__19_) );
  FA_X1 u5_mult_87_S2_29_18 ( .A(u5_mult_87_ab_29__18_), .B(
        u5_mult_87_CARRYB_28__18_), .CI(u5_mult_87_SUMB_28__19_), .CO(
        u5_mult_87_CARRYB_29__18_), .S(u5_mult_87_SUMB_29__18_) );
  FA_X1 u5_mult_87_S2_29_17 ( .A(u5_mult_87_ab_29__17_), .B(
        u5_mult_87_CARRYB_28__17_), .CI(u5_mult_87_SUMB_28__18_), .CO(
        u5_mult_87_CARRYB_29__17_), .S(u5_mult_87_SUMB_29__17_) );
  FA_X1 u5_mult_87_S2_29_16 ( .A(u5_mult_87_ab_29__16_), .B(
        u5_mult_87_CARRYB_28__16_), .CI(u5_mult_87_SUMB_28__17_), .CO(
        u5_mult_87_CARRYB_29__16_), .S(u5_mult_87_SUMB_29__16_) );
  FA_X1 u5_mult_87_S2_29_15 ( .A(u5_mult_87_ab_29__15_), .B(
        u5_mult_87_CARRYB_28__15_), .CI(u5_mult_87_SUMB_28__16_), .CO(
        u5_mult_87_CARRYB_29__15_), .S(u5_mult_87_SUMB_29__15_) );
  FA_X1 u5_mult_87_S2_29_14 ( .A(u5_mult_87_ab_29__14_), .B(
        u5_mult_87_CARRYB_28__14_), .CI(u5_mult_87_SUMB_28__15_), .CO(
        u5_mult_87_CARRYB_29__14_), .S(u5_mult_87_SUMB_29__14_) );
  FA_X1 u5_mult_87_S2_29_13 ( .A(u5_mult_87_ab_29__13_), .B(
        u5_mult_87_CARRYB_28__13_), .CI(u5_mult_87_SUMB_28__14_), .CO(
        u5_mult_87_CARRYB_29__13_), .S(u5_mult_87_SUMB_29__13_) );
  FA_X1 u5_mult_87_S2_29_12 ( .A(u5_mult_87_ab_29__12_), .B(
        u5_mult_87_CARRYB_28__12_), .CI(u5_mult_87_SUMB_28__13_), .CO(
        u5_mult_87_CARRYB_29__12_), .S(u5_mult_87_SUMB_29__12_) );
  FA_X1 u5_mult_87_S2_29_11 ( .A(u5_mult_87_ab_29__11_), .B(
        u5_mult_87_CARRYB_28__11_), .CI(u5_mult_87_SUMB_28__12_), .CO(
        u5_mult_87_CARRYB_29__11_), .S(u5_mult_87_SUMB_29__11_) );
  FA_X1 u5_mult_87_S2_29_10 ( .A(u5_mult_87_ab_29__10_), .B(
        u5_mult_87_CARRYB_28__10_), .CI(u5_mult_87_SUMB_28__11_), .CO(
        u5_mult_87_CARRYB_29__10_), .S(u5_mult_87_SUMB_29__10_) );
  FA_X1 u5_mult_87_S2_29_9 ( .A(u5_mult_87_ab_29__9_), .B(
        u5_mult_87_CARRYB_28__9_), .CI(u5_mult_87_SUMB_28__10_), .CO(
        u5_mult_87_CARRYB_29__9_), .S(u5_mult_87_SUMB_29__9_) );
  FA_X1 u5_mult_87_S2_29_8 ( .A(u5_mult_87_ab_29__8_), .B(
        u5_mult_87_CARRYB_28__8_), .CI(u5_mult_87_SUMB_28__9_), .CO(
        u5_mult_87_CARRYB_29__8_), .S(u5_mult_87_SUMB_29__8_) );
  FA_X1 u5_mult_87_S2_29_7 ( .A(u5_mult_87_ab_29__7_), .B(
        u5_mult_87_CARRYB_28__7_), .CI(u5_mult_87_SUMB_28__8_), .CO(
        u5_mult_87_CARRYB_29__7_), .S(u5_mult_87_SUMB_29__7_) );
  FA_X1 u5_mult_87_S2_29_6 ( .A(u5_mult_87_ab_29__6_), .B(
        u5_mult_87_CARRYB_28__6_), .CI(u5_mult_87_SUMB_28__7_), .CO(
        u5_mult_87_CARRYB_29__6_), .S(u5_mult_87_SUMB_29__6_) );
  FA_X1 u5_mult_87_S2_29_5 ( .A(u5_mult_87_ab_29__5_), .B(
        u5_mult_87_CARRYB_28__5_), .CI(u5_mult_87_SUMB_28__6_), .CO(
        u5_mult_87_CARRYB_29__5_), .S(u5_mult_87_SUMB_29__5_) );
  FA_X1 u5_mult_87_S2_29_4 ( .A(u5_mult_87_ab_29__4_), .B(
        u5_mult_87_CARRYB_28__4_), .CI(u5_mult_87_SUMB_28__5_), .CO(
        u5_mult_87_CARRYB_29__4_), .S(u5_mult_87_SUMB_29__4_) );
  FA_X1 u5_mult_87_S2_29_3 ( .A(u5_mult_87_ab_29__3_), .B(
        u5_mult_87_CARRYB_28__3_), .CI(u5_mult_87_SUMB_28__4_), .CO(
        u5_mult_87_CARRYB_29__3_), .S(u5_mult_87_SUMB_29__3_) );
  FA_X1 u5_mult_87_S2_29_2 ( .A(u5_mult_87_ab_29__2_), .B(
        u5_mult_87_CARRYB_28__2_), .CI(u5_mult_87_SUMB_28__3_), .CO(
        u5_mult_87_CARRYB_29__2_), .S(u5_mult_87_SUMB_29__2_) );
  FA_X1 u5_mult_87_S2_29_1 ( .A(u5_mult_87_ab_29__1_), .B(
        u5_mult_87_CARRYB_28__1_), .CI(u5_mult_87_SUMB_28__2_), .CO(
        u5_mult_87_CARRYB_29__1_), .S(u5_mult_87_SUMB_29__1_) );
  FA_X1 u5_mult_87_S1_29_0 ( .A(u5_mult_87_ab_29__0_), .B(
        u5_mult_87_CARRYB_28__0_), .CI(u5_mult_87_SUMB_28__1_), .CO(
        u5_mult_87_CARRYB_29__0_), .S(u5_N29) );
  FA_X1 u5_mult_87_S3_30_51 ( .A(u5_mult_87_ab_30__51_), .B(
        u5_mult_87_CARRYB_29__51_), .CI(u5_mult_87_ab_29__52_), .CO(
        u5_mult_87_CARRYB_30__51_), .S(u5_mult_87_SUMB_30__51_) );
  FA_X1 u5_mult_87_S2_30_50 ( .A(u5_mult_87_ab_30__50_), .B(
        u5_mult_87_CARRYB_29__50_), .CI(u5_mult_87_SUMB_29__51_), .CO(
        u5_mult_87_CARRYB_30__50_), .S(u5_mult_87_SUMB_30__50_) );
  FA_X1 u5_mult_87_S2_30_49 ( .A(u5_mult_87_ab_30__49_), .B(
        u5_mult_87_CARRYB_29__49_), .CI(u5_mult_87_SUMB_29__50_), .CO(
        u5_mult_87_CARRYB_30__49_), .S(u5_mult_87_SUMB_30__49_) );
  FA_X1 u5_mult_87_S2_30_48 ( .A(u5_mult_87_ab_30__48_), .B(
        u5_mult_87_CARRYB_29__48_), .CI(u5_mult_87_SUMB_29__49_), .CO(
        u5_mult_87_CARRYB_30__48_), .S(u5_mult_87_SUMB_30__48_) );
  FA_X1 u5_mult_87_S2_30_47 ( .A(u5_mult_87_ab_30__47_), .B(
        u5_mult_87_CARRYB_29__47_), .CI(u5_mult_87_SUMB_29__48_), .CO(
        u5_mult_87_CARRYB_30__47_), .S(u5_mult_87_SUMB_30__47_) );
  FA_X1 u5_mult_87_S2_30_46 ( .A(u5_mult_87_ab_30__46_), .B(
        u5_mult_87_CARRYB_29__46_), .CI(u5_mult_87_SUMB_29__47_), .CO(
        u5_mult_87_CARRYB_30__46_), .S(u5_mult_87_SUMB_30__46_) );
  FA_X1 u5_mult_87_S2_30_45 ( .A(u5_mult_87_ab_30__45_), .B(
        u5_mult_87_CARRYB_29__45_), .CI(u5_mult_87_SUMB_29__46_), .CO(
        u5_mult_87_CARRYB_30__45_), .S(u5_mult_87_SUMB_30__45_) );
  FA_X1 u5_mult_87_S2_30_44 ( .A(u5_mult_87_ab_30__44_), .B(
        u5_mult_87_CARRYB_29__44_), .CI(u5_mult_87_SUMB_29__45_), .CO(
        u5_mult_87_CARRYB_30__44_), .S(u5_mult_87_SUMB_30__44_) );
  FA_X1 u5_mult_87_S2_30_43 ( .A(u5_mult_87_ab_30__43_), .B(
        u5_mult_87_CARRYB_29__43_), .CI(u5_mult_87_SUMB_29__44_), .CO(
        u5_mult_87_CARRYB_30__43_), .S(u5_mult_87_SUMB_30__43_) );
  FA_X1 u5_mult_87_S2_30_42 ( .A(u5_mult_87_ab_30__42_), .B(
        u5_mult_87_CARRYB_29__42_), .CI(u5_mult_87_SUMB_29__43_), .CO(
        u5_mult_87_CARRYB_30__42_), .S(u5_mult_87_SUMB_30__42_) );
  FA_X1 u5_mult_87_S2_30_41 ( .A(u5_mult_87_ab_30__41_), .B(
        u5_mult_87_CARRYB_29__41_), .CI(u5_mult_87_SUMB_29__42_), .CO(
        u5_mult_87_CARRYB_30__41_), .S(u5_mult_87_SUMB_30__41_) );
  FA_X1 u5_mult_87_S2_30_40 ( .A(u5_mult_87_ab_30__40_), .B(
        u5_mult_87_CARRYB_29__40_), .CI(u5_mult_87_SUMB_29__41_), .CO(
        u5_mult_87_CARRYB_30__40_), .S(u5_mult_87_SUMB_30__40_) );
  FA_X1 u5_mult_87_S2_30_39 ( .A(u5_mult_87_ab_30__39_), .B(
        u5_mult_87_CARRYB_29__39_), .CI(u5_mult_87_SUMB_29__40_), .CO(
        u5_mult_87_CARRYB_30__39_), .S(u5_mult_87_SUMB_30__39_) );
  FA_X1 u5_mult_87_S2_30_38 ( .A(u5_mult_87_ab_30__38_), .B(
        u5_mult_87_CARRYB_29__38_), .CI(u5_mult_87_SUMB_29__39_), .CO(
        u5_mult_87_CARRYB_30__38_), .S(u5_mult_87_SUMB_30__38_) );
  FA_X1 u5_mult_87_S2_30_37 ( .A(u5_mult_87_ab_30__37_), .B(
        u5_mult_87_CARRYB_29__37_), .CI(u5_mult_87_SUMB_29__38_), .CO(
        u5_mult_87_CARRYB_30__37_), .S(u5_mult_87_SUMB_30__37_) );
  FA_X1 u5_mult_87_S2_30_36 ( .A(u5_mult_87_ab_30__36_), .B(
        u5_mult_87_CARRYB_29__36_), .CI(u5_mult_87_SUMB_29__37_), .CO(
        u5_mult_87_CARRYB_30__36_), .S(u5_mult_87_SUMB_30__36_) );
  FA_X1 u5_mult_87_S2_30_35 ( .A(u5_mult_87_ab_30__35_), .B(
        u5_mult_87_CARRYB_29__35_), .CI(u5_mult_87_SUMB_29__36_), .CO(
        u5_mult_87_CARRYB_30__35_), .S(u5_mult_87_SUMB_30__35_) );
  FA_X1 u5_mult_87_S2_30_34 ( .A(u5_mult_87_ab_30__34_), .B(
        u5_mult_87_CARRYB_29__34_), .CI(u5_mult_87_SUMB_29__35_), .CO(
        u5_mult_87_CARRYB_30__34_), .S(u5_mult_87_SUMB_30__34_) );
  FA_X1 u5_mult_87_S2_30_33 ( .A(u5_mult_87_ab_30__33_), .B(
        u5_mult_87_CARRYB_29__33_), .CI(u5_mult_87_SUMB_29__34_), .CO(
        u5_mult_87_CARRYB_30__33_), .S(u5_mult_87_SUMB_30__33_) );
  FA_X1 u5_mult_87_S2_30_32 ( .A(u5_mult_87_ab_30__32_), .B(
        u5_mult_87_CARRYB_29__32_), .CI(u5_mult_87_SUMB_29__33_), .CO(
        u5_mult_87_CARRYB_30__32_), .S(u5_mult_87_SUMB_30__32_) );
  FA_X1 u5_mult_87_S2_30_31 ( .A(u5_mult_87_ab_30__31_), .B(
        u5_mult_87_CARRYB_29__31_), .CI(u5_mult_87_SUMB_29__32_), .CO(
        u5_mult_87_CARRYB_30__31_), .S(u5_mult_87_SUMB_30__31_) );
  FA_X1 u5_mult_87_S2_30_30 ( .A(u5_mult_87_ab_30__30_), .B(
        u5_mult_87_CARRYB_29__30_), .CI(u5_mult_87_SUMB_29__31_), .CO(
        u5_mult_87_CARRYB_30__30_), .S(u5_mult_87_SUMB_30__30_) );
  FA_X1 u5_mult_87_S2_30_29 ( .A(u5_mult_87_ab_30__29_), .B(
        u5_mult_87_CARRYB_29__29_), .CI(u5_mult_87_SUMB_29__30_), .CO(
        u5_mult_87_CARRYB_30__29_), .S(u5_mult_87_SUMB_30__29_) );
  FA_X1 u5_mult_87_S2_30_28 ( .A(u5_mult_87_ab_30__28_), .B(
        u5_mult_87_CARRYB_29__28_), .CI(u5_mult_87_SUMB_29__29_), .CO(
        u5_mult_87_CARRYB_30__28_), .S(u5_mult_87_SUMB_30__28_) );
  FA_X1 u5_mult_87_S2_30_27 ( .A(u5_mult_87_ab_30__27_), .B(
        u5_mult_87_CARRYB_29__27_), .CI(u5_mult_87_SUMB_29__28_), .CO(
        u5_mult_87_CARRYB_30__27_), .S(u5_mult_87_SUMB_30__27_) );
  FA_X1 u5_mult_87_S2_30_26 ( .A(u5_mult_87_ab_30__26_), .B(
        u5_mult_87_CARRYB_29__26_), .CI(u5_mult_87_SUMB_29__27_), .CO(
        u5_mult_87_CARRYB_30__26_), .S(u5_mult_87_SUMB_30__26_) );
  FA_X1 u5_mult_87_S2_30_25 ( .A(u5_mult_87_ab_30__25_), .B(
        u5_mult_87_CARRYB_29__25_), .CI(u5_mult_87_SUMB_29__26_), .CO(
        u5_mult_87_CARRYB_30__25_), .S(u5_mult_87_SUMB_30__25_) );
  FA_X1 u5_mult_87_S2_30_24 ( .A(u5_mult_87_ab_30__24_), .B(
        u5_mult_87_CARRYB_29__24_), .CI(u5_mult_87_SUMB_29__25_), .CO(
        u5_mult_87_CARRYB_30__24_), .S(u5_mult_87_SUMB_30__24_) );
  FA_X1 u5_mult_87_S2_30_23 ( .A(u5_mult_87_ab_30__23_), .B(
        u5_mult_87_CARRYB_29__23_), .CI(u5_mult_87_SUMB_29__24_), .CO(
        u5_mult_87_CARRYB_30__23_), .S(u5_mult_87_SUMB_30__23_) );
  FA_X1 u5_mult_87_S2_30_22 ( .A(u5_mult_87_ab_30__22_), .B(
        u5_mult_87_CARRYB_29__22_), .CI(u5_mult_87_SUMB_29__23_), .CO(
        u5_mult_87_CARRYB_30__22_), .S(u5_mult_87_SUMB_30__22_) );
  FA_X1 u5_mult_87_S2_30_21 ( .A(u5_mult_87_ab_30__21_), .B(
        u5_mult_87_CARRYB_29__21_), .CI(u5_mult_87_SUMB_29__22_), .CO(
        u5_mult_87_CARRYB_30__21_), .S(u5_mult_87_SUMB_30__21_) );
  FA_X1 u5_mult_87_S2_30_20 ( .A(u5_mult_87_ab_30__20_), .B(
        u5_mult_87_CARRYB_29__20_), .CI(u5_mult_87_SUMB_29__21_), .CO(
        u5_mult_87_CARRYB_30__20_), .S(u5_mult_87_SUMB_30__20_) );
  FA_X1 u5_mult_87_S2_30_19 ( .A(u5_mult_87_ab_30__19_), .B(
        u5_mult_87_CARRYB_29__19_), .CI(u5_mult_87_SUMB_29__20_), .CO(
        u5_mult_87_CARRYB_30__19_), .S(u5_mult_87_SUMB_30__19_) );
  FA_X1 u5_mult_87_S2_30_18 ( .A(u5_mult_87_ab_30__18_), .B(
        u5_mult_87_CARRYB_29__18_), .CI(u5_mult_87_SUMB_29__19_), .CO(
        u5_mult_87_CARRYB_30__18_), .S(u5_mult_87_SUMB_30__18_) );
  FA_X1 u5_mult_87_S2_30_17 ( .A(u5_mult_87_ab_30__17_), .B(
        u5_mult_87_CARRYB_29__17_), .CI(u5_mult_87_SUMB_29__18_), .CO(
        u5_mult_87_CARRYB_30__17_), .S(u5_mult_87_SUMB_30__17_) );
  FA_X1 u5_mult_87_S2_30_16 ( .A(u5_mult_87_ab_30__16_), .B(
        u5_mult_87_CARRYB_29__16_), .CI(u5_mult_87_SUMB_29__17_), .CO(
        u5_mult_87_CARRYB_30__16_), .S(u5_mult_87_SUMB_30__16_) );
  FA_X1 u5_mult_87_S2_30_15 ( .A(u5_mult_87_ab_30__15_), .B(
        u5_mult_87_CARRYB_29__15_), .CI(u5_mult_87_SUMB_29__16_), .CO(
        u5_mult_87_CARRYB_30__15_), .S(u5_mult_87_SUMB_30__15_) );
  FA_X1 u5_mult_87_S2_30_14 ( .A(u5_mult_87_ab_30__14_), .B(
        u5_mult_87_CARRYB_29__14_), .CI(u5_mult_87_SUMB_29__15_), .CO(
        u5_mult_87_CARRYB_30__14_), .S(u5_mult_87_SUMB_30__14_) );
  FA_X1 u5_mult_87_S2_30_13 ( .A(u5_mult_87_ab_30__13_), .B(
        u5_mult_87_CARRYB_29__13_), .CI(u5_mult_87_SUMB_29__14_), .CO(
        u5_mult_87_CARRYB_30__13_), .S(u5_mult_87_SUMB_30__13_) );
  FA_X1 u5_mult_87_S2_30_12 ( .A(u5_mult_87_ab_30__12_), .B(
        u5_mult_87_CARRYB_29__12_), .CI(u5_mult_87_SUMB_29__13_), .CO(
        u5_mult_87_CARRYB_30__12_), .S(u5_mult_87_SUMB_30__12_) );
  FA_X1 u5_mult_87_S2_30_11 ( .A(u5_mult_87_ab_30__11_), .B(
        u5_mult_87_CARRYB_29__11_), .CI(u5_mult_87_SUMB_29__12_), .CO(
        u5_mult_87_CARRYB_30__11_), .S(u5_mult_87_SUMB_30__11_) );
  FA_X1 u5_mult_87_S2_30_10 ( .A(u5_mult_87_ab_30__10_), .B(
        u5_mult_87_CARRYB_29__10_), .CI(u5_mult_87_SUMB_29__11_), .CO(
        u5_mult_87_CARRYB_30__10_), .S(u5_mult_87_SUMB_30__10_) );
  FA_X1 u5_mult_87_S2_30_9 ( .A(u5_mult_87_ab_30__9_), .B(
        u5_mult_87_CARRYB_29__9_), .CI(u5_mult_87_SUMB_29__10_), .CO(
        u5_mult_87_CARRYB_30__9_), .S(u5_mult_87_SUMB_30__9_) );
  FA_X1 u5_mult_87_S2_30_8 ( .A(u5_mult_87_ab_30__8_), .B(
        u5_mult_87_CARRYB_29__8_), .CI(u5_mult_87_SUMB_29__9_), .CO(
        u5_mult_87_CARRYB_30__8_), .S(u5_mult_87_SUMB_30__8_) );
  FA_X1 u5_mult_87_S2_30_7 ( .A(u5_mult_87_ab_30__7_), .B(
        u5_mult_87_CARRYB_29__7_), .CI(u5_mult_87_SUMB_29__8_), .CO(
        u5_mult_87_CARRYB_30__7_), .S(u5_mult_87_SUMB_30__7_) );
  FA_X1 u5_mult_87_S2_30_6 ( .A(u5_mult_87_ab_30__6_), .B(
        u5_mult_87_CARRYB_29__6_), .CI(u5_mult_87_SUMB_29__7_), .CO(
        u5_mult_87_CARRYB_30__6_), .S(u5_mult_87_SUMB_30__6_) );
  FA_X1 u5_mult_87_S2_30_5 ( .A(u5_mult_87_ab_30__5_), .B(
        u5_mult_87_CARRYB_29__5_), .CI(u5_mult_87_SUMB_29__6_), .CO(
        u5_mult_87_CARRYB_30__5_), .S(u5_mult_87_SUMB_30__5_) );
  FA_X1 u5_mult_87_S2_30_4 ( .A(u5_mult_87_ab_30__4_), .B(
        u5_mult_87_CARRYB_29__4_), .CI(u5_mult_87_SUMB_29__5_), .CO(
        u5_mult_87_CARRYB_30__4_), .S(u5_mult_87_SUMB_30__4_) );
  FA_X1 u5_mult_87_S2_30_3 ( .A(u5_mult_87_ab_30__3_), .B(
        u5_mult_87_CARRYB_29__3_), .CI(u5_mult_87_SUMB_29__4_), .CO(
        u5_mult_87_CARRYB_30__3_), .S(u5_mult_87_SUMB_30__3_) );
  FA_X1 u5_mult_87_S2_30_2 ( .A(u5_mult_87_ab_30__2_), .B(
        u5_mult_87_CARRYB_29__2_), .CI(u5_mult_87_SUMB_29__3_), .CO(
        u5_mult_87_CARRYB_30__2_), .S(u5_mult_87_SUMB_30__2_) );
  FA_X1 u5_mult_87_S2_30_1 ( .A(u5_mult_87_ab_30__1_), .B(
        u5_mult_87_CARRYB_29__1_), .CI(u5_mult_87_SUMB_29__2_), .CO(
        u5_mult_87_CARRYB_30__1_), .S(u5_mult_87_SUMB_30__1_) );
  FA_X1 u5_mult_87_S1_30_0 ( .A(u5_mult_87_ab_30__0_), .B(
        u5_mult_87_CARRYB_29__0_), .CI(u5_mult_87_SUMB_29__1_), .CO(
        u5_mult_87_CARRYB_30__0_), .S(u5_N30) );
  FA_X1 u5_mult_87_S3_31_51 ( .A(u5_mult_87_ab_31__51_), .B(
        u5_mult_87_CARRYB_30__51_), .CI(u5_mult_87_ab_30__52_), .CO(
        u5_mult_87_CARRYB_31__51_), .S(u5_mult_87_SUMB_31__51_) );
  FA_X1 u5_mult_87_S2_31_50 ( .A(u5_mult_87_ab_31__50_), .B(
        u5_mult_87_CARRYB_30__50_), .CI(u5_mult_87_SUMB_30__51_), .CO(
        u5_mult_87_CARRYB_31__50_), .S(u5_mult_87_SUMB_31__50_) );
  FA_X1 u5_mult_87_S2_31_49 ( .A(u5_mult_87_ab_31__49_), .B(
        u5_mult_87_CARRYB_30__49_), .CI(u5_mult_87_SUMB_30__50_), .CO(
        u5_mult_87_CARRYB_31__49_), .S(u5_mult_87_SUMB_31__49_) );
  FA_X1 u5_mult_87_S2_31_48 ( .A(u5_mult_87_ab_31__48_), .B(
        u5_mult_87_CARRYB_30__48_), .CI(u5_mult_87_SUMB_30__49_), .CO(
        u5_mult_87_CARRYB_31__48_), .S(u5_mult_87_SUMB_31__48_) );
  FA_X1 u5_mult_87_S2_31_47 ( .A(u5_mult_87_ab_31__47_), .B(
        u5_mult_87_CARRYB_30__47_), .CI(u5_mult_87_SUMB_30__48_), .CO(
        u5_mult_87_CARRYB_31__47_), .S(u5_mult_87_SUMB_31__47_) );
  FA_X1 u5_mult_87_S2_31_46 ( .A(u5_mult_87_ab_31__46_), .B(
        u5_mult_87_CARRYB_30__46_), .CI(u5_mult_87_SUMB_30__47_), .CO(
        u5_mult_87_CARRYB_31__46_), .S(u5_mult_87_SUMB_31__46_) );
  FA_X1 u5_mult_87_S2_31_45 ( .A(u5_mult_87_ab_31__45_), .B(
        u5_mult_87_CARRYB_30__45_), .CI(u5_mult_87_SUMB_30__46_), .CO(
        u5_mult_87_CARRYB_31__45_), .S(u5_mult_87_SUMB_31__45_) );
  FA_X1 u5_mult_87_S2_31_44 ( .A(u5_mult_87_ab_31__44_), .B(
        u5_mult_87_CARRYB_30__44_), .CI(u5_mult_87_SUMB_30__45_), .CO(
        u5_mult_87_CARRYB_31__44_), .S(u5_mult_87_SUMB_31__44_) );
  FA_X1 u5_mult_87_S2_31_43 ( .A(u5_mult_87_ab_31__43_), .B(
        u5_mult_87_CARRYB_30__43_), .CI(u5_mult_87_SUMB_30__44_), .CO(
        u5_mult_87_CARRYB_31__43_), .S(u5_mult_87_SUMB_31__43_) );
  FA_X1 u5_mult_87_S2_31_42 ( .A(u5_mult_87_ab_31__42_), .B(
        u5_mult_87_CARRYB_30__42_), .CI(u5_mult_87_SUMB_30__43_), .CO(
        u5_mult_87_CARRYB_31__42_), .S(u5_mult_87_SUMB_31__42_) );
  FA_X1 u5_mult_87_S2_31_41 ( .A(u5_mult_87_ab_31__41_), .B(
        u5_mult_87_CARRYB_30__41_), .CI(u5_mult_87_SUMB_30__42_), .CO(
        u5_mult_87_CARRYB_31__41_), .S(u5_mult_87_SUMB_31__41_) );
  FA_X1 u5_mult_87_S2_31_40 ( .A(u5_mult_87_ab_31__40_), .B(
        u5_mult_87_CARRYB_30__40_), .CI(u5_mult_87_SUMB_30__41_), .CO(
        u5_mult_87_CARRYB_31__40_), .S(u5_mult_87_SUMB_31__40_) );
  FA_X1 u5_mult_87_S2_31_39 ( .A(u5_mult_87_ab_31__39_), .B(
        u5_mult_87_CARRYB_30__39_), .CI(u5_mult_87_SUMB_30__40_), .CO(
        u5_mult_87_CARRYB_31__39_), .S(u5_mult_87_SUMB_31__39_) );
  FA_X1 u5_mult_87_S2_31_38 ( .A(u5_mult_87_ab_31__38_), .B(
        u5_mult_87_CARRYB_30__38_), .CI(u5_mult_87_SUMB_30__39_), .CO(
        u5_mult_87_CARRYB_31__38_), .S(u5_mult_87_SUMB_31__38_) );
  FA_X1 u5_mult_87_S2_31_37 ( .A(u5_mult_87_ab_31__37_), .B(
        u5_mult_87_CARRYB_30__37_), .CI(u5_mult_87_SUMB_30__38_), .CO(
        u5_mult_87_CARRYB_31__37_), .S(u5_mult_87_SUMB_31__37_) );
  FA_X1 u5_mult_87_S2_31_36 ( .A(u5_mult_87_ab_31__36_), .B(
        u5_mult_87_CARRYB_30__36_), .CI(u5_mult_87_SUMB_30__37_), .CO(
        u5_mult_87_CARRYB_31__36_), .S(u5_mult_87_SUMB_31__36_) );
  FA_X1 u5_mult_87_S2_31_35 ( .A(u5_mult_87_ab_31__35_), .B(
        u5_mult_87_CARRYB_30__35_), .CI(u5_mult_87_SUMB_30__36_), .CO(
        u5_mult_87_CARRYB_31__35_), .S(u5_mult_87_SUMB_31__35_) );
  FA_X1 u5_mult_87_S2_31_34 ( .A(u5_mult_87_ab_31__34_), .B(
        u5_mult_87_CARRYB_30__34_), .CI(u5_mult_87_SUMB_30__35_), .CO(
        u5_mult_87_CARRYB_31__34_), .S(u5_mult_87_SUMB_31__34_) );
  FA_X1 u5_mult_87_S2_31_33 ( .A(u5_mult_87_ab_31__33_), .B(
        u5_mult_87_CARRYB_30__33_), .CI(u5_mult_87_SUMB_30__34_), .CO(
        u5_mult_87_CARRYB_31__33_), .S(u5_mult_87_SUMB_31__33_) );
  FA_X1 u5_mult_87_S2_31_32 ( .A(u5_mult_87_ab_31__32_), .B(
        u5_mult_87_CARRYB_30__32_), .CI(u5_mult_87_SUMB_30__33_), .CO(
        u5_mult_87_CARRYB_31__32_), .S(u5_mult_87_SUMB_31__32_) );
  FA_X1 u5_mult_87_S2_31_31 ( .A(u5_mult_87_ab_31__31_), .B(
        u5_mult_87_CARRYB_30__31_), .CI(u5_mult_87_SUMB_30__32_), .CO(
        u5_mult_87_CARRYB_31__31_), .S(u5_mult_87_SUMB_31__31_) );
  FA_X1 u5_mult_87_S2_31_30 ( .A(u5_mult_87_ab_31__30_), .B(
        u5_mult_87_CARRYB_30__30_), .CI(u5_mult_87_SUMB_30__31_), .CO(
        u5_mult_87_CARRYB_31__30_), .S(u5_mult_87_SUMB_31__30_) );
  FA_X1 u5_mult_87_S2_31_29 ( .A(u5_mult_87_ab_31__29_), .B(
        u5_mult_87_CARRYB_30__29_), .CI(u5_mult_87_SUMB_30__30_), .CO(
        u5_mult_87_CARRYB_31__29_), .S(u5_mult_87_SUMB_31__29_) );
  FA_X1 u5_mult_87_S2_31_28 ( .A(u5_mult_87_ab_31__28_), .B(
        u5_mult_87_CARRYB_30__28_), .CI(u5_mult_87_SUMB_30__29_), .CO(
        u5_mult_87_CARRYB_31__28_), .S(u5_mult_87_SUMB_31__28_) );
  FA_X1 u5_mult_87_S2_31_27 ( .A(u5_mult_87_ab_31__27_), .B(
        u5_mult_87_CARRYB_30__27_), .CI(u5_mult_87_SUMB_30__28_), .CO(
        u5_mult_87_CARRYB_31__27_), .S(u5_mult_87_SUMB_31__27_) );
  FA_X1 u5_mult_87_S2_31_26 ( .A(u5_mult_87_ab_31__26_), .B(
        u5_mult_87_CARRYB_30__26_), .CI(u5_mult_87_SUMB_30__27_), .CO(
        u5_mult_87_CARRYB_31__26_), .S(u5_mult_87_SUMB_31__26_) );
  FA_X1 u5_mult_87_S2_31_25 ( .A(u5_mult_87_ab_31__25_), .B(
        u5_mult_87_CARRYB_30__25_), .CI(u5_mult_87_SUMB_30__26_), .CO(
        u5_mult_87_CARRYB_31__25_), .S(u5_mult_87_SUMB_31__25_) );
  FA_X1 u5_mult_87_S2_31_24 ( .A(u5_mult_87_ab_31__24_), .B(
        u5_mult_87_CARRYB_30__24_), .CI(u5_mult_87_SUMB_30__25_), .CO(
        u5_mult_87_CARRYB_31__24_), .S(u5_mult_87_SUMB_31__24_) );
  FA_X1 u5_mult_87_S2_31_23 ( .A(u5_mult_87_ab_31__23_), .B(
        u5_mult_87_CARRYB_30__23_), .CI(u5_mult_87_SUMB_30__24_), .CO(
        u5_mult_87_CARRYB_31__23_), .S(u5_mult_87_SUMB_31__23_) );
  FA_X1 u5_mult_87_S2_31_22 ( .A(u5_mult_87_ab_31__22_), .B(
        u5_mult_87_CARRYB_30__22_), .CI(u5_mult_87_SUMB_30__23_), .CO(
        u5_mult_87_CARRYB_31__22_), .S(u5_mult_87_SUMB_31__22_) );
  FA_X1 u5_mult_87_S2_31_21 ( .A(u5_mult_87_ab_31__21_), .B(
        u5_mult_87_CARRYB_30__21_), .CI(u5_mult_87_SUMB_30__22_), .CO(
        u5_mult_87_CARRYB_31__21_), .S(u5_mult_87_SUMB_31__21_) );
  FA_X1 u5_mult_87_S2_31_20 ( .A(u5_mult_87_ab_31__20_), .B(
        u5_mult_87_CARRYB_30__20_), .CI(u5_mult_87_SUMB_30__21_), .CO(
        u5_mult_87_CARRYB_31__20_), .S(u5_mult_87_SUMB_31__20_) );
  FA_X1 u5_mult_87_S2_31_19 ( .A(u5_mult_87_ab_31__19_), .B(
        u5_mult_87_CARRYB_30__19_), .CI(u5_mult_87_SUMB_30__20_), .CO(
        u5_mult_87_CARRYB_31__19_), .S(u5_mult_87_SUMB_31__19_) );
  FA_X1 u5_mult_87_S2_31_18 ( .A(u5_mult_87_ab_31__18_), .B(
        u5_mult_87_CARRYB_30__18_), .CI(u5_mult_87_SUMB_30__19_), .CO(
        u5_mult_87_CARRYB_31__18_), .S(u5_mult_87_SUMB_31__18_) );
  FA_X1 u5_mult_87_S2_31_17 ( .A(u5_mult_87_ab_31__17_), .B(
        u5_mult_87_CARRYB_30__17_), .CI(u5_mult_87_SUMB_30__18_), .CO(
        u5_mult_87_CARRYB_31__17_), .S(u5_mult_87_SUMB_31__17_) );
  FA_X1 u5_mult_87_S2_31_16 ( .A(u5_mult_87_ab_31__16_), .B(
        u5_mult_87_CARRYB_30__16_), .CI(u5_mult_87_SUMB_30__17_), .CO(
        u5_mult_87_CARRYB_31__16_), .S(u5_mult_87_SUMB_31__16_) );
  FA_X1 u5_mult_87_S2_31_15 ( .A(u5_mult_87_ab_31__15_), .B(
        u5_mult_87_CARRYB_30__15_), .CI(u5_mult_87_SUMB_30__16_), .CO(
        u5_mult_87_CARRYB_31__15_), .S(u5_mult_87_SUMB_31__15_) );
  FA_X1 u5_mult_87_S2_31_14 ( .A(u5_mult_87_ab_31__14_), .B(
        u5_mult_87_CARRYB_30__14_), .CI(u5_mult_87_SUMB_30__15_), .CO(
        u5_mult_87_CARRYB_31__14_), .S(u5_mult_87_SUMB_31__14_) );
  FA_X1 u5_mult_87_S2_31_13 ( .A(u5_mult_87_ab_31__13_), .B(
        u5_mult_87_CARRYB_30__13_), .CI(u5_mult_87_SUMB_30__14_), .CO(
        u5_mult_87_CARRYB_31__13_), .S(u5_mult_87_SUMB_31__13_) );
  FA_X1 u5_mult_87_S2_31_12 ( .A(u5_mult_87_ab_31__12_), .B(
        u5_mult_87_CARRYB_30__12_), .CI(u5_mult_87_SUMB_30__13_), .CO(
        u5_mult_87_CARRYB_31__12_), .S(u5_mult_87_SUMB_31__12_) );
  FA_X1 u5_mult_87_S2_31_11 ( .A(u5_mult_87_ab_31__11_), .B(
        u5_mult_87_CARRYB_30__11_), .CI(u5_mult_87_SUMB_30__12_), .CO(
        u5_mult_87_CARRYB_31__11_), .S(u5_mult_87_SUMB_31__11_) );
  FA_X1 u5_mult_87_S2_31_10 ( .A(u5_mult_87_ab_31__10_), .B(
        u5_mult_87_CARRYB_30__10_), .CI(u5_mult_87_SUMB_30__11_), .CO(
        u5_mult_87_CARRYB_31__10_), .S(u5_mult_87_SUMB_31__10_) );
  FA_X1 u5_mult_87_S2_31_9 ( .A(u5_mult_87_ab_31__9_), .B(
        u5_mult_87_CARRYB_30__9_), .CI(u5_mult_87_SUMB_30__10_), .CO(
        u5_mult_87_CARRYB_31__9_), .S(u5_mult_87_SUMB_31__9_) );
  FA_X1 u5_mult_87_S2_31_8 ( .A(u5_mult_87_ab_31__8_), .B(
        u5_mult_87_CARRYB_30__8_), .CI(u5_mult_87_SUMB_30__9_), .CO(
        u5_mult_87_CARRYB_31__8_), .S(u5_mult_87_SUMB_31__8_) );
  FA_X1 u5_mult_87_S2_31_7 ( .A(u5_mult_87_ab_31__7_), .B(
        u5_mult_87_CARRYB_30__7_), .CI(u5_mult_87_SUMB_30__8_), .CO(
        u5_mult_87_CARRYB_31__7_), .S(u5_mult_87_SUMB_31__7_) );
  FA_X1 u5_mult_87_S2_31_6 ( .A(u5_mult_87_ab_31__6_), .B(
        u5_mult_87_CARRYB_30__6_), .CI(u5_mult_87_SUMB_30__7_), .CO(
        u5_mult_87_CARRYB_31__6_), .S(u5_mult_87_SUMB_31__6_) );
  FA_X1 u5_mult_87_S2_31_5 ( .A(u5_mult_87_ab_31__5_), .B(
        u5_mult_87_CARRYB_30__5_), .CI(u5_mult_87_SUMB_30__6_), .CO(
        u5_mult_87_CARRYB_31__5_), .S(u5_mult_87_SUMB_31__5_) );
  FA_X1 u5_mult_87_S2_31_4 ( .A(u5_mult_87_ab_31__4_), .B(
        u5_mult_87_CARRYB_30__4_), .CI(u5_mult_87_SUMB_30__5_), .CO(
        u5_mult_87_CARRYB_31__4_), .S(u5_mult_87_SUMB_31__4_) );
  FA_X1 u5_mult_87_S2_31_3 ( .A(u5_mult_87_ab_31__3_), .B(
        u5_mult_87_CARRYB_30__3_), .CI(u5_mult_87_SUMB_30__4_), .CO(
        u5_mult_87_CARRYB_31__3_), .S(u5_mult_87_SUMB_31__3_) );
  FA_X1 u5_mult_87_S2_31_2 ( .A(u5_mult_87_ab_31__2_), .B(
        u5_mult_87_CARRYB_30__2_), .CI(u5_mult_87_SUMB_30__3_), .CO(
        u5_mult_87_CARRYB_31__2_), .S(u5_mult_87_SUMB_31__2_) );
  FA_X1 u5_mult_87_S2_31_1 ( .A(u5_mult_87_ab_31__1_), .B(
        u5_mult_87_CARRYB_30__1_), .CI(u5_mult_87_SUMB_30__2_), .CO(
        u5_mult_87_CARRYB_31__1_), .S(u5_mult_87_SUMB_31__1_) );
  FA_X1 u5_mult_87_S1_31_0 ( .A(u5_mult_87_ab_31__0_), .B(
        u5_mult_87_CARRYB_30__0_), .CI(u5_mult_87_SUMB_30__1_), .CO(
        u5_mult_87_CARRYB_31__0_), .S(u5_N31) );
  FA_X1 u5_mult_87_S3_32_51 ( .A(u5_mult_87_ab_32__51_), .B(
        u5_mult_87_CARRYB_31__51_), .CI(u5_mult_87_ab_31__52_), .CO(
        u5_mult_87_CARRYB_32__51_), .S(u5_mult_87_SUMB_32__51_) );
  FA_X1 u5_mult_87_S2_32_50 ( .A(u5_mult_87_ab_32__50_), .B(
        u5_mult_87_CARRYB_31__50_), .CI(u5_mult_87_SUMB_31__51_), .CO(
        u5_mult_87_CARRYB_32__50_), .S(u5_mult_87_SUMB_32__50_) );
  FA_X1 u5_mult_87_S2_32_49 ( .A(u5_mult_87_ab_32__49_), .B(
        u5_mult_87_CARRYB_31__49_), .CI(u5_mult_87_SUMB_31__50_), .CO(
        u5_mult_87_CARRYB_32__49_), .S(u5_mult_87_SUMB_32__49_) );
  FA_X1 u5_mult_87_S2_32_48 ( .A(u5_mult_87_ab_32__48_), .B(
        u5_mult_87_CARRYB_31__48_), .CI(u5_mult_87_SUMB_31__49_), .CO(
        u5_mult_87_CARRYB_32__48_), .S(u5_mult_87_SUMB_32__48_) );
  FA_X1 u5_mult_87_S2_32_47 ( .A(u5_mult_87_ab_32__47_), .B(
        u5_mult_87_CARRYB_31__47_), .CI(u5_mult_87_SUMB_31__48_), .CO(
        u5_mult_87_CARRYB_32__47_), .S(u5_mult_87_SUMB_32__47_) );
  FA_X1 u5_mult_87_S2_32_46 ( .A(u5_mult_87_ab_32__46_), .B(
        u5_mult_87_CARRYB_31__46_), .CI(u5_mult_87_SUMB_31__47_), .CO(
        u5_mult_87_CARRYB_32__46_), .S(u5_mult_87_SUMB_32__46_) );
  FA_X1 u5_mult_87_S2_32_45 ( .A(u5_mult_87_ab_32__45_), .B(
        u5_mult_87_CARRYB_31__45_), .CI(u5_mult_87_SUMB_31__46_), .CO(
        u5_mult_87_CARRYB_32__45_), .S(u5_mult_87_SUMB_32__45_) );
  FA_X1 u5_mult_87_S2_32_44 ( .A(u5_mult_87_ab_32__44_), .B(
        u5_mult_87_CARRYB_31__44_), .CI(u5_mult_87_SUMB_31__45_), .CO(
        u5_mult_87_CARRYB_32__44_), .S(u5_mult_87_SUMB_32__44_) );
  FA_X1 u5_mult_87_S2_32_43 ( .A(u5_mult_87_ab_32__43_), .B(
        u5_mult_87_CARRYB_31__43_), .CI(u5_mult_87_SUMB_31__44_), .CO(
        u5_mult_87_CARRYB_32__43_), .S(u5_mult_87_SUMB_32__43_) );
  FA_X1 u5_mult_87_S2_32_42 ( .A(u5_mult_87_ab_32__42_), .B(
        u5_mult_87_CARRYB_31__42_), .CI(u5_mult_87_SUMB_31__43_), .CO(
        u5_mult_87_CARRYB_32__42_), .S(u5_mult_87_SUMB_32__42_) );
  FA_X1 u5_mult_87_S2_32_41 ( .A(u5_mult_87_ab_32__41_), .B(
        u5_mult_87_CARRYB_31__41_), .CI(u5_mult_87_SUMB_31__42_), .CO(
        u5_mult_87_CARRYB_32__41_), .S(u5_mult_87_SUMB_32__41_) );
  FA_X1 u5_mult_87_S2_32_40 ( .A(u5_mult_87_ab_32__40_), .B(
        u5_mult_87_CARRYB_31__40_), .CI(u5_mult_87_SUMB_31__41_), .CO(
        u5_mult_87_CARRYB_32__40_), .S(u5_mult_87_SUMB_32__40_) );
  FA_X1 u5_mult_87_S2_32_39 ( .A(u5_mult_87_ab_32__39_), .B(
        u5_mult_87_CARRYB_31__39_), .CI(u5_mult_87_SUMB_31__40_), .CO(
        u5_mult_87_CARRYB_32__39_), .S(u5_mult_87_SUMB_32__39_) );
  FA_X1 u5_mult_87_S2_32_38 ( .A(u5_mult_87_ab_32__38_), .B(
        u5_mult_87_CARRYB_31__38_), .CI(u5_mult_87_SUMB_31__39_), .CO(
        u5_mult_87_CARRYB_32__38_), .S(u5_mult_87_SUMB_32__38_) );
  FA_X1 u5_mult_87_S2_32_37 ( .A(u5_mult_87_ab_32__37_), .B(
        u5_mult_87_CARRYB_31__37_), .CI(u5_mult_87_SUMB_31__38_), .CO(
        u5_mult_87_CARRYB_32__37_), .S(u5_mult_87_SUMB_32__37_) );
  FA_X1 u5_mult_87_S2_32_36 ( .A(u5_mult_87_ab_32__36_), .B(
        u5_mult_87_CARRYB_31__36_), .CI(u5_mult_87_SUMB_31__37_), .CO(
        u5_mult_87_CARRYB_32__36_), .S(u5_mult_87_SUMB_32__36_) );
  FA_X1 u5_mult_87_S2_32_35 ( .A(u5_mult_87_ab_32__35_), .B(
        u5_mult_87_CARRYB_31__35_), .CI(u5_mult_87_SUMB_31__36_), .CO(
        u5_mult_87_CARRYB_32__35_), .S(u5_mult_87_SUMB_32__35_) );
  FA_X1 u5_mult_87_S2_32_34 ( .A(u5_mult_87_ab_32__34_), .B(
        u5_mult_87_CARRYB_31__34_), .CI(u5_mult_87_SUMB_31__35_), .CO(
        u5_mult_87_CARRYB_32__34_), .S(u5_mult_87_SUMB_32__34_) );
  FA_X1 u5_mult_87_S2_32_33 ( .A(u5_mult_87_ab_32__33_), .B(
        u5_mult_87_CARRYB_31__33_), .CI(u5_mult_87_SUMB_31__34_), .CO(
        u5_mult_87_CARRYB_32__33_), .S(u5_mult_87_SUMB_32__33_) );
  FA_X1 u5_mult_87_S2_32_32 ( .A(u5_mult_87_ab_32__32_), .B(
        u5_mult_87_CARRYB_31__32_), .CI(u5_mult_87_SUMB_31__33_), .CO(
        u5_mult_87_CARRYB_32__32_), .S(u5_mult_87_SUMB_32__32_) );
  FA_X1 u5_mult_87_S2_32_31 ( .A(u5_mult_87_ab_32__31_), .B(
        u5_mult_87_CARRYB_31__31_), .CI(u5_mult_87_SUMB_31__32_), .CO(
        u5_mult_87_CARRYB_32__31_), .S(u5_mult_87_SUMB_32__31_) );
  FA_X1 u5_mult_87_S2_32_30 ( .A(u5_mult_87_ab_32__30_), .B(
        u5_mult_87_CARRYB_31__30_), .CI(u5_mult_87_SUMB_31__31_), .CO(
        u5_mult_87_CARRYB_32__30_), .S(u5_mult_87_SUMB_32__30_) );
  FA_X1 u5_mult_87_S2_32_29 ( .A(u5_mult_87_ab_32__29_), .B(
        u5_mult_87_CARRYB_31__29_), .CI(u5_mult_87_SUMB_31__30_), .CO(
        u5_mult_87_CARRYB_32__29_), .S(u5_mult_87_SUMB_32__29_) );
  FA_X1 u5_mult_87_S2_32_28 ( .A(u5_mult_87_ab_32__28_), .B(
        u5_mult_87_CARRYB_31__28_), .CI(u5_mult_87_SUMB_31__29_), .CO(
        u5_mult_87_CARRYB_32__28_), .S(u5_mult_87_SUMB_32__28_) );
  FA_X1 u5_mult_87_S2_32_27 ( .A(u5_mult_87_ab_32__27_), .B(
        u5_mult_87_CARRYB_31__27_), .CI(u5_mult_87_SUMB_31__28_), .CO(
        u5_mult_87_CARRYB_32__27_), .S(u5_mult_87_SUMB_32__27_) );
  FA_X1 u5_mult_87_S2_32_26 ( .A(u5_mult_87_ab_32__26_), .B(
        u5_mult_87_CARRYB_31__26_), .CI(u5_mult_87_SUMB_31__27_), .CO(
        u5_mult_87_CARRYB_32__26_), .S(u5_mult_87_SUMB_32__26_) );
  FA_X1 u5_mult_87_S2_32_25 ( .A(u5_mult_87_ab_32__25_), .B(
        u5_mult_87_CARRYB_31__25_), .CI(u5_mult_87_SUMB_31__26_), .CO(
        u5_mult_87_CARRYB_32__25_), .S(u5_mult_87_SUMB_32__25_) );
  FA_X1 u5_mult_87_S2_32_24 ( .A(u5_mult_87_ab_32__24_), .B(
        u5_mult_87_CARRYB_31__24_), .CI(u5_mult_87_SUMB_31__25_), .CO(
        u5_mult_87_CARRYB_32__24_), .S(u5_mult_87_SUMB_32__24_) );
  FA_X1 u5_mult_87_S2_32_23 ( .A(u5_mult_87_ab_32__23_), .B(
        u5_mult_87_CARRYB_31__23_), .CI(u5_mult_87_SUMB_31__24_), .CO(
        u5_mult_87_CARRYB_32__23_), .S(u5_mult_87_SUMB_32__23_) );
  FA_X1 u5_mult_87_S2_32_22 ( .A(u5_mult_87_ab_32__22_), .B(
        u5_mult_87_CARRYB_31__22_), .CI(u5_mult_87_SUMB_31__23_), .CO(
        u5_mult_87_CARRYB_32__22_), .S(u5_mult_87_SUMB_32__22_) );
  FA_X1 u5_mult_87_S2_32_21 ( .A(u5_mult_87_ab_32__21_), .B(
        u5_mult_87_CARRYB_31__21_), .CI(u5_mult_87_SUMB_31__22_), .CO(
        u5_mult_87_CARRYB_32__21_), .S(u5_mult_87_SUMB_32__21_) );
  FA_X1 u5_mult_87_S2_32_20 ( .A(u5_mult_87_ab_32__20_), .B(
        u5_mult_87_CARRYB_31__20_), .CI(u5_mult_87_SUMB_31__21_), .CO(
        u5_mult_87_CARRYB_32__20_), .S(u5_mult_87_SUMB_32__20_) );
  FA_X1 u5_mult_87_S2_32_19 ( .A(u5_mult_87_ab_32__19_), .B(
        u5_mult_87_CARRYB_31__19_), .CI(u5_mult_87_SUMB_31__20_), .CO(
        u5_mult_87_CARRYB_32__19_), .S(u5_mult_87_SUMB_32__19_) );
  FA_X1 u5_mult_87_S2_32_18 ( .A(u5_mult_87_ab_32__18_), .B(
        u5_mult_87_CARRYB_31__18_), .CI(u5_mult_87_SUMB_31__19_), .CO(
        u5_mult_87_CARRYB_32__18_), .S(u5_mult_87_SUMB_32__18_) );
  FA_X1 u5_mult_87_S2_32_17 ( .A(u5_mult_87_ab_32__17_), .B(
        u5_mult_87_CARRYB_31__17_), .CI(u5_mult_87_SUMB_31__18_), .CO(
        u5_mult_87_CARRYB_32__17_), .S(u5_mult_87_SUMB_32__17_) );
  FA_X1 u5_mult_87_S2_32_16 ( .A(u5_mult_87_ab_32__16_), .B(
        u5_mult_87_CARRYB_31__16_), .CI(u5_mult_87_SUMB_31__17_), .CO(
        u5_mult_87_CARRYB_32__16_), .S(u5_mult_87_SUMB_32__16_) );
  FA_X1 u5_mult_87_S2_32_15 ( .A(u5_mult_87_ab_32__15_), .B(
        u5_mult_87_CARRYB_31__15_), .CI(u5_mult_87_SUMB_31__16_), .CO(
        u5_mult_87_CARRYB_32__15_), .S(u5_mult_87_SUMB_32__15_) );
  FA_X1 u5_mult_87_S2_32_14 ( .A(u5_mult_87_ab_32__14_), .B(
        u5_mult_87_CARRYB_31__14_), .CI(u5_mult_87_SUMB_31__15_), .CO(
        u5_mult_87_CARRYB_32__14_), .S(u5_mult_87_SUMB_32__14_) );
  FA_X1 u5_mult_87_S2_32_13 ( .A(u5_mult_87_ab_32__13_), .B(
        u5_mult_87_CARRYB_31__13_), .CI(u5_mult_87_SUMB_31__14_), .CO(
        u5_mult_87_CARRYB_32__13_), .S(u5_mult_87_SUMB_32__13_) );
  FA_X1 u5_mult_87_S2_32_12 ( .A(u5_mult_87_ab_32__12_), .B(
        u5_mult_87_CARRYB_31__12_), .CI(u5_mult_87_SUMB_31__13_), .CO(
        u5_mult_87_CARRYB_32__12_), .S(u5_mult_87_SUMB_32__12_) );
  FA_X1 u5_mult_87_S2_32_11 ( .A(u5_mult_87_ab_32__11_), .B(
        u5_mult_87_CARRYB_31__11_), .CI(u5_mult_87_SUMB_31__12_), .CO(
        u5_mult_87_CARRYB_32__11_), .S(u5_mult_87_SUMB_32__11_) );
  FA_X1 u5_mult_87_S2_32_10 ( .A(u5_mult_87_ab_32__10_), .B(
        u5_mult_87_CARRYB_31__10_), .CI(u5_mult_87_SUMB_31__11_), .CO(
        u5_mult_87_CARRYB_32__10_), .S(u5_mult_87_SUMB_32__10_) );
  FA_X1 u5_mult_87_S2_32_9 ( .A(u5_mult_87_ab_32__9_), .B(
        u5_mult_87_CARRYB_31__9_), .CI(u5_mult_87_SUMB_31__10_), .CO(
        u5_mult_87_CARRYB_32__9_), .S(u5_mult_87_SUMB_32__9_) );
  FA_X1 u5_mult_87_S2_32_8 ( .A(u5_mult_87_ab_32__8_), .B(
        u5_mult_87_CARRYB_31__8_), .CI(u5_mult_87_SUMB_31__9_), .CO(
        u5_mult_87_CARRYB_32__8_), .S(u5_mult_87_SUMB_32__8_) );
  FA_X1 u5_mult_87_S2_32_7 ( .A(u5_mult_87_ab_32__7_), .B(
        u5_mult_87_CARRYB_31__7_), .CI(u5_mult_87_SUMB_31__8_), .CO(
        u5_mult_87_CARRYB_32__7_), .S(u5_mult_87_SUMB_32__7_) );
  FA_X1 u5_mult_87_S2_32_6 ( .A(u5_mult_87_ab_32__6_), .B(
        u5_mult_87_CARRYB_31__6_), .CI(u5_mult_87_SUMB_31__7_), .CO(
        u5_mult_87_CARRYB_32__6_), .S(u5_mult_87_SUMB_32__6_) );
  FA_X1 u5_mult_87_S2_32_5 ( .A(u5_mult_87_ab_32__5_), .B(
        u5_mult_87_CARRYB_31__5_), .CI(u5_mult_87_SUMB_31__6_), .CO(
        u5_mult_87_CARRYB_32__5_), .S(u5_mult_87_SUMB_32__5_) );
  FA_X1 u5_mult_87_S2_32_4 ( .A(u5_mult_87_ab_32__4_), .B(
        u5_mult_87_CARRYB_31__4_), .CI(u5_mult_87_SUMB_31__5_), .CO(
        u5_mult_87_CARRYB_32__4_), .S(u5_mult_87_SUMB_32__4_) );
  FA_X1 u5_mult_87_S2_32_3 ( .A(u5_mult_87_ab_32__3_), .B(
        u5_mult_87_CARRYB_31__3_), .CI(u5_mult_87_SUMB_31__4_), .CO(
        u5_mult_87_CARRYB_32__3_), .S(u5_mult_87_SUMB_32__3_) );
  FA_X1 u5_mult_87_S2_32_2 ( .A(u5_mult_87_ab_32__2_), .B(
        u5_mult_87_CARRYB_31__2_), .CI(u5_mult_87_SUMB_31__3_), .CO(
        u5_mult_87_CARRYB_32__2_), .S(u5_mult_87_SUMB_32__2_) );
  FA_X1 u5_mult_87_S2_32_1 ( .A(u5_mult_87_ab_32__1_), .B(
        u5_mult_87_CARRYB_31__1_), .CI(u5_mult_87_SUMB_31__2_), .CO(
        u5_mult_87_CARRYB_32__1_), .S(u5_mult_87_SUMB_32__1_) );
  FA_X1 u5_mult_87_S1_32_0 ( .A(u5_mult_87_ab_32__0_), .B(
        u5_mult_87_CARRYB_31__0_), .CI(u5_mult_87_SUMB_31__1_), .CO(
        u5_mult_87_CARRYB_32__0_), .S(u5_N32) );
  FA_X1 u5_mult_87_S3_33_51 ( .A(u5_mult_87_ab_33__51_), .B(
        u5_mult_87_CARRYB_32__51_), .CI(u5_mult_87_ab_32__52_), .CO(
        u5_mult_87_CARRYB_33__51_), .S(u5_mult_87_SUMB_33__51_) );
  FA_X1 u5_mult_87_S2_33_50 ( .A(u5_mult_87_ab_33__50_), .B(
        u5_mult_87_CARRYB_32__50_), .CI(u5_mult_87_SUMB_32__51_), .CO(
        u5_mult_87_CARRYB_33__50_), .S(u5_mult_87_SUMB_33__50_) );
  FA_X1 u5_mult_87_S2_33_49 ( .A(u5_mult_87_ab_33__49_), .B(
        u5_mult_87_CARRYB_32__49_), .CI(u5_mult_87_SUMB_32__50_), .CO(
        u5_mult_87_CARRYB_33__49_), .S(u5_mult_87_SUMB_33__49_) );
  FA_X1 u5_mult_87_S2_33_48 ( .A(u5_mult_87_ab_33__48_), .B(
        u5_mult_87_CARRYB_32__48_), .CI(u5_mult_87_SUMB_32__49_), .CO(
        u5_mult_87_CARRYB_33__48_), .S(u5_mult_87_SUMB_33__48_) );
  FA_X1 u5_mult_87_S2_33_47 ( .A(u5_mult_87_ab_33__47_), .B(
        u5_mult_87_CARRYB_32__47_), .CI(u5_mult_87_SUMB_32__48_), .CO(
        u5_mult_87_CARRYB_33__47_), .S(u5_mult_87_SUMB_33__47_) );
  FA_X1 u5_mult_87_S2_33_46 ( .A(u5_mult_87_ab_33__46_), .B(
        u5_mult_87_CARRYB_32__46_), .CI(u5_mult_87_SUMB_32__47_), .CO(
        u5_mult_87_CARRYB_33__46_), .S(u5_mult_87_SUMB_33__46_) );
  FA_X1 u5_mult_87_S2_33_45 ( .A(u5_mult_87_ab_33__45_), .B(
        u5_mult_87_CARRYB_32__45_), .CI(u5_mult_87_SUMB_32__46_), .CO(
        u5_mult_87_CARRYB_33__45_), .S(u5_mult_87_SUMB_33__45_) );
  FA_X1 u5_mult_87_S2_33_44 ( .A(u5_mult_87_ab_33__44_), .B(
        u5_mult_87_CARRYB_32__44_), .CI(u5_mult_87_SUMB_32__45_), .CO(
        u5_mult_87_CARRYB_33__44_), .S(u5_mult_87_SUMB_33__44_) );
  FA_X1 u5_mult_87_S2_33_43 ( .A(u5_mult_87_ab_33__43_), .B(
        u5_mult_87_CARRYB_32__43_), .CI(u5_mult_87_SUMB_32__44_), .CO(
        u5_mult_87_CARRYB_33__43_), .S(u5_mult_87_SUMB_33__43_) );
  FA_X1 u5_mult_87_S2_33_42 ( .A(u5_mult_87_ab_33__42_), .B(
        u5_mult_87_CARRYB_32__42_), .CI(u5_mult_87_SUMB_32__43_), .CO(
        u5_mult_87_CARRYB_33__42_), .S(u5_mult_87_SUMB_33__42_) );
  FA_X1 u5_mult_87_S2_33_41 ( .A(u5_mult_87_ab_33__41_), .B(
        u5_mult_87_CARRYB_32__41_), .CI(u5_mult_87_SUMB_32__42_), .CO(
        u5_mult_87_CARRYB_33__41_), .S(u5_mult_87_SUMB_33__41_) );
  FA_X1 u5_mult_87_S2_33_40 ( .A(u5_mult_87_ab_33__40_), .B(
        u5_mult_87_CARRYB_32__40_), .CI(u5_mult_87_SUMB_32__41_), .CO(
        u5_mult_87_CARRYB_33__40_), .S(u5_mult_87_SUMB_33__40_) );
  FA_X1 u5_mult_87_S2_33_39 ( .A(u5_mult_87_ab_33__39_), .B(
        u5_mult_87_CARRYB_32__39_), .CI(u5_mult_87_SUMB_32__40_), .CO(
        u5_mult_87_CARRYB_33__39_), .S(u5_mult_87_SUMB_33__39_) );
  FA_X1 u5_mult_87_S2_33_38 ( .A(u5_mult_87_ab_33__38_), .B(
        u5_mult_87_CARRYB_32__38_), .CI(u5_mult_87_SUMB_32__39_), .CO(
        u5_mult_87_CARRYB_33__38_), .S(u5_mult_87_SUMB_33__38_) );
  FA_X1 u5_mult_87_S2_33_37 ( .A(u5_mult_87_ab_33__37_), .B(
        u5_mult_87_CARRYB_32__37_), .CI(u5_mult_87_SUMB_32__38_), .CO(
        u5_mult_87_CARRYB_33__37_), .S(u5_mult_87_SUMB_33__37_) );
  FA_X1 u5_mult_87_S2_33_36 ( .A(u5_mult_87_ab_33__36_), .B(
        u5_mult_87_CARRYB_32__36_), .CI(u5_mult_87_SUMB_32__37_), .CO(
        u5_mult_87_CARRYB_33__36_), .S(u5_mult_87_SUMB_33__36_) );
  FA_X1 u5_mult_87_S2_33_35 ( .A(u5_mult_87_ab_33__35_), .B(
        u5_mult_87_CARRYB_32__35_), .CI(u5_mult_87_SUMB_32__36_), .CO(
        u5_mult_87_CARRYB_33__35_), .S(u5_mult_87_SUMB_33__35_) );
  FA_X1 u5_mult_87_S2_33_34 ( .A(u5_mult_87_ab_33__34_), .B(
        u5_mult_87_CARRYB_32__34_), .CI(u5_mult_87_SUMB_32__35_), .CO(
        u5_mult_87_CARRYB_33__34_), .S(u5_mult_87_SUMB_33__34_) );
  FA_X1 u5_mult_87_S2_33_33 ( .A(u5_mult_87_ab_33__33_), .B(
        u5_mult_87_CARRYB_32__33_), .CI(u5_mult_87_SUMB_32__34_), .CO(
        u5_mult_87_CARRYB_33__33_), .S(u5_mult_87_SUMB_33__33_) );
  FA_X1 u5_mult_87_S2_33_32 ( .A(u5_mult_87_ab_33__32_), .B(
        u5_mult_87_CARRYB_32__32_), .CI(u5_mult_87_SUMB_32__33_), .CO(
        u5_mult_87_CARRYB_33__32_), .S(u5_mult_87_SUMB_33__32_) );
  FA_X1 u5_mult_87_S2_33_31 ( .A(u5_mult_87_ab_33__31_), .B(
        u5_mult_87_CARRYB_32__31_), .CI(u5_mult_87_SUMB_32__32_), .CO(
        u5_mult_87_CARRYB_33__31_), .S(u5_mult_87_SUMB_33__31_) );
  FA_X1 u5_mult_87_S2_33_30 ( .A(u5_mult_87_ab_33__30_), .B(
        u5_mult_87_CARRYB_32__30_), .CI(u5_mult_87_SUMB_32__31_), .CO(
        u5_mult_87_CARRYB_33__30_), .S(u5_mult_87_SUMB_33__30_) );
  FA_X1 u5_mult_87_S2_33_29 ( .A(u5_mult_87_ab_33__29_), .B(
        u5_mult_87_CARRYB_32__29_), .CI(u5_mult_87_SUMB_32__30_), .CO(
        u5_mult_87_CARRYB_33__29_), .S(u5_mult_87_SUMB_33__29_) );
  FA_X1 u5_mult_87_S2_33_28 ( .A(u5_mult_87_ab_33__28_), .B(
        u5_mult_87_CARRYB_32__28_), .CI(u5_mult_87_SUMB_32__29_), .CO(
        u5_mult_87_CARRYB_33__28_), .S(u5_mult_87_SUMB_33__28_) );
  FA_X1 u5_mult_87_S2_33_27 ( .A(u5_mult_87_ab_33__27_), .B(
        u5_mult_87_CARRYB_32__27_), .CI(u5_mult_87_SUMB_32__28_), .CO(
        u5_mult_87_CARRYB_33__27_), .S(u5_mult_87_SUMB_33__27_) );
  FA_X1 u5_mult_87_S2_33_26 ( .A(u5_mult_87_ab_33__26_), .B(
        u5_mult_87_CARRYB_32__26_), .CI(u5_mult_87_SUMB_32__27_), .CO(
        u5_mult_87_CARRYB_33__26_), .S(u5_mult_87_SUMB_33__26_) );
  FA_X1 u5_mult_87_S2_33_25 ( .A(u5_mult_87_ab_33__25_), .B(
        u5_mult_87_CARRYB_32__25_), .CI(u5_mult_87_SUMB_32__26_), .CO(
        u5_mult_87_CARRYB_33__25_), .S(u5_mult_87_SUMB_33__25_) );
  FA_X1 u5_mult_87_S2_33_24 ( .A(u5_mult_87_ab_33__24_), .B(
        u5_mult_87_CARRYB_32__24_), .CI(u5_mult_87_SUMB_32__25_), .CO(
        u5_mult_87_CARRYB_33__24_), .S(u5_mult_87_SUMB_33__24_) );
  FA_X1 u5_mult_87_S2_33_23 ( .A(u5_mult_87_ab_33__23_), .B(
        u5_mult_87_CARRYB_32__23_), .CI(u5_mult_87_SUMB_32__24_), .CO(
        u5_mult_87_CARRYB_33__23_), .S(u5_mult_87_SUMB_33__23_) );
  FA_X1 u5_mult_87_S2_33_22 ( .A(u5_mult_87_ab_33__22_), .B(
        u5_mult_87_CARRYB_32__22_), .CI(u5_mult_87_SUMB_32__23_), .CO(
        u5_mult_87_CARRYB_33__22_), .S(u5_mult_87_SUMB_33__22_) );
  FA_X1 u5_mult_87_S2_33_21 ( .A(u5_mult_87_ab_33__21_), .B(
        u5_mult_87_CARRYB_32__21_), .CI(u5_mult_87_SUMB_32__22_), .CO(
        u5_mult_87_CARRYB_33__21_), .S(u5_mult_87_SUMB_33__21_) );
  FA_X1 u5_mult_87_S2_33_20 ( .A(u5_mult_87_ab_33__20_), .B(
        u5_mult_87_CARRYB_32__20_), .CI(u5_mult_87_SUMB_32__21_), .CO(
        u5_mult_87_CARRYB_33__20_), .S(u5_mult_87_SUMB_33__20_) );
  FA_X1 u5_mult_87_S2_33_19 ( .A(u5_mult_87_ab_33__19_), .B(
        u5_mult_87_CARRYB_32__19_), .CI(u5_mult_87_SUMB_32__20_), .CO(
        u5_mult_87_CARRYB_33__19_), .S(u5_mult_87_SUMB_33__19_) );
  FA_X1 u5_mult_87_S2_33_18 ( .A(u5_mult_87_ab_33__18_), .B(
        u5_mult_87_CARRYB_32__18_), .CI(u5_mult_87_SUMB_32__19_), .CO(
        u5_mult_87_CARRYB_33__18_), .S(u5_mult_87_SUMB_33__18_) );
  FA_X1 u5_mult_87_S2_33_17 ( .A(u5_mult_87_ab_33__17_), .B(
        u5_mult_87_CARRYB_32__17_), .CI(u5_mult_87_SUMB_32__18_), .CO(
        u5_mult_87_CARRYB_33__17_), .S(u5_mult_87_SUMB_33__17_) );
  FA_X1 u5_mult_87_S2_33_16 ( .A(u5_mult_87_ab_33__16_), .B(
        u5_mult_87_CARRYB_32__16_), .CI(u5_mult_87_SUMB_32__17_), .CO(
        u5_mult_87_CARRYB_33__16_), .S(u5_mult_87_SUMB_33__16_) );
  FA_X1 u5_mult_87_S2_33_15 ( .A(u5_mult_87_ab_33__15_), .B(
        u5_mult_87_CARRYB_32__15_), .CI(u5_mult_87_SUMB_32__16_), .CO(
        u5_mult_87_CARRYB_33__15_), .S(u5_mult_87_SUMB_33__15_) );
  FA_X1 u5_mult_87_S2_33_14 ( .A(u5_mult_87_ab_33__14_), .B(
        u5_mult_87_CARRYB_32__14_), .CI(u5_mult_87_SUMB_32__15_), .CO(
        u5_mult_87_CARRYB_33__14_), .S(u5_mult_87_SUMB_33__14_) );
  FA_X1 u5_mult_87_S2_33_13 ( .A(u5_mult_87_ab_33__13_), .B(
        u5_mult_87_CARRYB_32__13_), .CI(u5_mult_87_SUMB_32__14_), .CO(
        u5_mult_87_CARRYB_33__13_), .S(u5_mult_87_SUMB_33__13_) );
  FA_X1 u5_mult_87_S2_33_12 ( .A(u5_mult_87_ab_33__12_), .B(
        u5_mult_87_CARRYB_32__12_), .CI(u5_mult_87_SUMB_32__13_), .CO(
        u5_mult_87_CARRYB_33__12_), .S(u5_mult_87_SUMB_33__12_) );
  FA_X1 u5_mult_87_S2_33_11 ( .A(u5_mult_87_ab_33__11_), .B(
        u5_mult_87_CARRYB_32__11_), .CI(u5_mult_87_SUMB_32__12_), .CO(
        u5_mult_87_CARRYB_33__11_), .S(u5_mult_87_SUMB_33__11_) );
  FA_X1 u5_mult_87_S2_33_10 ( .A(u5_mult_87_ab_33__10_), .B(
        u5_mult_87_CARRYB_32__10_), .CI(u5_mult_87_SUMB_32__11_), .CO(
        u5_mult_87_CARRYB_33__10_), .S(u5_mult_87_SUMB_33__10_) );
  FA_X1 u5_mult_87_S2_33_9 ( .A(u5_mult_87_ab_33__9_), .B(
        u5_mult_87_CARRYB_32__9_), .CI(u5_mult_87_SUMB_32__10_), .CO(
        u5_mult_87_CARRYB_33__9_), .S(u5_mult_87_SUMB_33__9_) );
  FA_X1 u5_mult_87_S2_33_8 ( .A(u5_mult_87_ab_33__8_), .B(
        u5_mult_87_CARRYB_32__8_), .CI(u5_mult_87_SUMB_32__9_), .CO(
        u5_mult_87_CARRYB_33__8_), .S(u5_mult_87_SUMB_33__8_) );
  FA_X1 u5_mult_87_S2_33_7 ( .A(u5_mult_87_ab_33__7_), .B(
        u5_mult_87_CARRYB_32__7_), .CI(u5_mult_87_SUMB_32__8_), .CO(
        u5_mult_87_CARRYB_33__7_), .S(u5_mult_87_SUMB_33__7_) );
  FA_X1 u5_mult_87_S2_33_6 ( .A(u5_mult_87_ab_33__6_), .B(
        u5_mult_87_CARRYB_32__6_), .CI(u5_mult_87_SUMB_32__7_), .CO(
        u5_mult_87_CARRYB_33__6_), .S(u5_mult_87_SUMB_33__6_) );
  FA_X1 u5_mult_87_S2_33_5 ( .A(u5_mult_87_ab_33__5_), .B(
        u5_mult_87_CARRYB_32__5_), .CI(u5_mult_87_SUMB_32__6_), .CO(
        u5_mult_87_CARRYB_33__5_), .S(u5_mult_87_SUMB_33__5_) );
  FA_X1 u5_mult_87_S2_33_4 ( .A(u5_mult_87_ab_33__4_), .B(
        u5_mult_87_CARRYB_32__4_), .CI(u5_mult_87_SUMB_32__5_), .CO(
        u5_mult_87_CARRYB_33__4_), .S(u5_mult_87_SUMB_33__4_) );
  FA_X1 u5_mult_87_S2_33_3 ( .A(u5_mult_87_ab_33__3_), .B(
        u5_mult_87_CARRYB_32__3_), .CI(u5_mult_87_SUMB_32__4_), .CO(
        u5_mult_87_CARRYB_33__3_), .S(u5_mult_87_SUMB_33__3_) );
  FA_X1 u5_mult_87_S2_33_2 ( .A(u5_mult_87_ab_33__2_), .B(
        u5_mult_87_CARRYB_32__2_), .CI(u5_mult_87_SUMB_32__3_), .CO(
        u5_mult_87_CARRYB_33__2_), .S(u5_mult_87_SUMB_33__2_) );
  FA_X1 u5_mult_87_S2_33_1 ( .A(u5_mult_87_ab_33__1_), .B(
        u5_mult_87_CARRYB_32__1_), .CI(u5_mult_87_SUMB_32__2_), .CO(
        u5_mult_87_CARRYB_33__1_), .S(u5_mult_87_SUMB_33__1_) );
  FA_X1 u5_mult_87_S1_33_0 ( .A(u5_mult_87_ab_33__0_), .B(
        u5_mult_87_CARRYB_32__0_), .CI(u5_mult_87_SUMB_32__1_), .CO(
        u5_mult_87_CARRYB_33__0_), .S(u5_N33) );
  FA_X1 u5_mult_87_S3_34_51 ( .A(u5_mult_87_ab_34__51_), .B(
        u5_mult_87_CARRYB_33__51_), .CI(u5_mult_87_ab_33__52_), .CO(
        u5_mult_87_CARRYB_34__51_), .S(u5_mult_87_SUMB_34__51_) );
  FA_X1 u5_mult_87_S2_34_50 ( .A(u5_mult_87_ab_34__50_), .B(
        u5_mult_87_CARRYB_33__50_), .CI(u5_mult_87_SUMB_33__51_), .CO(
        u5_mult_87_CARRYB_34__50_), .S(u5_mult_87_SUMB_34__50_) );
  FA_X1 u5_mult_87_S2_34_49 ( .A(u5_mult_87_ab_34__49_), .B(
        u5_mult_87_CARRYB_33__49_), .CI(u5_mult_87_SUMB_33__50_), .CO(
        u5_mult_87_CARRYB_34__49_), .S(u5_mult_87_SUMB_34__49_) );
  FA_X1 u5_mult_87_S2_34_48 ( .A(u5_mult_87_ab_34__48_), .B(
        u5_mult_87_CARRYB_33__48_), .CI(u5_mult_87_SUMB_33__49_), .CO(
        u5_mult_87_CARRYB_34__48_), .S(u5_mult_87_SUMB_34__48_) );
  FA_X1 u5_mult_87_S2_34_47 ( .A(u5_mult_87_ab_34__47_), .B(
        u5_mult_87_CARRYB_33__47_), .CI(u5_mult_87_SUMB_33__48_), .CO(
        u5_mult_87_CARRYB_34__47_), .S(u5_mult_87_SUMB_34__47_) );
  FA_X1 u5_mult_87_S2_34_46 ( .A(u5_mult_87_ab_34__46_), .B(
        u5_mult_87_CARRYB_33__46_), .CI(u5_mult_87_SUMB_33__47_), .CO(
        u5_mult_87_CARRYB_34__46_), .S(u5_mult_87_SUMB_34__46_) );
  FA_X1 u5_mult_87_S2_34_45 ( .A(u5_mult_87_ab_34__45_), .B(
        u5_mult_87_CARRYB_33__45_), .CI(u5_mult_87_SUMB_33__46_), .CO(
        u5_mult_87_CARRYB_34__45_), .S(u5_mult_87_SUMB_34__45_) );
  FA_X1 u5_mult_87_S2_34_44 ( .A(u5_mult_87_ab_34__44_), .B(
        u5_mult_87_CARRYB_33__44_), .CI(u5_mult_87_SUMB_33__45_), .CO(
        u5_mult_87_CARRYB_34__44_), .S(u5_mult_87_SUMB_34__44_) );
  FA_X1 u5_mult_87_S2_34_43 ( .A(u5_mult_87_ab_34__43_), .B(
        u5_mult_87_CARRYB_33__43_), .CI(u5_mult_87_SUMB_33__44_), .CO(
        u5_mult_87_CARRYB_34__43_), .S(u5_mult_87_SUMB_34__43_) );
  FA_X1 u5_mult_87_S2_34_42 ( .A(u5_mult_87_ab_34__42_), .B(
        u5_mult_87_CARRYB_33__42_), .CI(u5_mult_87_SUMB_33__43_), .CO(
        u5_mult_87_CARRYB_34__42_), .S(u5_mult_87_SUMB_34__42_) );
  FA_X1 u5_mult_87_S2_34_41 ( .A(u5_mult_87_ab_34__41_), .B(
        u5_mult_87_CARRYB_33__41_), .CI(u5_mult_87_SUMB_33__42_), .CO(
        u5_mult_87_CARRYB_34__41_), .S(u5_mult_87_SUMB_34__41_) );
  FA_X1 u5_mult_87_S2_34_40 ( .A(u5_mult_87_ab_34__40_), .B(
        u5_mult_87_CARRYB_33__40_), .CI(u5_mult_87_SUMB_33__41_), .CO(
        u5_mult_87_CARRYB_34__40_), .S(u5_mult_87_SUMB_34__40_) );
  FA_X1 u5_mult_87_S2_34_39 ( .A(u5_mult_87_ab_34__39_), .B(
        u5_mult_87_CARRYB_33__39_), .CI(u5_mult_87_SUMB_33__40_), .CO(
        u5_mult_87_CARRYB_34__39_), .S(u5_mult_87_SUMB_34__39_) );
  FA_X1 u5_mult_87_S2_34_38 ( .A(u5_mult_87_ab_34__38_), .B(
        u5_mult_87_CARRYB_33__38_), .CI(u5_mult_87_SUMB_33__39_), .CO(
        u5_mult_87_CARRYB_34__38_), .S(u5_mult_87_SUMB_34__38_) );
  FA_X1 u5_mult_87_S2_34_37 ( .A(u5_mult_87_ab_34__37_), .B(
        u5_mult_87_CARRYB_33__37_), .CI(u5_mult_87_SUMB_33__38_), .CO(
        u5_mult_87_CARRYB_34__37_), .S(u5_mult_87_SUMB_34__37_) );
  FA_X1 u5_mult_87_S2_34_36 ( .A(u5_mult_87_ab_34__36_), .B(
        u5_mult_87_CARRYB_33__36_), .CI(u5_mult_87_SUMB_33__37_), .CO(
        u5_mult_87_CARRYB_34__36_), .S(u5_mult_87_SUMB_34__36_) );
  FA_X1 u5_mult_87_S2_34_35 ( .A(u5_mult_87_ab_34__35_), .B(
        u5_mult_87_CARRYB_33__35_), .CI(u5_mult_87_SUMB_33__36_), .CO(
        u5_mult_87_CARRYB_34__35_), .S(u5_mult_87_SUMB_34__35_) );
  FA_X1 u5_mult_87_S2_34_34 ( .A(u5_mult_87_ab_34__34_), .B(
        u5_mult_87_CARRYB_33__34_), .CI(u5_mult_87_SUMB_33__35_), .CO(
        u5_mult_87_CARRYB_34__34_), .S(u5_mult_87_SUMB_34__34_) );
  FA_X1 u5_mult_87_S2_34_33 ( .A(u5_mult_87_ab_34__33_), .B(
        u5_mult_87_CARRYB_33__33_), .CI(u5_mult_87_SUMB_33__34_), .CO(
        u5_mult_87_CARRYB_34__33_), .S(u5_mult_87_SUMB_34__33_) );
  FA_X1 u5_mult_87_S2_34_32 ( .A(u5_mult_87_ab_34__32_), .B(
        u5_mult_87_CARRYB_33__32_), .CI(u5_mult_87_SUMB_33__33_), .CO(
        u5_mult_87_CARRYB_34__32_), .S(u5_mult_87_SUMB_34__32_) );
  FA_X1 u5_mult_87_S2_34_31 ( .A(u5_mult_87_ab_34__31_), .B(
        u5_mult_87_CARRYB_33__31_), .CI(u5_mult_87_SUMB_33__32_), .CO(
        u5_mult_87_CARRYB_34__31_), .S(u5_mult_87_SUMB_34__31_) );
  FA_X1 u5_mult_87_S2_34_30 ( .A(u5_mult_87_ab_34__30_), .B(
        u5_mult_87_CARRYB_33__30_), .CI(u5_mult_87_SUMB_33__31_), .CO(
        u5_mult_87_CARRYB_34__30_), .S(u5_mult_87_SUMB_34__30_) );
  FA_X1 u5_mult_87_S2_34_29 ( .A(u5_mult_87_ab_34__29_), .B(
        u5_mult_87_CARRYB_33__29_), .CI(u5_mult_87_SUMB_33__30_), .CO(
        u5_mult_87_CARRYB_34__29_), .S(u5_mult_87_SUMB_34__29_) );
  FA_X1 u5_mult_87_S2_34_28 ( .A(u5_mult_87_ab_34__28_), .B(
        u5_mult_87_CARRYB_33__28_), .CI(u5_mult_87_SUMB_33__29_), .CO(
        u5_mult_87_CARRYB_34__28_), .S(u5_mult_87_SUMB_34__28_) );
  FA_X1 u5_mult_87_S2_34_27 ( .A(u5_mult_87_ab_34__27_), .B(
        u5_mult_87_CARRYB_33__27_), .CI(u5_mult_87_SUMB_33__28_), .CO(
        u5_mult_87_CARRYB_34__27_), .S(u5_mult_87_SUMB_34__27_) );
  FA_X1 u5_mult_87_S2_34_26 ( .A(u5_mult_87_ab_34__26_), .B(
        u5_mult_87_CARRYB_33__26_), .CI(u5_mult_87_SUMB_33__27_), .CO(
        u5_mult_87_CARRYB_34__26_), .S(u5_mult_87_SUMB_34__26_) );
  FA_X1 u5_mult_87_S2_34_25 ( .A(u5_mult_87_ab_34__25_), .B(
        u5_mult_87_CARRYB_33__25_), .CI(u5_mult_87_SUMB_33__26_), .CO(
        u5_mult_87_CARRYB_34__25_), .S(u5_mult_87_SUMB_34__25_) );
  FA_X1 u5_mult_87_S2_34_24 ( .A(u5_mult_87_ab_34__24_), .B(
        u5_mult_87_CARRYB_33__24_), .CI(u5_mult_87_SUMB_33__25_), .CO(
        u5_mult_87_CARRYB_34__24_), .S(u5_mult_87_SUMB_34__24_) );
  FA_X1 u5_mult_87_S2_34_23 ( .A(u5_mult_87_ab_34__23_), .B(
        u5_mult_87_CARRYB_33__23_), .CI(u5_mult_87_SUMB_33__24_), .CO(
        u5_mult_87_CARRYB_34__23_), .S(u5_mult_87_SUMB_34__23_) );
  FA_X1 u5_mult_87_S2_34_22 ( .A(u5_mult_87_ab_34__22_), .B(
        u5_mult_87_CARRYB_33__22_), .CI(u5_mult_87_SUMB_33__23_), .CO(
        u5_mult_87_CARRYB_34__22_), .S(u5_mult_87_SUMB_34__22_) );
  FA_X1 u5_mult_87_S2_34_21 ( .A(u5_mult_87_ab_34__21_), .B(
        u5_mult_87_CARRYB_33__21_), .CI(u5_mult_87_SUMB_33__22_), .CO(
        u5_mult_87_CARRYB_34__21_), .S(u5_mult_87_SUMB_34__21_) );
  FA_X1 u5_mult_87_S2_34_20 ( .A(u5_mult_87_ab_34__20_), .B(
        u5_mult_87_CARRYB_33__20_), .CI(u5_mult_87_SUMB_33__21_), .CO(
        u5_mult_87_CARRYB_34__20_), .S(u5_mult_87_SUMB_34__20_) );
  FA_X1 u5_mult_87_S2_34_19 ( .A(u5_mult_87_ab_34__19_), .B(
        u5_mult_87_CARRYB_33__19_), .CI(u5_mult_87_SUMB_33__20_), .CO(
        u5_mult_87_CARRYB_34__19_), .S(u5_mult_87_SUMB_34__19_) );
  FA_X1 u5_mult_87_S2_34_18 ( .A(u5_mult_87_ab_34__18_), .B(
        u5_mult_87_CARRYB_33__18_), .CI(u5_mult_87_SUMB_33__19_), .CO(
        u5_mult_87_CARRYB_34__18_), .S(u5_mult_87_SUMB_34__18_) );
  FA_X1 u5_mult_87_S2_34_17 ( .A(u5_mult_87_ab_34__17_), .B(
        u5_mult_87_CARRYB_33__17_), .CI(u5_mult_87_SUMB_33__18_), .CO(
        u5_mult_87_CARRYB_34__17_), .S(u5_mult_87_SUMB_34__17_) );
  FA_X1 u5_mult_87_S2_34_16 ( .A(u5_mult_87_ab_34__16_), .B(
        u5_mult_87_CARRYB_33__16_), .CI(u5_mult_87_SUMB_33__17_), .CO(
        u5_mult_87_CARRYB_34__16_), .S(u5_mult_87_SUMB_34__16_) );
  FA_X1 u5_mult_87_S2_34_15 ( .A(u5_mult_87_ab_34__15_), .B(
        u5_mult_87_CARRYB_33__15_), .CI(u5_mult_87_SUMB_33__16_), .CO(
        u5_mult_87_CARRYB_34__15_), .S(u5_mult_87_SUMB_34__15_) );
  FA_X1 u5_mult_87_S2_34_14 ( .A(u5_mult_87_ab_34__14_), .B(
        u5_mult_87_CARRYB_33__14_), .CI(u5_mult_87_SUMB_33__15_), .CO(
        u5_mult_87_CARRYB_34__14_), .S(u5_mult_87_SUMB_34__14_) );
  FA_X1 u5_mult_87_S2_34_13 ( .A(u5_mult_87_ab_34__13_), .B(
        u5_mult_87_CARRYB_33__13_), .CI(u5_mult_87_SUMB_33__14_), .CO(
        u5_mult_87_CARRYB_34__13_), .S(u5_mult_87_SUMB_34__13_) );
  FA_X1 u5_mult_87_S2_34_12 ( .A(u5_mult_87_ab_34__12_), .B(
        u5_mult_87_CARRYB_33__12_), .CI(u5_mult_87_SUMB_33__13_), .CO(
        u5_mult_87_CARRYB_34__12_), .S(u5_mult_87_SUMB_34__12_) );
  FA_X1 u5_mult_87_S2_34_11 ( .A(u5_mult_87_ab_34__11_), .B(
        u5_mult_87_CARRYB_33__11_), .CI(u5_mult_87_SUMB_33__12_), .CO(
        u5_mult_87_CARRYB_34__11_), .S(u5_mult_87_SUMB_34__11_) );
  FA_X1 u5_mult_87_S2_34_10 ( .A(u5_mult_87_ab_34__10_), .B(
        u5_mult_87_CARRYB_33__10_), .CI(u5_mult_87_SUMB_33__11_), .CO(
        u5_mult_87_CARRYB_34__10_), .S(u5_mult_87_SUMB_34__10_) );
  FA_X1 u5_mult_87_S2_34_9 ( .A(u5_mult_87_ab_34__9_), .B(
        u5_mult_87_CARRYB_33__9_), .CI(u5_mult_87_SUMB_33__10_), .CO(
        u5_mult_87_CARRYB_34__9_), .S(u5_mult_87_SUMB_34__9_) );
  FA_X1 u5_mult_87_S2_34_8 ( .A(u5_mult_87_ab_34__8_), .B(
        u5_mult_87_CARRYB_33__8_), .CI(u5_mult_87_SUMB_33__9_), .CO(
        u5_mult_87_CARRYB_34__8_), .S(u5_mult_87_SUMB_34__8_) );
  FA_X1 u5_mult_87_S2_34_7 ( .A(u5_mult_87_ab_34__7_), .B(
        u5_mult_87_CARRYB_33__7_), .CI(u5_mult_87_SUMB_33__8_), .CO(
        u5_mult_87_CARRYB_34__7_), .S(u5_mult_87_SUMB_34__7_) );
  FA_X1 u5_mult_87_S2_34_6 ( .A(u5_mult_87_ab_34__6_), .B(
        u5_mult_87_CARRYB_33__6_), .CI(u5_mult_87_SUMB_33__7_), .CO(
        u5_mult_87_CARRYB_34__6_), .S(u5_mult_87_SUMB_34__6_) );
  FA_X1 u5_mult_87_S2_34_5 ( .A(u5_mult_87_ab_34__5_), .B(
        u5_mult_87_CARRYB_33__5_), .CI(u5_mult_87_SUMB_33__6_), .CO(
        u5_mult_87_CARRYB_34__5_), .S(u5_mult_87_SUMB_34__5_) );
  FA_X1 u5_mult_87_S2_34_4 ( .A(u5_mult_87_ab_34__4_), .B(
        u5_mult_87_CARRYB_33__4_), .CI(u5_mult_87_SUMB_33__5_), .CO(
        u5_mult_87_CARRYB_34__4_), .S(u5_mult_87_SUMB_34__4_) );
  FA_X1 u5_mult_87_S2_34_3 ( .A(u5_mult_87_ab_34__3_), .B(
        u5_mult_87_CARRYB_33__3_), .CI(u5_mult_87_SUMB_33__4_), .CO(
        u5_mult_87_CARRYB_34__3_), .S(u5_mult_87_SUMB_34__3_) );
  FA_X1 u5_mult_87_S2_34_2 ( .A(u5_mult_87_ab_34__2_), .B(
        u5_mult_87_CARRYB_33__2_), .CI(u5_mult_87_SUMB_33__3_), .CO(
        u5_mult_87_CARRYB_34__2_), .S(u5_mult_87_SUMB_34__2_) );
  FA_X1 u5_mult_87_S2_34_1 ( .A(u5_mult_87_ab_34__1_), .B(
        u5_mult_87_CARRYB_33__1_), .CI(u5_mult_87_SUMB_33__2_), .CO(
        u5_mult_87_CARRYB_34__1_), .S(u5_mult_87_SUMB_34__1_) );
  FA_X1 u5_mult_87_S1_34_0 ( .A(u5_mult_87_ab_34__0_), .B(
        u5_mult_87_CARRYB_33__0_), .CI(u5_mult_87_SUMB_33__1_), .CO(
        u5_mult_87_CARRYB_34__0_), .S(u5_N34) );
  FA_X1 u5_mult_87_S3_35_51 ( .A(u5_mult_87_ab_35__51_), .B(
        u5_mult_87_CARRYB_34__51_), .CI(u5_mult_87_ab_34__52_), .CO(
        u5_mult_87_CARRYB_35__51_), .S(u5_mult_87_SUMB_35__51_) );
  FA_X1 u5_mult_87_S2_35_50 ( .A(u5_mult_87_ab_35__50_), .B(
        u5_mult_87_CARRYB_34__50_), .CI(u5_mult_87_SUMB_34__51_), .CO(
        u5_mult_87_CARRYB_35__50_), .S(u5_mult_87_SUMB_35__50_) );
  FA_X1 u5_mult_87_S2_35_49 ( .A(u5_mult_87_ab_35__49_), .B(
        u5_mult_87_CARRYB_34__49_), .CI(u5_mult_87_SUMB_34__50_), .CO(
        u5_mult_87_CARRYB_35__49_), .S(u5_mult_87_SUMB_35__49_) );
  FA_X1 u5_mult_87_S2_35_48 ( .A(u5_mult_87_ab_35__48_), .B(
        u5_mult_87_CARRYB_34__48_), .CI(u5_mult_87_SUMB_34__49_), .CO(
        u5_mult_87_CARRYB_35__48_), .S(u5_mult_87_SUMB_35__48_) );
  FA_X1 u5_mult_87_S2_35_47 ( .A(u5_mult_87_ab_35__47_), .B(
        u5_mult_87_CARRYB_34__47_), .CI(u5_mult_87_SUMB_34__48_), .CO(
        u5_mult_87_CARRYB_35__47_), .S(u5_mult_87_SUMB_35__47_) );
  FA_X1 u5_mult_87_S2_35_46 ( .A(u5_mult_87_ab_35__46_), .B(
        u5_mult_87_CARRYB_34__46_), .CI(u5_mult_87_SUMB_34__47_), .CO(
        u5_mult_87_CARRYB_35__46_), .S(u5_mult_87_SUMB_35__46_) );
  FA_X1 u5_mult_87_S2_35_45 ( .A(u5_mult_87_ab_35__45_), .B(
        u5_mult_87_CARRYB_34__45_), .CI(u5_mult_87_SUMB_34__46_), .CO(
        u5_mult_87_CARRYB_35__45_), .S(u5_mult_87_SUMB_35__45_) );
  FA_X1 u5_mult_87_S2_35_44 ( .A(u5_mult_87_ab_35__44_), .B(
        u5_mult_87_CARRYB_34__44_), .CI(u5_mult_87_SUMB_34__45_), .CO(
        u5_mult_87_CARRYB_35__44_), .S(u5_mult_87_SUMB_35__44_) );
  FA_X1 u5_mult_87_S2_35_43 ( .A(u5_mult_87_ab_35__43_), .B(
        u5_mult_87_CARRYB_34__43_), .CI(u5_mult_87_SUMB_34__44_), .CO(
        u5_mult_87_CARRYB_35__43_), .S(u5_mult_87_SUMB_35__43_) );
  FA_X1 u5_mult_87_S2_35_42 ( .A(u5_mult_87_ab_35__42_), .B(
        u5_mult_87_CARRYB_34__42_), .CI(u5_mult_87_SUMB_34__43_), .CO(
        u5_mult_87_CARRYB_35__42_), .S(u5_mult_87_SUMB_35__42_) );
  FA_X1 u5_mult_87_S2_35_41 ( .A(u5_mult_87_ab_35__41_), .B(
        u5_mult_87_CARRYB_34__41_), .CI(u5_mult_87_SUMB_34__42_), .CO(
        u5_mult_87_CARRYB_35__41_), .S(u5_mult_87_SUMB_35__41_) );
  FA_X1 u5_mult_87_S2_35_40 ( .A(u5_mult_87_ab_35__40_), .B(
        u5_mult_87_CARRYB_34__40_), .CI(u5_mult_87_SUMB_34__41_), .CO(
        u5_mult_87_CARRYB_35__40_), .S(u5_mult_87_SUMB_35__40_) );
  FA_X1 u5_mult_87_S2_35_39 ( .A(u5_mult_87_ab_35__39_), .B(
        u5_mult_87_CARRYB_34__39_), .CI(u5_mult_87_SUMB_34__40_), .CO(
        u5_mult_87_CARRYB_35__39_), .S(u5_mult_87_SUMB_35__39_) );
  FA_X1 u5_mult_87_S2_35_38 ( .A(u5_mult_87_ab_35__38_), .B(
        u5_mult_87_CARRYB_34__38_), .CI(u5_mult_87_SUMB_34__39_), .CO(
        u5_mult_87_CARRYB_35__38_), .S(u5_mult_87_SUMB_35__38_) );
  FA_X1 u5_mult_87_S2_35_37 ( .A(u5_mult_87_ab_35__37_), .B(
        u5_mult_87_CARRYB_34__37_), .CI(u5_mult_87_SUMB_34__38_), .CO(
        u5_mult_87_CARRYB_35__37_), .S(u5_mult_87_SUMB_35__37_) );
  FA_X1 u5_mult_87_S2_35_36 ( .A(u5_mult_87_ab_35__36_), .B(
        u5_mult_87_CARRYB_34__36_), .CI(u5_mult_87_SUMB_34__37_), .CO(
        u5_mult_87_CARRYB_35__36_), .S(u5_mult_87_SUMB_35__36_) );
  FA_X1 u5_mult_87_S2_35_35 ( .A(u5_mult_87_ab_35__35_), .B(
        u5_mult_87_CARRYB_34__35_), .CI(u5_mult_87_SUMB_34__36_), .CO(
        u5_mult_87_CARRYB_35__35_), .S(u5_mult_87_SUMB_35__35_) );
  FA_X1 u5_mult_87_S2_35_34 ( .A(u5_mult_87_ab_35__34_), .B(
        u5_mult_87_CARRYB_34__34_), .CI(u5_mult_87_SUMB_34__35_), .CO(
        u5_mult_87_CARRYB_35__34_), .S(u5_mult_87_SUMB_35__34_) );
  FA_X1 u5_mult_87_S2_35_33 ( .A(u5_mult_87_ab_35__33_), .B(
        u5_mult_87_CARRYB_34__33_), .CI(u5_mult_87_SUMB_34__34_), .CO(
        u5_mult_87_CARRYB_35__33_), .S(u5_mult_87_SUMB_35__33_) );
  FA_X1 u5_mult_87_S2_35_32 ( .A(u5_mult_87_ab_35__32_), .B(
        u5_mult_87_CARRYB_34__32_), .CI(u5_mult_87_SUMB_34__33_), .CO(
        u5_mult_87_CARRYB_35__32_), .S(u5_mult_87_SUMB_35__32_) );
  FA_X1 u5_mult_87_S2_35_31 ( .A(u5_mult_87_ab_35__31_), .B(
        u5_mult_87_CARRYB_34__31_), .CI(u5_mult_87_SUMB_34__32_), .CO(
        u5_mult_87_CARRYB_35__31_), .S(u5_mult_87_SUMB_35__31_) );
  FA_X1 u5_mult_87_S2_35_30 ( .A(u5_mult_87_ab_35__30_), .B(
        u5_mult_87_CARRYB_34__30_), .CI(u5_mult_87_SUMB_34__31_), .CO(
        u5_mult_87_CARRYB_35__30_), .S(u5_mult_87_SUMB_35__30_) );
  FA_X1 u5_mult_87_S2_35_29 ( .A(u5_mult_87_ab_35__29_), .B(
        u5_mult_87_CARRYB_34__29_), .CI(u5_mult_87_SUMB_34__30_), .CO(
        u5_mult_87_CARRYB_35__29_), .S(u5_mult_87_SUMB_35__29_) );
  FA_X1 u5_mult_87_S2_35_28 ( .A(u5_mult_87_ab_35__28_), .B(
        u5_mult_87_CARRYB_34__28_), .CI(u5_mult_87_SUMB_34__29_), .CO(
        u5_mult_87_CARRYB_35__28_), .S(u5_mult_87_SUMB_35__28_) );
  FA_X1 u5_mult_87_S2_35_27 ( .A(u5_mult_87_ab_35__27_), .B(
        u5_mult_87_CARRYB_34__27_), .CI(u5_mult_87_SUMB_34__28_), .CO(
        u5_mult_87_CARRYB_35__27_), .S(u5_mult_87_SUMB_35__27_) );
  FA_X1 u5_mult_87_S2_35_26 ( .A(u5_mult_87_ab_35__26_), .B(
        u5_mult_87_CARRYB_34__26_), .CI(u5_mult_87_SUMB_34__27_), .CO(
        u5_mult_87_CARRYB_35__26_), .S(u5_mult_87_SUMB_35__26_) );
  FA_X1 u5_mult_87_S2_35_25 ( .A(u5_mult_87_ab_35__25_), .B(
        u5_mult_87_CARRYB_34__25_), .CI(u5_mult_87_SUMB_34__26_), .CO(
        u5_mult_87_CARRYB_35__25_), .S(u5_mult_87_SUMB_35__25_) );
  FA_X1 u5_mult_87_S2_35_24 ( .A(u5_mult_87_ab_35__24_), .B(
        u5_mult_87_CARRYB_34__24_), .CI(u5_mult_87_SUMB_34__25_), .CO(
        u5_mult_87_CARRYB_35__24_), .S(u5_mult_87_SUMB_35__24_) );
  FA_X1 u5_mult_87_S2_35_23 ( .A(u5_mult_87_ab_35__23_), .B(
        u5_mult_87_CARRYB_34__23_), .CI(u5_mult_87_SUMB_34__24_), .CO(
        u5_mult_87_CARRYB_35__23_), .S(u5_mult_87_SUMB_35__23_) );
  FA_X1 u5_mult_87_S2_35_22 ( .A(u5_mult_87_ab_35__22_), .B(
        u5_mult_87_CARRYB_34__22_), .CI(u5_mult_87_SUMB_34__23_), .CO(
        u5_mult_87_CARRYB_35__22_), .S(u5_mult_87_SUMB_35__22_) );
  FA_X1 u5_mult_87_S2_35_21 ( .A(u5_mult_87_ab_35__21_), .B(
        u5_mult_87_CARRYB_34__21_), .CI(u5_mult_87_SUMB_34__22_), .CO(
        u5_mult_87_CARRYB_35__21_), .S(u5_mult_87_SUMB_35__21_) );
  FA_X1 u5_mult_87_S2_35_20 ( .A(u5_mult_87_ab_35__20_), .B(
        u5_mult_87_CARRYB_34__20_), .CI(u5_mult_87_SUMB_34__21_), .CO(
        u5_mult_87_CARRYB_35__20_), .S(u5_mult_87_SUMB_35__20_) );
  FA_X1 u5_mult_87_S2_35_19 ( .A(u5_mult_87_ab_35__19_), .B(
        u5_mult_87_CARRYB_34__19_), .CI(u5_mult_87_SUMB_34__20_), .CO(
        u5_mult_87_CARRYB_35__19_), .S(u5_mult_87_SUMB_35__19_) );
  FA_X1 u5_mult_87_S2_35_18 ( .A(u5_mult_87_ab_35__18_), .B(
        u5_mult_87_CARRYB_34__18_), .CI(u5_mult_87_SUMB_34__19_), .CO(
        u5_mult_87_CARRYB_35__18_), .S(u5_mult_87_SUMB_35__18_) );
  FA_X1 u5_mult_87_S2_35_17 ( .A(u5_mult_87_ab_35__17_), .B(
        u5_mult_87_CARRYB_34__17_), .CI(u5_mult_87_SUMB_34__18_), .CO(
        u5_mult_87_CARRYB_35__17_), .S(u5_mult_87_SUMB_35__17_) );
  FA_X1 u5_mult_87_S2_35_16 ( .A(u5_mult_87_ab_35__16_), .B(
        u5_mult_87_CARRYB_34__16_), .CI(u5_mult_87_SUMB_34__17_), .CO(
        u5_mult_87_CARRYB_35__16_), .S(u5_mult_87_SUMB_35__16_) );
  FA_X1 u5_mult_87_S2_35_15 ( .A(u5_mult_87_ab_35__15_), .B(
        u5_mult_87_CARRYB_34__15_), .CI(u5_mult_87_SUMB_34__16_), .CO(
        u5_mult_87_CARRYB_35__15_), .S(u5_mult_87_SUMB_35__15_) );
  FA_X1 u5_mult_87_S2_35_14 ( .A(u5_mult_87_ab_35__14_), .B(
        u5_mult_87_CARRYB_34__14_), .CI(u5_mult_87_SUMB_34__15_), .CO(
        u5_mult_87_CARRYB_35__14_), .S(u5_mult_87_SUMB_35__14_) );
  FA_X1 u5_mult_87_S2_35_13 ( .A(u5_mult_87_ab_35__13_), .B(
        u5_mult_87_CARRYB_34__13_), .CI(u5_mult_87_SUMB_34__14_), .CO(
        u5_mult_87_CARRYB_35__13_), .S(u5_mult_87_SUMB_35__13_) );
  FA_X1 u5_mult_87_S2_35_12 ( .A(u5_mult_87_ab_35__12_), .B(
        u5_mult_87_CARRYB_34__12_), .CI(u5_mult_87_SUMB_34__13_), .CO(
        u5_mult_87_CARRYB_35__12_), .S(u5_mult_87_SUMB_35__12_) );
  FA_X1 u5_mult_87_S2_35_11 ( .A(u5_mult_87_ab_35__11_), .B(
        u5_mult_87_CARRYB_34__11_), .CI(u5_mult_87_SUMB_34__12_), .CO(
        u5_mult_87_CARRYB_35__11_), .S(u5_mult_87_SUMB_35__11_) );
  FA_X1 u5_mult_87_S2_35_10 ( .A(u5_mult_87_ab_35__10_), .B(
        u5_mult_87_CARRYB_34__10_), .CI(u5_mult_87_SUMB_34__11_), .CO(
        u5_mult_87_CARRYB_35__10_), .S(u5_mult_87_SUMB_35__10_) );
  FA_X1 u5_mult_87_S2_35_9 ( .A(u5_mult_87_ab_35__9_), .B(
        u5_mult_87_CARRYB_34__9_), .CI(u5_mult_87_SUMB_34__10_), .CO(
        u5_mult_87_CARRYB_35__9_), .S(u5_mult_87_SUMB_35__9_) );
  FA_X1 u5_mult_87_S2_35_8 ( .A(u5_mult_87_ab_35__8_), .B(
        u5_mult_87_CARRYB_34__8_), .CI(u5_mult_87_SUMB_34__9_), .CO(
        u5_mult_87_CARRYB_35__8_), .S(u5_mult_87_SUMB_35__8_) );
  FA_X1 u5_mult_87_S2_35_7 ( .A(u5_mult_87_ab_35__7_), .B(
        u5_mult_87_CARRYB_34__7_), .CI(u5_mult_87_SUMB_34__8_), .CO(
        u5_mult_87_CARRYB_35__7_), .S(u5_mult_87_SUMB_35__7_) );
  FA_X1 u5_mult_87_S2_35_6 ( .A(u5_mult_87_ab_35__6_), .B(
        u5_mult_87_CARRYB_34__6_), .CI(u5_mult_87_SUMB_34__7_), .CO(
        u5_mult_87_CARRYB_35__6_), .S(u5_mult_87_SUMB_35__6_) );
  FA_X1 u5_mult_87_S2_35_5 ( .A(u5_mult_87_ab_35__5_), .B(
        u5_mult_87_CARRYB_34__5_), .CI(u5_mult_87_SUMB_34__6_), .CO(
        u5_mult_87_CARRYB_35__5_), .S(u5_mult_87_SUMB_35__5_) );
  FA_X1 u5_mult_87_S2_35_4 ( .A(u5_mult_87_ab_35__4_), .B(
        u5_mult_87_CARRYB_34__4_), .CI(u5_mult_87_SUMB_34__5_), .CO(
        u5_mult_87_CARRYB_35__4_), .S(u5_mult_87_SUMB_35__4_) );
  FA_X1 u5_mult_87_S2_35_3 ( .A(u5_mult_87_ab_35__3_), .B(
        u5_mult_87_CARRYB_34__3_), .CI(u5_mult_87_SUMB_34__4_), .CO(
        u5_mult_87_CARRYB_35__3_), .S(u5_mult_87_SUMB_35__3_) );
  FA_X1 u5_mult_87_S2_35_2 ( .A(u5_mult_87_ab_35__2_), .B(
        u5_mult_87_CARRYB_34__2_), .CI(u5_mult_87_SUMB_34__3_), .CO(
        u5_mult_87_CARRYB_35__2_), .S(u5_mult_87_SUMB_35__2_) );
  FA_X1 u5_mult_87_S2_35_1 ( .A(u5_mult_87_ab_35__1_), .B(
        u5_mult_87_CARRYB_34__1_), .CI(u5_mult_87_SUMB_34__2_), .CO(
        u5_mult_87_CARRYB_35__1_), .S(u5_mult_87_SUMB_35__1_) );
  FA_X1 u5_mult_87_S1_35_0 ( .A(u5_mult_87_ab_35__0_), .B(
        u5_mult_87_CARRYB_34__0_), .CI(u5_mult_87_SUMB_34__1_), .CO(
        u5_mult_87_CARRYB_35__0_), .S(u5_N35) );
  FA_X1 u5_mult_87_S3_36_51 ( .A(u5_mult_87_ab_36__51_), .B(
        u5_mult_87_CARRYB_35__51_), .CI(u5_mult_87_ab_35__52_), .CO(
        u5_mult_87_CARRYB_36__51_), .S(u5_mult_87_SUMB_36__51_) );
  FA_X1 u5_mult_87_S2_36_50 ( .A(u5_mult_87_ab_36__50_), .B(
        u5_mult_87_CARRYB_35__50_), .CI(u5_mult_87_SUMB_35__51_), .CO(
        u5_mult_87_CARRYB_36__50_), .S(u5_mult_87_SUMB_36__50_) );
  FA_X1 u5_mult_87_S2_36_49 ( .A(u5_mult_87_ab_36__49_), .B(
        u5_mult_87_CARRYB_35__49_), .CI(u5_mult_87_SUMB_35__50_), .CO(
        u5_mult_87_CARRYB_36__49_), .S(u5_mult_87_SUMB_36__49_) );
  FA_X1 u5_mult_87_S2_36_48 ( .A(u5_mult_87_ab_36__48_), .B(
        u5_mult_87_CARRYB_35__48_), .CI(u5_mult_87_SUMB_35__49_), .CO(
        u5_mult_87_CARRYB_36__48_), .S(u5_mult_87_SUMB_36__48_) );
  FA_X1 u5_mult_87_S2_36_47 ( .A(u5_mult_87_ab_36__47_), .B(
        u5_mult_87_CARRYB_35__47_), .CI(u5_mult_87_SUMB_35__48_), .CO(
        u5_mult_87_CARRYB_36__47_), .S(u5_mult_87_SUMB_36__47_) );
  FA_X1 u5_mult_87_S2_36_46 ( .A(u5_mult_87_ab_36__46_), .B(
        u5_mult_87_CARRYB_35__46_), .CI(u5_mult_87_SUMB_35__47_), .CO(
        u5_mult_87_CARRYB_36__46_), .S(u5_mult_87_SUMB_36__46_) );
  FA_X1 u5_mult_87_S2_36_45 ( .A(u5_mult_87_ab_36__45_), .B(
        u5_mult_87_CARRYB_35__45_), .CI(u5_mult_87_SUMB_35__46_), .CO(
        u5_mult_87_CARRYB_36__45_), .S(u5_mult_87_SUMB_36__45_) );
  FA_X1 u5_mult_87_S2_36_44 ( .A(u5_mult_87_ab_36__44_), .B(
        u5_mult_87_CARRYB_35__44_), .CI(u5_mult_87_SUMB_35__45_), .CO(
        u5_mult_87_CARRYB_36__44_), .S(u5_mult_87_SUMB_36__44_) );
  FA_X1 u5_mult_87_S2_36_43 ( .A(u5_mult_87_ab_36__43_), .B(
        u5_mult_87_CARRYB_35__43_), .CI(u5_mult_87_SUMB_35__44_), .CO(
        u5_mult_87_CARRYB_36__43_), .S(u5_mult_87_SUMB_36__43_) );
  FA_X1 u5_mult_87_S2_36_42 ( .A(u5_mult_87_ab_36__42_), .B(
        u5_mult_87_CARRYB_35__42_), .CI(u5_mult_87_SUMB_35__43_), .CO(
        u5_mult_87_CARRYB_36__42_), .S(u5_mult_87_SUMB_36__42_) );
  FA_X1 u5_mult_87_S2_36_41 ( .A(u5_mult_87_ab_36__41_), .B(
        u5_mult_87_CARRYB_35__41_), .CI(u5_mult_87_SUMB_35__42_), .CO(
        u5_mult_87_CARRYB_36__41_), .S(u5_mult_87_SUMB_36__41_) );
  FA_X1 u5_mult_87_S2_36_40 ( .A(u5_mult_87_ab_36__40_), .B(
        u5_mult_87_CARRYB_35__40_), .CI(u5_mult_87_SUMB_35__41_), .CO(
        u5_mult_87_CARRYB_36__40_), .S(u5_mult_87_SUMB_36__40_) );
  FA_X1 u5_mult_87_S2_36_39 ( .A(u5_mult_87_ab_36__39_), .B(
        u5_mult_87_CARRYB_35__39_), .CI(u5_mult_87_SUMB_35__40_), .CO(
        u5_mult_87_CARRYB_36__39_), .S(u5_mult_87_SUMB_36__39_) );
  FA_X1 u5_mult_87_S2_36_38 ( .A(u5_mult_87_ab_36__38_), .B(
        u5_mult_87_CARRYB_35__38_), .CI(u5_mult_87_SUMB_35__39_), .CO(
        u5_mult_87_CARRYB_36__38_), .S(u5_mult_87_SUMB_36__38_) );
  FA_X1 u5_mult_87_S2_36_37 ( .A(u5_mult_87_ab_36__37_), .B(
        u5_mult_87_CARRYB_35__37_), .CI(u5_mult_87_SUMB_35__38_), .CO(
        u5_mult_87_CARRYB_36__37_), .S(u5_mult_87_SUMB_36__37_) );
  FA_X1 u5_mult_87_S2_36_36 ( .A(u5_mult_87_ab_36__36_), .B(
        u5_mult_87_CARRYB_35__36_), .CI(u5_mult_87_SUMB_35__37_), .CO(
        u5_mult_87_CARRYB_36__36_), .S(u5_mult_87_SUMB_36__36_) );
  FA_X1 u5_mult_87_S2_36_35 ( .A(u5_mult_87_ab_36__35_), .B(
        u5_mult_87_CARRYB_35__35_), .CI(u5_mult_87_SUMB_35__36_), .CO(
        u5_mult_87_CARRYB_36__35_), .S(u5_mult_87_SUMB_36__35_) );
  FA_X1 u5_mult_87_S2_36_34 ( .A(u5_mult_87_ab_36__34_), .B(
        u5_mult_87_CARRYB_35__34_), .CI(u5_mult_87_SUMB_35__35_), .CO(
        u5_mult_87_CARRYB_36__34_), .S(u5_mult_87_SUMB_36__34_) );
  FA_X1 u5_mult_87_S2_36_33 ( .A(u5_mult_87_ab_36__33_), .B(
        u5_mult_87_CARRYB_35__33_), .CI(u5_mult_87_SUMB_35__34_), .CO(
        u5_mult_87_CARRYB_36__33_), .S(u5_mult_87_SUMB_36__33_) );
  FA_X1 u5_mult_87_S2_36_32 ( .A(u5_mult_87_ab_36__32_), .B(
        u5_mult_87_CARRYB_35__32_), .CI(u5_mult_87_SUMB_35__33_), .CO(
        u5_mult_87_CARRYB_36__32_), .S(u5_mult_87_SUMB_36__32_) );
  FA_X1 u5_mult_87_S2_36_31 ( .A(u5_mult_87_ab_36__31_), .B(
        u5_mult_87_CARRYB_35__31_), .CI(u5_mult_87_SUMB_35__32_), .CO(
        u5_mult_87_CARRYB_36__31_), .S(u5_mult_87_SUMB_36__31_) );
  FA_X1 u5_mult_87_S2_36_30 ( .A(u5_mult_87_ab_36__30_), .B(
        u5_mult_87_CARRYB_35__30_), .CI(u5_mult_87_SUMB_35__31_), .CO(
        u5_mult_87_CARRYB_36__30_), .S(u5_mult_87_SUMB_36__30_) );
  FA_X1 u5_mult_87_S2_36_29 ( .A(u5_mult_87_ab_36__29_), .B(
        u5_mult_87_CARRYB_35__29_), .CI(u5_mult_87_SUMB_35__30_), .CO(
        u5_mult_87_CARRYB_36__29_), .S(u5_mult_87_SUMB_36__29_) );
  FA_X1 u5_mult_87_S2_36_28 ( .A(u5_mult_87_ab_36__28_), .B(
        u5_mult_87_CARRYB_35__28_), .CI(u5_mult_87_SUMB_35__29_), .CO(
        u5_mult_87_CARRYB_36__28_), .S(u5_mult_87_SUMB_36__28_) );
  FA_X1 u5_mult_87_S2_36_27 ( .A(u5_mult_87_ab_36__27_), .B(
        u5_mult_87_CARRYB_35__27_), .CI(u5_mult_87_SUMB_35__28_), .CO(
        u5_mult_87_CARRYB_36__27_), .S(u5_mult_87_SUMB_36__27_) );
  FA_X1 u5_mult_87_S2_36_26 ( .A(u5_mult_87_ab_36__26_), .B(
        u5_mult_87_CARRYB_35__26_), .CI(u5_mult_87_SUMB_35__27_), .CO(
        u5_mult_87_CARRYB_36__26_), .S(u5_mult_87_SUMB_36__26_) );
  FA_X1 u5_mult_87_S2_36_25 ( .A(u5_mult_87_ab_36__25_), .B(
        u5_mult_87_CARRYB_35__25_), .CI(u5_mult_87_SUMB_35__26_), .CO(
        u5_mult_87_CARRYB_36__25_), .S(u5_mult_87_SUMB_36__25_) );
  FA_X1 u5_mult_87_S2_36_24 ( .A(u5_mult_87_ab_36__24_), .B(
        u5_mult_87_CARRYB_35__24_), .CI(u5_mult_87_SUMB_35__25_), .CO(
        u5_mult_87_CARRYB_36__24_), .S(u5_mult_87_SUMB_36__24_) );
  FA_X1 u5_mult_87_S2_36_23 ( .A(u5_mult_87_ab_36__23_), .B(
        u5_mult_87_CARRYB_35__23_), .CI(u5_mult_87_SUMB_35__24_), .CO(
        u5_mult_87_CARRYB_36__23_), .S(u5_mult_87_SUMB_36__23_) );
  FA_X1 u5_mult_87_S2_36_22 ( .A(u5_mult_87_ab_36__22_), .B(
        u5_mult_87_CARRYB_35__22_), .CI(u5_mult_87_SUMB_35__23_), .CO(
        u5_mult_87_CARRYB_36__22_), .S(u5_mult_87_SUMB_36__22_) );
  FA_X1 u5_mult_87_S2_36_21 ( .A(u5_mult_87_ab_36__21_), .B(
        u5_mult_87_CARRYB_35__21_), .CI(u5_mult_87_SUMB_35__22_), .CO(
        u5_mult_87_CARRYB_36__21_), .S(u5_mult_87_SUMB_36__21_) );
  FA_X1 u5_mult_87_S2_36_20 ( .A(u5_mult_87_ab_36__20_), .B(
        u5_mult_87_CARRYB_35__20_), .CI(u5_mult_87_SUMB_35__21_), .CO(
        u5_mult_87_CARRYB_36__20_), .S(u5_mult_87_SUMB_36__20_) );
  FA_X1 u5_mult_87_S2_36_19 ( .A(u5_mult_87_ab_36__19_), .B(
        u5_mult_87_CARRYB_35__19_), .CI(u5_mult_87_SUMB_35__20_), .CO(
        u5_mult_87_CARRYB_36__19_), .S(u5_mult_87_SUMB_36__19_) );
  FA_X1 u5_mult_87_S2_36_18 ( .A(u5_mult_87_ab_36__18_), .B(
        u5_mult_87_CARRYB_35__18_), .CI(u5_mult_87_SUMB_35__19_), .CO(
        u5_mult_87_CARRYB_36__18_), .S(u5_mult_87_SUMB_36__18_) );
  FA_X1 u5_mult_87_S2_36_17 ( .A(u5_mult_87_ab_36__17_), .B(
        u5_mult_87_CARRYB_35__17_), .CI(u5_mult_87_SUMB_35__18_), .CO(
        u5_mult_87_CARRYB_36__17_), .S(u5_mult_87_SUMB_36__17_) );
  FA_X1 u5_mult_87_S2_36_16 ( .A(u5_mult_87_ab_36__16_), .B(
        u5_mult_87_CARRYB_35__16_), .CI(u5_mult_87_SUMB_35__17_), .CO(
        u5_mult_87_CARRYB_36__16_), .S(u5_mult_87_SUMB_36__16_) );
  FA_X1 u5_mult_87_S2_36_15 ( .A(u5_mult_87_ab_36__15_), .B(
        u5_mult_87_CARRYB_35__15_), .CI(u5_mult_87_SUMB_35__16_), .CO(
        u5_mult_87_CARRYB_36__15_), .S(u5_mult_87_SUMB_36__15_) );
  FA_X1 u5_mult_87_S2_36_14 ( .A(u5_mult_87_ab_36__14_), .B(
        u5_mult_87_CARRYB_35__14_), .CI(u5_mult_87_SUMB_35__15_), .CO(
        u5_mult_87_CARRYB_36__14_), .S(u5_mult_87_SUMB_36__14_) );
  FA_X1 u5_mult_87_S2_36_13 ( .A(u5_mult_87_ab_36__13_), .B(
        u5_mult_87_CARRYB_35__13_), .CI(u5_mult_87_SUMB_35__14_), .CO(
        u5_mult_87_CARRYB_36__13_), .S(u5_mult_87_SUMB_36__13_) );
  FA_X1 u5_mult_87_S2_36_12 ( .A(u5_mult_87_ab_36__12_), .B(
        u5_mult_87_CARRYB_35__12_), .CI(u5_mult_87_SUMB_35__13_), .CO(
        u5_mult_87_CARRYB_36__12_), .S(u5_mult_87_SUMB_36__12_) );
  FA_X1 u5_mult_87_S2_36_11 ( .A(u5_mult_87_ab_36__11_), .B(
        u5_mult_87_CARRYB_35__11_), .CI(u5_mult_87_SUMB_35__12_), .CO(
        u5_mult_87_CARRYB_36__11_), .S(u5_mult_87_SUMB_36__11_) );
  FA_X1 u5_mult_87_S2_36_10 ( .A(u5_mult_87_ab_36__10_), .B(
        u5_mult_87_CARRYB_35__10_), .CI(u5_mult_87_SUMB_35__11_), .CO(
        u5_mult_87_CARRYB_36__10_), .S(u5_mult_87_SUMB_36__10_) );
  FA_X1 u5_mult_87_S2_36_9 ( .A(u5_mult_87_ab_36__9_), .B(
        u5_mult_87_CARRYB_35__9_), .CI(u5_mult_87_SUMB_35__10_), .CO(
        u5_mult_87_CARRYB_36__9_), .S(u5_mult_87_SUMB_36__9_) );
  FA_X1 u5_mult_87_S2_36_8 ( .A(u5_mult_87_ab_36__8_), .B(
        u5_mult_87_CARRYB_35__8_), .CI(u5_mult_87_SUMB_35__9_), .CO(
        u5_mult_87_CARRYB_36__8_), .S(u5_mult_87_SUMB_36__8_) );
  FA_X1 u5_mult_87_S2_36_7 ( .A(u5_mult_87_ab_36__7_), .B(
        u5_mult_87_CARRYB_35__7_), .CI(u5_mult_87_SUMB_35__8_), .CO(
        u5_mult_87_CARRYB_36__7_), .S(u5_mult_87_SUMB_36__7_) );
  FA_X1 u5_mult_87_S2_36_6 ( .A(u5_mult_87_ab_36__6_), .B(
        u5_mult_87_CARRYB_35__6_), .CI(u5_mult_87_SUMB_35__7_), .CO(
        u5_mult_87_CARRYB_36__6_), .S(u5_mult_87_SUMB_36__6_) );
  FA_X1 u5_mult_87_S2_36_5 ( .A(u5_mult_87_ab_36__5_), .B(
        u5_mult_87_CARRYB_35__5_), .CI(u5_mult_87_SUMB_35__6_), .CO(
        u5_mult_87_CARRYB_36__5_), .S(u5_mult_87_SUMB_36__5_) );
  FA_X1 u5_mult_87_S2_36_4 ( .A(u5_mult_87_ab_36__4_), .B(
        u5_mult_87_CARRYB_35__4_), .CI(u5_mult_87_SUMB_35__5_), .CO(
        u5_mult_87_CARRYB_36__4_), .S(u5_mult_87_SUMB_36__4_) );
  FA_X1 u5_mult_87_S2_36_3 ( .A(u5_mult_87_ab_36__3_), .B(
        u5_mult_87_CARRYB_35__3_), .CI(u5_mult_87_SUMB_35__4_), .CO(
        u5_mult_87_CARRYB_36__3_), .S(u5_mult_87_SUMB_36__3_) );
  FA_X1 u5_mult_87_S2_36_2 ( .A(u5_mult_87_ab_36__2_), .B(
        u5_mult_87_CARRYB_35__2_), .CI(u5_mult_87_SUMB_35__3_), .CO(
        u5_mult_87_CARRYB_36__2_), .S(u5_mult_87_SUMB_36__2_) );
  FA_X1 u5_mult_87_S2_36_1 ( .A(u5_mult_87_ab_36__1_), .B(
        u5_mult_87_CARRYB_35__1_), .CI(u5_mult_87_SUMB_35__2_), .CO(
        u5_mult_87_CARRYB_36__1_), .S(u5_mult_87_SUMB_36__1_) );
  FA_X1 u5_mult_87_S1_36_0 ( .A(u5_mult_87_ab_36__0_), .B(
        u5_mult_87_CARRYB_35__0_), .CI(u5_mult_87_SUMB_35__1_), .CO(
        u5_mult_87_CARRYB_36__0_), .S(u5_N36) );
  FA_X1 u5_mult_87_S3_37_51 ( .A(u5_mult_87_ab_37__51_), .B(
        u5_mult_87_CARRYB_36__51_), .CI(u5_mult_87_ab_36__52_), .CO(
        u5_mult_87_CARRYB_37__51_), .S(u5_mult_87_SUMB_37__51_) );
  FA_X1 u5_mult_87_S2_37_50 ( .A(u5_mult_87_ab_37__50_), .B(
        u5_mult_87_CARRYB_36__50_), .CI(u5_mult_87_SUMB_36__51_), .CO(
        u5_mult_87_CARRYB_37__50_), .S(u5_mult_87_SUMB_37__50_) );
  FA_X1 u5_mult_87_S2_37_49 ( .A(u5_mult_87_ab_37__49_), .B(
        u5_mult_87_CARRYB_36__49_), .CI(u5_mult_87_SUMB_36__50_), .CO(
        u5_mult_87_CARRYB_37__49_), .S(u5_mult_87_SUMB_37__49_) );
  FA_X1 u5_mult_87_S2_37_48 ( .A(u5_mult_87_ab_37__48_), .B(
        u5_mult_87_CARRYB_36__48_), .CI(u5_mult_87_SUMB_36__49_), .CO(
        u5_mult_87_CARRYB_37__48_), .S(u5_mult_87_SUMB_37__48_) );
  FA_X1 u5_mult_87_S2_37_47 ( .A(u5_mult_87_ab_37__47_), .B(
        u5_mult_87_CARRYB_36__47_), .CI(u5_mult_87_SUMB_36__48_), .CO(
        u5_mult_87_CARRYB_37__47_), .S(u5_mult_87_SUMB_37__47_) );
  FA_X1 u5_mult_87_S2_37_46 ( .A(u5_mult_87_ab_37__46_), .B(
        u5_mult_87_CARRYB_36__46_), .CI(u5_mult_87_SUMB_36__47_), .CO(
        u5_mult_87_CARRYB_37__46_), .S(u5_mult_87_SUMB_37__46_) );
  FA_X1 u5_mult_87_S2_37_45 ( .A(u5_mult_87_ab_37__45_), .B(
        u5_mult_87_CARRYB_36__45_), .CI(u5_mult_87_SUMB_36__46_), .CO(
        u5_mult_87_CARRYB_37__45_), .S(u5_mult_87_SUMB_37__45_) );
  FA_X1 u5_mult_87_S2_37_44 ( .A(u5_mult_87_ab_37__44_), .B(
        u5_mult_87_CARRYB_36__44_), .CI(u5_mult_87_SUMB_36__45_), .CO(
        u5_mult_87_CARRYB_37__44_), .S(u5_mult_87_SUMB_37__44_) );
  FA_X1 u5_mult_87_S2_37_43 ( .A(u5_mult_87_ab_37__43_), .B(
        u5_mult_87_CARRYB_36__43_), .CI(u5_mult_87_SUMB_36__44_), .CO(
        u5_mult_87_CARRYB_37__43_), .S(u5_mult_87_SUMB_37__43_) );
  FA_X1 u5_mult_87_S2_37_42 ( .A(u5_mult_87_ab_37__42_), .B(
        u5_mult_87_CARRYB_36__42_), .CI(u5_mult_87_SUMB_36__43_), .CO(
        u5_mult_87_CARRYB_37__42_), .S(u5_mult_87_SUMB_37__42_) );
  FA_X1 u5_mult_87_S2_37_41 ( .A(u5_mult_87_ab_37__41_), .B(
        u5_mult_87_CARRYB_36__41_), .CI(u5_mult_87_SUMB_36__42_), .CO(
        u5_mult_87_CARRYB_37__41_), .S(u5_mult_87_SUMB_37__41_) );
  FA_X1 u5_mult_87_S2_37_40 ( .A(u5_mult_87_ab_37__40_), .B(
        u5_mult_87_CARRYB_36__40_), .CI(u5_mult_87_SUMB_36__41_), .CO(
        u5_mult_87_CARRYB_37__40_), .S(u5_mult_87_SUMB_37__40_) );
  FA_X1 u5_mult_87_S2_37_39 ( .A(u5_mult_87_ab_37__39_), .B(
        u5_mult_87_CARRYB_36__39_), .CI(u5_mult_87_SUMB_36__40_), .CO(
        u5_mult_87_CARRYB_37__39_), .S(u5_mult_87_SUMB_37__39_) );
  FA_X1 u5_mult_87_S2_37_38 ( .A(u5_mult_87_ab_37__38_), .B(
        u5_mult_87_CARRYB_36__38_), .CI(u5_mult_87_SUMB_36__39_), .CO(
        u5_mult_87_CARRYB_37__38_), .S(u5_mult_87_SUMB_37__38_) );
  FA_X1 u5_mult_87_S2_37_37 ( .A(u5_mult_87_ab_37__37_), .B(
        u5_mult_87_CARRYB_36__37_), .CI(u5_mult_87_SUMB_36__38_), .CO(
        u5_mult_87_CARRYB_37__37_), .S(u5_mult_87_SUMB_37__37_) );
  FA_X1 u5_mult_87_S2_37_36 ( .A(u5_mult_87_ab_37__36_), .B(
        u5_mult_87_CARRYB_36__36_), .CI(u5_mult_87_SUMB_36__37_), .CO(
        u5_mult_87_CARRYB_37__36_), .S(u5_mult_87_SUMB_37__36_) );
  FA_X1 u5_mult_87_S2_37_35 ( .A(u5_mult_87_ab_37__35_), .B(
        u5_mult_87_CARRYB_36__35_), .CI(u5_mult_87_SUMB_36__36_), .CO(
        u5_mult_87_CARRYB_37__35_), .S(u5_mult_87_SUMB_37__35_) );
  FA_X1 u5_mult_87_S2_37_34 ( .A(u5_mult_87_ab_37__34_), .B(
        u5_mult_87_CARRYB_36__34_), .CI(u5_mult_87_SUMB_36__35_), .CO(
        u5_mult_87_CARRYB_37__34_), .S(u5_mult_87_SUMB_37__34_) );
  FA_X1 u5_mult_87_S2_37_33 ( .A(u5_mult_87_ab_37__33_), .B(
        u5_mult_87_CARRYB_36__33_), .CI(u5_mult_87_SUMB_36__34_), .CO(
        u5_mult_87_CARRYB_37__33_), .S(u5_mult_87_SUMB_37__33_) );
  FA_X1 u5_mult_87_S2_37_32 ( .A(u5_mult_87_ab_37__32_), .B(
        u5_mult_87_CARRYB_36__32_), .CI(u5_mult_87_SUMB_36__33_), .CO(
        u5_mult_87_CARRYB_37__32_), .S(u5_mult_87_SUMB_37__32_) );
  FA_X1 u5_mult_87_S2_37_31 ( .A(u5_mult_87_ab_37__31_), .B(
        u5_mult_87_CARRYB_36__31_), .CI(u5_mult_87_SUMB_36__32_), .CO(
        u5_mult_87_CARRYB_37__31_), .S(u5_mult_87_SUMB_37__31_) );
  FA_X1 u5_mult_87_S2_37_30 ( .A(u5_mult_87_ab_37__30_), .B(
        u5_mult_87_CARRYB_36__30_), .CI(u5_mult_87_SUMB_36__31_), .CO(
        u5_mult_87_CARRYB_37__30_), .S(u5_mult_87_SUMB_37__30_) );
  FA_X1 u5_mult_87_S2_37_29 ( .A(u5_mult_87_ab_37__29_), .B(
        u5_mult_87_CARRYB_36__29_), .CI(u5_mult_87_SUMB_36__30_), .CO(
        u5_mult_87_CARRYB_37__29_), .S(u5_mult_87_SUMB_37__29_) );
  FA_X1 u5_mult_87_S2_37_28 ( .A(u5_mult_87_ab_37__28_), .B(
        u5_mult_87_CARRYB_36__28_), .CI(u5_mult_87_SUMB_36__29_), .CO(
        u5_mult_87_CARRYB_37__28_), .S(u5_mult_87_SUMB_37__28_) );
  FA_X1 u5_mult_87_S2_37_27 ( .A(u5_mult_87_ab_37__27_), .B(
        u5_mult_87_CARRYB_36__27_), .CI(u5_mult_87_SUMB_36__28_), .CO(
        u5_mult_87_CARRYB_37__27_), .S(u5_mult_87_SUMB_37__27_) );
  FA_X1 u5_mult_87_S2_37_26 ( .A(u5_mult_87_ab_37__26_), .B(
        u5_mult_87_CARRYB_36__26_), .CI(u5_mult_87_SUMB_36__27_), .CO(
        u5_mult_87_CARRYB_37__26_), .S(u5_mult_87_SUMB_37__26_) );
  FA_X1 u5_mult_87_S2_37_25 ( .A(u5_mult_87_ab_37__25_), .B(
        u5_mult_87_CARRYB_36__25_), .CI(u5_mult_87_SUMB_36__26_), .CO(
        u5_mult_87_CARRYB_37__25_), .S(u5_mult_87_SUMB_37__25_) );
  FA_X1 u5_mult_87_S2_37_24 ( .A(u5_mult_87_ab_37__24_), .B(
        u5_mult_87_CARRYB_36__24_), .CI(u5_mult_87_SUMB_36__25_), .CO(
        u5_mult_87_CARRYB_37__24_), .S(u5_mult_87_SUMB_37__24_) );
  FA_X1 u5_mult_87_S2_37_23 ( .A(u5_mult_87_ab_37__23_), .B(
        u5_mult_87_CARRYB_36__23_), .CI(u5_mult_87_SUMB_36__24_), .CO(
        u5_mult_87_CARRYB_37__23_), .S(u5_mult_87_SUMB_37__23_) );
  FA_X1 u5_mult_87_S2_37_22 ( .A(u5_mult_87_ab_37__22_), .B(
        u5_mult_87_CARRYB_36__22_), .CI(u5_mult_87_SUMB_36__23_), .CO(
        u5_mult_87_CARRYB_37__22_), .S(u5_mult_87_SUMB_37__22_) );
  FA_X1 u5_mult_87_S2_37_21 ( .A(u5_mult_87_ab_37__21_), .B(
        u5_mult_87_CARRYB_36__21_), .CI(u5_mult_87_SUMB_36__22_), .CO(
        u5_mult_87_CARRYB_37__21_), .S(u5_mult_87_SUMB_37__21_) );
  FA_X1 u5_mult_87_S2_37_20 ( .A(u5_mult_87_ab_37__20_), .B(
        u5_mult_87_CARRYB_36__20_), .CI(u5_mult_87_SUMB_36__21_), .CO(
        u5_mult_87_CARRYB_37__20_), .S(u5_mult_87_SUMB_37__20_) );
  FA_X1 u5_mult_87_S2_37_19 ( .A(u5_mult_87_ab_37__19_), .B(
        u5_mult_87_CARRYB_36__19_), .CI(u5_mult_87_SUMB_36__20_), .CO(
        u5_mult_87_CARRYB_37__19_), .S(u5_mult_87_SUMB_37__19_) );
  FA_X1 u5_mult_87_S2_37_18 ( .A(u5_mult_87_ab_37__18_), .B(
        u5_mult_87_CARRYB_36__18_), .CI(u5_mult_87_SUMB_36__19_), .CO(
        u5_mult_87_CARRYB_37__18_), .S(u5_mult_87_SUMB_37__18_) );
  FA_X1 u5_mult_87_S2_37_17 ( .A(u5_mult_87_ab_37__17_), .B(
        u5_mult_87_CARRYB_36__17_), .CI(u5_mult_87_SUMB_36__18_), .CO(
        u5_mult_87_CARRYB_37__17_), .S(u5_mult_87_SUMB_37__17_) );
  FA_X1 u5_mult_87_S2_37_16 ( .A(u5_mult_87_ab_37__16_), .B(
        u5_mult_87_CARRYB_36__16_), .CI(u5_mult_87_SUMB_36__17_), .CO(
        u5_mult_87_CARRYB_37__16_), .S(u5_mult_87_SUMB_37__16_) );
  FA_X1 u5_mult_87_S2_37_15 ( .A(u5_mult_87_ab_37__15_), .B(
        u5_mult_87_CARRYB_36__15_), .CI(u5_mult_87_SUMB_36__16_), .CO(
        u5_mult_87_CARRYB_37__15_), .S(u5_mult_87_SUMB_37__15_) );
  FA_X1 u5_mult_87_S2_37_14 ( .A(u5_mult_87_ab_37__14_), .B(
        u5_mult_87_CARRYB_36__14_), .CI(u5_mult_87_SUMB_36__15_), .CO(
        u5_mult_87_CARRYB_37__14_), .S(u5_mult_87_SUMB_37__14_) );
  FA_X1 u5_mult_87_S2_37_13 ( .A(u5_mult_87_ab_37__13_), .B(
        u5_mult_87_CARRYB_36__13_), .CI(u5_mult_87_SUMB_36__14_), .CO(
        u5_mult_87_CARRYB_37__13_), .S(u5_mult_87_SUMB_37__13_) );
  FA_X1 u5_mult_87_S2_37_12 ( .A(u5_mult_87_ab_37__12_), .B(
        u5_mult_87_CARRYB_36__12_), .CI(u5_mult_87_SUMB_36__13_), .CO(
        u5_mult_87_CARRYB_37__12_), .S(u5_mult_87_SUMB_37__12_) );
  FA_X1 u5_mult_87_S2_37_11 ( .A(u5_mult_87_ab_37__11_), .B(
        u5_mult_87_CARRYB_36__11_), .CI(u5_mult_87_SUMB_36__12_), .CO(
        u5_mult_87_CARRYB_37__11_), .S(u5_mult_87_SUMB_37__11_) );
  FA_X1 u5_mult_87_S2_37_10 ( .A(u5_mult_87_ab_37__10_), .B(
        u5_mult_87_CARRYB_36__10_), .CI(u5_mult_87_SUMB_36__11_), .CO(
        u5_mult_87_CARRYB_37__10_), .S(u5_mult_87_SUMB_37__10_) );
  FA_X1 u5_mult_87_S2_37_9 ( .A(u5_mult_87_ab_37__9_), .B(
        u5_mult_87_CARRYB_36__9_), .CI(u5_mult_87_SUMB_36__10_), .CO(
        u5_mult_87_CARRYB_37__9_), .S(u5_mult_87_SUMB_37__9_) );
  FA_X1 u5_mult_87_S2_37_8 ( .A(u5_mult_87_ab_37__8_), .B(
        u5_mult_87_CARRYB_36__8_), .CI(u5_mult_87_SUMB_36__9_), .CO(
        u5_mult_87_CARRYB_37__8_), .S(u5_mult_87_SUMB_37__8_) );
  FA_X1 u5_mult_87_S2_37_7 ( .A(u5_mult_87_ab_37__7_), .B(
        u5_mult_87_CARRYB_36__7_), .CI(u5_mult_87_SUMB_36__8_), .CO(
        u5_mult_87_CARRYB_37__7_), .S(u5_mult_87_SUMB_37__7_) );
  FA_X1 u5_mult_87_S2_37_6 ( .A(u5_mult_87_ab_37__6_), .B(
        u5_mult_87_CARRYB_36__6_), .CI(u5_mult_87_SUMB_36__7_), .CO(
        u5_mult_87_CARRYB_37__6_), .S(u5_mult_87_SUMB_37__6_) );
  FA_X1 u5_mult_87_S2_37_5 ( .A(u5_mult_87_ab_37__5_), .B(
        u5_mult_87_CARRYB_36__5_), .CI(u5_mult_87_SUMB_36__6_), .CO(
        u5_mult_87_CARRYB_37__5_), .S(u5_mult_87_SUMB_37__5_) );
  FA_X1 u5_mult_87_S2_37_4 ( .A(u5_mult_87_ab_37__4_), .B(
        u5_mult_87_CARRYB_36__4_), .CI(u5_mult_87_SUMB_36__5_), .CO(
        u5_mult_87_CARRYB_37__4_), .S(u5_mult_87_SUMB_37__4_) );
  FA_X1 u5_mult_87_S2_37_3 ( .A(u5_mult_87_ab_37__3_), .B(
        u5_mult_87_CARRYB_36__3_), .CI(u5_mult_87_SUMB_36__4_), .CO(
        u5_mult_87_CARRYB_37__3_), .S(u5_mult_87_SUMB_37__3_) );
  FA_X1 u5_mult_87_S2_37_2 ( .A(u5_mult_87_ab_37__2_), .B(
        u5_mult_87_CARRYB_36__2_), .CI(u5_mult_87_SUMB_36__3_), .CO(
        u5_mult_87_CARRYB_37__2_), .S(u5_mult_87_SUMB_37__2_) );
  FA_X1 u5_mult_87_S2_37_1 ( .A(u5_mult_87_ab_37__1_), .B(
        u5_mult_87_CARRYB_36__1_), .CI(u5_mult_87_SUMB_36__2_), .CO(
        u5_mult_87_CARRYB_37__1_), .S(u5_mult_87_SUMB_37__1_) );
  FA_X1 u5_mult_87_S1_37_0 ( .A(u5_mult_87_ab_37__0_), .B(
        u5_mult_87_CARRYB_36__0_), .CI(u5_mult_87_SUMB_36__1_), .CO(
        u5_mult_87_CARRYB_37__0_), .S(u5_N37) );
  FA_X1 u5_mult_87_S3_38_51 ( .A(u5_mult_87_ab_38__51_), .B(
        u5_mult_87_CARRYB_37__51_), .CI(u5_mult_87_ab_37__52_), .CO(
        u5_mult_87_CARRYB_38__51_), .S(u5_mult_87_SUMB_38__51_) );
  FA_X1 u5_mult_87_S2_38_50 ( .A(u5_mult_87_ab_38__50_), .B(
        u5_mult_87_CARRYB_37__50_), .CI(u5_mult_87_SUMB_37__51_), .CO(
        u5_mult_87_CARRYB_38__50_), .S(u5_mult_87_SUMB_38__50_) );
  FA_X1 u5_mult_87_S2_38_49 ( .A(u5_mult_87_ab_38__49_), .B(
        u5_mult_87_CARRYB_37__49_), .CI(u5_mult_87_SUMB_37__50_), .CO(
        u5_mult_87_CARRYB_38__49_), .S(u5_mult_87_SUMB_38__49_) );
  FA_X1 u5_mult_87_S2_38_48 ( .A(u5_mult_87_ab_38__48_), .B(
        u5_mult_87_CARRYB_37__48_), .CI(u5_mult_87_SUMB_37__49_), .CO(
        u5_mult_87_CARRYB_38__48_), .S(u5_mult_87_SUMB_38__48_) );
  FA_X1 u5_mult_87_S2_38_47 ( .A(u5_mult_87_ab_38__47_), .B(
        u5_mult_87_CARRYB_37__47_), .CI(u5_mult_87_SUMB_37__48_), .CO(
        u5_mult_87_CARRYB_38__47_), .S(u5_mult_87_SUMB_38__47_) );
  FA_X1 u5_mult_87_S2_38_46 ( .A(u5_mult_87_ab_38__46_), .B(
        u5_mult_87_CARRYB_37__46_), .CI(u5_mult_87_SUMB_37__47_), .CO(
        u5_mult_87_CARRYB_38__46_), .S(u5_mult_87_SUMB_38__46_) );
  FA_X1 u5_mult_87_S2_38_45 ( .A(u5_mult_87_ab_38__45_), .B(
        u5_mult_87_CARRYB_37__45_), .CI(u5_mult_87_SUMB_37__46_), .CO(
        u5_mult_87_CARRYB_38__45_), .S(u5_mult_87_SUMB_38__45_) );
  FA_X1 u5_mult_87_S2_38_44 ( .A(u5_mult_87_ab_38__44_), .B(
        u5_mult_87_CARRYB_37__44_), .CI(u5_mult_87_SUMB_37__45_), .CO(
        u5_mult_87_CARRYB_38__44_), .S(u5_mult_87_SUMB_38__44_) );
  FA_X1 u5_mult_87_S2_38_43 ( .A(u5_mult_87_ab_38__43_), .B(
        u5_mult_87_CARRYB_37__43_), .CI(u5_mult_87_SUMB_37__44_), .CO(
        u5_mult_87_CARRYB_38__43_), .S(u5_mult_87_SUMB_38__43_) );
  FA_X1 u5_mult_87_S2_38_42 ( .A(u5_mult_87_ab_38__42_), .B(
        u5_mult_87_CARRYB_37__42_), .CI(u5_mult_87_SUMB_37__43_), .CO(
        u5_mult_87_CARRYB_38__42_), .S(u5_mult_87_SUMB_38__42_) );
  FA_X1 u5_mult_87_S2_38_41 ( .A(u5_mult_87_ab_38__41_), .B(
        u5_mult_87_CARRYB_37__41_), .CI(u5_mult_87_SUMB_37__42_), .CO(
        u5_mult_87_CARRYB_38__41_), .S(u5_mult_87_SUMB_38__41_) );
  FA_X1 u5_mult_87_S2_38_40 ( .A(u5_mult_87_ab_38__40_), .B(
        u5_mult_87_CARRYB_37__40_), .CI(u5_mult_87_SUMB_37__41_), .CO(
        u5_mult_87_CARRYB_38__40_), .S(u5_mult_87_SUMB_38__40_) );
  FA_X1 u5_mult_87_S2_38_39 ( .A(u5_mult_87_ab_38__39_), .B(
        u5_mult_87_CARRYB_37__39_), .CI(u5_mult_87_SUMB_37__40_), .CO(
        u5_mult_87_CARRYB_38__39_), .S(u5_mult_87_SUMB_38__39_) );
  FA_X1 u5_mult_87_S2_38_38 ( .A(u5_mult_87_ab_38__38_), .B(
        u5_mult_87_CARRYB_37__38_), .CI(u5_mult_87_SUMB_37__39_), .CO(
        u5_mult_87_CARRYB_38__38_), .S(u5_mult_87_SUMB_38__38_) );
  FA_X1 u5_mult_87_S2_38_37 ( .A(u5_mult_87_ab_38__37_), .B(
        u5_mult_87_CARRYB_37__37_), .CI(u5_mult_87_SUMB_37__38_), .CO(
        u5_mult_87_CARRYB_38__37_), .S(u5_mult_87_SUMB_38__37_) );
  FA_X1 u5_mult_87_S2_38_36 ( .A(u5_mult_87_ab_38__36_), .B(
        u5_mult_87_CARRYB_37__36_), .CI(u5_mult_87_SUMB_37__37_), .CO(
        u5_mult_87_CARRYB_38__36_), .S(u5_mult_87_SUMB_38__36_) );
  FA_X1 u5_mult_87_S2_38_35 ( .A(u5_mult_87_ab_38__35_), .B(
        u5_mult_87_CARRYB_37__35_), .CI(u5_mult_87_SUMB_37__36_), .CO(
        u5_mult_87_CARRYB_38__35_), .S(u5_mult_87_SUMB_38__35_) );
  FA_X1 u5_mult_87_S2_38_34 ( .A(u5_mult_87_ab_38__34_), .B(
        u5_mult_87_CARRYB_37__34_), .CI(u5_mult_87_SUMB_37__35_), .CO(
        u5_mult_87_CARRYB_38__34_), .S(u5_mult_87_SUMB_38__34_) );
  FA_X1 u5_mult_87_S2_38_33 ( .A(u5_mult_87_ab_38__33_), .B(
        u5_mult_87_CARRYB_37__33_), .CI(u5_mult_87_SUMB_37__34_), .CO(
        u5_mult_87_CARRYB_38__33_), .S(u5_mult_87_SUMB_38__33_) );
  FA_X1 u5_mult_87_S2_38_32 ( .A(u5_mult_87_ab_38__32_), .B(
        u5_mult_87_CARRYB_37__32_), .CI(u5_mult_87_SUMB_37__33_), .CO(
        u5_mult_87_CARRYB_38__32_), .S(u5_mult_87_SUMB_38__32_) );
  FA_X1 u5_mult_87_S2_38_31 ( .A(u5_mult_87_ab_38__31_), .B(
        u5_mult_87_CARRYB_37__31_), .CI(u5_mult_87_SUMB_37__32_), .CO(
        u5_mult_87_CARRYB_38__31_), .S(u5_mult_87_SUMB_38__31_) );
  FA_X1 u5_mult_87_S2_38_30 ( .A(u5_mult_87_ab_38__30_), .B(
        u5_mult_87_CARRYB_37__30_), .CI(u5_mult_87_SUMB_37__31_), .CO(
        u5_mult_87_CARRYB_38__30_), .S(u5_mult_87_SUMB_38__30_) );
  FA_X1 u5_mult_87_S2_38_29 ( .A(u5_mult_87_ab_38__29_), .B(
        u5_mult_87_CARRYB_37__29_), .CI(u5_mult_87_SUMB_37__30_), .CO(
        u5_mult_87_CARRYB_38__29_), .S(u5_mult_87_SUMB_38__29_) );
  FA_X1 u5_mult_87_S2_38_28 ( .A(u5_mult_87_ab_38__28_), .B(
        u5_mult_87_CARRYB_37__28_), .CI(u5_mult_87_SUMB_37__29_), .CO(
        u5_mult_87_CARRYB_38__28_), .S(u5_mult_87_SUMB_38__28_) );
  FA_X1 u5_mult_87_S2_38_27 ( .A(u5_mult_87_ab_38__27_), .B(
        u5_mult_87_CARRYB_37__27_), .CI(u5_mult_87_SUMB_37__28_), .CO(
        u5_mult_87_CARRYB_38__27_), .S(u5_mult_87_SUMB_38__27_) );
  FA_X1 u5_mult_87_S2_38_26 ( .A(u5_mult_87_ab_38__26_), .B(
        u5_mult_87_CARRYB_37__26_), .CI(u5_mult_87_SUMB_37__27_), .CO(
        u5_mult_87_CARRYB_38__26_), .S(u5_mult_87_SUMB_38__26_) );
  FA_X1 u5_mult_87_S2_38_25 ( .A(u5_mult_87_ab_38__25_), .B(
        u5_mult_87_CARRYB_37__25_), .CI(u5_mult_87_SUMB_37__26_), .CO(
        u5_mult_87_CARRYB_38__25_), .S(u5_mult_87_SUMB_38__25_) );
  FA_X1 u5_mult_87_S2_38_24 ( .A(u5_mult_87_ab_38__24_), .B(
        u5_mult_87_CARRYB_37__24_), .CI(u5_mult_87_SUMB_37__25_), .CO(
        u5_mult_87_CARRYB_38__24_), .S(u5_mult_87_SUMB_38__24_) );
  FA_X1 u5_mult_87_S2_38_23 ( .A(u5_mult_87_ab_38__23_), .B(
        u5_mult_87_CARRYB_37__23_), .CI(u5_mult_87_SUMB_37__24_), .CO(
        u5_mult_87_CARRYB_38__23_), .S(u5_mult_87_SUMB_38__23_) );
  FA_X1 u5_mult_87_S2_38_22 ( .A(u5_mult_87_ab_38__22_), .B(
        u5_mult_87_CARRYB_37__22_), .CI(u5_mult_87_SUMB_37__23_), .CO(
        u5_mult_87_CARRYB_38__22_), .S(u5_mult_87_SUMB_38__22_) );
  FA_X1 u5_mult_87_S2_38_21 ( .A(u5_mult_87_ab_38__21_), .B(
        u5_mult_87_CARRYB_37__21_), .CI(u5_mult_87_SUMB_37__22_), .CO(
        u5_mult_87_CARRYB_38__21_), .S(u5_mult_87_SUMB_38__21_) );
  FA_X1 u5_mult_87_S2_38_20 ( .A(u5_mult_87_ab_38__20_), .B(
        u5_mult_87_CARRYB_37__20_), .CI(u5_mult_87_SUMB_37__21_), .CO(
        u5_mult_87_CARRYB_38__20_), .S(u5_mult_87_SUMB_38__20_) );
  FA_X1 u5_mult_87_S2_38_19 ( .A(u5_mult_87_ab_38__19_), .B(
        u5_mult_87_CARRYB_37__19_), .CI(u5_mult_87_SUMB_37__20_), .CO(
        u5_mult_87_CARRYB_38__19_), .S(u5_mult_87_SUMB_38__19_) );
  FA_X1 u5_mult_87_S2_38_18 ( .A(u5_mult_87_ab_38__18_), .B(
        u5_mult_87_CARRYB_37__18_), .CI(u5_mult_87_SUMB_37__19_), .CO(
        u5_mult_87_CARRYB_38__18_), .S(u5_mult_87_SUMB_38__18_) );
  FA_X1 u5_mult_87_S2_38_17 ( .A(u5_mult_87_ab_38__17_), .B(
        u5_mult_87_CARRYB_37__17_), .CI(u5_mult_87_SUMB_37__18_), .CO(
        u5_mult_87_CARRYB_38__17_), .S(u5_mult_87_SUMB_38__17_) );
  FA_X1 u5_mult_87_S2_38_16 ( .A(u5_mult_87_ab_38__16_), .B(
        u5_mult_87_CARRYB_37__16_), .CI(u5_mult_87_SUMB_37__17_), .CO(
        u5_mult_87_CARRYB_38__16_), .S(u5_mult_87_SUMB_38__16_) );
  FA_X1 u5_mult_87_S2_38_15 ( .A(u5_mult_87_ab_38__15_), .B(
        u5_mult_87_CARRYB_37__15_), .CI(u5_mult_87_SUMB_37__16_), .CO(
        u5_mult_87_CARRYB_38__15_), .S(u5_mult_87_SUMB_38__15_) );
  FA_X1 u5_mult_87_S2_38_14 ( .A(u5_mult_87_ab_38__14_), .B(
        u5_mult_87_CARRYB_37__14_), .CI(u5_mult_87_SUMB_37__15_), .CO(
        u5_mult_87_CARRYB_38__14_), .S(u5_mult_87_SUMB_38__14_) );
  FA_X1 u5_mult_87_S2_38_13 ( .A(u5_mult_87_ab_38__13_), .B(
        u5_mult_87_CARRYB_37__13_), .CI(u5_mult_87_SUMB_37__14_), .CO(
        u5_mult_87_CARRYB_38__13_), .S(u5_mult_87_SUMB_38__13_) );
  FA_X1 u5_mult_87_S2_38_12 ( .A(u5_mult_87_ab_38__12_), .B(
        u5_mult_87_CARRYB_37__12_), .CI(u5_mult_87_SUMB_37__13_), .CO(
        u5_mult_87_CARRYB_38__12_), .S(u5_mult_87_SUMB_38__12_) );
  FA_X1 u5_mult_87_S2_38_11 ( .A(u5_mult_87_ab_38__11_), .B(
        u5_mult_87_CARRYB_37__11_), .CI(u5_mult_87_SUMB_37__12_), .CO(
        u5_mult_87_CARRYB_38__11_), .S(u5_mult_87_SUMB_38__11_) );
  FA_X1 u5_mult_87_S2_38_10 ( .A(u5_mult_87_ab_38__10_), .B(
        u5_mult_87_CARRYB_37__10_), .CI(u5_mult_87_SUMB_37__11_), .CO(
        u5_mult_87_CARRYB_38__10_), .S(u5_mult_87_SUMB_38__10_) );
  FA_X1 u5_mult_87_S2_38_9 ( .A(u5_mult_87_ab_38__9_), .B(
        u5_mult_87_CARRYB_37__9_), .CI(u5_mult_87_SUMB_37__10_), .CO(
        u5_mult_87_CARRYB_38__9_), .S(u5_mult_87_SUMB_38__9_) );
  FA_X1 u5_mult_87_S2_38_8 ( .A(u5_mult_87_ab_38__8_), .B(
        u5_mult_87_CARRYB_37__8_), .CI(u5_mult_87_SUMB_37__9_), .CO(
        u5_mult_87_CARRYB_38__8_), .S(u5_mult_87_SUMB_38__8_) );
  FA_X1 u5_mult_87_S2_38_7 ( .A(u5_mult_87_ab_38__7_), .B(
        u5_mult_87_CARRYB_37__7_), .CI(u5_mult_87_SUMB_37__8_), .CO(
        u5_mult_87_CARRYB_38__7_), .S(u5_mult_87_SUMB_38__7_) );
  FA_X1 u5_mult_87_S2_38_6 ( .A(u5_mult_87_ab_38__6_), .B(
        u5_mult_87_CARRYB_37__6_), .CI(u5_mult_87_SUMB_37__7_), .CO(
        u5_mult_87_CARRYB_38__6_), .S(u5_mult_87_SUMB_38__6_) );
  FA_X1 u5_mult_87_S2_38_5 ( .A(u5_mult_87_ab_38__5_), .B(
        u5_mult_87_CARRYB_37__5_), .CI(u5_mult_87_SUMB_37__6_), .CO(
        u5_mult_87_CARRYB_38__5_), .S(u5_mult_87_SUMB_38__5_) );
  FA_X1 u5_mult_87_S2_38_4 ( .A(u5_mult_87_ab_38__4_), .B(
        u5_mult_87_CARRYB_37__4_), .CI(u5_mult_87_SUMB_37__5_), .CO(
        u5_mult_87_CARRYB_38__4_), .S(u5_mult_87_SUMB_38__4_) );
  FA_X1 u5_mult_87_S2_38_3 ( .A(u5_mult_87_ab_38__3_), .B(
        u5_mult_87_CARRYB_37__3_), .CI(u5_mult_87_SUMB_37__4_), .CO(
        u5_mult_87_CARRYB_38__3_), .S(u5_mult_87_SUMB_38__3_) );
  FA_X1 u5_mult_87_S2_38_2 ( .A(u5_mult_87_ab_38__2_), .B(
        u5_mult_87_CARRYB_37__2_), .CI(u5_mult_87_SUMB_37__3_), .CO(
        u5_mult_87_CARRYB_38__2_), .S(u5_mult_87_SUMB_38__2_) );
  FA_X1 u5_mult_87_S2_38_1 ( .A(u5_mult_87_ab_38__1_), .B(
        u5_mult_87_CARRYB_37__1_), .CI(u5_mult_87_SUMB_37__2_), .CO(
        u5_mult_87_CARRYB_38__1_), .S(u5_mult_87_SUMB_38__1_) );
  FA_X1 u5_mult_87_S1_38_0 ( .A(u5_mult_87_ab_38__0_), .B(
        u5_mult_87_CARRYB_37__0_), .CI(u5_mult_87_SUMB_37__1_), .CO(
        u5_mult_87_CARRYB_38__0_), .S(u5_N38) );
  FA_X1 u5_mult_87_S3_39_51 ( .A(u5_mult_87_ab_39__51_), .B(
        u5_mult_87_CARRYB_38__51_), .CI(u5_mult_87_ab_38__52_), .CO(
        u5_mult_87_CARRYB_39__51_), .S(u5_mult_87_SUMB_39__51_) );
  FA_X1 u5_mult_87_S2_39_50 ( .A(u5_mult_87_ab_39__50_), .B(
        u5_mult_87_CARRYB_38__50_), .CI(u5_mult_87_SUMB_38__51_), .CO(
        u5_mult_87_CARRYB_39__50_), .S(u5_mult_87_SUMB_39__50_) );
  FA_X1 u5_mult_87_S2_39_49 ( .A(u5_mult_87_ab_39__49_), .B(
        u5_mult_87_CARRYB_38__49_), .CI(u5_mult_87_SUMB_38__50_), .CO(
        u5_mult_87_CARRYB_39__49_), .S(u5_mult_87_SUMB_39__49_) );
  FA_X1 u5_mult_87_S2_39_48 ( .A(u5_mult_87_ab_39__48_), .B(
        u5_mult_87_CARRYB_38__48_), .CI(u5_mult_87_SUMB_38__49_), .CO(
        u5_mult_87_CARRYB_39__48_), .S(u5_mult_87_SUMB_39__48_) );
  FA_X1 u5_mult_87_S2_39_47 ( .A(u5_mult_87_ab_39__47_), .B(
        u5_mult_87_CARRYB_38__47_), .CI(u5_mult_87_SUMB_38__48_), .CO(
        u5_mult_87_CARRYB_39__47_), .S(u5_mult_87_SUMB_39__47_) );
  FA_X1 u5_mult_87_S2_39_46 ( .A(u5_mult_87_ab_39__46_), .B(
        u5_mult_87_CARRYB_38__46_), .CI(u5_mult_87_SUMB_38__47_), .CO(
        u5_mult_87_CARRYB_39__46_), .S(u5_mult_87_SUMB_39__46_) );
  FA_X1 u5_mult_87_S2_39_45 ( .A(u5_mult_87_ab_39__45_), .B(
        u5_mult_87_CARRYB_38__45_), .CI(u5_mult_87_SUMB_38__46_), .CO(
        u5_mult_87_CARRYB_39__45_), .S(u5_mult_87_SUMB_39__45_) );
  FA_X1 u5_mult_87_S2_39_44 ( .A(u5_mult_87_ab_39__44_), .B(
        u5_mult_87_CARRYB_38__44_), .CI(u5_mult_87_SUMB_38__45_), .CO(
        u5_mult_87_CARRYB_39__44_), .S(u5_mult_87_SUMB_39__44_) );
  FA_X1 u5_mult_87_S2_39_43 ( .A(u5_mult_87_ab_39__43_), .B(
        u5_mult_87_CARRYB_38__43_), .CI(u5_mult_87_SUMB_38__44_), .CO(
        u5_mult_87_CARRYB_39__43_), .S(u5_mult_87_SUMB_39__43_) );
  FA_X1 u5_mult_87_S2_39_42 ( .A(u5_mult_87_ab_39__42_), .B(
        u5_mult_87_CARRYB_38__42_), .CI(u5_mult_87_SUMB_38__43_), .CO(
        u5_mult_87_CARRYB_39__42_), .S(u5_mult_87_SUMB_39__42_) );
  FA_X1 u5_mult_87_S2_39_41 ( .A(u5_mult_87_ab_39__41_), .B(
        u5_mult_87_CARRYB_38__41_), .CI(u5_mult_87_SUMB_38__42_), .CO(
        u5_mult_87_CARRYB_39__41_), .S(u5_mult_87_SUMB_39__41_) );
  FA_X1 u5_mult_87_S2_39_40 ( .A(u5_mult_87_ab_39__40_), .B(
        u5_mult_87_CARRYB_38__40_), .CI(u5_mult_87_SUMB_38__41_), .CO(
        u5_mult_87_CARRYB_39__40_), .S(u5_mult_87_SUMB_39__40_) );
  FA_X1 u5_mult_87_S2_39_39 ( .A(u5_mult_87_ab_39__39_), .B(
        u5_mult_87_CARRYB_38__39_), .CI(u5_mult_87_SUMB_38__40_), .CO(
        u5_mult_87_CARRYB_39__39_), .S(u5_mult_87_SUMB_39__39_) );
  FA_X1 u5_mult_87_S2_39_38 ( .A(u5_mult_87_ab_39__38_), .B(
        u5_mult_87_CARRYB_38__38_), .CI(u5_mult_87_SUMB_38__39_), .CO(
        u5_mult_87_CARRYB_39__38_), .S(u5_mult_87_SUMB_39__38_) );
  FA_X1 u5_mult_87_S2_39_37 ( .A(u5_mult_87_ab_39__37_), .B(
        u5_mult_87_CARRYB_38__37_), .CI(u5_mult_87_SUMB_38__38_), .CO(
        u5_mult_87_CARRYB_39__37_), .S(u5_mult_87_SUMB_39__37_) );
  FA_X1 u5_mult_87_S2_39_36 ( .A(u5_mult_87_ab_39__36_), .B(
        u5_mult_87_CARRYB_38__36_), .CI(u5_mult_87_SUMB_38__37_), .CO(
        u5_mult_87_CARRYB_39__36_), .S(u5_mult_87_SUMB_39__36_) );
  FA_X1 u5_mult_87_S2_39_35 ( .A(u5_mult_87_ab_39__35_), .B(
        u5_mult_87_CARRYB_38__35_), .CI(u5_mult_87_SUMB_38__36_), .CO(
        u5_mult_87_CARRYB_39__35_), .S(u5_mult_87_SUMB_39__35_) );
  FA_X1 u5_mult_87_S2_39_34 ( .A(u5_mult_87_ab_39__34_), .B(
        u5_mult_87_CARRYB_38__34_), .CI(u5_mult_87_SUMB_38__35_), .CO(
        u5_mult_87_CARRYB_39__34_), .S(u5_mult_87_SUMB_39__34_) );
  FA_X1 u5_mult_87_S2_39_33 ( .A(u5_mult_87_ab_39__33_), .B(
        u5_mult_87_CARRYB_38__33_), .CI(u5_mult_87_SUMB_38__34_), .CO(
        u5_mult_87_CARRYB_39__33_), .S(u5_mult_87_SUMB_39__33_) );
  FA_X1 u5_mult_87_S2_39_32 ( .A(u5_mult_87_ab_39__32_), .B(
        u5_mult_87_CARRYB_38__32_), .CI(u5_mult_87_SUMB_38__33_), .CO(
        u5_mult_87_CARRYB_39__32_), .S(u5_mult_87_SUMB_39__32_) );
  FA_X1 u5_mult_87_S2_39_31 ( .A(u5_mult_87_ab_39__31_), .B(
        u5_mult_87_CARRYB_38__31_), .CI(u5_mult_87_SUMB_38__32_), .CO(
        u5_mult_87_CARRYB_39__31_), .S(u5_mult_87_SUMB_39__31_) );
  FA_X1 u5_mult_87_S2_39_30 ( .A(u5_mult_87_ab_39__30_), .B(
        u5_mult_87_CARRYB_38__30_), .CI(u5_mult_87_SUMB_38__31_), .CO(
        u5_mult_87_CARRYB_39__30_), .S(u5_mult_87_SUMB_39__30_) );
  FA_X1 u5_mult_87_S2_39_29 ( .A(u5_mult_87_ab_39__29_), .B(
        u5_mult_87_CARRYB_38__29_), .CI(u5_mult_87_SUMB_38__30_), .CO(
        u5_mult_87_CARRYB_39__29_), .S(u5_mult_87_SUMB_39__29_) );
  FA_X1 u5_mult_87_S2_39_28 ( .A(u5_mult_87_ab_39__28_), .B(
        u5_mult_87_CARRYB_38__28_), .CI(u5_mult_87_SUMB_38__29_), .CO(
        u5_mult_87_CARRYB_39__28_), .S(u5_mult_87_SUMB_39__28_) );
  FA_X1 u5_mult_87_S2_39_27 ( .A(u5_mult_87_ab_39__27_), .B(
        u5_mult_87_CARRYB_38__27_), .CI(u5_mult_87_SUMB_38__28_), .CO(
        u5_mult_87_CARRYB_39__27_), .S(u5_mult_87_SUMB_39__27_) );
  FA_X1 u5_mult_87_S2_39_26 ( .A(u5_mult_87_ab_39__26_), .B(
        u5_mult_87_CARRYB_38__26_), .CI(u5_mult_87_SUMB_38__27_), .CO(
        u5_mult_87_CARRYB_39__26_), .S(u5_mult_87_SUMB_39__26_) );
  FA_X1 u5_mult_87_S2_39_25 ( .A(u5_mult_87_ab_39__25_), .B(
        u5_mult_87_CARRYB_38__25_), .CI(u5_mult_87_SUMB_38__26_), .CO(
        u5_mult_87_CARRYB_39__25_), .S(u5_mult_87_SUMB_39__25_) );
  FA_X1 u5_mult_87_S2_39_24 ( .A(u5_mult_87_ab_39__24_), .B(
        u5_mult_87_CARRYB_38__24_), .CI(u5_mult_87_SUMB_38__25_), .CO(
        u5_mult_87_CARRYB_39__24_), .S(u5_mult_87_SUMB_39__24_) );
  FA_X1 u5_mult_87_S2_39_23 ( .A(u5_mult_87_ab_39__23_), .B(
        u5_mult_87_CARRYB_38__23_), .CI(u5_mult_87_SUMB_38__24_), .CO(
        u5_mult_87_CARRYB_39__23_), .S(u5_mult_87_SUMB_39__23_) );
  FA_X1 u5_mult_87_S2_39_22 ( .A(u5_mult_87_ab_39__22_), .B(
        u5_mult_87_CARRYB_38__22_), .CI(u5_mult_87_SUMB_38__23_), .CO(
        u5_mult_87_CARRYB_39__22_), .S(u5_mult_87_SUMB_39__22_) );
  FA_X1 u5_mult_87_S2_39_21 ( .A(u5_mult_87_ab_39__21_), .B(
        u5_mult_87_CARRYB_38__21_), .CI(u5_mult_87_SUMB_38__22_), .CO(
        u5_mult_87_CARRYB_39__21_), .S(u5_mult_87_SUMB_39__21_) );
  FA_X1 u5_mult_87_S2_39_20 ( .A(u5_mult_87_ab_39__20_), .B(
        u5_mult_87_CARRYB_38__20_), .CI(u5_mult_87_SUMB_38__21_), .CO(
        u5_mult_87_CARRYB_39__20_), .S(u5_mult_87_SUMB_39__20_) );
  FA_X1 u5_mult_87_S2_39_19 ( .A(u5_mult_87_ab_39__19_), .B(
        u5_mult_87_CARRYB_38__19_), .CI(u5_mult_87_SUMB_38__20_), .CO(
        u5_mult_87_CARRYB_39__19_), .S(u5_mult_87_SUMB_39__19_) );
  FA_X1 u5_mult_87_S2_39_18 ( .A(u5_mult_87_ab_39__18_), .B(
        u5_mult_87_CARRYB_38__18_), .CI(u5_mult_87_SUMB_38__19_), .CO(
        u5_mult_87_CARRYB_39__18_), .S(u5_mult_87_SUMB_39__18_) );
  FA_X1 u5_mult_87_S2_39_17 ( .A(u5_mult_87_ab_39__17_), .B(
        u5_mult_87_CARRYB_38__17_), .CI(u5_mult_87_SUMB_38__18_), .CO(
        u5_mult_87_CARRYB_39__17_), .S(u5_mult_87_SUMB_39__17_) );
  FA_X1 u5_mult_87_S2_39_16 ( .A(u5_mult_87_ab_39__16_), .B(
        u5_mult_87_CARRYB_38__16_), .CI(u5_mult_87_SUMB_38__17_), .CO(
        u5_mult_87_CARRYB_39__16_), .S(u5_mult_87_SUMB_39__16_) );
  FA_X1 u5_mult_87_S2_39_15 ( .A(u5_mult_87_ab_39__15_), .B(
        u5_mult_87_CARRYB_38__15_), .CI(u5_mult_87_SUMB_38__16_), .CO(
        u5_mult_87_CARRYB_39__15_), .S(u5_mult_87_SUMB_39__15_) );
  FA_X1 u5_mult_87_S2_39_14 ( .A(u5_mult_87_ab_39__14_), .B(
        u5_mult_87_CARRYB_38__14_), .CI(u5_mult_87_SUMB_38__15_), .CO(
        u5_mult_87_CARRYB_39__14_), .S(u5_mult_87_SUMB_39__14_) );
  FA_X1 u5_mult_87_S2_39_13 ( .A(u5_mult_87_ab_39__13_), .B(
        u5_mult_87_CARRYB_38__13_), .CI(u5_mult_87_SUMB_38__14_), .CO(
        u5_mult_87_CARRYB_39__13_), .S(u5_mult_87_SUMB_39__13_) );
  FA_X1 u5_mult_87_S2_39_12 ( .A(u5_mult_87_ab_39__12_), .B(
        u5_mult_87_CARRYB_38__12_), .CI(u5_mult_87_SUMB_38__13_), .CO(
        u5_mult_87_CARRYB_39__12_), .S(u5_mult_87_SUMB_39__12_) );
  FA_X1 u5_mult_87_S2_39_11 ( .A(u5_mult_87_ab_39__11_), .B(
        u5_mult_87_CARRYB_38__11_), .CI(u5_mult_87_SUMB_38__12_), .CO(
        u5_mult_87_CARRYB_39__11_), .S(u5_mult_87_SUMB_39__11_) );
  FA_X1 u5_mult_87_S2_39_10 ( .A(u5_mult_87_ab_39__10_), .B(
        u5_mult_87_CARRYB_38__10_), .CI(u5_mult_87_SUMB_38__11_), .CO(
        u5_mult_87_CARRYB_39__10_), .S(u5_mult_87_SUMB_39__10_) );
  FA_X1 u5_mult_87_S2_39_9 ( .A(u5_mult_87_ab_39__9_), .B(
        u5_mult_87_CARRYB_38__9_), .CI(u5_mult_87_SUMB_38__10_), .CO(
        u5_mult_87_CARRYB_39__9_), .S(u5_mult_87_SUMB_39__9_) );
  FA_X1 u5_mult_87_S2_39_8 ( .A(u5_mult_87_ab_39__8_), .B(
        u5_mult_87_CARRYB_38__8_), .CI(u5_mult_87_SUMB_38__9_), .CO(
        u5_mult_87_CARRYB_39__8_), .S(u5_mult_87_SUMB_39__8_) );
  FA_X1 u5_mult_87_S2_39_7 ( .A(u5_mult_87_ab_39__7_), .B(
        u5_mult_87_CARRYB_38__7_), .CI(u5_mult_87_SUMB_38__8_), .CO(
        u5_mult_87_CARRYB_39__7_), .S(u5_mult_87_SUMB_39__7_) );
  FA_X1 u5_mult_87_S2_39_6 ( .A(u5_mult_87_ab_39__6_), .B(
        u5_mult_87_CARRYB_38__6_), .CI(u5_mult_87_SUMB_38__7_), .CO(
        u5_mult_87_CARRYB_39__6_), .S(u5_mult_87_SUMB_39__6_) );
  FA_X1 u5_mult_87_S2_39_5 ( .A(u5_mult_87_ab_39__5_), .B(
        u5_mult_87_CARRYB_38__5_), .CI(u5_mult_87_SUMB_38__6_), .CO(
        u5_mult_87_CARRYB_39__5_), .S(u5_mult_87_SUMB_39__5_) );
  FA_X1 u5_mult_87_S2_39_4 ( .A(u5_mult_87_ab_39__4_), .B(
        u5_mult_87_CARRYB_38__4_), .CI(u5_mult_87_SUMB_38__5_), .CO(
        u5_mult_87_CARRYB_39__4_), .S(u5_mult_87_SUMB_39__4_) );
  FA_X1 u5_mult_87_S2_39_3 ( .A(u5_mult_87_ab_39__3_), .B(
        u5_mult_87_CARRYB_38__3_), .CI(u5_mult_87_SUMB_38__4_), .CO(
        u5_mult_87_CARRYB_39__3_), .S(u5_mult_87_SUMB_39__3_) );
  FA_X1 u5_mult_87_S2_39_2 ( .A(u5_mult_87_ab_39__2_), .B(
        u5_mult_87_CARRYB_38__2_), .CI(u5_mult_87_SUMB_38__3_), .CO(
        u5_mult_87_CARRYB_39__2_), .S(u5_mult_87_SUMB_39__2_) );
  FA_X1 u5_mult_87_S2_39_1 ( .A(u5_mult_87_ab_39__1_), .B(
        u5_mult_87_CARRYB_38__1_), .CI(u5_mult_87_SUMB_38__2_), .CO(
        u5_mult_87_CARRYB_39__1_), .S(u5_mult_87_SUMB_39__1_) );
  FA_X1 u5_mult_87_S1_39_0 ( .A(u5_mult_87_ab_39__0_), .B(
        u5_mult_87_CARRYB_38__0_), .CI(u5_mult_87_SUMB_38__1_), .CO(
        u5_mult_87_CARRYB_39__0_), .S(u5_N39) );
  FA_X1 u5_mult_87_S3_40_51 ( .A(u5_mult_87_ab_40__51_), .B(
        u5_mult_87_CARRYB_39__51_), .CI(u5_mult_87_ab_39__52_), .CO(
        u5_mult_87_CARRYB_40__51_), .S(u5_mult_87_SUMB_40__51_) );
  FA_X1 u5_mult_87_S2_40_50 ( .A(u5_mult_87_ab_40__50_), .B(
        u5_mult_87_CARRYB_39__50_), .CI(u5_mult_87_SUMB_39__51_), .CO(
        u5_mult_87_CARRYB_40__50_), .S(u5_mult_87_SUMB_40__50_) );
  FA_X1 u5_mult_87_S2_40_49 ( .A(u5_mult_87_ab_40__49_), .B(
        u5_mult_87_CARRYB_39__49_), .CI(u5_mult_87_SUMB_39__50_), .CO(
        u5_mult_87_CARRYB_40__49_), .S(u5_mult_87_SUMB_40__49_) );
  FA_X1 u5_mult_87_S2_40_48 ( .A(u5_mult_87_ab_40__48_), .B(
        u5_mult_87_CARRYB_39__48_), .CI(u5_mult_87_SUMB_39__49_), .CO(
        u5_mult_87_CARRYB_40__48_), .S(u5_mult_87_SUMB_40__48_) );
  FA_X1 u5_mult_87_S2_40_47 ( .A(u5_mult_87_ab_40__47_), .B(
        u5_mult_87_CARRYB_39__47_), .CI(u5_mult_87_SUMB_39__48_), .CO(
        u5_mult_87_CARRYB_40__47_), .S(u5_mult_87_SUMB_40__47_) );
  FA_X1 u5_mult_87_S2_40_46 ( .A(u5_mult_87_ab_40__46_), .B(
        u5_mult_87_CARRYB_39__46_), .CI(u5_mult_87_SUMB_39__47_), .CO(
        u5_mult_87_CARRYB_40__46_), .S(u5_mult_87_SUMB_40__46_) );
  FA_X1 u5_mult_87_S2_40_45 ( .A(u5_mult_87_ab_40__45_), .B(
        u5_mult_87_CARRYB_39__45_), .CI(u5_mult_87_SUMB_39__46_), .CO(
        u5_mult_87_CARRYB_40__45_), .S(u5_mult_87_SUMB_40__45_) );
  FA_X1 u5_mult_87_S2_40_44 ( .A(u5_mult_87_ab_40__44_), .B(
        u5_mult_87_CARRYB_39__44_), .CI(u5_mult_87_SUMB_39__45_), .CO(
        u5_mult_87_CARRYB_40__44_), .S(u5_mult_87_SUMB_40__44_) );
  FA_X1 u5_mult_87_S2_40_43 ( .A(u5_mult_87_ab_40__43_), .B(
        u5_mult_87_CARRYB_39__43_), .CI(u5_mult_87_SUMB_39__44_), .CO(
        u5_mult_87_CARRYB_40__43_), .S(u5_mult_87_SUMB_40__43_) );
  FA_X1 u5_mult_87_S2_40_42 ( .A(u5_mult_87_ab_40__42_), .B(
        u5_mult_87_CARRYB_39__42_), .CI(u5_mult_87_SUMB_39__43_), .CO(
        u5_mult_87_CARRYB_40__42_), .S(u5_mult_87_SUMB_40__42_) );
  FA_X1 u5_mult_87_S2_40_41 ( .A(u5_mult_87_ab_40__41_), .B(
        u5_mult_87_CARRYB_39__41_), .CI(u5_mult_87_SUMB_39__42_), .CO(
        u5_mult_87_CARRYB_40__41_), .S(u5_mult_87_SUMB_40__41_) );
  FA_X1 u5_mult_87_S2_40_40 ( .A(u5_mult_87_ab_40__40_), .B(
        u5_mult_87_CARRYB_39__40_), .CI(u5_mult_87_SUMB_39__41_), .CO(
        u5_mult_87_CARRYB_40__40_), .S(u5_mult_87_SUMB_40__40_) );
  FA_X1 u5_mult_87_S2_40_39 ( .A(u5_mult_87_ab_40__39_), .B(
        u5_mult_87_CARRYB_39__39_), .CI(u5_mult_87_SUMB_39__40_), .CO(
        u5_mult_87_CARRYB_40__39_), .S(u5_mult_87_SUMB_40__39_) );
  FA_X1 u5_mult_87_S2_40_38 ( .A(u5_mult_87_ab_40__38_), .B(
        u5_mult_87_CARRYB_39__38_), .CI(u5_mult_87_SUMB_39__39_), .CO(
        u5_mult_87_CARRYB_40__38_), .S(u5_mult_87_SUMB_40__38_) );
  FA_X1 u5_mult_87_S2_40_37 ( .A(u5_mult_87_ab_40__37_), .B(
        u5_mult_87_CARRYB_39__37_), .CI(u5_mult_87_SUMB_39__38_), .CO(
        u5_mult_87_CARRYB_40__37_), .S(u5_mult_87_SUMB_40__37_) );
  FA_X1 u5_mult_87_S2_40_36 ( .A(u5_mult_87_ab_40__36_), .B(
        u5_mult_87_CARRYB_39__36_), .CI(u5_mult_87_SUMB_39__37_), .CO(
        u5_mult_87_CARRYB_40__36_), .S(u5_mult_87_SUMB_40__36_) );
  FA_X1 u5_mult_87_S2_40_35 ( .A(u5_mult_87_ab_40__35_), .B(
        u5_mult_87_CARRYB_39__35_), .CI(u5_mult_87_SUMB_39__36_), .CO(
        u5_mult_87_CARRYB_40__35_), .S(u5_mult_87_SUMB_40__35_) );
  FA_X1 u5_mult_87_S2_40_34 ( .A(u5_mult_87_ab_40__34_), .B(
        u5_mult_87_CARRYB_39__34_), .CI(u5_mult_87_SUMB_39__35_), .CO(
        u5_mult_87_CARRYB_40__34_), .S(u5_mult_87_SUMB_40__34_) );
  FA_X1 u5_mult_87_S2_40_33 ( .A(u5_mult_87_ab_40__33_), .B(
        u5_mult_87_CARRYB_39__33_), .CI(u5_mult_87_SUMB_39__34_), .CO(
        u5_mult_87_CARRYB_40__33_), .S(u5_mult_87_SUMB_40__33_) );
  FA_X1 u5_mult_87_S2_40_32 ( .A(u5_mult_87_ab_40__32_), .B(
        u5_mult_87_CARRYB_39__32_), .CI(u5_mult_87_SUMB_39__33_), .CO(
        u5_mult_87_CARRYB_40__32_), .S(u5_mult_87_SUMB_40__32_) );
  FA_X1 u5_mult_87_S2_40_31 ( .A(u5_mult_87_ab_40__31_), .B(
        u5_mult_87_CARRYB_39__31_), .CI(u5_mult_87_SUMB_39__32_), .CO(
        u5_mult_87_CARRYB_40__31_), .S(u5_mult_87_SUMB_40__31_) );
  FA_X1 u5_mult_87_S2_40_30 ( .A(u5_mult_87_ab_40__30_), .B(
        u5_mult_87_CARRYB_39__30_), .CI(u5_mult_87_SUMB_39__31_), .CO(
        u5_mult_87_CARRYB_40__30_), .S(u5_mult_87_SUMB_40__30_) );
  FA_X1 u5_mult_87_S2_40_29 ( .A(u5_mult_87_ab_40__29_), .B(
        u5_mult_87_CARRYB_39__29_), .CI(u5_mult_87_SUMB_39__30_), .CO(
        u5_mult_87_CARRYB_40__29_), .S(u5_mult_87_SUMB_40__29_) );
  FA_X1 u5_mult_87_S2_40_28 ( .A(u5_mult_87_ab_40__28_), .B(
        u5_mult_87_CARRYB_39__28_), .CI(u5_mult_87_SUMB_39__29_), .CO(
        u5_mult_87_CARRYB_40__28_), .S(u5_mult_87_SUMB_40__28_) );
  FA_X1 u5_mult_87_S2_40_27 ( .A(u5_mult_87_ab_40__27_), .B(
        u5_mult_87_CARRYB_39__27_), .CI(u5_mult_87_SUMB_39__28_), .CO(
        u5_mult_87_CARRYB_40__27_), .S(u5_mult_87_SUMB_40__27_) );
  FA_X1 u5_mult_87_S2_40_26 ( .A(u5_mult_87_ab_40__26_), .B(
        u5_mult_87_CARRYB_39__26_), .CI(u5_mult_87_SUMB_39__27_), .CO(
        u5_mult_87_CARRYB_40__26_), .S(u5_mult_87_SUMB_40__26_) );
  FA_X1 u5_mult_87_S2_40_25 ( .A(u5_mult_87_ab_40__25_), .B(
        u5_mult_87_CARRYB_39__25_), .CI(u5_mult_87_SUMB_39__26_), .CO(
        u5_mult_87_CARRYB_40__25_), .S(u5_mult_87_SUMB_40__25_) );
  FA_X1 u5_mult_87_S2_40_24 ( .A(u5_mult_87_ab_40__24_), .B(
        u5_mult_87_CARRYB_39__24_), .CI(u5_mult_87_SUMB_39__25_), .CO(
        u5_mult_87_CARRYB_40__24_), .S(u5_mult_87_SUMB_40__24_) );
  FA_X1 u5_mult_87_S2_40_23 ( .A(u5_mult_87_ab_40__23_), .B(
        u5_mult_87_CARRYB_39__23_), .CI(u5_mult_87_SUMB_39__24_), .CO(
        u5_mult_87_CARRYB_40__23_), .S(u5_mult_87_SUMB_40__23_) );
  FA_X1 u5_mult_87_S2_40_22 ( .A(u5_mult_87_ab_40__22_), .B(
        u5_mult_87_CARRYB_39__22_), .CI(u5_mult_87_SUMB_39__23_), .CO(
        u5_mult_87_CARRYB_40__22_), .S(u5_mult_87_SUMB_40__22_) );
  FA_X1 u5_mult_87_S2_40_21 ( .A(u5_mult_87_ab_40__21_), .B(
        u5_mult_87_CARRYB_39__21_), .CI(u5_mult_87_SUMB_39__22_), .CO(
        u5_mult_87_CARRYB_40__21_), .S(u5_mult_87_SUMB_40__21_) );
  FA_X1 u5_mult_87_S2_40_20 ( .A(u5_mult_87_ab_40__20_), .B(
        u5_mult_87_CARRYB_39__20_), .CI(u5_mult_87_SUMB_39__21_), .CO(
        u5_mult_87_CARRYB_40__20_), .S(u5_mult_87_SUMB_40__20_) );
  FA_X1 u5_mult_87_S2_40_19 ( .A(u5_mult_87_ab_40__19_), .B(
        u5_mult_87_CARRYB_39__19_), .CI(u5_mult_87_SUMB_39__20_), .CO(
        u5_mult_87_CARRYB_40__19_), .S(u5_mult_87_SUMB_40__19_) );
  FA_X1 u5_mult_87_S2_40_18 ( .A(u5_mult_87_ab_40__18_), .B(
        u5_mult_87_CARRYB_39__18_), .CI(u5_mult_87_SUMB_39__19_), .CO(
        u5_mult_87_CARRYB_40__18_), .S(u5_mult_87_SUMB_40__18_) );
  FA_X1 u5_mult_87_S2_40_17 ( .A(u5_mult_87_ab_40__17_), .B(
        u5_mult_87_CARRYB_39__17_), .CI(u5_mult_87_SUMB_39__18_), .CO(
        u5_mult_87_CARRYB_40__17_), .S(u5_mult_87_SUMB_40__17_) );
  FA_X1 u5_mult_87_S2_40_16 ( .A(u5_mult_87_ab_40__16_), .B(
        u5_mult_87_CARRYB_39__16_), .CI(u5_mult_87_SUMB_39__17_), .CO(
        u5_mult_87_CARRYB_40__16_), .S(u5_mult_87_SUMB_40__16_) );
  FA_X1 u5_mult_87_S2_40_15 ( .A(u5_mult_87_ab_40__15_), .B(
        u5_mult_87_CARRYB_39__15_), .CI(u5_mult_87_SUMB_39__16_), .CO(
        u5_mult_87_CARRYB_40__15_), .S(u5_mult_87_SUMB_40__15_) );
  FA_X1 u5_mult_87_S2_40_14 ( .A(u5_mult_87_ab_40__14_), .B(
        u5_mult_87_CARRYB_39__14_), .CI(u5_mult_87_SUMB_39__15_), .CO(
        u5_mult_87_CARRYB_40__14_), .S(u5_mult_87_SUMB_40__14_) );
  FA_X1 u5_mult_87_S2_40_13 ( .A(u5_mult_87_ab_40__13_), .B(
        u5_mult_87_CARRYB_39__13_), .CI(u5_mult_87_SUMB_39__14_), .CO(
        u5_mult_87_CARRYB_40__13_), .S(u5_mult_87_SUMB_40__13_) );
  FA_X1 u5_mult_87_S2_40_12 ( .A(u5_mult_87_ab_40__12_), .B(
        u5_mult_87_CARRYB_39__12_), .CI(u5_mult_87_SUMB_39__13_), .CO(
        u5_mult_87_CARRYB_40__12_), .S(u5_mult_87_SUMB_40__12_) );
  FA_X1 u5_mult_87_S2_40_11 ( .A(u5_mult_87_ab_40__11_), .B(
        u5_mult_87_CARRYB_39__11_), .CI(u5_mult_87_SUMB_39__12_), .CO(
        u5_mult_87_CARRYB_40__11_), .S(u5_mult_87_SUMB_40__11_) );
  FA_X1 u5_mult_87_S2_40_10 ( .A(u5_mult_87_ab_40__10_), .B(
        u5_mult_87_CARRYB_39__10_), .CI(u5_mult_87_SUMB_39__11_), .CO(
        u5_mult_87_CARRYB_40__10_), .S(u5_mult_87_SUMB_40__10_) );
  FA_X1 u5_mult_87_S2_40_9 ( .A(u5_mult_87_ab_40__9_), .B(
        u5_mult_87_CARRYB_39__9_), .CI(u5_mult_87_SUMB_39__10_), .CO(
        u5_mult_87_CARRYB_40__9_), .S(u5_mult_87_SUMB_40__9_) );
  FA_X1 u5_mult_87_S2_40_8 ( .A(u5_mult_87_ab_40__8_), .B(
        u5_mult_87_CARRYB_39__8_), .CI(u5_mult_87_SUMB_39__9_), .CO(
        u5_mult_87_CARRYB_40__8_), .S(u5_mult_87_SUMB_40__8_) );
  FA_X1 u5_mult_87_S2_40_7 ( .A(u5_mult_87_ab_40__7_), .B(
        u5_mult_87_CARRYB_39__7_), .CI(u5_mult_87_SUMB_39__8_), .CO(
        u5_mult_87_CARRYB_40__7_), .S(u5_mult_87_SUMB_40__7_) );
  FA_X1 u5_mult_87_S2_40_6 ( .A(u5_mult_87_ab_40__6_), .B(
        u5_mult_87_CARRYB_39__6_), .CI(u5_mult_87_SUMB_39__7_), .CO(
        u5_mult_87_CARRYB_40__6_), .S(u5_mult_87_SUMB_40__6_) );
  FA_X1 u5_mult_87_S2_40_5 ( .A(u5_mult_87_ab_40__5_), .B(
        u5_mult_87_CARRYB_39__5_), .CI(u5_mult_87_SUMB_39__6_), .CO(
        u5_mult_87_CARRYB_40__5_), .S(u5_mult_87_SUMB_40__5_) );
  FA_X1 u5_mult_87_S2_40_4 ( .A(u5_mult_87_ab_40__4_), .B(
        u5_mult_87_CARRYB_39__4_), .CI(u5_mult_87_SUMB_39__5_), .CO(
        u5_mult_87_CARRYB_40__4_), .S(u5_mult_87_SUMB_40__4_) );
  FA_X1 u5_mult_87_S2_40_3 ( .A(u5_mult_87_ab_40__3_), .B(
        u5_mult_87_CARRYB_39__3_), .CI(u5_mult_87_SUMB_39__4_), .CO(
        u5_mult_87_CARRYB_40__3_), .S(u5_mult_87_SUMB_40__3_) );
  FA_X1 u5_mult_87_S2_40_2 ( .A(u5_mult_87_ab_40__2_), .B(
        u5_mult_87_CARRYB_39__2_), .CI(u5_mult_87_SUMB_39__3_), .CO(
        u5_mult_87_CARRYB_40__2_), .S(u5_mult_87_SUMB_40__2_) );
  FA_X1 u5_mult_87_S2_40_1 ( .A(u5_mult_87_ab_40__1_), .B(
        u5_mult_87_CARRYB_39__1_), .CI(u5_mult_87_SUMB_39__2_), .CO(
        u5_mult_87_CARRYB_40__1_), .S(u5_mult_87_SUMB_40__1_) );
  FA_X1 u5_mult_87_S1_40_0 ( .A(u5_mult_87_ab_40__0_), .B(
        u5_mult_87_CARRYB_39__0_), .CI(u5_mult_87_SUMB_39__1_), .CO(
        u5_mult_87_CARRYB_40__0_), .S(u5_N40) );
  FA_X1 u5_mult_87_S3_41_51 ( .A(u5_mult_87_ab_41__51_), .B(
        u5_mult_87_CARRYB_40__51_), .CI(u5_mult_87_ab_40__52_), .CO(
        u5_mult_87_CARRYB_41__51_), .S(u5_mult_87_SUMB_41__51_) );
  FA_X1 u5_mult_87_S2_41_50 ( .A(u5_mult_87_ab_41__50_), .B(
        u5_mult_87_CARRYB_40__50_), .CI(u5_mult_87_SUMB_40__51_), .CO(
        u5_mult_87_CARRYB_41__50_), .S(u5_mult_87_SUMB_41__50_) );
  FA_X1 u5_mult_87_S2_41_49 ( .A(u5_mult_87_ab_41__49_), .B(
        u5_mult_87_CARRYB_40__49_), .CI(u5_mult_87_SUMB_40__50_), .CO(
        u5_mult_87_CARRYB_41__49_), .S(u5_mult_87_SUMB_41__49_) );
  FA_X1 u5_mult_87_S2_41_48 ( .A(u5_mult_87_ab_41__48_), .B(
        u5_mult_87_CARRYB_40__48_), .CI(u5_mult_87_SUMB_40__49_), .CO(
        u5_mult_87_CARRYB_41__48_), .S(u5_mult_87_SUMB_41__48_) );
  FA_X1 u5_mult_87_S2_41_47 ( .A(u5_mult_87_ab_41__47_), .B(
        u5_mult_87_CARRYB_40__47_), .CI(u5_mult_87_SUMB_40__48_), .CO(
        u5_mult_87_CARRYB_41__47_), .S(u5_mult_87_SUMB_41__47_) );
  FA_X1 u5_mult_87_S2_41_46 ( .A(u5_mult_87_ab_41__46_), .B(
        u5_mult_87_CARRYB_40__46_), .CI(u5_mult_87_SUMB_40__47_), .CO(
        u5_mult_87_CARRYB_41__46_), .S(u5_mult_87_SUMB_41__46_) );
  FA_X1 u5_mult_87_S2_41_45 ( .A(u5_mult_87_ab_41__45_), .B(
        u5_mult_87_CARRYB_40__45_), .CI(u5_mult_87_SUMB_40__46_), .CO(
        u5_mult_87_CARRYB_41__45_), .S(u5_mult_87_SUMB_41__45_) );
  FA_X1 u5_mult_87_S2_41_44 ( .A(u5_mult_87_ab_41__44_), .B(
        u5_mult_87_CARRYB_40__44_), .CI(u5_mult_87_SUMB_40__45_), .CO(
        u5_mult_87_CARRYB_41__44_), .S(u5_mult_87_SUMB_41__44_) );
  FA_X1 u5_mult_87_S2_41_43 ( .A(u5_mult_87_ab_41__43_), .B(
        u5_mult_87_CARRYB_40__43_), .CI(u5_mult_87_SUMB_40__44_), .CO(
        u5_mult_87_CARRYB_41__43_), .S(u5_mult_87_SUMB_41__43_) );
  FA_X1 u5_mult_87_S2_41_42 ( .A(u5_mult_87_ab_41__42_), .B(
        u5_mult_87_CARRYB_40__42_), .CI(u5_mult_87_SUMB_40__43_), .CO(
        u5_mult_87_CARRYB_41__42_), .S(u5_mult_87_SUMB_41__42_) );
  FA_X1 u5_mult_87_S2_41_41 ( .A(u5_mult_87_ab_41__41_), .B(
        u5_mult_87_CARRYB_40__41_), .CI(u5_mult_87_SUMB_40__42_), .CO(
        u5_mult_87_CARRYB_41__41_), .S(u5_mult_87_SUMB_41__41_) );
  FA_X1 u5_mult_87_S2_41_40 ( .A(u5_mult_87_ab_41__40_), .B(
        u5_mult_87_CARRYB_40__40_), .CI(u5_mult_87_SUMB_40__41_), .CO(
        u5_mult_87_CARRYB_41__40_), .S(u5_mult_87_SUMB_41__40_) );
  FA_X1 u5_mult_87_S2_41_39 ( .A(u5_mult_87_ab_41__39_), .B(
        u5_mult_87_CARRYB_40__39_), .CI(u5_mult_87_SUMB_40__40_), .CO(
        u5_mult_87_CARRYB_41__39_), .S(u5_mult_87_SUMB_41__39_) );
  FA_X1 u5_mult_87_S2_41_38 ( .A(u5_mult_87_ab_41__38_), .B(
        u5_mult_87_CARRYB_40__38_), .CI(u5_mult_87_SUMB_40__39_), .CO(
        u5_mult_87_CARRYB_41__38_), .S(u5_mult_87_SUMB_41__38_) );
  FA_X1 u5_mult_87_S2_41_37 ( .A(u5_mult_87_ab_41__37_), .B(
        u5_mult_87_CARRYB_40__37_), .CI(u5_mult_87_SUMB_40__38_), .CO(
        u5_mult_87_CARRYB_41__37_), .S(u5_mult_87_SUMB_41__37_) );
  FA_X1 u5_mult_87_S2_41_36 ( .A(u5_mult_87_ab_41__36_), .B(
        u5_mult_87_CARRYB_40__36_), .CI(u5_mult_87_SUMB_40__37_), .CO(
        u5_mult_87_CARRYB_41__36_), .S(u5_mult_87_SUMB_41__36_) );
  FA_X1 u5_mult_87_S2_41_35 ( .A(u5_mult_87_ab_41__35_), .B(
        u5_mult_87_CARRYB_40__35_), .CI(u5_mult_87_SUMB_40__36_), .CO(
        u5_mult_87_CARRYB_41__35_), .S(u5_mult_87_SUMB_41__35_) );
  FA_X1 u5_mult_87_S2_41_34 ( .A(u5_mult_87_ab_41__34_), .B(
        u5_mult_87_CARRYB_40__34_), .CI(u5_mult_87_SUMB_40__35_), .CO(
        u5_mult_87_CARRYB_41__34_), .S(u5_mult_87_SUMB_41__34_) );
  FA_X1 u5_mult_87_S2_41_33 ( .A(u5_mult_87_ab_41__33_), .B(
        u5_mult_87_CARRYB_40__33_), .CI(u5_mult_87_SUMB_40__34_), .CO(
        u5_mult_87_CARRYB_41__33_), .S(u5_mult_87_SUMB_41__33_) );
  FA_X1 u5_mult_87_S2_41_32 ( .A(u5_mult_87_ab_41__32_), .B(
        u5_mult_87_CARRYB_40__32_), .CI(u5_mult_87_SUMB_40__33_), .CO(
        u5_mult_87_CARRYB_41__32_), .S(u5_mult_87_SUMB_41__32_) );
  FA_X1 u5_mult_87_S2_41_31 ( .A(u5_mult_87_ab_41__31_), .B(
        u5_mult_87_CARRYB_40__31_), .CI(u5_mult_87_SUMB_40__32_), .CO(
        u5_mult_87_CARRYB_41__31_), .S(u5_mult_87_SUMB_41__31_) );
  FA_X1 u5_mult_87_S2_41_30 ( .A(u5_mult_87_ab_41__30_), .B(
        u5_mult_87_CARRYB_40__30_), .CI(u5_mult_87_SUMB_40__31_), .CO(
        u5_mult_87_CARRYB_41__30_), .S(u5_mult_87_SUMB_41__30_) );
  FA_X1 u5_mult_87_S2_41_29 ( .A(u5_mult_87_ab_41__29_), .B(
        u5_mult_87_CARRYB_40__29_), .CI(u5_mult_87_SUMB_40__30_), .CO(
        u5_mult_87_CARRYB_41__29_), .S(u5_mult_87_SUMB_41__29_) );
  FA_X1 u5_mult_87_S2_41_28 ( .A(u5_mult_87_ab_41__28_), .B(
        u5_mult_87_CARRYB_40__28_), .CI(u5_mult_87_SUMB_40__29_), .CO(
        u5_mult_87_CARRYB_41__28_), .S(u5_mult_87_SUMB_41__28_) );
  FA_X1 u5_mult_87_S2_41_27 ( .A(u5_mult_87_ab_41__27_), .B(
        u5_mult_87_CARRYB_40__27_), .CI(u5_mult_87_SUMB_40__28_), .CO(
        u5_mult_87_CARRYB_41__27_), .S(u5_mult_87_SUMB_41__27_) );
  FA_X1 u5_mult_87_S2_41_26 ( .A(u5_mult_87_ab_41__26_), .B(
        u5_mult_87_CARRYB_40__26_), .CI(u5_mult_87_SUMB_40__27_), .CO(
        u5_mult_87_CARRYB_41__26_), .S(u5_mult_87_SUMB_41__26_) );
  FA_X1 u5_mult_87_S2_41_25 ( .A(u5_mult_87_ab_41__25_), .B(
        u5_mult_87_CARRYB_40__25_), .CI(u5_mult_87_SUMB_40__26_), .CO(
        u5_mult_87_CARRYB_41__25_), .S(u5_mult_87_SUMB_41__25_) );
  FA_X1 u5_mult_87_S2_41_24 ( .A(u5_mult_87_ab_41__24_), .B(
        u5_mult_87_CARRYB_40__24_), .CI(u5_mult_87_SUMB_40__25_), .CO(
        u5_mult_87_CARRYB_41__24_), .S(u5_mult_87_SUMB_41__24_) );
  FA_X1 u5_mult_87_S2_41_23 ( .A(u5_mult_87_ab_41__23_), .B(
        u5_mult_87_CARRYB_40__23_), .CI(u5_mult_87_SUMB_40__24_), .CO(
        u5_mult_87_CARRYB_41__23_), .S(u5_mult_87_SUMB_41__23_) );
  FA_X1 u5_mult_87_S2_41_22 ( .A(u5_mult_87_ab_41__22_), .B(
        u5_mult_87_CARRYB_40__22_), .CI(u5_mult_87_SUMB_40__23_), .CO(
        u5_mult_87_CARRYB_41__22_), .S(u5_mult_87_SUMB_41__22_) );
  FA_X1 u5_mult_87_S2_41_21 ( .A(u5_mult_87_ab_41__21_), .B(
        u5_mult_87_CARRYB_40__21_), .CI(u5_mult_87_SUMB_40__22_), .CO(
        u5_mult_87_CARRYB_41__21_), .S(u5_mult_87_SUMB_41__21_) );
  FA_X1 u5_mult_87_S2_41_20 ( .A(u5_mult_87_ab_41__20_), .B(
        u5_mult_87_CARRYB_40__20_), .CI(u5_mult_87_SUMB_40__21_), .CO(
        u5_mult_87_CARRYB_41__20_), .S(u5_mult_87_SUMB_41__20_) );
  FA_X1 u5_mult_87_S2_41_19 ( .A(u5_mult_87_ab_41__19_), .B(
        u5_mult_87_CARRYB_40__19_), .CI(u5_mult_87_SUMB_40__20_), .CO(
        u5_mult_87_CARRYB_41__19_), .S(u5_mult_87_SUMB_41__19_) );
  FA_X1 u5_mult_87_S2_41_18 ( .A(u5_mult_87_ab_41__18_), .B(
        u5_mult_87_CARRYB_40__18_), .CI(u5_mult_87_SUMB_40__19_), .CO(
        u5_mult_87_CARRYB_41__18_), .S(u5_mult_87_SUMB_41__18_) );
  FA_X1 u5_mult_87_S2_41_17 ( .A(u5_mult_87_ab_41__17_), .B(
        u5_mult_87_CARRYB_40__17_), .CI(u5_mult_87_SUMB_40__18_), .CO(
        u5_mult_87_CARRYB_41__17_), .S(u5_mult_87_SUMB_41__17_) );
  FA_X1 u5_mult_87_S2_41_16 ( .A(u5_mult_87_ab_41__16_), .B(
        u5_mult_87_CARRYB_40__16_), .CI(u5_mult_87_SUMB_40__17_), .CO(
        u5_mult_87_CARRYB_41__16_), .S(u5_mult_87_SUMB_41__16_) );
  FA_X1 u5_mult_87_S2_41_15 ( .A(u5_mult_87_ab_41__15_), .B(
        u5_mult_87_CARRYB_40__15_), .CI(u5_mult_87_SUMB_40__16_), .CO(
        u5_mult_87_CARRYB_41__15_), .S(u5_mult_87_SUMB_41__15_) );
  FA_X1 u5_mult_87_S2_41_14 ( .A(u5_mult_87_ab_41__14_), .B(
        u5_mult_87_CARRYB_40__14_), .CI(u5_mult_87_SUMB_40__15_), .CO(
        u5_mult_87_CARRYB_41__14_), .S(u5_mult_87_SUMB_41__14_) );
  FA_X1 u5_mult_87_S2_41_13 ( .A(u5_mult_87_ab_41__13_), .B(
        u5_mult_87_CARRYB_40__13_), .CI(u5_mult_87_SUMB_40__14_), .CO(
        u5_mult_87_CARRYB_41__13_), .S(u5_mult_87_SUMB_41__13_) );
  FA_X1 u5_mult_87_S2_41_12 ( .A(u5_mult_87_ab_41__12_), .B(
        u5_mult_87_CARRYB_40__12_), .CI(u5_mult_87_SUMB_40__13_), .CO(
        u5_mult_87_CARRYB_41__12_), .S(u5_mult_87_SUMB_41__12_) );
  FA_X1 u5_mult_87_S2_41_11 ( .A(u5_mult_87_ab_41__11_), .B(
        u5_mult_87_CARRYB_40__11_), .CI(u5_mult_87_SUMB_40__12_), .CO(
        u5_mult_87_CARRYB_41__11_), .S(u5_mult_87_SUMB_41__11_) );
  FA_X1 u5_mult_87_S2_41_10 ( .A(u5_mult_87_ab_41__10_), .B(
        u5_mult_87_CARRYB_40__10_), .CI(u5_mult_87_SUMB_40__11_), .CO(
        u5_mult_87_CARRYB_41__10_), .S(u5_mult_87_SUMB_41__10_) );
  FA_X1 u5_mult_87_S2_41_9 ( .A(u5_mult_87_ab_41__9_), .B(
        u5_mult_87_CARRYB_40__9_), .CI(u5_mult_87_SUMB_40__10_), .CO(
        u5_mult_87_CARRYB_41__9_), .S(u5_mult_87_SUMB_41__9_) );
  FA_X1 u5_mult_87_S2_41_8 ( .A(u5_mult_87_ab_41__8_), .B(
        u5_mult_87_CARRYB_40__8_), .CI(u5_mult_87_SUMB_40__9_), .CO(
        u5_mult_87_CARRYB_41__8_), .S(u5_mult_87_SUMB_41__8_) );
  FA_X1 u5_mult_87_S2_41_7 ( .A(u5_mult_87_ab_41__7_), .B(
        u5_mult_87_CARRYB_40__7_), .CI(u5_mult_87_SUMB_40__8_), .CO(
        u5_mult_87_CARRYB_41__7_), .S(u5_mult_87_SUMB_41__7_) );
  FA_X1 u5_mult_87_S2_41_6 ( .A(u5_mult_87_ab_41__6_), .B(
        u5_mult_87_CARRYB_40__6_), .CI(u5_mult_87_SUMB_40__7_), .CO(
        u5_mult_87_CARRYB_41__6_), .S(u5_mult_87_SUMB_41__6_) );
  FA_X1 u5_mult_87_S2_41_5 ( .A(u5_mult_87_ab_41__5_), .B(
        u5_mult_87_CARRYB_40__5_), .CI(u5_mult_87_SUMB_40__6_), .CO(
        u5_mult_87_CARRYB_41__5_), .S(u5_mult_87_SUMB_41__5_) );
  FA_X1 u5_mult_87_S2_41_4 ( .A(u5_mult_87_ab_41__4_), .B(
        u5_mult_87_CARRYB_40__4_), .CI(u5_mult_87_SUMB_40__5_), .CO(
        u5_mult_87_CARRYB_41__4_), .S(u5_mult_87_SUMB_41__4_) );
  FA_X1 u5_mult_87_S2_41_3 ( .A(u5_mult_87_ab_41__3_), .B(
        u5_mult_87_CARRYB_40__3_), .CI(u5_mult_87_SUMB_40__4_), .CO(
        u5_mult_87_CARRYB_41__3_), .S(u5_mult_87_SUMB_41__3_) );
  FA_X1 u5_mult_87_S2_41_2 ( .A(u5_mult_87_ab_41__2_), .B(
        u5_mult_87_CARRYB_40__2_), .CI(u5_mult_87_SUMB_40__3_), .CO(
        u5_mult_87_CARRYB_41__2_), .S(u5_mult_87_SUMB_41__2_) );
  FA_X1 u5_mult_87_S2_41_1 ( .A(u5_mult_87_ab_41__1_), .B(
        u5_mult_87_CARRYB_40__1_), .CI(u5_mult_87_SUMB_40__2_), .CO(
        u5_mult_87_CARRYB_41__1_), .S(u5_mult_87_SUMB_41__1_) );
  FA_X1 u5_mult_87_S1_41_0 ( .A(u5_mult_87_ab_41__0_), .B(
        u5_mult_87_CARRYB_40__0_), .CI(u5_mult_87_SUMB_40__1_), .CO(
        u5_mult_87_CARRYB_41__0_), .S(u5_N41) );
  FA_X1 u5_mult_87_S3_42_51 ( .A(u5_mult_87_ab_42__51_), .B(
        u5_mult_87_CARRYB_41__51_), .CI(u5_mult_87_ab_41__52_), .CO(
        u5_mult_87_CARRYB_42__51_), .S(u5_mult_87_SUMB_42__51_) );
  FA_X1 u5_mult_87_S2_42_50 ( .A(u5_mult_87_ab_42__50_), .B(
        u5_mult_87_CARRYB_41__50_), .CI(u5_mult_87_SUMB_41__51_), .CO(
        u5_mult_87_CARRYB_42__50_), .S(u5_mult_87_SUMB_42__50_) );
  FA_X1 u5_mult_87_S2_42_49 ( .A(u5_mult_87_ab_42__49_), .B(
        u5_mult_87_CARRYB_41__49_), .CI(u5_mult_87_SUMB_41__50_), .CO(
        u5_mult_87_CARRYB_42__49_), .S(u5_mult_87_SUMB_42__49_) );
  FA_X1 u5_mult_87_S2_42_48 ( .A(u5_mult_87_ab_42__48_), .B(
        u5_mult_87_CARRYB_41__48_), .CI(u5_mult_87_SUMB_41__49_), .CO(
        u5_mult_87_CARRYB_42__48_), .S(u5_mult_87_SUMB_42__48_) );
  FA_X1 u5_mult_87_S2_42_47 ( .A(u5_mult_87_ab_42__47_), .B(
        u5_mult_87_CARRYB_41__47_), .CI(u5_mult_87_SUMB_41__48_), .CO(
        u5_mult_87_CARRYB_42__47_), .S(u5_mult_87_SUMB_42__47_) );
  FA_X1 u5_mult_87_S2_42_46 ( .A(u5_mult_87_ab_42__46_), .B(
        u5_mult_87_CARRYB_41__46_), .CI(u5_mult_87_SUMB_41__47_), .CO(
        u5_mult_87_CARRYB_42__46_), .S(u5_mult_87_SUMB_42__46_) );
  FA_X1 u5_mult_87_S2_42_45 ( .A(u5_mult_87_ab_42__45_), .B(
        u5_mult_87_CARRYB_41__45_), .CI(u5_mult_87_SUMB_41__46_), .CO(
        u5_mult_87_CARRYB_42__45_), .S(u5_mult_87_SUMB_42__45_) );
  FA_X1 u5_mult_87_S2_42_44 ( .A(u5_mult_87_ab_42__44_), .B(
        u5_mult_87_CARRYB_41__44_), .CI(u5_mult_87_SUMB_41__45_), .CO(
        u5_mult_87_CARRYB_42__44_), .S(u5_mult_87_SUMB_42__44_) );
  FA_X1 u5_mult_87_S2_42_43 ( .A(u5_mult_87_ab_42__43_), .B(
        u5_mult_87_CARRYB_41__43_), .CI(u5_mult_87_SUMB_41__44_), .CO(
        u5_mult_87_CARRYB_42__43_), .S(u5_mult_87_SUMB_42__43_) );
  FA_X1 u5_mult_87_S2_42_42 ( .A(u5_mult_87_ab_42__42_), .B(
        u5_mult_87_CARRYB_41__42_), .CI(u5_mult_87_SUMB_41__43_), .CO(
        u5_mult_87_CARRYB_42__42_), .S(u5_mult_87_SUMB_42__42_) );
  FA_X1 u5_mult_87_S2_42_41 ( .A(u5_mult_87_ab_42__41_), .B(
        u5_mult_87_CARRYB_41__41_), .CI(u5_mult_87_SUMB_41__42_), .CO(
        u5_mult_87_CARRYB_42__41_), .S(u5_mult_87_SUMB_42__41_) );
  FA_X1 u5_mult_87_S2_42_40 ( .A(u5_mult_87_ab_42__40_), .B(
        u5_mult_87_CARRYB_41__40_), .CI(u5_mult_87_SUMB_41__41_), .CO(
        u5_mult_87_CARRYB_42__40_), .S(u5_mult_87_SUMB_42__40_) );
  FA_X1 u5_mult_87_S2_42_39 ( .A(u5_mult_87_ab_42__39_), .B(
        u5_mult_87_CARRYB_41__39_), .CI(u5_mult_87_SUMB_41__40_), .CO(
        u5_mult_87_CARRYB_42__39_), .S(u5_mult_87_SUMB_42__39_) );
  FA_X1 u5_mult_87_S2_42_38 ( .A(u5_mult_87_ab_42__38_), .B(
        u5_mult_87_CARRYB_41__38_), .CI(u5_mult_87_SUMB_41__39_), .CO(
        u5_mult_87_CARRYB_42__38_), .S(u5_mult_87_SUMB_42__38_) );
  FA_X1 u5_mult_87_S2_42_37 ( .A(u5_mult_87_ab_42__37_), .B(
        u5_mult_87_CARRYB_41__37_), .CI(u5_mult_87_SUMB_41__38_), .CO(
        u5_mult_87_CARRYB_42__37_), .S(u5_mult_87_SUMB_42__37_) );
  FA_X1 u5_mult_87_S2_42_36 ( .A(u5_mult_87_ab_42__36_), .B(
        u5_mult_87_CARRYB_41__36_), .CI(u5_mult_87_SUMB_41__37_), .CO(
        u5_mult_87_CARRYB_42__36_), .S(u5_mult_87_SUMB_42__36_) );
  FA_X1 u5_mult_87_S2_42_35 ( .A(u5_mult_87_ab_42__35_), .B(
        u5_mult_87_CARRYB_41__35_), .CI(u5_mult_87_SUMB_41__36_), .CO(
        u5_mult_87_CARRYB_42__35_), .S(u5_mult_87_SUMB_42__35_) );
  FA_X1 u5_mult_87_S2_42_34 ( .A(u5_mult_87_ab_42__34_), .B(
        u5_mult_87_CARRYB_41__34_), .CI(u5_mult_87_SUMB_41__35_), .CO(
        u5_mult_87_CARRYB_42__34_), .S(u5_mult_87_SUMB_42__34_) );
  FA_X1 u5_mult_87_S2_42_33 ( .A(u5_mult_87_ab_42__33_), .B(
        u5_mult_87_CARRYB_41__33_), .CI(u5_mult_87_SUMB_41__34_), .CO(
        u5_mult_87_CARRYB_42__33_), .S(u5_mult_87_SUMB_42__33_) );
  FA_X1 u5_mult_87_S2_42_32 ( .A(u5_mult_87_ab_42__32_), .B(
        u5_mult_87_CARRYB_41__32_), .CI(u5_mult_87_SUMB_41__33_), .CO(
        u5_mult_87_CARRYB_42__32_), .S(u5_mult_87_SUMB_42__32_) );
  FA_X1 u5_mult_87_S2_42_31 ( .A(u5_mult_87_ab_42__31_), .B(
        u5_mult_87_CARRYB_41__31_), .CI(u5_mult_87_SUMB_41__32_), .CO(
        u5_mult_87_CARRYB_42__31_), .S(u5_mult_87_SUMB_42__31_) );
  FA_X1 u5_mult_87_S2_42_30 ( .A(u5_mult_87_ab_42__30_), .B(
        u5_mult_87_CARRYB_41__30_), .CI(u5_mult_87_SUMB_41__31_), .CO(
        u5_mult_87_CARRYB_42__30_), .S(u5_mult_87_SUMB_42__30_) );
  FA_X1 u5_mult_87_S2_42_29 ( .A(u5_mult_87_ab_42__29_), .B(
        u5_mult_87_CARRYB_41__29_), .CI(u5_mult_87_SUMB_41__30_), .CO(
        u5_mult_87_CARRYB_42__29_), .S(u5_mult_87_SUMB_42__29_) );
  FA_X1 u5_mult_87_S2_42_28 ( .A(u5_mult_87_ab_42__28_), .B(
        u5_mult_87_CARRYB_41__28_), .CI(u5_mult_87_SUMB_41__29_), .CO(
        u5_mult_87_CARRYB_42__28_), .S(u5_mult_87_SUMB_42__28_) );
  FA_X1 u5_mult_87_S2_42_27 ( .A(u5_mult_87_ab_42__27_), .B(
        u5_mult_87_CARRYB_41__27_), .CI(u5_mult_87_SUMB_41__28_), .CO(
        u5_mult_87_CARRYB_42__27_), .S(u5_mult_87_SUMB_42__27_) );
  FA_X1 u5_mult_87_S2_42_26 ( .A(u5_mult_87_ab_42__26_), .B(
        u5_mult_87_CARRYB_41__26_), .CI(u5_mult_87_SUMB_41__27_), .CO(
        u5_mult_87_CARRYB_42__26_), .S(u5_mult_87_SUMB_42__26_) );
  FA_X1 u5_mult_87_S2_42_25 ( .A(u5_mult_87_ab_42__25_), .B(
        u5_mult_87_CARRYB_41__25_), .CI(u5_mult_87_SUMB_41__26_), .CO(
        u5_mult_87_CARRYB_42__25_), .S(u5_mult_87_SUMB_42__25_) );
  FA_X1 u5_mult_87_S2_42_24 ( .A(u5_mult_87_ab_42__24_), .B(
        u5_mult_87_CARRYB_41__24_), .CI(u5_mult_87_SUMB_41__25_), .CO(
        u5_mult_87_CARRYB_42__24_), .S(u5_mult_87_SUMB_42__24_) );
  FA_X1 u5_mult_87_S2_42_23 ( .A(u5_mult_87_ab_42__23_), .B(
        u5_mult_87_CARRYB_41__23_), .CI(u5_mult_87_SUMB_41__24_), .CO(
        u5_mult_87_CARRYB_42__23_), .S(u5_mult_87_SUMB_42__23_) );
  FA_X1 u5_mult_87_S2_42_22 ( .A(u5_mult_87_ab_42__22_), .B(
        u5_mult_87_CARRYB_41__22_), .CI(u5_mult_87_SUMB_41__23_), .CO(
        u5_mult_87_CARRYB_42__22_), .S(u5_mult_87_SUMB_42__22_) );
  FA_X1 u5_mult_87_S2_42_21 ( .A(u5_mult_87_ab_42__21_), .B(
        u5_mult_87_CARRYB_41__21_), .CI(u5_mult_87_SUMB_41__22_), .CO(
        u5_mult_87_CARRYB_42__21_), .S(u5_mult_87_SUMB_42__21_) );
  FA_X1 u5_mult_87_S2_42_20 ( .A(u5_mult_87_ab_42__20_), .B(
        u5_mult_87_CARRYB_41__20_), .CI(u5_mult_87_SUMB_41__21_), .CO(
        u5_mult_87_CARRYB_42__20_), .S(u5_mult_87_SUMB_42__20_) );
  FA_X1 u5_mult_87_S2_42_19 ( .A(u5_mult_87_ab_42__19_), .B(
        u5_mult_87_CARRYB_41__19_), .CI(u5_mult_87_SUMB_41__20_), .CO(
        u5_mult_87_CARRYB_42__19_), .S(u5_mult_87_SUMB_42__19_) );
  FA_X1 u5_mult_87_S2_42_18 ( .A(u5_mult_87_ab_42__18_), .B(
        u5_mult_87_CARRYB_41__18_), .CI(u5_mult_87_SUMB_41__19_), .CO(
        u5_mult_87_CARRYB_42__18_), .S(u5_mult_87_SUMB_42__18_) );
  FA_X1 u5_mult_87_S2_42_17 ( .A(u5_mult_87_ab_42__17_), .B(
        u5_mult_87_CARRYB_41__17_), .CI(u5_mult_87_SUMB_41__18_), .CO(
        u5_mult_87_CARRYB_42__17_), .S(u5_mult_87_SUMB_42__17_) );
  FA_X1 u5_mult_87_S2_42_16 ( .A(u5_mult_87_ab_42__16_), .B(
        u5_mult_87_CARRYB_41__16_), .CI(u5_mult_87_SUMB_41__17_), .CO(
        u5_mult_87_CARRYB_42__16_), .S(u5_mult_87_SUMB_42__16_) );
  FA_X1 u5_mult_87_S2_42_15 ( .A(u5_mult_87_ab_42__15_), .B(
        u5_mult_87_CARRYB_41__15_), .CI(u5_mult_87_SUMB_41__16_), .CO(
        u5_mult_87_CARRYB_42__15_), .S(u5_mult_87_SUMB_42__15_) );
  FA_X1 u5_mult_87_S2_42_14 ( .A(u5_mult_87_ab_42__14_), .B(
        u5_mult_87_CARRYB_41__14_), .CI(u5_mult_87_SUMB_41__15_), .CO(
        u5_mult_87_CARRYB_42__14_), .S(u5_mult_87_SUMB_42__14_) );
  FA_X1 u5_mult_87_S2_42_13 ( .A(u5_mult_87_ab_42__13_), .B(
        u5_mult_87_CARRYB_41__13_), .CI(u5_mult_87_SUMB_41__14_), .CO(
        u5_mult_87_CARRYB_42__13_), .S(u5_mult_87_SUMB_42__13_) );
  FA_X1 u5_mult_87_S2_42_12 ( .A(u5_mult_87_ab_42__12_), .B(
        u5_mult_87_CARRYB_41__12_), .CI(u5_mult_87_SUMB_41__13_), .CO(
        u5_mult_87_CARRYB_42__12_), .S(u5_mult_87_SUMB_42__12_) );
  FA_X1 u5_mult_87_S2_42_11 ( .A(u5_mult_87_ab_42__11_), .B(
        u5_mult_87_CARRYB_41__11_), .CI(u5_mult_87_SUMB_41__12_), .CO(
        u5_mult_87_CARRYB_42__11_), .S(u5_mult_87_SUMB_42__11_) );
  FA_X1 u5_mult_87_S2_42_10 ( .A(u5_mult_87_ab_42__10_), .B(
        u5_mult_87_CARRYB_41__10_), .CI(u5_mult_87_SUMB_41__11_), .CO(
        u5_mult_87_CARRYB_42__10_), .S(u5_mult_87_SUMB_42__10_) );
  FA_X1 u5_mult_87_S2_42_9 ( .A(u5_mult_87_ab_42__9_), .B(
        u5_mult_87_CARRYB_41__9_), .CI(u5_mult_87_SUMB_41__10_), .CO(
        u5_mult_87_CARRYB_42__9_), .S(u5_mult_87_SUMB_42__9_) );
  FA_X1 u5_mult_87_S2_42_8 ( .A(u5_mult_87_ab_42__8_), .B(
        u5_mult_87_CARRYB_41__8_), .CI(u5_mult_87_SUMB_41__9_), .CO(
        u5_mult_87_CARRYB_42__8_), .S(u5_mult_87_SUMB_42__8_) );
  FA_X1 u5_mult_87_S2_42_7 ( .A(u5_mult_87_ab_42__7_), .B(
        u5_mult_87_CARRYB_41__7_), .CI(u5_mult_87_SUMB_41__8_), .CO(
        u5_mult_87_CARRYB_42__7_), .S(u5_mult_87_SUMB_42__7_) );
  FA_X1 u5_mult_87_S2_42_6 ( .A(u5_mult_87_ab_42__6_), .B(
        u5_mult_87_CARRYB_41__6_), .CI(u5_mult_87_SUMB_41__7_), .CO(
        u5_mult_87_CARRYB_42__6_), .S(u5_mult_87_SUMB_42__6_) );
  FA_X1 u5_mult_87_S2_42_5 ( .A(u5_mult_87_ab_42__5_), .B(
        u5_mult_87_CARRYB_41__5_), .CI(u5_mult_87_SUMB_41__6_), .CO(
        u5_mult_87_CARRYB_42__5_), .S(u5_mult_87_SUMB_42__5_) );
  FA_X1 u5_mult_87_S2_42_4 ( .A(u5_mult_87_ab_42__4_), .B(
        u5_mult_87_CARRYB_41__4_), .CI(u5_mult_87_SUMB_41__5_), .CO(
        u5_mult_87_CARRYB_42__4_), .S(u5_mult_87_SUMB_42__4_) );
  FA_X1 u5_mult_87_S2_42_3 ( .A(u5_mult_87_ab_42__3_), .B(
        u5_mult_87_CARRYB_41__3_), .CI(u5_mult_87_SUMB_41__4_), .CO(
        u5_mult_87_CARRYB_42__3_), .S(u5_mult_87_SUMB_42__3_) );
  FA_X1 u5_mult_87_S2_42_2 ( .A(u5_mult_87_ab_42__2_), .B(
        u5_mult_87_CARRYB_41__2_), .CI(u5_mult_87_SUMB_41__3_), .CO(
        u5_mult_87_CARRYB_42__2_), .S(u5_mult_87_SUMB_42__2_) );
  FA_X1 u5_mult_87_S2_42_1 ( .A(u5_mult_87_ab_42__1_), .B(
        u5_mult_87_CARRYB_41__1_), .CI(u5_mult_87_SUMB_41__2_), .CO(
        u5_mult_87_CARRYB_42__1_), .S(u5_mult_87_SUMB_42__1_) );
  FA_X1 u5_mult_87_S1_42_0 ( .A(u5_mult_87_ab_42__0_), .B(
        u5_mult_87_CARRYB_41__0_), .CI(u5_mult_87_SUMB_41__1_), .CO(
        u5_mult_87_CARRYB_42__0_), .S(u5_N42) );
  FA_X1 u5_mult_87_S3_43_51 ( .A(u5_mult_87_ab_43__51_), .B(
        u5_mult_87_CARRYB_42__51_), .CI(u5_mult_87_ab_42__52_), .CO(
        u5_mult_87_CARRYB_43__51_), .S(u5_mult_87_SUMB_43__51_) );
  FA_X1 u5_mult_87_S2_43_50 ( .A(u5_mult_87_ab_43__50_), .B(
        u5_mult_87_CARRYB_42__50_), .CI(u5_mult_87_SUMB_42__51_), .CO(
        u5_mult_87_CARRYB_43__50_), .S(u5_mult_87_SUMB_43__50_) );
  FA_X1 u5_mult_87_S2_43_49 ( .A(u5_mult_87_ab_43__49_), .B(
        u5_mult_87_CARRYB_42__49_), .CI(u5_mult_87_SUMB_42__50_), .CO(
        u5_mult_87_CARRYB_43__49_), .S(u5_mult_87_SUMB_43__49_) );
  FA_X1 u5_mult_87_S2_43_48 ( .A(u5_mult_87_ab_43__48_), .B(
        u5_mult_87_CARRYB_42__48_), .CI(u5_mult_87_SUMB_42__49_), .CO(
        u5_mult_87_CARRYB_43__48_), .S(u5_mult_87_SUMB_43__48_) );
  FA_X1 u5_mult_87_S2_43_47 ( .A(u5_mult_87_ab_43__47_), .B(
        u5_mult_87_CARRYB_42__47_), .CI(u5_mult_87_SUMB_42__48_), .CO(
        u5_mult_87_CARRYB_43__47_), .S(u5_mult_87_SUMB_43__47_) );
  FA_X1 u5_mult_87_S2_43_46 ( .A(u5_mult_87_ab_43__46_), .B(
        u5_mult_87_CARRYB_42__46_), .CI(u5_mult_87_SUMB_42__47_), .CO(
        u5_mult_87_CARRYB_43__46_), .S(u5_mult_87_SUMB_43__46_) );
  FA_X1 u5_mult_87_S2_43_45 ( .A(u5_mult_87_ab_43__45_), .B(
        u5_mult_87_CARRYB_42__45_), .CI(u5_mult_87_SUMB_42__46_), .CO(
        u5_mult_87_CARRYB_43__45_), .S(u5_mult_87_SUMB_43__45_) );
  FA_X1 u5_mult_87_S2_43_44 ( .A(u5_mult_87_ab_43__44_), .B(
        u5_mult_87_CARRYB_42__44_), .CI(u5_mult_87_SUMB_42__45_), .CO(
        u5_mult_87_CARRYB_43__44_), .S(u5_mult_87_SUMB_43__44_) );
  FA_X1 u5_mult_87_S2_43_43 ( .A(u5_mult_87_ab_43__43_), .B(
        u5_mult_87_CARRYB_42__43_), .CI(u5_mult_87_SUMB_42__44_), .CO(
        u5_mult_87_CARRYB_43__43_), .S(u5_mult_87_SUMB_43__43_) );
  FA_X1 u5_mult_87_S2_43_42 ( .A(u5_mult_87_ab_43__42_), .B(
        u5_mult_87_CARRYB_42__42_), .CI(u5_mult_87_SUMB_42__43_), .CO(
        u5_mult_87_CARRYB_43__42_), .S(u5_mult_87_SUMB_43__42_) );
  FA_X1 u5_mult_87_S2_43_41 ( .A(u5_mult_87_ab_43__41_), .B(
        u5_mult_87_CARRYB_42__41_), .CI(u5_mult_87_SUMB_42__42_), .CO(
        u5_mult_87_CARRYB_43__41_), .S(u5_mult_87_SUMB_43__41_) );
  FA_X1 u5_mult_87_S2_43_40 ( .A(u5_mult_87_ab_43__40_), .B(
        u5_mult_87_CARRYB_42__40_), .CI(u5_mult_87_SUMB_42__41_), .CO(
        u5_mult_87_CARRYB_43__40_), .S(u5_mult_87_SUMB_43__40_) );
  FA_X1 u5_mult_87_S2_43_39 ( .A(u5_mult_87_ab_43__39_), .B(
        u5_mult_87_CARRYB_42__39_), .CI(u5_mult_87_SUMB_42__40_), .CO(
        u5_mult_87_CARRYB_43__39_), .S(u5_mult_87_SUMB_43__39_) );
  FA_X1 u5_mult_87_S2_43_38 ( .A(u5_mult_87_ab_43__38_), .B(
        u5_mult_87_CARRYB_42__38_), .CI(u5_mult_87_SUMB_42__39_), .CO(
        u5_mult_87_CARRYB_43__38_), .S(u5_mult_87_SUMB_43__38_) );
  FA_X1 u5_mult_87_S2_43_37 ( .A(u5_mult_87_ab_43__37_), .B(
        u5_mult_87_CARRYB_42__37_), .CI(u5_mult_87_SUMB_42__38_), .CO(
        u5_mult_87_CARRYB_43__37_), .S(u5_mult_87_SUMB_43__37_) );
  FA_X1 u5_mult_87_S2_43_36 ( .A(u5_mult_87_ab_43__36_), .B(
        u5_mult_87_CARRYB_42__36_), .CI(u5_mult_87_SUMB_42__37_), .CO(
        u5_mult_87_CARRYB_43__36_), .S(u5_mult_87_SUMB_43__36_) );
  FA_X1 u5_mult_87_S2_43_35 ( .A(u5_mult_87_ab_43__35_), .B(
        u5_mult_87_CARRYB_42__35_), .CI(u5_mult_87_SUMB_42__36_), .CO(
        u5_mult_87_CARRYB_43__35_), .S(u5_mult_87_SUMB_43__35_) );
  FA_X1 u5_mult_87_S2_43_34 ( .A(u5_mult_87_ab_43__34_), .B(
        u5_mult_87_CARRYB_42__34_), .CI(u5_mult_87_SUMB_42__35_), .CO(
        u5_mult_87_CARRYB_43__34_), .S(u5_mult_87_SUMB_43__34_) );
  FA_X1 u5_mult_87_S2_43_33 ( .A(u5_mult_87_ab_43__33_), .B(
        u5_mult_87_CARRYB_42__33_), .CI(u5_mult_87_SUMB_42__34_), .CO(
        u5_mult_87_CARRYB_43__33_), .S(u5_mult_87_SUMB_43__33_) );
  FA_X1 u5_mult_87_S2_43_32 ( .A(u5_mult_87_ab_43__32_), .B(
        u5_mult_87_CARRYB_42__32_), .CI(u5_mult_87_SUMB_42__33_), .CO(
        u5_mult_87_CARRYB_43__32_), .S(u5_mult_87_SUMB_43__32_) );
  FA_X1 u5_mult_87_S2_43_31 ( .A(u5_mult_87_ab_43__31_), .B(
        u5_mult_87_CARRYB_42__31_), .CI(u5_mult_87_SUMB_42__32_), .CO(
        u5_mult_87_CARRYB_43__31_), .S(u5_mult_87_SUMB_43__31_) );
  FA_X1 u5_mult_87_S2_43_30 ( .A(u5_mult_87_ab_43__30_), .B(
        u5_mult_87_CARRYB_42__30_), .CI(u5_mult_87_SUMB_42__31_), .CO(
        u5_mult_87_CARRYB_43__30_), .S(u5_mult_87_SUMB_43__30_) );
  FA_X1 u5_mult_87_S2_43_29 ( .A(u5_mult_87_ab_43__29_), .B(
        u5_mult_87_CARRYB_42__29_), .CI(u5_mult_87_SUMB_42__30_), .CO(
        u5_mult_87_CARRYB_43__29_), .S(u5_mult_87_SUMB_43__29_) );
  FA_X1 u5_mult_87_S2_43_28 ( .A(u5_mult_87_ab_43__28_), .B(
        u5_mult_87_CARRYB_42__28_), .CI(u5_mult_87_SUMB_42__29_), .CO(
        u5_mult_87_CARRYB_43__28_), .S(u5_mult_87_SUMB_43__28_) );
  FA_X1 u5_mult_87_S2_43_27 ( .A(u5_mult_87_ab_43__27_), .B(
        u5_mult_87_CARRYB_42__27_), .CI(u5_mult_87_SUMB_42__28_), .CO(
        u5_mult_87_CARRYB_43__27_), .S(u5_mult_87_SUMB_43__27_) );
  FA_X1 u5_mult_87_S2_43_26 ( .A(u5_mult_87_ab_43__26_), .B(
        u5_mult_87_CARRYB_42__26_), .CI(u5_mult_87_SUMB_42__27_), .CO(
        u5_mult_87_CARRYB_43__26_), .S(u5_mult_87_SUMB_43__26_) );
  FA_X1 u5_mult_87_S2_43_25 ( .A(u5_mult_87_ab_43__25_), .B(
        u5_mult_87_CARRYB_42__25_), .CI(u5_mult_87_SUMB_42__26_), .CO(
        u5_mult_87_CARRYB_43__25_), .S(u5_mult_87_SUMB_43__25_) );
  FA_X1 u5_mult_87_S2_43_24 ( .A(u5_mult_87_ab_43__24_), .B(
        u5_mult_87_CARRYB_42__24_), .CI(u5_mult_87_SUMB_42__25_), .CO(
        u5_mult_87_CARRYB_43__24_), .S(u5_mult_87_SUMB_43__24_) );
  FA_X1 u5_mult_87_S2_43_23 ( .A(u5_mult_87_ab_43__23_), .B(
        u5_mult_87_CARRYB_42__23_), .CI(u5_mult_87_SUMB_42__24_), .CO(
        u5_mult_87_CARRYB_43__23_), .S(u5_mult_87_SUMB_43__23_) );
  FA_X1 u5_mult_87_S2_43_22 ( .A(u5_mult_87_ab_43__22_), .B(
        u5_mult_87_CARRYB_42__22_), .CI(u5_mult_87_SUMB_42__23_), .CO(
        u5_mult_87_CARRYB_43__22_), .S(u5_mult_87_SUMB_43__22_) );
  FA_X1 u5_mult_87_S2_43_21 ( .A(u5_mult_87_ab_43__21_), .B(
        u5_mult_87_CARRYB_42__21_), .CI(u5_mult_87_SUMB_42__22_), .CO(
        u5_mult_87_CARRYB_43__21_), .S(u5_mult_87_SUMB_43__21_) );
  FA_X1 u5_mult_87_S2_43_20 ( .A(u5_mult_87_ab_43__20_), .B(
        u5_mult_87_CARRYB_42__20_), .CI(u5_mult_87_SUMB_42__21_), .CO(
        u5_mult_87_CARRYB_43__20_), .S(u5_mult_87_SUMB_43__20_) );
  FA_X1 u5_mult_87_S2_43_19 ( .A(u5_mult_87_ab_43__19_), .B(
        u5_mult_87_CARRYB_42__19_), .CI(u5_mult_87_SUMB_42__20_), .CO(
        u5_mult_87_CARRYB_43__19_), .S(u5_mult_87_SUMB_43__19_) );
  FA_X1 u5_mult_87_S2_43_18 ( .A(u5_mult_87_ab_43__18_), .B(
        u5_mult_87_CARRYB_42__18_), .CI(u5_mult_87_SUMB_42__19_), .CO(
        u5_mult_87_CARRYB_43__18_), .S(u5_mult_87_SUMB_43__18_) );
  FA_X1 u5_mult_87_S2_43_17 ( .A(u5_mult_87_ab_43__17_), .B(
        u5_mult_87_CARRYB_42__17_), .CI(u5_mult_87_SUMB_42__18_), .CO(
        u5_mult_87_CARRYB_43__17_), .S(u5_mult_87_SUMB_43__17_) );
  FA_X1 u5_mult_87_S2_43_16 ( .A(u5_mult_87_ab_43__16_), .B(
        u5_mult_87_CARRYB_42__16_), .CI(u5_mult_87_SUMB_42__17_), .CO(
        u5_mult_87_CARRYB_43__16_), .S(u5_mult_87_SUMB_43__16_) );
  FA_X1 u5_mult_87_S2_43_15 ( .A(u5_mult_87_ab_43__15_), .B(
        u5_mult_87_CARRYB_42__15_), .CI(u5_mult_87_SUMB_42__16_), .CO(
        u5_mult_87_CARRYB_43__15_), .S(u5_mult_87_SUMB_43__15_) );
  FA_X1 u5_mult_87_S2_43_14 ( .A(u5_mult_87_ab_43__14_), .B(
        u5_mult_87_CARRYB_42__14_), .CI(u5_mult_87_SUMB_42__15_), .CO(
        u5_mult_87_CARRYB_43__14_), .S(u5_mult_87_SUMB_43__14_) );
  FA_X1 u5_mult_87_S2_43_13 ( .A(u5_mult_87_ab_43__13_), .B(
        u5_mult_87_CARRYB_42__13_), .CI(u5_mult_87_SUMB_42__14_), .CO(
        u5_mult_87_CARRYB_43__13_), .S(u5_mult_87_SUMB_43__13_) );
  FA_X1 u5_mult_87_S2_43_12 ( .A(u5_mult_87_ab_43__12_), .B(
        u5_mult_87_CARRYB_42__12_), .CI(u5_mult_87_SUMB_42__13_), .CO(
        u5_mult_87_CARRYB_43__12_), .S(u5_mult_87_SUMB_43__12_) );
  FA_X1 u5_mult_87_S2_43_11 ( .A(u5_mult_87_ab_43__11_), .B(
        u5_mult_87_CARRYB_42__11_), .CI(u5_mult_87_SUMB_42__12_), .CO(
        u5_mult_87_CARRYB_43__11_), .S(u5_mult_87_SUMB_43__11_) );
  FA_X1 u5_mult_87_S2_43_10 ( .A(u5_mult_87_ab_43__10_), .B(
        u5_mult_87_CARRYB_42__10_), .CI(u5_mult_87_SUMB_42__11_), .CO(
        u5_mult_87_CARRYB_43__10_), .S(u5_mult_87_SUMB_43__10_) );
  FA_X1 u5_mult_87_S2_43_9 ( .A(u5_mult_87_ab_43__9_), .B(
        u5_mult_87_CARRYB_42__9_), .CI(u5_mult_87_SUMB_42__10_), .CO(
        u5_mult_87_CARRYB_43__9_), .S(u5_mult_87_SUMB_43__9_) );
  FA_X1 u5_mult_87_S2_43_8 ( .A(u5_mult_87_ab_43__8_), .B(
        u5_mult_87_CARRYB_42__8_), .CI(u5_mult_87_SUMB_42__9_), .CO(
        u5_mult_87_CARRYB_43__8_), .S(u5_mult_87_SUMB_43__8_) );
  FA_X1 u5_mult_87_S2_43_7 ( .A(u5_mult_87_ab_43__7_), .B(
        u5_mult_87_CARRYB_42__7_), .CI(u5_mult_87_SUMB_42__8_), .CO(
        u5_mult_87_CARRYB_43__7_), .S(u5_mult_87_SUMB_43__7_) );
  FA_X1 u5_mult_87_S2_43_6 ( .A(u5_mult_87_ab_43__6_), .B(
        u5_mult_87_CARRYB_42__6_), .CI(u5_mult_87_SUMB_42__7_), .CO(
        u5_mult_87_CARRYB_43__6_), .S(u5_mult_87_SUMB_43__6_) );
  FA_X1 u5_mult_87_S2_43_5 ( .A(u5_mult_87_ab_43__5_), .B(
        u5_mult_87_CARRYB_42__5_), .CI(u5_mult_87_SUMB_42__6_), .CO(
        u5_mult_87_CARRYB_43__5_), .S(u5_mult_87_SUMB_43__5_) );
  FA_X1 u5_mult_87_S2_43_4 ( .A(u5_mult_87_ab_43__4_), .B(
        u5_mult_87_CARRYB_42__4_), .CI(u5_mult_87_SUMB_42__5_), .CO(
        u5_mult_87_CARRYB_43__4_), .S(u5_mult_87_SUMB_43__4_) );
  FA_X1 u5_mult_87_S2_43_3 ( .A(u5_mult_87_ab_43__3_), .B(
        u5_mult_87_CARRYB_42__3_), .CI(u5_mult_87_SUMB_42__4_), .CO(
        u5_mult_87_CARRYB_43__3_), .S(u5_mult_87_SUMB_43__3_) );
  FA_X1 u5_mult_87_S2_43_2 ( .A(u5_mult_87_ab_43__2_), .B(
        u5_mult_87_CARRYB_42__2_), .CI(u5_mult_87_SUMB_42__3_), .CO(
        u5_mult_87_CARRYB_43__2_), .S(u5_mult_87_SUMB_43__2_) );
  FA_X1 u5_mult_87_S2_43_1 ( .A(u5_mult_87_ab_43__1_), .B(
        u5_mult_87_CARRYB_42__1_), .CI(u5_mult_87_SUMB_42__2_), .CO(
        u5_mult_87_CARRYB_43__1_), .S(u5_mult_87_SUMB_43__1_) );
  FA_X1 u5_mult_87_S1_43_0 ( .A(u5_mult_87_ab_43__0_), .B(
        u5_mult_87_CARRYB_42__0_), .CI(u5_mult_87_SUMB_42__1_), .CO(
        u5_mult_87_CARRYB_43__0_), .S(u5_N43) );
  FA_X1 u5_mult_87_S3_44_51 ( .A(u5_mult_87_ab_44__51_), .B(
        u5_mult_87_CARRYB_43__51_), .CI(u5_mult_87_ab_43__52_), .CO(
        u5_mult_87_CARRYB_44__51_), .S(u5_mult_87_SUMB_44__51_) );
  FA_X1 u5_mult_87_S2_44_50 ( .A(u5_mult_87_ab_44__50_), .B(
        u5_mult_87_CARRYB_43__50_), .CI(u5_mult_87_SUMB_43__51_), .CO(
        u5_mult_87_CARRYB_44__50_), .S(u5_mult_87_SUMB_44__50_) );
  FA_X1 u5_mult_87_S2_44_49 ( .A(u5_mult_87_ab_44__49_), .B(
        u5_mult_87_CARRYB_43__49_), .CI(u5_mult_87_SUMB_43__50_), .CO(
        u5_mult_87_CARRYB_44__49_), .S(u5_mult_87_SUMB_44__49_) );
  FA_X1 u5_mult_87_S2_44_48 ( .A(u5_mult_87_ab_44__48_), .B(
        u5_mult_87_CARRYB_43__48_), .CI(u5_mult_87_SUMB_43__49_), .CO(
        u5_mult_87_CARRYB_44__48_), .S(u5_mult_87_SUMB_44__48_) );
  FA_X1 u5_mult_87_S2_44_47 ( .A(u5_mult_87_ab_44__47_), .B(
        u5_mult_87_CARRYB_43__47_), .CI(u5_mult_87_SUMB_43__48_), .CO(
        u5_mult_87_CARRYB_44__47_), .S(u5_mult_87_SUMB_44__47_) );
  FA_X1 u5_mult_87_S2_44_46 ( .A(u5_mult_87_ab_44__46_), .B(
        u5_mult_87_CARRYB_43__46_), .CI(u5_mult_87_SUMB_43__47_), .CO(
        u5_mult_87_CARRYB_44__46_), .S(u5_mult_87_SUMB_44__46_) );
  FA_X1 u5_mult_87_S2_44_45 ( .A(u5_mult_87_ab_44__45_), .B(
        u5_mult_87_CARRYB_43__45_), .CI(u5_mult_87_SUMB_43__46_), .CO(
        u5_mult_87_CARRYB_44__45_), .S(u5_mult_87_SUMB_44__45_) );
  FA_X1 u5_mult_87_S2_44_44 ( .A(u5_mult_87_ab_44__44_), .B(
        u5_mult_87_CARRYB_43__44_), .CI(u5_mult_87_SUMB_43__45_), .CO(
        u5_mult_87_CARRYB_44__44_), .S(u5_mult_87_SUMB_44__44_) );
  FA_X1 u5_mult_87_S2_44_43 ( .A(u5_mult_87_ab_44__43_), .B(
        u5_mult_87_CARRYB_43__43_), .CI(u5_mult_87_SUMB_43__44_), .CO(
        u5_mult_87_CARRYB_44__43_), .S(u5_mult_87_SUMB_44__43_) );
  FA_X1 u5_mult_87_S2_44_42 ( .A(u5_mult_87_ab_44__42_), .B(
        u5_mult_87_CARRYB_43__42_), .CI(u5_mult_87_SUMB_43__43_), .CO(
        u5_mult_87_CARRYB_44__42_), .S(u5_mult_87_SUMB_44__42_) );
  FA_X1 u5_mult_87_S2_44_41 ( .A(u5_mult_87_ab_44__41_), .B(
        u5_mult_87_CARRYB_43__41_), .CI(u5_mult_87_SUMB_43__42_), .CO(
        u5_mult_87_CARRYB_44__41_), .S(u5_mult_87_SUMB_44__41_) );
  FA_X1 u5_mult_87_S2_44_40 ( .A(u5_mult_87_ab_44__40_), .B(
        u5_mult_87_CARRYB_43__40_), .CI(u5_mult_87_SUMB_43__41_), .CO(
        u5_mult_87_CARRYB_44__40_), .S(u5_mult_87_SUMB_44__40_) );
  FA_X1 u5_mult_87_S2_44_39 ( .A(u5_mult_87_ab_44__39_), .B(
        u5_mult_87_CARRYB_43__39_), .CI(u5_mult_87_SUMB_43__40_), .CO(
        u5_mult_87_CARRYB_44__39_), .S(u5_mult_87_SUMB_44__39_) );
  FA_X1 u5_mult_87_S2_44_38 ( .A(u5_mult_87_ab_44__38_), .B(
        u5_mult_87_CARRYB_43__38_), .CI(u5_mult_87_SUMB_43__39_), .CO(
        u5_mult_87_CARRYB_44__38_), .S(u5_mult_87_SUMB_44__38_) );
  FA_X1 u5_mult_87_S2_44_37 ( .A(u5_mult_87_ab_44__37_), .B(
        u5_mult_87_CARRYB_43__37_), .CI(u5_mult_87_SUMB_43__38_), .CO(
        u5_mult_87_CARRYB_44__37_), .S(u5_mult_87_SUMB_44__37_) );
  FA_X1 u5_mult_87_S2_44_36 ( .A(u5_mult_87_ab_44__36_), .B(
        u5_mult_87_CARRYB_43__36_), .CI(u5_mult_87_SUMB_43__37_), .CO(
        u5_mult_87_CARRYB_44__36_), .S(u5_mult_87_SUMB_44__36_) );
  FA_X1 u5_mult_87_S2_44_35 ( .A(u5_mult_87_ab_44__35_), .B(
        u5_mult_87_CARRYB_43__35_), .CI(u5_mult_87_SUMB_43__36_), .CO(
        u5_mult_87_CARRYB_44__35_), .S(u5_mult_87_SUMB_44__35_) );
  FA_X1 u5_mult_87_S2_44_34 ( .A(u5_mult_87_ab_44__34_), .B(
        u5_mult_87_CARRYB_43__34_), .CI(u5_mult_87_SUMB_43__35_), .CO(
        u5_mult_87_CARRYB_44__34_), .S(u5_mult_87_SUMB_44__34_) );
  FA_X1 u5_mult_87_S2_44_33 ( .A(u5_mult_87_ab_44__33_), .B(
        u5_mult_87_CARRYB_43__33_), .CI(u5_mult_87_SUMB_43__34_), .CO(
        u5_mult_87_CARRYB_44__33_), .S(u5_mult_87_SUMB_44__33_) );
  FA_X1 u5_mult_87_S2_44_32 ( .A(u5_mult_87_ab_44__32_), .B(
        u5_mult_87_CARRYB_43__32_), .CI(u5_mult_87_SUMB_43__33_), .CO(
        u5_mult_87_CARRYB_44__32_), .S(u5_mult_87_SUMB_44__32_) );
  FA_X1 u5_mult_87_S2_44_31 ( .A(u5_mult_87_ab_44__31_), .B(
        u5_mult_87_CARRYB_43__31_), .CI(u5_mult_87_SUMB_43__32_), .CO(
        u5_mult_87_CARRYB_44__31_), .S(u5_mult_87_SUMB_44__31_) );
  FA_X1 u5_mult_87_S2_44_30 ( .A(u5_mult_87_ab_44__30_), .B(
        u5_mult_87_CARRYB_43__30_), .CI(u5_mult_87_SUMB_43__31_), .CO(
        u5_mult_87_CARRYB_44__30_), .S(u5_mult_87_SUMB_44__30_) );
  FA_X1 u5_mult_87_S2_44_29 ( .A(u5_mult_87_ab_44__29_), .B(
        u5_mult_87_CARRYB_43__29_), .CI(u5_mult_87_SUMB_43__30_), .CO(
        u5_mult_87_CARRYB_44__29_), .S(u5_mult_87_SUMB_44__29_) );
  FA_X1 u5_mult_87_S2_44_28 ( .A(u5_mult_87_ab_44__28_), .B(
        u5_mult_87_CARRYB_43__28_), .CI(u5_mult_87_SUMB_43__29_), .CO(
        u5_mult_87_CARRYB_44__28_), .S(u5_mult_87_SUMB_44__28_) );
  FA_X1 u5_mult_87_S2_44_27 ( .A(u5_mult_87_ab_44__27_), .B(
        u5_mult_87_CARRYB_43__27_), .CI(u5_mult_87_SUMB_43__28_), .CO(
        u5_mult_87_CARRYB_44__27_), .S(u5_mult_87_SUMB_44__27_) );
  FA_X1 u5_mult_87_S2_44_26 ( .A(u5_mult_87_ab_44__26_), .B(
        u5_mult_87_CARRYB_43__26_), .CI(u5_mult_87_SUMB_43__27_), .CO(
        u5_mult_87_CARRYB_44__26_), .S(u5_mult_87_SUMB_44__26_) );
  FA_X1 u5_mult_87_S2_44_25 ( .A(u5_mult_87_ab_44__25_), .B(
        u5_mult_87_CARRYB_43__25_), .CI(u5_mult_87_SUMB_43__26_), .CO(
        u5_mult_87_CARRYB_44__25_), .S(u5_mult_87_SUMB_44__25_) );
  FA_X1 u5_mult_87_S2_44_24 ( .A(u5_mult_87_ab_44__24_), .B(
        u5_mult_87_CARRYB_43__24_), .CI(u5_mult_87_SUMB_43__25_), .CO(
        u5_mult_87_CARRYB_44__24_), .S(u5_mult_87_SUMB_44__24_) );
  FA_X1 u5_mult_87_S2_44_23 ( .A(u5_mult_87_ab_44__23_), .B(
        u5_mult_87_CARRYB_43__23_), .CI(u5_mult_87_SUMB_43__24_), .CO(
        u5_mult_87_CARRYB_44__23_), .S(u5_mult_87_SUMB_44__23_) );
  FA_X1 u5_mult_87_S2_44_22 ( .A(u5_mult_87_ab_44__22_), .B(
        u5_mult_87_CARRYB_43__22_), .CI(u5_mult_87_SUMB_43__23_), .CO(
        u5_mult_87_CARRYB_44__22_), .S(u5_mult_87_SUMB_44__22_) );
  FA_X1 u5_mult_87_S2_44_21 ( .A(u5_mult_87_ab_44__21_), .B(
        u5_mult_87_CARRYB_43__21_), .CI(u5_mult_87_SUMB_43__22_), .CO(
        u5_mult_87_CARRYB_44__21_), .S(u5_mult_87_SUMB_44__21_) );
  FA_X1 u5_mult_87_S2_44_20 ( .A(u5_mult_87_ab_44__20_), .B(
        u5_mult_87_CARRYB_43__20_), .CI(u5_mult_87_SUMB_43__21_), .CO(
        u5_mult_87_CARRYB_44__20_), .S(u5_mult_87_SUMB_44__20_) );
  FA_X1 u5_mult_87_S2_44_19 ( .A(u5_mult_87_ab_44__19_), .B(
        u5_mult_87_CARRYB_43__19_), .CI(u5_mult_87_SUMB_43__20_), .CO(
        u5_mult_87_CARRYB_44__19_), .S(u5_mult_87_SUMB_44__19_) );
  FA_X1 u5_mult_87_S2_44_18 ( .A(u5_mult_87_ab_44__18_), .B(
        u5_mult_87_CARRYB_43__18_), .CI(u5_mult_87_SUMB_43__19_), .CO(
        u5_mult_87_CARRYB_44__18_), .S(u5_mult_87_SUMB_44__18_) );
  FA_X1 u5_mult_87_S2_44_17 ( .A(u5_mult_87_ab_44__17_), .B(
        u5_mult_87_CARRYB_43__17_), .CI(u5_mult_87_SUMB_43__18_), .CO(
        u5_mult_87_CARRYB_44__17_), .S(u5_mult_87_SUMB_44__17_) );
  FA_X1 u5_mult_87_S2_44_16 ( .A(u5_mult_87_ab_44__16_), .B(
        u5_mult_87_CARRYB_43__16_), .CI(u5_mult_87_SUMB_43__17_), .CO(
        u5_mult_87_CARRYB_44__16_), .S(u5_mult_87_SUMB_44__16_) );
  FA_X1 u5_mult_87_S2_44_15 ( .A(u5_mult_87_ab_44__15_), .B(
        u5_mult_87_CARRYB_43__15_), .CI(u5_mult_87_SUMB_43__16_), .CO(
        u5_mult_87_CARRYB_44__15_), .S(u5_mult_87_SUMB_44__15_) );
  FA_X1 u5_mult_87_S2_44_14 ( .A(u5_mult_87_ab_44__14_), .B(
        u5_mult_87_CARRYB_43__14_), .CI(u5_mult_87_SUMB_43__15_), .CO(
        u5_mult_87_CARRYB_44__14_), .S(u5_mult_87_SUMB_44__14_) );
  FA_X1 u5_mult_87_S2_44_13 ( .A(u5_mult_87_ab_44__13_), .B(
        u5_mult_87_CARRYB_43__13_), .CI(u5_mult_87_SUMB_43__14_), .CO(
        u5_mult_87_CARRYB_44__13_), .S(u5_mult_87_SUMB_44__13_) );
  FA_X1 u5_mult_87_S2_44_12 ( .A(u5_mult_87_ab_44__12_), .B(
        u5_mult_87_CARRYB_43__12_), .CI(u5_mult_87_SUMB_43__13_), .CO(
        u5_mult_87_CARRYB_44__12_), .S(u5_mult_87_SUMB_44__12_) );
  FA_X1 u5_mult_87_S2_44_11 ( .A(u5_mult_87_ab_44__11_), .B(
        u5_mult_87_CARRYB_43__11_), .CI(u5_mult_87_SUMB_43__12_), .CO(
        u5_mult_87_CARRYB_44__11_), .S(u5_mult_87_SUMB_44__11_) );
  FA_X1 u5_mult_87_S2_44_10 ( .A(u5_mult_87_ab_44__10_), .B(
        u5_mult_87_CARRYB_43__10_), .CI(u5_mult_87_SUMB_43__11_), .CO(
        u5_mult_87_CARRYB_44__10_), .S(u5_mult_87_SUMB_44__10_) );
  FA_X1 u5_mult_87_S2_44_9 ( .A(u5_mult_87_ab_44__9_), .B(
        u5_mult_87_CARRYB_43__9_), .CI(u5_mult_87_SUMB_43__10_), .CO(
        u5_mult_87_CARRYB_44__9_), .S(u5_mult_87_SUMB_44__9_) );
  FA_X1 u5_mult_87_S2_44_8 ( .A(u5_mult_87_ab_44__8_), .B(
        u5_mult_87_CARRYB_43__8_), .CI(u5_mult_87_SUMB_43__9_), .CO(
        u5_mult_87_CARRYB_44__8_), .S(u5_mult_87_SUMB_44__8_) );
  FA_X1 u5_mult_87_S2_44_7 ( .A(u5_mult_87_ab_44__7_), .B(
        u5_mult_87_CARRYB_43__7_), .CI(u5_mult_87_SUMB_43__8_), .CO(
        u5_mult_87_CARRYB_44__7_), .S(u5_mult_87_SUMB_44__7_) );
  FA_X1 u5_mult_87_S2_44_6 ( .A(u5_mult_87_ab_44__6_), .B(
        u5_mult_87_CARRYB_43__6_), .CI(u5_mult_87_SUMB_43__7_), .CO(
        u5_mult_87_CARRYB_44__6_), .S(u5_mult_87_SUMB_44__6_) );
  FA_X1 u5_mult_87_S2_44_5 ( .A(u5_mult_87_ab_44__5_), .B(
        u5_mult_87_CARRYB_43__5_), .CI(u5_mult_87_SUMB_43__6_), .CO(
        u5_mult_87_CARRYB_44__5_), .S(u5_mult_87_SUMB_44__5_) );
  FA_X1 u5_mult_87_S2_44_4 ( .A(u5_mult_87_ab_44__4_), .B(
        u5_mult_87_CARRYB_43__4_), .CI(u5_mult_87_SUMB_43__5_), .CO(
        u5_mult_87_CARRYB_44__4_), .S(u5_mult_87_SUMB_44__4_) );
  FA_X1 u5_mult_87_S2_44_3 ( .A(u5_mult_87_ab_44__3_), .B(
        u5_mult_87_CARRYB_43__3_), .CI(u5_mult_87_SUMB_43__4_), .CO(
        u5_mult_87_CARRYB_44__3_), .S(u5_mult_87_SUMB_44__3_) );
  FA_X1 u5_mult_87_S2_44_2 ( .A(u5_mult_87_ab_44__2_), .B(
        u5_mult_87_CARRYB_43__2_), .CI(u5_mult_87_SUMB_43__3_), .CO(
        u5_mult_87_CARRYB_44__2_), .S(u5_mult_87_SUMB_44__2_) );
  FA_X1 u5_mult_87_S2_44_1 ( .A(u5_mult_87_ab_44__1_), .B(
        u5_mult_87_CARRYB_43__1_), .CI(u5_mult_87_SUMB_43__2_), .CO(
        u5_mult_87_CARRYB_44__1_), .S(u5_mult_87_SUMB_44__1_) );
  FA_X1 u5_mult_87_S1_44_0 ( .A(u5_mult_87_ab_44__0_), .B(
        u5_mult_87_CARRYB_43__0_), .CI(u5_mult_87_SUMB_43__1_), .CO(
        u5_mult_87_CARRYB_44__0_), .S(u5_N44) );
  FA_X1 u5_mult_87_S3_45_51 ( .A(u5_mult_87_ab_45__51_), .B(
        u5_mult_87_CARRYB_44__51_), .CI(u5_mult_87_ab_44__52_), .CO(
        u5_mult_87_CARRYB_45__51_), .S(u5_mult_87_SUMB_45__51_) );
  FA_X1 u5_mult_87_S2_45_50 ( .A(u5_mult_87_ab_45__50_), .B(
        u5_mult_87_CARRYB_44__50_), .CI(u5_mult_87_SUMB_44__51_), .CO(
        u5_mult_87_CARRYB_45__50_), .S(u5_mult_87_SUMB_45__50_) );
  FA_X1 u5_mult_87_S2_45_49 ( .A(u5_mult_87_ab_45__49_), .B(
        u5_mult_87_CARRYB_44__49_), .CI(u5_mult_87_SUMB_44__50_), .CO(
        u5_mult_87_CARRYB_45__49_), .S(u5_mult_87_SUMB_45__49_) );
  FA_X1 u5_mult_87_S2_45_48 ( .A(u5_mult_87_ab_45__48_), .B(
        u5_mult_87_CARRYB_44__48_), .CI(u5_mult_87_SUMB_44__49_), .CO(
        u5_mult_87_CARRYB_45__48_), .S(u5_mult_87_SUMB_45__48_) );
  FA_X1 u5_mult_87_S2_45_47 ( .A(u5_mult_87_ab_45__47_), .B(
        u5_mult_87_CARRYB_44__47_), .CI(u5_mult_87_SUMB_44__48_), .CO(
        u5_mult_87_CARRYB_45__47_), .S(u5_mult_87_SUMB_45__47_) );
  FA_X1 u5_mult_87_S2_45_46 ( .A(u5_mult_87_ab_45__46_), .B(
        u5_mult_87_CARRYB_44__46_), .CI(u5_mult_87_SUMB_44__47_), .CO(
        u5_mult_87_CARRYB_45__46_), .S(u5_mult_87_SUMB_45__46_) );
  FA_X1 u5_mult_87_S2_45_45 ( .A(u5_mult_87_ab_45__45_), .B(
        u5_mult_87_CARRYB_44__45_), .CI(u5_mult_87_SUMB_44__46_), .CO(
        u5_mult_87_CARRYB_45__45_), .S(u5_mult_87_SUMB_45__45_) );
  FA_X1 u5_mult_87_S2_45_44 ( .A(u5_mult_87_ab_45__44_), .B(
        u5_mult_87_CARRYB_44__44_), .CI(u5_mult_87_SUMB_44__45_), .CO(
        u5_mult_87_CARRYB_45__44_), .S(u5_mult_87_SUMB_45__44_) );
  FA_X1 u5_mult_87_S2_45_43 ( .A(u5_mult_87_ab_45__43_), .B(
        u5_mult_87_CARRYB_44__43_), .CI(u5_mult_87_SUMB_44__44_), .CO(
        u5_mult_87_CARRYB_45__43_), .S(u5_mult_87_SUMB_45__43_) );
  FA_X1 u5_mult_87_S2_45_42 ( .A(u5_mult_87_ab_45__42_), .B(
        u5_mult_87_CARRYB_44__42_), .CI(u5_mult_87_SUMB_44__43_), .CO(
        u5_mult_87_CARRYB_45__42_), .S(u5_mult_87_SUMB_45__42_) );
  FA_X1 u5_mult_87_S2_45_41 ( .A(u5_mult_87_ab_45__41_), .B(
        u5_mult_87_CARRYB_44__41_), .CI(u5_mult_87_SUMB_44__42_), .CO(
        u5_mult_87_CARRYB_45__41_), .S(u5_mult_87_SUMB_45__41_) );
  FA_X1 u5_mult_87_S2_45_40 ( .A(u5_mult_87_ab_45__40_), .B(
        u5_mult_87_CARRYB_44__40_), .CI(u5_mult_87_SUMB_44__41_), .CO(
        u5_mult_87_CARRYB_45__40_), .S(u5_mult_87_SUMB_45__40_) );
  FA_X1 u5_mult_87_S2_45_39 ( .A(u5_mult_87_ab_45__39_), .B(
        u5_mult_87_CARRYB_44__39_), .CI(u5_mult_87_SUMB_44__40_), .CO(
        u5_mult_87_CARRYB_45__39_), .S(u5_mult_87_SUMB_45__39_) );
  FA_X1 u5_mult_87_S2_45_38 ( .A(u5_mult_87_ab_45__38_), .B(
        u5_mult_87_CARRYB_44__38_), .CI(u5_mult_87_SUMB_44__39_), .CO(
        u5_mult_87_CARRYB_45__38_), .S(u5_mult_87_SUMB_45__38_) );
  FA_X1 u5_mult_87_S2_45_37 ( .A(u5_mult_87_ab_45__37_), .B(
        u5_mult_87_CARRYB_44__37_), .CI(u5_mult_87_SUMB_44__38_), .CO(
        u5_mult_87_CARRYB_45__37_), .S(u5_mult_87_SUMB_45__37_) );
  FA_X1 u5_mult_87_S2_45_36 ( .A(u5_mult_87_ab_45__36_), .B(
        u5_mult_87_CARRYB_44__36_), .CI(u5_mult_87_SUMB_44__37_), .CO(
        u5_mult_87_CARRYB_45__36_), .S(u5_mult_87_SUMB_45__36_) );
  FA_X1 u5_mult_87_S2_45_35 ( .A(u5_mult_87_ab_45__35_), .B(
        u5_mult_87_CARRYB_44__35_), .CI(u5_mult_87_SUMB_44__36_), .CO(
        u5_mult_87_CARRYB_45__35_), .S(u5_mult_87_SUMB_45__35_) );
  FA_X1 u5_mult_87_S2_45_34 ( .A(u5_mult_87_ab_45__34_), .B(
        u5_mult_87_CARRYB_44__34_), .CI(u5_mult_87_SUMB_44__35_), .CO(
        u5_mult_87_CARRYB_45__34_), .S(u5_mult_87_SUMB_45__34_) );
  FA_X1 u5_mult_87_S2_45_33 ( .A(u5_mult_87_ab_45__33_), .B(
        u5_mult_87_CARRYB_44__33_), .CI(u5_mult_87_SUMB_44__34_), .CO(
        u5_mult_87_CARRYB_45__33_), .S(u5_mult_87_SUMB_45__33_) );
  FA_X1 u5_mult_87_S2_45_32 ( .A(u5_mult_87_ab_45__32_), .B(
        u5_mult_87_CARRYB_44__32_), .CI(u5_mult_87_SUMB_44__33_), .CO(
        u5_mult_87_CARRYB_45__32_), .S(u5_mult_87_SUMB_45__32_) );
  FA_X1 u5_mult_87_S2_45_31 ( .A(u5_mult_87_ab_45__31_), .B(
        u5_mult_87_CARRYB_44__31_), .CI(u5_mult_87_SUMB_44__32_), .CO(
        u5_mult_87_CARRYB_45__31_), .S(u5_mult_87_SUMB_45__31_) );
  FA_X1 u5_mult_87_S2_45_30 ( .A(u5_mult_87_ab_45__30_), .B(
        u5_mult_87_CARRYB_44__30_), .CI(u5_mult_87_SUMB_44__31_), .CO(
        u5_mult_87_CARRYB_45__30_), .S(u5_mult_87_SUMB_45__30_) );
  FA_X1 u5_mult_87_S2_45_29 ( .A(u5_mult_87_ab_45__29_), .B(
        u5_mult_87_CARRYB_44__29_), .CI(u5_mult_87_SUMB_44__30_), .CO(
        u5_mult_87_CARRYB_45__29_), .S(u5_mult_87_SUMB_45__29_) );
  FA_X1 u5_mult_87_S2_45_28 ( .A(u5_mult_87_ab_45__28_), .B(
        u5_mult_87_CARRYB_44__28_), .CI(u5_mult_87_SUMB_44__29_), .CO(
        u5_mult_87_CARRYB_45__28_), .S(u5_mult_87_SUMB_45__28_) );
  FA_X1 u5_mult_87_S2_45_27 ( .A(u5_mult_87_ab_45__27_), .B(
        u5_mult_87_CARRYB_44__27_), .CI(u5_mult_87_SUMB_44__28_), .CO(
        u5_mult_87_CARRYB_45__27_), .S(u5_mult_87_SUMB_45__27_) );
  FA_X1 u5_mult_87_S2_45_26 ( .A(u5_mult_87_ab_45__26_), .B(
        u5_mult_87_CARRYB_44__26_), .CI(u5_mult_87_SUMB_44__27_), .CO(
        u5_mult_87_CARRYB_45__26_), .S(u5_mult_87_SUMB_45__26_) );
  FA_X1 u5_mult_87_S2_45_25 ( .A(u5_mult_87_ab_45__25_), .B(
        u5_mult_87_CARRYB_44__25_), .CI(u5_mult_87_SUMB_44__26_), .CO(
        u5_mult_87_CARRYB_45__25_), .S(u5_mult_87_SUMB_45__25_) );
  FA_X1 u5_mult_87_S2_45_24 ( .A(u5_mult_87_ab_45__24_), .B(
        u5_mult_87_CARRYB_44__24_), .CI(u5_mult_87_SUMB_44__25_), .CO(
        u5_mult_87_CARRYB_45__24_), .S(u5_mult_87_SUMB_45__24_) );
  FA_X1 u5_mult_87_S2_45_23 ( .A(u5_mult_87_ab_45__23_), .B(
        u5_mult_87_CARRYB_44__23_), .CI(u5_mult_87_SUMB_44__24_), .CO(
        u5_mult_87_CARRYB_45__23_), .S(u5_mult_87_SUMB_45__23_) );
  FA_X1 u5_mult_87_S2_45_22 ( .A(u5_mult_87_ab_45__22_), .B(
        u5_mult_87_CARRYB_44__22_), .CI(u5_mult_87_SUMB_44__23_), .CO(
        u5_mult_87_CARRYB_45__22_), .S(u5_mult_87_SUMB_45__22_) );
  FA_X1 u5_mult_87_S2_45_21 ( .A(u5_mult_87_ab_45__21_), .B(
        u5_mult_87_CARRYB_44__21_), .CI(u5_mult_87_SUMB_44__22_), .CO(
        u5_mult_87_CARRYB_45__21_), .S(u5_mult_87_SUMB_45__21_) );
  FA_X1 u5_mult_87_S2_45_20 ( .A(u5_mult_87_ab_45__20_), .B(
        u5_mult_87_CARRYB_44__20_), .CI(u5_mult_87_SUMB_44__21_), .CO(
        u5_mult_87_CARRYB_45__20_), .S(u5_mult_87_SUMB_45__20_) );
  FA_X1 u5_mult_87_S2_45_19 ( .A(u5_mult_87_ab_45__19_), .B(
        u5_mult_87_CARRYB_44__19_), .CI(u5_mult_87_SUMB_44__20_), .CO(
        u5_mult_87_CARRYB_45__19_), .S(u5_mult_87_SUMB_45__19_) );
  FA_X1 u5_mult_87_S2_45_18 ( .A(u5_mult_87_ab_45__18_), .B(
        u5_mult_87_CARRYB_44__18_), .CI(u5_mult_87_SUMB_44__19_), .CO(
        u5_mult_87_CARRYB_45__18_), .S(u5_mult_87_SUMB_45__18_) );
  FA_X1 u5_mult_87_S2_45_17 ( .A(u5_mult_87_ab_45__17_), .B(
        u5_mult_87_CARRYB_44__17_), .CI(u5_mult_87_SUMB_44__18_), .CO(
        u5_mult_87_CARRYB_45__17_), .S(u5_mult_87_SUMB_45__17_) );
  FA_X1 u5_mult_87_S2_45_16 ( .A(u5_mult_87_ab_45__16_), .B(
        u5_mult_87_CARRYB_44__16_), .CI(u5_mult_87_SUMB_44__17_), .CO(
        u5_mult_87_CARRYB_45__16_), .S(u5_mult_87_SUMB_45__16_) );
  FA_X1 u5_mult_87_S2_45_15 ( .A(u5_mult_87_ab_45__15_), .B(
        u5_mult_87_CARRYB_44__15_), .CI(u5_mult_87_SUMB_44__16_), .CO(
        u5_mult_87_CARRYB_45__15_), .S(u5_mult_87_SUMB_45__15_) );
  FA_X1 u5_mult_87_S2_45_14 ( .A(u5_mult_87_ab_45__14_), .B(
        u5_mult_87_CARRYB_44__14_), .CI(u5_mult_87_SUMB_44__15_), .CO(
        u5_mult_87_CARRYB_45__14_), .S(u5_mult_87_SUMB_45__14_) );
  FA_X1 u5_mult_87_S2_45_13 ( .A(u5_mult_87_ab_45__13_), .B(
        u5_mult_87_CARRYB_44__13_), .CI(u5_mult_87_SUMB_44__14_), .CO(
        u5_mult_87_CARRYB_45__13_), .S(u5_mult_87_SUMB_45__13_) );
  FA_X1 u5_mult_87_S2_45_12 ( .A(u5_mult_87_ab_45__12_), .B(
        u5_mult_87_CARRYB_44__12_), .CI(u5_mult_87_SUMB_44__13_), .CO(
        u5_mult_87_CARRYB_45__12_), .S(u5_mult_87_SUMB_45__12_) );
  FA_X1 u5_mult_87_S2_45_11 ( .A(u5_mult_87_ab_45__11_), .B(
        u5_mult_87_CARRYB_44__11_), .CI(u5_mult_87_SUMB_44__12_), .CO(
        u5_mult_87_CARRYB_45__11_), .S(u5_mult_87_SUMB_45__11_) );
  FA_X1 u5_mult_87_S2_45_10 ( .A(u5_mult_87_ab_45__10_), .B(
        u5_mult_87_CARRYB_44__10_), .CI(u5_mult_87_SUMB_44__11_), .CO(
        u5_mult_87_CARRYB_45__10_), .S(u5_mult_87_SUMB_45__10_) );
  FA_X1 u5_mult_87_S2_45_9 ( .A(u5_mult_87_ab_45__9_), .B(
        u5_mult_87_CARRYB_44__9_), .CI(u5_mult_87_SUMB_44__10_), .CO(
        u5_mult_87_CARRYB_45__9_), .S(u5_mult_87_SUMB_45__9_) );
  FA_X1 u5_mult_87_S2_45_8 ( .A(u5_mult_87_ab_45__8_), .B(
        u5_mult_87_CARRYB_44__8_), .CI(u5_mult_87_SUMB_44__9_), .CO(
        u5_mult_87_CARRYB_45__8_), .S(u5_mult_87_SUMB_45__8_) );
  FA_X1 u5_mult_87_S2_45_7 ( .A(u5_mult_87_ab_45__7_), .B(
        u5_mult_87_CARRYB_44__7_), .CI(u5_mult_87_SUMB_44__8_), .CO(
        u5_mult_87_CARRYB_45__7_), .S(u5_mult_87_SUMB_45__7_) );
  FA_X1 u5_mult_87_S2_45_6 ( .A(u5_mult_87_ab_45__6_), .B(
        u5_mult_87_CARRYB_44__6_), .CI(u5_mult_87_SUMB_44__7_), .CO(
        u5_mult_87_CARRYB_45__6_), .S(u5_mult_87_SUMB_45__6_) );
  FA_X1 u5_mult_87_S2_45_5 ( .A(u5_mult_87_ab_45__5_), .B(
        u5_mult_87_CARRYB_44__5_), .CI(u5_mult_87_SUMB_44__6_), .CO(
        u5_mult_87_CARRYB_45__5_), .S(u5_mult_87_SUMB_45__5_) );
  FA_X1 u5_mult_87_S2_45_4 ( .A(u5_mult_87_ab_45__4_), .B(
        u5_mult_87_CARRYB_44__4_), .CI(u5_mult_87_SUMB_44__5_), .CO(
        u5_mult_87_CARRYB_45__4_), .S(u5_mult_87_SUMB_45__4_) );
  FA_X1 u5_mult_87_S2_45_3 ( .A(u5_mult_87_ab_45__3_), .B(
        u5_mult_87_CARRYB_44__3_), .CI(u5_mult_87_SUMB_44__4_), .CO(
        u5_mult_87_CARRYB_45__3_), .S(u5_mult_87_SUMB_45__3_) );
  FA_X1 u5_mult_87_S2_45_2 ( .A(u5_mult_87_ab_45__2_), .B(
        u5_mult_87_CARRYB_44__2_), .CI(u5_mult_87_SUMB_44__3_), .CO(
        u5_mult_87_CARRYB_45__2_), .S(u5_mult_87_SUMB_45__2_) );
  FA_X1 u5_mult_87_S2_45_1 ( .A(u5_mult_87_ab_45__1_), .B(
        u5_mult_87_CARRYB_44__1_), .CI(u5_mult_87_SUMB_44__2_), .CO(
        u5_mult_87_CARRYB_45__1_), .S(u5_mult_87_SUMB_45__1_) );
  FA_X1 u5_mult_87_S1_45_0 ( .A(u5_mult_87_ab_45__0_), .B(
        u5_mult_87_CARRYB_44__0_), .CI(u5_mult_87_SUMB_44__1_), .CO(
        u5_mult_87_CARRYB_45__0_), .S(u5_N45) );
  FA_X1 u5_mult_87_S3_46_51 ( .A(u5_mult_87_ab_46__51_), .B(
        u5_mult_87_CARRYB_45__51_), .CI(u5_mult_87_ab_45__52_), .CO(
        u5_mult_87_CARRYB_46__51_), .S(u5_mult_87_SUMB_46__51_) );
  FA_X1 u5_mult_87_S2_46_50 ( .A(u5_mult_87_ab_46__50_), .B(
        u5_mult_87_CARRYB_45__50_), .CI(u5_mult_87_SUMB_45__51_), .CO(
        u5_mult_87_CARRYB_46__50_), .S(u5_mult_87_SUMB_46__50_) );
  FA_X1 u5_mult_87_S2_46_49 ( .A(u5_mult_87_ab_46__49_), .B(
        u5_mult_87_CARRYB_45__49_), .CI(u5_mult_87_SUMB_45__50_), .CO(
        u5_mult_87_CARRYB_46__49_), .S(u5_mult_87_SUMB_46__49_) );
  FA_X1 u5_mult_87_S2_46_48 ( .A(u5_mult_87_ab_46__48_), .B(
        u5_mult_87_CARRYB_45__48_), .CI(u5_mult_87_SUMB_45__49_), .CO(
        u5_mult_87_CARRYB_46__48_), .S(u5_mult_87_SUMB_46__48_) );
  FA_X1 u5_mult_87_S2_46_47 ( .A(u5_mult_87_ab_46__47_), .B(
        u5_mult_87_CARRYB_45__47_), .CI(u5_mult_87_SUMB_45__48_), .CO(
        u5_mult_87_CARRYB_46__47_), .S(u5_mult_87_SUMB_46__47_) );
  FA_X1 u5_mult_87_S2_46_46 ( .A(u5_mult_87_ab_46__46_), .B(
        u5_mult_87_CARRYB_45__46_), .CI(u5_mult_87_SUMB_45__47_), .CO(
        u5_mult_87_CARRYB_46__46_), .S(u5_mult_87_SUMB_46__46_) );
  FA_X1 u5_mult_87_S2_46_45 ( .A(u5_mult_87_ab_46__45_), .B(
        u5_mult_87_CARRYB_45__45_), .CI(u5_mult_87_SUMB_45__46_), .CO(
        u5_mult_87_CARRYB_46__45_), .S(u5_mult_87_SUMB_46__45_) );
  FA_X1 u5_mult_87_S2_46_44 ( .A(u5_mult_87_ab_46__44_), .B(
        u5_mult_87_CARRYB_45__44_), .CI(u5_mult_87_SUMB_45__45_), .CO(
        u5_mult_87_CARRYB_46__44_), .S(u5_mult_87_SUMB_46__44_) );
  FA_X1 u5_mult_87_S2_46_43 ( .A(u5_mult_87_ab_46__43_), .B(
        u5_mult_87_CARRYB_45__43_), .CI(u5_mult_87_SUMB_45__44_), .CO(
        u5_mult_87_CARRYB_46__43_), .S(u5_mult_87_SUMB_46__43_) );
  FA_X1 u5_mult_87_S2_46_42 ( .A(u5_mult_87_ab_46__42_), .B(
        u5_mult_87_CARRYB_45__42_), .CI(u5_mult_87_SUMB_45__43_), .CO(
        u5_mult_87_CARRYB_46__42_), .S(u5_mult_87_SUMB_46__42_) );
  FA_X1 u5_mult_87_S2_46_41 ( .A(u5_mult_87_ab_46__41_), .B(
        u5_mult_87_CARRYB_45__41_), .CI(u5_mult_87_SUMB_45__42_), .CO(
        u5_mult_87_CARRYB_46__41_), .S(u5_mult_87_SUMB_46__41_) );
  FA_X1 u5_mult_87_S2_46_40 ( .A(u5_mult_87_ab_46__40_), .B(
        u5_mult_87_CARRYB_45__40_), .CI(u5_mult_87_SUMB_45__41_), .CO(
        u5_mult_87_CARRYB_46__40_), .S(u5_mult_87_SUMB_46__40_) );
  FA_X1 u5_mult_87_S2_46_39 ( .A(u5_mult_87_ab_46__39_), .B(
        u5_mult_87_CARRYB_45__39_), .CI(u5_mult_87_SUMB_45__40_), .CO(
        u5_mult_87_CARRYB_46__39_), .S(u5_mult_87_SUMB_46__39_) );
  FA_X1 u5_mult_87_S2_46_38 ( .A(u5_mult_87_ab_46__38_), .B(
        u5_mult_87_CARRYB_45__38_), .CI(u5_mult_87_SUMB_45__39_), .CO(
        u5_mult_87_CARRYB_46__38_), .S(u5_mult_87_SUMB_46__38_) );
  FA_X1 u5_mult_87_S2_46_37 ( .A(u5_mult_87_ab_46__37_), .B(
        u5_mult_87_CARRYB_45__37_), .CI(u5_mult_87_SUMB_45__38_), .CO(
        u5_mult_87_CARRYB_46__37_), .S(u5_mult_87_SUMB_46__37_) );
  FA_X1 u5_mult_87_S2_46_36 ( .A(u5_mult_87_ab_46__36_), .B(
        u5_mult_87_CARRYB_45__36_), .CI(u5_mult_87_SUMB_45__37_), .CO(
        u5_mult_87_CARRYB_46__36_), .S(u5_mult_87_SUMB_46__36_) );
  FA_X1 u5_mult_87_S2_46_35 ( .A(u5_mult_87_ab_46__35_), .B(
        u5_mult_87_CARRYB_45__35_), .CI(u5_mult_87_SUMB_45__36_), .CO(
        u5_mult_87_CARRYB_46__35_), .S(u5_mult_87_SUMB_46__35_) );
  FA_X1 u5_mult_87_S2_46_34 ( .A(u5_mult_87_ab_46__34_), .B(
        u5_mult_87_CARRYB_45__34_), .CI(u5_mult_87_SUMB_45__35_), .CO(
        u5_mult_87_CARRYB_46__34_), .S(u5_mult_87_SUMB_46__34_) );
  FA_X1 u5_mult_87_S2_46_33 ( .A(u5_mult_87_ab_46__33_), .B(
        u5_mult_87_CARRYB_45__33_), .CI(u5_mult_87_SUMB_45__34_), .CO(
        u5_mult_87_CARRYB_46__33_), .S(u5_mult_87_SUMB_46__33_) );
  FA_X1 u5_mult_87_S2_46_32 ( .A(u5_mult_87_ab_46__32_), .B(
        u5_mult_87_CARRYB_45__32_), .CI(u5_mult_87_SUMB_45__33_), .CO(
        u5_mult_87_CARRYB_46__32_), .S(u5_mult_87_SUMB_46__32_) );
  FA_X1 u5_mult_87_S2_46_31 ( .A(u5_mult_87_ab_46__31_), .B(
        u5_mult_87_CARRYB_45__31_), .CI(u5_mult_87_SUMB_45__32_), .CO(
        u5_mult_87_CARRYB_46__31_), .S(u5_mult_87_SUMB_46__31_) );
  FA_X1 u5_mult_87_S2_46_30 ( .A(u5_mult_87_ab_46__30_), .B(
        u5_mult_87_CARRYB_45__30_), .CI(u5_mult_87_SUMB_45__31_), .CO(
        u5_mult_87_CARRYB_46__30_), .S(u5_mult_87_SUMB_46__30_) );
  FA_X1 u5_mult_87_S2_46_29 ( .A(u5_mult_87_ab_46__29_), .B(
        u5_mult_87_CARRYB_45__29_), .CI(u5_mult_87_SUMB_45__30_), .CO(
        u5_mult_87_CARRYB_46__29_), .S(u5_mult_87_SUMB_46__29_) );
  FA_X1 u5_mult_87_S2_46_28 ( .A(u5_mult_87_ab_46__28_), .B(
        u5_mult_87_CARRYB_45__28_), .CI(u5_mult_87_SUMB_45__29_), .CO(
        u5_mult_87_CARRYB_46__28_), .S(u5_mult_87_SUMB_46__28_) );
  FA_X1 u5_mult_87_S2_46_27 ( .A(u5_mult_87_ab_46__27_), .B(
        u5_mult_87_CARRYB_45__27_), .CI(u5_mult_87_SUMB_45__28_), .CO(
        u5_mult_87_CARRYB_46__27_), .S(u5_mult_87_SUMB_46__27_) );
  FA_X1 u5_mult_87_S2_46_26 ( .A(u5_mult_87_ab_46__26_), .B(
        u5_mult_87_CARRYB_45__26_), .CI(u5_mult_87_SUMB_45__27_), .CO(
        u5_mult_87_CARRYB_46__26_), .S(u5_mult_87_SUMB_46__26_) );
  FA_X1 u5_mult_87_S2_46_25 ( .A(u5_mult_87_ab_46__25_), .B(
        u5_mult_87_CARRYB_45__25_), .CI(u5_mult_87_SUMB_45__26_), .CO(
        u5_mult_87_CARRYB_46__25_), .S(u5_mult_87_SUMB_46__25_) );
  FA_X1 u5_mult_87_S2_46_24 ( .A(u5_mult_87_ab_46__24_), .B(
        u5_mult_87_CARRYB_45__24_), .CI(u5_mult_87_SUMB_45__25_), .CO(
        u5_mult_87_CARRYB_46__24_), .S(u5_mult_87_SUMB_46__24_) );
  FA_X1 u5_mult_87_S2_46_23 ( .A(u5_mult_87_ab_46__23_), .B(
        u5_mult_87_CARRYB_45__23_), .CI(u5_mult_87_SUMB_45__24_), .CO(
        u5_mult_87_CARRYB_46__23_), .S(u5_mult_87_SUMB_46__23_) );
  FA_X1 u5_mult_87_S2_46_22 ( .A(u5_mult_87_ab_46__22_), .B(
        u5_mult_87_CARRYB_45__22_), .CI(u5_mult_87_SUMB_45__23_), .CO(
        u5_mult_87_CARRYB_46__22_), .S(u5_mult_87_SUMB_46__22_) );
  FA_X1 u5_mult_87_S2_46_21 ( .A(u5_mult_87_ab_46__21_), .B(
        u5_mult_87_CARRYB_45__21_), .CI(u5_mult_87_SUMB_45__22_), .CO(
        u5_mult_87_CARRYB_46__21_), .S(u5_mult_87_SUMB_46__21_) );
  FA_X1 u5_mult_87_S2_46_20 ( .A(u5_mult_87_ab_46__20_), .B(
        u5_mult_87_CARRYB_45__20_), .CI(u5_mult_87_SUMB_45__21_), .CO(
        u5_mult_87_CARRYB_46__20_), .S(u5_mult_87_SUMB_46__20_) );
  FA_X1 u5_mult_87_S2_46_19 ( .A(u5_mult_87_ab_46__19_), .B(
        u5_mult_87_CARRYB_45__19_), .CI(u5_mult_87_SUMB_45__20_), .CO(
        u5_mult_87_CARRYB_46__19_), .S(u5_mult_87_SUMB_46__19_) );
  FA_X1 u5_mult_87_S2_46_18 ( .A(u5_mult_87_ab_46__18_), .B(
        u5_mult_87_CARRYB_45__18_), .CI(u5_mult_87_SUMB_45__19_), .CO(
        u5_mult_87_CARRYB_46__18_), .S(u5_mult_87_SUMB_46__18_) );
  FA_X1 u5_mult_87_S2_46_17 ( .A(u5_mult_87_ab_46__17_), .B(
        u5_mult_87_CARRYB_45__17_), .CI(u5_mult_87_SUMB_45__18_), .CO(
        u5_mult_87_CARRYB_46__17_), .S(u5_mult_87_SUMB_46__17_) );
  FA_X1 u5_mult_87_S2_46_16 ( .A(u5_mult_87_ab_46__16_), .B(
        u5_mult_87_CARRYB_45__16_), .CI(u5_mult_87_SUMB_45__17_), .CO(
        u5_mult_87_CARRYB_46__16_), .S(u5_mult_87_SUMB_46__16_) );
  FA_X1 u5_mult_87_S2_46_15 ( .A(u5_mult_87_ab_46__15_), .B(
        u5_mult_87_CARRYB_45__15_), .CI(u5_mult_87_SUMB_45__16_), .CO(
        u5_mult_87_CARRYB_46__15_), .S(u5_mult_87_SUMB_46__15_) );
  FA_X1 u5_mult_87_S2_46_14 ( .A(u5_mult_87_ab_46__14_), .B(
        u5_mult_87_CARRYB_45__14_), .CI(u5_mult_87_SUMB_45__15_), .CO(
        u5_mult_87_CARRYB_46__14_), .S(u5_mult_87_SUMB_46__14_) );
  FA_X1 u5_mult_87_S2_46_13 ( .A(u5_mult_87_ab_46__13_), .B(
        u5_mult_87_CARRYB_45__13_), .CI(u5_mult_87_SUMB_45__14_), .CO(
        u5_mult_87_CARRYB_46__13_), .S(u5_mult_87_SUMB_46__13_) );
  FA_X1 u5_mult_87_S2_46_12 ( .A(u5_mult_87_ab_46__12_), .B(
        u5_mult_87_CARRYB_45__12_), .CI(u5_mult_87_SUMB_45__13_), .CO(
        u5_mult_87_CARRYB_46__12_), .S(u5_mult_87_SUMB_46__12_) );
  FA_X1 u5_mult_87_S2_46_11 ( .A(u5_mult_87_ab_46__11_), .B(
        u5_mult_87_CARRYB_45__11_), .CI(u5_mult_87_SUMB_45__12_), .CO(
        u5_mult_87_CARRYB_46__11_), .S(u5_mult_87_SUMB_46__11_) );
  FA_X1 u5_mult_87_S2_46_10 ( .A(u5_mult_87_ab_46__10_), .B(
        u5_mult_87_CARRYB_45__10_), .CI(u5_mult_87_SUMB_45__11_), .CO(
        u5_mult_87_CARRYB_46__10_), .S(u5_mult_87_SUMB_46__10_) );
  FA_X1 u5_mult_87_S2_46_9 ( .A(u5_mult_87_ab_46__9_), .B(
        u5_mult_87_CARRYB_45__9_), .CI(u5_mult_87_SUMB_45__10_), .CO(
        u5_mult_87_CARRYB_46__9_), .S(u5_mult_87_SUMB_46__9_) );
  FA_X1 u5_mult_87_S2_46_8 ( .A(u5_mult_87_ab_46__8_), .B(
        u5_mult_87_CARRYB_45__8_), .CI(u5_mult_87_SUMB_45__9_), .CO(
        u5_mult_87_CARRYB_46__8_), .S(u5_mult_87_SUMB_46__8_) );
  FA_X1 u5_mult_87_S2_46_7 ( .A(u5_mult_87_ab_46__7_), .B(
        u5_mult_87_CARRYB_45__7_), .CI(u5_mult_87_SUMB_45__8_), .CO(
        u5_mult_87_CARRYB_46__7_), .S(u5_mult_87_SUMB_46__7_) );
  FA_X1 u5_mult_87_S2_46_6 ( .A(u5_mult_87_ab_46__6_), .B(
        u5_mult_87_CARRYB_45__6_), .CI(u5_mult_87_SUMB_45__7_), .CO(
        u5_mult_87_CARRYB_46__6_), .S(u5_mult_87_SUMB_46__6_) );
  FA_X1 u5_mult_87_S2_46_5 ( .A(u5_mult_87_ab_46__5_), .B(
        u5_mult_87_CARRYB_45__5_), .CI(u5_mult_87_SUMB_45__6_), .CO(
        u5_mult_87_CARRYB_46__5_), .S(u5_mult_87_SUMB_46__5_) );
  FA_X1 u5_mult_87_S2_46_4 ( .A(u5_mult_87_ab_46__4_), .B(
        u5_mult_87_CARRYB_45__4_), .CI(u5_mult_87_SUMB_45__5_), .CO(
        u5_mult_87_CARRYB_46__4_), .S(u5_mult_87_SUMB_46__4_) );
  FA_X1 u5_mult_87_S2_46_3 ( .A(u5_mult_87_ab_46__3_), .B(
        u5_mult_87_CARRYB_45__3_), .CI(u5_mult_87_SUMB_45__4_), .CO(
        u5_mult_87_CARRYB_46__3_), .S(u5_mult_87_SUMB_46__3_) );
  FA_X1 u5_mult_87_S2_46_2 ( .A(u5_mult_87_ab_46__2_), .B(
        u5_mult_87_CARRYB_45__2_), .CI(u5_mult_87_SUMB_45__3_), .CO(
        u5_mult_87_CARRYB_46__2_), .S(u5_mult_87_SUMB_46__2_) );
  FA_X1 u5_mult_87_S2_46_1 ( .A(u5_mult_87_ab_46__1_), .B(
        u5_mult_87_CARRYB_45__1_), .CI(u5_mult_87_SUMB_45__2_), .CO(
        u5_mult_87_CARRYB_46__1_), .S(u5_mult_87_SUMB_46__1_) );
  FA_X1 u5_mult_87_S1_46_0 ( .A(u5_mult_87_ab_46__0_), .B(
        u5_mult_87_CARRYB_45__0_), .CI(u5_mult_87_SUMB_45__1_), .CO(
        u5_mult_87_CARRYB_46__0_), .S(u5_N46) );
  FA_X1 u5_mult_87_S3_47_51 ( .A(u5_mult_87_ab_47__51_), .B(
        u5_mult_87_CARRYB_46__51_), .CI(u5_mult_87_ab_46__52_), .CO(
        u5_mult_87_CARRYB_47__51_), .S(u5_mult_87_SUMB_47__51_) );
  FA_X1 u5_mult_87_S2_47_50 ( .A(u5_mult_87_ab_47__50_), .B(
        u5_mult_87_CARRYB_46__50_), .CI(u5_mult_87_SUMB_46__51_), .CO(
        u5_mult_87_CARRYB_47__50_), .S(u5_mult_87_SUMB_47__50_) );
  FA_X1 u5_mult_87_S2_47_49 ( .A(u5_mult_87_ab_47__49_), .B(
        u5_mult_87_CARRYB_46__49_), .CI(u5_mult_87_SUMB_46__50_), .CO(
        u5_mult_87_CARRYB_47__49_), .S(u5_mult_87_SUMB_47__49_) );
  FA_X1 u5_mult_87_S2_47_48 ( .A(u5_mult_87_ab_47__48_), .B(
        u5_mult_87_CARRYB_46__48_), .CI(u5_mult_87_SUMB_46__49_), .CO(
        u5_mult_87_CARRYB_47__48_), .S(u5_mult_87_SUMB_47__48_) );
  FA_X1 u5_mult_87_S2_47_47 ( .A(u5_mult_87_ab_47__47_), .B(
        u5_mult_87_CARRYB_46__47_), .CI(u5_mult_87_SUMB_46__48_), .CO(
        u5_mult_87_CARRYB_47__47_), .S(u5_mult_87_SUMB_47__47_) );
  FA_X1 u5_mult_87_S2_47_46 ( .A(u5_mult_87_ab_47__46_), .B(
        u5_mult_87_CARRYB_46__46_), .CI(u5_mult_87_SUMB_46__47_), .CO(
        u5_mult_87_CARRYB_47__46_), .S(u5_mult_87_SUMB_47__46_) );
  FA_X1 u5_mult_87_S2_47_45 ( .A(u5_mult_87_ab_47__45_), .B(
        u5_mult_87_CARRYB_46__45_), .CI(u5_mult_87_SUMB_46__46_), .CO(
        u5_mult_87_CARRYB_47__45_), .S(u5_mult_87_SUMB_47__45_) );
  FA_X1 u5_mult_87_S2_47_44 ( .A(u5_mult_87_ab_47__44_), .B(
        u5_mult_87_CARRYB_46__44_), .CI(u5_mult_87_SUMB_46__45_), .CO(
        u5_mult_87_CARRYB_47__44_), .S(u5_mult_87_SUMB_47__44_) );
  FA_X1 u5_mult_87_S2_47_43 ( .A(u5_mult_87_ab_47__43_), .B(
        u5_mult_87_CARRYB_46__43_), .CI(u5_mult_87_SUMB_46__44_), .CO(
        u5_mult_87_CARRYB_47__43_), .S(u5_mult_87_SUMB_47__43_) );
  FA_X1 u5_mult_87_S2_47_42 ( .A(u5_mult_87_ab_47__42_), .B(
        u5_mult_87_CARRYB_46__42_), .CI(u5_mult_87_SUMB_46__43_), .CO(
        u5_mult_87_CARRYB_47__42_), .S(u5_mult_87_SUMB_47__42_) );
  FA_X1 u5_mult_87_S2_47_41 ( .A(u5_mult_87_ab_47__41_), .B(
        u5_mult_87_CARRYB_46__41_), .CI(u5_mult_87_SUMB_46__42_), .CO(
        u5_mult_87_CARRYB_47__41_), .S(u5_mult_87_SUMB_47__41_) );
  FA_X1 u5_mult_87_S2_47_40 ( .A(u5_mult_87_ab_47__40_), .B(
        u5_mult_87_CARRYB_46__40_), .CI(u5_mult_87_SUMB_46__41_), .CO(
        u5_mult_87_CARRYB_47__40_), .S(u5_mult_87_SUMB_47__40_) );
  FA_X1 u5_mult_87_S2_47_39 ( .A(u5_mult_87_ab_47__39_), .B(
        u5_mult_87_CARRYB_46__39_), .CI(u5_mult_87_SUMB_46__40_), .CO(
        u5_mult_87_CARRYB_47__39_), .S(u5_mult_87_SUMB_47__39_) );
  FA_X1 u5_mult_87_S2_47_38 ( .A(u5_mult_87_ab_47__38_), .B(
        u5_mult_87_CARRYB_46__38_), .CI(u5_mult_87_SUMB_46__39_), .CO(
        u5_mult_87_CARRYB_47__38_), .S(u5_mult_87_SUMB_47__38_) );
  FA_X1 u5_mult_87_S2_47_37 ( .A(u5_mult_87_ab_47__37_), .B(
        u5_mult_87_CARRYB_46__37_), .CI(u5_mult_87_SUMB_46__38_), .CO(
        u5_mult_87_CARRYB_47__37_), .S(u5_mult_87_SUMB_47__37_) );
  FA_X1 u5_mult_87_S2_47_36 ( .A(u5_mult_87_ab_47__36_), .B(
        u5_mult_87_CARRYB_46__36_), .CI(u5_mult_87_SUMB_46__37_), .CO(
        u5_mult_87_CARRYB_47__36_), .S(u5_mult_87_SUMB_47__36_) );
  FA_X1 u5_mult_87_S2_47_35 ( .A(u5_mult_87_ab_47__35_), .B(
        u5_mult_87_CARRYB_46__35_), .CI(u5_mult_87_SUMB_46__36_), .CO(
        u5_mult_87_CARRYB_47__35_), .S(u5_mult_87_SUMB_47__35_) );
  FA_X1 u5_mult_87_S2_47_34 ( .A(u5_mult_87_ab_47__34_), .B(
        u5_mult_87_CARRYB_46__34_), .CI(u5_mult_87_SUMB_46__35_), .CO(
        u5_mult_87_CARRYB_47__34_), .S(u5_mult_87_SUMB_47__34_) );
  FA_X1 u5_mult_87_S2_47_33 ( .A(u5_mult_87_ab_47__33_), .B(
        u5_mult_87_CARRYB_46__33_), .CI(u5_mult_87_SUMB_46__34_), .CO(
        u5_mult_87_CARRYB_47__33_), .S(u5_mult_87_SUMB_47__33_) );
  FA_X1 u5_mult_87_S2_47_32 ( .A(u5_mult_87_ab_47__32_), .B(
        u5_mult_87_CARRYB_46__32_), .CI(u5_mult_87_SUMB_46__33_), .CO(
        u5_mult_87_CARRYB_47__32_), .S(u5_mult_87_SUMB_47__32_) );
  FA_X1 u5_mult_87_S2_47_31 ( .A(u5_mult_87_ab_47__31_), .B(
        u5_mult_87_CARRYB_46__31_), .CI(u5_mult_87_SUMB_46__32_), .CO(
        u5_mult_87_CARRYB_47__31_), .S(u5_mult_87_SUMB_47__31_) );
  FA_X1 u5_mult_87_S2_47_30 ( .A(u5_mult_87_ab_47__30_), .B(
        u5_mult_87_CARRYB_46__30_), .CI(u5_mult_87_SUMB_46__31_), .CO(
        u5_mult_87_CARRYB_47__30_), .S(u5_mult_87_SUMB_47__30_) );
  FA_X1 u5_mult_87_S2_47_29 ( .A(u5_mult_87_ab_47__29_), .B(
        u5_mult_87_CARRYB_46__29_), .CI(u5_mult_87_SUMB_46__30_), .CO(
        u5_mult_87_CARRYB_47__29_), .S(u5_mult_87_SUMB_47__29_) );
  FA_X1 u5_mult_87_S2_47_28 ( .A(u5_mult_87_ab_47__28_), .B(
        u5_mult_87_CARRYB_46__28_), .CI(u5_mult_87_SUMB_46__29_), .CO(
        u5_mult_87_CARRYB_47__28_), .S(u5_mult_87_SUMB_47__28_) );
  FA_X1 u5_mult_87_S2_47_27 ( .A(u5_mult_87_ab_47__27_), .B(
        u5_mult_87_CARRYB_46__27_), .CI(u5_mult_87_SUMB_46__28_), .CO(
        u5_mult_87_CARRYB_47__27_), .S(u5_mult_87_SUMB_47__27_) );
  FA_X1 u5_mult_87_S2_47_26 ( .A(u5_mult_87_ab_47__26_), .B(
        u5_mult_87_CARRYB_46__26_), .CI(u5_mult_87_SUMB_46__27_), .CO(
        u5_mult_87_CARRYB_47__26_), .S(u5_mult_87_SUMB_47__26_) );
  FA_X1 u5_mult_87_S2_47_25 ( .A(u5_mult_87_ab_47__25_), .B(
        u5_mult_87_CARRYB_46__25_), .CI(u5_mult_87_SUMB_46__26_), .CO(
        u5_mult_87_CARRYB_47__25_), .S(u5_mult_87_SUMB_47__25_) );
  FA_X1 u5_mult_87_S2_47_24 ( .A(u5_mult_87_ab_47__24_), .B(
        u5_mult_87_CARRYB_46__24_), .CI(u5_mult_87_SUMB_46__25_), .CO(
        u5_mult_87_CARRYB_47__24_), .S(u5_mult_87_SUMB_47__24_) );
  FA_X1 u5_mult_87_S2_47_23 ( .A(u5_mult_87_ab_47__23_), .B(
        u5_mult_87_CARRYB_46__23_), .CI(u5_mult_87_SUMB_46__24_), .CO(
        u5_mult_87_CARRYB_47__23_), .S(u5_mult_87_SUMB_47__23_) );
  FA_X1 u5_mult_87_S2_47_22 ( .A(u5_mult_87_ab_47__22_), .B(
        u5_mult_87_CARRYB_46__22_), .CI(u5_mult_87_SUMB_46__23_), .CO(
        u5_mult_87_CARRYB_47__22_), .S(u5_mult_87_SUMB_47__22_) );
  FA_X1 u5_mult_87_S2_47_21 ( .A(u5_mult_87_ab_47__21_), .B(
        u5_mult_87_CARRYB_46__21_), .CI(u5_mult_87_SUMB_46__22_), .CO(
        u5_mult_87_CARRYB_47__21_), .S(u5_mult_87_SUMB_47__21_) );
  FA_X1 u5_mult_87_S2_47_20 ( .A(u5_mult_87_ab_47__20_), .B(
        u5_mult_87_CARRYB_46__20_), .CI(u5_mult_87_SUMB_46__21_), .CO(
        u5_mult_87_CARRYB_47__20_), .S(u5_mult_87_SUMB_47__20_) );
  FA_X1 u5_mult_87_S2_47_19 ( .A(u5_mult_87_ab_47__19_), .B(
        u5_mult_87_CARRYB_46__19_), .CI(u5_mult_87_SUMB_46__20_), .CO(
        u5_mult_87_CARRYB_47__19_), .S(u5_mult_87_SUMB_47__19_) );
  FA_X1 u5_mult_87_S2_47_18 ( .A(u5_mult_87_ab_47__18_), .B(
        u5_mult_87_CARRYB_46__18_), .CI(u5_mult_87_SUMB_46__19_), .CO(
        u5_mult_87_CARRYB_47__18_), .S(u5_mult_87_SUMB_47__18_) );
  FA_X1 u5_mult_87_S2_47_17 ( .A(u5_mult_87_ab_47__17_), .B(
        u5_mult_87_CARRYB_46__17_), .CI(u5_mult_87_SUMB_46__18_), .CO(
        u5_mult_87_CARRYB_47__17_), .S(u5_mult_87_SUMB_47__17_) );
  FA_X1 u5_mult_87_S2_47_16 ( .A(u5_mult_87_ab_47__16_), .B(
        u5_mult_87_CARRYB_46__16_), .CI(u5_mult_87_SUMB_46__17_), .CO(
        u5_mult_87_CARRYB_47__16_), .S(u5_mult_87_SUMB_47__16_) );
  FA_X1 u5_mult_87_S2_47_15 ( .A(u5_mult_87_ab_47__15_), .B(
        u5_mult_87_CARRYB_46__15_), .CI(u5_mult_87_SUMB_46__16_), .CO(
        u5_mult_87_CARRYB_47__15_), .S(u5_mult_87_SUMB_47__15_) );
  FA_X1 u5_mult_87_S2_47_14 ( .A(u5_mult_87_ab_47__14_), .B(
        u5_mult_87_CARRYB_46__14_), .CI(u5_mult_87_SUMB_46__15_), .CO(
        u5_mult_87_CARRYB_47__14_), .S(u5_mult_87_SUMB_47__14_) );
  FA_X1 u5_mult_87_S2_47_13 ( .A(u5_mult_87_ab_47__13_), .B(
        u5_mult_87_CARRYB_46__13_), .CI(u5_mult_87_SUMB_46__14_), .CO(
        u5_mult_87_CARRYB_47__13_), .S(u5_mult_87_SUMB_47__13_) );
  FA_X1 u5_mult_87_S2_47_12 ( .A(u5_mult_87_ab_47__12_), .B(
        u5_mult_87_CARRYB_46__12_), .CI(u5_mult_87_SUMB_46__13_), .CO(
        u5_mult_87_CARRYB_47__12_), .S(u5_mult_87_SUMB_47__12_) );
  FA_X1 u5_mult_87_S2_47_11 ( .A(u5_mult_87_ab_47__11_), .B(
        u5_mult_87_CARRYB_46__11_), .CI(u5_mult_87_SUMB_46__12_), .CO(
        u5_mult_87_CARRYB_47__11_), .S(u5_mult_87_SUMB_47__11_) );
  FA_X1 u5_mult_87_S2_47_10 ( .A(u5_mult_87_ab_47__10_), .B(
        u5_mult_87_CARRYB_46__10_), .CI(u5_mult_87_SUMB_46__11_), .CO(
        u5_mult_87_CARRYB_47__10_), .S(u5_mult_87_SUMB_47__10_) );
  FA_X1 u5_mult_87_S2_47_9 ( .A(u5_mult_87_ab_47__9_), .B(
        u5_mult_87_CARRYB_46__9_), .CI(u5_mult_87_SUMB_46__10_), .CO(
        u5_mult_87_CARRYB_47__9_), .S(u5_mult_87_SUMB_47__9_) );
  FA_X1 u5_mult_87_S2_47_8 ( .A(u5_mult_87_ab_47__8_), .B(
        u5_mult_87_CARRYB_46__8_), .CI(u5_mult_87_SUMB_46__9_), .CO(
        u5_mult_87_CARRYB_47__8_), .S(u5_mult_87_SUMB_47__8_) );
  FA_X1 u5_mult_87_S2_47_7 ( .A(u5_mult_87_ab_47__7_), .B(
        u5_mult_87_CARRYB_46__7_), .CI(u5_mult_87_SUMB_46__8_), .CO(
        u5_mult_87_CARRYB_47__7_), .S(u5_mult_87_SUMB_47__7_) );
  FA_X1 u5_mult_87_S2_47_6 ( .A(u5_mult_87_ab_47__6_), .B(
        u5_mult_87_CARRYB_46__6_), .CI(u5_mult_87_SUMB_46__7_), .CO(
        u5_mult_87_CARRYB_47__6_), .S(u5_mult_87_SUMB_47__6_) );
  FA_X1 u5_mult_87_S2_47_5 ( .A(u5_mult_87_ab_47__5_), .B(
        u5_mult_87_CARRYB_46__5_), .CI(u5_mult_87_SUMB_46__6_), .CO(
        u5_mult_87_CARRYB_47__5_), .S(u5_mult_87_SUMB_47__5_) );
  FA_X1 u5_mult_87_S2_47_4 ( .A(u5_mult_87_ab_47__4_), .B(
        u5_mult_87_CARRYB_46__4_), .CI(u5_mult_87_SUMB_46__5_), .CO(
        u5_mult_87_CARRYB_47__4_), .S(u5_mult_87_SUMB_47__4_) );
  FA_X1 u5_mult_87_S2_47_3 ( .A(u5_mult_87_ab_47__3_), .B(
        u5_mult_87_CARRYB_46__3_), .CI(u5_mult_87_SUMB_46__4_), .CO(
        u5_mult_87_CARRYB_47__3_), .S(u5_mult_87_SUMB_47__3_) );
  FA_X1 u5_mult_87_S2_47_2 ( .A(u5_mult_87_ab_47__2_), .B(
        u5_mult_87_CARRYB_46__2_), .CI(u5_mult_87_SUMB_46__3_), .CO(
        u5_mult_87_CARRYB_47__2_), .S(u5_mult_87_SUMB_47__2_) );
  FA_X1 u5_mult_87_S2_47_1 ( .A(u5_mult_87_ab_47__1_), .B(
        u5_mult_87_CARRYB_46__1_), .CI(u5_mult_87_SUMB_46__2_), .CO(
        u5_mult_87_CARRYB_47__1_), .S(u5_mult_87_SUMB_47__1_) );
  FA_X1 u5_mult_87_S1_47_0 ( .A(u5_mult_87_ab_47__0_), .B(
        u5_mult_87_CARRYB_46__0_), .CI(u5_mult_87_SUMB_46__1_), .CO(
        u5_mult_87_CARRYB_47__0_), .S(u5_N47) );
  FA_X1 u5_mult_87_S3_48_51 ( .A(u5_mult_87_ab_48__51_), .B(
        u5_mult_87_CARRYB_47__51_), .CI(u5_mult_87_ab_47__52_), .CO(
        u5_mult_87_CARRYB_48__51_), .S(u5_mult_87_SUMB_48__51_) );
  FA_X1 u5_mult_87_S2_48_50 ( .A(u5_mult_87_ab_48__50_), .B(
        u5_mult_87_CARRYB_47__50_), .CI(u5_mult_87_SUMB_47__51_), .CO(
        u5_mult_87_CARRYB_48__50_), .S(u5_mult_87_SUMB_48__50_) );
  FA_X1 u5_mult_87_S2_48_49 ( .A(u5_mult_87_ab_48__49_), .B(
        u5_mult_87_CARRYB_47__49_), .CI(u5_mult_87_SUMB_47__50_), .CO(
        u5_mult_87_CARRYB_48__49_), .S(u5_mult_87_SUMB_48__49_) );
  FA_X1 u5_mult_87_S2_48_48 ( .A(u5_mult_87_ab_48__48_), .B(
        u5_mult_87_CARRYB_47__48_), .CI(u5_mult_87_SUMB_47__49_), .CO(
        u5_mult_87_CARRYB_48__48_), .S(u5_mult_87_SUMB_48__48_) );
  FA_X1 u5_mult_87_S2_48_47 ( .A(u5_mult_87_ab_48__47_), .B(
        u5_mult_87_CARRYB_47__47_), .CI(u5_mult_87_SUMB_47__48_), .CO(
        u5_mult_87_CARRYB_48__47_), .S(u5_mult_87_SUMB_48__47_) );
  FA_X1 u5_mult_87_S2_48_46 ( .A(u5_mult_87_ab_48__46_), .B(
        u5_mult_87_CARRYB_47__46_), .CI(u5_mult_87_SUMB_47__47_), .CO(
        u5_mult_87_CARRYB_48__46_), .S(u5_mult_87_SUMB_48__46_) );
  FA_X1 u5_mult_87_S2_48_45 ( .A(u5_mult_87_ab_48__45_), .B(
        u5_mult_87_CARRYB_47__45_), .CI(u5_mult_87_SUMB_47__46_), .CO(
        u5_mult_87_CARRYB_48__45_), .S(u5_mult_87_SUMB_48__45_) );
  FA_X1 u5_mult_87_S2_48_44 ( .A(u5_mult_87_ab_48__44_), .B(
        u5_mult_87_CARRYB_47__44_), .CI(u5_mult_87_SUMB_47__45_), .CO(
        u5_mult_87_CARRYB_48__44_), .S(u5_mult_87_SUMB_48__44_) );
  FA_X1 u5_mult_87_S2_48_43 ( .A(u5_mult_87_ab_48__43_), .B(
        u5_mult_87_CARRYB_47__43_), .CI(u5_mult_87_SUMB_47__44_), .CO(
        u5_mult_87_CARRYB_48__43_), .S(u5_mult_87_SUMB_48__43_) );
  FA_X1 u5_mult_87_S2_48_42 ( .A(u5_mult_87_ab_48__42_), .B(
        u5_mult_87_CARRYB_47__42_), .CI(u5_mult_87_SUMB_47__43_), .CO(
        u5_mult_87_CARRYB_48__42_), .S(u5_mult_87_SUMB_48__42_) );
  FA_X1 u5_mult_87_S2_48_41 ( .A(u5_mult_87_ab_48__41_), .B(
        u5_mult_87_CARRYB_47__41_), .CI(u5_mult_87_SUMB_47__42_), .CO(
        u5_mult_87_CARRYB_48__41_), .S(u5_mult_87_SUMB_48__41_) );
  FA_X1 u5_mult_87_S2_48_40 ( .A(u5_mult_87_ab_48__40_), .B(
        u5_mult_87_CARRYB_47__40_), .CI(u5_mult_87_SUMB_47__41_), .CO(
        u5_mult_87_CARRYB_48__40_), .S(u5_mult_87_SUMB_48__40_) );
  FA_X1 u5_mult_87_S2_48_39 ( .A(u5_mult_87_ab_48__39_), .B(
        u5_mult_87_CARRYB_47__39_), .CI(u5_mult_87_SUMB_47__40_), .CO(
        u5_mult_87_CARRYB_48__39_), .S(u5_mult_87_SUMB_48__39_) );
  FA_X1 u5_mult_87_S2_48_38 ( .A(u5_mult_87_ab_48__38_), .B(
        u5_mult_87_CARRYB_47__38_), .CI(u5_mult_87_SUMB_47__39_), .CO(
        u5_mult_87_CARRYB_48__38_), .S(u5_mult_87_SUMB_48__38_) );
  FA_X1 u5_mult_87_S2_48_37 ( .A(u5_mult_87_ab_48__37_), .B(
        u5_mult_87_CARRYB_47__37_), .CI(u5_mult_87_SUMB_47__38_), .CO(
        u5_mult_87_CARRYB_48__37_), .S(u5_mult_87_SUMB_48__37_) );
  FA_X1 u5_mult_87_S2_48_36 ( .A(u5_mult_87_ab_48__36_), .B(
        u5_mult_87_CARRYB_47__36_), .CI(u5_mult_87_SUMB_47__37_), .CO(
        u5_mult_87_CARRYB_48__36_), .S(u5_mult_87_SUMB_48__36_) );
  FA_X1 u5_mult_87_S2_48_35 ( .A(u5_mult_87_ab_48__35_), .B(
        u5_mult_87_CARRYB_47__35_), .CI(u5_mult_87_SUMB_47__36_), .CO(
        u5_mult_87_CARRYB_48__35_), .S(u5_mult_87_SUMB_48__35_) );
  FA_X1 u5_mult_87_S2_48_34 ( .A(u5_mult_87_ab_48__34_), .B(
        u5_mult_87_CARRYB_47__34_), .CI(u5_mult_87_SUMB_47__35_), .CO(
        u5_mult_87_CARRYB_48__34_), .S(u5_mult_87_SUMB_48__34_) );
  FA_X1 u5_mult_87_S2_48_33 ( .A(u5_mult_87_ab_48__33_), .B(
        u5_mult_87_CARRYB_47__33_), .CI(u5_mult_87_SUMB_47__34_), .CO(
        u5_mult_87_CARRYB_48__33_), .S(u5_mult_87_SUMB_48__33_) );
  FA_X1 u5_mult_87_S2_48_32 ( .A(u5_mult_87_ab_48__32_), .B(
        u5_mult_87_CARRYB_47__32_), .CI(u5_mult_87_SUMB_47__33_), .CO(
        u5_mult_87_CARRYB_48__32_), .S(u5_mult_87_SUMB_48__32_) );
  FA_X1 u5_mult_87_S2_48_31 ( .A(u5_mult_87_ab_48__31_), .B(
        u5_mult_87_CARRYB_47__31_), .CI(u5_mult_87_SUMB_47__32_), .CO(
        u5_mult_87_CARRYB_48__31_), .S(u5_mult_87_SUMB_48__31_) );
  FA_X1 u5_mult_87_S2_48_30 ( .A(u5_mult_87_ab_48__30_), .B(
        u5_mult_87_CARRYB_47__30_), .CI(u5_mult_87_SUMB_47__31_), .CO(
        u5_mult_87_CARRYB_48__30_), .S(u5_mult_87_SUMB_48__30_) );
  FA_X1 u5_mult_87_S2_48_29 ( .A(u5_mult_87_ab_48__29_), .B(
        u5_mult_87_CARRYB_47__29_), .CI(u5_mult_87_SUMB_47__30_), .CO(
        u5_mult_87_CARRYB_48__29_), .S(u5_mult_87_SUMB_48__29_) );
  FA_X1 u5_mult_87_S2_48_28 ( .A(u5_mult_87_ab_48__28_), .B(
        u5_mult_87_CARRYB_47__28_), .CI(u5_mult_87_SUMB_47__29_), .CO(
        u5_mult_87_CARRYB_48__28_), .S(u5_mult_87_SUMB_48__28_) );
  FA_X1 u5_mult_87_S2_48_27 ( .A(u5_mult_87_ab_48__27_), .B(
        u5_mult_87_CARRYB_47__27_), .CI(u5_mult_87_SUMB_47__28_), .CO(
        u5_mult_87_CARRYB_48__27_), .S(u5_mult_87_SUMB_48__27_) );
  FA_X1 u5_mult_87_S2_48_26 ( .A(u5_mult_87_ab_48__26_), .B(
        u5_mult_87_CARRYB_47__26_), .CI(u5_mult_87_SUMB_47__27_), .CO(
        u5_mult_87_CARRYB_48__26_), .S(u5_mult_87_SUMB_48__26_) );
  FA_X1 u5_mult_87_S2_48_25 ( .A(u5_mult_87_ab_48__25_), .B(
        u5_mult_87_CARRYB_47__25_), .CI(u5_mult_87_SUMB_47__26_), .CO(
        u5_mult_87_CARRYB_48__25_), .S(u5_mult_87_SUMB_48__25_) );
  FA_X1 u5_mult_87_S2_48_24 ( .A(u5_mult_87_ab_48__24_), .B(
        u5_mult_87_CARRYB_47__24_), .CI(u5_mult_87_SUMB_47__25_), .CO(
        u5_mult_87_CARRYB_48__24_), .S(u5_mult_87_SUMB_48__24_) );
  FA_X1 u5_mult_87_S2_48_23 ( .A(u5_mult_87_ab_48__23_), .B(
        u5_mult_87_CARRYB_47__23_), .CI(u5_mult_87_SUMB_47__24_), .CO(
        u5_mult_87_CARRYB_48__23_), .S(u5_mult_87_SUMB_48__23_) );
  FA_X1 u5_mult_87_S2_48_22 ( .A(u5_mult_87_ab_48__22_), .B(
        u5_mult_87_CARRYB_47__22_), .CI(u5_mult_87_SUMB_47__23_), .CO(
        u5_mult_87_CARRYB_48__22_), .S(u5_mult_87_SUMB_48__22_) );
  FA_X1 u5_mult_87_S2_48_21 ( .A(u5_mult_87_ab_48__21_), .B(
        u5_mult_87_CARRYB_47__21_), .CI(u5_mult_87_SUMB_47__22_), .CO(
        u5_mult_87_CARRYB_48__21_), .S(u5_mult_87_SUMB_48__21_) );
  FA_X1 u5_mult_87_S2_48_20 ( .A(u5_mult_87_ab_48__20_), .B(
        u5_mult_87_CARRYB_47__20_), .CI(u5_mult_87_SUMB_47__21_), .CO(
        u5_mult_87_CARRYB_48__20_), .S(u5_mult_87_SUMB_48__20_) );
  FA_X1 u5_mult_87_S2_48_19 ( .A(u5_mult_87_ab_48__19_), .B(
        u5_mult_87_CARRYB_47__19_), .CI(u5_mult_87_SUMB_47__20_), .CO(
        u5_mult_87_CARRYB_48__19_), .S(u5_mult_87_SUMB_48__19_) );
  FA_X1 u5_mult_87_S2_48_18 ( .A(u5_mult_87_ab_48__18_), .B(
        u5_mult_87_CARRYB_47__18_), .CI(u5_mult_87_SUMB_47__19_), .CO(
        u5_mult_87_CARRYB_48__18_), .S(u5_mult_87_SUMB_48__18_) );
  FA_X1 u5_mult_87_S2_48_17 ( .A(u5_mult_87_ab_48__17_), .B(
        u5_mult_87_CARRYB_47__17_), .CI(u5_mult_87_SUMB_47__18_), .CO(
        u5_mult_87_CARRYB_48__17_), .S(u5_mult_87_SUMB_48__17_) );
  FA_X1 u5_mult_87_S2_48_16 ( .A(u5_mult_87_ab_48__16_), .B(
        u5_mult_87_CARRYB_47__16_), .CI(u5_mult_87_SUMB_47__17_), .CO(
        u5_mult_87_CARRYB_48__16_), .S(u5_mult_87_SUMB_48__16_) );
  FA_X1 u5_mult_87_S2_48_15 ( .A(u5_mult_87_ab_48__15_), .B(
        u5_mult_87_CARRYB_47__15_), .CI(u5_mult_87_SUMB_47__16_), .CO(
        u5_mult_87_CARRYB_48__15_), .S(u5_mult_87_SUMB_48__15_) );
  FA_X1 u5_mult_87_S2_48_14 ( .A(u5_mult_87_ab_48__14_), .B(
        u5_mult_87_CARRYB_47__14_), .CI(u5_mult_87_SUMB_47__15_), .CO(
        u5_mult_87_CARRYB_48__14_), .S(u5_mult_87_SUMB_48__14_) );
  FA_X1 u5_mult_87_S2_48_13 ( .A(u5_mult_87_ab_48__13_), .B(
        u5_mult_87_CARRYB_47__13_), .CI(u5_mult_87_SUMB_47__14_), .CO(
        u5_mult_87_CARRYB_48__13_), .S(u5_mult_87_SUMB_48__13_) );
  FA_X1 u5_mult_87_S2_48_12 ( .A(u5_mult_87_ab_48__12_), .B(
        u5_mult_87_CARRYB_47__12_), .CI(u5_mult_87_SUMB_47__13_), .CO(
        u5_mult_87_CARRYB_48__12_), .S(u5_mult_87_SUMB_48__12_) );
  FA_X1 u5_mult_87_S2_48_11 ( .A(u5_mult_87_ab_48__11_), .B(
        u5_mult_87_CARRYB_47__11_), .CI(u5_mult_87_SUMB_47__12_), .CO(
        u5_mult_87_CARRYB_48__11_), .S(u5_mult_87_SUMB_48__11_) );
  FA_X1 u5_mult_87_S2_48_10 ( .A(u5_mult_87_ab_48__10_), .B(
        u5_mult_87_CARRYB_47__10_), .CI(u5_mult_87_SUMB_47__11_), .CO(
        u5_mult_87_CARRYB_48__10_), .S(u5_mult_87_SUMB_48__10_) );
  FA_X1 u5_mult_87_S2_48_9 ( .A(u5_mult_87_ab_48__9_), .B(
        u5_mult_87_CARRYB_47__9_), .CI(u5_mult_87_SUMB_47__10_), .CO(
        u5_mult_87_CARRYB_48__9_), .S(u5_mult_87_SUMB_48__9_) );
  FA_X1 u5_mult_87_S2_48_8 ( .A(u5_mult_87_ab_48__8_), .B(
        u5_mult_87_CARRYB_47__8_), .CI(u5_mult_87_SUMB_47__9_), .CO(
        u5_mult_87_CARRYB_48__8_), .S(u5_mult_87_SUMB_48__8_) );
  FA_X1 u5_mult_87_S2_48_7 ( .A(u5_mult_87_ab_48__7_), .B(
        u5_mult_87_CARRYB_47__7_), .CI(u5_mult_87_SUMB_47__8_), .CO(
        u5_mult_87_CARRYB_48__7_), .S(u5_mult_87_SUMB_48__7_) );
  FA_X1 u5_mult_87_S2_48_6 ( .A(u5_mult_87_ab_48__6_), .B(
        u5_mult_87_CARRYB_47__6_), .CI(u5_mult_87_SUMB_47__7_), .CO(
        u5_mult_87_CARRYB_48__6_), .S(u5_mult_87_SUMB_48__6_) );
  FA_X1 u5_mult_87_S2_48_5 ( .A(u5_mult_87_ab_48__5_), .B(
        u5_mult_87_CARRYB_47__5_), .CI(u5_mult_87_SUMB_47__6_), .CO(
        u5_mult_87_CARRYB_48__5_), .S(u5_mult_87_SUMB_48__5_) );
  FA_X1 u5_mult_87_S2_48_4 ( .A(u5_mult_87_ab_48__4_), .B(
        u5_mult_87_CARRYB_47__4_), .CI(u5_mult_87_SUMB_47__5_), .CO(
        u5_mult_87_CARRYB_48__4_), .S(u5_mult_87_SUMB_48__4_) );
  FA_X1 u5_mult_87_S2_48_3 ( .A(u5_mult_87_ab_48__3_), .B(
        u5_mult_87_CARRYB_47__3_), .CI(u5_mult_87_SUMB_47__4_), .CO(
        u5_mult_87_CARRYB_48__3_), .S(u5_mult_87_SUMB_48__3_) );
  FA_X1 u5_mult_87_S2_48_2 ( .A(u5_mult_87_ab_48__2_), .B(
        u5_mult_87_CARRYB_47__2_), .CI(u5_mult_87_SUMB_47__3_), .CO(
        u5_mult_87_CARRYB_48__2_), .S(u5_mult_87_SUMB_48__2_) );
  FA_X1 u5_mult_87_S2_48_1 ( .A(u5_mult_87_ab_48__1_), .B(
        u5_mult_87_CARRYB_47__1_), .CI(u5_mult_87_SUMB_47__2_), .CO(
        u5_mult_87_CARRYB_48__1_), .S(u5_mult_87_SUMB_48__1_) );
  FA_X1 u5_mult_87_S1_48_0 ( .A(u5_mult_87_ab_48__0_), .B(
        u5_mult_87_CARRYB_47__0_), .CI(u5_mult_87_SUMB_47__1_), .CO(
        u5_mult_87_CARRYB_48__0_), .S(u5_N48) );
  FA_X1 u5_mult_87_S3_49_51 ( .A(u5_mult_87_ab_49__51_), .B(
        u5_mult_87_CARRYB_48__51_), .CI(u5_mult_87_ab_48__52_), .CO(
        u5_mult_87_CARRYB_49__51_), .S(u5_mult_87_SUMB_49__51_) );
  FA_X1 u5_mult_87_S2_49_50 ( .A(u5_mult_87_ab_49__50_), .B(
        u5_mult_87_CARRYB_48__50_), .CI(u5_mult_87_SUMB_48__51_), .CO(
        u5_mult_87_CARRYB_49__50_), .S(u5_mult_87_SUMB_49__50_) );
  FA_X1 u5_mult_87_S2_49_49 ( .A(u5_mult_87_ab_49__49_), .B(
        u5_mult_87_CARRYB_48__49_), .CI(u5_mult_87_SUMB_48__50_), .CO(
        u5_mult_87_CARRYB_49__49_), .S(u5_mult_87_SUMB_49__49_) );
  FA_X1 u5_mult_87_S2_49_48 ( .A(u5_mult_87_ab_49__48_), .B(
        u5_mult_87_CARRYB_48__48_), .CI(u5_mult_87_SUMB_48__49_), .CO(
        u5_mult_87_CARRYB_49__48_), .S(u5_mult_87_SUMB_49__48_) );
  FA_X1 u5_mult_87_S2_49_47 ( .A(u5_mult_87_ab_49__47_), .B(
        u5_mult_87_CARRYB_48__47_), .CI(u5_mult_87_SUMB_48__48_), .CO(
        u5_mult_87_CARRYB_49__47_), .S(u5_mult_87_SUMB_49__47_) );
  FA_X1 u5_mult_87_S2_49_46 ( .A(u5_mult_87_ab_49__46_), .B(
        u5_mult_87_CARRYB_48__46_), .CI(u5_mult_87_SUMB_48__47_), .CO(
        u5_mult_87_CARRYB_49__46_), .S(u5_mult_87_SUMB_49__46_) );
  FA_X1 u5_mult_87_S2_49_45 ( .A(u5_mult_87_ab_49__45_), .B(
        u5_mult_87_CARRYB_48__45_), .CI(u5_mult_87_SUMB_48__46_), .CO(
        u5_mult_87_CARRYB_49__45_), .S(u5_mult_87_SUMB_49__45_) );
  FA_X1 u5_mult_87_S2_49_44 ( .A(u5_mult_87_ab_49__44_), .B(
        u5_mult_87_CARRYB_48__44_), .CI(u5_mult_87_SUMB_48__45_), .CO(
        u5_mult_87_CARRYB_49__44_), .S(u5_mult_87_SUMB_49__44_) );
  FA_X1 u5_mult_87_S2_49_43 ( .A(u5_mult_87_ab_49__43_), .B(
        u5_mult_87_CARRYB_48__43_), .CI(u5_mult_87_SUMB_48__44_), .CO(
        u5_mult_87_CARRYB_49__43_), .S(u5_mult_87_SUMB_49__43_) );
  FA_X1 u5_mult_87_S2_49_42 ( .A(u5_mult_87_ab_49__42_), .B(
        u5_mult_87_CARRYB_48__42_), .CI(u5_mult_87_SUMB_48__43_), .CO(
        u5_mult_87_CARRYB_49__42_), .S(u5_mult_87_SUMB_49__42_) );
  FA_X1 u5_mult_87_S2_49_41 ( .A(u5_mult_87_ab_49__41_), .B(
        u5_mult_87_CARRYB_48__41_), .CI(u5_mult_87_SUMB_48__42_), .CO(
        u5_mult_87_CARRYB_49__41_), .S(u5_mult_87_SUMB_49__41_) );
  FA_X1 u5_mult_87_S2_49_40 ( .A(u5_mult_87_ab_49__40_), .B(
        u5_mult_87_CARRYB_48__40_), .CI(u5_mult_87_SUMB_48__41_), .CO(
        u5_mult_87_CARRYB_49__40_), .S(u5_mult_87_SUMB_49__40_) );
  FA_X1 u5_mult_87_S2_49_39 ( .A(u5_mult_87_ab_49__39_), .B(
        u5_mult_87_CARRYB_48__39_), .CI(u5_mult_87_SUMB_48__40_), .CO(
        u5_mult_87_CARRYB_49__39_), .S(u5_mult_87_SUMB_49__39_) );
  FA_X1 u5_mult_87_S2_49_38 ( .A(u5_mult_87_ab_49__38_), .B(
        u5_mult_87_CARRYB_48__38_), .CI(u5_mult_87_SUMB_48__39_), .CO(
        u5_mult_87_CARRYB_49__38_), .S(u5_mult_87_SUMB_49__38_) );
  FA_X1 u5_mult_87_S2_49_37 ( .A(u5_mult_87_ab_49__37_), .B(
        u5_mult_87_CARRYB_48__37_), .CI(u5_mult_87_SUMB_48__38_), .CO(
        u5_mult_87_CARRYB_49__37_), .S(u5_mult_87_SUMB_49__37_) );
  FA_X1 u5_mult_87_S2_49_36 ( .A(u5_mult_87_ab_49__36_), .B(
        u5_mult_87_CARRYB_48__36_), .CI(u5_mult_87_SUMB_48__37_), .CO(
        u5_mult_87_CARRYB_49__36_), .S(u5_mult_87_SUMB_49__36_) );
  FA_X1 u5_mult_87_S2_49_35 ( .A(u5_mult_87_ab_49__35_), .B(
        u5_mult_87_CARRYB_48__35_), .CI(u5_mult_87_SUMB_48__36_), .CO(
        u5_mult_87_CARRYB_49__35_), .S(u5_mult_87_SUMB_49__35_) );
  FA_X1 u5_mult_87_S2_49_34 ( .A(u5_mult_87_ab_49__34_), .B(
        u5_mult_87_CARRYB_48__34_), .CI(u5_mult_87_SUMB_48__35_), .CO(
        u5_mult_87_CARRYB_49__34_), .S(u5_mult_87_SUMB_49__34_) );
  FA_X1 u5_mult_87_S2_49_33 ( .A(u5_mult_87_ab_49__33_), .B(
        u5_mult_87_CARRYB_48__33_), .CI(u5_mult_87_SUMB_48__34_), .CO(
        u5_mult_87_CARRYB_49__33_), .S(u5_mult_87_SUMB_49__33_) );
  FA_X1 u5_mult_87_S2_49_32 ( .A(u5_mult_87_ab_49__32_), .B(
        u5_mult_87_CARRYB_48__32_), .CI(u5_mult_87_SUMB_48__33_), .CO(
        u5_mult_87_CARRYB_49__32_), .S(u5_mult_87_SUMB_49__32_) );
  FA_X1 u5_mult_87_S2_49_31 ( .A(u5_mult_87_ab_49__31_), .B(
        u5_mult_87_CARRYB_48__31_), .CI(u5_mult_87_SUMB_48__32_), .CO(
        u5_mult_87_CARRYB_49__31_), .S(u5_mult_87_SUMB_49__31_) );
  FA_X1 u5_mult_87_S2_49_30 ( .A(u5_mult_87_ab_49__30_), .B(
        u5_mult_87_CARRYB_48__30_), .CI(u5_mult_87_SUMB_48__31_), .CO(
        u5_mult_87_CARRYB_49__30_), .S(u5_mult_87_SUMB_49__30_) );
  FA_X1 u5_mult_87_S2_49_29 ( .A(u5_mult_87_ab_49__29_), .B(
        u5_mult_87_CARRYB_48__29_), .CI(u5_mult_87_SUMB_48__30_), .CO(
        u5_mult_87_CARRYB_49__29_), .S(u5_mult_87_SUMB_49__29_) );
  FA_X1 u5_mult_87_S2_49_28 ( .A(u5_mult_87_ab_49__28_), .B(
        u5_mult_87_CARRYB_48__28_), .CI(u5_mult_87_SUMB_48__29_), .CO(
        u5_mult_87_CARRYB_49__28_), .S(u5_mult_87_SUMB_49__28_) );
  FA_X1 u5_mult_87_S2_49_27 ( .A(u5_mult_87_ab_49__27_), .B(
        u5_mult_87_CARRYB_48__27_), .CI(u5_mult_87_SUMB_48__28_), .CO(
        u5_mult_87_CARRYB_49__27_), .S(u5_mult_87_SUMB_49__27_) );
  FA_X1 u5_mult_87_S2_49_26 ( .A(u5_mult_87_ab_49__26_), .B(
        u5_mult_87_CARRYB_48__26_), .CI(u5_mult_87_SUMB_48__27_), .CO(
        u5_mult_87_CARRYB_49__26_), .S(u5_mult_87_SUMB_49__26_) );
  FA_X1 u5_mult_87_S2_49_25 ( .A(u5_mult_87_ab_49__25_), .B(
        u5_mult_87_CARRYB_48__25_), .CI(u5_mult_87_SUMB_48__26_), .CO(
        u5_mult_87_CARRYB_49__25_), .S(u5_mult_87_SUMB_49__25_) );
  FA_X1 u5_mult_87_S2_49_24 ( .A(u5_mult_87_ab_49__24_), .B(
        u5_mult_87_CARRYB_48__24_), .CI(u5_mult_87_SUMB_48__25_), .CO(
        u5_mult_87_CARRYB_49__24_), .S(u5_mult_87_SUMB_49__24_) );
  FA_X1 u5_mult_87_S2_49_23 ( .A(u5_mult_87_ab_49__23_), .B(
        u5_mult_87_CARRYB_48__23_), .CI(u5_mult_87_SUMB_48__24_), .CO(
        u5_mult_87_CARRYB_49__23_), .S(u5_mult_87_SUMB_49__23_) );
  FA_X1 u5_mult_87_S2_49_22 ( .A(u5_mult_87_ab_49__22_), .B(
        u5_mult_87_CARRYB_48__22_), .CI(u5_mult_87_SUMB_48__23_), .CO(
        u5_mult_87_CARRYB_49__22_), .S(u5_mult_87_SUMB_49__22_) );
  FA_X1 u5_mult_87_S2_49_21 ( .A(u5_mult_87_ab_49__21_), .B(
        u5_mult_87_CARRYB_48__21_), .CI(u5_mult_87_SUMB_48__22_), .CO(
        u5_mult_87_CARRYB_49__21_), .S(u5_mult_87_SUMB_49__21_) );
  FA_X1 u5_mult_87_S2_49_20 ( .A(u5_mult_87_ab_49__20_), .B(
        u5_mult_87_CARRYB_48__20_), .CI(u5_mult_87_SUMB_48__21_), .CO(
        u5_mult_87_CARRYB_49__20_), .S(u5_mult_87_SUMB_49__20_) );
  FA_X1 u5_mult_87_S2_49_19 ( .A(u5_mult_87_ab_49__19_), .B(
        u5_mult_87_CARRYB_48__19_), .CI(u5_mult_87_SUMB_48__20_), .CO(
        u5_mult_87_CARRYB_49__19_), .S(u5_mult_87_SUMB_49__19_) );
  FA_X1 u5_mult_87_S2_49_18 ( .A(u5_mult_87_ab_49__18_), .B(
        u5_mult_87_CARRYB_48__18_), .CI(u5_mult_87_SUMB_48__19_), .CO(
        u5_mult_87_CARRYB_49__18_), .S(u5_mult_87_SUMB_49__18_) );
  FA_X1 u5_mult_87_S2_49_17 ( .A(u5_mult_87_ab_49__17_), .B(
        u5_mult_87_CARRYB_48__17_), .CI(u5_mult_87_SUMB_48__18_), .CO(
        u5_mult_87_CARRYB_49__17_), .S(u5_mult_87_SUMB_49__17_) );
  FA_X1 u5_mult_87_S2_49_16 ( .A(u5_mult_87_ab_49__16_), .B(
        u5_mult_87_CARRYB_48__16_), .CI(u5_mult_87_SUMB_48__17_), .CO(
        u5_mult_87_CARRYB_49__16_), .S(u5_mult_87_SUMB_49__16_) );
  FA_X1 u5_mult_87_S2_49_15 ( .A(u5_mult_87_ab_49__15_), .B(
        u5_mult_87_CARRYB_48__15_), .CI(u5_mult_87_SUMB_48__16_), .CO(
        u5_mult_87_CARRYB_49__15_), .S(u5_mult_87_SUMB_49__15_) );
  FA_X1 u5_mult_87_S2_49_14 ( .A(u5_mult_87_ab_49__14_), .B(
        u5_mult_87_CARRYB_48__14_), .CI(u5_mult_87_SUMB_48__15_), .CO(
        u5_mult_87_CARRYB_49__14_), .S(u5_mult_87_SUMB_49__14_) );
  FA_X1 u5_mult_87_S2_49_13 ( .A(u5_mult_87_ab_49__13_), .B(
        u5_mult_87_CARRYB_48__13_), .CI(u5_mult_87_SUMB_48__14_), .CO(
        u5_mult_87_CARRYB_49__13_), .S(u5_mult_87_SUMB_49__13_) );
  FA_X1 u5_mult_87_S2_49_12 ( .A(u5_mult_87_ab_49__12_), .B(
        u5_mult_87_CARRYB_48__12_), .CI(u5_mult_87_SUMB_48__13_), .CO(
        u5_mult_87_CARRYB_49__12_), .S(u5_mult_87_SUMB_49__12_) );
  FA_X1 u5_mult_87_S2_49_11 ( .A(u5_mult_87_ab_49__11_), .B(
        u5_mult_87_CARRYB_48__11_), .CI(u5_mult_87_SUMB_48__12_), .CO(
        u5_mult_87_CARRYB_49__11_), .S(u5_mult_87_SUMB_49__11_) );
  FA_X1 u5_mult_87_S2_49_10 ( .A(u5_mult_87_ab_49__10_), .B(
        u5_mult_87_CARRYB_48__10_), .CI(u5_mult_87_SUMB_48__11_), .CO(
        u5_mult_87_CARRYB_49__10_), .S(u5_mult_87_SUMB_49__10_) );
  FA_X1 u5_mult_87_S2_49_9 ( .A(u5_mult_87_ab_49__9_), .B(
        u5_mult_87_CARRYB_48__9_), .CI(u5_mult_87_SUMB_48__10_), .CO(
        u5_mult_87_CARRYB_49__9_), .S(u5_mult_87_SUMB_49__9_) );
  FA_X1 u5_mult_87_S2_49_8 ( .A(u5_mult_87_ab_49__8_), .B(
        u5_mult_87_CARRYB_48__8_), .CI(u5_mult_87_SUMB_48__9_), .CO(
        u5_mult_87_CARRYB_49__8_), .S(u5_mult_87_SUMB_49__8_) );
  FA_X1 u5_mult_87_S2_49_7 ( .A(u5_mult_87_ab_49__7_), .B(
        u5_mult_87_CARRYB_48__7_), .CI(u5_mult_87_SUMB_48__8_), .CO(
        u5_mult_87_CARRYB_49__7_), .S(u5_mult_87_SUMB_49__7_) );
  FA_X1 u5_mult_87_S2_49_6 ( .A(u5_mult_87_ab_49__6_), .B(
        u5_mult_87_CARRYB_48__6_), .CI(u5_mult_87_SUMB_48__7_), .CO(
        u5_mult_87_CARRYB_49__6_), .S(u5_mult_87_SUMB_49__6_) );
  FA_X1 u5_mult_87_S2_49_5 ( .A(u5_mult_87_ab_49__5_), .B(
        u5_mult_87_CARRYB_48__5_), .CI(u5_mult_87_SUMB_48__6_), .CO(
        u5_mult_87_CARRYB_49__5_), .S(u5_mult_87_SUMB_49__5_) );
  FA_X1 u5_mult_87_S2_49_4 ( .A(u5_mult_87_ab_49__4_), .B(
        u5_mult_87_CARRYB_48__4_), .CI(u5_mult_87_SUMB_48__5_), .CO(
        u5_mult_87_CARRYB_49__4_), .S(u5_mult_87_SUMB_49__4_) );
  FA_X1 u5_mult_87_S2_49_3 ( .A(u5_mult_87_ab_49__3_), .B(
        u5_mult_87_CARRYB_48__3_), .CI(u5_mult_87_SUMB_48__4_), .CO(
        u5_mult_87_CARRYB_49__3_), .S(u5_mult_87_SUMB_49__3_) );
  FA_X1 u5_mult_87_S2_49_2 ( .A(u5_mult_87_ab_49__2_), .B(
        u5_mult_87_CARRYB_48__2_), .CI(u5_mult_87_SUMB_48__3_), .CO(
        u5_mult_87_CARRYB_49__2_), .S(u5_mult_87_SUMB_49__2_) );
  FA_X1 u5_mult_87_S2_49_1 ( .A(u5_mult_87_ab_49__1_), .B(
        u5_mult_87_CARRYB_48__1_), .CI(u5_mult_87_SUMB_48__2_), .CO(
        u5_mult_87_CARRYB_49__1_), .S(u5_mult_87_SUMB_49__1_) );
  FA_X1 u5_mult_87_S1_49_0 ( .A(u5_mult_87_ab_49__0_), .B(
        u5_mult_87_CARRYB_48__0_), .CI(u5_mult_87_SUMB_48__1_), .CO(
        u5_mult_87_CARRYB_49__0_), .S(u5_N49) );
  FA_X1 u5_mult_87_S3_50_51 ( .A(u5_mult_87_ab_50__51_), .B(
        u5_mult_87_CARRYB_49__51_), .CI(u5_mult_87_ab_49__52_), .CO(
        u5_mult_87_CARRYB_50__51_), .S(u5_mult_87_SUMB_50__51_) );
  FA_X1 u5_mult_87_S2_50_50 ( .A(u5_mult_87_ab_50__50_), .B(
        u5_mult_87_CARRYB_49__50_), .CI(u5_mult_87_SUMB_49__51_), .CO(
        u5_mult_87_CARRYB_50__50_), .S(u5_mult_87_SUMB_50__50_) );
  FA_X1 u5_mult_87_S2_50_49 ( .A(u5_mult_87_ab_50__49_), .B(
        u5_mult_87_CARRYB_49__49_), .CI(u5_mult_87_SUMB_49__50_), .CO(
        u5_mult_87_CARRYB_50__49_), .S(u5_mult_87_SUMB_50__49_) );
  FA_X1 u5_mult_87_S2_50_48 ( .A(u5_mult_87_ab_50__48_), .B(
        u5_mult_87_CARRYB_49__48_), .CI(u5_mult_87_SUMB_49__49_), .CO(
        u5_mult_87_CARRYB_50__48_), .S(u5_mult_87_SUMB_50__48_) );
  FA_X1 u5_mult_87_S2_50_47 ( .A(u5_mult_87_ab_50__47_), .B(
        u5_mult_87_CARRYB_49__47_), .CI(u5_mult_87_SUMB_49__48_), .CO(
        u5_mult_87_CARRYB_50__47_), .S(u5_mult_87_SUMB_50__47_) );
  FA_X1 u5_mult_87_S2_50_46 ( .A(u5_mult_87_ab_50__46_), .B(
        u5_mult_87_CARRYB_49__46_), .CI(u5_mult_87_SUMB_49__47_), .CO(
        u5_mult_87_CARRYB_50__46_), .S(u5_mult_87_SUMB_50__46_) );
  FA_X1 u5_mult_87_S2_50_45 ( .A(u5_mult_87_ab_50__45_), .B(
        u5_mult_87_CARRYB_49__45_), .CI(u5_mult_87_SUMB_49__46_), .CO(
        u5_mult_87_CARRYB_50__45_), .S(u5_mult_87_SUMB_50__45_) );
  FA_X1 u5_mult_87_S2_50_44 ( .A(u5_mult_87_ab_50__44_), .B(
        u5_mult_87_CARRYB_49__44_), .CI(u5_mult_87_SUMB_49__45_), .CO(
        u5_mult_87_CARRYB_50__44_), .S(u5_mult_87_SUMB_50__44_) );
  FA_X1 u5_mult_87_S2_50_43 ( .A(u5_mult_87_ab_50__43_), .B(
        u5_mult_87_CARRYB_49__43_), .CI(u5_mult_87_SUMB_49__44_), .CO(
        u5_mult_87_CARRYB_50__43_), .S(u5_mult_87_SUMB_50__43_) );
  FA_X1 u5_mult_87_S2_50_42 ( .A(u5_mult_87_ab_50__42_), .B(
        u5_mult_87_CARRYB_49__42_), .CI(u5_mult_87_SUMB_49__43_), .CO(
        u5_mult_87_CARRYB_50__42_), .S(u5_mult_87_SUMB_50__42_) );
  FA_X1 u5_mult_87_S2_50_41 ( .A(u5_mult_87_ab_50__41_), .B(
        u5_mult_87_CARRYB_49__41_), .CI(u5_mult_87_SUMB_49__42_), .CO(
        u5_mult_87_CARRYB_50__41_), .S(u5_mult_87_SUMB_50__41_) );
  FA_X1 u5_mult_87_S2_50_40 ( .A(u5_mult_87_ab_50__40_), .B(
        u5_mult_87_CARRYB_49__40_), .CI(u5_mult_87_SUMB_49__41_), .CO(
        u5_mult_87_CARRYB_50__40_), .S(u5_mult_87_SUMB_50__40_) );
  FA_X1 u5_mult_87_S2_50_39 ( .A(u5_mult_87_ab_50__39_), .B(
        u5_mult_87_CARRYB_49__39_), .CI(u5_mult_87_SUMB_49__40_), .CO(
        u5_mult_87_CARRYB_50__39_), .S(u5_mult_87_SUMB_50__39_) );
  FA_X1 u5_mult_87_S2_50_38 ( .A(u5_mult_87_ab_50__38_), .B(
        u5_mult_87_CARRYB_49__38_), .CI(u5_mult_87_SUMB_49__39_), .CO(
        u5_mult_87_CARRYB_50__38_), .S(u5_mult_87_SUMB_50__38_) );
  FA_X1 u5_mult_87_S2_50_37 ( .A(u5_mult_87_ab_50__37_), .B(
        u5_mult_87_CARRYB_49__37_), .CI(u5_mult_87_SUMB_49__38_), .CO(
        u5_mult_87_CARRYB_50__37_), .S(u5_mult_87_SUMB_50__37_) );
  FA_X1 u5_mult_87_S2_50_36 ( .A(u5_mult_87_ab_50__36_), .B(
        u5_mult_87_CARRYB_49__36_), .CI(u5_mult_87_SUMB_49__37_), .CO(
        u5_mult_87_CARRYB_50__36_), .S(u5_mult_87_SUMB_50__36_) );
  FA_X1 u5_mult_87_S2_50_35 ( .A(u5_mult_87_ab_50__35_), .B(
        u5_mult_87_CARRYB_49__35_), .CI(u5_mult_87_SUMB_49__36_), .CO(
        u5_mult_87_CARRYB_50__35_), .S(u5_mult_87_SUMB_50__35_) );
  FA_X1 u5_mult_87_S2_50_34 ( .A(u5_mult_87_ab_50__34_), .B(
        u5_mult_87_CARRYB_49__34_), .CI(u5_mult_87_SUMB_49__35_), .CO(
        u5_mult_87_CARRYB_50__34_), .S(u5_mult_87_SUMB_50__34_) );
  FA_X1 u5_mult_87_S2_50_33 ( .A(u5_mult_87_ab_50__33_), .B(
        u5_mult_87_CARRYB_49__33_), .CI(u5_mult_87_SUMB_49__34_), .CO(
        u5_mult_87_CARRYB_50__33_), .S(u5_mult_87_SUMB_50__33_) );
  FA_X1 u5_mult_87_S2_50_32 ( .A(u5_mult_87_ab_50__32_), .B(
        u5_mult_87_CARRYB_49__32_), .CI(u5_mult_87_SUMB_49__33_), .CO(
        u5_mult_87_CARRYB_50__32_), .S(u5_mult_87_SUMB_50__32_) );
  FA_X1 u5_mult_87_S2_50_31 ( .A(u5_mult_87_ab_50__31_), .B(
        u5_mult_87_CARRYB_49__31_), .CI(u5_mult_87_SUMB_49__32_), .CO(
        u5_mult_87_CARRYB_50__31_), .S(u5_mult_87_SUMB_50__31_) );
  FA_X1 u5_mult_87_S2_50_30 ( .A(u5_mult_87_ab_50__30_), .B(
        u5_mult_87_CARRYB_49__30_), .CI(u5_mult_87_SUMB_49__31_), .CO(
        u5_mult_87_CARRYB_50__30_), .S(u5_mult_87_SUMB_50__30_) );
  FA_X1 u5_mult_87_S2_50_29 ( .A(u5_mult_87_ab_50__29_), .B(
        u5_mult_87_CARRYB_49__29_), .CI(u5_mult_87_SUMB_49__30_), .CO(
        u5_mult_87_CARRYB_50__29_), .S(u5_mult_87_SUMB_50__29_) );
  FA_X1 u5_mult_87_S2_50_28 ( .A(u5_mult_87_ab_50__28_), .B(
        u5_mult_87_CARRYB_49__28_), .CI(u5_mult_87_SUMB_49__29_), .CO(
        u5_mult_87_CARRYB_50__28_), .S(u5_mult_87_SUMB_50__28_) );
  FA_X1 u5_mult_87_S2_50_27 ( .A(u5_mult_87_ab_50__27_), .B(
        u5_mult_87_CARRYB_49__27_), .CI(u5_mult_87_SUMB_49__28_), .CO(
        u5_mult_87_CARRYB_50__27_), .S(u5_mult_87_SUMB_50__27_) );
  FA_X1 u5_mult_87_S2_50_26 ( .A(u5_mult_87_ab_50__26_), .B(
        u5_mult_87_CARRYB_49__26_), .CI(u5_mult_87_SUMB_49__27_), .CO(
        u5_mult_87_CARRYB_50__26_), .S(u5_mult_87_SUMB_50__26_) );
  FA_X1 u5_mult_87_S2_50_25 ( .A(u5_mult_87_ab_50__25_), .B(
        u5_mult_87_CARRYB_49__25_), .CI(u5_mult_87_SUMB_49__26_), .CO(
        u5_mult_87_CARRYB_50__25_), .S(u5_mult_87_SUMB_50__25_) );
  FA_X1 u5_mult_87_S2_50_24 ( .A(u5_mult_87_ab_50__24_), .B(
        u5_mult_87_CARRYB_49__24_), .CI(u5_mult_87_SUMB_49__25_), .CO(
        u5_mult_87_CARRYB_50__24_), .S(u5_mult_87_SUMB_50__24_) );
  FA_X1 u5_mult_87_S2_50_23 ( .A(u5_mult_87_ab_50__23_), .B(
        u5_mult_87_CARRYB_49__23_), .CI(u5_mult_87_SUMB_49__24_), .CO(
        u5_mult_87_CARRYB_50__23_), .S(u5_mult_87_SUMB_50__23_) );
  FA_X1 u5_mult_87_S2_50_22 ( .A(u5_mult_87_ab_50__22_), .B(
        u5_mult_87_CARRYB_49__22_), .CI(u5_mult_87_SUMB_49__23_), .CO(
        u5_mult_87_CARRYB_50__22_), .S(u5_mult_87_SUMB_50__22_) );
  FA_X1 u5_mult_87_S2_50_21 ( .A(u5_mult_87_ab_50__21_), .B(
        u5_mult_87_CARRYB_49__21_), .CI(u5_mult_87_SUMB_49__22_), .CO(
        u5_mult_87_CARRYB_50__21_), .S(u5_mult_87_SUMB_50__21_) );
  FA_X1 u5_mult_87_S2_50_20 ( .A(u5_mult_87_ab_50__20_), .B(
        u5_mult_87_CARRYB_49__20_), .CI(u5_mult_87_SUMB_49__21_), .CO(
        u5_mult_87_CARRYB_50__20_), .S(u5_mult_87_SUMB_50__20_) );
  FA_X1 u5_mult_87_S2_50_19 ( .A(u5_mult_87_ab_50__19_), .B(
        u5_mult_87_CARRYB_49__19_), .CI(u5_mult_87_SUMB_49__20_), .CO(
        u5_mult_87_CARRYB_50__19_), .S(u5_mult_87_SUMB_50__19_) );
  FA_X1 u5_mult_87_S2_50_18 ( .A(u5_mult_87_ab_50__18_), .B(
        u5_mult_87_CARRYB_49__18_), .CI(u5_mult_87_SUMB_49__19_), .CO(
        u5_mult_87_CARRYB_50__18_), .S(u5_mult_87_SUMB_50__18_) );
  FA_X1 u5_mult_87_S2_50_17 ( .A(u5_mult_87_ab_50__17_), .B(
        u5_mult_87_CARRYB_49__17_), .CI(u5_mult_87_SUMB_49__18_), .CO(
        u5_mult_87_CARRYB_50__17_), .S(u5_mult_87_SUMB_50__17_) );
  FA_X1 u5_mult_87_S2_50_16 ( .A(u5_mult_87_ab_50__16_), .B(
        u5_mult_87_CARRYB_49__16_), .CI(u5_mult_87_SUMB_49__17_), .CO(
        u5_mult_87_CARRYB_50__16_), .S(u5_mult_87_SUMB_50__16_) );
  FA_X1 u5_mult_87_S2_50_15 ( .A(u5_mult_87_ab_50__15_), .B(
        u5_mult_87_CARRYB_49__15_), .CI(u5_mult_87_SUMB_49__16_), .CO(
        u5_mult_87_CARRYB_50__15_), .S(u5_mult_87_SUMB_50__15_) );
  FA_X1 u5_mult_87_S2_50_14 ( .A(u5_mult_87_ab_50__14_), .B(
        u5_mult_87_CARRYB_49__14_), .CI(u5_mult_87_SUMB_49__15_), .CO(
        u5_mult_87_CARRYB_50__14_), .S(u5_mult_87_SUMB_50__14_) );
  FA_X1 u5_mult_87_S2_50_13 ( .A(u5_mult_87_ab_50__13_), .B(
        u5_mult_87_CARRYB_49__13_), .CI(u5_mult_87_SUMB_49__14_), .CO(
        u5_mult_87_CARRYB_50__13_), .S(u5_mult_87_SUMB_50__13_) );
  FA_X1 u5_mult_87_S2_50_12 ( .A(u5_mult_87_ab_50__12_), .B(
        u5_mult_87_CARRYB_49__12_), .CI(u5_mult_87_SUMB_49__13_), .CO(
        u5_mult_87_CARRYB_50__12_), .S(u5_mult_87_SUMB_50__12_) );
  FA_X1 u5_mult_87_S2_50_11 ( .A(u5_mult_87_ab_50__11_), .B(
        u5_mult_87_CARRYB_49__11_), .CI(u5_mult_87_SUMB_49__12_), .CO(
        u5_mult_87_CARRYB_50__11_), .S(u5_mult_87_SUMB_50__11_) );
  FA_X1 u5_mult_87_S2_50_10 ( .A(u5_mult_87_ab_50__10_), .B(
        u5_mult_87_CARRYB_49__10_), .CI(u5_mult_87_SUMB_49__11_), .CO(
        u5_mult_87_CARRYB_50__10_), .S(u5_mult_87_SUMB_50__10_) );
  FA_X1 u5_mult_87_S2_50_9 ( .A(u5_mult_87_ab_50__9_), .B(
        u5_mult_87_CARRYB_49__9_), .CI(u5_mult_87_SUMB_49__10_), .CO(
        u5_mult_87_CARRYB_50__9_), .S(u5_mult_87_SUMB_50__9_) );
  FA_X1 u5_mult_87_S2_50_8 ( .A(u5_mult_87_ab_50__8_), .B(
        u5_mult_87_CARRYB_49__8_), .CI(u5_mult_87_SUMB_49__9_), .CO(
        u5_mult_87_CARRYB_50__8_), .S(u5_mult_87_SUMB_50__8_) );
  FA_X1 u5_mult_87_S2_50_7 ( .A(u5_mult_87_ab_50__7_), .B(
        u5_mult_87_CARRYB_49__7_), .CI(u5_mult_87_SUMB_49__8_), .CO(
        u5_mult_87_CARRYB_50__7_), .S(u5_mult_87_SUMB_50__7_) );
  FA_X1 u5_mult_87_S2_50_6 ( .A(u5_mult_87_ab_50__6_), .B(
        u5_mult_87_CARRYB_49__6_), .CI(u5_mult_87_SUMB_49__7_), .CO(
        u5_mult_87_CARRYB_50__6_), .S(u5_mult_87_SUMB_50__6_) );
  FA_X1 u5_mult_87_S2_50_5 ( .A(u5_mult_87_ab_50__5_), .B(
        u5_mult_87_CARRYB_49__5_), .CI(u5_mult_87_SUMB_49__6_), .CO(
        u5_mult_87_CARRYB_50__5_), .S(u5_mult_87_SUMB_50__5_) );
  FA_X1 u5_mult_87_S2_50_4 ( .A(u5_mult_87_ab_50__4_), .B(
        u5_mult_87_CARRYB_49__4_), .CI(u5_mult_87_SUMB_49__5_), .CO(
        u5_mult_87_CARRYB_50__4_), .S(u5_mult_87_SUMB_50__4_) );
  FA_X1 u5_mult_87_S2_50_3 ( .A(u5_mult_87_ab_50__3_), .B(
        u5_mult_87_CARRYB_49__3_), .CI(u5_mult_87_SUMB_49__4_), .CO(
        u5_mult_87_CARRYB_50__3_), .S(u5_mult_87_SUMB_50__3_) );
  FA_X1 u5_mult_87_S2_50_2 ( .A(u5_mult_87_ab_50__2_), .B(
        u5_mult_87_CARRYB_49__2_), .CI(u5_mult_87_SUMB_49__3_), .CO(
        u5_mult_87_CARRYB_50__2_), .S(u5_mult_87_SUMB_50__2_) );
  FA_X1 u5_mult_87_S2_50_1 ( .A(u5_mult_87_ab_50__1_), .B(
        u5_mult_87_CARRYB_49__1_), .CI(u5_mult_87_SUMB_49__2_), .CO(
        u5_mult_87_CARRYB_50__1_), .S(u5_mult_87_SUMB_50__1_) );
  FA_X1 u5_mult_87_S1_50_0 ( .A(u5_mult_87_ab_50__0_), .B(
        u5_mult_87_CARRYB_49__0_), .CI(u5_mult_87_SUMB_49__1_), .CO(
        u5_mult_87_CARRYB_50__0_), .S(u5_N50) );
  FA_X1 u5_mult_87_S3_51_51 ( .A(u5_mult_87_ab_51__51_), .B(
        u5_mult_87_CARRYB_50__51_), .CI(u5_mult_87_ab_50__52_), .CO(
        u5_mult_87_CARRYB_51__51_), .S(u5_mult_87_SUMB_51__51_) );
  FA_X1 u5_mult_87_S2_51_50 ( .A(u5_mult_87_ab_51__50_), .B(
        u5_mult_87_CARRYB_50__50_), .CI(u5_mult_87_SUMB_50__51_), .CO(
        u5_mult_87_CARRYB_51__50_), .S(u5_mult_87_SUMB_51__50_) );
  FA_X1 u5_mult_87_S2_51_49 ( .A(u5_mult_87_ab_51__49_), .B(
        u5_mult_87_CARRYB_50__49_), .CI(u5_mult_87_SUMB_50__50_), .CO(
        u5_mult_87_CARRYB_51__49_), .S(u5_mult_87_SUMB_51__49_) );
  FA_X1 u5_mult_87_S2_51_48 ( .A(u5_mult_87_ab_51__48_), .B(
        u5_mult_87_CARRYB_50__48_), .CI(u5_mult_87_SUMB_50__49_), .CO(
        u5_mult_87_CARRYB_51__48_), .S(u5_mult_87_SUMB_51__48_) );
  FA_X1 u5_mult_87_S2_51_47 ( .A(u5_mult_87_ab_51__47_), .B(
        u5_mult_87_CARRYB_50__47_), .CI(u5_mult_87_SUMB_50__48_), .CO(
        u5_mult_87_CARRYB_51__47_), .S(u5_mult_87_SUMB_51__47_) );
  FA_X1 u5_mult_87_S2_51_46 ( .A(u5_mult_87_ab_51__46_), .B(
        u5_mult_87_CARRYB_50__46_), .CI(u5_mult_87_SUMB_50__47_), .CO(
        u5_mult_87_CARRYB_51__46_), .S(u5_mult_87_SUMB_51__46_) );
  FA_X1 u5_mult_87_S2_51_45 ( .A(u5_mult_87_ab_51__45_), .B(
        u5_mult_87_CARRYB_50__45_), .CI(u5_mult_87_SUMB_50__46_), .CO(
        u5_mult_87_CARRYB_51__45_), .S(u5_mult_87_SUMB_51__45_) );
  FA_X1 u5_mult_87_S2_51_44 ( .A(u5_mult_87_ab_51__44_), .B(
        u5_mult_87_CARRYB_50__44_), .CI(u5_mult_87_SUMB_50__45_), .CO(
        u5_mult_87_CARRYB_51__44_), .S(u5_mult_87_SUMB_51__44_) );
  FA_X1 u5_mult_87_S2_51_43 ( .A(u5_mult_87_ab_51__43_), .B(
        u5_mult_87_CARRYB_50__43_), .CI(u5_mult_87_SUMB_50__44_), .CO(
        u5_mult_87_CARRYB_51__43_), .S(u5_mult_87_SUMB_51__43_) );
  FA_X1 u5_mult_87_S2_51_42 ( .A(u5_mult_87_ab_51__42_), .B(
        u5_mult_87_CARRYB_50__42_), .CI(u5_mult_87_SUMB_50__43_), .CO(
        u5_mult_87_CARRYB_51__42_), .S(u5_mult_87_SUMB_51__42_) );
  FA_X1 u5_mult_87_S2_51_41 ( .A(u5_mult_87_ab_51__41_), .B(
        u5_mult_87_CARRYB_50__41_), .CI(u5_mult_87_SUMB_50__42_), .CO(
        u5_mult_87_CARRYB_51__41_), .S(u5_mult_87_SUMB_51__41_) );
  FA_X1 u5_mult_87_S2_51_40 ( .A(u5_mult_87_ab_51__40_), .B(
        u5_mult_87_CARRYB_50__40_), .CI(u5_mult_87_SUMB_50__41_), .CO(
        u5_mult_87_CARRYB_51__40_), .S(u5_mult_87_SUMB_51__40_) );
  FA_X1 u5_mult_87_S2_51_39 ( .A(u5_mult_87_ab_51__39_), .B(
        u5_mult_87_CARRYB_50__39_), .CI(u5_mult_87_SUMB_50__40_), .CO(
        u5_mult_87_CARRYB_51__39_), .S(u5_mult_87_SUMB_51__39_) );
  FA_X1 u5_mult_87_S2_51_38 ( .A(u5_mult_87_ab_51__38_), .B(
        u5_mult_87_CARRYB_50__38_), .CI(u5_mult_87_SUMB_50__39_), .CO(
        u5_mult_87_CARRYB_51__38_), .S(u5_mult_87_SUMB_51__38_) );
  FA_X1 u5_mult_87_S2_51_37 ( .A(u5_mult_87_ab_51__37_), .B(
        u5_mult_87_CARRYB_50__37_), .CI(u5_mult_87_SUMB_50__38_), .CO(
        u5_mult_87_CARRYB_51__37_), .S(u5_mult_87_SUMB_51__37_) );
  FA_X1 u5_mult_87_S2_51_36 ( .A(u5_mult_87_ab_51__36_), .B(
        u5_mult_87_CARRYB_50__36_), .CI(u5_mult_87_SUMB_50__37_), .CO(
        u5_mult_87_CARRYB_51__36_), .S(u5_mult_87_SUMB_51__36_) );
  FA_X1 u5_mult_87_S2_51_35 ( .A(u5_mult_87_ab_51__35_), .B(
        u5_mult_87_CARRYB_50__35_), .CI(u5_mult_87_SUMB_50__36_), .CO(
        u5_mult_87_CARRYB_51__35_), .S(u5_mult_87_SUMB_51__35_) );
  FA_X1 u5_mult_87_S2_51_34 ( .A(u5_mult_87_ab_51__34_), .B(
        u5_mult_87_CARRYB_50__34_), .CI(u5_mult_87_SUMB_50__35_), .CO(
        u5_mult_87_CARRYB_51__34_), .S(u5_mult_87_SUMB_51__34_) );
  FA_X1 u5_mult_87_S2_51_33 ( .A(u5_mult_87_ab_51__33_), .B(
        u5_mult_87_CARRYB_50__33_), .CI(u5_mult_87_SUMB_50__34_), .CO(
        u5_mult_87_CARRYB_51__33_), .S(u5_mult_87_SUMB_51__33_) );
  FA_X1 u5_mult_87_S2_51_32 ( .A(u5_mult_87_ab_51__32_), .B(
        u5_mult_87_CARRYB_50__32_), .CI(u5_mult_87_SUMB_50__33_), .CO(
        u5_mult_87_CARRYB_51__32_), .S(u5_mult_87_SUMB_51__32_) );
  FA_X1 u5_mult_87_S2_51_31 ( .A(u5_mult_87_ab_51__31_), .B(
        u5_mult_87_CARRYB_50__31_), .CI(u5_mult_87_SUMB_50__32_), .CO(
        u5_mult_87_CARRYB_51__31_), .S(u5_mult_87_SUMB_51__31_) );
  FA_X1 u5_mult_87_S2_51_30 ( .A(u5_mult_87_ab_51__30_), .B(
        u5_mult_87_CARRYB_50__30_), .CI(u5_mult_87_SUMB_50__31_), .CO(
        u5_mult_87_CARRYB_51__30_), .S(u5_mult_87_SUMB_51__30_) );
  FA_X1 u5_mult_87_S2_51_29 ( .A(u5_mult_87_ab_51__29_), .B(
        u5_mult_87_CARRYB_50__29_), .CI(u5_mult_87_SUMB_50__30_), .CO(
        u5_mult_87_CARRYB_51__29_), .S(u5_mult_87_SUMB_51__29_) );
  FA_X1 u5_mult_87_S2_51_28 ( .A(u5_mult_87_ab_51__28_), .B(
        u5_mult_87_CARRYB_50__28_), .CI(u5_mult_87_SUMB_50__29_), .CO(
        u5_mult_87_CARRYB_51__28_), .S(u5_mult_87_SUMB_51__28_) );
  FA_X1 u5_mult_87_S2_51_27 ( .A(u5_mult_87_ab_51__27_), .B(
        u5_mult_87_CARRYB_50__27_), .CI(u5_mult_87_SUMB_50__28_), .CO(
        u5_mult_87_CARRYB_51__27_), .S(u5_mult_87_SUMB_51__27_) );
  FA_X1 u5_mult_87_S2_51_26 ( .A(u5_mult_87_ab_51__26_), .B(
        u5_mult_87_CARRYB_50__26_), .CI(u5_mult_87_SUMB_50__27_), .CO(
        u5_mult_87_CARRYB_51__26_), .S(u5_mult_87_SUMB_51__26_) );
  FA_X1 u5_mult_87_S2_51_25 ( .A(u5_mult_87_ab_51__25_), .B(
        u5_mult_87_CARRYB_50__25_), .CI(u5_mult_87_SUMB_50__26_), .CO(
        u5_mult_87_CARRYB_51__25_), .S(u5_mult_87_SUMB_51__25_) );
  FA_X1 u5_mult_87_S2_51_24 ( .A(u5_mult_87_ab_51__24_), .B(
        u5_mult_87_CARRYB_50__24_), .CI(u5_mult_87_SUMB_50__25_), .CO(
        u5_mult_87_CARRYB_51__24_), .S(u5_mult_87_SUMB_51__24_) );
  FA_X1 u5_mult_87_S2_51_23 ( .A(u5_mult_87_ab_51__23_), .B(
        u5_mult_87_CARRYB_50__23_), .CI(u5_mult_87_SUMB_50__24_), .CO(
        u5_mult_87_CARRYB_51__23_), .S(u5_mult_87_SUMB_51__23_) );
  FA_X1 u5_mult_87_S2_51_22 ( .A(u5_mult_87_ab_51__22_), .B(
        u5_mult_87_CARRYB_50__22_), .CI(u5_mult_87_SUMB_50__23_), .CO(
        u5_mult_87_CARRYB_51__22_), .S(u5_mult_87_SUMB_51__22_) );
  FA_X1 u5_mult_87_S2_51_21 ( .A(u5_mult_87_ab_51__21_), .B(
        u5_mult_87_CARRYB_50__21_), .CI(u5_mult_87_SUMB_50__22_), .CO(
        u5_mult_87_CARRYB_51__21_), .S(u5_mult_87_SUMB_51__21_) );
  FA_X1 u5_mult_87_S2_51_20 ( .A(u5_mult_87_ab_51__20_), .B(
        u5_mult_87_CARRYB_50__20_), .CI(u5_mult_87_SUMB_50__21_), .CO(
        u5_mult_87_CARRYB_51__20_), .S(u5_mult_87_SUMB_51__20_) );
  FA_X1 u5_mult_87_S2_51_19 ( .A(u5_mult_87_ab_51__19_), .B(
        u5_mult_87_CARRYB_50__19_), .CI(u5_mult_87_SUMB_50__20_), .CO(
        u5_mult_87_CARRYB_51__19_), .S(u5_mult_87_SUMB_51__19_) );
  FA_X1 u5_mult_87_S2_51_18 ( .A(u5_mult_87_ab_51__18_), .B(
        u5_mult_87_CARRYB_50__18_), .CI(u5_mult_87_SUMB_50__19_), .CO(
        u5_mult_87_CARRYB_51__18_), .S(u5_mult_87_SUMB_51__18_) );
  FA_X1 u5_mult_87_S2_51_17 ( .A(u5_mult_87_ab_51__17_), .B(
        u5_mult_87_CARRYB_50__17_), .CI(u5_mult_87_SUMB_50__18_), .CO(
        u5_mult_87_CARRYB_51__17_), .S(u5_mult_87_SUMB_51__17_) );
  FA_X1 u5_mult_87_S2_51_16 ( .A(u5_mult_87_ab_51__16_), .B(
        u5_mult_87_CARRYB_50__16_), .CI(u5_mult_87_SUMB_50__17_), .CO(
        u5_mult_87_CARRYB_51__16_), .S(u5_mult_87_SUMB_51__16_) );
  FA_X1 u5_mult_87_S2_51_15 ( .A(u5_mult_87_ab_51__15_), .B(
        u5_mult_87_CARRYB_50__15_), .CI(u5_mult_87_SUMB_50__16_), .CO(
        u5_mult_87_CARRYB_51__15_), .S(u5_mult_87_SUMB_51__15_) );
  FA_X1 u5_mult_87_S2_51_14 ( .A(u5_mult_87_ab_51__14_), .B(
        u5_mult_87_CARRYB_50__14_), .CI(u5_mult_87_SUMB_50__15_), .CO(
        u5_mult_87_CARRYB_51__14_), .S(u5_mult_87_SUMB_51__14_) );
  FA_X1 u5_mult_87_S2_51_13 ( .A(u5_mult_87_ab_51__13_), .B(
        u5_mult_87_CARRYB_50__13_), .CI(u5_mult_87_SUMB_50__14_), .CO(
        u5_mult_87_CARRYB_51__13_), .S(u5_mult_87_SUMB_51__13_) );
  FA_X1 u5_mult_87_S2_51_12 ( .A(u5_mult_87_ab_51__12_), .B(
        u5_mult_87_CARRYB_50__12_), .CI(u5_mult_87_SUMB_50__13_), .CO(
        u5_mult_87_CARRYB_51__12_), .S(u5_mult_87_SUMB_51__12_) );
  FA_X1 u5_mult_87_S2_51_11 ( .A(u5_mult_87_ab_51__11_), .B(
        u5_mult_87_CARRYB_50__11_), .CI(u5_mult_87_SUMB_50__12_), .CO(
        u5_mult_87_CARRYB_51__11_), .S(u5_mult_87_SUMB_51__11_) );
  FA_X1 u5_mult_87_S2_51_10 ( .A(u5_mult_87_ab_51__10_), .B(
        u5_mult_87_CARRYB_50__10_), .CI(u5_mult_87_SUMB_50__11_), .CO(
        u5_mult_87_CARRYB_51__10_), .S(u5_mult_87_SUMB_51__10_) );
  FA_X1 u5_mult_87_S2_51_9 ( .A(u5_mult_87_ab_51__9_), .B(
        u5_mult_87_CARRYB_50__9_), .CI(u5_mult_87_SUMB_50__10_), .CO(
        u5_mult_87_CARRYB_51__9_), .S(u5_mult_87_SUMB_51__9_) );
  FA_X1 u5_mult_87_S2_51_8 ( .A(u5_mult_87_ab_51__8_), .B(
        u5_mult_87_CARRYB_50__8_), .CI(u5_mult_87_SUMB_50__9_), .CO(
        u5_mult_87_CARRYB_51__8_), .S(u5_mult_87_SUMB_51__8_) );
  FA_X1 u5_mult_87_S2_51_7 ( .A(u5_mult_87_ab_51__7_), .B(
        u5_mult_87_CARRYB_50__7_), .CI(u5_mult_87_SUMB_50__8_), .CO(
        u5_mult_87_CARRYB_51__7_), .S(u5_mult_87_SUMB_51__7_) );
  FA_X1 u5_mult_87_S2_51_6 ( .A(u5_mult_87_ab_51__6_), .B(
        u5_mult_87_CARRYB_50__6_), .CI(u5_mult_87_SUMB_50__7_), .CO(
        u5_mult_87_CARRYB_51__6_), .S(u5_mult_87_SUMB_51__6_) );
  FA_X1 u5_mult_87_S2_51_5 ( .A(u5_mult_87_ab_51__5_), .B(
        u5_mult_87_CARRYB_50__5_), .CI(u5_mult_87_SUMB_50__6_), .CO(
        u5_mult_87_CARRYB_51__5_), .S(u5_mult_87_SUMB_51__5_) );
  FA_X1 u5_mult_87_S2_51_4 ( .A(u5_mult_87_ab_51__4_), .B(
        u5_mult_87_CARRYB_50__4_), .CI(u5_mult_87_SUMB_50__5_), .CO(
        u5_mult_87_CARRYB_51__4_), .S(u5_mult_87_SUMB_51__4_) );
  FA_X1 u5_mult_87_S2_51_3 ( .A(u5_mult_87_ab_51__3_), .B(
        u5_mult_87_CARRYB_50__3_), .CI(u5_mult_87_SUMB_50__4_), .CO(
        u5_mult_87_CARRYB_51__3_), .S(u5_mult_87_SUMB_51__3_) );
  FA_X1 u5_mult_87_S2_51_2 ( .A(u5_mult_87_ab_51__2_), .B(
        u5_mult_87_CARRYB_50__2_), .CI(u5_mult_87_SUMB_50__3_), .CO(
        u5_mult_87_CARRYB_51__2_), .S(u5_mult_87_SUMB_51__2_) );
  FA_X1 u5_mult_87_S2_51_1 ( .A(u5_mult_87_ab_51__1_), .B(
        u5_mult_87_CARRYB_50__1_), .CI(u5_mult_87_SUMB_50__2_), .CO(
        u5_mult_87_CARRYB_51__1_), .S(u5_mult_87_SUMB_51__1_) );
  FA_X1 u5_mult_87_S1_51_0 ( .A(u5_mult_87_ab_51__0_), .B(
        u5_mult_87_CARRYB_50__0_), .CI(u5_mult_87_SUMB_50__1_), .CO(
        u5_mult_87_CARRYB_51__0_), .S(u5_N51) );
  FA_X1 u5_mult_87_S5_51 ( .A(u5_mult_87_ab_52__51_), .B(
        u5_mult_87_CARRYB_51__51_), .CI(u5_mult_87_ab_51__52_), .CO(
        u5_mult_87_CARRYB_52__51_), .S(u5_mult_87_SUMB_52__51_) );
  FA_X1 u5_mult_87_S4_50 ( .A(u5_mult_87_ab_52__50_), .B(
        u5_mult_87_CARRYB_51__50_), .CI(u5_mult_87_SUMB_51__51_), .CO(
        u5_mult_87_CARRYB_52__50_), .S(u5_mult_87_SUMB_52__50_) );
  FA_X1 u5_mult_87_S4_49 ( .A(u5_mult_87_ab_52__49_), .B(
        u5_mult_87_CARRYB_51__49_), .CI(u5_mult_87_SUMB_51__50_), .CO(
        u5_mult_87_CARRYB_52__49_), .S(u5_mult_87_SUMB_52__49_) );
  FA_X1 u5_mult_87_S4_48 ( .A(u5_mult_87_ab_52__48_), .B(
        u5_mult_87_CARRYB_51__48_), .CI(u5_mult_87_SUMB_51__49_), .CO(
        u5_mult_87_CARRYB_52__48_), .S(u5_mult_87_SUMB_52__48_) );
  FA_X1 u5_mult_87_S4_47 ( .A(u5_mult_87_ab_52__47_), .B(
        u5_mult_87_CARRYB_51__47_), .CI(u5_mult_87_SUMB_51__48_), .CO(
        u5_mult_87_CARRYB_52__47_), .S(u5_mult_87_SUMB_52__47_) );
  FA_X1 u5_mult_87_S4_46 ( .A(u5_mult_87_ab_52__46_), .B(
        u5_mult_87_CARRYB_51__46_), .CI(u5_mult_87_SUMB_51__47_), .CO(
        u5_mult_87_CARRYB_52__46_), .S(u5_mult_87_SUMB_52__46_) );
  FA_X1 u5_mult_87_S4_45 ( .A(u5_mult_87_ab_52__45_), .B(
        u5_mult_87_CARRYB_51__45_), .CI(u5_mult_87_SUMB_51__46_), .CO(
        u5_mult_87_CARRYB_52__45_), .S(u5_mult_87_SUMB_52__45_) );
  FA_X1 u5_mult_87_S4_44 ( .A(u5_mult_87_ab_52__44_), .B(
        u5_mult_87_CARRYB_51__44_), .CI(u5_mult_87_SUMB_51__45_), .CO(
        u5_mult_87_CARRYB_52__44_), .S(u5_mult_87_SUMB_52__44_) );
  FA_X1 u5_mult_87_S4_43 ( .A(u5_mult_87_ab_52__43_), .B(
        u5_mult_87_CARRYB_51__43_), .CI(u5_mult_87_SUMB_51__44_), .CO(
        u5_mult_87_CARRYB_52__43_), .S(u5_mult_87_SUMB_52__43_) );
  FA_X1 u5_mult_87_S4_42 ( .A(u5_mult_87_ab_52__42_), .B(
        u5_mult_87_CARRYB_51__42_), .CI(u5_mult_87_SUMB_51__43_), .CO(
        u5_mult_87_CARRYB_52__42_), .S(u5_mult_87_SUMB_52__42_) );
  FA_X1 u5_mult_87_S4_41 ( .A(u5_mult_87_ab_52__41_), .B(
        u5_mult_87_CARRYB_51__41_), .CI(u5_mult_87_SUMB_51__42_), .CO(
        u5_mult_87_CARRYB_52__41_), .S(u5_mult_87_SUMB_52__41_) );
  FA_X1 u5_mult_87_S4_40 ( .A(u5_mult_87_ab_52__40_), .B(
        u5_mult_87_CARRYB_51__40_), .CI(u5_mult_87_SUMB_51__41_), .CO(
        u5_mult_87_CARRYB_52__40_), .S(u5_mult_87_SUMB_52__40_) );
  FA_X1 u5_mult_87_S4_39 ( .A(u5_mult_87_ab_52__39_), .B(
        u5_mult_87_CARRYB_51__39_), .CI(u5_mult_87_SUMB_51__40_), .CO(
        u5_mult_87_CARRYB_52__39_), .S(u5_mult_87_SUMB_52__39_) );
  FA_X1 u5_mult_87_S4_38 ( .A(u5_mult_87_ab_52__38_), .B(
        u5_mult_87_CARRYB_51__38_), .CI(u5_mult_87_SUMB_51__39_), .CO(
        u5_mult_87_CARRYB_52__38_), .S(u5_mult_87_SUMB_52__38_) );
  FA_X1 u5_mult_87_S4_37 ( .A(u5_mult_87_ab_52__37_), .B(
        u5_mult_87_CARRYB_51__37_), .CI(u5_mult_87_SUMB_51__38_), .CO(
        u5_mult_87_CARRYB_52__37_), .S(u5_mult_87_SUMB_52__37_) );
  FA_X1 u5_mult_87_S4_36 ( .A(u5_mult_87_ab_52__36_), .B(
        u5_mult_87_CARRYB_51__36_), .CI(u5_mult_87_SUMB_51__37_), .CO(
        u5_mult_87_CARRYB_52__36_), .S(u5_mult_87_SUMB_52__36_) );
  FA_X1 u5_mult_87_S4_35 ( .A(u5_mult_87_ab_52__35_), .B(
        u5_mult_87_CARRYB_51__35_), .CI(u5_mult_87_SUMB_51__36_), .CO(
        u5_mult_87_CARRYB_52__35_), .S(u5_mult_87_SUMB_52__35_) );
  FA_X1 u5_mult_87_S4_34 ( .A(u5_mult_87_ab_52__34_), .B(
        u5_mult_87_CARRYB_51__34_), .CI(u5_mult_87_SUMB_51__35_), .CO(
        u5_mult_87_CARRYB_52__34_), .S(u5_mult_87_SUMB_52__34_) );
  FA_X1 u5_mult_87_S4_33 ( .A(u5_mult_87_ab_52__33_), .B(
        u5_mult_87_CARRYB_51__33_), .CI(u5_mult_87_SUMB_51__34_), .CO(
        u5_mult_87_CARRYB_52__33_), .S(u5_mult_87_SUMB_52__33_) );
  FA_X1 u5_mult_87_S4_32 ( .A(u5_mult_87_ab_52__32_), .B(
        u5_mult_87_CARRYB_51__32_), .CI(u5_mult_87_SUMB_51__33_), .CO(
        u5_mult_87_CARRYB_52__32_), .S(u5_mult_87_SUMB_52__32_) );
  FA_X1 u5_mult_87_S4_31 ( .A(u5_mult_87_ab_52__31_), .B(
        u5_mult_87_CARRYB_51__31_), .CI(u5_mult_87_SUMB_51__32_), .CO(
        u5_mult_87_CARRYB_52__31_), .S(u5_mult_87_SUMB_52__31_) );
  FA_X1 u5_mult_87_S4_30 ( .A(u5_mult_87_ab_52__30_), .B(
        u5_mult_87_CARRYB_51__30_), .CI(u5_mult_87_SUMB_51__31_), .CO(
        u5_mult_87_CARRYB_52__30_), .S(u5_mult_87_SUMB_52__30_) );
  FA_X1 u5_mult_87_S4_29 ( .A(u5_mult_87_ab_52__29_), .B(
        u5_mult_87_CARRYB_51__29_), .CI(u5_mult_87_SUMB_51__30_), .CO(
        u5_mult_87_CARRYB_52__29_), .S(u5_mult_87_SUMB_52__29_) );
  FA_X1 u5_mult_87_S4_28 ( .A(u5_mult_87_ab_52__28_), .B(
        u5_mult_87_CARRYB_51__28_), .CI(u5_mult_87_SUMB_51__29_), .CO(
        u5_mult_87_CARRYB_52__28_), .S(u5_mult_87_SUMB_52__28_) );
  FA_X1 u5_mult_87_S4_27 ( .A(u5_mult_87_ab_52__27_), .B(
        u5_mult_87_CARRYB_51__27_), .CI(u5_mult_87_SUMB_51__28_), .CO(
        u5_mult_87_CARRYB_52__27_), .S(u5_mult_87_SUMB_52__27_) );
  FA_X1 u5_mult_87_S4_26 ( .A(u5_mult_87_ab_52__26_), .B(
        u5_mult_87_CARRYB_51__26_), .CI(u5_mult_87_SUMB_51__27_), .CO(
        u5_mult_87_CARRYB_52__26_), .S(u5_mult_87_SUMB_52__26_) );
  FA_X1 u5_mult_87_S4_25 ( .A(u5_mult_87_ab_52__25_), .B(
        u5_mult_87_CARRYB_51__25_), .CI(u5_mult_87_SUMB_51__26_), .CO(
        u5_mult_87_CARRYB_52__25_), .S(u5_mult_87_SUMB_52__25_) );
  FA_X1 u5_mult_87_S4_24 ( .A(u5_mult_87_ab_52__24_), .B(
        u5_mult_87_CARRYB_51__24_), .CI(u5_mult_87_SUMB_51__25_), .CO(
        u5_mult_87_CARRYB_52__24_), .S(u5_mult_87_SUMB_52__24_) );
  FA_X1 u5_mult_87_S4_23 ( .A(u5_mult_87_ab_52__23_), .B(
        u5_mult_87_CARRYB_51__23_), .CI(u5_mult_87_SUMB_51__24_), .CO(
        u5_mult_87_CARRYB_52__23_), .S(u5_mult_87_SUMB_52__23_) );
  FA_X1 u5_mult_87_S4_22 ( .A(u5_mult_87_ab_52__22_), .B(
        u5_mult_87_CARRYB_51__22_), .CI(u5_mult_87_SUMB_51__23_), .CO(
        u5_mult_87_CARRYB_52__22_), .S(u5_mult_87_SUMB_52__22_) );
  FA_X1 u5_mult_87_S4_21 ( .A(u5_mult_87_ab_52__21_), .B(
        u5_mult_87_CARRYB_51__21_), .CI(u5_mult_87_SUMB_51__22_), .CO(
        u5_mult_87_CARRYB_52__21_), .S(u5_mult_87_SUMB_52__21_) );
  FA_X1 u5_mult_87_S4_20 ( .A(u5_mult_87_ab_52__20_), .B(
        u5_mult_87_CARRYB_51__20_), .CI(u5_mult_87_SUMB_51__21_), .CO(
        u5_mult_87_CARRYB_52__20_), .S(u5_mult_87_SUMB_52__20_) );
  FA_X1 u5_mult_87_S4_19 ( .A(u5_mult_87_ab_52__19_), .B(
        u5_mult_87_CARRYB_51__19_), .CI(u5_mult_87_SUMB_51__20_), .CO(
        u5_mult_87_CARRYB_52__19_), .S(u5_mult_87_SUMB_52__19_) );
  FA_X1 u5_mult_87_S4_18 ( .A(u5_mult_87_ab_52__18_), .B(
        u5_mult_87_CARRYB_51__18_), .CI(u5_mult_87_SUMB_51__19_), .CO(
        u5_mult_87_CARRYB_52__18_), .S(u5_mult_87_SUMB_52__18_) );
  FA_X1 u5_mult_87_S4_17 ( .A(u5_mult_87_ab_52__17_), .B(
        u5_mult_87_CARRYB_51__17_), .CI(u5_mult_87_SUMB_51__18_), .CO(
        u5_mult_87_CARRYB_52__17_), .S(u5_mult_87_SUMB_52__17_) );
  FA_X1 u5_mult_87_S4_16 ( .A(u5_mult_87_ab_52__16_), .B(
        u5_mult_87_CARRYB_51__16_), .CI(u5_mult_87_SUMB_51__17_), .CO(
        u5_mult_87_CARRYB_52__16_), .S(u5_mult_87_SUMB_52__16_) );
  FA_X1 u5_mult_87_S4_15 ( .A(u5_mult_87_ab_52__15_), .B(
        u5_mult_87_CARRYB_51__15_), .CI(u5_mult_87_SUMB_51__16_), .CO(
        u5_mult_87_CARRYB_52__15_), .S(u5_mult_87_SUMB_52__15_) );
  FA_X1 u5_mult_87_S4_14 ( .A(u5_mult_87_ab_52__14_), .B(
        u5_mult_87_CARRYB_51__14_), .CI(u5_mult_87_SUMB_51__15_), .CO(
        u5_mult_87_CARRYB_52__14_), .S(u5_mult_87_SUMB_52__14_) );
  FA_X1 u5_mult_87_S4_13 ( .A(u5_mult_87_ab_52__13_), .B(
        u5_mult_87_CARRYB_51__13_), .CI(u5_mult_87_SUMB_51__14_), .CO(
        u5_mult_87_CARRYB_52__13_), .S(u5_mult_87_SUMB_52__13_) );
  FA_X1 u5_mult_87_S4_12 ( .A(u5_mult_87_ab_52__12_), .B(
        u5_mult_87_CARRYB_51__12_), .CI(u5_mult_87_SUMB_51__13_), .CO(
        u5_mult_87_CARRYB_52__12_), .S(u5_mult_87_SUMB_52__12_) );
  FA_X1 u5_mult_87_S4_11 ( .A(u5_mult_87_ab_52__11_), .B(
        u5_mult_87_CARRYB_51__11_), .CI(u5_mult_87_SUMB_51__12_), .CO(
        u5_mult_87_CARRYB_52__11_), .S(u5_mult_87_SUMB_52__11_) );
  FA_X1 u5_mult_87_S4_10 ( .A(u5_mult_87_ab_52__10_), .B(
        u5_mult_87_CARRYB_51__10_), .CI(u5_mult_87_SUMB_51__11_), .CO(
        u5_mult_87_CARRYB_52__10_), .S(u5_mult_87_SUMB_52__10_) );
  FA_X1 u5_mult_87_S4_9 ( .A(u5_mult_87_ab_52__9_), .B(
        u5_mult_87_CARRYB_51__9_), .CI(u5_mult_87_SUMB_51__10_), .CO(
        u5_mult_87_CARRYB_52__9_), .S(u5_mult_87_SUMB_52__9_) );
  FA_X1 u5_mult_87_S4_8 ( .A(u5_mult_87_ab_52__8_), .B(
        u5_mult_87_CARRYB_51__8_), .CI(u5_mult_87_SUMB_51__9_), .CO(
        u5_mult_87_CARRYB_52__8_), .S(u5_mult_87_SUMB_52__8_) );
  FA_X1 u5_mult_87_S4_7 ( .A(u5_mult_87_ab_52__7_), .B(
        u5_mult_87_CARRYB_51__7_), .CI(u5_mult_87_SUMB_51__8_), .CO(
        u5_mult_87_CARRYB_52__7_), .S(u5_mult_87_SUMB_52__7_) );
  FA_X1 u5_mult_87_S4_6 ( .A(u5_mult_87_ab_52__6_), .B(
        u5_mult_87_CARRYB_51__6_), .CI(u5_mult_87_SUMB_51__7_), .CO(
        u5_mult_87_CARRYB_52__6_), .S(u5_mult_87_SUMB_52__6_) );
  FA_X1 u5_mult_87_S4_5 ( .A(u5_mult_87_ab_52__5_), .B(
        u5_mult_87_CARRYB_51__5_), .CI(u5_mult_87_SUMB_51__6_), .CO(
        u5_mult_87_CARRYB_52__5_), .S(u5_mult_87_SUMB_52__5_) );
  FA_X1 u5_mult_87_S4_4 ( .A(u5_mult_87_ab_52__4_), .B(
        u5_mult_87_CARRYB_51__4_), .CI(u5_mult_87_SUMB_51__5_), .CO(
        u5_mult_87_CARRYB_52__4_), .S(u5_mult_87_SUMB_52__4_) );
  FA_X1 u5_mult_87_S4_3 ( .A(u5_mult_87_ab_52__3_), .B(
        u5_mult_87_CARRYB_51__3_), .CI(u5_mult_87_SUMB_51__4_), .CO(
        u5_mult_87_CARRYB_52__3_), .S(u5_mult_87_SUMB_52__3_) );
  FA_X1 u5_mult_87_S4_2 ( .A(u5_mult_87_ab_52__2_), .B(
        u5_mult_87_CARRYB_51__2_), .CI(u5_mult_87_SUMB_51__3_), .CO(
        u5_mult_87_CARRYB_52__2_), .S(u5_mult_87_SUMB_52__2_) );
  FA_X1 u5_mult_87_S4_1 ( .A(u5_mult_87_ab_52__1_), .B(
        u5_mult_87_CARRYB_51__1_), .CI(u5_mult_87_SUMB_51__2_), .CO(
        u5_mult_87_CARRYB_52__1_), .S(u5_mult_87_SUMB_52__1_) );
  FA_X1 u5_mult_87_S4_0 ( .A(u5_mult_87_ab_52__0_), .B(
        u5_mult_87_CARRYB_51__0_), .CI(u5_mult_87_SUMB_51__1_), .CO(
        u5_mult_87_CARRYB_52__0_), .S(u5_N52) );
  NOR2_X1 u5_mult_87_FS_1_U383 ( .A1(u5_mult_87_n205), .A2(u5_mult_87_n103), 
        .ZN(u5_mult_87_FS_1_n284) );
  NOR2_X1 u5_mult_87_FS_1_U382 ( .A1(u5_mult_87_n204), .A2(u5_mult_87_n102), 
        .ZN(u5_mult_87_FS_1_n84) );
  NAND2_X1 u5_mult_87_FS_1_U381 ( .A1(u5_mult_87_n189), .A2(u5_mult_87_n96), 
        .ZN(u5_mult_87_FS_1_n89) );
  NAND2_X1 u5_mult_87_FS_1_U380 ( .A1(u5_mult_87_n204), .A2(u5_mult_87_n102), 
        .ZN(u5_mult_87_FS_1_n85) );
  OAI21_X1 u5_mult_87_FS_1_U379 ( .B1(u5_mult_87_FS_1_n84), .B2(
        u5_mult_87_FS_1_n89), .A(u5_mult_87_FS_1_n85), .ZN(
        u5_mult_87_FS_1_n331) );
  NAND2_X1 u5_mult_87_FS_1_U378 ( .A1(u5_mult_87_n205), .A2(u5_mult_87_n103), 
        .ZN(u5_mult_87_FS_1_n86) );
  AOI21_X1 u5_mult_87_FS_1_U377 ( .B1(u5_mult_87_FS_1_n9), .B2(
        u5_mult_87_FS_1_n331), .A(u5_mult_87_FS_1_n8), .ZN(
        u5_mult_87_FS_1_n282) );
  NOR2_X1 u5_mult_87_FS_1_U376 ( .A1(u5_mult_87_n95), .A2(u5_mult_87_n206), 
        .ZN(u5_mult_87_FS_1_n79) );
  NOR2_X1 u5_mult_87_FS_1_U375 ( .A1(u5_mult_87_n187), .A2(u5_mult_87_n90), 
        .ZN(u5_mult_87_FS_1_n139) );
  NOR2_X1 u5_mult_87_FS_1_U374 ( .A1(u5_mult_87_n203), .A2(u5_mult_87_n89), 
        .ZN(u5_mult_87_FS_1_n132) );
  NOR2_X1 u5_mult_87_FS_1_U373 ( .A1(u5_mult_87_n193), .A2(u5_mult_87_n62), 
        .ZN(u5_mult_87_FS_1_n134) );
  NOR2_X1 u5_mult_87_FS_1_U372 ( .A1(u5_mult_87_n186), .A2(u5_mult_87_n88), 
        .ZN(u5_mult_87_FS_1_n136) );
  NOR4_X1 u5_mult_87_FS_1_U371 ( .A1(u5_mult_87_FS_1_n139), .A2(
        u5_mult_87_FS_1_n132), .A3(u5_mult_87_FS_1_n134), .A4(
        u5_mult_87_FS_1_n136), .ZN(u5_mult_87_FS_1_n125) );
  NOR2_X1 u5_mult_87_FS_1_U370 ( .A1(u5_mult_87_n202), .A2(u5_mult_87_n87), 
        .ZN(u5_mult_87_FS_1_n121) );
  NOR2_X1 u5_mult_87_FS_1_U369 ( .A1(u5_mult_87_n201), .A2(u5_mult_87_n101), 
        .ZN(u5_mult_87_FS_1_n111) );
  NOR2_X1 u5_mult_87_FS_1_U368 ( .A1(u5_mult_87_n200), .A2(u5_mult_87_n86), 
        .ZN(u5_mult_87_FS_1_n114) );
  NOR2_X1 u5_mult_87_FS_1_U367 ( .A1(u5_mult_87_n199), .A2(u5_mult_87_n85), 
        .ZN(u5_mult_87_FS_1_n118) );
  NOR4_X1 u5_mult_87_FS_1_U366 ( .A1(u5_mult_87_FS_1_n121), .A2(
        u5_mult_87_FS_1_n111), .A3(u5_mult_87_FS_1_n114), .A4(
        u5_mult_87_FS_1_n118), .ZN(u5_mult_87_FS_1_n293) );
  NOR2_X1 u5_mult_87_FS_1_U365 ( .A1(u5_mult_87_n198), .A2(u5_mult_87_n100), 
        .ZN(u5_mult_87_FS_1_n105) );
  NOR2_X1 u5_mult_87_FS_1_U364 ( .A1(u5_mult_87_n197), .A2(u5_mult_87_n99), 
        .ZN(u5_mult_87_FS_1_n300) );
  NOR2_X1 u5_mult_87_FS_1_U363 ( .A1(u5_mult_87_n192), .A2(u5_mult_87_n94), 
        .ZN(u5_mult_87_FS_1_n99) );
  NOR2_X1 u5_mult_87_FS_1_U362 ( .A1(u5_mult_87_n196), .A2(u5_mult_87_n98), 
        .ZN(u5_mult_87_FS_1_n101) );
  NOR4_X1 u5_mult_87_FS_1_U361 ( .A1(u5_mult_87_FS_1_n105), .A2(
        u5_mult_87_FS_1_n300), .A3(u5_mult_87_FS_1_n99), .A4(
        u5_mult_87_FS_1_n101), .ZN(u5_mult_87_FS_1_n287) );
  NOR2_X1 u5_mult_87_FS_1_U360 ( .A1(u5_mult_87_n185), .A2(u5_mult_87_n84), 
        .ZN(u5_mult_87_FS_1_n153) );
  NOR2_X1 u5_mult_87_FS_1_U359 ( .A1(u5_mult_87_n184), .A2(u5_mult_87_n83), 
        .ZN(u5_mult_87_FS_1_n206) );
  NOR2_X1 u5_mult_87_FS_1_U358 ( .A1(u5_mult_87_n183), .A2(u5_mult_87_n82), 
        .ZN(u5_mult_87_FS_1_n199) );
  NOR2_X1 u5_mult_87_FS_1_U357 ( .A1(u5_mult_87_n162), .A2(u5_mult_87_n61), 
        .ZN(u5_mult_87_FS_1_n201) );
  NOR2_X1 u5_mult_87_FS_1_U356 ( .A1(u5_mult_87_n182), .A2(u5_mult_87_n81), 
        .ZN(u5_mult_87_FS_1_n203) );
  NOR4_X1 u5_mult_87_FS_1_U355 ( .A1(u5_mult_87_FS_1_n206), .A2(
        u5_mult_87_FS_1_n199), .A3(u5_mult_87_FS_1_n201), .A4(
        u5_mult_87_FS_1_n203), .ZN(u5_mult_87_FS_1_n192) );
  NOR2_X1 u5_mult_87_FS_1_U354 ( .A1(u5_mult_87_n181), .A2(u5_mult_87_n80), 
        .ZN(u5_mult_87_FS_1_n188) );
  NOR2_X1 u5_mult_87_FS_1_U353 ( .A1(u5_mult_87_n180), .A2(u5_mult_87_n79), 
        .ZN(u5_mult_87_FS_1_n178) );
  NOR2_X1 u5_mult_87_FS_1_U352 ( .A1(u5_mult_87_n179), .A2(u5_mult_87_n78), 
        .ZN(u5_mult_87_FS_1_n181) );
  NOR2_X1 u5_mult_87_FS_1_U351 ( .A1(u5_mult_87_n178), .A2(u5_mult_87_n77), 
        .ZN(u5_mult_87_FS_1_n185) );
  NOR4_X1 u5_mult_87_FS_1_U350 ( .A1(u5_mult_87_FS_1_n188), .A2(
        u5_mult_87_FS_1_n178), .A3(u5_mult_87_FS_1_n181), .A4(
        u5_mult_87_FS_1_n185), .ZN(u5_mult_87_FS_1_n310) );
  NOR2_X1 u5_mult_87_FS_1_U349 ( .A1(u5_mult_87_n177), .A2(u5_mult_87_n76), 
        .ZN(u5_mult_87_FS_1_n172) );
  NOR2_X1 u5_mult_87_FS_1_U348 ( .A1(u5_mult_87_n176), .A2(u5_mult_87_n75), 
        .ZN(u5_mult_87_FS_1_n317) );
  NOR2_X1 u5_mult_87_FS_1_U347 ( .A1(u5_mult_87_n161), .A2(u5_mult_87_n60), 
        .ZN(u5_mult_87_FS_1_n166) );
  NOR2_X1 u5_mult_87_FS_1_U346 ( .A1(u5_mult_87_n175), .A2(u5_mult_87_n74), 
        .ZN(u5_mult_87_FS_1_n168) );
  NOR4_X1 u5_mult_87_FS_1_U345 ( .A1(u5_mult_87_FS_1_n172), .A2(
        u5_mult_87_FS_1_n317), .A3(u5_mult_87_FS_1_n166), .A4(
        u5_mult_87_FS_1_n168), .ZN(u5_mult_87_FS_1_n304) );
  NOR2_X1 u5_mult_87_FS_1_U344 ( .A1(u5_mult_87_n174), .A2(u5_mult_87_n73), 
        .ZN(u5_mult_87_FS_1_n220) );
  OR2_X1 u5_mult_87_FS_1_U343 ( .A1(u5_mult_87_n158), .A2(u5_mult_87_n63), 
        .ZN(u5_mult_87_FS_1_n231) );
  NOR2_X1 u5_mult_87_FS_1_U342 ( .A1(u5_mult_87_n173), .A2(u5_mult_87_n72), 
        .ZN(u5_mult_87_FS_1_n234) );
  NAND2_X1 u5_mult_87_FS_1_U341 ( .A1(u5_mult_87_n172), .A2(u5_mult_87_n71), 
        .ZN(u5_mult_87_FS_1_n241) );
  NAND2_X1 u5_mult_87_FS_1_U340 ( .A1(u5_mult_87_n173), .A2(u5_mult_87_n72), 
        .ZN(u5_mult_87_FS_1_n235) );
  OAI21_X1 u5_mult_87_FS_1_U339 ( .B1(u5_mult_87_FS_1_n234), .B2(
        u5_mult_87_FS_1_n241), .A(u5_mult_87_FS_1_n235), .ZN(
        u5_mult_87_FS_1_n330) );
  NAND2_X1 u5_mult_87_FS_1_U338 ( .A1(u5_mult_87_n158), .A2(u5_mult_87_n63), 
        .ZN(u5_mult_87_FS_1_n236) );
  AOI21_X1 u5_mult_87_FS_1_U337 ( .B1(u5_mult_87_FS_1_n231), .B2(
        u5_mult_87_FS_1_n330), .A(u5_mult_87_FS_1_n62), .ZN(
        u5_mult_87_FS_1_n319) );
  NOR2_X1 u5_mult_87_FS_1_U336 ( .A1(u5_mult_87_n171), .A2(u5_mult_87_n70), 
        .ZN(u5_mult_87_FS_1_n320) );
  NAND2_X1 u5_mult_87_FS_1_U335 ( .A1(u5_mult_87_n171), .A2(u5_mult_87_n70), 
        .ZN(u5_mult_87_FS_1_n229) );
  NOR2_X1 u5_mult_87_FS_1_U334 ( .A1(u5_mult_87_n160), .A2(u5_mult_87_n4), 
        .ZN(u5_mult_87_FS_1_n248) );
  NOR2_X1 u5_mult_87_FS_1_U333 ( .A1(u5_mult_87_n170), .A2(u5_mult_87_n10), 
        .ZN(u5_mult_87_FS_1_n250) );
  NAND2_X1 u5_mult_87_FS_1_U332 ( .A1(u5_mult_87_n169), .A2(u5_mult_87_n9), 
        .ZN(u5_mult_87_FS_1_n256) );
  NAND2_X1 u5_mult_87_FS_1_U331 ( .A1(u5_mult_87_n170), .A2(u5_mult_87_n10), 
        .ZN(u5_mult_87_FS_1_n251) );
  OAI21_X1 u5_mult_87_FS_1_U330 ( .B1(u5_mult_87_FS_1_n250), .B2(
        u5_mult_87_FS_1_n256), .A(u5_mult_87_FS_1_n251), .ZN(
        u5_mult_87_FS_1_n329) );
  AND2_X1 u5_mult_87_FS_1_U329 ( .A1(u5_mult_87_n160), .A2(u5_mult_87_n4), 
        .ZN(u5_mult_87_FS_1_n245) );
  AOI21_X1 u5_mult_87_FS_1_U328 ( .B1(u5_mult_87_FS_1_n67), .B2(
        u5_mult_87_FS_1_n329), .A(u5_mult_87_FS_1_n245), .ZN(
        u5_mult_87_FS_1_n323) );
  NOR2_X1 u5_mult_87_FS_1_U327 ( .A1(u5_mult_87_n168), .A2(u5_mult_87_n69), 
        .ZN(u5_mult_87_FS_1_n324) );
  NOR2_X1 u5_mult_87_FS_1_U326 ( .A1(u5_mult_87_n107), .A2(u5_mult_87_n8), 
        .ZN(u5_mult_87_FS_1_n262) );
  NOR2_X1 u5_mult_87_FS_1_U325 ( .A1(u5_mult_87_n106), .A2(u5_mult_87_n7), 
        .ZN(u5_mult_87_FS_1_n265) );
  NAND2_X1 u5_mult_87_FS_1_U324 ( .A1(u5_mult_87_n105), .A2(u5_mult_87_n5), 
        .ZN(u5_mult_87_FS_1_n268) );
  NAND2_X1 u5_mult_87_FS_1_U323 ( .A1(u5_mult_87_n106), .A2(u5_mult_87_n7), 
        .ZN(u5_mult_87_FS_1_n267) );
  OAI21_X1 u5_mult_87_FS_1_U322 ( .B1(u5_mult_87_FS_1_n265), .B2(
        u5_mult_87_FS_1_n268), .A(u5_mult_87_FS_1_n267), .ZN(
        u5_mult_87_FS_1_n328) );
  NAND2_X1 u5_mult_87_FS_1_U321 ( .A1(u5_mult_87_n107), .A2(u5_mult_87_n8), 
        .ZN(u5_mult_87_FS_1_n263) );
  AOI21_X1 u5_mult_87_FS_1_U320 ( .B1(u5_mult_87_FS_1_n73), .B2(
        u5_mult_87_FS_1_n328), .A(u5_mult_87_FS_1_n72), .ZN(
        u5_mult_87_FS_1_n327) );
  NOR2_X1 u5_mult_87_FS_1_U319 ( .A1(u5_mult_87_n167), .A2(u5_mult_87_n6), 
        .ZN(u5_mult_87_FS_1_n259) );
  NAND2_X1 u5_mult_87_FS_1_U318 ( .A1(u5_mult_87_n167), .A2(u5_mult_87_n6), 
        .ZN(u5_mult_87_FS_1_n260) );
  NAND3_X1 u5_mult_87_FS_1_U317 ( .A1(u5_mult_87_FS_1_n66), .A2(
        u5_mult_87_FS_1_n253), .A3(u5_mult_87_FS_1_n67), .ZN(
        u5_mult_87_FS_1_n325) );
  NOR2_X1 u5_mult_87_FS_1_U316 ( .A1(u5_mult_87_n169), .A2(u5_mult_87_n9), 
        .ZN(u5_mult_87_FS_1_n255) );
  NAND2_X1 u5_mult_87_FS_1_U315 ( .A1(u5_mult_87_FS_1_n69), .A2(
        u5_mult_87_FS_1_n68), .ZN(u5_mult_87_FS_1_n326) );
  NAND2_X1 u5_mult_87_FS_1_U314 ( .A1(u5_mult_87_n168), .A2(u5_mult_87_n69), 
        .ZN(u5_mult_87_FS_1_n246) );
  OAI221_X1 u5_mult_87_FS_1_U313 ( .B1(u5_mult_87_FS_1_n323), .B2(
        u5_mult_87_FS_1_n324), .C1(u5_mult_87_FS_1_n325), .C2(
        u5_mult_87_FS_1_n326), .A(u5_mult_87_FS_1_n246), .ZN(
        u5_mult_87_FS_1_n322) );
  NOR2_X1 u5_mult_87_FS_1_U312 ( .A1(u5_mult_87_n172), .A2(u5_mult_87_n71), 
        .ZN(u5_mult_87_FS_1_n240) );
  NOR2_X1 u5_mult_87_FS_1_U311 ( .A1(u5_mult_87_FS_1_n65), .A2(
        u5_mult_87_FS_1_n240), .ZN(u5_mult_87_FS_1_n238) );
  NAND4_X1 u5_mult_87_FS_1_U310 ( .A1(u5_mult_87_FS_1_n238), .A2(
        u5_mult_87_FS_1_n63), .A3(u5_mult_87_FS_1_n231), .A4(
        u5_mult_87_FS_1_n61), .ZN(u5_mult_87_FS_1_n321) );
  OAI211_X1 u5_mult_87_FS_1_U309 ( .C1(u5_mult_87_FS_1_n319), .C2(
        u5_mult_87_FS_1_n320), .A(u5_mult_87_FS_1_n229), .B(
        u5_mult_87_FS_1_n321), .ZN(u5_mult_87_FS_1_n226) );
  NOR2_X1 u5_mult_87_FS_1_U308 ( .A1(u5_mult_87_n166), .A2(u5_mult_87_n68), 
        .ZN(u5_mult_87_FS_1_n216) );
  NOR2_X1 u5_mult_87_FS_1_U307 ( .A1(u5_mult_87_n165), .A2(u5_mult_87_n67), 
        .ZN(u5_mult_87_FS_1_n213) );
  NOR2_X1 u5_mult_87_FS_1_U306 ( .A1(u5_mult_87_n164), .A2(u5_mult_87_n66), 
        .ZN(u5_mult_87_FS_1_n223) );
  OR2_X1 u5_mult_87_FS_1_U305 ( .A1(u5_mult_87_FS_1_n213), .A2(
        u5_mult_87_FS_1_n223), .ZN(u5_mult_87_FS_1_n318) );
  NOR4_X1 u5_mult_87_FS_1_U304 ( .A1(u5_mult_87_FS_1_n220), .A2(
        u5_mult_87_FS_1_n60), .A3(u5_mult_87_FS_1_n216), .A4(
        u5_mult_87_FS_1_n318), .ZN(u5_mult_87_FS_1_n210) );
  NAND4_X1 u5_mult_87_FS_1_U303 ( .A1(u5_mult_87_FS_1_n192), .A2(
        u5_mult_87_FS_1_n310), .A3(u5_mult_87_FS_1_n304), .A4(
        u5_mult_87_FS_1_n210), .ZN(u5_mult_87_FS_1_n302) );
  NAND2_X1 u5_mult_87_FS_1_U302 ( .A1(u5_mult_87_n176), .A2(u5_mult_87_n75), 
        .ZN(u5_mult_87_FS_1_n164) );
  NAND2_X1 u5_mult_87_FS_1_U301 ( .A1(u5_mult_87_n177), .A2(u5_mult_87_n76), 
        .ZN(u5_mult_87_FS_1_n174) );
  NAND2_X1 u5_mult_87_FS_1_U300 ( .A1(u5_mult_87_n175), .A2(u5_mult_87_n74), 
        .ZN(u5_mult_87_FS_1_n169) );
  OAI21_X1 u5_mult_87_FS_1_U299 ( .B1(u5_mult_87_FS_1_n174), .B2(
        u5_mult_87_FS_1_n168), .A(u5_mult_87_FS_1_n169), .ZN(
        u5_mult_87_FS_1_n316) );
  AND2_X1 u5_mult_87_FS_1_U298 ( .A1(u5_mult_87_n161), .A2(u5_mult_87_n60), 
        .ZN(u5_mult_87_FS_1_n163) );
  AOI21_X1 u5_mult_87_FS_1_U297 ( .B1(u5_mult_87_FS_1_n316), .B2(
        u5_mult_87_FS_1_n37), .A(u5_mult_87_FS_1_n163), .ZN(
        u5_mult_87_FS_1_n315) );
  NAND2_X1 u5_mult_87_FS_1_U296 ( .A1(u5_mult_87_n164), .A2(u5_mult_87_n66), 
        .ZN(u5_mult_87_FS_1_n224) );
  NAND2_X1 u5_mult_87_FS_1_U295 ( .A1(u5_mult_87_n174), .A2(u5_mult_87_n73), 
        .ZN(u5_mult_87_FS_1_n222) );
  OAI21_X1 u5_mult_87_FS_1_U294 ( .B1(u5_mult_87_FS_1_n220), .B2(
        u5_mult_87_FS_1_n224), .A(u5_mult_87_FS_1_n222), .ZN(
        u5_mult_87_FS_1_n314) );
  NAND2_X1 u5_mult_87_FS_1_U293 ( .A1(u5_mult_87_n166), .A2(u5_mult_87_n68), 
        .ZN(u5_mult_87_FS_1_n217) );
  AOI21_X1 u5_mult_87_FS_1_U292 ( .B1(u5_mult_87_FS_1_n56), .B2(
        u5_mult_87_FS_1_n314), .A(u5_mult_87_FS_1_n55), .ZN(
        u5_mult_87_FS_1_n313) );
  NAND2_X1 u5_mult_87_FS_1_U291 ( .A1(u5_mult_87_n165), .A2(u5_mult_87_n67), 
        .ZN(u5_mult_87_FS_1_n214) );
  OAI21_X1 u5_mult_87_FS_1_U290 ( .B1(u5_mult_87_FS_1_n313), .B2(
        u5_mult_87_FS_1_n213), .A(u5_mult_87_FS_1_n214), .ZN(
        u5_mult_87_FS_1_n209) );
  NAND2_X1 u5_mult_87_FS_1_U289 ( .A1(u5_mult_87_n184), .A2(u5_mult_87_n83), 
        .ZN(u5_mult_87_FS_1_n208) );
  NAND2_X1 u5_mult_87_FS_1_U288 ( .A1(u5_mult_87_n182), .A2(u5_mult_87_n81), 
        .ZN(u5_mult_87_FS_1_n204) );
  OAI21_X1 u5_mult_87_FS_1_U287 ( .B1(u5_mult_87_FS_1_n203), .B2(
        u5_mult_87_FS_1_n208), .A(u5_mult_87_FS_1_n204), .ZN(
        u5_mult_87_FS_1_n312) );
  AND2_X1 u5_mult_87_FS_1_U286 ( .A1(u5_mult_87_n162), .A2(u5_mult_87_n61), 
        .ZN(u5_mult_87_FS_1_n197) );
  AOI21_X1 u5_mult_87_FS_1_U285 ( .B1(u5_mult_87_FS_1_n50), .B2(
        u5_mult_87_FS_1_n312), .A(u5_mult_87_FS_1_n197), .ZN(
        u5_mult_87_FS_1_n311) );
  NAND2_X1 u5_mult_87_FS_1_U284 ( .A1(u5_mult_87_n183), .A2(u5_mult_87_n82), 
        .ZN(u5_mult_87_FS_1_n198) );
  OAI21_X1 u5_mult_87_FS_1_U283 ( .B1(u5_mult_87_FS_1_n311), .B2(
        u5_mult_87_FS_1_n199), .A(u5_mult_87_FS_1_n198), .ZN(
        u5_mult_87_FS_1_n193) );
  AOI21_X1 u5_mult_87_FS_1_U282 ( .B1(u5_mult_87_FS_1_n192), .B2(
        u5_mult_87_FS_1_n209), .A(u5_mult_87_FS_1_n193), .ZN(
        u5_mult_87_FS_1_n306) );
  NAND2_X1 u5_mult_87_FS_1_U281 ( .A1(u5_mult_87_n181), .A2(u5_mult_87_n80), 
        .ZN(u5_mult_87_FS_1_n189) );
  NAND2_X1 u5_mult_87_FS_1_U280 ( .A1(u5_mult_87_n178), .A2(u5_mult_87_n77), 
        .ZN(u5_mult_87_FS_1_n187) );
  OAI21_X1 u5_mult_87_FS_1_U279 ( .B1(u5_mult_87_FS_1_n185), .B2(
        u5_mult_87_FS_1_n189), .A(u5_mult_87_FS_1_n187), .ZN(
        u5_mult_87_FS_1_n309) );
  NAND2_X1 u5_mult_87_FS_1_U278 ( .A1(u5_mult_87_n179), .A2(u5_mult_87_n78), 
        .ZN(u5_mult_87_FS_1_n182) );
  AOI21_X1 u5_mult_87_FS_1_U277 ( .B1(u5_mult_87_FS_1_n45), .B2(
        u5_mult_87_FS_1_n309), .A(u5_mult_87_FS_1_n44), .ZN(
        u5_mult_87_FS_1_n308) );
  NAND2_X1 u5_mult_87_FS_1_U276 ( .A1(u5_mult_87_n180), .A2(u5_mult_87_n79), 
        .ZN(u5_mult_87_FS_1_n179) );
  OAI21_X1 u5_mult_87_FS_1_U275 ( .B1(u5_mult_87_FS_1_n308), .B2(
        u5_mult_87_FS_1_n178), .A(u5_mult_87_FS_1_n179), .ZN(
        u5_mult_87_FS_1_n307) );
  OAI21_X1 u5_mult_87_FS_1_U274 ( .B1(u5_mult_87_FS_1_n306), .B2(
        u5_mult_87_FS_1_n43), .A(u5_mult_87_FS_1_n41), .ZN(
        u5_mult_87_FS_1_n305) );
  AOI22_X1 u5_mult_87_FS_1_U273 ( .A1(u5_mult_87_FS_1_n35), .A2(
        u5_mult_87_FS_1_n36), .B1(u5_mult_87_FS_1_n304), .B2(
        u5_mult_87_FS_1_n305), .ZN(u5_mult_87_FS_1_n303) );
  NAND3_X1 u5_mult_87_FS_1_U272 ( .A1(u5_mult_87_FS_1_n302), .A2(
        u5_mult_87_FS_1_n164), .A3(u5_mult_87_FS_1_n303), .ZN(
        u5_mult_87_FS_1_n156) );
  NOR2_X1 u5_mult_87_FS_1_U271 ( .A1(u5_mult_87_n159), .A2(u5_mult_87_n59), 
        .ZN(u5_mult_87_FS_1_n151) );
  NOR2_X1 u5_mult_87_FS_1_U270 ( .A1(u5_mult_87_n195), .A2(u5_mult_87_n65), 
        .ZN(u5_mult_87_FS_1_n149) );
  NOR2_X1 u5_mult_87_FS_1_U269 ( .A1(u5_mult_87_n163), .A2(u5_mult_87_n64), 
        .ZN(u5_mult_87_FS_1_n157) );
  NOR2_X1 u5_mult_87_FS_1_U268 ( .A1(u5_mult_87_FS_1_n149), .A2(
        u5_mult_87_FS_1_n157), .ZN(u5_mult_87_FS_1_n301) );
  AND4_X1 u5_mult_87_FS_1_U267 ( .A1(u5_mult_87_FS_1_n32), .A2(
        u5_mult_87_FS_1_n156), .A3(u5_mult_87_FS_1_n31), .A4(
        u5_mult_87_FS_1_n301), .ZN(u5_mult_87_FS_1_n143) );
  NAND4_X1 u5_mult_87_FS_1_U266 ( .A1(u5_mult_87_FS_1_n125), .A2(
        u5_mult_87_FS_1_n293), .A3(u5_mult_87_FS_1_n287), .A4(
        u5_mult_87_FS_1_n143), .ZN(u5_mult_87_FS_1_n285) );
  NAND2_X1 u5_mult_87_FS_1_U265 ( .A1(u5_mult_87_n197), .A2(u5_mult_87_n99), 
        .ZN(u5_mult_87_FS_1_n97) );
  NAND2_X1 u5_mult_87_FS_1_U264 ( .A1(u5_mult_87_n198), .A2(u5_mult_87_n100), 
        .ZN(u5_mult_87_FS_1_n107) );
  NAND2_X1 u5_mult_87_FS_1_U263 ( .A1(u5_mult_87_n196), .A2(u5_mult_87_n98), 
        .ZN(u5_mult_87_FS_1_n102) );
  OAI21_X1 u5_mult_87_FS_1_U262 ( .B1(u5_mult_87_FS_1_n107), .B2(
        u5_mult_87_FS_1_n101), .A(u5_mult_87_FS_1_n102), .ZN(
        u5_mult_87_FS_1_n299) );
  AND2_X1 u5_mult_87_FS_1_U261 ( .A1(u5_mult_87_n192), .A2(u5_mult_87_n94), 
        .ZN(u5_mult_87_FS_1_n96) );
  AOI21_X1 u5_mult_87_FS_1_U260 ( .B1(u5_mult_87_FS_1_n299), .B2(
        u5_mult_87_FS_1_n13), .A(u5_mult_87_FS_1_n96), .ZN(
        u5_mult_87_FS_1_n298) );
  NAND2_X1 u5_mult_87_FS_1_U259 ( .A1(u5_mult_87_n163), .A2(u5_mult_87_n64), 
        .ZN(u5_mult_87_FS_1_n159) );
  NAND2_X1 u5_mult_87_FS_1_U258 ( .A1(u5_mult_87_n185), .A2(u5_mult_87_n84), 
        .ZN(u5_mult_87_FS_1_n154) );
  OAI21_X1 u5_mult_87_FS_1_U257 ( .B1(u5_mult_87_FS_1_n153), .B2(
        u5_mult_87_FS_1_n159), .A(u5_mult_87_FS_1_n154), .ZN(
        u5_mult_87_FS_1_n297) );
  AND2_X1 u5_mult_87_FS_1_U256 ( .A1(u5_mult_87_n159), .A2(u5_mult_87_n59), 
        .ZN(u5_mult_87_FS_1_n147) );
  AOI21_X1 u5_mult_87_FS_1_U255 ( .B1(u5_mult_87_FS_1_n31), .B2(
        u5_mult_87_FS_1_n297), .A(u5_mult_87_FS_1_n147), .ZN(
        u5_mult_87_FS_1_n296) );
  NAND2_X1 u5_mult_87_FS_1_U254 ( .A1(u5_mult_87_n195), .A2(u5_mult_87_n65), 
        .ZN(u5_mult_87_FS_1_n148) );
  OAI21_X1 u5_mult_87_FS_1_U253 ( .B1(u5_mult_87_FS_1_n296), .B2(
        u5_mult_87_FS_1_n149), .A(u5_mult_87_FS_1_n148), .ZN(
        u5_mult_87_FS_1_n142) );
  NAND2_X1 u5_mult_87_FS_1_U252 ( .A1(u5_mult_87_n187), .A2(u5_mult_87_n90), 
        .ZN(u5_mult_87_FS_1_n141) );
  NAND2_X1 u5_mult_87_FS_1_U251 ( .A1(u5_mult_87_n186), .A2(u5_mult_87_n88), 
        .ZN(u5_mult_87_FS_1_n137) );
  OAI21_X1 u5_mult_87_FS_1_U250 ( .B1(u5_mult_87_FS_1_n136), .B2(
        u5_mult_87_FS_1_n141), .A(u5_mult_87_FS_1_n137), .ZN(
        u5_mult_87_FS_1_n295) );
  AND2_X1 u5_mult_87_FS_1_U249 ( .A1(u5_mult_87_n193), .A2(u5_mult_87_n62), 
        .ZN(u5_mult_87_FS_1_n130) );
  AOI21_X1 u5_mult_87_FS_1_U248 ( .B1(u5_mult_87_FS_1_n26), .B2(
        u5_mult_87_FS_1_n295), .A(u5_mult_87_FS_1_n130), .ZN(
        u5_mult_87_FS_1_n294) );
  NAND2_X1 u5_mult_87_FS_1_U247 ( .A1(u5_mult_87_n203), .A2(u5_mult_87_n89), 
        .ZN(u5_mult_87_FS_1_n131) );
  OAI21_X1 u5_mult_87_FS_1_U246 ( .B1(u5_mult_87_FS_1_n294), .B2(
        u5_mult_87_FS_1_n132), .A(u5_mult_87_FS_1_n131), .ZN(
        u5_mult_87_FS_1_n126) );
  AOI21_X1 u5_mult_87_FS_1_U245 ( .B1(u5_mult_87_FS_1_n125), .B2(
        u5_mult_87_FS_1_n142), .A(u5_mult_87_FS_1_n126), .ZN(
        u5_mult_87_FS_1_n289) );
  NAND2_X1 u5_mult_87_FS_1_U244 ( .A1(u5_mult_87_n202), .A2(u5_mult_87_n87), 
        .ZN(u5_mult_87_FS_1_n122) );
  NAND2_X1 u5_mult_87_FS_1_U243 ( .A1(u5_mult_87_n199), .A2(u5_mult_87_n85), 
        .ZN(u5_mult_87_FS_1_n120) );
  OAI21_X1 u5_mult_87_FS_1_U242 ( .B1(u5_mult_87_FS_1_n118), .B2(
        u5_mult_87_FS_1_n122), .A(u5_mult_87_FS_1_n120), .ZN(
        u5_mult_87_FS_1_n292) );
  NAND2_X1 u5_mult_87_FS_1_U241 ( .A1(u5_mult_87_n200), .A2(u5_mult_87_n86), 
        .ZN(u5_mult_87_FS_1_n115) );
  AOI21_X1 u5_mult_87_FS_1_U240 ( .B1(u5_mult_87_FS_1_n21), .B2(
        u5_mult_87_FS_1_n292), .A(u5_mult_87_FS_1_n20), .ZN(
        u5_mult_87_FS_1_n291) );
  NAND2_X1 u5_mult_87_FS_1_U239 ( .A1(u5_mult_87_n201), .A2(u5_mult_87_n101), 
        .ZN(u5_mult_87_FS_1_n112) );
  OAI21_X1 u5_mult_87_FS_1_U238 ( .B1(u5_mult_87_FS_1_n291), .B2(
        u5_mult_87_FS_1_n111), .A(u5_mult_87_FS_1_n112), .ZN(
        u5_mult_87_FS_1_n290) );
  OAI21_X1 u5_mult_87_FS_1_U237 ( .B1(u5_mult_87_FS_1_n289), .B2(
        u5_mult_87_FS_1_n19), .A(u5_mult_87_FS_1_n17), .ZN(
        u5_mult_87_FS_1_n288) );
  AOI22_X1 u5_mult_87_FS_1_U236 ( .A1(u5_mult_87_FS_1_n11), .A2(
        u5_mult_87_FS_1_n12), .B1(u5_mult_87_FS_1_n287), .B2(
        u5_mult_87_FS_1_n288), .ZN(u5_mult_87_FS_1_n286) );
  NAND3_X1 u5_mult_87_FS_1_U235 ( .A1(u5_mult_87_FS_1_n285), .A2(
        u5_mult_87_FS_1_n97), .A3(u5_mult_87_FS_1_n286), .ZN(
        u5_mult_87_FS_1_n91) );
  OR2_X1 u5_mult_87_FS_1_U234 ( .A1(u5_mult_87_n189), .A2(u5_mult_87_n96), 
        .ZN(u5_mult_87_FS_1_n92) );
  NAND2_X1 u5_mult_87_FS_1_U233 ( .A1(u5_mult_87_FS_1_n91), .A2(
        u5_mult_87_FS_1_n92), .ZN(u5_mult_87_FS_1_n88) );
  OR4_X1 u5_mult_87_FS_1_U232 ( .A1(u5_mult_87_FS_1_n88), .A2(
        u5_mult_87_FS_1_n84), .A3(u5_mult_87_FS_1_n284), .A4(
        u5_mult_87_FS_1_n79), .ZN(u5_mult_87_FS_1_n283) );
  NAND2_X1 u5_mult_87_FS_1_U231 ( .A1(u5_mult_87_n206), .A2(u5_mult_87_n95), 
        .ZN(u5_mult_87_FS_1_n80) );
  OAI211_X1 u5_mult_87_FS_1_U230 ( .C1(u5_mult_87_FS_1_n282), .C2(
        u5_mult_87_FS_1_n79), .A(u5_mult_87_FS_1_n283), .B(u5_mult_87_FS_1_n80), .ZN(u5_mult_87_FS_1_n278) );
  NOR2_X1 u5_mult_87_FS_1_U229 ( .A1(u5_mult_87_n191), .A2(u5_mult_87_n93), 
        .ZN(u5_mult_87_FS_1_n280) );
  AND2_X1 u5_mult_87_FS_1_U228 ( .A1(u5_mult_87_n191), .A2(u5_mult_87_n93), 
        .ZN(u5_mult_87_FS_1_n279) );
  NOR2_X1 u5_mult_87_FS_1_U227 ( .A1(u5_mult_87_FS_1_n280), .A2(
        u5_mult_87_FS_1_n279), .ZN(u5_mult_87_FS_1_n281) );
  XOR2_X1 u5_mult_87_FS_1_U226 ( .A(u5_mult_87_FS_1_n278), .B(
        u5_mult_87_FS_1_n281), .Z(u5_N102) );
  NAND2_X1 u5_mult_87_FS_1_U225 ( .A1(u5_mult_87_n194), .A2(u5_mult_87_n97), 
        .ZN(u5_mult_87_FS_1_n276) );
  NOR2_X1 u5_mult_87_FS_1_U224 ( .A1(u5_mult_87_n194), .A2(u5_mult_87_n97), 
        .ZN(u5_mult_87_FS_1_n274) );
  NAND2_X1 u5_mult_87_FS_1_U223 ( .A1(u5_mult_87_FS_1_n276), .A2(
        u5_mult_87_FS_1_n5), .ZN(u5_mult_87_FS_1_n277) );
  AOI21_X1 u5_mult_87_FS_1_U222 ( .B1(u5_mult_87_FS_1_n6), .B2(
        u5_mult_87_FS_1_n278), .A(u5_mult_87_FS_1_n279), .ZN(
        u5_mult_87_FS_1_n275) );
  XOR2_X1 u5_mult_87_FS_1_U221 ( .A(u5_mult_87_FS_1_n277), .B(
        u5_mult_87_FS_1_n275), .Z(u5_N103) );
  OAI21_X1 u5_mult_87_FS_1_U220 ( .B1(u5_mult_87_FS_1_n274), .B2(
        u5_mult_87_FS_1_n275), .A(u5_mult_87_FS_1_n276), .ZN(
        u5_mult_87_FS_1_n270) );
  NOR2_X1 u5_mult_87_FS_1_U219 ( .A1(u5_mult_87_n190), .A2(u5_mult_87_n92), 
        .ZN(u5_mult_87_FS_1_n272) );
  AND2_X1 u5_mult_87_FS_1_U218 ( .A1(u5_mult_87_n190), .A2(u5_mult_87_n92), 
        .ZN(u5_mult_87_FS_1_n271) );
  NOR2_X1 u5_mult_87_FS_1_U217 ( .A1(u5_mult_87_FS_1_n272), .A2(
        u5_mult_87_FS_1_n271), .ZN(u5_mult_87_FS_1_n273) );
  XOR2_X1 u5_mult_87_FS_1_U216 ( .A(u5_mult_87_FS_1_n270), .B(
        u5_mult_87_FS_1_n273), .Z(u5_N104) );
  AOI21_X1 u5_mult_87_FS_1_U215 ( .B1(u5_mult_87_FS_1_n270), .B2(
        u5_mult_87_FS_1_n4), .A(u5_mult_87_FS_1_n271), .ZN(
        u5_mult_87_FS_1_n269) );
  XOR2_X1 u5_mult_87_FS_1_U214 ( .A(u5_mult_87_FS_1_n3), .B(
        u5_mult_87_FS_1_n269), .Z(u5_N105) );
  NOR2_X1 u5_mult_87_FS_1_U213 ( .A1(u5_mult_87_FS_1_n74), .A2(
        u5_mult_87_FS_1_n265), .ZN(u5_mult_87_FS_1_n266) );
  XOR2_X1 u5_mult_87_FS_1_U212 ( .A(u5_mult_87_FS_1_n76), .B(
        u5_mult_87_FS_1_n266), .Z(u5_N55) );
  NAND2_X1 u5_mult_87_FS_1_U211 ( .A1(u5_mult_87_FS_1_n73), .A2(
        u5_mult_87_FS_1_n263), .ZN(u5_mult_87_FS_1_n264) );
  AOI21_X1 u5_mult_87_FS_1_U210 ( .B1(u5_mult_87_FS_1_n76), .B2(
        u5_mult_87_FS_1_n75), .A(u5_mult_87_FS_1_n74), .ZN(
        u5_mult_87_FS_1_n261) );
  XOR2_X1 u5_mult_87_FS_1_U209 ( .A(u5_mult_87_FS_1_n264), .B(
        u5_mult_87_FS_1_n261), .Z(u5_N56) );
  OAI21_X1 u5_mult_87_FS_1_U208 ( .B1(u5_mult_87_FS_1_n261), .B2(
        u5_mult_87_FS_1_n262), .A(u5_mult_87_FS_1_n263), .ZN(
        u5_mult_87_FS_1_n257) );
  NOR2_X1 u5_mult_87_FS_1_U207 ( .A1(u5_mult_87_FS_1_n71), .A2(
        u5_mult_87_FS_1_n259), .ZN(u5_mult_87_FS_1_n258) );
  XOR2_X1 u5_mult_87_FS_1_U206 ( .A(u5_mult_87_FS_1_n257), .B(
        u5_mult_87_FS_1_n258), .Z(u5_N57) );
  NOR2_X1 u5_mult_87_FS_1_U205 ( .A1(u5_mult_87_FS_1_n255), .A2(
        u5_mult_87_FS_1_n70), .ZN(u5_mult_87_FS_1_n254) );
  XOR2_X1 u5_mult_87_FS_1_U204 ( .A(u5_mult_87_FS_1_n253), .B(
        u5_mult_87_FS_1_n254), .Z(u5_N58) );
  NAND2_X1 u5_mult_87_FS_1_U203 ( .A1(u5_mult_87_FS_1_n68), .A2(
        u5_mult_87_FS_1_n251), .ZN(u5_mult_87_FS_1_n252) );
  AOI21_X1 u5_mult_87_FS_1_U202 ( .B1(u5_mult_87_FS_1_n69), .B2(
        u5_mult_87_FS_1_n253), .A(u5_mult_87_FS_1_n70), .ZN(
        u5_mult_87_FS_1_n249) );
  XOR2_X1 u5_mult_87_FS_1_U201 ( .A(u5_mult_87_FS_1_n252), .B(
        u5_mult_87_FS_1_n249), .Z(u5_N59) );
  OAI21_X1 u5_mult_87_FS_1_U200 ( .B1(u5_mult_87_FS_1_n249), .B2(
        u5_mult_87_FS_1_n250), .A(u5_mult_87_FS_1_n251), .ZN(
        u5_mult_87_FS_1_n244) );
  NOR2_X1 u5_mult_87_FS_1_U199 ( .A1(u5_mult_87_FS_1_n245), .A2(
        u5_mult_87_FS_1_n248), .ZN(u5_mult_87_FS_1_n247) );
  XOR2_X1 u5_mult_87_FS_1_U198 ( .A(u5_mult_87_FS_1_n244), .B(
        u5_mult_87_FS_1_n247), .Z(u5_N60) );
  NAND2_X1 u5_mult_87_FS_1_U197 ( .A1(u5_mult_87_FS_1_n66), .A2(
        u5_mult_87_FS_1_n246), .ZN(u5_mult_87_FS_1_n242) );
  AOI21_X1 u5_mult_87_FS_1_U196 ( .B1(u5_mult_87_FS_1_n67), .B2(
        u5_mult_87_FS_1_n244), .A(u5_mult_87_FS_1_n245), .ZN(
        u5_mult_87_FS_1_n243) );
  XOR2_X1 u5_mult_87_FS_1_U195 ( .A(u5_mult_87_FS_1_n242), .B(
        u5_mult_87_FS_1_n243), .Z(u5_N61) );
  NOR2_X1 u5_mult_87_FS_1_U194 ( .A1(u5_mult_87_FS_1_n240), .A2(
        u5_mult_87_FS_1_n64), .ZN(u5_mult_87_FS_1_n239) );
  XNOR2_X1 u5_mult_87_FS_1_U193 ( .A(u5_mult_87_FS_1_n65), .B(
        u5_mult_87_FS_1_n239), .ZN(u5_N62) );
  NOR2_X1 u5_mult_87_FS_1_U192 ( .A1(u5_mult_87_FS_1_n238), .A2(
        u5_mult_87_FS_1_n64), .ZN(u5_mult_87_FS_1_n233) );
  AND2_X1 u5_mult_87_FS_1_U191 ( .A1(u5_mult_87_FS_1_n235), .A2(
        u5_mult_87_FS_1_n63), .ZN(u5_mult_87_FS_1_n237) );
  XNOR2_X1 u5_mult_87_FS_1_U190 ( .A(u5_mult_87_FS_1_n233), .B(
        u5_mult_87_FS_1_n237), .ZN(u5_N63) );
  NAND2_X1 u5_mult_87_FS_1_U189 ( .A1(u5_mult_87_FS_1_n231), .A2(
        u5_mult_87_FS_1_n236), .ZN(u5_mult_87_FS_1_n232) );
  OAI21_X1 u5_mult_87_FS_1_U188 ( .B1(u5_mult_87_FS_1_n233), .B2(
        u5_mult_87_FS_1_n234), .A(u5_mult_87_FS_1_n235), .ZN(
        u5_mult_87_FS_1_n230) );
  XNOR2_X1 u5_mult_87_FS_1_U187 ( .A(u5_mult_87_FS_1_n232), .B(
        u5_mult_87_FS_1_n230), .ZN(u5_N64) );
  AOI21_X1 u5_mult_87_FS_1_U186 ( .B1(u5_mult_87_FS_1_n230), .B2(
        u5_mult_87_FS_1_n231), .A(u5_mult_87_FS_1_n62), .ZN(
        u5_mult_87_FS_1_n227) );
  AND2_X1 u5_mult_87_FS_1_U185 ( .A1(u5_mult_87_FS_1_n229), .A2(
        u5_mult_87_FS_1_n61), .ZN(u5_mult_87_FS_1_n228) );
  XNOR2_X1 u5_mult_87_FS_1_U184 ( .A(u5_mult_87_FS_1_n227), .B(
        u5_mult_87_FS_1_n228), .ZN(u5_N65) );
  NAND2_X1 u5_mult_87_FS_1_U183 ( .A1(u5_mult_87_FS_1_n224), .A2(
        u5_mult_87_FS_1_n59), .ZN(u5_mult_87_FS_1_n225) );
  XNOR2_X1 u5_mult_87_FS_1_U182 ( .A(u5_mult_87_FS_1_n225), .B(
        u5_mult_87_FS_1_n226), .ZN(u5_N66) );
  OAI21_X1 u5_mult_87_FS_1_U181 ( .B1(u5_mult_87_FS_1_n223), .B2(
        u5_mult_87_FS_1_n60), .A(u5_mult_87_FS_1_n224), .ZN(
        u5_mult_87_FS_1_n219) );
  NOR2_X1 u5_mult_87_FS_1_U180 ( .A1(u5_mult_87_FS_1_n57), .A2(
        u5_mult_87_FS_1_n220), .ZN(u5_mult_87_FS_1_n221) );
  XOR2_X1 u5_mult_87_FS_1_U179 ( .A(u5_mult_87_FS_1_n219), .B(
        u5_mult_87_FS_1_n221), .Z(u5_N67) );
  AOI21_X1 u5_mult_87_FS_1_U178 ( .B1(u5_mult_87_FS_1_n219), .B2(
        u5_mult_87_FS_1_n58), .A(u5_mult_87_FS_1_n57), .ZN(
        u5_mult_87_FS_1_n215) );
  NOR2_X1 u5_mult_87_FS_1_U177 ( .A1(u5_mult_87_FS_1_n55), .A2(
        u5_mult_87_FS_1_n216), .ZN(u5_mult_87_FS_1_n218) );
  XNOR2_X1 u5_mult_87_FS_1_U176 ( .A(u5_mult_87_FS_1_n215), .B(
        u5_mult_87_FS_1_n218), .ZN(u5_N68) );
  OAI21_X1 u5_mult_87_FS_1_U175 ( .B1(u5_mult_87_FS_1_n215), .B2(
        u5_mult_87_FS_1_n216), .A(u5_mult_87_FS_1_n217), .ZN(
        u5_mult_87_FS_1_n211) );
  NOR2_X1 u5_mult_87_FS_1_U174 ( .A1(u5_mult_87_FS_1_n54), .A2(
        u5_mult_87_FS_1_n213), .ZN(u5_mult_87_FS_1_n212) );
  XOR2_X1 u5_mult_87_FS_1_U173 ( .A(u5_mult_87_FS_1_n211), .B(
        u5_mult_87_FS_1_n212), .Z(u5_N69) );
  OR2_X1 u5_mult_87_FS_1_U172 ( .A1(u5_mult_87_FS_1_n209), .A2(
        u5_mult_87_FS_1_n210), .ZN(u5_mult_87_FS_1_n191) );
  NOR2_X1 u5_mult_87_FS_1_U171 ( .A1(u5_mult_87_FS_1_n206), .A2(
        u5_mult_87_FS_1_n52), .ZN(u5_mult_87_FS_1_n207) );
  XOR2_X1 u5_mult_87_FS_1_U170 ( .A(u5_mult_87_FS_1_n191), .B(
        u5_mult_87_FS_1_n207), .Z(u5_N70) );
  NAND2_X1 u5_mult_87_FS_1_U169 ( .A1(u5_mult_87_FS_1_n51), .A2(
        u5_mult_87_FS_1_n204), .ZN(u5_mult_87_FS_1_n205) );
  AOI21_X1 u5_mult_87_FS_1_U168 ( .B1(u5_mult_87_FS_1_n53), .B2(
        u5_mult_87_FS_1_n191), .A(u5_mult_87_FS_1_n52), .ZN(
        u5_mult_87_FS_1_n202) );
  XOR2_X1 u5_mult_87_FS_1_U167 ( .A(u5_mult_87_FS_1_n205), .B(
        u5_mult_87_FS_1_n202), .Z(u5_N71) );
  OAI21_X1 u5_mult_87_FS_1_U166 ( .B1(u5_mult_87_FS_1_n202), .B2(
        u5_mult_87_FS_1_n203), .A(u5_mult_87_FS_1_n204), .ZN(
        u5_mult_87_FS_1_n196) );
  NOR2_X1 u5_mult_87_FS_1_U165 ( .A1(u5_mult_87_FS_1_n197), .A2(
        u5_mult_87_FS_1_n201), .ZN(u5_mult_87_FS_1_n200) );
  XOR2_X1 u5_mult_87_FS_1_U164 ( .A(u5_mult_87_FS_1_n196), .B(
        u5_mult_87_FS_1_n200), .Z(u5_N72) );
  NAND2_X1 u5_mult_87_FS_1_U163 ( .A1(u5_mult_87_FS_1_n49), .A2(
        u5_mult_87_FS_1_n198), .ZN(u5_mult_87_FS_1_n194) );
  AOI21_X1 u5_mult_87_FS_1_U162 ( .B1(u5_mult_87_FS_1_n50), .B2(
        u5_mult_87_FS_1_n196), .A(u5_mult_87_FS_1_n197), .ZN(
        u5_mult_87_FS_1_n195) );
  XOR2_X1 u5_mult_87_FS_1_U161 ( .A(u5_mult_87_FS_1_n194), .B(
        u5_mult_87_FS_1_n195), .Z(u5_N73) );
  NAND2_X1 u5_mult_87_FS_1_U160 ( .A1(u5_mult_87_FS_1_n189), .A2(
        u5_mult_87_FS_1_n48), .ZN(u5_mult_87_FS_1_n190) );
  AOI21_X1 u5_mult_87_FS_1_U159 ( .B1(u5_mult_87_FS_1_n191), .B2(
        u5_mult_87_FS_1_n192), .A(u5_mult_87_FS_1_n193), .ZN(
        u5_mult_87_FS_1_n175) );
  XOR2_X1 u5_mult_87_FS_1_U158 ( .A(u5_mult_87_FS_1_n190), .B(
        u5_mult_87_FS_1_n175), .Z(u5_N74) );
  OAI21_X1 u5_mult_87_FS_1_U157 ( .B1(u5_mult_87_FS_1_n188), .B2(
        u5_mult_87_FS_1_n175), .A(u5_mult_87_FS_1_n189), .ZN(
        u5_mult_87_FS_1_n184) );
  NOR2_X1 u5_mult_87_FS_1_U156 ( .A1(u5_mult_87_FS_1_n46), .A2(
        u5_mult_87_FS_1_n185), .ZN(u5_mult_87_FS_1_n186) );
  XOR2_X1 u5_mult_87_FS_1_U155 ( .A(u5_mult_87_FS_1_n184), .B(
        u5_mult_87_FS_1_n186), .Z(u5_N75) );
  AOI21_X1 u5_mult_87_FS_1_U154 ( .B1(u5_mult_87_FS_1_n184), .B2(
        u5_mult_87_FS_1_n47), .A(u5_mult_87_FS_1_n46), .ZN(
        u5_mult_87_FS_1_n180) );
  NOR2_X1 u5_mult_87_FS_1_U153 ( .A1(u5_mult_87_FS_1_n44), .A2(
        u5_mult_87_FS_1_n181), .ZN(u5_mult_87_FS_1_n183) );
  XNOR2_X1 u5_mult_87_FS_1_U152 ( .A(u5_mult_87_FS_1_n180), .B(
        u5_mult_87_FS_1_n183), .ZN(u5_N76) );
  OAI21_X1 u5_mult_87_FS_1_U151 ( .B1(u5_mult_87_FS_1_n180), .B2(
        u5_mult_87_FS_1_n181), .A(u5_mult_87_FS_1_n182), .ZN(
        u5_mult_87_FS_1_n176) );
  NOR2_X1 u5_mult_87_FS_1_U150 ( .A1(u5_mult_87_FS_1_n42), .A2(
        u5_mult_87_FS_1_n178), .ZN(u5_mult_87_FS_1_n177) );
  XOR2_X1 u5_mult_87_FS_1_U149 ( .A(u5_mult_87_FS_1_n176), .B(
        u5_mult_87_FS_1_n177), .Z(u5_N77) );
  OAI21_X1 u5_mult_87_FS_1_U148 ( .B1(u5_mult_87_FS_1_n175), .B2(
        u5_mult_87_FS_1_n43), .A(u5_mult_87_FS_1_n41), .ZN(
        u5_mult_87_FS_1_n171) );
  NOR2_X1 u5_mult_87_FS_1_U147 ( .A1(u5_mult_87_FS_1_n172), .A2(
        u5_mult_87_FS_1_n39), .ZN(u5_mult_87_FS_1_n173) );
  XOR2_X1 u5_mult_87_FS_1_U146 ( .A(u5_mult_87_FS_1_n171), .B(
        u5_mult_87_FS_1_n173), .Z(u5_N78) );
  NAND2_X1 u5_mult_87_FS_1_U145 ( .A1(u5_mult_87_FS_1_n38), .A2(
        u5_mult_87_FS_1_n169), .ZN(u5_mult_87_FS_1_n170) );
  AOI21_X1 u5_mult_87_FS_1_U144 ( .B1(u5_mult_87_FS_1_n40), .B2(
        u5_mult_87_FS_1_n171), .A(u5_mult_87_FS_1_n39), .ZN(
        u5_mult_87_FS_1_n167) );
  XOR2_X1 u5_mult_87_FS_1_U143 ( .A(u5_mult_87_FS_1_n170), .B(
        u5_mult_87_FS_1_n167), .Z(u5_N79) );
  OAI21_X1 u5_mult_87_FS_1_U142 ( .B1(u5_mult_87_FS_1_n167), .B2(
        u5_mult_87_FS_1_n168), .A(u5_mult_87_FS_1_n169), .ZN(
        u5_mult_87_FS_1_n162) );
  NOR2_X1 u5_mult_87_FS_1_U141 ( .A1(u5_mult_87_FS_1_n163), .A2(
        u5_mult_87_FS_1_n166), .ZN(u5_mult_87_FS_1_n165) );
  XOR2_X1 u5_mult_87_FS_1_U140 ( .A(u5_mult_87_FS_1_n162), .B(
        u5_mult_87_FS_1_n165), .Z(u5_N80) );
  NAND2_X1 u5_mult_87_FS_1_U139 ( .A1(u5_mult_87_FS_1_n35), .A2(
        u5_mult_87_FS_1_n164), .ZN(u5_mult_87_FS_1_n160) );
  AOI21_X1 u5_mult_87_FS_1_U138 ( .B1(u5_mult_87_FS_1_n37), .B2(
        u5_mult_87_FS_1_n162), .A(u5_mult_87_FS_1_n163), .ZN(
        u5_mult_87_FS_1_n161) );
  XOR2_X1 u5_mult_87_FS_1_U137 ( .A(u5_mult_87_FS_1_n160), .B(
        u5_mult_87_FS_1_n161), .Z(u5_N81) );
  NOR2_X1 u5_mult_87_FS_1_U136 ( .A1(u5_mult_87_FS_1_n157), .A2(
        u5_mult_87_FS_1_n33), .ZN(u5_mult_87_FS_1_n158) );
  XOR2_X1 u5_mult_87_FS_1_U135 ( .A(u5_mult_87_FS_1_n156), .B(
        u5_mult_87_FS_1_n158), .Z(u5_N82) );
  NAND2_X1 u5_mult_87_FS_1_U134 ( .A1(u5_mult_87_FS_1_n32), .A2(
        u5_mult_87_FS_1_n154), .ZN(u5_mult_87_FS_1_n155) );
  AOI21_X1 u5_mult_87_FS_1_U133 ( .B1(u5_mult_87_FS_1_n34), .B2(
        u5_mult_87_FS_1_n156), .A(u5_mult_87_FS_1_n33), .ZN(
        u5_mult_87_FS_1_n152) );
  XOR2_X1 u5_mult_87_FS_1_U132 ( .A(u5_mult_87_FS_1_n155), .B(
        u5_mult_87_FS_1_n152), .Z(u5_N83) );
  OAI21_X1 u5_mult_87_FS_1_U131 ( .B1(u5_mult_87_FS_1_n152), .B2(
        u5_mult_87_FS_1_n153), .A(u5_mult_87_FS_1_n154), .ZN(
        u5_mult_87_FS_1_n146) );
  NOR2_X1 u5_mult_87_FS_1_U130 ( .A1(u5_mult_87_FS_1_n147), .A2(
        u5_mult_87_FS_1_n151), .ZN(u5_mult_87_FS_1_n150) );
  XOR2_X1 u5_mult_87_FS_1_U129 ( .A(u5_mult_87_FS_1_n146), .B(
        u5_mult_87_FS_1_n150), .Z(u5_N84) );
  NAND2_X1 u5_mult_87_FS_1_U128 ( .A1(u5_mult_87_FS_1_n30), .A2(
        u5_mult_87_FS_1_n148), .ZN(u5_mult_87_FS_1_n144) );
  AOI21_X1 u5_mult_87_FS_1_U127 ( .B1(u5_mult_87_FS_1_n31), .B2(
        u5_mult_87_FS_1_n146), .A(u5_mult_87_FS_1_n147), .ZN(
        u5_mult_87_FS_1_n145) );
  XOR2_X1 u5_mult_87_FS_1_U126 ( .A(u5_mult_87_FS_1_n144), .B(
        u5_mult_87_FS_1_n145), .Z(u5_N85) );
  OR2_X1 u5_mult_87_FS_1_U125 ( .A1(u5_mult_87_FS_1_n142), .A2(
        u5_mult_87_FS_1_n143), .ZN(u5_mult_87_FS_1_n124) );
  NOR2_X1 u5_mult_87_FS_1_U124 ( .A1(u5_mult_87_FS_1_n139), .A2(
        u5_mult_87_FS_1_n28), .ZN(u5_mult_87_FS_1_n140) );
  XOR2_X1 u5_mult_87_FS_1_U123 ( .A(u5_mult_87_FS_1_n124), .B(
        u5_mult_87_FS_1_n140), .Z(u5_N86) );
  NAND2_X1 u5_mult_87_FS_1_U122 ( .A1(u5_mult_87_FS_1_n27), .A2(
        u5_mult_87_FS_1_n137), .ZN(u5_mult_87_FS_1_n138) );
  AOI21_X1 u5_mult_87_FS_1_U121 ( .B1(u5_mult_87_FS_1_n29), .B2(
        u5_mult_87_FS_1_n124), .A(u5_mult_87_FS_1_n28), .ZN(
        u5_mult_87_FS_1_n135) );
  XOR2_X1 u5_mult_87_FS_1_U120 ( .A(u5_mult_87_FS_1_n138), .B(
        u5_mult_87_FS_1_n135), .Z(u5_N87) );
  OAI21_X1 u5_mult_87_FS_1_U119 ( .B1(u5_mult_87_FS_1_n135), .B2(
        u5_mult_87_FS_1_n136), .A(u5_mult_87_FS_1_n137), .ZN(
        u5_mult_87_FS_1_n129) );
  NOR2_X1 u5_mult_87_FS_1_U118 ( .A1(u5_mult_87_FS_1_n130), .A2(
        u5_mult_87_FS_1_n134), .ZN(u5_mult_87_FS_1_n133) );
  XOR2_X1 u5_mult_87_FS_1_U117 ( .A(u5_mult_87_FS_1_n129), .B(
        u5_mult_87_FS_1_n133), .Z(u5_N88) );
  NAND2_X1 u5_mult_87_FS_1_U116 ( .A1(u5_mult_87_FS_1_n25), .A2(
        u5_mult_87_FS_1_n131), .ZN(u5_mult_87_FS_1_n127) );
  AOI21_X1 u5_mult_87_FS_1_U115 ( .B1(u5_mult_87_FS_1_n26), .B2(
        u5_mult_87_FS_1_n129), .A(u5_mult_87_FS_1_n130), .ZN(
        u5_mult_87_FS_1_n128) );
  XOR2_X1 u5_mult_87_FS_1_U114 ( .A(u5_mult_87_FS_1_n127), .B(
        u5_mult_87_FS_1_n128), .Z(u5_N89) );
  NAND2_X1 u5_mult_87_FS_1_U113 ( .A1(u5_mult_87_FS_1_n122), .A2(
        u5_mult_87_FS_1_n24), .ZN(u5_mult_87_FS_1_n123) );
  AOI21_X1 u5_mult_87_FS_1_U112 ( .B1(u5_mult_87_FS_1_n124), .B2(
        u5_mult_87_FS_1_n125), .A(u5_mult_87_FS_1_n126), .ZN(
        u5_mult_87_FS_1_n108) );
  XOR2_X1 u5_mult_87_FS_1_U111 ( .A(u5_mult_87_FS_1_n123), .B(
        u5_mult_87_FS_1_n108), .Z(u5_N90) );
  OAI21_X1 u5_mult_87_FS_1_U110 ( .B1(u5_mult_87_FS_1_n121), .B2(
        u5_mult_87_FS_1_n108), .A(u5_mult_87_FS_1_n122), .ZN(
        u5_mult_87_FS_1_n117) );
  NOR2_X1 u5_mult_87_FS_1_U109 ( .A1(u5_mult_87_FS_1_n22), .A2(
        u5_mult_87_FS_1_n118), .ZN(u5_mult_87_FS_1_n119) );
  XOR2_X1 u5_mult_87_FS_1_U108 ( .A(u5_mult_87_FS_1_n117), .B(
        u5_mult_87_FS_1_n119), .Z(u5_N91) );
  NAND2_X1 u5_mult_87_FS_1_U107 ( .A1(u5_mult_87_FS_1_n21), .A2(
        u5_mult_87_FS_1_n115), .ZN(u5_mult_87_FS_1_n116) );
  AOI21_X1 u5_mult_87_FS_1_U106 ( .B1(u5_mult_87_FS_1_n117), .B2(
        u5_mult_87_FS_1_n23), .A(u5_mult_87_FS_1_n22), .ZN(
        u5_mult_87_FS_1_n113) );
  XOR2_X1 u5_mult_87_FS_1_U105 ( .A(u5_mult_87_FS_1_n116), .B(
        u5_mult_87_FS_1_n113), .Z(u5_N92) );
  OAI21_X1 u5_mult_87_FS_1_U104 ( .B1(u5_mult_87_FS_1_n113), .B2(
        u5_mult_87_FS_1_n114), .A(u5_mult_87_FS_1_n115), .ZN(
        u5_mult_87_FS_1_n109) );
  NOR2_X1 u5_mult_87_FS_1_U103 ( .A1(u5_mult_87_FS_1_n18), .A2(
        u5_mult_87_FS_1_n111), .ZN(u5_mult_87_FS_1_n110) );
  XOR2_X1 u5_mult_87_FS_1_U102 ( .A(u5_mult_87_FS_1_n109), .B(
        u5_mult_87_FS_1_n110), .Z(u5_N93) );
  OAI21_X1 u5_mult_87_FS_1_U101 ( .B1(u5_mult_87_FS_1_n108), .B2(
        u5_mult_87_FS_1_n19), .A(u5_mult_87_FS_1_n17), .ZN(
        u5_mult_87_FS_1_n104) );
  NOR2_X1 u5_mult_87_FS_1_U100 ( .A1(u5_mult_87_FS_1_n105), .A2(
        u5_mult_87_FS_1_n15), .ZN(u5_mult_87_FS_1_n106) );
  XOR2_X1 u5_mult_87_FS_1_U99 ( .A(u5_mult_87_FS_1_n104), .B(
        u5_mult_87_FS_1_n106), .Z(u5_N94) );
  NAND2_X1 u5_mult_87_FS_1_U98 ( .A1(u5_mult_87_FS_1_n14), .A2(
        u5_mult_87_FS_1_n102), .ZN(u5_mult_87_FS_1_n103) );
  AOI21_X1 u5_mult_87_FS_1_U97 ( .B1(u5_mult_87_FS_1_n16), .B2(
        u5_mult_87_FS_1_n104), .A(u5_mult_87_FS_1_n15), .ZN(
        u5_mult_87_FS_1_n100) );
  XOR2_X1 u5_mult_87_FS_1_U96 ( .A(u5_mult_87_FS_1_n103), .B(
        u5_mult_87_FS_1_n100), .Z(u5_N95) );
  OAI21_X1 u5_mult_87_FS_1_U95 ( .B1(u5_mult_87_FS_1_n100), .B2(
        u5_mult_87_FS_1_n101), .A(u5_mult_87_FS_1_n102), .ZN(
        u5_mult_87_FS_1_n95) );
  NOR2_X1 u5_mult_87_FS_1_U94 ( .A1(u5_mult_87_FS_1_n96), .A2(
        u5_mult_87_FS_1_n99), .ZN(u5_mult_87_FS_1_n98) );
  XOR2_X1 u5_mult_87_FS_1_U93 ( .A(u5_mult_87_FS_1_n95), .B(
        u5_mult_87_FS_1_n98), .Z(u5_N96) );
  NAND2_X1 u5_mult_87_FS_1_U92 ( .A1(u5_mult_87_FS_1_n11), .A2(
        u5_mult_87_FS_1_n97), .ZN(u5_mult_87_FS_1_n93) );
  AOI21_X1 u5_mult_87_FS_1_U91 ( .B1(u5_mult_87_FS_1_n13), .B2(
        u5_mult_87_FS_1_n95), .A(u5_mult_87_FS_1_n96), .ZN(u5_mult_87_FS_1_n94) );
  XOR2_X1 u5_mult_87_FS_1_U90 ( .A(u5_mult_87_FS_1_n93), .B(
        u5_mult_87_FS_1_n94), .Z(u5_N97) );
  NAND2_X1 u5_mult_87_FS_1_U89 ( .A1(u5_mult_87_FS_1_n89), .A2(
        u5_mult_87_FS_1_n92), .ZN(u5_mult_87_FS_1_n90) );
  XNOR2_X1 u5_mult_87_FS_1_U88 ( .A(u5_mult_87_FS_1_n90), .B(
        u5_mult_87_FS_1_n91), .ZN(u5_N98) );
  NAND2_X1 u5_mult_87_FS_1_U87 ( .A1(u5_mult_87_FS_1_n10), .A2(
        u5_mult_87_FS_1_n85), .ZN(u5_mult_87_FS_1_n87) );
  AND2_X1 u5_mult_87_FS_1_U86 ( .A1(u5_mult_87_FS_1_n88), .A2(
        u5_mult_87_FS_1_n89), .ZN(u5_mult_87_FS_1_n83) );
  XOR2_X1 u5_mult_87_FS_1_U85 ( .A(u5_mult_87_FS_1_n87), .B(
        u5_mult_87_FS_1_n83), .Z(u5_N99) );
  NAND2_X1 u5_mult_87_FS_1_U84 ( .A1(u5_mult_87_FS_1_n9), .A2(
        u5_mult_87_FS_1_n86), .ZN(u5_mult_87_FS_1_n82) );
  OAI21_X1 u5_mult_87_FS_1_U83 ( .B1(u5_mult_87_FS_1_n83), .B2(
        u5_mult_87_FS_1_n84), .A(u5_mult_87_FS_1_n85), .ZN(u5_mult_87_FS_1_n81) );
  XNOR2_X1 u5_mult_87_FS_1_U82 ( .A(u5_mult_87_FS_1_n82), .B(
        u5_mult_87_FS_1_n81), .ZN(u5_N100) );
  AOI21_X1 u5_mult_87_FS_1_U81 ( .B1(u5_mult_87_FS_1_n81), .B2(
        u5_mult_87_FS_1_n9), .A(u5_mult_87_FS_1_n8), .ZN(u5_mult_87_FS_1_n77)
         );
  NOR2_X1 u5_mult_87_FS_1_U80 ( .A1(u5_mult_87_FS_1_n79), .A2(
        u5_mult_87_FS_1_n7), .ZN(u5_mult_87_FS_1_n78) );
  XNOR2_X1 u5_mult_87_FS_1_U79 ( .A(u5_mult_87_FS_1_n77), .B(
        u5_mult_87_FS_1_n78), .ZN(u5_N101) );
  INV_X4 u5_mult_87_FS_1_U78 ( .A(u5_mult_87_FS_1_n268), .ZN(
        u5_mult_87_FS_1_n76) );
  INV_X4 u5_mult_87_FS_1_U77 ( .A(u5_mult_87_FS_1_n265), .ZN(
        u5_mult_87_FS_1_n75) );
  INV_X4 u5_mult_87_FS_1_U76 ( .A(u5_mult_87_FS_1_n267), .ZN(
        u5_mult_87_FS_1_n74) );
  INV_X4 u5_mult_87_FS_1_U75 ( .A(u5_mult_87_FS_1_n262), .ZN(
        u5_mult_87_FS_1_n73) );
  INV_X4 u5_mult_87_FS_1_U74 ( .A(u5_mult_87_FS_1_n263), .ZN(
        u5_mult_87_FS_1_n72) );
  INV_X4 u5_mult_87_FS_1_U73 ( .A(u5_mult_87_FS_1_n260), .ZN(
        u5_mult_87_FS_1_n71) );
  INV_X4 u5_mult_87_FS_1_U72 ( .A(u5_mult_87_FS_1_n256), .ZN(
        u5_mult_87_FS_1_n70) );
  INV_X4 u5_mult_87_FS_1_U71 ( .A(u5_mult_87_FS_1_n255), .ZN(
        u5_mult_87_FS_1_n69) );
  INV_X4 u5_mult_87_FS_1_U70 ( .A(u5_mult_87_FS_1_n250), .ZN(
        u5_mult_87_FS_1_n68) );
  INV_X4 u5_mult_87_FS_1_U69 ( .A(u5_mult_87_FS_1_n248), .ZN(
        u5_mult_87_FS_1_n67) );
  INV_X4 u5_mult_87_FS_1_U68 ( .A(u5_mult_87_FS_1_n324), .ZN(
        u5_mult_87_FS_1_n66) );
  INV_X4 u5_mult_87_FS_1_U67 ( .A(u5_mult_87_FS_1_n322), .ZN(
        u5_mult_87_FS_1_n65) );
  INV_X4 u5_mult_87_FS_1_U66 ( .A(u5_mult_87_FS_1_n241), .ZN(
        u5_mult_87_FS_1_n64) );
  INV_X4 u5_mult_87_FS_1_U65 ( .A(u5_mult_87_FS_1_n234), .ZN(
        u5_mult_87_FS_1_n63) );
  INV_X4 u5_mult_87_FS_1_U64 ( .A(u5_mult_87_FS_1_n236), .ZN(
        u5_mult_87_FS_1_n62) );
  INV_X4 u5_mult_87_FS_1_U63 ( .A(u5_mult_87_FS_1_n320), .ZN(
        u5_mult_87_FS_1_n61) );
  INV_X4 u5_mult_87_FS_1_U62 ( .A(u5_mult_87_FS_1_n226), .ZN(
        u5_mult_87_FS_1_n60) );
  INV_X4 u5_mult_87_FS_1_U61 ( .A(u5_mult_87_FS_1_n223), .ZN(
        u5_mult_87_FS_1_n59) );
  INV_X4 u5_mult_87_FS_1_U60 ( .A(u5_mult_87_FS_1_n220), .ZN(
        u5_mult_87_FS_1_n58) );
  INV_X4 u5_mult_87_FS_1_U59 ( .A(u5_mult_87_FS_1_n222), .ZN(
        u5_mult_87_FS_1_n57) );
  INV_X4 u5_mult_87_FS_1_U58 ( .A(u5_mult_87_FS_1_n216), .ZN(
        u5_mult_87_FS_1_n56) );
  INV_X4 u5_mult_87_FS_1_U57 ( .A(u5_mult_87_FS_1_n217), .ZN(
        u5_mult_87_FS_1_n55) );
  INV_X4 u5_mult_87_FS_1_U56 ( .A(u5_mult_87_FS_1_n214), .ZN(
        u5_mult_87_FS_1_n54) );
  INV_X4 u5_mult_87_FS_1_U55 ( .A(u5_mult_87_FS_1_n206), .ZN(
        u5_mult_87_FS_1_n53) );
  INV_X4 u5_mult_87_FS_1_U54 ( .A(u5_mult_87_FS_1_n208), .ZN(
        u5_mult_87_FS_1_n52) );
  INV_X4 u5_mult_87_FS_1_U53 ( .A(u5_mult_87_FS_1_n203), .ZN(
        u5_mult_87_FS_1_n51) );
  INV_X4 u5_mult_87_FS_1_U52 ( .A(u5_mult_87_FS_1_n201), .ZN(
        u5_mult_87_FS_1_n50) );
  INV_X4 u5_mult_87_FS_1_U51 ( .A(u5_mult_87_FS_1_n199), .ZN(
        u5_mult_87_FS_1_n49) );
  INV_X4 u5_mult_87_FS_1_U50 ( .A(u5_mult_87_FS_1_n188), .ZN(
        u5_mult_87_FS_1_n48) );
  INV_X4 u5_mult_87_FS_1_U49 ( .A(u5_mult_87_FS_1_n185), .ZN(
        u5_mult_87_FS_1_n47) );
  INV_X4 u5_mult_87_FS_1_U48 ( .A(u5_mult_87_FS_1_n187), .ZN(
        u5_mult_87_FS_1_n46) );
  INV_X4 u5_mult_87_FS_1_U47 ( .A(u5_mult_87_FS_1_n181), .ZN(
        u5_mult_87_FS_1_n45) );
  INV_X4 u5_mult_87_FS_1_U46 ( .A(u5_mult_87_FS_1_n182), .ZN(
        u5_mult_87_FS_1_n44) );
  INV_X4 u5_mult_87_FS_1_U45 ( .A(u5_mult_87_FS_1_n310), .ZN(
        u5_mult_87_FS_1_n43) );
  INV_X4 u5_mult_87_FS_1_U44 ( .A(u5_mult_87_FS_1_n179), .ZN(
        u5_mult_87_FS_1_n42) );
  INV_X4 u5_mult_87_FS_1_U43 ( .A(u5_mult_87_FS_1_n307), .ZN(
        u5_mult_87_FS_1_n41) );
  INV_X4 u5_mult_87_FS_1_U42 ( .A(u5_mult_87_FS_1_n172), .ZN(
        u5_mult_87_FS_1_n40) );
  INV_X4 u5_mult_87_FS_1_U41 ( .A(u5_mult_87_FS_1_n174), .ZN(
        u5_mult_87_FS_1_n39) );
  INV_X4 u5_mult_87_FS_1_U40 ( .A(u5_mult_87_FS_1_n168), .ZN(
        u5_mult_87_FS_1_n38) );
  INV_X4 u5_mult_87_FS_1_U39 ( .A(u5_mult_87_FS_1_n166), .ZN(
        u5_mult_87_FS_1_n37) );
  INV_X4 u5_mult_87_FS_1_U38 ( .A(u5_mult_87_FS_1_n315), .ZN(
        u5_mult_87_FS_1_n36) );
  INV_X4 u5_mult_87_FS_1_U37 ( .A(u5_mult_87_FS_1_n317), .ZN(
        u5_mult_87_FS_1_n35) );
  INV_X4 u5_mult_87_FS_1_U36 ( .A(u5_mult_87_FS_1_n157), .ZN(
        u5_mult_87_FS_1_n34) );
  INV_X4 u5_mult_87_FS_1_U35 ( .A(u5_mult_87_FS_1_n159), .ZN(
        u5_mult_87_FS_1_n33) );
  INV_X4 u5_mult_87_FS_1_U34 ( .A(u5_mult_87_FS_1_n153), .ZN(
        u5_mult_87_FS_1_n32) );
  INV_X4 u5_mult_87_FS_1_U33 ( .A(u5_mult_87_FS_1_n151), .ZN(
        u5_mult_87_FS_1_n31) );
  INV_X4 u5_mult_87_FS_1_U32 ( .A(u5_mult_87_FS_1_n149), .ZN(
        u5_mult_87_FS_1_n30) );
  INV_X4 u5_mult_87_FS_1_U31 ( .A(u5_mult_87_FS_1_n139), .ZN(
        u5_mult_87_FS_1_n29) );
  INV_X4 u5_mult_87_FS_1_U30 ( .A(u5_mult_87_FS_1_n141), .ZN(
        u5_mult_87_FS_1_n28) );
  INV_X4 u5_mult_87_FS_1_U29 ( .A(u5_mult_87_FS_1_n136), .ZN(
        u5_mult_87_FS_1_n27) );
  INV_X4 u5_mult_87_FS_1_U28 ( .A(u5_mult_87_FS_1_n134), .ZN(
        u5_mult_87_FS_1_n26) );
  INV_X4 u5_mult_87_FS_1_U27 ( .A(u5_mult_87_FS_1_n132), .ZN(
        u5_mult_87_FS_1_n25) );
  INV_X4 u5_mult_87_FS_1_U26 ( .A(u5_mult_87_FS_1_n121), .ZN(
        u5_mult_87_FS_1_n24) );
  INV_X4 u5_mult_87_FS_1_U25 ( .A(u5_mult_87_FS_1_n118), .ZN(
        u5_mult_87_FS_1_n23) );
  INV_X4 u5_mult_87_FS_1_U24 ( .A(u5_mult_87_FS_1_n120), .ZN(
        u5_mult_87_FS_1_n22) );
  INV_X4 u5_mult_87_FS_1_U23 ( .A(u5_mult_87_FS_1_n114), .ZN(
        u5_mult_87_FS_1_n21) );
  INV_X4 u5_mult_87_FS_1_U22 ( .A(u5_mult_87_FS_1_n115), .ZN(
        u5_mult_87_FS_1_n20) );
  INV_X4 u5_mult_87_FS_1_U21 ( .A(u5_mult_87_FS_1_n293), .ZN(
        u5_mult_87_FS_1_n19) );
  INV_X4 u5_mult_87_FS_1_U20 ( .A(u5_mult_87_FS_1_n112), .ZN(
        u5_mult_87_FS_1_n18) );
  INV_X4 u5_mult_87_FS_1_U19 ( .A(u5_mult_87_FS_1_n290), .ZN(
        u5_mult_87_FS_1_n17) );
  INV_X4 u5_mult_87_FS_1_U18 ( .A(u5_mult_87_FS_1_n105), .ZN(
        u5_mult_87_FS_1_n16) );
  INV_X4 u5_mult_87_FS_1_U17 ( .A(u5_mult_87_FS_1_n107), .ZN(
        u5_mult_87_FS_1_n15) );
  INV_X4 u5_mult_87_FS_1_U16 ( .A(u5_mult_87_FS_1_n101), .ZN(
        u5_mult_87_FS_1_n14) );
  INV_X4 u5_mult_87_FS_1_U15 ( .A(u5_mult_87_FS_1_n99), .ZN(
        u5_mult_87_FS_1_n13) );
  INV_X4 u5_mult_87_FS_1_U14 ( .A(u5_mult_87_FS_1_n298), .ZN(
        u5_mult_87_FS_1_n12) );
  INV_X4 u5_mult_87_FS_1_U13 ( .A(u5_mult_87_FS_1_n300), .ZN(
        u5_mult_87_FS_1_n11) );
  INV_X4 u5_mult_87_FS_1_U12 ( .A(u5_mult_87_FS_1_n84), .ZN(
        u5_mult_87_FS_1_n10) );
  INV_X4 u5_mult_87_FS_1_U11 ( .A(u5_mult_87_FS_1_n284), .ZN(
        u5_mult_87_FS_1_n9) );
  INV_X4 u5_mult_87_FS_1_U10 ( .A(u5_mult_87_FS_1_n86), .ZN(u5_mult_87_FS_1_n8) );
  INV_X4 u5_mult_87_FS_1_U9 ( .A(u5_mult_87_FS_1_n80), .ZN(u5_mult_87_FS_1_n7)
         );
  INV_X4 u5_mult_87_FS_1_U8 ( .A(u5_mult_87_FS_1_n280), .ZN(u5_mult_87_FS_1_n6) );
  INV_X4 u5_mult_87_FS_1_U7 ( .A(u5_mult_87_FS_1_n274), .ZN(u5_mult_87_FS_1_n5) );
  INV_X4 u5_mult_87_FS_1_U6 ( .A(u5_mult_87_FS_1_n272), .ZN(u5_mult_87_FS_1_n4) );
  INV_X4 u5_mult_87_FS_1_U5 ( .A(u5_mult_87_n208), .ZN(u5_mult_87_FS_1_n3) );
  OR2_X4 u5_mult_87_FS_1_U4 ( .A1(u5_mult_87_n105), .A2(u5_mult_87_n5), .ZN(
        u5_mult_87_FS_1_n2) );
  AND2_X4 u5_mult_87_FS_1_U3 ( .A1(u5_mult_87_FS_1_n268), .A2(
        u5_mult_87_FS_1_n2), .ZN(u5_N54) );
  OAI21_X2 u5_mult_87_FS_1_U2 ( .B1(u5_mult_87_FS_1_n327), .B2(
        u5_mult_87_FS_1_n259), .A(u5_mult_87_FS_1_n260), .ZN(
        u5_mult_87_FS_1_n253) );
endmodule

