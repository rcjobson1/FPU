`define BIT_SIZE 15 
`define EXP_SIZE 4
`define MANT_SIZE 9 
`define BIAS 15
`define EXP_SHIFT 3
