`timescale 1ns / 100ps
    module test;

    ////////////////////////////////////////////////////////////////////////
    // Parameters
    // 64 bit = 0
    // 32 bit = 1
    // 16 bit = 2
    parameter
      FPU_TYPE = 2,
      BIT_SIZE = 16 * 2**(2 - FPU_TYPE) - 1,
      EXP_SIZE = 11 - (3*FPU_TYPE) - 1,
      MANT_SIZE = BIT_SIZE  - EXP_SIZE - 2,
      BIAS = 2**(10-(3*FPU_TYPE)) - 1;

    ////////////////////////////////////////////////////////////////////////

    initial begin
      $dumpfile("CPU_16.vcd");
      $dumpvars(0,test);
    end
    event		error_event;
    reg clk = 0;
    always #10 clk = !clk;
    reg [1:0] fpu_rmode = 0; //round to nearest even
    reg [15:0] opa, opb;
    reg [2:0] fpu_op;
    wire [15:0] out;
    wire snan, qnan, inf, ine, overflow, underflow, div_by_zero, zero;

    fpu #(.BIT_SIZE(BIT_SIZE), .EXP_SIZE(EXP_SIZE), .MANT_SIZE(MANT_SIZE), .BIAS(BIAS) ) u0(clk, fpu_rmode, fpu_op, opa, opb, out, snan, qnan, inf, ine, overflow, underflow, div_by_zero, zero);

    always #1800 $finish;
initial begin
#40 fpu_op <= 1;
opa <= 16'hf0cd;
opb <= 16'h6119;

#40 fpu_op <= 2;
opa <= 16'h75c8;
opb <= 16'h9a15;

#40 fpu_op <= 0;
opa <= 16'hc401;
opb <= 16'h38af;

#40 fpu_op <= 2;
opa <= 16'hdbd8;
opb <= 16'h96a9;

#40 fpu_op <= 0;
opa <= 16'hd686;
opb <= 16'h217;

#40 fpu_op <= 0;
opa <= 16'h576;
opb <= 16'h4cbe;

#40 fpu_op <= 2;
opa <= 16'hff54;
opb <= 16'hcc1e;

#40 fpu_op <= 1;
opa <= 16'hd4d1;
opb <= 16'h7efb;

#40 fpu_op <= 0;
opa <= 16'hddc2;
opb <= 16'hce3d;

#40 fpu_op <= 0;
opa <= 16'h1dbb;
opb <= 16'hd63d;

end
endmodule