
module fpu_DW01_ash_1 ( A, DATA_TC, SH, SH_TC, B );
  input [29:0] A;
  input [4:0] SH;
  output [29:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][27] , \ML_int[1][24] , \ML_int[1][22] , \ML_int[1][21] ,
         \ML_int[1][20] , \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] ,
         \ML_int[1][16] , \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] ,
         \ML_int[1][12] , \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] ,
         \ML_int[1][8] , \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] ,
         \ML_int[1][4] , \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] ,
         \ML_int[1][0] , \ML_int[2][27] , \ML_int[2][26] , \ML_int[2][25] ,
         \ML_int[2][24] , \ML_int[2][23] , \ML_int[2][22] , \ML_int[2][21] ,
         \ML_int[2][20] , \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] ,
         \ML_int[2][16] , \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] ,
         \ML_int[2][12] , \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] ,
         \ML_int[2][8] , \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] ,
         \ML_int[2][4] , \ML_int[2][3] , \ML_int[2][2] , \ML_int[3][27] ,
         \ML_int[3][26] , \ML_int[3][25] , \ML_int[3][24] , \ML_int[3][23] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] ,
         \ML_int[3][8] , \ML_int[3][7] , \ML_int[3][3] , \ML_int[3][2] ,
         \ML_int[3][1] , \ML_int[3][0] , \ML_int[4][27] , \ML_int[4][26] ,
         \ML_int[4][25] , \ML_int[4][24] , \ML_int[4][23] , \ML_int[4][11] ,
         \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] , \ML_int[4][7] ,
         \ML_int[5][27] , \ML_int[5][26] , \ML_int[5][25] , \ML_int[5][24] ,
         \ML_int[5][23] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36;
  assign B[27] = \ML_int[5][27] ;
  assign B[26] = \ML_int[5][26] ;
  assign B[25] = \ML_int[5][25] ;
  assign B[24] = \ML_int[5][24] ;
  assign B[23] = \ML_int[5][23] ;

  MUX2_X2 M1_4_27 ( .A(\ML_int[4][27] ), .B(\ML_int[4][11] ), .S(SH[4]), .Z(
        \ML_int[5][27] ) );
  MUX2_X2 M1_4_26 ( .A(\ML_int[4][26] ), .B(\ML_int[4][10] ), .S(SH[4]), .Z(
        \ML_int[5][26] ) );
  MUX2_X2 M1_4_23 ( .A(\ML_int[4][23] ), .B(\ML_int[4][7] ), .S(SH[4]), .Z(
        \ML_int[5][23] ) );
  MUX2_X2 M1_3_27 ( .A(\ML_int[3][27] ), .B(\ML_int[3][19] ), .S(SH[3]), .Z(
        \ML_int[4][27] ) );
  MUX2_X2 M1_3_26 ( .A(\ML_int[3][26] ), .B(\ML_int[3][18] ), .S(SH[3]), .Z(
        \ML_int[4][26] ) );
  MUX2_X2 M1_3_23 ( .A(\ML_int[3][23] ), .B(\ML_int[3][15] ), .S(SH[3]), .Z(
        \ML_int[4][23] ) );
  MUX2_X2 M1_3_11 ( .A(\ML_int[3][11] ), .B(\ML_int[3][3] ), .S(SH[3]), .Z(
        \ML_int[4][11] ) );
  MUX2_X2 M1_3_10 ( .A(\ML_int[3][10] ), .B(\ML_int[3][2] ), .S(SH[3]), .Z(
        \ML_int[4][10] ) );
  MUX2_X2 M1_3_9 ( .A(\ML_int[3][9] ), .B(\ML_int[3][1] ), .S(SH[3]), .Z(
        \ML_int[4][9] ) );
  MUX2_X2 M1_2_27 ( .A(\ML_int[2][27] ), .B(\ML_int[2][23] ), .S(n28), .Z(
        \ML_int[3][27] ) );
  MUX2_X2 M1_2_26 ( .A(\ML_int[2][26] ), .B(\ML_int[2][22] ), .S(n28), .Z(
        \ML_int[3][26] ) );
  MUX2_X2 M1_2_25 ( .A(\ML_int[2][25] ), .B(\ML_int[2][21] ), .S(n28), .Z(
        \ML_int[3][25] ) );
  MUX2_X2 M1_2_24 ( .A(\ML_int[2][24] ), .B(\ML_int[2][20] ), .S(n28), .Z(
        \ML_int[3][24] ) );
  MUX2_X2 M1_2_23 ( .A(\ML_int[2][23] ), .B(\ML_int[2][19] ), .S(n28), .Z(
        \ML_int[3][23] ) );
  MUX2_X2 M1_2_19 ( .A(\ML_int[2][19] ), .B(\ML_int[2][15] ), .S(n28), .Z(
        \ML_int[3][19] ) );
  MUX2_X2 M1_2_18 ( .A(\ML_int[2][18] ), .B(\ML_int[2][14] ), .S(n28), .Z(
        \ML_int[3][18] ) );
  MUX2_X2 M1_2_15 ( .A(\ML_int[2][15] ), .B(\ML_int[2][11] ), .S(n28), .Z(
        \ML_int[3][15] ) );
  MUX2_X2 M1_2_11 ( .A(\ML_int[2][11] ), .B(\ML_int[2][7] ), .S(n28), .Z(
        \ML_int[3][11] ) );
  MUX2_X2 M1_2_10 ( .A(\ML_int[2][10] ), .B(\ML_int[2][6] ), .S(n28), .Z(
        \ML_int[3][10] ) );
  MUX2_X2 M1_2_9 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S(n28), .Z(
        \ML_int[3][9] ) );
  MUX2_X2 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(n28), .Z(
        \ML_int[3][8] ) );
  MUX2_X2 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(n28), .Z(
        \ML_int[3][7] ) );
  MUX2_X2 M1_1_27 ( .A(\ML_int[1][27] ), .B(\ML_int[1][27] ), .S(n32), .Z(
        \ML_int[2][27] ) );
  MUX2_X2 M1_1_26 ( .A(\ML_int[1][27] ), .B(\ML_int[1][24] ), .S(n32), .Z(
        \ML_int[2][26] ) );
  MUX2_X2 M1_1_23 ( .A(\ML_int[1][27] ), .B(\ML_int[1][21] ), .S(n32), .Z(
        \ML_int[2][23] ) );
  MUX2_X2 M1_1_22 ( .A(\ML_int[1][22] ), .B(\ML_int[1][20] ), .S(n32), .Z(
        \ML_int[2][22] ) );
  MUX2_X2 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S(n32), .Z(
        \ML_int[2][21] ) );
  MUX2_X2 M1_1_19 ( .A(\ML_int[1][19] ), .B(\ML_int[1][17] ), .S(n32), .Z(
        \ML_int[2][19] ) );
  MUX2_X2 M1_1_18 ( .A(\ML_int[1][18] ), .B(\ML_int[1][16] ), .S(n32), .Z(
        \ML_int[2][18] ) );
  MUX2_X2 M1_1_17 ( .A(\ML_int[1][17] ), .B(\ML_int[1][15] ), .S(n32), .Z(
        \ML_int[2][17] ) );
  MUX2_X2 M1_1_16 ( .A(\ML_int[1][16] ), .B(\ML_int[1][14] ), .S(n33), .Z(
        \ML_int[2][16] ) );
  MUX2_X2 M1_1_15 ( .A(\ML_int[1][15] ), .B(\ML_int[1][13] ), .S(n33), .Z(
        \ML_int[2][15] ) );
  MUX2_X2 M1_1_14 ( .A(\ML_int[1][14] ), .B(\ML_int[1][12] ), .S(n33), .Z(
        \ML_int[2][14] ) );
  MUX2_X2 M1_1_11 ( .A(\ML_int[1][11] ), .B(\ML_int[1][9] ), .S(n33), .Z(
        \ML_int[2][11] ) );
  MUX2_X2 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S(n33), .Z(
        \ML_int[2][10] ) );
  MUX2_X2 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S(n33), .Z(
        \ML_int[2][9] ) );
  MUX2_X2 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S(n33), .Z(
        \ML_int[2][8] ) );
  MUX2_X2 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S(n33), .Z(
        \ML_int[2][7] ) );
  MUX2_X2 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(n34), .Z(
        \ML_int[2][3] ) );
  MUX2_X2 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S(n34), .Z(
        \ML_int[2][2] ) );
  MUX2_X2 M1_0_24 ( .A(A[24]), .B(A[23]), .S(n30), .Z(\ML_int[1][24] ) );
  MUX2_X2 M1_0_22 ( .A(A[22]), .B(A[21]), .S(n30), .Z(\ML_int[1][22] ) );
  MUX2_X2 M1_0_21 ( .A(A[21]), .B(A[20]), .S(n30), .Z(\ML_int[1][21] ) );
  MUX2_X2 M1_0_20 ( .A(A[20]), .B(A[19]), .S(n30), .Z(\ML_int[1][20] ) );
  MUX2_X2 M1_0_19 ( .A(A[19]), .B(A[18]), .S(n30), .Z(\ML_int[1][19] ) );
  MUX2_X2 M1_0_18 ( .A(A[18]), .B(A[17]), .S(n30), .Z(\ML_int[1][18] ) );
  MUX2_X2 M1_0_17 ( .A(A[17]), .B(A[16]), .S(n30), .Z(\ML_int[1][17] ) );
  MUX2_X2 M1_0_16 ( .A(A[16]), .B(A[15]), .S(n30), .Z(\ML_int[1][16] ) );
  MUX2_X2 M1_0_15 ( .A(A[15]), .B(A[14]), .S(n30), .Z(\ML_int[1][15] ) );
  MUX2_X2 M1_0_14 ( .A(A[14]), .B(A[13]), .S(n30), .Z(\ML_int[1][14] ) );
  MUX2_X2 M1_0_13 ( .A(A[13]), .B(A[12]), .S(n30), .Z(\ML_int[1][13] ) );
  MUX2_X2 M1_0_12 ( .A(A[12]), .B(A[11]), .S(n30), .Z(\ML_int[1][12] ) );
  MUX2_X2 M1_0_11 ( .A(A[11]), .B(A[10]), .S(n29), .Z(\ML_int[1][11] ) );
  MUX2_X2 M1_0_10 ( .A(A[10]), .B(A[9]), .S(n29), .Z(\ML_int[1][10] ) );
  MUX2_X2 M1_0_9 ( .A(A[9]), .B(A[8]), .S(n29), .Z(\ML_int[1][9] ) );
  MUX2_X2 M1_0_8 ( .A(A[8]), .B(A[7]), .S(n29), .Z(\ML_int[1][8] ) );
  MUX2_X2 M1_0_7 ( .A(A[7]), .B(A[6]), .S(n29), .Z(\ML_int[1][7] ) );
  MUX2_X2 M1_0_6 ( .A(A[6]), .B(A[5]), .S(n29), .Z(\ML_int[1][6] ) );
  MUX2_X2 M1_0_4 ( .A(A[4]), .B(A[3]), .S(n29), .Z(\ML_int[1][4] ) );
  MUX2_X2 M1_0_3 ( .A(A[3]), .B(A[2]), .S(n29), .Z(\ML_int[1][3] ) );
  MUX2_X2 M1_0_2 ( .A(A[2]), .B(A[1]), .S(n29), .Z(\ML_int[1][2] ) );
  MUX2_X2 M1_0_1 ( .A(A[1]), .B(A[0]), .S(n29), .Z(\ML_int[1][1] ) );
  MUX2_X1 M1_2_16 ( .A(\ML_int[2][16] ), .B(\ML_int[2][12] ), .S(n28), .Z(
        \ML_int[3][16] ) );
  MUX2_X1 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S(n33), .Z(
        \ML_int[2][6] ) );
  MUX2_X2 M1_2_17 ( .A(\ML_int[2][17] ), .B(\ML_int[2][13] ), .S(n28), .Z(
        \ML_int[3][17] ) );
  MUX2_X2 M1_0_27 ( .A(A[27]), .B(A[26]), .S(n30), .Z(\ML_int[1][27] ) );
  NAND2_X1 U3 ( .A1(A[5]), .A2(n4), .ZN(n5) );
  NAND2_X4 U4 ( .A1(n25), .A2(n26), .ZN(\ML_int[5][25] ) );
  NAND2_X1 U5 ( .A1(\ML_int[1][3] ), .A2(n1), .ZN(n2) );
  NAND2_X2 U6 ( .A1(\ML_int[1][5] ), .A2(n35), .ZN(n3) );
  NAND2_X2 U7 ( .A1(n2), .A2(n3), .ZN(\ML_int[2][5] ) );
  INV_X1 U8 ( .A(n35), .ZN(n1) );
  NAND2_X1 U9 ( .A1(A[4]), .A2(n29), .ZN(n6) );
  NAND2_X2 U10 ( .A1(n5), .A2(n6), .ZN(\ML_int[1][5] ) );
  INV_X1 U11 ( .A(n29), .ZN(n4) );
  INV_X16 U12 ( .A(n31), .ZN(n30) );
  INV_X16 U13 ( .A(n31), .ZN(n29) );
  INV_X4 U14 ( .A(SH[0]), .ZN(n31) );
  INV_X4 U15 ( .A(n33), .ZN(n21) );
  INV_X4 U16 ( .A(SH[4]), .ZN(n24) );
  INV_X8 U17 ( .A(n27), .ZN(n28) );
  INV_X4 U18 ( .A(SH[2]), .ZN(n27) );
  NAND2_X4 U19 ( .A1(\ML_int[4][25] ), .A2(n24), .ZN(n25) );
  MUX2_X2 U20 ( .A(\ML_int[1][22] ), .B(\ML_int[1][24] ), .S(n21), .Z(
        \ML_int[2][24] ) );
  INV_X8 U21 ( .A(n35), .ZN(n32) );
  OAI21_X2 U22 ( .B1(n7), .B2(SH[3]), .A(n10), .ZN(\ML_int[4][25] ) );
  INV_X4 U23 ( .A(\ML_int[3][25] ), .ZN(n7) );
  NAND2_X2 U24 ( .A1(\ML_int[3][8] ), .A2(n16), .ZN(n8) );
  NAND2_X2 U25 ( .A1(\ML_int[3][0] ), .A2(SH[3]), .ZN(n9) );
  NAND2_X2 U26 ( .A1(n8), .A2(n9), .ZN(\ML_int[4][8] ) );
  NAND2_X4 U27 ( .A1(n17), .A2(n18), .ZN(\ML_int[4][24] ) );
  NAND2_X2 U28 ( .A1(\ML_int[3][16] ), .A2(SH[3]), .ZN(n18) );
  NAND2_X4 U29 ( .A1(\ML_int[4][8] ), .A2(SH[4]), .ZN(n20) );
  NAND2_X4 U30 ( .A1(n19), .A2(n20), .ZN(\ML_int[5][24] ) );
  NAND2_X4 U31 ( .A1(\ML_int[3][24] ), .A2(n16), .ZN(n17) );
  INV_X4 U32 ( .A(n35), .ZN(n34) );
  NAND2_X2 U33 ( .A1(\ML_int[4][9] ), .A2(SH[4]), .ZN(n26) );
  NAND2_X2 U34 ( .A1(\ML_int[3][17] ), .A2(SH[3]), .ZN(n10) );
  NAND2_X1 U35 ( .A1(\ML_int[1][13] ), .A2(n21), .ZN(n11) );
  NAND2_X1 U36 ( .A1(\ML_int[1][11] ), .A2(n33), .ZN(n12) );
  NAND2_X2 U37 ( .A1(n11), .A2(n12), .ZN(\ML_int[2][13] ) );
  NAND2_X1 U38 ( .A1(\ML_int[1][27] ), .A2(n13), .ZN(n14) );
  NAND2_X1 U39 ( .A1(\ML_int[1][27] ), .A2(n32), .ZN(n15) );
  NAND2_X2 U40 ( .A1(n14), .A2(n15), .ZN(\ML_int[2][25] ) );
  INV_X1 U41 ( .A(n32), .ZN(n13) );
  INV_X1 U42 ( .A(SH[3]), .ZN(n16) );
  NAND2_X4 U43 ( .A1(\ML_int[4][24] ), .A2(n24), .ZN(n19) );
  MUX2_X2 U44 ( .A(\ML_int[1][2] ), .B(\ML_int[1][4] ), .S(n35), .Z(
        \ML_int[2][4] ) );
  NAND2_X1 U45 ( .A1(\ML_int[1][12] ), .A2(n21), .ZN(n22) );
  NAND2_X1 U46 ( .A1(\ML_int[1][10] ), .A2(n33), .ZN(n23) );
  NAND2_X2 U47 ( .A1(n22), .A2(n23), .ZN(\ML_int[2][12] ) );
  MUX2_X2 U48 ( .A(\ML_int[1][18] ), .B(\ML_int[1][20] ), .S(n13), .Z(
        \ML_int[2][20] ) );
  INV_X32 U49 ( .A(n35), .ZN(n33) );
  INV_X32 U50 ( .A(SH[1]), .ZN(n35) );
  AND2_X1 U51 ( .A1(\ML_int[3][7] ), .A2(n16), .ZN(\ML_int[4][7] ) );
  AND2_X1 U52 ( .A1(\ML_int[2][3] ), .A2(n27), .ZN(\ML_int[3][3] ) );
  AND2_X1 U53 ( .A1(\ML_int[2][2] ), .A2(n27), .ZN(\ML_int[3][2] ) );
  AND2_X1 U54 ( .A1(\ML_int[1][1] ), .A2(n36), .ZN(\ML_int[3][1] ) );
  AND2_X1 U55 ( .A1(n36), .A2(\ML_int[1][0] ), .ZN(\ML_int[3][0] ) );
  NOR2_X1 U56 ( .A1(n32), .A2(n28), .ZN(n36) );
  AND2_X1 U57 ( .A1(A[0]), .A2(n31), .ZN(\ML_int[1][0] ) );
endmodule


module fpu_DW01_sub_7 ( A, B, CI, DIFF, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;
  wire   [14:1] carry;

  FA_X1 U2_13 ( .A(A[13]), .B(n18), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FA_X1 U2_12 ( .A(A[12]), .B(n17), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FA_X1 U2_11 ( .A(A[11]), .B(n16), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FA_X1 U2_10 ( .A(A[10]), .B(n15), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FA_X1 U2_9 ( .A(A[9]), .B(n14), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FA_X1 U2_8 ( .A(A[8]), .B(n13), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FA_X1 U2_7 ( .A(A[7]), .B(n12), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FA_X1 U2_6 ( .A(A[6]), .B(n11), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA_X1 U2_5 ( .A(A[5]), .B(n10), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n9), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_3 ( .A(A[3]), .B(n8), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA_X1 U2_2 ( .A(A[2]), .B(n7), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA_X1 U2_1 ( .A(A[1]), .B(n6), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  INV_X1 U1 ( .A(n3), .ZN(n1) );
  NAND2_X4 U2 ( .A1(n2), .A2(n3), .ZN(carry[1]) );
  XNOR2_X2 U3 ( .A(n5), .B(n1), .ZN(DIFF[0]) );
  INV_X4 U4 ( .A(n5), .ZN(n2) );
  INV_X4 U5 ( .A(A[0]), .ZN(n3) );
  INV_X4 U6 ( .A(carry[14]), .ZN(DIFF[14]) );
  INV_X4 U7 ( .A(B[0]), .ZN(n5) );
  INV_X4 U8 ( .A(B[1]), .ZN(n6) );
  INV_X4 U9 ( .A(B[2]), .ZN(n7) );
  INV_X4 U10 ( .A(B[3]), .ZN(n8) );
  INV_X4 U11 ( .A(B[4]), .ZN(n9) );
  INV_X4 U12 ( .A(B[5]), .ZN(n10) );
  INV_X4 U13 ( .A(B[6]), .ZN(n11) );
  INV_X4 U14 ( .A(B[7]), .ZN(n12) );
  INV_X4 U15 ( .A(B[8]), .ZN(n13) );
  INV_X4 U16 ( .A(B[9]), .ZN(n14) );
  INV_X4 U17 ( .A(B[10]), .ZN(n15) );
  INV_X4 U18 ( .A(B[11]), .ZN(n16) );
  INV_X4 U19 ( .A(B[12]), .ZN(n17) );
  INV_X4 U20 ( .A(B[13]), .ZN(n18) );
endmodule


module fpu_DW01_add_5 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n4;
  wire   [13:1] carry;

  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(SUM[14]), .S(SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  BUF_X32 U1 ( .A(A[0]), .Z(n1) );
  BUF_X32 U2 ( .A(B[0]), .Z(n2) );
  XOR2_X1 U3 ( .A(n2), .B(n1), .Z(SUM[0]) );
  NAND2_X2 U4 ( .A1(B[0]), .A2(A[0]), .ZN(n4) );
  INV_X4 U5 ( .A(n4), .ZN(carry[1]) );
endmodule


module fpu_DW01_ash_2 ( A, DATA_TC, SH, SH_TC, B );
  input [10:0] A;
  input [3:0] SH;
  output [10:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] , \ML_int[1][7] ,
         \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] , \ML_int[1][3] ,
         \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] , \ML_int[2][10] ,
         \ML_int[2][9] , \ML_int[2][8] , \ML_int[2][7] , \ML_int[2][6] ,
         \ML_int[2][5] , \ML_int[2][4] , \ML_int[2][3] , \ML_int[2][2] ,
         \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] , \ML_int[3][7] ,
         \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] , \ML_int[3][2] ,
         \ML_int[3][1] , \ML_int[3][0] , \ML_int[4][10] , \ML_int[4][9] ,
         \ML_int[4][8] , \ML_int[4][7] , \ML_int[4][6] , \ML_int[4][5] ,
         \ML_int[4][4] , \ML_int[4][3] , \ML_int[4][2] , \ML_int[4][1] ,
         \ML_int[4][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;
  assign B[10] = \ML_int[4][10] ;
  assign B[9] = \ML_int[4][9] ;
  assign B[8] = \ML_int[4][8] ;
  assign B[7] = \ML_int[4][7] ;
  assign B[6] = \ML_int[4][6] ;
  assign B[5] = \ML_int[4][5] ;
  assign B[4] = \ML_int[4][4] ;
  assign B[3] = \ML_int[4][3] ;
  assign B[2] = \ML_int[4][2] ;
  assign B[1] = \ML_int[4][1] ;
  assign B[0] = \ML_int[4][0] ;

  MUX2_X2 M1_3_10 ( .A(\ML_int[3][10] ), .B(\ML_int[3][2] ), .S(SH[3]), .Z(
        \ML_int[4][10] ) );
  MUX2_X2 M1_3_9 ( .A(\ML_int[3][9] ), .B(\ML_int[3][1] ), .S(SH[3]), .Z(
        \ML_int[4][9] ) );
  MUX2_X2 M1_3_8 ( .A(\ML_int[3][8] ), .B(\ML_int[3][0] ), .S(SH[3]), .Z(
        \ML_int[4][8] ) );
  MUX2_X2 M1_2_10 ( .A(\ML_int[2][10] ), .B(\ML_int[2][6] ), .S(SH[2]), .Z(
        \ML_int[3][10] ) );
  MUX2_X2 M1_2_9 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S(SH[2]), .Z(
        \ML_int[3][9] ) );
  MUX2_X2 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(SH[2]), .Z(
        \ML_int[3][8] ) );
  MUX2_X2 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(SH[2]), .Z(
        \ML_int[3][7] ) );
  MUX2_X2 M1_2_6 ( .A(\ML_int[2][6] ), .B(\ML_int[2][2] ), .S(SH[2]), .Z(
        \ML_int[3][6] ) );
  MUX2_X2 M1_2_5 ( .A(\ML_int[2][5] ), .B(n4), .S(SH[2]), .Z(\ML_int[3][5] )
         );
  MUX2_X2 M1_2_4 ( .A(\ML_int[2][4] ), .B(n2), .S(SH[2]), .Z(\ML_int[3][4] )
         );
  MUX2_X2 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S(SH[1]), .Z(
        \ML_int[2][10] ) );
  MUX2_X2 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S(SH[1]), .Z(
        \ML_int[2][9] ) );
  MUX2_X2 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S(SH[1]), .Z(
        \ML_int[2][8] ) );
  MUX2_X2 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S(SH[1]), .Z(
        \ML_int[2][7] ) );
  MUX2_X2 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S(SH[1]), .Z(
        \ML_int[2][6] ) );
  MUX2_X2 M1_1_5 ( .A(\ML_int[1][5] ), .B(\ML_int[1][3] ), .S(SH[1]), .Z(
        \ML_int[2][5] ) );
  MUX2_X2 M1_1_4 ( .A(\ML_int[1][4] ), .B(\ML_int[1][2] ), .S(SH[1]), .Z(
        \ML_int[2][4] ) );
  MUX2_X2 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(SH[1]), .Z(
        \ML_int[2][3] ) );
  MUX2_X2 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S(SH[1]), .Z(
        \ML_int[2][2] ) );
  MUX2_X2 M1_0_10 ( .A(A[10]), .B(A[9]), .S(SH[0]), .Z(\ML_int[1][10] ) );
  MUX2_X2 M1_0_9 ( .A(A[9]), .B(A[8]), .S(SH[0]), .Z(\ML_int[1][9] ) );
  MUX2_X2 M1_0_8 ( .A(A[8]), .B(A[7]), .S(SH[0]), .Z(\ML_int[1][8] ) );
  MUX2_X2 M1_0_7 ( .A(A[7]), .B(A[6]), .S(SH[0]), .Z(\ML_int[1][7] ) );
  MUX2_X2 M1_0_6 ( .A(A[6]), .B(A[5]), .S(SH[0]), .Z(\ML_int[1][6] ) );
  MUX2_X2 M1_0_5 ( .A(A[5]), .B(A[4]), .S(SH[0]), .Z(\ML_int[1][5] ) );
  MUX2_X2 M1_0_4 ( .A(A[4]), .B(A[3]), .S(SH[0]), .Z(\ML_int[1][4] ) );
  MUX2_X2 M1_0_3 ( .A(A[3]), .B(A[2]), .S(SH[0]), .Z(\ML_int[1][3] ) );
  MUX2_X2 M1_0_2 ( .A(A[2]), .B(A[1]), .S(SH[0]), .Z(\ML_int[1][2] ) );
  MUX2_X2 M1_0_1 ( .A(A[1]), .B(A[0]), .S(SH[0]), .Z(\ML_int[1][1] ) );
  AND2_X2 U3 ( .A1(A[0]), .A2(n1), .ZN(\ML_int[1][0] ) );
  INV_X4 U4 ( .A(SH[0]), .ZN(n1) );
  INV_X4 U5 ( .A(n11), .ZN(n2) );
  INV_X4 U6 ( .A(\ML_int[2][2] ), .ZN(n3) );
  INV_X4 U7 ( .A(n10), .ZN(n4) );
  INV_X4 U8 ( .A(\ML_int[2][3] ), .ZN(n5) );
  INV_X4 U9 ( .A(SH[3]), .ZN(n6) );
  INV_X4 U10 ( .A(SH[2]), .ZN(n7) );
  INV_X4 U11 ( .A(SH[1]), .ZN(n8) );
  AND2_X1 U12 ( .A1(\ML_int[3][7] ), .A2(n6), .ZN(\ML_int[4][7] ) );
  AND2_X1 U13 ( .A1(\ML_int[3][6] ), .A2(n6), .ZN(\ML_int[4][6] ) );
  AND2_X1 U14 ( .A1(\ML_int[3][5] ), .A2(n6), .ZN(\ML_int[4][5] ) );
  AND2_X1 U15 ( .A1(\ML_int[3][4] ), .A2(n6), .ZN(\ML_int[4][4] ) );
  NOR2_X1 U16 ( .A1(n5), .A2(n9), .ZN(\ML_int[4][3] ) );
  NOR2_X1 U17 ( .A1(n9), .A2(n3), .ZN(\ML_int[4][2] ) );
  NOR2_X1 U18 ( .A1(n9), .A2(n10), .ZN(\ML_int[4][1] ) );
  NOR2_X1 U19 ( .A1(n9), .A2(n11), .ZN(\ML_int[4][0] ) );
  NAND2_X1 U20 ( .A1(n7), .A2(n6), .ZN(n9) );
  NOR2_X1 U21 ( .A1(SH[2]), .A2(n3), .ZN(\ML_int[3][2] ) );
  NOR2_X1 U22 ( .A1(SH[2]), .A2(n10), .ZN(\ML_int[3][1] ) );
  NOR2_X1 U23 ( .A1(SH[2]), .A2(n11), .ZN(\ML_int[3][0] ) );
  NAND2_X1 U24 ( .A1(\ML_int[1][1] ), .A2(n8), .ZN(n10) );
  NAND2_X1 U25 ( .A1(\ML_int[1][0] ), .A2(n8), .ZN(n11) );
endmodule


module fpu_DW01_add_11 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   \A[9] , \A[8] , \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] ,
         \A[1] , \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83;
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign SUM[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign SUM[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign SUM[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  AND2_X2 U2 ( .A1(A[10]), .A2(B[10]), .ZN(n1) );
  NAND4_X2 U3 ( .A1(n46), .A2(n39), .A3(n78), .A4(n53), .ZN(n52) );
  INV_X4 U4 ( .A(A[11]), .ZN(n83) );
  INV_X4 U5 ( .A(n71), .ZN(n53) );
  AOI21_X2 U6 ( .B1(n23), .B2(n18), .A(n24), .ZN(n22) );
  AOI21_X2 U7 ( .B1(n62), .B2(n46), .A(n63), .ZN(n56) );
  INV_X4 U8 ( .A(n45), .ZN(n78) );
  OR2_X2 U9 ( .A1(n45), .A2(n71), .ZN(n2) );
  OR2_X2 U10 ( .A1(n25), .A2(n26), .ZN(n3) );
  OR2_X1 U11 ( .A1(n80), .A2(n71), .ZN(n4) );
  NOR2_X2 U12 ( .A1(n1), .A2(n48), .ZN(SUM[10]) );
  NOR2_X1 U13 ( .A1(A[10]), .A2(B[10]), .ZN(n48) );
  NAND2_X4 U14 ( .A1(n50), .A2(n51), .ZN(n72) );
  NAND2_X4 U15 ( .A1(n47), .A2(n49), .ZN(n35) );
  NAND2_X4 U16 ( .A1(n50), .A2(n51), .ZN(n49) );
  NAND2_X4 U17 ( .A1(n35), .A2(n36), .ZN(n31) );
  XNOR2_X1 U18 ( .A(n31), .B(n34), .ZN(SUM[16]) );
  INV_X8 U19 ( .A(n31), .ZN(n7) );
  NAND2_X4 U20 ( .A1(n82), .A2(n83), .ZN(n79) );
  NAND2_X1 U21 ( .A1(n51), .A2(n79), .ZN(n81) );
  NOR3_X2 U22 ( .A1(n44), .A2(n40), .A3(n45), .ZN(n37) );
  NOR2_X2 U23 ( .A1(n45), .A2(n69), .ZN(n68) );
  NAND2_X4 U24 ( .A1(n73), .A2(n74), .ZN(n46) );
  INV_X4 U25 ( .A(B[19]), .ZN(n5) );
  XNOR2_X2 U26 ( .A(n6), .B(n5), .ZN(SUM[19]) );
  OAI21_X4 U27 ( .B1(n7), .B2(n8), .A(n9), .ZN(n6) );
  AOI21_X4 U28 ( .B1(n10), .B2(n11), .A(n12), .ZN(n9) );
  INV_X4 U29 ( .A(n13), .ZN(n12) );
  NAND2_X2 U30 ( .A1(n14), .A2(n15), .ZN(n11) );
  NAND2_X2 U31 ( .A1(n10), .A2(n16), .ZN(n8) );
  INV_X4 U32 ( .A(n17), .ZN(n10) );
  NAND2_X2 U33 ( .A1(n18), .A2(n19), .ZN(n17) );
  XNOR2_X2 U34 ( .A(n21), .B(n20), .ZN(SUM[18]) );
  OAI21_X4 U35 ( .B1(n7), .B2(n3), .A(n22), .ZN(n21) );
  INV_X4 U36 ( .A(n14), .ZN(n24) );
  INV_X4 U37 ( .A(n15), .ZN(n23) );
  INV_X4 U38 ( .A(n18), .ZN(n25) );
  NAND2_X2 U39 ( .A1(n19), .A2(n13), .ZN(n20) );
  NAND2_X2 U40 ( .A1(B[18]), .A2(A[18]), .ZN(n13) );
  NAND2_X2 U41 ( .A1(n27), .A2(n28), .ZN(n19) );
  INV_X4 U42 ( .A(A[18]), .ZN(n28) );
  INV_X4 U43 ( .A(B[18]), .ZN(n27) );
  XNOR2_X2 U44 ( .A(n30), .B(n29), .ZN(SUM[17]) );
  OAI21_X4 U45 ( .B1(n7), .B2(n26), .A(n15), .ZN(n30) );
  INV_X4 U46 ( .A(n16), .ZN(n26) );
  NAND2_X2 U47 ( .A1(n14), .A2(n18), .ZN(n29) );
  NAND2_X2 U48 ( .A1(n32), .A2(n33), .ZN(n18) );
  INV_X4 U49 ( .A(A[17]), .ZN(n33) );
  INV_X4 U50 ( .A(B[17]), .ZN(n32) );
  NAND2_X2 U51 ( .A1(B[17]), .A2(A[17]), .ZN(n14) );
  OAI21_X4 U52 ( .B1(n37), .B2(n38), .A(n39), .ZN(n36) );
  OAI211_X2 U53 ( .C1(n40), .C2(n41), .A(n42), .B(n43), .ZN(n38) );
  NAND2_X2 U54 ( .A1(A[13]), .A2(B[13]), .ZN(n41) );
  INV_X4 U55 ( .A(n46), .ZN(n40) );
  NAND2_X2 U56 ( .A1(B[12]), .A2(A[12]), .ZN(n44) );
  INV_X4 U57 ( .A(n52), .ZN(n47) );
  NAND2_X2 U58 ( .A1(n16), .A2(n15), .ZN(n34) );
  NAND2_X2 U59 ( .A1(B[16]), .A2(A[16]), .ZN(n15) );
  NAND2_X2 U60 ( .A1(n54), .A2(n55), .ZN(n16) );
  INV_X4 U61 ( .A(A[16]), .ZN(n55) );
  INV_X4 U62 ( .A(B[16]), .ZN(n54) );
  XNOR2_X2 U63 ( .A(n56), .B(n57), .ZN(SUM[15]) );
  NOR2_X4 U64 ( .A1(n58), .A2(n59), .ZN(n57) );
  INV_X4 U65 ( .A(n42), .ZN(n59) );
  NAND2_X2 U66 ( .A1(B[15]), .A2(A[15]), .ZN(n42) );
  INV_X4 U67 ( .A(n39), .ZN(n58) );
  NAND2_X2 U68 ( .A1(n60), .A2(n61), .ZN(n39) );
  INV_X4 U69 ( .A(A[15]), .ZN(n61) );
  INV_X4 U70 ( .A(B[15]), .ZN(n60) );
  INV_X4 U71 ( .A(n43), .ZN(n63) );
  XNOR2_X2 U72 ( .A(n62), .B(n64), .ZN(SUM[14]) );
  OAI21_X4 U73 ( .B1(n65), .B2(n2), .A(n66), .ZN(n62) );
  NOR2_X4 U74 ( .A1(n67), .A2(n68), .ZN(n66) );
  INV_X4 U75 ( .A(n70), .ZN(n67) );
  INV_X4 U76 ( .A(n72), .ZN(n65) );
  NAND2_X2 U77 ( .A1(n46), .A2(n43), .ZN(n64) );
  NAND2_X2 U78 ( .A1(B[14]), .A2(A[14]), .ZN(n43) );
  INV_X4 U79 ( .A(A[14]), .ZN(n74) );
  INV_X4 U80 ( .A(B[14]), .ZN(n73) );
  XNOR2_X2 U81 ( .A(n76), .B(n75), .ZN(SUM[13]) );
  NAND2_X2 U82 ( .A1(n77), .A2(n69), .ZN(n76) );
  NAND2_X2 U83 ( .A1(n72), .A2(n53), .ZN(n77) );
  NAND2_X2 U84 ( .A1(n78), .A2(n70), .ZN(n75) );
  NAND2_X2 U85 ( .A1(B[13]), .A2(A[13]), .ZN(n70) );
  NOR2_X4 U86 ( .A1(A[13]), .A2(B[13]), .ZN(n45) );
  XNOR2_X2 U87 ( .A(n72), .B(n4), .ZN(SUM[12]) );
  NAND3_X4 U88 ( .A1(n79), .A2(B[10]), .A3(A[10]), .ZN(n50) );
  NOR2_X4 U89 ( .A1(A[12]), .A2(B[12]), .ZN(n71) );
  INV_X4 U90 ( .A(n69), .ZN(n80) );
  NAND2_X2 U91 ( .A1(B[12]), .A2(A[12]), .ZN(n69) );
  XNOR2_X2 U92 ( .A(n1), .B(n81), .ZN(SUM[11]) );
  NAND2_X2 U93 ( .A1(A[11]), .A2(B[11]), .ZN(n51) );
  INV_X4 U94 ( .A(B[11]), .ZN(n82) );
endmodule


module fpu_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [10:0] A;
  input [10:0] B;
  output [21:0] PRODUCT;
  input TC;
  wire   \ab[10][10] , \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] ,
         \ab[10][5] , \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] ,
         \ab[10][0] , \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] ,
         \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] ,
         \ab[9][1] , \ab[9][0] , \ab[8][10] , \ab[8][9] , \ab[8][8] ,
         \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] , \ab[8][3] ,
         \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][10] , \ab[7][9] ,
         \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] , \ab[7][4] ,
         \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] , \ab[6][10] ,
         \ab[6][9] , \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] ,
         \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] ,
         \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] ,
         \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] ,
         \ab[5][0] , \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] ,
         \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] ,
         \ab[4][1] , \ab[4][0] , \ab[3][10] , \ab[3][9] , \ab[3][8] ,
         \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][10] , \ab[2][9] ,
         \ab[2][8] , \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] ,
         \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] , \ab[1][10] ,
         \ab[1][9] , \ab[1][8] , \ab[1][7] , \ab[1][6] , \ab[1][5] ,
         \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[1][0] ,
         \ab[0][9] , \ab[0][8] , \ab[0][7] , \ab[0][6] , \ab[0][5] ,
         \ab[0][4] , \ab[0][3] , \ab[0][2] , \ab[0][1] , \CARRYB[10][9] ,
         \CARRYB[10][8] , \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] ,
         \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] ,
         \CARRYB[10][0] , \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] ,
         \CARRYB[9][6] , \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] ,
         \CARRYB[9][2] , \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][9] ,
         \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] ,
         \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] ,
         \CARRYB[8][0] , \CARRYB[7][9] , \CARRYB[7][8] , \CARRYB[7][7] ,
         \CARRYB[7][6] , \CARRYB[7][5] , \CARRYB[7][4] , \CARRYB[7][3] ,
         \CARRYB[7][2] , \CARRYB[7][1] , \CARRYB[7][0] , \CARRYB[6][9] ,
         \CARRYB[6][8] , \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] ,
         \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] ,
         \CARRYB[6][0] , \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] ,
         \CARRYB[5][6] , \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] ,
         \CARRYB[5][2] , \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][9] ,
         \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] ,
         \CARRYB[4][0] , \CARRYB[3][9] , \CARRYB[3][8] , \CARRYB[3][7] ,
         \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][4] , \CARRYB[3][3] ,
         \CARRYB[3][2] , \CARRYB[3][1] , \CARRYB[3][0] , \CARRYB[2][9] ,
         \CARRYB[2][8] , \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \CARRYB[1][9] , \CARRYB[1][8] , \CARRYB[1][7] ,
         \CARRYB[1][6] , \CARRYB[1][5] , \CARRYB[1][4] , \CARRYB[1][3] ,
         \CARRYB[1][2] , \CARRYB[1][1] , \CARRYB[1][0] , \SUMB[10][9] ,
         \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] , \SUMB[10][5] ,
         \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] , \SUMB[10][1] ,
         \SUMB[10][0] , \SUMB[9][9] , \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] ,
         \SUMB[9][5] , \SUMB[9][4] , \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] ,
         \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] ,
         \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][9] ,
         \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] , \SUMB[7][4] ,
         \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][9] , \SUMB[6][8] ,
         \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] , \SUMB[6][4] , \SUMB[6][3] ,
         \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] ,
         \SUMB[5][6] , \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] ,
         \SUMB[5][1] , \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][9] ,
         \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] ,
         \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][9] , \SUMB[1][8] ,
         \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] ,
         \SUMB[1][2] , \SUMB[1][1] , n3, n4, n5, n6, n7, n8, n9, n10, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69;
  wire   [19:16] CLA_CARRY;
  wire   [19:2] CLA_SUM;

  FA_X1 S4_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\SUMB[10][0] ) );
  FA_X1 S4_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA_X1 S4_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA_X1 S4_3 ( .A(\CARRYB[9][3] ), .B(\ab[10][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA_X1 S4_4 ( .A(\CARRYB[9][4] ), .B(\ab[10][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA_X1 S4_5 ( .A(\CARRYB[9][5] ), .B(\ab[10][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA_X1 S4_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA_X1 S4_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA_X1 S4_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA_X1 S5_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\ab[9][10] ), .CO(
        \CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA_X1 S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(CLA_SUM[9]) );
  FA_X1 S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA_X1 S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA_X1 S2_9_3 ( .A(\CARRYB[8][3] ), .B(\ab[9][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA_X1 S2_9_4 ( .A(\CARRYB[8][4] ), .B(\ab[9][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA_X1 S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA_X1 S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA_X1 S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA_X1 S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA_X1 S3_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\ab[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA_X1 S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(CLA_SUM[8]) );
  FA_X1 S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA_X1 S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA_X1 S2_8_3 ( .A(\CARRYB[7][3] ), .B(\ab[8][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA_X1 S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA_X1 S2_8_5 ( .A(\CARRYB[7][5] ), .B(\ab[8][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA_X1 S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA_X1 S2_8_7 ( .A(\ab[8][7] ), .B(\SUMB[7][8] ), .CI(\CARRYB[7][7] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA_X1 S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA_X1 S3_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\ab[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA_X1 S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(CLA_SUM[7]) );
  FA_X1 S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA_X1 S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA_X1 S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA_X1 S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA_X1 S2_7_5 ( .A(\CARRYB[6][5] ), .B(\ab[7][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA_X1 S2_7_6 ( .A(\CARRYB[6][6] ), .B(\ab[7][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA_X1 S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA_X1 S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA_X1 S3_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\ab[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA_X1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(CLA_SUM[6]) );
  FA_X1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA_X1 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA_X1 S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA_X1 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA_X1 S2_6_5 ( .A(\CARRYB[5][5] ), .B(\ab[6][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA_X1 S2_6_6 ( .A(\CARRYB[5][6] ), .B(\ab[6][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA_X1 S2_6_7 ( .A(\ab[6][7] ), .B(\SUMB[5][8] ), .CI(\CARRYB[5][7] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA_X1 S2_6_8 ( .A(\CARRYB[5][8] ), .B(\ab[6][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA_X1 S3_6_9 ( .A(\ab[6][9] ), .B(\ab[5][10] ), .CI(\CARRYB[5][9] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA_X1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(CLA_SUM[5]) );
  FA_X1 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA_X1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA_X1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA_X1 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA_X1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA_X1 S2_5_6 ( .A(\CARRYB[4][6] ), .B(\ab[5][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA_X1 S2_5_7 ( .A(\CARRYB[4][7] ), .B(\ab[5][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA_X1 S2_5_8 ( .A(\CARRYB[4][8] ), .B(\ab[5][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA_X1 S3_5_9 ( .A(\ab[5][9] ), .B(\ab[4][10] ), .CI(\CARRYB[4][9] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA_X1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(CLA_SUM[4]) );
  FA_X1 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA_X1 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA_X1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA_X1 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA_X1 S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA_X1 S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA_X1 S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA_X1 S2_4_8 ( .A(\SUMB[3][9] ), .B(\ab[4][8] ), .CI(\CARRYB[3][8] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA_X1 S3_4_9 ( .A(\ab[4][9] ), .B(\ab[3][10] ), .CI(\CARRYB[3][9] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA_X1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(CLA_SUM[3]) );
  FA_X1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA_X1 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA_X1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA_X1 S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA_X1 S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA_X1 S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA_X1 S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA_X1 S2_3_8 ( .A(\CARRYB[2][8] ), .B(\ab[3][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA_X1 S3_3_9 ( .A(\ab[3][9] ), .B(\ab[2][10] ), .CI(\CARRYB[2][9] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA_X1 S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(CLA_SUM[2]) );
  FA_X1 S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FA_X1 S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FA_X1 S2_2_3 ( .A(\ab[2][3] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FA_X1 S2_2_4 ( .A(\ab[2][4] ), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FA_X1 S2_2_5 ( .A(\ab[2][5] ), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FA_X1 S2_2_6 ( .A(\ab[2][6] ), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FA_X1 S2_2_7 ( .A(\ab[2][7] ), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FA_X1 S2_2_8 ( .A(\ab[2][8] ), .B(\CARRYB[1][8] ), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FA_X1 S3_2_9 ( .A(\CARRYB[1][9] ), .B(\ab[2][9] ), .CI(\ab[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  fpu_DW01_add_11 FS_1 ( .A({1'b0, n8, CLA_SUM[19:11], \SUMB[10][0] , 
        CLA_SUM[9:2]}), .B({n12, CLA_CARRY, n9, n5, n6, n10, n7, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM(
        PRODUCT[21:2]) );
  INV_X1 U2 ( .A(n56), .ZN(n3) );
  INV_X4 U3 ( .A(n3), .ZN(n4) );
  INV_X8 U4 ( .A(B[8]), .ZN(n56) );
  NOR2_X2 U5 ( .A1(n55), .A2(n53), .ZN(\ab[6][9] ) );
  INV_X16 U6 ( .A(B[9]), .ZN(n55) );
  NAND2_X4 U7 ( .A1(\ab[0][9] ), .A2(\ab[1][8] ), .ZN(n44) );
  NOR2_X1 U8 ( .A1(n61), .A2(n54), .ZN(\ab[7][3] ) );
  INV_X8 U9 ( .A(B[2]), .ZN(n62) );
  NOR2_X1 U10 ( .A1(n63), .A2(n54), .ZN(\ab[7][1] ) );
  INV_X8 U11 ( .A(B[0]), .ZN(n65) );
  NOR2_X1 U12 ( .A1(n59), .A2(n50), .ZN(\ab[3][5] ) );
  INV_X8 U13 ( .A(B[4]), .ZN(n60) );
  NOR2_X1 U14 ( .A1(n61), .A2(n52), .ZN(\ab[5][3] ) );
  NOR2_X1 U15 ( .A1(n69), .A2(n61), .ZN(\ab[8][3] ) );
  NOR2_X1 U16 ( .A1(n69), .A2(n62), .ZN(\ab[8][2] ) );
  INV_X8 U17 ( .A(B[1]), .ZN(n63) );
  NOR2_X1 U18 ( .A1(n69), .A2(n65), .ZN(\ab[8][0] ) );
  NOR2_X2 U19 ( .A1(n57), .A2(n52), .ZN(\ab[5][7] ) );
  NOR2_X2 U20 ( .A1(n58), .A2(n52), .ZN(\ab[5][6] ) );
  NOR2_X2 U21 ( .A1(n59), .A2(n52), .ZN(\ab[5][5] ) );
  NOR2_X1 U22 ( .A1(n69), .A2(n4), .ZN(\ab[8][8] ) );
  NOR2_X2 U23 ( .A1(n69), .A2(n57), .ZN(\ab[8][7] ) );
  NOR2_X2 U24 ( .A1(n69), .A2(n58), .ZN(\ab[8][6] ) );
  NOR2_X2 U25 ( .A1(n69), .A2(n59), .ZN(\ab[8][5] ) );
  NOR2_X1 U26 ( .A1(n60), .A2(n51), .ZN(\ab[4][4] ) );
  INV_X8 U27 ( .A(B[7]), .ZN(n57) );
  INV_X8 U28 ( .A(B[6]), .ZN(n58) );
  INV_X8 U29 ( .A(B[5]), .ZN(n59) );
  NOR2_X1 U30 ( .A1(n69), .A2(n60), .ZN(\ab[8][4] ) );
  NOR2_X1 U31 ( .A1(n61), .A2(n51), .ZN(\ab[4][3] ) );
  NOR2_X1 U32 ( .A1(n68), .A2(n62), .ZN(\ab[9][2] ) );
  NOR2_X1 U33 ( .A1(n62), .A2(n51), .ZN(\ab[4][2] ) );
  NOR2_X1 U34 ( .A1(n69), .A2(n63), .ZN(\ab[8][1] ) );
  NOR2_X1 U35 ( .A1(n63), .A2(n51), .ZN(\ab[4][1] ) );
  NOR2_X1 U36 ( .A1(n65), .A2(n54), .ZN(\ab[7][0] ) );
  NOR2_X1 U37 ( .A1(n65), .A2(n51), .ZN(\ab[4][0] ) );
  NOR2_X1 U38 ( .A1(n57), .A2(n50), .ZN(\ab[3][7] ) );
  NOR2_X1 U39 ( .A1(n57), .A2(n53), .ZN(\ab[6][7] ) );
  NOR2_X1 U40 ( .A1(n58), .A2(n53), .ZN(\ab[6][6] ) );
  NOR2_X1 U41 ( .A1(n58), .A2(n50), .ZN(\ab[3][6] ) );
  NOR2_X1 U42 ( .A1(n59), .A2(n53), .ZN(\ab[6][5] ) );
  NOR2_X1 U43 ( .A1(n68), .A2(n4), .ZN(\ab[9][8] ) );
  NOR2_X1 U44 ( .A1(n68), .A2(n57), .ZN(\ab[9][7] ) );
  NOR2_X1 U45 ( .A1(n68), .A2(n58), .ZN(\ab[9][6] ) );
  NOR2_X1 U46 ( .A1(n68), .A2(n59), .ZN(\ab[9][5] ) );
  NOR2_X1 U47 ( .A1(n68), .A2(n60), .ZN(\ab[9][4] ) );
  NOR2_X1 U48 ( .A1(n60), .A2(n52), .ZN(\ab[5][4] ) );
  NOR2_X1 U49 ( .A1(n68), .A2(n61), .ZN(\ab[9][3] ) );
  NOR2_X1 U50 ( .A1(n61), .A2(n50), .ZN(\ab[3][3] ) );
  NOR2_X1 U51 ( .A1(n62), .A2(n54), .ZN(\ab[7][2] ) );
  NOR2_X1 U52 ( .A1(n62), .A2(n50), .ZN(\ab[3][2] ) );
  NOR2_X1 U53 ( .A1(n67), .A2(n63), .ZN(\ab[10][1] ) );
  INV_X4 U54 ( .A(A[9]), .ZN(n68) );
  NOR2_X1 U55 ( .A1(n63), .A2(n53), .ZN(\ab[6][1] ) );
  NOR2_X1 U56 ( .A1(n63), .A2(n50), .ZN(\ab[3][1] ) );
  INV_X8 U57 ( .A(A[2]), .ZN(n49) );
  NOR2_X1 U58 ( .A1(n67), .A2(n65), .ZN(\ab[10][0] ) );
  NOR2_X1 U59 ( .A1(n65), .A2(n53), .ZN(\ab[6][0] ) );
  NOR2_X1 U60 ( .A1(n65), .A2(n50), .ZN(\ab[3][0] ) );
  NOR2_X1 U61 ( .A1(n57), .A2(n51), .ZN(\ab[4][7] ) );
  NOR2_X1 U62 ( .A1(n58), .A2(n51), .ZN(\ab[4][6] ) );
  NOR2_X1 U63 ( .A1(n57), .A2(n54), .ZN(\ab[7][7] ) );
  NOR2_X1 U64 ( .A1(n58), .A2(n54), .ZN(\ab[7][6] ) );
  NOR2_X1 U65 ( .A1(n59), .A2(n54), .ZN(\ab[7][5] ) );
  NOR2_X1 U66 ( .A1(n59), .A2(n51), .ZN(\ab[4][5] ) );
  NOR2_X1 U67 ( .A1(n60), .A2(n54), .ZN(\ab[7][4] ) );
  NOR2_X1 U68 ( .A1(n60), .A2(n50), .ZN(\ab[3][4] ) );
  INV_X4 U69 ( .A(B[10]), .ZN(n64) );
  NOR2_X1 U70 ( .A1(n67), .A2(n4), .ZN(\ab[10][8] ) );
  NOR2_X1 U71 ( .A1(n67), .A2(n57), .ZN(\ab[10][7] ) );
  NOR2_X1 U72 ( .A1(n67), .A2(n58), .ZN(\ab[10][6] ) );
  NOR2_X1 U73 ( .A1(n67), .A2(n59), .ZN(\ab[10][5] ) );
  NOR2_X1 U74 ( .A1(n67), .A2(n60), .ZN(\ab[10][4] ) );
  NOR2_X1 U75 ( .A1(n67), .A2(n61), .ZN(\ab[10][3] ) );
  NOR2_X1 U76 ( .A1(n61), .A2(n53), .ZN(\ab[6][3] ) );
  NOR2_X1 U77 ( .A1(n67), .A2(n62), .ZN(\ab[10][2] ) );
  NOR2_X1 U78 ( .A1(n62), .A2(n52), .ZN(\ab[5][2] ) );
  INV_X4 U79 ( .A(A[8]), .ZN(n69) );
  INV_X1 U80 ( .A(A[10]), .ZN(n67) );
  NOR2_X1 U81 ( .A1(n68), .A2(n63), .ZN(\ab[9][1] ) );
  INV_X8 U82 ( .A(A[7]), .ZN(n54) );
  NOR2_X1 U83 ( .A1(n63), .A2(n52), .ZN(\ab[5][1] ) );
  NOR2_X1 U84 ( .A1(n68), .A2(n65), .ZN(\ab[9][0] ) );
  NOR2_X1 U85 ( .A1(n65), .A2(n52), .ZN(\ab[5][0] ) );
  NOR2_X1 U86 ( .A1(n65), .A2(n49), .ZN(\ab[2][0] ) );
  AND2_X4 U87 ( .A1(\SUMB[10][4] ), .A2(\CARRYB[10][3] ), .ZN(n5) );
  AND2_X4 U88 ( .A1(\CARRYB[10][2] ), .A2(\SUMB[10][3] ), .ZN(n6) );
  AND2_X4 U89 ( .A1(\SUMB[10][1] ), .A2(\CARRYB[10][0] ), .ZN(n7) );
  XOR2_X2 U90 ( .A(\CARRYB[10][9] ), .B(\ab[10][10] ), .Z(n8) );
  AND2_X4 U91 ( .A1(\SUMB[10][5] ), .A2(\CARRYB[10][4] ), .ZN(n9) );
  AND2_X4 U92 ( .A1(\SUMB[10][2] ), .A2(\CARRYB[10][1] ), .ZN(n10) );
  XOR2_X1 U93 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Z(PRODUCT[1]) );
  AND2_X2 U94 ( .A1(\ab[10][10] ), .A2(\CARRYB[10][9] ), .ZN(n12) );
  NOR2_X2 U95 ( .A1(n58), .A2(n48), .ZN(\ab[1][6] ) );
  NOR2_X1 U96 ( .A1(n66), .A2(n65), .ZN(PRODUCT[0]) );
  NOR2_X2 U97 ( .A1(n55), .A2(n51), .ZN(\ab[4][9] ) );
  NOR2_X2 U98 ( .A1(n55), .A2(n52), .ZN(\ab[5][9] ) );
  NOR2_X2 U99 ( .A1(n66), .A2(n56), .ZN(\ab[0][8] ) );
  NOR2_X2 U100 ( .A1(n66), .A2(n58), .ZN(\ab[0][6] ) );
  NOR2_X2 U101 ( .A1(n57), .A2(n48), .ZN(\ab[1][7] ) );
  NOR2_X2 U102 ( .A1(n57), .A2(n49), .ZN(\ab[2][7] ) );
  NOR2_X2 U103 ( .A1(n14), .A2(n49), .ZN(\ab[2][10] ) );
  NOR2_X2 U104 ( .A1(n58), .A2(n49), .ZN(\ab[2][6] ) );
  NOR2_X2 U105 ( .A1(n59), .A2(n49), .ZN(\ab[2][5] ) );
  NOR2_X2 U106 ( .A1(n60), .A2(n49), .ZN(\ab[2][4] ) );
  NOR2_X2 U107 ( .A1(n61), .A2(n49), .ZN(\ab[2][3] ) );
  NOR2_X2 U108 ( .A1(n62), .A2(n49), .ZN(\ab[2][2] ) );
  NOR2_X2 U109 ( .A1(n63), .A2(n49), .ZN(\ab[2][1] ) );
  INV_X2 U110 ( .A(n16), .ZN(CLA_SUM[11]) );
  NOR2_X4 U111 ( .A1(n14), .A2(n48), .ZN(\ab[1][10] ) );
  NOR2_X1 U112 ( .A1(n67), .A2(n55), .ZN(\ab[10][9] ) );
  NOR2_X1 U113 ( .A1(n55), .A2(n50), .ZN(\ab[3][9] ) );
  NOR2_X1 U114 ( .A1(n55), .A2(n49), .ZN(\ab[2][9] ) );
  NOR2_X2 U115 ( .A1(n66), .A2(n57), .ZN(\ab[0][7] ) );
  NOR2_X2 U116 ( .A1(n66), .A2(n60), .ZN(\ab[0][4] ) );
  NOR2_X2 U117 ( .A1(n66), .A2(n59), .ZN(\ab[0][5] ) );
  NOR2_X2 U118 ( .A1(n66), .A2(n61), .ZN(\ab[0][3] ) );
  NOR2_X2 U119 ( .A1(n66), .A2(n62), .ZN(\ab[0][2] ) );
  NOR2_X2 U120 ( .A1(n66), .A2(n63), .ZN(\ab[0][1] ) );
  NOR2_X2 U121 ( .A1(n56), .A2(n49), .ZN(\ab[2][8] ) );
  NOR2_X2 U122 ( .A1(n56), .A2(n50), .ZN(\ab[3][8] ) );
  NOR2_X2 U123 ( .A1(n56), .A2(n51), .ZN(\ab[4][8] ) );
  NOR2_X2 U124 ( .A1(n56), .A2(n52), .ZN(\ab[5][8] ) );
  NOR2_X2 U125 ( .A1(n56), .A2(n53), .ZN(\ab[6][8] ) );
  NOR2_X1 U126 ( .A1(n4), .A2(n54), .ZN(\ab[7][8] ) );
  INV_X8 U127 ( .A(n13), .ZN(n14) );
  INV_X2 U128 ( .A(n64), .ZN(n13) );
  NOR2_X1 U129 ( .A1(n55), .A2(n54), .ZN(\ab[7][9] ) );
  NOR2_X1 U130 ( .A1(n69), .A2(n55), .ZN(\ab[8][9] ) );
  NOR2_X1 U131 ( .A1(n68), .A2(n55), .ZN(\ab[9][9] ) );
  NOR2_X1 U132 ( .A1(n65), .A2(n48), .ZN(\ab[1][0] ) );
  NOR2_X1 U133 ( .A1(n63), .A2(n48), .ZN(\ab[1][1] ) );
  NOR2_X1 U134 ( .A1(n62), .A2(n48), .ZN(\ab[1][2] ) );
  NOR2_X1 U135 ( .A1(n61), .A2(n48), .ZN(\ab[1][3] ) );
  NOR2_X1 U136 ( .A1(n60), .A2(n48), .ZN(\ab[1][4] ) );
  NOR2_X1 U137 ( .A1(n59), .A2(n48), .ZN(\ab[1][5] ) );
  NOR2_X1 U138 ( .A1(n67), .A2(n14), .ZN(\ab[10][10] ) );
  NOR2_X1 U139 ( .A1(n68), .A2(n14), .ZN(\ab[9][10] ) );
  NOR2_X1 U140 ( .A1(n69), .A2(n14), .ZN(\ab[8][10] ) );
  NOR2_X1 U141 ( .A1(n14), .A2(n54), .ZN(\ab[7][10] ) );
  NOR2_X1 U142 ( .A1(n14), .A2(n53), .ZN(\ab[6][10] ) );
  NOR2_X1 U143 ( .A1(n14), .A2(n52), .ZN(\ab[5][10] ) );
  NOR2_X1 U144 ( .A1(n14), .A2(n51), .ZN(\ab[4][10] ) );
  NOR2_X1 U145 ( .A1(n14), .A2(n50), .ZN(\ab[3][10] ) );
  NOR2_X4 U146 ( .A1(n64), .A2(n66), .ZN(n15) );
  XNOR2_X1 U147 ( .A(\SUMB[10][1] ), .B(\CARRYB[10][0] ), .ZN(n16) );
  INV_X8 U148 ( .A(n17), .ZN(CLA_SUM[12]) );
  XNOR2_X2 U149 ( .A(\SUMB[10][3] ), .B(\CARRYB[10][2] ), .ZN(n18) );
  XNOR2_X2 U150 ( .A(\SUMB[10][2] ), .B(\CARRYB[10][1] ), .ZN(n17) );
  INV_X4 U151 ( .A(n18), .ZN(CLA_SUM[13]) );
  XNOR2_X2 U152 ( .A(\SUMB[10][4] ), .B(\CARRYB[10][3] ), .ZN(n19) );
  INV_X4 U153 ( .A(n19), .ZN(CLA_SUM[14]) );
  XNOR2_X2 U154 ( .A(\SUMB[10][5] ), .B(\CARRYB[10][4] ), .ZN(n20) );
  INV_X4 U155 ( .A(n20), .ZN(CLA_SUM[15]) );
  NAND2_X2 U156 ( .A1(\SUMB[10][6] ), .A2(\CARRYB[10][5] ), .ZN(n21) );
  INV_X4 U157 ( .A(n21), .ZN(CLA_CARRY[16]) );
  XNOR2_X2 U158 ( .A(\CARRYB[10][5] ), .B(\SUMB[10][6] ), .ZN(n22) );
  INV_X4 U159 ( .A(n22), .ZN(CLA_SUM[16]) );
  NAND2_X2 U160 ( .A1(\SUMB[10][7] ), .A2(\CARRYB[10][6] ), .ZN(n23) );
  INV_X4 U161 ( .A(n23), .ZN(CLA_CARRY[17]) );
  XNOR2_X2 U162 ( .A(\CARRYB[10][6] ), .B(\SUMB[10][7] ), .ZN(n24) );
  INV_X4 U163 ( .A(n24), .ZN(CLA_SUM[17]) );
  NAND2_X2 U164 ( .A1(\SUMB[10][8] ), .A2(\CARRYB[10][7] ), .ZN(n25) );
  INV_X4 U165 ( .A(n25), .ZN(CLA_CARRY[18]) );
  XNOR2_X2 U166 ( .A(\CARRYB[10][7] ), .B(\SUMB[10][8] ), .ZN(n26) );
  INV_X4 U167 ( .A(n26), .ZN(CLA_SUM[18]) );
  NAND2_X2 U168 ( .A1(\SUMB[10][9] ), .A2(\CARRYB[10][8] ), .ZN(n27) );
  INV_X4 U169 ( .A(n27), .ZN(CLA_CARRY[19]) );
  XNOR2_X2 U170 ( .A(\CARRYB[10][8] ), .B(\SUMB[10][9] ), .ZN(n28) );
  INV_X4 U171 ( .A(n28), .ZN(CLA_SUM[19]) );
  NAND2_X2 U172 ( .A1(\ab[0][1] ), .A2(\ab[1][0] ), .ZN(n29) );
  INV_X4 U173 ( .A(n29), .ZN(\CARRYB[1][0] ) );
  NAND2_X2 U174 ( .A1(\ab[0][2] ), .A2(\ab[1][1] ), .ZN(n30) );
  INV_X4 U175 ( .A(n30), .ZN(\CARRYB[1][1] ) );
  XNOR2_X2 U176 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .ZN(n31) );
  INV_X4 U177 ( .A(n31), .ZN(\SUMB[1][1] ) );
  NAND2_X2 U178 ( .A1(\ab[0][3] ), .A2(\ab[1][2] ), .ZN(n32) );
  INV_X4 U179 ( .A(n32), .ZN(\CARRYB[1][2] ) );
  XNOR2_X2 U180 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .ZN(n33) );
  INV_X4 U181 ( .A(n33), .ZN(\SUMB[1][2] ) );
  NAND2_X2 U182 ( .A1(\ab[0][4] ), .A2(\ab[1][3] ), .ZN(n34) );
  INV_X4 U183 ( .A(n34), .ZN(\CARRYB[1][3] ) );
  XNOR2_X2 U184 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .ZN(n35) );
  INV_X4 U185 ( .A(n35), .ZN(\SUMB[1][3] ) );
  NAND2_X2 U186 ( .A1(\ab[0][5] ), .A2(\ab[1][4] ), .ZN(n36) );
  INV_X4 U187 ( .A(n36), .ZN(\CARRYB[1][4] ) );
  XNOR2_X2 U188 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .ZN(n37) );
  INV_X4 U189 ( .A(n37), .ZN(\SUMB[1][4] ) );
  NAND2_X2 U190 ( .A1(\ab[0][6] ), .A2(\ab[1][5] ), .ZN(n38) );
  INV_X4 U191 ( .A(n38), .ZN(\CARRYB[1][5] ) );
  XNOR2_X2 U192 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .ZN(n39) );
  INV_X4 U193 ( .A(n39), .ZN(\SUMB[1][5] ) );
  NAND2_X2 U194 ( .A1(\ab[0][7] ), .A2(\ab[1][6] ), .ZN(n40) );
  INV_X4 U195 ( .A(n40), .ZN(\CARRYB[1][6] ) );
  XNOR2_X2 U196 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .ZN(n41) );
  INV_X4 U197 ( .A(n41), .ZN(\SUMB[1][6] ) );
  NAND2_X2 U198 ( .A1(\ab[0][8] ), .A2(\ab[1][7] ), .ZN(n42) );
  INV_X4 U199 ( .A(n42), .ZN(\CARRYB[1][7] ) );
  XNOR2_X2 U200 ( .A(\ab[0][8] ), .B(\ab[1][7] ), .ZN(n43) );
  INV_X4 U201 ( .A(n43), .ZN(\SUMB[1][7] ) );
  INV_X4 U202 ( .A(n44), .ZN(\CARRYB[1][8] ) );
  XNOR2_X2 U203 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .ZN(n45) );
  INV_X4 U204 ( .A(n45), .ZN(\SUMB[1][8] ) );
  NAND2_X2 U205 ( .A1(n15), .A2(\ab[1][9] ), .ZN(n46) );
  INV_X4 U206 ( .A(n46), .ZN(\CARRYB[1][9] ) );
  XNOR2_X2 U207 ( .A(n15), .B(\ab[1][9] ), .ZN(n47) );
  INV_X4 U208 ( .A(n47), .ZN(\SUMB[1][9] ) );
  INV_X16 U209 ( .A(A[0]), .ZN(n66) );
  INV_X16 U210 ( .A(A[1]), .ZN(n48) );
  INV_X16 U211 ( .A(B[3]), .ZN(n61) );
  INV_X16 U212 ( .A(A[3]), .ZN(n50) );
  INV_X16 U213 ( .A(A[4]), .ZN(n51) );
  INV_X16 U214 ( .A(A[5]), .ZN(n52) );
  INV_X16 U215 ( .A(A[6]), .ZN(n53) );
  NOR2_X4 U216 ( .A1(n55), .A2(n48), .ZN(\ab[1][9] ) );
  NOR2_X4 U217 ( .A1(n66), .A2(n55), .ZN(\ab[0][9] ) );
  NOR2_X4 U218 ( .A1(n56), .A2(n48), .ZN(\ab[1][8] ) );
  NOR2_X4 U219 ( .A1(n60), .A2(n53), .ZN(\ab[6][4] ) );
  NOR2_X4 U220 ( .A1(n62), .A2(n53), .ZN(\ab[6][2] ) );
endmodule


module fpu_DW01_inc_5 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  XOR2_X1 U2 ( .A(n4), .B(A[1]), .Z(SUM[1]) );
  NAND3_X4 U3 ( .A1(A[8]), .A2(A[7]), .A3(A[9]), .ZN(n30) );
  AND3_X4 U4 ( .A1(A[4]), .A2(A[5]), .A3(n11), .ZN(n2) );
  INV_X1 U5 ( .A(A[0]), .ZN(n3) );
  INV_X4 U6 ( .A(n3), .ZN(n4) );
  NAND4_X1 U7 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(n19) );
  INV_X4 U8 ( .A(n4), .ZN(SUM[0]) );
  NAND2_X4 U9 ( .A1(A[4]), .A2(A[3]), .ZN(n29) );
  INV_X2 U10 ( .A(A[3]), .ZN(n22) );
  NAND2_X1 U11 ( .A1(n2), .A2(A[6]), .ZN(n15) );
  INV_X1 U12 ( .A(A[6]), .ZN(n16) );
  NAND2_X4 U13 ( .A1(n26), .A2(n27), .ZN(n25) );
  NOR2_X4 U14 ( .A1(n28), .A2(n29), .ZN(n27) );
  INV_X8 U15 ( .A(n25), .ZN(SUM[10]) );
  CLKBUF_X2 U16 ( .A(A[2]), .Z(n5) );
  INV_X2 U17 ( .A(A[4]), .ZN(n20) );
  INV_X1 U18 ( .A(A[9]), .ZN(n7) );
  XNOR2_X1 U19 ( .A(A[7]), .B(n15), .ZN(SUM[7]) );
  NOR2_X2 U20 ( .A1(n23), .A2(n24), .ZN(n21) );
  INV_X1 U21 ( .A(A[8]), .ZN(n9) );
  NAND3_X2 U22 ( .A1(A[0]), .A2(A[2]), .A3(A[1]), .ZN(n28) );
  NOR2_X2 U23 ( .A1(n13), .A2(n14), .ZN(n12) );
  NOR2_X2 U24 ( .A1(n8), .A2(n9), .ZN(n6) );
  INV_X1 U25 ( .A(A[5]), .ZN(n18) );
  NAND2_X1 U26 ( .A1(A[6]), .A2(A[5]), .ZN(n31) );
  NAND2_X1 U27 ( .A1(A[7]), .A2(A[6]), .ZN(n13) );
  NOR2_X1 U28 ( .A1(n19), .A2(n20), .ZN(n17) );
  NAND2_X1 U29 ( .A1(A[4]), .A2(A[5]), .ZN(n14) );
  NAND2_X1 U30 ( .A1(A[1]), .A2(n4), .ZN(n24) );
  NOR2_X2 U31 ( .A1(n30), .A2(n31), .ZN(n26) );
  XNOR2_X2 U32 ( .A(n6), .B(n7), .ZN(SUM[9]) );
  XNOR2_X2 U33 ( .A(n10), .B(n9), .ZN(SUM[8]) );
  INV_X4 U34 ( .A(n8), .ZN(n10) );
  NAND2_X2 U35 ( .A1(n11), .A2(n12), .ZN(n8) );
  XNOR2_X2 U36 ( .A(n2), .B(n16), .ZN(SUM[6]) );
  XNOR2_X2 U37 ( .A(n17), .B(n18), .ZN(SUM[5]) );
  XNOR2_X2 U38 ( .A(n11), .B(n20), .ZN(SUM[4]) );
  INV_X4 U39 ( .A(n19), .ZN(n11) );
  XNOR2_X2 U40 ( .A(n21), .B(n22), .ZN(SUM[3]) );
  INV_X4 U41 ( .A(A[2]), .ZN(n23) );
  XNOR2_X2 U42 ( .A(n5), .B(n24), .ZN(SUM[2]) );
endmodule


module fpu_DW_rash_2 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [2:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   n2, n3, n4, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170;

  OAI211_X2 U3 ( .C1(SH[2]), .C2(n152), .A(1'b1), .B(n153), .ZN(B[10]) );
  OAI211_X2 U4 ( .C1(SH[2]), .C2(n138), .A(1'b1), .B(n139), .ZN(B[11]) );
  OAI211_X2 U5 ( .C1(n132), .C2(SH[2]), .A(1'b1), .B(n133), .ZN(B[12]) );
  NAND2_X2 U6 ( .A1(n118), .A2(n119), .ZN(B[13]) );
  OAI21_X4 U7 ( .B1(n94), .B2(n112), .A(n113), .ZN(B[14]) );
  OAI211_X2 U8 ( .C1(n94), .C2(n106), .A(1'b1), .B(n107), .ZN(B[15]) );
  OAI211_X2 U9 ( .C1(SH[2]), .C2(n96), .A(1'b1), .B(n97), .ZN(B[16]) );
  OAI211_X2 U10 ( .C1(n74), .C2(n94), .A(1'b1), .B(n95), .ZN(B[17]) );
  NAND2_X2 U11 ( .A1(n79), .A2(n80), .ZN(B[1]) );
  INV_X4 U12 ( .A(n76), .ZN(B[20]) );
  INV_X4 U13 ( .A(n72), .ZN(B[21]) );
  NAND2_X2 U14 ( .A1(n65), .A2(n66), .ZN(B[2]) );
  NAND2_X2 U15 ( .A1(n55), .A2(n56), .ZN(B[3]) );
  AOI21_X1 U16 ( .B1(A[19]), .B2(n20), .A(n105), .ZN(n135) );
  AOI21_X1 U17 ( .B1(A[15]), .B2(n20), .A(n2), .ZN(n100) );
  AND2_X2 U18 ( .A1(n92), .A2(n25), .ZN(B[18]) );
  INV_X4 U19 ( .A(SH[1]), .ZN(n19) );
  INV_X4 U20 ( .A(SH[0]), .ZN(n22) );
  INV_X4 U21 ( .A(n17), .ZN(n16) );
  AND2_X2 U22 ( .A1(A[14]), .A2(n22), .ZN(n2) );
  AND2_X2 U23 ( .A1(A[16]), .A2(n54), .ZN(n3) );
  AND2_X2 U24 ( .A1(A[10]), .A2(n22), .ZN(n4) );
  AND2_X2 U25 ( .A1(n90), .A2(n25), .ZN(B[19]) );
  NAND2_X1 U26 ( .A1(A[7]), .A2(n84), .ZN(n159) );
  NAND2_X1 U27 ( .A1(A[7]), .A2(n15), .ZN(n146) );
  INV_X1 U28 ( .A(A[4]), .ZN(n71) );
  NAND2_X1 U29 ( .A1(A[4]), .A2(n14), .ZN(n169) );
  NAND2_X1 U30 ( .A1(A[14]), .A2(n54), .ZN(n156) );
  NAND2_X1 U31 ( .A1(A[14]), .A2(n84), .ZN(n121) );
  NAND2_X1 U32 ( .A1(A[18]), .A2(n14), .ZN(n116) );
  NAND2_X1 U33 ( .A1(A[18]), .A2(n84), .ZN(n125) );
  NAND2_X1 U34 ( .A1(A[18]), .A2(n22), .ZN(n136) );
  INV_X4 U35 ( .A(SH[2]), .ZN(n94) );
  NAND2_X2 U36 ( .A1(n49), .A2(n50), .ZN(B[4]) );
  NAND2_X2 U37 ( .A1(n46), .A2(n47), .ZN(B[5]) );
  NAND2_X2 U38 ( .A1(n41), .A2(n42), .ZN(B[6]) );
  NAND2_X2 U39 ( .A1(n36), .A2(n37), .ZN(B[7]) );
  NAND2_X2 U40 ( .A1(n30), .A2(n31), .ZN(B[8]) );
  NAND2_X2 U41 ( .A1(n23), .A2(n24), .ZN(B[9]) );
  NAND2_X2 U42 ( .A1(n98), .A2(n99), .ZN(n77) );
  NAND2_X2 U49 ( .A1(n54), .A2(n12), .ZN(n74) );
  INV_X4 U50 ( .A(n17), .ZN(n12) );
  NOR2_X4 U51 ( .A1(n21), .A2(n13), .ZN(n111) );
  INV_X4 U52 ( .A(n16), .ZN(n13) );
  NAND2_X1 U53 ( .A1(A[19]), .A2(n84), .ZN(n115) );
  NAND2_X1 U54 ( .A1(A[19]), .A2(n15), .ZN(n110) );
  NAND2_X1 U55 ( .A1(A[6]), .A2(n15), .ZN(n160) );
  NAND2_X1 U56 ( .A1(A[6]), .A2(n84), .ZN(n82) );
  INV_X1 U57 ( .A(A[6]), .ZN(n64) );
  NAND2_X1 U58 ( .A1(A[10]), .A2(n84), .ZN(n129) );
  NAND2_X1 U59 ( .A1(n15), .A2(A[10]), .ZN(n164) );
  NAND2_X1 U60 ( .A1(A[20]), .A2(n15), .ZN(n99) );
  NAND2_X1 U61 ( .A1(A[17]), .A2(n15), .ZN(n126) );
  NAND2_X1 U62 ( .A1(A[17]), .A2(n84), .ZN(n103) );
  NAND2_X1 U63 ( .A1(A[5]), .A2(n84), .ZN(n168) );
  NAND2_X1 U64 ( .A1(A[5]), .A2(n54), .ZN(n83) );
  NAND2_X1 U65 ( .A1(A[20]), .A2(n84), .ZN(n109) );
  INV_X2 U66 ( .A(A[21]), .ZN(n17) );
  OAI21_X2 U67 ( .B1(n135), .B2(n19), .A(n103), .ZN(n134) );
  AOI21_X1 U68 ( .B1(A[11]), .B2(n20), .A(n4), .ZN(n51) );
  NAND2_X1 U69 ( .A1(A[11]), .A2(n14), .ZN(n150) );
  NAND2_X1 U70 ( .A1(A[11]), .A2(n84), .ZN(n163) );
  NAND2_X1 U71 ( .A1(A[9]), .A2(n84), .ZN(n52) );
  NAND2_X1 U72 ( .A1(A[9]), .A2(n14), .ZN(n130) );
  NAND2_X1 U73 ( .A1(A[8]), .A2(n14), .ZN(n53) );
  NAND2_X1 U74 ( .A1(A[8]), .A2(n84), .ZN(n145) );
  INV_X16 U75 ( .A(SH[2]), .ZN(n25) );
  NOR2_X4 U76 ( .A1(n18), .A2(n20), .ZN(n14) );
  NOR2_X4 U77 ( .A1(n18), .A2(n20), .ZN(n15) );
  INV_X8 U78 ( .A(n58), .ZN(n84) );
  INV_X8 U79 ( .A(n94), .ZN(n27) );
  INV_X32 U80 ( .A(n19), .ZN(n18) );
  INV_X32 U81 ( .A(n22), .ZN(n20) );
  INV_X32 U82 ( .A(n22), .ZN(n21) );
  NAND2_X2 U83 ( .A1(n25), .A2(n26), .ZN(n24) );
  NAND2_X2 U84 ( .A1(n27), .A2(n28), .ZN(n23) );
  NAND2_X2 U85 ( .A1(n32), .A2(n25), .ZN(n31) );
  NAND2_X2 U86 ( .A1(n27), .A2(n33), .ZN(n30) );
  NAND2_X2 U87 ( .A1(n38), .A2(n25), .ZN(n37) );
  NAND2_X2 U88 ( .A1(n27), .A2(n39), .ZN(n36) );
  NAND2_X2 U89 ( .A1(n43), .A2(n25), .ZN(n42) );
  NAND2_X2 U90 ( .A1(n27), .A2(n44), .ZN(n41) );
  NAND2_X2 U91 ( .A1(n25), .A2(n29), .ZN(n47) );
  NAND2_X2 U92 ( .A1(n27), .A2(n26), .ZN(n46) );
  NAND2_X2 U93 ( .A1(n27), .A2(n32), .ZN(n50) );
  OAI211_X2 U94 ( .C1(n51), .C2(n19), .A(n52), .B(n53), .ZN(n32) );
  NAND2_X2 U95 ( .A1(n34), .A2(n25), .ZN(n49) );
  NAND2_X2 U96 ( .A1(n27), .A2(n38), .ZN(n56) );
  NAND2_X2 U97 ( .A1(n60), .A2(n25), .ZN(n55) );
  INV_X4 U98 ( .A(n35), .ZN(n60) );
  MUX2_X2 U99 ( .A(n61), .B(n62), .S(n18), .Z(n35) );
  MUX2_X2 U100 ( .A(n63), .B(n64), .S(n20), .Z(n62) );
  NAND2_X2 U101 ( .A1(n68), .A2(n25), .ZN(n66) );
  INV_X4 U102 ( .A(n40), .ZN(n68) );
  MUX2_X2 U103 ( .A(n69), .B(n70), .S(n18), .Z(n40) );
  MUX2_X2 U104 ( .A(n71), .B(n63), .S(n21), .Z(n70) );
  INV_X4 U105 ( .A(A[5]), .ZN(n63) );
  NAND2_X2 U106 ( .A1(n27), .A2(n43), .ZN(n65) );
  NAND2_X2 U107 ( .A1(n73), .A2(n25), .ZN(n72) );
  INV_X4 U108 ( .A(n74), .ZN(n73) );
  NAND2_X2 U109 ( .A1(n77), .A2(n25), .ZN(n76) );
  NAND2_X2 U110 ( .A1(n27), .A2(n29), .ZN(n80) );
  NAND3_X2 U111 ( .A1(n81), .A2(n82), .A3(n83), .ZN(n29) );
  NAND2_X2 U112 ( .A1(n85), .A2(n18), .ZN(n81) );
  MUX2_X2 U113 ( .A(A[7]), .B(A[8]), .S(n21), .Z(n85) );
  NAND2_X2 U114 ( .A1(n86), .A2(n25), .ZN(n79) );
  INV_X4 U115 ( .A(n45), .ZN(n86) );
  MUX2_X2 U116 ( .A(n57), .B(n61), .S(n18), .Z(n45) );
  MUX2_X2 U117 ( .A(n87), .B(n71), .S(n21), .Z(n61) );
  MUX2_X2 U118 ( .A(n88), .B(n89), .S(n21), .Z(n57) );
  NAND2_X2 U119 ( .A1(n75), .A2(n25), .ZN(n95) );
  NAND2_X2 U120 ( .A1(n27), .A2(n77), .ZN(n97) );
  NAND2_X2 U121 ( .A1(n16), .A2(n84), .ZN(n98) );
  OAI211_X2 U122 ( .C1(n100), .C2(n19), .A(n101), .B(n102), .ZN(n33) );
  NAND2_X2 U123 ( .A1(A[12]), .A2(n14), .ZN(n102) );
  INV_X4 U124 ( .A(n78), .ZN(n96) );
  OAI211_X2 U125 ( .C1(n135), .C2(n19), .A(n103), .B(n104), .ZN(n78) );
  NAND2_X2 U126 ( .A1(A[16]), .A2(n54), .ZN(n104) );
  NAND2_X2 U127 ( .A1(n91), .A2(n25), .ZN(n107) );
  INV_X4 U128 ( .A(n90), .ZN(n106) );
  NAND3_X2 U129 ( .A1(n108), .A2(n109), .A3(n110), .ZN(n90) );
  NAND2_X2 U130 ( .A1(n111), .A2(n18), .ZN(n108) );
  NAND2_X2 U131 ( .A1(n93), .A2(n25), .ZN(n113) );
  INV_X4 U132 ( .A(n92), .ZN(n112) );
  NAND3_X2 U133 ( .A1(n114), .A2(n115), .A3(n116), .ZN(n92) );
  NAND2_X2 U134 ( .A1(n117), .A2(n18), .ZN(n114) );
  MUX2_X2 U135 ( .A(A[20]), .B(n16), .S(n21), .Z(n117) );
  NAND2_X2 U136 ( .A1(n25), .A2(n28), .ZN(n119) );
  NAND3_X2 U137 ( .A1(n120), .A2(n121), .A3(n122), .ZN(n28) );
  NAND2_X2 U138 ( .A1(A[13]), .A2(n54), .ZN(n122) );
  NAND2_X2 U139 ( .A1(n123), .A2(n18), .ZN(n120) );
  MUX2_X2 U140 ( .A(A[15]), .B(A[16]), .S(n21), .Z(n123) );
  NAND2_X2 U141 ( .A1(n27), .A2(n75), .ZN(n118) );
  NAND3_X2 U142 ( .A1(n124), .A2(n125), .A3(n126), .ZN(n75) );
  NAND2_X2 U143 ( .A1(n127), .A2(n18), .ZN(n124) );
  MUX2_X2 U144 ( .A(A[19]), .B(A[20]), .S(n21), .Z(n127) );
  NAND3_X2 U145 ( .A1(n128), .A2(n129), .A3(n130), .ZN(n26) );
  NAND2_X2 U146 ( .A1(n131), .A2(n18), .ZN(n128) );
  MUX2_X2 U147 ( .A(A[11]), .B(A[12]), .S(n21), .Z(n131) );
  OAI21_X4 U148 ( .B1(n134), .B2(n3), .A(n27), .ZN(n133) );
  INV_X4 U149 ( .A(n136), .ZN(n105) );
  INV_X4 U150 ( .A(n137), .ZN(n132) );
  OAI211_X2 U151 ( .C1(n100), .C2(n19), .A(n101), .B(n102), .ZN(n137) );
  NAND2_X2 U152 ( .A1(A[13]), .A2(n84), .ZN(n101) );
  NAND2_X2 U153 ( .A1(n27), .A2(n91), .ZN(n139) );
  NAND3_X2 U154 ( .A1(n140), .A2(n141), .A3(n142), .ZN(n91) );
  NAND2_X2 U155 ( .A1(A[15]), .A2(n54), .ZN(n142) );
  NAND2_X2 U156 ( .A1(A[16]), .A2(n84), .ZN(n141) );
  NAND2_X2 U157 ( .A1(n143), .A2(n18), .ZN(n140) );
  MUX2_X2 U158 ( .A(A[17]), .B(A[18]), .S(n20), .Z(n143) );
  NAND3_X2 U159 ( .A1(n144), .A2(n145), .A3(n146), .ZN(n38) );
  NAND2_X2 U160 ( .A1(n147), .A2(n18), .ZN(n144) );
  MUX2_X2 U161 ( .A(A[9]), .B(A[10]), .S(n21), .Z(n147) );
  INV_X4 U162 ( .A(n39), .ZN(n138) );
  NAND3_X2 U163 ( .A1(n148), .A2(n149), .A3(n150), .ZN(n39) );
  NAND2_X2 U164 ( .A1(A[12]), .A2(n84), .ZN(n149) );
  NAND2_X2 U165 ( .A1(n151), .A2(n18), .ZN(n148) );
  MUX2_X2 U166 ( .A(A[13]), .B(A[14]), .S(n20), .Z(n151) );
  NAND2_X2 U167 ( .A1(n27), .A2(n93), .ZN(n153) );
  NAND3_X2 U168 ( .A1(n154), .A2(n155), .A3(n156), .ZN(n93) );
  NAND2_X2 U169 ( .A1(A[15]), .A2(n84), .ZN(n155) );
  NAND2_X2 U170 ( .A1(n157), .A2(n18), .ZN(n154) );
  MUX2_X2 U171 ( .A(A[16]), .B(A[17]), .S(n21), .Z(n157) );
  NAND3_X2 U172 ( .A1(n158), .A2(n159), .A3(n160), .ZN(n43) );
  NAND2_X2 U173 ( .A1(n161), .A2(n18), .ZN(n158) );
  MUX2_X2 U174 ( .A(A[8]), .B(A[9]), .S(n20), .Z(n161) );
  INV_X4 U175 ( .A(n44), .ZN(n152) );
  NAND3_X2 U176 ( .A1(n162), .A2(n163), .A3(n164), .ZN(n44) );
  NAND2_X2 U177 ( .A1(n165), .A2(n18), .ZN(n162) );
  MUX2_X2 U178 ( .A(A[12]), .B(A[13]), .S(n20), .Z(n165) );
  OAI21_X4 U179 ( .B1(SH[2]), .B2(n48), .A(n166), .ZN(B[0]) );
  NAND2_X2 U180 ( .A1(n27), .A2(n34), .ZN(n166) );
  NAND3_X2 U181 ( .A1(n167), .A2(n168), .A3(n169), .ZN(n34) );
  NOR2_X4 U182 ( .A1(n18), .A2(n20), .ZN(n54) );
  NAND2_X2 U183 ( .A1(n21), .A2(n19), .ZN(n58) );
  NAND2_X2 U184 ( .A1(n170), .A2(n18), .ZN(n167) );
  MUX2_X2 U185 ( .A(A[6]), .B(A[7]), .S(n20), .Z(n170) );
  MUX2_X2 U186 ( .A(n67), .B(n69), .S(n18), .Z(n48) );
  MUX2_X2 U187 ( .A(n89), .B(n87), .S(n20), .Z(n69) );
  INV_X4 U188 ( .A(A[3]), .ZN(n87) );
  INV_X4 U189 ( .A(A[2]), .ZN(n89) );
  MUX2_X2 U190 ( .A(n59), .B(n88), .S(n21), .Z(n67) );
  INV_X4 U191 ( .A(A[1]), .ZN(n88) );
  INV_X4 U192 ( .A(A[0]), .ZN(n59) );
endmodule


module fpu_DW01_ash_4 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [2:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][20] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][0] , \ML_int[2][20] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][16] , \ML_int[2][15] ,
         \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][11] , \ML_int[2][9] ,
         \ML_int[2][8] , \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] ,
         \ML_int[2][4] , \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] ,
         \ML_int[2][0] , net85895, net85899, net85903, net88351, net88458,
         net88600, net88672, net88766, net88778, net88783, net88852, net88861,
         net88908, net88921, net88980, net88998, net89007, net89012, net89040,
         net89046, net89052, net89050, net89170, net89236, net89240, net89257,
         net89339, net89358, net89354, net89420, net89441, net89694, net89773,
         net90992, net91003, net91001, net91017, net91147, net91155, net91202,
         net91269, net91311, net91388, net91392, net91526, net99829, net99836,
         net99835, \ML_int[1][15] , net99764, net89357, net88995, net88994,
         net88993, net88992, net88991, net88990, net85898, net85894,
         \ML_int[2][21] , \ML_int[2][17] , \ML_int[1][21] , \ML_int[1][19] ,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100
;

  MUX2_X2 M1_2_10 ( .A(n16), .B(\ML_int[2][6] ), .S(net85895), .Z(B[10]) );
  MUX2_X2 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(net85895), .Z(
        B[8]) );
  MUX2_X2 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(net85895), .Z(
        B[7]) );
  MUX2_X2 M1_2_5 ( .A(\ML_int[2][5] ), .B(\ML_int[2][1] ), .S(net85895), .Z(
        B[5]) );
  MUX2_X2 M1_0_20 ( .A(A[20]), .B(A[19]), .S(net88600), .Z(\ML_int[1][20] ) );
  MUX2_X2 M1_0_11 ( .A(A[11]), .B(A[10]), .S(net85903), .Z(\ML_int[1][11] ) );
  MUX2_X2 M1_0_9 ( .A(A[9]), .B(A[8]), .S(net88672), .Z(\ML_int[1][9] ) );
  MUX2_X2 M1_0_14 ( .A(A[14]), .B(A[13]), .S(net88672), .Z(\ML_int[1][14] ) );
  MUX2_X2 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S(net85899), 
        .Z(\ML_int[2][21] ) );
  MUX2_X2 M0_0_0 ( .A(A[0]), .B(1'b0), .S(net88672), .Z(\ML_int[1][0] ) );
  NAND2_X2 U3 ( .A1(net99764), .A2(net88990), .ZN(net88991) );
  NAND2_X2 U4 ( .A1(A[19]), .A2(net89357), .ZN(n10) );
  NAND2_X2 U5 ( .A1(\ML_int[1][5] ), .A2(net88766), .ZN(n18) );
  NAND2_X4 U6 ( .A1(n77), .A2(n78), .ZN(n1) );
  NAND2_X1 U7 ( .A1(n77), .A2(n78), .ZN(n16) );
  NAND2_X1 U8 ( .A1(\ML_int[2][11] ), .A2(net89236), .ZN(n53) );
  NAND2_X2 U9 ( .A1(n63), .A2(n64), .ZN(n2) );
  NAND2_X2 U10 ( .A1(A[11]), .A2(n4), .ZN(n64) );
  NAND2_X2 U11 ( .A1(\ML_int[1][7] ), .A2(net89012), .ZN(n27) );
  NAND2_X1 U12 ( .A1(A[21]), .A2(net89257), .ZN(n11) );
  NAND2_X1 U13 ( .A1(\ML_int[1][20] ), .A2(net91392), .ZN(n83) );
  NAND2_X2 U14 ( .A1(\ML_int[1][6] ), .A2(net89046), .ZN(n61) );
  NAND2_X2 U15 ( .A1(n24), .A2(n25), .ZN(\ML_int[2][14] ) );
  INV_X4 U16 ( .A(net88600), .ZN(n3) );
  INV_X4 U17 ( .A(n3), .ZN(n4) );
  NAND2_X2 U18 ( .A1(A[3]), .A2(net85903), .ZN(n62) );
  INV_X1 U19 ( .A(n76), .ZN(n5) );
  INV_X4 U20 ( .A(net85895), .ZN(net88351) );
  INV_X4 U21 ( .A(net88351), .ZN(net88861) );
  NAND2_X4 U22 ( .A1(net88458), .A2(n2), .ZN(n96) );
  NOR2_X2 U23 ( .A1(n40), .A2(net85898), .ZN(n8) );
  INV_X1 U24 ( .A(A[9]), .ZN(n46) );
  NAND2_X2 U25 ( .A1(\ML_int[1][10] ), .A2(net85899), .ZN(n97) );
  NAND2_X2 U26 ( .A1(\ML_int[1][6] ), .A2(net85899), .ZN(n57) );
  NAND2_X2 U27 ( .A1(n33), .A2(n34), .ZN(\ML_int[2][13] ) );
  NAND2_X2 U28 ( .A1(n22), .A2(n23), .ZN(\ML_int[2][9] ) );
  INV_X1 U29 ( .A(A[0]), .ZN(n42) );
  INV_X1 U30 ( .A(A[1]), .ZN(n41) );
  INV_X8 U31 ( .A(net85895), .ZN(net91311) );
  NAND2_X2 U32 ( .A1(n60), .A2(n61), .ZN(\ML_int[2][6] ) );
  NAND2_X2 U33 ( .A1(\ML_int[1][4] ), .A2(net89354), .ZN(n60) );
  NAND2_X2 U34 ( .A1(\ML_int[2][8] ), .A2(net88861), .ZN(n87) );
  NAND2_X2 U35 ( .A1(net88351), .A2(n17), .ZN(n88) );
  NAND2_X2 U36 ( .A1(\ML_int[2][7] ), .A2(net88861), .ZN(n52) );
  NAND2_X2 U37 ( .A1(n70), .A2(n69), .ZN(B[13]) );
  NAND2_X2 U38 ( .A1(net88600), .A2(A[18]), .ZN(net89773) );
  INV_X8 U39 ( .A(net88600), .ZN(net89257) );
  INV_X8 U40 ( .A(n13), .ZN(net85903) );
  NAND2_X2 U41 ( .A1(n31), .A2(n32), .ZN(\ML_int[2][18] ) );
  NAND2_X4 U42 ( .A1(n48), .A2(n49), .ZN(B[15]) );
  NAND2_X4 U43 ( .A1(\ML_int[1][3] ), .A2(net89007), .ZN(n75) );
  NAND2_X2 U44 ( .A1(\ML_int[1][3] ), .A2(net85899), .ZN(n19) );
  NAND2_X1 U45 ( .A1(A[20]), .A2(net85903), .ZN(n12) );
  NAND2_X4 U46 ( .A1(n36), .A2(n37), .ZN(B[19]) );
  NAND2_X2 U47 ( .A1(\ML_int[2][15] ), .A2(net85895), .ZN(n37) );
  NAND2_X2 U48 ( .A1(\ML_int[1][8] ), .A2(net89441), .ZN(n56) );
  NAND2_X4 U49 ( .A1(n73), .A2(net89040), .ZN(B[17]) );
  NAND2_X4 U50 ( .A1(\ML_int[2][17] ), .A2(net88778), .ZN(net89040) );
  NAND2_X4 U51 ( .A1(n95), .A2(n94), .ZN(\ML_int[2][16] ) );
  MUX2_X2 U52 ( .A(A[18]), .B(A[17]), .S(net88600), .Z(n6) );
  NAND2_X4 U53 ( .A1(n47), .A2(net88908), .ZN(n82) );
  NAND2_X2 U54 ( .A1(\ML_int[1][15] ), .A2(net85899), .ZN(net88992) );
  NAND2_X2 U55 ( .A1(\ML_int[1][15] ), .A2(net88766), .ZN(net88783) );
  NAND2_X2 U56 ( .A1(net99836), .A2(net89050), .ZN(n72) );
  INV_X4 U57 ( .A(net99835), .ZN(net99836) );
  NAND2_X4 U58 ( .A1(n17), .A2(net85895), .ZN(n29) );
  NAND2_X4 U59 ( .A1(n97), .A2(n96), .ZN(n17) );
  NOR2_X4 U60 ( .A1(n100), .A2(net85899), .ZN(\ML_int[2][0] ) );
  INV_X4 U61 ( .A(\ML_int[1][0] ), .ZN(n100) );
  INV_X2 U62 ( .A(net85899), .ZN(net89046) );
  OAI21_X1 U63 ( .B1(n5), .B2(n9), .A(net85894), .ZN(n7) );
  INV_X2 U64 ( .A(n7), .ZN(B[3]) );
  INV_X4 U65 ( .A(n8), .ZN(n76) );
  INV_X1 U66 ( .A(n75), .ZN(n9) );
  AND2_X2 U67 ( .A1(\ML_int[2][1] ), .A2(net85894), .ZN(B[1]) );
  NAND2_X4 U68 ( .A1(net88994), .A2(net88995), .ZN(B[21]) );
  NAND2_X4 U69 ( .A1(\ML_int[2][17] ), .A2(net85895), .ZN(net88995) );
  INV_X32 U70 ( .A(net85894), .ZN(net85895) );
  INV_X8 U71 ( .A(SH[2]), .ZN(net85894) );
  NAND2_X4 U72 ( .A1(\ML_int[2][21] ), .A2(net88993), .ZN(net88994) );
  INV_X1 U73 ( .A(net85895), .ZN(net88993) );
  INV_X32 U74 ( .A(net85898), .ZN(net85899) );
  INV_X8 U75 ( .A(SH[1]), .ZN(net85898) );
  NAND2_X2 U76 ( .A1(n12), .A2(n11), .ZN(\ML_int[1][21] ) );
  INV_X2 U77 ( .A(net89257), .ZN(net91526) );
  NAND2_X1 U78 ( .A1(A[13]), .A2(net89257), .ZN(net91001) );
  INV_X16 U79 ( .A(n13), .ZN(net88600) );
  INV_X16 U80 ( .A(SH[0]), .ZN(n13) );
  INV_X16 U81 ( .A(n13), .ZN(net88672) );
  NAND2_X4 U82 ( .A1(net88991), .A2(net88992), .ZN(\ML_int[2][17] ) );
  INV_X1 U83 ( .A(net85899), .ZN(net88990) );
  NAND2_X4 U84 ( .A1(net89773), .A2(n10), .ZN(\ML_int[1][19] ) );
  INV_X1 U85 ( .A(\ML_int[1][19] ), .ZN(net99835) );
  INV_X4 U86 ( .A(net85903), .ZN(net89357) );
  NAND2_X1 U87 ( .A1(A[2]), .A2(net89357), .ZN(net91147) );
  NAND2_X1 U88 ( .A1(A[4]), .A2(net89357), .ZN(net89358) );
  MUX2_X2 U89 ( .A(A[17]), .B(A[16]), .S(net88672), .Z(net99764) );
  NAND2_X2 U90 ( .A1(net85899), .A2(net99764), .ZN(net89052) );
  MUX2_X2 U91 ( .A(A[16]), .B(A[15]), .S(net88600), .Z(net99829) );
  NAND2_X4 U92 ( .A1(n14), .A2(n15), .ZN(\ML_int[1][15] ) );
  NAND2_X1 U93 ( .A1(A[14]), .A2(net88600), .ZN(n15) );
  NAND2_X2 U94 ( .A1(A[15]), .A2(net89257), .ZN(n14) );
  NAND2_X1 U95 ( .A1(A[3]), .A2(net89257), .ZN(net89170) );
  NAND2_X4 U96 ( .A1(\ML_int[2][13] ), .A2(net88980), .ZN(n73) );
  NAND2_X2 U97 ( .A1(\ML_int[2][14] ), .A2(net89420), .ZN(n58) );
  INV_X1 U98 ( .A(net85899), .ZN(net88908) );
  NAND2_X4 U99 ( .A1(\ML_int[2][14] ), .A2(net88980), .ZN(n79) );
  NAND2_X4 U100 ( .A1(n1), .A2(net85895), .ZN(n59) );
  NAND2_X4 U101 ( .A1(\ML_int[2][11] ), .A2(net88980), .ZN(n48) );
  NAND2_X4 U102 ( .A1(n81), .A2(n82), .ZN(\ML_int[2][11] ) );
  INV_X4 U103 ( .A(net85895), .ZN(net88778) );
  NAND2_X4 U104 ( .A1(n59), .A2(n58), .ZN(B[14]) );
  INV_X1 U105 ( .A(A[10]), .ZN(n45) );
  NAND2_X2 U106 ( .A1(net85899), .A2(net99829), .ZN(n32) );
  NAND2_X2 U107 ( .A1(n85), .A2(n86), .ZN(\ML_int[1][6] ) );
  NAND2_X1 U108 ( .A1(A[8]), .A2(net89257), .ZN(n54) );
  NAND2_X2 U109 ( .A1(n62), .A2(net89358), .ZN(\ML_int[1][4] ) );
  NAND2_X1 U110 ( .A1(A[2]), .A2(net85903), .ZN(n71) );
  NAND2_X2 U111 ( .A1(n54), .A2(n55), .ZN(\ML_int[1][8] ) );
  NAND2_X2 U112 ( .A1(n18), .A2(n19), .ZN(\ML_int[2][5] ) );
  NAND2_X2 U113 ( .A1(\ML_int[2][5] ), .A2(net85895), .ZN(n51) );
  NAND2_X1 U114 ( .A1(A[4]), .A2(net88600), .ZN(n68) );
  INV_X2 U115 ( .A(net88908), .ZN(net88921) );
  INV_X2 U116 ( .A(net89046), .ZN(net89354) );
  INV_X2 U117 ( .A(net89012), .ZN(net91202) );
  NAND2_X4 U118 ( .A1(\ML_int[2][19] ), .A2(net91003), .ZN(n36) );
  NAND2_X2 U119 ( .A1(\ML_int[2][15] ), .A2(net88351), .ZN(n49) );
  NAND2_X4 U120 ( .A1(n91), .A2(net88783), .ZN(\ML_int[2][15] ) );
  NAND2_X2 U121 ( .A1(\ML_int[1][11] ), .A2(net85899), .ZN(n34) );
  NAND2_X2 U122 ( .A1(\ML_int[1][9] ), .A2(net88921), .ZN(n81) );
  NAND2_X2 U123 ( .A1(n74), .A2(net91392), .ZN(n20) );
  NAND2_X1 U124 ( .A1(\ML_int[1][0] ), .A2(net85899), .ZN(n21) );
  NAND2_X2 U125 ( .A1(n20), .A2(n21), .ZN(\ML_int[2][2] ) );
  INV_X1 U126 ( .A(net85899), .ZN(net91392) );
  NOR2_X1 U127 ( .A1(net85895), .A2(n99), .ZN(B[0]) );
  NOR2_X1 U128 ( .A1(n98), .A2(net85895), .ZN(B[2]) );
  NAND2_X2 U129 ( .A1(\ML_int[1][9] ), .A2(net91388), .ZN(n22) );
  NAND2_X2 U130 ( .A1(\ML_int[1][7] ), .A2(net85899), .ZN(n23) );
  INV_X1 U131 ( .A(net85899), .ZN(net91388) );
  NAND2_X2 U132 ( .A1(\ML_int[2][9] ), .A2(net85895), .ZN(n70) );
  NAND2_X2 U133 ( .A1(\ML_int[2][9] ), .A2(net89694), .ZN(n50) );
  NAND2_X1 U134 ( .A1(A[6]), .A2(n4), .ZN(n93) );
  NAND2_X1 U135 ( .A1(\ML_int[1][12] ), .A2(net85899), .ZN(n25) );
  NAND2_X2 U136 ( .A1(\ML_int[1][14] ), .A2(net91269), .ZN(n24) );
  NAND2_X2 U137 ( .A1(n6), .A2(net91017), .ZN(n31) );
  NAND2_X2 U138 ( .A1(\ML_int[1][14] ), .A2(net91202), .ZN(n94) );
  MUX2_X2 U139 ( .A(\ML_int[2][0] ), .B(\ML_int[2][4] ), .S(net91311), .Z(B[4]) );
  NAND2_X4 U140 ( .A1(\ML_int[2][16] ), .A2(net91155), .ZN(n28) );
  NAND2_X1 U141 ( .A1(A[7]), .A2(net89257), .ZN(n92) );
  INV_X1 U142 ( .A(net85899), .ZN(net91269) );
  NAND2_X2 U143 ( .A1(\ML_int[2][16] ), .A2(net85895), .ZN(n39) );
  NAND2_X4 U144 ( .A1(\ML_int[2][18] ), .A2(net88778), .ZN(n80) );
  NAND2_X4 U145 ( .A1(n80), .A2(n79), .ZN(B[18]) );
  NAND2_X1 U146 ( .A1(\ML_int[1][5] ), .A2(net91202), .ZN(n26) );
  NAND2_X2 U147 ( .A1(n26), .A2(n27), .ZN(\ML_int[2][7] ) );
  NAND2_X2 U148 ( .A1(n92), .A2(n93), .ZN(\ML_int[1][7] ) );
  INV_X1 U149 ( .A(net85899), .ZN(net89012) );
  NAND2_X4 U150 ( .A1(n29), .A2(n28), .ZN(B[16]) );
  INV_X1 U151 ( .A(net85895), .ZN(net91155) );
  NAND2_X1 U152 ( .A1(A[1]), .A2(net88600), .ZN(n30) );
  NAND2_X2 U153 ( .A1(net91147), .A2(n30), .ZN(\ML_int[1][2] ) );
  NAND2_X2 U154 ( .A1(net99829), .A2(net91388), .ZN(n95) );
  NAND2_X1 U155 ( .A1(A[5]), .A2(net88600), .ZN(n86) );
  INV_X1 U156 ( .A(net85899), .ZN(net91017) );
  NAND2_X2 U157 ( .A1(n43), .A2(net91269), .ZN(n33) );
  NAND2_X2 U158 ( .A1(\ML_int[2][13] ), .A2(net89240), .ZN(n69) );
  NAND2_X1 U159 ( .A1(A[12]), .A2(net91526), .ZN(n35) );
  NAND2_X2 U160 ( .A1(net91001), .A2(n35), .ZN(\ML_int[1][13] ) );
  INV_X1 U161 ( .A(net85895), .ZN(net91003) );
  NAND2_X2 U162 ( .A1(\ML_int[1][13] ), .A2(net88921), .ZN(n91) );
  NAND2_X2 U163 ( .A1(\ML_int[2][20] ), .A2(net90992), .ZN(n38) );
  NAND2_X2 U164 ( .A1(n38), .A2(n39), .ZN(B[20]) );
  INV_X1 U165 ( .A(net85895), .ZN(net90992) );
  NAND2_X2 U166 ( .A1(\ML_int[1][2] ), .A2(net85899), .ZN(n66) );
  MUX2_X2 U167 ( .A(n41), .B(n42), .S(net88600), .Z(n40) );
  MUX2_X2 U168 ( .A(A[13]), .B(A[12]), .S(net88600), .Z(n43) );
  MUX2_X2 U169 ( .A(n45), .B(n46), .S(net88672), .Z(n44) );
  INV_X4 U170 ( .A(n44), .ZN(\ML_int[1][10] ) );
  INV_X1 U171 ( .A(\ML_int[2][0] ), .ZN(n99) );
  MUX2_X2 U172 ( .A(A[11]), .B(A[10]), .S(net85903), .Z(n47) );
  NAND2_X2 U173 ( .A1(n75), .A2(n76), .ZN(\ML_int[2][3] ) );
  NAND2_X2 U174 ( .A1(n50), .A2(n51), .ZN(B[9]) );
  INV_X1 U175 ( .A(net85895), .ZN(net89694) );
  NAND2_X1 U176 ( .A1(\ML_int[2][6] ), .A2(net88852), .ZN(n89) );
  NAND2_X2 U177 ( .A1(\ML_int[2][2] ), .A2(net85895), .ZN(n90) );
  NAND2_X4 U178 ( .A1(n52), .A2(n53), .ZN(B[11]) );
  INV_X1 U179 ( .A(net85895), .ZN(net89236) );
  NAND2_X1 U180 ( .A1(A[7]), .A2(net85903), .ZN(n55) );
  NAND2_X4 U181 ( .A1(n56), .A2(n57), .ZN(\ML_int[2][8] ) );
  INV_X1 U182 ( .A(net85899), .ZN(net89441) );
  NAND2_X2 U183 ( .A1(\ML_int[1][8] ), .A2(net85899), .ZN(n78) );
  INV_X1 U184 ( .A(net85895), .ZN(net89420) );
  INV_X2 U185 ( .A(\ML_int[2][2] ), .ZN(n98) );
  NAND2_X4 U186 ( .A1(\ML_int[1][4] ), .A2(net89339), .ZN(n65) );
  NAND2_X2 U187 ( .A1(n6), .A2(net85899), .ZN(n84) );
  NAND2_X2 U188 ( .A1(A[12]), .A2(net89357), .ZN(n63) );
  NAND2_X2 U189 ( .A1(n63), .A2(n64), .ZN(\ML_int[1][12] ) );
  NAND2_X2 U190 ( .A1(n65), .A2(n66), .ZN(\ML_int[2][4] ) );
  INV_X1 U191 ( .A(net85899), .ZN(net89339) );
  NAND2_X1 U192 ( .A1(A[5]), .A2(net89257), .ZN(n67) );
  NAND2_X2 U193 ( .A1(n67), .A2(n68), .ZN(\ML_int[1][5] ) );
  NOR2_X2 U194 ( .A1(net85899), .A2(n40), .ZN(\ML_int[2][1] ) );
  INV_X1 U195 ( .A(net85895), .ZN(net89240) );
  NAND2_X2 U196 ( .A1(net89170), .A2(n71), .ZN(\ML_int[1][3] ) );
  NAND2_X2 U197 ( .A1(n72), .A2(net89052), .ZN(\ML_int[2][19] ) );
  INV_X1 U198 ( .A(net85899), .ZN(net89050) );
  MUX2_X2 U199 ( .A(A[2]), .B(A[1]), .S(net85903), .Z(n74) );
  INV_X1 U200 ( .A(net85899), .ZN(net89007) );
  NAND2_X2 U201 ( .A1(\ML_int[1][10] ), .A2(net88998), .ZN(n77) );
  INV_X1 U202 ( .A(net85899), .ZN(net88998) );
  INV_X4 U203 ( .A(net88778), .ZN(net88980) );
  NAND2_X2 U204 ( .A1(n83), .A2(n84), .ZN(\ML_int[2][20] ) );
  NAND2_X1 U205 ( .A1(A[6]), .A2(net89257), .ZN(n85) );
  NAND2_X4 U206 ( .A1(n87), .A2(n88), .ZN(B[12]) );
  NAND2_X2 U207 ( .A1(n90), .A2(n89), .ZN(B[6]) );
  INV_X1 U208 ( .A(net85895), .ZN(net88852) );
  INV_X1 U209 ( .A(net85899), .ZN(net88766) );
  INV_X1 U210 ( .A(net85899), .ZN(net88458) );
endmodule


module fpu_DW01_sub_23 ( A, B, CI, DIFF, CO );
  input [6:0] A;
  input [6:0] B;
  output [6:0] DIFF;
  input CI;
  output CO;
  wire   net64864, net64862, net64843, net64841, net64840, net85706, net89571,
         net89670, net89739, net64871, net90964, net90963, net90960, net90954,
         net90950, net90938, net90300, net64870, net64847, net64863, net64848,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;
  assign net85706 = A[1];

  OAI21_X2 U3 ( .B1(net64840), .B2(net64841), .A(net64864), .ZN(n17) );
  INV_X4 U4 ( .A(n23), .ZN(n19) );
  NAND2_X2 U5 ( .A1(net89739), .A2(net64843), .ZN(net64864) );
  NAND2_X1 U6 ( .A1(n1), .A2(n4), .ZN(net90938) );
  INV_X1 U7 ( .A(n9), .ZN(net89739) );
  INV_X8 U8 ( .A(A[2]), .ZN(net64843) );
  NAND2_X1 U9 ( .A1(net89571), .A2(n8), .ZN(net64841) );
  INV_X4 U10 ( .A(net85706), .ZN(n1) );
  NOR2_X4 U11 ( .A1(n2), .A2(n1), .ZN(n3) );
  AOI21_X4 U12 ( .B1(net64863), .B2(net90300), .A(n3), .ZN(net64870) );
  NAND2_X2 U13 ( .A1(n2), .A2(n1), .ZN(net64863) );
  INV_X8 U14 ( .A(net64848), .ZN(n2) );
  BUF_X32 U15 ( .A(n2), .Z(n4) );
  INV_X8 U16 ( .A(B[1]), .ZN(net64848) );
  NAND2_X1 U17 ( .A1(net85706), .A2(net64848), .ZN(net89571) );
  NOR2_X1 U18 ( .A1(net85706), .A2(net64848), .ZN(net64847) );
  XNOR2_X2 U19 ( .A(B[1]), .B(net85706), .ZN(net90964) );
  XNOR2_X2 U20 ( .A(net64870), .B(net64871), .ZN(DIFF[2]) );
  INV_X8 U21 ( .A(net90954), .ZN(net90300) );
  NAND3_X1 U22 ( .A1(net90938), .A2(net90300), .A3(net64864), .ZN(net64862) );
  INV_X4 U23 ( .A(net90950), .ZN(net90954) );
  NOR2_X2 U24 ( .A1(net64847), .A2(net90954), .ZN(net64840) );
  XNOR2_X2 U25 ( .A(net90954), .B(net90964), .ZN(DIFF[1]) );
  NAND2_X4 U26 ( .A1(B[0]), .A2(n5), .ZN(net90950) );
  NAND2_X2 U27 ( .A1(net90950), .A2(net90963), .ZN(DIFF[0]) );
  INV_X4 U28 ( .A(A[0]), .ZN(n5) );
  INV_X4 U29 ( .A(B[0]), .ZN(net90960) );
  NAND2_X2 U30 ( .A1(A[0]), .A2(net90960), .ZN(net90963) );
  NOR2_X4 U31 ( .A1(n7), .A2(n6), .ZN(net64871) );
  NOR2_X4 U32 ( .A1(n9), .A2(A[2]), .ZN(n6) );
  INV_X8 U33 ( .A(B[2]), .ZN(n9) );
  NAND2_X4 U34 ( .A1(n9), .A2(A[2]), .ZN(n8) );
  INV_X8 U35 ( .A(n8), .ZN(n7) );
  NOR2_X2 U36 ( .A1(n22), .A2(B[4]), .ZN(n10) );
  INV_X4 U37 ( .A(n10), .ZN(n21) );
  NAND2_X4 U38 ( .A1(n24), .A2(n25), .ZN(n16) );
  INV_X4 U39 ( .A(n15), .ZN(n11) );
  NAND2_X1 U40 ( .A1(n22), .A2(B[4]), .ZN(n25) );
  INV_X4 U41 ( .A(B[3]), .ZN(n35) );
  NAND2_X1 U42 ( .A1(n29), .A2(n24), .ZN(n28) );
  INV_X1 U43 ( .A(net89571), .ZN(net89670) );
  NAND2_X2 U44 ( .A1(n15), .A2(A[5]), .ZN(n13) );
  NAND2_X4 U45 ( .A1(n11), .A2(n12), .ZN(n14) );
  NAND2_X4 U46 ( .A1(n14), .A2(n13), .ZN(DIFF[5]) );
  INV_X4 U47 ( .A(A[5]), .ZN(n12) );
  AOI21_X1 U48 ( .B1(n34), .B2(net89670), .A(n7), .ZN(n33) );
  NAND2_X1 U49 ( .A1(n25), .A2(n21), .ZN(n26) );
  NAND2_X4 U50 ( .A1(n35), .A2(A[3]), .ZN(n23) );
  NAND2_X2 U51 ( .A1(B[4]), .A2(n22), .ZN(n20) );
  NAND2_X1 U52 ( .A1(n24), .A2(n23), .ZN(n31) );
  NAND2_X1 U53 ( .A1(n28), .A2(n23), .ZN(n27) );
  NAND2_X1 U54 ( .A1(net64843), .A2(net89739), .ZN(n34) );
  OAI21_X4 U55 ( .B1(n17), .B2(n16), .A(n18), .ZN(n15) );
  AOI21_X4 U56 ( .B1(n19), .B2(n20), .A(n10), .ZN(n18) );
  XNOR2_X2 U57 ( .A(n26), .B(n27), .ZN(DIFF[4]) );
  INV_X4 U58 ( .A(A[4]), .ZN(n22) );
  INV_X4 U59 ( .A(n30), .ZN(DIFF[3]) );
  XNOR2_X2 U60 ( .A(n31), .B(n32), .ZN(n30) );
  INV_X4 U61 ( .A(n29), .ZN(n32) );
  NAND2_X2 U62 ( .A1(n33), .A2(net64862), .ZN(n29) );
  NAND2_X2 U63 ( .A1(n36), .A2(B[3]), .ZN(n24) );
  INV_X4 U64 ( .A(A[3]), .ZN(n36) );
endmodule


module fpu_DW_rash_11 ( A, DATA_TC, SH, SH_TC, B );
  input [13:0] A;
  input [3:0] SH;
  output [13:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140;

  NAND2_X2 U3 ( .A1(A[9]), .A2(n130), .ZN(n129) );
  NAND2_X2 U4 ( .A1(A[8]), .A2(n130), .ZN(n103) );
  NAND2_X2 U5 ( .A1(n130), .A2(A[4]), .ZN(n99) );
  NAND2_X2 U6 ( .A1(A[11]), .A2(n130), .ZN(n112) );
  NAND2_X2 U7 ( .A1(A[7]), .A2(n130), .ZN(n118) );
  INV_X8 U8 ( .A(n131), .ZN(n130) );
  NAND2_X4 U9 ( .A1(A[10]), .A2(n69), .ZN(n89) );
  NAND2_X4 U10 ( .A1(n34), .A2(n35), .ZN(B[5]) );
  NOR2_X2 U11 ( .A1(n73), .A2(n74), .ZN(n63) );
  NOR2_X1 U12 ( .A1(n32), .A2(n14), .ZN(n53) );
  NOR2_X1 U13 ( .A1(n15), .A2(n12), .ZN(n132) );
  NAND2_X2 U14 ( .A1(A[5]), .A2(n130), .ZN(n137) );
  NOR2_X2 U15 ( .A1(n21), .A2(n12), .ZN(n41) );
  NOR2_X1 U16 ( .A1(n20), .A2(n14), .ZN(n17) );
  NOR2_X1 U17 ( .A1(n19), .A2(n12), .ZN(n18) );
  NOR3_X2 U18 ( .A1(n59), .A2(SH[2]), .A3(n2), .ZN(n58) );
  NOR2_X2 U19 ( .A1(n9), .A2(n10), .ZN(n6) );
  NOR2_X1 U20 ( .A1(n13), .A2(n14), .ZN(n9) );
  NOR2_X1 U21 ( .A1(n13), .A2(n12), .ZN(n72) );
  NOR2_X1 U22 ( .A1(n5), .A2(n12), .ZN(n54) );
  NOR2_X2 U23 ( .A1(n132), .A2(n133), .ZN(n123) );
  INV_X4 U24 ( .A(SH[3]), .ZN(n134) );
  AND2_X2 U25 ( .A1(SH[0]), .A2(SH[1]), .ZN(n1) );
  AND2_X2 U26 ( .A1(n27), .A2(n8), .ZN(n2) );
  OR2_X4 U27 ( .A1(n19), .A2(n14), .ZN(n3) );
  AND2_X2 U28 ( .A1(A[7]), .A2(n69), .ZN(n4) );
  AND3_X4 U29 ( .A1(n121), .A2(n122), .A3(n120), .ZN(n5) );
  NOR2_X2 U30 ( .A1(n20), .A2(n12), .ZN(B[12]) );
  NOR2_X1 U31 ( .A1(n33), .A2(n12), .ZN(B[10]) );
  NAND2_X4 U32 ( .A1(n36), .A2(n64), .ZN(n35) );
  OAI21_X2 U33 ( .B1(n7), .B2(SH[3]), .A(n37), .ZN(n36) );
  NOR2_X2 U34 ( .A1(n11), .A2(n44), .ZN(n59) );
  NOR2_X1 U35 ( .A1(n11), .A2(n14), .ZN(n38) );
  NOR2_X1 U36 ( .A1(n11), .A2(n12), .ZN(n10) );
  AND4_X4 U37 ( .A1(n75), .A2(n76), .A3(n77), .A4(n78), .ZN(n11) );
  NAND2_X1 U38 ( .A1(n27), .A2(n28), .ZN(n22) );
  NAND3_X2 U39 ( .A1(n45), .A2(n46), .A3(n47), .ZN(B[3]) );
  INV_X1 U40 ( .A(SH[0]), .ZN(n140) );
  NAND3_X2 U41 ( .A1(n89), .A2(n90), .A3(n91), .ZN(n88) );
  NAND3_X2 U42 ( .A1(n107), .A2(n108), .A3(n106), .ZN(n26) );
  NAND2_X2 U43 ( .A1(A[6]), .A2(n130), .ZN(n84) );
  NOR2_X4 U44 ( .A1(SH[1]), .A2(SH[0]), .ZN(n24) );
  NAND2_X2 U45 ( .A1(A[5]), .A2(n24), .ZN(n82) );
  NAND2_X2 U46 ( .A1(A[12]), .A2(n24), .ZN(n87) );
  NOR2_X2 U47 ( .A1(SH[2]), .A2(SH[3]), .ZN(n27) );
  NOR2_X1 U48 ( .A1(n21), .A2(n14), .ZN(n133) );
  AND4_X4 U49 ( .A1(n135), .A2(n136), .A3(n137), .A4(n138), .ZN(n21) );
  NAND2_X1 U50 ( .A1(n130), .A2(A[3]), .ZN(n121) );
  INV_X2 U51 ( .A(SH[1]), .ZN(n70) );
  NAND2_X1 U52 ( .A1(n87), .A2(n86), .ZN(n127) );
  NOR2_X2 U53 ( .A1(n7), .A2(SH[3]), .ZN(n65) );
  INV_X1 U54 ( .A(n24), .ZN(n73) );
  NAND2_X2 U55 ( .A1(SH[0]), .A2(n70), .ZN(n131) );
  NAND2_X1 U56 ( .A1(A[6]), .A2(n24), .ZN(n116) );
  NAND2_X1 U57 ( .A1(A[10]), .A2(n24), .ZN(n110) );
  NAND2_X1 U58 ( .A1(A[3]), .A2(n24), .ZN(n97) );
  NAND2_X1 U59 ( .A1(A[7]), .A2(n24), .ZN(n101) );
  NAND2_X1 U60 ( .A1(A[9]), .A2(n24), .ZN(n75) );
  NAND2_X1 U61 ( .A1(A[4]), .A2(n24), .ZN(n135) );
  NAND2_X4 U62 ( .A1(A[8]), .A2(n24), .ZN(n95) );
  NAND3_X1 U63 ( .A1(SH[1]), .A2(SH[0]), .A3(A[8]), .ZN(n83) );
  NAND3_X1 U64 ( .A1(A[13]), .A2(n70), .A3(SH[0]), .ZN(n86) );
  INV_X4 U65 ( .A(n6), .ZN(B[9]) );
  NAND2_X2 U66 ( .A1(n66), .A2(n67), .ZN(n8) );
  NAND2_X2 U67 ( .A1(n86), .A2(n87), .ZN(n43) );
  INV_X4 U68 ( .A(n96), .ZN(B[11]) );
  NAND2_X2 U69 ( .A1(n51), .A2(n52), .ZN(B[2]) );
  NAND3_X4 U70 ( .A1(n3), .A2(n40), .A3(n39), .ZN(B[4]) );
  NAND2_X2 U71 ( .A1(n22), .A2(n23), .ZN(B[7]) );
  INV_X4 U72 ( .A(n29), .ZN(B[6]) );
  INV_X4 U73 ( .A(n16), .ZN(B[8]) );
  INV_X4 U74 ( .A(n37), .ZN(n60) );
  NAND2_X2 U75 ( .A1(n1), .A2(A[3]), .ZN(n15) );
  INV_X4 U76 ( .A(n72), .ZN(n71) );
  INV_X4 U77 ( .A(n48), .ZN(n47) );
  NAND2_X4 U78 ( .A1(SH[2]), .A2(n134), .ZN(n14) );
  INV_X8 U79 ( .A(n139), .ZN(n69) );
  NAND2_X4 U80 ( .A1(SH[1]), .A2(SH[0]), .ZN(n68) );
  INV_X8 U81 ( .A(n27), .ZN(n12) );
  NOR2_X4 U82 ( .A1(n17), .A2(n18), .ZN(n16) );
  NAND2_X2 U83 ( .A1(n25), .A2(n26), .ZN(n23) );
  INV_X4 U84 ( .A(n14), .ZN(n25) );
  NOR2_X4 U85 ( .A1(n30), .A2(n31), .ZN(n29) );
  NOR2_X4 U86 ( .A1(n32), .A2(n12), .ZN(n31) );
  NOR2_X4 U87 ( .A1(n33), .A2(n14), .ZN(n30) );
  INV_X4 U88 ( .A(n38), .ZN(n34) );
  INV_X4 U89 ( .A(n41), .ZN(n40) );
  NAND2_X2 U90 ( .A1(n42), .A2(n43), .ZN(n39) );
  INV_X4 U91 ( .A(n44), .ZN(n42) );
  NOR2_X4 U92 ( .A1(n49), .A2(n44), .ZN(n48) );
  INV_X4 U93 ( .A(n26), .ZN(n49) );
  NAND2_X2 U94 ( .A1(n25), .A2(n28), .ZN(n46) );
  NAND2_X2 U95 ( .A1(n27), .A2(n50), .ZN(n45) );
  NOR2_X4 U96 ( .A1(n53), .A2(n54), .ZN(n52) );
  NAND2_X2 U97 ( .A1(n42), .A2(n55), .ZN(n51) );
  AOI21_X4 U98 ( .B1(n56), .B2(n57), .A(n58), .ZN(B[1]) );
  NOR2_X4 U99 ( .A1(n59), .A2(n60), .ZN(n57) );
  NAND2_X2 U100 ( .A1(n62), .A2(n63), .ZN(n37) );
  NAND2_X2 U101 ( .A1(n62), .A2(n64), .ZN(n44) );
  NOR2_X4 U102 ( .A1(n2), .A2(n65), .ZN(n56) );
  NAND2_X2 U103 ( .A1(A[4]), .A2(n61), .ZN(n67) );
  INV_X4 U104 ( .A(n68), .ZN(n61) );
  NAND2_X2 U105 ( .A1(A[3]), .A2(n69), .ZN(n66) );
  INV_X4 U106 ( .A(n71), .ZN(B[13]) );
  INV_X4 U107 ( .A(n63), .ZN(n13) );
  INV_X4 U108 ( .A(A[13]), .ZN(n74) );
  NAND2_X2 U109 ( .A1(A[11]), .A2(n69), .ZN(n78) );
  NAND2_X2 U110 ( .A1(A[10]), .A2(n130), .ZN(n77) );
  NAND2_X2 U111 ( .A1(A[12]), .A2(n79), .ZN(n76) );
  INV_X4 U112 ( .A(n68), .ZN(n79) );
  NOR3_X4 U113 ( .A1(n4), .A2(n80), .A3(n81), .ZN(n7) );
  NAND2_X2 U114 ( .A1(n82), .A2(n83), .ZN(n81) );
  INV_X4 U115 ( .A(n84), .ZN(n80) );
  INV_X4 U116 ( .A(n43), .ZN(n20) );
  INV_X4 U117 ( .A(n88), .ZN(n19) );
  NOR2_X4 U118 ( .A1(n92), .A2(n93), .ZN(n91) );
  NOR2_X4 U119 ( .A1(n68), .A2(n94), .ZN(n93) );
  INV_X4 U120 ( .A(A[11]), .ZN(n94) );
  INV_X4 U121 ( .A(n95), .ZN(n92) );
  NAND2_X2 U122 ( .A1(A[9]), .A2(n130), .ZN(n90) );
  NAND4_X2 U123 ( .A1(n97), .A2(n98), .A3(n99), .A4(n100), .ZN(n50) );
  NAND2_X2 U124 ( .A1(A[5]), .A2(n69), .ZN(n100) );
  NAND2_X2 U125 ( .A1(A[6]), .A2(n61), .ZN(n98) );
  NAND4_X2 U126 ( .A1(n101), .A2(n102), .A3(n103), .A4(n104), .ZN(n28) );
  NAND2_X2 U127 ( .A1(A[9]), .A2(n69), .ZN(n104) );
  NAND2_X2 U128 ( .A1(A[10]), .A2(n105), .ZN(n102) );
  INV_X4 U129 ( .A(n68), .ZN(n105) );
  NAND2_X2 U130 ( .A1(n27), .A2(n26), .ZN(n96) );
  NAND2_X2 U131 ( .A1(A[13]), .A2(n69), .ZN(n108) );
  NAND2_X2 U132 ( .A1(A[12]), .A2(n130), .ZN(n107) );
  NAND2_X2 U133 ( .A1(A[11]), .A2(n24), .ZN(n106) );
  INV_X4 U134 ( .A(n55), .ZN(n33) );
  NAND4_X2 U135 ( .A1(n110), .A2(n111), .A3(n112), .A4(n113), .ZN(n55) );
  NAND2_X2 U136 ( .A1(A[12]), .A2(n69), .ZN(n113) );
  NAND2_X2 U137 ( .A1(A[13]), .A2(n114), .ZN(n111) );
  INV_X4 U138 ( .A(n68), .ZN(n114) );
  INV_X4 U139 ( .A(n115), .ZN(n32) );
  NAND4_X2 U140 ( .A1(n116), .A2(n117), .A3(n118), .A4(n119), .ZN(n115) );
  NAND2_X2 U141 ( .A1(A[8]), .A2(n69), .ZN(n119) );
  NAND2_X2 U142 ( .A1(A[9]), .A2(n61), .ZN(n117) );
  INV_X4 U143 ( .A(SH[2]), .ZN(n64) );
  NAND2_X2 U144 ( .A1(A[4]), .A2(n69), .ZN(n122) );
  NAND2_X2 U145 ( .A1(A[5]), .A2(n114), .ZN(n120) );
  NAND2_X2 U146 ( .A1(n123), .A2(n124), .ZN(B[0]) );
  NAND2_X2 U147 ( .A1(n125), .A2(n62), .ZN(n124) );
  INV_X4 U148 ( .A(n134), .ZN(n62) );
  MUX2_X2 U149 ( .A(n126), .B(n127), .S(SH[2]), .Z(n125) );
  NAND4_X2 U150 ( .A1(n128), .A2(n129), .A3(n89), .A4(n95), .ZN(n126) );
  NAND2_X2 U151 ( .A1(A[11]), .A2(n105), .ZN(n128) );
  NAND2_X2 U152 ( .A1(A[6]), .A2(n69), .ZN(n138) );
  NAND2_X2 U153 ( .A1(SH[1]), .A2(n140), .ZN(n139) );
  NAND2_X2 U154 ( .A1(A[7]), .A2(n79), .ZN(n136) );
endmodule


module fpu ( clk, rmode, fpu_op, opa, opb, out, inf, snan, qnan, ine, overflow, 
        underflow, zero, div_by_zero );
  input [1:0] rmode;
  input [2:0] fpu_op;
  input [15:0] opa;
  input [15:0] opb;
  output [15:0] out;
  input clk;
  output inf, snan, qnan, ine, overflow, underflow, zero, div_by_zero;
  wire   snan_d, opa_nan, opb_nan, opa_00, opb_00, opa_inf, opb_inf, opa_dn,
         opb_dn, sign_fasu, nan_sign_d, result_zero_sign_d, fasu_op,
         sign_fasu_r, sign_mul, sign_exe, inf_mul, sign_mul_r, sign_exe_r, N34,
         N44, N56, N65, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77,
         N96, N97, N98, N99, N100, N106, N110, N111, N112, N113, N114, N115,
         N116, \fract_i2f[7] , N138, N139, N140, N141, N150, N151, N179, N180,
         N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191,
         N192, N193, N194, N195, N196, opas_r1, opas_r2, sign, N216,
         fasu_op_r1, N220, N221, N222, N223, N224, N225, N226, N227, N228,
         N229, N230, N231, N232, N233, N234, N254, N278, N281, N283, N285,
         N290, N291, N292, N296, \u0/N17 , \u0/N16 , \u0/expb_00 ,
         \u0/expa_00 , \u0/N11 , \u0/N10 , \u0/N7 , \u0/N6 , \u0/N5 , \u0/N4 ,
         \u0/infb_f_r , \u0/infa_f_r , \u0/expb_ff , \u0/expa_ff , \u1/N133 ,
         \u1/fracta_eq_fractb , \u1/N124 , \u1/fracta_lt_fractb , \u1/N123 ,
         \u1/N122 , \u1/add_r , \u1/signa_r , \u1/sign_d ,
         \u1/adj_op_out_sft[0] , \u1/adj_op_out_sft[1] ,
         \u1/adj_op_out_sft[2] , \u1/adj_op_out_sft[3] ,
         \u1/adj_op_out_sft[4] , \u1/adj_op_out_sft[5] ,
         \u1/adj_op_out_sft[6] , \u1/adj_op_out_sft[7] ,
         \u1/adj_op_out_sft[8] , \u1/adj_op_out_sft[9] ,
         \u1/adj_op_out_sft[10] , \u1/adj_op_out_sft[11] ,
         \u1/adj_op_out_sft[12] , \u1/adj_op_out_sft[13] ,
         \u1/exp_diff_sft[0] , \u1/adj_op[9] , \u1/N39 , \u1/N38 , \u1/N37 ,
         \u1/N36 , \u1/N35 , \u2/N73 , \u2/sign_d , \u2/N66 ,
         \u2/exp_ovf_d[0] , \u2/exp_ovf_d[1] , \u2/N44 , \u2/N43 , \u2/N42 ,
         \u2/N41 , \u2/N40 , \u2/N37 , \u2/N34 , \u2/N33 , \u2/N32 , \u2/N31 ,
         \u2/exp_tmp4[0] , \u2/exp_tmp4[1] , \u2/exp_tmp4[2] ,
         \u2/exp_tmp4[3] , \u2/exp_tmp4[4] , \u2/exp_tmp3[1] ,
         \u2/exp_tmp3[2] , \u2/exp_tmp3[3] , \u2/exp_tmp3[4] , \u2/N29 ,
         \u2/N28 , \u2/N27 , \u2/N26 , \u2/N25 , \u2/N23 , \u2/N22 , \u2/N21 ,
         \u2/N20 , \u2/N19 , \u2/N17 , \u2/N16 , \u2/N15 , \u2/N14 , \u2/N13 ,
         \u2/N12 , \u2/N11 , \u2/N10 , \u2/N9 , \u2/N8 , \u2/N7 , \u2/N6 ,
         \u3/N32 , \u3/N31 , \u3/N30 , \u3/N29 , \u3/N28 , \u3/N27 , \u3/N26 ,
         \u3/N25 , \u3/N24 , \u3/N23 , \u3/N22 , \u3/N21 , \u3/N20 , \u3/N19 ,
         \u3/N18 , \u3/N17 , \u3/N16 , \u3/N15 , \u3/N14 , \u3/N13 , \u3/N12 ,
         \u3/N11 , \u3/N10 , \u3/N9 , \u3/N8 , \u3/N7 , \u3/N6 , \u3/N5 ,
         \u3/N4 , \u3/N3 , \u5/N21 , \u5/N20 , \u5/N19 , \u5/N18 , \u5/N17 ,
         \u5/N16 , \u5/N15 , \u5/N14 , \u5/N13 , \u5/N12 , \u5/N11 , \u5/N10 ,
         \u5/N9 , \u5/N8 , \u5/N7 , \u5/N6 , \u5/N5 , \u5/N4 , \u5/N3 ,
         \u5/N2 , \u5/N1 , \u5/N0 , \u6/N23 , \u6/N22 , \u6/N21 , \u6/N20 ,
         \u6/N19 , \u6/N18 , \u6/N17 , \u6/N16 , \u6/N15 , \u6/N14 , \u6/N13 ,
         \u6/N10 , \u6/N9 , \u6/N8 , \u6/N7 , \u6/N6 , \u6/N5 , \u6/N4 ,
         \u6/N3 , \u6/N2 , \u6/N1 , \u6/N0 , \u4/N656 , \u4/N655 , \u4/N653 ,
         \u4/div_exp3[1] , \u4/fi_ldz_mi1[2] , \u4/fi_ldz_mi1[3] , \u4/N433 ,
         \u4/N432 , \u4/N431 , \u4/N430 , \u4/N429 , \u4/N428 , \u4/N427 ,
         \u4/N426 , \u4/N425 , \u4/N424 , \u4/N423 , \u4/N422 , \u4/N421 ,
         \u4/N420 , \u4/N419 , \u4/N418 , \u4/N417 , \u4/N416 , \u4/N415 ,
         \u4/N414 , \u4/N413 , \u4/N412 , \u4/N409 , \u4/N408 , \u4/N407 ,
         \u4/N406 , \u4/N405 , \u4/N404 , \u4/N403 , \u4/N402 , \u4/N401 ,
         \u4/N400 , \u4/N399 , \u4/N398 , \u4/N397 , \u4/N396 , \u4/N395 ,
         \u4/N394 , \u4/N393 , \u4/N392 , \u4/N391 , \u4/N390 , \u4/N389 ,
         \u4/N388 , \u4/N386 , \u4/exp_in_pl1[2] , \u4/exp_in_pl1[3] ,
         \u4/exp_in_pl1[4] , \u4/exp_in_pl1[5] , \u4/f2i_shft[2] ,
         \u4/f2i_shft[3] , \u4/f2i_shft[4] , \u4/div_shft2[0] ,
         \u4/fract_out_pl1[0] , \u4/fract_out_pl1[1] , \u4/fract_out_pl1[2] ,
         \u4/fract_out_pl1[3] , \u4/fract_out_pl1[4] , \u4/fract_out_pl1[5] ,
         \u4/fract_out_pl1[6] , \u4/fract_out_pl1[7] , \u4/fract_out_pl1[8] ,
         \u4/fract_out_pl1[9] , \u4/fract_out_pl1[10] , \u4/exp_next_mi[0] ,
         \u4/exp_next_mi[1] , \u4/exp_next_mi[2] , \u4/exp_next_mi[3] ,
         \u4/exp_next_mi[4] , \u4/exp_next_mi[5] , \u4/fract_out[1] ,
         \u4/fract_out[5] , \u4/exp_out[2] , n845, n851, n872, n888, n1521,
         net10316, \u2/lt_130/A[0] , \u2/lt_130/A[1] , \u2/lt_130/A[2] ,
         \u2/lt_130/A[3] , \u2/gt_140/B[5] , net11677, net11676, net11675,
         net11671, net11670, net11627, net11582, net11576, net11567, net11566,
         net11564, net11562, net11560, net11558, net11555, net11485,
         \u4/sub_409/net10540 , \u2/add_113/A[0] , \u2/add_113/A[1] ,
         \u2/add_113/A[2] , \u2/add_113/A[3] , \u2/add_113/A[4] ,
         \u2/sub_111/carry[2] , \u2/sub_111/carry[3] , \u2/sub_111/carry[4] ,
         \u2/sub_111/carry[5] , \u2/add_111/carry[2] , \u2/add_111/carry[3] ,
         \u2/add_111/carry[4] , \u2/add_111/carry[5] , net15448, net15944,
         net30297, net33278, net60630, net76048, net76254, net76619, net76645,
         net76672, net76926, net77045, net77073, net77161, net77637, net77815,
         net83296, net83361, net83364, net83368, net83402, net83403, net83407,
         net83408, net83414, net83419, net83421, net83423, net83427, net83429,
         net83432, net83438, net83439, net83736, net83747, net83754, net83765,
         net83779, net83780, net83781, net83787, net83791, net83800, net83802,
         net83806, net83807, net83811, net83812, net83820, net83821, net83827,
         net83833, net83836, net83844, net83849, net83853, net83855, net83856,
         net83860, net83861, net83862, net83863, net83864, net83868, net83869,
         net83871, net83874, net83875, net83876, net83878, net83883, net83906,
         net83913, net83925, net83927, net83933, net83934, net83936, net83940,
         net83941, net83942, net83945, net83946, net83950, net83951, net83959,
         net83963, net83967, net83968, net83969, net83971, net83972, net83973,
         net83975, net83987, net83990, net83993, net83994, net83995, net84003,
         net84010, net84012, net84015, net84021, net84024, net84044, net84047,
         net84048, net84050, net84055, net84059, net84060, net84069, net84070,
         net84072, net84073, net84076, net84079, net84080, net84081, net84083,
         net84095, net84096, net84103, net84107, net84115, net84118, net84119,
         net84128, net84133, net84134, net84135, net84136, net84138, net84146,
         net84148, net84149, net84150, net84151, net84157, net84159, net84160,
         net84165, net84166, net84167, net84168, net84169, net84191, net84199,
         net84200, net84211, net84214, net84215, net84216, net84218, net84220,
         net84236, net84249, net84253, net84254, net84263, net84265, net84266,
         net84276, net84277, net84278, net84279, net84280, net84290, net84297,
         net84298, net84299, net84305, net84310, net84312, net84314, net84315,
         net84322, net84326, net84327, net84329, net84332, net84333, net84334,
         net84341, net84343, net84344, net84347, net84352, net84366, net84368,
         net84371, net84373, net84374, net84381, net84398, net84402, net84403,
         net84421, net84445, net84448, net84449, net84450, net84453, net84458,
         net84465, net84468, net84469, net84474, net84475, net84480, net84482,
         net84487, net84488, net84490, net84498, net84500, net84501, net84502,
         net84506, net84511, net84520, net84522, net84523, net84524, net84531,
         net84532, net84548, net84549, net84550, net84551, net84552, net84555,
         net84561, net84564, net84565, net84568, net84571, net84579, net84590,
         net84591, net84595, net84598, net84599, net84600, net84601, net84602,
         net84604, net84605, net84609, net84610, net84611, net84614, net84615,
         net84617, net84619, net84624, net84625, net84626, net84629, net84632,
         net84633, net84637, net84639, net84642, net84643, net84644, net84645,
         net84647, net84648, net84649, net84652, net84655, net84656, net84659,
         net84660, net84661, net84662, net84663, net84664, net84667, net84668,
         net84669, net84672, net84675, net84684, net84702, net84722, net84749,
         net84753, net84754, net84755, net84758, net84761, net84762, net84763,
         net84764, net84765, net84766, net84767, net84768, net84774, net84775,
         net84777, net84778, net84783, net84784, net84810, net84814, net84822,
         net84823, net84839, net84840, net84842, net84847, net84848, net84853,
         net84856, net84858, net84867, net84869, net84870, net84884, net84886,
         net84887, net84890, net84900, net84901, net84906, net84907, net84911,
         net84912, net84915, net84916, net84921, net84953, net84968, net84975,
         net84982, net84983, net84990, net84992, net84995, net84996, net85004,
         net85006, net85010, net85015, net85027, net85030, net85032, net85037,
         net85038, net85039, net85040, net85041, net85043, net85045, net85046,
         net85051, net85059, net85060, net85061, net85067, net85068, net85069,
         net85071, net85076, net85080, net85091, net85093, net85095, net85096,
         net85099, net85103, net85104, net85105, net85111, net85112, net85113,
         net85114, net85115, net85116, net85123, net85124, net85126, net85127,
         net85131, net85136, net85137, net85140, net85141, net85144, net85150,
         net85164, net85168, net85169, net85170, net85171, net85176, net85178,
         net85182, net85191, net85192, net85194, net85195, net85196, net85197,
         net85200, net85203, net85204, net85205, net85206, net85207, net85210,
         net85211, net85212, net85213, net85216, net85220, net85224, net85227,
         net85232, net85234, net85247, net85257, net85263, net85280, net85281,
         net85285, net85292, net85310, net85313, net85316, net85320, net85331,
         net85336, net85351, net85361, net85365, net85369, net85373, net85374,
         net85393, net85676, net85674, net85712, net85710, net85722, net85720,
         net85718, net85716, net85738, net85736, net85732, net85730, net85728,
         net85752, net85748, net85746, net85744, net85778, net85788, net85786,
         net85794, net85790, net85828, net85832, net85842, net85847, net85854,
         net85853, net85974, net85998, net86004, net86006, net86010, net86016,
         net86038, net86037, net86061, net86090, net86096, net86106, net86113,
         net86112, net86125, net86169, net86263, net88287, net88293, net88292,
         net88319, net88421, net88427, net88440, net88500, net88503, net88510,
         net88545, net88566, net88585, net88618, net88695, net88699, net88721,
         net88877, net88896, net88950, net88972, net89029, net89078, net89121,
         net89120, net89129, net89250, net89266, net89314, net89412, net89411,
         net89485, net89537, net89543, net89546, net89624, net89677, net89681,
         net89680, net89679, net89692, net89716, net89741, net89753, net89819,
         net89817, net89863, net89862, net89919, net89924, net89926, net89933,
         net89943, net89948, net89964, net89965, net89975, net89987, net89998,
         net90007, net90026, net90031, net90037, net90047, net90064, net90074,
         net90080, net90115, net90122, net90124, net90126, net90144, net90207,
         net90211, net90210, net90217, net90252, net90268, net90287, net90290,
         net90292, net90299, net90302, net86262, net85081, net91047, net91057,
         net91056, net91059, net91070, net91069, net91075, net91095, net91112,
         net91128, net91159, net91299, net91298, net91325, net91512, net91542,
         net91548, net91555, net83406, net85166, net85160, net85157, net85155,
         net85135, net85125, net85120, net85133, net85107, net84830, net90035,
         net85337, net85335, net85162, net85147, net84910, net91467, net90997,
         net84994, net89447, net89446, net83420, net90072, net85165, net85042,
         net84909, net88895, net84452, net89856, net99868, net99874, net85272,
         net85270, net85265, net85264, net85254, net85253, net85252, net85251,
         net85250, net85189, net85163, net85684, net85261, net85187, net91177,
         net85033, net84984, net84673, net91109, net88551, net85239, net85215,
         net85214, net85177, net85098, net85087, net84503, net85260, net90215,
         net89935, net88605, net86027, net86026, net85290, net85283, net85240,
         net84969, net84960, net84957, net90019, net89300, net88636, net85360,
         net85357, net85159, net85158, net85097, net85089, net85085, net110929,
         net110951, net99862, net85079, net85190, net85188, net85184, net85083,
         net86060, net85317, net76872, net84213, net84071, net83870, net91353,
         net86171, net86015, net84677, net84394, net84393, net84387, net84386,
         net91015, net84882, \u4/fract_out[8] , \u4/fract_out[3] , net84845,
         net84844, net84456, net84110, net85199, net85193, net85185, net85143,
         net85142, net84043, net84033, net84029, net84028, net84026, net85342,
         net86174, net84414, net84075, net85020, net85018, net84974, net85021,
         net84913, net84895, net89073, net84484, net84409, net84401, net84390,
         \u4/fract_out[6] , net84113, net89595, net84553, net84473, net84770,
         net84678, net84573, net84519, net84518, net90110, net88332, net85297,
         net85296, net85186, net85161, net85048, net84030, net84027, net89917,
         net89077, net89076, net86160, net84408, net84385, net84372, net89372,
         net85017, net84967, net84956, net85384, net85248, net85180, net85179,
         net85084, net85082, net85077, net84757, net76352, net84584, net85975,
         net85678, net85387, net85349, net85181, net85174, net85128, net85108,
         net84301, net91511, net91404, net84576, net84575, net84574, net88374,
         net84206, net84204, net84202, net84201, net84085, net84074, net91375,
         net89842, net89224, net89055, net89054, net85831, net84963, net84950,
         net84948, net99831, net84651, net84554, net84483, net89615, net86165,
         net85827, net83974, net83813, net84854, net84846, net84566, net84064,
         net84052, net84051, net84025, net83819, \u4/fract_out[7] ,
         \u4/fract_out[4] , net91150, net84908, net84836, net84829, net84811,
         net84808, net84769, net84586, net84572, net84570, net84569, net89664,
         net89663, net84683, net84679, net84676, net84674, net84472, net84471,
         net84451, net86067, net83394, net83393, net84606, net83395, net89736,
         net89658, net89657, net88646, net83398, \u4/exp_out[4] , net85742,
         net85740, net85726, net85724, net85323, net85028, net84588, net91144,
         net90079, net85846, net85756, net85754, net84658, net84657, net84654,
         net84014, \u4/f2i_shft[1] , net83417, net83416, net83392, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1539, n1541, n1543, n1546, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1718,
         n1719, n1720, n1721, n1722, n1723, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1736, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1969, n1970, n1971, n1972, n1973, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323;
  wire   [15:10] opa_r;
  wire   [15:10] opb_r;
  wire   [1:0] rmode_r1;
  wire   [1:0] rmode_r2;
  wire   [1:0] rmode_r3;
  wire   [2:0] fpu_op_r1;
  wire   [2:0] fpu_op_r2;
  wire   [13:0] fracta;
  wire   [13:0] fractb;
  wire   [9:0] fracta_mul;
  wire   [1:0] exp_ovf;
  wire   [2:0] underflow_fmul_d;
  wire   [14:1] fract_out_q;
  wire   [21:0] prod;
  wire   [22:0] quo;
  wire   [3:0] div_opa_ldz_r1;
  wire   [3:0] div_opa_ldz_r2;
  wire   [4:1] exp_r;
  wire   [11:4] opa_r1;
  wire   [10:9] fract_denorm;
  wire   [2:1] underflow_fmul_r;
  wire   [13:0] \u1/fractb_s ;
  wire   [13:0] \u1/fracta_s ;
  wire   [2:1] \u2/underflow_d ;
  wire   [21:0] \u5/prod1 ;
  wire   [23:0] \u6/remainder ;
  wire   [23:0] \u6/quo1 ;
  wire   [27:23] \u4/exp_f2i_1 ;
  wire   [2:0] \u4/shift_left ;
  wire   [4:0] \u4/shift_right ;
  wire   [4:3] \u4/add_407/carry ;
  wire   [4:2] \u2/add_115/carry ;
  wire   [4:2] \u2/add_113/carry ;
  wire   [4:1] \u2/add_110/carry ;
  wire   [5:1] \u2/sub_110/carry ;
  wire   [20:8] \sub_435_3/carry ;
  wire   [10:2] \sub_435_b0/carry ;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45;

  OR2_X2 \u4/C1739  ( .A1(\u4/N655 ), .A2(net30297), .ZN(\u4/N656 ) );
  OR2_X2 \u4/C1742  ( .A1(net85842), .A2(n2997), .ZN(\u4/N653 ) );
  OR2_X2 \u4/C1935  ( .A1(\u4/shift_right [4]), .A2(\u4/shift_right [3]), .ZN(
        \u4/N386 ) );
  AOI22_X2 U16 ( .A1(\u4/div_exp3[1] ), .A2(net15944), .B1(n3009), .B2(
        net77815), .ZN(n845) );
  OAI211_X2 U18 ( .C1(net89919), .C2(n3010), .A(n851), .B(n1669), .ZN(
        \u4/exp_out[2] ) );
  OAI221_X2 U100 ( .B1(net83296), .B2(n872), .C1(n888), .C2(net85794), .A(
        n1664), .ZN(\u4/shift_right [0]) );
  DFF_X2 \opa_r_reg[15]  ( .D(opa[15]), .CK(clk), .Q(opa_r[15]), .QN(n1569) );
  DFF_X2 \opa_r_reg[14]  ( .D(opa[14]), .CK(clk), .Q(opa_r[14]), .QN(n1594) );
  DFF_X2 \opa_r_reg[13]  ( .D(opa[13]), .CK(clk), .Q(opa_r[13]), .QN(n1560) );
  DFF_X2 \opa_r_reg[12]  ( .D(opa[12]), .CK(clk), .Q(opa_r[12]), .QN(n1573) );
  DFF_X2 \opa_r_reg[11]  ( .D(opa[11]), .CK(clk), .Q(opa_r[11]), .QN(n1725) );
  DFF_X2 \opa_r_reg[10]  ( .D(opa[10]), .CK(clk), .Q(opa_r[10]), .QN(n1723) );
  DFF_X2 \opa_r_reg[9]  ( .D(opa[9]), .CK(clk), .Q(fracta_mul[9]), .QN(n3120)
         );
  DFF_X2 \opa_r_reg[8]  ( .D(opa[8]), .CK(clk), .Q(fracta_mul[8]), .QN(n3119)
         );
  DFF_X2 \opa_r_reg[7]  ( .D(opa[7]), .CK(clk), .Q(fracta_mul[7]), .QN(n3118)
         );
  DFF_X2 \opa_r_reg[6]  ( .D(opa[6]), .CK(clk), .Q(fracta_mul[6]), .QN(n3117)
         );
  DFF_X2 \opa_r_reg[5]  ( .D(opa[5]), .CK(clk), .Q(fracta_mul[5]), .QN(n3116)
         );
  DFF_X2 \opa_r_reg[4]  ( .D(opa[4]), .CK(clk), .Q(fracta_mul[4]), .QN(n3115)
         );
  DFF_X2 \opa_r_reg[3]  ( .D(opa[3]), .CK(clk), .Q(fracta_mul[3]), .QN(n3114)
         );
  DFF_X2 \opa_r_reg[2]  ( .D(opa[2]), .CK(clk), .Q(fracta_mul[2]), .QN(n3113)
         );
  DFF_X2 \opa_r_reg[1]  ( .D(opa[1]), .CK(clk), .Q(fracta_mul[1]), .QN(n3112)
         );
  DFF_X2 \opa_r_reg[0]  ( .D(opa[0]), .CK(clk), .Q(fracta_mul[0]), .QN(n3111)
         );
  DFF_X2 \opb_r_reg[15]  ( .D(opb[15]), .CK(clk), .Q(opb_r[15]), .QN(n1686) );
  DFF_X2 \opb_r_reg[14]  ( .D(opb[14]), .CK(clk), .Q(opb_r[14]), .QN(n1734) );
  DFF_X2 \opb_r_reg[13]  ( .D(opb[13]), .CK(clk), .Q(opb_r[13]), .QN(n1728) );
  DFF_X2 \opb_r_reg[12]  ( .D(opb[12]), .CK(clk), .Q(opb_r[12]), .QN(n1727) );
  DFF_X2 \opb_r_reg[11]  ( .D(opb[11]), .CK(clk), .Q(opb_r[11]), .QN(n1730) );
  DFF_X2 \opb_r_reg[10]  ( .D(opb[10]), .CK(clk), .Q(opb_r[10]), .QN(n1726) );
  DFF_X2 \opb_r_reg[9]  ( .D(opb[9]), .CK(clk), .Q(\u6/N9 ), .QN(n3110) );
  DFF_X2 \opb_r_reg[8]  ( .D(opb[8]), .CK(clk), .Q(\u6/N8 ), .QN(n3109) );
  DFF_X2 \opb_r_reg[7]  ( .D(opb[7]), .CK(clk), .Q(\u6/N7 ), .QN(n3108) );
  DFF_X2 \opb_r_reg[6]  ( .D(opb[6]), .CK(clk), .Q(\u6/N6 ), .QN(n3107) );
  DFF_X2 \opb_r_reg[5]  ( .D(opb[5]), .CK(clk), .Q(\u6/N5 ), .QN(n3106) );
  DFF_X2 \opb_r_reg[4]  ( .D(opb[4]), .CK(clk), .Q(\u6/N4 ), .QN(n3105) );
  DFF_X2 \opb_r_reg[3]  ( .D(opb[3]), .CK(clk), .Q(\u6/N3 ), .QN(n3104) );
  DFF_X2 \opb_r_reg[2]  ( .D(opb[2]), .CK(clk), .Q(\u6/N2 ), .QN(n3103) );
  DFF_X2 \opb_r_reg[1]  ( .D(opb[1]), .CK(clk), .Q(\u6/N1 ), .QN(n3102) );
  DFF_X2 \opb_r_reg[0]  ( .D(opb[0]), .CK(clk), .Q(\u6/N0 ), .QN(n3101) );
  DFF_X2 \rmode_r1_reg[1]  ( .D(rmode[1]), .CK(clk), .Q(rmode_r1[1]) );
  DFF_X2 \rmode_r1_reg[0]  ( .D(rmode[0]), .CK(clk), .Q(rmode_r1[0]) );
  DFF_X2 \rmode_r2_reg[1]  ( .D(rmode_r1[1]), .CK(clk), .Q(rmode_r2[1]) );
  DFF_X2 \rmode_r2_reg[0]  ( .D(rmode_r1[0]), .CK(clk), .Q(rmode_r2[0]) );
  DFF_X2 \rmode_r3_reg[1]  ( .D(rmode_r2[1]), .CK(clk), .Q(rmode_r3[1]), .QN(
        n1768) );
  DFF_X2 \rmode_r3_reg[0]  ( .D(rmode_r2[0]), .CK(clk), .Q(rmode_r3[0]), .QN(
        n1614) );
  DFF_X2 \fpu_op_r1_reg[2]  ( .D(fpu_op[2]), .CK(clk), .Q(fpu_op_r1[2]), .QN(
        n3100) );
  DFF_X2 \fpu_op_r1_reg[1]  ( .D(fpu_op[1]), .CK(clk), .Q(fpu_op_r1[1]) );
  DFF_X2 \fpu_op_r1_reg[0]  ( .D(fpu_op[0]), .CK(clk), .Q(fpu_op_r1[0]), .QN(
        n3317) );
  DFF_X2 \fpu_op_r2_reg[2]  ( .D(fpu_op_r1[2]), .CK(clk), .Q(fpu_op_r2[2]), 
        .QN(n3099) );
  DFF_X2 \fpu_op_r2_reg[1]  ( .D(fpu_op_r1[1]), .CK(clk), .Q(fpu_op_r2[1]), 
        .QN(n3098) );
  DFF_X2 \fpu_op_r2_reg[0]  ( .D(fpu_op_r1[0]), .CK(clk), .Q(fpu_op_r2[0]), 
        .QN(n3097) );
  DFF_X2 \fpu_op_r3_reg[2]  ( .D(fpu_op_r2[2]), .CK(clk), .Q(net86090), .QN(
        net11677) );
  DFF_X2 \fpu_op_r3_reg[1]  ( .D(fpu_op_r2[1]), .CK(clk), .Q(net86006), .QN(
        net11676) );
  DFF_X2 \fpu_op_r3_reg[0]  ( .D(fpu_op_r2[0]), .CK(clk), .Q(net88695), .QN(
        net11675) );
  DFF_X2 \div_opa_ldz_r1_reg[3]  ( .D(N34), .CK(clk), .Q(div_opa_ldz_r1[3]) );
  DFF_X2 \div_opa_ldz_r1_reg[2]  ( .D(N44), .CK(clk), .Q(div_opa_ldz_r1[2]) );
  DFF_X2 \div_opa_ldz_r1_reg[1]  ( .D(N56), .CK(clk), .Q(div_opa_ldz_r1[1]) );
  DFF_X2 \div_opa_ldz_r1_reg[0]  ( .D(N65), .CK(clk), .Q(div_opa_ldz_r1[0]) );
  DFF_X2 \div_opa_ldz_r2_reg[3]  ( .D(div_opa_ldz_r1[3]), .CK(clk), .Q(
        div_opa_ldz_r2[3]), .QN(n1663) );
  DFF_X2 \div_opa_ldz_r2_reg[2]  ( .D(div_opa_ldz_r1[2]), .CK(clk), .Q(
        div_opa_ldz_r2[2]), .QN(n3096) );
  DFF_X2 \div_opa_ldz_r2_reg[1]  ( .D(div_opa_ldz_r1[1]), .CK(clk), .Q(
        div_opa_ldz_r2[1]), .QN(net11671) );
  DFF_X2 \div_opa_ldz_r2_reg[0]  ( .D(div_opa_ldz_r1[0]), .CK(clk), .Q(
        div_opa_ldz_r2[0]), .QN(net11670) );
  DFF_X2 \opa_r1_reg[14]  ( .D(opa_r[14]), .CK(clk), .QN(n1635) );
  DFF_X2 \opa_r1_reg[13]  ( .D(opa_r[13]), .CK(clk), .QN(n1636) );
  DFF_X2 \opa_r1_reg[12]  ( .D(opa_r[12]), .CK(clk), .QN(n1637) );
  DFF_X2 \opa_r1_reg[11]  ( .D(opa_r[11]), .CK(clk), .Q(opa_r1[11]), .QN(n1672) );
  DFF_X2 \opa_r1_reg[10]  ( .D(opa_r[10]), .CK(clk), .Q(opa_r1[10]), .QN(n1673) );
  DFF_X2 \opa_r1_reg[9]  ( .D(fracta_mul[9]), .CK(clk), .QN(n1624) );
  DFF_X2 \opa_r1_reg[8]  ( .D(fracta_mul[8]), .CK(clk), .QN(n1625) );
  DFF_X2 \opa_r1_reg[7]  ( .D(fracta_mul[7]), .CK(clk), .QN(n1626) );
  DFF_X2 \opa_r1_reg[6]  ( .D(fracta_mul[6]), .CK(clk), .QN(n1627) );
  DFF_X2 \opa_r1_reg[5]  ( .D(fracta_mul[5]), .CK(clk), .Q(opa_r1[5]), .QN(
        n1678) );
  DFF_X2 \opa_r1_reg[4]  ( .D(fracta_mul[4]), .CK(clk), .Q(opa_r1[4]), .QN(
        n1679) );
  DFF_X2 \opa_r1_reg[3]  ( .D(fracta_mul[3]), .CK(clk), .QN(n1674) );
  DFF_X2 \opa_r1_reg[2]  ( .D(fracta_mul[2]), .CK(clk), .QN(n1675) );
  DFF_X2 \opa_r1_reg[1]  ( .D(fracta_mul[1]), .CK(clk), .QN(n1676) );
  DFF_X2 \opa_r1_reg[0]  ( .D(fracta_mul[0]), .CK(clk), .Q(N106), .QN(n1680)
         );
  DFF_X2 opas_r1_reg ( .D(opa_r[15]), .CK(clk), .Q(opas_r1) );
  DFF_X2 opas_r2_reg ( .D(opas_r1), .CK(clk), .Q(opas_r2), .QN(n1608) );
  DFF_X2 \u0/fractb_00_reg  ( .D(n3316), .CK(clk), .QN(n3095) );
  DFF_X2 \u0/fracta_00_reg  ( .D(n3314), .CK(clk), .QN(n3094) );
  DFF_X2 \u0/expb_00_reg  ( .D(n3013), .CK(clk), .Q(\u0/expb_00 ), .QN(n3093)
         );
  DFF_X2 \u0/opb_dn_reg  ( .D(\u0/expb_00 ), .CK(clk), .Q(opb_dn), .QN(
        net85974) );
  DFF_X2 \u0/opb_00_reg  ( .D(\u0/N17 ), .CK(clk), .Q(opb_00), .QN(n1570) );
  DFF_X2 \u0/expa_00_reg  ( .D(n3012), .CK(clk), .Q(\u0/expa_00 ), .QN(n3092)
         );
  DFF_X2 \u0/opa_dn_reg  ( .D(\u0/expa_00 ), .CK(clk), .Q(opa_dn), .QN(n1641)
         );
  DFF_X2 \u0/opa_00_reg  ( .D(\u0/N16 ), .CK(clk), .Q(opa_00), .QN(n1615) );
  DFF_X2 \u0/opb_nan_reg  ( .D(\u0/N11 ), .CK(clk), .Q(opb_nan), .QN(n1684) );
  DFF_X2 \u0/opa_nan_reg  ( .D(\u0/N10 ), .CK(clk), .Q(opa_nan), .QN(n1681) );
  DFF_X2 opa_nan_r_reg ( .D(N291), .CK(clk), .QN(n3091) );
  DFF_X2 \u0/snan_r_b_reg  ( .D(\u0/N5 ), .CK(clk), .QN(n3090) );
  DFF_X2 \u0/qnan_r_b_reg  ( .D(\u6/N9 ), .CK(clk), .QN(n3089) );
  DFF_X2 \u0/snan_r_a_reg  ( .D(\u0/N4 ), .CK(clk), .QN(n3088) );
  DFF_X2 \u0/qnan_r_a_reg  ( .D(fracta_mul[9]), .CK(clk), .QN(n3087) );
  DFF_X2 \u0/infb_f_r_reg  ( .D(n3316), .CK(clk), .Q(\u0/infb_f_r ) );
  DFF_X2 \u0/infa_f_r_reg  ( .D(n3314), .CK(clk), .Q(\u0/infa_f_r ) );
  DFF_X2 \u0/expb_ff_reg  ( .D(n3315), .CK(clk), .Q(\u0/expb_ff ), .QN(n1677)
         );
  DFF_X2 \u0/opb_inf_reg  ( .D(n3322), .CK(clk), .Q(opb_inf), .QN(n1595) );
  DFF_X2 \u0/expa_ff_reg  ( .D(n3312), .CK(clk), .Q(\u0/expa_ff ), .QN(n1591)
         );
  DFF_X2 \u0/snan_reg  ( .D(n3320), .CK(clk), .Q(snan_d), .QN(n3086) );
  DFF_X2 snan_reg ( .D(snan_d), .CK(clk), .Q(snan) );
  DFF_X2 \u0/qnan_reg  ( .D(n3321), .CK(clk), .QN(n3085) );
  DFF_X2 \u0/opa_inf_reg  ( .D(n3323), .CK(clk), .Q(opa_inf), .QN(n1572) );
  DFF_X2 div_by_zero_reg ( .D(N292), .CK(clk), .Q(div_by_zero) );
  DFF_X2 \u0/inf_reg  ( .D(\u0/N7 ), .CK(clk), .Q(n1576) );
  DFF_X2 \u0/ind_reg  ( .D(\u0/N6 ), .CK(clk), .Q(n1611) );
  DFF_X2 \u1/fasu_op_reg  ( .D(n3299), .CK(clk), .Q(fasu_op), .QN(n3084) );
  DFF_X2 fasu_op_r1_reg ( .D(fasu_op), .CK(clk), .Q(fasu_op_r1) );
  DFF_X2 fasu_op_r2_reg ( .D(fasu_op_r1), .CK(clk), .QN(net11627) );
  DFF_X2 qnan_reg ( .D(N283), .CK(clk), .Q(qnan) );
  DFF_X2 \u1/fracta_eq_fractb_reg  ( .D(\u1/N124 ), .CK(clk), .Q(
        \u1/fracta_eq_fractb ) );
  DFF_X2 \u1/fracta_lt_fractb_reg  ( .D(\u1/N123 ), .CK(clk), .Q(
        \u1/fracta_lt_fractb ), .QN(n1683) );
  DFF_X2 \u1/add_r_reg  ( .D(n3317), .CK(clk), .Q(\u1/add_r ) );
  DFF_X2 \u1/signb_r_reg  ( .D(opb_r[15]), .CK(clk), .QN(n1671) );
  DFF_X2 \u1/signa_r_reg  ( .D(opa_r[15]), .CK(clk), .Q(\u1/signa_r ), .QN(
        n1682) );
  DFF_X2 \u1/result_zero_sign_reg  ( .D(\u1/N122 ), .CK(clk), .Q(
        result_zero_sign_d) );
  DFF_X2 \u1/nan_sign_reg  ( .D(\u1/N133 ), .CK(clk), .Q(nan_sign_d) );
  DFF_X2 sign_fasu_r_reg ( .D(sign_fasu), .CK(clk), .Q(sign_fasu_r), .QN(n1685) );
  DFF_X2 \u1/fractb_out_reg[4]  ( .D(\u1/fractb_s [4]), .CK(clk), .Q(fractb[4]) );
  DFF_X2 \u1/fracta_out_reg[0]  ( .D(\u1/fracta_s [0]), .CK(clk), .Q(fracta[0]) );
  DFF_X2 \u1/fracta_out_reg[2]  ( .D(\u1/fracta_s [2]), .CK(clk), .Q(fracta[2]) );
  DFF_X2 \u1/fracta_out_reg[3]  ( .D(\u1/fracta_s [3]), .CK(clk), .Q(fracta[3]) );
  DFF_X2 \u1/fracta_out_reg[4]  ( .D(\u1/fracta_s [4]), .CK(clk), .Q(fracta[4]) );
  DFF_X2 \u1/fracta_out_reg[13]  ( .D(\u1/fracta_s [13]), .CK(clk), .Q(
        fracta[13]) );
  DFF_X2 \fract_out_q_reg[1]  ( .D(n3297), .CK(clk), .Q(fract_out_q[1]) );
  DFF_X2 \fract_out_q_reg[2]  ( .D(n3296), .CK(clk), .Q(fract_out_q[2]) );
  DFF_X2 \fract_out_q_reg[3]  ( .D(n3295), .CK(clk), .Q(fract_out_q[3]) );
  DFF_X2 \fract_out_q_reg[4]  ( .D(n3294), .CK(clk), .Q(fract_out_q[4]) );
  DFF_X2 \fract_out_q_reg[5]  ( .D(n3293), .CK(clk), .Q(fract_out_q[5]) );
  DFF_X2 \fract_out_q_reg[6]  ( .D(n3292), .CK(clk), .Q(fract_out_q[6]) );
  DFF_X2 \fract_out_q_reg[7]  ( .D(n3291), .CK(clk), .Q(fract_out_q[7]) );
  DFF_X2 \fract_out_q_reg[8]  ( .D(n3290), .CK(clk), .Q(fract_out_q[8]) );
  DFF_X2 \fract_out_q_reg[9]  ( .D(n3289), .CK(clk), .Q(fract_out_q[9]) );
  DFF_X2 \fract_out_q_reg[13]  ( .D(n3285), .CK(clk), .Q(fract_out_q[13]) );
  DFF_X2 \u1/exp_dn_out_reg[0]  ( .D(\u1/N35 ), .CK(clk), .QN(n3083) );
  DFF_X2 \u1/exp_dn_out_reg[1]  ( .D(\u1/N36 ), .CK(clk), .QN(n3082) );
  DFF_X2 \u1/exp_dn_out_reg[2]  ( .D(\u1/N37 ), .CK(clk), .QN(n3081) );
  DFF_X2 \u1/exp_dn_out_reg[3]  ( .D(\u1/N38 ), .CK(clk), .QN(n3080) );
  DFF_X2 \u1/exp_dn_out_reg[4]  ( .D(\u1/N39 ), .CK(clk), .QN(n3079) );
  DFF_X2 \u2/sign_exe_reg  ( .D(\u2/N73 ), .CK(clk), .Q(sign_exe) );
  DFF_X2 sign_exe_r_reg ( .D(sign_exe), .CK(clk), .Q(sign_exe_r), .QN(n1617)
         );
  DFF_X2 \u2/sign_reg  ( .D(\u2/sign_d ), .CK(clk), .Q(sign_mul) );
  DFF_X2 sign_mul_r_reg ( .D(sign_mul), .CK(clk), .Q(sign_mul_r), .QN(n1644)
         );
  DFF_X2 sign_reg ( .D(N216), .CK(clk), .Q(sign), .QN(net86016) );
  DFF_X2 \fract_i2f_reg[20]  ( .D(N195), .CK(clk), .Q(n1609) );
  DFF_X2 \fract_i2f_reg[18]  ( .D(N193), .CK(clk), .QN(n3078) );
  DFF_X2 \fract_i2f_reg[16]  ( .D(N191), .CK(clk), .QN(n3077) );
  DFF_X2 \fract_i2f_reg[14]  ( .D(N189), .CK(clk), .QN(n3076) );
  DFF_X2 \fract_i2f_reg[13]  ( .D(N188), .CK(clk), .QN(n3075) );
  DFF_X2 \fract_i2f_reg[10]  ( .D(N185), .CK(clk), .QN(net11582) );
  DFF_X2 \fract_i2f_reg[8]  ( .D(N183), .CK(clk), .QN(n3074) );
  DFF_X2 \fract_i2f_reg[7]  ( .D(N182), .CK(clk), .Q(\fract_i2f[7] ) );
  DFF_X2 \fract_i2f_reg[4]  ( .D(N179), .CK(clk), .QN(net11576) );
  DFF_X2 \fract_i2f_reg[3]  ( .D(n3281), .CK(clk), .QN(n3073) );
  DFF_X2 \fract_i2f_reg[1]  ( .D(n3283), .CK(clk), .QN(n3072) );
  DFF_X2 \u2/inf_reg  ( .D(\u2/N66 ), .CK(clk), .Q(inf_mul) );
  DFF_X2 inf_mul_r_reg ( .D(inf_mul), .CK(clk), .Q(n1631), .QN(n3071) );
  DFF_X2 \u2/underflow_reg[0]  ( .D(n1655), .CK(clk), .Q(underflow_fmul_d[0])
         );
  DFF_X2 \underflow_fmul_r_reg[0]  ( .D(underflow_fmul_d[0]), .CK(clk), .Q(
        n1612) );
  DFF_X2 \u2/underflow_reg[1]  ( .D(\u2/underflow_d [1]), .CK(clk), .Q(
        underflow_fmul_d[1]) );
  DFF_X2 \underflow_fmul_r_reg[1]  ( .D(underflow_fmul_d[1]), .CK(clk), .Q(
        underflow_fmul_r[1]) );
  DFF_X2 \u2/underflow_reg[2]  ( .D(\u2/underflow_d [2]), .CK(clk), .Q(
        underflow_fmul_d[2]) );
  DFF_X2 \underflow_fmul_r_reg[2]  ( .D(underflow_fmul_d[2]), .CK(clk), .Q(
        underflow_fmul_r[2]) );
  DFF_X2 \u2/exp_ovf_reg[0]  ( .D(\u2/exp_ovf_d[0] ), .CK(clk), .Q(exp_ovf[0])
         );
  DFF_X2 \exp_ovf_r_reg[0]  ( .D(exp_ovf[0]), .CK(clk), .Q(n1596), .QN(
        net11567) );
  DFF_X2 \u2/exp_ovf_reg[1]  ( .D(\u2/exp_ovf_d[1] ), .CK(clk), .Q(exp_ovf[1])
         );
  DFF_X2 \exp_ovf_r_reg[1]  ( .D(exp_ovf[1]), .CK(clk), .Q(n1571), .QN(
        net11566) );
  DFF_X2 \u2/exp_out_reg[0]  ( .D(\u2/N40 ), .CK(clk), .QN(n3070) );
  DFF_X2 \exp_r_reg[0]  ( .D(N96), .CK(clk), .Q(\u4/div_shft2[0] ), .QN(
        net11564) );
  DFF_X2 \u2/exp_out_reg[1]  ( .D(\u2/N41 ), .CK(clk), .QN(n3069) );
  DFF_X2 \exp_r_reg[1]  ( .D(N97), .CK(clk), .Q(exp_r[1]), .QN(net11562) );
  DFF_X2 \u2/exp_out_reg[2]  ( .D(\u2/N42 ), .CK(clk), .QN(n3068) );
  DFF_X2 \exp_r_reg[2]  ( .D(N98), .CK(clk), .Q(exp_r[2]), .QN(net11560) );
  DFF_X2 \u2/exp_out_reg[3]  ( .D(\u2/N43 ), .CK(clk), .QN(n3067) );
  DFF_X2 \exp_r_reg[3]  ( .D(N99), .CK(clk), .Q(exp_r[3]), .QN(net11558) );
  DFF_X2 \u2/exp_out_reg[4]  ( .D(\u2/N44 ), .CK(clk), .QN(n3066) );
  DFF_X2 inf_mul2_reg ( .D(N296), .CK(clk), .QN(n3065) );
  DFF_X2 \exp_r_reg[4]  ( .D(N100), .CK(clk), .Q(exp_r[4]), .QN(net11555) );
  DFF_X2 \u5/prod1_reg[0]  ( .D(\u5/N0 ), .CK(clk), .Q(\u5/prod1 [0]) );
  DFF_X2 \u5/prod_reg[0]  ( .D(\u5/prod1 [0]), .CK(clk), .Q(prod[0]) );
  DFF_X2 \u5/prod1_reg[1]  ( .D(\u5/N1 ), .CK(clk), .Q(\u5/prod1 [1]) );
  DFF_X2 \u5/prod_reg[1]  ( .D(\u5/prod1 [1]), .CK(clk), .Q(prod[1]) );
  DFF_X2 \u5/prod1_reg[2]  ( .D(\u5/N2 ), .CK(clk), .Q(\u5/prod1 [2]) );
  DFF_X2 \u5/prod_reg[2]  ( .D(\u5/prod1 [2]), .CK(clk), .Q(prod[2]) );
  DFF_X2 \u5/prod1_reg[3]  ( .D(\u5/N3 ), .CK(clk), .Q(\u5/prod1 [3]) );
  DFF_X2 \u5/prod_reg[3]  ( .D(\u5/prod1 [3]), .CK(clk), .Q(prod[3]), .QN(
        net89543) );
  DFF_X2 \u5/prod1_reg[4]  ( .D(\u5/N4 ), .CK(clk), .Q(\u5/prod1 [4]) );
  DFF_X2 \u5/prod_reg[4]  ( .D(\u5/prod1 [4]), .CK(clk), .Q(prod[4]), .QN(
        net88972) );
  DFF_X2 \u5/prod1_reg[5]  ( .D(\u5/N5 ), .CK(clk), .Q(\u5/prod1 [5]) );
  DFF_X2 \u5/prod_reg[5]  ( .D(\u5/prod1 [5]), .CK(clk), .Q(prod[5]) );
  DFF_X2 \u5/prod1_reg[6]  ( .D(\u5/N6 ), .CK(clk), .Q(\u5/prod1 [6]) );
  DFF_X2 \u5/prod_reg[6]  ( .D(\u5/prod1 [6]), .CK(clk), .Q(prod[6]) );
  DFF_X2 \u5/prod1_reg[7]  ( .D(\u5/N7 ), .CK(clk), .Q(\u5/prod1 [7]) );
  DFF_X2 \u5/prod_reg[7]  ( .D(\u5/prod1 [7]), .CK(clk), .Q(prod[7]), .QN(
        n1604) );
  DFF_X2 \u5/prod_reg[8]  ( .D(\u5/prod1 [8]), .CK(clk), .Q(prod[8]) );
  DFF_X2 \u5/prod1_reg[9]  ( .D(\u5/N9 ), .CK(clk), .Q(\u5/prod1 [9]) );
  DFF_X2 \u5/prod_reg[9]  ( .D(\u5/prod1 [9]), .CK(clk), .Q(prod[9]) );
  DFF_X2 \u5/prod_reg[10]  ( .D(\u5/prod1 [10]), .CK(clk), .Q(prod[10]) );
  DFF_X2 \u5/prod_reg[11]  ( .D(\u5/prod1 [11]), .CK(clk), .Q(prod[11]) );
  DFF_X2 \u5/prod1_reg[12]  ( .D(\u5/N12 ), .CK(clk), .Q(\u5/prod1 [12]) );
  DFF_X2 \u5/prod_reg[12]  ( .D(\u5/prod1 [12]), .CK(clk), .Q(prod[12]) );
  DFF_X2 \u5/prod_reg[13]  ( .D(\u5/prod1 [13]), .CK(clk), .Q(prod[13]) );
  DFF_X2 \u5/prod1_reg[14]  ( .D(\u5/N14 ), .CK(clk), .Q(\u5/prod1 [14]) );
  DFF_X2 \u5/prod_reg[14]  ( .D(\u5/prod1 [14]), .CK(clk), .Q(prod[14]) );
  DFF_X2 \u5/prod1_reg[15]  ( .D(\u5/N15 ), .CK(clk), .Q(\u5/prod1 [15]) );
  DFF_X2 \u5/prod_reg[15]  ( .D(\u5/prod1 [15]), .CK(clk), .Q(prod[15]) );
  DFF_X2 \u5/prod1_reg[16]  ( .D(\u5/N16 ), .CK(clk), .Q(\u5/prod1 [16]) );
  DFF_X2 \u5/prod_reg[16]  ( .D(\u5/prod1 [16]), .CK(clk), .Q(prod[16]) );
  DFF_X2 \u5/prod_reg[17]  ( .D(\u5/prod1 [17]), .CK(clk), .Q(prod[17]) );
  DFF_X2 \u5/prod1_reg[18]  ( .D(\u5/N18 ), .CK(clk), .Q(\u5/prod1 [18]) );
  DFF_X2 \u5/prod_reg[18]  ( .D(\u5/prod1 [18]), .CK(clk), .Q(prod[18]) );
  DFF_X2 \u5/prod1_reg[19]  ( .D(\u5/N19 ), .CK(clk), .Q(\u5/prod1 [19]) );
  DFF_X2 \u5/prod_reg[19]  ( .D(\u5/prod1 [19]), .CK(clk), .Q(prod[19]) );
  DFF_X2 \u5/prod1_reg[20]  ( .D(\u5/N20 ), .CK(clk), .Q(\u5/prod1 [20]) );
  DFF_X2 \u5/prod_reg[20]  ( .D(\u5/prod1 [20]), .CK(clk), .Q(prod[20]) );
  DFF_X2 \u5/prod1_reg[21]  ( .D(\u5/N21 ), .CK(clk), .Q(\u5/prod1 [21]) );
  DFF_X2 \u5/prod_reg[21]  ( .D(\u5/prod1 [21]), .CK(clk), .Q(prod[21]) );
  DFF_X2 \u6/remainder_reg[0]  ( .D(\u6/N0 ), .CK(clk), .Q(\u6/remainder [0])
         );
  DFF_X2 \u6/rem_reg[0]  ( .D(\u6/remainder [0]), .CK(clk), .QN(n1568) );
  DFF_X2 \u6/remainder_reg[1]  ( .D(\u6/N1 ), .CK(clk), .Q(\u6/remainder [1])
         );
  DFF_X2 \u6/rem_reg[1]  ( .D(\u6/remainder [1]), .CK(clk), .QN(n3064) );
  DFF_X2 \u6/remainder_reg[2]  ( .D(\u6/N2 ), .CK(clk), .Q(\u6/remainder [2])
         );
  DFF_X2 \u6/rem_reg[2]  ( .D(\u6/remainder [2]), .CK(clk), .QN(n3063) );
  DFF_X2 \u6/remainder_reg[3]  ( .D(\u6/N3 ), .CK(clk), .Q(\u6/remainder [3])
         );
  DFF_X2 \u6/rem_reg[3]  ( .D(\u6/remainder [3]), .CK(clk), .QN(n3062) );
  DFF_X2 \u6/remainder_reg[4]  ( .D(\u6/N4 ), .CK(clk), .Q(\u6/remainder [4])
         );
  DFF_X2 \u6/rem_reg[4]  ( .D(\u6/remainder [4]), .CK(clk), .QN(n1587) );
  DFF_X2 \u6/remainder_reg[5]  ( .D(\u6/N5 ), .CK(clk), .Q(\u6/remainder [5])
         );
  DFF_X2 \u6/rem_reg[5]  ( .D(\u6/remainder [5]), .CK(clk), .QN(n1620) );
  DFF_X2 \u6/remainder_reg[6]  ( .D(\u6/N6 ), .CK(clk), .Q(\u6/remainder [6])
         );
  DFF_X2 \u6/rem_reg[6]  ( .D(\u6/remainder [6]), .CK(clk), .QN(n1584) );
  DFF_X2 \u6/remainder_reg[7]  ( .D(\u6/N7 ), .CK(clk), .Q(\u6/remainder [7])
         );
  DFF_X2 \u6/rem_reg[7]  ( .D(\u6/remainder [7]), .CK(clk), .QN(n3061) );
  DFF_X2 \u6/remainder_reg[8]  ( .D(\u6/N8 ), .CK(clk), .Q(\u6/remainder [8])
         );
  DFF_X2 \u6/rem_reg[8]  ( .D(\u6/remainder [8]), .CK(clk), .QN(n3060) );
  DFF_X2 \u6/remainder_reg[9]  ( .D(\u6/N9 ), .CK(clk), .Q(\u6/remainder [9])
         );
  DFF_X2 \u6/rem_reg[9]  ( .D(\u6/remainder [9]), .CK(clk), .QN(n3059) );
  DFF_X2 \u6/remainder_reg[10]  ( .D(n1731), .CK(clk), .Q(\u6/remainder [10])
         );
  DFF_X2 \u6/rem_reg[10]  ( .D(\u6/remainder [10]), .CK(clk), .QN(n1616) );
  DFF_X2 \u6/remainder_reg[13]  ( .D(\u6/N13 ), .CK(clk), .Q(
        \u6/remainder [13]) );
  DFF_X2 \u6/rem_reg[13]  ( .D(\u6/remainder [13]), .CK(clk), .QN(n3058) );
  DFF_X2 \u6/remainder_reg[14]  ( .D(\u6/N14 ), .CK(clk), .Q(
        \u6/remainder [14]) );
  DFF_X2 \u6/rem_reg[14]  ( .D(\u6/remainder [14]), .CK(clk), .QN(n3057) );
  DFF_X2 \u6/remainder_reg[15]  ( .D(\u6/N15 ), .CK(clk), .Q(
        \u6/remainder [15]) );
  DFF_X2 \u6/rem_reg[15]  ( .D(\u6/remainder [15]), .CK(clk), .QN(n1566) );
  DFF_X2 \u6/remainder_reg[16]  ( .D(\u6/N16 ), .CK(clk), .Q(
        \u6/remainder [16]) );
  DFF_X2 \u6/rem_reg[16]  ( .D(\u6/remainder [16]), .CK(clk), .QN(n1585) );
  DFF_X2 \u6/remainder_reg[17]  ( .D(\u6/N17 ), .CK(clk), .Q(
        \u6/remainder [17]) );
  DFF_X2 \u6/rem_reg[17]  ( .D(\u6/remainder [17]), .CK(clk), .QN(n1618) );
  DFF_X2 \u6/remainder_reg[18]  ( .D(\u6/N18 ), .CK(clk), .Q(
        \u6/remainder [18]) );
  DFF_X2 \u6/rem_reg[18]  ( .D(\u6/remainder [18]), .CK(clk), .QN(n3056) );
  DFF_X2 \u6/remainder_reg[19]  ( .D(\u6/N19 ), .CK(clk), .Q(
        \u6/remainder [19]) );
  DFF_X2 \u6/rem_reg[19]  ( .D(\u6/remainder [19]), .CK(clk), .QN(n3055) );
  DFF_X2 \u6/remainder_reg[20]  ( .D(\u6/N20 ), .CK(clk), .Q(
        \u6/remainder [20]) );
  DFF_X2 \u6/rem_reg[20]  ( .D(\u6/remainder [20]), .CK(clk), .QN(n1567) );
  DFF_X2 \u6/remainder_reg[21]  ( .D(\u6/N21 ), .CK(clk), .Q(
        \u6/remainder [21]) );
  DFF_X2 \u6/rem_reg[21]  ( .D(\u6/remainder [21]), .CK(clk), .QN(n1586) );
  DFF_X2 \u6/remainder_reg[22]  ( .D(\u6/N22 ), .CK(clk), .Q(
        \u6/remainder [22]) );
  DFF_X2 \u6/rem_reg[22]  ( .D(\u6/remainder [22]), .CK(clk), .QN(n1619) );
  DFF_X2 \u6/remainder_reg[23]  ( .D(\u6/N23 ), .CK(clk), .Q(
        \u6/remainder [23]) );
  DFF_X2 \u6/rem_reg[23]  ( .D(\u6/remainder [23]), .CK(clk), .QN(n3054) );
  DFF_X2 \u6/quo1_reg[0]  ( .D(\u6/N0 ), .CK(clk), .Q(\u6/quo1 [0]) );
  DFF_X2 \u6/quo_reg[0]  ( .D(\u6/quo1 [0]), .CK(clk), .Q(quo[0]) );
  DFF_X2 \u6/quo1_reg[1]  ( .D(\u6/N1 ), .CK(clk), .Q(\u6/quo1 [1]) );
  DFF_X2 \u6/quo_reg[1]  ( .D(\u6/quo1 [1]), .CK(clk), .Q(quo[1]) );
  DFF_X2 \u6/quo1_reg[2]  ( .D(\u6/N2 ), .CK(clk), .Q(\u6/quo1 [2]) );
  DFF_X2 \u6/quo_reg[2]  ( .D(\u6/quo1 [2]), .CK(clk), .Q(quo[2]), .QN(n1642)
         );
  DFF_X2 \u6/quo1_reg[3]  ( .D(\u6/N3 ), .CK(clk), .Q(\u6/quo1 [3]) );
  DFF_X2 \u6/quo_reg[3]  ( .D(\u6/quo1 [3]), .CK(clk), .Q(quo[3]) );
  DFF_X2 \u6/quo1_reg[4]  ( .D(\u6/N4 ), .CK(clk), .Q(\u6/quo1 [4]) );
  DFF_X2 \u6/quo_reg[4]  ( .D(\u6/quo1 [4]), .CK(clk), .Q(quo[4]) );
  DFF_X2 \u6/quo1_reg[5]  ( .D(\u6/N5 ), .CK(clk), .Q(\u6/quo1 [5]) );
  DFF_X2 \u6/quo_reg[5]  ( .D(\u6/quo1 [5]), .CK(clk), .Q(quo[5]), .QN(n1650)
         );
  DFF_X2 \u6/quo1_reg[6]  ( .D(\u6/N6 ), .CK(clk), .Q(\u6/quo1 [6]) );
  DFF_X2 \u6/quo_reg[6]  ( .D(\u6/quo1 [6]), .CK(clk), .Q(quo[6]) );
  DFF_X2 \u6/quo1_reg[7]  ( .D(\u6/N7 ), .CK(clk), .Q(\u6/quo1 [7]) );
  DFF_X2 \u6/quo_reg[7]  ( .D(\u6/quo1 [7]), .CK(clk), .Q(quo[7]) );
  DFF_X2 \u6/quo1_reg[8]  ( .D(\u6/N8 ), .CK(clk), .Q(\u6/quo1 [8]) );
  DFF_X2 \u6/quo_reg[8]  ( .D(\u6/quo1 [8]), .CK(clk), .Q(quo[8]) );
  DFF_X2 \u6/quo1_reg[9]  ( .D(\u6/N9 ), .CK(clk), .Q(\u6/quo1 [9]) );
  DFF_X2 \u6/quo_reg[9]  ( .D(\u6/quo1 [9]), .CK(clk), .Q(quo[9]), .QN(n1937)
         );
  DFF_X2 \u6/quo1_reg[10]  ( .D(n1731), .CK(clk), .Q(\u6/quo1 [10]) );
  DFF_X2 \u6/quo_reg[10]  ( .D(\u6/quo1 [10]), .CK(clk), .Q(quo[10]) );
  DFF_X2 \u6/quo1_reg[13]  ( .D(\u6/N13 ), .CK(clk), .Q(\u6/quo1 [13]) );
  DFF_X2 \u6/quo_reg[13]  ( .D(\u6/quo1 [13]), .CK(clk), .Q(quo[13]), .QN(
        net86061) );
  DFF_X2 \u6/quo1_reg[14]  ( .D(\u6/N14 ), .CK(clk), .Q(\u6/quo1 [14]) );
  DFF_X2 \u6/quo_reg[14]  ( .D(\u6/quo1 [14]), .CK(clk), .Q(quo[14]) );
  DFF_X2 \u6/quo1_reg[15]  ( .D(\u6/N15 ), .CK(clk), .Q(\u6/quo1 [15]) );
  DFF_X2 \u6/quo_reg[15]  ( .D(\u6/quo1 [15]), .CK(clk), .Q(quo[15]) );
  DFF_X2 \u6/quo1_reg[16]  ( .D(\u6/N16 ), .CK(clk), .Q(\u6/quo1 [16]) );
  DFF_X2 \u6/quo_reg[16]  ( .D(\u6/quo1 [16]), .CK(clk), .Q(quo[16]) );
  DFF_X2 \u6/quo1_reg[17]  ( .D(\u6/N17 ), .CK(clk), .Q(\u6/quo1 [17]) );
  DFF_X2 \u6/quo_reg[17]  ( .D(\u6/quo1 [17]), .CK(clk), .Q(quo[17]) );
  DFF_X2 \u6/quo1_reg[18]  ( .D(\u6/N18 ), .CK(clk), .Q(\u6/quo1 [18]) );
  DFF_X2 \u6/quo_reg[18]  ( .D(\u6/quo1 [18]), .CK(clk), .Q(quo[18]) );
  DFF_X2 \u6/quo1_reg[19]  ( .D(\u6/N19 ), .CK(clk), .Q(\u6/quo1 [19]) );
  DFF_X2 \u6/quo_reg[19]  ( .D(\u6/quo1 [19]), .CK(clk), .Q(quo[19]) );
  DFF_X2 \u6/quo1_reg[20]  ( .D(\u6/N20 ), .CK(clk), .Q(\u6/quo1 [20]) );
  DFF_X2 \u6/quo_reg[20]  ( .D(\u6/quo1 [20]), .CK(clk), .Q(quo[20]) );
  DFF_X2 \u6/quo1_reg[21]  ( .D(\u6/N21 ), .CK(clk), .Q(\u6/quo1 [21]) );
  DFF_X2 \u6/quo_reg[21]  ( .D(\u6/quo1 [21]), .CK(clk), .Q(quo[21]) );
  DFF_X2 \u6/quo1_reg[22]  ( .D(\u6/N22 ), .CK(clk), .Q(\u6/quo1 [22]) );
  DFF_X2 \u6/quo_reg[22]  ( .D(\u6/quo1 [22]), .CK(clk), .Q(quo[22]) );
  DFF_X2 \out_reg[13]  ( .D(N233), .CK(clk), .Q(out[13]) );
  DFF_X2 \out_reg[14]  ( .D(N234), .CK(clk), .Q(out[14]) );
  DFF_X2 \u6/quo1_reg[23]  ( .D(\u6/N23 ), .CK(clk), .Q(\u6/quo1 [23]) );
  DFF_X2 \u6/quo_reg[23]  ( .D(\u6/quo1 [23]), .CK(clk), .QN(net11485) );
  fpu_DW01_ash_1 \u4/sll_479  ( .A({net85786, net85786, net85786, net85786, 
        net85786, net85786, net85786, net85786, net85786, net86263, net77045, 
        net77161, n3003, net76254, net89624, n3002, n3004, net76672, n3005, 
        fract_denorm, net76926, net77073, net77637, net90292, net10316, n3001, 
        net76048, net90080, n3319}), .DATA_TC(1'b0), .SH({\u4/f2i_shft[4] , 
        \u4/f2i_shft[3] , \u4/f2i_shft[2] , net85710, net11564}), .SH_TC(1'b0), 
        .B({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, \u4/exp_f2i_1 , 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24}) );
  fpu_DW01_sub_7 \u3/sub_59  ( .A({1'b0, fracta}), .B({1'b0, fractb}), .CI(
        1'b0), .DIFF({\u3/N32 , \u3/N31 , \u3/N30 , \u3/N29 , \u3/N28 , 
        \u3/N27 , \u3/N26 , \u3/N25 , \u3/N24 , \u3/N23 , \u3/N22 , \u3/N21 , 
        \u3/N20 , \u3/N19 , \u3/N18 }) );
  fpu_DW01_add_5 \u3/add_59  ( .A({1'b0, fracta}), .B({1'b0, fractb}), .CI(
        1'b0), .SUM({\u3/N17 , \u3/N16 , \u3/N15 , \u3/N14 , \u3/N13 , 
        \u3/N12 , \u3/N11 , \u3/N10 , \u3/N9 , \u3/N8 , \u3/N7 , \u3/N6 , 
        \u3/N5 , \u3/N4 , \u3/N3 }) );
  fpu_DW01_ash_2 sll_385 ( .A({n3313, fracta_mul}), .DATA_TC(1'b0), .SH({N34, 
        N44, N56, N65}), .SH_TC(1'b0), .B({N77, N76, N75, N74, N73, N72, N71, 
        N70, N69, N68, N67}) );
  fpu_DW02_mult_0 \u5/mult_78  ( .A({n3313, fracta_mul[9:3], n2848, n3014, 
        n3015}), .B({\u6/N10 , \u6/N9 , \u6/N8 , \u6/N7 , \u6/N6 , \u6/N5 , 
        \u6/N4 , \u6/N3 , \u6/N2 , \u6/N1 , \u6/N0 }), .TC(1'b0), .PRODUCT({
        \u5/N21 , \u5/N20 , \u5/N19 , \u5/N18 , \u5/N17 , \u5/N16 , \u5/N15 , 
        \u5/N14 , \u5/N13 , \u5/N12 , \u5/N11 , \u5/N10 , \u5/N9 , \u5/N8 , 
        \u5/N7 , \u5/N6 , \u5/N5 , \u5/N4 , \u5/N3 , \u5/N2 , \u5/N1 , \u5/N0 }) );
  HA_X1 \u2/add_115/U1_1_1  ( .A(\u2/exp_tmp4[1] ), .B(\u2/exp_tmp4[0] ), .CO(
        \u2/add_115/carry [2]), .S(\u2/N31 ) );
  HA_X1 \u2/add_115/U1_1_2  ( .A(\u2/exp_tmp4[2] ), .B(\u2/add_115/carry [2]), 
        .CO(\u2/add_115/carry [3]), .S(\u2/N32 ) );
  HA_X1 \u2/add_115/U1_1_3  ( .A(\u2/exp_tmp4[3] ), .B(\u2/add_115/carry [3]), 
        .CO(\u2/add_115/carry [4]), .S(\u2/N33 ) );
  HA_X1 \u2/add_113/U1_1_1  ( .A(\u2/add_113/A[1] ), .B(\u2/add_113/A[0] ), 
        .CO(\u2/add_113/carry [2]), .S(\u2/exp_tmp3[1] ) );
  HA_X1 \u2/add_113/U1_1_2  ( .A(\u2/add_113/A[2] ), .B(\u2/add_113/carry [2]), 
        .CO(\u2/add_113/carry [3]), .S(\u2/exp_tmp3[2] ) );
  HA_X1 \u2/add_113/U1_1_3  ( .A(\u2/add_113/A[3] ), .B(\u2/add_113/carry [3]), 
        .CO(\u2/add_113/carry [4]), .S(\u2/exp_tmp3[3] ) );
  FA_X1 \u2/add_110/U1_1  ( .A(opa_r[11]), .B(opb_r[11]), .CI(
        \u2/add_110/carry [1]), .CO(\u2/add_110/carry [2]), .S(\u2/N13 ) );
  FA_X1 \u2/add_110/U1_2  ( .A(opa_r[12]), .B(opb_r[12]), .CI(
        \u2/add_110/carry [2]), .CO(\u2/add_110/carry [3]), .S(\u2/N14 ) );
  FA_X1 \u2/add_110/U1_3  ( .A(opa_r[13]), .B(opb_r[13]), .CI(
        \u2/add_110/carry [3]), .CO(\u2/add_110/carry [4]), .S(\u2/N15 ) );
  FA_X1 \u2/add_110/U1_4  ( .A(opa_r[14]), .B(n1733), .CI(
        \u2/add_110/carry [4]), .CO(\u2/N17 ), .S(\u2/N16 ) );
  FA_X1 \u2/sub_110/U2_1  ( .A(opa_r[11]), .B(n3016), .CI(
        \u2/sub_110/carry [1]), .CO(\u2/sub_110/carry [2]), .S(\u2/N7 ) );
  FA_X1 \u2/sub_110/U2_2  ( .A(opa_r[12]), .B(n2799), .CI(
        \u2/sub_110/carry [2]), .CO(\u2/sub_110/carry [3]), .S(\u2/N8 ) );
  FA_X1 \u2/sub_110/U2_3  ( .A(opa_r[13]), .B(n3017), .CI(
        \u2/sub_110/carry [3]), .CO(\u2/sub_110/carry [4]), .S(\u2/N9 ) );
  FA_X1 \u2/sub_110/U2_4  ( .A(opa_r[14]), .B(n1541), .CI(
        \u2/sub_110/carry [4]), .CO(\u2/sub_110/carry [5]), .S(\u2/N10 ) );
  fpu_DW01_inc_5 \u4/add_393  ( .A({1'b0, net91299, net90252, 
        \u4/fract_out[7] , net91512, n1528, net89933, net99874, n3006, n1920, 
        net60630}), .SUM({\u4/fract_out_pl1[10] , \u4/fract_out_pl1[9] , 
        \u4/fract_out_pl1[8] , \u4/fract_out_pl1[7] , \u4/fract_out_pl1[6] , 
        \u4/fract_out_pl1[5] , \u4/fract_out_pl1[4] , \u4/fract_out_pl1[3] , 
        \u4/fract_out_pl1[2] , \u4/fract_out_pl1[1] , \u4/fract_out_pl1[0] })
         );
  fpu_DW_rash_2 \u4/srl_450  ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, net85786, net86263, net91070, net90115, n3003, 
        net86004, net89624, n3002, n3004, net90007, n3005, fract_denorm[10], 
        net90211, net90037, n1883, net90290, n2998, net10316, n3001, n2999, 
        n1926, n3319}), .DATA_TC(1'b0), .SH(\u4/shift_right [2:0]), .SH_TC(
        1'b0), .B({SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, \u4/N409 , 
        \u4/N408 , \u4/N407 , \u4/N406 , \u4/N405 , \u4/N404 , \u4/N403 , 
        \u4/N402 , \u4/N401 , \u4/N400 , \u4/N399 , \u4/N398 , \u4/N397 , 
        \u4/N396 , \u4/N395 , \u4/N394 , \u4/N393 , \u4/N392 , \u4/N391 , 
        \u4/N390 , \u4/N389 , \u4/N388 }) );
  fpu_DW01_ash_4 \u4/sll_451  ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, net85786, net86263, net91070, net90115, n3003, 
        net86004, net89624, n3002, n3004, net90007, n3005, fract_denorm[10], 
        net90211, net90037, n1883, net90290, n2998, net10316, n3001, n2999, 
        n3000, n3319}), .DATA_TC(1'b0), .SH(\u4/shift_left ), .SH_TC(1'b0), 
        .B({SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, \u4/N433 , 
        \u4/N432 , \u4/N431 , \u4/N430 , \u4/N429 , \u4/N428 , \u4/N427 , 
        \u4/N426 , \u4/N425 , \u4/N424 , \u4/N423 , \u4/N422 , \u4/N421 , 
        \u4/N420 , \u4/N419 , \u4/N418 , \u4/N417 , \u4/N416 , \u4/N415 , 
        \u4/N414 , \u4/N413 , \u4/N412 }) );
  fpu_DW01_sub_23 \u4/sub_467  ( .A({1'b0, \u4/exp_in_pl1[5] , 
        \u4/exp_in_pl1[4] , \u4/exp_in_pl1[3] , \u4/exp_in_pl1[2] , net85712, 
        net15448}), .B({1'b0, 1'b0, n3008, \u4/fi_ldz_mi1[3] , 
        \u4/fi_ldz_mi1[2] , net33278, net89965}), .CI(1'b0), .DIFF({
        SYNOPSYS_UNCONNECTED__45, \u4/exp_next_mi[5] , \u4/exp_next_mi[4] , 
        \u4/exp_next_mi[3] , \u4/exp_next_mi[2] , \u4/exp_next_mi[1] , 
        \u4/exp_next_mi[0] }) );
  fpu_DW_rash_11 \u1/srl_146  ( .A({n1521, \u1/adj_op[9] , n3303, n3304, n3305, 
        n3306, n3307, n3308, n3309, n3310, n3311, 1'b0, 1'b0, 1'b0}), 
        .DATA_TC(1'b0), .SH({n3302, n3301, n3300, n1718}), .SH_TC(1'b0), .B({
        \u1/adj_op_out_sft[13] , \u1/adj_op_out_sft[12] , 
        \u1/adj_op_out_sft[11] , \u1/adj_op_out_sft[10] , 
        \u1/adj_op_out_sft[9] , \u1/adj_op_out_sft[8] , \u1/adj_op_out_sft[7] , 
        \u1/adj_op_out_sft[6] , \u1/adj_op_out_sft[5] , \u1/adj_op_out_sft[4] , 
        \u1/adj_op_out_sft[3] , \u1/adj_op_out_sft[2] , \u1/adj_op_out_sft[1] , 
        \u1/adj_op_out_sft[0] }) );
  DFF_X1 inf_reg ( .D(N285), .CK(clk), .Q(inf) );
  DFF_X1 \out_reg[4]  ( .D(N224), .CK(clk), .Q(out[4]) );
  DFF_X1 \out_reg[3]  ( .D(N223), .CK(clk), .Q(out[3]) );
  DFF_X1 \out_reg[2]  ( .D(N222), .CK(clk), .Q(out[2]) );
  DFF_X1 \out_reg[1]  ( .D(N221), .CK(clk), .Q(out[1]) );
  DFF_X1 \out_reg[5]  ( .D(N225), .CK(clk), .Q(out[5]) );
  DFF_X1 zero_reg ( .D(N290), .CK(clk), .Q(zero) );
  DFF_X1 ine_reg ( .D(n3007), .CK(clk), .Q(ine) );
  DFF_X1 underflow_reg ( .D(N281), .CK(clk), .Q(underflow) );
  DFF_X1 \out_reg[15]  ( .D(N254), .CK(clk), .Q(out[15]) );
  DFF_X2 \fract_i2f_reg[9]  ( .D(N184), .CK(clk), .QN(net90064) );
  DFF_X1 overflow_reg ( .D(N278), .CK(clk), .Q(overflow) );
  DFF_X1 \out_reg[6]  ( .D(N226), .CK(clk), .Q(out[6]) );
  DFF_X1 \out_reg[7]  ( .D(N227), .CK(clk), .Q(out[7]) );
  DFF_X1 \out_reg[8]  ( .D(N228), .CK(clk), .Q(out[8]) );
  DFF_X1 \out_reg[9]  ( .D(N229), .CK(clk), .Q(out[9]) );
  DFF_X1 \out_reg[12]  ( .D(N232), .CK(clk), .Q(out[12]) );
  DFF_X1 \u5/prod1_reg[13]  ( .D(\u5/N13 ), .CK(clk), .Q(\u5/prod1 [13]) );
  DFF_X1 \u5/prod1_reg[11]  ( .D(\u5/N11 ), .CK(clk), .Q(\u5/prod1 [11]) );
  DFF_X1 \u1/fracta_out_reg[5]  ( .D(\u1/fracta_s [5]), .CK(clk), .Q(fracta[5]) );
  DFF_X1 \u1/fractb_out_reg[13]  ( .D(\u1/fractb_s [13]), .CK(clk), .Q(
        fractb[13]) );
  DFF_X1 \u1/fractb_out_reg[10]  ( .D(\u1/fractb_s [10]), .CK(clk), .Q(
        fractb[10]) );
  DFF_X1 \u1/fractb_out_reg[6]  ( .D(\u1/fractb_s [6]), .CK(clk), .Q(fractb[6]) );
  DFF_X1 \u1/fractb_out_reg[9]  ( .D(\u1/fractb_s [9]), .CK(clk), .Q(fractb[9]) );
  DFF_X1 \u1/fractb_out_reg[11]  ( .D(\u1/fractb_s [11]), .CK(clk), .Q(
        fractb[11]) );
  DFF_X1 \u1/fracta_out_reg[1]  ( .D(\u1/fracta_s [1]), .CK(clk), .Q(fracta[1]) );
  DFF_X1 \u1/fractb_out_reg[8]  ( .D(\u1/fractb_s [8]), .CK(clk), .Q(fractb[8]) );
  DFF_X1 \u1/fracta_out_reg[6]  ( .D(\u1/fracta_s [6]), .CK(clk), .Q(fracta[6]) );
  DFF_X1 \u1/fractb_out_reg[5]  ( .D(\u1/fractb_s [5]), .CK(clk), .Q(fractb[5]) );
  DFF_X1 \u1/fractb_out_reg[2]  ( .D(\u1/fractb_s [2]), .CK(clk), .Q(fractb[2]) );
  DFF_X1 \u1/fractb_out_reg[1]  ( .D(\u1/fractb_s [1]), .CK(clk), .Q(fractb[1]) );
  DFF_X1 \u1/fractb_out_reg[7]  ( .D(\u1/fractb_s [7]), .CK(clk), .Q(fractb[7]) );
  DFF_X1 \u1/fractb_out_reg[3]  ( .D(\u1/fractb_s [3]), .CK(clk), .Q(fractb[3]) );
  DFF_X1 \u1/sign_reg  ( .D(\u1/sign_d ), .CK(clk), .Q(sign_fasu) );
  DFF_X1 \u1/fracta_out_reg[9]  ( .D(\u1/fracta_s [9]), .CK(clk), .Q(fracta[9]) );
  DFF_X1 \u1/fracta_out_reg[10]  ( .D(\u1/fracta_s [10]), .CK(clk), .Q(
        fracta[10]) );
  DFF_X1 \u1/fracta_out_reg[12]  ( .D(\u1/fracta_s [12]), .CK(clk), .Q(
        fracta[12]) );
  DFF_X1 \u1/fracta_out_reg[8]  ( .D(\u1/fracta_s [8]), .CK(clk), .Q(fracta[8]) );
  DFF_X1 \u1/fractb_out_reg[12]  ( .D(\u1/fractb_s [12]), .CK(clk), .Q(
        fractb[12]) );
  DFF_X1 \u1/fracta_out_reg[11]  ( .D(\u1/fracta_s [11]), .CK(clk), .Q(
        fracta[11]) );
  DFF_X1 \u1/fracta_out_reg[7]  ( .D(\u1/fracta_s [7]), .CK(clk), .Q(fracta[7]) );
  DFF_X1 \fract_out_q_reg[14]  ( .D(n3284), .CK(clk), .Q(fract_out_q[14]) );
  DFF_X1 \u5/prod1_reg[10]  ( .D(\u5/N10 ), .CK(clk), .Q(\u5/prod1 [10]) );
  DFF_X1 \fract_out_q_reg[11]  ( .D(n3287), .CK(clk), .Q(fract_out_q[11]) );
  DFF_X1 \fract_out_q_reg[10]  ( .D(n3288), .CK(clk), .Q(fract_out_q[10]) );
  DFF_X1 \u5/prod1_reg[8]  ( .D(\u5/N8 ), .CK(clk), .Q(\u5/prod1 [8]) );
  DFF_X1 \fract_i2f_reg[2]  ( .D(n3282), .CK(clk), .Q(n1668) );
  DFF_X1 \fract_i2f_reg[15]  ( .D(N190), .CK(clk), .Q(n1667) );
  DFF_X1 \fract_i2f_reg[0]  ( .D(n3318), .CK(clk), .Q(n1660) );
  DFF_X1 \fract_i2f_reg[11]  ( .D(N186), .CK(clk), .Q(n1659) );
  DFF_X1 \fract_i2f_reg[12]  ( .D(N187), .CK(clk), .Q(n1658) );
  DFF_X1 \fract_i2f_reg[6]  ( .D(N181), .CK(clk), .Q(n1657) );
  DFF_X1 \fract_out_q_reg[0]  ( .D(n3298), .CK(clk), .Q(n1656) );
  DFF_X1 \fract_i2f_reg[5]  ( .D(N180), .CK(clk), .Q(n1652) );
  DFF_X1 \fract_i2f_reg[21]  ( .D(N196), .CK(clk), .Q(n1643) );
  DFF_X1 \fract_i2f_reg[17]  ( .D(N192), .CK(clk), .Q(n1634) );
  DFF_X1 \fract_i2f_reg[19]  ( .D(N194), .CK(clk), .Q(n1633) );
  DFF_X1 \out_reg[0]  ( .D(N220), .CK(clk), .Q(out[0]) );
  DFF_X1 \out_reg[11]  ( .D(N231), .CK(clk), .Q(out[11]) );
  DFF_X1 \out_reg[10]  ( .D(N230), .CK(clk), .Q(out[10]) );
  DFF_X1 \u5/prod1_reg[17]  ( .D(\u5/N17 ), .CK(clk), .Q(\u5/prod1 [17]) );
  DFF_X2 \u1/fractb_out_reg[0]  ( .D(\u1/fractb_s [0]), .CK(clk), .Q(fractb[0]) );
  DFF_X1 \fract_out_q_reg[12]  ( .D(n3286), .CK(clk), .Q(fract_out_q[12]) );
  INV_X4 U1188 ( .A(net85292), .ZN(net90110) );
  INV_X4 U1189 ( .A(net85292), .ZN(net85160) );
  INV_X4 U1190 ( .A(net85263), .ZN(net85357) );
  NAND4_X2 U1191 ( .A1(net85260), .A2(n1743), .A3(net85263), .A4(1'b1), .ZN(
        net85187) );
  NAND2_X2 U1192 ( .A1(net85349), .A2(n1839), .ZN(n1838) );
  NAND2_X2 U1193 ( .A1(n3058), .A2(n3057), .ZN(n2177) );
  NAND2_X2 U1194 ( .A1(n1616), .A2(n1584), .ZN(n2173) );
  INV_X4 U1195 ( .A(net83963), .ZN(n2213) );
  INV_X4 U1196 ( .A(exp_r[4]), .ZN(n2115) );
  NAND2_X2 U1197 ( .A1(fract_out_q[13]), .A2(net83780), .ZN(net91059) );
  NAND2_X2 U1198 ( .A1(net83780), .A2(fract_out_q[13]), .ZN(net85247) );
  INV_X4 U1199 ( .A(exp_r[4]), .ZN(n2288) );
  INV_X4 U1200 ( .A(net91112), .ZN(n2200) );
  NAND2_X2 U1201 ( .A1(n2214), .A2(n2213), .ZN(net84722) );
  OAI211_X2 U1202 ( .C1(n2117), .C2(1'b0), .A(n2115), .B(n2114), .ZN(n2634) );
  NOR2_X1 U1203 ( .A1(n2099), .A2(n1527), .ZN(n1524) );
  NOR2_X2 U1204 ( .A1(n1524), .A2(n1525), .ZN(n1552) );
  AND2_X2 U1205 ( .A1(n1526), .A2(n1549), .ZN(n1525) );
  INV_X4 U1206 ( .A(n1825), .ZN(n1526) );
  OR2_X4 U1207 ( .A1(net88293), .A2(n1825), .ZN(n1527) );
  OAI21_X4 U1208 ( .B1(net84778), .B2(n2161), .A(n2160), .ZN(n1528) );
  INV_X8 U1209 ( .A(\u4/fract_out[6] ), .ZN(net84113) );
  INV_X8 U1210 ( .A(net91299), .ZN(net84118) );
  INV_X2 U1211 ( .A(n1752), .ZN(net91298) );
  NOR2_X4 U1212 ( .A1(\u4/fract_out[1] ), .A2(\u4/fract_out[4] ), .ZN(n1798)
         );
  NAND2_X4 U1213 ( .A1(n1873), .A2(net83959), .ZN(n1745) );
  NAND2_X2 U1214 ( .A1(net84069), .A2(net84070), .ZN(net84055) );
  NAND2_X2 U1215 ( .A1(net84071), .A2(net84072), .ZN(net83860) );
  INV_X2 U1216 ( .A(net83860), .ZN(net84070) );
  OAI21_X2 U1217 ( .B1(n2627), .B2(net83860), .A(net83861), .ZN(n2708) );
  INV_X2 U1218 ( .A(n2453), .ZN(n2455) );
  AOI21_X2 U1219 ( .B1(n2695), .B2(n2694), .A(n2615), .ZN(n2616) );
  OAI21_X4 U1220 ( .B1(net84575), .B2(net84574), .A(net84576), .ZN(n1529) );
  OAI21_X2 U1221 ( .B1(net84575), .B2(net84574), .A(net84576), .ZN(net91511)
         );
  OAI211_X2 U1222 ( .C1(net91015), .C2(net85018), .A(net85020), .B(net85021), 
        .ZN(n1530) );
  NOR2_X2 U1223 ( .A1(net84374), .A2(net84373), .ZN(n1536) );
  INV_X1 U1224 ( .A(n2625), .ZN(n1531) );
  INV_X2 U1225 ( .A(net84373), .ZN(n1532) );
  INV_X4 U1226 ( .A(n1532), .ZN(n1533) );
  NOR3_X2 U1227 ( .A1(n2359), .A2(n2360), .A3(n1597), .ZN(net84373) );
  INV_X2 U1228 ( .A(n1749), .ZN(n1534) );
  INV_X2 U1229 ( .A(n1534), .ZN(n1535) );
  NOR2_X4 U1230 ( .A1(net84372), .A2(n1537), .ZN(net86174) );
  INV_X4 U1231 ( .A(n1536), .ZN(n1537) );
  INV_X4 U1232 ( .A(n2926), .ZN(n2924) );
  NAND2_X4 U1233 ( .A1(opa_r[12]), .A2(n2799), .ZN(n2773) );
  INV_X4 U1234 ( .A(n2809), .ZN(n1539) );
  INV_X2 U1235 ( .A(n2817), .ZN(n2806) );
  OAI21_X2 U1236 ( .B1(n2820), .B2(n2818), .A(n2817), .ZN(n2822) );
  AOI211_X4 U1237 ( .C1(n2894), .C2(n2893), .A(n2892), .B(n2891), .ZN(n2903)
         );
  NOR2_X1 U1238 ( .A1(opa_r[14]), .A2(opb_r[14]), .ZN(n2815) );
  NOR2_X2 U1239 ( .A1(\u1/adj_op_out_sft[13] ), .A2(n2791), .ZN(n2928) );
  NOR2_X1 U1240 ( .A1(opa_r[13]), .A2(opa_r[14]), .ZN(n1984) );
  INV_X4 U1241 ( .A(n1733), .ZN(n1541) );
  NAND2_X4 U1242 ( .A1(n1734), .A2(n1730), .ZN(n1729) );
  BUF_X32 U1243 ( .A(n1728), .Z(n1543) );
  AND2_X2 U1244 ( .A1(fracta_mul[0]), .A2(n3045), .ZN(n3022) );
  OAI21_X4 U1245 ( .B1(net84211), .B2(n2339), .A(net91542), .ZN(net84169) );
  NAND2_X4 U1246 ( .A1(n2527), .A2(n2526), .ZN(net84060) );
  INV_X2 U1247 ( .A(net83736), .ZN(net83856) );
  NAND2_X4 U1248 ( .A1(net83871), .A2(n1736), .ZN(N230) );
  NAND2_X4 U1249 ( .A1(n2457), .A2(n2458), .ZN(n2520) );
  NAND2_X2 U1250 ( .A1(n2433), .A2(n2707), .ZN(N234) );
  BUF_X4 U1251 ( .A(net83765), .Z(n1546) );
  INV_X8 U1252 ( .A(net83765), .ZN(net83800) );
  INV_X8 U1253 ( .A(n2460), .ZN(n2528) );
  NAND3_X4 U1254 ( .A1(n1832), .A2(net84253), .A3(net84254), .ZN(net84096) );
  AOI21_X4 U1255 ( .B1(n2705), .B2(n2704), .A(n2703), .ZN(N278) );
  INV_X8 U1256 ( .A(n2618), .ZN(n2656) );
  AND3_X2 U1257 ( .A1(n2656), .A2(n1742), .A3(net83806), .ZN(N290) );
  BUF_X32 U1258 ( .A(n1751), .Z(n1548) );
  INV_X8 U1259 ( .A(net84138), .ZN(net84211) );
  OAI21_X1 U1260 ( .B1(n1548), .B2(net83429), .A(n2963), .ZN(n3010) );
  NAND2_X4 U1261 ( .A1(n1746), .A2(net84472), .ZN(n1597) );
  INV_X2 U1262 ( .A(n1747), .ZN(n1746) );
  OAI211_X1 U1263 ( .C1(n1554), .C2(net84312), .A(net85842), .B(net84133), 
        .ZN(n1842) );
  NAND4_X1 U1264 ( .A1(net91511), .A2(n1749), .A3(net84128), .A4(n1580), .ZN(
        n2359) );
  INV_X16 U1265 ( .A(net85853), .ZN(net86067) );
  NAND2_X4 U1266 ( .A1(net85317), .A2(net86067), .ZN(n1878) );
  INV_X8 U1267 ( .A(n2065), .ZN(n2043) );
  AOI22_X4 U1268 ( .A1(net89998), .A2(n1609), .B1(net85077), .B2(prod[20]), 
        .ZN(net90019) );
  NAND2_X4 U1269 ( .A1(n1896), .A2(net85071), .ZN(net90080) );
  NOR2_X4 U1270 ( .A1(net85752), .A2(net85730), .ZN(n2015) );
  INV_X4 U1271 ( .A(net77637), .ZN(net84910) );
  INV_X8 U1272 ( .A(net84910), .ZN(net90290) );
  INV_X8 U1273 ( .A(net85331), .ZN(net85203) );
  OR2_X4 U1274 ( .A1(net85832), .A2(net86037), .ZN(n1549) );
  AND2_X2 U1275 ( .A1(n2653), .A2(net86038), .ZN(n1550) );
  AND2_X4 U1276 ( .A1(net85107), .A2(net85108), .ZN(n1551) );
  INV_X8 U1277 ( .A(n2139), .ZN(n1940) );
  OAI21_X4 U1278 ( .B1(net84754), .B2(net84755), .A(n1905), .ZN(n1761) );
  INV_X1 U1279 ( .A(net83945), .ZN(net84672) );
  INV_X2 U1280 ( .A(net84672), .ZN(net88500) );
  INV_X16 U1281 ( .A(net91404), .ZN(net84150) );
  INV_X8 U1282 ( .A(net84995), .ZN(net85015) );
  INV_X8 U1283 ( .A(net84994), .ZN(net89753) );
  AND2_X2 U1284 ( .A1(net83959), .A2(n1593), .ZN(n1553) );
  INV_X8 U1285 ( .A(net91298), .ZN(net91299) );
  NAND2_X4 U1286 ( .A1(net84366), .A2(net84453), .ZN(n2437) );
  AND2_X4 U1287 ( .A1(net84474), .A2(net84475), .ZN(n1554) );
  AND2_X2 U1288 ( .A1(n1754), .A2(n2170), .ZN(n1555) );
  NAND2_X4 U1289 ( .A1(net84133), .A2(n2437), .ZN(n2490) );
  INV_X16 U1290 ( .A(net84135), .ZN(net84133) );
  INV_X1 U1291 ( .A(net83875), .ZN(net84085) );
  NAND2_X4 U1292 ( .A1(net84136), .A2(rmode_r3[1]), .ZN(n2496) );
  AOI21_X4 U1293 ( .B1(net86174), .B2(net84075), .A(net84206), .ZN(net84204)
         );
  NAND2_X1 U1294 ( .A1(net89856), .A2(net85041), .ZN(net10316) );
  INV_X16 U1295 ( .A(net85097), .ZN(net85089) );
  NAND2_X4 U1296 ( .A1(net84757), .A2(net84758), .ZN(net91555) );
  NAND2_X2 U1297 ( .A1(net84757), .A2(net84758), .ZN(net84301) );
  NAND3_X2 U1298 ( .A1(net85730), .A2(net85716), .A3(fract_out_q[4]), .ZN(
        n2068) );
  NOR2_X4 U1299 ( .A1(net11576), .A2(net85718), .ZN(n1556) );
  NAND3_X2 U1300 ( .A1(n2070), .A2(n2068), .A3(n2069), .ZN(net85197) );
  INV_X4 U1301 ( .A(n2070), .ZN(n2071) );
  NAND2_X2 U1302 ( .A1(net85144), .A2(n2053), .ZN(n1954) );
  OAI21_X1 U1303 ( .B1(n2055), .B2(net89677), .A(net85105), .ZN(n2057) );
  INV_X8 U1304 ( .A(n1912), .ZN(n1909) );
  AND2_X4 U1305 ( .A1(net86090), .A2(n1893), .ZN(n1891) );
  INV_X16 U1306 ( .A(net85010), .ZN(net83959) );
  BUF_X16 U1307 ( .A(net85095), .Z(net89078) );
  NOR2_X4 U1308 ( .A1(\u4/N656 ), .A2(n1571), .ZN(net85010) );
  BUF_X16 U1309 ( .A(net84609), .Z(net90122) );
  INV_X8 U1310 ( .A(n1792), .ZN(net89657) );
  NOR2_X4 U1311 ( .A1(\u4/exp_out[2] ), .A2(\u4/N653 ), .ZN(n1787) );
  INV_X2 U1312 ( .A(net86112), .ZN(net85038) );
  NAND2_X2 U1313 ( .A1(n1652), .A2(net85720), .ZN(net86096) );
  NOR2_X4 U1314 ( .A1(net76619), .A2(net85204), .ZN(n2047) );
  NAND2_X2 U1315 ( .A1(net85043), .A2(net85042), .ZN(net76619) );
  XNOR2_X1 U1316 ( .A(net84668), .B(net84610), .ZN(net84667) );
  INV_X4 U1317 ( .A(net85082), .ZN(net88618) );
  INV_X8 U1318 ( .A(net84299), .ZN(net88877) );
  NAND2_X4 U1319 ( .A1(net88895), .A2(n1777), .ZN(n1776) );
  NAND2_X2 U1320 ( .A1(n1794), .A2(net89658), .ZN(net83395) );
  NAND2_X2 U1321 ( .A1(net88646), .A2(n1792), .ZN(net89658) );
  NAND2_X2 U1322 ( .A1(n1951), .A2(n1950), .ZN(n1557) );
  INV_X8 U1323 ( .A(n2383), .ZN(n2385) );
  INV_X8 U1324 ( .A(net85720), .ZN(net88319) );
  INV_X2 U1325 ( .A(\u4/N424 ), .ZN(net84830) );
  NAND2_X4 U1326 ( .A1(\u4/N424 ), .A2(net84522), .ZN(n1869) );
  OAI21_X2 U1327 ( .B1(net84761), .B2(net85712), .A(net84610), .ZN(n1781) );
  NAND3_X1 U1328 ( .A1(net85712), .A2(n2099), .A3(net86038), .ZN(n2090) );
  NOR2_X1 U1329 ( .A1(rmode_r3[0]), .A2(net85847), .ZN(n2279) );
  AOI21_X2 U1330 ( .B1(n2221), .B2(n2261), .A(n2220), .ZN(n2224) );
  AOI21_X2 U1331 ( .B1(net83941), .B2(n1813), .A(n1814), .ZN(n1812) );
  NOR2_X2 U1332 ( .A1(net84206), .A2(net83864), .ZN(n1833) );
  NOR2_X1 U1333 ( .A1(n1720), .A2(n2948), .ZN(n2851) );
  OAI21_X1 U1334 ( .B1(net83849), .B2(n1596), .A(net83439), .ZN(n1906) );
  NAND3_X2 U1335 ( .A1(net84524), .A2(net84518), .A3(net84519), .ZN(net84458)
         );
  NAND3_X2 U1336 ( .A1(n2300), .A2(n2299), .A3(n2298), .ZN(net84524) );
  NOR2_X1 U1337 ( .A1(net85794), .A2(net83439), .ZN(n2299) );
  NOR2_X2 U1338 ( .A1(n2084), .A2(n2083), .ZN(n2085) );
  NAND2_X1 U1339 ( .A1(net89372), .A2(net85832), .ZN(net84160) );
  NOR2_X1 U1340 ( .A1(n2415), .A2(net83878), .ZN(n2325) );
  NOR2_X1 U1341 ( .A1(net11560), .A2(net84167), .ZN(n2562) );
  NAND3_X2 U1342 ( .A1(net84518), .A2(net85790), .A3(net84519), .ZN(net83946)
         );
  AOI21_X2 U1343 ( .B1(n2127), .B2(net85790), .A(n2126), .ZN(n2129) );
  NOR2_X1 U1344 ( .A1(n2306), .A2(n2991), .ZN(n2126) );
  NAND2_X2 U1345 ( .A1(n1842), .A2(net84385), .ZN(n1845) );
  INV_X4 U1346 ( .A(net86015), .ZN(net84394) );
  NAND3_X2 U1347 ( .A1(n2857), .A2(n2856), .A3(n2855), .ZN(n2864) );
  NOR2_X2 U1348 ( .A1(n2904), .A2(n2937), .ZN(n2908) );
  INV_X4 U1349 ( .A(n2190), .ZN(n2054) );
  NOR2_X1 U1350 ( .A1(net11671), .A2(net83993), .ZN(n2207) );
  NAND2_X2 U1351 ( .A1(n2498), .A2(net84128), .ZN(n2499) );
  NOR3_X1 U1352 ( .A1(n2472), .A2(n2471), .A3(n2470), .ZN(n2473) );
  NAND3_X1 U1353 ( .A1(net84343), .A2(net85790), .A3(n2317), .ZN(n2318) );
  AOI21_X1 U1354 ( .B1(n2316), .B2(net85790), .A(n2315), .ZN(n2319) );
  NAND2_X2 U1355 ( .A1(n2372), .A2(n2374), .ZN(n1932) );
  NOR2_X2 U1356 ( .A1(net83791), .A2(n1576), .ZN(net83747) );
  INV_X4 U1357 ( .A(net11567), .ZN(net85827) );
  NAND3_X2 U1358 ( .A1(n1984), .A2(n1573), .A3(n1983), .ZN(n3313) );
  INV_X4 U1359 ( .A(n1911), .ZN(n1910) );
  NOR2_X1 U1360 ( .A1(\u4/exp_in_pl1[3] ), .A2(n2551), .ZN(n2195) );
  NOR2_X2 U1361 ( .A1(n2943), .A2(n2890), .ZN(n2891) );
  NOR2_X1 U1362 ( .A1(net83995), .A2(net83974), .ZN(net83971) );
  AOI21_X1 U1363 ( .B1(n2562), .B2(net85832), .A(net83968), .ZN(n2563) );
  NAND3_X1 U1364 ( .A1(n2141), .A2(n872), .A3(n2140), .ZN(n2142) );
  NOR2_X2 U1365 ( .A1(n2263), .A2(n2243), .ZN(n2150) );
  NOR2_X2 U1366 ( .A1(n2573), .A2(n2546), .ZN(n2547) );
  NAND3_X2 U1367 ( .A1(n2181), .A2(n2180), .A3(n2179), .ZN(n2548) );
  NOR2_X2 U1368 ( .A1(n2172), .A2(n2171), .ZN(n2181) );
  NOR2_X2 U1369 ( .A1(n2174), .A2(n2173), .ZN(n2180) );
  NOR2_X2 U1370 ( .A1(n2469), .A2(n2486), .ZN(n2470) );
  AOI21_X1 U1371 ( .B1(n2305), .B2(net83927), .A(net83969), .ZN(n2312) );
  NAND3_X1 U1372 ( .A1(net83813), .A2(net84501), .A3(net84498), .ZN(net84500)
         );
  NOR2_X2 U1373 ( .A1(net86169), .A2(net84220), .ZN(n2321) );
  AOI211_X2 U1374 ( .C1(\u4/exp_next_mi[3] ), .C2(net84157), .A(net84220), .B(
        net83878), .ZN(n1877) );
  OAI21_X2 U1375 ( .B1(n2121), .B2(n2132), .A(n2120), .ZN(n2281) );
  NOR2_X1 U1376 ( .A1(prod[20]), .A2(n2650), .ZN(n2652) );
  NAND3_X1 U1377 ( .A1(net83940), .A2(net83941), .A3(net83936), .ZN(n2601) );
  NOR2_X1 U1378 ( .A1(n2573), .A2(net83950), .ZN(n2574) );
  NOR2_X2 U1379 ( .A1(n1613), .A2(n1575), .ZN(n2353) );
  OAI21_X1 U1380 ( .B1(n2876), .B2(n2863), .A(n2862), .ZN(n2865) );
  NOR2_X2 U1381 ( .A1(n2928), .A2(n2929), .ZN(n2917) );
  NOR2_X2 U1382 ( .A1(n1927), .A2(n3319), .ZN(net84912) );
  OAI21_X2 U1383 ( .B1(n2105), .B2(n2104), .A(n2103), .ZN(n2106) );
  NAND2_X1 U1384 ( .A1(net84672), .A2(net84673), .ZN(net84602) );
  OAI21_X1 U1385 ( .B1(net83427), .B2(net84600), .A(net83408), .ZN(net84598)
         );
  NOR2_X1 U1386 ( .A1(net83438), .A2(net83427), .ZN(net84599) );
  NOR2_X2 U1387 ( .A1(n1822), .A2(n1823), .ZN(n1824) );
  NOR2_X2 U1388 ( .A1(n1859), .A2(n1617), .ZN(n1858) );
  NOR3_X2 U1389 ( .A1(net84043), .A2(n1561), .A3(net84033), .ZN(n1861) );
  NAND3_X2 U1390 ( .A1(opa_inf), .A2(opb_inf), .A3(sign_exe_r), .ZN(net84047)
         );
  AOI21_X2 U1391 ( .B1(net85778), .B2(net84326), .A(n2303), .ZN(n2158) );
  NAND4_X2 U1392 ( .A1(n2523), .A2(n2527), .A3(n2526), .A4(n2524), .ZN(n2502)
         );
  NOR2_X2 U1393 ( .A1(opa_inf), .A2(opb_00), .ZN(n2376) );
  NOR2_X1 U1394 ( .A1(net84076), .A2(n2531), .ZN(net84073) );
  NOR2_X2 U1395 ( .A1(n3143), .A2(n2767), .ZN(n2730) );
  NOR2_X1 U1396 ( .A1(net83849), .A2(net83933), .ZN(n2114) );
  OAI21_X1 U1397 ( .B1(div_opa_ldz_r2[3]), .B2(net83968), .A(n2292), .ZN(n2285) );
  OAI21_X1 U1398 ( .B1(net83968), .B2(n2225), .A(exp_r[4]), .ZN(n2227) );
  AOI211_X2 U1399 ( .C1(n2258), .C2(n2257), .A(n2256), .B(net83423), .ZN(n2267) );
  AOI21_X1 U1400 ( .B1(n2255), .B2(net84639), .A(net83408), .ZN(n2256) );
  OAI21_X1 U1401 ( .B1(net11555), .B2(net83849), .A(net85828), .ZN(n2597) );
  OAI21_X2 U1402 ( .B1(n2700), .B2(net86010), .A(n2699), .ZN(n2701) );
  NOR2_X2 U1403 ( .A1(n1574), .A2(n1629), .ZN(n2700) );
  INV_X16 U1404 ( .A(net85846), .ZN(net85847) );
  NAND3_X2 U1405 ( .A1(n2538), .A2(n2537), .A3(n2536), .ZN(n2540) );
  NAND3_X2 U1406 ( .A1(n1575), .A2(net84021), .A3(n2535), .ZN(n2537) );
  NOR2_X2 U1407 ( .A1(n3143), .A2(n2833), .ZN(n2759) );
  NOR2_X2 U1408 ( .A1(net84249), .A2(net83791), .ZN(n2430) );
  NOR2_X2 U1409 ( .A1(n2889), .A2(n2896), .ZN(n1993) );
  INV_X8 U1410 ( .A(net85832), .ZN(net85778) );
  NOR3_X2 U1411 ( .A1(net84643), .A2(net84445), .A3(n1852), .ZN(net84645) );
  NAND2_X2 U1412 ( .A1(net84654), .A2(n1788), .ZN(net90079) );
  NOR2_X1 U1413 ( .A1(net83993), .A2(net83994), .ZN(n2560) );
  AOI21_X2 U1414 ( .B1(n2297), .B2(n2296), .A(n2295), .ZN(n2298) );
  INV_X4 U1415 ( .A(net86006), .ZN(net85732) );
  INV_X4 U1416 ( .A(net85071), .ZN(net85211) );
  NOR2_X2 U1417 ( .A1(n1642), .A2(opb_dn), .ZN(n1760) );
  NOR2_X2 U1418 ( .A1(net85847), .A2(n2077), .ZN(n2079) );
  OAI21_X2 U1419 ( .B1(n2260), .B2(n2195), .A(n2194), .ZN(n2202) );
  OAI21_X2 U1420 ( .B1(n2241), .B2(n2240), .A(n2239), .ZN(n2245) );
  NOR2_X2 U1421 ( .A1(n2238), .A2(n2263), .ZN(n2240) );
  NOR3_X1 U1422 ( .A1(n2019), .A2(net84290), .A3(net84305), .ZN(
        \u4/exp_in_pl1[5] ) );
  NAND3_X2 U1423 ( .A1(n1620), .A2(n1587), .A3(n1568), .ZN(n2174) );
  NAND3_X2 U1424 ( .A1(n1619), .A2(n1586), .A3(n1567), .ZN(n2171) );
  NAND3_X2 U1425 ( .A1(n1618), .A2(n1585), .A3(n1566), .ZN(n2172) );
  NAND3_X1 U1426 ( .A1(net83942), .A2(n1817), .A3(net84858), .ZN(n1813) );
  NOR2_X2 U1427 ( .A1(n2836), .A2(n2835), .ZN(n2838) );
  NOR2_X1 U1428 ( .A1(net11670), .A2(net85832), .ZN(n2208) );
  NOR2_X2 U1429 ( .A1(net85137), .A2(net77161), .ZN(net85136) );
  INV_X8 U1430 ( .A(net85196), .ZN(n1865) );
  INV_X4 U1431 ( .A(net85360), .ZN(net85159) );
  NOR2_X2 U1432 ( .A1(net83969), .A2(n2561), .ZN(n2569) );
  AOI21_X2 U1433 ( .B1(net84133), .B2(net84134), .A(net84128), .ZN(n2495) );
  NOR2_X1 U1434 ( .A1(net11560), .A2(n2461), .ZN(n2463) );
  NOR2_X1 U1435 ( .A1(n2466), .A2(n2482), .ZN(n2471) );
  OAI21_X2 U1436 ( .B1(net84884), .B2(n1571), .A(n2145), .ZN(net84853) );
  OAI21_X1 U1437 ( .B1(n2580), .B2(net84675), .A(net85794), .ZN(n2145) );
  NOR2_X1 U1438 ( .A1(net84886), .A2(n1596), .ZN(net84884) );
  AOI21_X1 U1439 ( .B1(n2314), .B2(n2313), .A(net84468), .ZN(n2315) );
  OAI21_X1 U1440 ( .B1(net83933), .B2(net83963), .A(net84465), .ZN(n2313) );
  NAND2_X2 U1441 ( .A1(n2339), .A2(net84421), .ZN(n2498) );
  NOR2_X2 U1442 ( .A1(n2409), .A2(n2408), .ZN(n2410) );
  AOI21_X2 U1443 ( .B1(n2403), .B2(n2444), .A(n2402), .ZN(n2412) );
  NOR2_X1 U1444 ( .A1(\u4/exp_in_pl1[3] ), .A2(n2401), .ZN(n2402) );
  NOR2_X1 U1445 ( .A1(net11555), .A2(n1571), .ZN(net84278) );
  NAND3_X1 U1446 ( .A1(n2304), .A2(net85832), .A3(net83963), .ZN(net83927) );
  NOR2_X1 U1447 ( .A1(opa_dn), .A2(net88427), .ZN(net84506) );
  NAND3_X2 U1448 ( .A1(n2859), .A2(n2862), .A3(n2858), .ZN(n2866) );
  NOR2_X2 U1449 ( .A1(opb_r[11]), .A2(n1725), .ZN(n2771) );
  NOR2_X2 U1450 ( .A1(n2204), .A2(n2203), .ZN(n2212) );
  NOR2_X1 U1451 ( .A1(n3096), .A2(net83994), .ZN(n2203) );
  NOR2_X1 U1452 ( .A1(n1663), .A2(net83968), .ZN(n2204) );
  NOR2_X1 U1453 ( .A1(net11558), .A2(n2209), .ZN(n2210) );
  NAND3_X2 U1454 ( .A1(n2184), .A2(n2183), .A3(n2182), .ZN(n2301) );
  NAND3_X2 U1455 ( .A1(net83934), .A2(n1853), .A3(net83936), .ZN(net83836) );
  NOR2_X2 U1456 ( .A1(n2425), .A2(n2387), .ZN(n2389) );
  NOR3_X2 U1457 ( .A1(n2458), .A2(n2343), .A3(n2342), .ZN(n2344) );
  AOI21_X2 U1458 ( .B1(n1583), .B2(n2418), .A(net85794), .ZN(net84265) );
  OAI21_X2 U1459 ( .B1(net84465), .B2(n2324), .A(n2323), .ZN(net84080) );
  NOR2_X1 U1460 ( .A1(net84468), .A2(net84343), .ZN(n2323) );
  NOR3_X2 U1461 ( .A1(net84469), .A2(net83927), .A3(n2322), .ZN(n2324) );
  AOI21_X2 U1462 ( .B1(n2362), .B2(net84368), .A(n1768), .ZN(n2371) );
  OAI21_X2 U1463 ( .B1(n1628), .B2(n2368), .A(n2367), .ZN(n2369) );
  NAND3_X1 U1464 ( .A1(net85828), .A2(net85790), .A3(n1571), .ZN(n1835) );
  OAI21_X2 U1465 ( .B1(n2100), .B2(n2076), .A(n2102), .ZN(n2108) );
  INV_X4 U1466 ( .A(net89411), .ZN(net89412) );
  INV_X4 U1467 ( .A(net89446), .ZN(net89447) );
  NOR2_X1 U1468 ( .A1(net83968), .A2(n1663), .ZN(n2113) );
  OAI21_X2 U1469 ( .B1(n2284), .B2(n2283), .A(n2282), .ZN(n2292) );
  NOR2_X1 U1470 ( .A1(div_opa_ldz_r2[2]), .A2(exp_r[2]), .ZN(n2283) );
  NOR2_X1 U1471 ( .A1(n2266), .A2(net83427), .ZN(net84617) );
  NOR2_X1 U1472 ( .A1(net84445), .A2(net83402), .ZN(n2258) );
  NOR2_X1 U1473 ( .A1(net84632), .A2(net83403), .ZN(n2257) );
  AOI211_X1 U1474 ( .C1(net84823), .C2(net11566), .A(net84571), .B(net85790), 
        .ZN(n2169) );
  NOR2_X1 U1475 ( .A1(net11555), .A2(net84279), .ZN(net84823) );
  NOR2_X1 U1476 ( .A1(n2307), .A2(net88427), .ZN(net84664) );
  NAND2_X2 U1477 ( .A1(\u1/adj_op_out_sft[1] ), .A2(n2791), .ZN(n2923) );
  NOR2_X2 U1478 ( .A1(n1561), .A2(n1581), .ZN(net84064) );
  NOR2_X2 U1479 ( .A1(net83791), .A2(n1631), .ZN(n2653) );
  NOR3_X1 U1480 ( .A1(prod[17]), .A2(prod[18]), .A3(prod[19]), .ZN(n2651) );
  OAI21_X2 U1481 ( .B1(n2591), .B2(n2590), .A(n2619), .ZN(n2592) );
  NOR2_X2 U1482 ( .A1(n2589), .A2(n2588), .ZN(n2590) );
  NOR3_X2 U1483 ( .A1(n1605), .A2(n2603), .A3(n2602), .ZN(n2607) );
  NOR2_X2 U1484 ( .A1(opa_inf), .A2(net83791), .ZN(n2535) );
  NOR2_X2 U1485 ( .A1(net83791), .A2(n2698), .ZN(n2534) );
  NOR2_X2 U1486 ( .A1(net84326), .A2(net84327), .ZN(n2384) );
  NAND3_X1 U1487 ( .A1(net84465), .A2(net84343), .A3(net85790), .ZN(n2320) );
  INV_X4 U1488 ( .A(n2770), .ZN(n2784) );
  INV_X2 U1489 ( .A(\u1/adj_op_out_sft[4] ), .ZN(n1721) );
  NOR2_X1 U1490 ( .A1(net85794), .A2(n1570), .ZN(n2428) );
  INV_X4 U1491 ( .A(net83419), .ZN(n1783) );
  OAI21_X1 U1492 ( .B1(n2973), .B2(n2972), .A(n2971), .ZN(n2974) );
  AOI21_X1 U1493 ( .B1(n2270), .B2(net84604), .A(net83403), .ZN(n2274) );
  NOR2_X1 U1494 ( .A1(n1852), .A2(net84579), .ZN(n1851) );
  NOR2_X2 U1495 ( .A1(net84913), .A2(n1608), .ZN(net84906) );
  NOR2_X2 U1496 ( .A1(result_zero_sign_d), .A2(n1803), .ZN(n1807) );
  AOI21_X2 U1497 ( .B1(n1561), .B2(n1860), .A(n1861), .ZN(n1855) );
  NOR2_X1 U1498 ( .A1(net84048), .A2(n1863), .ZN(net84028) );
  OAI21_X1 U1499 ( .B1(net85794), .B2(n2376), .A(net83779), .ZN(n2377) );
  INV_X4 U1500 ( .A(n2666), .ZN(n2670) );
  OAI21_X2 U1501 ( .B1(net83791), .B2(n2662), .A(n2661), .ZN(n2669) );
  OAI21_X2 U1502 ( .B1(n2660), .B2(n2659), .A(n1561), .ZN(n2661) );
  NOR2_X2 U1503 ( .A1(opb_inf), .A2(n1572), .ZN(n2660) );
  NOR2_X2 U1504 ( .A1(opa_00), .A2(n1570), .ZN(n2659) );
  NAND2_X2 U1505 ( .A1(n3192), .A2(n3174), .ZN(n3159) );
  NAND2_X2 U1506 ( .A1(n3188), .A2(n3165), .ZN(n3180) );
  NAND2_X2 U1507 ( .A1(n3174), .A2(n3165), .ZN(n3181) );
  NAND2_X2 U1508 ( .A1(n1653), .A2(n3182), .ZN(n3175) );
  NOR3_X2 U1509 ( .A1(n1990), .A2(n2895), .A3(n1989), .ZN(n2959) );
  NOR2_X1 U1510 ( .A1(n1725), .A2(n1723), .ZN(n1987) );
  NOR2_X1 U1511 ( .A1(n1541), .A2(n3017), .ZN(n1986) );
  NOR2_X1 U1512 ( .A1(net83402), .A2(net83403), .ZN(net83394) );
  INV_X8 U1513 ( .A(\u4/f2i_shft[1] ), .ZN(net85712) );
  OAI21_X2 U1514 ( .B1(n2986), .B2(n2976), .A(n2975), .ZN(n2977) );
  NOR2_X1 U1515 ( .A1(\u4/sub_409/net10540 ), .A2(div_opa_ldz_r2[3]), .ZN(
        n2976) );
  NOR2_X1 U1516 ( .A1(net84445), .A2(net84643), .ZN(n2268) );
  OAI211_X2 U1517 ( .C1(net83754), .C2(net83819), .A(net83820), .B(n1546), 
        .ZN(net83802) );
  NOR2_X1 U1518 ( .A1(net85847), .A2(net83791), .ZN(n2539) );
  NOR2_X2 U1519 ( .A1(n2737), .A2(n2736), .ZN(n2741) );
  NOR2_X2 U1520 ( .A1(n2744), .A2(n2743), .ZN(n2747) );
  NOR2_X2 U1521 ( .A1(n2749), .A2(n2748), .ZN(n2752) );
  NOR2_X2 U1522 ( .A1(n2756), .A2(n2755), .ZN(n2762) );
  NOR2_X2 U1523 ( .A1(n3121), .A2(n2765), .ZN(\u2/underflow_d [2]) );
  NOR2_X2 U1524 ( .A1(n2957), .A2(net86010), .ZN(N283) );
  NOR2_X2 U1525 ( .A1(n3156), .A2(fracta_mul[9]), .ZN(\u0/N4 ) );
  NOR2_X2 U1526 ( .A1(n2959), .A2(n2958), .ZN(\u0/N5 ) );
  INV_X1 U1527 ( .A(n3313), .ZN(n3012) );
  OAI21_X2 U1528 ( .B1(n1999), .B2(fracta_mul[8]), .A(n3120), .ZN(N65) );
  AOI21_X2 U1529 ( .B1(n3117), .B2(n1998), .A(fracta_mul[7]), .ZN(n1999) );
  OAI21_X2 U1530 ( .B1(n1997), .B2(n2896), .A(n3116), .ZN(n1998) );
  AOI21_X1 U1531 ( .B1(n3113), .B2(fracta_mul[1]), .A(n2889), .ZN(n1997) );
  OAI21_X2 U1532 ( .B1(n1995), .B2(n1994), .A(n3120), .ZN(n1996) );
  AOI21_X2 U1533 ( .B1(n1993), .B2(n1992), .A(n1991), .ZN(n1995) );
  NOR2_X2 U1534 ( .A1(n2961), .A2(n2960), .ZN(n888) );
  NOR2_X1 U1535 ( .A1(net83438), .A2(n2989), .ZN(n2961) );
  NOR2_X1 U1536 ( .A1(n2962), .A2(net83432), .ZN(n2963) );
  OAI21_X1 U1537 ( .B1(n872), .B2(n2996), .A(n2995), .ZN(\u4/shift_right [3])
         );
  AOI21_X1 U1538 ( .B1(n2994), .B2(net85790), .A(n2993), .ZN(n2995) );
  NOR2_X1 U1539 ( .A1(n2992), .A2(n2991), .ZN(n2993) );
  OAI21_X1 U1540 ( .B1(n872), .B2(net84393), .A(net83368), .ZN(
        \u4/shift_right [4]) );
  AOI21_X1 U1541 ( .B1(n2984), .B2(net85790), .A(n2983), .ZN(net83368) );
  NOR2_X1 U1542 ( .A1(n2982), .A2(n2991), .ZN(n2983) );
  INV_X4 U1543 ( .A(net84030), .ZN(net84027) );
  NAND2_X1 U1544 ( .A1(n2695), .A2(n2676), .ZN(n2677) );
  NAND2_X1 U1545 ( .A1(n2695), .A2(n2682), .ZN(n2684) );
  NAND2_X2 U1546 ( .A1(n1944), .A2(n2695), .ZN(n2668) );
  AND2_X2 U1547 ( .A1(n1749), .A2(net84128), .ZN(n1603) );
  INV_X8 U1548 ( .A(n1748), .ZN(n1749) );
  INV_X4 U1549 ( .A(n2520), .ZN(n2522) );
  NOR3_X2 U1550 ( .A1(n1809), .A2(n1810), .A3(n1811), .ZN(net84051) );
  OAI21_X4 U1551 ( .B1(n2529), .B2(net84083), .A(n1685), .ZN(net84050) );
  NAND2_X1 U1552 ( .A1(n2433), .A2(n1531), .ZN(N232) );
  NAND2_X4 U1553 ( .A1(n1751), .A2(net84409), .ZN(n1748) );
  INV_X4 U1554 ( .A(net84401), .ZN(n1751) );
  NAND2_X4 U1555 ( .A1(net91375), .A2(n1552), .ZN(net84950) );
  NAND2_X2 U1556 ( .A1(net84468), .A2(net84588), .ZN(net84584) );
  OAI22_X2 U1557 ( .A1(n2513), .A2(n2510), .B1(net89485), .B2(n1961), .ZN(
        n2678) );
  AOI21_X2 U1558 ( .B1(net84071), .B2(net84072), .A(net84206), .ZN(n1834) );
  NOR3_X2 U1559 ( .A1(n2595), .A2(n2594), .A3(n2593), .ZN(n2610) );
  INV_X8 U1560 ( .A(net83853), .ZN(net83906) );
  INV_X1 U1561 ( .A(net89657), .ZN(net89919) );
  OAI21_X1 U1562 ( .B1(n2702), .B2(net85794), .A(n2701), .ZN(n2703) );
  NAND3_X2 U1563 ( .A1(n2657), .A2(net83802), .A3(n2658), .ZN(N281) );
  NAND3_X2 U1564 ( .A1(n2656), .A2(net83806), .A3(n2655), .ZN(n2657) );
  AOI21_X2 U1565 ( .B1(n2647), .B2(n2646), .A(n2645), .ZN(n2658) );
  NAND2_X2 U1566 ( .A1(net83395), .A2(net83394), .ZN(net83393) );
  INV_X4 U1567 ( .A(net89054), .ZN(net89055) );
  INV_X4 U1568 ( .A(net84554), .ZN(net84575) );
  BUF_X8 U1569 ( .A(n1535), .Z(net91542) );
  NAND2_X2 U1570 ( .A1(net84329), .A2(net86171), .ZN(net84136) );
  NAND2_X2 U1571 ( .A1(net84329), .A2(rmode_r3[1]), .ZN(n2383) );
  OAI21_X2 U1572 ( .B1(sign), .B2(net84401), .A(net84403), .ZN(net84329) );
  NOR3_X4 U1573 ( .A1(n2709), .A2(n2626), .A3(n2625), .ZN(n2647) );
  NAND2_X4 U1574 ( .A1(net84026), .A2(net84025), .ZN(N254) );
  NAND2_X2 U1575 ( .A1(net84483), .A2(n1654), .ZN(net84554) );
  NAND4_X4 U1576 ( .A1(net90035), .A2(net84912), .A3(net84911), .A4(net84910), 
        .ZN(net84561) );
  INV_X4 U1577 ( .A(net85114), .ZN(net85113) );
  NAND4_X2 U1578 ( .A1(net89943), .A2(n1910), .A3(net85131), .A4(net85180), 
        .ZN(net85114) );
  AND4_X4 U1579 ( .A1(n1636), .A2(n1635), .A3(n1637), .A4(n3193), .ZN(n1558)
         );
  XNOR2_X2 U1580 ( .A(n1676), .B(n1680), .ZN(n1559) );
  INV_X1 U1581 ( .A(n2924), .ZN(n1977) );
  INV_X16 U1582 ( .A(n2926), .ZN(n1975) );
  AND2_X2 U1583 ( .A1(net83779), .A2(net85790), .ZN(n1561) );
  XNOR2_X2 U1584 ( .A(n1625), .B(\sub_435_3/carry [14]), .ZN(n1562) );
  AND2_X2 U1585 ( .A1(\u1/adj_op_out_sft[2] ), .A2(n2791), .ZN(n1563) );
  XNOR2_X2 U1586 ( .A(n1674), .B(\sub_435_b0/carry [3]), .ZN(n1564) );
  XNOR2_X2 U1587 ( .A(n1675), .B(\sub_435_b0/carry [2]), .ZN(n1565) );
  AND2_X4 U1588 ( .A1(net83747), .A2(n1570), .ZN(n1574) );
  AND2_X2 U1589 ( .A1(opb_inf), .A2(net85790), .ZN(n1575) );
  XNOR2_X2 U1590 ( .A(n1624), .B(\sub_435_3/carry [15]), .ZN(n1577) );
  XNOR2_X2 U1591 ( .A(n1637), .B(\sub_435_3/carry [18]), .ZN(n1578) );
  XOR2_X1 U1592 ( .A(div_opa_ldz_r2[3]), .B(net83968), .Z(n1579) );
  AND2_X4 U1593 ( .A1(net84475), .A2(net84150), .ZN(n1580) );
  OR2_X4 U1594 ( .A1(net83791), .A2(n1611), .ZN(n1581) );
  INV_X4 U1595 ( .A(net84079), .ZN(net84157) );
  OR2_X4 U1596 ( .A1(n1731), .A2(n3316), .ZN(n1582) );
  AND2_X2 U1597 ( .A1(n2417), .A2(n2416), .ZN(n1583) );
  AND2_X2 U1598 ( .A1(net84081), .A2(net91404), .ZN(n1588) );
  AND2_X2 U1599 ( .A1(n2187), .A2(net88500), .ZN(n1589) );
  AND2_X2 U1600 ( .A1(\u1/adj_op_out_sft[2] ), .A2(n2793), .ZN(n1590) );
  INV_X2 U1601 ( .A(net85832), .ZN(net15448) );
  INV_X4 U1602 ( .A(net85831), .ZN(net85832) );
  NAND2_X2 U1603 ( .A1(net89863), .A2(net85126), .ZN(n2276) );
  INV_X2 U1604 ( .A(n1977), .ZN(n1976) );
  INV_X8 U1605 ( .A(net91375), .ZN(net89842) );
  XNOR2_X2 U1606 ( .A(n2133), .B(n2100), .ZN(n1592) );
  INV_X4 U1607 ( .A(opb_r[12]), .ZN(n2799) );
  AND2_X2 U1608 ( .A1(n2226), .A2(net84236), .ZN(n1593) );
  INV_X2 U1609 ( .A(\u4/N404 ), .ZN(n1800) );
  XNOR2_X2 U1610 ( .A(n1672), .B(\sub_435_3/carry [17]), .ZN(n1598) );
  XNOR2_X2 U1611 ( .A(n1673), .B(\sub_435_3/carry [16]), .ZN(n1599) );
  XNOR2_X2 U1612 ( .A(n1626), .B(\sub_435_3/carry [13]), .ZN(n1600) );
  XNOR2_X2 U1613 ( .A(n1627), .B(\sub_435_3/carry [12]), .ZN(n1601) );
  XNOR2_X2 U1614 ( .A(n1678), .B(\sub_435_3/carry [11]), .ZN(n1602) );
  AND2_X4 U1615 ( .A1(n2575), .A2(net88500), .ZN(n1605) );
  AND3_X4 U1616 ( .A1(net83941), .A2(net83942), .A3(net84488), .ZN(n1606) );
  AND2_X4 U1617 ( .A1(net84265), .A2(net84266), .ZN(n1607) );
  NAND2_X1 U1618 ( .A1(n1821), .A2(net84015), .ZN(net84651) );
  INV_X4 U1619 ( .A(net84651), .ZN(net84649) );
  CLKBUF_X2 U1620 ( .A(n1761), .Z(net89537) );
  AND2_X2 U1621 ( .A1(n2545), .A2(net83946), .ZN(n1610) );
  AND2_X2 U1622 ( .A1(net86038), .A2(opb_00), .ZN(n1613) );
  INV_X4 U1623 ( .A(n2276), .ZN(n1930) );
  INV_X4 U1624 ( .A(net85140), .ZN(net88566) );
  INV_X2 U1625 ( .A(n2938), .ZN(n2904) );
  OR2_X2 U1626 ( .A1(net84984), .A2(net83933), .ZN(n1621) );
  XNOR2_X2 U1627 ( .A(n1689), .B(n3021), .ZN(n1622) );
  NAND2_X2 U1628 ( .A1(n1757), .A2(net89615), .ZN(n1623) );
  AND2_X2 U1629 ( .A1(n2482), .A2(n2486), .ZN(n1628) );
  AND2_X4 U1630 ( .A1(net83747), .A2(net90287), .ZN(n1629) );
  XOR2_X2 U1631 ( .A(\u2/exp_tmp4[3] ), .B(n3020), .Z(n1630) );
  AND2_X2 U1632 ( .A1(n2425), .A2(net85790), .ZN(n1632) );
  AND2_X2 U1633 ( .A1(net84482), .A2(net84551), .ZN(n1638) );
  OR2_X2 U1634 ( .A1(n2488), .A2(n2489), .ZN(n1639) );
  AND2_X2 U1635 ( .A1(net84673), .A2(net85794), .ZN(n1640) );
  INV_X4 U1636 ( .A(n3124), .ZN(n3136) );
  NAND3_X2 U1637 ( .A1(fpu_op_r1[0]), .A2(fpu_op_r1[1]), .A3(n3100), .ZN(n3124) );
  AND2_X2 U1638 ( .A1(\u1/adj_op_out_sft[1] ), .A2(n1976), .ZN(n1645) );
  AND2_X2 U1639 ( .A1(n2565), .A2(net11558), .ZN(n1646) );
  AND2_X2 U1640 ( .A1(net85786), .A2(net85712), .ZN(n1647) );
  AND3_X4 U1641 ( .A1(n2338), .A2(n2494), .A3(n2490), .ZN(n1648) );
  AND2_X2 U1642 ( .A1(n2928), .A2(n2929), .ZN(n1649) );
  AND2_X4 U1643 ( .A1(n1550), .A2(n1612), .ZN(n1651) );
  NAND2_X2 U1644 ( .A1(\sub_435_b0/carry [10]), .A2(n1558), .ZN(n1653) );
  NAND2_X1 U1645 ( .A1(net89073), .A2(net84568), .ZN(n1654) );
  AND3_X4 U1646 ( .A1(n3132), .A2(n3131), .A3(n2767), .ZN(n1655) );
  INV_X4 U1647 ( .A(net84984), .ZN(net85006) );
  AND4_X4 U1648 ( .A1(n1769), .A2(n1770), .A3(n1771), .A4(net84118), .ZN(n1661) );
  AND3_X4 U1649 ( .A1(n2565), .A2(net83963), .A3(n2564), .ZN(n1662) );
  OR2_X4 U1650 ( .A1(n2991), .A2(net85832), .ZN(n1664) );
  AND2_X2 U1651 ( .A1(\u4/exp_f2i_1 [26]), .A2(n1606), .ZN(n1665) );
  NAND2_X2 U1652 ( .A1(\sub_435_3/carry [20]), .A2(n1635), .ZN(n1666) );
  NAND3_X2 U1653 ( .A1(n2872), .A2(n2854), .A3(n2853), .ZN(n2869) );
  AND2_X2 U1654 ( .A1(net83393), .A2(net83392), .ZN(n1669) );
  OR2_X4 U1655 ( .A1(underflow_fmul_r[1]), .A2(n1612), .ZN(n1670) );
  NAND3_X2 U1656 ( .A1(n2169), .A2(n2168), .A3(n2322), .ZN(net84774) );
  NAND2_X2 U1657 ( .A1(n3085), .A2(n3086), .ZN(net83791) );
  XNOR2_X1 U1658 ( .A(net83968), .B(\u4/add_407/carry [3]), .ZN(n1687) );
  XNOR2_X1 U1659 ( .A(exp_r[4]), .B(\u4/add_407/carry [4]), .ZN(n1688) );
  NAND3_X1 U1660 ( .A1(n3134), .A2(n3136), .A3(n2833), .ZN(n2757) );
  MUX2_X2 U1661 ( .A(\u2/N29 ), .B(\u2/N23 ), .S(n3136), .Z(n3134) );
  NAND3_X2 U1662 ( .A1(n2733), .A2(n2734), .A3(n2735), .ZN(\u2/N44 ) );
  NOR2_X2 U1663 ( .A1(n3142), .A2(n2754), .ZN(n2755) );
  NOR2_X2 U1664 ( .A1(n3141), .A2(n2754), .ZN(n2748) );
  NOR2_X2 U1665 ( .A1(n3140), .A2(n2754), .ZN(n2743) );
  NOR2_X2 U1666 ( .A1(n3139), .A2(n2754), .ZN(n2736) );
  NOR2_X2 U1667 ( .A1(n3138), .A2(n2754), .ZN(n2731) );
  INV_X2 U1668 ( .A(n3143), .ZN(\u2/exp_ovf_d[1] ) );
  INV_X2 U1669 ( .A(\u2/lt_130/A[3] ), .ZN(\u2/exp_tmp4[3] ) );
  OR2_X2 U1670 ( .A1(\u2/lt_130/A[3] ), .A2(\u2/add_111/carry[3] ), .ZN(
        \u2/add_111/carry[4] ) );
  AND2_X2 U1671 ( .A1(\u2/sub_111/carry[3] ), .A2(\u2/lt_130/A[3] ), .ZN(
        \u2/sub_111/carry[4] ) );
  MUX2_X2 U1672 ( .A(\u2/N15 ), .B(\u2/N9 ), .S(n3136), .Z(\u2/lt_130/A[3] )
         );
  MUX2_X2 U1673 ( .A(\u2/N10 ), .B(\u2/N16 ), .S(n3124), .Z(n1689) );
  OR2_X2 U1674 ( .A1(n1689), .A2(\u2/sub_111/carry[4] ), .ZN(
        \u2/sub_111/carry[5] ) );
  AND2_X2 U1675 ( .A1(\u2/add_111/carry[4] ), .A2(\u2/exp_tmp4[4] ), .ZN(
        \u2/add_111/carry[5] ) );
  NOR2_X1 U1676 ( .A1(n2753), .A2(n1622), .ZN(n2732) );
  NOR2_X2 U1677 ( .A1(n2753), .A2(n1630), .ZN(n2737) );
  NOR2_X2 U1678 ( .A1(n2753), .A2(n2742), .ZN(n2744) );
  NOR2_X2 U1679 ( .A1(n2753), .A2(n3018), .ZN(n2749) );
  NOR2_X2 U1680 ( .A1(n2753), .A2(\u2/exp_tmp4[0] ), .ZN(n2756) );
  NAND2_X4 U1681 ( .A1(n2730), .A2(n3124), .ZN(n2753) );
  NOR2_X2 U1682 ( .A1(n2732), .A2(n2731), .ZN(n2735) );
  MUX2_X2 U1683 ( .A(\u2/N10 ), .B(\u2/N16 ), .S(n3124), .Z(\u2/exp_tmp4[4] )
         );
  NOR4_X2 U1684 ( .A1(n3138), .A2(n3136), .A3(opa_r[14]), .A4(n1733), .ZN(
        n3144) );
  NOR2_X4 U1685 ( .A1(n3134), .A2(n3144), .ZN(n3143) );
  NOR3_X1 U1686 ( .A1(n2785), .A2(n2783), .A3(n2784), .ZN(n2786) );
  INV_X8 U1687 ( .A(n2954), .ZN(n1980) );
  INV_X8 U1688 ( .A(n2875), .ZN(n1718) );
  INV_X4 U1689 ( .A(n2875), .ZN(\u1/exp_diff_sft[0] ) );
  AOI21_X2 U1690 ( .B1(n2868), .B2(n2867), .A(n2874), .ZN(n2880) );
  INV_X2 U1691 ( .A(n1718), .ZN(n1719) );
  NOR2_X1 U1692 ( .A1(n1594), .A2(n1560), .ZN(n1988) );
  NOR2_X2 U1693 ( .A1(n2763), .A2(n1594), .ZN(\u2/exp_ovf_d[0] ) );
  NAND2_X2 U1694 ( .A1(opb_r[12]), .A2(n1573), .ZN(n2770) );
  NAND2_X4 U1695 ( .A1(n2822), .A2(n2821), .ZN(n2823) );
  MUX2_X2 U1696 ( .A(n1721), .B(n3102), .S(n1976), .Z(n1720) );
  INV_X4 U1697 ( .A(n1720), .ZN(n2947) );
  OAI21_X4 U1698 ( .B1(n2836), .B2(n2829), .A(n1722), .ZN(n3301) );
  CLKBUF_X2 U1699 ( .A(n2837), .Z(n1722) );
  INV_X4 U1700 ( .A(n3300), .ZN(n2876) );
  NAND2_X1 U1701 ( .A1(n2866), .A2(n3300), .ZN(n2867) );
  AOI21_X1 U1702 ( .B1(n2870), .B2(n2857), .A(n3302), .ZN(n2878) );
  NAND2_X4 U1703 ( .A1(n2837), .A2(n2838), .ZN(n2875) );
  NAND2_X1 U1704 ( .A1(opa_r[14]), .A2(n1734), .ZN(n2789) );
  NAND2_X4 U1705 ( .A1(n1594), .A2(opb_r[14]), .ZN(n2780) );
  NOR2_X2 U1706 ( .A1(opb_r[10]), .A2(n1723), .ZN(n2772) );
  NAND3_X1 U1707 ( .A1(opa_r[12]), .A2(n1988), .A3(n1987), .ZN(n3158) );
  OAI211_X4 U1708 ( .C1(n2883), .C2(n2950), .A(n2925), .B(n2923), .ZN(n2886)
         );
  NOR2_X2 U1709 ( .A1(n2887), .A2(n2945), .ZN(n2892) );
  OAI211_X4 U1710 ( .C1(n2886), .C2(n1563), .A(n2885), .B(n2884), .ZN(n2893)
         );
  OAI211_X4 U1711 ( .C1(n2903), .C2(n2902), .A(n2901), .B(n2900), .ZN(n2909)
         );
  INV_X8 U1712 ( .A(n2791), .ZN(n2793) );
  MUX2_X1 U1713 ( .A(n2878), .B(n2877), .S(n2876), .Z(n2879) );
  NOR2_X2 U1714 ( .A1(opa_r[10]), .A2(opa_r[11]), .ZN(n1983) );
  NAND2_X4 U1715 ( .A1(n2790), .A2(n2789), .ZN(n2926) );
  INV_X1 U1716 ( .A(fracta_mul[1]), .ZN(n3049) );
  INV_X16 U1717 ( .A(n1980), .ZN(n1979) );
  NOR2_X1 U1718 ( .A1(n3016), .A2(n1726), .ZN(n1985) );
  OR2_X4 U1719 ( .A1(n1726), .A2(opa_r[10]), .ZN(\u2/sub_110/carry [1]) );
  AND2_X2 U1720 ( .A1(n1727), .A2(n1728), .ZN(n1981) );
  NOR2_X1 U1721 ( .A1(n2779), .A2(n2791), .ZN(n2787) );
  NOR2_X1 U1722 ( .A1(n2927), .A2(n2791), .ZN(n2953) );
  NAND2_X4 U1723 ( .A1(n2882), .A2(n2791), .ZN(n2925) );
  AOI21_X1 U1724 ( .B1(n1718), .B2(n2865), .A(n2864), .ZN(n2868) );
  NAND2_X1 U1725 ( .A1(n1718), .A2(n3308), .ZN(n2870) );
  INV_X4 U1726 ( .A(n1729), .ZN(n1982) );
  NAND3_X1 U1727 ( .A1(n1982), .A2(n1726), .A3(n1981), .ZN(n1731) );
  NAND3_X2 U1728 ( .A1(n1982), .A2(n1726), .A3(n1981), .ZN(\u6/N10 ) );
  NAND2_X1 U1729 ( .A1(opb_r[10]), .A2(n1723), .ZN(n2781) );
  AND2_X2 U1730 ( .A1(opa_r[10]), .A2(opb_r[10]), .ZN(\u2/add_110/carry [1])
         );
  INV_X1 U1731 ( .A(opb_r[14]), .ZN(n1732) );
  INV_X4 U1732 ( .A(n1732), .ZN(n1733) );
  INV_X1 U1733 ( .A(n1731), .ZN(n3013) );
  NOR2_X1 U1734 ( .A1(n3313), .A2(n1731), .ZN(n2836) );
  NOR2_X1 U1735 ( .A1(opa_r[14]), .A2(n1731), .ZN(n2768) );
  OAI22_X1 U1736 ( .A1(n3130), .A2(n1731), .B1(n3129), .B2(n3313), .ZN(n2765)
         );
  NAND2_X1 U1737 ( .A1(n3313), .A2(n1731), .ZN(n2833) );
  NOR2_X1 U1738 ( .A1(opb_r[13]), .A2(n1560), .ZN(n2778) );
  NAND2_X1 U1739 ( .A1(opb_r[13]), .A2(n1560), .ZN(n2769) );
  NAND3_X1 U1740 ( .A1(opb_r[12]), .A2(n1986), .A3(n1985), .ZN(n3157) );
  NOR2_X1 U1741 ( .A1(opa_r[14]), .A2(n1733), .ZN(n2766) );
  INV_X1 U1742 ( .A(opb_r[13]), .ZN(n3017) );
  AOI21_X2 U1743 ( .B1(net83863), .B2(net83862), .A(net83864), .ZN(n2627) );
  INV_X8 U1744 ( .A(n2708), .ZN(n2665) );
  INV_X4 U1745 ( .A(n2707), .ZN(n2626) );
  AND2_X2 U1746 ( .A1(n2623), .A2(n2433), .ZN(n1736) );
  AOI211_X4 U1747 ( .C1(n2337), .C2(n1925), .A(n2335), .B(n2334), .ZN(n2348)
         );
  NAND3_X2 U1748 ( .A1(net84315), .A2(net84263), .A3(net84366), .ZN(n2419) );
  OAI211_X1 U1749 ( .C1(n2422), .C2(n2421), .A(n1597), .B(net84263), .ZN(n2423) );
  NAND2_X4 U1750 ( .A1(n2358), .A2(n2357), .ZN(net84263) );
  OAI21_X2 U1751 ( .B1(n2596), .B2(n2326), .A(n2325), .ZN(n2329) );
  INV_X2 U1752 ( .A(n2596), .ZN(n2613) );
  OR3_X4 U1753 ( .A1(n2540), .A2(net84012), .A3(n2539), .ZN(n1742) );
  NAND2_X4 U1754 ( .A1(n2524), .A2(n2523), .ZN(net84059) );
  NAND3_X4 U1755 ( .A1(fract_out_q[5]), .A2(net85730), .A3(net85718), .ZN(
        n2023) );
  OAI21_X4 U1756 ( .B1(net88618), .B2(net89546), .A(net84758), .ZN(n1900) );
  NAND3_X4 U1757 ( .A1(net85227), .A2(n1744), .A3(net85678), .ZN(net85061) );
  INV_X32 U1758 ( .A(net85754), .ZN(net85752) );
  INV_X4 U1759 ( .A(net84677), .ZN(net86171) );
  INV_X8 U1760 ( .A(\u4/fract_out_pl1[10] ), .ZN(net84677) );
  NAND2_X2 U1761 ( .A1(net83863), .A2(net83862), .ZN(net83870) );
  INV_X8 U1762 ( .A(net85290), .ZN(net85240) );
  OAI21_X4 U1763 ( .B1(n2672), .B2(n2673), .A(n2671), .ZN(N285) );
  INV_X2 U1764 ( .A(n1915), .ZN(n2365) );
  NAND3_X2 U1765 ( .A1(n1915), .A2(n2425), .A3(net85794), .ZN(net84079) );
  NAND3_X2 U1766 ( .A1(n1915), .A2(n2566), .A3(n1632), .ZN(n2486) );
  NAND3_X2 U1767 ( .A1(n2555), .A2(n1915), .A3(n1632), .ZN(n2482) );
  INV_X8 U1768 ( .A(n2997), .ZN(n2996) );
  NAND2_X4 U1769 ( .A1(n2456), .A2(n2997), .ZN(net84072) );
  NAND2_X4 U1770 ( .A1(n2358), .A2(n2357), .ZN(n2997) );
  NOR2_X4 U1771 ( .A1(net84055), .A2(n1806), .ZN(n1805) );
  NAND2_X1 U1772 ( .A1(n2433), .A2(n2689), .ZN(n2690) );
  NAND2_X4 U1773 ( .A1(net89595), .A2(net84584), .ZN(net84553) );
  INV_X8 U1774 ( .A(net84553), .ZN(net84574) );
  OAI211_X4 U1775 ( .C1(n1841), .C2(n1843), .A(net84149), .B(net85842), .ZN(
        n1840) );
  INV_X32 U1776 ( .A(n1960), .ZN(n1961) );
  NAND2_X4 U1777 ( .A1(net83934), .A2(net84571), .ZN(net84648) );
  NAND2_X4 U1778 ( .A1(net84552), .A2(n1638), .ZN(n2356) );
  NOR2_X2 U1779 ( .A1(net85736), .A2(net85720), .ZN(net85297) );
  XNOR2_X2 U1780 ( .A(net84136), .B(net30297), .ZN(n2370) );
  INV_X1 U1781 ( .A(net85998), .ZN(net90217) );
  NAND3_X2 U1782 ( .A1(n1942), .A2(quo[1]), .A3(net85684), .ZN(n1743) );
  NAND3_X2 U1783 ( .A1(n1894), .A2(quo[1]), .A3(net85684), .ZN(net85261) );
  OAI21_X4 U1784 ( .B1(net85373), .B2(net85676), .A(net85374), .ZN(n1914) );
  NAND2_X4 U1785 ( .A1(net89129), .A2(quo[7]), .ZN(net85373) );
  INV_X4 U1786 ( .A(net85748), .ZN(n1744) );
  NOR2_X1 U1787 ( .A1(net84060), .A2(net83875), .ZN(n1804) );
  INV_X1 U1788 ( .A(net84471), .ZN(n1747) );
  AOI21_X4 U1789 ( .B1(n2355), .B2(net84214), .A(n2354), .ZN(n2374) );
  NAND3_X1 U1790 ( .A1(net85847), .A2(n2588), .A3(net83861), .ZN(n2354) );
  INV_X4 U1791 ( .A(net86171), .ZN(net91353) );
  NAND3_X4 U1792 ( .A1(net84343), .A2(net86171), .A3(net84334), .ZN(net84371)
         );
  NOR2_X2 U1793 ( .A1(n2350), .A2(n2349), .ZN(n2355) );
  OAI21_X4 U1794 ( .B1(net90047), .B2(n1623), .A(n1756), .ZN(net85021) );
  INV_X8 U1795 ( .A(net86165), .ZN(net90047) );
  NOR2_X1 U1796 ( .A1(n2541), .A2(n2441), .ZN(net83862) );
  NAND2_X1 U1797 ( .A1(n1849), .A2(net88721), .ZN(n1750) );
  OAI22_X4 U1798 ( .A1(net84322), .A2(n1961), .B1(n1928), .B2(n2386), .ZN(
        n2515) );
  OAI22_X4 U1799 ( .A1(net89716), .A2(n1961), .B1(n1928), .B2(n2508), .ZN(
        n2685) );
  INV_X4 U1800 ( .A(net84523), .ZN(n1766) );
  NOR3_X4 U1801 ( .A1(n2678), .A2(n2676), .A3(n2680), .ZN(n2517) );
  NAND2_X4 U1802 ( .A1(net84846), .A2(n1753), .ZN(n1752) );
  OR2_X2 U1803 ( .A1(net84778), .A2(net84845), .ZN(n1753) );
  NAND2_X2 U1804 ( .A1(\u4/N426 ), .A2(net84522), .ZN(n1754) );
  NAND2_X4 U1805 ( .A1(\u4/N426 ), .A2(net84522), .ZN(n1899) );
  NAND2_X1 U1806 ( .A1(div_opa_ldz_r2[1]), .A2(net84901), .ZN(n2103) );
  INV_X16 U1807 ( .A(net84982), .ZN(net83933) );
  NAND2_X4 U1808 ( .A1(net11555), .A2(net85033), .ZN(net84982) );
  INV_X8 U1809 ( .A(net83421), .ZN(\u4/exp_in_pl1[2] ) );
  NAND2_X2 U1810 ( .A1(net88636), .A2(net85089), .ZN(n1755) );
  INV_X8 U1811 ( .A(net86026), .ZN(net88636) );
  INV_X1 U1812 ( .A(net84895), .ZN(n1757) );
  INV_X1 U1813 ( .A(net85790), .ZN(n1758) );
  NAND2_X1 U1814 ( .A1(n1757), .A2(n1758), .ZN(n1756) );
  NAND2_X4 U1815 ( .A1(net85296), .A2(n1759), .ZN(net85161) );
  NAND2_X2 U1816 ( .A1(n2001), .A2(n1760), .ZN(n1759) );
  INV_X16 U1817 ( .A(n1880), .ZN(n1879) );
  BUF_X32 U1818 ( .A(net84909), .Z(net90035) );
  NAND4_X4 U1819 ( .A1(net85061), .A2(n2043), .A3(n2067), .A4(n2066), .ZN(
        n3004) );
  AOI21_X2 U1820 ( .B1(net90302), .B2(net89372), .A(net83407), .ZN(net84502)
         );
  INV_X2 U1821 ( .A(net89965), .ZN(net89372) );
  INV_X2 U1822 ( .A(net84755), .ZN(net89121) );
  OAI22_X4 U1823 ( .A1(n1928), .A2(n2506), .B1(net84118), .B2(n1961), .ZN(
        n2691) );
  OAI22_X4 U1824 ( .A1(net84103), .A2(n1961), .B1(n1928), .B2(n2512), .ZN(
        n2674) );
  OAI22_X4 U1825 ( .A1(n1555), .A2(n1961), .B1(n2513), .B2(n2509), .ZN(n2676)
         );
  NAND2_X2 U1826 ( .A1(net84199), .A2(net84200), .ZN(n2457) );
  AOI21_X4 U1827 ( .B1(n1580), .B2(n1529), .A(net84390), .ZN(n1762) );
  AOI211_X2 U1828 ( .C1(net85842), .C2(net84386), .A(net84387), .B(n1762), 
        .ZN(net84199) );
  INV_X1 U1829 ( .A(net84808), .ZN(n1771) );
  INV_X8 U1830 ( .A(net84014), .ZN(net85846) );
  NAND2_X4 U1831 ( .A1(net85028), .A2(n1744), .ZN(net84014) );
  BUF_X16 U1832 ( .A(net84570), .Z(net89029) );
  INV_X2 U1833 ( .A(net84059), .ZN(n1808) );
  NAND4_X1 U1834 ( .A1(n2164), .A2(n2166), .A3(n2167), .A4(n2165), .ZN(n1763)
         );
  INV_X4 U1835 ( .A(net84565), .ZN(n1764) );
  NAND4_X2 U1836 ( .A1(n2165), .A2(n2166), .A3(n2167), .A4(n2164), .ZN(
        net84523) );
  INV_X4 U1837 ( .A(n1763), .ZN(net84565) );
  INV_X4 U1838 ( .A(net84472), .ZN(net89664) );
  NAND2_X4 U1839 ( .A1(net84674), .A2(net83429), .ZN(net84472) );
  INV_X4 U1840 ( .A(net83787), .ZN(net83819) );
  NAND4_X2 U1841 ( .A1(net84569), .A2(net84648), .A3(net99831), .A4(net84649), 
        .ZN(net84644) );
  NAND2_X4 U1842 ( .A1(net84381), .A2(n1554), .ZN(net30297) );
  OAI21_X4 U1843 ( .B1(net84574), .B2(net84575), .A(net84576), .ZN(net84381)
         );
  NAND3_X2 U1844 ( .A1(net84554), .A2(net84553), .A3(net84403), .ZN(net84552)
         );
  OAI21_X4 U1845 ( .B1(net91375), .B2(net85017), .A(net84967), .ZN(net84870)
         );
  NAND2_X4 U1846 ( .A1(n2520), .A2(n2459), .ZN(n2460) );
  INV_X1 U1847 ( .A(n2521), .ZN(n2459) );
  OAI21_X4 U1848 ( .B1(n2528), .B2(n2502), .A(net83861), .ZN(net84010) );
  NAND2_X4 U1849 ( .A1(n2351), .A2(net84149), .ZN(net84214) );
  OAI21_X4 U1850 ( .B1(n1766), .B2(n1765), .A(net84649), .ZN(net84573) );
  INV_X1 U1851 ( .A(net91325), .ZN(n1765) );
  NOR2_X2 U1852 ( .A1(net89664), .A2(net84676), .ZN(net89663) );
  AOI21_X2 U1853 ( .B1(net84070), .B2(net84069), .A(sign_fasu_r), .ZN(n1810)
         );
  INV_X4 U1854 ( .A(net83868), .ZN(net84069) );
  NAND4_X1 U1855 ( .A1(net84150), .A2(net84081), .A3(n2478), .A4(net84169), 
        .ZN(n2345) );
  INV_X8 U1856 ( .A(net84220), .ZN(net84081) );
  NAND3_X1 U1857 ( .A1(net83950), .A2(n2302), .A3(\u4/fract_out_pl1[10] ), 
        .ZN(net84398) );
  INV_X8 U1858 ( .A(net84458), .ZN(net83950) );
  OAI21_X4 U1859 ( .B1(net89663), .B2(\u4/exp_out[4] ), .A(net84014), .ZN(
        net84588) );
  NAND3_X2 U1860 ( .A1(n1767), .A2(net85337), .A3(net85210), .ZN(n3001) );
  INV_X1 U1861 ( .A(net85336), .ZN(n1767) );
  NAND2_X4 U1862 ( .A1(n1951), .A2(n1950), .ZN(net84753) );
  NAND3_X4 U1863 ( .A1(n1768), .A2(n2365), .A3(rmode_r3[0]), .ZN(net84135) );
  AND2_X2 U1864 ( .A1(n1764), .A2(net84522), .ZN(n1823) );
  AOI211_X4 U1865 ( .C1(sign), .C2(net84403), .A(net84480), .B(net84675), .ZN(
        net84409) );
  INV_X1 U1866 ( .A(net84456), .ZN(n1769) );
  INV_X1 U1867 ( .A(\u4/fract_out[8] ), .ZN(n1770) );
  INV_X4 U1868 ( .A(net84676), .ZN(net84471) );
  NAND2_X4 U1869 ( .A1(n1772), .A2(net89842), .ZN(net89224) );
  INV_X1 U1870 ( .A(net84956), .ZN(n1772) );
  AOI21_X4 U1871 ( .B1(net84588), .B2(net84468), .A(n1824), .ZN(net84483) );
  INV_X8 U1872 ( .A(net84015), .ZN(net84468) );
  AOI211_X4 U1873 ( .C1(\u4/exp_f2i_1 [25]), .C2(n1606), .A(net83406), .B(
        n1773), .ZN(net83392) );
  OAI21_X4 U1874 ( .B1(n1774), .B2(n1775), .A(n1776), .ZN(n1773) );
  NOR2_X1 U1875 ( .A1(net88427), .A2(net83403), .ZN(n1777) );
  INV_X8 U1876 ( .A(opb_dn), .ZN(net88427) );
  NAND2_X2 U1877 ( .A1(net83416), .A2(net83417), .ZN(n1775) );
  INV_X4 U1878 ( .A(net83403), .ZN(net83417) );
  AOI211_X2 U1879 ( .C1(net83417), .C2(net84615), .A(n1665), .B(net84617), 
        .ZN(net84614) );
  AOI211_X4 U1880 ( .C1(net84655), .C2(net83417), .A(net84656), .B(net84657), 
        .ZN(net84654) );
  INV_X4 U1881 ( .A(net84611), .ZN(net83416) );
  NAND2_X2 U1882 ( .A1(net83416), .A2(net84667), .ZN(net84660) );
  NAND2_X2 U1883 ( .A1(net83416), .A2(net84629), .ZN(net84625) );
  NAND2_X4 U1884 ( .A1(n1785), .A2(n1786), .ZN(n1774) );
  NAND2_X4 U1885 ( .A1(n1783), .A2(n1784), .ZN(n1786) );
  INV_X8 U1886 ( .A(n1778), .ZN(n1784) );
  INV_X2 U1887 ( .A(n1784), .ZN(net90268) );
  INV_X8 U1888 ( .A(n1780), .ZN(n1778) );
  NAND2_X2 U1889 ( .A1(n1778), .A2(net83419), .ZN(n1785) );
  OAI21_X4 U1890 ( .B1(net85710), .B2(n1779), .A(n1781), .ZN(n1780) );
  NAND2_X4 U1891 ( .A1(net85313), .A2(n1782), .ZN(\u4/f2i_shft[1] ) );
  INV_X4 U1892 ( .A(net85030), .ZN(n1782) );
  INV_X4 U1893 ( .A(net84761), .ZN(n1779) );
  NOR2_X1 U1894 ( .A1(net89924), .A2(n1779), .ZN(net83987) );
  XNOR2_X2 U1895 ( .A(n1779), .B(net85710), .ZN(net84668) );
  INV_X32 U1896 ( .A(net85712), .ZN(net85710) );
  NAND2_X2 U1897 ( .A1(n1787), .A2(net91144), .ZN(\u4/N655 ) );
  INV_X4 U1898 ( .A(net90079), .ZN(net91144) );
  BUF_X32 U1899 ( .A(net90079), .Z(net91404) );
  NOR2_X4 U1900 ( .A1(n1789), .A2(n1790), .ZN(n1788) );
  NAND2_X4 U1901 ( .A1(n845), .A2(net84637), .ZN(n1790) );
  NOR2_X4 U1902 ( .A1(n1791), .A2(net83945), .ZN(n1789) );
  OR2_X4 U1903 ( .A1(net85788), .A2(net83951), .ZN(n1791) );
  INV_X16 U1904 ( .A(net76872), .ZN(net85788) );
  INV_X4 U1905 ( .A(net84658), .ZN(net84657) );
  NAND2_X4 U1906 ( .A1(\u4/exp_f2i_1 [24]), .A2(n1606), .ZN(net84658) );
  INV_X4 U1907 ( .A(net85847), .ZN(net83941) );
  AOI22_X1 U1908 ( .A1(n1574), .A2(n1744), .B1(n1550), .B2(n1670), .ZN(
        net83827) );
  INV_X1 U1909 ( .A(n1744), .ZN(net90287) );
  INV_X16 U1910 ( .A(net85752), .ZN(net85746) );
  INV_X32 U1911 ( .A(net85752), .ZN(net85744) );
  INV_X16 U1912 ( .A(net85756), .ZN(net85754) );
  INV_X4 U1913 ( .A(net11675), .ZN(net85756) );
  INV_X4 U1914 ( .A(net85323), .ZN(net85028) );
  NAND2_X1 U1915 ( .A1(net85028), .A2(net91548), .ZN(net84341) );
  NAND2_X4 U1916 ( .A1(net85028), .A2(n1643), .ZN(net85320) );
  NAND2_X4 U1917 ( .A1(net85730), .A2(net85722), .ZN(net85323) );
  INV_X16 U1918 ( .A(net85724), .ZN(net85722) );
  INV_X16 U1919 ( .A(net85726), .ZN(net85724) );
  INV_X16 U1920 ( .A(net85724), .ZN(net85720) );
  INV_X4 U1921 ( .A(net11677), .ZN(net85726) );
  INV_X16 U1922 ( .A(net85738), .ZN(net85730) );
  INV_X32 U1923 ( .A(net85740), .ZN(net85738) );
  INV_X16 U1924 ( .A(net85742), .ZN(net85740) );
  INV_X8 U1925 ( .A(net85740), .ZN(net85736) );
  INV_X4 U1926 ( .A(net11676), .ZN(net85742) );
  NAND2_X4 U1927 ( .A1(net84471), .A2(net84472), .ZN(\u4/exp_out[4] ) );
  NAND2_X4 U1928 ( .A1(net89657), .A2(net89736), .ZN(n1794) );
  NAND2_X4 U1929 ( .A1(n1793), .A2(net83398), .ZN(net89736) );
  INV_X4 U1930 ( .A(net89736), .ZN(net88646) );
  INV_X4 U1931 ( .A(net84606), .ZN(net83398) );
  AOI21_X2 U1932 ( .B1(net84663), .B2(net83398), .A(net84664), .ZN(net84662)
         );
  NOR3_X1 U1933 ( .A1(net85790), .A2(net83398), .A3(net83951), .ZN(net84591)
         );
  NAND3_X1 U1934 ( .A1(net89919), .A2(net84766), .A3(net83398), .ZN(net84642)
         );
  AOI21_X4 U1935 ( .B1(\u4/exp_next_mi[1] ), .B2(net85788), .A(n1647), .ZN(
        n1793) );
  INV_X32 U1936 ( .A(net85788), .ZN(net85786) );
  AOI22_X4 U1937 ( .A1(\u4/exp_in_pl1[2] ), .A2(net85786), .B1(
        \u4/exp_next_mi[2] ), .B2(net85788), .ZN(n1792) );
  NAND2_X1 U1938 ( .A1(\u4/exp_in_pl1[2] ), .A2(net110951), .ZN(net84298) );
  NOR2_X1 U1939 ( .A1(\u4/exp_in_pl1[2] ), .A2(net110951), .ZN(net84297) );
  NAND3_X1 U1940 ( .A1(net77815), .A2(net84606), .A3(net84633), .ZN(net84661)
         );
  NOR2_X1 U1941 ( .A1(net83402), .A2(net84606), .ZN(net84605) );
  BUF_X32 U1942 ( .A(\u4/exp_next_mi[1] ), .Z(net89692) );
  NAND2_X2 U1943 ( .A1(\u4/exp_next_mi[1] ), .A2(net85788), .ZN(net91056) );
  INV_X4 U1944 ( .A(net85313), .ZN(net85316) );
  XNOR2_X2 U1945 ( .A(net85313), .B(net11560), .ZN(net83421) );
  NOR2_X1 U1946 ( .A1(net85030), .A2(net11560), .ZN(net84916) );
  BUF_X32 U1947 ( .A(\u4/exp_next_mi[2] ), .Z(net89948) );
  MUX2_X2 U1948 ( .A(\u4/exp_next_mi[0] ), .B(net85778), .S(net76872), .Z(
        net84606) );
  NAND2_X1 U1949 ( .A1(net85712), .A2(net76872), .ZN(net91057) );
  BUF_X32 U1950 ( .A(\u4/exp_out[2] ), .Z(net86169) );
  NAND2_X2 U1951 ( .A1(net83849), .A2(net84236), .ZN(net83402) );
  INV_X8 U1952 ( .A(net83813), .ZN(net83849) );
  NAND2_X2 U1953 ( .A1(net84669), .A2(net86067), .ZN(net83403) );
  INV_X4 U1954 ( .A(net84452), .ZN(net84674) );
  OAI21_X4 U1955 ( .B1(net84678), .B2(net84677), .A(net84451), .ZN(net84676)
         );
  INV_X4 U1956 ( .A(net84679), .ZN(net84451) );
  NAND2_X2 U1957 ( .A1(net84451), .A2(net84452), .ZN(net84450) );
  OAI21_X2 U1958 ( .B1(net85794), .B2(net83995), .A(n1795), .ZN(net84679) );
  AOI21_X2 U1959 ( .B1(\u4/exp_f2i_1 [27]), .B2(n1606), .A(n1796), .ZN(n1795)
         );
  NAND2_X1 U1960 ( .A1(n1797), .A2(net84637), .ZN(n1796) );
  NAND3_X1 U1961 ( .A1(net84639), .A2(net83990), .A3(net84683), .ZN(n1797) );
  INV_X4 U1962 ( .A(net83408), .ZN(net84683) );
  NAND2_X1 U1963 ( .A1(net84683), .A2(net90302), .ZN(net84659) );
  NAND2_X4 U1964 ( .A1(net84586), .A2(net84569), .ZN(net84769) );
  OAI21_X4 U1965 ( .B1(net84769), .B2(net84573), .A(net84770), .ZN(net84678)
         );
  NAND3_X2 U1966 ( .A1(net84570), .A2(net84572), .A3(net84571), .ZN(net84586)
         );
  INV_X4 U1967 ( .A(net84829), .ZN(net84571) );
  NAND2_X2 U1968 ( .A1(net83936), .A2(n1571), .ZN(net84829) );
  NOR4_X4 U1969 ( .A1(net84808), .A2(\u4/fract_out[8] ), .A3(n1752), .A4(
        net84456), .ZN(net84572) );
  INV_X4 U1970 ( .A(net84811), .ZN(net84570) );
  NAND3_X2 U1971 ( .A1(n1798), .A2(n1799), .A3(n1801), .ZN(net84811) );
  INV_X4 U1972 ( .A(net84814), .ZN(n1801) );
  NOR2_X4 U1973 ( .A1(\u4/fract_out[5] ), .A2(n1924), .ZN(n1799) );
  NAND2_X2 U1974 ( .A1(net89819), .A2(net84842), .ZN(\u4/fract_out[7] ) );
  NAND2_X4 U1975 ( .A1(net84836), .A2(n1802), .ZN(\u4/fract_out[4] ) );
  NAND2_X2 U1976 ( .A1(net91150), .A2(\u4/N404 ), .ZN(n1802) );
  OAI21_X4 U1977 ( .B1(net84778), .B2(n1800), .A(net84836), .ZN(net89933) );
  INV_X1 U1978 ( .A(net84778), .ZN(net91150) );
  NAND2_X4 U1979 ( .A1(\u4/N428 ), .A2(net84522), .ZN(net84836) );
  INV_X16 U1980 ( .A(net84566), .ZN(net84522) );
  NAND2_X4 U1981 ( .A1(net84774), .A2(net84775), .ZN(net84569) );
  NAND3_X1 U1982 ( .A1(net89073), .A2(net84568), .A3(net84569), .ZN(net84484)
         );
  NAND2_X4 U1983 ( .A1(net84908), .A2(net91112), .ZN(net83936) );
  INV_X4 U1984 ( .A(net84561), .ZN(net84908) );
  NAND2_X4 U1985 ( .A1(net84110), .A2(net84113), .ZN(net84808) );
  NAND4_X2 U1986 ( .A1(n1750), .A2(net84050), .A3(net84051), .A4(net84052), 
        .ZN(net84025) );
  NAND4_X2 U1987 ( .A1(net84024), .A2(n1804), .A3(n1805), .A4(net83819), .ZN(
        net84052) );
  NOR2_X4 U1988 ( .A1(sign_fasu_r), .A2(net83819), .ZN(n1809) );
  NAND2_X2 U1989 ( .A1(net84024), .A2(net83819), .ZN(net83883) );
  NAND2_X2 U1990 ( .A1(n1807), .A2(n1808), .ZN(n1806) );
  INV_X4 U1991 ( .A(net83747), .ZN(n1803) );
  NOR2_X1 U1992 ( .A1(net84015), .A2(n1803), .ZN(net84012) );
  NAND2_X2 U1993 ( .A1(net84064), .A2(net84044), .ZN(n1811) );
  NAND2_X2 U1994 ( .A1(nan_sign_d), .A2(n1581), .ZN(net84043) );
  NAND2_X2 U1995 ( .A1(net11627), .A2(n1611), .ZN(net83781) );
  INV_X32 U1996 ( .A(net85794), .ZN(net85790) );
  INV_X16 U1997 ( .A(net86067), .ZN(net85794) );
  NAND2_X2 U1998 ( .A1(net84619), .A2(net86067), .ZN(net83427) );
  INV_X4 U1999 ( .A(net83791), .ZN(net83779) );
  NAND2_X4 U2000 ( .A1(\u4/N433 ), .A2(net84522), .ZN(net84846) );
  NAND3_X2 U2001 ( .A1(net84847), .A2(net84848), .A3(n1812), .ZN(net84566) );
  NOR2_X1 U2002 ( .A1(net84565), .A2(net84566), .ZN(net84555) );
  OAI21_X4 U2003 ( .B1(net84830), .B2(net84566), .A(net84810), .ZN(net60630)
         );
  NAND2_X2 U2004 ( .A1(net84564), .A2(net84566), .ZN(net84519) );
  NAND2_X2 U2005 ( .A1(n1815), .A2(net84853), .ZN(n1814) );
  NAND2_X2 U2006 ( .A1(net84854), .A2(n1816), .ZN(n1815) );
  NAND2_X2 U2007 ( .A1(net11555), .A2(net11558), .ZN(n1816) );
  INV_X2 U2008 ( .A(net84856), .ZN(net84854) );
  INV_X4 U2009 ( .A(\u4/f2i_shft[4] ), .ZN(n1817) );
  NAND2_X1 U2010 ( .A1(n1818), .A2(net83439), .ZN(net89615) );
  OAI21_X1 U2011 ( .B1(net85828), .B2(net83849), .A(net83974), .ZN(n1818) );
  INV_X32 U2012 ( .A(net85827), .ZN(net85828) );
  INV_X4 U2013 ( .A(\u4/N656 ), .ZN(net86165) );
  NAND2_X2 U2014 ( .A1(net90997), .A2(net86165), .ZN(net110929) );
  NOR2_X4 U2015 ( .A1(net86165), .A2(n1621), .ZN(net91177) );
  NAND2_X4 U2016 ( .A1(net83813), .A2(n1571), .ZN(net83439) );
  NAND2_X2 U2017 ( .A1(net83849), .A2(n1571), .ZN(net83974) );
  OAI21_X4 U2018 ( .B1(net83973), .B2(net83974), .A(net83975), .ZN(net83972)
         );
  NAND2_X2 U2019 ( .A1(n1641), .A2(net88427), .ZN(net83813) );
  OAI211_X1 U2020 ( .C1(net83811), .C2(net83812), .A(net86038), .B(net83813), 
        .ZN(net83807) );
  NAND2_X1 U2021 ( .A1(opa_dn), .A2(net85676), .ZN(net84669) );
  NAND2_X2 U2022 ( .A1(opa_dn), .A2(net84722), .ZN(net84611) );
  NOR2_X4 U2023 ( .A1(net85718), .A2(net11582), .ZN(n1819) );
  AOI21_X4 U2024 ( .B1(net85297), .B2(fract_out_q[3]), .A(n1819), .ZN(net85296) );
  INV_X32 U2025 ( .A(net85720), .ZN(net85718) );
  AND2_X2 U2026 ( .A1(net99831), .A2(net84649), .ZN(net89073) );
  NAND2_X1 U2027 ( .A1(net91325), .A2(n1763), .ZN(net99831) );
  NAND2_X4 U2028 ( .A1(net84483), .A2(net84484), .ZN(net84401) );
  INV_X4 U2029 ( .A(n1820), .ZN(n1822) );
  AOI21_X1 U2030 ( .B1(net84518), .B2(net84519), .A(net84015), .ZN(n1820) );
  NAND3_X2 U2031 ( .A1(net84571), .A2(net83849), .A3(net85794), .ZN(n1821) );
  NAND3_X4 U2032 ( .A1(net84948), .A2(net89224), .A3(net84950), .ZN(
        \u4/shift_left [0]) );
  NOR2_X4 U2033 ( .A1(net85832), .A2(net84867), .ZN(n1825) );
  INV_X1 U2034 ( .A(\u4/div_shft2[0] ), .ZN(net85831) );
  NAND4_X2 U2035 ( .A1(net11562), .A2(net85831), .A3(net11558), .A4(net11560), 
        .ZN(net84279) );
  NOR2_X4 U2036 ( .A1(net88292), .A2(n1549), .ZN(net84953) );
  INV_X8 U2037 ( .A(net88287), .ZN(net86037) );
  NAND4_X1 U2038 ( .A1(net84996), .A2(net11566), .A3(net85788), .A4(net91375), 
        .ZN(net84990) );
  BUF_X32 U2039 ( .A(\u4/exp_next_mi[5] ), .Z(net91375) );
  NOR2_X4 U2040 ( .A1(net84957), .A2(net89055), .ZN(net84948) );
  NOR2_X4 U2041 ( .A1(n1827), .A2(n1826), .ZN(net89054) );
  NOR2_X2 U2042 ( .A1(net85778), .A2(net84856), .ZN(n1826) );
  NAND2_X4 U2043 ( .A1(net84960), .A2(n1828), .ZN(n1827) );
  NAND2_X4 U2044 ( .A1(net85015), .A2(net84963), .ZN(n1828) );
  INV_X4 U2045 ( .A(net11670), .ZN(net84963) );
  NAND2_X4 U2046 ( .A1(net84202), .A2(net88374), .ZN(net84201) );
  INV_X8 U2047 ( .A(net84201), .ZN(net88721) );
  NAND2_X4 U2048 ( .A1(net83875), .A2(n1829), .ZN(net88374) );
  INV_X8 U2049 ( .A(n1830), .ZN(n1829) );
  NAND3_X4 U2050 ( .A1(n1829), .A2(net83874), .A3(net83875), .ZN(net83871) );
  NAND2_X4 U2051 ( .A1(n1832), .A2(net83861), .ZN(n1830) );
  INV_X4 U2052 ( .A(net84206), .ZN(net83861) );
  NAND2_X2 U2053 ( .A1(net84085), .A2(net83736), .ZN(net84083) );
  AOI211_X4 U2054 ( .C1(n1833), .C2(net83870), .A(n1834), .B(net84204), .ZN(
        net84202) );
  NAND3_X4 U2055 ( .A1(net84074), .A2(n1607), .A3(net84200), .ZN(n1832) );
  NAND2_X4 U2056 ( .A1(n1832), .A2(n1831), .ZN(net83853) );
  AOI21_X2 U2057 ( .B1(n1607), .B2(net84003), .A(net83878), .ZN(n1831) );
  NOR3_X4 U2058 ( .A1(net84372), .A2(n1533), .A3(net84374), .ZN(net84074) );
  NAND2_X2 U2059 ( .A1(net84414), .A2(n1835), .ZN(net84206) );
  NAND2_X2 U2060 ( .A1(n1580), .A2(n1529), .ZN(net84138) );
  INV_X4 U2061 ( .A(net84473), .ZN(net84576) );
  NAND2_X2 U2062 ( .A1(net84474), .A2(net84475), .ZN(net84453) );
  NAND2_X2 U2063 ( .A1(n1554), .A2(net84473), .ZN(net84315) );
  XNOR2_X2 U2064 ( .A(net91555), .B(net11671), .ZN(net84763) );
  AOI22_X4 U2065 ( .A1(net85080), .A2(net85079), .B1(net85081), .B2(net91555), 
        .ZN(net33278) );
  INV_X8 U2066 ( .A(net85174), .ZN(net84758) );
  NAND2_X4 U2067 ( .A1(n1836), .A2(net85108), .ZN(net85174) );
  INV_X8 U2068 ( .A(net85178), .ZN(net85108) );
  NAND2_X2 U2069 ( .A1(net85108), .A2(net84550), .ZN(net85127) );
  NAND3_X4 U2070 ( .A1(net85112), .A2(net85113), .A3(net85108), .ZN(net85111)
         );
  NAND3_X4 U2071 ( .A1(net85176), .A2(net86262), .A3(net85128), .ZN(n1836) );
  INV_X8 U2072 ( .A(net85181), .ZN(net85128) );
  NAND2_X1 U2073 ( .A1(net85128), .A2(net86262), .ZN(net85115) );
  NAND2_X2 U2074 ( .A1(net86262), .A2(net85128), .ZN(net85133) );
  NAND4_X4 U2075 ( .A1(net85128), .A2(net86262), .A3(net85179), .A4(net85180), 
        .ZN(net85084) );
  NAND2_X4 U2076 ( .A1(n1837), .A2(net85220), .ZN(net85181) );
  INV_X8 U2077 ( .A(n1838), .ZN(n1837) );
  NAND2_X4 U2078 ( .A1(net85220), .A2(n1837), .ZN(net77045) );
  NAND3_X4 U2079 ( .A1(net85076), .A2(net85676), .A3(quo[21]), .ZN(n1839) );
  INV_X16 U2080 ( .A(net85678), .ZN(net85676) );
  INV_X16 U2081 ( .A(net85975), .ZN(net85678) );
  INV_X16 U2082 ( .A(net85678), .ZN(net85674) );
  NAND3_X4 U2083 ( .A1(net85342), .A2(quo[3]), .A3(net85678), .ZN(net85051) );
  INV_X4 U2084 ( .A(net85974), .ZN(net85975) );
  INV_X8 U2085 ( .A(net85975), .ZN(net85684) );
  INV_X8 U2086 ( .A(net85351), .ZN(net85076) );
  NAND2_X4 U2087 ( .A1(fract_out_q[12]), .A2(net83780), .ZN(net85349) );
  INV_X8 U2088 ( .A(net85387), .ZN(net83780) );
  NAND2_X4 U2089 ( .A1(net85998), .A2(net85718), .ZN(net85387) );
  NAND2_X4 U2090 ( .A1(net85083), .A2(net85082), .ZN(net84757) );
  INV_X2 U2091 ( .A(net84757), .ZN(net89411) );
  INV_X8 U2092 ( .A(net85084), .ZN(net85082) );
  INV_X8 U2093 ( .A(net76645), .ZN(net85180) );
  INV_X4 U2094 ( .A(n1909), .ZN(net89624) );
  INV_X4 U2095 ( .A(net76254), .ZN(net85179) );
  INV_X1 U2096 ( .A(net85179), .ZN(net86004) );
  INV_X8 U2097 ( .A(net76352), .ZN(net86262) );
  NAND3_X2 U2098 ( .A1(net85247), .A2(net90019), .A3(net85248), .ZN(net76352)
         );
  NAND3_X2 U2099 ( .A1(net85076), .A2(net85676), .A3(quo[22]), .ZN(net85248)
         );
  INV_X4 U2100 ( .A(net85384), .ZN(net85077) );
  NAND2_X2 U2101 ( .A1(net85738), .A2(net85748), .ZN(net85384) );
  INV_X16 U2102 ( .A(net85752), .ZN(net85748) );
  OAI21_X4 U2103 ( .B1(net84974), .B2(net84975), .A(net89372), .ZN(net84956)
         );
  OAI211_X4 U2104 ( .C1(net84967), .C2(net84956), .A(net84968), .B(net84969), 
        .ZN(net84957) );
  NAND2_X4 U2105 ( .A1(\u4/exp_next_mi[5] ), .A2(net85788), .ZN(net84983) );
  INV_X2 U2106 ( .A(n1530), .ZN(net84967) );
  INV_X1 U2107 ( .A(net84975), .ZN(net85017) );
  MUX2_X2 U2108 ( .A(net84598), .B(net84599), .S(net89965), .Z(net84595) );
  NAND2_X1 U2109 ( .A1(net89965), .A2(net85778), .ZN(net84166) );
  NAND2_X4 U2110 ( .A1(net89917), .A2(net89077), .ZN(net84372) );
  INV_X4 U2111 ( .A(net89076), .ZN(net89077) );
  NAND2_X4 U2112 ( .A1(n1840), .A2(n1846), .ZN(net89076) );
  INV_X4 U2113 ( .A(n1845), .ZN(n1846) );
  OAI211_X2 U2114 ( .C1(net86169), .C2(net84408), .A(net84409), .B(net85842), 
        .ZN(net84385) );
  INV_X16 U2115 ( .A(net86160), .ZN(net85842) );
  INV_X8 U2116 ( .A(n1597), .ZN(net86160) );
  INV_X4 U2117 ( .A(net84445), .ZN(net84408) );
  NOR2_X4 U2118 ( .A1(net84408), .A2(net84642), .ZN(net84765) );
  OAI211_X2 U2119 ( .C1(net84408), .C2(net84624), .A(net84625), .B(net84626), 
        .ZN(net84615) );
  INV_X4 U2120 ( .A(n1844), .ZN(n1843) );
  OAI211_X1 U2121 ( .C1(n1841), .C2(n1843), .A(net84421), .B(net85842), .ZN(
        net89975) );
  NOR2_X1 U2122 ( .A1(n1554), .A2(net84312), .ZN(n1844) );
  INV_X4 U2123 ( .A(net84263), .ZN(n1841) );
  NOR3_X2 U2124 ( .A1(net84312), .A2(n1841), .A3(net84314), .ZN(net84276) );
  AOI211_X4 U2125 ( .C1(net84386), .C2(net85842), .A(net84387), .B(n1762), 
        .ZN(net89917) );
  NAND2_X4 U2126 ( .A1(net88721), .A2(n1849), .ZN(net84030) );
  AOI22_X4 U2127 ( .A1(net84027), .A2(net84028), .B1(net84030), .B2(net84029), 
        .ZN(net84026) );
  INV_X4 U2128 ( .A(n1848), .ZN(n1849) );
  NAND2_X4 U2129 ( .A1(net84010), .A2(n1847), .ZN(n1848) );
  NOR2_X4 U2130 ( .A1(net83787), .A2(net85847), .ZN(n1847) );
  NAND2_X4 U2131 ( .A1(net88332), .A2(net85048), .ZN(net85186) );
  NOR3_X4 U2132 ( .A1(net86027), .A2(net85186), .A3(net85285), .ZN(net88605)
         );
  OAI211_X4 U2133 ( .C1(net85186), .C2(net85187), .A(net85143), .B(net85142), 
        .ZN(net85185) );
  INV_X4 U2134 ( .A(net90110), .ZN(net85048) );
  INV_X8 U2135 ( .A(net85161), .ZN(net88332) );
  NAND4_X4 U2136 ( .A1(net88332), .A2(net85159), .A3(net85158), .A4(net85157), 
        .ZN(net85155) );
  OR2_X4 U2137 ( .A1(net85161), .A2(net90110), .ZN(fract_denorm[10]) );
  NAND2_X2 U2138 ( .A1(net84522), .A2(n1764), .ZN(net88950) );
  NAND2_X2 U2139 ( .A1(net84564), .A2(n1850), .ZN(net84518) );
  INV_X2 U2140 ( .A(\u4/N423 ), .ZN(n1850) );
  NOR2_X4 U2141 ( .A1(net84783), .A2(net84519), .ZN(net84777) );
  NAND2_X2 U2142 ( .A1(net86037), .A2(net85854), .ZN(net84015) );
  NOR2_X4 U2143 ( .A1(net84452), .A2(net84490), .ZN(net84770) );
  NAND2_X2 U2144 ( .A1(net84448), .A2(net84764), .ZN(net84452) );
  NAND2_X1 U2145 ( .A1(n1851), .A2(\u4/fract_out_pl1[10] ), .ZN(net84473) );
  INV_X4 U2146 ( .A(net84449), .ZN(n1852) );
  AND2_X2 U2147 ( .A1(net84774), .A2(net84775), .ZN(net89595) );
  INV_X4 U2148 ( .A(net84579), .ZN(net84590) );
  NAND2_X2 U2149 ( .A1(net84448), .A2(net84449), .ZN(net83432) );
  BUF_X32 U2150 ( .A(net84113), .Z(net89716) );
  NAND2_X4 U2151 ( .A1(net84839), .A2(net84840), .ZN(\u4/fract_out[6] ) );
  INV_X8 U2152 ( .A(\u4/fract_out[3] ), .ZN(net84110) );
  INV_X4 U2153 ( .A(net84110), .ZN(net99874) );
  NAND2_X4 U2154 ( .A1(n1749), .A2(net85842), .ZN(net84390) );
  INV_X1 U2155 ( .A(n1535), .ZN(net89987) );
  OAI22_X2 U2156 ( .A1(net84402), .A2(net86016), .B1(n1751), .B2(net84402), 
        .ZN(net86015) );
  INV_X4 U2157 ( .A(net84675), .ZN(n1853) );
  NOR2_X1 U2158 ( .A1(net84480), .A2(n1853), .ZN(net84551) );
  NAND2_X2 U2159 ( .A1(net85828), .A2(n1853), .ZN(net83429) );
  OAI211_X4 U2160 ( .C1(net91015), .C2(net85018), .A(net85020), .B(net85021), 
        .ZN(net84974) );
  INV_X4 U2161 ( .A(net84913), .ZN(net84895) );
  NAND2_X2 U2162 ( .A1(net84895), .A2(net83936), .ZN(net83408) );
  NAND2_X2 U2163 ( .A1(net83951), .A2(net85847), .ZN(net84913) );
  NAND2_X4 U2164 ( .A1(net91177), .A2(net85786), .ZN(net85020) );
  AOI21_X1 U2165 ( .B1(net84822), .B2(net85786), .A(n1571), .ZN(net85018) );
  NAND2_X1 U2166 ( .A1(net84081), .A2(net86174), .ZN(net84347) );
  NAND3_X2 U2167 ( .A1(net84073), .A2(net86174), .A3(net84075), .ZN(net83868)
         );
  NAND2_X2 U2168 ( .A1(n1854), .A2(net83963), .ZN(net84075) );
  INV_X4 U2169 ( .A(net11555), .ZN(net83963) );
  INV_X4 U2170 ( .A(net84168), .ZN(n1854) );
  INV_X4 U2171 ( .A(net84333), .ZN(net84414) );
  OAI21_X2 U2172 ( .B1(net84901), .B2(net84168), .A(net84169), .ZN(net84151)
         );
  NOR2_X4 U2173 ( .A1(net85778), .A2(net84168), .ZN(net84352) );
  OAI21_X4 U2174 ( .B1(net11558), .B2(net84168), .A(net84214), .ZN(net84213)
         );
  NOR2_X4 U2175 ( .A1(net84332), .A2(net84333), .ZN(net84095) );
  NOR2_X4 U2176 ( .A1(net85744), .A2(net85998), .ZN(net85342) );
  INV_X32 U2177 ( .A(net85738), .ZN(net85998) );
  NAND2_X2 U2178 ( .A1(n1855), .A2(n1856), .ZN(net84029) );
  NAND2_X2 U2179 ( .A1(net84033), .A2(n1857), .ZN(n1856) );
  XNOR2_X2 U2180 ( .A(n1858), .B(n1644), .ZN(n1857) );
  INV_X4 U2181 ( .A(net83925), .ZN(n1859) );
  INV_X4 U2182 ( .A(net84044), .ZN(net84033) );
  MUX2_X2 U2183 ( .A(n1862), .B(net84047), .S(sign_mul_r), .Z(n1860) );
  NAND2_X2 U2184 ( .A1(net84047), .A2(net84021), .ZN(n1862) );
  NAND2_X2 U2185 ( .A1(net83779), .A2(opas_r2), .ZN(n1863) );
  OAI211_X4 U2186 ( .C1(net85182), .C2(n1866), .A(net85184), .B(net85185), 
        .ZN(net85083) );
  NOR3_X4 U2187 ( .A1(net85197), .A2(net85199), .A3(n1867), .ZN(net85142) );
  INV_X8 U2188 ( .A(n1864), .ZN(n1867) );
  NOR3_X4 U2189 ( .A1(net85197), .A2(net85199), .A3(n1867), .ZN(n1868) );
  NOR3_X4 U2190 ( .A1(net85234), .A2(n1867), .A3(net88699), .ZN(net85232) );
  INV_X2 U2191 ( .A(n1867), .ZN(net88440) );
  NAND3_X4 U2192 ( .A1(net85369), .A2(quo[13]), .A3(net85674), .ZN(n1864) );
  INV_X4 U2193 ( .A(net85051), .ZN(net85199) );
  INV_X2 U2194 ( .A(net85199), .ZN(net88421) );
  INV_X8 U2195 ( .A(net85193), .ZN(net85143) );
  NAND3_X2 U2196 ( .A1(net85188), .A2(net85143), .A3(n1868), .ZN(n1866) );
  NAND2_X2 U2197 ( .A1(n1868), .A2(net85143), .ZN(net84549) );
  NAND3_X4 U2198 ( .A1(n1865), .A2(net85195), .A3(net85194), .ZN(net85193) );
  INV_X8 U2199 ( .A(n1865), .ZN(net90215) );
  NAND2_X1 U2200 ( .A1(n1865), .A2(net85059), .ZN(net76672) );
  BUF_X32 U2201 ( .A(net84110), .Z(net89485) );
  OAI21_X4 U2202 ( .B1(net84778), .B2(n1870), .A(n1871), .ZN(\u4/fract_out[3] ) );
  NAND2_X4 U2203 ( .A1(\u4/N427 ), .A2(net84522), .ZN(n1871) );
  INV_X4 U2204 ( .A(\u4/N403 ), .ZN(n1870) );
  NAND2_X4 U2205 ( .A1(net84844), .A2(net89250), .ZN(\u4/fract_out[8] ) );
  NAND2_X4 U2206 ( .A1(\u4/N432 ), .A2(net84522), .ZN(net84844) );
  INV_X4 U2207 ( .A(\u4/N409 ), .ZN(net84845) );
  NAND2_X4 U2208 ( .A1(n1869), .A2(net84810), .ZN(net84456) );
  INV_X1 U2209 ( .A(net84456), .ZN(net84322) );
  NAND2_X2 U2210 ( .A1(net84839), .A2(net84840), .ZN(net91512) );
  NAND2_X2 U2211 ( .A1(net84844), .A2(net89250), .ZN(net90252) );
  NAND2_X4 U2212 ( .A1(net84882), .A2(n1872), .ZN(net84778) );
  INV_X4 U2213 ( .A(\u4/N386 ), .ZN(n1872) );
  INV_X4 U2214 ( .A(net84853), .ZN(net84882) );
  NAND2_X4 U2215 ( .A1(n1873), .A2(net83959), .ZN(net91015) );
  OAI21_X4 U2216 ( .B1(n1745), .B2(net85027), .A(net90207), .ZN(net84975) );
  AND2_X2 U2217 ( .A1(net86038), .A2(n1593), .ZN(n1873) );
  NAND3_X2 U2218 ( .A1(net84394), .A2(n1874), .A3(n1875), .ZN(net84386) );
  AOI22_X1 U2219 ( .A1(rmode_r3[1]), .A2(net91353), .B1(net84343), .B2(
        net84398), .ZN(n1875) );
  INV_X4 U2220 ( .A(net84326), .ZN(net84343) );
  NAND2_X2 U2221 ( .A1(net84133), .A2(net84134), .ZN(n1874) );
  NOR3_X4 U2222 ( .A1(net84135), .A2(net84148), .A3(net84393), .ZN(net84387)
         );
  INV_X4 U2223 ( .A(n1597), .ZN(net84393) );
  INV_X4 U2224 ( .A(net83870), .ZN(net83869) );
  NOR2_X4 U2225 ( .A1(n1876), .A2(net84213), .ZN(net84071) );
  NAND4_X2 U2226 ( .A1(net84215), .A2(net84216), .A3(n1877), .A4(net84218), 
        .ZN(n1876) );
  INV_X4 U2227 ( .A(net84080), .ZN(net83878) );
  NAND3_X4 U2228 ( .A1(n1879), .A2(n1878), .A3(net85216), .ZN(net76872) );
  INV_X4 U2229 ( .A(net86060), .ZN(net85317) );
  MUX2_X2 U2230 ( .A(net11485), .B(net86061), .S(net85974), .Z(net86060) );
  NAND3_X4 U2231 ( .A1(n1878), .A2(net85216), .A3(n1879), .ZN(net85178) );
  NAND2_X4 U2232 ( .A1(net85320), .A2(n1881), .ZN(n1880) );
  NAND2_X4 U2233 ( .A1(fract_out_q[14]), .A2(net83780), .ZN(n1881) );
  INV_X8 U2234 ( .A(net85083), .ZN(net89546) );
  NOR2_X2 U2235 ( .A1(net85140), .A2(net85141), .ZN(net85184) );
  NOR2_X4 U2236 ( .A1(net85190), .A2(net85189), .ZN(net85188) );
  NAND3_X2 U2237 ( .A1(net85191), .A2(net86106), .A3(net85192), .ZN(net85190)
         );
  INV_X8 U2238 ( .A(net85150), .ZN(net85192) );
  INV_X4 U2239 ( .A(net99862), .ZN(net85079) );
  OAI21_X4 U2240 ( .B1(net89546), .B2(net88618), .A(net84758), .ZN(net99862)
         );
  OAI21_X2 U2241 ( .B1(net90047), .B2(net84867), .A(net85847), .ZN(n1885) );
  NOR2_X1 U2242 ( .A1(n2151), .A2(net110929), .ZN(n2152) );
  INV_X2 U2243 ( .A(n2632), .ZN(n2633) );
  NOR2_X2 U2244 ( .A1(net83933), .A2(n2632), .ZN(n2582) );
  INV_X4 U2245 ( .A(net77073), .ZN(n1882) );
  INV_X4 U2246 ( .A(n1882), .ZN(n1883) );
  INV_X2 U2247 ( .A(net85115), .ZN(net85112) );
  INV_X4 U2248 ( .A(net88877), .ZN(net110951) );
  INV_X1 U2249 ( .A(net85080), .ZN(net90026) );
  INV_X4 U2250 ( .A(net110929), .ZN(net91467) );
  NAND2_X4 U2251 ( .A1(net88636), .A2(net85089), .ZN(net85085) );
  NAND3_X4 U2252 ( .A1(net85085), .A2(net85215), .A3(net85087), .ZN(net84503)
         );
  AND3_X4 U2253 ( .A1(n1755), .A2(net88551), .A3(net85087), .ZN(net89965) );
  INV_X4 U2254 ( .A(net85089), .ZN(net91109) );
  NAND3_X2 U2255 ( .A1(net85089), .A2(net89935), .A3(net88605), .ZN(net85214)
         );
  OAI21_X4 U2256 ( .B1(n1884), .B2(fract_denorm[9]), .A(net89300), .ZN(
        net85097) );
  INV_X4 U2257 ( .A(net76926), .ZN(n1884) );
  INV_X4 U2258 ( .A(n1884), .ZN(net90037) );
  NAND2_X4 U2259 ( .A1(net85159), .A2(net85158), .ZN(fract_denorm[9]) );
  INV_X8 U2260 ( .A(fract_denorm[9]), .ZN(net90210) );
  INV_X4 U2261 ( .A(net85357), .ZN(net85158) );
  NAND2_X4 U2262 ( .A1(net85260), .A2(net85261), .ZN(net85360) );
  AND3_X4 U2263 ( .A1(net91059), .A2(net90019), .A3(net85248), .ZN(net89300)
         );
  OAI211_X4 U2264 ( .C1(net85137), .C2(net85240), .A(net89300), .B(net85177), 
        .ZN(net85239) );
  NAND2_X4 U2265 ( .A1(net89753), .A2(net84600), .ZN(net84960) );
  NAND2_X2 U2266 ( .A1(n1885), .A2(net85778), .ZN(net84969) );
  NAND2_X4 U2267 ( .A1(net88605), .A2(net89935), .ZN(net86026) );
  OAI211_X4 U2268 ( .C1(net86026), .C2(net91109), .A(net88551), .B(net85087), 
        .ZN(net85081) );
  NAND2_X4 U2269 ( .A1(net85283), .A2(net85240), .ZN(net86027) );
  NAND4_X2 U2270 ( .A1(net85168), .A2(net85171), .A3(net85169), .A4(net85170), 
        .ZN(net85290) );
  NOR3_X4 U2271 ( .A1(n1887), .A2(net90215), .A3(net85060), .ZN(net85283) );
  NAND4_X4 U2272 ( .A1(net85068), .A2(n1886), .A3(net85067), .A4(net85069), 
        .ZN(n1887) );
  NOR2_X4 U2273 ( .A1(n1888), .A2(net85310), .ZN(n1886) );
  INV_X4 U2274 ( .A(n1889), .ZN(n1888) );
  NOR2_X4 U2275 ( .A1(n1888), .A2(net85310), .ZN(net90144) );
  NAND3_X2 U2276 ( .A1(net85736), .A2(net85744), .A3(prod[14]), .ZN(n1889) );
  OAI221_X4 U2277 ( .B1(net85250), .B2(net85251), .C1(net85252), .C2(net85253), 
        .A(net85254), .ZN(net89935) );
  NOR2_X4 U2278 ( .A1(n1890), .A2(n1891), .ZN(net85260) );
  INV_X2 U2279 ( .A(net90064), .ZN(n1893) );
  INV_X4 U2280 ( .A(n1892), .ZN(n1890) );
  NAND3_X2 U2281 ( .A1(net85998), .A2(net85716), .A3(fract_out_q[2]), .ZN(
        n1892) );
  INV_X32 U2282 ( .A(net85722), .ZN(net85716) );
  XNOR2_X2 U2283 ( .A(net84503), .B(net84762), .ZN(net84609) );
  NAND2_X4 U2284 ( .A1(net84503), .A2(div_opa_ldz_r2[0]), .ZN(net84755) );
  INV_X8 U2285 ( .A(net84503), .ZN(net85080) );
  NAND3_X4 U2286 ( .A1(net84503), .A2(net89412), .A3(net89447), .ZN(net84684)
         );
  NAND2_X4 U2287 ( .A1(net85099), .A2(net85098), .ZN(net85215) );
  NAND3_X2 U2288 ( .A1(net85215), .A2(net85214), .A3(net85087), .ZN(net85213)
         );
  INV_X8 U2289 ( .A(net85239), .ZN(net85098) );
  NAND2_X4 U2290 ( .A1(net85098), .A2(net85099), .ZN(net88551) );
  INV_X8 U2291 ( .A(net85285), .ZN(net85177) );
  NAND2_X4 U2292 ( .A1(net85177), .A2(net89943), .ZN(net85176) );
  AOI21_X4 U2293 ( .B1(net77045), .B2(net86262), .A(net85178), .ZN(net85087)
         );
  INV_X2 U2294 ( .A(net91177), .ZN(net90207) );
  NAND2_X2 U2295 ( .A1(net84468), .A2(net84673), .ZN(net84984) );
  INV_X4 U2296 ( .A(net83951), .ZN(net84673) );
  NAND3_X1 U2297 ( .A1(net85786), .A2(net84915), .A3(net84673), .ZN(net84887)
         );
  INV_X4 U2298 ( .A(net84279), .ZN(net85033) );
  NAND3_X4 U2299 ( .A1(net84278), .A2(net84279), .A3(net84280), .ZN(net84277)
         );
  INV_X16 U2300 ( .A(net86037), .ZN(net86038) );
  NOR2_X4 U2301 ( .A1(net85187), .A2(net85189), .ZN(net85254) );
  NOR2_X4 U2302 ( .A1(net85744), .A2(net85728), .ZN(n1894) );
  INV_X16 U2303 ( .A(net85738), .ZN(net85728) );
  NAND2_X4 U2304 ( .A1(net85265), .A2(net85264), .ZN(net85253) );
  INV_X4 U2305 ( .A(net85251), .ZN(net85264) );
  INV_X2 U2306 ( .A(net85163), .ZN(net85265) );
  AOI21_X4 U2307 ( .B1(net85270), .B2(net90080), .A(net85272), .ZN(net85252)
         );
  INV_X8 U2308 ( .A(net85212), .ZN(n1896) );
  CLKBUF_X3 U2309 ( .A(n1896), .Z(net89266) );
  NOR2_X4 U2310 ( .A1(net85039), .A2(net86112), .ZN(net85270) );
  INV_X4 U2311 ( .A(net90292), .ZN(net85250) );
  NAND3_X2 U2312 ( .A1(net85205), .A2(net85280), .A3(net85281), .ZN(net85251)
         );
  NAND3_X4 U2313 ( .A1(n1895), .A2(net85046), .A3(net85045), .ZN(net85189) );
  INV_X8 U2314 ( .A(n1897), .ZN(n1895) );
  NAND3_X2 U2315 ( .A1(n1895), .A2(net85045), .A3(net85046), .ZN(net77073) );
  OAI21_X4 U2316 ( .B1(n1604), .B2(net90031), .A(net85257), .ZN(n1897) );
  OAI21_X4 U2317 ( .B1(n1604), .B2(net90031), .A(net85257), .ZN(net99868) );
  NAND2_X4 U2318 ( .A1(net89856), .A2(net85041), .ZN(net85163) );
  NOR3_X4 U2319 ( .A1(net85163), .A2(net90072), .A3(net85165), .ZN(net84909)
         );
  NAND2_X4 U2320 ( .A1(n1898), .A2(net85210), .ZN(net85272) );
  AOI211_X4 U2321 ( .C1(net85207), .C2(net85206), .A(net89314), .B(net85272), 
        .ZN(net85200) );
  INV_X1 U2322 ( .A(net85272), .ZN(net85162) );
  NOR2_X4 U2323 ( .A1(net85335), .A2(net85336), .ZN(n1898) );
  NAND2_X4 U2324 ( .A1(n2088), .A2(net84990), .ZN(n2093) );
  AOI22_X4 U2325 ( .A1(net85015), .A2(net84992), .B1(net89753), .B2(n1592), 
        .ZN(n2088) );
  INV_X4 U2326 ( .A(net85213), .ZN(net85116) );
  NAND2_X4 U2327 ( .A1(\fract_i2f[7] ), .A2(net85720), .ZN(net85257) );
  INV_X2 U2328 ( .A(net88695), .ZN(net91548) );
  NOR3_X2 U2329 ( .A1(\u4/N414 ), .A2(\u4/N413 ), .A3(\u4/N412 ), .ZN(n2167)
         );
  NAND2_X2 U2330 ( .A1(net91159), .A2(net84870), .ZN(n2097) );
  NAND2_X2 U2331 ( .A1(n1947), .A2(net85131), .ZN(n2055) );
  NOR2_X4 U2332 ( .A1(n1901), .A2(n1556), .ZN(net89856) );
  INV_X8 U2333 ( .A(n1903), .ZN(n1901) );
  NOR2_X4 U2334 ( .A1(n1901), .A2(n1902), .ZN(net85040) );
  NAND3_X4 U2335 ( .A1(net85736), .A2(net85744), .A3(n1904), .ZN(n1903) );
  INV_X4 U2336 ( .A(net88972), .ZN(n1904) );
  NOR2_X4 U2337 ( .A1(net11576), .A2(net85718), .ZN(n1902) );
  INV_X4 U2338 ( .A(net84643), .ZN(net84448) );
  XNOR2_X2 U2339 ( .A(net88896), .B(net84511), .ZN(net88895) );
  BUF_X32 U2340 ( .A(net88895), .Z(net89679) );
  NAND3_X2 U2341 ( .A1(net84910), .A2(net85162), .A3(net84909), .ZN(net85147)
         );
  INV_X4 U2342 ( .A(net85042), .ZN(net85165) );
  INV_X1 U2343 ( .A(net85165), .ZN(net90074) );
  NAND2_X2 U2344 ( .A1(net85393), .A2(net86096), .ZN(net90072) );
  INV_X1 U2345 ( .A(net90072), .ZN(net88585) );
  NAND3_X4 U2346 ( .A1(net85361), .A2(quo[7]), .A3(net85674), .ZN(net85042) );
  NAND2_X4 U2347 ( .A1(net85043), .A2(net85042), .ZN(net90292) );
  NAND2_X4 U2348 ( .A1(net85040), .A2(net85041), .ZN(net89314) );
  NAND2_X4 U2349 ( .A1(net85393), .A2(net86096), .ZN(net85164) );
  NAND3_X2 U2350 ( .A1(net85361), .A2(quo[8]), .A3(net85684), .ZN(net85168) );
  XNOR2_X2 U2351 ( .A(n1761), .B(net84753), .ZN(net83420) );
  INV_X4 U2352 ( .A(net83420), .ZN(net88503) );
  XNOR2_X2 U2353 ( .A(n1761), .B(n1557), .ZN(net90299) );
  NAND3_X2 U2354 ( .A1(net89412), .A2(div_opa_ldz_r2[1]), .A3(net89447), .ZN(
        n1905) );
  INV_X2 U2355 ( .A(net84758), .ZN(net89446) );
  NAND2_X4 U2356 ( .A1(net91467), .A2(net84982), .ZN(net84994) );
  NAND2_X4 U2357 ( .A1(net91467), .A2(net83933), .ZN(net84995) );
  NOR2_X1 U2358 ( .A1(net85854), .A2(n1907), .ZN(net90997) );
  INV_X4 U2359 ( .A(n1906), .ZN(n1907) );
  NAND2_X2 U2360 ( .A1(n1571), .A2(n1596), .ZN(net83844) );
  NAND4_X4 U2361 ( .A1(net85135), .A2(net85147), .A3(net85126), .A4(net85125), 
        .ZN(net85120) );
  INV_X8 U2362 ( .A(net85337), .ZN(net85335) );
  NAND3_X4 U2363 ( .A1(net85736), .A2(net85746), .A3(n1908), .ZN(net85337) );
  INV_X4 U2364 ( .A(net89543), .ZN(n1908) );
  NAND2_X4 U2365 ( .A1(net85203), .A2(net85205), .ZN(net77637) );
  NAND2_X4 U2366 ( .A1(net85032), .A2(n1551), .ZN(net90126) );
  NAND2_X2 U2367 ( .A1(n1551), .A2(net85032), .ZN(net85093) );
  NAND2_X4 U2368 ( .A1(net85032), .A2(n1551), .ZN(net84299) );
  INV_X4 U2369 ( .A(net85133), .ZN(net85107) );
  NAND3_X2 U2370 ( .A1(net85104), .A2(net85105), .A3(net85107), .ZN(net85095)
         );
  INV_X8 U2371 ( .A(net85120), .ZN(net85144) );
  INV_X8 U2372 ( .A(net85155), .ZN(net85125) );
  INV_X1 U2373 ( .A(net85125), .ZN(net89862) );
  INV_X4 U2374 ( .A(net85160), .ZN(net85157) );
  INV_X8 U2375 ( .A(net85166), .ZN(net85135) );
  OAI211_X4 U2376 ( .C1(net84549), .C2(net85124), .A(net85135), .B(net85136), 
        .ZN(net85105) );
  NAND2_X4 U2377 ( .A1(n1909), .A2(n1910), .ZN(net85166) );
  NAND4_X2 U2378 ( .A1(net85168), .A2(net85171), .A3(net85170), .A4(net85169), 
        .ZN(n1911) );
  NAND2_X4 U2379 ( .A1(net85224), .A2(n1913), .ZN(n1912) );
  INV_X8 U2380 ( .A(n1914), .ZN(n1913) );
  NAND2_X4 U2381 ( .A1(net85224), .A2(n1913), .ZN(net76645) );
  NOR2_X4 U2382 ( .A1(net83407), .A2(net83408), .ZN(net83406) );
  INV_X8 U2383 ( .A(net76048), .ZN(net85207) );
  INV_X8 U2384 ( .A(net84301), .ZN(net91159) );
  INV_X1 U2385 ( .A(net85144), .ZN(net89677) );
  AOI211_X4 U2386 ( .C1(net88950), .C2(n1610), .A(net84322), .B(n1916), .ZN(
        n1915) );
  OR2_X2 U2387 ( .A1(net83927), .A2(net84458), .ZN(n1916) );
  NAND3_X2 U2388 ( .A1(net84199), .A2(net89975), .A3(net84200), .ZN(net83863)
         );
  AOI21_X2 U2389 ( .B1(n2346), .B2(n2345), .A(n2344), .ZN(n2347) );
  OR2_X4 U2390 ( .A1(n2099), .A2(net88293), .ZN(n1917) );
  INV_X4 U2391 ( .A(n1571), .ZN(net88293) );
  NOR2_X1 U2392 ( .A1(net11560), .A2(net84856), .ZN(n2078) );
  NOR2_X2 U2393 ( .A1(net84901), .A2(net84856), .ZN(n2091) );
  NOR2_X2 U2394 ( .A1(n1662), .A2(n2567), .ZN(n2568) );
  NAND3_X2 U2395 ( .A1(net83849), .A2(n2554), .A3(n2553), .ZN(n2556) );
  NAND2_X4 U2396 ( .A1(net83861), .A2(net84220), .ZN(n2623) );
  NAND3_X2 U2397 ( .A1(n2436), .A2(n2435), .A3(n2623), .ZN(n2373) );
  OAI21_X4 U2398 ( .B1(n2501), .B2(n2500), .A(n2499), .ZN(n2523) );
  NAND3_X1 U2399 ( .A1(net85342), .A2(quo[0]), .A3(net85684), .ZN(net86106) );
  INV_X16 U2400 ( .A(net86262), .ZN(net86263) );
  NAND2_X2 U2401 ( .A1(n1900), .A2(net85116), .ZN(n1948) );
  NAND3_X2 U2402 ( .A1(quo[10]), .A2(net85752), .A3(net85738), .ZN(n1918) );
  NOR2_X4 U2403 ( .A1(net85744), .A2(net85728), .ZN(n1942) );
  NAND2_X1 U2404 ( .A1(net89266), .A2(net85071), .ZN(n3000) );
  NOR2_X2 U2405 ( .A1(net77815), .A2(net83402), .ZN(net84663) );
  NOR2_X4 U2406 ( .A1(net85730), .A2(net88695), .ZN(n2005) );
  NAND2_X4 U2407 ( .A1(n1754), .A2(n2170), .ZN(n3006) );
  NAND2_X4 U2408 ( .A1(net89819), .A2(net84842), .ZN(n1924) );
  NAND2_X4 U2409 ( .A1(\u4/N431 ), .A2(net84522), .ZN(net84842) );
  NOR3_X4 U2410 ( .A1(\u4/N416 ), .A2(\u4/N417 ), .A3(\u4/N415 ), .ZN(n2166)
         );
  NAND2_X4 U2411 ( .A1(n2162), .A2(n1952), .ZN(\u4/fract_out[1] ) );
  NAND2_X4 U2412 ( .A1(\u4/N429 ), .A2(net84522), .ZN(n2160) );
  INV_X2 U2413 ( .A(net84299), .ZN(net89681) );
  NAND2_X4 U2414 ( .A1(n3096), .A2(net90126), .ZN(n1950) );
  NAND4_X2 U2415 ( .A1(n2491), .A2(n2496), .A3(n1588), .A4(n2477), .ZN(n2480)
         );
  NOR2_X2 U2416 ( .A1(n2707), .A2(net83800), .ZN(n2664) );
  AND2_X2 U2417 ( .A1(net84522), .A2(net84774), .ZN(net91325) );
  NOR2_X4 U2418 ( .A1(div_opa_ldz_r2[1]), .A2(net91159), .ZN(net84754) );
  NAND2_X2 U2419 ( .A1(net85722), .A2(n1657), .ZN(net85281) );
  NOR2_X1 U2420 ( .A1(net88618), .A2(net89546), .ZN(n2056) );
  NOR2_X2 U2421 ( .A1(net85137), .A2(net76645), .ZN(n2045) );
  NAND2_X2 U2422 ( .A1(net89029), .A2(n1661), .ZN(net84652) );
  NAND4_X4 U2423 ( .A1(n2709), .A2(net88319), .A3(n2665), .A4(net83779), .ZN(
        n2666) );
  AOI21_X2 U2424 ( .B1(net84211), .B2(net84128), .A(net89987), .ZN(n2453) );
  NAND2_X4 U2425 ( .A1(net85116), .A2(n1900), .ZN(n2139) );
  NAND2_X4 U2426 ( .A1(\u4/N430 ), .A2(net84522), .ZN(net84839) );
  INV_X8 U2427 ( .A(net91128), .ZN(net83407) );
  CLKBUF_X3 U2428 ( .A(net84702), .Z(net91128) );
  NOR2_X4 U2429 ( .A1(net99868), .A2(n2049), .ZN(n2051) );
  NAND2_X2 U2430 ( .A1(net85720), .A2(n1658), .ZN(n2022) );
  NAND2_X1 U2431 ( .A1(net85720), .A2(n1667), .ZN(net85374) );
  AND2_X2 U2432 ( .A1(net84869), .A2(n2054), .ZN(net91112) );
  OAI21_X4 U2433 ( .B1(n2216), .B2(n2250), .A(n2215), .ZN(net84511) );
  NOR2_X4 U2434 ( .A1(net85710), .A2(net89964), .ZN(n2216) );
  AOI22_X4 U2435 ( .A1(n2018), .A2(net85684), .B1(n2017), .B2(fract_out_q[10]), 
        .ZN(n2038) );
  NAND4_X4 U2436 ( .A1(n2051), .A2(n1970), .A3(net85045), .A4(net85046), .ZN(
        n2052) );
  NAND2_X1 U2437 ( .A1(net85722), .A2(n1668), .ZN(n2029) );
  NAND2_X2 U2438 ( .A1(net85722), .A2(n1659), .ZN(n2069) );
  NAND2_X4 U2439 ( .A1(net89680), .A2(net89681), .ZN(n1935) );
  INV_X1 U2440 ( .A(net83407), .ZN(net91095) );
  AND4_X4 U2441 ( .A1(net85061), .A2(n2043), .A3(n2067), .A4(n2066), .ZN(n1971) );
  INV_X1 U2442 ( .A(net86263), .ZN(net84601) );
  INV_X4 U2443 ( .A(net90031), .ZN(net86125) );
  NAND2_X4 U2444 ( .A1(net85144), .A2(n2053), .ZN(net85104) );
  NOR2_X4 U2445 ( .A1(n2035), .A2(net89998), .ZN(net88287) );
  BUF_X8 U2446 ( .A(net83780), .Z(net91075) );
  INV_X4 U2447 ( .A(net77045), .ZN(net91069) );
  INV_X8 U2448 ( .A(net91069), .ZN(net91070) );
  NAND2_X4 U2449 ( .A1(net84749), .A2(n2190), .ZN(n2443) );
  NAND3_X4 U2450 ( .A1(n1930), .A2(net85123), .A3(net84531), .ZN(n2190) );
  NAND2_X4 U2451 ( .A1(net85091), .A2(net85095), .ZN(n1972) );
  NAND4_X2 U2452 ( .A1(net85192), .A2(net85191), .A3(n1969), .A4(n2050), .ZN(
        net76926) );
  NAND2_X4 U2453 ( .A1(net91056), .A2(net91057), .ZN(net77815) );
  BUF_X32 U2454 ( .A(\u4/fi_ldz_mi1[3] ), .Z(n1919) );
  INV_X4 U2455 ( .A(n2448), .ZN(\u4/fi_ldz_mi1[3] ) );
  NAND3_X1 U2456 ( .A1(n2040), .A2(quo[0]), .A3(net85684), .ZN(n1970) );
  XNOR2_X1 U2457 ( .A(net91112), .B(n2410), .ZN(n2411) );
  BUF_X32 U2458 ( .A(net84869), .Z(net91047) );
  NAND2_X2 U2459 ( .A1(net84953), .A2(n2099), .ZN(net84968) );
  NAND2_X4 U2460 ( .A1(n2162), .A2(n1952), .ZN(n1920) );
  NAND2_X4 U2461 ( .A1(net85778), .A2(net90026), .ZN(n2250) );
  NAND2_X2 U2462 ( .A1(net84600), .A2(net90026), .ZN(n2968) );
  INV_X2 U2463 ( .A(net85081), .ZN(net85096) );
  NAND2_X2 U2464 ( .A1(n2009), .A2(prod[15]), .ZN(n2008) );
  INV_X4 U2465 ( .A(net84310), .ZN(net90302) );
  NOR3_X4 U2466 ( .A1(n1937), .A2(net85748), .A3(net85998), .ZN(n2018) );
  NOR2_X4 U2467 ( .A1(net85748), .A2(net85730), .ZN(n2040) );
  INV_X8 U2468 ( .A(net90210), .ZN(net90211) );
  INV_X4 U2469 ( .A(n1918), .ZN(n1921) );
  NAND3_X2 U2470 ( .A1(net85369), .A2(quo[20]), .A3(net85674), .ZN(n2027) );
  NAND2_X2 U2471 ( .A1(n2047), .A2(net85203), .ZN(n2048) );
  NOR2_X1 U2472 ( .A1(net84672), .A2(net85004), .ZN(n2154) );
  OAI21_X1 U2473 ( .B1(n2154), .B2(net84867), .A(n2153), .ZN(n2157) );
  NOR3_X1 U2474 ( .A1(net83421), .A2(net84867), .A3(n2154), .ZN(n2084) );
  NOR2_X1 U2475 ( .A1(n2580), .A2(n2579), .ZN(n2581) );
  NAND3_X2 U2476 ( .A1(n2095), .A2(net85006), .A3(n2094), .ZN(n2096) );
  OAI21_X2 U2477 ( .B1(net91095), .B2(n2219), .A(n2218), .ZN(n2261) );
  NOR2_X4 U2478 ( .A1(net85744), .A2(net85998), .ZN(n1922) );
  NAND2_X4 U2479 ( .A1(net84609), .A2(net85832), .ZN(net84610) );
  NAND3_X2 U2480 ( .A1(net84662), .A2(net84661), .A3(net84660), .ZN(net84655)
         );
  NAND2_X4 U2481 ( .A1(net83969), .A2(net85853), .ZN(n872) );
  NAND2_X4 U2482 ( .A1(net84236), .A2(net85853), .ZN(n2991) );
  NAND3_X4 U2483 ( .A1(net85736), .A2(net85752), .A3(net85716), .ZN(net85853)
         );
  INV_X4 U2484 ( .A(net85192), .ZN(net90124) );
  INV_X1 U2485 ( .A(net85131), .ZN(net90115) );
  INV_X8 U2486 ( .A(net77161), .ZN(net85131) );
  INV_X8 U2487 ( .A(net11562), .ZN(net83993) );
  INV_X1 U2488 ( .A(exp_r[1]), .ZN(net84901) );
  INV_X1 U2489 ( .A(exp_r[1]), .ZN(net84167) );
  NOR2_X4 U2490 ( .A1(net85744), .A2(net85730), .ZN(n2001) );
  NOR2_X2 U2491 ( .A1(n3077), .A2(net85716), .ZN(n2003) );
  OAI21_X2 U2492 ( .B1(net88319), .B2(n2607), .A(n2606), .ZN(n2614) );
  NAND3_X2 U2493 ( .A1(net85998), .A2(net85716), .A3(fract_out_q[9]), .ZN(
        net85169) );
  NOR3_X4 U2494 ( .A1(n2052), .A2(net90124), .A3(n1921), .ZN(net85126) );
  NOR2_X4 U2495 ( .A1(net85744), .A2(net85728), .ZN(n2016) );
  NAND3_X2 U2496 ( .A1(n2098), .A2(n2097), .A3(n2096), .ZN(\u4/shift_left [1])
         );
  INV_X2 U2497 ( .A(net84684), .ZN(net89680) );
  INV_X1 U2498 ( .A(net89964), .ZN(net84310) );
  INV_X2 U2499 ( .A(net84549), .ZN(net85123) );
  NOR2_X1 U2500 ( .A1(net84548), .A2(net84549), .ZN(n2300) );
  NAND3_X1 U2501 ( .A1(net84322), .A2(net88950), .A3(n1610), .ZN(n2302) );
  NAND3_X1 U2502 ( .A1(net83946), .A2(net88950), .A3(n2574), .ZN(n2575) );
  NAND2_X4 U2503 ( .A1(net85738), .A2(net85748), .ZN(net90031) );
  NAND3_X2 U2504 ( .A1(n2034), .A2(quo[10]), .A3(net85684), .ZN(n1923) );
  INV_X2 U2505 ( .A(net89933), .ZN(net84107) );
  BUF_X4 U2506 ( .A(net76672), .Z(net90007) );
  INV_X8 U2507 ( .A(net85718), .ZN(net89998) );
  NOR2_X2 U2508 ( .A1(net85114), .A2(net85115), .ZN(net84550) );
  NAND3_X1 U2509 ( .A1(n2321), .A2(n2474), .A3(n2498), .ZN(n1925) );
  NAND3_X2 U2510 ( .A1(net89029), .A2(net84571), .A3(n1661), .ZN(net84568) );
  NAND2_X4 U2511 ( .A1(net84684), .A2(n1948), .ZN(net89964) );
  NAND3_X2 U2512 ( .A1(n2068), .A2(n2070), .A3(n2069), .ZN(net85234) );
  OAI22_X4 U2513 ( .A1(net84107), .A2(n1961), .B1(n2513), .B2(n2511), .ZN(
        n2680) );
  NOR2_X4 U2514 ( .A1(net85744), .A2(net85730), .ZN(n2024) );
  NOR2_X4 U2515 ( .A1(net85744), .A2(net85728), .ZN(net85361) );
  INV_X2 U2516 ( .A(n1924), .ZN(n2503) );
  OAI21_X2 U2517 ( .B1(n2143), .B2(net84890), .A(n2142), .ZN(n2144) );
  NOR2_X1 U2518 ( .A1(net84191), .A2(net84079), .ZN(n2472) );
  NAND2_X1 U2519 ( .A1(net89266), .A2(net85071), .ZN(n1926) );
  NAND2_X1 U2520 ( .A1(net89266), .A2(net85071), .ZN(n1927) );
  NOR3_X1 U2521 ( .A1(net84146), .A2(net84312), .A3(net86016), .ZN(n2362) );
  NAND3_X1 U2522 ( .A1(n2478), .A2(net84150), .A3(net84081), .ZN(n2479) );
  AND3_X4 U2523 ( .A1(n2036), .A2(n2038), .A3(n2037), .ZN(net89943) );
  OAI21_X4 U2524 ( .B1(n2385), .B2(n2384), .A(net84095), .ZN(n1928) );
  BUF_X32 U2525 ( .A(\u4/fi_ldz_mi1[2] ), .Z(n1929) );
  BUF_X32 U2526 ( .A(n845), .Z(net89926) );
  INV_X1 U2527 ( .A(net88503), .ZN(net89924) );
  INV_X1 U2528 ( .A(n1919), .ZN(n1931) );
  INV_X2 U2529 ( .A(net89862), .ZN(net89863) );
  NAND2_X4 U2530 ( .A1(opas_r2), .A2(net83936), .ZN(n2159) );
  NAND2_X4 U2531 ( .A1(net85194), .A2(net85195), .ZN(net85060) );
  NAND2_X4 U2532 ( .A1(net89817), .A2(\u4/N407 ), .ZN(net89819) );
  INV_X1 U2533 ( .A(net84778), .ZN(net89817) );
  INV_X1 U2534 ( .A(\u4/fract_out[1] ), .ZN(net84103) );
  NOR2_X4 U2535 ( .A1(\u4/N421 ), .A2(\u4/N422 ), .ZN(n2164) );
  INV_X4 U2536 ( .A(net84763), .ZN(net89120) );
  XNOR2_X2 U2537 ( .A(net84702), .B(n2306), .ZN(net88896) );
  NOR2_X4 U2538 ( .A1(net84151), .A2(n1639), .ZN(n2527) );
  NOR2_X1 U2539 ( .A1(n2483), .A2(n2482), .ZN(n2489) );
  OAI21_X1 U2540 ( .B1(n2487), .B2(n2486), .A(n2485), .ZN(n2488) );
  NAND3_X2 U2541 ( .A1(net84315), .A2(net84263), .A3(net84366), .ZN(n2596) );
  NAND2_X4 U2542 ( .A1(n2341), .A2(n2340), .ZN(n2521) );
  NAND2_X4 U2543 ( .A1(n2330), .A2(n2416), .ZN(n2341) );
  INV_X1 U2544 ( .A(net89753), .ZN(net89741) );
  INV_X8 U2545 ( .A(net30297), .ZN(net83296) );
  NAND2_X1 U2546 ( .A1(n2433), .A2(n2515), .ZN(n2434) );
  NOR2_X4 U2547 ( .A1(n2515), .A2(n2674), .ZN(n2516) );
  NAND2_X2 U2548 ( .A1(net84421), .A2(n2360), .ZN(n2361) );
  NAND2_X4 U2549 ( .A1(n2356), .A2(net84371), .ZN(net84149) );
  NAND2_X2 U2550 ( .A1(net84010), .A2(net88721), .ZN(n2618) );
  INV_X4 U2551 ( .A(n2706), .ZN(n2625) );
  NAND3_X2 U2552 ( .A1(net84347), .A2(n2373), .A3(n1933), .ZN(n2375) );
  INV_X4 U2553 ( .A(n1932), .ZN(n1933) );
  NAND2_X1 U2554 ( .A1(net83878), .A2(n2623), .ZN(n2372) );
  NAND2_X4 U2555 ( .A1(n2336), .A2(n2454), .ZN(n2333) );
  NOR2_X1 U2556 ( .A1(n2706), .A2(net83736), .ZN(n2663) );
  NAND2_X2 U2557 ( .A1(net84684), .A2(net90126), .ZN(n1934) );
  NAND2_X4 U2558 ( .A1(n1935), .A2(n1934), .ZN(net84702) );
  NAND2_X2 U2559 ( .A1(net84755), .A2(net84763), .ZN(n1945) );
  NOR3_X1 U2560 ( .A1(n2080), .A2(n2079), .A3(n2078), .ZN(n2086) );
  INV_X1 U2561 ( .A(net89679), .ZN(net83414) );
  INV_X1 U2562 ( .A(net90047), .ZN(net85004) );
  NOR2_X1 U2563 ( .A1(net90268), .A2(net83421), .ZN(n2188) );
  NOR2_X4 U2564 ( .A1(net85998), .A2(net85752), .ZN(n1936) );
  NAND2_X2 U2565 ( .A1(\u4/N423 ), .A2(net84522), .ZN(n2275) );
  NAND2_X4 U2566 ( .A1(n1949), .A2(net88877), .ZN(n1951) );
  OAI21_X2 U2567 ( .B1(n2468), .B2(net84297), .A(net84298), .ZN(n2444) );
  INV_X1 U2568 ( .A(n2253), .ZN(n2254) );
  INV_X2 U2569 ( .A(n2196), .ZN(n2199) );
  NAND2_X1 U2570 ( .A1(n2401), .A2(n2222), .ZN(n2223) );
  NOR2_X4 U2571 ( .A1(net85744), .A2(net85998), .ZN(net85369) );
  OAI21_X1 U2572 ( .B1(net85676), .B2(n2572), .A(n2571), .ZN(n2629) );
  NAND2_X1 U2573 ( .A1(net85676), .A2(n2309), .ZN(net84626) );
  AOI22_X1 U2574 ( .A1(net83416), .A2(n2269), .B1(net85676), .B2(n2366), .ZN(
        n2270) );
  NAND3_X1 U2575 ( .A1(net85076), .A2(net85676), .A3(quo[2]), .ZN(n2063) );
  INV_X4 U2576 ( .A(net85365), .ZN(net85224) );
  INV_X4 U2577 ( .A(net85676), .ZN(net86113) );
  AOI21_X4 U2578 ( .B1(net89078), .B2(n1940), .A(net83990), .ZN(n3008) );
  NOR2_X2 U2579 ( .A1(n3078), .A2(net85716), .ZN(n2012) );
  OAI21_X4 U2580 ( .B1(n2670), .B2(n2669), .A(n2668), .ZN(n2672) );
  NAND4_X2 U2581 ( .A1(net90144), .A2(net85067), .A3(net85068), .A4(net85069), 
        .ZN(n3002) );
  NOR2_X2 U2582 ( .A1(net85730), .A2(n1650), .ZN(net85227) );
  NAND2_X4 U2583 ( .A1(\u4/N425 ), .A2(net84522), .ZN(n2162) );
  NAND2_X1 U2584 ( .A1(n2695), .A2(n2674), .ZN(n2675) );
  NOR2_X2 U2585 ( .A1(n1768), .A2(net84329), .ZN(n2382) );
  NAND2_X1 U2586 ( .A1(net84371), .A2(net83296), .ZN(n1938) );
  NAND2_X1 U2587 ( .A1(n1648), .A2(net30297), .ZN(n1939) );
  NAND2_X2 U2588 ( .A1(n1938), .A2(n1939), .ZN(n2435) );
  AOI21_X2 U2589 ( .B1(n2675), .B2(n1546), .A(n2683), .ZN(N221) );
  NAND3_X2 U2590 ( .A1(n2425), .A2(net85842), .A3(n2365), .ZN(n2461) );
  INV_X8 U2591 ( .A(net85164), .ZN(net85043) );
  INV_X1 U2592 ( .A(net90252), .ZN(net84119) );
  NOR2_X4 U2593 ( .A1(net85998), .A2(net85752), .ZN(n2039) );
  AOI21_X1 U2594 ( .B1(net91047), .B2(net84870), .A(n2152), .ZN(net84847) );
  NOR2_X1 U2595 ( .A1(n2234), .A2(net89741), .ZN(n2080) );
  NAND2_X2 U2596 ( .A1(net91150), .A2(\u4/N408 ), .ZN(net89250) );
  NAND3_X2 U2597 ( .A1(n2087), .A2(n2086), .A3(n2085), .ZN(\u4/shift_left [2])
         );
  NAND2_X4 U2598 ( .A1(n2356), .A2(net84371), .ZN(net84421) );
  AOI21_X2 U2599 ( .B1(n2644), .B2(n2643), .A(net83827), .ZN(n2645) );
  NAND3_X2 U2600 ( .A1(n2321), .A2(n2474), .A3(n2498), .ZN(n2336) );
  NAND2_X1 U2601 ( .A1(n2667), .A2(net83787), .ZN(n1943) );
  INV_X4 U2602 ( .A(n1943), .ZN(n1944) );
  NAND2_X1 U2603 ( .A1(net91542), .A2(net84138), .ZN(n2497) );
  NAND3_X2 U2604 ( .A1(net85790), .A2(net85010), .A3(net83849), .ZN(net84856)
         );
  NAND3_X2 U2605 ( .A1(net85716), .A2(n1656), .A3(net85728), .ZN(net85045) );
  AOI21_X2 U2606 ( .B1(n2681), .B2(n1546), .A(n2683), .ZN(N224) );
  AOI21_X2 U2607 ( .B1(n2677), .B2(n1546), .A(n2683), .ZN(N222) );
  AOI21_X2 U2608 ( .B1(n2679), .B2(n1546), .A(n2683), .ZN(N223) );
  AOI21_X2 U2609 ( .B1(n2684), .B2(n1546), .A(n2683), .ZN(N225) );
  NAND4_X4 U2610 ( .A1(net85061), .A2(n2043), .A3(n2067), .A4(n2066), .ZN(
        net85141) );
  INV_X1 U2611 ( .A(net85205), .ZN(net85204) );
  NAND2_X4 U2612 ( .A1(net85037), .A2(net85038), .ZN(n2999) );
  NOR2_X4 U2613 ( .A1(net85744), .A2(net85732), .ZN(net89129) );
  NAND2_X4 U2614 ( .A1(net89120), .A2(net89121), .ZN(n1946) );
  NAND2_X4 U2615 ( .A1(n1945), .A2(n1946), .ZN(net84761) );
  INV_X4 U2616 ( .A(n2035), .ZN(n1955) );
  NAND2_X4 U2617 ( .A1(net85194), .A2(net85195), .ZN(n2041) );
  NAND2_X2 U2618 ( .A1(n2621), .A2(n2620), .ZN(n3007) );
  NOR2_X2 U2619 ( .A1(n2616), .A2(n2617), .ZN(n2621) );
  NAND2_X4 U2620 ( .A1(net84421), .A2(net83296), .ZN(n2491) );
  OAI22_X4 U2621 ( .A1(n2186), .A2(net84777), .B1(net84778), .B2(n2185), .ZN(
        net84775) );
  AND3_X4 U2622 ( .A1(n2036), .A2(n2037), .A3(n2038), .ZN(n1947) );
  INV_X8 U2623 ( .A(n1947), .ZN(n3003) );
  OAI21_X2 U2624 ( .B1(n2233), .B2(n2968), .A(n2232), .ZN(n2965) );
  OAI21_X1 U2625 ( .B1(net85832), .B2(net90122), .A(net84610), .ZN(n2269) );
  OAI21_X2 U2626 ( .B1(n2422), .B2(net84502), .A(n2421), .ZN(net84469) );
  NAND4_X2 U2627 ( .A1(net85171), .A2(net85168), .A3(net85169), .A4(net85170), 
        .ZN(net76254) );
  NAND2_X2 U2628 ( .A1(net90299), .A2(net83421), .ZN(n1958) );
  INV_X4 U2629 ( .A(n3096), .ZN(n1949) );
  NAND2_X4 U2630 ( .A1(net90074), .A2(net88585), .ZN(n2998) );
  NAND4_X4 U2631 ( .A1(n2519), .A2(n2518), .A3(n2517), .A4(n2516), .ZN(
        net83787) );
  NAND2_X4 U2632 ( .A1(n1899), .A2(n2170), .ZN(net84814) );
  OR2_X4 U2633 ( .A1(net84778), .A2(n2163), .ZN(n1952) );
  NAND3_X2 U2634 ( .A1(n2040), .A2(quo[10]), .A3(net85684), .ZN(n2025) );
  NAND2_X4 U2635 ( .A1(n2462), .A2(n2363), .ZN(net84168) );
  INV_X8 U2636 ( .A(net85051), .ZN(net88699) );
  NOR3_X1 U2637 ( .A1(prod[0]), .A2(prod[10]), .A3(prod[1]), .ZN(n2648) );
  INV_X1 U2638 ( .A(n1528), .ZN(net84115) );
  NAND2_X4 U2639 ( .A1(net88503), .A2(\u4/exp_in_pl1[2] ), .ZN(n1959) );
  NAND2_X1 U2640 ( .A1(net84983), .A2(net84822), .ZN(n2579) );
  INV_X16 U2641 ( .A(net84858), .ZN(\u4/f2i_shft[3] ) );
  NAND2_X4 U2642 ( .A1(n2029), .A2(n2030), .ZN(net85039) );
  NAND2_X4 U2643 ( .A1(n1956), .A2(net88566), .ZN(n1957) );
  NAND2_X4 U2644 ( .A1(n1957), .A2(n2045), .ZN(net85099) );
  INV_X4 U2645 ( .A(n2046), .ZN(n1956) );
  NOR2_X4 U2646 ( .A1(n2044), .A2(net85141), .ZN(n2046) );
  OAI21_X1 U2647 ( .B1(n2192), .B2(net110951), .A(n2191), .ZN(n2196) );
  NAND2_X4 U2648 ( .A1(n1959), .A2(n1958), .ZN(net83419) );
  XNOR2_X1 U2649 ( .A(net84167), .B(net90302), .ZN(n2481) );
  NAND2_X1 U2650 ( .A1(net90302), .A2(net84167), .ZN(n2393) );
  NAND2_X1 U2651 ( .A1(net84511), .A2(n2217), .ZN(n2218) );
  NOR2_X1 U2652 ( .A1(net84511), .A2(n2217), .ZN(n2219) );
  NOR2_X1 U2653 ( .A1(n1592), .A2(net89964), .ZN(n2233) );
  NAND2_X1 U2654 ( .A1(n1592), .A2(net89964), .ZN(n2232) );
  XNOR2_X1 U2655 ( .A(net89964), .B(net85710), .ZN(n2251) );
  INV_X1 U2656 ( .A(net85207), .ZN(net88545) );
  NAND2_X4 U2657 ( .A1(net83993), .A2(net83967), .ZN(net85313) );
  NOR2_X2 U2658 ( .A1(net85211), .A2(net85212), .ZN(net85206) );
  INV_X1 U2659 ( .A(net91159), .ZN(net88510) );
  INV_X1 U2660 ( .A(net89948), .ZN(net84191) );
  NOR2_X4 U2661 ( .A1(net85738), .A2(net85722), .ZN(n2017) );
  AOI21_X2 U2662 ( .B1(n2398), .B2(n2449), .A(n2397), .ZN(n2399) );
  NAND2_X4 U2663 ( .A1(n2005), .A2(prod[2]), .ZN(n2030) );
  NOR3_X1 U2664 ( .A1(prod[14]), .A2(prod[15]), .A3(prod[16]), .ZN(n2649) );
  NOR2_X1 U2665 ( .A1(n3001), .A2(net88545), .ZN(net84911) );
  NAND3_X2 U2666 ( .A1(n2006), .A2(n2007), .A3(n2008), .ZN(net85365) );
  NAND2_X1 U2667 ( .A1(n1919), .A2(net84305), .ZN(n2398) );
  NOR2_X1 U2668 ( .A1(n1919), .A2(net84305), .ZN(n2397) );
  NOR2_X1 U2669 ( .A1(net84601), .A2(net84602), .ZN(n2273) );
  NOR2_X1 U2670 ( .A1(net83414), .A2(n2307), .ZN(n2308) );
  NAND2_X4 U2671 ( .A1(n2061), .A2(n2405), .ZN(\u4/f2i_shft[4] ) );
  NAND3_X2 U2672 ( .A1(n2075), .A2(net84290), .A3(net84305), .ZN(n2226) );
  NAND2_X4 U2673 ( .A1(net11566), .A2(net83933), .ZN(net84236) );
  NOR2_X2 U2674 ( .A1(net85730), .A2(net85752), .ZN(n2009) );
  AND2_X2 U2675 ( .A1(exp_r[2]), .A2(net83993), .ZN(\u4/add_407/carry [3]) );
  AOI22_X1 U2676 ( .A1(n2393), .A2(net84166), .B1(net84310), .B2(net83993), 
        .ZN(n2465) );
  XOR2_X1 U2677 ( .A(exp_r[2]), .B(net83993), .Z(n2119) );
  NOR2_X1 U2678 ( .A1(div_opa_ldz_r2[1]), .A2(net83993), .ZN(n2121) );
  NAND2_X1 U2679 ( .A1(net83993), .A2(div_opa_ldz_r2[1]), .ZN(n2120) );
  NAND2_X1 U2680 ( .A1(net83993), .A2(net11671), .ZN(n2102) );
  XNOR2_X1 U2681 ( .A(div_opa_ldz_r2[1]), .B(net83993), .ZN(n2133) );
  NAND2_X1 U2682 ( .A1(net85030), .A2(net11560), .ZN(n2225) );
  NAND3_X4 U2683 ( .A1(n2074), .A2(net88440), .A3(net88421), .ZN(n3005) );
  OAI211_X1 U2684 ( .C1(net83987), .C2(n2551), .A(n2550), .B(net83990), .ZN(
        n2557) );
  OAI21_X1 U2685 ( .B1(n2364), .B2(n2443), .A(net83990), .ZN(n2566) );
  NAND2_X1 U2686 ( .A1(n2223), .A2(net83990), .ZN(n2242) );
  NAND3_X2 U2687 ( .A1(net85736), .A2(net85746), .A3(prod[1]), .ZN(n2032) );
  NAND3_X2 U2688 ( .A1(net85744), .A2(net85736), .A3(prod[18]), .ZN(n2011) );
  NAND3_X2 U2689 ( .A1(net85746), .A2(net85736), .A3(prod[13]), .ZN(n2042) );
  NAND3_X2 U2690 ( .A1(net85998), .A2(net85716), .A3(fract_out_q[6]), .ZN(
        n2066) );
  NOR2_X2 U2691 ( .A1(net85744), .A2(net85728), .ZN(n2033) );
  NOR2_X2 U2692 ( .A1(net91548), .A2(net85728), .ZN(n2034) );
  NOR2_X2 U2693 ( .A1(net85748), .A2(net85728), .ZN(n2014) );
  NAND3_X2 U2694 ( .A1(net85998), .A2(net85716), .A3(fract_out_q[7]), .ZN(
        net85069) );
  NAND3_X2 U2695 ( .A1(net85998), .A2(net85716), .A3(fract_out_q[11]), .ZN(
        n2026) );
  NAND2_X2 U2696 ( .A1(fract_out_q[8]), .A2(n2017), .ZN(n2007) );
  AND3_X4 U2697 ( .A1(n2426), .A2(net85794), .A3(net88500), .ZN(n2392) );
  NAND2_X1 U2698 ( .A1(net86169), .A2(net91404), .ZN(net84312) );
  OAI21_X1 U2699 ( .B1(net88500), .B2(net84887), .A(n2144), .ZN(
        \u4/shift_right [1]) );
  NAND3_X1 U2700 ( .A1(net90047), .A2(net84982), .A3(net84983), .ZN(n2094) );
  NOR2_X4 U2701 ( .A1(n2099), .A2(net88293), .ZN(net88292) );
  INV_X1 U2702 ( .A(n2068), .ZN(n2073) );
  AOI22_X1 U2703 ( .A1(n2400), .A2(net84160), .B1(net88510), .B2(net85712), 
        .ZN(n2468) );
  NAND2_X1 U2706 ( .A1(net90126), .A2(net84684), .ZN(n2222) );
  NOR2_X1 U2707 ( .A1(net110951), .A2(net84684), .ZN(n2253) );
  NOR2_X2 U2708 ( .A1(n3076), .A2(net85718), .ZN(net85310) );
  AOI21_X2 U2709 ( .B1(n2664), .B2(n2663), .A(n2669), .ZN(n2673) );
  NAND4_X4 U2710 ( .A1(n2598), .A2(net83844), .A3(net83855), .A4(net83906), 
        .ZN(n2702) );
  XNOR2_X1 U2711 ( .A(n1931), .B(net83968), .ZN(n2450) );
  NAND2_X4 U2712 ( .A1(net84869), .A2(n2054), .ZN(net83990) );
  INV_X1 U2713 ( .A(fract_denorm[10]), .ZN(net84532) );
  AOI22_X4 U2714 ( .A1(net89998), .A2(n1633), .B1(prod[19]), .B2(net86125), 
        .ZN(net85220) );
  AOI21_X1 U2715 ( .B1(net90268), .B2(net83421), .A(net89924), .ZN(n2189) );
  NOR2_X1 U2716 ( .A1(\u4/fract_out_pl1[10] ), .A2(net83429), .ZN(n2962) );
  INV_X8 U2717 ( .A(n2514), .ZN(n1960) );
  OAI21_X2 U2718 ( .B1(net83754), .B2(n2693), .A(n2692), .ZN(N229) );
  OAI21_X2 U2719 ( .B1(net83754), .B2(n2690), .A(n2692), .ZN(N228) );
  OAI21_X2 U2720 ( .B1(net83754), .B2(n2688), .A(n2692), .ZN(N227) );
  OAI21_X2 U2721 ( .B1(net83754), .B2(n2686), .A(n2692), .ZN(N226) );
  OAI21_X2 U2722 ( .B1(net83754), .B2(n2434), .A(n2692), .ZN(N220) );
  NAND2_X4 U2723 ( .A1(n2702), .A2(net85790), .ZN(n2609) );
  AOI21_X4 U2724 ( .B1(n2609), .B2(n2610), .A(n2608), .ZN(n2617) );
  NAND2_X1 U2725 ( .A1(net84421), .A2(net30297), .ZN(n2478) );
  NAND2_X1 U2726 ( .A1(net84421), .A2(net84150), .ZN(n2493) );
  NOR2_X2 U2727 ( .A1(net83853), .A2(n2628), .ZN(n2642) );
  AOI21_X2 U2728 ( .B1(n1648), .B2(n2496), .A(n2996), .ZN(n2350) );
  NAND4_X1 U2729 ( .A1(n2496), .A2(n2491), .A3(net84081), .A4(net86169), .ZN(
        n2337) );
  NAND2_X4 U2730 ( .A1(net84983), .A2(net84982), .ZN(n2081) );
  NAND3_X2 U2731 ( .A1(net85116), .A2(n2057), .A3(n2056), .ZN(n2059) );
  INV_X1 U2732 ( .A(net86169), .ZN(net84128) );
  INV_X2 U2733 ( .A(net85060), .ZN(net85059) );
  INV_X1 U2734 ( .A(n1929), .ZN(n2394) );
  NAND2_X1 U2735 ( .A1(exp_r[2]), .A2(n2394), .ZN(n2395) );
  NOR2_X1 U2736 ( .A1(exp_r[2]), .A2(n2394), .ZN(n2396) );
  INV_X8 U2737 ( .A(net85103), .ZN(net85032) );
  NAND2_X4 U2738 ( .A1(n1954), .A2(net85105), .ZN(net85103) );
  NAND2_X4 U2739 ( .A1(net85738), .A2(net85752), .ZN(net85351) );
  NAND2_X1 U2740 ( .A1(opa_00), .A2(net84015), .ZN(n2352) );
  OAI21_X2 U2741 ( .B1(n2378), .B2(n2377), .A(net84341), .ZN(n2380) );
  OAI21_X2 U2742 ( .B1(n2429), .B2(n2428), .A(opa_00), .ZN(n2431) );
  NAND2_X4 U2743 ( .A1(net85738), .A2(net85748), .ZN(n2035) );
  OAI211_X1 U2744 ( .C1(n2276), .C2(net84561), .A(net11555), .B(n1608), .ZN(
        n2277) );
  NAND3_X2 U2745 ( .A1(fract_out_q[1]), .A2(net85716), .A3(net85732), .ZN(
        n1969) );
  INV_X4 U2746 ( .A(n1969), .ZN(n2049) );
  NAND2_X4 U2747 ( .A1(n2015), .A2(prod[10]), .ZN(net85292) );
  NOR2_X4 U2748 ( .A1(n2031), .A2(net86113), .ZN(net86112) );
  NAND2_X4 U2749 ( .A1(n1921), .A2(net85676), .ZN(net85191) );
  NAND3_X2 U2750 ( .A1(n2034), .A2(quo[0]), .A3(net85684), .ZN(n2050) );
  NAND2_X4 U2751 ( .A1(n2039), .A2(prod[11]), .ZN(n2070) );
  OAI211_X4 U2752 ( .C1(n2031), .C2(net85684), .A(n2030), .B(n2029), .ZN(
        net76048) );
  NAND4_X4 U2753 ( .A1(n2028), .A2(n2027), .A3(n2026), .A4(n2025), .ZN(
        net85285) );
  NAND2_X4 U2754 ( .A1(net85280), .A2(net85281), .ZN(net85331) );
  NAND2_X4 U2755 ( .A1(n2033), .A2(quo[4]), .ZN(n2031) );
  NAND3_X1 U2756 ( .A1(net88319), .A2(n1744), .A3(net90217), .ZN(net85854) );
  NAND2_X4 U2757 ( .A1(n2015), .A2(prod[9]), .ZN(net85263) );
  NAND3_X4 U2758 ( .A1(net85076), .A2(net85674), .A3(quo[18]), .ZN(net85170)
         );
  NAND2_X4 U2759 ( .A1(n1936), .A2(prod[6]), .ZN(net85280) );
  NAND2_X4 U2760 ( .A1(n1973), .A2(net85096), .ZN(n2060) );
  INV_X4 U2761 ( .A(n1972), .ZN(n1973) );
  NAND2_X4 U2762 ( .A1(n1971), .A2(net88566), .ZN(net85124) );
  NAND2_X4 U2763 ( .A1(n2436), .A2(n2435), .ZN(net83875) );
  NAND2_X1 U2764 ( .A1(rmode_r3[1]), .A2(net84403), .ZN(net84402) );
  NAND3_X2 U2765 ( .A1(n2656), .A2(n2619), .A3(net83806), .ZN(n2620) );
  INV_X1 U2766 ( .A(net88319), .ZN(net86010) );
  NAND3_X2 U2767 ( .A1(net85744), .A2(net86006), .A3(prod[16]), .ZN(n2002) );
  XNOR2_X1 U2768 ( .A(net89681), .B(net83421), .ZN(n2467) );
  AOI22_X1 U2769 ( .A1(net85015), .A2(n1949), .B1(net89681), .B2(net84870), 
        .ZN(n2087) );
  AOI22_X4 U2770 ( .A1(net89998), .A2(n1634), .B1(n1955), .B2(prod[17]), .ZN(
        n2036) );
  NAND3_X2 U2771 ( .A1(net85736), .A2(net85746), .A3(prod[8]), .ZN(n2010) );
  NAND3_X2 U2772 ( .A1(net85746), .A2(net85736), .A3(prod[5]), .ZN(net85393)
         );
  INV_X2 U2773 ( .A(n2695), .ZN(n2696) );
  NAND2_X1 U2774 ( .A1(n2695), .A2(n2678), .ZN(n2679) );
  NAND2_X1 U2775 ( .A1(n2695), .A2(n2680), .ZN(n2681) );
  NOR2_X1 U2776 ( .A1(net86037), .A2(n1595), .ZN(n2429) );
  NOR2_X1 U2777 ( .A1(net86037), .A2(net83925), .ZN(n2587) );
  NOR2_X1 U2778 ( .A1(net86037), .A2(n2585), .ZN(n2378) );
  NOR2_X1 U2779 ( .A1(net86037), .A2(net85710), .ZN(net84996) );
  NAND4_X4 U2780 ( .A1(n2028), .A2(n2026), .A3(n2027), .A4(n1923), .ZN(
        net77161) );
  NAND3_X2 U2781 ( .A1(n2036), .A2(n2037), .A3(n2038), .ZN(net85137) );
  NAND2_X1 U2782 ( .A1(net84983), .A2(n1553), .ZN(n2082) );
  XNOR2_X1 U2783 ( .A(n1929), .B(net11560), .ZN(n2464) );
  NAND2_X1 U2784 ( .A1(n2613), .A2(net85842), .ZN(n2694) );
  NAND3_X1 U2785 ( .A1(n2597), .A2(net85842), .A3(n2613), .ZN(n2598) );
  NAND3_X1 U2786 ( .A1(n2425), .A2(net11566), .A3(net85842), .ZN(n2418) );
  XNOR2_X1 U2787 ( .A(net91159), .B(net85710), .ZN(n2484) );
  NAND2_X1 U2788 ( .A1(net91159), .A2(net85710), .ZN(n2400) );
  NOR2_X1 U2789 ( .A1(net89681), .A2(net91159), .ZN(n2364) );
  NOR2_X1 U2790 ( .A1(div_opa_ldz_r2[2]), .A2(net89537), .ZN(n2192) );
  NAND2_X1 U2791 ( .A1(div_opa_ldz_r2[2]), .A2(net89537), .ZN(n2191) );
  AOI22_X4 U2792 ( .A1(net83800), .A2(n2433), .B1(n2683), .B2(n2956), .ZN(
        n2692) );
  NAND3_X1 U2793 ( .A1(net11566), .A2(net85786), .A3(n2327), .ZN(n2543) );
  NAND2_X1 U2794 ( .A1(\u4/exp_in_pl1[5] ), .A2(net85786), .ZN(net84822) );
  NOR3_X1 U2795 ( .A1(net83849), .A2(net83959), .A3(n2566), .ZN(n2567) );
  NOR2_X1 U2796 ( .A1(net83968), .A2(net83959), .ZN(n2553) );
  NAND2_X4 U2797 ( .A1(n2081), .A2(net84468), .ZN(net83945) );
  NAND2_X4 U2798 ( .A1(n2611), .A2(n2612), .ZN(n2695) );
  NAND2_X1 U2799 ( .A1(\u4/exp_next_mi[0] ), .A2(net84157), .ZN(n2367) );
  AOI21_X1 U2800 ( .B1(net86038), .B2(n2698), .A(net85790), .ZN(n2704) );
  NAND4_X1 U2801 ( .A1(net86038), .A2(n1572), .A3(n1595), .A4(n2534), .ZN(
        n2538) );
  NAND2_X4 U2802 ( .A1(net83871), .A2(n2623), .ZN(n2709) );
  NAND2_X1 U2803 ( .A1(net83779), .A2(net86038), .ZN(net84044) );
  NAND4_X1 U2804 ( .A1(n2584), .A2(net83927), .A3(n2583), .A4(net86038), .ZN(
        n2639) );
  NAND3_X1 U2805 ( .A1(n1574), .A2(net86038), .A3(n1615), .ZN(n2605) );
  NAND2_X1 U2806 ( .A1(net86038), .A2(n2579), .ZN(n2187) );
  NAND2_X1 U2807 ( .A1(net86038), .A2(n1571), .ZN(net84675) );
  NAND2_X4 U2808 ( .A1(net88287), .A2(prod[21]), .ZN(net85216) );
  NAND2_X1 U2809 ( .A1(\u4/fract_out_pl1[10] ), .A2(rmode_r3[1]), .ZN(net84480) );
  NAND3_X1 U2810 ( .A1(n1917), .A2(n2082), .A3(net86038), .ZN(n2153) );
  NAND2_X4 U2811 ( .A1(net84096), .A2(net84095), .ZN(net83765) );
  INV_X32 U2812 ( .A(n1980), .ZN(n1978) );
  INV_X4 U2813 ( .A(opb_r[11]), .ZN(n3016) );
  INV_X4 U2814 ( .A(n3112), .ZN(n3014) );
  INV_X4 U2815 ( .A(n3111), .ZN(n3015) );
  NAND4_X2 U2816 ( .A1(n3103), .A2(n3104), .A3(n3101), .A4(n3102), .ZN(n1990)
         );
  INV_X4 U2817 ( .A(n3105), .ZN(n2895) );
  NAND4_X2 U2818 ( .A1(n3109), .A2(n3107), .A3(n3108), .A4(n3106), .ZN(n1989)
         );
  NAND2_X2 U2819 ( .A1(n2959), .A2(n3110), .ZN(n3130) );
  INV_X4 U2820 ( .A(n3114), .ZN(n2889) );
  INV_X4 U2821 ( .A(n3115), .ZN(n2896) );
  NAND2_X2 U2822 ( .A1(n3113), .A2(n3112), .ZN(n1992) );
  NAND2_X2 U2823 ( .A1(n3117), .A2(n3116), .ZN(n1991) );
  NAND2_X2 U2824 ( .A1(n3119), .A2(n3118), .ZN(n1994) );
  INV_X4 U2825 ( .A(n1996), .ZN(N56) );
  INV_X4 U2826 ( .A(N77), .ZN(n2000) );
  NAND2_X2 U2827 ( .A1(n2000), .A2(n3012), .ZN(\u6/N23 ) );
  NOR2_X4 U2828 ( .A1(exp_r[1]), .A2(\u4/div_shft2[0] ), .ZN(net85030) );
  INV_X4 U2829 ( .A(n2002), .ZN(n2004) );
  NOR2_X4 U2830 ( .A1(n2004), .A2(n2003), .ZN(net85171) );
  NAND3_X2 U2831 ( .A1(n2040), .A2(quo[17]), .A3(net85674), .ZN(n2006) );
  OAI21_X4 U2832 ( .B1(n3074), .B2(net88319), .A(n2010), .ZN(net85150) );
  INV_X4 U2833 ( .A(n2011), .ZN(n2013) );
  NOR2_X4 U2834 ( .A1(n2013), .A2(n2012), .ZN(n2028) );
  NOR2_X4 U2835 ( .A1(n3073), .A2(net85716), .ZN(net85336) );
  NAND3_X4 U2836 ( .A1(n1894), .A2(quo[5]), .A3(net85676), .ZN(net85210) );
  NAND3_X4 U2837 ( .A1(n1922), .A2(quo[8]), .A3(net85674), .ZN(net85205) );
  NAND3_X2 U2838 ( .A1(net85076), .A2(net85676), .A3(quo[19]), .ZN(n2037) );
  NAND2_X2 U2839 ( .A1(net85316), .A2(exp_r[2]), .ZN(n2019) );
  INV_X4 U2840 ( .A(exp_r[4]), .ZN(net84290) );
  INV_X4 U2841 ( .A(exp_r[3]), .ZN(net84305) );
  NAND2_X2 U2842 ( .A1(exp_r[3]), .A2(net84290), .ZN(n2404) );
  INV_X4 U2843 ( .A(n2019), .ZN(n2406) );
  MUX2_X2 U2844 ( .A(net84290), .B(n2404), .S(n2406), .Z(n2020) );
  NAND2_X2 U2845 ( .A1(exp_r[4]), .A2(net84305), .ZN(n2405) );
  NAND2_X2 U2846 ( .A1(n2020), .A2(n2405), .ZN(\u4/exp_in_pl1[4] ) );
  XNOR2_X2 U2847 ( .A(net83968), .B(n2406), .ZN(n2442) );
  INV_X4 U2848 ( .A(n2442), .ZN(\u4/exp_in_pl1[3] ) );
  NAND3_X4 U2850 ( .A1(quo[6]), .A2(net85684), .A3(net85076), .ZN(net85067) );
  NAND3_X4 U2851 ( .A1(n2024), .A2(quo[16]), .A3(net85676), .ZN(net85068) );
  NAND3_X4 U2852 ( .A1(net85736), .A2(prod[12]), .A3(net85744), .ZN(n2021) );
  NAND3_X4 U2853 ( .A1(n2023), .A2(n2022), .A3(n2021), .ZN(net85196) );
  NAND3_X4 U2854 ( .A1(net89129), .A2(quo[4]), .A3(net88427), .ZN(net85194) );
  NAND3_X4 U2855 ( .A1(n1942), .A2(quo[14]), .A3(net85676), .ZN(net85195) );
  OAI21_X4 U2856 ( .B1(n3072), .B2(net88319), .A(n2032), .ZN(net85212) );
  NAND3_X4 U2857 ( .A1(n2001), .A2(quo[3]), .A3(net85674), .ZN(net85071) );
  NAND3_X4 U2858 ( .A1(n2016), .A2(quo[6]), .A3(net85674), .ZN(net85041) );
  NAND3_X4 U2859 ( .A1(n2014), .A2(quo[9]), .A3(net85676), .ZN(net85046) );
  NOR3_X4 U2860 ( .A1(net85232), .A2(n2041), .A3(net85196), .ZN(n2044) );
  NAND3_X4 U2861 ( .A1(n2024), .A2(quo[15]), .A3(net85676), .ZN(n2067) );
  OAI21_X4 U2862 ( .B1(n3075), .B2(net88319), .A(n2042), .ZN(n2065) );
  NAND4_X2 U2863 ( .A1(net90144), .A2(net85068), .A3(net85069), .A4(net85067), 
        .ZN(net85140) );
  NOR2_X4 U2864 ( .A1(net85200), .A2(n2048), .ZN(net85182) );
  INV_X4 U2865 ( .A(n2055), .ZN(n2053) );
  INV_X4 U2866 ( .A(net85127), .ZN(net84869) );
  INV_X4 U2867 ( .A(net85124), .ZN(net84531) );
  INV_X4 U2868 ( .A(net85111), .ZN(net84749) );
  NAND2_X2 U2869 ( .A1(net84749), .A2(n2190), .ZN(n2058) );
  XNOR2_X2 U2870 ( .A(n2059), .B(n2058), .ZN(n2448) );
  OAI21_X4 U2871 ( .B1(net89546), .B2(net88618), .A(net84758), .ZN(net85091)
         );
  OAI21_X4 U2872 ( .B1(n1940), .B2(net85093), .A(n2060), .ZN(
        \u4/fi_ldz_mi1[2] ) );
  MUX2_X2 U2873 ( .A(net84290), .B(n2404), .S(net84916), .Z(n2061) );
  NAND2_X2 U2874 ( .A1(prod[0]), .A2(net86125), .ZN(n2064) );
  NAND2_X2 U2875 ( .A1(net89998), .A2(n1660), .ZN(n2062) );
  NAND3_X4 U2876 ( .A1(n2064), .A2(n2063), .A3(n2062), .ZN(n3319) );
  INV_X4 U2877 ( .A(n2069), .ZN(n2072) );
  NOR3_X4 U2878 ( .A1(n2073), .A2(n2072), .A3(n2071), .ZN(n2074) );
  INV_X4 U2879 ( .A(net85039), .ZN(net85037) );
  XNOR2_X2 U2880 ( .A(exp_r[2]), .B(net85030), .ZN(\u4/f2i_shft[2] ) );
  INV_X4 U2881 ( .A(net84822), .ZN(net85027) );
  INV_X4 U2882 ( .A(n2225), .ZN(n2075) );
  NAND3_X4 U2883 ( .A1(net83959), .A2(n2226), .A3(net84236), .ZN(n2099) );
  NAND2_X2 U2884 ( .A1(net84341), .A2(net85847), .ZN(net83951) );
  XNOR2_X2 U2885 ( .A(div_opa_ldz_r2[2]), .B(exp_r[2]), .ZN(n2122) );
  INV_X4 U2886 ( .A(div_opa_ldz_r2[0]), .ZN(net84762) );
  NOR2_X4 U2887 ( .A1(net85832), .A2(net84762), .ZN(n2100) );
  INV_X4 U2888 ( .A(n2103), .ZN(n2076) );
  XNOR2_X2 U2889 ( .A(n2122), .B(n2108), .ZN(n2234) );
  INV_X4 U2890 ( .A(\u4/f2i_shft[2] ), .ZN(n2077) );
  NAND2_X2 U2891 ( .A1(net85006), .A2(net84982), .ZN(net84867) );
  NOR2_X4 U2892 ( .A1(net83421), .A2(n2153), .ZN(n2083) );
  INV_X4 U2893 ( .A(net11671), .ZN(net84992) );
  NAND2_X2 U2894 ( .A1(net83941), .A2(net85710), .ZN(n2089) );
  NAND2_X2 U2895 ( .A1(n2090), .A2(n2089), .ZN(n2092) );
  NOR3_X4 U2896 ( .A1(n2093), .A2(n2092), .A3(n2091), .ZN(n2098) );
  NAND2_X2 U2897 ( .A1(net85710), .A2(net84982), .ZN(n2095) );
  NAND2_X2 U2898 ( .A1(net85832), .A2(net84762), .ZN(n2131) );
  INV_X4 U2899 ( .A(n2100), .ZN(n2101) );
  NAND2_X2 U2900 ( .A1(n2131), .A2(n2101), .ZN(net84600) );
  INV_X4 U2901 ( .A(net84236), .ZN(net83969) );
  INV_X4 U2902 ( .A(n2102), .ZN(n2105) );
  INV_X4 U2903 ( .A(n2131), .ZN(n2104) );
  INV_X4 U2904 ( .A(n2106), .ZN(n2972) );
  INV_X4 U2905 ( .A(n2122), .ZN(n2107) );
  XNOR2_X2 U2906 ( .A(n2972), .B(n2107), .ZN(n2125) );
  INV_X4 U2907 ( .A(n2108), .ZN(n2110) );
  NAND2_X2 U2908 ( .A1(div_opa_ldz_r2[2]), .A2(net11560), .ZN(n2971) );
  INV_X4 U2909 ( .A(n2971), .ZN(n2109) );
  NAND2_X2 U2910 ( .A1(exp_r[2]), .A2(n3096), .ZN(n2970) );
  OAI21_X4 U2911 ( .B1(n2110), .B2(n2109), .A(n2970), .ZN(n2111) );
  INV_X4 U2912 ( .A(n2111), .ZN(n2146) );
  NAND2_X2 U2913 ( .A1(net83968), .A2(n1663), .ZN(n2112) );
  OAI21_X4 U2914 ( .B1(n2146), .B2(n2113), .A(n2112), .ZN(n2148) );
  INV_X4 U2915 ( .A(n2148), .ZN(n2117) );
  INV_X4 U2916 ( .A(n2634), .ZN(n2118) );
  NAND2_X2 U2917 ( .A1(n2118), .A2(net83439), .ZN(n2989) );
  NAND2_X2 U2918 ( .A1(n2634), .A2(net83439), .ZN(net83361) );
  INV_X4 U2919 ( .A(net83361), .ZN(net84886) );
  NAND2_X2 U2920 ( .A1(net84886), .A2(n2119), .ZN(n2124) );
  INV_X4 U2921 ( .A(net83439), .ZN(net83364) );
  NAND2_X2 U2922 ( .A1(div_opa_ldz_r2[0]), .A2(net85832), .ZN(n2132) );
  XNOR2_X2 U2923 ( .A(n2122), .B(n2281), .ZN(n2289) );
  NAND2_X2 U2924 ( .A1(net83364), .A2(n2289), .ZN(n2123) );
  OAI211_X2 U2925 ( .C1(n2125), .C2(n2989), .A(n2124), .B(n2123), .ZN(n2127)
         );
  INV_X4 U2926 ( .A(net84916), .ZN(net84921) );
  NAND2_X2 U2927 ( .A1(net84921), .A2(n2225), .ZN(n2217) );
  INV_X4 U2928 ( .A(n2217), .ZN(n2306) );
  INV_X4 U2929 ( .A(n872), .ZN(net84915) );
  NAND2_X2 U2930 ( .A1(net86169), .A2(net84915), .ZN(n2128) );
  NAND2_X2 U2931 ( .A1(n2129), .A2(n2128), .ZN(\u4/shift_right [2]) );
  XNOR2_X2 U2932 ( .A(net83968), .B(net84916), .ZN(net84858) );
  INV_X4 U2933 ( .A(n2991), .ZN(n2130) );
  NAND2_X2 U2934 ( .A1(n2130), .A2(net85710), .ZN(n2140) );
  INV_X4 U2935 ( .A(net83936), .ZN(net84907) );
  NAND2_X2 U2936 ( .A1(net84906), .A2(net84907), .ZN(net84637) );
  XNOR2_X2 U2937 ( .A(n2133), .B(n2131), .ZN(n2137) );
  XNOR2_X2 U2938 ( .A(n2133), .B(n2132), .ZN(n2290) );
  INV_X4 U2939 ( .A(n2290), .ZN(n2134) );
  NAND2_X2 U2940 ( .A1(net83364), .A2(n2134), .ZN(n2136) );
  INV_X4 U2941 ( .A(net83361), .ZN(net84900) );
  NAND2_X2 U2942 ( .A1(net84900), .A2(net84901), .ZN(n2135) );
  OAI211_X2 U2943 ( .C1(n2989), .C2(n2137), .A(n2136), .B(n2135), .ZN(n2138)
         );
  NAND2_X2 U2944 ( .A1(net85790), .A2(n2138), .ZN(n2141) );
  NAND4_X2 U2945 ( .A1(n2140), .A2(net84637), .A3(n2141), .A4(net84659), .ZN(
        n2143) );
  INV_X4 U2946 ( .A(net89926), .ZN(net84890) );
  INV_X4 U2947 ( .A(n2226), .ZN(n2580) );
  XNOR2_X2 U2948 ( .A(n2146), .B(n1579), .ZN(n2147) );
  INV_X4 U2949 ( .A(n2147), .ZN(n2263) );
  XNOR2_X2 U2950 ( .A(n2288), .B(n2148), .ZN(n2149) );
  INV_X4 U2951 ( .A(n2149), .ZN(n2243) );
  MUX2_X2 U2952 ( .A(n2150), .B(n1663), .S(net83933), .Z(n2151) );
  INV_X4 U2953 ( .A(\u4/exp_in_pl1[4] ), .ZN(n2155) );
  NAND2_X2 U2954 ( .A1(n2442), .A2(n2155), .ZN(n2156) );
  NAND2_X2 U2955 ( .A1(n2157), .A2(n2156), .ZN(net84848) );
  NAND2_X2 U2956 ( .A1(rmode_r3[1]), .A2(rmode_r3[0]), .ZN(n2248) );
  NAND2_X2 U2957 ( .A1(n1614), .A2(n1768), .ZN(net84326) );
  INV_X4 U2958 ( .A(net11558), .ZN(net83968) );
  NAND2_X2 U2959 ( .A1(n2562), .A2(net83968), .ZN(n2303) );
  NOR2_X4 U2960 ( .A1(n2158), .A2(net83963), .ZN(net84048) );
  OAI21_X4 U2961 ( .B1(n2159), .B2(n2248), .A(net84048), .ZN(net83942) );
  INV_X4 U2962 ( .A(net84778), .ZN(net84520) );
  NAND2_X2 U2963 ( .A1(\u4/N406 ), .A2(net84520), .ZN(net84840) );
  INV_X4 U2964 ( .A(\u4/N405 ), .ZN(n2161) );
  OAI21_X4 U2965 ( .B1(net84778), .B2(n2161), .A(n2160), .ZN(\u4/fract_out[5] ) );
  NAND2_X2 U2966 ( .A1(\u4/N402 ), .A2(net84520), .ZN(n2170) );
  INV_X4 U2967 ( .A(\u4/N401 ), .ZN(n2163) );
  NAND2_X2 U2968 ( .A1(\u4/N400 ), .A2(net84520), .ZN(net84810) );
  NOR3_X4 U2969 ( .A1(\u4/N419 ), .A2(\u4/N420 ), .A3(\u4/N418 ), .ZN(n2165)
         );
  NAND2_X2 U2970 ( .A1(net85828), .A2(n2579), .ZN(n2168) );
  NAND2_X2 U2971 ( .A1(net85828), .A2(net11566), .ZN(n2322) );
  NAND2_X2 U2972 ( .A1(\u4/N399 ), .A2(net84520), .ZN(net84564) );
  INV_X4 U2973 ( .A(net84564), .ZN(net84784) );
  NAND3_X2 U2974 ( .A1(n3055), .A2(n3056), .A3(n3054), .ZN(n2178) );
  NAND3_X2 U2975 ( .A1(n3060), .A2(n3061), .A3(n3059), .ZN(n2176) );
  NAND3_X2 U2976 ( .A1(n3063), .A2(n3064), .A3(n3062), .ZN(n2175) );
  NOR4_X2 U2977 ( .A1(n2178), .A2(n2177), .A3(n2176), .A4(n2175), .ZN(n2179)
         );
  NAND2_X2 U2978 ( .A1(n2548), .A2(net85790), .ZN(net83913) );
  INV_X4 U2979 ( .A(net83913), .ZN(net84783) );
  NOR3_X4 U2980 ( .A1(\u4/N423 ), .A2(net84783), .A3(net84784), .ZN(n2186) );
  NOR3_X4 U2981 ( .A1(\u4/N390 ), .A2(\u4/N392 ), .A3(\u4/N388 ), .ZN(n2184)
         );
  NOR4_X2 U2982 ( .A1(\u4/N394 ), .A2(\u4/N395 ), .A3(\u4/N389 ), .A4(
        \u4/N391 ), .ZN(n2183) );
  NOR4_X2 U2983 ( .A1(\u4/N398 ), .A2(\u4/N396 ), .A3(\u4/N393 ), .A4(
        \u4/N397 ), .ZN(n2182) );
  INV_X4 U2984 ( .A(n2301), .ZN(n2185) );
  NAND2_X2 U2985 ( .A1(n1640), .A2(n1589), .ZN(net84643) );
  MUX2_X2 U2986 ( .A(\u4/exp_in_pl1[4] ), .B(\u4/exp_next_mi[4] ), .S(net85788), .Z(net84764) );
  NAND2_X2 U2987 ( .A1(rmode_r3[1]), .A2(net86016), .ZN(net84490) );
  INV_X4 U2988 ( .A(net83402), .ZN(net84633) );
  INV_X4 U2989 ( .A(\u4/exp_next_mi[3] ), .ZN(net84768) );
  MUX2_X2 U2990 ( .A(n2442), .B(net84768), .S(net85788), .Z(net84445) );
  MUX2_X2 U2991 ( .A(net85712), .B(net89692), .S(net85788), .Z(net84767) );
  INV_X4 U2992 ( .A(net84767), .ZN(net84766) );
  XOR2_X2 U2993 ( .A(net84764), .B(net84765), .Z(n2231) );
  NOR2_X4 U2994 ( .A1(n2189), .A2(n2188), .ZN(n2260) );
  XNOR2_X2 U2995 ( .A(n2443), .B(div_opa_ldz_r2[3]), .ZN(n2193) );
  XNOR2_X2 U2996 ( .A(n2193), .B(n2196), .ZN(n2551) );
  NAND2_X2 U2997 ( .A1(\u4/exp_in_pl1[3] ), .A2(n2551), .ZN(n2194) );
  INV_X4 U2998 ( .A(n2443), .ZN(n2401) );
  NOR2_X4 U2999 ( .A1(div_opa_ldz_r2[3]), .A2(n2401), .ZN(n2198) );
  NAND2_X2 U3000 ( .A1(n2401), .A2(div_opa_ldz_r2[3]), .ZN(n2197) );
  OAI21_X4 U3001 ( .B1(n2199), .B2(n2198), .A(n2197), .ZN(n2549) );
  XNOR2_X2 U3002 ( .A(n2549), .B(n2200), .ZN(n2552) );
  XNOR2_X2 U3003 ( .A(n2552), .B(\u4/exp_in_pl1[4] ), .ZN(n2201) );
  XNOR2_X2 U3004 ( .A(n2202), .B(n2201), .ZN(n2229) );
  INV_X4 U3005 ( .A(net11560), .ZN(net83994) );
  INV_X4 U3006 ( .A(net11564), .ZN(net83967) );
  NAND2_X2 U3007 ( .A1(n3096), .A2(net83994), .ZN(n2206) );
  NAND2_X2 U3008 ( .A1(net11671), .A2(net83993), .ZN(n2205) );
  OAI211_X2 U3009 ( .C1(n2208), .C2(n2207), .A(n2206), .B(n2205), .ZN(n2211)
         );
  INV_X4 U3010 ( .A(n1663), .ZN(n2209) );
  AOI21_X2 U3011 ( .B1(n2212), .B2(n2211), .A(n2210), .ZN(n2214) );
  XNOR2_X2 U3012 ( .A(n2222), .B(n2443), .ZN(n2422) );
  XNOR2_X2 U3013 ( .A(n2225), .B(net84305), .ZN(n2992) );
  NAND2_X2 U3014 ( .A1(n2422), .A2(n2992), .ZN(n2221) );
  NAND2_X2 U3015 ( .A1(net89964), .A2(net85710), .ZN(n2215) );
  NOR2_X4 U3016 ( .A1(n2422), .A2(n2992), .ZN(n2220) );
  XNOR2_X2 U3017 ( .A(n2224), .B(n2242), .ZN(n2228) );
  NAND2_X2 U3018 ( .A1(n2227), .A2(n2226), .ZN(n2981) );
  XNOR2_X2 U3019 ( .A(n2228), .B(n2981), .ZN(n2311) );
  OAI22_X2 U3020 ( .A1(n2229), .A2(net84611), .B1(n2311), .B2(net88427), .ZN(
        n2230) );
  AOI21_X2 U3021 ( .B1(net84633), .B2(n2231), .A(n2230), .ZN(n2247) );
  INV_X4 U3022 ( .A(n2965), .ZN(n2237) );
  INV_X4 U3023 ( .A(n2234), .ZN(n2964) );
  NOR2_X4 U3024 ( .A1(net83407), .A2(n2964), .ZN(n2236) );
  NAND2_X2 U3025 ( .A1(n2964), .A2(net83407), .ZN(n2235) );
  OAI21_X4 U3026 ( .B1(n2237), .B2(n2236), .A(n2235), .ZN(n2264) );
  INV_X4 U3027 ( .A(n2264), .ZN(n2241) );
  INV_X4 U3028 ( .A(n2422), .ZN(n2238) );
  NAND2_X2 U3029 ( .A1(n2263), .A2(n2238), .ZN(n2239) );
  INV_X4 U3030 ( .A(n2242), .ZN(n2421) );
  XNOR2_X2 U3031 ( .A(n2243), .B(n2421), .ZN(n2244) );
  XNOR2_X2 U3032 ( .A(n2245), .B(n2244), .ZN(n2246) );
  INV_X4 U3033 ( .A(net84669), .ZN(net84619) );
  MUX2_X2 U3034 ( .A(n2247), .B(n2246), .S(net84619), .Z(net83995) );
  INV_X4 U3035 ( .A(n2248), .ZN(n2249) );
  NAND4_X2 U3036 ( .A1(n2249), .A2(opas_r2), .A3(net83936), .A4(net84048), 
        .ZN(net84488) );
  NAND2_X2 U3037 ( .A1(n2401), .A2(n2253), .ZN(net84639) );
  XNOR2_X2 U3038 ( .A(n2251), .B(n2250), .ZN(n2307) );
  INV_X4 U3039 ( .A(net84659), .ZN(net84656) );
  INV_X4 U3040 ( .A(net84652), .ZN(net83934) );
  INV_X4 U3041 ( .A(net83429), .ZN(net84647) );
  NAND2_X2 U3042 ( .A1(net84647), .A2(net84490), .ZN(net84449) );
  INV_X4 U3043 ( .A(n2962), .ZN(n2252) );
  NAND3_X4 U3044 ( .A1(net84644), .A2(net84645), .A3(n2252), .ZN(n2358) );
  INV_X4 U3045 ( .A(net84642), .ZN(net84632) );
  NAND2_X2 U3046 ( .A1(n2254), .A2(n2443), .ZN(n2255) );
  INV_X4 U3047 ( .A(net84637), .ZN(net83423) );
  NAND2_X2 U3048 ( .A1(net84632), .A2(net84633), .ZN(net84624) );
  XNOR2_X2 U3049 ( .A(n2551), .B(n2442), .ZN(n2259) );
  XNOR2_X2 U3050 ( .A(n2260), .B(n2259), .ZN(net84629) );
  XNOR2_X2 U3051 ( .A(n2422), .B(n2992), .ZN(n2262) );
  XNOR2_X2 U3052 ( .A(n2262), .B(n2261), .ZN(n2309) );
  XNOR2_X2 U3053 ( .A(n2263), .B(n2422), .ZN(n2265) );
  XNOR2_X2 U3054 ( .A(n2265), .B(n2264), .ZN(n2266) );
  NAND2_X2 U3055 ( .A1(n2267), .A2(net84614), .ZN(n2331) );
  OAI21_X4 U3056 ( .B1(n2268), .B2(n2331), .A(net83429), .ZN(n2357) );
  NAND2_X2 U3057 ( .A1(net84160), .A2(net84166), .ZN(n2366) );
  INV_X4 U3058 ( .A(net84605), .ZN(net84604) );
  INV_X4 U3059 ( .A(net84600), .ZN(net83438) );
  NAND2_X2 U3060 ( .A1(\u4/exp_f2i_1 [23]), .A2(n1606), .ZN(n2271) );
  INV_X4 U3061 ( .A(n2271), .ZN(n2272) );
  NOR4_X2 U3062 ( .A1(n2274), .A2(n2273), .A3(net84595), .A4(n2272), .ZN(
        net84474) );
  NAND2_X2 U3063 ( .A1(net84591), .A2(n1589), .ZN(net84579) );
  NAND2_X2 U3064 ( .A1(net84590), .A2(net83429), .ZN(net84475) );
  NAND2_X2 U3065 ( .A1(n2275), .A2(net84564), .ZN(n2546) );
  INV_X4 U3066 ( .A(n2546), .ZN(n2278) );
  NAND2_X2 U3067 ( .A1(n2278), .A2(n2277), .ZN(n2280) );
  OAI21_X4 U3068 ( .B1(net84555), .B2(n2280), .A(n2279), .ZN(net84403) );
  NAND2_X2 U3069 ( .A1(sign), .A2(net84403), .ZN(net84482) );
  INV_X4 U3070 ( .A(net84550), .ZN(net84548) );
  NAND2_X2 U3071 ( .A1(net83968), .A2(div_opa_ldz_r2[3]), .ZN(n2286) );
  INV_X4 U3072 ( .A(n2281), .ZN(n2284) );
  NAND2_X2 U3073 ( .A1(exp_r[2]), .A2(div_opa_ldz_r2[2]), .ZN(n2282) );
  NAND2_X2 U3074 ( .A1(n2286), .A2(n2285), .ZN(n2287) );
  XNOR2_X2 U3075 ( .A(n2288), .B(n2287), .ZN(n2978) );
  INV_X4 U3076 ( .A(n2978), .ZN(n2297) );
  INV_X4 U3077 ( .A(n2289), .ZN(n2291) );
  NAND2_X2 U3078 ( .A1(n2291), .A2(n2290), .ZN(n2294) );
  INV_X4 U3079 ( .A(n2292), .ZN(n2293) );
  XNOR2_X2 U3080 ( .A(n1579), .B(n2293), .ZN(n2987) );
  NAND2_X2 U3081 ( .A1(n2294), .A2(n2987), .ZN(n2296) );
  NAND2_X2 U3082 ( .A1(net84531), .A2(net84532), .ZN(n2295) );
  NAND2_X2 U3083 ( .A1(net84520), .A2(n2301), .ZN(n2545) );
  NAND2_X2 U3084 ( .A1(net83950), .A2(n2302), .ZN(net84327) );
  INV_X4 U3085 ( .A(net84327), .ZN(net84334) );
  INV_X4 U3086 ( .A(n2322), .ZN(n2305) );
  INV_X4 U3087 ( .A(n2303), .ZN(n2304) );
  NAND3_X2 U3088 ( .A1(n2309), .A2(n2366), .A3(n2308), .ZN(n2310) );
  NAND3_X4 U3089 ( .A1(n2311), .A2(n2310), .A3(net84506), .ZN(n2420) );
  INV_X4 U3090 ( .A(net84469), .ZN(net84501) );
  INV_X4 U3091 ( .A(net83927), .ZN(net84498) );
  OAI21_X4 U3092 ( .B1(n2312), .B2(n2420), .A(net84500), .ZN(n2316) );
  NAND2_X2 U3093 ( .A1(net84498), .A2(net85794), .ZN(n2314) );
  INV_X4 U3094 ( .A(net83844), .ZN(net84465) );
  INV_X4 U3095 ( .A(n2420), .ZN(n2317) );
  OAI21_X4 U3096 ( .B1(n2319), .B2(net84490), .A(n2318), .ZN(net84332) );
  INV_X4 U3097 ( .A(net84332), .ZN(net83855) );
  INV_X4 U3098 ( .A(net84488), .ZN(net84487) );
  NAND2_X2 U3099 ( .A1(net84487), .A2(net83941), .ZN(n2600) );
  NAND3_X4 U3100 ( .A1(net83855), .A2(n2600), .A3(n2320), .ZN(net84220) );
  NAND2_X2 U3101 ( .A1(n1603), .A2(net84211), .ZN(n2474) );
  NOR2_X4 U3102 ( .A1(net83296), .A2(net84150), .ZN(n2339) );
  INV_X4 U3103 ( .A(net84312), .ZN(net84366) );
  NAND2_X2 U3104 ( .A1(n2437), .A2(n2420), .ZN(n2424) );
  NAND2_X2 U3105 ( .A1(rmode_r3[0]), .A2(n1768), .ZN(n2588) );
  INV_X4 U3106 ( .A(n2588), .ZN(n2425) );
  NAND2_X2 U3107 ( .A1(n2425), .A2(n1597), .ZN(n2326) );
  NOR2_X4 U3108 ( .A1(n2420), .A2(n2588), .ZN(n2415) );
  OAI21_X4 U3109 ( .B1(net85828), .B2(net83927), .A(n2420), .ZN(n2327) );
  INV_X4 U3110 ( .A(n2543), .ZN(n2328) );
  AOI211_X4 U3111 ( .C1(net83969), .C2(n2424), .A(n2329), .B(n2328), .ZN(n2458) );
  INV_X4 U3112 ( .A(n2329), .ZN(n2330) );
  NAND2_X2 U3113 ( .A1(sign), .A2(rmode_r3[1]), .ZN(n2416) );
  NAND2_X2 U3114 ( .A1(net84080), .A2(net85794), .ZN(n2340) );
  NOR2_X4 U3115 ( .A1(n2458), .A2(n2521), .ZN(n2335) );
  NAND2_X2 U3116 ( .A1(net84343), .A2(net84398), .ZN(n2494) );
  NAND2_X2 U3117 ( .A1(net84450), .A2(net85847), .ZN(net84134) );
  INV_X4 U3118 ( .A(net84134), .ZN(net84368) );
  INV_X4 U3119 ( .A(n2331), .ZN(n2332) );
  OAI21_X4 U3120 ( .B1(net84445), .B2(net83432), .A(n2332), .ZN(net84148) );
  NAND2_X2 U3121 ( .A1(net84368), .A2(net84148), .ZN(n2388) );
  NAND3_X4 U3122 ( .A1(n2490), .A2(n2494), .A3(n2338), .ZN(n2454) );
  INV_X4 U3123 ( .A(n2333), .ZN(n2334) );
  NAND2_X2 U3124 ( .A1(net84133), .A2(n2388), .ZN(n2338) );
  NAND4_X2 U3125 ( .A1(n1648), .A2(n2496), .A3(n1588), .A4(n2491), .ZN(n2346)
         );
  INV_X4 U3126 ( .A(n2340), .ZN(n2343) );
  INV_X4 U3127 ( .A(n2341), .ZN(n2342) );
  NOR2_X4 U3128 ( .A1(n2348), .A2(n2347), .ZN(n2612) );
  NAND3_X4 U3129 ( .A1(n1603), .A2(n2996), .A3(net84211), .ZN(net84218) );
  NAND2_X2 U3130 ( .A1(net84081), .A2(net84218), .ZN(n2349) );
  INV_X4 U3131 ( .A(n2437), .ZN(n2426) );
  XNOR2_X2 U3132 ( .A(n2996), .B(n2426), .ZN(n2351) );
  NAND2_X2 U3133 ( .A1(n2353), .A2(n2352), .ZN(net84333) );
  NAND2_X2 U3134 ( .A1(n2358), .A2(n2357), .ZN(n2360) );
  NOR3_X4 U3135 ( .A1(n2361), .A2(n2437), .A3(n1597), .ZN(net84374) );
  INV_X4 U3136 ( .A(n2419), .ZN(n2462) );
  INV_X4 U3137 ( .A(n2461), .ZN(n2363) );
  INV_X4 U3138 ( .A(n2566), .ZN(n2555) );
  INV_X4 U3139 ( .A(n2366), .ZN(n2368) );
  AOI211_X4 U3140 ( .C1(n2370), .C2(n2371), .A(net84352), .B(n2369), .ZN(n2436) );
  INV_X4 U3141 ( .A(n2375), .ZN(n2611) );
  NAND2_X2 U3142 ( .A1(n2611), .A2(n2612), .ZN(net84344) );
  INV_X4 U3143 ( .A(net84344), .ZN(net83754) );
  NAND2_X2 U3144 ( .A1(n3065), .A2(n3071), .ZN(n2698) );
  NAND2_X2 U3145 ( .A1(net84343), .A2(n2698), .ZN(n2585) );
  NAND2_X2 U3146 ( .A1(n1640), .A2(n1576), .ZN(n2379) );
  NAND2_X2 U3147 ( .A1(n2380), .A2(n2379), .ZN(n2683) );
  OAI21_X4 U3148 ( .B1(net84334), .B2(net84326), .A(n2588), .ZN(n2381) );
  OAI21_X4 U3149 ( .B1(n2382), .B2(n2381), .A(net84095), .ZN(n2514) );
  OAI21_X4 U3150 ( .B1(n2385), .B2(n2384), .A(net84095), .ZN(n2513) );
  INV_X4 U3151 ( .A(\u4/fract_out_pl1[0] ), .ZN(n2386) );
  INV_X4 U3152 ( .A(n2416), .ZN(n2387) );
  NOR2_X4 U3153 ( .A1(n2389), .A2(n2388), .ZN(n2391) );
  INV_X4 U3154 ( .A(n2600), .ZN(n2390) );
  AOI211_X4 U3155 ( .C1(n2392), .C2(n2391), .A(net83878), .B(n2390), .ZN(
        net84253) );
  INV_X4 U3156 ( .A(net84315), .ZN(net84314) );
  OAI21_X4 U3157 ( .B1(n2465), .B2(n2396), .A(n2395), .ZN(n2449) );
  XNOR2_X2 U3158 ( .A(exp_r[4]), .B(n2399), .ZN(n2414) );
  NAND2_X2 U3159 ( .A1(\u4/exp_in_pl1[3] ), .A2(n2401), .ZN(n2403) );
  INV_X4 U3160 ( .A(n2404), .ZN(n2409) );
  INV_X4 U3161 ( .A(n2405), .ZN(n2407) );
  MUX2_X2 U3162 ( .A(n2407), .B(net84290), .S(n2406), .Z(n2408) );
  XNOR2_X2 U3163 ( .A(n2412), .B(n2411), .ZN(n2413) );
  OAI22_X2 U3164 ( .A1(n2414), .A2(n2482), .B1(n2413), .B2(n2486), .ZN(
        net84076) );
  INV_X4 U3165 ( .A(net84076), .ZN(net84280) );
  NOR2_X4 U3166 ( .A1(net84276), .A2(net84277), .ZN(net84200) );
  INV_X4 U3167 ( .A(n2415), .ZN(n2417) );
  NAND2_X2 U3168 ( .A1(n1583), .A2(n2419), .ZN(net84266) );
  NAND2_X2 U3169 ( .A1(net84265), .A2(net84266), .ZN(net83864) );
  INV_X4 U3170 ( .A(net83864), .ZN(net83876) );
  INV_X4 U3171 ( .A(n2420), .ZN(n2438) );
  INV_X4 U3172 ( .A(n2423), .ZN(n2439) );
  OAI211_X2 U3173 ( .C1(n2438), .C2(n2439), .A(n2424), .B(net83969), .ZN(n2427) );
  OAI21_X4 U3174 ( .B1(n2438), .B2(n2426), .A(n2425), .ZN(n2542) );
  NAND3_X2 U3175 ( .A1(n2427), .A2(n2542), .A3(n2543), .ZN(n2622) );
  NAND2_X2 U3176 ( .A1(net83876), .A2(n2622), .ZN(net84254) );
  INV_X4 U3177 ( .A(n2683), .ZN(n2433) );
  NAND2_X2 U3178 ( .A1(opa_inf), .A2(n1613), .ZN(n2432) );
  INV_X4 U3179 ( .A(net83781), .ZN(net84249) );
  NAND3_X2 U3180 ( .A1(n2432), .A2(n2431), .A3(n2430), .ZN(n2956) );
  AOI21_X4 U3181 ( .B1(n2439), .B2(n2426), .A(n2438), .ZN(n2440) );
  NOR2_X4 U3182 ( .A1(n2440), .A2(net84236), .ZN(n2541) );
  NAND2_X2 U3183 ( .A1(n2543), .A2(n2542), .ZN(n2441) );
  INV_X4 U3184 ( .A(n2486), .ZN(n2447) );
  XNOR2_X2 U3185 ( .A(n2443), .B(n2442), .ZN(n2445) );
  XNOR2_X2 U3186 ( .A(n2445), .B(n2444), .ZN(n2446) );
  NAND2_X2 U3187 ( .A1(n2447), .A2(n2446), .ZN(net84215) );
  INV_X4 U3188 ( .A(n2482), .ZN(n2452) );
  XNOR2_X2 U3189 ( .A(n2450), .B(n2449), .ZN(n2451) );
  NAND2_X2 U3190 ( .A1(n2452), .A2(n2451), .ZN(net84216) );
  INV_X4 U3191 ( .A(n2454), .ZN(n2477) );
  NAND3_X2 U3192 ( .A1(n2455), .A2(n2496), .A3(n2477), .ZN(n2456) );
  NAND2_X2 U3193 ( .A1(n2463), .A2(n2462), .ZN(n2475) );
  XNOR2_X2 U3194 ( .A(n2465), .B(n2464), .ZN(n2466) );
  XNOR2_X2 U3195 ( .A(n2468), .B(n2467), .ZN(n2469) );
  NAND4_X2 U3196 ( .A1(n2475), .A2(n2474), .A3(net84081), .A4(n2473), .ZN(
        n2476) );
  INV_X4 U3197 ( .A(n2476), .ZN(n2524) );
  NAND2_X2 U3198 ( .A1(n2480), .A2(n2479), .ZN(n2526) );
  INV_X4 U3199 ( .A(net84166), .ZN(net84165) );
  XNOR2_X2 U3200 ( .A(n2481), .B(net84165), .ZN(n2483) );
  INV_X4 U3201 ( .A(net84160), .ZN(net84159) );
  XNOR2_X2 U3202 ( .A(n2484), .B(net84159), .ZN(n2487) );
  NAND2_X2 U3203 ( .A1(net89692), .A2(net84157), .ZN(n2485) );
  INV_X4 U3204 ( .A(net84148), .ZN(net84146) );
  NAND2_X2 U3205 ( .A1(net84146), .A2(net84133), .ZN(n2492) );
  NAND4_X2 U3206 ( .A1(n2493), .A2(n2492), .A3(n2491), .A4(n2490), .ZN(n2501)
         );
  NAND4_X2 U3207 ( .A1(n2497), .A2(n2496), .A3(n2495), .A4(n2494), .ZN(n2500)
         );
  INV_X4 U3208 ( .A(\u4/fract_out_pl1[7] ), .ZN(n2504) );
  OAI22_X2 U3209 ( .A1(n1928), .A2(n2504), .B1(n2503), .B2(n1961), .ZN(n2687)
         );
  INV_X4 U3210 ( .A(\u4/fract_out_pl1[8] ), .ZN(n2505) );
  OAI22_X2 U3211 ( .A1(net84119), .A2(n1961), .B1(n2513), .B2(n2505), .ZN(
        n2689) );
  INV_X4 U3212 ( .A(\u4/fract_out_pl1[9] ), .ZN(n2506) );
  NOR3_X4 U3213 ( .A1(n2687), .A2(n2689), .A3(n2691), .ZN(n2519) );
  INV_X4 U3214 ( .A(\u4/fract_out_pl1[5] ), .ZN(n2507) );
  OAI22_X2 U3215 ( .A1(net84115), .A2(n1961), .B1(n2513), .B2(n2507), .ZN(
        n2682) );
  INV_X4 U3216 ( .A(\u4/fract_out_pl1[6] ), .ZN(n2508) );
  NOR2_X4 U3217 ( .A1(n2682), .A2(n2685), .ZN(n2518) );
  INV_X4 U3218 ( .A(\u4/fract_out_pl1[2] ), .ZN(n2509) );
  INV_X4 U3219 ( .A(\u4/fract_out_pl1[3] ), .ZN(n2510) );
  INV_X4 U3220 ( .A(\u4/fract_out_pl1[4] ), .ZN(n2511) );
  INV_X4 U3221 ( .A(\u4/fract_out_pl1[1] ), .ZN(n2512) );
  NAND2_X2 U3222 ( .A1(net84095), .A2(net84096), .ZN(net84024) );
  NOR2_X4 U3223 ( .A1(n2522), .A2(n2521), .ZN(n2525) );
  OAI21_X4 U3224 ( .B1(n2525), .B2(net84059), .A(net83861), .ZN(n2706) );
  NAND3_X2 U3225 ( .A1(net83747), .A2(net84024), .A3(n2706), .ZN(n2529) );
  OAI21_X4 U3226 ( .B1(n2528), .B2(net84060), .A(net83861), .ZN(net83736) );
  INV_X4 U3227 ( .A(\u4/exp_next_mi[4] ), .ZN(n2530) );
  OAI211_X2 U3228 ( .C1(n2530), .C2(net84079), .A(net84080), .B(net84081), 
        .ZN(n2531) );
  NAND2_X2 U3229 ( .A1(opa_00), .A2(opb_00), .ZN(net84021) );
  NAND2_X2 U3230 ( .A1(opa_00), .A2(opb_inf), .ZN(n2533) );
  NAND2_X2 U3231 ( .A1(opa_inf), .A2(opb_00), .ZN(n2532) );
  NAND2_X2 U3232 ( .A1(n2533), .A2(n2532), .ZN(net83925) );
  NAND3_X2 U3233 ( .A1(n1561), .A2(n1570), .A3(n1595), .ZN(n2536) );
  INV_X4 U3234 ( .A(n2541), .ZN(n2544) );
  NAND3_X2 U3235 ( .A1(n2544), .A2(n2543), .A3(n2542), .ZN(net84003) );
  INV_X4 U3236 ( .A(n2545), .ZN(n2573) );
  NAND2_X2 U3237 ( .A1(n2547), .A2(net88950), .ZN(n2583) );
  INV_X4 U3238 ( .A(n2583), .ZN(n2572) );
  INV_X4 U3239 ( .A(n2548), .ZN(n2570) );
  INV_X4 U3240 ( .A(net83995), .ZN(net83973) );
  INV_X4 U3241 ( .A(n2549), .ZN(n2550) );
  INV_X4 U3242 ( .A(n2552), .ZN(n2554) );
  NAND2_X2 U3243 ( .A1(n2555), .A2(net83364), .ZN(n2558) );
  OAI21_X4 U3244 ( .B1(n2557), .B2(n2556), .A(n2558), .ZN(n2559) );
  INV_X4 U3245 ( .A(n2558), .ZN(n2565) );
  AOI21_X4 U3246 ( .B1(n2560), .B2(n2559), .A(n1646), .ZN(net83975) );
  MUX2_X2 U3247 ( .A(net83971), .B(net83972), .S(net11555), .Z(n2561) );
  INV_X4 U3248 ( .A(n2563), .ZN(n2564) );
  OAI21_X4 U3249 ( .B1(n2570), .B2(n2569), .A(n2568), .ZN(n2630) );
  NAND2_X2 U3250 ( .A1(net85828), .A2(n2630), .ZN(n2571) );
  NAND2_X2 U3251 ( .A1(n2629), .A2(net85790), .ZN(n2578) );
  NAND2_X2 U3252 ( .A1(n2583), .A2(net83951), .ZN(n2599) );
  INV_X4 U3253 ( .A(net83942), .ZN(net83940) );
  INV_X4 U3254 ( .A(n2601), .ZN(n2576) );
  NOR2_X4 U3255 ( .A1(n1605), .A2(n2576), .ZN(n2577) );
  NAND4_X2 U3256 ( .A1(net83906), .A2(n2578), .A3(n2599), .A4(n2577), .ZN(
        n2595) );
  NAND2_X2 U3257 ( .A1(net90047), .A2(net11566), .ZN(n2632) );
  NAND2_X2 U3258 ( .A1(n2582), .A2(n2581), .ZN(n2584) );
  NAND2_X2 U3259 ( .A1(net83836), .A2(n2639), .ZN(n2594) );
  NAND3_X2 U3260 ( .A1(n2585), .A2(n1572), .A3(n1595), .ZN(n2586) );
  NAND2_X2 U3261 ( .A1(n2587), .A2(n2586), .ZN(n2662) );
  INV_X4 U3262 ( .A(n2662), .ZN(n2591) );
  INV_X4 U3263 ( .A(n2698), .ZN(n2589) );
  INV_X4 U3264 ( .A(n2605), .ZN(n2619) );
  NAND3_X2 U3265 ( .A1(n2592), .A2(n2600), .A3(net83913), .ZN(n2593) );
  INV_X4 U3266 ( .A(n2599), .ZN(n2603) );
  NAND2_X2 U3267 ( .A1(n2601), .A2(n2600), .ZN(n2602) );
  NAND2_X2 U3268 ( .A1(net83747), .A2(net91075), .ZN(n2699) );
  NAND2_X2 U3269 ( .A1(n1574), .A2(net85790), .ZN(n2604) );
  AND3_X2 U3270 ( .A1(n2605), .A2(n2699), .A3(n2604), .ZN(n2606) );
  INV_X4 U3271 ( .A(n2614), .ZN(n2608) );
  NAND2_X2 U3272 ( .A1(n2614), .A2(net85794), .ZN(n2615) );
  INV_X4 U3273 ( .A(net83883), .ZN(net83806) );
  AOI21_X2 U3274 ( .B1(net83876), .B2(n2622), .A(net83878), .ZN(net83874) );
  NOR2_X4 U3275 ( .A1(net83869), .A2(net83864), .ZN(n2624) );
  OAI21_X4 U3276 ( .B1(n2624), .B2(net83868), .A(net83861), .ZN(n2707) );
  NAND2_X2 U3277 ( .A1(underflow_fmul_r[2]), .A2(n1550), .ZN(net83821) );
  NOR3_X4 U3278 ( .A1(net83856), .A2(n2665), .A3(net83821), .ZN(n2646) );
  NAND2_X2 U3279 ( .A1(net83855), .A2(net85790), .ZN(n2628) );
  INV_X4 U3280 ( .A(n2629), .ZN(n2638) );
  INV_X4 U3281 ( .A(n2630), .ZN(n2631) );
  MUX2_X2 U3282 ( .A(net83849), .B(n2631), .S(net85828), .Z(n2635) );
  NAND3_X2 U3283 ( .A1(n2635), .A2(n2634), .A3(n2633), .ZN(n2636) );
  NAND2_X2 U3284 ( .A1(n2636), .A2(net83844), .ZN(n2637) );
  NOR2_X4 U3285 ( .A1(n2638), .A2(n2637), .ZN(n2641) );
  INV_X4 U3286 ( .A(n2639), .ZN(n2640) );
  AOI21_X4 U3287 ( .B1(n2642), .B2(n2641), .A(n2640), .ZN(n2644) );
  INV_X4 U3288 ( .A(net83836), .ZN(net83833) );
  NOR2_X4 U3289 ( .A1(net83833), .A2(n1651), .ZN(n2643) );
  INV_X4 U3290 ( .A(net83821), .ZN(net83820) );
  NAND2_X2 U3291 ( .A1(n2649), .A2(n2648), .ZN(net83811) );
  INV_X4 U3292 ( .A(n3170), .ZN(n2650) );
  NAND4_X2 U3293 ( .A1(n3172), .A2(n3171), .A3(n2652), .A4(n2651), .ZN(
        net83812) );
  INV_X4 U3294 ( .A(n2653), .ZN(n2654) );
  NOR3_X2 U3295 ( .A1(net83807), .A2(net86016), .A3(n2654), .ZN(n2655) );
  INV_X4 U3296 ( .A(n2669), .ZN(n2667) );
  NAND4_X2 U3297 ( .A1(net83779), .A2(net91075), .A3(net83781), .A4(n1576), 
        .ZN(n2671) );
  NAND2_X2 U3298 ( .A1(n2433), .A2(n2685), .ZN(n2686) );
  NAND2_X2 U3299 ( .A1(n2433), .A2(n2687), .ZN(n2688) );
  NAND2_X2 U3300 ( .A1(n2433), .A2(n2691), .ZN(n2693) );
  INV_X4 U3301 ( .A(n2694), .ZN(n2697) );
  NOR2_X4 U3302 ( .A1(n2697), .A2(n2696), .ZN(n2705) );
  NAND2_X2 U3303 ( .A1(net83736), .A2(n2433), .ZN(N231) );
  NAND2_X2 U3304 ( .A1(n2708), .A2(n2433), .ZN(N233) );
  INV_X4 U3305 ( .A(N76), .ZN(n2710) );
  MUX2_X2 U3306 ( .A(n3120), .B(n2710), .S(n3012), .Z(n2711) );
  INV_X4 U3307 ( .A(n2711), .ZN(\u6/N22 ) );
  INV_X4 U3308 ( .A(N75), .ZN(n2712) );
  MUX2_X2 U3309 ( .A(n3119), .B(n2712), .S(n3012), .Z(n2713) );
  INV_X4 U3310 ( .A(n2713), .ZN(\u6/N21 ) );
  INV_X4 U3311 ( .A(N74), .ZN(n2714) );
  MUX2_X2 U3312 ( .A(n3118), .B(n2714), .S(n3012), .Z(n2715) );
  INV_X4 U3313 ( .A(n2715), .ZN(\u6/N20 ) );
  INV_X4 U3314 ( .A(N73), .ZN(n2716) );
  MUX2_X2 U3315 ( .A(n3117), .B(n2716), .S(n3012), .Z(n2717) );
  INV_X4 U3316 ( .A(n2717), .ZN(\u6/N19 ) );
  INV_X4 U3317 ( .A(N72), .ZN(n2718) );
  MUX2_X2 U3318 ( .A(n3116), .B(n2718), .S(n3012), .Z(n2719) );
  INV_X4 U3319 ( .A(n2719), .ZN(\u6/N18 ) );
  INV_X4 U3320 ( .A(N71), .ZN(n2720) );
  MUX2_X2 U3321 ( .A(n3115), .B(n2720), .S(n3012), .Z(n2721) );
  INV_X4 U3322 ( .A(n2721), .ZN(\u6/N17 ) );
  INV_X4 U3323 ( .A(N70), .ZN(n2722) );
  MUX2_X2 U3324 ( .A(n3114), .B(n2722), .S(n3012), .Z(n2723) );
  INV_X4 U3325 ( .A(n2723), .ZN(\u6/N16 ) );
  INV_X4 U3326 ( .A(N69), .ZN(n2724) );
  MUX2_X2 U3327 ( .A(n3113), .B(n2724), .S(n3012), .Z(n2725) );
  INV_X4 U3328 ( .A(n2725), .ZN(\u6/N15 ) );
  INV_X4 U3329 ( .A(N68), .ZN(n2726) );
  MUX2_X2 U3330 ( .A(n3112), .B(n2726), .S(n3012), .Z(n2727) );
  INV_X4 U3331 ( .A(n2727), .ZN(\u6/N14 ) );
  INV_X4 U3332 ( .A(N67), .ZN(n2728) );
  MUX2_X2 U3333 ( .A(n3111), .B(n2728), .S(n3012), .Z(n2729) );
  INV_X4 U3334 ( .A(n2729), .ZN(\u6/N13 ) );
  INV_X4 U3335 ( .A(n2833), .ZN(n2767) );
  NAND2_X2 U3336 ( .A1(n3143), .A2(n2767), .ZN(n2754) );
  NAND2_X2 U3337 ( .A1(\u2/N34 ), .A2(n2738), .ZN(n2734) );
  NOR2_X4 U3338 ( .A1(\u2/exp_ovf_d[1] ), .A2(n2767), .ZN(n2758) );
  AOI22_X2 U3339 ( .A1(n2759), .A2(n1689), .B1(\u2/exp_tmp3[4] ), .B2(n2758), 
        .ZN(n2733) );
  INV_X4 U3340 ( .A(n2757), .ZN(n2738) );
  NAND2_X2 U3341 ( .A1(\u2/N33 ), .A2(n2738), .ZN(n2740) );
  AOI22_X2 U3342 ( .A1(\u2/exp_tmp4[3] ), .A2(n2759), .B1(\u2/exp_tmp3[3] ), 
        .B2(n2758), .ZN(n2739) );
  NAND3_X4 U3343 ( .A1(n2741), .A2(n2740), .A3(n2739), .ZN(\u2/N43 ) );
  INV_X4 U3344 ( .A(\u2/N37 ), .ZN(n2742) );
  NAND2_X2 U3345 ( .A1(\u2/N32 ), .A2(n2738), .ZN(n2746) );
  AOI22_X2 U3346 ( .A1(\u2/exp_tmp4[2] ), .A2(n2759), .B1(\u2/exp_tmp3[2] ), 
        .B2(n2758), .ZN(n2745) );
  NAND3_X4 U3347 ( .A1(n2747), .A2(n2746), .A3(n2745), .ZN(\u2/N42 ) );
  NAND2_X2 U3348 ( .A1(\u2/N31 ), .A2(n2738), .ZN(n2751) );
  AOI22_X2 U3349 ( .A1(\u2/exp_tmp4[1] ), .A2(n2759), .B1(\u2/exp_tmp3[1] ), 
        .B2(n2758), .ZN(n2750) );
  NAND3_X4 U3350 ( .A1(n2752), .A2(n2751), .A3(n2750), .ZN(\u2/N41 ) );
  NAND2_X2 U3351 ( .A1(\u2/lt_130/A[0] ), .A2(n2738), .ZN(n2761) );
  AOI22_X2 U3352 ( .A1(\u2/exp_tmp4[0] ), .A2(n2759), .B1(n3142), .B2(n2758), 
        .ZN(n2760) );
  NAND3_X4 U3353 ( .A1(n2762), .A2(n2761), .A3(n2760), .ZN(\u2/N40 ) );
  MUX2_X2 U3354 ( .A(n3124), .B(n3133), .S(n1733), .Z(n2763) );
  NAND2_X2 U3355 ( .A1(n3129), .A2(n3012), .ZN(n2764) );
  OAI211_X2 U3356 ( .C1(n2766), .C2(n2765), .A(n1582), .B(n2764), .ZN(
        \u2/underflow_d [1]) );
  MUX2_X2 U3357 ( .A(n2768), .B(n3135), .S(n3124), .Z(\u2/N66 ) );
  INV_X4 U3358 ( .A(n2769), .ZN(n2779) );
  NAND2_X2 U3359 ( .A1(opb_r[11]), .A2(n1725), .ZN(n2782) );
  AOI21_X4 U3360 ( .B1(n2772), .B2(n2782), .A(n2771), .ZN(n2774) );
  OAI21_X4 U3361 ( .B1(n2784), .B2(n2774), .A(n2773), .ZN(n2777) );
  INV_X4 U3362 ( .A(n2780), .ZN(n2775) );
  NOR2_X4 U3363 ( .A1(n2775), .A2(n2779), .ZN(n2776) );
  OAI21_X4 U3364 ( .B1(n2777), .B2(n2778), .A(n2776), .ZN(n2790) );
  NAND2_X2 U3365 ( .A1(n2781), .A2(n2780), .ZN(n2785) );
  INV_X4 U3366 ( .A(n2782), .ZN(n2783) );
  NAND4_X2 U3367 ( .A1(\u1/N124 ), .A2(n3145), .A3(n2787), .A4(n2786), .ZN(
        n2792) );
  INV_X4 U3368 ( .A(n2815), .ZN(n2788) );
  AND2_X2 U3369 ( .A1(n2792), .A2(n2788), .ZN(\u1/N39 ) );
  MUX2_X2 U3370 ( .A(n1560), .B(n1543), .S(n1975), .Z(n2819) );
  AND2_X2 U3371 ( .A1(n2792), .A2(n2818), .ZN(\u1/N38 ) );
  MUX2_X2 U3372 ( .A(n1573), .B(n2799), .S(n1975), .Z(n2811) );
  INV_X4 U3373 ( .A(n2811), .ZN(n2800) );
  AND2_X2 U3374 ( .A1(n2792), .A2(n2800), .ZN(\u1/N37 ) );
  MUX2_X2 U3375 ( .A(n1725), .B(n3016), .S(n1975), .Z(n2807) );
  INV_X4 U3376 ( .A(n2807), .ZN(n2796) );
  AND2_X2 U3377 ( .A1(n2792), .A2(n2796), .ZN(\u1/N36 ) );
  NAND2_X2 U3378 ( .A1(n2790), .A2(n2789), .ZN(n2791) );
  MUX2_X2 U3379 ( .A(n1723), .B(n1726), .S(n1975), .Z(n2794) );
  INV_X4 U3380 ( .A(n2794), .ZN(n2832) );
  AND2_X2 U3381 ( .A1(n2792), .A2(n2832), .ZN(\u1/N35 ) );
  MUX2_X2 U3382 ( .A(\u3/N17 ), .B(\u3/N32 ), .S(n3084), .Z(n3284) );
  MUX2_X2 U3383 ( .A(\u3/N16 ), .B(\u3/N31 ), .S(n3084), .Z(n3285) );
  MUX2_X2 U3384 ( .A(\u3/N15 ), .B(\u3/N30 ), .S(n3084), .Z(n3286) );
  MUX2_X2 U3385 ( .A(\u3/N14 ), .B(\u3/N29 ), .S(n3084), .Z(n3287) );
  MUX2_X2 U3386 ( .A(\u3/N13 ), .B(\u3/N28 ), .S(n3084), .Z(n3288) );
  MUX2_X2 U3387 ( .A(\u3/N12 ), .B(\u3/N27 ), .S(n3084), .Z(n3289) );
  MUX2_X2 U3388 ( .A(\u3/N11 ), .B(\u3/N26 ), .S(n3084), .Z(n3290) );
  MUX2_X2 U3389 ( .A(\u3/N10 ), .B(\u3/N25 ), .S(n3084), .Z(n3291) );
  MUX2_X2 U3390 ( .A(\u3/N9 ), .B(\u3/N24 ), .S(n3084), .Z(n3292) );
  MUX2_X2 U3391 ( .A(\u3/N8 ), .B(\u3/N23 ), .S(n3084), .Z(n3293) );
  MUX2_X2 U3392 ( .A(\u3/N7 ), .B(\u3/N22 ), .S(n3084), .Z(n3294) );
  MUX2_X2 U3393 ( .A(\u3/N6 ), .B(\u3/N21 ), .S(n3084), .Z(n3295) );
  MUX2_X2 U3394 ( .A(\u3/N5 ), .B(\u3/N20 ), .S(n3084), .Z(n3296) );
  MUX2_X2 U3395 ( .A(\u3/N4 ), .B(\u3/N19 ), .S(n3084), .Z(n3297) );
  MUX2_X2 U3396 ( .A(\u3/N3 ), .B(\u3/N18 ), .S(n3084), .Z(n3298) );
  MUX2_X2 U3397 ( .A(n1731), .B(n3313), .S(n2793), .Z(n1521) );
  INV_X4 U3398 ( .A(n3110), .ZN(n2958) );
  MUX2_X2 U3399 ( .A(n2958), .B(fracta_mul[9]), .S(n2793), .Z(\u1/adj_op[9] )
         );
  INV_X4 U3400 ( .A(n3109), .ZN(n2911) );
  MUX2_X2 U3401 ( .A(n2911), .B(fracta_mul[8]), .S(n1975), .Z(n3303) );
  INV_X4 U3402 ( .A(n3108), .ZN(n2905) );
  MUX2_X2 U3403 ( .A(n2905), .B(fracta_mul[7]), .S(n1975), .Z(n3304) );
  INV_X4 U3404 ( .A(n3107), .ZN(n2844) );
  INV_X4 U3405 ( .A(n3117), .ZN(n2843) );
  MUX2_X2 U3406 ( .A(n2844), .B(n2843), .S(n1975), .Z(n3305) );
  INV_X4 U3407 ( .A(n3106), .ZN(n2841) );
  INV_X4 U3408 ( .A(n3116), .ZN(n2842) );
  MUX2_X2 U3409 ( .A(n2841), .B(n2842), .S(n1975), .Z(n3306) );
  MUX2_X2 U3410 ( .A(n2895), .B(n2896), .S(n1975), .Z(n3307) );
  INV_X4 U3411 ( .A(n3104), .ZN(n2888) );
  MUX2_X2 U3412 ( .A(n2888), .B(n2889), .S(n1975), .Z(n3308) );
  INV_X4 U3413 ( .A(n3103), .ZN(n2847) );
  INV_X4 U3414 ( .A(n3113), .ZN(n2848) );
  MUX2_X2 U3415 ( .A(n2847), .B(n2848), .S(n2924), .Z(n3309) );
  INV_X4 U3416 ( .A(n3102), .ZN(n2846) );
  MUX2_X2 U3417 ( .A(n2846), .B(n3014), .S(n2924), .Z(n3310) );
  INV_X4 U3418 ( .A(n3101), .ZN(n2852) );
  MUX2_X2 U3419 ( .A(n2852), .B(n3015), .S(n2924), .Z(n3311) );
  MUX2_X2 U3420 ( .A(n1726), .B(n1723), .S(n1975), .Z(n2831) );
  INV_X4 U3421 ( .A(n2831), .ZN(n2795) );
  OAI21_X4 U3422 ( .B1(n2795), .B2(n2833), .A(n2794), .ZN(n2809) );
  MUX2_X2 U3423 ( .A(n3016), .B(n1725), .S(n1975), .Z(n2808) );
  NOR2_X4 U3424 ( .A1(n2808), .A2(n2796), .ZN(n2798) );
  NAND2_X2 U3425 ( .A1(n2796), .A2(n2808), .ZN(n2797) );
  OAI21_X4 U3426 ( .B1(n1539), .B2(n2798), .A(n2797), .ZN(n2813) );
  INV_X4 U3427 ( .A(n2813), .ZN(n2803) );
  MUX2_X2 U3428 ( .A(n2799), .B(n1573), .S(n2924), .Z(n2812) );
  NOR2_X4 U3429 ( .A1(n2812), .A2(n2800), .ZN(n2802) );
  NAND2_X2 U3430 ( .A1(n2800), .A2(n2812), .ZN(n2801) );
  OAI21_X4 U3431 ( .B1(n2803), .B2(n2802), .A(n2801), .ZN(n2817) );
  MUX2_X2 U3432 ( .A(n1543), .B(n1560), .S(n2924), .Z(n2820) );
  INV_X4 U3433 ( .A(n2820), .ZN(n2804) );
  XNOR2_X2 U3434 ( .A(n2804), .B(n2819), .ZN(n2805) );
  XNOR2_X2 U3435 ( .A(n2806), .B(n2805), .ZN(n2828) );
  XNOR2_X2 U3436 ( .A(n2808), .B(n2807), .ZN(n2810) );
  XNOR2_X2 U3437 ( .A(n2810), .B(n2809), .ZN(n2830) );
  XNOR2_X2 U3438 ( .A(n2812), .B(n2811), .ZN(n2814) );
  XNOR2_X2 U3439 ( .A(n2813), .B(n2814), .ZN(n2829) );
  NOR3_X4 U3440 ( .A1(n2828), .A2(n2830), .A3(n2829), .ZN(n2827) );
  MUX2_X2 U3441 ( .A(opb_r[14]), .B(opa_r[14]), .S(n2924), .Z(n2816) );
  NOR2_X4 U3442 ( .A1(n2816), .A2(n2815), .ZN(n2824) );
  INV_X4 U3443 ( .A(n2819), .ZN(n2818) );
  NAND2_X2 U3444 ( .A1(n2818), .A2(n2820), .ZN(n2821) );
  XNOR2_X2 U3445 ( .A(n2823), .B(n2824), .ZN(n2826) );
  INV_X4 U3446 ( .A(n2836), .ZN(n2825) );
  OAI21_X4 U3447 ( .B1(n2827), .B2(n2826), .A(n2825), .ZN(n2837) );
  OAI21_X4 U3448 ( .B1(n2836), .B2(n2828), .A(n2837), .ZN(n3302) );
  OAI21_X4 U3449 ( .B1(n2836), .B2(n2830), .A(n2837), .ZN(n3300) );
  XNOR2_X2 U3450 ( .A(n2832), .B(n2831), .ZN(n2834) );
  XNOR2_X2 U3451 ( .A(n2834), .B(n2833), .ZN(n2835) );
  MUX2_X2 U3452 ( .A(\u1/adj_op_out_sft[13] ), .B(n1731), .S(n1976), .Z(n2929)
         );
  INV_X4 U3453 ( .A(n2929), .ZN(n2839) );
  NAND2_X2 U3454 ( .A1(n2839), .A2(n2928), .ZN(\u1/fracta_s [13]) );
  MUX2_X2 U3455 ( .A(\u1/adj_op_out_sft[12] ), .B(n2958), .S(n1976), .Z(n2931)
         );
  MUX2_X2 U3456 ( .A(fracta_mul[9]), .B(\u1/adj_op_out_sft[12] ), .S(n1976), 
        .Z(n2932) );
  INV_X4 U3457 ( .A(n2932), .ZN(n2840) );
  NAND2_X2 U3458 ( .A1(n2840), .A2(n2931), .ZN(n2919) );
  MUX2_X2 U3459 ( .A(\u1/adj_op_out_sft[8] ), .B(n2841), .S(n1976), .Z(n2939)
         );
  MUX2_X2 U3460 ( .A(n2842), .B(\u1/adj_op_out_sft[8] ), .S(n1976), .Z(n2940)
         );
  INV_X4 U3461 ( .A(n2940), .ZN(n2845) );
  MUX2_X2 U3462 ( .A(n2843), .B(\u1/adj_op_out_sft[9] ), .S(n1976), .Z(n2938)
         );
  MUX2_X2 U3463 ( .A(\u1/adj_op_out_sft[9] ), .B(n2844), .S(n1976), .Z(n2937)
         );
  AOI22_X2 U3464 ( .A1(n2939), .A2(n2845), .B1(n2904), .B2(n2937), .ZN(n2910)
         );
  MUX2_X2 U3465 ( .A(n3014), .B(\u1/adj_op_out_sft[4] ), .S(n1976), .Z(n2948)
         );
  MUX2_X2 U3466 ( .A(\u1/adj_op_out_sft[5] ), .B(n2847), .S(n1976), .Z(n2945)
         );
  INV_X4 U3467 ( .A(n2945), .ZN(n2849) );
  MUX2_X2 U3468 ( .A(fracta_mul[2]), .B(\u1/adj_op_out_sft[5] ), .S(n1976), 
        .Z(n2946) );
  NOR2_X4 U3469 ( .A1(n2849), .A2(n2946), .ZN(n2850) );
  NOR2_X4 U3470 ( .A1(n2851), .A2(n2850), .ZN(n2894) );
  MUX2_X2 U3471 ( .A(\u1/adj_op_out_sft[3] ), .B(n2852), .S(n1976), .Z(n2949)
         );
  INV_X4 U3472 ( .A(n2949), .ZN(n2883) );
  MUX2_X2 U3473 ( .A(fracta_mul[0]), .B(\u1/adj_op_out_sft[3] ), .S(n1976), 
        .Z(n2950) );
  INV_X4 U3474 ( .A(n3311), .ZN(n2872) );
  INV_X4 U3475 ( .A(n3310), .ZN(n2854) );
  INV_X4 U3476 ( .A(n3309), .ZN(n2853) );
  INV_X4 U3477 ( .A(n2869), .ZN(n2857) );
  INV_X4 U3478 ( .A(n3308), .ZN(n2856) );
  INV_X4 U3479 ( .A(n3307), .ZN(n2855) );
  INV_X4 U3480 ( .A(n2864), .ZN(n2859) );
  INV_X4 U3481 ( .A(n3306), .ZN(n2862) );
  INV_X4 U3482 ( .A(n3305), .ZN(n2858) );
  INV_X4 U3483 ( .A(n2866), .ZN(n2861) );
  INV_X4 U3484 ( .A(n3304), .ZN(n2860) );
  NAND2_X2 U3485 ( .A1(n2861), .A2(n2860), .ZN(n2871) );
  INV_X4 U3486 ( .A(n2871), .ZN(n2863) );
  INV_X4 U3487 ( .A(n3302), .ZN(n2874) );
  AOI211_X4 U3488 ( .C1(\u1/exp_diff_sft[0] ), .C2(\u1/adj_op[9] ), .A(n3303), 
        .B(n2871), .ZN(n2873) );
  OAI221_X2 U3489 ( .B1(n2854), .B2(n1719), .C1(n2874), .C2(n2873), .A(n2872), 
        .ZN(n2877) );
  MUX2_X2 U3490 ( .A(n2880), .B(n2879), .S(n3301), .Z(n2881) );
  NOR2_X4 U3491 ( .A1(\u1/adj_op_out_sft[0] ), .A2(n2881), .ZN(n2927) );
  INV_X4 U3492 ( .A(n2927), .ZN(n2882) );
  NAND2_X2 U3493 ( .A1(n1720), .A2(n2948), .ZN(n2885) );
  NAND2_X2 U3494 ( .A1(n2883), .A2(n2950), .ZN(n2884) );
  INV_X4 U3495 ( .A(n2946), .ZN(n2887) );
  MUX2_X2 U3496 ( .A(\u1/adj_op_out_sft[6] ), .B(n2888), .S(n1976), .Z(n2943)
         );
  MUX2_X2 U3497 ( .A(n2889), .B(\u1/adj_op_out_sft[6] ), .S(n1976), .Z(n2944)
         );
  INV_X4 U3498 ( .A(n2944), .ZN(n2890) );
  MUX2_X2 U3499 ( .A(\u1/adj_op_out_sft[7] ), .B(n2895), .S(n1976), .Z(n2941)
         );
  INV_X4 U3500 ( .A(n2941), .ZN(n2899) );
  MUX2_X2 U3501 ( .A(n2896), .B(\u1/adj_op_out_sft[7] ), .S(n1976), .Z(n2942)
         );
  INV_X4 U3502 ( .A(n2943), .ZN(n2897) );
  OAI22_X2 U3503 ( .A1(n2899), .A2(n2942), .B1(n2944), .B2(n2897), .ZN(n2902)
         );
  INV_X4 U3504 ( .A(n2939), .ZN(n2898) );
  NAND2_X2 U3505 ( .A1(n2940), .A2(n2898), .ZN(n2901) );
  NAND2_X2 U3506 ( .A1(n2899), .A2(n2942), .ZN(n2900) );
  MUX2_X2 U3507 ( .A(\u1/adj_op_out_sft[10] ), .B(n2905), .S(n1976), .Z(n2935)
         );
  MUX2_X2 U3508 ( .A(fracta_mul[7]), .B(\u1/adj_op_out_sft[10] ), .S(n1976), 
        .Z(n2936) );
  INV_X4 U3509 ( .A(n2936), .ZN(n2906) );
  NOR2_X4 U3510 ( .A1(n2935), .A2(n2906), .ZN(n2907) );
  AOI211_X4 U3511 ( .C1(n2909), .C2(n2910), .A(n2908), .B(n2907), .ZN(n2916)
         );
  MUX2_X2 U3512 ( .A(fracta_mul[8]), .B(\u1/adj_op_out_sft[11] ), .S(n1976), 
        .Z(n2934) );
  MUX2_X2 U3513 ( .A(\u1/adj_op_out_sft[11] ), .B(n2911), .S(n1976), .Z(n2933)
         );
  INV_X4 U3514 ( .A(n2933), .ZN(n2913) );
  INV_X4 U3515 ( .A(n2935), .ZN(n2912) );
  OAI22_X2 U3516 ( .A1(n2934), .A2(n2913), .B1(n2936), .B2(n2912), .ZN(n2915)
         );
  NAND2_X2 U3517 ( .A1(n2934), .A2(n2913), .ZN(n2914) );
  OAI21_X4 U3518 ( .B1(n2916), .B2(n2915), .A(n2914), .ZN(n2918) );
  AOI21_X4 U3519 ( .B1(n2918), .B2(n2919), .A(n2917), .ZN(n2922) );
  INV_X4 U3520 ( .A(n2931), .ZN(n2920) );
  NAND2_X2 U3521 ( .A1(n2920), .A2(n2932), .ZN(n2921) );
  AOI21_X4 U3522 ( .B1(n2922), .B2(n2921), .A(n1649), .ZN(n2954) );
  MUX2_X2 U3523 ( .A(n2931), .B(n2932), .S(n1979), .Z(\u1/fracta_s [12]) );
  MUX2_X2 U3524 ( .A(n2933), .B(n2934), .S(n1979), .Z(\u1/fracta_s [11]) );
  MUX2_X2 U3525 ( .A(n2935), .B(n2936), .S(n1979), .Z(\u1/fracta_s [10]) );
  MUX2_X2 U3526 ( .A(n2937), .B(n2938), .S(n1979), .Z(\u1/fracta_s [9]) );
  MUX2_X2 U3527 ( .A(n2939), .B(n2940), .S(n1979), .Z(\u1/fracta_s [8]) );
  MUX2_X2 U3528 ( .A(n2941), .B(n2942), .S(n1979), .Z(\u1/fracta_s [7]) );
  MUX2_X2 U3529 ( .A(n2943), .B(n2944), .S(n1978), .Z(\u1/fracta_s [6]) );
  MUX2_X2 U3530 ( .A(n2945), .B(n2946), .S(n1978), .Z(\u1/fracta_s [5]) );
  MUX2_X2 U3531 ( .A(n2947), .B(n2948), .S(n1979), .Z(\u1/fracta_s [4]) );
  MUX2_X2 U3532 ( .A(n2949), .B(n2950), .S(n1979), .Z(\u1/fracta_s [3]) );
  MUX2_X2 U3533 ( .A(n1563), .B(n1590), .S(n1979), .Z(\u1/fracta_s [2]) );
  INV_X4 U3534 ( .A(n2923), .ZN(n2951) );
  MUX2_X2 U3535 ( .A(n2951), .B(n1645), .S(n1978), .Z(\u1/fracta_s [1]) );
  INV_X4 U3536 ( .A(n2925), .ZN(n2952) );
  MUX2_X2 U3537 ( .A(n2952), .B(n2953), .S(n1978), .Z(\u1/fracta_s [0]) );
  INV_X4 U3538 ( .A(n2928), .ZN(n2930) );
  MUX2_X2 U3539 ( .A(n2930), .B(n2929), .S(n1978), .Z(\u1/fractb_s [13]) );
  MUX2_X2 U3540 ( .A(n2932), .B(n2931), .S(n1979), .Z(\u1/fractb_s [12]) );
  MUX2_X2 U3541 ( .A(n2934), .B(n2933), .S(n1978), .Z(\u1/fractb_s [11]) );
  MUX2_X2 U3542 ( .A(n2936), .B(n2935), .S(n1978), .Z(\u1/fractb_s [10]) );
  MUX2_X2 U3543 ( .A(n2938), .B(n2937), .S(n1978), .Z(\u1/fractb_s [9]) );
  MUX2_X2 U3544 ( .A(n2940), .B(n2939), .S(n1978), .Z(\u1/fractb_s [8]) );
  MUX2_X2 U3545 ( .A(n2942), .B(n2941), .S(n1978), .Z(\u1/fractb_s [7]) );
  MUX2_X2 U3546 ( .A(n2944), .B(n2943), .S(n1978), .Z(\u1/fractb_s [6]) );
  MUX2_X2 U3547 ( .A(n2946), .B(n2945), .S(n1978), .Z(\u1/fractb_s [5]) );
  MUX2_X2 U3548 ( .A(n2948), .B(n2947), .S(n1978), .Z(\u1/fractb_s [4]) );
  MUX2_X2 U3549 ( .A(n2950), .B(n2949), .S(n1978), .Z(\u1/fractb_s [3]) );
  MUX2_X2 U3550 ( .A(n1590), .B(n1563), .S(n1978), .Z(\u1/fractb_s [2]) );
  MUX2_X2 U3551 ( .A(n1645), .B(n2951), .S(n1978), .Z(\u1/fractb_s [1]) );
  MUX2_X2 U3552 ( .A(n2953), .B(n2952), .S(n1978), .Z(\u1/fractb_s [0]) );
  XNOR2_X2 U3553 ( .A(n3317), .B(opb_r[15]), .ZN(n2955) );
  MUX2_X2 U3554 ( .A(n2955), .B(opa_r[15]), .S(n1978), .Z(\u1/sign_d ) );
  INV_X4 U3555 ( .A(n2956), .ZN(n2957) );
  INV_X4 U3556 ( .A(n3158), .ZN(n3312) );
  INV_X4 U3557 ( .A(n3157), .ZN(n3315) );
  OAI22_X2 U3558 ( .A1(net85778), .A2(net83361), .B1(net83438), .B2(net83439), 
        .ZN(n2960) );
  INV_X4 U3559 ( .A(net83427), .ZN(net15944) );
  XNOR2_X2 U3560 ( .A(net83407), .B(n2964), .ZN(n2966) );
  XNOR2_X2 U3561 ( .A(n2966), .B(n2965), .ZN(n2967) );
  AOI21_X4 U3562 ( .B1(net15944), .B2(n2967), .A(net83423), .ZN(n851) );
  INV_X4 U3563 ( .A(n2968), .ZN(n2969) );
  FA_X1 U3564 ( .A(n1592), .B(n2969), .CI(net89964), .S(\u4/div_exp3[1] ) );
  INV_X4 U3565 ( .A(n3010), .ZN(n3009) );
  INV_X4 U3566 ( .A(n2970), .ZN(n2973) );
  INV_X4 U3567 ( .A(n2974), .ZN(n2986) );
  NAND2_X2 U3568 ( .A1(\u4/sub_409/net10540 ), .A2(div_opa_ldz_r2[3]), .ZN(
        n2975) );
  XNOR2_X2 U3569 ( .A(net11555), .B(n2977), .ZN(n2980) );
  NAND2_X2 U3570 ( .A1(net83364), .A2(n2978), .ZN(n2979) );
  OAI221_X2 U3571 ( .B1(n2980), .B2(n2989), .C1(net83361), .C2(n1688), .A(
        n2979), .ZN(n2984) );
  INV_X4 U3572 ( .A(n2981), .ZN(n2982) );
  XNOR2_X2 U3573 ( .A(\u4/sub_409/net10540 ), .B(div_opa_ldz_r2[3]), .ZN(n2985) );
  XNOR2_X2 U3574 ( .A(n2986), .B(n2985), .ZN(n2990) );
  NAND2_X2 U3575 ( .A1(net83364), .A2(n2987), .ZN(n2988) );
  OAI221_X2 U3576 ( .B1(n2990), .B2(n2989), .C1(net83361), .C2(n1687), .A(
        n2988), .ZN(n2994) );
  AND2_X1 U3577 ( .A1(net83968), .A2(\u4/add_407/carry [3]), .ZN(
        \u4/add_407/carry [4]) );
  XOR2_X1 U3578 ( .A(\u2/gt_140/B[5] ), .B(\u2/add_111/carry[5] ), .Z(\u2/N23 ) );
  XOR2_X1 U3579 ( .A(\u2/exp_tmp4[4] ), .B(\u2/add_111/carry[4] ), .Z(\u2/N22 ) );
  XNOR2_X1 U3580 ( .A(\u2/add_111/carry[3] ), .B(\u2/lt_130/A[3] ), .ZN(
        \u2/N21 ) );
  OR2_X1 U3581 ( .A1(\u2/lt_130/A[2] ), .A2(\u2/add_111/carry[2] ), .ZN(
        \u2/add_111/carry[3] ) );
  XNOR2_X1 U3582 ( .A(\u2/add_111/carry[2] ), .B(\u2/lt_130/A[2] ), .ZN(
        \u2/N20 ) );
  OR2_X1 U3583 ( .A1(\u2/lt_130/A[1] ), .A2(\u2/lt_130/A[0] ), .ZN(
        \u2/add_111/carry[2] ) );
  XNOR2_X1 U3584 ( .A(\u2/lt_130/A[0] ), .B(\u2/lt_130/A[1] ), .ZN(\u2/N19 )
         );
  XNOR2_X1 U3585 ( .A(\u2/gt_140/B[5] ), .B(\u2/sub_111/carry[5] ), .ZN(
        \u2/N29 ) );
  XNOR2_X1 U3586 ( .A(\u2/sub_111/carry[4] ), .B(\u2/exp_tmp4[4] ), .ZN(
        \u2/N28 ) );
  XOR2_X1 U3587 ( .A(\u2/lt_130/A[3] ), .B(\u2/sub_111/carry[3] ), .Z(\u2/N27 ) );
  AND2_X1 U3588 ( .A1(\u2/sub_111/carry[2] ), .A2(\u2/lt_130/A[2] ), .ZN(
        \u2/sub_111/carry[3] ) );
  XOR2_X1 U3589 ( .A(\u2/lt_130/A[2] ), .B(\u2/sub_111/carry[2] ), .Z(\u2/N26 ) );
  AND2_X1 U3590 ( .A1(\u2/lt_130/A[0] ), .A2(\u2/lt_130/A[1] ), .ZN(
        \u2/sub_111/carry[2] ) );
  XOR2_X1 U3591 ( .A(\u2/lt_130/A[1] ), .B(\u2/lt_130/A[0] ), .Z(\u2/N25 ) );
  XOR2_X1 U3592 ( .A(opb_r[10]), .B(opa_r[10]), .Z(\u2/N12 ) );
  XNOR2_X1 U3593 ( .A(n1726), .B(opa_r[10]), .ZN(\u2/N6 ) );
  XOR2_X1 U3594 ( .A(n1635), .B(\sub_435_3/carry [20]), .Z(N151) );
  AND2_X1 U3595 ( .A1(\sub_435_3/carry [19]), .A2(n1636), .ZN(
        \sub_435_3/carry [20]) );
  XOR2_X1 U3596 ( .A(n1636), .B(\sub_435_3/carry [19]), .Z(N150) );
  AND2_X1 U3597 ( .A1(\sub_435_3/carry [18]), .A2(n1637), .ZN(
        \sub_435_3/carry [19]) );
  AND2_X1 U3598 ( .A1(\sub_435_3/carry [17]), .A2(n1672), .ZN(
        \sub_435_3/carry [18]) );
  AND2_X1 U3599 ( .A1(\sub_435_3/carry [16]), .A2(n1673), .ZN(
        \sub_435_3/carry [17]) );
  AND2_X1 U3600 ( .A1(\sub_435_3/carry [15]), .A2(n1624), .ZN(
        \sub_435_3/carry [16]) );
  AND2_X1 U3601 ( .A1(\sub_435_3/carry [14]), .A2(n1625), .ZN(
        \sub_435_3/carry [15]) );
  AND2_X1 U3602 ( .A1(\sub_435_3/carry [13]), .A2(n1626), .ZN(
        \sub_435_3/carry [14]) );
  AND2_X1 U3603 ( .A1(\sub_435_3/carry [12]), .A2(n1627), .ZN(
        \sub_435_3/carry [13]) );
  AND2_X1 U3604 ( .A1(\sub_435_3/carry [11]), .A2(n1678), .ZN(
        \sub_435_3/carry [12]) );
  AND2_X1 U3605 ( .A1(\sub_435_3/carry [10]), .A2(n1679), .ZN(
        \sub_435_3/carry [11]) );
  XOR2_X1 U3606 ( .A(n1679), .B(\sub_435_3/carry [10]), .Z(N141) );
  AND2_X1 U3607 ( .A1(\sub_435_3/carry [9]), .A2(n1674), .ZN(
        \sub_435_3/carry [10]) );
  XOR2_X1 U3608 ( .A(n1674), .B(\sub_435_3/carry [9]), .Z(N140) );
  AND2_X1 U3609 ( .A1(\sub_435_3/carry [8]), .A2(n1675), .ZN(
        \sub_435_3/carry [9]) );
  XOR2_X1 U3610 ( .A(n1675), .B(\sub_435_3/carry [8]), .Z(N139) );
  AND2_X1 U3611 ( .A1(n1680), .A2(n1676), .ZN(\sub_435_3/carry [8]) );
  XOR2_X1 U3612 ( .A(n1676), .B(n1680), .Z(N138) );
  XOR2_X1 U3613 ( .A(n1558), .B(\sub_435_b0/carry [10]), .Z(N116) );
  AND2_X1 U3614 ( .A1(\sub_435_b0/carry [9]), .A2(n1624), .ZN(
        \sub_435_b0/carry [10]) );
  XOR2_X1 U3615 ( .A(n1624), .B(\sub_435_b0/carry [9]), .Z(N115) );
  AND2_X1 U3616 ( .A1(\sub_435_b0/carry [8]), .A2(n1625), .ZN(
        \sub_435_b0/carry [9]) );
  XOR2_X1 U3617 ( .A(n1625), .B(\sub_435_b0/carry [8]), .Z(N114) );
  AND2_X1 U3618 ( .A1(\sub_435_b0/carry [7]), .A2(n1626), .ZN(
        \sub_435_b0/carry [8]) );
  XOR2_X1 U3619 ( .A(n1626), .B(\sub_435_b0/carry [7]), .Z(N113) );
  AND2_X1 U3620 ( .A1(\sub_435_b0/carry [6]), .A2(n1627), .ZN(
        \sub_435_b0/carry [7]) );
  XOR2_X1 U3621 ( .A(n1627), .B(\sub_435_b0/carry [6]), .Z(N112) );
  AND2_X1 U3622 ( .A1(\sub_435_b0/carry [5]), .A2(n1678), .ZN(
        \sub_435_b0/carry [6]) );
  XOR2_X1 U3623 ( .A(n1678), .B(\sub_435_b0/carry [5]), .Z(N111) );
  AND2_X1 U3624 ( .A1(\sub_435_b0/carry [4]), .A2(n1679), .ZN(
        \sub_435_b0/carry [5]) );
  XOR2_X1 U3625 ( .A(n1679), .B(\sub_435_b0/carry [4]), .Z(N110) );
  AND2_X1 U3626 ( .A1(\sub_435_b0/carry [3]), .A2(n1674), .ZN(
        \sub_435_b0/carry [4]) );
  AND2_X1 U3627 ( .A1(\sub_435_b0/carry [2]), .A2(n1675), .ZN(
        \sub_435_b0/carry [3]) );
  AND2_X1 U3628 ( .A1(n1680), .A2(n1676), .ZN(\sub_435_b0/carry [2]) );
  INV_X4 U3629 ( .A(\u2/sub_110/carry [5]), .ZN(\u2/N11 ) );
  XOR2_X1 U3630 ( .A(\u2/add_113/carry [4]), .B(\u2/add_113/A[4] ), .Z(
        \u2/exp_tmp3[4] ) );
  INV_X4 U3631 ( .A(\u2/lt_130/A[0] ), .ZN(\u2/exp_tmp4[0] ) );
  INV_X4 U3632 ( .A(\u2/lt_130/A[1] ), .ZN(\u2/exp_tmp4[1] ) );
  INV_X4 U3633 ( .A(\u2/lt_130/A[2] ), .ZN(\u2/exp_tmp4[2] ) );
  XOR2_X1 U3634 ( .A(\u2/add_115/carry [4]), .B(n1689), .Z(\u2/N34 ) );
  NOR2_X1 U3635 ( .A1(\u2/exp_tmp4[1] ), .A2(\u2/exp_tmp4[0] ), .ZN(n3019) );
  AOI21_X1 U3636 ( .B1(\u2/exp_tmp4[0] ), .B2(\u2/exp_tmp4[1] ), .A(n3019), 
        .ZN(n3018) );
  NAND2_X1 U3637 ( .A1(n3019), .A2(\u2/lt_130/A[2] ), .ZN(n3020) );
  OAI21_X1 U3638 ( .B1(n3019), .B2(\u2/lt_130/A[2] ), .A(n3020), .ZN(\u2/N37 )
         );
  NOR2_X1 U3639 ( .A1(\u2/exp_tmp4[3] ), .A2(n3020), .ZN(n3021) );
  INV_X4 U3640 ( .A(net83968), .ZN(\u4/sub_409/net10540 ) );
  OAI22_X1 U3641 ( .A1(fracta_mul[1]), .A2(n3022), .B1(n3022), .B2(n3046), 
        .ZN(n3024) );
  NAND2_X1 U3642 ( .A1(fracta_mul[7]), .A2(n3108), .ZN(n3025) );
  NAND2_X1 U3643 ( .A1(fracta_mul[5]), .A2(n3106), .ZN(n3033) );
  NAND2_X1 U3644 ( .A1(fracta_mul[6]), .A2(n3107), .ZN(n3034) );
  AND2_X1 U3645 ( .A1(n3033), .A2(n3034), .ZN(n3023) );
  OR2_X1 U3646 ( .A1(n3119), .A2(\u6/N8 ), .ZN(n3026) );
  NAND4_X1 U3647 ( .A1(n3024), .A2(n3025), .A3(n3023), .A4(n3026), .ZN(n3044)
         );
  NAND2_X1 U3648 ( .A1(fracta_mul[9]), .A2(n3110), .ZN(n3040) );
  AND2_X1 U3649 ( .A1(n3026), .A2(n3025), .ZN(n3037) );
  NAND2_X1 U3650 ( .A1(fracta_mul[4]), .A2(n3105), .ZN(n3042) );
  NAND2_X1 U3651 ( .A1(fracta_mul[3]), .A2(n3104), .ZN(n3041) );
  NOR2_X1 U3652 ( .A1(n3045), .A2(fracta_mul[0]), .ZN(n3028) );
  OAI21_X1 U3653 ( .B1(fracta_mul[1]), .B2(n3048), .A(n3046), .ZN(n3027) );
  NAND2_X1 U3654 ( .A1(fracta_mul[2]), .A2(n3047), .ZN(n3039) );
  OAI211_X1 U3655 ( .C1(n3028), .C2(n3049), .A(n3027), .B(n3039), .ZN(n3029)
         );
  OAI221_X1 U3656 ( .B1(fracta_mul[2]), .B2(n3047), .C1(fracta_mul[3]), .C2(
        n3104), .A(n3029), .ZN(n3030) );
  NAND3_X1 U3657 ( .A1(n3042), .A2(n3041), .A3(n3030), .ZN(n3031) );
  OAI221_X1 U3658 ( .B1(fracta_mul[4]), .B2(n3105), .C1(fracta_mul[5]), .C2(
        n3106), .A(n3031), .ZN(n3032) );
  NAND3_X1 U3659 ( .A1(n3034), .A2(n3033), .A3(n3032), .ZN(n3035) );
  OAI221_X1 U3660 ( .B1(fracta_mul[6]), .B2(n3107), .C1(fracta_mul[7]), .C2(
        n3108), .A(n3035), .ZN(n3036) );
  AOI22_X1 U3661 ( .A1(\u6/N8 ), .A2(n3119), .B1(n3037), .B2(n3036), .ZN(n3038) );
  OAI22_X1 U3662 ( .A1(fracta_mul[9]), .A2(n3110), .B1(n3052), .B2(n3038), 
        .ZN(\u1/N123 ) );
  NAND3_X1 U3663 ( .A1(n3040), .A2(n3053), .A3(n3039), .ZN(n3043) );
  NOR4_X1 U3664 ( .A1(n3044), .A2(n3043), .A3(n3050), .A4(n3051), .ZN(
        \u1/N124 ) );
  INV_X4 U3665 ( .A(\u6/N0 ), .ZN(n3045) );
  INV_X4 U3666 ( .A(\u6/N1 ), .ZN(n3046) );
  INV_X4 U3667 ( .A(\u6/N2 ), .ZN(n3047) );
  INV_X4 U3668 ( .A(n3028), .ZN(n3048) );
  INV_X4 U3669 ( .A(n3041), .ZN(n3050) );
  INV_X4 U3670 ( .A(n3042), .ZN(n3051) );
  INV_X4 U3671 ( .A(n3040), .ZN(n3052) );
  INV_X4 U3672 ( .A(\u1/N123 ), .ZN(n3053) );
  MUX2_X1 U3673 ( .A(n3122), .B(n3123), .S(n3124), .Z(n3121) );
  NAND4_X1 U3674 ( .A1(\u2/N15 ), .A2(\u2/N14 ), .A3(n3125), .A4(\u2/N13 ), 
        .ZN(n3123) );
  NOR2_X1 U3675 ( .A1(\u2/N16 ), .A2(n3126), .ZN(n3125) );
  INV_X1 U3676 ( .A(\u2/N12 ), .ZN(n3126) );
  NAND4_X1 U3677 ( .A1(\u2/N9 ), .A2(\u2/N8 ), .A3(n3127), .A4(\u2/N7 ), .ZN(
        n3122) );
  NOR2_X1 U3678 ( .A1(\u2/N10 ), .A2(n3128), .ZN(n3127) );
  INV_X1 U3679 ( .A(\u2/N6 ), .ZN(n3128) );
  NAND2_X1 U3680 ( .A1(n3134), .A2(n3124), .ZN(n3133) );
  NOR2_X1 U3681 ( .A1(n1686), .A2(n1569), .ZN(\u2/N73 ) );
  NOR2_X1 U3682 ( .A1(n3131), .A2(n3132), .ZN(n3135) );
  INV_X1 U3683 ( .A(\u2/gt_140/B[5] ), .ZN(n3132) );
  MUX2_X1 U3684 ( .A(\u2/N17 ), .B(\u2/N11 ), .S(n3136), .Z(\u2/gt_140/B[5] )
         );
  NOR2_X1 U3685 ( .A1(n1689), .A2(n3137), .ZN(n3131) );
  AND4_X1 U3686 ( .A1(\u2/lt_130/A[3] ), .A2(\u2/lt_130/A[2] ), .A3(
        \u2/lt_130/A[0] ), .A4(\u2/lt_130/A[1] ), .ZN(n3137) );
  MUX2_X1 U3687 ( .A(\u2/N13 ), .B(\u2/N7 ), .S(n3136), .Z(\u2/lt_130/A[1] )
         );
  MUX2_X1 U3688 ( .A(\u2/N12 ), .B(\u2/N6 ), .S(n3136), .Z(\u2/lt_130/A[0] )
         );
  MUX2_X1 U3689 ( .A(\u2/N14 ), .B(\u2/N8 ), .S(n3136), .Z(\u2/lt_130/A[2] )
         );
  INV_X1 U3690 ( .A(\u2/add_113/A[3] ), .ZN(n3139) );
  INV_X1 U3691 ( .A(\u2/add_113/A[2] ), .ZN(n3140) );
  INV_X1 U3692 ( .A(\u2/add_113/A[1] ), .ZN(n3141) );
  INV_X1 U3693 ( .A(\u2/add_113/A[4] ), .ZN(n3138) );
  INV_X1 U3694 ( .A(\u2/add_113/A[0] ), .ZN(n3142) );
  OAI21_X1 U3695 ( .B1(n3146), .B2(n1671), .A(n3147), .ZN(\u1/N133 ) );
  OAI21_X1 U3696 ( .B1(n3148), .B2(n1684), .A(\u1/signa_r ), .ZN(n3147) );
  NOR3_X1 U3697 ( .A1(n1681), .A2(\u1/fracta_lt_fractb ), .A3(
        \u1/fracta_eq_fractb ), .ZN(n3148) );
  AOI21_X1 U3698 ( .B1(opb_nan), .B2(n3149), .A(\u1/signa_r ), .ZN(n3146) );
  OAI21_X1 U3699 ( .B1(\u1/fracta_eq_fractb ), .B2(n1683), .A(opa_nan), .ZN(
        n3149) );
  OAI22_X1 U3700 ( .A1(n1682), .A2(n3150), .B1(n3151), .B2(n3152), .ZN(
        \u1/N122 ) );
  XNOR2_X1 U3701 ( .A(n1671), .B(\u1/add_r ), .ZN(n3152) );
  NOR2_X1 U3702 ( .A1(n3153), .A2(\u1/signa_r ), .ZN(n3151) );
  NAND2_X1 U3703 ( .A1(n3154), .A2(n3155), .ZN(\u0/N7 ) );
  NOR2_X1 U3704 ( .A1(n3155), .A2(n3154), .ZN(\u0/N6 ) );
  NOR2_X1 U3705 ( .A1(n3093), .A2(n3095), .ZN(\u0/N17 ) );
  NOR2_X1 U3706 ( .A1(n3092), .A2(n3094), .ZN(\u0/N16 ) );
  NOR2_X1 U3707 ( .A1(n3316), .A2(n3157), .ZN(\u0/N11 ) );
  NOR2_X1 U3708 ( .A1(n3314), .A2(n3158), .ZN(\u0/N10 ) );
  OAI22_X1 U3709 ( .A1(n3159), .A2(n1674), .B1(n3160), .B2(n1564), .ZN(n3281)
         );
  OAI22_X1 U3710 ( .A1(n3159), .A2(n1675), .B1(n3160), .B2(n1565), .ZN(n3282)
         );
  OAI22_X1 U3711 ( .A1(n3159), .A2(n1676), .B1(n3160), .B2(n1559), .ZN(n3283)
         );
  MUX2_X1 U3712 ( .A(\u2/N22 ), .B(\u2/N28 ), .S(n3124), .Z(\u2/add_113/A[4] )
         );
  MUX2_X1 U3713 ( .A(\u2/N21 ), .B(\u2/N27 ), .S(n3124), .Z(\u2/add_113/A[3] )
         );
  MUX2_X1 U3714 ( .A(\u2/N26 ), .B(\u2/N20 ), .S(n3136), .Z(\u2/add_113/A[2] )
         );
  MUX2_X1 U3715 ( .A(\u2/N19 ), .B(\u2/N25 ), .S(n3124), .Z(\u2/add_113/A[1] )
         );
  MUX2_X1 U3716 ( .A(\u2/exp_tmp4[0] ), .B(\u2/exp_tmp4[0] ), .S(n3136), .Z(
        \u2/add_113/A[0] ) );
  INV_X1 U3717 ( .A(n3145), .ZN(n3299) );
  XOR2_X1 U3718 ( .A(fpu_op_r1[0]), .B(\u2/sign_d ), .Z(n3145) );
  XNOR2_X1 U3719 ( .A(n1569), .B(opb_r[15]), .ZN(\u2/sign_d ) );
  INV_X1 U3720 ( .A(n3129), .ZN(n3314) );
  NAND2_X1 U3721 ( .A1(n3120), .A2(n3156), .ZN(n3129) );
  AND4_X1 U3722 ( .A1(n3118), .A2(n3113), .A3(n3119), .A4(n3161), .ZN(n3156)
         );
  NOR3_X1 U3723 ( .A1(n3014), .A2(n3162), .A3(n3015), .ZN(n3161) );
  INV_X1 U3724 ( .A(n3130), .ZN(n3316) );
  OAI22_X1 U3725 ( .A1(n3159), .A2(n1680), .B1(n3160), .B2(n1680), .ZN(n3318)
         );
  OAI22_X1 U3726 ( .A1(n1677), .A2(n3090), .B1(n1591), .B2(n3088), .ZN(n3320)
         );
  OAI22_X1 U3727 ( .A1(n1677), .A2(n3089), .B1(n1591), .B2(n3087), .ZN(n3321)
         );
  INV_X1 U3728 ( .A(n3154), .ZN(n3322) );
  NAND2_X1 U3729 ( .A1(\u0/infb_f_r ), .A2(\u0/expb_ff ), .ZN(n3154) );
  INV_X1 U3730 ( .A(n3155), .ZN(n3323) );
  NAND2_X1 U3731 ( .A1(\u0/infa_f_r ), .A2(\u0/expa_ff ), .ZN(n3155) );
  OAI222_X1 U3732 ( .A1(n3080), .A2(n3163), .B1(n3067), .B2(n3164), .C1(n3165), 
        .C2(n1636), .ZN(N99) );
  OAI222_X1 U3733 ( .A1(n3081), .A2(n3163), .B1(n3166), .B2(n1637), .C1(n3098), 
        .C2(n3068), .ZN(N98) );
  OAI222_X1 U3734 ( .A1(n3082), .A2(n3163), .B1(n3166), .B2(n1672), .C1(n3098), 
        .C2(n3069), .ZN(N97) );
  OAI222_X1 U3735 ( .A1(n3083), .A2(n3163), .B1(n3166), .B2(n1673), .C1(n3098), 
        .C2(n3070), .ZN(N96) );
  NOR2_X1 U3736 ( .A1(n3167), .A2(n3168), .ZN(N44) );
  INV_X1 U3737 ( .A(n3162), .ZN(n3167) );
  NOR2_X1 U3738 ( .A1(n3162), .A2(n3168), .ZN(N34) );
  NAND3_X1 U3739 ( .A1(n3119), .A2(n3118), .A3(n3120), .ZN(n3168) );
  NAND4_X1 U3740 ( .A1(n3117), .A2(n3116), .A3(n3115), .A4(n3114), .ZN(n3162)
         );
  NOR4_X1 U3741 ( .A1(n3169), .A2(n3068), .A3(n3070), .A4(n3069), .ZN(N296) );
  OR2_X1 U3742 ( .A1(n3066), .A2(n3067), .ZN(n3169) );
  NOR4_X1 U3743 ( .A1(opa_inf), .A2(opa_00), .A3(n3091), .A4(n1570), .ZN(N292)
         );
  NOR3_X1 U3744 ( .A1(n3164), .A2(opa_nan), .A3(n3097), .ZN(N291) );
  NOR3_X1 U3745 ( .A1(prod[11]), .A2(prod[13]), .A3(prod[12]), .ZN(n3170) );
  NOR4_X1 U3746 ( .A1(n3173), .A2(prod[4]), .A3(prod[6]), .A4(prod[5]), .ZN(
        n3172) );
  OR3_X1 U3747 ( .A1(prod[8]), .A2(prod[9]), .A3(prod[7]), .ZN(n3173) );
  NOR3_X1 U3748 ( .A1(prod[21]), .A2(prod[3]), .A3(prod[2]), .ZN(n3171) );
  XNOR2_X1 U3749 ( .A(n3174), .B(n3153), .ZN(N216) );
  INV_X1 U3750 ( .A(n3150), .ZN(n3153) );
  NAND2_X1 U3751 ( .A1(rmode_r2[1]), .A2(rmode_r2[0]), .ZN(n3150) );
  NAND2_X1 U3752 ( .A1(n3175), .A2(n3176), .ZN(N196) );
  NAND2_X1 U3753 ( .A1(n1666), .A2(n3177), .ZN(n3176) );
  NAND2_X1 U3754 ( .A1(n3175), .A2(n3178), .ZN(N195) );
  NAND2_X1 U3755 ( .A1(N151), .A2(n3177), .ZN(n3178) );
  NAND2_X1 U3756 ( .A1(n3175), .A2(n3179), .ZN(N194) );
  NAND2_X1 U3757 ( .A1(N150), .A2(n3177), .ZN(n3179) );
  OAI221_X1 U3758 ( .B1(n3180), .B2(n1578), .C1(n3181), .C2(n1635), .A(n3175), 
        .ZN(N193) );
  OAI221_X1 U3759 ( .B1(n3180), .B2(n1598), .C1(n1636), .C2(n3181), .A(n3175), 
        .ZN(N192) );
  OAI221_X1 U3760 ( .B1(n3180), .B2(n1599), .C1(n1637), .C2(n3181), .A(n3175), 
        .ZN(N191) );
  OAI221_X1 U3761 ( .B1(n3180), .B2(n1577), .C1(n1672), .C2(n3181), .A(n3175), 
        .ZN(N190) );
  OAI221_X1 U3762 ( .B1(n3180), .B2(n1562), .C1(n1673), .C2(n3181), .A(n3175), 
        .ZN(N189) );
  OAI221_X1 U3763 ( .B1(n3180), .B2(n1600), .C1(n3181), .C2(n1624), .A(n3175), 
        .ZN(N188) );
  OAI221_X1 U3764 ( .B1(n3180), .B2(n1601), .C1(n3181), .C2(n1625), .A(n3175), 
        .ZN(N187) );
  OAI221_X1 U3765 ( .B1(n3180), .B2(n1602), .C1(n3181), .C2(n1626), .A(n3175), 
        .ZN(N186) );
  OAI221_X1 U3766 ( .B1(n1558), .B2(n3159), .C1(n3181), .C2(n1627), .A(n3183), 
        .ZN(N185) );
  AOI22_X1 U3767 ( .A1(N141), .A2(n3177), .B1(N116), .B2(n3182), .ZN(n3183) );
  OAI221_X1 U3768 ( .B1(n3159), .B2(n1624), .C1(n3181), .C2(n1678), .A(n3184), 
        .ZN(N184) );
  AOI22_X1 U3769 ( .A1(N140), .A2(n3177), .B1(N115), .B2(n3182), .ZN(n3184) );
  OAI221_X1 U3770 ( .B1(n3159), .B2(n1625), .C1(n3181), .C2(n1679), .A(n3185), 
        .ZN(N183) );
  AOI22_X1 U3771 ( .A1(N139), .A2(n3177), .B1(N114), .B2(n3182), .ZN(n3185) );
  OAI221_X1 U3772 ( .B1(n3159), .B2(n1626), .C1(n1674), .C2(n3181), .A(n3186), 
        .ZN(N182) );
  AOI22_X1 U3773 ( .A1(N138), .A2(n3177), .B1(N113), .B2(n3182), .ZN(n3186) );
  OAI221_X1 U3774 ( .B1(n3159), .B2(n1627), .C1(n1675), .C2(n3181), .A(n3187), 
        .ZN(N181) );
  AOI22_X1 U3775 ( .A1(n3177), .A2(N106), .B1(N112), .B2(n3182), .ZN(n3187) );
  INV_X1 U3776 ( .A(n3180), .ZN(n3177) );
  OAI21_X1 U3777 ( .B1(n1676), .B2(n3181), .A(n3189), .ZN(N180) );
  AOI22_X1 U3778 ( .A1(N111), .A2(n3182), .B1(opa_r1[5]), .B2(n3190), .ZN(
        n3189) );
  OAI21_X1 U3779 ( .B1(n1680), .B2(n3181), .A(n3191), .ZN(N179) );
  AOI22_X1 U3780 ( .A1(N110), .A2(n3182), .B1(opa_r1[4]), .B2(n3190), .ZN(
        n3191) );
  INV_X1 U3781 ( .A(n3159), .ZN(n3190) );
  INV_X1 U3782 ( .A(n3160), .ZN(n3182) );
  NAND2_X1 U3783 ( .A1(n3192), .A2(n3188), .ZN(n3160) );
  INV_X1 U3784 ( .A(n3188), .ZN(n3174) );
  MUX2_X1 U3785 ( .A(sign_fasu), .B(sign_mul), .S(fpu_op_r2[1]), .Z(n3188) );
  NOR2_X1 U3786 ( .A1(opa_r1[11]), .A2(opa_r1[10]), .ZN(n3193) );
  OAI222_X1 U3787 ( .A1(n3079), .A2(n3163), .B1(n3066), .B2(n3164), .C1(n3165), 
        .C2(n1635), .ZN(N100) );
  INV_X1 U3788 ( .A(n3192), .ZN(n3165) );
  NOR2_X1 U3789 ( .A1(fpu_op_r2[1]), .A2(n3166), .ZN(n3192) );
  OR2_X1 U3790 ( .A1(n3097), .A2(n3099), .ZN(n3166) );
  NAND2_X1 U3791 ( .A1(n3099), .A2(fpu_op_r2[1]), .ZN(n3164) );
  NAND2_X1 U3792 ( .A1(n3099), .A2(n3098), .ZN(n3163) );
endmodule

