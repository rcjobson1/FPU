
<<<<<<< HEAD
module fpu_DW01_ash_1 ( A, DATA_TC, SH, SH_TC, B );
  input [29:0] A;
  input [4:0] SH;
  output [29:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][27] , \ML_int[1][24] , \ML_int[1][22] , \ML_int[1][21] ,
=======
module fpu_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;
  wire   [10:1] carry;

  FA_X1 U2_6 ( .A(A[6]), .B(n12), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA_X1 U2_5 ( .A(A[5]), .B(n11), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n10), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_3 ( .A(A[3]), .B(n9), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA_X1 U2_2 ( .A(A[2]), .B(n8), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA_X1 U2_1 ( .A(A[1]), .B(n13), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  XNOR2_X2 U1 ( .A(A[10]), .B(carry[10]), .ZN(DIFF[10]) );
  NAND2_X2 U2 ( .A1(n1), .A2(n2), .ZN(carry[8]) );
  XNOR2_X2 U3 ( .A(A[7]), .B(carry[7]), .ZN(DIFF[7]) );
  INV_X4 U4 ( .A(A[7]), .ZN(n1) );
  INV_X4 U5 ( .A(carry[7]), .ZN(n2) );
  NAND2_X2 U6 ( .A1(n3), .A2(n4), .ZN(carry[9]) );
  XNOR2_X2 U7 ( .A(A[8]), .B(carry[8]), .ZN(DIFF[8]) );
  INV_X4 U8 ( .A(A[8]), .ZN(n3) );
  INV_X4 U9 ( .A(carry[8]), .ZN(n4) );
  NAND2_X2 U10 ( .A1(n5), .A2(n6), .ZN(carry[10]) );
  XNOR2_X2 U11 ( .A(A[9]), .B(carry[9]), .ZN(DIFF[9]) );
  INV_X4 U12 ( .A(A[9]), .ZN(n5) );
  INV_X4 U13 ( .A(carry[9]), .ZN(n6) );
  NAND2_X2 U14 ( .A1(B[0]), .A2(n7), .ZN(carry[1]) );
  XNOR2_X2 U15 ( .A(n14), .B(A[0]), .ZN(DIFF[0]) );
  INV_X4 U16 ( .A(A[0]), .ZN(n7) );
  INV_X4 U17 ( .A(B[2]), .ZN(n8) );
  INV_X4 U18 ( .A(B[3]), .ZN(n9) );
  INV_X4 U19 ( .A(B[4]), .ZN(n10) );
  INV_X4 U20 ( .A(B[5]), .ZN(n11) );
  INV_X4 U21 ( .A(B[6]), .ZN(n12) );
  INV_X4 U22 ( .A(B[1]), .ZN(n13) );
  INV_X4 U23 ( .A(B[0]), .ZN(n14) );
endmodule


module fpu_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;
  wire   [10:1] carry;

  FA_X1 U2_6 ( .A(A[6]), .B(n8), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA_X1 U2_5 ( .A(A[5]), .B(n9), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n10), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_3 ( .A(A[3]), .B(n11), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA_X1 U2_2 ( .A(A[2]), .B(n12), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA_X1 U2_1 ( .A(A[1]), .B(n13), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  XNOR2_X2 U1 ( .A(A[10]), .B(carry[10]), .ZN(DIFF[10]) );
  NAND2_X2 U2 ( .A1(n1), .A2(n2), .ZN(carry[8]) );
  XNOR2_X2 U3 ( .A(A[7]), .B(carry[7]), .ZN(DIFF[7]) );
  INV_X4 U4 ( .A(A[7]), .ZN(n1) );
  INV_X4 U5 ( .A(carry[7]), .ZN(n2) );
  NAND2_X2 U6 ( .A1(n3), .A2(n4), .ZN(carry[9]) );
  XNOR2_X2 U7 ( .A(A[8]), .B(carry[8]), .ZN(DIFF[8]) );
  INV_X4 U8 ( .A(A[8]), .ZN(n3) );
  INV_X4 U9 ( .A(carry[8]), .ZN(n4) );
  NAND2_X2 U10 ( .A1(n5), .A2(n6), .ZN(carry[10]) );
  XNOR2_X2 U11 ( .A(A[9]), .B(carry[9]), .ZN(DIFF[9]) );
  INV_X4 U12 ( .A(A[9]), .ZN(n5) );
  INV_X4 U13 ( .A(carry[9]), .ZN(n6) );
  NAND2_X2 U14 ( .A1(B[0]), .A2(n7), .ZN(carry[1]) );
  XNOR2_X2 U15 ( .A(n14), .B(A[0]), .ZN(DIFF[0]) );
  INV_X4 U16 ( .A(A[0]), .ZN(n7) );
  INV_X4 U17 ( .A(B[6]), .ZN(n8) );
  INV_X4 U18 ( .A(B[5]), .ZN(n9) );
  INV_X4 U19 ( .A(B[4]), .ZN(n10) );
  INV_X4 U20 ( .A(B[3]), .ZN(n11) );
  INV_X4 U21 ( .A(B[2]), .ZN(n12) );
  INV_X4 U22 ( .A(B[1]), .ZN(n13) );
  INV_X4 U23 ( .A(B[0]), .ZN(n14) );
endmodule


module fpu_DW01_inc_0 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HA_X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(carry[10]), .B(A[10]), .Z(SUM[10]) );
  INV_X1 U2 ( .A(A[0]), .ZN(SUM[0]) );
endmodule


module fpu_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [105:0] A;
  input [8:0] SH;
  output [105:0] B;
  input DATA_TC, SH_TC;
  wire   \temp_int_SH[5] , \ML_int[1][105] , \ML_int[1][104] ,
         \ML_int[1][103] , \ML_int[1][102] , \ML_int[1][101] ,
         \ML_int[1][100] , \ML_int[1][99] , \ML_int[1][98] , \ML_int[1][97] ,
         \ML_int[1][96] , \ML_int[1][95] , \ML_int[1][94] , \ML_int[1][93] ,
         \ML_int[1][92] , \ML_int[1][91] , \ML_int[1][90] , \ML_int[1][89] ,
         \ML_int[1][88] , \ML_int[1][87] , \ML_int[1][86] , \ML_int[1][85] ,
         \ML_int[1][84] , \ML_int[1][83] , \ML_int[1][82] , \ML_int[1][81] ,
         \ML_int[1][80] , \ML_int[1][79] , \ML_int[1][78] , \ML_int[1][77] ,
         \ML_int[1][76] , \ML_int[1][75] , \ML_int[1][74] , \ML_int[1][73] ,
         \ML_int[1][72] , \ML_int[1][71] , \ML_int[1][70] , \ML_int[1][69] ,
         \ML_int[1][68] , \ML_int[1][67] , \ML_int[1][66] , \ML_int[1][65] ,
         \ML_int[1][64] , \ML_int[1][63] , \ML_int[1][62] , \ML_int[1][61] ,
         \ML_int[1][60] , \ML_int[1][59] , \ML_int[1][58] , \ML_int[1][57] ,
         \ML_int[1][56] , \ML_int[1][55] , \ML_int[1][54] , \ML_int[1][53] ,
         \ML_int[1][52] , \ML_int[1][51] , \ML_int[1][50] , \ML_int[1][49] ,
         \ML_int[1][48] , \ML_int[1][47] , \ML_int[1][46] , \ML_int[1][45] ,
         \ML_int[1][44] , \ML_int[1][43] , \ML_int[1][42] , \ML_int[1][41] ,
         \ML_int[1][40] , \ML_int[1][39] , \ML_int[1][38] , \ML_int[1][37] ,
         \ML_int[1][36] , \ML_int[1][35] , \ML_int[1][34] , \ML_int[1][33] ,
         \ML_int[1][32] , \ML_int[1][31] , \ML_int[1][30] , \ML_int[1][29] ,
         \ML_int[1][28] , \ML_int[1][27] , \ML_int[1][26] , \ML_int[1][25] ,
         \ML_int[1][24] , \ML_int[1][23] , \ML_int[1][22] , \ML_int[1][21] ,
         \ML_int[1][20] , \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] ,
         \ML_int[1][16] , \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] ,
         \ML_int[1][12] , \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] ,
         \ML_int[1][8] , \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] ,
         \ML_int[1][4] , \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] ,
         \ML_int[1][0] , \ML_int[2][105] , \ML_int[2][104] , \ML_int[2][103] ,
         \ML_int[2][102] , \ML_int[2][101] , \ML_int[2][100] , \ML_int[2][99] ,
         \ML_int[2][98] , \ML_int[2][97] , \ML_int[2][96] , \ML_int[2][95] ,
         \ML_int[2][94] , \ML_int[2][93] , \ML_int[2][92] , \ML_int[2][91] ,
         \ML_int[2][90] , \ML_int[2][89] , \ML_int[2][88] , \ML_int[2][87] ,
         \ML_int[2][86] , \ML_int[2][85] , \ML_int[2][84] , \ML_int[2][83] ,
         \ML_int[2][82] , \ML_int[2][81] , \ML_int[2][80] , \ML_int[2][79] ,
         \ML_int[2][78] , \ML_int[2][77] , \ML_int[2][76] , \ML_int[2][75] ,
         \ML_int[2][74] , \ML_int[2][73] , \ML_int[2][72] , \ML_int[2][71] ,
         \ML_int[2][70] , \ML_int[2][69] , \ML_int[2][68] , \ML_int[2][67] ,
         \ML_int[2][66] , \ML_int[2][65] , \ML_int[2][64] , \ML_int[2][63] ,
         \ML_int[2][62] , \ML_int[2][61] , \ML_int[2][60] , \ML_int[2][59] ,
         \ML_int[2][58] , \ML_int[2][57] , \ML_int[2][56] , \ML_int[2][55] ,
         \ML_int[2][54] , \ML_int[2][53] , \ML_int[2][52] , \ML_int[2][51] ,
         \ML_int[2][50] , \ML_int[2][49] , \ML_int[2][48] , \ML_int[2][47] ,
         \ML_int[2][46] , \ML_int[2][45] , \ML_int[2][44] , \ML_int[2][43] ,
         \ML_int[2][42] , \ML_int[2][41] , \ML_int[2][40] , \ML_int[2][39] ,
         \ML_int[2][38] , \ML_int[2][37] , \ML_int[2][36] , \ML_int[2][35] ,
         \ML_int[2][34] , \ML_int[2][33] , \ML_int[2][32] , \ML_int[2][31] ,
         \ML_int[2][30] , \ML_int[2][29] , \ML_int[2][28] , \ML_int[2][27] ,
         \ML_int[2][26] , \ML_int[2][25] , \ML_int[2][24] , \ML_int[2][23] ,
         \ML_int[2][22] , \ML_int[2][21] , \ML_int[2][20] , \ML_int[2][19] ,
         \ML_int[2][18] , \ML_int[2][17] , \ML_int[2][16] , \ML_int[2][15] ,
         \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] , \ML_int[2][11] ,
         \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] , \ML_int[2][7] ,
         \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] , \ML_int[2][3] ,
         \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] , \ML_int[3][105] ,
         \ML_int[3][104] , \ML_int[3][103] , \ML_int[3][102] ,
         \ML_int[3][101] , \ML_int[3][100] , \ML_int[3][99] , \ML_int[3][98] ,
         \ML_int[3][97] , \ML_int[3][96] , \ML_int[3][95] , \ML_int[3][94] ,
         \ML_int[3][93] , \ML_int[3][92] , \ML_int[3][91] , \ML_int[3][90] ,
         \ML_int[3][89] , \ML_int[3][88] , \ML_int[3][87] , \ML_int[3][86] ,
         \ML_int[3][85] , \ML_int[3][84] , \ML_int[3][83] , \ML_int[3][82] ,
         \ML_int[3][81] , \ML_int[3][80] , \ML_int[3][79] , \ML_int[3][78] ,
         \ML_int[3][77] , \ML_int[3][76] , \ML_int[3][75] , \ML_int[3][74] ,
         \ML_int[3][73] , \ML_int[3][72] , \ML_int[3][71] , \ML_int[3][70] ,
         \ML_int[3][69] , \ML_int[3][68] , \ML_int[3][67] , \ML_int[3][66] ,
         \ML_int[3][65] , \ML_int[3][64] , \ML_int[3][63] , \ML_int[3][62] ,
         \ML_int[3][61] , \ML_int[3][60] , \ML_int[3][59] , \ML_int[3][58] ,
         \ML_int[3][57] , \ML_int[3][56] , \ML_int[3][55] , \ML_int[3][54] ,
         \ML_int[3][53] , \ML_int[3][52] , \ML_int[3][51] , \ML_int[3][50] ,
         \ML_int[3][49] , \ML_int[3][48] , \ML_int[3][47] , \ML_int[3][46] ,
         \ML_int[3][45] , \ML_int[3][44] , \ML_int[3][43] , \ML_int[3][42] ,
         \ML_int[3][41] , \ML_int[3][40] , \ML_int[3][39] , \ML_int[3][38] ,
         \ML_int[3][37] , \ML_int[3][36] , \ML_int[3][35] , \ML_int[3][34] ,
         \ML_int[3][33] , \ML_int[3][32] , \ML_int[3][31] , \ML_int[3][30] ,
         \ML_int[3][29] , \ML_int[3][28] , \ML_int[3][27] , \ML_int[3][26] ,
         \ML_int[3][25] , \ML_int[3][24] , \ML_int[3][23] , \ML_int[3][22] ,
         \ML_int[3][21] , \ML_int[3][20] , \ML_int[3][19] , \ML_int[3][18] ,
         \ML_int[3][17] , \ML_int[3][16] , \ML_int[3][15] , \ML_int[3][14] ,
         \ML_int[3][13] , \ML_int[3][12] , \ML_int[3][11] , \ML_int[3][10] ,
         \ML_int[3][9] , \ML_int[3][8] , \ML_int[3][7] , \ML_int[3][6] ,
         \ML_int[3][5] , \ML_int[3][4] , \ML_int[3][3] , \ML_int[3][2] ,
         \ML_int[3][1] , \ML_int[3][0] , \ML_int[4][105] , \ML_int[4][104] ,
         \ML_int[4][103] , \ML_int[4][102] , \ML_int[4][101] ,
         \ML_int[4][100] , \ML_int[4][99] , \ML_int[4][98] , \ML_int[4][97] ,
         \ML_int[4][96] , \ML_int[4][95] , \ML_int[4][94] , \ML_int[4][93] ,
         \ML_int[4][92] , \ML_int[4][91] , \ML_int[4][90] , \ML_int[4][89] ,
         \ML_int[4][88] , \ML_int[4][87] , \ML_int[4][86] , \ML_int[4][85] ,
         \ML_int[4][84] , \ML_int[4][83] , \ML_int[4][82] , \ML_int[4][81] ,
         \ML_int[4][80] , \ML_int[4][79] , \ML_int[4][78] , \ML_int[4][77] ,
         \ML_int[4][76] , \ML_int[4][75] , \ML_int[4][74] , \ML_int[4][73] ,
         \ML_int[4][72] , \ML_int[4][71] , \ML_int[4][70] , \ML_int[4][69] ,
         \ML_int[4][68] , \ML_int[4][67] , \ML_int[4][66] , \ML_int[4][65] ,
         \ML_int[4][64] , \ML_int[4][63] , \ML_int[4][62] , \ML_int[4][61] ,
         \ML_int[4][60] , \ML_int[4][59] , \ML_int[4][58] , \ML_int[4][57] ,
         \ML_int[4][56] , \ML_int[4][55] , \ML_int[4][54] , \ML_int[4][53] ,
         \ML_int[4][52] , \ML_int[4][51] , \ML_int[4][50] , \ML_int[4][49] ,
         \ML_int[4][48] , \ML_int[4][47] , \ML_int[4][46] , \ML_int[4][45] ,
         \ML_int[4][44] , \ML_int[4][43] , \ML_int[4][42] , \ML_int[4][41] ,
         \ML_int[4][40] , \ML_int[4][39] , \ML_int[4][38] , \ML_int[4][37] ,
         \ML_int[4][36] , \ML_int[4][35] , \ML_int[4][34] , \ML_int[4][33] ,
         \ML_int[4][32] , \ML_int[4][31] , \ML_int[4][30] , \ML_int[4][29] ,
         \ML_int[4][28] , \ML_int[4][27] , \ML_int[4][26] , \ML_int[4][25] ,
         \ML_int[4][24] , \ML_int[4][23] , \ML_int[4][22] , \ML_int[4][21] ,
         \ML_int[4][20] , \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] ,
         \ML_int[4][16] , \ML_int[4][15] , \ML_int[4][14] , \ML_int[4][13] ,
         \ML_int[4][12] , \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] ,
         \ML_int[4][8] , \ML_int[4][7] , \ML_int[4][6] , \ML_int[4][5] ,
         \ML_int[4][4] , \ML_int[4][3] , \ML_int[4][2] , \ML_int[4][1] ,
         \ML_int[4][0] , \ML_int[5][105] , \ML_int[5][104] , \ML_int[5][103] ,
         \ML_int[5][102] , \ML_int[5][101] , \ML_int[5][100] , \ML_int[5][99] ,
         \ML_int[5][98] , \ML_int[5][97] , \ML_int[5][96] , \ML_int[5][95] ,
         \ML_int[5][94] , \ML_int[5][93] , \ML_int[5][92] , \ML_int[5][91] ,
         \ML_int[5][90] , \ML_int[5][89] , \ML_int[5][88] , \ML_int[5][87] ,
         \ML_int[5][86] , \ML_int[5][85] , \ML_int[5][84] , \ML_int[5][83] ,
         \ML_int[5][82] , \ML_int[5][81] , \ML_int[5][80] , \ML_int[5][79] ,
         \ML_int[5][78] , \ML_int[5][77] , \ML_int[5][76] , \ML_int[5][75] ,
         \ML_int[5][74] , \ML_int[5][73] , \ML_int[5][72] , \ML_int[5][71] ,
         \ML_int[5][70] , \ML_int[5][69] , \ML_int[5][68] , \ML_int[5][67] ,
         \ML_int[5][66] , \ML_int[5][65] , \ML_int[5][64] , \ML_int[5][63] ,
         \ML_int[5][62] , \ML_int[5][61] , \ML_int[5][60] , \ML_int[5][59] ,
         \ML_int[5][58] , \ML_int[5][57] , \ML_int[5][56] , \ML_int[5][55] ,
         \ML_int[5][54] , \ML_int[5][53] , \ML_int[5][52] , \ML_int[5][51] ,
         \ML_int[5][50] , \ML_int[5][49] , \ML_int[5][48] , \ML_int[5][47] ,
         \ML_int[5][46] , \ML_int[5][45] , \ML_int[5][44] , \ML_int[5][43] ,
         \ML_int[5][42] , \ML_int[5][41] , \ML_int[5][40] , \ML_int[5][39] ,
         \ML_int[5][38] , \ML_int[5][37] , \ML_int[5][36] , \ML_int[5][35] ,
         \ML_int[5][34] , \ML_int[5][33] , \ML_int[5][32] , \ML_int[5][31] ,
         \ML_int[5][30] , \ML_int[5][29] , \ML_int[5][28] , \ML_int[5][27] ,
         \ML_int[5][26] , \ML_int[5][25] , \ML_int[5][24] , \ML_int[5][23] ,
         \ML_int[5][22] , \ML_int[5][21] , \ML_int[5][20] , \ML_int[5][19] ,
         \ML_int[5][18] , \ML_int[5][17] , \ML_int[5][16] , \ML_int[5][15] ,
         \ML_int[5][14] , \ML_int[5][13] , \ML_int[5][12] , \ML_int[5][11] ,
         \ML_int[5][10] , \ML_int[5][9] , \ML_int[5][8] , \ML_int[5][7] ,
         \ML_int[5][6] , \ML_int[5][5] , \ML_int[5][4] , \ML_int[5][3] ,
         \ML_int[5][2] , \ML_int[5][1] , \ML_int[5][0] , \ML_int[6][105] ,
         \ML_int[6][104] , \ML_int[6][103] , \ML_int[6][102] ,
         \ML_int[6][101] , \ML_int[6][100] , \ML_int[6][99] , \ML_int[6][98] ,
         \ML_int[6][97] , \ML_int[6][96] , \ML_int[6][95] , \ML_int[6][94] ,
         \ML_int[6][93] , \ML_int[6][92] , \ML_int[6][91] , \ML_int[6][90] ,
         \ML_int[6][89] , \ML_int[6][88] , \ML_int[6][87] , \ML_int[6][86] ,
         \ML_int[6][85] , \ML_int[6][84] , \ML_int[6][83] , \ML_int[6][82] ,
         \ML_int[6][81] , \ML_int[6][80] , \ML_int[6][79] , \ML_int[6][78] ,
         \ML_int[6][77] , \ML_int[6][76] , \ML_int[6][75] , \ML_int[6][74] ,
         \ML_int[6][73] , \ML_int[6][72] , \ML_int[6][71] , \ML_int[6][70] ,
         \ML_int[6][69] , \ML_int[6][68] , \ML_int[6][67] , \ML_int[6][66] ,
         \ML_int[6][65] , \ML_int[6][64] , \ML_int[6][63] , \ML_int[6][62] ,
         \ML_int[6][61] , \ML_int[6][60] , \ML_int[6][59] , \ML_int[6][58] ,
         \ML_int[6][57] , \ML_int[6][56] , \ML_int[6][55] , \ML_int[6][54] ,
         \ML_int[6][53] , \ML_int[6][52] , \ML_int[6][51] , \ML_int[6][50] ,
         \ML_int[6][49] , \ML_int[6][48] , \ML_int[6][47] , \ML_int[6][46] ,
         \ML_int[6][45] , \ML_int[6][44] , \ML_int[6][43] , \ML_int[6][42] ,
         \ML_int[6][41] , \ML_int[6][40] , \ML_int[6][39] , \ML_int[6][38] ,
         \ML_int[6][37] , \ML_int[6][36] , \ML_int[6][35] , \ML_int[6][34] ,
         \ML_int[6][33] , \ML_int[6][32] , \ML_int[6][31] , \ML_int[6][30] ,
         \ML_int[6][29] , \ML_int[6][28] , \ML_int[6][27] , \ML_int[6][26] ,
         \ML_int[6][25] , \ML_int[6][24] , \ML_int[6][23] , \ML_int[6][22] ,
         \ML_int[6][21] , \ML_int[6][20] , \ML_int[6][19] , \ML_int[6][18] ,
         \ML_int[6][17] , \ML_int[6][16] , \ML_int[6][15] , \ML_int[6][14] ,
         \ML_int[6][13] , \ML_int[6][12] , \ML_int[6][11] , \ML_int[6][10] ,
         \ML_int[6][9] , \ML_int[6][8] , \ML_int[6][7] , \ML_int[6][6] ,
         \ML_int[6][5] , \ML_int[6][4] , \ML_int[6][3] , \ML_int[6][2] ,
         \ML_int[6][1] , \ML_int[6][0] , \ML_int[7][105] , \ML_int[7][104] ,
         \ML_int[7][103] , \ML_int[7][102] , \ML_int[7][101] ,
         \ML_int[7][100] , \ML_int[7][99] , \ML_int[7][98] , \ML_int[7][97] ,
         \ML_int[7][96] , \ML_int[7][95] , \ML_int[7][94] , \ML_int[7][93] ,
         \ML_int[7][92] , \ML_int[7][91] , \ML_int[7][90] , \ML_int[7][89] ,
         \ML_int[7][88] , \ML_int[7][87] , \ML_int[7][86] , \ML_int[7][85] ,
         \ML_int[7][84] , \ML_int[7][83] , \ML_int[7][82] , \ML_int[7][81] ,
         \ML_int[7][80] , \ML_int[7][79] , \ML_int[7][78] , \ML_int[7][77] ,
         \ML_int[7][76] , \ML_int[7][75] , \ML_int[7][74] , \ML_int[7][73] ,
         \ML_int[7][72] , \ML_int[7][71] , \ML_int[7][70] , \ML_int[7][69] ,
         \ML_int[7][68] , \ML_int[7][67] , \ML_int[7][66] , \ML_int[7][65] ,
         \ML_int[7][64] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88;
  wire   [6:0] SHMAG;

  MUX2_X2 M1_6_105 ( .A(\ML_int[6][105] ), .B(\ML_int[6][41] ), .S(n38), .Z(
        \ML_int[7][105] ) );
  MUX2_X2 M1_6_104 ( .A(\ML_int[6][104] ), .B(\ML_int[6][40] ), .S(n38), .Z(
        \ML_int[7][104] ) );
  MUX2_X2 M1_6_103 ( .A(\ML_int[6][103] ), .B(\ML_int[6][39] ), .S(n38), .Z(
        \ML_int[7][103] ) );
  MUX2_X2 M1_6_102 ( .A(\ML_int[6][102] ), .B(\ML_int[6][38] ), .S(n38), .Z(
        \ML_int[7][102] ) );
  MUX2_X2 M1_6_101 ( .A(\ML_int[6][101] ), .B(\ML_int[6][37] ), .S(n38), .Z(
        \ML_int[7][101] ) );
  MUX2_X2 M1_6_100 ( .A(\ML_int[6][100] ), .B(\ML_int[6][36] ), .S(n38), .Z(
        \ML_int[7][100] ) );
  MUX2_X2 M1_6_99 ( .A(\ML_int[6][99] ), .B(\ML_int[6][35] ), .S(n38), .Z(
        \ML_int[7][99] ) );
  MUX2_X2 M1_6_98 ( .A(\ML_int[6][98] ), .B(\ML_int[6][34] ), .S(n38), .Z(
        \ML_int[7][98] ) );
  MUX2_X2 M1_6_97 ( .A(\ML_int[6][97] ), .B(\ML_int[6][33] ), .S(n38), .Z(
        \ML_int[7][97] ) );
  MUX2_X2 M1_6_96 ( .A(\ML_int[6][96] ), .B(\ML_int[6][32] ), .S(n38), .Z(
        \ML_int[7][96] ) );
  MUX2_X2 M1_6_95 ( .A(\ML_int[6][95] ), .B(\ML_int[6][31] ), .S(n38), .Z(
        \ML_int[7][95] ) );
  MUX2_X2 M1_6_94 ( .A(\ML_int[6][94] ), .B(\ML_int[6][30] ), .S(n37), .Z(
        \ML_int[7][94] ) );
  MUX2_X2 M1_6_93 ( .A(\ML_int[6][93] ), .B(\ML_int[6][29] ), .S(n37), .Z(
        \ML_int[7][93] ) );
  MUX2_X2 M1_6_92 ( .A(\ML_int[6][92] ), .B(\ML_int[6][28] ), .S(n37), .Z(
        \ML_int[7][92] ) );
  MUX2_X2 M1_6_91 ( .A(\ML_int[6][91] ), .B(\ML_int[6][27] ), .S(n37), .Z(
        \ML_int[7][91] ) );
  MUX2_X2 M1_6_90 ( .A(\ML_int[6][90] ), .B(\ML_int[6][26] ), .S(n37), .Z(
        \ML_int[7][90] ) );
  MUX2_X2 M1_6_89 ( .A(\ML_int[6][89] ), .B(\ML_int[6][25] ), .S(n37), .Z(
        \ML_int[7][89] ) );
  MUX2_X2 M1_6_88 ( .A(\ML_int[6][88] ), .B(\ML_int[6][24] ), .S(n37), .Z(
        \ML_int[7][88] ) );
  MUX2_X2 M1_6_87 ( .A(\ML_int[6][87] ), .B(\ML_int[6][23] ), .S(n37), .Z(
        \ML_int[7][87] ) );
  MUX2_X2 M1_6_86 ( .A(\ML_int[6][86] ), .B(\ML_int[6][22] ), .S(n37), .Z(
        \ML_int[7][86] ) );
  MUX2_X2 M1_6_85 ( .A(\ML_int[6][85] ), .B(\ML_int[6][21] ), .S(n37), .Z(
        \ML_int[7][85] ) );
  MUX2_X2 M1_6_84 ( .A(\ML_int[6][84] ), .B(\ML_int[6][20] ), .S(n38), .Z(
        \ML_int[7][84] ) );
  MUX2_X2 M1_6_83 ( .A(\ML_int[6][83] ), .B(\ML_int[6][19] ), .S(n38), .Z(
        \ML_int[7][83] ) );
  MUX2_X2 M1_6_82 ( .A(\ML_int[6][82] ), .B(\ML_int[6][18] ), .S(n38), .Z(
        \ML_int[7][82] ) );
  MUX2_X2 M1_6_81 ( .A(\ML_int[6][81] ), .B(\ML_int[6][17] ), .S(n38), .Z(
        \ML_int[7][81] ) );
  MUX2_X2 M1_6_80 ( .A(\ML_int[6][80] ), .B(\ML_int[6][16] ), .S(n38), .Z(
        \ML_int[7][80] ) );
  MUX2_X2 M1_6_79 ( .A(\ML_int[6][79] ), .B(\ML_int[6][15] ), .S(n38), .Z(
        \ML_int[7][79] ) );
  MUX2_X2 M1_6_78 ( .A(\ML_int[6][78] ), .B(\ML_int[6][14] ), .S(n38), .Z(
        \ML_int[7][78] ) );
  MUX2_X2 M1_6_77 ( .A(\ML_int[6][77] ), .B(\ML_int[6][13] ), .S(n38), .Z(
        \ML_int[7][77] ) );
  MUX2_X2 M1_6_76 ( .A(\ML_int[6][76] ), .B(\ML_int[6][12] ), .S(n38), .Z(
        \ML_int[7][76] ) );
  MUX2_X2 M1_6_75 ( .A(\ML_int[6][75] ), .B(\ML_int[6][11] ), .S(n38), .Z(
        \ML_int[7][75] ) );
  MUX2_X2 M1_6_74 ( .A(\ML_int[6][74] ), .B(\ML_int[6][10] ), .S(n37), .Z(
        \ML_int[7][74] ) );
  MUX2_X2 M1_6_73 ( .A(\ML_int[6][73] ), .B(\ML_int[6][9] ), .S(n37), .Z(
        \ML_int[7][73] ) );
  MUX2_X2 M1_6_72 ( .A(\ML_int[6][72] ), .B(\ML_int[6][8] ), .S(n38), .Z(
        \ML_int[7][72] ) );
  MUX2_X2 M1_6_71 ( .A(\ML_int[6][71] ), .B(\ML_int[6][7] ), .S(n38), .Z(
        \ML_int[7][71] ) );
  MUX2_X2 M1_6_70 ( .A(\ML_int[6][70] ), .B(\ML_int[6][6] ), .S(n38), .Z(
        \ML_int[7][70] ) );
  MUX2_X2 M1_6_69 ( .A(\ML_int[6][69] ), .B(\ML_int[6][5] ), .S(n38), .Z(
        \ML_int[7][69] ) );
  MUX2_X2 M1_6_68 ( .A(\ML_int[6][68] ), .B(\ML_int[6][4] ), .S(n38), .Z(
        \ML_int[7][68] ) );
  MUX2_X2 M1_6_67 ( .A(\ML_int[6][67] ), .B(\ML_int[6][3] ), .S(n38), .Z(
        \ML_int[7][67] ) );
  MUX2_X2 M1_6_66 ( .A(\ML_int[6][66] ), .B(\ML_int[6][2] ), .S(n38), .Z(
        \ML_int[7][66] ) );
  MUX2_X2 M1_6_65 ( .A(\ML_int[6][65] ), .B(\ML_int[6][1] ), .S(n38), .Z(
        \ML_int[7][65] ) );
  MUX2_X2 M1_6_64 ( .A(\ML_int[6][64] ), .B(\ML_int[6][0] ), .S(n37), .Z(
        \ML_int[7][64] ) );
  MUX2_X2 M1_5_105 ( .A(\ML_int[5][105] ), .B(\ML_int[5][73] ), .S(n43), .Z(
        \ML_int[6][105] ) );
  MUX2_X2 M1_5_104 ( .A(\ML_int[5][104] ), .B(\ML_int[5][72] ), .S(n43), .Z(
        \ML_int[6][104] ) );
  MUX2_X2 M1_5_103 ( .A(\ML_int[5][103] ), .B(\ML_int[5][71] ), .S(n43), .Z(
        \ML_int[6][103] ) );
  MUX2_X2 M1_5_102 ( .A(\ML_int[5][102] ), .B(\ML_int[5][70] ), .S(n43), .Z(
        \ML_int[6][102] ) );
  MUX2_X2 M1_5_101 ( .A(\ML_int[5][101] ), .B(\ML_int[5][69] ), .S(n43), .Z(
        \ML_int[6][101] ) );
  MUX2_X2 M1_5_100 ( .A(\ML_int[5][100] ), .B(\ML_int[5][68] ), .S(n43), .Z(
        \ML_int[6][100] ) );
  MUX2_X2 M1_5_99 ( .A(\ML_int[5][99] ), .B(\ML_int[5][67] ), .S(n43), .Z(
        \ML_int[6][99] ) );
  MUX2_X2 M1_5_98 ( .A(\ML_int[5][98] ), .B(\ML_int[5][66] ), .S(n43), .Z(
        \ML_int[6][98] ) );
  MUX2_X2 M1_5_97 ( .A(\ML_int[5][97] ), .B(\ML_int[5][65] ), .S(n43), .Z(
        \ML_int[6][97] ) );
  MUX2_X2 M1_5_96 ( .A(\ML_int[5][96] ), .B(\ML_int[5][64] ), .S(n43), .Z(
        \ML_int[6][96] ) );
  MUX2_X2 M1_5_95 ( .A(\ML_int[5][95] ), .B(\ML_int[5][63] ), .S(n43), .Z(
        \ML_int[6][95] ) );
  MUX2_X2 M1_5_94 ( .A(\ML_int[5][94] ), .B(\ML_int[5][62] ), .S(n43), .Z(
        \ML_int[6][94] ) );
  MUX2_X2 M1_5_93 ( .A(\ML_int[5][93] ), .B(\ML_int[5][61] ), .S(n43), .Z(
        \ML_int[6][93] ) );
  MUX2_X2 M1_5_92 ( .A(\ML_int[5][92] ), .B(\ML_int[5][60] ), .S(n43), .Z(
        \ML_int[6][92] ) );
  MUX2_X2 M1_5_91 ( .A(\ML_int[5][91] ), .B(\ML_int[5][59] ), .S(n47), .Z(
        \ML_int[6][91] ) );
  MUX2_X2 M1_5_90 ( .A(\ML_int[5][90] ), .B(\ML_int[5][58] ), .S(n47), .Z(
        \ML_int[6][90] ) );
  MUX2_X2 M1_5_89 ( .A(\ML_int[5][89] ), .B(\ML_int[5][57] ), .S(n47), .Z(
        \ML_int[6][89] ) );
  MUX2_X2 M1_5_88 ( .A(\ML_int[5][88] ), .B(\ML_int[5][56] ), .S(n47), .Z(
        \ML_int[6][88] ) );
  MUX2_X2 M1_5_87 ( .A(\ML_int[5][87] ), .B(\ML_int[5][55] ), .S(n47), .Z(
        \ML_int[6][87] ) );
  MUX2_X2 M1_5_86 ( .A(\ML_int[5][86] ), .B(\ML_int[5][54] ), .S(n47), .Z(
        \ML_int[6][86] ) );
  MUX2_X2 M1_5_85 ( .A(\ML_int[5][85] ), .B(\ML_int[5][53] ), .S(n47), .Z(
        \ML_int[6][85] ) );
  MUX2_X2 M1_5_84 ( .A(\ML_int[5][84] ), .B(\ML_int[5][52] ), .S(n47), .Z(
        \ML_int[6][84] ) );
  MUX2_X2 M1_5_83 ( .A(\ML_int[5][83] ), .B(\ML_int[5][51] ), .S(n47), .Z(
        \ML_int[6][83] ) );
  MUX2_X2 M1_5_82 ( .A(\ML_int[5][82] ), .B(\ML_int[5][50] ), .S(n47), .Z(
        \ML_int[6][82] ) );
  MUX2_X2 M1_5_81 ( .A(\ML_int[5][81] ), .B(\ML_int[5][49] ), .S(n47), .Z(
        \ML_int[6][81] ) );
  MUX2_X2 M1_5_80 ( .A(\ML_int[5][80] ), .B(\ML_int[5][48] ), .S(n47), .Z(
        \ML_int[6][80] ) );
  MUX2_X2 M1_5_79 ( .A(\ML_int[5][79] ), .B(\ML_int[5][47] ), .S(n47), .Z(
        \ML_int[6][79] ) );
  MUX2_X2 M1_5_78 ( .A(\ML_int[5][78] ), .B(\ML_int[5][46] ), .S(n47), .Z(
        \ML_int[6][78] ) );
  MUX2_X2 M1_5_77 ( .A(\ML_int[5][77] ), .B(\ML_int[5][45] ), .S(n47), .Z(
        \ML_int[6][77] ) );
  MUX2_X2 M1_5_76 ( .A(\ML_int[5][76] ), .B(\ML_int[5][44] ), .S(n47), .Z(
        \ML_int[6][76] ) );
  MUX2_X2 M1_5_75 ( .A(\ML_int[5][75] ), .B(\ML_int[5][43] ), .S(n47), .Z(
        \ML_int[6][75] ) );
  MUX2_X2 M1_5_74 ( .A(\ML_int[5][74] ), .B(\ML_int[5][42] ), .S(n47), .Z(
        \ML_int[6][74] ) );
  MUX2_X2 M1_5_73 ( .A(\ML_int[5][73] ), .B(\ML_int[5][41] ), .S(n46), .Z(
        \ML_int[6][73] ) );
  MUX2_X2 M1_5_72 ( .A(\ML_int[5][72] ), .B(\ML_int[5][40] ), .S(n46), .Z(
        \ML_int[6][72] ) );
  MUX2_X2 M1_5_71 ( .A(\ML_int[5][71] ), .B(\ML_int[5][39] ), .S(n46), .Z(
        \ML_int[6][71] ) );
  MUX2_X2 M1_5_70 ( .A(\ML_int[5][70] ), .B(\ML_int[5][38] ), .S(n46), .Z(
        \ML_int[6][70] ) );
  MUX2_X2 M1_5_69 ( .A(\ML_int[5][69] ), .B(\ML_int[5][37] ), .S(n46), .Z(
        \ML_int[6][69] ) );
  MUX2_X2 M1_5_68 ( .A(\ML_int[5][68] ), .B(\ML_int[5][36] ), .S(n46), .Z(
        \ML_int[6][68] ) );
  MUX2_X2 M1_5_67 ( .A(\ML_int[5][67] ), .B(\ML_int[5][35] ), .S(n46), .Z(
        \ML_int[6][67] ) );
  MUX2_X2 M1_5_66 ( .A(\ML_int[5][66] ), .B(\ML_int[5][34] ), .S(n46), .Z(
        \ML_int[6][66] ) );
  MUX2_X2 M1_5_65 ( .A(\ML_int[5][65] ), .B(\ML_int[5][33] ), .S(n46), .Z(
        \ML_int[6][65] ) );
  MUX2_X2 M1_5_64 ( .A(\ML_int[5][64] ), .B(\ML_int[5][32] ), .S(n46), .Z(
        \ML_int[6][64] ) );
  MUX2_X2 M1_5_63 ( .A(\ML_int[5][63] ), .B(\ML_int[5][31] ), .S(n46), .Z(
        \ML_int[6][63] ) );
  MUX2_X2 M1_5_62 ( .A(\ML_int[5][62] ), .B(\ML_int[5][30] ), .S(n46), .Z(
        \ML_int[6][62] ) );
  MUX2_X2 M1_5_61 ( .A(\ML_int[5][61] ), .B(\ML_int[5][29] ), .S(n46), .Z(
        \ML_int[6][61] ) );
  MUX2_X2 M1_5_60 ( .A(\ML_int[5][60] ), .B(\ML_int[5][28] ), .S(n46), .Z(
        \ML_int[6][60] ) );
  MUX2_X2 M1_5_59 ( .A(\ML_int[5][59] ), .B(\ML_int[5][27] ), .S(n46), .Z(
        \ML_int[6][59] ) );
  MUX2_X2 M1_5_58 ( .A(\ML_int[5][58] ), .B(\ML_int[5][26] ), .S(n46), .Z(
        \ML_int[6][58] ) );
  MUX2_X2 M1_5_57 ( .A(\ML_int[5][57] ), .B(\ML_int[5][25] ), .S(n46), .Z(
        \ML_int[6][57] ) );
  MUX2_X2 M1_5_56 ( .A(\ML_int[5][56] ), .B(\ML_int[5][24] ), .S(n46), .Z(
        \ML_int[6][56] ) );
  MUX2_X2 M1_5_55 ( .A(\ML_int[5][55] ), .B(\ML_int[5][23] ), .S(n45), .Z(
        \ML_int[6][55] ) );
  MUX2_X2 M1_5_54 ( .A(\ML_int[5][54] ), .B(\ML_int[5][22] ), .S(n45), .Z(
        \ML_int[6][54] ) );
  MUX2_X2 M1_5_53 ( .A(\ML_int[5][53] ), .B(\ML_int[5][21] ), .S(n45), .Z(
        \ML_int[6][53] ) );
  MUX2_X2 M1_5_52 ( .A(\ML_int[5][52] ), .B(\ML_int[5][20] ), .S(n45), .Z(
        \ML_int[6][52] ) );
  MUX2_X2 M1_5_51 ( .A(\ML_int[5][51] ), .B(\ML_int[5][19] ), .S(n45), .Z(
        \ML_int[6][51] ) );
  MUX2_X2 M1_5_50 ( .A(\ML_int[5][50] ), .B(\ML_int[5][18] ), .S(n45), .Z(
        \ML_int[6][50] ) );
  MUX2_X2 M1_5_49 ( .A(\ML_int[5][49] ), .B(\ML_int[5][17] ), .S(n45), .Z(
        \ML_int[6][49] ) );
  MUX2_X2 M1_5_48 ( .A(\ML_int[5][48] ), .B(\ML_int[5][16] ), .S(n45), .Z(
        \ML_int[6][48] ) );
  MUX2_X2 M1_5_47 ( .A(\ML_int[5][47] ), .B(\ML_int[5][15] ), .S(n45), .Z(
        \ML_int[6][47] ) );
  MUX2_X2 M1_5_46 ( .A(\ML_int[5][46] ), .B(\ML_int[5][14] ), .S(n45), .Z(
        \ML_int[6][46] ) );
  MUX2_X2 M1_5_45 ( .A(\ML_int[5][45] ), .B(\ML_int[5][13] ), .S(n45), .Z(
        \ML_int[6][45] ) );
  MUX2_X2 M1_5_44 ( .A(\ML_int[5][44] ), .B(\ML_int[5][12] ), .S(n45), .Z(
        \ML_int[6][44] ) );
  MUX2_X2 M1_5_43 ( .A(\ML_int[5][43] ), .B(\ML_int[5][11] ), .S(n45), .Z(
        \ML_int[6][43] ) );
  MUX2_X2 M1_5_42 ( .A(\ML_int[5][42] ), .B(\ML_int[5][10] ), .S(n45), .Z(
        \ML_int[6][42] ) );
  MUX2_X2 M1_5_41 ( .A(\ML_int[5][41] ), .B(\ML_int[5][9] ), .S(n45), .Z(
        \ML_int[6][41] ) );
  MUX2_X2 M1_5_40 ( .A(\ML_int[5][40] ), .B(\ML_int[5][8] ), .S(n45), .Z(
        \ML_int[6][40] ) );
  MUX2_X2 M1_5_39 ( .A(\ML_int[5][39] ), .B(\ML_int[5][7] ), .S(n45), .Z(
        \ML_int[6][39] ) );
  MUX2_X2 M1_5_38 ( .A(\ML_int[5][38] ), .B(\ML_int[5][6] ), .S(n45), .Z(
        \ML_int[6][38] ) );
  MUX2_X2 M1_5_37 ( .A(\ML_int[5][37] ), .B(\ML_int[5][5] ), .S(n44), .Z(
        \ML_int[6][37] ) );
  MUX2_X2 M1_5_36 ( .A(\ML_int[5][36] ), .B(\ML_int[5][4] ), .S(n44), .Z(
        \ML_int[6][36] ) );
  MUX2_X2 M1_5_35 ( .A(\ML_int[5][35] ), .B(\ML_int[5][3] ), .S(n44), .Z(
        \ML_int[6][35] ) );
  MUX2_X2 M1_5_34 ( .A(\ML_int[5][34] ), .B(\ML_int[5][2] ), .S(n44), .Z(
        \ML_int[6][34] ) );
  MUX2_X2 M1_5_33 ( .A(\ML_int[5][33] ), .B(\ML_int[5][1] ), .S(n44), .Z(
        \ML_int[6][33] ) );
  MUX2_X2 M1_5_32 ( .A(\ML_int[5][32] ), .B(\ML_int[5][0] ), .S(n44), .Z(
        \ML_int[6][32] ) );
  MUX2_X2 M1_4_105 ( .A(\ML_int[4][105] ), .B(\ML_int[4][89] ), .S(n29), .Z(
        \ML_int[5][105] ) );
  MUX2_X2 M1_4_104 ( .A(\ML_int[4][104] ), .B(\ML_int[4][88] ), .S(n29), .Z(
        \ML_int[5][104] ) );
  MUX2_X2 M1_4_103 ( .A(\ML_int[4][103] ), .B(\ML_int[4][87] ), .S(n28), .Z(
        \ML_int[5][103] ) );
  MUX2_X2 M1_4_102 ( .A(\ML_int[4][102] ), .B(\ML_int[4][86] ), .S(n29), .Z(
        \ML_int[5][102] ) );
  MUX2_X2 M1_4_101 ( .A(\ML_int[4][101] ), .B(\ML_int[4][85] ), .S(n29), .Z(
        \ML_int[5][101] ) );
  MUX2_X2 M1_4_100 ( .A(\ML_int[4][100] ), .B(\ML_int[4][84] ), .S(n29), .Z(
        \ML_int[5][100] ) );
  MUX2_X2 M1_4_99 ( .A(\ML_int[4][99] ), .B(\ML_int[4][83] ), .S(n29), .Z(
        \ML_int[5][99] ) );
  MUX2_X2 M1_4_98 ( .A(\ML_int[4][98] ), .B(\ML_int[4][82] ), .S(n29), .Z(
        \ML_int[5][98] ) );
  MUX2_X2 M1_4_97 ( .A(\ML_int[4][97] ), .B(\ML_int[4][81] ), .S(n29), .Z(
        \ML_int[5][97] ) );
  MUX2_X2 M1_4_96 ( .A(\ML_int[4][96] ), .B(\ML_int[4][80] ), .S(n29), .Z(
        \ML_int[5][96] ) );
  MUX2_X2 M1_4_95 ( .A(\ML_int[4][95] ), .B(\ML_int[4][79] ), .S(n29), .Z(
        \ML_int[5][95] ) );
  MUX2_X2 M1_4_94 ( .A(\ML_int[4][94] ), .B(\ML_int[4][78] ), .S(n29), .Z(
        \ML_int[5][94] ) );
  MUX2_X2 M1_4_93 ( .A(\ML_int[4][93] ), .B(\ML_int[4][77] ), .S(n29), .Z(
        \ML_int[5][93] ) );
  MUX2_X2 M1_4_92 ( .A(\ML_int[4][92] ), .B(\ML_int[4][76] ), .S(n27), .Z(
        \ML_int[5][92] ) );
  MUX2_X2 M1_4_91 ( .A(\ML_int[4][91] ), .B(\ML_int[4][75] ), .S(n28), .Z(
        \ML_int[5][91] ) );
  MUX2_X2 M1_4_90 ( .A(\ML_int[4][90] ), .B(\ML_int[4][74] ), .S(n27), .Z(
        \ML_int[5][90] ) );
  MUX2_X2 M1_4_89 ( .A(\ML_int[4][89] ), .B(\ML_int[4][73] ), .S(n28), .Z(
        \ML_int[5][89] ) );
  MUX2_X2 M1_4_88 ( .A(\ML_int[4][88] ), .B(\ML_int[4][72] ), .S(n27), .Z(
        \ML_int[5][88] ) );
  MUX2_X2 M1_4_87 ( .A(\ML_int[4][87] ), .B(\ML_int[4][71] ), .S(n27), .Z(
        \ML_int[5][87] ) );
  MUX2_X2 M1_4_86 ( .A(\ML_int[4][86] ), .B(\ML_int[4][70] ), .S(n27), .Z(
        \ML_int[5][86] ) );
  MUX2_X2 M1_4_85 ( .A(\ML_int[4][85] ), .B(\ML_int[4][69] ), .S(n27), .Z(
        \ML_int[5][85] ) );
  MUX2_X2 M1_4_84 ( .A(\ML_int[4][84] ), .B(\ML_int[4][68] ), .S(n27), .Z(
        \ML_int[5][84] ) );
  MUX2_X2 M1_4_83 ( .A(\ML_int[4][83] ), .B(\ML_int[4][67] ), .S(n27), .Z(
        \ML_int[5][83] ) );
  MUX2_X2 M1_4_82 ( .A(\ML_int[4][82] ), .B(\ML_int[4][66] ), .S(n27), .Z(
        \ML_int[5][82] ) );
  MUX2_X2 M1_4_81 ( .A(\ML_int[4][81] ), .B(\ML_int[4][65] ), .S(n30), .Z(
        \ML_int[5][81] ) );
  MUX2_X2 M1_4_80 ( .A(\ML_int[4][80] ), .B(\ML_int[4][64] ), .S(n30), .Z(
        \ML_int[5][80] ) );
  MUX2_X2 M1_4_79 ( .A(\ML_int[4][79] ), .B(\ML_int[4][63] ), .S(n31), .Z(
        \ML_int[5][79] ) );
  MUX2_X2 M1_4_78 ( .A(\ML_int[4][78] ), .B(\ML_int[4][62] ), .S(n31), .Z(
        \ML_int[5][78] ) );
  MUX2_X2 M1_4_77 ( .A(\ML_int[4][77] ), .B(\ML_int[4][61] ), .S(n31), .Z(
        \ML_int[5][77] ) );
  MUX2_X2 M1_4_76 ( .A(\ML_int[4][76] ), .B(\ML_int[4][60] ), .S(n31), .Z(
        \ML_int[5][76] ) );
  MUX2_X2 M1_4_75 ( .A(\ML_int[4][75] ), .B(\ML_int[4][59] ), .S(n31), .Z(
        \ML_int[5][75] ) );
  MUX2_X2 M1_4_74 ( .A(\ML_int[4][74] ), .B(\ML_int[4][58] ), .S(n31), .Z(
        \ML_int[5][74] ) );
  MUX2_X2 M1_4_73 ( .A(\ML_int[4][73] ), .B(\ML_int[4][57] ), .S(n31), .Z(
        \ML_int[5][73] ) );
  MUX2_X2 M1_4_72 ( .A(\ML_int[4][72] ), .B(\ML_int[4][56] ), .S(n31), .Z(
        \ML_int[5][72] ) );
  MUX2_X2 M1_4_71 ( .A(\ML_int[4][71] ), .B(\ML_int[4][55] ), .S(n31), .Z(
        \ML_int[5][71] ) );
  MUX2_X2 M1_4_70 ( .A(\ML_int[4][70] ), .B(\ML_int[4][54] ), .S(n30), .Z(
        \ML_int[5][70] ) );
  MUX2_X2 M1_4_69 ( .A(\ML_int[4][69] ), .B(\ML_int[4][53] ), .S(n30), .Z(
        \ML_int[5][69] ) );
  MUX2_X2 M1_4_68 ( .A(\ML_int[4][68] ), .B(\ML_int[4][52] ), .S(n30), .Z(
        \ML_int[5][68] ) );
  MUX2_X2 M1_4_67 ( .A(\ML_int[4][67] ), .B(\ML_int[4][51] ), .S(n30), .Z(
        \ML_int[5][67] ) );
  MUX2_X2 M1_4_66 ( .A(\ML_int[4][66] ), .B(\ML_int[4][50] ), .S(n30), .Z(
        \ML_int[5][66] ) );
  MUX2_X2 M1_4_65 ( .A(\ML_int[4][65] ), .B(\ML_int[4][49] ), .S(n30), .Z(
        \ML_int[5][65] ) );
  MUX2_X2 M1_4_64 ( .A(\ML_int[4][64] ), .B(\ML_int[4][48] ), .S(n30), .Z(
        \ML_int[5][64] ) );
  MUX2_X2 M1_4_63 ( .A(\ML_int[4][63] ), .B(\ML_int[4][47] ), .S(n30), .Z(
        \ML_int[5][63] ) );
  MUX2_X2 M1_4_62 ( .A(\ML_int[4][62] ), .B(\ML_int[4][46] ), .S(n30), .Z(
        \ML_int[5][62] ) );
  MUX2_X2 M1_4_61 ( .A(\ML_int[4][61] ), .B(\ML_int[4][45] ), .S(n30), .Z(
        \ML_int[5][61] ) );
  MUX2_X2 M1_4_60 ( .A(\ML_int[4][60] ), .B(\ML_int[4][44] ), .S(n30), .Z(
        \ML_int[5][60] ) );
  MUX2_X2 M1_4_59 ( .A(\ML_int[4][59] ), .B(\ML_int[4][43] ), .S(n29), .Z(
        \ML_int[5][59] ) );
  MUX2_X2 M1_4_58 ( .A(\ML_int[4][58] ), .B(\ML_int[4][42] ), .S(n29), .Z(
        \ML_int[5][58] ) );
  MUX2_X2 M1_4_57 ( .A(\ML_int[4][57] ), .B(\ML_int[4][41] ), .S(n29), .Z(
        \ML_int[5][57] ) );
  MUX2_X2 M1_4_56 ( .A(\ML_int[4][56] ), .B(\ML_int[4][40] ), .S(n29), .Z(
        \ML_int[5][56] ) );
  MUX2_X2 M1_4_55 ( .A(\ML_int[4][55] ), .B(\ML_int[4][39] ), .S(n29), .Z(
        \ML_int[5][55] ) );
  MUX2_X2 M1_4_54 ( .A(\ML_int[4][54] ), .B(\ML_int[4][38] ), .S(n29), .Z(
        \ML_int[5][54] ) );
  MUX2_X2 M1_4_53 ( .A(\ML_int[4][53] ), .B(\ML_int[4][37] ), .S(n30), .Z(
        \ML_int[5][53] ) );
  MUX2_X2 M1_4_52 ( .A(\ML_int[4][52] ), .B(\ML_int[4][36] ), .S(n30), .Z(
        \ML_int[5][52] ) );
  MUX2_X2 M1_4_51 ( .A(\ML_int[4][51] ), .B(\ML_int[4][35] ), .S(n30), .Z(
        \ML_int[5][51] ) );
  MUX2_X2 M1_4_50 ( .A(\ML_int[4][50] ), .B(\ML_int[4][34] ), .S(n30), .Z(
        \ML_int[5][50] ) );
  MUX2_X2 M1_4_49 ( .A(\ML_int[4][49] ), .B(\ML_int[4][33] ), .S(n30), .Z(
        \ML_int[5][49] ) );
  MUX2_X2 M1_4_48 ( .A(\ML_int[4][48] ), .B(\ML_int[4][32] ), .S(n32), .Z(
        \ML_int[5][48] ) );
  MUX2_X2 M1_4_47 ( .A(\ML_int[4][47] ), .B(\ML_int[4][31] ), .S(n32), .Z(
        \ML_int[5][47] ) );
  MUX2_X2 M1_4_46 ( .A(\ML_int[4][46] ), .B(\ML_int[4][30] ), .S(n32), .Z(
        \ML_int[5][46] ) );
  MUX2_X2 M1_4_45 ( .A(\ML_int[4][45] ), .B(\ML_int[4][29] ), .S(n32), .Z(
        \ML_int[5][45] ) );
  MUX2_X2 M1_4_44 ( .A(\ML_int[4][44] ), .B(\ML_int[4][28] ), .S(n32), .Z(
        \ML_int[5][44] ) );
  MUX2_X2 M1_4_43 ( .A(\ML_int[4][43] ), .B(\ML_int[4][27] ), .S(n27), .Z(
        \ML_int[5][43] ) );
  MUX2_X2 M1_4_42 ( .A(\ML_int[4][42] ), .B(\ML_int[4][26] ), .S(n27), .Z(
        \ML_int[5][42] ) );
  MUX2_X2 M1_4_41 ( .A(\ML_int[4][41] ), .B(\ML_int[4][25] ), .S(n27), .Z(
        \ML_int[5][41] ) );
  MUX2_X2 M1_4_40 ( .A(\ML_int[4][40] ), .B(\ML_int[4][24] ), .S(n27), .Z(
        \ML_int[5][40] ) );
  MUX2_X2 M1_4_39 ( .A(\ML_int[4][39] ), .B(\ML_int[4][23] ), .S(n27), .Z(
        \ML_int[5][39] ) );
  MUX2_X2 M1_4_38 ( .A(\ML_int[4][38] ), .B(\ML_int[4][22] ), .S(n28), .Z(
        \ML_int[5][38] ) );
  MUX2_X2 M1_4_37 ( .A(\ML_int[4][37] ), .B(\ML_int[4][21] ), .S(n32), .Z(
        \ML_int[5][37] ) );
  MUX2_X2 M1_4_36 ( .A(\ML_int[4][36] ), .B(\ML_int[4][20] ), .S(n32), .Z(
        \ML_int[5][36] ) );
  MUX2_X2 M1_4_35 ( .A(\ML_int[4][35] ), .B(\ML_int[4][19] ), .S(n32), .Z(
        \ML_int[5][35] ) );
  MUX2_X2 M1_4_34 ( .A(\ML_int[4][34] ), .B(\ML_int[4][18] ), .S(n32), .Z(
        \ML_int[5][34] ) );
  MUX2_X2 M1_4_33 ( .A(\ML_int[4][33] ), .B(\ML_int[4][17] ), .S(n32), .Z(
        \ML_int[5][33] ) );
  MUX2_X2 M1_4_32 ( .A(\ML_int[4][32] ), .B(\ML_int[4][16] ), .S(n32), .Z(
        \ML_int[5][32] ) );
  MUX2_X2 M1_4_31 ( .A(\ML_int[4][31] ), .B(\ML_int[4][15] ), .S(n32), .Z(
        \ML_int[5][31] ) );
  MUX2_X2 M1_4_30 ( .A(\ML_int[4][30] ), .B(\ML_int[4][14] ), .S(n32), .Z(
        \ML_int[5][30] ) );
  MUX2_X2 M1_4_29 ( .A(\ML_int[4][29] ), .B(\ML_int[4][13] ), .S(n32), .Z(
        \ML_int[5][29] ) );
  MUX2_X2 M1_4_28 ( .A(\ML_int[4][28] ), .B(\ML_int[4][12] ), .S(n32), .Z(
        \ML_int[5][28] ) );
  MUX2_X2 M1_4_27 ( .A(\ML_int[4][27] ), .B(\ML_int[4][11] ), .S(n32), .Z(
        \ML_int[5][27] ) );
  MUX2_X2 M1_4_26 ( .A(\ML_int[4][26] ), .B(\ML_int[4][10] ), .S(n31), .Z(
        \ML_int[5][26] ) );
  MUX2_X2 M1_4_25 ( .A(\ML_int[4][25] ), .B(\ML_int[4][9] ), .S(n31), .Z(
        \ML_int[5][25] ) );
  MUX2_X2 M1_4_24 ( .A(\ML_int[4][24] ), .B(\ML_int[4][8] ), .S(n31), .Z(
        \ML_int[5][24] ) );
  MUX2_X2 M1_4_23 ( .A(\ML_int[4][23] ), .B(\ML_int[4][7] ), .S(n31), .Z(
        \ML_int[5][23] ) );
  MUX2_X2 M1_4_22 ( .A(\ML_int[4][22] ), .B(\ML_int[4][6] ), .S(n31), .Z(
        \ML_int[5][22] ) );
  MUX2_X2 M1_4_21 ( .A(\ML_int[4][21] ), .B(\ML_int[4][5] ), .S(n31), .Z(
        \ML_int[5][21] ) );
  MUX2_X2 M1_4_20 ( .A(\ML_int[4][20] ), .B(\ML_int[4][4] ), .S(n31), .Z(
        \ML_int[5][20] ) );
  MUX2_X2 M1_4_19 ( .A(\ML_int[4][19] ), .B(\ML_int[4][3] ), .S(n31), .Z(
        \ML_int[5][19] ) );
  MUX2_X2 M1_4_18 ( .A(\ML_int[4][18] ), .B(\ML_int[4][2] ), .S(n31), .Z(
        \ML_int[5][18] ) );
  MUX2_X2 M1_4_17 ( .A(\ML_int[4][17] ), .B(\ML_int[4][1] ), .S(n32), .Z(
        \ML_int[5][17] ) );
  MUX2_X2 M1_4_16 ( .A(\ML_int[4][16] ), .B(\ML_int[4][0] ), .S(n32), .Z(
        \ML_int[5][16] ) );
  MUX2_X2 M1_3_105 ( .A(\ML_int[3][105] ), .B(\ML_int[3][97] ), .S(n18), .Z(
        \ML_int[4][105] ) );
  MUX2_X2 M1_3_104 ( .A(\ML_int[3][104] ), .B(\ML_int[3][96] ), .S(n18), .Z(
        \ML_int[4][104] ) );
  MUX2_X2 M1_3_103 ( .A(\ML_int[3][103] ), .B(\ML_int[3][95] ), .S(n18), .Z(
        \ML_int[4][103] ) );
  MUX2_X2 M1_3_102 ( .A(\ML_int[3][102] ), .B(\ML_int[3][94] ), .S(n18), .Z(
        \ML_int[4][102] ) );
  MUX2_X2 M1_3_101 ( .A(\ML_int[3][101] ), .B(\ML_int[3][93] ), .S(n18), .Z(
        \ML_int[4][101] ) );
  MUX2_X2 M1_3_100 ( .A(\ML_int[3][100] ), .B(\ML_int[3][92] ), .S(n18), .Z(
        \ML_int[4][100] ) );
  MUX2_X2 M1_3_99 ( .A(\ML_int[3][99] ), .B(\ML_int[3][91] ), .S(n18), .Z(
        \ML_int[4][99] ) );
  MUX2_X2 M1_3_98 ( .A(\ML_int[3][98] ), .B(\ML_int[3][90] ), .S(n18), .Z(
        \ML_int[4][98] ) );
  MUX2_X2 M1_3_97 ( .A(\ML_int[3][97] ), .B(\ML_int[3][89] ), .S(n19), .Z(
        \ML_int[4][97] ) );
  MUX2_X2 M1_3_96 ( .A(\ML_int[3][96] ), .B(\ML_int[3][88] ), .S(n19), .Z(
        \ML_int[4][96] ) );
  MUX2_X2 M1_3_95 ( .A(\ML_int[3][95] ), .B(\ML_int[3][87] ), .S(n18), .Z(
        \ML_int[4][95] ) );
  MUX2_X2 M1_3_94 ( .A(\ML_int[3][94] ), .B(\ML_int[3][86] ), .S(n18), .Z(
        \ML_int[4][94] ) );
  MUX2_X2 M1_3_93 ( .A(\ML_int[3][93] ), .B(\ML_int[3][85] ), .S(n18), .Z(
        \ML_int[4][93] ) );
  MUX2_X2 M1_3_92 ( .A(\ML_int[3][92] ), .B(\ML_int[3][84] ), .S(n18), .Z(
        \ML_int[4][92] ) );
  MUX2_X2 M1_3_91 ( .A(\ML_int[3][91] ), .B(\ML_int[3][83] ), .S(n18), .Z(
        \ML_int[4][91] ) );
  MUX2_X2 M1_3_90 ( .A(\ML_int[3][90] ), .B(\ML_int[3][82] ), .S(n18), .Z(
        \ML_int[4][90] ) );
  MUX2_X2 M1_3_89 ( .A(\ML_int[3][89] ), .B(\ML_int[3][81] ), .S(n18), .Z(
        \ML_int[4][89] ) );
  MUX2_X2 M1_3_88 ( .A(\ML_int[3][88] ), .B(\ML_int[3][80] ), .S(n18), .Z(
        \ML_int[4][88] ) );
  MUX2_X2 M1_3_87 ( .A(\ML_int[3][87] ), .B(\ML_int[3][79] ), .S(n18), .Z(
        \ML_int[4][87] ) );
  MUX2_X2 M1_3_86 ( .A(\ML_int[3][86] ), .B(\ML_int[3][78] ), .S(n18), .Z(
        \ML_int[4][86] ) );
  MUX2_X2 M1_3_85 ( .A(\ML_int[3][85] ), .B(\ML_int[3][77] ), .S(n18), .Z(
        \ML_int[4][85] ) );
  MUX2_X2 M1_3_84 ( .A(\ML_int[3][84] ), .B(\ML_int[3][76] ), .S(n18), .Z(
        \ML_int[4][84] ) );
  MUX2_X2 M1_3_83 ( .A(\ML_int[3][83] ), .B(\ML_int[3][75] ), .S(n18), .Z(
        \ML_int[4][83] ) );
  MUX2_X2 M1_3_82 ( .A(\ML_int[3][82] ), .B(\ML_int[3][74] ), .S(n18), .Z(
        \ML_int[4][82] ) );
  MUX2_X2 M1_3_81 ( .A(\ML_int[3][81] ), .B(\ML_int[3][73] ), .S(n18), .Z(
        \ML_int[4][81] ) );
  MUX2_X2 M1_3_80 ( .A(\ML_int[3][80] ), .B(\ML_int[3][72] ), .S(n18), .Z(
        \ML_int[4][80] ) );
  MUX2_X2 M1_3_79 ( .A(\ML_int[3][79] ), .B(\ML_int[3][71] ), .S(n18), .Z(
        \ML_int[4][79] ) );
  MUX2_X2 M1_3_78 ( .A(\ML_int[3][78] ), .B(\ML_int[3][70] ), .S(n18), .Z(
        \ML_int[4][78] ) );
  MUX2_X2 M1_3_77 ( .A(\ML_int[3][77] ), .B(\ML_int[3][69] ), .S(n18), .Z(
        \ML_int[4][77] ) );
  MUX2_X2 M1_3_76 ( .A(\ML_int[3][76] ), .B(\ML_int[3][68] ), .S(n18), .Z(
        \ML_int[4][76] ) );
  MUX2_X2 M1_3_75 ( .A(\ML_int[3][75] ), .B(\ML_int[3][67] ), .S(n18), .Z(
        \ML_int[4][75] ) );
  MUX2_X2 M1_3_74 ( .A(\ML_int[3][74] ), .B(\ML_int[3][66] ), .S(n18), .Z(
        \ML_int[4][74] ) );
  MUX2_X2 M1_3_73 ( .A(\ML_int[3][73] ), .B(\ML_int[3][65] ), .S(n20), .Z(
        \ML_int[4][73] ) );
  MUX2_X2 M1_3_72 ( .A(\ML_int[3][72] ), .B(\ML_int[3][64] ), .S(n20), .Z(
        \ML_int[4][72] ) );
  MUX2_X2 M1_3_71 ( .A(\ML_int[3][71] ), .B(\ML_int[3][63] ), .S(n20), .Z(
        \ML_int[4][71] ) );
  MUX2_X2 M1_3_70 ( .A(\ML_int[3][70] ), .B(\ML_int[3][62] ), .S(n20), .Z(
        \ML_int[4][70] ) );
  MUX2_X2 M1_3_69 ( .A(\ML_int[3][69] ), .B(\ML_int[3][61] ), .S(n20), .Z(
        \ML_int[4][69] ) );
  MUX2_X2 M1_3_68 ( .A(\ML_int[3][68] ), .B(\ML_int[3][60] ), .S(n20), .Z(
        \ML_int[4][68] ) );
  MUX2_X2 M1_3_67 ( .A(\ML_int[3][67] ), .B(\ML_int[3][59] ), .S(n20), .Z(
        \ML_int[4][67] ) );
  MUX2_X2 M1_3_66 ( .A(\ML_int[3][66] ), .B(\ML_int[3][58] ), .S(n20), .Z(
        \ML_int[4][66] ) );
  MUX2_X2 M1_3_65 ( .A(\ML_int[3][65] ), .B(\ML_int[3][57] ), .S(n20), .Z(
        \ML_int[4][65] ) );
  MUX2_X2 M1_3_64 ( .A(\ML_int[3][64] ), .B(\ML_int[3][56] ), .S(n20), .Z(
        \ML_int[4][64] ) );
  MUX2_X2 M1_3_63 ( .A(\ML_int[3][63] ), .B(\ML_int[3][55] ), .S(n20), .Z(
        \ML_int[4][63] ) );
  MUX2_X2 M1_3_62 ( .A(\ML_int[3][62] ), .B(\ML_int[3][54] ), .S(n19), .Z(
        \ML_int[4][62] ) );
  MUX2_X2 M1_3_61 ( .A(\ML_int[3][61] ), .B(\ML_int[3][53] ), .S(n19), .Z(
        \ML_int[4][61] ) );
  MUX2_X2 M1_3_60 ( .A(\ML_int[3][60] ), .B(\ML_int[3][52] ), .S(n19), .Z(
        \ML_int[4][60] ) );
  MUX2_X2 M1_3_59 ( .A(\ML_int[3][59] ), .B(\ML_int[3][51] ), .S(n19), .Z(
        \ML_int[4][59] ) );
  MUX2_X2 M1_3_58 ( .A(\ML_int[3][58] ), .B(\ML_int[3][50] ), .S(n19), .Z(
        \ML_int[4][58] ) );
  MUX2_X2 M1_3_57 ( .A(\ML_int[3][57] ), .B(\ML_int[3][49] ), .S(n20), .Z(
        \ML_int[4][57] ) );
  MUX2_X2 M1_3_56 ( .A(\ML_int[3][56] ), .B(\ML_int[3][48] ), .S(n20), .Z(
        \ML_int[4][56] ) );
  MUX2_X2 M1_3_55 ( .A(\ML_int[3][55] ), .B(\ML_int[3][47] ), .S(n20), .Z(
        \ML_int[4][55] ) );
  MUX2_X2 M1_3_54 ( .A(\ML_int[3][54] ), .B(\ML_int[3][46] ), .S(n20), .Z(
        \ML_int[4][54] ) );
  MUX2_X2 M1_3_53 ( .A(\ML_int[3][53] ), .B(\ML_int[3][45] ), .S(n20), .Z(
        \ML_int[4][53] ) );
  MUX2_X2 M1_3_52 ( .A(\ML_int[3][52] ), .B(\ML_int[3][44] ), .S(n20), .Z(
        \ML_int[4][52] ) );
  MUX2_X2 M1_3_51 ( .A(\ML_int[3][51] ), .B(\ML_int[3][43] ), .S(n19), .Z(
        \ML_int[4][51] ) );
  MUX2_X2 M1_3_50 ( .A(\ML_int[3][50] ), .B(\ML_int[3][42] ), .S(n19), .Z(
        \ML_int[4][50] ) );
  MUX2_X2 M1_3_49 ( .A(\ML_int[3][49] ), .B(\ML_int[3][41] ), .S(n19), .Z(
        \ML_int[4][49] ) );
  MUX2_X2 M1_3_48 ( .A(\ML_int[3][48] ), .B(\ML_int[3][40] ), .S(n19), .Z(
        \ML_int[4][48] ) );
  MUX2_X2 M1_3_47 ( .A(\ML_int[3][47] ), .B(\ML_int[3][39] ), .S(n19), .Z(
        \ML_int[4][47] ) );
  MUX2_X2 M1_3_46 ( .A(\ML_int[3][46] ), .B(\ML_int[3][38] ), .S(n19), .Z(
        \ML_int[4][46] ) );
  MUX2_X2 M1_3_45 ( .A(\ML_int[3][45] ), .B(\ML_int[3][37] ), .S(n19), .Z(
        \ML_int[4][45] ) );
  MUX2_X2 M1_3_44 ( .A(\ML_int[3][44] ), .B(\ML_int[3][36] ), .S(n19), .Z(
        \ML_int[4][44] ) );
  MUX2_X2 M1_3_43 ( .A(\ML_int[3][43] ), .B(\ML_int[3][35] ), .S(n19), .Z(
        \ML_int[4][43] ) );
  MUX2_X2 M1_3_42 ( .A(\ML_int[3][42] ), .B(\ML_int[3][34] ), .S(n19), .Z(
        \ML_int[4][42] ) );
  MUX2_X2 M1_3_41 ( .A(\ML_int[3][41] ), .B(\ML_int[3][33] ), .S(n19), .Z(
        \ML_int[4][41] ) );
  MUX2_X2 M1_3_40 ( .A(\ML_int[3][40] ), .B(\ML_int[3][32] ), .S(n19), .Z(
        \ML_int[4][40] ) );
  MUX2_X2 M1_3_39 ( .A(\ML_int[3][39] ), .B(\ML_int[3][31] ), .S(n20), .Z(
        \ML_int[4][39] ) );
  MUX2_X2 M1_3_38 ( .A(\ML_int[3][38] ), .B(\ML_int[3][30] ), .S(n24), .Z(
        \ML_int[4][38] ) );
  MUX2_X2 M1_3_37 ( .A(\ML_int[3][37] ), .B(\ML_int[3][29] ), .S(n18), .Z(
        \ML_int[4][37] ) );
  MUX2_X2 M1_3_36 ( .A(\ML_int[3][36] ), .B(\ML_int[3][28] ), .S(n18), .Z(
        \ML_int[4][36] ) );
  MUX2_X2 M1_3_35 ( .A(\ML_int[3][35] ), .B(\ML_int[3][27] ), .S(n18), .Z(
        \ML_int[4][35] ) );
  MUX2_X2 M1_3_34 ( .A(\ML_int[3][34] ), .B(\ML_int[3][26] ), .S(n18), .Z(
        \ML_int[4][34] ) );
  MUX2_X2 M1_3_33 ( .A(\ML_int[3][33] ), .B(\ML_int[3][25] ), .S(n18), .Z(
        \ML_int[4][33] ) );
  MUX2_X2 M1_3_32 ( .A(\ML_int[3][32] ), .B(\ML_int[3][24] ), .S(n18), .Z(
        \ML_int[4][32] ) );
  MUX2_X2 M1_3_31 ( .A(\ML_int[3][31] ), .B(\ML_int[3][23] ), .S(n18), .Z(
        \ML_int[4][31] ) );
  MUX2_X2 M1_3_30 ( .A(\ML_int[3][30] ), .B(\ML_int[3][22] ), .S(n18), .Z(
        \ML_int[4][30] ) );
  MUX2_X2 M1_3_29 ( .A(\ML_int[3][29] ), .B(\ML_int[3][21] ), .S(n21), .Z(
        \ML_int[4][29] ) );
  MUX2_X2 M1_3_28 ( .A(\ML_int[3][28] ), .B(\ML_int[3][20] ), .S(n21), .Z(
        \ML_int[4][28] ) );
  MUX2_X2 M1_3_27 ( .A(\ML_int[3][27] ), .B(\ML_int[3][19] ), .S(n21), .Z(
        \ML_int[4][27] ) );
  MUX2_X2 M1_3_26 ( .A(\ML_int[3][26] ), .B(\ML_int[3][18] ), .S(n21), .Z(
        \ML_int[4][26] ) );
  MUX2_X2 M1_3_25 ( .A(\ML_int[3][25] ), .B(\ML_int[3][17] ), .S(n21), .Z(
        \ML_int[4][25] ) );
  MUX2_X2 M1_3_24 ( .A(\ML_int[3][24] ), .B(\ML_int[3][16] ), .S(n21), .Z(
        \ML_int[4][24] ) );
  MUX2_X2 M1_3_23 ( .A(\ML_int[3][23] ), .B(\ML_int[3][15] ), .S(n21), .Z(
        \ML_int[4][23] ) );
  MUX2_X2 M1_3_22 ( .A(\ML_int[3][22] ), .B(\ML_int[3][14] ), .S(n21), .Z(
        \ML_int[4][22] ) );
  MUX2_X2 M1_3_21 ( .A(\ML_int[3][21] ), .B(\ML_int[3][13] ), .S(n18), .Z(
        \ML_int[4][21] ) );
  MUX2_X2 M1_3_20 ( .A(\ML_int[3][20] ), .B(\ML_int[3][12] ), .S(n18), .Z(
        \ML_int[4][20] ) );
  MUX2_X2 M1_3_19 ( .A(\ML_int[3][19] ), .B(\ML_int[3][11] ), .S(n18), .Z(
        \ML_int[4][19] ) );
  MUX2_X2 M1_3_18 ( .A(\ML_int[3][18] ), .B(\ML_int[3][10] ), .S(n20), .Z(
        \ML_int[4][18] ) );
  MUX2_X2 M1_3_17 ( .A(\ML_int[3][17] ), .B(\ML_int[3][9] ), .S(n21), .Z(
        \ML_int[4][17] ) );
  MUX2_X2 M1_3_16 ( .A(\ML_int[3][16] ), .B(\ML_int[3][8] ), .S(n21), .Z(
        \ML_int[4][16] ) );
  MUX2_X2 M1_3_15 ( .A(\ML_int[3][15] ), .B(\ML_int[3][7] ), .S(n21), .Z(
        \ML_int[4][15] ) );
  MUX2_X2 M1_3_14 ( .A(\ML_int[3][14] ), .B(\ML_int[3][6] ), .S(n21), .Z(
        \ML_int[4][14] ) );
  MUX2_X2 M1_3_13 ( .A(\ML_int[3][13] ), .B(\ML_int[3][5] ), .S(n21), .Z(
        \ML_int[4][13] ) );
  MUX2_X2 M1_3_12 ( .A(\ML_int[3][12] ), .B(\ML_int[3][4] ), .S(n21), .Z(
        \ML_int[4][12] ) );
  MUX2_X2 M1_3_11 ( .A(\ML_int[3][11] ), .B(\ML_int[3][3] ), .S(n21), .Z(
        \ML_int[4][11] ) );
  MUX2_X2 M1_3_10 ( .A(\ML_int[3][10] ), .B(\ML_int[3][2] ), .S(n21), .Z(
        \ML_int[4][10] ) );
  MUX2_X2 M1_3_9 ( .A(\ML_int[3][9] ), .B(\ML_int[3][1] ), .S(n21), .Z(
        \ML_int[4][9] ) );
  MUX2_X2 M1_3_8 ( .A(\ML_int[3][8] ), .B(\ML_int[3][0] ), .S(n21), .Z(
        \ML_int[4][8] ) );
  MUX2_X2 M1_2_105 ( .A(\ML_int[2][105] ), .B(\ML_int[2][101] ), .S(n15), .Z(
        \ML_int[3][105] ) );
  MUX2_X2 M1_2_104 ( .A(\ML_int[2][104] ), .B(\ML_int[2][100] ), .S(n15), .Z(
        \ML_int[3][104] ) );
  MUX2_X2 M1_2_103 ( .A(\ML_int[2][103] ), .B(\ML_int[2][99] ), .S(n15), .Z(
        \ML_int[3][103] ) );
  MUX2_X2 M1_2_102 ( .A(\ML_int[2][102] ), .B(\ML_int[2][98] ), .S(n15), .Z(
        \ML_int[3][102] ) );
  MUX2_X2 M1_2_101 ( .A(\ML_int[2][101] ), .B(\ML_int[2][97] ), .S(n15), .Z(
        \ML_int[3][101] ) );
  MUX2_X2 M1_2_100 ( .A(\ML_int[2][100] ), .B(\ML_int[2][96] ), .S(n15), .Z(
        \ML_int[3][100] ) );
  MUX2_X2 M1_2_99 ( .A(\ML_int[2][99] ), .B(\ML_int[2][95] ), .S(n15), .Z(
        \ML_int[3][99] ) );
  MUX2_X2 M1_2_98 ( .A(\ML_int[2][98] ), .B(\ML_int[2][94] ), .S(n15), .Z(
        \ML_int[3][98] ) );
  MUX2_X2 M1_2_97 ( .A(\ML_int[2][97] ), .B(\ML_int[2][93] ), .S(n15), .Z(
        \ML_int[3][97] ) );
  MUX2_X2 M1_2_96 ( .A(\ML_int[2][96] ), .B(\ML_int[2][92] ), .S(n15), .Z(
        \ML_int[3][96] ) );
  MUX2_X2 M1_2_95 ( .A(\ML_int[2][95] ), .B(\ML_int[2][91] ), .S(n15), .Z(
        \ML_int[3][95] ) );
  MUX2_X2 M1_2_94 ( .A(\ML_int[2][94] ), .B(\ML_int[2][90] ), .S(n15), .Z(
        \ML_int[3][94] ) );
  MUX2_X2 M1_2_93 ( .A(\ML_int[2][93] ), .B(\ML_int[2][89] ), .S(n15), .Z(
        \ML_int[3][93] ) );
  MUX2_X2 M1_2_92 ( .A(\ML_int[2][92] ), .B(\ML_int[2][88] ), .S(n15), .Z(
        \ML_int[3][92] ) );
  MUX2_X2 M1_2_91 ( .A(\ML_int[2][91] ), .B(\ML_int[2][87] ), .S(n17), .Z(
        \ML_int[3][91] ) );
  MUX2_X2 M1_2_90 ( .A(\ML_int[2][90] ), .B(\ML_int[2][86] ), .S(n17), .Z(
        \ML_int[3][90] ) );
  MUX2_X2 M1_2_89 ( .A(\ML_int[2][89] ), .B(\ML_int[2][85] ), .S(n17), .Z(
        \ML_int[3][89] ) );
  MUX2_X2 M1_2_88 ( .A(\ML_int[2][88] ), .B(\ML_int[2][84] ), .S(n17), .Z(
        \ML_int[3][88] ) );
  MUX2_X2 M1_2_87 ( .A(\ML_int[2][87] ), .B(\ML_int[2][83] ), .S(n17), .Z(
        \ML_int[3][87] ) );
  MUX2_X2 M1_2_86 ( .A(\ML_int[2][86] ), .B(\ML_int[2][82] ), .S(n17), .Z(
        \ML_int[3][86] ) );
  MUX2_X2 M1_2_85 ( .A(\ML_int[2][85] ), .B(\ML_int[2][81] ), .S(n17), .Z(
        \ML_int[3][85] ) );
  MUX2_X2 M1_2_84 ( .A(\ML_int[2][84] ), .B(\ML_int[2][80] ), .S(n15), .Z(
        \ML_int[3][84] ) );
  MUX2_X2 M1_2_83 ( .A(\ML_int[2][83] ), .B(\ML_int[2][79] ), .S(n15), .Z(
        \ML_int[3][83] ) );
  MUX2_X2 M1_2_82 ( .A(\ML_int[2][82] ), .B(\ML_int[2][78] ), .S(n15), .Z(
        \ML_int[3][82] ) );
  MUX2_X2 M1_2_81 ( .A(\ML_int[2][81] ), .B(\ML_int[2][77] ), .S(n15), .Z(
        \ML_int[3][81] ) );
  MUX2_X2 M1_2_80 ( .A(\ML_int[2][80] ), .B(\ML_int[2][76] ), .S(n15), .Z(
        \ML_int[3][80] ) );
  MUX2_X2 M1_2_79 ( .A(\ML_int[2][79] ), .B(\ML_int[2][75] ), .S(n15), .Z(
        \ML_int[3][79] ) );
  MUX2_X2 M1_2_78 ( .A(\ML_int[2][78] ), .B(\ML_int[2][74] ), .S(n15), .Z(
        \ML_int[3][78] ) );
  MUX2_X2 M1_2_77 ( .A(\ML_int[2][77] ), .B(\ML_int[2][73] ), .S(n15), .Z(
        \ML_int[3][77] ) );
  MUX2_X2 M1_2_76 ( .A(\ML_int[2][76] ), .B(\ML_int[2][72] ), .S(n15), .Z(
        \ML_int[3][76] ) );
  MUX2_X2 M1_2_75 ( .A(\ML_int[2][75] ), .B(\ML_int[2][71] ), .S(n15), .Z(
        \ML_int[3][75] ) );
  MUX2_X2 M1_2_74 ( .A(\ML_int[2][74] ), .B(\ML_int[2][70] ), .S(n15), .Z(
        \ML_int[3][74] ) );
  MUX2_X2 M1_2_73 ( .A(\ML_int[2][73] ), .B(\ML_int[2][69] ), .S(n15), .Z(
        \ML_int[3][73] ) );
  MUX2_X2 M1_2_72 ( .A(\ML_int[2][72] ), .B(\ML_int[2][68] ), .S(n16), .Z(
        \ML_int[3][72] ) );
  MUX2_X2 M1_2_71 ( .A(\ML_int[2][71] ), .B(\ML_int[2][67] ), .S(n17), .Z(
        \ML_int[3][71] ) );
  MUX2_X2 M1_2_70 ( .A(\ML_int[2][70] ), .B(\ML_int[2][66] ), .S(n14), .Z(
        \ML_int[3][70] ) );
  MUX2_X2 M1_2_69 ( .A(\ML_int[2][69] ), .B(\ML_int[2][65] ), .S(n14), .Z(
        \ML_int[3][69] ) );
  MUX2_X2 M1_2_68 ( .A(\ML_int[2][68] ), .B(\ML_int[2][64] ), .S(n15), .Z(
        \ML_int[3][68] ) );
  MUX2_X2 M1_2_67 ( .A(\ML_int[2][67] ), .B(\ML_int[2][63] ), .S(n15), .Z(
        \ML_int[3][67] ) );
  MUX2_X2 M1_2_66 ( .A(\ML_int[2][66] ), .B(\ML_int[2][62] ), .S(n15), .Z(
        \ML_int[3][66] ) );
  MUX2_X2 M1_2_65 ( .A(\ML_int[2][65] ), .B(\ML_int[2][61] ), .S(n15), .Z(
        \ML_int[3][65] ) );
  MUX2_X2 M1_2_64 ( .A(\ML_int[2][64] ), .B(\ML_int[2][60] ), .S(n15), .Z(
        \ML_int[3][64] ) );
  MUX2_X2 M1_2_63 ( .A(\ML_int[2][63] ), .B(\ML_int[2][59] ), .S(n15), .Z(
        \ML_int[3][63] ) );
  MUX2_X2 M1_2_62 ( .A(\ML_int[2][62] ), .B(\ML_int[2][58] ), .S(n15), .Z(
        \ML_int[3][62] ) );
  MUX2_X2 M1_2_61 ( .A(\ML_int[2][61] ), .B(\ML_int[2][57] ), .S(n15), .Z(
        \ML_int[3][61] ) );
  MUX2_X2 M1_2_60 ( .A(\ML_int[2][60] ), .B(\ML_int[2][56] ), .S(n15), .Z(
        \ML_int[3][60] ) );
  MUX2_X2 M1_2_59 ( .A(\ML_int[2][59] ), .B(\ML_int[2][55] ), .S(n15), .Z(
        \ML_int[3][59] ) );
  MUX2_X2 M1_2_58 ( .A(\ML_int[2][58] ), .B(\ML_int[2][54] ), .S(n14), .Z(
        \ML_int[3][58] ) );
  MUX2_X2 M1_2_57 ( .A(\ML_int[2][57] ), .B(\ML_int[2][53] ), .S(n14), .Z(
        \ML_int[3][57] ) );
  MUX2_X2 M1_2_56 ( .A(\ML_int[2][56] ), .B(\ML_int[2][52] ), .S(n14), .Z(
        \ML_int[3][56] ) );
  MUX2_X2 M1_2_55 ( .A(\ML_int[2][55] ), .B(\ML_int[2][51] ), .S(n14), .Z(
        \ML_int[3][55] ) );
  MUX2_X2 M1_2_54 ( .A(\ML_int[2][54] ), .B(\ML_int[2][50] ), .S(n14), .Z(
        \ML_int[3][54] ) );
  MUX2_X2 M1_2_53 ( .A(\ML_int[2][53] ), .B(\ML_int[2][49] ), .S(n14), .Z(
        \ML_int[3][53] ) );
  MUX2_X2 M1_2_52 ( .A(\ML_int[2][52] ), .B(\ML_int[2][48] ), .S(n14), .Z(
        \ML_int[3][52] ) );
  MUX2_X2 M1_2_51 ( .A(\ML_int[2][51] ), .B(\ML_int[2][47] ), .S(n14), .Z(
        \ML_int[3][51] ) );
  MUX2_X2 M1_2_50 ( .A(\ML_int[2][50] ), .B(\ML_int[2][46] ), .S(n14), .Z(
        \ML_int[3][50] ) );
  MUX2_X2 M1_2_49 ( .A(\ML_int[2][49] ), .B(\ML_int[2][45] ), .S(n14), .Z(
        \ML_int[3][49] ) );
  MUX2_X2 M1_2_48 ( .A(\ML_int[2][48] ), .B(\ML_int[2][44] ), .S(n14), .Z(
        \ML_int[3][48] ) );
  MUX2_X2 M1_2_47 ( .A(\ML_int[2][47] ), .B(\ML_int[2][43] ), .S(n16), .Z(
        \ML_int[3][47] ) );
  MUX2_X2 M1_2_46 ( .A(\ML_int[2][46] ), .B(\ML_int[2][42] ), .S(n16), .Z(
        \ML_int[3][46] ) );
  MUX2_X2 M1_2_45 ( .A(\ML_int[2][45] ), .B(\ML_int[2][41] ), .S(n16), .Z(
        \ML_int[3][45] ) );
  MUX2_X2 M1_2_44 ( .A(\ML_int[2][44] ), .B(\ML_int[2][40] ), .S(n16), .Z(
        \ML_int[3][44] ) );
  MUX2_X2 M1_2_43 ( .A(\ML_int[2][43] ), .B(\ML_int[2][39] ), .S(n16), .Z(
        \ML_int[3][43] ) );
  MUX2_X2 M1_2_42 ( .A(\ML_int[2][42] ), .B(\ML_int[2][38] ), .S(n16), .Z(
        \ML_int[3][42] ) );
  MUX2_X2 M1_2_41 ( .A(\ML_int[2][41] ), .B(\ML_int[2][37] ), .S(n16), .Z(
        \ML_int[3][41] ) );
  MUX2_X2 M1_2_40 ( .A(\ML_int[2][40] ), .B(\ML_int[2][36] ), .S(n16), .Z(
        \ML_int[3][40] ) );
  MUX2_X2 M1_2_39 ( .A(\ML_int[2][39] ), .B(\ML_int[2][35] ), .S(n16), .Z(
        \ML_int[3][39] ) );
  MUX2_X2 M1_2_38 ( .A(\ML_int[2][38] ), .B(\ML_int[2][34] ), .S(n16), .Z(
        \ML_int[3][38] ) );
  MUX2_X2 M1_2_37 ( .A(\ML_int[2][37] ), .B(\ML_int[2][33] ), .S(n16), .Z(
        \ML_int[3][37] ) );
  MUX2_X2 M1_2_36 ( .A(\ML_int[2][36] ), .B(\ML_int[2][32] ), .S(n15), .Z(
        \ML_int[3][36] ) );
  MUX2_X2 M1_2_35 ( .A(\ML_int[2][35] ), .B(\ML_int[2][31] ), .S(n15), .Z(
        \ML_int[3][35] ) );
  MUX2_X2 M1_2_34 ( .A(\ML_int[2][34] ), .B(\ML_int[2][30] ), .S(n15), .Z(
        \ML_int[3][34] ) );
  MUX2_X2 M1_2_33 ( .A(\ML_int[2][33] ), .B(\ML_int[2][29] ), .S(n17), .Z(
        \ML_int[3][33] ) );
  MUX2_X2 M1_2_32 ( .A(\ML_int[2][32] ), .B(\ML_int[2][28] ), .S(n16), .Z(
        \ML_int[3][32] ) );
  MUX2_X2 M1_2_31 ( .A(\ML_int[2][31] ), .B(\ML_int[2][27] ), .S(n16), .Z(
        \ML_int[3][31] ) );
  MUX2_X2 M1_2_30 ( .A(\ML_int[2][30] ), .B(\ML_int[2][26] ), .S(n16), .Z(
        \ML_int[3][30] ) );
  MUX2_X2 M1_2_29 ( .A(\ML_int[2][29] ), .B(\ML_int[2][25] ), .S(n16), .Z(
        \ML_int[3][29] ) );
  MUX2_X2 M1_2_28 ( .A(\ML_int[2][28] ), .B(\ML_int[2][24] ), .S(n16), .Z(
        \ML_int[3][28] ) );
  MUX2_X2 M1_2_27 ( .A(\ML_int[2][27] ), .B(\ML_int[2][23] ), .S(n16), .Z(
        \ML_int[3][27] ) );
  MUX2_X2 M1_2_26 ( .A(\ML_int[2][26] ), .B(\ML_int[2][22] ), .S(n16), .Z(
        \ML_int[3][26] ) );
  MUX2_X2 M1_2_25 ( .A(\ML_int[2][25] ), .B(\ML_int[2][21] ), .S(n16), .Z(
        \ML_int[3][25] ) );
  MUX2_X2 M1_2_24 ( .A(\ML_int[2][24] ), .B(\ML_int[2][20] ), .S(n17), .Z(
        \ML_int[3][24] ) );
  MUX2_X2 M1_2_23 ( .A(\ML_int[2][23] ), .B(\ML_int[2][19] ), .S(n14), .Z(
        \ML_int[3][23] ) );
  MUX2_X2 M1_2_22 ( .A(\ML_int[2][22] ), .B(\ML_int[2][18] ), .S(n17), .Z(
        \ML_int[3][22] ) );
  MUX2_X2 M1_2_21 ( .A(\ML_int[2][21] ), .B(\ML_int[2][17] ), .S(n15), .Z(
        \ML_int[3][21] ) );
  MUX2_X2 M1_2_20 ( .A(\ML_int[2][20] ), .B(\ML_int[2][16] ), .S(n15), .Z(
        \ML_int[3][20] ) );
  MUX2_X2 M1_2_19 ( .A(\ML_int[2][19] ), .B(\ML_int[2][15] ), .S(n15), .Z(
        \ML_int[3][19] ) );
  MUX2_X2 M1_2_18 ( .A(\ML_int[2][18] ), .B(\ML_int[2][14] ), .S(n15), .Z(
        \ML_int[3][18] ) );
  MUX2_X2 M1_2_17 ( .A(\ML_int[2][17] ), .B(\ML_int[2][13] ), .S(n17), .Z(
        \ML_int[3][17] ) );
  MUX2_X2 M1_2_16 ( .A(\ML_int[2][16] ), .B(\ML_int[2][12] ), .S(n17), .Z(
        \ML_int[3][16] ) );
  MUX2_X2 M1_2_15 ( .A(\ML_int[2][15] ), .B(\ML_int[2][11] ), .S(n14), .Z(
        \ML_int[3][15] ) );
  MUX2_X2 M1_2_14 ( .A(\ML_int[2][14] ), .B(\ML_int[2][10] ), .S(n17), .Z(
        \ML_int[3][14] ) );
  MUX2_X2 M1_2_13 ( .A(\ML_int[2][13] ), .B(\ML_int[2][9] ), .S(n17), .Z(
        \ML_int[3][13] ) );
  MUX2_X2 M1_2_12 ( .A(\ML_int[2][12] ), .B(\ML_int[2][8] ), .S(n17), .Z(
        \ML_int[3][12] ) );
  MUX2_X2 M1_2_11 ( .A(\ML_int[2][11] ), .B(\ML_int[2][7] ), .S(n17), .Z(
        \ML_int[3][11] ) );
  MUX2_X2 M1_2_10 ( .A(\ML_int[2][10] ), .B(\ML_int[2][6] ), .S(n17), .Z(
        \ML_int[3][10] ) );
  MUX2_X2 M1_2_9 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S(n17), .Z(
        \ML_int[3][9] ) );
  MUX2_X2 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(n17), .Z(
        \ML_int[3][8] ) );
  MUX2_X2 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(n17), .Z(
        \ML_int[3][7] ) );
  MUX2_X2 M1_2_6 ( .A(\ML_int[2][6] ), .B(\ML_int[2][2] ), .S(n17), .Z(
        \ML_int[3][6] ) );
  MUX2_X2 M1_2_5 ( .A(\ML_int[2][5] ), .B(\ML_int[2][1] ), .S(n17), .Z(
        \ML_int[3][5] ) );
  MUX2_X2 M1_2_4 ( .A(\ML_int[2][4] ), .B(\ML_int[2][0] ), .S(n17), .Z(
        \ML_int[3][4] ) );
  MUX2_X2 M1_1_105 ( .A(\ML_int[1][105] ), .B(\ML_int[1][103] ), .S(n11), .Z(
        \ML_int[2][105] ) );
  MUX2_X2 M1_1_104 ( .A(\ML_int[1][104] ), .B(\ML_int[1][102] ), .S(n11), .Z(
        \ML_int[2][104] ) );
  MUX2_X2 M1_1_103 ( .A(\ML_int[1][103] ), .B(\ML_int[1][101] ), .S(n11), .Z(
        \ML_int[2][103] ) );
  MUX2_X2 M1_1_102 ( .A(\ML_int[1][102] ), .B(\ML_int[1][100] ), .S(n11), .Z(
        \ML_int[2][102] ) );
  MUX2_X2 M1_1_101 ( .A(\ML_int[1][101] ), .B(\ML_int[1][99] ), .S(n11), .Z(
        \ML_int[2][101] ) );
  MUX2_X2 M1_1_100 ( .A(\ML_int[1][100] ), .B(\ML_int[1][98] ), .S(n11), .Z(
        \ML_int[2][100] ) );
  MUX2_X2 M1_1_99 ( .A(\ML_int[1][99] ), .B(\ML_int[1][97] ), .S(n11), .Z(
        \ML_int[2][99] ) );
  MUX2_X2 M1_1_98 ( .A(\ML_int[1][98] ), .B(\ML_int[1][96] ), .S(n11), .Z(
        \ML_int[2][98] ) );
  MUX2_X2 M1_1_97 ( .A(\ML_int[1][97] ), .B(\ML_int[1][95] ), .S(n11), .Z(
        \ML_int[2][97] ) );
  MUX2_X2 M1_1_96 ( .A(\ML_int[1][96] ), .B(\ML_int[1][94] ), .S(n11), .Z(
        \ML_int[2][96] ) );
  MUX2_X2 M1_1_95 ( .A(\ML_int[1][95] ), .B(\ML_int[1][93] ), .S(n11), .Z(
        \ML_int[2][95] ) );
  MUX2_X2 M1_1_94 ( .A(\ML_int[1][94] ), .B(\ML_int[1][92] ), .S(n11), .Z(
        \ML_int[2][94] ) );
  MUX2_X2 M1_1_93 ( .A(\ML_int[1][93] ), .B(\ML_int[1][91] ), .S(n11), .Z(
        \ML_int[2][93] ) );
  MUX2_X2 M1_1_92 ( .A(\ML_int[1][92] ), .B(\ML_int[1][90] ), .S(n11), .Z(
        \ML_int[2][92] ) );
  MUX2_X2 M1_1_91 ( .A(\ML_int[1][91] ), .B(\ML_int[1][89] ), .S(n11), .Z(
        \ML_int[2][91] ) );
  MUX2_X2 M1_1_90 ( .A(\ML_int[1][90] ), .B(\ML_int[1][88] ), .S(n11), .Z(
        \ML_int[2][90] ) );
  MUX2_X2 M1_1_89 ( .A(\ML_int[1][89] ), .B(\ML_int[1][87] ), .S(n12), .Z(
        \ML_int[2][89] ) );
  MUX2_X2 M1_1_88 ( .A(\ML_int[1][88] ), .B(\ML_int[1][86] ), .S(n13), .Z(
        \ML_int[2][88] ) );
  MUX2_X2 M1_1_87 ( .A(\ML_int[1][87] ), .B(\ML_int[1][85] ), .S(n12), .Z(
        \ML_int[2][87] ) );
  MUX2_X2 M1_1_86 ( .A(\ML_int[1][86] ), .B(\ML_int[1][84] ), .S(n13), .Z(
        \ML_int[2][86] ) );
  MUX2_X2 M1_1_85 ( .A(\ML_int[1][85] ), .B(\ML_int[1][83] ), .S(n12), .Z(
        \ML_int[2][85] ) );
  MUX2_X2 M1_1_84 ( .A(\ML_int[1][84] ), .B(\ML_int[1][82] ), .S(n11), .Z(
        \ML_int[2][84] ) );
  MUX2_X2 M1_1_83 ( .A(\ML_int[1][83] ), .B(\ML_int[1][81] ), .S(n11), .Z(
        \ML_int[2][83] ) );
  MUX2_X2 M1_1_82 ( .A(\ML_int[1][82] ), .B(\ML_int[1][80] ), .S(n11), .Z(
        \ML_int[2][82] ) );
  MUX2_X2 M1_1_81 ( .A(\ML_int[1][81] ), .B(\ML_int[1][79] ), .S(n11), .Z(
        \ML_int[2][81] ) );
  MUX2_X2 M1_1_80 ( .A(\ML_int[1][80] ), .B(\ML_int[1][78] ), .S(n11), .Z(
        \ML_int[2][80] ) );
  MUX2_X2 M1_1_79 ( .A(\ML_int[1][79] ), .B(\ML_int[1][77] ), .S(n11), .Z(
        \ML_int[2][79] ) );
  MUX2_X2 M1_1_78 ( .A(\ML_int[1][78] ), .B(\ML_int[1][76] ), .S(n11), .Z(
        \ML_int[2][78] ) );
  MUX2_X2 M1_1_77 ( .A(\ML_int[1][77] ), .B(\ML_int[1][75] ), .S(n11), .Z(
        \ML_int[2][77] ) );
  MUX2_X2 M1_1_76 ( .A(\ML_int[1][76] ), .B(\ML_int[1][74] ), .S(n11), .Z(
        \ML_int[2][76] ) );
  MUX2_X2 M1_1_75 ( .A(\ML_int[1][75] ), .B(\ML_int[1][73] ), .S(n11), .Z(
        \ML_int[2][75] ) );
  MUX2_X2 M1_1_74 ( .A(\ML_int[1][74] ), .B(\ML_int[1][72] ), .S(n11), .Z(
        \ML_int[2][74] ) );
  MUX2_X2 M1_1_73 ( .A(\ML_int[1][73] ), .B(\ML_int[1][71] ), .S(n11), .Z(
        \ML_int[2][73] ) );
  MUX2_X2 M1_1_72 ( .A(\ML_int[1][72] ), .B(\ML_int[1][70] ), .S(n11), .Z(
        \ML_int[2][72] ) );
  MUX2_X2 M1_1_71 ( .A(\ML_int[1][71] ), .B(\ML_int[1][69] ), .S(n11), .Z(
        \ML_int[2][71] ) );
  MUX2_X2 M1_1_70 ( .A(\ML_int[1][70] ), .B(\ML_int[1][68] ), .S(n12), .Z(
        \ML_int[2][70] ) );
  MUX2_X2 M1_1_69 ( .A(\ML_int[1][69] ), .B(\ML_int[1][67] ), .S(n12), .Z(
        \ML_int[2][69] ) );
  MUX2_X2 M1_1_68 ( .A(\ML_int[1][68] ), .B(\ML_int[1][66] ), .S(n12), .Z(
        \ML_int[2][68] ) );
  MUX2_X2 M1_1_67 ( .A(\ML_int[1][67] ), .B(\ML_int[1][65] ), .S(n10), .Z(
        \ML_int[2][67] ) );
  MUX2_X2 M1_1_66 ( .A(\ML_int[1][66] ), .B(\ML_int[1][64] ), .S(n11), .Z(
        \ML_int[2][66] ) );
  MUX2_X2 M1_1_65 ( .A(\ML_int[1][65] ), .B(\ML_int[1][63] ), .S(n11), .Z(
        \ML_int[2][65] ) );
  MUX2_X2 M1_1_64 ( .A(\ML_int[1][64] ), .B(\ML_int[1][62] ), .S(n11), .Z(
        \ML_int[2][64] ) );
  MUX2_X2 M1_1_63 ( .A(\ML_int[1][63] ), .B(\ML_int[1][61] ), .S(n11), .Z(
        \ML_int[2][63] ) );
  MUX2_X2 M1_1_62 ( .A(\ML_int[1][62] ), .B(\ML_int[1][60] ), .S(n11), .Z(
        \ML_int[2][62] ) );
  MUX2_X2 M1_1_61 ( .A(\ML_int[1][61] ), .B(\ML_int[1][59] ), .S(n11), .Z(
        \ML_int[2][61] ) );
  MUX2_X2 M1_1_60 ( .A(\ML_int[1][60] ), .B(\ML_int[1][58] ), .S(n11), .Z(
        \ML_int[2][60] ) );
  MUX2_X2 M1_1_59 ( .A(\ML_int[1][59] ), .B(\ML_int[1][57] ), .S(n11), .Z(
        \ML_int[2][59] ) );
  MUX2_X2 M1_1_58 ( .A(\ML_int[1][58] ), .B(\ML_int[1][56] ), .S(n11), .Z(
        \ML_int[2][58] ) );
  MUX2_X2 M1_1_57 ( .A(\ML_int[1][57] ), .B(\ML_int[1][55] ), .S(n11), .Z(
        \ML_int[2][57] ) );
  MUX2_X2 M1_1_56 ( .A(\ML_int[1][56] ), .B(\ML_int[1][54] ), .S(n10), .Z(
        \ML_int[2][56] ) );
  MUX2_X2 M1_1_55 ( .A(\ML_int[1][55] ), .B(\ML_int[1][53] ), .S(n10), .Z(
        \ML_int[2][55] ) );
  MUX2_X2 M1_1_54 ( .A(\ML_int[1][54] ), .B(\ML_int[1][52] ), .S(n10), .Z(
        \ML_int[2][54] ) );
  MUX2_X2 M1_1_53 ( .A(\ML_int[1][53] ), .B(\ML_int[1][51] ), .S(n10), .Z(
        \ML_int[2][53] ) );
  MUX2_X2 M1_1_52 ( .A(\ML_int[1][52] ), .B(\ML_int[1][50] ), .S(n10), .Z(
        \ML_int[2][52] ) );
  MUX2_X2 M1_1_51 ( .A(\ML_int[1][51] ), .B(\ML_int[1][49] ), .S(n10), .Z(
        \ML_int[2][51] ) );
  MUX2_X2 M1_1_50 ( .A(\ML_int[1][50] ), .B(\ML_int[1][48] ), .S(n10), .Z(
        \ML_int[2][50] ) );
  MUX2_X2 M1_1_49 ( .A(\ML_int[1][49] ), .B(\ML_int[1][47] ), .S(n10), .Z(
        \ML_int[2][49] ) );
  MUX2_X2 M1_1_48 ( .A(\ML_int[1][48] ), .B(\ML_int[1][46] ), .S(n10), .Z(
        \ML_int[2][48] ) );
  MUX2_X2 M1_1_47 ( .A(\ML_int[1][47] ), .B(\ML_int[1][45] ), .S(n10), .Z(
        \ML_int[2][47] ) );
  MUX2_X2 M1_1_46 ( .A(\ML_int[1][46] ), .B(\ML_int[1][44] ), .S(n10), .Z(
        \ML_int[2][46] ) );
  MUX2_X2 M1_1_45 ( .A(\ML_int[1][45] ), .B(\ML_int[1][43] ), .S(n13), .Z(
        \ML_int[2][45] ) );
  MUX2_X2 M1_1_44 ( .A(\ML_int[1][44] ), .B(\ML_int[1][42] ), .S(n13), .Z(
        \ML_int[2][44] ) );
  MUX2_X2 M1_1_43 ( .A(\ML_int[1][43] ), .B(\ML_int[1][41] ), .S(n13), .Z(
        \ML_int[2][43] ) );
  MUX2_X2 M1_1_42 ( .A(\ML_int[1][42] ), .B(\ML_int[1][40] ), .S(n13), .Z(
        \ML_int[2][42] ) );
  MUX2_X2 M1_1_41 ( .A(\ML_int[1][41] ), .B(\ML_int[1][39] ), .S(n13), .Z(
        \ML_int[2][41] ) );
  MUX2_X2 M1_1_40 ( .A(\ML_int[1][40] ), .B(\ML_int[1][38] ), .S(n13), .Z(
        \ML_int[2][40] ) );
  MUX2_X2 M1_1_39 ( .A(\ML_int[1][39] ), .B(\ML_int[1][37] ), .S(n13), .Z(
        \ML_int[2][39] ) );
  MUX2_X2 M1_1_38 ( .A(\ML_int[1][38] ), .B(\ML_int[1][36] ), .S(n13), .Z(
        \ML_int[2][38] ) );
  MUX2_X2 M1_1_37 ( .A(\ML_int[1][37] ), .B(\ML_int[1][35] ), .S(n13), .Z(
        \ML_int[2][37] ) );
  MUX2_X2 M1_1_36 ( .A(\ML_int[1][36] ), .B(\ML_int[1][34] ), .S(n13), .Z(
        \ML_int[2][36] ) );
  MUX2_X2 M1_1_35 ( .A(\ML_int[1][35] ), .B(\ML_int[1][33] ), .S(n13), .Z(
        \ML_int[2][35] ) );
  MUX2_X2 M1_1_34 ( .A(\ML_int[1][34] ), .B(\ML_int[1][32] ), .S(n12), .Z(
        \ML_int[2][34] ) );
  MUX2_X2 M1_1_33 ( .A(\ML_int[1][33] ), .B(\ML_int[1][31] ), .S(n12), .Z(
        \ML_int[2][33] ) );
  MUX2_X2 M1_1_32 ( .A(\ML_int[1][32] ), .B(\ML_int[1][30] ), .S(n12), .Z(
        \ML_int[2][32] ) );
  MUX2_X2 M1_1_31 ( .A(\ML_int[1][31] ), .B(\ML_int[1][29] ), .S(n12), .Z(
        \ML_int[2][31] ) );
  MUX2_X2 M1_1_30 ( .A(\ML_int[1][30] ), .B(\ML_int[1][28] ), .S(n13), .Z(
        \ML_int[2][30] ) );
  MUX2_X2 M1_1_29 ( .A(\ML_int[1][29] ), .B(\ML_int[1][27] ), .S(n13), .Z(
        \ML_int[2][29] ) );
  MUX2_X2 M1_1_28 ( .A(\ML_int[1][28] ), .B(\ML_int[1][26] ), .S(n13), .Z(
        \ML_int[2][28] ) );
  MUX2_X2 M1_1_27 ( .A(\ML_int[1][27] ), .B(\ML_int[1][25] ), .S(n13), .Z(
        \ML_int[2][27] ) );
  MUX2_X2 M1_1_26 ( .A(\ML_int[1][26] ), .B(\ML_int[1][24] ), .S(n13), .Z(
        \ML_int[2][26] ) );
  MUX2_X2 M1_1_25 ( .A(\ML_int[1][25] ), .B(\ML_int[1][23] ), .S(n13), .Z(
        \ML_int[2][25] ) );
  MUX2_X2 M1_1_24 ( .A(\ML_int[1][24] ), .B(\ML_int[1][22] ), .S(n13), .Z(
        \ML_int[2][24] ) );
  MUX2_X2 M1_1_23 ( .A(\ML_int[1][23] ), .B(\ML_int[1][21] ), .S(n12), .Z(
        \ML_int[2][23] ) );
  MUX2_X2 M1_1_22 ( .A(\ML_int[1][22] ), .B(\ML_int[1][20] ), .S(n12), .Z(
        \ML_int[2][22] ) );
  MUX2_X2 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S(n12), .Z(
        \ML_int[2][21] ) );
  MUX2_X2 M1_1_20 ( .A(\ML_int[1][20] ), .B(\ML_int[1][18] ), .S(n12), .Z(
        \ML_int[2][20] ) );
  MUX2_X2 M1_1_19 ( .A(\ML_int[1][19] ), .B(\ML_int[1][17] ), .S(n12), .Z(
        \ML_int[2][19] ) );
  MUX2_X2 M1_1_18 ( .A(\ML_int[1][18] ), .B(\ML_int[1][16] ), .S(n12), .Z(
        \ML_int[2][18] ) );
  MUX2_X2 M1_1_17 ( .A(\ML_int[1][17] ), .B(\ML_int[1][15] ), .S(n12), .Z(
        \ML_int[2][17] ) );
  MUX2_X2 M1_1_16 ( .A(\ML_int[1][16] ), .B(\ML_int[1][14] ), .S(n12), .Z(
        \ML_int[2][16] ) );
  MUX2_X2 M1_1_15 ( .A(\ML_int[1][15] ), .B(\ML_int[1][13] ), .S(n12), .Z(
        \ML_int[2][15] ) );
  MUX2_X2 M1_1_14 ( .A(\ML_int[1][14] ), .B(\ML_int[1][12] ), .S(n12), .Z(
        \ML_int[2][14] ) );
  MUX2_X2 M1_1_13 ( .A(\ML_int[1][13] ), .B(\ML_int[1][11] ), .S(n12), .Z(
        \ML_int[2][13] ) );
  MUX2_X2 M1_1_12 ( .A(\ML_int[1][12] ), .B(\ML_int[1][10] ), .S(n10), .Z(
        \ML_int[2][12] ) );
  MUX2_X2 M1_1_11 ( .A(\ML_int[1][11] ), .B(\ML_int[1][9] ), .S(n10), .Z(
        \ML_int[2][11] ) );
  MUX2_X2 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S(n12), .Z(
        \ML_int[2][10] ) );
  MUX2_X2 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S(n12), .Z(
        \ML_int[2][9] ) );
  MUX2_X2 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S(n12), .Z(
        \ML_int[2][8] ) );
  MUX2_X2 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S(n10), .Z(
        \ML_int[2][7] ) );
  MUX2_X2 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S(n10), .Z(
        \ML_int[2][6] ) );
  MUX2_X2 M1_1_5 ( .A(\ML_int[1][5] ), .B(\ML_int[1][3] ), .S(n12), .Z(
        \ML_int[2][5] ) );
  MUX2_X2 M1_1_4 ( .A(\ML_int[1][4] ), .B(\ML_int[1][2] ), .S(n12), .Z(
        \ML_int[2][4] ) );
  MUX2_X2 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(n10), .Z(
        \ML_int[2][3] ) );
  MUX2_X2 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S(n10), .Z(
        \ML_int[2][2] ) );
  MUX2_X2 M1_0_105 ( .A(A[105]), .B(A[104]), .S(n8), .Z(\ML_int[1][105] ) );
  MUX2_X2 M1_0_104 ( .A(A[104]), .B(A[103]), .S(n8), .Z(\ML_int[1][104] ) );
  MUX2_X2 M1_0_103 ( .A(A[103]), .B(A[102]), .S(n8), .Z(\ML_int[1][103] ) );
  MUX2_X2 M1_0_102 ( .A(A[102]), .B(A[101]), .S(n8), .Z(\ML_int[1][102] ) );
  MUX2_X2 M1_0_101 ( .A(A[101]), .B(A[100]), .S(n8), .Z(\ML_int[1][101] ) );
  MUX2_X2 M1_0_100 ( .A(A[100]), .B(A[99]), .S(n8), .Z(\ML_int[1][100] ) );
  MUX2_X2 M1_0_99 ( .A(A[99]), .B(A[98]), .S(n8), .Z(\ML_int[1][99] ) );
  MUX2_X2 M1_0_98 ( .A(A[98]), .B(A[97]), .S(n8), .Z(\ML_int[1][98] ) );
  MUX2_X2 M1_0_97 ( .A(A[97]), .B(A[96]), .S(n8), .Z(\ML_int[1][97] ) );
  MUX2_X2 M1_0_96 ( .A(A[96]), .B(A[95]), .S(n8), .Z(\ML_int[1][96] ) );
  MUX2_X2 M1_0_95 ( .A(A[95]), .B(A[94]), .S(n8), .Z(\ML_int[1][95] ) );
  MUX2_X2 M1_0_94 ( .A(A[94]), .B(A[93]), .S(n8), .Z(\ML_int[1][94] ) );
  MUX2_X2 M1_0_93 ( .A(A[93]), .B(A[92]), .S(n8), .Z(\ML_int[1][93] ) );
  MUX2_X2 M1_0_92 ( .A(A[92]), .B(A[91]), .S(n8), .Z(\ML_int[1][92] ) );
  MUX2_X2 M1_0_91 ( .A(A[91]), .B(A[90]), .S(n8), .Z(\ML_int[1][91] ) );
  MUX2_X2 M1_0_90 ( .A(A[90]), .B(A[89]), .S(n8), .Z(\ML_int[1][90] ) );
  MUX2_X2 M1_0_89 ( .A(A[89]), .B(A[88]), .S(n8), .Z(\ML_int[1][89] ) );
  MUX2_X2 M1_0_88 ( .A(A[88]), .B(A[87]), .S(n6), .Z(\ML_int[1][88] ) );
  MUX2_X2 M1_0_87 ( .A(A[87]), .B(A[86]), .S(n6), .Z(\ML_int[1][87] ) );
  MUX2_X2 M1_0_86 ( .A(A[86]), .B(A[85]), .S(n6), .Z(\ML_int[1][86] ) );
  MUX2_X2 M1_0_85 ( .A(A[85]), .B(A[84]), .S(n6), .Z(\ML_int[1][85] ) );
  MUX2_X2 M1_0_84 ( .A(A[84]), .B(A[83]), .S(n6), .Z(\ML_int[1][84] ) );
  MUX2_X2 M1_0_83 ( .A(A[83]), .B(A[82]), .S(n6), .Z(\ML_int[1][83] ) );
  MUX2_X2 M1_0_82 ( .A(A[82]), .B(A[81]), .S(n6), .Z(\ML_int[1][82] ) );
  MUX2_X2 M1_0_81 ( .A(A[81]), .B(A[80]), .S(n8), .Z(\ML_int[1][81] ) );
  MUX2_X2 M1_0_80 ( .A(A[80]), .B(A[79]), .S(n8), .Z(\ML_int[1][80] ) );
  MUX2_X2 M1_0_79 ( .A(A[79]), .B(A[78]), .S(n8), .Z(\ML_int[1][79] ) );
  MUX2_X2 M1_0_78 ( .A(A[78]), .B(A[77]), .S(n8), .Z(\ML_int[1][78] ) );
  MUX2_X2 M1_0_77 ( .A(A[77]), .B(A[76]), .S(n8), .Z(\ML_int[1][77] ) );
  MUX2_X2 M1_0_76 ( .A(A[76]), .B(A[75]), .S(n8), .Z(\ML_int[1][76] ) );
  MUX2_X2 M1_0_75 ( .A(A[75]), .B(A[74]), .S(n8), .Z(\ML_int[1][75] ) );
  MUX2_X2 M1_0_74 ( .A(A[74]), .B(A[73]), .S(n8), .Z(\ML_int[1][74] ) );
  MUX2_X2 M1_0_73 ( .A(A[73]), .B(A[72]), .S(n8), .Z(\ML_int[1][73] ) );
  MUX2_X2 M1_0_72 ( .A(A[72]), .B(A[71]), .S(n8), .Z(\ML_int[1][72] ) );
  MUX2_X2 M1_0_71 ( .A(A[71]), .B(A[70]), .S(n8), .Z(\ML_int[1][71] ) );
  MUX2_X2 M1_0_70 ( .A(A[70]), .B(A[69]), .S(n8), .Z(\ML_int[1][70] ) );
  MUX2_X2 M1_0_69 ( .A(A[69]), .B(A[68]), .S(n9), .Z(\ML_int[1][69] ) );
  MUX2_X2 M1_0_68 ( .A(A[68]), .B(A[67]), .S(n9), .Z(\ML_int[1][68] ) );
  MUX2_X2 M1_0_67 ( .A(A[67]), .B(A[66]), .S(n9), .Z(\ML_int[1][67] ) );
  MUX2_X2 M1_0_66 ( .A(A[66]), .B(A[65]), .S(n7), .Z(\ML_int[1][66] ) );
  MUX2_X2 M1_0_65 ( .A(A[65]), .B(A[64]), .S(n8), .Z(\ML_int[1][65] ) );
  MUX2_X2 M1_0_64 ( .A(A[64]), .B(A[63]), .S(n8), .Z(\ML_int[1][64] ) );
  MUX2_X2 M1_0_63 ( .A(A[63]), .B(A[62]), .S(n8), .Z(\ML_int[1][63] ) );
  MUX2_X2 M1_0_62 ( .A(A[62]), .B(A[61]), .S(n8), .Z(\ML_int[1][62] ) );
  MUX2_X2 M1_0_61 ( .A(A[61]), .B(A[60]), .S(n8), .Z(\ML_int[1][61] ) );
  MUX2_X2 M1_0_60 ( .A(A[60]), .B(A[59]), .S(n8), .Z(\ML_int[1][60] ) );
  MUX2_X2 M1_0_59 ( .A(A[59]), .B(A[58]), .S(n8), .Z(\ML_int[1][59] ) );
  MUX2_X2 M1_0_58 ( .A(A[58]), .B(A[57]), .S(n8), .Z(\ML_int[1][58] ) );
  MUX2_X2 M1_0_57 ( .A(A[57]), .B(A[56]), .S(n8), .Z(\ML_int[1][57] ) );
  MUX2_X2 M1_0_56 ( .A(A[56]), .B(A[55]), .S(n8), .Z(\ML_int[1][56] ) );
  MUX2_X2 M1_0_55 ( .A(A[55]), .B(A[54]), .S(n7), .Z(\ML_int[1][55] ) );
  MUX2_X2 M1_0_54 ( .A(A[54]), .B(A[53]), .S(n7), .Z(\ML_int[1][54] ) );
  MUX2_X2 M1_0_53 ( .A(A[53]), .B(A[52]), .S(n7), .Z(\ML_int[1][53] ) );
  MUX2_X2 M1_0_52 ( .A(A[52]), .B(A[51]), .S(n7), .Z(\ML_int[1][52] ) );
  MUX2_X2 M1_0_51 ( .A(A[51]), .B(A[50]), .S(n7), .Z(\ML_int[1][51] ) );
  MUX2_X2 M1_0_50 ( .A(A[50]), .B(A[49]), .S(n7), .Z(\ML_int[1][50] ) );
  MUX2_X2 M1_0_49 ( .A(A[49]), .B(A[48]), .S(n7), .Z(\ML_int[1][49] ) );
  MUX2_X2 M1_0_48 ( .A(A[48]), .B(A[47]), .S(n7), .Z(\ML_int[1][48] ) );
  MUX2_X2 M1_0_47 ( .A(A[47]), .B(A[46]), .S(n7), .Z(\ML_int[1][47] ) );
  MUX2_X2 M1_0_46 ( .A(A[46]), .B(A[45]), .S(n7), .Z(\ML_int[1][46] ) );
  MUX2_X2 M1_0_45 ( .A(A[45]), .B(A[44]), .S(n7), .Z(\ML_int[1][45] ) );
  MUX2_X2 M1_0_44 ( .A(A[44]), .B(A[43]), .S(n9), .Z(\ML_int[1][44] ) );
  MUX2_X2 M1_0_43 ( .A(A[43]), .B(A[42]), .S(n9), .Z(\ML_int[1][43] ) );
  MUX2_X2 M1_0_42 ( .A(A[42]), .B(A[41]), .S(n9), .Z(\ML_int[1][42] ) );
  MUX2_X2 M1_0_41 ( .A(A[41]), .B(A[40]), .S(n9), .Z(\ML_int[1][41] ) );
  MUX2_X2 M1_0_40 ( .A(A[40]), .B(A[39]), .S(n9), .Z(\ML_int[1][40] ) );
  MUX2_X2 M1_0_39 ( .A(A[39]), .B(A[38]), .S(n9), .Z(\ML_int[1][39] ) );
  MUX2_X2 M1_0_38 ( .A(A[38]), .B(A[37]), .S(n9), .Z(\ML_int[1][38] ) );
  MUX2_X2 M1_0_37 ( .A(A[37]), .B(A[36]), .S(n9), .Z(\ML_int[1][37] ) );
  MUX2_X2 M1_0_36 ( .A(A[36]), .B(A[35]), .S(n9), .Z(\ML_int[1][36] ) );
  MUX2_X2 M1_0_35 ( .A(A[35]), .B(A[34]), .S(n9), .Z(\ML_int[1][35] ) );
  MUX2_X2 M1_0_34 ( .A(A[34]), .B(A[33]), .S(n9), .Z(\ML_int[1][34] ) );
  MUX2_X2 M1_0_33 ( .A(A[33]), .B(A[32]), .S(n9), .Z(\ML_int[1][33] ) );
  MUX2_X2 M1_0_32 ( .A(A[32]), .B(A[31]), .S(n9), .Z(\ML_int[1][32] ) );
  MUX2_X2 M1_0_31 ( .A(A[31]), .B(A[30]), .S(n9), .Z(\ML_int[1][31] ) );
  MUX2_X2 M1_0_30 ( .A(A[30]), .B(A[29]), .S(n9), .Z(\ML_int[1][30] ) );
  MUX2_X2 M1_0_29 ( .A(A[29]), .B(A[28]), .S(n9), .Z(\ML_int[1][29] ) );
  MUX2_X2 M1_0_28 ( .A(A[28]), .B(A[27]), .S(n9), .Z(\ML_int[1][28] ) );
  MUX2_X2 M1_0_27 ( .A(A[27]), .B(A[26]), .S(n9), .Z(\ML_int[1][27] ) );
  MUX2_X2 M1_0_26 ( .A(A[26]), .B(A[25]), .S(n9), .Z(\ML_int[1][26] ) );
  MUX2_X2 M1_0_25 ( .A(A[25]), .B(A[24]), .S(n9), .Z(\ML_int[1][25] ) );
  MUX2_X2 M1_0_24 ( .A(A[24]), .B(A[23]), .S(n9), .Z(\ML_int[1][24] ) );
  MUX2_X2 M1_0_23 ( .A(A[23]), .B(A[22]), .S(n9), .Z(\ML_int[1][23] ) );
  MUX2_X2 M1_0_22 ( .A(A[22]), .B(A[21]), .S(n9), .Z(\ML_int[1][22] ) );
  MUX2_X2 M1_0_21 ( .A(A[21]), .B(A[20]), .S(n9), .Z(\ML_int[1][21] ) );
  MUX2_X2 M1_0_20 ( .A(A[20]), .B(A[19]), .S(n9), .Z(\ML_int[1][20] ) );
  MUX2_X2 M1_0_19 ( .A(A[19]), .B(A[18]), .S(n9), .Z(\ML_int[1][19] ) );
  MUX2_X2 M1_0_18 ( .A(A[18]), .B(A[17]), .S(n9), .Z(\ML_int[1][18] ) );
  MUX2_X2 M1_0_17 ( .A(A[17]), .B(A[16]), .S(n9), .Z(\ML_int[1][17] ) );
  MUX2_X2 M1_0_16 ( .A(A[16]), .B(A[15]), .S(n9), .Z(\ML_int[1][16] ) );
  MUX2_X2 M1_0_15 ( .A(A[15]), .B(A[14]), .S(n9), .Z(\ML_int[1][15] ) );
  MUX2_X2 M1_0_14 ( .A(A[14]), .B(A[13]), .S(n9), .Z(\ML_int[1][14] ) );
  MUX2_X2 M1_0_13 ( .A(A[13]), .B(A[12]), .S(n9), .Z(\ML_int[1][13] ) );
  MUX2_X2 M1_0_12 ( .A(A[12]), .B(A[11]), .S(n9), .Z(\ML_int[1][12] ) );
  MUX2_X2 M1_0_11 ( .A(A[11]), .B(A[10]), .S(n6), .Z(\ML_int[1][11] ) );
  MUX2_X2 M1_0_10 ( .A(A[10]), .B(A[9]), .S(n7), .Z(\ML_int[1][10] ) );
  MUX2_X2 M1_0_9 ( .A(A[9]), .B(A[8]), .S(n6), .Z(\ML_int[1][9] ) );
  MUX2_X2 M1_0_8 ( .A(A[8]), .B(A[7]), .S(n6), .Z(\ML_int[1][8] ) );
  MUX2_X2 M1_0_7 ( .A(A[7]), .B(A[6]), .S(n6), .Z(\ML_int[1][7] ) );
  MUX2_X2 M1_0_6 ( .A(A[6]), .B(A[5]), .S(n6), .Z(\ML_int[1][6] ) );
  MUX2_X2 M1_0_5 ( .A(A[5]), .B(A[4]), .S(n6), .Z(\ML_int[1][5] ) );
  MUX2_X2 M1_0_4 ( .A(A[4]), .B(A[3]), .S(n6), .Z(\ML_int[1][4] ) );
  MUX2_X2 M1_0_3 ( .A(A[3]), .B(A[2]), .S(n6), .Z(\ML_int[1][3] ) );
  MUX2_X2 M1_0_2 ( .A(A[2]), .B(A[1]), .S(n6), .Z(\ML_int[1][2] ) );
  MUX2_X2 M1_0_1 ( .A(A[1]), .B(A[0]), .S(n6), .Z(\ML_int[1][1] ) );
  INV_X4 U3 ( .A(n22), .ZN(n21) );
  INV_X4 U4 ( .A(SHMAG[4]), .ZN(n36) );
  INV_X4 U5 ( .A(\temp_int_SH[5] ), .ZN(n51) );
  INV_X4 U6 ( .A(n33), .ZN(n32) );
  INV_X4 U7 ( .A(n33), .ZN(n31) );
  INV_X4 U8 ( .A(n34), .ZN(n30) );
  INV_X4 U9 ( .A(n49), .ZN(n45) );
  INV_X4 U10 ( .A(n48), .ZN(n46) );
  INV_X4 U11 ( .A(n34), .ZN(n29) );
  INV_X4 U12 ( .A(n24), .ZN(n22) );
  INV_X4 U13 ( .A(SHMAG[3]), .ZN(n24) );
  INV_X4 U14 ( .A(n22), .ZN(n20) );
  INV_X4 U15 ( .A(n23), .ZN(n19) );
  INV_X4 U16 ( .A(n42), .ZN(n41) );
  INV_X4 U17 ( .A(n28), .ZN(n26) );
  INV_X4 U18 ( .A(n50), .ZN(n49) );
  INV_X4 U19 ( .A(n48), .ZN(n47) );
  INV_X4 U20 ( .A(n51), .ZN(n50) );
  INV_X4 U21 ( .A(n36), .ZN(n34) );
  INV_X4 U22 ( .A(SHMAG[2]), .ZN(n16) );
  INV_X4 U23 ( .A(SHMAG[2]), .ZN(n17) );
  INV_X4 U24 ( .A(SHMAG[1]), .ZN(n12) );
  INV_X4 U25 ( .A(SHMAG[1]), .ZN(n13) );
  INV_X4 U26 ( .A(SHMAG[1]), .ZN(n10) );
  INV_X4 U27 ( .A(n43), .ZN(n40) );
  NOR2_X2 U28 ( .A1(n37), .A2(SH[8]), .ZN(n1) );
  INV_X4 U29 ( .A(SHMAG[0]), .ZN(n9) );
  INV_X4 U30 ( .A(n36), .ZN(n33) );
  INV_X4 U31 ( .A(n49), .ZN(n44) );
  INV_X4 U32 ( .A(n47), .ZN(n39) );
  INV_X4 U33 ( .A(SHMAG[0]), .ZN(n6) );
  INV_X4 U34 ( .A(n36), .ZN(n35) );
  INV_X4 U35 ( .A(SHMAG[2]), .ZN(n14) );
  INV_X4 U36 ( .A(SH[8]), .ZN(n2) );
  INV_X4 U37 ( .A(SH[8]), .ZN(n3) );
  INV_X4 U38 ( .A(SHMAG[0]), .ZN(n7) );
  INV_X4 U39 ( .A(SHMAG[1]), .ZN(n11) );
  INV_X4 U40 ( .A(n23), .ZN(n18) );
  INV_X4 U41 ( .A(n27), .ZN(n25) );
  INV_X4 U42 ( .A(SHMAG[6]), .ZN(n37) );
  INV_X4 U43 ( .A(SHMAG[6]), .ZN(n38) );
  INV_X4 U44 ( .A(SHMAG[0]), .ZN(n8) );
  INV_X4 U45 ( .A(n24), .ZN(n23) );
  INV_X4 U46 ( .A(n35), .ZN(n27) );
  INV_X4 U47 ( .A(n39), .ZN(n42) );
  INV_X4 U48 ( .A(SHMAG[2]), .ZN(n15) );
  INV_X4 U49 ( .A(n35), .ZN(n28) );
  INV_X4 U50 ( .A(n50), .ZN(n48) );
  INV_X4 U51 ( .A(n39), .ZN(n43) );
  INV_X4 U52 ( .A(n1), .ZN(n4) );
  INV_X4 U53 ( .A(n1), .ZN(n5) );
  NOR2_X1 U54 ( .A1(n4), .A2(n52), .ZN(B[9]) );
  AND2_X1 U55 ( .A1(\ML_int[7][99] ), .A2(n2), .ZN(B[99]) );
  AND2_X1 U56 ( .A1(\ML_int[7][98] ), .A2(n2), .ZN(B[98]) );
  AND2_X1 U57 ( .A1(\ML_int[7][97] ), .A2(n2), .ZN(B[97]) );
  AND2_X1 U58 ( .A1(\ML_int[7][96] ), .A2(n2), .ZN(B[96]) );
  AND2_X1 U59 ( .A1(\ML_int[7][95] ), .A2(n2), .ZN(B[95]) );
  AND2_X1 U60 ( .A1(\ML_int[7][94] ), .A2(n2), .ZN(B[94]) );
  AND2_X1 U61 ( .A1(\ML_int[7][93] ), .A2(n2), .ZN(B[93]) );
  AND2_X1 U62 ( .A1(\ML_int[7][92] ), .A2(n2), .ZN(B[92]) );
  AND2_X1 U63 ( .A1(\ML_int[7][91] ), .A2(n2), .ZN(B[91]) );
  AND2_X1 U64 ( .A1(\ML_int[7][90] ), .A2(n2), .ZN(B[90]) );
  NOR2_X1 U65 ( .A1(n4), .A2(n54), .ZN(B[8]) );
  AND2_X1 U66 ( .A1(\ML_int[7][89] ), .A2(n2), .ZN(B[89]) );
  AND2_X1 U67 ( .A1(\ML_int[7][88] ), .A2(n53), .ZN(B[88]) );
  AND2_X1 U68 ( .A1(\ML_int[7][87] ), .A2(n53), .ZN(B[87]) );
  AND2_X1 U69 ( .A1(\ML_int[7][86] ), .A2(n53), .ZN(B[86]) );
  AND2_X1 U70 ( .A1(\ML_int[7][85] ), .A2(n53), .ZN(B[85]) );
  AND2_X1 U71 ( .A1(\ML_int[7][84] ), .A2(n53), .ZN(B[84]) );
  AND2_X1 U72 ( .A1(\ML_int[7][83] ), .A2(n53), .ZN(B[83]) );
  AND2_X1 U73 ( .A1(\ML_int[7][82] ), .A2(n53), .ZN(B[82]) );
  AND2_X1 U74 ( .A1(\ML_int[7][81] ), .A2(n53), .ZN(B[81]) );
  AND2_X1 U75 ( .A1(\ML_int[7][80] ), .A2(n53), .ZN(B[80]) );
  NOR2_X1 U76 ( .A1(n5), .A2(n55), .ZN(B[7]) );
  AND2_X1 U77 ( .A1(\ML_int[7][79] ), .A2(n53), .ZN(B[79]) );
  AND2_X1 U78 ( .A1(\ML_int[7][78] ), .A2(n53), .ZN(B[78]) );
  AND2_X1 U79 ( .A1(\ML_int[7][77] ), .A2(n53), .ZN(B[77]) );
  AND2_X1 U80 ( .A1(\ML_int[7][76] ), .A2(n53), .ZN(B[76]) );
  AND2_X1 U81 ( .A1(\ML_int[7][75] ), .A2(n53), .ZN(B[75]) );
  AND2_X1 U82 ( .A1(\ML_int[7][74] ), .A2(n53), .ZN(B[74]) );
  AND2_X1 U83 ( .A1(\ML_int[7][73] ), .A2(n53), .ZN(B[73]) );
  AND2_X1 U84 ( .A1(\ML_int[7][72] ), .A2(n53), .ZN(B[72]) );
  AND2_X1 U85 ( .A1(\ML_int[7][71] ), .A2(n53), .ZN(B[71]) );
  AND2_X1 U86 ( .A1(\ML_int[7][70] ), .A2(n53), .ZN(B[70]) );
  NOR2_X1 U87 ( .A1(n4), .A2(n56), .ZN(B[6]) );
  AND2_X1 U88 ( .A1(\ML_int[7][69] ), .A2(n2), .ZN(B[69]) );
  AND2_X1 U89 ( .A1(\ML_int[7][68] ), .A2(n2), .ZN(B[68]) );
  AND2_X1 U90 ( .A1(\ML_int[7][67] ), .A2(n3), .ZN(B[67]) );
  AND2_X1 U91 ( .A1(\ML_int[7][66] ), .A2(n3), .ZN(B[66]) );
  AND2_X1 U92 ( .A1(\ML_int[7][65] ), .A2(n3), .ZN(B[65]) );
  AND2_X1 U93 ( .A1(\ML_int[7][64] ), .A2(n3), .ZN(B[64]) );
  AND2_X1 U94 ( .A1(\ML_int[6][63] ), .A2(n1), .ZN(B[63]) );
  AND2_X1 U95 ( .A1(\ML_int[6][62] ), .A2(n1), .ZN(B[62]) );
  AND2_X1 U96 ( .A1(\ML_int[6][61] ), .A2(n1), .ZN(B[61]) );
  AND2_X1 U97 ( .A1(\ML_int[6][60] ), .A2(n1), .ZN(B[60]) );
  NOR2_X1 U98 ( .A1(n4), .A2(n57), .ZN(B[5]) );
  AND2_X1 U99 ( .A1(\ML_int[6][59] ), .A2(n1), .ZN(B[59]) );
  AND2_X1 U100 ( .A1(\ML_int[6][58] ), .A2(n1), .ZN(B[58]) );
  AND2_X1 U101 ( .A1(\ML_int[6][57] ), .A2(n1), .ZN(B[57]) );
  AND2_X1 U102 ( .A1(\ML_int[6][56] ), .A2(n1), .ZN(B[56]) );
  AND2_X1 U103 ( .A1(\ML_int[6][55] ), .A2(n1), .ZN(B[55]) );
  AND2_X1 U104 ( .A1(\ML_int[6][54] ), .A2(n1), .ZN(B[54]) );
  AND2_X1 U105 ( .A1(\ML_int[6][53] ), .A2(n1), .ZN(B[53]) );
  AND2_X1 U106 ( .A1(\ML_int[6][52] ), .A2(n1), .ZN(B[52]) );
  AND2_X1 U107 ( .A1(\ML_int[6][51] ), .A2(n1), .ZN(B[51]) );
  AND2_X1 U108 ( .A1(\ML_int[6][50] ), .A2(n1), .ZN(B[50]) );
  NOR2_X1 U109 ( .A1(n4), .A2(n58), .ZN(B[4]) );
  AND2_X1 U110 ( .A1(\ML_int[6][49] ), .A2(n1), .ZN(B[49]) );
  AND2_X1 U111 ( .A1(\ML_int[6][48] ), .A2(n1), .ZN(B[48]) );
  AND2_X1 U112 ( .A1(\ML_int[6][47] ), .A2(n1), .ZN(B[47]) );
  AND2_X1 U113 ( .A1(\ML_int[6][46] ), .A2(n1), .ZN(B[46]) );
  AND2_X1 U114 ( .A1(\ML_int[6][45] ), .A2(n1), .ZN(B[45]) );
  AND2_X1 U115 ( .A1(\ML_int[6][44] ), .A2(n1), .ZN(B[44]) );
  AND2_X1 U116 ( .A1(\ML_int[6][43] ), .A2(n1), .ZN(B[43]) );
  AND2_X1 U117 ( .A1(\ML_int[6][42] ), .A2(n1), .ZN(B[42]) );
  AND2_X1 U118 ( .A1(\ML_int[6][41] ), .A2(n1), .ZN(B[41]) );
  AND2_X1 U119 ( .A1(\ML_int[6][40] ), .A2(n1), .ZN(B[40]) );
  NOR2_X1 U120 ( .A1(n4), .A2(n59), .ZN(B[3]) );
  AND2_X1 U121 ( .A1(\ML_int[6][39] ), .A2(n1), .ZN(B[39]) );
  AND2_X1 U122 ( .A1(\ML_int[6][38] ), .A2(n1), .ZN(B[38]) );
  AND2_X1 U123 ( .A1(\ML_int[6][37] ), .A2(n1), .ZN(B[37]) );
  AND2_X1 U124 ( .A1(\ML_int[6][36] ), .A2(n1), .ZN(B[36]) );
  AND2_X1 U125 ( .A1(\ML_int[6][35] ), .A2(n1), .ZN(B[35]) );
  AND2_X1 U126 ( .A1(\ML_int[6][34] ), .A2(n1), .ZN(B[34]) );
  AND2_X1 U127 ( .A1(\ML_int[6][33] ), .A2(n1), .ZN(B[33]) );
  AND2_X1 U128 ( .A1(\ML_int[6][32] ), .A2(n1), .ZN(B[32]) );
  NOR2_X1 U129 ( .A1(n5), .A2(n60), .ZN(B[31]) );
  NOR2_X1 U130 ( .A1(n4), .A2(n61), .ZN(B[30]) );
  NOR2_X1 U131 ( .A1(n4), .A2(n62), .ZN(B[2]) );
  NOR2_X1 U132 ( .A1(n5), .A2(n63), .ZN(B[29]) );
  NOR2_X1 U133 ( .A1(n5), .A2(n64), .ZN(B[28]) );
  NOR2_X1 U134 ( .A1(n5), .A2(n65), .ZN(B[27]) );
  NOR2_X1 U135 ( .A1(n5), .A2(n66), .ZN(B[26]) );
  NOR2_X1 U136 ( .A1(n5), .A2(n67), .ZN(B[25]) );
  NOR2_X1 U137 ( .A1(n5), .A2(n68), .ZN(B[24]) );
  NOR2_X1 U138 ( .A1(n5), .A2(n69), .ZN(B[23]) );
  NOR2_X1 U139 ( .A1(n5), .A2(n70), .ZN(B[22]) );
  NOR2_X1 U140 ( .A1(n5), .A2(n71), .ZN(B[21]) );
  NOR2_X1 U141 ( .A1(n5), .A2(n72), .ZN(B[20]) );
  NOR2_X1 U142 ( .A1(n5), .A2(n73), .ZN(B[1]) );
  NOR2_X1 U143 ( .A1(n4), .A2(n74), .ZN(B[19]) );
  NOR2_X1 U144 ( .A1(n4), .A2(n75), .ZN(B[18]) );
  NOR2_X1 U145 ( .A1(n4), .A2(n76), .ZN(B[17]) );
  NOR2_X1 U146 ( .A1(n4), .A2(n77), .ZN(B[16]) );
  NOR2_X1 U147 ( .A1(n4), .A2(n78), .ZN(B[15]) );
  NOR2_X1 U148 ( .A1(n4), .A2(n79), .ZN(B[14]) );
  NOR2_X1 U149 ( .A1(n4), .A2(n80), .ZN(B[13]) );
  NOR2_X1 U150 ( .A1(n4), .A2(n81), .ZN(B[12]) );
  NOR2_X1 U151 ( .A1(n4), .A2(n82), .ZN(B[11]) );
  NOR2_X1 U152 ( .A1(n4), .A2(n83), .ZN(B[10]) );
  AND2_X1 U153 ( .A1(\ML_int[7][105] ), .A2(n3), .ZN(B[105]) );
  AND2_X1 U154 ( .A1(\ML_int[7][104] ), .A2(n3), .ZN(B[104]) );
  AND2_X1 U155 ( .A1(\ML_int[7][103] ), .A2(n3), .ZN(B[103]) );
  AND2_X1 U156 ( .A1(\ML_int[7][102] ), .A2(n3), .ZN(B[102]) );
  AND2_X1 U157 ( .A1(\ML_int[7][101] ), .A2(n3), .ZN(B[101]) );
  AND2_X1 U158 ( .A1(\ML_int[7][100] ), .A2(n3), .ZN(B[100]) );
  NOR2_X1 U159 ( .A1(n4), .A2(n84), .ZN(B[0]) );
  AOI21_X1 U160 ( .B1(SH[6]), .B2(n85), .A(n86), .ZN(SHMAG[6]) );
  INV_X1 U161 ( .A(n52), .ZN(\ML_int[6][9] ) );
  NAND2_X1 U162 ( .A1(\ML_int[5][9] ), .A2(n41), .ZN(n52) );
  INV_X1 U163 ( .A(n54), .ZN(\ML_int[6][8] ) );
  NAND2_X1 U164 ( .A1(\ML_int[5][8] ), .A2(n41), .ZN(n54) );
  INV_X1 U165 ( .A(n55), .ZN(\ML_int[6][7] ) );
  NAND2_X1 U166 ( .A1(\ML_int[5][7] ), .A2(n41), .ZN(n55) );
  INV_X1 U167 ( .A(n56), .ZN(\ML_int[6][6] ) );
  NAND2_X1 U168 ( .A1(\ML_int[5][6] ), .A2(n41), .ZN(n56) );
  INV_X1 U169 ( .A(n57), .ZN(\ML_int[6][5] ) );
  NAND2_X1 U170 ( .A1(\ML_int[5][5] ), .A2(n41), .ZN(n57) );
  INV_X1 U171 ( .A(n58), .ZN(\ML_int[6][4] ) );
  NAND2_X1 U172 ( .A1(\ML_int[5][4] ), .A2(n41), .ZN(n58) );
  INV_X1 U173 ( .A(n59), .ZN(\ML_int[6][3] ) );
  NAND2_X1 U174 ( .A1(\ML_int[5][3] ), .A2(n41), .ZN(n59) );
  INV_X1 U175 ( .A(n60), .ZN(\ML_int[6][31] ) );
  NAND2_X1 U176 ( .A1(\ML_int[5][31] ), .A2(n41), .ZN(n60) );
  INV_X1 U177 ( .A(n61), .ZN(\ML_int[6][30] ) );
  NAND2_X1 U178 ( .A1(\ML_int[5][30] ), .A2(n41), .ZN(n61) );
  INV_X1 U179 ( .A(n62), .ZN(\ML_int[6][2] ) );
  NAND2_X1 U180 ( .A1(\ML_int[5][2] ), .A2(n41), .ZN(n62) );
  INV_X1 U181 ( .A(n63), .ZN(\ML_int[6][29] ) );
  NAND2_X1 U182 ( .A1(\ML_int[5][29] ), .A2(n41), .ZN(n63) );
  INV_X1 U183 ( .A(n64), .ZN(\ML_int[6][28] ) );
  NAND2_X1 U184 ( .A1(\ML_int[5][28] ), .A2(n41), .ZN(n64) );
  INV_X1 U185 ( .A(n65), .ZN(\ML_int[6][27] ) );
  NAND2_X1 U186 ( .A1(\ML_int[5][27] ), .A2(n41), .ZN(n65) );
  INV_X1 U187 ( .A(n66), .ZN(\ML_int[6][26] ) );
  NAND2_X1 U188 ( .A1(\ML_int[5][26] ), .A2(n41), .ZN(n66) );
  INV_X1 U189 ( .A(n67), .ZN(\ML_int[6][25] ) );
  NAND2_X1 U190 ( .A1(\ML_int[5][25] ), .A2(n40), .ZN(n67) );
  INV_X1 U191 ( .A(n68), .ZN(\ML_int[6][24] ) );
  NAND2_X1 U192 ( .A1(\ML_int[5][24] ), .A2(n40), .ZN(n68) );
  INV_X1 U193 ( .A(n69), .ZN(\ML_int[6][23] ) );
  NAND2_X1 U194 ( .A1(\ML_int[5][23] ), .A2(n40), .ZN(n69) );
  INV_X1 U195 ( .A(n70), .ZN(\ML_int[6][22] ) );
  NAND2_X1 U196 ( .A1(\ML_int[5][22] ), .A2(n40), .ZN(n70) );
  INV_X1 U197 ( .A(n71), .ZN(\ML_int[6][21] ) );
  NAND2_X1 U198 ( .A1(\ML_int[5][21] ), .A2(n40), .ZN(n71) );
  INV_X1 U199 ( .A(n72), .ZN(\ML_int[6][20] ) );
  NAND2_X1 U200 ( .A1(\ML_int[5][20] ), .A2(n40), .ZN(n72) );
  INV_X1 U201 ( .A(n73), .ZN(\ML_int[6][1] ) );
  NAND2_X1 U202 ( .A1(\ML_int[5][1] ), .A2(n41), .ZN(n73) );
  INV_X1 U203 ( .A(n74), .ZN(\ML_int[6][19] ) );
  NAND2_X1 U204 ( .A1(\ML_int[5][19] ), .A2(n40), .ZN(n74) );
  INV_X1 U205 ( .A(n75), .ZN(\ML_int[6][18] ) );
  NAND2_X1 U206 ( .A1(\ML_int[5][18] ), .A2(n40), .ZN(n75) );
  INV_X1 U207 ( .A(n76), .ZN(\ML_int[6][17] ) );
  NAND2_X1 U208 ( .A1(\ML_int[5][17] ), .A2(n40), .ZN(n76) );
  INV_X1 U209 ( .A(n77), .ZN(\ML_int[6][16] ) );
  NAND2_X1 U210 ( .A1(\ML_int[5][16] ), .A2(n40), .ZN(n77) );
  INV_X1 U211 ( .A(n78), .ZN(\ML_int[6][15] ) );
  NAND2_X1 U212 ( .A1(\ML_int[5][15] ), .A2(n40), .ZN(n78) );
  INV_X1 U213 ( .A(n79), .ZN(\ML_int[6][14] ) );
  NAND2_X1 U214 ( .A1(\ML_int[5][14] ), .A2(n40), .ZN(n79) );
  INV_X1 U215 ( .A(n80), .ZN(\ML_int[6][13] ) );
  NAND2_X1 U216 ( .A1(\ML_int[5][13] ), .A2(n39), .ZN(n80) );
  INV_X1 U217 ( .A(n81), .ZN(\ML_int[6][12] ) );
  NAND2_X1 U218 ( .A1(\ML_int[5][12] ), .A2(n40), .ZN(n81) );
  INV_X1 U219 ( .A(n82), .ZN(\ML_int[6][11] ) );
  NAND2_X1 U220 ( .A1(\ML_int[5][11] ), .A2(n39), .ZN(n82) );
  INV_X1 U221 ( .A(n83), .ZN(\ML_int[6][10] ) );
  NAND2_X1 U222 ( .A1(\ML_int[5][10] ), .A2(n39), .ZN(n83) );
  INV_X1 U223 ( .A(n84), .ZN(\ML_int[6][0] ) );
  NAND2_X1 U224 ( .A1(\ML_int[5][0] ), .A2(n39), .ZN(n84) );
  NAND2_X1 U225 ( .A1(n87), .A2(n88), .ZN(\temp_int_SH[5] ) );
  NAND2_X1 U226 ( .A1(SH[5]), .A2(n85), .ZN(n88) );
  AND2_X1 U227 ( .A1(\ML_int[4][9] ), .A2(n26), .ZN(\ML_int[5][9] ) );
  AND2_X1 U228 ( .A1(\ML_int[4][8] ), .A2(n26), .ZN(\ML_int[5][8] ) );
  AND2_X1 U229 ( .A1(\ML_int[4][7] ), .A2(n26), .ZN(\ML_int[5][7] ) );
  AND2_X1 U230 ( .A1(\ML_int[4][6] ), .A2(n26), .ZN(\ML_int[5][6] ) );
  AND2_X1 U231 ( .A1(\ML_int[4][5] ), .A2(n26), .ZN(\ML_int[5][5] ) );
  AND2_X1 U232 ( .A1(\ML_int[4][4] ), .A2(n26), .ZN(\ML_int[5][4] ) );
  AND2_X1 U233 ( .A1(\ML_int[4][3] ), .A2(n26), .ZN(\ML_int[5][3] ) );
  AND2_X1 U234 ( .A1(\ML_int[4][2] ), .A2(n26), .ZN(\ML_int[5][2] ) );
  AND2_X1 U235 ( .A1(\ML_int[4][1] ), .A2(n35), .ZN(\ML_int[5][1] ) );
  AND2_X1 U236 ( .A1(\ML_int[4][15] ), .A2(n25), .ZN(\ML_int[5][15] ) );
  AND2_X1 U237 ( .A1(\ML_int[4][14] ), .A2(n25), .ZN(\ML_int[5][14] ) );
  AND2_X1 U238 ( .A1(\ML_int[4][13] ), .A2(n25), .ZN(\ML_int[5][13] ) );
  AND2_X1 U239 ( .A1(\ML_int[4][12] ), .A2(n25), .ZN(\ML_int[5][12] ) );
  AND2_X1 U240 ( .A1(\ML_int[4][11] ), .A2(n25), .ZN(\ML_int[5][11] ) );
  AND2_X1 U241 ( .A1(\ML_int[4][10] ), .A2(n25), .ZN(\ML_int[5][10] ) );
  AND2_X1 U242 ( .A1(\ML_int[4][0] ), .A2(n35), .ZN(\ML_int[5][0] ) );
  AOI21_X1 U243 ( .B1(SH[4]), .B2(n85), .A(n86), .ZN(SHMAG[4]) );
  AND2_X1 U244 ( .A1(\ML_int[3][7] ), .A2(n23), .ZN(\ML_int[4][7] ) );
  AND2_X1 U245 ( .A1(\ML_int[3][6] ), .A2(n23), .ZN(\ML_int[4][6] ) );
  AND2_X1 U246 ( .A1(\ML_int[3][5] ), .A2(n23), .ZN(\ML_int[4][5] ) );
  AND2_X1 U247 ( .A1(\ML_int[3][4] ), .A2(n23), .ZN(\ML_int[4][4] ) );
  AND2_X1 U248 ( .A1(\ML_int[3][3] ), .A2(n23), .ZN(\ML_int[4][3] ) );
  AND2_X1 U249 ( .A1(\ML_int[3][2] ), .A2(n23), .ZN(\ML_int[4][2] ) );
  AND2_X1 U250 ( .A1(\ML_int[3][1] ), .A2(n23), .ZN(\ML_int[4][1] ) );
  AND2_X1 U251 ( .A1(\ML_int[3][0] ), .A2(n23), .ZN(\ML_int[4][0] ) );
  AOI21_X1 U252 ( .B1(SH[3]), .B2(n85), .A(n86), .ZN(SHMAG[3]) );
  AND2_X1 U253 ( .A1(\ML_int[2][3] ), .A2(SHMAG[2]), .ZN(\ML_int[3][3] ) );
  AND2_X1 U254 ( .A1(\ML_int[2][2] ), .A2(SHMAG[2]), .ZN(\ML_int[3][2] ) );
  AND2_X1 U255 ( .A1(\ML_int[2][1] ), .A2(SHMAG[2]), .ZN(\ML_int[3][1] ) );
  AND2_X1 U256 ( .A1(\ML_int[2][0] ), .A2(SHMAG[2]), .ZN(\ML_int[3][0] ) );
  AOI21_X1 U257 ( .B1(SH[2]), .B2(n85), .A(n86), .ZN(SHMAG[2]) );
  AND2_X1 U258 ( .A1(\ML_int[1][1] ), .A2(SHMAG[1]), .ZN(\ML_int[2][1] ) );
  AND2_X1 U259 ( .A1(\ML_int[1][0] ), .A2(SHMAG[1]), .ZN(\ML_int[2][0] ) );
  AOI21_X1 U260 ( .B1(SH[1]), .B2(n85), .A(n86), .ZN(SHMAG[1]) );
  AND2_X1 U261 ( .A1(A[0]), .A2(SHMAG[0]), .ZN(\ML_int[1][0] ) );
  AOI21_X1 U262 ( .B1(SH[0]), .B2(n85), .A(n86), .ZN(SHMAG[0]) );
  INV_X1 U263 ( .A(n87), .ZN(n86) );
  NAND2_X1 U264 ( .A1(SH[7]), .A2(n3), .ZN(n87) );
  OR2_X1 U265 ( .A1(n2), .A2(SH[7]), .ZN(n85) );
  INV_X1 U266 ( .A(SH[8]), .ZN(n53) );
endmodule


module fpu_DW_rash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [105:0] A;
  input [8:0] SH;
  output [105:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879;

  INV_X4 U3 ( .A(n2), .ZN(n34) );
  INV_X4 U4 ( .A(n51), .ZN(n53) );
  INV_X4 U5 ( .A(n54), .ZN(n50) );
  INV_X4 U6 ( .A(n53), .ZN(n48) );
  INV_X4 U7 ( .A(n53), .ZN(n49) );
  INV_X4 U8 ( .A(n34), .ZN(n30) );
  NAND2_X2 U9 ( .A1(n801), .A2(n392), .ZN(n179) );
  NAND2_X2 U10 ( .A1(n801), .A2(SH[4]), .ZN(n177) );
  INV_X4 U11 ( .A(n33), .ZN(n32) );
  NAND2_X2 U12 ( .A1(n266), .A2(SH[4]), .ZN(n242) );
  NAND2_X2 U13 ( .A1(n266), .A2(n392), .ZN(n238) );
  INV_X4 U14 ( .A(n2), .ZN(n35) );
  INV_X4 U15 ( .A(n53), .ZN(n47) );
  INV_X4 U16 ( .A(SH[4]), .ZN(n392) );
  NOR2_X2 U17 ( .A1(n383), .A2(n238), .ZN(n408) );
  NAND2_X2 U18 ( .A1(n26), .A2(n794), .ZN(n168) );
  NAND2_X2 U19 ( .A1(n794), .A2(n23), .ZN(n170) );
  NOR2_X2 U20 ( .A1(n242), .A2(n174), .ZN(n171) );
  NOR2_X2 U21 ( .A1(n174), .A2(SH[8]), .ZN(n210) );
  OR2_X4 U22 ( .A1(n879), .A2(n878), .ZN(n1) );
  NAND2_X4 U23 ( .A1(n878), .A2(SH[0]), .ZN(n2) );
  OR2_X4 U24 ( .A1(SH[2]), .A2(n833), .ZN(n3) );
  OR2_X4 U25 ( .A1(n299), .A2(SH[4]), .ZN(n4) );
  INV_X4 U26 ( .A(n31), .ZN(n33) );
  AND2_X4 U27 ( .A1(n386), .A2(SH[4]), .ZN(n5) );
  INV_X4 U28 ( .A(n41), .ZN(n36) );
  INV_X4 U29 ( .A(n34), .ZN(n31) );
  INV_X4 U30 ( .A(n35), .ZN(n29) );
  INV_X4 U31 ( .A(n396), .ZN(n55) );
  NOR2_X2 U32 ( .A1(SH[0]), .A2(n878), .ZN(n396) );
  NAND2_X2 U33 ( .A1(n878), .A2(n879), .ZN(n6) );
  INV_X4 U34 ( .A(n1), .ZN(n44) );
  INV_X4 U35 ( .A(n396), .ZN(n54) );
  INV_X4 U36 ( .A(n181), .ZN(n7) );
  INV_X4 U37 ( .A(n19), .ZN(n15) );
  INV_X4 U38 ( .A(n18), .ZN(n17) );
  INV_X4 U39 ( .A(n1), .ZN(n45) );
  INV_X4 U40 ( .A(n55), .ZN(n52) );
  INV_X4 U41 ( .A(n55), .ZN(n51) );
  INV_X4 U42 ( .A(n7), .ZN(n8) );
  INV_X4 U43 ( .A(n393), .ZN(n19) );
  INV_X4 U44 ( .A(n409), .ZN(n58) );
  INV_X4 U45 ( .A(n58), .ZN(n56) );
  INV_X4 U46 ( .A(n1), .ZN(n46) );
  INV_X4 U47 ( .A(n1), .ZN(n43) );
  INV_X4 U48 ( .A(n394), .ZN(n24) );
  INV_X4 U49 ( .A(n41), .ZN(n38) );
  INV_X4 U50 ( .A(n1), .ZN(n42) );
  INV_X4 U51 ( .A(n24), .ZN(n21) );
  INV_X4 U52 ( .A(n393), .ZN(n18) );
  INV_X4 U53 ( .A(n6), .ZN(n41) );
  INV_X4 U54 ( .A(n58), .ZN(n57) );
  INV_X4 U55 ( .A(n3), .ZN(n25) );
  INV_X4 U56 ( .A(n4), .ZN(n13) );
  INV_X4 U57 ( .A(n312), .ZN(n11) );
  INV_X4 U58 ( .A(n18), .ZN(n16) );
  INV_X4 U59 ( .A(n24), .ZN(n23) );
  INV_X4 U60 ( .A(n24), .ZN(n22) );
  INV_X4 U61 ( .A(n24), .ZN(n20) );
  INV_X4 U62 ( .A(n3), .ZN(n28) );
  INV_X4 U63 ( .A(n3), .ZN(n27) );
  INV_X4 U64 ( .A(n3), .ZN(n26) );
  INV_X4 U65 ( .A(n41), .ZN(n40) );
  INV_X4 U66 ( .A(n41), .ZN(n37) );
  INV_X4 U67 ( .A(n41), .ZN(n39) );
  INV_X4 U68 ( .A(n11), .ZN(n12) );
  INV_X4 U69 ( .A(n5), .ZN(n10) );
  INV_X4 U70 ( .A(n5), .ZN(n9) );
  INV_X4 U71 ( .A(n409), .ZN(n59) );
  INV_X4 U72 ( .A(n4), .ZN(n14) );
  AND2_X4 U73 ( .A1(n409), .A2(n794), .ZN(n164) );
  AND2_X4 U74 ( .A1(n16), .A2(n794), .ZN(n162) );
  INV_X4 U75 ( .A(n859), .ZN(n174) );
  INV_X4 U76 ( .A(n376), .ZN(n383) );
  INV_X4 U77 ( .A(A[2]), .ZN(n60) );
  INV_X4 U78 ( .A(A[3]), .ZN(n61) );
  INV_X4 U79 ( .A(A[4]), .ZN(n62) );
  INV_X4 U80 ( .A(A[5]), .ZN(n63) );
  INV_X4 U81 ( .A(A[6]), .ZN(n64) );
  INV_X4 U82 ( .A(A[7]), .ZN(n65) );
  INV_X4 U83 ( .A(A[8]), .ZN(n66) );
  INV_X4 U84 ( .A(A[91]), .ZN(n67) );
  INV_X4 U85 ( .A(A[92]), .ZN(n68) );
  INV_X4 U86 ( .A(A[93]), .ZN(n69) );
  INV_X4 U87 ( .A(A[94]), .ZN(n70) );
  INV_X4 U88 ( .A(A[96]), .ZN(n71) );
  INV_X4 U89 ( .A(A[97]), .ZN(n72) );
  INV_X4 U90 ( .A(A[95]), .ZN(n73) );
  INV_X4 U91 ( .A(A[90]), .ZN(n74) );
  INV_X4 U92 ( .A(A[99]), .ZN(n75) );
  INV_X4 U93 ( .A(A[101]), .ZN(n76) );
  INV_X4 U94 ( .A(A[102]), .ZN(n77) );
  INV_X4 U95 ( .A(A[100]), .ZN(n78) );
  INV_X4 U96 ( .A(A[98]), .ZN(n79) );
  INV_X4 U97 ( .A(A[49]), .ZN(n80) );
  INV_X4 U98 ( .A(A[53]), .ZN(n81) );
  INV_X4 U99 ( .A(A[54]), .ZN(n82) );
  INV_X4 U100 ( .A(A[56]), .ZN(n83) );
  INV_X4 U101 ( .A(A[57]), .ZN(n84) );
  INV_X4 U102 ( .A(A[55]), .ZN(n85) );
  INV_X4 U103 ( .A(A[83]), .ZN(n86) );
  INV_X4 U104 ( .A(A[84]), .ZN(n87) );
  INV_X4 U105 ( .A(A[85]), .ZN(n88) );
  INV_X4 U106 ( .A(A[86]), .ZN(n89) );
  INV_X4 U107 ( .A(A[88]), .ZN(n90) );
  INV_X4 U108 ( .A(A[89]), .ZN(n91) );
  INV_X4 U109 ( .A(A[87]), .ZN(n92) );
  INV_X4 U110 ( .A(A[75]), .ZN(n93) );
  INV_X4 U111 ( .A(A[76]), .ZN(n94) );
  INV_X4 U112 ( .A(A[77]), .ZN(n95) );
  INV_X4 U113 ( .A(A[78]), .ZN(n96) );
  INV_X4 U114 ( .A(A[80]), .ZN(n97) );
  INV_X4 U115 ( .A(A[81]), .ZN(n98) );
  INV_X4 U116 ( .A(A[79]), .ZN(n99) );
  INV_X4 U117 ( .A(A[59]), .ZN(n100) );
  INV_X4 U118 ( .A(A[60]), .ZN(n101) );
  INV_X4 U119 ( .A(A[61]), .ZN(n102) );
  INV_X4 U120 ( .A(A[62]), .ZN(n103) );
  INV_X4 U121 ( .A(A[64]), .ZN(n104) );
  INV_X4 U122 ( .A(A[65]), .ZN(n105) );
  INV_X4 U123 ( .A(A[63]), .ZN(n106) );
  INV_X4 U124 ( .A(A[67]), .ZN(n107) );
  INV_X4 U125 ( .A(A[68]), .ZN(n108) );
  INV_X4 U126 ( .A(A[69]), .ZN(n109) );
  INV_X4 U127 ( .A(A[70]), .ZN(n110) );
  INV_X4 U128 ( .A(A[72]), .ZN(n111) );
  INV_X4 U129 ( .A(A[73]), .ZN(n112) );
  INV_X4 U130 ( .A(A[71]), .ZN(n113) );
  INV_X4 U131 ( .A(A[52]), .ZN(n114) );
  INV_X4 U132 ( .A(A[58]), .ZN(n115) );
  INV_X4 U133 ( .A(A[66]), .ZN(n116) );
  INV_X4 U134 ( .A(A[82]), .ZN(n117) );
  INV_X4 U135 ( .A(A[74]), .ZN(n118) );
  INV_X4 U136 ( .A(A[51]), .ZN(n119) );
  INV_X4 U137 ( .A(A[50]), .ZN(n120) );
  INV_X4 U138 ( .A(A[43]), .ZN(n121) );
  INV_X4 U139 ( .A(A[44]), .ZN(n122) );
  INV_X4 U140 ( .A(A[45]), .ZN(n123) );
  INV_X4 U141 ( .A(A[46]), .ZN(n124) );
  INV_X4 U142 ( .A(A[48]), .ZN(n125) );
  INV_X4 U143 ( .A(A[47]), .ZN(n126) );
  INV_X4 U144 ( .A(A[11]), .ZN(n127) );
  INV_X4 U145 ( .A(A[12]), .ZN(n128) );
  INV_X4 U146 ( .A(A[13]), .ZN(n129) );
  INV_X4 U147 ( .A(A[14]), .ZN(n130) );
  INV_X4 U148 ( .A(A[16]), .ZN(n131) );
  INV_X4 U149 ( .A(A[17]), .ZN(n132) );
  INV_X4 U150 ( .A(A[15]), .ZN(n133) );
  INV_X4 U151 ( .A(A[19]), .ZN(n134) );
  INV_X4 U152 ( .A(A[21]), .ZN(n135) );
  INV_X4 U153 ( .A(A[22]), .ZN(n136) );
  INV_X4 U154 ( .A(A[24]), .ZN(n137) );
  INV_X4 U155 ( .A(A[25]), .ZN(n138) );
  INV_X4 U156 ( .A(A[23]), .ZN(n139) );
  INV_X4 U157 ( .A(A[27]), .ZN(n140) );
  INV_X4 U158 ( .A(A[28]), .ZN(n141) );
  INV_X4 U159 ( .A(A[29]), .ZN(n142) );
  INV_X4 U160 ( .A(A[30]), .ZN(n143) );
  INV_X4 U161 ( .A(A[32]), .ZN(n144) );
  INV_X4 U162 ( .A(A[33]), .ZN(n145) );
  INV_X4 U163 ( .A(A[31]), .ZN(n146) );
  INV_X4 U164 ( .A(A[35]), .ZN(n147) );
  INV_X4 U165 ( .A(A[36]), .ZN(n148) );
  INV_X4 U166 ( .A(A[37]), .ZN(n149) );
  INV_X4 U167 ( .A(A[38]), .ZN(n150) );
  INV_X4 U168 ( .A(A[40]), .ZN(n151) );
  INV_X4 U169 ( .A(A[41]), .ZN(n152) );
  INV_X4 U170 ( .A(A[39]), .ZN(n153) );
  INV_X4 U171 ( .A(A[34]), .ZN(n154) );
  INV_X4 U172 ( .A(A[26]), .ZN(n155) );
  INV_X4 U173 ( .A(A[18]), .ZN(n156) );
  INV_X4 U174 ( .A(A[10]), .ZN(n157) );
  INV_X4 U175 ( .A(A[9]), .ZN(n158) );
  INV_X4 U176 ( .A(A[42]), .ZN(n159) );
  AOI21_X1 U177 ( .B1(n160), .B2(n161), .A(SH[8]), .ZN(B[9]) );
  AOI221_X1 U178 ( .B1(n162), .B2(n163), .C1(n164), .C2(n165), .A(n166), .ZN(
        n161) );
  OAI22_X1 U179 ( .A1(n167), .A2(n168), .B1(n169), .B2(n170), .ZN(n166) );
  AOI221_X1 U180 ( .B1(n171), .B2(n172), .C1(n173), .C2(n174), .A(n175), .ZN(
        n160) );
  OAI22_X1 U181 ( .A1(n176), .A2(n177), .B1(n178), .B2(n179), .ZN(n175) );
  NOR2_X1 U182 ( .A1(n180), .A2(n8), .ZN(B[99]) );
  NOR2_X1 U183 ( .A1(n182), .A2(n8), .ZN(B[98]) );
  NOR2_X1 U184 ( .A1(n183), .A2(n8), .ZN(B[97]) );
  NOR2_X1 U185 ( .A1(n184), .A2(n8), .ZN(B[96]) );
  NOR2_X1 U186 ( .A1(n185), .A2(n8), .ZN(B[95]) );
  NOR2_X1 U187 ( .A1(n186), .A2(n8), .ZN(B[94]) );
  NOR2_X1 U188 ( .A1(n187), .A2(n8), .ZN(B[93]) );
  NOR2_X1 U189 ( .A1(n188), .A2(n8), .ZN(B[92]) );
  NOR2_X1 U190 ( .A1(n189), .A2(n8), .ZN(B[91]) );
  NOR2_X1 U191 ( .A1(n190), .A2(n8), .ZN(B[90]) );
  AOI21_X1 U192 ( .B1(n191), .B2(n192), .A(SH[8]), .ZN(B[8]) );
  AOI221_X1 U193 ( .B1(n162), .B2(n193), .C1(n164), .C2(n194), .A(n195), .ZN(
        n192) );
  OAI22_X1 U194 ( .A1(n196), .A2(n168), .B1(n197), .B2(n170), .ZN(n195) );
  AOI221_X1 U195 ( .B1(n171), .B2(n198), .C1(n199), .C2(n174), .A(n200), .ZN(
        n191) );
  OAI22_X1 U196 ( .A1(n201), .A2(n177), .B1(n202), .B2(n179), .ZN(n200) );
  NOR2_X1 U197 ( .A1(n203), .A2(n204), .ZN(B[89]) );
  NOR2_X1 U198 ( .A1(n205), .A2(n204), .ZN(B[88]) );
  NOR2_X1 U199 ( .A1(n206), .A2(n204), .ZN(B[87]) );
  NOR2_X1 U200 ( .A1(n207), .A2(n204), .ZN(B[86]) );
  NOR2_X1 U201 ( .A1(n208), .A2(n204), .ZN(B[85]) );
  AND2_X1 U202 ( .A1(n209), .A2(n210), .ZN(B[84]) );
  NOR2_X1 U203 ( .A1(n211), .A2(n212), .ZN(B[83]) );
  NOR2_X1 U204 ( .A1(n213), .A2(n212), .ZN(B[82]) );
  NOR2_X1 U205 ( .A1(n214), .A2(n212), .ZN(B[81]) );
  NOR2_X1 U206 ( .A1(n215), .A2(n212), .ZN(B[80]) );
  AOI21_X1 U207 ( .B1(n216), .B2(n217), .A(SH[8]), .ZN(B[7]) );
  AOI221_X1 U208 ( .B1(n218), .B2(n219), .C1(n220), .C2(n221), .A(n222), .ZN(
        n217) );
  INV_X1 U209 ( .A(n223), .ZN(n222) );
  AOI22_X1 U210 ( .A1(n224), .A2(n164), .B1(n225), .B2(n162), .ZN(n223) );
  AOI221_X1 U211 ( .B1(n171), .B2(n226), .C1(n227), .C2(n174), .A(n228), .ZN(
        n216) );
  OAI22_X1 U212 ( .A1(n229), .A2(n177), .B1(n230), .B2(n179), .ZN(n228) );
  AND2_X1 U213 ( .A1(n231), .A2(n210), .ZN(B[79]) );
  AND2_X1 U214 ( .A1(n232), .A2(n210), .ZN(B[78]) );
  AND2_X1 U215 ( .A1(n233), .A2(n210), .ZN(B[77]) );
  AND2_X1 U216 ( .A1(n234), .A2(n210), .ZN(B[76]) );
  AND2_X1 U217 ( .A1(n235), .A2(n210), .ZN(B[75]) );
  AND2_X1 U218 ( .A1(n236), .A2(n210), .ZN(B[74]) );
  AND2_X1 U219 ( .A1(n173), .A2(n210), .ZN(B[73]) );
  OAI222_X1 U220 ( .A1(n237), .A2(n238), .B1(n239), .B2(n240), .C1(n241), .C2(
        n242), .ZN(n173) );
  AND2_X1 U221 ( .A1(n199), .A2(n210), .ZN(B[72]) );
  OAI222_X1 U222 ( .A1(n243), .A2(n238), .B1(n244), .B2(n239), .C1(n245), .C2(
        n242), .ZN(n199) );
  AND2_X1 U223 ( .A1(n227), .A2(n210), .ZN(B[71]) );
  OAI222_X1 U224 ( .A1(n246), .A2(n238), .B1(n247), .B2(n239), .C1(n248), .C2(
        n242), .ZN(n227) );
  AND2_X1 U225 ( .A1(n249), .A2(n210), .ZN(B[70]) );
  AOI21_X1 U226 ( .B1(n250), .B2(n251), .A(SH[8]), .ZN(B[6]) );
  AOI221_X1 U227 ( .B1(n218), .B2(n252), .C1(n220), .C2(n253), .A(n254), .ZN(
        n251) );
  INV_X1 U228 ( .A(n255), .ZN(n254) );
  AOI22_X1 U229 ( .A1(n256), .A2(n164), .B1(n257), .B2(n162), .ZN(n255) );
  AOI221_X1 U230 ( .B1(n171), .B2(n258), .C1(n249), .C2(n174), .A(n259), .ZN(
        n250) );
  OAI22_X1 U231 ( .A1(n260), .A2(n177), .B1(n261), .B2(n179), .ZN(n259) );
  OAI222_X1 U232 ( .A1(n262), .A2(n238), .B1(n263), .B2(n239), .C1(n264), .C2(
        n242), .ZN(n249) );
  OR2_X1 U233 ( .A1(n265), .A2(n266), .ZN(n239) );
  AND2_X1 U234 ( .A1(n267), .A2(n210), .ZN(B[69]) );
  AND2_X1 U235 ( .A1(n268), .A2(n210), .ZN(B[68]) );
  NOR2_X1 U236 ( .A1(n269), .A2(n212), .ZN(B[67]) );
  NOR2_X1 U237 ( .A1(n270), .A2(n212), .ZN(B[66]) );
  NOR2_X1 U238 ( .A1(n271), .A2(n212), .ZN(B[65]) );
  NOR2_X1 U239 ( .A1(n272), .A2(n212), .ZN(B[64]) );
  INV_X1 U240 ( .A(n210), .ZN(n212) );
  OAI222_X1 U241 ( .A1(n273), .A2(n9), .B1(n185), .B2(n4), .C1(n274), .C2(n181), .ZN(B[63]) );
  OAI222_X1 U242 ( .A1(n275), .A2(n9), .B1(n186), .B2(n4), .C1(n276), .C2(n181), .ZN(B[62]) );
  OAI222_X1 U243 ( .A1(n277), .A2(n9), .B1(n187), .B2(n4), .C1(n278), .C2(n8), 
        .ZN(B[61]) );
  OAI222_X1 U244 ( .A1(n279), .A2(n9), .B1(n188), .B2(n4), .C1(n280), .C2(n8), 
        .ZN(B[60]) );
  AOI21_X1 U245 ( .B1(n281), .B2(n282), .A(SH[8]), .ZN(B[5]) );
  AOI221_X1 U246 ( .B1(n218), .B2(n283), .C1(n220), .C2(n163), .A(n284), .ZN(
        n282) );
  INV_X1 U247 ( .A(n285), .ZN(n284) );
  AOI22_X1 U248 ( .A1(n286), .A2(n164), .B1(n165), .B2(n162), .ZN(n285) );
  AOI221_X1 U249 ( .B1(n171), .B2(n287), .C1(n267), .C2(n174), .A(n288), .ZN(
        n281) );
  OAI22_X1 U250 ( .A1(n289), .A2(n177), .B1(n290), .B2(n179), .ZN(n288) );
  OAI222_X1 U251 ( .A1(n291), .A2(n238), .B1(n292), .B2(n293), .C1(n294), .C2(
        n242), .ZN(n267) );
  OAI222_X1 U252 ( .A1(n295), .A2(n9), .B1(n189), .B2(n4), .C1(n296), .C2(n8), 
        .ZN(B[59]) );
  OAI222_X1 U253 ( .A1(n297), .A2(n10), .B1(n190), .B2(n4), .C1(n298), .C2(n8), 
        .ZN(B[58]) );
  OAI222_X1 U254 ( .A1(n176), .A2(n181), .B1(n237), .B2(n9), .C1(n203), .C2(
        n299), .ZN(B[57]) );
  INV_X1 U255 ( .A(n300), .ZN(n203) );
  INV_X1 U256 ( .A(n301), .ZN(n237) );
  OAI222_X1 U257 ( .A1(n201), .A2(n181), .B1(n243), .B2(n9), .C1(n205), .C2(
        n299), .ZN(B[56]) );
  INV_X1 U258 ( .A(n302), .ZN(n205) );
  INV_X1 U259 ( .A(n303), .ZN(n243) );
  OAI222_X1 U260 ( .A1(n229), .A2(n181), .B1(n246), .B2(n10), .C1(n206), .C2(
        n299), .ZN(B[55]) );
  INV_X1 U261 ( .A(n304), .ZN(n206) );
  INV_X1 U262 ( .A(n305), .ZN(n246) );
  OAI222_X1 U263 ( .A1(n260), .A2(n181), .B1(n262), .B2(n10), .C1(n207), .C2(
        n299), .ZN(B[54]) );
  INV_X1 U264 ( .A(n306), .ZN(n207) );
  INV_X1 U265 ( .A(n307), .ZN(n262) );
  OAI222_X1 U266 ( .A1(n289), .A2(n181), .B1(n291), .B2(n9), .C1(n208), .C2(
        n299), .ZN(B[53]) );
  INV_X1 U267 ( .A(n308), .ZN(n291) );
  OAI221_X1 U268 ( .B1(n309), .B2(n9), .C1(n310), .C2(n8), .A(n311), .ZN(B[52]) );
  AOI22_X1 U269 ( .A1(n12), .A2(n313), .B1(n14), .B2(n314), .ZN(n311) );
  OAI221_X1 U270 ( .B1(n315), .B2(n9), .C1(n316), .C2(n8), .A(n317), .ZN(B[51]) );
  AOI22_X1 U271 ( .A1(n12), .A2(n318), .B1(n14), .B2(n319), .ZN(n317) );
  OAI221_X1 U272 ( .B1(n320), .B2(n9), .C1(n321), .C2(n8), .A(n322), .ZN(B[50]) );
  AOI22_X1 U273 ( .A1(n12), .A2(n323), .B1(n14), .B2(n324), .ZN(n322) );
  AOI21_X1 U274 ( .B1(n325), .B2(n326), .A(SH[8]), .ZN(B[4]) );
  AOI221_X1 U275 ( .B1(n218), .B2(n327), .C1(n220), .C2(n193), .A(n328), .ZN(
        n326) );
  INV_X1 U276 ( .A(n329), .ZN(n328) );
  AOI22_X1 U277 ( .A1(n330), .A2(n164), .B1(n194), .B2(n162), .ZN(n329) );
  INV_X1 U278 ( .A(n168), .ZN(n220) );
  INV_X1 U279 ( .A(n170), .ZN(n218) );
  AOI221_X1 U280 ( .B1(n171), .B2(n331), .C1(n268), .C2(n174), .A(n332), .ZN(
        n325) );
  OAI22_X1 U281 ( .A1(n310), .A2(n177), .B1(n333), .B2(n179), .ZN(n332) );
  OAI222_X1 U282 ( .A1(n309), .A2(n238), .B1(n334), .B2(n293), .C1(n335), .C2(
        n242), .ZN(n268) );
  INV_X1 U283 ( .A(n336), .ZN(n293) );
  INV_X1 U284 ( .A(n337), .ZN(n309) );
  OAI221_X1 U285 ( .B1(n338), .B2(n9), .C1(n339), .C2(n8), .A(n340), .ZN(B[49]) );
  AOI22_X1 U286 ( .A1(n12), .A2(n341), .B1(n14), .B2(n342), .ZN(n340) );
  OAI221_X1 U287 ( .B1(n343), .B2(n9), .C1(n344), .C2(n8), .A(n345), .ZN(B[48]) );
  AOI22_X1 U288 ( .A1(n12), .A2(n346), .B1(n14), .B2(n347), .ZN(n345) );
  OAI221_X1 U289 ( .B1(n185), .B2(n11), .C1(n273), .C2(n4), .A(n348), .ZN(
        B[47]) );
  INV_X1 U290 ( .A(n349), .ZN(n348) );
  OAI22_X1 U291 ( .A1(n9), .A2(n274), .B1(n8), .B2(n350), .ZN(n349) );
  OAI221_X1 U292 ( .B1(n186), .B2(n11), .C1(n275), .C2(n4), .A(n351), .ZN(
        B[46]) );
  INV_X1 U293 ( .A(n352), .ZN(n351) );
  OAI22_X1 U294 ( .A1(n9), .A2(n276), .B1(n8), .B2(n353), .ZN(n352) );
  INV_X1 U295 ( .A(n354), .ZN(B[45]) );
  AOI221_X1 U296 ( .B1(n355), .B2(n312), .C1(n356), .C2(n14), .A(n357), .ZN(
        n354) );
  OAI22_X1 U297 ( .A1(n9), .A2(n278), .B1(n8), .B2(n358), .ZN(n357) );
  INV_X1 U298 ( .A(n359), .ZN(B[44]) );
  AOI221_X1 U299 ( .B1(n360), .B2(n312), .C1(n361), .C2(n14), .A(n362), .ZN(
        n359) );
  OAI22_X1 U300 ( .A1(n9), .A2(n280), .B1(n8), .B2(n363), .ZN(n362) );
  INV_X1 U301 ( .A(n364), .ZN(B[43]) );
  AOI221_X1 U302 ( .B1(n365), .B2(n312), .C1(n366), .C2(n14), .A(n367), .ZN(
        n364) );
  OAI22_X1 U303 ( .A1(n10), .A2(n296), .B1(n8), .B2(n368), .ZN(n367) );
  INV_X1 U304 ( .A(n369), .ZN(B[42]) );
  AOI221_X1 U305 ( .B1(n370), .B2(n312), .C1(n371), .C2(n14), .A(n372), .ZN(
        n369) );
  OAI22_X1 U306 ( .A1(n9), .A2(n298), .B1(n8), .B2(n373), .ZN(n372) );
  OAI221_X1 U307 ( .B1(n176), .B2(n9), .C1(n178), .C2(n8), .A(n374), .ZN(B[41]) );
  AOI222_X1 U308 ( .A1(n14), .A2(n301), .B1(n375), .B2(n376), .C1(n312), .C2(
        n377), .ZN(n374) );
  INV_X1 U309 ( .A(n241), .ZN(n377) );
  OAI221_X1 U310 ( .B1(n201), .B2(n9), .C1(n202), .C2(n8), .A(n378), .ZN(B[40]) );
  AOI222_X1 U311 ( .A1(n13), .A2(n303), .B1(n379), .B2(n380), .C1(n12), .C2(
        n381), .ZN(n378) );
  INV_X1 U312 ( .A(n382), .ZN(n201) );
  OAI221_X1 U313 ( .B1(n269), .B2(n383), .C1(n316), .C2(n11), .A(n384), .ZN(
        B[3]) );
  AOI22_X1 U314 ( .A1(n14), .A2(n385), .B1(n386), .B2(n387), .ZN(n384) );
  OAI21_X1 U315 ( .B1(n388), .B2(n265), .A(n389), .ZN(n387) );
  MUX2_X1 U316 ( .A(n390), .B(n391), .S(n392), .Z(n389) );
  AOI222_X1 U317 ( .A1(n15), .A2(n224), .B1(n21), .B2(n221), .C1(n25), .C2(
        n225), .ZN(n391) );
  OAI221_X1 U318 ( .B1(n31), .B2(n66), .C1(n39), .C2(n65), .A(n395), .ZN(n224)
         );
  AOI22_X1 U319 ( .A1(A[10]), .A2(n44), .B1(A[9]), .B2(n47), .ZN(n395) );
  AOI221_X1 U320 ( .B1(A[6]), .B2(n42), .C1(A[5]), .C2(n47), .A(n397), .ZN(
        n388) );
  OAI22_X1 U321 ( .A1(n36), .A2(n61), .B1(n29), .B2(n62), .ZN(n397) );
  INV_X1 U322 ( .A(n398), .ZN(n385) );
  AOI222_X1 U323 ( .A1(n399), .A2(n400), .B1(n318), .B2(n336), .C1(n319), .C2(
        n401), .ZN(n269) );
  OAI221_X1 U324 ( .B1(n229), .B2(n9), .C1(n230), .C2(n8), .A(n402), .ZN(B[39]) );
  AOI222_X1 U325 ( .A1(n13), .A2(n305), .B1(n379), .B2(n403), .C1(n12), .C2(
        n404), .ZN(n402) );
  INV_X1 U326 ( .A(n248), .ZN(n404) );
  OAI221_X1 U327 ( .B1(n260), .B2(n9), .C1(n261), .C2(n8), .A(n405), .ZN(B[38]) );
  AOI222_X1 U328 ( .A1(n14), .A2(n307), .B1(n379), .B2(n406), .C1(n12), .C2(
        n407), .ZN(n405) );
  INV_X1 U329 ( .A(n264), .ZN(n407) );
  AND2_X1 U330 ( .A1(n408), .A2(n409), .ZN(n379) );
  OAI221_X1 U331 ( .B1(n289), .B2(n9), .C1(n290), .C2(n8), .A(n410), .ZN(B[37]) );
  AOI222_X1 U332 ( .A1(n14), .A2(n308), .B1(n408), .B2(n411), .C1(n12), .C2(
        n412), .ZN(n410) );
  INV_X1 U333 ( .A(n294), .ZN(n412) );
  INV_X1 U334 ( .A(n292), .ZN(n411) );
  OAI221_X1 U335 ( .B1(n310), .B2(n9), .C1(n333), .C2(n8), .A(n413), .ZN(B[36]) );
  AOI222_X1 U336 ( .A1(n13), .A2(n337), .B1(n12), .B2(n314), .C1(n408), .C2(
        n313), .ZN(n413) );
  INV_X1 U337 ( .A(n334), .ZN(n313) );
  OAI221_X1 U338 ( .B1(n316), .B2(n9), .C1(n398), .C2(n8), .A(n414), .ZN(B[35]) );
  AOI222_X1 U339 ( .A1(n13), .A2(n399), .B1(n12), .B2(n319), .C1(n408), .C2(
        n318), .ZN(n414) );
  OAI221_X1 U340 ( .B1(n321), .B2(n9), .C1(n415), .C2(n8), .A(n416), .ZN(B[34]) );
  AOI222_X1 U341 ( .A1(n14), .A2(n417), .B1(n12), .B2(n324), .C1(n408), .C2(
        n323), .ZN(n416) );
  OAI221_X1 U342 ( .B1(n339), .B2(n9), .C1(n418), .C2(n8), .A(n419), .ZN(B[33]) );
  AOI222_X1 U343 ( .A1(n14), .A2(n420), .B1(n12), .B2(n342), .C1(n408), .C2(
        n341), .ZN(n419) );
  OAI221_X1 U344 ( .B1(n344), .B2(n9), .C1(n421), .C2(n8), .A(n422), .ZN(B[32]) );
  AOI222_X1 U345 ( .A1(n13), .A2(n423), .B1(n12), .B2(n347), .C1(n408), .C2(
        n346), .ZN(n422) );
  OAI221_X1 U346 ( .B1(n350), .B2(n9), .C1(n424), .C2(n8), .A(n425), .ZN(B[31]) );
  AOI222_X1 U347 ( .A1(n14), .A2(n426), .B1(n12), .B2(n427), .C1(n408), .C2(
        n428), .ZN(n425) );
  INV_X1 U348 ( .A(n185), .ZN(n428) );
  OAI221_X1 U349 ( .B1(n353), .B2(n10), .C1(n429), .C2(n8), .A(n430), .ZN(
        B[30]) );
  AOI222_X1 U350 ( .A1(n13), .A2(n431), .B1(n12), .B2(n432), .C1(n408), .C2(
        n433), .ZN(n430) );
  INV_X1 U351 ( .A(n186), .ZN(n433) );
  INV_X1 U352 ( .A(n276), .ZN(n431) );
  OAI221_X1 U353 ( .B1(n270), .B2(n383), .C1(n321), .C2(n11), .A(n434), .ZN(
        B[2]) );
  AOI22_X1 U354 ( .A1(n14), .A2(n435), .B1(n386), .B2(n436), .ZN(n434) );
  OAI21_X1 U355 ( .B1(n437), .B2(n265), .A(n438), .ZN(n436) );
  MUX2_X1 U356 ( .A(n439), .B(n440), .S(n392), .Z(n438) );
  AOI222_X1 U357 ( .A1(n15), .A2(n256), .B1(n21), .B2(n253), .C1(n25), .C2(
        n257), .ZN(n440) );
  OAI221_X1 U358 ( .B1(n29), .B2(n65), .C1(n36), .C2(n64), .A(n441), .ZN(n256)
         );
  AOI22_X1 U359 ( .A1(A[9]), .A2(n42), .B1(A[8]), .B2(n47), .ZN(n441) );
  AOI221_X1 U360 ( .B1(A[5]), .B2(n42), .C1(A[4]), .C2(n47), .A(n442), .ZN(
        n437) );
  OAI22_X1 U361 ( .A1(n36), .A2(n60), .B1(n29), .B2(n61), .ZN(n442) );
  INV_X1 U362 ( .A(n415), .ZN(n435) );
  AOI222_X1 U363 ( .A1(n417), .A2(n400), .B1(n323), .B2(n336), .C1(n324), .C2(
        n401), .ZN(n270) );
  OAI221_X1 U364 ( .B1(n358), .B2(n10), .C1(n443), .C2(n8), .A(n444), .ZN(
        B[29]) );
  AOI222_X1 U365 ( .A1(n13), .A2(n445), .B1(n12), .B2(n356), .C1(n408), .C2(
        n355), .ZN(n444) );
  INV_X1 U366 ( .A(n187), .ZN(n355) );
  INV_X1 U367 ( .A(n278), .ZN(n445) );
  OAI221_X1 U368 ( .B1(n363), .B2(n10), .C1(n446), .C2(n8), .A(n447), .ZN(
        B[28]) );
  AOI222_X1 U369 ( .A1(n13), .A2(n448), .B1(n12), .B2(n361), .C1(n408), .C2(
        n360), .ZN(n447) );
  OAI221_X1 U370 ( .B1(n368), .B2(n10), .C1(n449), .C2(n8), .A(n450), .ZN(
        B[27]) );
  AOI222_X1 U371 ( .A1(n13), .A2(n451), .B1(n12), .B2(n366), .C1(n408), .C2(
        n365), .ZN(n450) );
  INV_X1 U372 ( .A(n189), .ZN(n365) );
  INV_X1 U373 ( .A(n296), .ZN(n451) );
  OAI221_X1 U374 ( .B1(n373), .B2(n10), .C1(n452), .C2(n8), .A(n453), .ZN(
        B[26]) );
  AOI222_X1 U375 ( .A1(n13), .A2(n454), .B1(n12), .B2(n371), .C1(n408), .C2(
        n370), .ZN(n453) );
  INV_X1 U376 ( .A(n190), .ZN(n370) );
  INV_X1 U377 ( .A(n298), .ZN(n454) );
  OAI221_X1 U378 ( .B1(n178), .B2(n10), .C1(n455), .C2(n8), .A(n456), .ZN(
        B[25]) );
  AOI222_X1 U379 ( .A1(n13), .A2(n457), .B1(n458), .B2(n300), .C1(n312), .C2(
        n301), .ZN(n456) );
  OAI221_X1 U380 ( .B1(n459), .B2(n18), .C1(n460), .C2(n59), .A(n461), .ZN(
        n301) );
  AOI22_X1 U381 ( .A1(n20), .A2(n462), .B1(n25), .B2(n463), .ZN(n461) );
  OAI22_X1 U382 ( .A1(n241), .A2(SH[4]), .B1(n240), .B2(n464), .ZN(n300) );
  AOI221_X1 U383 ( .B1(n465), .B2(n15), .C1(n466), .C2(n56), .A(n467), .ZN(
        n241) );
  INV_X1 U384 ( .A(n468), .ZN(n467) );
  AOI22_X1 U385 ( .A1(n22), .A2(n469), .B1(n28), .B2(n470), .ZN(n468) );
  INV_X1 U386 ( .A(n176), .ZN(n457) );
  AOI221_X1 U387 ( .B1(n471), .B2(n17), .C1(n472), .C2(n56), .A(n473), .ZN(
        n176) );
  INV_X1 U388 ( .A(n474), .ZN(n473) );
  AOI22_X1 U389 ( .A1(n21), .A2(n475), .B1(n25), .B2(n476), .ZN(n474) );
  INV_X1 U390 ( .A(n172), .ZN(n455) );
  OAI221_X1 U391 ( .B1(n477), .B2(n18), .C1(n478), .C2(n59), .A(n479), .ZN(
        n172) );
  AOI22_X1 U392 ( .A1(n21), .A2(n480), .B1(n25), .B2(n481), .ZN(n479) );
  INV_X1 U393 ( .A(n482), .ZN(n477) );
  AOI221_X1 U394 ( .B1(n483), .B2(n15), .C1(n484), .C2(n56), .A(n485), .ZN(
        n178) );
  INV_X1 U395 ( .A(n486), .ZN(n485) );
  AOI22_X1 U396 ( .A1(n21), .A2(n487), .B1(n26), .B2(n488), .ZN(n486) );
  OAI221_X1 U397 ( .B1(n202), .B2(n10), .C1(n489), .C2(n8), .A(n490), .ZN(
        B[24]) );
  AOI222_X1 U398 ( .A1(n13), .A2(n382), .B1(n458), .B2(n302), .C1(n312), .C2(
        n303), .ZN(n490) );
  OAI221_X1 U399 ( .B1(n491), .B2(n18), .C1(n492), .C2(n59), .A(n493), .ZN(
        n303) );
  AOI22_X1 U400 ( .A1(n21), .A2(n494), .B1(n26), .B2(n495), .ZN(n493) );
  OAI22_X1 U401 ( .A1(SH[4]), .A2(n245), .B1(n244), .B2(n464), .ZN(n302) );
  INV_X1 U402 ( .A(n381), .ZN(n245) );
  OAI221_X1 U403 ( .B1(n496), .B2(n18), .C1(n497), .C2(n59), .A(n498), .ZN(
        n381) );
  AOI22_X1 U404 ( .A1(n23), .A2(n499), .B1(n27), .B2(n500), .ZN(n498) );
  OAI221_X1 U405 ( .B1(n501), .B2(n18), .C1(n502), .C2(n59), .A(n503), .ZN(
        n382) );
  AOI22_X1 U406 ( .A1(n21), .A2(n504), .B1(n26), .B2(n505), .ZN(n503) );
  INV_X1 U407 ( .A(n506), .ZN(n502) );
  INV_X1 U408 ( .A(n198), .ZN(n489) );
  OAI221_X1 U409 ( .B1(n507), .B2(n18), .C1(n508), .C2(n59), .A(n509), .ZN(
        n198) );
  AOI22_X1 U410 ( .A1(n22), .A2(n510), .B1(n26), .B2(n511), .ZN(n509) );
  INV_X1 U411 ( .A(n512), .ZN(n507) );
  AOI221_X1 U412 ( .B1(n513), .B2(n17), .C1(n514), .C2(n56), .A(n515), .ZN(
        n202) );
  INV_X1 U413 ( .A(n516), .ZN(n515) );
  AOI22_X1 U414 ( .A1(n21), .A2(n517), .B1(n26), .B2(n518), .ZN(n516) );
  OAI221_X1 U415 ( .B1(n230), .B2(n9), .C1(n519), .C2(n8), .A(n520), .ZN(B[23]) );
  AOI222_X1 U416 ( .A1(n13), .A2(n521), .B1(n458), .B2(n304), .C1(n312), .C2(
        n305), .ZN(n520) );
  OAI221_X1 U417 ( .B1(n522), .B2(n18), .C1(n523), .C2(n59), .A(n524), .ZN(
        n305) );
  AOI22_X1 U418 ( .A1(n22), .A2(n525), .B1(n28), .B2(n526), .ZN(n524) );
  OAI22_X1 U419 ( .A1(SH[4]), .A2(n248), .B1(n247), .B2(n464), .ZN(n304) );
  AOI221_X1 U420 ( .B1(n527), .B2(n15), .C1(n528), .C2(n56), .A(n529), .ZN(
        n248) );
  INV_X1 U421 ( .A(n530), .ZN(n529) );
  AOI22_X1 U422 ( .A1(n394), .A2(n531), .B1(n25), .B2(n532), .ZN(n530) );
  INV_X1 U423 ( .A(n229), .ZN(n521) );
  AOI221_X1 U424 ( .B1(n533), .B2(n15), .C1(n534), .C2(n56), .A(n535), .ZN(
        n229) );
  INV_X1 U425 ( .A(n536), .ZN(n535) );
  AOI22_X1 U426 ( .A1(n21), .A2(n537), .B1(n25), .B2(n538), .ZN(n536) );
  INV_X1 U427 ( .A(n226), .ZN(n519) );
  OAI221_X1 U428 ( .B1(n539), .B2(n18), .C1(n540), .C2(n59), .A(n541), .ZN(
        n226) );
  AOI22_X1 U429 ( .A1(n21), .A2(n542), .B1(n28), .B2(n543), .ZN(n541) );
  AOI221_X1 U430 ( .B1(n544), .B2(n17), .C1(n545), .C2(n57), .A(n546), .ZN(
        n230) );
  INV_X1 U431 ( .A(n547), .ZN(n546) );
  AOI22_X1 U432 ( .A1(n21), .A2(n548), .B1(n28), .B2(n549), .ZN(n547) );
  OAI221_X1 U433 ( .B1(n261), .B2(n10), .C1(n550), .C2(n8), .A(n551), .ZN(
        B[22]) );
  AOI222_X1 U434 ( .A1(n13), .A2(n552), .B1(n458), .B2(n306), .C1(n312), .C2(
        n307), .ZN(n551) );
  OAI221_X1 U435 ( .B1(n553), .B2(n18), .C1(n554), .C2(n59), .A(n555), .ZN(
        n307) );
  AOI22_X1 U436 ( .A1(n20), .A2(n556), .B1(n28), .B2(n557), .ZN(n555) );
  OAI22_X1 U437 ( .A1(SH[4]), .A2(n264), .B1(n263), .B2(n464), .ZN(n306) );
  NAND2_X1 U438 ( .A1(n409), .A2(SH[4]), .ZN(n464) );
  AOI221_X1 U439 ( .B1(n558), .B2(n15), .C1(n559), .C2(n409), .A(n560), .ZN(
        n264) );
  INV_X1 U440 ( .A(n561), .ZN(n560) );
  AOI22_X1 U441 ( .A1(n394), .A2(n562), .B1(n25), .B2(n563), .ZN(n561) );
  INV_X1 U442 ( .A(n260), .ZN(n552) );
  AOI221_X1 U443 ( .B1(n564), .B2(n15), .C1(n565), .C2(n57), .A(n566), .ZN(
        n260) );
  INV_X1 U444 ( .A(n567), .ZN(n566) );
  AOI22_X1 U445 ( .A1(n20), .A2(n568), .B1(n25), .B2(n569), .ZN(n567) );
  INV_X1 U446 ( .A(n258), .ZN(n550) );
  OAI221_X1 U447 ( .B1(n570), .B2(n18), .C1(n571), .C2(n58), .A(n572), .ZN(
        n258) );
  AOI22_X1 U448 ( .A1(n21), .A2(n573), .B1(n26), .B2(n574), .ZN(n572) );
  AOI221_X1 U449 ( .B1(n575), .B2(n17), .C1(n576), .C2(n57), .A(n577), .ZN(
        n261) );
  INV_X1 U450 ( .A(n578), .ZN(n577) );
  AOI22_X1 U451 ( .A1(n21), .A2(n579), .B1(n26), .B2(n580), .ZN(n578) );
  OAI221_X1 U452 ( .B1(n290), .B2(n9), .C1(n581), .C2(n8), .A(n582), .ZN(B[21]) );
  AOI222_X1 U453 ( .A1(n13), .A2(n583), .B1(n458), .B2(n584), .C1(n312), .C2(
        n308), .ZN(n582) );
  OAI221_X1 U454 ( .B1(n460), .B2(n18), .C1(n585), .C2(n59), .A(n586), .ZN(
        n308) );
  AOI22_X1 U455 ( .A1(n20), .A2(n463), .B1(n28), .B2(n587), .ZN(n586) );
  INV_X1 U456 ( .A(n475), .ZN(n585) );
  INV_X1 U457 ( .A(n588), .ZN(n460) );
  INV_X1 U458 ( .A(n208), .ZN(n584) );
  MUX2_X1 U459 ( .A(n292), .B(n294), .S(n392), .Z(n208) );
  AOI221_X1 U460 ( .B1(n466), .B2(n16), .C1(n462), .C2(n57), .A(n589), .ZN(
        n294) );
  INV_X1 U461 ( .A(n590), .ZN(n589) );
  AOI22_X1 U462 ( .A1(n20), .A2(n470), .B1(n26), .B2(n465), .ZN(n590) );
  AND2_X1 U463 ( .A1(n376), .A2(n266), .ZN(n458) );
  INV_X1 U464 ( .A(n289), .ZN(n583) );
  AOI221_X1 U465 ( .B1(n472), .B2(n16), .C1(n487), .C2(n57), .A(n591), .ZN(
        n289) );
  INV_X1 U466 ( .A(n592), .ZN(n591) );
  AOI22_X1 U467 ( .A1(n20), .A2(n476), .B1(n26), .B2(n471), .ZN(n592) );
  INV_X1 U468 ( .A(n287), .ZN(n581) );
  OAI221_X1 U469 ( .B1(n478), .B2(n18), .C1(n169), .C2(n59), .A(n593), .ZN(
        n287) );
  AOI22_X1 U470 ( .A1(n20), .A2(n481), .B1(n26), .B2(n482), .ZN(n593) );
  AOI221_X1 U471 ( .B1(n484), .B2(n17), .C1(n480), .C2(n57), .A(n594), .ZN(
        n290) );
  INV_X1 U472 ( .A(n595), .ZN(n594) );
  AOI22_X1 U473 ( .A1(n20), .A2(n488), .B1(n26), .B2(n483), .ZN(n595) );
  OAI221_X1 U474 ( .B1(n333), .B2(n10), .C1(n596), .C2(n8), .A(n597), .ZN(
        B[20]) );
  AOI222_X1 U475 ( .A1(n13), .A2(n598), .B1(n376), .B2(n209), .C1(n312), .C2(
        n337), .ZN(n597) );
  OAI221_X1 U476 ( .B1(n492), .B2(n18), .C1(n599), .C2(n59), .A(n600), .ZN(
        n337) );
  AOI22_X1 U477 ( .A1(n20), .A2(n495), .B1(n26), .B2(n601), .ZN(n600) );
  INV_X1 U478 ( .A(n602), .ZN(n492) );
  OAI22_X1 U479 ( .A1(n334), .A2(n242), .B1(n335), .B2(n238), .ZN(n209) );
  INV_X1 U480 ( .A(n314), .ZN(n335) );
  OAI221_X1 U481 ( .B1(n497), .B2(n18), .C1(n603), .C2(n59), .A(n604), .ZN(
        n314) );
  AOI22_X1 U482 ( .A1(n20), .A2(n500), .B1(n26), .B2(n605), .ZN(n604) );
  INV_X1 U483 ( .A(n606), .ZN(n497) );
  INV_X1 U484 ( .A(n310), .ZN(n598) );
  AOI221_X1 U485 ( .B1(n506), .B2(n16), .C1(n517), .C2(n57), .A(n607), .ZN(
        n310) );
  INV_X1 U486 ( .A(n608), .ZN(n607) );
  AOI22_X1 U487 ( .A1(n20), .A2(n505), .B1(n26), .B2(n609), .ZN(n608) );
  INV_X1 U488 ( .A(n331), .ZN(n596) );
  OAI221_X1 U489 ( .B1(n508), .B2(n18), .C1(n197), .C2(n59), .A(n610), .ZN(
        n331) );
  AOI22_X1 U490 ( .A1(n20), .A2(n511), .B1(n28), .B2(n512), .ZN(n610) );
  AOI221_X1 U491 ( .B1(n514), .B2(n17), .C1(n510), .C2(n57), .A(n611), .ZN(
        n333) );
  INV_X1 U492 ( .A(n612), .ZN(n611) );
  AOI22_X1 U493 ( .A1(n20), .A2(n518), .B1(n28), .B2(n513), .ZN(n612) );
  OAI221_X1 U494 ( .B1(n271), .B2(n383), .C1(n339), .C2(n11), .A(n613), .ZN(
        B[1]) );
  AOI22_X1 U495 ( .A1(n14), .A2(n614), .B1(n386), .B2(n615), .ZN(n613) );
  OAI21_X1 U496 ( .B1(n616), .B2(n265), .A(n617), .ZN(n615) );
  MUX2_X1 U497 ( .A(n618), .B(n619), .S(n392), .Z(n617) );
  AOI222_X1 U498 ( .A1(n15), .A2(n286), .B1(n21), .B2(n163), .C1(n25), .C2(
        n165), .ZN(n619) );
  OAI221_X1 U499 ( .B1(n30), .B2(n157), .C1(n36), .C2(n158), .A(n620), .ZN(
        n165) );
  AOI22_X1 U500 ( .A1(A[12]), .A2(n42), .B1(A[11]), .B2(n47), .ZN(n620) );
  OAI221_X1 U501 ( .B1(n30), .B2(n64), .C1(n36), .C2(n63), .A(n621), .ZN(n286)
         );
  AOI22_X1 U502 ( .A1(A[8]), .A2(n42), .B1(A[7]), .B2(n47), .ZN(n621) );
  AOI221_X1 U503 ( .B1(A[4]), .B2(n42), .C1(A[3]), .C2(n47), .A(n622), .ZN(
        n616) );
  INV_X1 U504 ( .A(n623), .ZN(n622) );
  AOI22_X1 U505 ( .A1(n41), .A2(A[1]), .B1(n35), .B2(A[2]), .ZN(n623) );
  INV_X1 U506 ( .A(n418), .ZN(n614) );
  AOI222_X1 U507 ( .A1(n420), .A2(n400), .B1(n341), .B2(n336), .C1(n342), .C2(
        n401), .ZN(n271) );
  INV_X1 U508 ( .A(n338), .ZN(n420) );
  OAI221_X1 U509 ( .B1(n398), .B2(n9), .C1(n390), .C2(n8), .A(n624), .ZN(B[19]) );
  INV_X1 U510 ( .A(n625), .ZN(n624) );
  OAI222_X1 U511 ( .A1(n4), .A2(n316), .B1(n383), .B2(n211), .C1(n11), .C2(
        n315), .ZN(n625) );
  INV_X1 U512 ( .A(n399), .ZN(n315) );
  OAI221_X1 U513 ( .B1(n523), .B2(n18), .C1(n626), .C2(n59), .A(n627), .ZN(
        n399) );
  AOI22_X1 U514 ( .A1(n20), .A2(n526), .B1(n26), .B2(n628), .ZN(n627) );
  INV_X1 U515 ( .A(n629), .ZN(n523) );
  AOI22_X1 U516 ( .A1(n318), .A2(n401), .B1(n319), .B2(n400), .ZN(n211) );
  OAI221_X1 U517 ( .B1(n630), .B2(n18), .C1(n631), .C2(n59), .A(n632), .ZN(
        n319) );
  AOI22_X1 U518 ( .A1(n20), .A2(n532), .B1(n26), .B2(n527), .ZN(n632) );
  INV_X1 U519 ( .A(n528), .ZN(n630) );
  INV_X1 U520 ( .A(n180), .ZN(n318) );
  AOI22_X1 U521 ( .A1(n531), .A2(n409), .B1(n403), .B2(n16), .ZN(n180) );
  AOI221_X1 U522 ( .B1(n534), .B2(n17), .C1(n548), .C2(n57), .A(n633), .ZN(
        n316) );
  INV_X1 U523 ( .A(n634), .ZN(n633) );
  AOI22_X1 U524 ( .A1(n21), .A2(n538), .B1(n26), .B2(n533), .ZN(n634) );
  INV_X1 U525 ( .A(n635), .ZN(n390) );
  OAI221_X1 U526 ( .B1(n540), .B2(n18), .C1(n636), .C2(n59), .A(n637), .ZN(
        n635) );
  AOI22_X1 U527 ( .A1(n21), .A2(n543), .B1(n28), .B2(n638), .ZN(n637) );
  AOI221_X1 U528 ( .B1(n545), .B2(n16), .C1(n542), .C2(n57), .A(n639), .ZN(
        n398) );
  INV_X1 U529 ( .A(n640), .ZN(n639) );
  AOI22_X1 U530 ( .A1(n21), .A2(n549), .B1(n26), .B2(n544), .ZN(n640) );
  OAI221_X1 U531 ( .B1(n415), .B2(n10), .C1(n439), .C2(n8), .A(n641), .ZN(
        B[18]) );
  INV_X1 U532 ( .A(n642), .ZN(n641) );
  OAI222_X1 U533 ( .A1(n4), .A2(n321), .B1(n383), .B2(n213), .C1(n11), .C2(
        n320), .ZN(n642) );
  INV_X1 U534 ( .A(n417), .ZN(n320) );
  OAI221_X1 U535 ( .B1(n554), .B2(n18), .C1(n643), .C2(n59), .A(n644), .ZN(
        n417) );
  AOI22_X1 U536 ( .A1(n21), .A2(n557), .B1(n26), .B2(n645), .ZN(n644) );
  INV_X1 U537 ( .A(n568), .ZN(n643) );
  INV_X1 U538 ( .A(n646), .ZN(n554) );
  AOI22_X1 U539 ( .A1(n323), .A2(n401), .B1(n324), .B2(n400), .ZN(n213) );
  OAI221_X1 U540 ( .B1(n647), .B2(n18), .C1(n648), .C2(n59), .A(n649), .ZN(
        n324) );
  AOI22_X1 U541 ( .A1(n21), .A2(n563), .B1(n26), .B2(n558), .ZN(n649) );
  INV_X1 U542 ( .A(n559), .ZN(n647) );
  INV_X1 U543 ( .A(n182), .ZN(n323) );
  AOI22_X1 U544 ( .A1(n562), .A2(n409), .B1(n406), .B2(n16), .ZN(n182) );
  AOI221_X1 U545 ( .B1(n565), .B2(n16), .C1(n579), .C2(n57), .A(n650), .ZN(
        n321) );
  INV_X1 U546 ( .A(n651), .ZN(n650) );
  AOI22_X1 U547 ( .A1(n21), .A2(n569), .B1(n26), .B2(n564), .ZN(n651) );
  INV_X1 U548 ( .A(n652), .ZN(n439) );
  OAI221_X1 U549 ( .B1(n571), .B2(n18), .C1(n653), .C2(n58), .A(n654), .ZN(
        n652) );
  AOI22_X1 U550 ( .A1(n21), .A2(n574), .B1(n26), .B2(n655), .ZN(n654) );
  AOI221_X1 U551 ( .B1(n576), .B2(n16), .C1(n573), .C2(n57), .A(n656), .ZN(
        n415) );
  INV_X1 U552 ( .A(n657), .ZN(n656) );
  AOI22_X1 U553 ( .A1(n21), .A2(n580), .B1(n26), .B2(n575), .ZN(n657) );
  OAI221_X1 U554 ( .B1(n418), .B2(n10), .C1(n618), .C2(n8), .A(n658), .ZN(
        B[17]) );
  INV_X1 U555 ( .A(n659), .ZN(n658) );
  OAI222_X1 U556 ( .A1(n4), .A2(n339), .B1(n383), .B2(n214), .C1(n11), .C2(
        n338), .ZN(n659) );
  AOI221_X1 U557 ( .B1(n475), .B2(n16), .C1(n476), .C2(n57), .A(n660), .ZN(
        n338) );
  INV_X1 U558 ( .A(n661), .ZN(n660) );
  AOI22_X1 U559 ( .A1(n21), .A2(n587), .B1(n26), .B2(n588), .ZN(n661) );
  AOI22_X1 U560 ( .A1(n341), .A2(n401), .B1(n342), .B2(n400), .ZN(n214) );
  OAI221_X1 U561 ( .B1(n662), .B2(n18), .C1(n663), .C2(n58), .A(n664), .ZN(
        n342) );
  AOI22_X1 U562 ( .A1(n21), .A2(n465), .B1(n26), .B2(n466), .ZN(n664) );
  INV_X1 U563 ( .A(n462), .ZN(n662) );
  INV_X1 U564 ( .A(n183), .ZN(n341) );
  AOI222_X1 U565 ( .A1(n469), .A2(n15), .B1(n25), .B2(n665), .C1(n470), .C2(
        n56), .ZN(n183) );
  AOI221_X1 U566 ( .B1(n487), .B2(n16), .C1(n488), .C2(n57), .A(n666), .ZN(
        n339) );
  INV_X1 U567 ( .A(n667), .ZN(n666) );
  AOI22_X1 U568 ( .A1(n21), .A2(n471), .B1(n26), .B2(n472), .ZN(n667) );
  INV_X1 U569 ( .A(n668), .ZN(n618) );
  OAI221_X1 U570 ( .B1(n169), .B2(n18), .C1(n167), .C2(n58), .A(n669), .ZN(
        n668) );
  AOI22_X1 U571 ( .A1(n21), .A2(n482), .B1(n26), .B2(n670), .ZN(n669) );
  INV_X1 U572 ( .A(n283), .ZN(n167) );
  AOI221_X1 U573 ( .B1(n480), .B2(n16), .C1(n481), .C2(n57), .A(n671), .ZN(
        n418) );
  INV_X1 U574 ( .A(n672), .ZN(n671) );
  AOI22_X1 U575 ( .A1(n21), .A2(n483), .B1(n26), .B2(n484), .ZN(n672) );
  OAI221_X1 U576 ( .B1(n421), .B2(n9), .C1(n673), .C2(n8), .A(n674), .ZN(B[16]) );
  INV_X1 U577 ( .A(n675), .ZN(n674) );
  OAI222_X1 U578 ( .A1(n4), .A2(n344), .B1(n383), .B2(n215), .C1(n11), .C2(
        n343), .ZN(n675) );
  INV_X1 U579 ( .A(n423), .ZN(n343) );
  AOI22_X1 U580 ( .A1(n346), .A2(n401), .B1(n347), .B2(n400), .ZN(n215) );
  AOI21_X1 U581 ( .B1(n676), .B2(n677), .A(SH[8]), .ZN(B[15]) );
  AOI221_X1 U582 ( .B1(n162), .B2(n219), .C1(n164), .C2(n221), .A(n678), .ZN(
        n677) );
  OAI22_X1 U583 ( .A1(n540), .A2(n168), .B1(n539), .B2(n170), .ZN(n678) );
  INV_X1 U584 ( .A(n638), .ZN(n539) );
  INV_X1 U585 ( .A(n636), .ZN(n219) );
  AOI221_X1 U586 ( .B1(n171), .B2(n679), .C1(n231), .C2(n174), .A(n680), .ZN(
        n676) );
  OAI22_X1 U587 ( .A1(n274), .A2(n177), .B1(n350), .B2(n179), .ZN(n680) );
  AOI221_X1 U588 ( .B1(n548), .B2(n16), .C1(n549), .C2(n57), .A(n681), .ZN(
        n350) );
  INV_X1 U589 ( .A(n682), .ZN(n681) );
  AOI22_X1 U590 ( .A1(n20), .A2(n533), .B1(n26), .B2(n534), .ZN(n682) );
  INV_X1 U591 ( .A(n426), .ZN(n274) );
  OAI221_X1 U592 ( .B1(n626), .B2(n18), .C1(n683), .C2(n58), .A(n684), .ZN(
        n426) );
  AOI22_X1 U593 ( .A1(n20), .A2(n628), .B1(n27), .B2(n629), .ZN(n684) );
  INV_X1 U594 ( .A(n538), .ZN(n683) );
  INV_X1 U595 ( .A(n537), .ZN(n626) );
  OAI22_X1 U596 ( .A1(n185), .A2(n242), .B1(n273), .B2(n238), .ZN(n231) );
  INV_X1 U597 ( .A(n427), .ZN(n273) );
  OAI221_X1 U598 ( .B1(n631), .B2(n19), .C1(n685), .C2(n58), .A(n686), .ZN(
        n427) );
  AOI22_X1 U599 ( .A1(n20), .A2(n527), .B1(n27), .B2(n528), .ZN(n686) );
  INV_X1 U600 ( .A(n525), .ZN(n631) );
  AOI222_X1 U601 ( .A1(n531), .A2(n15), .B1(n403), .B2(n25), .C1(n532), .C2(
        n56), .ZN(n185) );
  INV_X1 U602 ( .A(n424), .ZN(n679) );
  AOI221_X1 U603 ( .B1(n542), .B2(n16), .C1(n543), .C2(n57), .A(n687), .ZN(
        n424) );
  INV_X1 U604 ( .A(n688), .ZN(n687) );
  AOI22_X1 U605 ( .A1(n21), .A2(n544), .B1(n27), .B2(n545), .ZN(n688) );
  AOI21_X1 U606 ( .B1(n689), .B2(n690), .A(SH[8]), .ZN(B[14]) );
  AOI221_X1 U607 ( .B1(n162), .B2(n252), .C1(n164), .C2(n253), .A(n691), .ZN(
        n690) );
  OAI22_X1 U608 ( .A1(n571), .A2(n168), .B1(n570), .B2(n170), .ZN(n691) );
  INV_X1 U609 ( .A(n655), .ZN(n570) );
  AOI221_X1 U610 ( .B1(n171), .B2(n692), .C1(n232), .C2(n174), .A(n693), .ZN(
        n689) );
  OAI22_X1 U611 ( .A1(n276), .A2(n177), .B1(n353), .B2(n179), .ZN(n693) );
  AOI221_X1 U612 ( .B1(n579), .B2(n17), .C1(n580), .C2(n57), .A(n694), .ZN(
        n353) );
  INV_X1 U613 ( .A(n695), .ZN(n694) );
  AOI22_X1 U614 ( .A1(n20), .A2(n564), .B1(n27), .B2(n565), .ZN(n695) );
  AOI221_X1 U615 ( .B1(n568), .B2(n17), .C1(n569), .C2(n57), .A(n696), .ZN(
        n276) );
  INV_X1 U616 ( .A(n697), .ZN(n696) );
  AOI22_X1 U617 ( .A1(n20), .A2(n645), .B1(n27), .B2(n646), .ZN(n697) );
  OAI22_X1 U618 ( .A1(n186), .A2(n242), .B1(n275), .B2(n238), .ZN(n232) );
  INV_X1 U619 ( .A(n432), .ZN(n275) );
  OAI221_X1 U620 ( .B1(n648), .B2(n19), .C1(n698), .C2(n58), .A(n699), .ZN(
        n432) );
  AOI22_X1 U621 ( .A1(n20), .A2(n558), .B1(n27), .B2(n559), .ZN(n699) );
  INV_X1 U622 ( .A(n556), .ZN(n648) );
  AOI222_X1 U623 ( .A1(n562), .A2(n15), .B1(n406), .B2(n25), .C1(n563), .C2(
        n56), .ZN(n186) );
  INV_X1 U624 ( .A(n429), .ZN(n692) );
  AOI221_X1 U625 ( .B1(n573), .B2(n17), .C1(n574), .C2(n57), .A(n700), .ZN(
        n429) );
  INV_X1 U626 ( .A(n701), .ZN(n700) );
  AOI22_X1 U627 ( .A1(n21), .A2(n575), .B1(n27), .B2(n576), .ZN(n701) );
  AOI21_X1 U628 ( .B1(n702), .B2(n703), .A(SH[8]), .ZN(B[13]) );
  AOI221_X1 U629 ( .B1(n162), .B2(n283), .C1(n164), .C2(n163), .A(n704), .ZN(
        n703) );
  OAI22_X1 U630 ( .A1(n169), .A2(n168), .B1(n478), .B2(n170), .ZN(n704) );
  INV_X1 U631 ( .A(n670), .ZN(n478) );
  OAI221_X1 U632 ( .B1(n29), .B2(n155), .C1(n36), .C2(n138), .A(n705), .ZN(
        n670) );
  AOI22_X1 U633 ( .A1(A[28]), .A2(n42), .B1(A[27]), .B2(n47), .ZN(n705) );
  AOI221_X1 U634 ( .B1(n35), .B2(A[22]), .C1(n41), .C2(A[21]), .A(n706), .ZN(
        n169) );
  OAI22_X1 U635 ( .A1(n137), .A2(n1), .B1(n139), .B2(n54), .ZN(n706) );
  OAI221_X1 U636 ( .B1(n30), .B2(n130), .C1(n36), .C2(n129), .A(n707), .ZN(
        n163) );
  AOI22_X1 U637 ( .A1(A[16]), .A2(n42), .B1(A[15]), .B2(n47), .ZN(n707) );
  OAI221_X1 U638 ( .B1(n30), .B2(n156), .C1(n36), .C2(n132), .A(n708), .ZN(
        n283) );
  AOI22_X1 U639 ( .A1(A[20]), .A2(n42), .B1(A[19]), .B2(n47), .ZN(n708) );
  AOI221_X1 U640 ( .B1(n171), .B2(n709), .C1(n233), .C2(n174), .A(n710), .ZN(
        n702) );
  OAI22_X1 U641 ( .A1(n278), .A2(n177), .B1(n358), .B2(n179), .ZN(n710) );
  AOI221_X1 U642 ( .B1(n488), .B2(n17), .C1(n483), .C2(n57), .A(n711), .ZN(
        n358) );
  INV_X1 U643 ( .A(n712), .ZN(n711) );
  AOI22_X1 U644 ( .A1(n21), .A2(n472), .B1(n27), .B2(n487), .ZN(n712) );
  OAI221_X1 U645 ( .B1(n30), .B2(n82), .C1(n36), .C2(n81), .A(n713), .ZN(n487)
         );
  AOI22_X1 U646 ( .A1(A[56]), .A2(n42), .B1(A[55]), .B2(n47), .ZN(n713) );
  OAI221_X1 U647 ( .B1(n30), .B2(n115), .C1(n36), .C2(n84), .A(n714), .ZN(n472) );
  AOI22_X1 U648 ( .A1(A[60]), .A2(n42), .B1(A[59]), .B2(n48), .ZN(n714) );
  OAI221_X1 U649 ( .B1(n30), .B2(n124), .C1(n36), .C2(n123), .A(n715), .ZN(
        n483) );
  AOI22_X1 U650 ( .A1(A[48]), .A2(n45), .B1(A[47]), .B2(n48), .ZN(n715) );
  OAI221_X1 U651 ( .B1(n29), .B2(n120), .C1(n37), .C2(n80), .A(n716), .ZN(n488) );
  AOI22_X1 U652 ( .A1(A[52]), .A2(n45), .B1(A[51]), .B2(n48), .ZN(n716) );
  AOI221_X1 U653 ( .B1(n476), .B2(n17), .C1(n471), .C2(n57), .A(n717), .ZN(
        n278) );
  INV_X1 U654 ( .A(n718), .ZN(n717) );
  AOI22_X1 U655 ( .A1(n20), .A2(n588), .B1(n27), .B2(n475), .ZN(n718) );
  OAI221_X1 U656 ( .B1(n29), .B2(n110), .C1(n37), .C2(n109), .A(n719), .ZN(
        n475) );
  AOI22_X1 U657 ( .A1(A[72]), .A2(n45), .B1(A[71]), .B2(n48), .ZN(n719) );
  OAI221_X1 U658 ( .B1(n29), .B2(n118), .C1(n37), .C2(n112), .A(n720), .ZN(
        n588) );
  AOI22_X1 U659 ( .A1(A[76]), .A2(n42), .B1(A[75]), .B2(n48), .ZN(n720) );
  OAI221_X1 U660 ( .B1(n29), .B2(n103), .C1(n37), .C2(n102), .A(n721), .ZN(
        n471) );
  AOI22_X1 U661 ( .A1(A[64]), .A2(n45), .B1(A[63]), .B2(n48), .ZN(n721) );
  OAI221_X1 U662 ( .B1(n29), .B2(n116), .C1(n37), .C2(n105), .A(n722), .ZN(
        n476) );
  AOI22_X1 U663 ( .A1(A[68]), .A2(n45), .B1(A[67]), .B2(n48), .ZN(n722) );
  OAI22_X1 U664 ( .A1(n187), .A2(n242), .B1(n277), .B2(n238), .ZN(n233) );
  INV_X1 U665 ( .A(n356), .ZN(n277) );
  OAI221_X1 U666 ( .B1(n663), .B2(n19), .C1(n459), .C2(n59), .A(n723), .ZN(
        n356) );
  AOI22_X1 U667 ( .A1(n22), .A2(n466), .B1(n27), .B2(n462), .ZN(n723) );
  OAI221_X1 U668 ( .B1(n29), .B2(n89), .C1(n37), .C2(n88), .A(n724), .ZN(n462)
         );
  AOI22_X1 U669 ( .A1(A[88]), .A2(n45), .B1(A[87]), .B2(n48), .ZN(n724) );
  OAI221_X1 U670 ( .B1(n29), .B2(n74), .C1(n37), .C2(n91), .A(n725), .ZN(n466)
         );
  AOI22_X1 U671 ( .A1(A[92]), .A2(n45), .B1(A[91]), .B2(n48), .ZN(n725) );
  INV_X1 U672 ( .A(n587), .ZN(n459) );
  OAI221_X1 U673 ( .B1(n29), .B2(n96), .C1(n37), .C2(n95), .A(n726), .ZN(n587)
         );
  AOI22_X1 U674 ( .A1(A[80]), .A2(n45), .B1(A[79]), .B2(n48), .ZN(n726) );
  INV_X1 U675 ( .A(n463), .ZN(n663) );
  OAI221_X1 U676 ( .B1(n29), .B2(n117), .C1(n37), .C2(n98), .A(n727), .ZN(n463) );
  AOI22_X1 U677 ( .A1(A[84]), .A2(n45), .B1(A[83]), .B2(n48), .ZN(n727) );
  AOI222_X1 U678 ( .A1(n465), .A2(n56), .B1(n470), .B2(n16), .C1(n728), .C2(
        n729), .ZN(n187) );
  OAI221_X1 U679 ( .B1(n29), .B2(n79), .C1(n37), .C2(n72), .A(n730), .ZN(n470)
         );
  AOI22_X1 U680 ( .A1(A[100]), .A2(n45), .B1(A[99]), .B2(n48), .ZN(n730) );
  OAI221_X1 U681 ( .B1(n29), .B2(n70), .C1(n37), .C2(n69), .A(n731), .ZN(n465)
         );
  AOI22_X1 U682 ( .A1(A[96]), .A2(n42), .B1(A[95]), .B2(n49), .ZN(n731) );
  INV_X1 U683 ( .A(n443), .ZN(n709) );
  AOI221_X1 U684 ( .B1(n481), .B2(n17), .C1(n482), .C2(n57), .A(n732), .ZN(
        n443) );
  INV_X1 U685 ( .A(n733), .ZN(n732) );
  AOI22_X1 U686 ( .A1(n22), .A2(n484), .B1(n27), .B2(n480), .ZN(n733) );
  OAI221_X1 U687 ( .B1(n29), .B2(n150), .C1(n36), .C2(n149), .A(n734), .ZN(
        n480) );
  AOI22_X1 U688 ( .A1(A[40]), .A2(n43), .B1(A[39]), .B2(n49), .ZN(n734) );
  OAI221_X1 U689 ( .B1(n30), .B2(n159), .C1(n36), .C2(n152), .A(n735), .ZN(
        n484) );
  AOI22_X1 U690 ( .A1(A[44]), .A2(n43), .B1(A[43]), .B2(n49), .ZN(n735) );
  OAI221_X1 U691 ( .B1(n29), .B2(n143), .C1(n37), .C2(n142), .A(n736), .ZN(
        n482) );
  AOI22_X1 U692 ( .A1(A[32]), .A2(n43), .B1(A[31]), .B2(n49), .ZN(n736) );
  OAI221_X1 U693 ( .B1(n29), .B2(n154), .C1(n37), .C2(n145), .A(n737), .ZN(
        n481) );
  AOI22_X1 U694 ( .A1(A[36]), .A2(n43), .B1(A[35]), .B2(n49), .ZN(n737) );
  AOI21_X1 U695 ( .B1(n738), .B2(n739), .A(SH[8]), .ZN(B[12]) );
  AOI221_X1 U696 ( .B1(n162), .B2(n327), .C1(n164), .C2(n193), .A(n740), .ZN(
        n739) );
  OAI22_X1 U697 ( .A1(n197), .A2(n168), .B1(n508), .B2(n170), .ZN(n740) );
  INV_X1 U698 ( .A(n741), .ZN(n508) );
  AOI221_X1 U699 ( .B1(n171), .B2(n742), .C1(n234), .C2(n174), .A(n743), .ZN(
        n738) );
  OAI22_X1 U700 ( .A1(n280), .A2(n177), .B1(n363), .B2(n179), .ZN(n743) );
  AOI221_X1 U701 ( .B1(n518), .B2(n17), .C1(n513), .C2(n57), .A(n744), .ZN(
        n363) );
  INV_X1 U702 ( .A(n745), .ZN(n744) );
  AOI22_X1 U703 ( .A1(n22), .A2(n506), .B1(n28), .B2(n517), .ZN(n745) );
  INV_X1 U704 ( .A(n448), .ZN(n280) );
  OAI221_X1 U705 ( .B1(n746), .B2(n19), .C1(n501), .C2(n59), .A(n747), .ZN(
        n448) );
  AOI22_X1 U706 ( .A1(n22), .A2(n602), .B1(n28), .B2(n504), .ZN(n747) );
  INV_X1 U707 ( .A(n609), .ZN(n501) );
  OAI22_X1 U708 ( .A1(n188), .A2(n242), .B1(n279), .B2(n238), .ZN(n234) );
  INV_X1 U709 ( .A(n361), .ZN(n279) );
  OAI221_X1 U710 ( .B1(n748), .B2(n19), .C1(n491), .C2(n59), .A(n749), .ZN(
        n361) );
  AOI22_X1 U711 ( .A1(n22), .A2(n606), .B1(n28), .B2(n494), .ZN(n749) );
  INV_X1 U712 ( .A(n601), .ZN(n491) );
  INV_X1 U713 ( .A(n360), .ZN(n188) );
  OAI221_X1 U714 ( .B1(n750), .B2(n19), .C1(n496), .C2(n59), .A(n751), .ZN(
        n360) );
  AOI22_X1 U715 ( .A1(n22), .A2(n380), .B1(n28), .B2(n499), .ZN(n751) );
  INV_X1 U716 ( .A(n605), .ZN(n496) );
  INV_X1 U717 ( .A(n500), .ZN(n750) );
  INV_X1 U718 ( .A(n446), .ZN(n742) );
  AOI221_X1 U719 ( .B1(n511), .B2(n17), .C1(n512), .C2(n57), .A(n752), .ZN(
        n446) );
  INV_X1 U720 ( .A(n753), .ZN(n752) );
  AOI22_X1 U721 ( .A1(n22), .A2(n514), .B1(n28), .B2(n510), .ZN(n753) );
  AOI21_X1 U722 ( .B1(n754), .B2(n755), .A(SH[8]), .ZN(B[11]) );
  AOI221_X1 U723 ( .B1(n162), .B2(n221), .C1(n164), .C2(n225), .A(n756), .ZN(
        n755) );
  OAI22_X1 U724 ( .A1(n636), .A2(n168), .B1(n540), .B2(n170), .ZN(n756) );
  AOI221_X1 U725 ( .B1(A[24]), .B2(n35), .C1(A[23]), .C2(n41), .A(n757), .ZN(
        n540) );
  OAI22_X1 U726 ( .A1(n155), .A2(n1), .B1(n138), .B2(n54), .ZN(n757) );
  AOI221_X1 U727 ( .B1(n35), .B2(A[20]), .C1(n41), .C2(A[19]), .A(n758), .ZN(
        n636) );
  OAI22_X1 U728 ( .A1(n136), .A2(n1), .B1(n135), .B2(n54), .ZN(n758) );
  OAI221_X1 U729 ( .B1(n30), .B2(n128), .C1(n36), .C2(n127), .A(n759), .ZN(
        n225) );
  AOI22_X1 U730 ( .A1(A[14]), .A2(n43), .B1(A[13]), .B2(n49), .ZN(n759) );
  OAI221_X1 U731 ( .B1(n30), .B2(n131), .C1(n39), .C2(n133), .A(n760), .ZN(
        n221) );
  AOI22_X1 U732 ( .A1(A[18]), .A2(n43), .B1(A[17]), .B2(n49), .ZN(n760) );
  AOI221_X1 U733 ( .B1(n171), .B2(n761), .C1(n235), .C2(n174), .A(n762), .ZN(
        n754) );
  OAI22_X1 U734 ( .A1(n296), .A2(n177), .B1(n368), .B2(n179), .ZN(n762) );
  AOI221_X1 U735 ( .B1(n549), .B2(n17), .C1(n544), .C2(n57), .A(n763), .ZN(
        n368) );
  INV_X1 U736 ( .A(n764), .ZN(n763) );
  AOI22_X1 U737 ( .A1(n22), .A2(n534), .B1(n28), .B2(n548), .ZN(n764) );
  OAI221_X1 U738 ( .B1(n30), .B2(n114), .C1(n36), .C2(n119), .A(n765), .ZN(
        n548) );
  AOI22_X1 U739 ( .A1(A[54]), .A2(n43), .B1(A[53]), .B2(n49), .ZN(n765) );
  OAI221_X1 U740 ( .B1(n29), .B2(n83), .C1(n37), .C2(n85), .A(n766), .ZN(n534)
         );
  AOI22_X1 U741 ( .A1(A[58]), .A2(n43), .B1(A[57]), .B2(n49), .ZN(n766) );
  OAI221_X1 U742 ( .B1(n29), .B2(n122), .C1(n37), .C2(n121), .A(n767), .ZN(
        n544) );
  AOI22_X1 U743 ( .A1(A[46]), .A2(n43), .B1(A[45]), .B2(n49), .ZN(n767) );
  OAI221_X1 U744 ( .B1(n29), .B2(n125), .C1(n37), .C2(n126), .A(n768), .ZN(
        n549) );
  AOI22_X1 U745 ( .A1(A[50]), .A2(n43), .B1(A[49]), .B2(n49), .ZN(n768) );
  AOI221_X1 U746 ( .B1(n538), .B2(n16), .C1(n533), .C2(n57), .A(n769), .ZN(
        n296) );
  INV_X1 U747 ( .A(n770), .ZN(n769) );
  AOI22_X1 U748 ( .A1(n22), .A2(n629), .B1(n28), .B2(n537), .ZN(n770) );
  OAI221_X1 U749 ( .B1(n30), .B2(n108), .C1(n37), .C2(n107), .A(n771), .ZN(
        n537) );
  AOI22_X1 U750 ( .A1(A[70]), .A2(n43), .B1(A[69]), .B2(n49), .ZN(n771) );
  OAI221_X1 U751 ( .B1(n29), .B2(n111), .C1(n38), .C2(n113), .A(n772), .ZN(
        n629) );
  AOI22_X1 U752 ( .A1(A[74]), .A2(n43), .B1(A[73]), .B2(n47), .ZN(n772) );
  OAI221_X1 U753 ( .B1(n30), .B2(n101), .C1(n38), .C2(n100), .A(n773), .ZN(
        n533) );
  AOI22_X1 U754 ( .A1(A[62]), .A2(n42), .B1(A[61]), .B2(n47), .ZN(n773) );
  OAI221_X1 U755 ( .B1(n30), .B2(n104), .C1(n38), .C2(n106), .A(n774), .ZN(
        n538) );
  AOI22_X1 U756 ( .A1(A[66]), .A2(n45), .B1(A[65]), .B2(n49), .ZN(n774) );
  OAI22_X1 U757 ( .A1(n189), .A2(n242), .B1(n295), .B2(n238), .ZN(n235) );
  INV_X1 U758 ( .A(n366), .ZN(n295) );
  OAI221_X1 U759 ( .B1(n685), .B2(n19), .C1(n522), .C2(n59), .A(n775), .ZN(
        n366) );
  AOI22_X1 U760 ( .A1(n22), .A2(n528), .B1(n28), .B2(n525), .ZN(n775) );
  OAI221_X1 U761 ( .B1(n30), .B2(n87), .C1(n38), .C2(n86), .A(n776), .ZN(n525)
         );
  AOI22_X1 U762 ( .A1(A[86]), .A2(n43), .B1(A[85]), .B2(n47), .ZN(n776) );
  OAI221_X1 U763 ( .B1(n30), .B2(n90), .C1(n38), .C2(n92), .A(n777), .ZN(n528)
         );
  AOI22_X1 U764 ( .A1(A[90]), .A2(n45), .B1(A[89]), .B2(n49), .ZN(n777) );
  INV_X1 U765 ( .A(n628), .ZN(n522) );
  OAI221_X1 U766 ( .B1(n30), .B2(n94), .C1(n38), .C2(n93), .A(n778), .ZN(n628)
         );
  AOI22_X1 U767 ( .A1(A[78]), .A2(n45), .B1(A[77]), .B2(n51), .ZN(n778) );
  INV_X1 U768 ( .A(n526), .ZN(n685) );
  OAI221_X1 U769 ( .B1(n30), .B2(n97), .C1(n38), .C2(n99), .A(n779), .ZN(n526)
         );
  AOI22_X1 U770 ( .A1(A[82]), .A2(n45), .B1(A[81]), .B2(n47), .ZN(n779) );
  AOI221_X1 U771 ( .B1(n532), .B2(n17), .C1(n527), .C2(n57), .A(n780), .ZN(
        n189) );
  INV_X1 U772 ( .A(n781), .ZN(n780) );
  AOI22_X1 U773 ( .A1(n22), .A2(n403), .B1(n28), .B2(n531), .ZN(n781) );
  OAI221_X1 U774 ( .B1(n30), .B2(n78), .C1(n38), .C2(n75), .A(n782), .ZN(n531)
         );
  AOI22_X1 U775 ( .A1(A[102]), .A2(n44), .B1(A[101]), .B2(n51), .ZN(n782) );
  INV_X1 U776 ( .A(n247), .ZN(n403) );
  OAI221_X1 U777 ( .B1(n30), .B2(n68), .C1(n38), .C2(n67), .A(n783), .ZN(n527)
         );
  AOI22_X1 U778 ( .A1(A[94]), .A2(n45), .B1(A[93]), .B2(n48), .ZN(n783) );
  OAI221_X1 U779 ( .B1(n30), .B2(n71), .C1(n38), .C2(n73), .A(n784), .ZN(n532)
         );
  AOI22_X1 U780 ( .A1(A[98]), .A2(n44), .B1(A[97]), .B2(n52), .ZN(n784) );
  INV_X1 U781 ( .A(n449), .ZN(n761) );
  AOI221_X1 U782 ( .B1(n543), .B2(n16), .C1(n638), .C2(n57), .A(n785), .ZN(
        n449) );
  INV_X1 U783 ( .A(n786), .ZN(n785) );
  AOI22_X1 U784 ( .A1(n22), .A2(n545), .B1(n28), .B2(n542), .ZN(n786) );
  OAI221_X1 U785 ( .B1(n30), .B2(n148), .C1(n38), .C2(n147), .A(n787), .ZN(
        n542) );
  AOI22_X1 U786 ( .A1(A[38]), .A2(n45), .B1(A[37]), .B2(n47), .ZN(n787) );
  OAI221_X1 U787 ( .B1(n30), .B2(n151), .C1(n39), .C2(n153), .A(n788), .ZN(
        n545) );
  AOI22_X1 U788 ( .A1(A[42]), .A2(n43), .B1(A[41]), .B2(n47), .ZN(n788) );
  OAI221_X1 U789 ( .B1(n31), .B2(n141), .C1(n39), .C2(n140), .A(n789), .ZN(
        n638) );
  AOI22_X1 U790 ( .A1(A[30]), .A2(n44), .B1(A[29]), .B2(n47), .ZN(n789) );
  OAI221_X1 U791 ( .B1(n31), .B2(n144), .C1(n39), .C2(n146), .A(n790), .ZN(
        n543) );
  AOI22_X1 U792 ( .A1(A[34]), .A2(n44), .B1(A[33]), .B2(n47), .ZN(n790) );
  AOI21_X1 U793 ( .B1(n791), .B2(n792), .A(SH[8]), .ZN(B[10]) );
  AOI221_X1 U794 ( .B1(n162), .B2(n253), .C1(n164), .C2(n257), .A(n793), .ZN(
        n792) );
  OAI22_X1 U795 ( .A1(n653), .A2(n168), .B1(n571), .B2(n170), .ZN(n793) );
  AOI221_X1 U796 ( .B1(A[23]), .B2(n35), .C1(A[22]), .C2(n41), .A(n795), .ZN(
        n571) );
  OAI22_X1 U797 ( .A1(n138), .A2(n1), .B1(n54), .B2(n137), .ZN(n795) );
  INV_X1 U798 ( .A(n252), .ZN(n653) );
  OAI221_X1 U799 ( .B1(n31), .B2(n134), .C1(n39), .C2(n156), .A(n796), .ZN(
        n252) );
  AOI22_X1 U800 ( .A1(A[21]), .A2(n44), .B1(A[20]), .B2(n47), .ZN(n796) );
  OAI221_X1 U801 ( .B1(n31), .B2(n127), .C1(n39), .C2(n157), .A(n797), .ZN(
        n257) );
  AOI22_X1 U802 ( .A1(A[13]), .A2(n44), .B1(A[12]), .B2(n47), .ZN(n797) );
  OAI221_X1 U803 ( .B1(n31), .B2(n133), .C1(n39), .C2(n130), .A(n798), .ZN(
        n253) );
  AOI22_X1 U804 ( .A1(A[17]), .A2(n44), .B1(A[16]), .B2(n47), .ZN(n798) );
  NOR2_X1 U805 ( .A1(n238), .A2(n174), .ZN(n794) );
  AOI221_X1 U806 ( .B1(n171), .B2(n799), .C1(n236), .C2(n174), .A(n800), .ZN(
        n791) );
  OAI22_X1 U807 ( .A1(n298), .A2(n177), .B1(n373), .B2(n179), .ZN(n800) );
  AOI221_X1 U808 ( .B1(n580), .B2(n16), .C1(n575), .C2(n57), .A(n802), .ZN(
        n373) );
  INV_X1 U809 ( .A(n803), .ZN(n802) );
  AOI22_X1 U810 ( .A1(n23), .A2(n565), .B1(n26), .B2(n579), .ZN(n803) );
  OAI221_X1 U811 ( .B1(n31), .B2(n119), .C1(n39), .C2(n120), .A(n804), .ZN(
        n579) );
  AOI22_X1 U812 ( .A1(A[53]), .A2(n44), .B1(A[52]), .B2(n47), .ZN(n804) );
  OAI221_X1 U813 ( .B1(n31), .B2(n85), .C1(n39), .C2(n82), .A(n805), .ZN(n565)
         );
  AOI22_X1 U814 ( .A1(A[57]), .A2(n44), .B1(A[56]), .B2(n47), .ZN(n805) );
  OAI221_X1 U815 ( .B1(n31), .B2(n121), .C1(n39), .C2(n159), .A(n806), .ZN(
        n575) );
  AOI22_X1 U816 ( .A1(A[45]), .A2(n44), .B1(A[44]), .B2(n47), .ZN(n806) );
  OAI221_X1 U817 ( .B1(n31), .B2(n126), .C1(n39), .C2(n124), .A(n807), .ZN(
        n580) );
  AOI22_X1 U818 ( .A1(A[49]), .A2(n44), .B1(A[48]), .B2(n47), .ZN(n807) );
  AOI221_X1 U819 ( .B1(n569), .B2(n17), .C1(n564), .C2(n57), .A(n808), .ZN(
        n298) );
  INV_X1 U820 ( .A(n809), .ZN(n808) );
  AOI22_X1 U821 ( .A1(n23), .A2(n646), .B1(n27), .B2(n568), .ZN(n809) );
  OAI221_X1 U822 ( .B1(n31), .B2(n107), .C1(n39), .C2(n116), .A(n810), .ZN(
        n568) );
  AOI22_X1 U823 ( .A1(A[69]), .A2(n44), .B1(A[68]), .B2(n49), .ZN(n810) );
  OAI221_X1 U824 ( .B1(n30), .B2(n113), .C1(n36), .C2(n110), .A(n811), .ZN(
        n646) );
  AOI22_X1 U825 ( .A1(A[73]), .A2(n44), .B1(A[72]), .B2(n51), .ZN(n811) );
  OAI221_X1 U826 ( .B1(n29), .B2(n100), .C1(n36), .C2(n115), .A(n812), .ZN(
        n564) );
  AOI22_X1 U827 ( .A1(A[61]), .A2(n44), .B1(A[60]), .B2(n50), .ZN(n812) );
  OAI221_X1 U828 ( .B1(n32), .B2(n106), .C1(n40), .C2(n103), .A(n813), .ZN(
        n569) );
  AOI22_X1 U829 ( .A1(A[65]), .A2(n43), .B1(A[64]), .B2(n50), .ZN(n813) );
  OAI22_X1 U830 ( .A1(n190), .A2(n242), .B1(n297), .B2(n238), .ZN(n236) );
  INV_X1 U831 ( .A(n371), .ZN(n297) );
  OAI221_X1 U832 ( .B1(n698), .B2(n19), .C1(n553), .C2(n59), .A(n814), .ZN(
        n371) );
  AOI22_X1 U833 ( .A1(n23), .A2(n559), .B1(n28), .B2(n556), .ZN(n814) );
  OAI221_X1 U834 ( .B1(n30), .B2(n86), .C1(n36), .C2(n117), .A(n815), .ZN(n556) );
  AOI22_X1 U835 ( .A1(A[85]), .A2(n42), .B1(A[84]), .B2(n50), .ZN(n815) );
  OAI221_X1 U836 ( .B1(n29), .B2(n92), .C1(n39), .C2(n89), .A(n816), .ZN(n559)
         );
  AOI22_X1 U837 ( .A1(A[89]), .A2(n46), .B1(A[88]), .B2(n50), .ZN(n816) );
  INV_X1 U838 ( .A(n645), .ZN(n553) );
  OAI221_X1 U839 ( .B1(n29), .B2(n93), .C1(n36), .C2(n118), .A(n817), .ZN(n645) );
  AOI22_X1 U840 ( .A1(A[77]), .A2(n45), .B1(A[76]), .B2(n50), .ZN(n817) );
  INV_X1 U841 ( .A(n557), .ZN(n698) );
  OAI221_X1 U842 ( .B1(n29), .B2(n99), .C1(n37), .C2(n96), .A(n818), .ZN(n557)
         );
  AOI22_X1 U843 ( .A1(A[81]), .A2(n43), .B1(A[80]), .B2(n50), .ZN(n818) );
  AOI221_X1 U844 ( .B1(n563), .B2(n16), .C1(n558), .C2(n57), .A(n819), .ZN(
        n190) );
  INV_X1 U845 ( .A(n820), .ZN(n819) );
  AOI22_X1 U846 ( .A1(n23), .A2(n406), .B1(n28), .B2(n562), .ZN(n820) );
  OAI221_X1 U847 ( .B1(n2), .B2(n75), .C1(n6), .C2(n79), .A(n821), .ZN(n562)
         );
  AOI22_X1 U848 ( .A1(A[101]), .A2(n46), .B1(A[100]), .B2(n50), .ZN(n821) );
  INV_X1 U849 ( .A(n263), .ZN(n406) );
  OAI221_X1 U850 ( .B1(n32), .B2(n67), .C1(n40), .C2(n74), .A(n822), .ZN(n558)
         );
  AOI22_X1 U851 ( .A1(A[93]), .A2(n44), .B1(A[92]), .B2(n50), .ZN(n822) );
  OAI221_X1 U852 ( .B1(n2), .B2(n73), .C1(n6), .C2(n70), .A(n823), .ZN(n563)
         );
  AOI22_X1 U853 ( .A1(A[97]), .A2(n46), .B1(A[96]), .B2(n50), .ZN(n823) );
  INV_X1 U854 ( .A(n452), .ZN(n799) );
  AOI221_X1 U855 ( .B1(n574), .B2(n16), .C1(n655), .C2(n409), .A(n824), .ZN(
        n452) );
  INV_X1 U856 ( .A(n825), .ZN(n824) );
  AOI22_X1 U857 ( .A1(n23), .A2(n576), .B1(n26), .B2(n573), .ZN(n825) );
  OAI221_X1 U858 ( .B1(n30), .B2(n147), .C1(n40), .C2(n154), .A(n826), .ZN(
        n573) );
  AOI22_X1 U859 ( .A1(A[37]), .A2(n42), .B1(A[36]), .B2(n50), .ZN(n826) );
  OAI221_X1 U860 ( .B1(n32), .B2(n153), .C1(n40), .C2(n150), .A(n827), .ZN(
        n576) );
  AOI22_X1 U861 ( .A1(A[41]), .A2(n43), .B1(A[40]), .B2(n50), .ZN(n827) );
  OAI221_X1 U862 ( .B1(n32), .B2(n140), .C1(n40), .C2(n155), .A(n828), .ZN(
        n655) );
  AOI22_X1 U863 ( .A1(A[29]), .A2(n42), .B1(A[28]), .B2(n50), .ZN(n828) );
  OAI221_X1 U864 ( .B1(n32), .B2(n146), .C1(n40), .C2(n143), .A(n829), .ZN(
        n574) );
  AOI22_X1 U865 ( .A1(A[33]), .A2(n43), .B1(A[32]), .B2(n51), .ZN(n829) );
  AND2_X1 U866 ( .A1(n210), .A2(n375), .ZN(B[105]) );
  NOR3_X1 U867 ( .A1(n58), .A2(n238), .A3(n240), .ZN(n375) );
  NOR2_X1 U868 ( .A1(n244), .A2(n830), .ZN(B[104]) );
  NOR2_X1 U869 ( .A1(n247), .A2(n830), .ZN(B[103]) );
  AOI222_X1 U870 ( .A1(n35), .A2(A[104]), .B1(n47), .B2(A[105]), .C1(n41), 
        .C2(A[103]), .ZN(n247) );
  NOR2_X1 U871 ( .A1(n263), .A2(n830), .ZN(B[102]) );
  OR2_X1 U872 ( .A1(n181), .A2(n59), .ZN(n830) );
  AOI221_X1 U873 ( .B1(n35), .B2(A[103]), .C1(n41), .C2(A[102]), .A(n831), 
        .ZN(n263) );
  INV_X1 U874 ( .A(n832), .ZN(n831) );
  AOI22_X1 U875 ( .A1(A[105]), .A2(n45), .B1(A[104]), .B2(n51), .ZN(n832) );
  NOR2_X1 U876 ( .A1(n181), .A2(n292), .ZN(B[101]) );
  NAND2_X1 U877 ( .A1(n833), .A2(n729), .ZN(n292) );
  MUX2_X1 U878 ( .A(n665), .B(n469), .S(n834), .Z(n729) );
  OAI221_X1 U879 ( .B1(n32), .B2(n77), .C1(n40), .C2(n76), .A(n835), .ZN(n469)
         );
  AOI22_X1 U880 ( .A1(A[104]), .A2(n45), .B1(A[103]), .B2(n51), .ZN(n835) );
  INV_X1 U881 ( .A(n240), .ZN(n665) );
  NAND2_X1 U882 ( .A1(A[105]), .A2(n41), .ZN(n240) );
  NOR2_X1 U883 ( .A1(n334), .A2(n8), .ZN(B[100]) );
  NAND2_X1 U884 ( .A1(n386), .A2(n392), .ZN(n181) );
  AOI22_X1 U885 ( .A1(n499), .A2(n409), .B1(n380), .B2(n16), .ZN(n334) );
  OAI221_X1 U886 ( .B1(n272), .B2(n383), .C1(n344), .C2(n11), .A(n836), .ZN(
        B[0]) );
  AOI22_X1 U887 ( .A1(n14), .A2(n837), .B1(n386), .B2(n838), .ZN(n836) );
  OAI21_X1 U888 ( .B1(n839), .B2(n265), .A(n840), .ZN(n838) );
  MUX2_X1 U889 ( .A(n673), .B(n841), .S(n392), .Z(n840) );
  AOI222_X1 U890 ( .A1(n15), .A2(n330), .B1(n21), .B2(n193), .C1(n25), .C2(
        n194), .ZN(n841) );
  OAI221_X1 U891 ( .B1(n32), .B2(n158), .C1(n40), .C2(n66), .A(n842), .ZN(n194) );
  AOI22_X1 U892 ( .A1(A[11]), .A2(n45), .B1(A[10]), .B2(n51), .ZN(n842) );
  OAI221_X1 U893 ( .B1(n32), .B2(n129), .C1(n40), .C2(n128), .A(n843), .ZN(
        n193) );
  AOI22_X1 U894 ( .A1(A[15]), .A2(n45), .B1(A[14]), .B2(n51), .ZN(n843) );
  OAI221_X1 U895 ( .B1(n32), .B2(n63), .C1(n40), .C2(n62), .A(n844), .ZN(n330)
         );
  AOI22_X1 U896 ( .A1(A[7]), .A2(n45), .B1(A[6]), .B2(n51), .ZN(n844) );
  INV_X1 U897 ( .A(n845), .ZN(n673) );
  OAI221_X1 U898 ( .B1(n197), .B2(n19), .C1(n196), .C2(n58), .A(n846), .ZN(
        n845) );
  AOI22_X1 U899 ( .A1(n23), .A2(n512), .B1(n26), .B2(n741), .ZN(n846) );
  OAI221_X1 U900 ( .B1(n32), .B2(n138), .C1(n137), .C2(n36), .A(n847), .ZN(
        n741) );
  AOI22_X1 U901 ( .A1(A[27]), .A2(n45), .B1(A[26]), .B2(n51), .ZN(n847) );
  OAI221_X1 U902 ( .B1(n32), .B2(n142), .C1(n40), .C2(n141), .A(n848), .ZN(
        n512) );
  AOI22_X1 U903 ( .A1(A[31]), .A2(n45), .B1(A[30]), .B2(n51), .ZN(n848) );
  INV_X1 U904 ( .A(n327), .ZN(n196) );
  OAI221_X1 U905 ( .B1(n32), .B2(n132), .C1(n40), .C2(n131), .A(n849), .ZN(
        n327) );
  AOI22_X1 U906 ( .A1(A[19]), .A2(n45), .B1(A[18]), .B2(n51), .ZN(n849) );
  AOI221_X1 U907 ( .B1(n35), .B2(A[21]), .C1(n41), .C2(A[20]), .A(n850), .ZN(
        n197) );
  OAI22_X1 U908 ( .A1(n139), .A2(n1), .B1(n136), .B2(n54), .ZN(n850) );
  NAND2_X1 U909 ( .A1(n409), .A2(n392), .ZN(n265) );
  AOI221_X1 U910 ( .B1(A[1]), .B2(n35), .C1(A[0]), .C2(n41), .A(n851), .ZN(
        n839) );
  OAI22_X1 U911 ( .A1(n54), .A2(n60), .B1(n1), .B2(n61), .ZN(n851) );
  INV_X1 U912 ( .A(n204), .ZN(n386) );
  NAND2_X1 U913 ( .A1(n210), .A2(n266), .ZN(n204) );
  INV_X1 U914 ( .A(n421), .ZN(n837) );
  AOI221_X1 U915 ( .B1(n510), .B2(n16), .C1(n511), .C2(n409), .A(n852), .ZN(
        n421) );
  INV_X1 U916 ( .A(n853), .ZN(n852) );
  AOI22_X1 U917 ( .A1(n23), .A2(n513), .B1(n26), .B2(n514), .ZN(n853) );
  OAI221_X1 U918 ( .B1(n32), .B2(n152), .C1(n40), .C2(n151), .A(n854), .ZN(
        n514) );
  AOI22_X1 U919 ( .A1(A[43]), .A2(n45), .B1(A[42]), .B2(n51), .ZN(n854) );
  OAI221_X1 U920 ( .B1(n30), .B2(n123), .C1(n36), .C2(n122), .A(n855), .ZN(
        n513) );
  AOI22_X1 U921 ( .A1(A[47]), .A2(n45), .B1(A[46]), .B2(n51), .ZN(n855) );
  OAI221_X1 U922 ( .B1(n30), .B2(n145), .C1(n36), .C2(n144), .A(n856), .ZN(
        n511) );
  AOI22_X1 U923 ( .A1(A[35]), .A2(n45), .B1(A[34]), .B2(n51), .ZN(n856) );
  OAI221_X1 U924 ( .B1(n30), .B2(n149), .C1(n36), .C2(n148), .A(n857), .ZN(
        n510) );
  AOI22_X1 U925 ( .A1(A[39]), .A2(n45), .B1(A[38]), .B2(n52), .ZN(n857) );
  NOR2_X1 U926 ( .A1(n299), .A2(n392), .ZN(n312) );
  NAND2_X1 U927 ( .A1(n801), .A2(n858), .ZN(n299) );
  INV_X1 U928 ( .A(SH[8]), .ZN(n858) );
  NOR2_X1 U929 ( .A1(n174), .A2(n266), .ZN(n801) );
  AOI221_X1 U930 ( .B1(n517), .B2(n17), .C1(n518), .C2(n56), .A(n860), .ZN(
        n344) );
  INV_X1 U931 ( .A(n861), .ZN(n860) );
  AOI22_X1 U932 ( .A1(n23), .A2(n609), .B1(n26), .B2(n506), .ZN(n861) );
  OAI221_X1 U933 ( .B1(n30), .B2(n84), .C1(n36), .C2(n83), .A(n862), .ZN(n506)
         );
  AOI22_X1 U934 ( .A1(A[59]), .A2(n43), .B1(A[58]), .B2(n52), .ZN(n862) );
  OAI221_X1 U935 ( .B1(n30), .B2(n102), .C1(n36), .C2(n101), .A(n863), .ZN(
        n609) );
  AOI22_X1 U936 ( .A1(A[63]), .A2(n42), .B1(A[62]), .B2(n52), .ZN(n863) );
  OAI221_X1 U937 ( .B1(n30), .B2(n80), .C1(n36), .C2(n125), .A(n864), .ZN(n518) );
  AOI22_X1 U938 ( .A1(A[51]), .A2(n43), .B1(A[50]), .B2(n52), .ZN(n864) );
  OAI221_X1 U939 ( .B1(n30), .B2(n81), .C1(n36), .C2(n114), .A(n865), .ZN(n517) );
  AOI22_X1 U940 ( .A1(A[55]), .A2(n42), .B1(A[54]), .B2(n52), .ZN(n865) );
  NOR2_X1 U941 ( .A1(n859), .A2(SH[8]), .ZN(n376) );
  NOR2_X1 U942 ( .A1(SH[6]), .A2(SH[7]), .ZN(n859) );
  AOI222_X1 U943 ( .A1(n423), .A2(n400), .B1(n346), .B2(n336), .C1(n347), .C2(
        n401), .ZN(n272) );
  INV_X1 U944 ( .A(n242), .ZN(n401) );
  OAI221_X1 U945 ( .B1(n603), .B2(n19), .C1(n748), .C2(n58), .A(n866), .ZN(
        n347) );
  AOI22_X1 U946 ( .A1(n23), .A2(n605), .B1(n26), .B2(n606), .ZN(n866) );
  OAI221_X1 U947 ( .B1(n29), .B2(n91), .C1(n36), .C2(n90), .A(n867), .ZN(n606)
         );
  AOI22_X1 U948 ( .A1(A[91]), .A2(n46), .B1(A[90]), .B2(n52), .ZN(n867) );
  OAI221_X1 U949 ( .B1(n29), .B2(n69), .C1(n39), .C2(n68), .A(n868), .ZN(n605)
         );
  AOI22_X1 U950 ( .A1(A[95]), .A2(n46), .B1(A[94]), .B2(n52), .ZN(n868) );
  INV_X1 U951 ( .A(n495), .ZN(n748) );
  OAI221_X1 U952 ( .B1(n30), .B2(n98), .C1(n36), .C2(n97), .A(n869), .ZN(n495)
         );
  AOI22_X1 U953 ( .A1(A[83]), .A2(n42), .B1(A[82]), .B2(n52), .ZN(n869) );
  INV_X1 U954 ( .A(n494), .ZN(n603) );
  OAI221_X1 U955 ( .B1(n30), .B2(n88), .C1(n36), .C2(n87), .A(n870), .ZN(n494)
         );
  AOI22_X1 U956 ( .A1(A[87]), .A2(n42), .B1(A[86]), .B2(n52), .ZN(n870) );
  NOR2_X1 U957 ( .A1(SH[4]), .A2(n266), .ZN(n336) );
  INV_X1 U958 ( .A(n184), .ZN(n346) );
  AOI222_X1 U959 ( .A1(n499), .A2(n15), .B1(n380), .B2(n25), .C1(n500), .C2(
        n56), .ZN(n184) );
  OAI221_X1 U960 ( .B1(n29), .B2(n72), .C1(n40), .C2(n71), .A(n871), .ZN(n500)
         );
  AOI22_X1 U961 ( .A1(A[99]), .A2(n46), .B1(A[98]), .B2(n52), .ZN(n871) );
  INV_X1 U962 ( .A(n244), .ZN(n380) );
  AOI22_X1 U963 ( .A1(n41), .A2(A[104]), .B1(n35), .B2(A[105]), .ZN(n244) );
  OAI221_X1 U964 ( .B1(n29), .B2(n76), .C1(n37), .C2(n78), .A(n872), .ZN(n499)
         );
  AOI22_X1 U965 ( .A1(A[103]), .A2(n46), .B1(A[102]), .B2(n52), .ZN(n872) );
  INV_X1 U966 ( .A(n238), .ZN(n400) );
  NOR2_X1 U967 ( .A1(SH[5]), .A2(SH[7]), .ZN(n266) );
  OAI221_X1 U968 ( .B1(n599), .B2(n18), .C1(n746), .C2(n59), .A(n873), .ZN(
        n423) );
  AOI22_X1 U969 ( .A1(n21), .A2(n601), .B1(n26), .B2(n602), .ZN(n873) );
  OAI221_X1 U970 ( .B1(n29), .B2(n112), .C1(n36), .C2(n111), .A(n874), .ZN(
        n602) );
  AOI22_X1 U971 ( .A1(A[75]), .A2(n42), .B1(A[74]), .B2(n52), .ZN(n874) );
  OAI221_X1 U972 ( .B1(n30), .B2(n95), .C1(n39), .C2(n94), .A(n875), .ZN(n601)
         );
  AOI22_X1 U973 ( .A1(A[79]), .A2(n43), .B1(A[78]), .B2(n49), .ZN(n875) );
  NOR2_X1 U974 ( .A1(n834), .A2(n833), .ZN(n394) );
  NOR2_X1 U975 ( .A1(n728), .A2(SH[2]), .ZN(n409) );
  INV_X1 U976 ( .A(n505), .ZN(n746) );
  OAI221_X1 U977 ( .B1(n29), .B2(n105), .C1(n36), .C2(n104), .A(n876), .ZN(
        n505) );
  AOI22_X1 U978 ( .A1(A[67]), .A2(n42), .B1(A[66]), .B2(n47), .ZN(n876) );
  NOR2_X1 U979 ( .A1(n728), .A2(n834), .ZN(n393) );
  INV_X1 U980 ( .A(SH[2]), .ZN(n834) );
  INV_X1 U981 ( .A(n833), .ZN(n728) );
  NOR2_X1 U982 ( .A1(SH[3]), .A2(SH[7]), .ZN(n833) );
  INV_X1 U983 ( .A(n504), .ZN(n599) );
  OAI221_X1 U984 ( .B1(n30), .B2(n109), .C1(n36), .C2(n108), .A(n877), .ZN(
        n504) );
  AOI22_X1 U985 ( .A1(A[71]), .A2(n42), .B1(A[70]), .B2(n47), .ZN(n877) );
  INV_X1 U986 ( .A(SH[0]), .ZN(n879) );
  NOR2_X1 U987 ( .A1(SH[1]), .A2(SH[7]), .ZN(n878) );
endmodule


module fpu_DW01_ash_1 ( A, DATA_TC, SH, SH_TC, B );
  input [117:0] A;
  input [10:0] SH;
  output [117:0] B;
  input DATA_TC, SH_TC;
  wire   \temp_int_SH[4] , \temp_int_SH[3] , \temp_int_SH[0] ,
         \MR_int[1][113] , \ML_int[1][113] , \ML_int[1][112] ,
         \ML_int[1][111] , \ML_int[1][110] , \ML_int[1][109] ,
         \ML_int[1][108] , \ML_int[1][107] , \ML_int[1][106] ,
         \ML_int[1][105] , \ML_int[1][104] , \ML_int[1][103] ,
         \ML_int[1][102] , \ML_int[1][101] , \ML_int[1][100] , \ML_int[1][99] ,
         \ML_int[1][98] , \ML_int[1][97] , \ML_int[1][96] , \ML_int[1][95] ,
         \ML_int[1][94] , \ML_int[1][93] , \ML_int[1][92] , \ML_int[1][91] ,
         \ML_int[1][90] , \ML_int[1][89] , \ML_int[1][88] , \ML_int[1][87] ,
         \ML_int[1][86] , \ML_int[1][85] , \ML_int[1][84] , \ML_int[1][83] ,
         \ML_int[1][82] , \ML_int[1][81] , \ML_int[1][80] , \ML_int[1][79] ,
         \ML_int[1][78] , \ML_int[1][77] , \ML_int[1][76] , \ML_int[1][75] ,
         \ML_int[1][74] , \ML_int[1][73] , \ML_int[1][72] , \ML_int[1][71] ,
         \ML_int[1][70] , \ML_int[1][69] , \ML_int[1][68] , \ML_int[1][67] ,
         \ML_int[1][66] , \ML_int[1][65] , \ML_int[1][64] , \ML_int[1][63] ,
         \ML_int[1][62] , \ML_int[1][61] , \ML_int[1][60] , \ML_int[1][59] ,
         \ML_int[1][58] , \ML_int[1][57] , \ML_int[1][56] , \ML_int[1][55] ,
         \ML_int[1][54] , \ML_int[1][53] , \ML_int[1][52] , \ML_int[1][51] ,
         \ML_int[1][50] , \ML_int[1][49] , \ML_int[1][48] , \ML_int[1][47] ,
         \ML_int[1][46] , \ML_int[1][45] , \ML_int[1][44] , \ML_int[1][43] ,
         \ML_int[1][42] , \ML_int[1][41] , \ML_int[1][40] , \ML_int[1][39] ,
         \ML_int[1][38] , \ML_int[1][37] , \ML_int[1][36] , \ML_int[1][35] ,
         \ML_int[1][34] , \ML_int[1][33] , \ML_int[1][32] , \ML_int[1][31] ,
         \ML_int[1][30] , \ML_int[1][29] , \ML_int[1][28] , \ML_int[1][27] ,
         \ML_int[1][26] , \ML_int[1][25] , \ML_int[1][24] , \ML_int[1][23] ,
         \ML_int[1][22] , \ML_int[1][21] , \ML_int[1][20] , \ML_int[1][19] ,
         \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] , \ML_int[1][15] ,
         \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] , \ML_int[1][11] ,
         \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] , \ML_int[1][7] ,
         \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] , \ML_int[1][3] ,
         \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] , \ML_int[2][114] ,
         \ML_int[2][113] , \ML_int[2][112] , \ML_int[2][111] ,
         \ML_int[2][110] , \ML_int[2][109] , \ML_int[2][108] ,
         \ML_int[2][107] , \ML_int[2][106] , \ML_int[2][105] ,
         \ML_int[2][104] , \ML_int[2][103] , \ML_int[2][102] ,
         \ML_int[2][101] , \ML_int[2][100] , \ML_int[2][99] , \ML_int[2][98] ,
         \ML_int[2][97] , \ML_int[2][96] , \ML_int[2][95] , \ML_int[2][94] ,
         \ML_int[2][93] , \ML_int[2][92] , \ML_int[2][91] , \ML_int[2][90] ,
         \ML_int[2][89] , \ML_int[2][88] , \ML_int[2][87] , \ML_int[2][86] ,
         \ML_int[2][85] , \ML_int[2][84] , \ML_int[2][83] , \ML_int[2][82] ,
         \ML_int[2][81] , \ML_int[2][80] , \ML_int[2][79] , \ML_int[2][78] ,
         \ML_int[2][77] , \ML_int[2][76] , \ML_int[2][75] , \ML_int[2][74] ,
         \ML_int[2][73] , \ML_int[2][72] , \ML_int[2][71] , \ML_int[2][70] ,
         \ML_int[2][69] , \ML_int[2][68] , \ML_int[2][67] , \ML_int[2][66] ,
         \ML_int[2][65] , \ML_int[2][64] , \ML_int[2][63] , \ML_int[2][62] ,
         \ML_int[2][61] , \ML_int[2][60] , \ML_int[2][59] , \ML_int[2][58] ,
         \ML_int[2][57] , \ML_int[2][56] , \ML_int[2][55] , \ML_int[2][54] ,
         \ML_int[2][53] , \ML_int[2][52] , \ML_int[2][51] , \ML_int[2][50] ,
         \ML_int[2][49] , \ML_int[2][48] , \ML_int[2][47] , \ML_int[2][46] ,
         \ML_int[2][45] , \ML_int[2][44] , \ML_int[2][43] , \ML_int[2][42] ,
         \ML_int[2][41] , \ML_int[2][40] , \ML_int[2][39] , \ML_int[2][38] ,
         \ML_int[2][37] , \ML_int[2][36] , \ML_int[2][35] , \ML_int[2][34] ,
         \ML_int[2][33] , \ML_int[2][32] , \ML_int[2][31] , \ML_int[2][30] ,
         \ML_int[2][29] , \ML_int[2][28] , \ML_int[2][27] , \ML_int[2][26] ,
         \ML_int[2][25] , \ML_int[2][24] , \ML_int[2][23] , \ML_int[2][22] ,
         \ML_int[2][21] , \ML_int[2][20] , \ML_int[2][19] , \ML_int[2][18] ,
         \ML_int[2][17] , \ML_int[2][16] , \ML_int[2][15] , \ML_int[2][14] ,
         \ML_int[2][13] , \ML_int[2][12] , \ML_int[2][11] , \ML_int[2][10] ,
         \ML_int[2][9] , \ML_int[2][8] , \ML_int[2][7] , \ML_int[2][6] ,
         \ML_int[2][5] , \ML_int[2][4] , \ML_int[2][3] , \ML_int[2][2] ,
         \ML_int[3][116] , \ML_int[3][115] , \ML_int[3][114] ,
         \ML_int[3][113] , \ML_int[3][112] , \ML_int[3][111] ,
         \ML_int[3][110] , \ML_int[3][109] , \ML_int[3][108] ,
         \ML_int[3][107] , \ML_int[3][106] , \ML_int[3][105] ,
         \ML_int[3][104] , \ML_int[3][103] , \ML_int[3][102] ,
         \ML_int[3][101] , \ML_int[3][100] , \ML_int[3][99] , \ML_int[3][98] ,
         \ML_int[3][97] , \ML_int[3][96] , \ML_int[3][95] , \ML_int[3][94] ,
         \ML_int[3][93] , \ML_int[3][92] , \ML_int[3][91] , \ML_int[3][90] ,
         \ML_int[3][89] , \ML_int[3][88] , \ML_int[3][87] , \ML_int[3][86] ,
         \ML_int[3][85] , \ML_int[3][84] , \ML_int[3][83] , \ML_int[3][82] ,
         \ML_int[3][81] , \ML_int[3][80] , \ML_int[3][79] , \ML_int[3][78] ,
         \ML_int[3][77] , \ML_int[3][76] , \ML_int[3][75] , \ML_int[3][74] ,
         \ML_int[3][73] , \ML_int[3][72] , \ML_int[3][71] , \ML_int[3][70] ,
         \ML_int[3][69] , \ML_int[3][68] , \ML_int[3][67] , \ML_int[3][66] ,
         \ML_int[3][65] , \ML_int[3][64] , \ML_int[3][63] , \ML_int[3][62] ,
         \ML_int[3][61] , \ML_int[3][60] , \ML_int[3][59] , \ML_int[3][58] ,
         \ML_int[3][57] , \ML_int[3][56] , \ML_int[3][55] , \ML_int[3][54] ,
         \ML_int[3][53] , \ML_int[3][52] , \ML_int[3][51] , \ML_int[3][50] ,
         \ML_int[3][49] , \ML_int[3][48] , \ML_int[3][47] , \ML_int[3][46] ,
         \ML_int[3][45] , \ML_int[3][44] , \ML_int[3][43] , \ML_int[3][42] ,
         \ML_int[3][41] , \ML_int[3][40] , \ML_int[3][39] , \ML_int[3][38] ,
         \ML_int[3][37] , \ML_int[3][36] , \ML_int[3][35] , \ML_int[3][34] ,
         \ML_int[3][33] , \ML_int[3][32] , \ML_int[3][31] , \ML_int[3][30] ,
         \ML_int[3][29] , \ML_int[3][28] , \ML_int[3][27] , \ML_int[3][26] ,
         \ML_int[3][25] , \ML_int[3][24] , \ML_int[3][23] , \ML_int[3][22] ,
         \ML_int[3][21] , \ML_int[3][20] , \ML_int[3][19] , \ML_int[3][18] ,
         \ML_int[3][17] , \ML_int[3][16] , \ML_int[3][15] , \ML_int[3][14] ,
         \ML_int[3][13] , \ML_int[3][12] , \ML_int[3][11] , \ML_int[3][10] ,
         \ML_int[3][9] , \ML_int[3][8] , \ML_int[3][7] , \ML_int[3][6] ,
         \ML_int[3][5] , \ML_int[3][4] , \ML_int[4][117] , \ML_int[4][116] ,
         \ML_int[4][115] , \ML_int[4][114] , \ML_int[4][113] ,
         \ML_int[4][112] , \ML_int[4][111] , \ML_int[4][110] ,
         \ML_int[4][109] , \ML_int[4][108] , \ML_int[4][107] ,
         \ML_int[4][101] , \ML_int[4][100] , \ML_int[4][99] , \ML_int[4][98] ,
         \ML_int[4][97] , \ML_int[4][96] , \ML_int[4][95] , \ML_int[4][94] ,
         \ML_int[4][93] , \ML_int[4][92] , \ML_int[4][91] , \ML_int[4][85] ,
         \ML_int[4][84] , \ML_int[4][83] , \ML_int[4][82] , \ML_int[4][81] ,
         \ML_int[4][80] , \ML_int[4][79] , \ML_int[4][78] , \ML_int[4][77] ,
         \ML_int[4][76] , \ML_int[4][75] , \ML_int[4][69] , \ML_int[4][68] ,
         \ML_int[4][67] , \ML_int[4][66] , \ML_int[4][65] , \ML_int[4][64] ,
         \ML_int[4][63] , \ML_int[4][62] , \ML_int[4][61] , \ML_int[4][60] ,
         \ML_int[4][59] , \ML_int[4][53] , \ML_int[4][52] , \ML_int[4][51] ,
         \ML_int[4][50] , \ML_int[4][49] , \ML_int[4][48] , \ML_int[4][47] ,
         \ML_int[4][46] , \ML_int[4][45] , \ML_int[4][44] , \ML_int[4][43] ,
         \ML_int[4][37] , \ML_int[4][36] , \ML_int[4][35] , \ML_int[4][34] ,
         \ML_int[4][33] , \ML_int[4][32] , \ML_int[4][31] , \ML_int[4][30] ,
         \ML_int[4][29] , \ML_int[4][28] , \ML_int[4][27] , \ML_int[4][21] ,
         \ML_int[4][20] , \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] ,
         \ML_int[4][16] , \ML_int[4][15] , \ML_int[4][14] , \ML_int[4][13] ,
         \ML_int[4][12] , \ML_int[4][11] , \ML_int[4][5] , \ML_int[4][4] ,
         \ML_int[4][3] , \ML_int[4][2] , \ML_int[4][1] , \ML_int[4][0] ,
         \ML_int[5][117] , \ML_int[5][116] , \ML_int[5][115] ,
         \ML_int[5][114] , \ML_int[5][113] , \ML_int[5][112] ,
         \ML_int[5][111] , \ML_int[5][110] , \ML_int[5][109] ,
         \ML_int[5][108] , \ML_int[5][107] , \ML_int[5][85] , \ML_int[5][84] ,
         \ML_int[5][83] , \ML_int[5][82] , \ML_int[5][81] , \ML_int[5][80] ,
         \ML_int[5][79] , \ML_int[5][78] , \ML_int[5][77] , \ML_int[5][76] ,
         \ML_int[5][75] , \ML_int[5][53] , \ML_int[5][52] , \ML_int[5][51] ,
         \ML_int[5][50] , \ML_int[5][49] , \ML_int[5][48] , \ML_int[5][47] ,
         \ML_int[5][46] , \ML_int[5][45] , \ML_int[5][44] , \ML_int[5][43] ,
         \ML_int[5][21] , \ML_int[5][20] , \ML_int[5][19] , \ML_int[5][18] ,
         \ML_int[5][17] , \ML_int[5][16] , \ML_int[5][15] , \ML_int[5][14] ,
         \ML_int[5][13] , \ML_int[5][12] , \ML_int[5][11] , \ML_int[6][117] ,
         \ML_int[6][116] , \ML_int[6][115] , \ML_int[6][114] ,
         \ML_int[6][113] , \ML_int[6][112] , \ML_int[6][111] ,
         \ML_int[6][110] , \ML_int[6][109] , \ML_int[6][108] ,
         \ML_int[6][107] , \ML_int[6][53] , \ML_int[6][52] , \ML_int[6][51] ,
         \ML_int[6][50] , \ML_int[6][49] , \ML_int[6][48] , \ML_int[6][47] ,
         \ML_int[6][46] , \ML_int[6][45] , \ML_int[6][44] , \ML_int[6][43] ,
         \ML_int[7][117] , \ML_int[7][116] , \ML_int[7][115] ,
         \ML_int[7][114] , \ML_int[7][113] , \ML_int[7][112] ,
         \ML_int[7][111] , \ML_int[7][110] , \ML_int[7][109] ,
         \ML_int[7][108] , \ML_int[7][107] , \ML_int[8][117] ,
         \ML_int[8][116] , \ML_int[8][115] , \ML_int[8][114] ,
         \ML_int[8][113] , \ML_int[8][112] , \ML_int[8][111] ,
         \ML_int[8][110] , \ML_int[8][109] , \ML_int[8][108] ,
         \ML_int[8][107] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57;
  wire   [6:5] SHMAG;
  assign B[117] = \ML_int[8][117] ;
  assign B[116] = \ML_int[8][116] ;
  assign B[115] = \ML_int[8][115] ;
  assign B[114] = \ML_int[8][114] ;
  assign B[113] = \ML_int[8][113] ;
  assign B[112] = \ML_int[8][112] ;
  assign B[111] = \ML_int[8][111] ;
  assign B[110] = \ML_int[8][110] ;
  assign B[109] = \ML_int[8][109] ;
  assign B[108] = \ML_int[8][108] ;
  assign B[107] = \ML_int[8][107] ;

  MUX2_X2 M1_6_117 ( .A(\ML_int[6][117] ), .B(\ML_int[6][53] ), .S(n42), .Z(
        \ML_int[7][117] ) );
  MUX2_X2 M1_6_116 ( .A(\ML_int[6][116] ), .B(\ML_int[6][52] ), .S(n42), .Z(
        \ML_int[7][116] ) );
  MUX2_X2 M1_6_115 ( .A(\ML_int[6][115] ), .B(\ML_int[6][51] ), .S(n42), .Z(
        \ML_int[7][115] ) );
  MUX2_X2 M1_6_114 ( .A(\ML_int[6][114] ), .B(\ML_int[6][50] ), .S(n42), .Z(
        \ML_int[7][114] ) );
  MUX2_X2 M1_6_113 ( .A(\ML_int[6][113] ), .B(\ML_int[6][49] ), .S(n42), .Z(
        \ML_int[7][113] ) );
  MUX2_X2 M1_6_112 ( .A(\ML_int[6][112] ), .B(\ML_int[6][48] ), .S(n42), .Z(
        \ML_int[7][112] ) );
  MUX2_X2 M1_6_111 ( .A(\ML_int[6][111] ), .B(\ML_int[6][47] ), .S(n42), .Z(
        \ML_int[7][111] ) );
  MUX2_X2 M1_6_110 ( .A(\ML_int[6][110] ), .B(\ML_int[6][46] ), .S(n42), .Z(
        \ML_int[7][110] ) );
  MUX2_X2 M1_6_109 ( .A(\ML_int[6][109] ), .B(\ML_int[6][45] ), .S(n42), .Z(
        \ML_int[7][109] ) );
  MUX2_X2 M1_6_108 ( .A(\ML_int[6][108] ), .B(\ML_int[6][44] ), .S(n42), .Z(
        \ML_int[7][108] ) );
  MUX2_X2 M1_6_107 ( .A(\ML_int[6][107] ), .B(\ML_int[6][43] ), .S(n42), .Z(
        \ML_int[7][107] ) );
  MUX2_X2 M1_5_117 ( .A(\ML_int[5][117] ), .B(\ML_int[5][85] ), .S(n41), .Z(
        \ML_int[6][117] ) );
  MUX2_X2 M1_5_116 ( .A(\ML_int[5][116] ), .B(\ML_int[5][84] ), .S(n41), .Z(
        \ML_int[6][116] ) );
  MUX2_X2 M1_5_115 ( .A(\ML_int[5][115] ), .B(\ML_int[5][83] ), .S(n41), .Z(
        \ML_int[6][115] ) );
  MUX2_X2 M1_5_114 ( .A(\ML_int[5][114] ), .B(\ML_int[5][82] ), .S(n41), .Z(
        \ML_int[6][114] ) );
  MUX2_X2 M1_5_113 ( .A(\ML_int[5][113] ), .B(\ML_int[5][81] ), .S(n41), .Z(
        \ML_int[6][113] ) );
  MUX2_X2 M1_5_112 ( .A(\ML_int[5][112] ), .B(\ML_int[5][80] ), .S(n41), .Z(
        \ML_int[6][112] ) );
  MUX2_X2 M1_5_111 ( .A(\ML_int[5][111] ), .B(\ML_int[5][79] ), .S(n41), .Z(
        \ML_int[6][111] ) );
  MUX2_X2 M1_5_110 ( .A(\ML_int[5][110] ), .B(\ML_int[5][78] ), .S(n41), .Z(
        \ML_int[6][110] ) );
  MUX2_X2 M1_5_109 ( .A(\ML_int[5][109] ), .B(\ML_int[5][77] ), .S(n41), .Z(
        \ML_int[6][109] ) );
  MUX2_X2 M1_5_108 ( .A(\ML_int[5][108] ), .B(\ML_int[5][76] ), .S(n41), .Z(
        \ML_int[6][108] ) );
  MUX2_X2 M1_5_107 ( .A(\ML_int[5][107] ), .B(\ML_int[5][75] ), .S(n41), .Z(
        \ML_int[6][107] ) );
  MUX2_X2 M1_5_53 ( .A(\ML_int[5][53] ), .B(\ML_int[5][21] ), .S(n41), .Z(
        \ML_int[6][53] ) );
  MUX2_X2 M1_5_52 ( .A(\ML_int[5][52] ), .B(\ML_int[5][20] ), .S(n41), .Z(
        \ML_int[6][52] ) );
  MUX2_X2 M1_5_51 ( .A(\ML_int[5][51] ), .B(\ML_int[5][19] ), .S(n41), .Z(
        \ML_int[6][51] ) );
  MUX2_X2 M1_5_50 ( .A(\ML_int[5][50] ), .B(\ML_int[5][18] ), .S(n41), .Z(
        \ML_int[6][50] ) );
  MUX2_X2 M1_5_49 ( .A(\ML_int[5][49] ), .B(\ML_int[5][17] ), .S(n41), .Z(
        \ML_int[6][49] ) );
  MUX2_X2 M1_5_48 ( .A(\ML_int[5][48] ), .B(\ML_int[5][16] ), .S(n41), .Z(
        \ML_int[6][48] ) );
  MUX2_X2 M1_5_47 ( .A(\ML_int[5][47] ), .B(\ML_int[5][15] ), .S(n41), .Z(
        \ML_int[6][47] ) );
  MUX2_X2 M1_5_46 ( .A(\ML_int[5][46] ), .B(\ML_int[5][14] ), .S(n41), .Z(
        \ML_int[6][46] ) );
  MUX2_X2 M1_5_45 ( .A(\ML_int[5][45] ), .B(\ML_int[5][13] ), .S(n41), .Z(
        \ML_int[6][45] ) );
  MUX2_X2 M1_5_44 ( .A(\ML_int[5][44] ), .B(\ML_int[5][12] ), .S(n41), .Z(
        \ML_int[6][44] ) );
  MUX2_X2 M1_5_43 ( .A(\ML_int[5][43] ), .B(\ML_int[5][11] ), .S(n41), .Z(
        \ML_int[6][43] ) );
  MUX2_X2 M1_4_117 ( .A(\ML_int[4][117] ), .B(\ML_int[4][101] ), .S(n36), .Z(
        \ML_int[5][117] ) );
  MUX2_X2 M1_4_116 ( .A(\ML_int[4][116] ), .B(\ML_int[4][100] ), .S(n35), .Z(
        \ML_int[5][116] ) );
  MUX2_X2 M1_4_115 ( .A(\ML_int[4][115] ), .B(\ML_int[4][99] ), .S(n36), .Z(
        \ML_int[5][115] ) );
  MUX2_X2 M1_4_114 ( .A(\ML_int[4][114] ), .B(\ML_int[4][98] ), .S(n35), .Z(
        \ML_int[5][114] ) );
  MUX2_X2 M1_4_113 ( .A(\ML_int[4][113] ), .B(\ML_int[4][97] ), .S(n35), .Z(
        \ML_int[5][113] ) );
  MUX2_X2 M1_4_112 ( .A(\ML_int[4][112] ), .B(\ML_int[4][96] ), .S(n36), .Z(
        \ML_int[5][112] ) );
  MUX2_X2 M1_4_111 ( .A(\ML_int[4][111] ), .B(\ML_int[4][95] ), .S(n36), .Z(
        \ML_int[5][111] ) );
  MUX2_X2 M1_4_110 ( .A(\ML_int[4][110] ), .B(\ML_int[4][94] ), .S(n36), .Z(
        \ML_int[5][110] ) );
  MUX2_X2 M1_4_109 ( .A(\ML_int[4][109] ), .B(\ML_int[4][93] ), .S(n36), .Z(
        \ML_int[5][109] ) );
  MUX2_X2 M1_4_108 ( .A(\ML_int[4][108] ), .B(\ML_int[4][92] ), .S(n36), .Z(
        \ML_int[5][108] ) );
  MUX2_X2 M1_4_107 ( .A(\ML_int[4][107] ), .B(\ML_int[4][91] ), .S(n36), .Z(
        \ML_int[5][107] ) );
  MUX2_X2 M1_4_85 ( .A(\ML_int[4][85] ), .B(\ML_int[4][69] ), .S(n36), .Z(
        \ML_int[5][85] ) );
  MUX2_X2 M1_4_84 ( .A(\ML_int[4][84] ), .B(\ML_int[4][68] ), .S(n36), .Z(
        \ML_int[5][84] ) );
  MUX2_X2 M1_4_83 ( .A(\ML_int[4][83] ), .B(\ML_int[4][67] ), .S(n36), .Z(
        \ML_int[5][83] ) );
  MUX2_X2 M1_4_82 ( .A(\ML_int[4][82] ), .B(\ML_int[4][66] ), .S(n36), .Z(
        \ML_int[5][82] ) );
  MUX2_X2 M1_4_81 ( .A(\ML_int[4][81] ), .B(\ML_int[4][65] ), .S(n36), .Z(
        \ML_int[5][81] ) );
  MUX2_X2 M1_4_80 ( .A(\ML_int[4][80] ), .B(\ML_int[4][64] ), .S(n36), .Z(
        \ML_int[5][80] ) );
  MUX2_X2 M1_4_79 ( .A(\ML_int[4][79] ), .B(\ML_int[4][63] ), .S(n35), .Z(
        \ML_int[5][79] ) );
  MUX2_X2 M1_4_78 ( .A(\ML_int[4][78] ), .B(\ML_int[4][62] ), .S(n35), .Z(
        \ML_int[5][78] ) );
  MUX2_X2 M1_4_77 ( .A(\ML_int[4][77] ), .B(\ML_int[4][61] ), .S(n35), .Z(
        \ML_int[5][77] ) );
  MUX2_X2 M1_4_76 ( .A(\ML_int[4][76] ), .B(\ML_int[4][60] ), .S(n35), .Z(
        \ML_int[5][76] ) );
  MUX2_X2 M1_4_75 ( .A(\ML_int[4][75] ), .B(\ML_int[4][59] ), .S(n35), .Z(
        \ML_int[5][75] ) );
  MUX2_X2 M1_4_53 ( .A(\ML_int[4][53] ), .B(\ML_int[4][37] ), .S(n35), .Z(
        \ML_int[5][53] ) );
  MUX2_X2 M1_4_52 ( .A(\ML_int[4][52] ), .B(\ML_int[4][36] ), .S(n35), .Z(
        \ML_int[5][52] ) );
  MUX2_X2 M1_4_51 ( .A(\ML_int[4][51] ), .B(\ML_int[4][35] ), .S(n35), .Z(
        \ML_int[5][51] ) );
  MUX2_X2 M1_4_50 ( .A(\ML_int[4][50] ), .B(\ML_int[4][34] ), .S(n35), .Z(
        \ML_int[5][50] ) );
  MUX2_X2 M1_4_49 ( .A(\ML_int[4][49] ), .B(\ML_int[4][33] ), .S(n35), .Z(
        \ML_int[5][49] ) );
  MUX2_X2 M1_4_48 ( .A(\ML_int[4][48] ), .B(\ML_int[4][32] ), .S(n35), .Z(
        \ML_int[5][48] ) );
  MUX2_X2 M1_4_47 ( .A(\ML_int[4][47] ), .B(\ML_int[4][31] ), .S(
        \temp_int_SH[4] ), .Z(\ML_int[5][47] ) );
  MUX2_X2 M1_4_46 ( .A(\ML_int[4][46] ), .B(\ML_int[4][30] ), .S(
        \temp_int_SH[4] ), .Z(\ML_int[5][46] ) );
  MUX2_X2 M1_4_45 ( .A(\ML_int[4][45] ), .B(\ML_int[4][29] ), .S(
        \temp_int_SH[4] ), .Z(\ML_int[5][45] ) );
  MUX2_X2 M1_4_44 ( .A(\ML_int[4][44] ), .B(\ML_int[4][28] ), .S(
        \temp_int_SH[4] ), .Z(\ML_int[5][44] ) );
  MUX2_X2 M1_4_43 ( .A(\ML_int[4][43] ), .B(\ML_int[4][27] ), .S(
        \temp_int_SH[4] ), .Z(\ML_int[5][43] ) );
  MUX2_X2 M1_4_21 ( .A(\ML_int[4][21] ), .B(\ML_int[4][5] ), .S(
        \temp_int_SH[4] ), .Z(\ML_int[5][21] ) );
  MUX2_X2 M1_4_20 ( .A(\ML_int[4][20] ), .B(\ML_int[4][4] ), .S(
        \temp_int_SH[4] ), .Z(\ML_int[5][20] ) );
  MUX2_X2 M1_4_19 ( .A(\ML_int[4][19] ), .B(\ML_int[4][3] ), .S(n35), .Z(
        \ML_int[5][19] ) );
  MUX2_X2 M1_4_18 ( .A(\ML_int[4][18] ), .B(\ML_int[4][2] ), .S(n36), .Z(
        \ML_int[5][18] ) );
  MUX2_X2 M1_4_17 ( .A(\ML_int[4][17] ), .B(\ML_int[4][1] ), .S(n35), .Z(
        \ML_int[5][17] ) );
  MUX2_X2 M1_4_16 ( .A(\ML_int[4][16] ), .B(\ML_int[4][0] ), .S(n35), .Z(
        \ML_int[5][16] ) );
  MUX2_X2 M1_3_117 ( .A(n5), .B(\ML_int[3][109] ), .S(n30), .Z(
        \ML_int[4][117] ) );
  MUX2_X2 M1_3_116 ( .A(\ML_int[3][116] ), .B(\ML_int[3][108] ), .S(n30), .Z(
        \ML_int[4][116] ) );
  MUX2_X2 M1_3_115 ( .A(\ML_int[3][115] ), .B(\ML_int[3][107] ), .S(n30), .Z(
        \ML_int[4][115] ) );
  MUX2_X2 M1_3_114 ( .A(\ML_int[3][114] ), .B(\ML_int[3][106] ), .S(n30), .Z(
        \ML_int[4][114] ) );
  MUX2_X2 M1_3_113 ( .A(\ML_int[3][113] ), .B(\ML_int[3][105] ), .S(n30), .Z(
        \ML_int[4][113] ) );
  MUX2_X2 M1_3_112 ( .A(\ML_int[3][112] ), .B(\ML_int[3][104] ), .S(n30), .Z(
        \ML_int[4][112] ) );
  MUX2_X2 M1_3_111 ( .A(\ML_int[3][111] ), .B(\ML_int[3][103] ), .S(n30), .Z(
        \ML_int[4][111] ) );
  MUX2_X2 M1_3_110 ( .A(\ML_int[3][110] ), .B(\ML_int[3][102] ), .S(n30), .Z(
        \ML_int[4][110] ) );
  MUX2_X2 M1_3_109 ( .A(\ML_int[3][109] ), .B(\ML_int[3][101] ), .S(n30), .Z(
        \ML_int[4][109] ) );
  MUX2_X2 M1_3_108 ( .A(\ML_int[3][108] ), .B(\ML_int[3][100] ), .S(n30), .Z(
        \ML_int[4][108] ) );
  MUX2_X2 M1_3_107 ( .A(\ML_int[3][107] ), .B(\ML_int[3][99] ), .S(n30), .Z(
        \ML_int[4][107] ) );
  MUX2_X2 M1_3_101 ( .A(\ML_int[3][101] ), .B(\ML_int[3][93] ), .S(n32), .Z(
        \ML_int[4][101] ) );
  MUX2_X2 M1_3_100 ( .A(\ML_int[3][100] ), .B(\ML_int[3][92] ), .S(n32), .Z(
        \ML_int[4][100] ) );
  MUX2_X2 M1_3_99 ( .A(\ML_int[3][99] ), .B(\ML_int[3][91] ), .S(n32), .Z(
        \ML_int[4][99] ) );
  MUX2_X2 M1_3_98 ( .A(\ML_int[3][98] ), .B(\ML_int[3][90] ), .S(n32), .Z(
        \ML_int[4][98] ) );
  MUX2_X2 M1_3_97 ( .A(\ML_int[3][97] ), .B(\ML_int[3][89] ), .S(n32), .Z(
        \ML_int[4][97] ) );
  MUX2_X2 M1_3_96 ( .A(\ML_int[3][96] ), .B(\ML_int[3][88] ), .S(n32), .Z(
        \ML_int[4][96] ) );
  MUX2_X2 M1_3_95 ( .A(\ML_int[3][95] ), .B(\ML_int[3][87] ), .S(n32), .Z(
        \ML_int[4][95] ) );
  MUX2_X2 M1_3_94 ( .A(\ML_int[3][94] ), .B(\ML_int[3][86] ), .S(n32), .Z(
        \ML_int[4][94] ) );
  MUX2_X2 M1_3_93 ( .A(\ML_int[3][93] ), .B(\ML_int[3][85] ), .S(n32), .Z(
        \ML_int[4][93] ) );
  MUX2_X2 M1_3_92 ( .A(\ML_int[3][92] ), .B(\ML_int[3][84] ), .S(n32), .Z(
        \ML_int[4][92] ) );
  MUX2_X2 M1_3_91 ( .A(\ML_int[3][91] ), .B(\ML_int[3][83] ), .S(n32), .Z(
        \ML_int[4][91] ) );
  MUX2_X2 M1_3_85 ( .A(\ML_int[3][85] ), .B(\ML_int[3][77] ), .S(n30), .Z(
        \ML_int[4][85] ) );
  MUX2_X2 M1_3_84 ( .A(\ML_int[3][84] ), .B(\ML_int[3][76] ), .S(n32), .Z(
        \ML_int[4][84] ) );
  MUX2_X2 M1_3_83 ( .A(\ML_int[3][83] ), .B(\ML_int[3][75] ), .S(
        \temp_int_SH[3] ), .Z(\ML_int[4][83] ) );
  MUX2_X2 M1_3_82 ( .A(\ML_int[3][82] ), .B(\ML_int[3][74] ), .S(n32), .Z(
        \ML_int[4][82] ) );
  MUX2_X2 M1_3_81 ( .A(\ML_int[3][81] ), .B(\ML_int[3][73] ), .S(n30), .Z(
        \ML_int[4][81] ) );
  MUX2_X2 M1_3_80 ( .A(\ML_int[3][80] ), .B(\ML_int[3][72] ), .S(
        \temp_int_SH[3] ), .Z(\ML_int[4][80] ) );
  MUX2_X2 M1_3_79 ( .A(\ML_int[3][79] ), .B(\ML_int[3][71] ), .S(n31), .Z(
        \ML_int[4][79] ) );
  MUX2_X2 M1_3_78 ( .A(\ML_int[3][78] ), .B(\ML_int[3][70] ), .S(
        \temp_int_SH[3] ), .Z(\ML_int[4][78] ) );
  MUX2_X2 M1_3_77 ( .A(\ML_int[3][77] ), .B(\ML_int[3][69] ), .S(n30), .Z(
        \ML_int[4][77] ) );
  MUX2_X2 M1_3_76 ( .A(\ML_int[3][76] ), .B(\ML_int[3][68] ), .S(n32), .Z(
        \ML_int[4][76] ) );
  MUX2_X2 M1_3_75 ( .A(\ML_int[3][75] ), .B(\ML_int[3][67] ), .S(n30), .Z(
        \ML_int[4][75] ) );
  MUX2_X2 M1_3_69 ( .A(\ML_int[3][69] ), .B(\ML_int[3][61] ), .S(n31), .Z(
        \ML_int[4][69] ) );
  MUX2_X2 M1_3_68 ( .A(\ML_int[3][68] ), .B(\ML_int[3][60] ), .S(n31), .Z(
        \ML_int[4][68] ) );
  MUX2_X2 M1_3_67 ( .A(\ML_int[3][67] ), .B(\ML_int[3][59] ), .S(n31), .Z(
        \ML_int[4][67] ) );
  MUX2_X2 M1_3_66 ( .A(\ML_int[3][66] ), .B(\ML_int[3][58] ), .S(n31), .Z(
        \ML_int[4][66] ) );
  MUX2_X2 M1_3_65 ( .A(\ML_int[3][65] ), .B(\ML_int[3][57] ), .S(n31), .Z(
        \ML_int[4][65] ) );
  MUX2_X2 M1_3_64 ( .A(\ML_int[3][64] ), .B(\ML_int[3][56] ), .S(n31), .Z(
        \ML_int[4][64] ) );
  MUX2_X2 M1_3_63 ( .A(\ML_int[3][63] ), .B(\ML_int[3][55] ), .S(n31), .Z(
        \ML_int[4][63] ) );
  MUX2_X2 M1_3_62 ( .A(\ML_int[3][62] ), .B(\ML_int[3][54] ), .S(n31), .Z(
        \ML_int[4][62] ) );
  MUX2_X2 M1_3_61 ( .A(\ML_int[3][61] ), .B(\ML_int[3][53] ), .S(n31), .Z(
        \ML_int[4][61] ) );
  MUX2_X2 M1_3_60 ( .A(\ML_int[3][60] ), .B(\ML_int[3][52] ), .S(n31), .Z(
        \ML_int[4][60] ) );
  MUX2_X2 M1_3_59 ( .A(\ML_int[3][59] ), .B(\ML_int[3][51] ), .S(n31), .Z(
        \ML_int[4][59] ) );
  MUX2_X2 M1_3_53 ( .A(\ML_int[3][53] ), .B(\ML_int[3][45] ), .S(n31), .Z(
        \ML_int[4][53] ) );
  MUX2_X2 M1_3_52 ( .A(\ML_int[3][52] ), .B(\ML_int[3][44] ), .S(n32), .Z(
        \ML_int[4][52] ) );
  MUX2_X2 M1_3_51 ( .A(\ML_int[3][51] ), .B(\ML_int[3][43] ), .S(n31), .Z(
        \ML_int[4][51] ) );
  MUX2_X2 M1_3_50 ( .A(\ML_int[3][50] ), .B(\ML_int[3][42] ), .S(n32), .Z(
        \ML_int[4][50] ) );
  MUX2_X2 M1_3_49 ( .A(\ML_int[3][49] ), .B(\ML_int[3][41] ), .S(n30), .Z(
        \ML_int[4][49] ) );
  MUX2_X2 M1_3_48 ( .A(\ML_int[3][48] ), .B(\ML_int[3][40] ), .S(
        \temp_int_SH[3] ), .Z(\ML_int[4][48] ) );
  MUX2_X2 M1_3_47 ( .A(\ML_int[3][47] ), .B(\ML_int[3][39] ), .S(n30), .Z(
        \ML_int[4][47] ) );
  MUX2_X2 M1_3_46 ( .A(\ML_int[3][46] ), .B(\ML_int[3][38] ), .S(
        \temp_int_SH[3] ), .Z(\ML_int[4][46] ) );
  MUX2_X2 M1_3_45 ( .A(\ML_int[3][45] ), .B(\ML_int[3][37] ), .S(n31), .Z(
        \ML_int[4][45] ) );
  MUX2_X2 M1_3_44 ( .A(\ML_int[3][44] ), .B(\ML_int[3][36] ), .S(n32), .Z(
        \ML_int[4][44] ) );
  MUX2_X2 M1_3_43 ( .A(\ML_int[3][43] ), .B(\ML_int[3][35] ), .S(n31), .Z(
        \ML_int[4][43] ) );
  MUX2_X2 M1_3_37 ( .A(\ML_int[3][37] ), .B(\ML_int[3][29] ), .S(n32), .Z(
        \ML_int[4][37] ) );
  MUX2_X2 M1_3_36 ( .A(\ML_int[3][36] ), .B(\ML_int[3][28] ), .S(n32), .Z(
        \ML_int[4][36] ) );
  MUX2_X2 M1_3_35 ( .A(\ML_int[3][35] ), .B(\ML_int[3][27] ), .S(n30), .Z(
        \ML_int[4][35] ) );
  MUX2_X2 M1_3_34 ( .A(\ML_int[3][34] ), .B(\ML_int[3][26] ), .S(n32), .Z(
        \ML_int[4][34] ) );
  MUX2_X2 M1_3_33 ( .A(\ML_int[3][33] ), .B(\ML_int[3][25] ), .S(
        \temp_int_SH[3] ), .Z(\ML_int[4][33] ) );
  MUX2_X2 M1_3_32 ( .A(\ML_int[3][32] ), .B(\ML_int[3][24] ), .S(
        \temp_int_SH[3] ), .Z(\ML_int[4][32] ) );
  MUX2_X2 M1_3_31 ( .A(\ML_int[3][31] ), .B(\ML_int[3][23] ), .S(
        \temp_int_SH[3] ), .Z(\ML_int[4][31] ) );
  MUX2_X2 M1_3_30 ( .A(\ML_int[3][30] ), .B(\ML_int[3][22] ), .S(
        \temp_int_SH[3] ), .Z(\ML_int[4][30] ) );
  MUX2_X2 M1_3_29 ( .A(\ML_int[3][29] ), .B(\ML_int[3][21] ), .S(n32), .Z(
        \ML_int[4][29] ) );
  MUX2_X2 M1_3_28 ( .A(\ML_int[3][28] ), .B(\ML_int[3][20] ), .S(n32), .Z(
        \ML_int[4][28] ) );
  MUX2_X2 M1_3_27 ( .A(\ML_int[3][27] ), .B(\ML_int[3][19] ), .S(n32), .Z(
        \ML_int[4][27] ) );
  MUX2_X2 M1_3_21 ( .A(\ML_int[3][21] ), .B(\ML_int[3][13] ), .S(n32), .Z(
        \ML_int[4][21] ) );
  MUX2_X2 M1_3_20 ( .A(\ML_int[3][20] ), .B(\ML_int[3][12] ), .S(n32), .Z(
        \ML_int[4][20] ) );
  MUX2_X2 M1_3_19 ( .A(\ML_int[3][19] ), .B(\ML_int[3][11] ), .S(n30), .Z(
        \ML_int[4][19] ) );
  MUX2_X2 M1_3_18 ( .A(\ML_int[3][18] ), .B(\ML_int[3][10] ), .S(n32), .Z(
        \ML_int[4][18] ) );
  MUX2_X2 M1_3_17 ( .A(\ML_int[3][17] ), .B(\ML_int[3][9] ), .S(
        \temp_int_SH[3] ), .Z(\ML_int[4][17] ) );
  MUX2_X2 M1_3_16 ( .A(\ML_int[3][16] ), .B(\ML_int[3][8] ), .S(
        \temp_int_SH[3] ), .Z(\ML_int[4][16] ) );
  MUX2_X2 M1_3_15 ( .A(\ML_int[3][15] ), .B(\ML_int[3][7] ), .S(
        \temp_int_SH[3] ), .Z(\ML_int[4][15] ) );
  MUX2_X2 M1_3_14 ( .A(\ML_int[3][14] ), .B(\ML_int[3][6] ), .S(n32), .Z(
        \ML_int[4][14] ) );
  MUX2_X2 M1_3_13 ( .A(\ML_int[3][13] ), .B(\ML_int[3][5] ), .S(n32), .Z(
        \ML_int[4][13] ) );
  MUX2_X2 M1_3_12 ( .A(\ML_int[3][12] ), .B(\ML_int[3][4] ), .S(n32), .Z(
        \ML_int[4][12] ) );
  MUX2_X2 M1_3_11 ( .A(\ML_int[3][11] ), .B(n40), .S(n32), .Z(\ML_int[4][11] )
         );
  MUX2_X2 M1_2_116 ( .A(n4), .B(\ML_int[2][112] ), .S(n29), .Z(
        \ML_int[3][116] ) );
  MUX2_X2 M1_2_115 ( .A(n3), .B(\ML_int[2][111] ), .S(n29), .Z(
        \ML_int[3][115] ) );
  MUX2_X2 M1_2_114 ( .A(\ML_int[2][114] ), .B(\ML_int[2][110] ), .S(n29), .Z(
        \ML_int[3][114] ) );
  MUX2_X2 M1_2_113 ( .A(\ML_int[2][113] ), .B(\ML_int[2][109] ), .S(n29), .Z(
        \ML_int[3][113] ) );
  MUX2_X2 M1_2_112 ( .A(\ML_int[2][112] ), .B(\ML_int[2][108] ), .S(n29), .Z(
        \ML_int[3][112] ) );
  MUX2_X2 M1_2_111 ( .A(\ML_int[2][111] ), .B(\ML_int[2][107] ), .S(n29), .Z(
        \ML_int[3][111] ) );
  MUX2_X2 M1_2_110 ( .A(\ML_int[2][110] ), .B(\ML_int[2][106] ), .S(n29), .Z(
        \ML_int[3][110] ) );
  MUX2_X2 M1_2_109 ( .A(\ML_int[2][109] ), .B(\ML_int[2][105] ), .S(n29), .Z(
        \ML_int[3][109] ) );
  MUX2_X2 M1_2_108 ( .A(\ML_int[2][108] ), .B(\ML_int[2][104] ), .S(n29), .Z(
        \ML_int[3][108] ) );
  MUX2_X2 M1_2_107 ( .A(\ML_int[2][107] ), .B(\ML_int[2][103] ), .S(n29), .Z(
        \ML_int[3][107] ) );
  MUX2_X2 M1_2_106 ( .A(\ML_int[2][106] ), .B(\ML_int[2][102] ), .S(n29), .Z(
        \ML_int[3][106] ) );
  MUX2_X2 M1_2_105 ( .A(\ML_int[2][105] ), .B(\ML_int[2][101] ), .S(n29), .Z(
        \ML_int[3][105] ) );
  MUX2_X2 M1_2_104 ( .A(\ML_int[2][104] ), .B(\ML_int[2][100] ), .S(n29), .Z(
        \ML_int[3][104] ) );
  MUX2_X2 M1_2_103 ( .A(\ML_int[2][103] ), .B(\ML_int[2][99] ), .S(n29), .Z(
        \ML_int[3][103] ) );
  MUX2_X2 M1_2_102 ( .A(\ML_int[2][102] ), .B(\ML_int[2][98] ), .S(n28), .Z(
        \ML_int[3][102] ) );
  MUX2_X2 M1_2_101 ( .A(\ML_int[2][101] ), .B(\ML_int[2][97] ), .S(n28), .Z(
        \ML_int[3][101] ) );
  MUX2_X2 M1_2_100 ( .A(\ML_int[2][100] ), .B(\ML_int[2][96] ), .S(n28), .Z(
        \ML_int[3][100] ) );
  MUX2_X2 M1_2_99 ( .A(\ML_int[2][99] ), .B(\ML_int[2][95] ), .S(n28), .Z(
        \ML_int[3][99] ) );
  MUX2_X2 M1_2_98 ( .A(\ML_int[2][98] ), .B(\ML_int[2][94] ), .S(n28), .Z(
        \ML_int[3][98] ) );
  MUX2_X2 M1_2_97 ( .A(\ML_int[2][97] ), .B(\ML_int[2][93] ), .S(n28), .Z(
        \ML_int[3][97] ) );
  MUX2_X2 M1_2_96 ( .A(\ML_int[2][96] ), .B(\ML_int[2][92] ), .S(n28), .Z(
        \ML_int[3][96] ) );
  MUX2_X2 M1_2_95 ( .A(\ML_int[2][95] ), .B(\ML_int[2][91] ), .S(n28), .Z(
        \ML_int[3][95] ) );
  MUX2_X2 M1_2_94 ( .A(\ML_int[2][94] ), .B(\ML_int[2][90] ), .S(n28), .Z(
        \ML_int[3][94] ) );
  MUX2_X2 M1_2_93 ( .A(\ML_int[2][93] ), .B(\ML_int[2][89] ), .S(n28), .Z(
        \ML_int[3][93] ) );
  MUX2_X2 M1_2_92 ( .A(\ML_int[2][92] ), .B(\ML_int[2][88] ), .S(n28), .Z(
        \ML_int[3][92] ) );
  MUX2_X2 M1_2_91 ( .A(\ML_int[2][91] ), .B(\ML_int[2][87] ), .S(n27), .Z(
        \ML_int[3][91] ) );
  MUX2_X2 M1_2_90 ( .A(\ML_int[2][90] ), .B(\ML_int[2][86] ), .S(n27), .Z(
        \ML_int[3][90] ) );
  MUX2_X2 M1_2_89 ( .A(\ML_int[2][89] ), .B(\ML_int[2][85] ), .S(n27), .Z(
        \ML_int[3][89] ) );
  MUX2_X2 M1_2_88 ( .A(\ML_int[2][88] ), .B(\ML_int[2][84] ), .S(n27), .Z(
        \ML_int[3][88] ) );
  MUX2_X2 M1_2_87 ( .A(\ML_int[2][87] ), .B(\ML_int[2][83] ), .S(n27), .Z(
        \ML_int[3][87] ) );
  MUX2_X2 M1_2_86 ( .A(\ML_int[2][86] ), .B(\ML_int[2][82] ), .S(n27), .Z(
        \ML_int[3][86] ) );
  MUX2_X2 M1_2_85 ( .A(\ML_int[2][85] ), .B(\ML_int[2][81] ), .S(n27), .Z(
        \ML_int[3][85] ) );
  MUX2_X2 M1_2_84 ( .A(\ML_int[2][84] ), .B(\ML_int[2][80] ), .S(n27), .Z(
        \ML_int[3][84] ) );
  MUX2_X2 M1_2_83 ( .A(\ML_int[2][83] ), .B(\ML_int[2][79] ), .S(n27), .Z(
        \ML_int[3][83] ) );
  MUX2_X2 M1_2_82 ( .A(\ML_int[2][82] ), .B(\ML_int[2][78] ), .S(n27), .Z(
        \ML_int[3][82] ) );
  MUX2_X2 M1_2_81 ( .A(\ML_int[2][81] ), .B(\ML_int[2][77] ), .S(n27), .Z(
        \ML_int[3][81] ) );
  MUX2_X2 M1_2_80 ( .A(\ML_int[2][80] ), .B(\ML_int[2][76] ), .S(n27), .Z(
        \ML_int[3][80] ) );
  MUX2_X2 M1_2_79 ( .A(\ML_int[2][79] ), .B(\ML_int[2][75] ), .S(n27), .Z(
        \ML_int[3][79] ) );
  MUX2_X2 M1_2_78 ( .A(\ML_int[2][78] ), .B(\ML_int[2][74] ), .S(n27), .Z(
        \ML_int[3][78] ) );
  MUX2_X2 M1_2_77 ( .A(\ML_int[2][77] ), .B(\ML_int[2][73] ), .S(n27), .Z(
        \ML_int[3][77] ) );
  MUX2_X2 M1_2_76 ( .A(\ML_int[2][76] ), .B(\ML_int[2][72] ), .S(n27), .Z(
        \ML_int[3][76] ) );
  MUX2_X2 M1_2_75 ( .A(\ML_int[2][75] ), .B(\ML_int[2][71] ), .S(n27), .Z(
        \ML_int[3][75] ) );
  MUX2_X2 M1_2_74 ( .A(\ML_int[2][74] ), .B(\ML_int[2][70] ), .S(n27), .Z(
        \ML_int[3][74] ) );
  MUX2_X2 M1_2_73 ( .A(\ML_int[2][73] ), .B(\ML_int[2][69] ), .S(n27), .Z(
        \ML_int[3][73] ) );
  MUX2_X2 M1_2_72 ( .A(\ML_int[2][72] ), .B(\ML_int[2][68] ), .S(n27), .Z(
        \ML_int[3][72] ) );
  MUX2_X2 M1_2_71 ( .A(\ML_int[2][71] ), .B(\ML_int[2][67] ), .S(n27), .Z(
        \ML_int[3][71] ) );
  MUX2_X2 M1_2_70 ( .A(\ML_int[2][70] ), .B(\ML_int[2][66] ), .S(n27), .Z(
        \ML_int[3][70] ) );
  MUX2_X2 M1_2_69 ( .A(\ML_int[2][69] ), .B(\ML_int[2][65] ), .S(n24), .Z(
        \ML_int[3][69] ) );
  MUX2_X2 M1_2_68 ( .A(\ML_int[2][68] ), .B(\ML_int[2][64] ), .S(n23), .Z(
        \ML_int[3][68] ) );
  MUX2_X2 M1_2_67 ( .A(\ML_int[2][67] ), .B(\ML_int[2][63] ), .S(n28), .Z(
        \ML_int[3][67] ) );
  MUX2_X2 M1_2_66 ( .A(\ML_int[2][66] ), .B(\ML_int[2][62] ), .S(n25), .Z(
        \ML_int[3][66] ) );
  MUX2_X2 M1_2_65 ( .A(\ML_int[2][65] ), .B(\ML_int[2][61] ), .S(n25), .Z(
        \ML_int[3][65] ) );
  MUX2_X2 M1_2_64 ( .A(\ML_int[2][64] ), .B(\ML_int[2][60] ), .S(n28), .Z(
        \ML_int[3][64] ) );
  MUX2_X2 M1_2_63 ( .A(\ML_int[2][63] ), .B(\ML_int[2][59] ), .S(n26), .Z(
        \ML_int[3][63] ) );
  MUX2_X2 M1_2_62 ( .A(\ML_int[2][62] ), .B(\ML_int[2][58] ), .S(n25), .Z(
        \ML_int[3][62] ) );
  MUX2_X2 M1_2_61 ( .A(\ML_int[2][61] ), .B(\ML_int[2][57] ), .S(n28), .Z(
        \ML_int[3][61] ) );
  MUX2_X2 M1_2_60 ( .A(\ML_int[2][60] ), .B(\ML_int[2][56] ), .S(n26), .Z(
        \ML_int[3][60] ) );
  MUX2_X2 M1_2_59 ( .A(\ML_int[2][59] ), .B(\ML_int[2][55] ), .S(n28), .Z(
        \ML_int[3][59] ) );
  MUX2_X2 M1_2_58 ( .A(\ML_int[2][58] ), .B(\ML_int[2][54] ), .S(n26), .Z(
        \ML_int[3][58] ) );
  MUX2_X2 M1_2_57 ( .A(\ML_int[2][57] ), .B(\ML_int[2][53] ), .S(n26), .Z(
        \ML_int[3][57] ) );
  MUX2_X2 M1_2_56 ( .A(\ML_int[2][56] ), .B(\ML_int[2][52] ), .S(n26), .Z(
        \ML_int[3][56] ) );
  MUX2_X2 M1_2_55 ( .A(\ML_int[2][55] ), .B(\ML_int[2][51] ), .S(n26), .Z(
        \ML_int[3][55] ) );
  MUX2_X2 M1_2_54 ( .A(\ML_int[2][54] ), .B(\ML_int[2][50] ), .S(n26), .Z(
        \ML_int[3][54] ) );
  MUX2_X2 M1_2_53 ( .A(\ML_int[2][53] ), .B(\ML_int[2][49] ), .S(n26), .Z(
        \ML_int[3][53] ) );
  MUX2_X2 M1_2_52 ( .A(\ML_int[2][52] ), .B(\ML_int[2][48] ), .S(n26), .Z(
        \ML_int[3][52] ) );
  MUX2_X2 M1_2_51 ( .A(\ML_int[2][51] ), .B(\ML_int[2][47] ), .S(n26), .Z(
        \ML_int[3][51] ) );
  MUX2_X2 M1_2_50 ( .A(\ML_int[2][50] ), .B(\ML_int[2][46] ), .S(n26), .Z(
        \ML_int[3][50] ) );
  MUX2_X2 M1_2_49 ( .A(\ML_int[2][49] ), .B(\ML_int[2][45] ), .S(n26), .Z(
        \ML_int[3][49] ) );
  MUX2_X2 M1_2_48 ( .A(\ML_int[2][48] ), .B(\ML_int[2][44] ), .S(n26), .Z(
        \ML_int[3][48] ) );
  MUX2_X2 M1_2_47 ( .A(\ML_int[2][47] ), .B(\ML_int[2][43] ), .S(n25), .Z(
        \ML_int[3][47] ) );
  MUX2_X2 M1_2_46 ( .A(\ML_int[2][46] ), .B(\ML_int[2][42] ), .S(n25), .Z(
        \ML_int[3][46] ) );
  MUX2_X2 M1_2_45 ( .A(\ML_int[2][45] ), .B(\ML_int[2][41] ), .S(n25), .Z(
        \ML_int[3][45] ) );
  MUX2_X2 M1_2_44 ( .A(\ML_int[2][44] ), .B(\ML_int[2][40] ), .S(n25), .Z(
        \ML_int[3][44] ) );
  MUX2_X2 M1_2_43 ( .A(\ML_int[2][43] ), .B(\ML_int[2][39] ), .S(n25), .Z(
        \ML_int[3][43] ) );
  MUX2_X2 M1_2_42 ( .A(\ML_int[2][42] ), .B(\ML_int[2][38] ), .S(n25), .Z(
        \ML_int[3][42] ) );
  MUX2_X2 M1_2_41 ( .A(\ML_int[2][41] ), .B(\ML_int[2][37] ), .S(n25), .Z(
        \ML_int[3][41] ) );
  MUX2_X2 M1_2_40 ( .A(\ML_int[2][40] ), .B(\ML_int[2][36] ), .S(n25), .Z(
        \ML_int[3][40] ) );
  MUX2_X2 M1_2_39 ( .A(\ML_int[2][39] ), .B(\ML_int[2][35] ), .S(n25), .Z(
        \ML_int[3][39] ) );
  MUX2_X2 M1_2_38 ( .A(\ML_int[2][38] ), .B(\ML_int[2][34] ), .S(n25), .Z(
        \ML_int[3][38] ) );
  MUX2_X2 M1_2_37 ( .A(\ML_int[2][37] ), .B(\ML_int[2][33] ), .S(n25), .Z(
        \ML_int[3][37] ) );
  MUX2_X2 M1_2_36 ( .A(\ML_int[2][36] ), .B(\ML_int[2][32] ), .S(n29), .Z(
        \ML_int[3][36] ) );
  MUX2_X2 M1_2_35 ( .A(\ML_int[2][35] ), .B(\ML_int[2][31] ), .S(n28), .Z(
        \ML_int[3][35] ) );
  MUX2_X2 M1_2_34 ( .A(\ML_int[2][34] ), .B(\ML_int[2][30] ), .S(n25), .Z(
        \ML_int[3][34] ) );
  MUX2_X2 M1_2_33 ( .A(\ML_int[2][33] ), .B(\ML_int[2][29] ), .S(n29), .Z(
        \ML_int[3][33] ) );
  MUX2_X2 M1_2_32 ( .A(\ML_int[2][32] ), .B(\ML_int[2][28] ), .S(n29), .Z(
        \ML_int[3][32] ) );
  MUX2_X2 M1_2_31 ( .A(\ML_int[2][31] ), .B(\ML_int[2][27] ), .S(n29), .Z(
        \ML_int[3][31] ) );
  MUX2_X2 M1_2_30 ( .A(\ML_int[2][30] ), .B(\ML_int[2][26] ), .S(n29), .Z(
        \ML_int[3][30] ) );
  MUX2_X2 M1_2_29 ( .A(\ML_int[2][29] ), .B(\ML_int[2][25] ), .S(n29), .Z(
        \ML_int[3][29] ) );
  MUX2_X2 M1_2_28 ( .A(\ML_int[2][28] ), .B(\ML_int[2][24] ), .S(n29), .Z(
        \ML_int[3][28] ) );
  MUX2_X2 M1_2_27 ( .A(\ML_int[2][27] ), .B(\ML_int[2][23] ), .S(n24), .Z(
        \ML_int[3][27] ) );
  MUX2_X2 M1_2_26 ( .A(\ML_int[2][26] ), .B(\ML_int[2][22] ), .S(n23), .Z(
        \ML_int[3][26] ) );
  MUX2_X2 M1_2_25 ( .A(\ML_int[2][25] ), .B(\ML_int[2][21] ), .S(n24), .Z(
        \ML_int[3][25] ) );
  MUX2_X2 M1_2_24 ( .A(\ML_int[2][24] ), .B(\ML_int[2][20] ), .S(n24), .Z(
        \ML_int[3][24] ) );
  MUX2_X2 M1_2_23 ( .A(\ML_int[2][23] ), .B(\ML_int[2][19] ), .S(n24), .Z(
        \ML_int[3][23] ) );
  MUX2_X2 M1_2_22 ( .A(\ML_int[2][22] ), .B(\ML_int[2][18] ), .S(n24), .Z(
        \ML_int[3][22] ) );
  MUX2_X2 M1_2_21 ( .A(\ML_int[2][21] ), .B(\ML_int[2][17] ), .S(n24), .Z(
        \ML_int[3][21] ) );
  MUX2_X2 M1_2_20 ( .A(\ML_int[2][20] ), .B(\ML_int[2][16] ), .S(n24), .Z(
        \ML_int[3][20] ) );
  MUX2_X2 M1_2_19 ( .A(\ML_int[2][19] ), .B(\ML_int[2][15] ), .S(n24), .Z(
        \ML_int[3][19] ) );
  MUX2_X2 M1_2_18 ( .A(\ML_int[2][18] ), .B(\ML_int[2][14] ), .S(n24), .Z(
        \ML_int[3][18] ) );
  MUX2_X2 M1_2_17 ( .A(\ML_int[2][17] ), .B(\ML_int[2][13] ), .S(n24), .Z(
        \ML_int[3][17] ) );
  MUX2_X2 M1_2_16 ( .A(\ML_int[2][16] ), .B(\ML_int[2][12] ), .S(n24), .Z(
        \ML_int[3][16] ) );
  MUX2_X2 M1_2_15 ( .A(\ML_int[2][15] ), .B(\ML_int[2][11] ), .S(n24), .Z(
        \ML_int[3][15] ) );
  MUX2_X2 M1_2_14 ( .A(\ML_int[2][14] ), .B(\ML_int[2][10] ), .S(n23), .Z(
        \ML_int[3][14] ) );
  MUX2_X2 M1_2_13 ( .A(\ML_int[2][13] ), .B(\ML_int[2][9] ), .S(n23), .Z(
        \ML_int[3][13] ) );
  MUX2_X2 M1_2_12 ( .A(\ML_int[2][12] ), .B(\ML_int[2][8] ), .S(n23), .Z(
        \ML_int[3][12] ) );
  MUX2_X2 M1_2_11 ( .A(\ML_int[2][11] ), .B(\ML_int[2][7] ), .S(n23), .Z(
        \ML_int[3][11] ) );
  MUX2_X2 M1_2_10 ( .A(\ML_int[2][10] ), .B(\ML_int[2][6] ), .S(n23), .Z(
        \ML_int[3][10] ) );
  MUX2_X2 M1_2_9 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S(n23), .Z(
        \ML_int[3][9] ) );
  MUX2_X2 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(n23), .Z(
        \ML_int[3][8] ) );
  MUX2_X2 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(n23), .Z(
        \ML_int[3][7] ) );
  MUX2_X2 M1_2_6 ( .A(\ML_int[2][6] ), .B(\ML_int[2][2] ), .S(n23), .Z(
        \ML_int[3][6] ) );
  MUX2_X2 M1_2_5 ( .A(\ML_int[2][5] ), .B(n39), .S(n23), .Z(\ML_int[3][5] ) );
  MUX2_X2 M1_2_4 ( .A(\ML_int[2][4] ), .B(n37), .S(n23), .Z(\ML_int[3][4] ) );
  MUX2_X2 M1_1_114 ( .A(\MR_int[1][113] ), .B(\ML_int[1][112] ), .S(n22), .Z(
        \ML_int[2][114] ) );
  MUX2_X2 M1_1_113 ( .A(\ML_int[1][113] ), .B(\ML_int[1][111] ), .S(n21), .Z(
        \ML_int[2][113] ) );
  MUX2_X2 M1_1_112 ( .A(\ML_int[1][112] ), .B(\ML_int[1][110] ), .S(n19), .Z(
        \ML_int[2][112] ) );
  MUX2_X2 M1_1_111 ( .A(\ML_int[1][111] ), .B(\ML_int[1][109] ), .S(n22), .Z(
        \ML_int[2][111] ) );
  MUX2_X2 M1_1_110 ( .A(\ML_int[1][110] ), .B(\ML_int[1][108] ), .S(n22), .Z(
        \ML_int[2][110] ) );
  MUX2_X2 M1_1_109 ( .A(\ML_int[1][109] ), .B(\ML_int[1][107] ), .S(n22), .Z(
        \ML_int[2][109] ) );
  MUX2_X2 M1_1_108 ( .A(\ML_int[1][108] ), .B(\ML_int[1][106] ), .S(n22), .Z(
        \ML_int[2][108] ) );
  MUX2_X2 M1_1_107 ( .A(\ML_int[1][107] ), .B(\ML_int[1][105] ), .S(n22), .Z(
        \ML_int[2][107] ) );
  MUX2_X2 M1_1_106 ( .A(\ML_int[1][106] ), .B(\ML_int[1][104] ), .S(n22), .Z(
        \ML_int[2][106] ) );
  MUX2_X2 M1_1_105 ( .A(\ML_int[1][105] ), .B(\ML_int[1][103] ), .S(n22), .Z(
        \ML_int[2][105] ) );
  MUX2_X2 M1_1_104 ( .A(\ML_int[1][104] ), .B(\ML_int[1][102] ), .S(n22), .Z(
        \ML_int[2][104] ) );
  MUX2_X2 M1_1_103 ( .A(\ML_int[1][103] ), .B(\ML_int[1][101] ), .S(n22), .Z(
        \ML_int[2][103] ) );
  MUX2_X2 M1_1_102 ( .A(\ML_int[1][102] ), .B(\ML_int[1][100] ), .S(n22), .Z(
        \ML_int[2][102] ) );
  MUX2_X2 M1_1_101 ( .A(\ML_int[1][101] ), .B(\ML_int[1][99] ), .S(n22), .Z(
        \ML_int[2][101] ) );
  MUX2_X2 M1_1_100 ( .A(\ML_int[1][100] ), .B(\ML_int[1][98] ), .S(n21), .Z(
        \ML_int[2][100] ) );
  MUX2_X2 M1_1_99 ( .A(\ML_int[1][99] ), .B(\ML_int[1][97] ), .S(n21), .Z(
        \ML_int[2][99] ) );
  MUX2_X2 M1_1_98 ( .A(\ML_int[1][98] ), .B(\ML_int[1][96] ), .S(n21), .Z(
        \ML_int[2][98] ) );
  MUX2_X2 M1_1_97 ( .A(\ML_int[1][97] ), .B(\ML_int[1][95] ), .S(n21), .Z(
        \ML_int[2][97] ) );
  MUX2_X2 M1_1_96 ( .A(\ML_int[1][96] ), .B(\ML_int[1][94] ), .S(n21), .Z(
        \ML_int[2][96] ) );
  MUX2_X2 M1_1_95 ( .A(\ML_int[1][95] ), .B(\ML_int[1][93] ), .S(n21), .Z(
        \ML_int[2][95] ) );
  MUX2_X2 M1_1_94 ( .A(\ML_int[1][94] ), .B(\ML_int[1][92] ), .S(n21), .Z(
        \ML_int[2][94] ) );
  MUX2_X2 M1_1_93 ( .A(\ML_int[1][93] ), .B(\ML_int[1][91] ), .S(n21), .Z(
        \ML_int[2][93] ) );
  MUX2_X2 M1_1_92 ( .A(\ML_int[1][92] ), .B(\ML_int[1][90] ), .S(n21), .Z(
        \ML_int[2][92] ) );
  MUX2_X2 M1_1_91 ( .A(\ML_int[1][91] ), .B(\ML_int[1][89] ), .S(n21), .Z(
        \ML_int[2][91] ) );
  MUX2_X2 M1_1_90 ( .A(\ML_int[1][90] ), .B(\ML_int[1][88] ), .S(n21), .Z(
        \ML_int[2][90] ) );
  MUX2_X2 M1_1_89 ( .A(\ML_int[1][89] ), .B(\ML_int[1][87] ), .S(n20), .Z(
        \ML_int[2][89] ) );
  MUX2_X2 M1_1_88 ( .A(\ML_int[1][88] ), .B(\ML_int[1][86] ), .S(n20), .Z(
        \ML_int[2][88] ) );
  MUX2_X2 M1_1_87 ( .A(\ML_int[1][87] ), .B(\ML_int[1][85] ), .S(n20), .Z(
        \ML_int[2][87] ) );
  MUX2_X2 M1_1_86 ( .A(\ML_int[1][86] ), .B(\ML_int[1][84] ), .S(n20), .Z(
        \ML_int[2][86] ) );
  MUX2_X2 M1_1_85 ( .A(\ML_int[1][85] ), .B(\ML_int[1][83] ), .S(n20), .Z(
        \ML_int[2][85] ) );
  MUX2_X2 M1_1_84 ( .A(\ML_int[1][84] ), .B(\ML_int[1][82] ), .S(n20), .Z(
        \ML_int[2][84] ) );
  MUX2_X2 M1_1_83 ( .A(\ML_int[1][83] ), .B(\ML_int[1][81] ), .S(n20), .Z(
        \ML_int[2][83] ) );
  MUX2_X2 M1_1_82 ( .A(\ML_int[1][82] ), .B(\ML_int[1][80] ), .S(n20), .Z(
        \ML_int[2][82] ) );
  MUX2_X2 M1_1_81 ( .A(\ML_int[1][81] ), .B(\ML_int[1][79] ), .S(n20), .Z(
        \ML_int[2][81] ) );
  MUX2_X2 M1_1_80 ( .A(\ML_int[1][80] ), .B(\ML_int[1][78] ), .S(n20), .Z(
        \ML_int[2][80] ) );
  MUX2_X2 M1_1_79 ( .A(\ML_int[1][79] ), .B(\ML_int[1][77] ), .S(n20), .Z(
        \ML_int[2][79] ) );
  MUX2_X2 M1_1_78 ( .A(\ML_int[1][78] ), .B(\ML_int[1][76] ), .S(n19), .Z(
        \ML_int[2][78] ) );
  MUX2_X2 M1_1_77 ( .A(\ML_int[1][77] ), .B(\ML_int[1][75] ), .S(n19), .Z(
        \ML_int[2][77] ) );
  MUX2_X2 M1_1_76 ( .A(\ML_int[1][76] ), .B(\ML_int[1][74] ), .S(n19), .Z(
        \ML_int[2][76] ) );
  MUX2_X2 M1_1_75 ( .A(\ML_int[1][75] ), .B(\ML_int[1][73] ), .S(n19), .Z(
        \ML_int[2][75] ) );
  MUX2_X2 M1_1_74 ( .A(\ML_int[1][74] ), .B(\ML_int[1][72] ), .S(n19), .Z(
        \ML_int[2][74] ) );
  MUX2_X2 M1_1_73 ( .A(\ML_int[1][73] ), .B(\ML_int[1][71] ), .S(n19), .Z(
        \ML_int[2][73] ) );
  MUX2_X2 M1_1_72 ( .A(\ML_int[1][72] ), .B(\ML_int[1][70] ), .S(n19), .Z(
        \ML_int[2][72] ) );
  MUX2_X2 M1_1_71 ( .A(\ML_int[1][71] ), .B(\ML_int[1][69] ), .S(n19), .Z(
        \ML_int[2][71] ) );
  MUX2_X2 M1_1_70 ( .A(\ML_int[1][70] ), .B(\ML_int[1][68] ), .S(n19), .Z(
        \ML_int[2][70] ) );
  MUX2_X2 M1_1_69 ( .A(\ML_int[1][69] ), .B(\ML_int[1][67] ), .S(n19), .Z(
        \ML_int[2][69] ) );
  MUX2_X2 M1_1_68 ( .A(\ML_int[1][68] ), .B(\ML_int[1][66] ), .S(n19), .Z(
        \ML_int[2][68] ) );
  MUX2_X2 M1_1_67 ( .A(\ML_int[1][67] ), .B(\ML_int[1][65] ), .S(n18), .Z(
        \ML_int[2][67] ) );
  MUX2_X2 M1_1_66 ( .A(\ML_int[1][66] ), .B(\ML_int[1][64] ), .S(n18), .Z(
        \ML_int[2][66] ) );
  MUX2_X2 M1_1_65 ( .A(\ML_int[1][65] ), .B(\ML_int[1][63] ), .S(n18), .Z(
        \ML_int[2][65] ) );
  MUX2_X2 M1_1_64 ( .A(\ML_int[1][64] ), .B(\ML_int[1][62] ), .S(n18), .Z(
        \ML_int[2][64] ) );
  MUX2_X2 M1_1_63 ( .A(\ML_int[1][63] ), .B(\ML_int[1][61] ), .S(n18), .Z(
        \ML_int[2][63] ) );
  MUX2_X2 M1_1_62 ( .A(\ML_int[1][62] ), .B(\ML_int[1][60] ), .S(n18), .Z(
        \ML_int[2][62] ) );
  MUX2_X2 M1_1_61 ( .A(\ML_int[1][61] ), .B(\ML_int[1][59] ), .S(n18), .Z(
        \ML_int[2][61] ) );
  MUX2_X2 M1_1_60 ( .A(\ML_int[1][60] ), .B(\ML_int[1][58] ), .S(n18), .Z(
        \ML_int[2][60] ) );
  MUX2_X2 M1_1_59 ( .A(\ML_int[1][59] ), .B(\ML_int[1][57] ), .S(n18), .Z(
        \ML_int[2][59] ) );
  MUX2_X2 M1_1_58 ( .A(\ML_int[1][58] ), .B(\ML_int[1][56] ), .S(n18), .Z(
        \ML_int[2][58] ) );
  MUX2_X2 M1_1_57 ( .A(\ML_int[1][57] ), .B(\ML_int[1][55] ), .S(n18), .Z(
        \ML_int[2][57] ) );
  MUX2_X2 M1_1_56 ( .A(\ML_int[1][56] ), .B(\ML_int[1][54] ), .S(n20), .Z(
        \ML_int[2][56] ) );
  MUX2_X2 M1_1_55 ( .A(\ML_int[1][55] ), .B(\ML_int[1][53] ), .S(n19), .Z(
        \ML_int[2][55] ) );
  MUX2_X2 M1_1_54 ( .A(\ML_int[1][54] ), .B(\ML_int[1][52] ), .S(n16), .Z(
        \ML_int[2][54] ) );
  MUX2_X2 M1_1_53 ( .A(\ML_int[1][53] ), .B(\ML_int[1][51] ), .S(n20), .Z(
        \ML_int[2][53] ) );
  MUX2_X2 M1_1_52 ( .A(\ML_int[1][52] ), .B(\ML_int[1][50] ), .S(n20), .Z(
        \ML_int[2][52] ) );
  MUX2_X2 M1_1_51 ( .A(\ML_int[1][51] ), .B(\ML_int[1][49] ), .S(n20), .Z(
        \ML_int[2][51] ) );
  MUX2_X2 M1_1_50 ( .A(\ML_int[1][50] ), .B(\ML_int[1][48] ), .S(n20), .Z(
        \ML_int[2][50] ) );
  MUX2_X2 M1_1_49 ( .A(\ML_int[1][49] ), .B(\ML_int[1][47] ), .S(n20), .Z(
        \ML_int[2][49] ) );
  MUX2_X2 M1_1_48 ( .A(\ML_int[1][48] ), .B(\ML_int[1][46] ), .S(n20), .Z(
        \ML_int[2][48] ) );
  MUX2_X2 M1_1_47 ( .A(\ML_int[1][47] ), .B(\ML_int[1][45] ), .S(n20), .Z(
        \ML_int[2][47] ) );
  MUX2_X2 M1_1_46 ( .A(\ML_int[1][46] ), .B(\ML_int[1][44] ), .S(n20), .Z(
        \ML_int[2][46] ) );
  MUX2_X2 M1_1_45 ( .A(\ML_int[1][45] ), .B(\ML_int[1][43] ), .S(n17), .Z(
        \ML_int[2][45] ) );
  MUX2_X2 M1_1_44 ( .A(\ML_int[1][44] ), .B(\ML_int[1][42] ), .S(n17), .Z(
        \ML_int[2][44] ) );
  MUX2_X2 M1_1_43 ( .A(\ML_int[1][43] ), .B(\ML_int[1][41] ), .S(n17), .Z(
        \ML_int[2][43] ) );
  MUX2_X2 M1_1_42 ( .A(\ML_int[1][42] ), .B(\ML_int[1][40] ), .S(n17), .Z(
        \ML_int[2][42] ) );
  MUX2_X2 M1_1_41 ( .A(\ML_int[1][41] ), .B(\ML_int[1][39] ), .S(n17), .Z(
        \ML_int[2][41] ) );
  MUX2_X2 M1_1_40 ( .A(\ML_int[1][40] ), .B(\ML_int[1][38] ), .S(n17), .Z(
        \ML_int[2][40] ) );
  MUX2_X2 M1_1_39 ( .A(\ML_int[1][39] ), .B(\ML_int[1][37] ), .S(n17), .Z(
        \ML_int[2][39] ) );
  MUX2_X2 M1_1_38 ( .A(\ML_int[1][38] ), .B(\ML_int[1][36] ), .S(n17), .Z(
        \ML_int[2][38] ) );
  MUX2_X2 M1_1_37 ( .A(\ML_int[1][37] ), .B(\ML_int[1][35] ), .S(n17), .Z(
        \ML_int[2][37] ) );
  MUX2_X2 M1_1_36 ( .A(\ML_int[1][36] ), .B(\ML_int[1][34] ), .S(n17), .Z(
        \ML_int[2][36] ) );
  MUX2_X2 M1_1_35 ( .A(\ML_int[1][35] ), .B(\ML_int[1][33] ), .S(n17), .Z(
        \ML_int[2][35] ) );
  MUX2_X2 M1_1_34 ( .A(\ML_int[1][34] ), .B(\ML_int[1][32] ), .S(n16), .Z(
        \ML_int[2][34] ) );
  MUX2_X2 M1_1_33 ( .A(\ML_int[1][33] ), .B(\ML_int[1][31] ), .S(n16), .Z(
        \ML_int[2][33] ) );
  MUX2_X2 M1_1_32 ( .A(\ML_int[1][32] ), .B(\ML_int[1][30] ), .S(n16), .Z(
        \ML_int[2][32] ) );
  MUX2_X2 M1_1_31 ( .A(\ML_int[1][31] ), .B(\ML_int[1][29] ), .S(n16), .Z(
        \ML_int[2][31] ) );
  MUX2_X2 M1_1_30 ( .A(\ML_int[1][30] ), .B(\ML_int[1][28] ), .S(n16), .Z(
        \ML_int[2][30] ) );
  MUX2_X2 M1_1_29 ( .A(\ML_int[1][29] ), .B(\ML_int[1][27] ), .S(n16), .Z(
        \ML_int[2][29] ) );
  MUX2_X2 M1_1_28 ( .A(\ML_int[1][28] ), .B(\ML_int[1][26] ), .S(n16), .Z(
        \ML_int[2][28] ) );
  MUX2_X2 M1_1_27 ( .A(\ML_int[1][27] ), .B(\ML_int[1][25] ), .S(n16), .Z(
        \ML_int[2][27] ) );
  MUX2_X2 M1_1_26 ( .A(\ML_int[1][26] ), .B(\ML_int[1][24] ), .S(n16), .Z(
        \ML_int[2][26] ) );
  MUX2_X2 M1_1_25 ( .A(\ML_int[1][25] ), .B(\ML_int[1][23] ), .S(n16), .Z(
        \ML_int[2][25] ) );
  MUX2_X2 M1_1_24 ( .A(\ML_int[1][24] ), .B(\ML_int[1][22] ), .S(n16), .Z(
        \ML_int[2][24] ) );
  MUX2_X2 M1_1_23 ( .A(\ML_int[1][23] ), .B(\ML_int[1][21] ), .S(n15), .Z(
        \ML_int[2][23] ) );
  MUX2_X2 M1_1_22 ( .A(\ML_int[1][22] ), .B(\ML_int[1][20] ), .S(n15), .Z(
        \ML_int[2][22] ) );
  MUX2_X2 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S(n19), .Z(
        \ML_int[2][21] ) );
  MUX2_X2 M1_1_20 ( .A(\ML_int[1][20] ), .B(\ML_int[1][18] ), .S(n16), .Z(
        \ML_int[2][20] ) );
  MUX2_X2 M1_1_19 ( .A(\ML_int[1][19] ), .B(\ML_int[1][17] ), .S(n18), .Z(
        \ML_int[2][19] ) );
  MUX2_X2 M1_1_18 ( .A(\ML_int[1][18] ), .B(\ML_int[1][16] ), .S(n16), .Z(
        \ML_int[2][18] ) );
  MUX2_X2 M1_1_17 ( .A(\ML_int[1][17] ), .B(\ML_int[1][15] ), .S(n20), .Z(
        \ML_int[2][17] ) );
  MUX2_X2 M1_1_16 ( .A(\ML_int[1][16] ), .B(\ML_int[1][14] ), .S(n18), .Z(
        \ML_int[2][16] ) );
  MUX2_X2 M1_1_15 ( .A(\ML_int[1][15] ), .B(\ML_int[1][13] ), .S(n20), .Z(
        \ML_int[2][15] ) );
  MUX2_X2 M1_1_14 ( .A(\ML_int[1][14] ), .B(\ML_int[1][12] ), .S(n17), .Z(
        \ML_int[2][14] ) );
  MUX2_X2 M1_1_13 ( .A(\ML_int[1][13] ), .B(\ML_int[1][11] ), .S(n17), .Z(
        \ML_int[2][13] ) );
  MUX2_X2 M1_1_12 ( .A(\ML_int[1][12] ), .B(\ML_int[1][10] ), .S(n15), .Z(
        \ML_int[2][12] ) );
  MUX2_X2 M1_1_11 ( .A(\ML_int[1][11] ), .B(\ML_int[1][9] ), .S(n15), .Z(
        \ML_int[2][11] ) );
  MUX2_X2 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S(n15), .Z(
        \ML_int[2][10] ) );
  MUX2_X2 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S(n15), .Z(
        \ML_int[2][9] ) );
  MUX2_X2 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S(n15), .Z(
        \ML_int[2][8] ) );
  MUX2_X2 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S(n15), .Z(
        \ML_int[2][7] ) );
  MUX2_X2 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S(n15), .Z(
        \ML_int[2][6] ) );
  MUX2_X2 M1_1_5 ( .A(\ML_int[1][5] ), .B(\ML_int[1][3] ), .S(n15), .Z(
        \ML_int[2][5] ) );
  MUX2_X2 M1_1_4 ( .A(\ML_int[1][4] ), .B(\ML_int[1][2] ), .S(n15), .Z(
        \ML_int[2][4] ) );
  MUX2_X2 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(n15), .Z(
        \ML_int[2][3] ) );
  MUX2_X2 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S(n15), .Z(
        \ML_int[2][2] ) );
  MUX2_X2 M1_0_113 ( .A(A[113]), .B(A[112]), .S(n6), .Z(\ML_int[1][113] ) );
  MUX2_X2 M1_0_112 ( .A(A[112]), .B(A[111]), .S(n6), .Z(\ML_int[1][112] ) );
  MUX2_X2 M1_0_111 ( .A(A[111]), .B(A[110]), .S(n6), .Z(\ML_int[1][111] ) );
  MUX2_X2 M1_0_110 ( .A(A[110]), .B(A[109]), .S(n6), .Z(\ML_int[1][110] ) );
  MUX2_X2 M1_0_109 ( .A(A[109]), .B(A[108]), .S(n6), .Z(\ML_int[1][109] ) );
  MUX2_X2 M1_0_108 ( .A(A[108]), .B(A[107]), .S(n6), .Z(\ML_int[1][108] ) );
  MUX2_X2 M1_0_107 ( .A(A[107]), .B(A[106]), .S(n6), .Z(\ML_int[1][107] ) );
  MUX2_X2 M1_0_106 ( .A(A[106]), .B(A[105]), .S(n6), .Z(\ML_int[1][106] ) );
  MUX2_X2 M1_0_105 ( .A(A[105]), .B(A[104]), .S(n6), .Z(\ML_int[1][105] ) );
  MUX2_X2 M1_0_104 ( .A(A[104]), .B(A[103]), .S(n6), .Z(\ML_int[1][104] ) );
  MUX2_X2 M1_0_103 ( .A(A[103]), .B(A[102]), .S(n6), .Z(\ML_int[1][103] ) );
  MUX2_X2 M1_0_102 ( .A(A[102]), .B(A[101]), .S(n8), .Z(\ML_int[1][102] ) );
  MUX2_X2 M1_0_101 ( .A(A[101]), .B(A[100]), .S(n13), .Z(\ML_int[1][101] ) );
  MUX2_X2 M1_0_100 ( .A(A[100]), .B(A[99]), .S(n13), .Z(\ML_int[1][100] ) );
  MUX2_X2 M1_0_99 ( .A(A[99]), .B(A[98]), .S(n6), .Z(\ML_int[1][99] ) );
  MUX2_X2 M1_0_98 ( .A(A[98]), .B(A[97]), .S(n8), .Z(\ML_int[1][98] ) );
  MUX2_X2 M1_0_97 ( .A(A[97]), .B(A[96]), .S(n6), .Z(\ML_int[1][97] ) );
  MUX2_X2 M1_0_96 ( .A(A[96]), .B(A[95]), .S(n8), .Z(\ML_int[1][96] ) );
  MUX2_X2 M1_0_95 ( .A(A[95]), .B(A[94]), .S(n8), .Z(\ML_int[1][95] ) );
  MUX2_X2 M1_0_94 ( .A(A[94]), .B(A[93]), .S(n6), .Z(\ML_int[1][94] ) );
  MUX2_X2 M1_0_93 ( .A(A[93]), .B(A[92]), .S(n13), .Z(\ML_int[1][93] ) );
  MUX2_X2 M1_0_92 ( .A(A[92]), .B(A[91]), .S(n13), .Z(\ML_int[1][92] ) );
  MUX2_X2 M1_0_91 ( .A(A[91]), .B(A[90]), .S(n12), .Z(\ML_int[1][91] ) );
  MUX2_X2 M1_0_90 ( .A(A[90]), .B(A[89]), .S(n12), .Z(\ML_int[1][90] ) );
  MUX2_X2 M1_0_89 ( .A(A[89]), .B(A[88]), .S(n9), .Z(\ML_int[1][89] ) );
  MUX2_X2 M1_0_88 ( .A(A[88]), .B(A[87]), .S(n13), .Z(\ML_int[1][88] ) );
  MUX2_X2 M1_0_87 ( .A(A[87]), .B(A[86]), .S(n13), .Z(\ML_int[1][87] ) );
  MUX2_X2 M1_0_86 ( .A(A[86]), .B(A[85]), .S(n13), .Z(\ML_int[1][86] ) );
  MUX2_X2 M1_0_85 ( .A(A[85]), .B(A[84]), .S(n12), .Z(\ML_int[1][85] ) );
  MUX2_X2 M1_0_84 ( .A(A[84]), .B(A[83]), .S(n12), .Z(\ML_int[1][84] ) );
  MUX2_X2 M1_0_83 ( .A(A[83]), .B(A[82]), .S(n9), .Z(\ML_int[1][83] ) );
  MUX2_X2 M1_0_82 ( .A(A[82]), .B(A[81]), .S(n9), .Z(\ML_int[1][82] ) );
  MUX2_X2 M1_0_81 ( .A(A[81]), .B(A[80]), .S(n13), .Z(\ML_int[1][81] ) );
  MUX2_X2 M1_0_80 ( .A(A[80]), .B(A[79]), .S(n8), .Z(\ML_int[1][80] ) );
  MUX2_X2 M1_0_79 ( .A(A[79]), .B(A[78]), .S(n8), .Z(\ML_int[1][79] ) );
  MUX2_X2 M1_0_78 ( .A(A[78]), .B(A[77]), .S(n13), .Z(\ML_int[1][78] ) );
  MUX2_X2 M1_0_77 ( .A(A[77]), .B(A[76]), .S(n8), .Z(\ML_int[1][77] ) );
  MUX2_X2 M1_0_76 ( .A(A[76]), .B(A[75]), .S(n13), .Z(\ML_int[1][76] ) );
  MUX2_X2 M1_0_75 ( .A(A[75]), .B(A[74]), .S(n8), .Z(\ML_int[1][75] ) );
  MUX2_X2 M1_0_74 ( .A(A[74]), .B(A[73]), .S(n8), .Z(\ML_int[1][74] ) );
  MUX2_X2 M1_0_73 ( .A(A[73]), .B(A[72]), .S(n8), .Z(\ML_int[1][73] ) );
  MUX2_X2 M1_0_72 ( .A(A[72]), .B(A[71]), .S(n8), .Z(\ML_int[1][72] ) );
  MUX2_X2 M1_0_71 ( .A(A[71]), .B(A[70]), .S(n8), .Z(\ML_int[1][71] ) );
  MUX2_X2 M1_0_70 ( .A(A[70]), .B(A[69]), .S(n8), .Z(\ML_int[1][70] ) );
  MUX2_X2 M1_0_69 ( .A(A[69]), .B(A[68]), .S(n12), .Z(\ML_int[1][69] ) );
  MUX2_X2 M1_0_68 ( .A(A[68]), .B(A[67]), .S(n12), .Z(\ML_int[1][68] ) );
  MUX2_X2 M1_0_67 ( .A(A[67]), .B(A[66]), .S(n13), .Z(\ML_int[1][67] ) );
  MUX2_X2 M1_0_66 ( .A(A[66]), .B(A[65]), .S(n8), .Z(\ML_int[1][66] ) );
  MUX2_X2 M1_0_65 ( .A(A[65]), .B(A[64]), .S(n13), .Z(\ML_int[1][65] ) );
  MUX2_X2 M1_0_64 ( .A(A[64]), .B(A[63]), .S(n9), .Z(\ML_int[1][64] ) );
  MUX2_X2 M1_0_63 ( .A(A[63]), .B(A[62]), .S(n12), .Z(\ML_int[1][63] ) );
  MUX2_X2 M1_0_62 ( .A(A[62]), .B(A[61]), .S(n12), .Z(\ML_int[1][62] ) );
  MUX2_X2 M1_0_61 ( .A(A[61]), .B(A[60]), .S(n13), .Z(\ML_int[1][61] ) );
  MUX2_X2 M1_0_60 ( .A(A[60]), .B(A[59]), .S(n12), .Z(\ML_int[1][60] ) );
  MUX2_X2 M1_0_59 ( .A(A[59]), .B(A[58]), .S(n9), .Z(\ML_int[1][59] ) );
  MUX2_X2 M1_0_58 ( .A(A[58]), .B(A[57]), .S(n7), .Z(\ML_int[1][58] ) );
  MUX2_X2 M1_0_57 ( .A(A[57]), .B(A[56]), .S(n7), .Z(\ML_int[1][57] ) );
  MUX2_X2 M1_0_56 ( .A(A[56]), .B(A[55]), .S(n7), .Z(\ML_int[1][56] ) );
  MUX2_X2 M1_0_55 ( .A(A[55]), .B(A[54]), .S(n7), .Z(\ML_int[1][55] ) );
  MUX2_X2 M1_0_54 ( .A(A[54]), .B(A[53]), .S(n7), .Z(\ML_int[1][54] ) );
  MUX2_X2 M1_0_53 ( .A(A[53]), .B(A[52]), .S(n7), .Z(\ML_int[1][53] ) );
  MUX2_X2 M1_0_52 ( .A(A[52]), .B(A[51]), .S(n7), .Z(\ML_int[1][52] ) );
  MUX2_X2 M1_0_51 ( .A(A[51]), .B(A[50]), .S(n7), .Z(\ML_int[1][51] ) );
  MUX2_X2 M1_0_50 ( .A(A[50]), .B(A[49]), .S(n7), .Z(\ML_int[1][50] ) );
  MUX2_X2 M1_0_49 ( .A(A[49]), .B(A[48]), .S(n7), .Z(\ML_int[1][49] ) );
  MUX2_X2 M1_0_48 ( .A(A[48]), .B(A[47]), .S(n7), .Z(\ML_int[1][48] ) );
  MUX2_X2 M1_0_47 ( .A(A[47]), .B(A[46]), .S(n13), .Z(\ML_int[1][47] ) );
  MUX2_X2 M1_0_46 ( .A(A[46]), .B(A[45]), .S(n6), .Z(\ML_int[1][46] ) );
  MUX2_X2 M1_0_45 ( .A(A[45]), .B(A[44]), .S(n13), .Z(\ML_int[1][45] ) );
  MUX2_X2 M1_0_44 ( .A(A[44]), .B(A[43]), .S(n13), .Z(\ML_int[1][44] ) );
  MUX2_X2 M1_0_43 ( .A(A[43]), .B(A[42]), .S(n6), .Z(\ML_int[1][43] ) );
  MUX2_X2 M1_0_42 ( .A(A[42]), .B(A[41]), .S(n6), .Z(\ML_int[1][42] ) );
  MUX2_X2 M1_0_41 ( .A(A[41]), .B(A[40]), .S(n13), .Z(\ML_int[1][41] ) );
  MUX2_X2 M1_0_40 ( .A(A[40]), .B(A[39]), .S(n13), .Z(\ML_int[1][40] ) );
  MUX2_X2 M1_0_39 ( .A(A[39]), .B(A[38]), .S(n13), .Z(\ML_int[1][39] ) );
  MUX2_X2 M1_0_38 ( .A(A[38]), .B(A[37]), .S(n13), .Z(\ML_int[1][38] ) );
  MUX2_X2 M1_0_37 ( .A(A[37]), .B(A[36]), .S(n13), .Z(\ML_int[1][37] ) );
  MUX2_X2 M1_0_36 ( .A(A[36]), .B(A[35]), .S(n8), .Z(\ML_int[1][36] ) );
  MUX2_X2 M1_0_35 ( .A(A[35]), .B(A[34]), .S(n8), .Z(\ML_int[1][35] ) );
  MUX2_X2 M1_0_34 ( .A(A[34]), .B(A[33]), .S(n8), .Z(\ML_int[1][34] ) );
  MUX2_X2 M1_0_33 ( .A(A[33]), .B(A[32]), .S(n8), .Z(\ML_int[1][33] ) );
  MUX2_X2 M1_0_32 ( .A(A[32]), .B(A[31]), .S(n8), .Z(\ML_int[1][32] ) );
  MUX2_X2 M1_0_31 ( .A(A[31]), .B(A[30]), .S(n8), .Z(\ML_int[1][31] ) );
  MUX2_X2 M1_0_30 ( .A(A[30]), .B(A[29]), .S(n8), .Z(\ML_int[1][30] ) );
  MUX2_X2 M1_0_29 ( .A(A[29]), .B(A[28]), .S(n8), .Z(\ML_int[1][29] ) );
  MUX2_X2 M1_0_28 ( .A(A[28]), .B(A[27]), .S(n8), .Z(\ML_int[1][28] ) );
  MUX2_X2 M1_0_27 ( .A(A[27]), .B(A[26]), .S(n8), .Z(\ML_int[1][27] ) );
  MUX2_X2 M1_0_26 ( .A(A[26]), .B(A[25]), .S(n8), .Z(\ML_int[1][26] ) );
  MUX2_X2 M1_0_25 ( .A(A[25]), .B(A[24]), .S(n7), .Z(\ML_int[1][25] ) );
  MUX2_X2 M1_0_24 ( .A(A[24]), .B(A[23]), .S(n13), .Z(\ML_int[1][24] ) );
  MUX2_X2 M1_0_23 ( .A(A[23]), .B(A[22]), .S(n7), .Z(\ML_int[1][23] ) );
  MUX2_X2 M1_0_22 ( .A(A[22]), .B(A[21]), .S(n7), .Z(\ML_int[1][22] ) );
  MUX2_X2 M1_0_21 ( .A(A[21]), .B(A[20]), .S(n7), .Z(\ML_int[1][21] ) );
  MUX2_X2 M1_0_20 ( .A(A[20]), .B(A[19]), .S(n7), .Z(\ML_int[1][20] ) );
  MUX2_X2 M1_0_19 ( .A(A[19]), .B(A[18]), .S(n7), .Z(\ML_int[1][19] ) );
  MUX2_X2 M1_0_18 ( .A(A[18]), .B(A[17]), .S(n7), .Z(\ML_int[1][18] ) );
  MUX2_X2 M1_0_17 ( .A(A[17]), .B(A[16]), .S(n7), .Z(\ML_int[1][17] ) );
  MUX2_X2 M1_0_16 ( .A(A[16]), .B(A[15]), .S(n13), .Z(\ML_int[1][16] ) );
  MUX2_X2 M1_0_15 ( .A(A[15]), .B(A[14]), .S(n6), .Z(\ML_int[1][15] ) );
  MUX2_X2 M1_0_14 ( .A(A[14]), .B(A[13]), .S(n9), .Z(\ML_int[1][14] ) );
  MUX2_X2 M1_0_13 ( .A(A[13]), .B(A[12]), .S(n9), .Z(\ML_int[1][13] ) );
  MUX2_X2 M1_0_12 ( .A(A[12]), .B(A[11]), .S(n9), .Z(\ML_int[1][12] ) );
  MUX2_X2 M1_0_11 ( .A(A[11]), .B(A[10]), .S(n9), .Z(\ML_int[1][11] ) );
  MUX2_X2 M1_0_10 ( .A(A[10]), .B(A[9]), .S(n9), .Z(\ML_int[1][10] ) );
  MUX2_X2 M1_0_9 ( .A(A[9]), .B(A[8]), .S(n9), .Z(\ML_int[1][9] ) );
  MUX2_X2 M1_0_8 ( .A(A[8]), .B(A[7]), .S(n9), .Z(\ML_int[1][8] ) );
  MUX2_X2 M1_0_7 ( .A(A[7]), .B(A[6]), .S(n9), .Z(\ML_int[1][7] ) );
  MUX2_X2 M1_0_6 ( .A(A[6]), .B(A[5]), .S(n9), .Z(\ML_int[1][6] ) );
  MUX2_X2 M1_0_5 ( .A(A[5]), .B(A[4]), .S(n9), .Z(\ML_int[1][5] ) );
  MUX2_X2 M1_0_4 ( .A(A[4]), .B(A[3]), .S(n9), .Z(\ML_int[1][4] ) );
  MUX2_X2 M1_0_3 ( .A(A[3]), .B(A[2]), .S(n13), .Z(\ML_int[1][3] ) );
  MUX2_X2 M1_0_2 ( .A(A[2]), .B(A[1]), .S(n13), .Z(\ML_int[1][2] ) );
  MUX2_X2 M1_0_1 ( .A(A[1]), .B(A[0]), .S(n13), .Z(\ML_int[1][1] ) );
  AND2_X4 U3 ( .A1(n46), .A2(n54), .ZN(n1) );
  AND2_X4 U4 ( .A1(n46), .A2(n53), .ZN(n2) );
  INV_X4 U5 ( .A(\temp_int_SH[0] ), .ZN(n14) );
  INV_X4 U6 ( .A(n2), .ZN(n27) );
  INV_X4 U7 ( .A(n10), .ZN(n7) );
  INV_X4 U8 ( .A(\temp_int_SH[0] ), .ZN(n10) );
  INV_X4 U9 ( .A(n10), .ZN(n9) );
  INV_X4 U10 ( .A(n14), .ZN(n12) );
  INV_X4 U11 ( .A(n14), .ZN(n8) );
  INV_X4 U12 ( .A(n2), .ZN(n26) );
  INV_X4 U13 ( .A(n11), .ZN(n6) );
  INV_X4 U14 ( .A(n1), .ZN(n16) );
  INV_X4 U15 ( .A(n1), .ZN(n19) );
  INV_X4 U16 ( .A(n1), .ZN(n20) );
  AND2_X4 U17 ( .A1(n19), .A2(\ML_int[1][113] ), .ZN(n3) );
  INV_X4 U18 ( .A(\temp_int_SH[3] ), .ZN(n33) );
  INV_X4 U19 ( .A(n33), .ZN(n31) );
  INV_X4 U20 ( .A(n33), .ZN(n30) );
  INV_X4 U21 ( .A(n1), .ZN(n15) );
  INV_X4 U22 ( .A(n1), .ZN(n18) );
  INV_X4 U23 ( .A(n1), .ZN(n17) );
  INV_X4 U24 ( .A(\temp_int_SH[4] ), .ZN(n34) );
  INV_X4 U25 ( .A(n12), .ZN(n11) );
  INV_X4 U26 ( .A(n2), .ZN(n25) );
  INV_X4 U27 ( .A(n2), .ZN(n29) );
  INV_X4 U28 ( .A(n2), .ZN(n23) );
  INV_X4 U29 ( .A(n2), .ZN(n24) );
  INV_X4 U30 ( .A(n2), .ZN(n28) );
  INV_X4 U31 ( .A(n33), .ZN(n32) );
  INV_X4 U32 ( .A(n34), .ZN(n35) );
  INV_X4 U33 ( .A(n34), .ZN(n36) );
  INV_X4 U34 ( .A(n1), .ZN(n22) );
  INV_X4 U35 ( .A(n1), .ZN(n21) );
  INV_X4 U36 ( .A(n14), .ZN(n13) );
  AND2_X4 U37 ( .A1(n15), .A2(\MR_int[1][113] ), .ZN(n4) );
  AND2_X4 U38 ( .A1(n29), .A2(\ML_int[2][113] ), .ZN(n5) );
  INV_X4 U39 ( .A(n51), .ZN(n37) );
  INV_X4 U40 ( .A(\ML_int[2][2] ), .ZN(n38) );
  INV_X4 U41 ( .A(n50), .ZN(n39) );
  INV_X4 U42 ( .A(n48), .ZN(n40) );
  INV_X4 U43 ( .A(SHMAG[5]), .ZN(n41) );
  INV_X4 U44 ( .A(SHMAG[6]), .ZN(n42) );
  INV_X4 U45 ( .A(n46), .ZN(n43) );
  INV_X4 U46 ( .A(SH[10]), .ZN(n44) );
  OAI21_X1 U47 ( .B1(SH[6]), .B2(n43), .A(n45), .ZN(SHMAG[6]) );
  OAI21_X1 U48 ( .B1(SH[5]), .B2(n43), .A(n45), .ZN(SHMAG[5]) );
  AND2_X1 U49 ( .A1(\ML_int[7][117] ), .A2(n44), .ZN(\ML_int[8][117] ) );
  AND2_X1 U50 ( .A1(\ML_int[7][116] ), .A2(n44), .ZN(\ML_int[8][116] ) );
  AND2_X1 U51 ( .A1(\ML_int[7][115] ), .A2(n44), .ZN(\ML_int[8][115] ) );
  AND2_X1 U52 ( .A1(\ML_int[7][114] ), .A2(n44), .ZN(\ML_int[8][114] ) );
  AND2_X1 U53 ( .A1(\ML_int[7][113] ), .A2(n44), .ZN(\ML_int[8][113] ) );
  AND2_X1 U54 ( .A1(\ML_int[7][112] ), .A2(n44), .ZN(\ML_int[8][112] ) );
  AND2_X1 U55 ( .A1(\ML_int[7][111] ), .A2(n44), .ZN(\ML_int[8][111] ) );
  AND2_X1 U56 ( .A1(\ML_int[7][110] ), .A2(n44), .ZN(\ML_int[8][110] ) );
  AND2_X1 U57 ( .A1(\ML_int[7][109] ), .A2(n44), .ZN(\ML_int[8][109] ) );
  AND2_X1 U58 ( .A1(\ML_int[7][108] ), .A2(n44), .ZN(\ML_int[8][108] ) );
  AND2_X1 U59 ( .A1(\ML_int[7][107] ), .A2(n44), .ZN(\ML_int[8][107] ) );
  AND2_X1 U60 ( .A1(\ML_int[4][15] ), .A2(n34), .ZN(\ML_int[5][15] ) );
  AND2_X1 U61 ( .A1(\ML_int[4][14] ), .A2(n34), .ZN(\ML_int[5][14] ) );
  AND2_X1 U62 ( .A1(\ML_int[4][13] ), .A2(n34), .ZN(\ML_int[5][13] ) );
  AND2_X1 U63 ( .A1(\ML_int[4][12] ), .A2(n34), .ZN(\ML_int[5][12] ) );
  AND2_X1 U64 ( .A1(\ML_int[4][11] ), .A2(n34), .ZN(\ML_int[5][11] ) );
  NAND2_X1 U65 ( .A1(n46), .A2(n47), .ZN(\temp_int_SH[4] ) );
  NAND2_X1 U66 ( .A1(SH[4]), .A2(n45), .ZN(n47) );
  AND2_X1 U67 ( .A1(\ML_int[3][5] ), .A2(n33), .ZN(\ML_int[4][5] ) );
  AND2_X1 U68 ( .A1(\ML_int[3][4] ), .A2(n33), .ZN(\ML_int[4][4] ) );
  NOR2_X1 U69 ( .A1(n30), .A2(n48), .ZN(\ML_int[4][3] ) );
  NOR2_X1 U70 ( .A1(n38), .A2(n49), .ZN(\ML_int[4][2] ) );
  NOR2_X1 U71 ( .A1(n49), .A2(n50), .ZN(\ML_int[4][1] ) );
  NOR2_X1 U72 ( .A1(n49), .A2(n51), .ZN(\ML_int[4][0] ) );
  NAND2_X1 U73 ( .A1(n2), .A2(n33), .ZN(n49) );
  NAND2_X1 U74 ( .A1(n46), .A2(n52), .ZN(\temp_int_SH[3] ) );
  NAND2_X1 U75 ( .A1(SH[3]), .A2(n45), .ZN(n52) );
  NAND2_X1 U76 ( .A1(\ML_int[2][3] ), .A2(n2), .ZN(n48) );
  NAND2_X1 U77 ( .A1(SH[2]), .A2(n45), .ZN(n53) );
  NAND2_X1 U78 ( .A1(\ML_int[1][1] ), .A2(n1), .ZN(n50) );
  NAND2_X1 U79 ( .A1(\ML_int[1][0] ), .A2(n1), .ZN(n51) );
  NAND2_X1 U80 ( .A1(SH[1]), .A2(n45), .ZN(n54) );
  AND2_X1 U81 ( .A1(A[113]), .A2(n6), .ZN(\MR_int[1][113] ) );
  AND2_X1 U82 ( .A1(A[0]), .A2(n11), .ZN(\ML_int[1][0] ) );
  NAND2_X1 U83 ( .A1(n46), .A2(n55), .ZN(\temp_int_SH[0] ) );
  NAND2_X1 U84 ( .A1(SH[0]), .A2(n45), .ZN(n55) );
  NAND2_X1 U85 ( .A1(SH[10]), .A2(n56), .ZN(n45) );
  NAND3_X1 U86 ( .A1(SH[8]), .A2(SH[7]), .A3(SH[9]), .ZN(n56) );
  NAND2_X1 U87 ( .A1(n57), .A2(n44), .ZN(n46) );
  OR3_X1 U88 ( .A1(SH[8]), .A2(SH[9]), .A3(SH[7]), .ZN(n57) );
endmodule


module fpu_DW01_sub_4 ( A, B, CI, DIFF, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
;
  wire   [11:1] carry;

  FA_X1 U2_6 ( .A(A[6]), .B(n14), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA_X1 U2_5 ( .A(A[5]), .B(n13), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n12), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_3 ( .A(A[3]), .B(n11), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA_X1 U2_2 ( .A(A[2]), .B(n10), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA_X1 U2_1 ( .A(A[1]), .B(n15), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  NAND2_X2 U1 ( .A1(n1), .A2(n2), .ZN(carry[11]) );
  XNOR2_X2 U2 ( .A(A[10]), .B(carry[10]), .ZN(DIFF[10]) );
  INV_X4 U3 ( .A(A[10]), .ZN(n1) );
  INV_X4 U4 ( .A(carry[10]), .ZN(n2) );
  XNOR2_X2 U5 ( .A(A[11]), .B(carry[11]), .ZN(DIFF[11]) );
  NAND2_X2 U6 ( .A1(n3), .A2(n4), .ZN(carry[8]) );
  XNOR2_X2 U7 ( .A(A[7]), .B(carry[7]), .ZN(DIFF[7]) );
  INV_X4 U8 ( .A(A[7]), .ZN(n3) );
  INV_X4 U9 ( .A(carry[7]), .ZN(n4) );
  NAND2_X2 U10 ( .A1(n5), .A2(n6), .ZN(carry[9]) );
  XNOR2_X2 U11 ( .A(A[8]), .B(carry[8]), .ZN(DIFF[8]) );
  INV_X4 U12 ( .A(A[8]), .ZN(n5) );
  INV_X4 U13 ( .A(carry[8]), .ZN(n6) );
  NAND2_X2 U14 ( .A1(n7), .A2(n8), .ZN(carry[10]) );
  XNOR2_X2 U15 ( .A(A[9]), .B(carry[9]), .ZN(DIFF[9]) );
  INV_X4 U16 ( .A(A[9]), .ZN(n7) );
  INV_X4 U17 ( .A(carry[9]), .ZN(n8) );
  NAND2_X2 U18 ( .A1(B[0]), .A2(n9), .ZN(carry[1]) );
  XNOR2_X2 U19 ( .A(n16), .B(A[0]), .ZN(DIFF[0]) );
  INV_X4 U20 ( .A(A[0]), .ZN(n9) );
  INV_X4 U21 ( .A(B[2]), .ZN(n10) );
  INV_X4 U22 ( .A(B[3]), .ZN(n11) );
  INV_X4 U23 ( .A(B[4]), .ZN(n12) );
  INV_X4 U24 ( .A(B[5]), .ZN(n13) );
  INV_X4 U25 ( .A(B[6]), .ZN(n14) );
  INV_X4 U26 ( .A(B[1]), .ZN(n15) );
  INV_X4 U27 ( .A(B[0]), .ZN(n16) );
endmodule


module fpu_DW01_sub_5 ( A, B, CI, DIFF, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;
  wire   [10:1] carry;

  FA_X1 U2_6 ( .A(A[6]), .B(n8), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA_X1 U2_5 ( .A(A[5]), .B(n9), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n10), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_3 ( .A(A[3]), .B(n11), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA_X1 U2_2 ( .A(A[2]), .B(n12), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA_X1 U2_1 ( .A(A[1]), .B(n13), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  XNOR2_X2 U1 ( .A(A[10]), .B(carry[10]), .ZN(DIFF[10]) );
  NAND2_X2 U2 ( .A1(n1), .A2(n2), .ZN(carry[8]) );
  XNOR2_X2 U3 ( .A(A[7]), .B(carry[7]), .ZN(DIFF[7]) );
  INV_X4 U4 ( .A(A[7]), .ZN(n1) );
  INV_X4 U5 ( .A(carry[7]), .ZN(n2) );
  NAND2_X2 U6 ( .A1(n3), .A2(n4), .ZN(carry[9]) );
  XNOR2_X2 U7 ( .A(A[8]), .B(carry[8]), .ZN(DIFF[8]) );
  INV_X4 U8 ( .A(A[8]), .ZN(n3) );
  INV_X4 U9 ( .A(carry[8]), .ZN(n4) );
  NAND2_X2 U10 ( .A1(n5), .A2(n6), .ZN(carry[10]) );
  XNOR2_X2 U11 ( .A(A[9]), .B(carry[9]), .ZN(DIFF[9]) );
  INV_X4 U12 ( .A(A[9]), .ZN(n5) );
  INV_X4 U13 ( .A(carry[9]), .ZN(n6) );
  NAND2_X2 U14 ( .A1(B[0]), .A2(n7), .ZN(carry[1]) );
  XNOR2_X2 U15 ( .A(n14), .B(A[0]), .ZN(DIFF[0]) );
  INV_X4 U16 ( .A(A[0]), .ZN(n7) );
  INV_X4 U17 ( .A(B[6]), .ZN(n8) );
  INV_X4 U18 ( .A(B[5]), .ZN(n9) );
  INV_X4 U19 ( .A(B[4]), .ZN(n10) );
  INV_X4 U20 ( .A(B[3]), .ZN(n11) );
  INV_X4 U21 ( .A(B[2]), .ZN(n12) );
  INV_X4 U22 ( .A(B[1]), .ZN(n13) );
  INV_X4 U23 ( .A(B[0]), .ZN(n14) );
endmodule


module fpu_DW01_add_0 ( A, B, CI, SUM, CO );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  input CI;
  output CO;
  wire   n3, n5;
  wire   [5:2] carry;

  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X2 U1 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  XOR2_X2 U2 ( .A(B[6]), .B(n5), .Z(SUM[6]) );
  AND2_X4 U3 ( .A1(B[0]), .A2(A[0]), .ZN(n3) );
  XOR2_X2 U4 ( .A(B[5]), .B(carry[5]), .Z(SUM[5]) );
  AND2_X4 U5 ( .A1(B[5]), .A2(carry[5]), .ZN(n5) );
endmodule


module fpu_DW01_inc_1 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [10:2] carry;

  HA_X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(SUM[11]), .S(SUM[10]) );
  HA_X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV_X4 U1 ( .A(A[0]), .ZN(SUM[0]) );
endmodule


module fpu_DW01_add_1 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n4, n5, n6;
  wire   [8:2] carry;

  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n4), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X2 U1 ( .A(A[9]), .B(n5), .Z(SUM[9]) );
  XOR2_X2 U2 ( .A(A[10]), .B(n6), .Z(SUM[10]) );
  XOR2_X2 U3 ( .A(A[8]), .B(carry[8]), .Z(SUM[8]) );
  AND2_X4 U4 ( .A1(B[0]), .A2(A[0]), .ZN(n4) );
  AND2_X4 U5 ( .A1(A[8]), .A2(carry[8]), .ZN(n5) );
  AND2_X4 U6 ( .A1(A[9]), .A2(n5), .ZN(n6) );
  XOR2_X2 U7 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module fpu_DW01_inc_2 ( A, SUM );
  input [52:0] A;
  output [52:0] SUM;

  wire   [51:2] carry;

  HA_X1 U1_1_51 ( .A(A[51]), .B(carry[51]), .CO(SUM[52]), .S(SUM[51]) );
  HA_X1 U1_1_50 ( .A(A[50]), .B(carry[50]), .CO(carry[51]), .S(SUM[50]) );
  HA_X1 U1_1_49 ( .A(A[49]), .B(carry[49]), .CO(carry[50]), .S(SUM[49]) );
  HA_X1 U1_1_48 ( .A(A[48]), .B(carry[48]), .CO(carry[49]), .S(SUM[48]) );
  HA_X1 U1_1_47 ( .A(A[47]), .B(carry[47]), .CO(carry[48]), .S(SUM[47]) );
  HA_X1 U1_1_46 ( .A(A[46]), .B(carry[46]), .CO(carry[47]), .S(SUM[46]) );
  HA_X1 U1_1_45 ( .A(A[45]), .B(carry[45]), .CO(carry[46]), .S(SUM[45]) );
  HA_X1 U1_1_44 ( .A(A[44]), .B(carry[44]), .CO(carry[45]), .S(SUM[44]) );
  HA_X1 U1_1_43 ( .A(A[43]), .B(carry[43]), .CO(carry[44]), .S(SUM[43]) );
  HA_X1 U1_1_42 ( .A(A[42]), .B(carry[42]), .CO(carry[43]), .S(SUM[42]) );
  HA_X1 U1_1_41 ( .A(A[41]), .B(carry[41]), .CO(carry[42]), .S(SUM[41]) );
  HA_X1 U1_1_40 ( .A(A[40]), .B(carry[40]), .CO(carry[41]), .S(SUM[40]) );
  HA_X1 U1_1_39 ( .A(A[39]), .B(carry[39]), .CO(carry[40]), .S(SUM[39]) );
  HA_X1 U1_1_38 ( .A(A[38]), .B(carry[38]), .CO(carry[39]), .S(SUM[38]) );
  HA_X1 U1_1_37 ( .A(A[37]), .B(carry[37]), .CO(carry[38]), .S(SUM[37]) );
  HA_X1 U1_1_36 ( .A(A[36]), .B(carry[36]), .CO(carry[37]), .S(SUM[36]) );
  HA_X1 U1_1_35 ( .A(A[35]), .B(carry[35]), .CO(carry[36]), .S(SUM[35]) );
  HA_X1 U1_1_34 ( .A(A[34]), .B(carry[34]), .CO(carry[35]), .S(SUM[34]) );
  HA_X1 U1_1_33 ( .A(A[33]), .B(carry[33]), .CO(carry[34]), .S(SUM[33]) );
  HA_X1 U1_1_32 ( .A(A[32]), .B(carry[32]), .CO(carry[33]), .S(SUM[32]) );
  HA_X1 U1_1_31 ( .A(A[31]), .B(carry[31]), .CO(carry[32]), .S(SUM[31]) );
  HA_X1 U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  HA_X1 U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  HA_X1 U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  HA_X1 U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  HA_X1 U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  HA_X1 U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  HA_X1 U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  HA_X1 U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  HA_X1 U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  HA_X1 U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  HA_X1 U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  HA_X1 U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  HA_X1 U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  HA_X1 U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  HA_X1 U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  HA_X1 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  HA_X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  HA_X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  HA_X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  HA_X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  HA_X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  HA_X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[0]), .ZN(SUM[0]) );
endmodule


module fpu_DW01_sub_9 ( A, B, CI, DIFF, CO );
  input [56:0] A;
  input [56:0] B;
  output [56:0] DIFF;
  input CI;
  output CO;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58;
  wire   [56:1] carry;

  FA_X1 U2_55 ( .A(A[55]), .B(n58), .CI(carry[55]), .CO(carry[56]), .S(
        DIFF[55]) );
  FA_X1 U2_54 ( .A(A[54]), .B(n57), .CI(carry[54]), .CO(carry[55]), .S(
        DIFF[54]) );
  FA_X1 U2_53 ( .A(A[53]), .B(n56), .CI(carry[53]), .CO(carry[54]), .S(
        DIFF[53]) );
  FA_X1 U2_52 ( .A(A[52]), .B(n55), .CI(carry[52]), .CO(carry[53]), .S(
        DIFF[52]) );
  FA_X1 U2_51 ( .A(A[51]), .B(n54), .CI(carry[51]), .CO(carry[52]), .S(
        DIFF[51]) );
  FA_X1 U2_50 ( .A(A[50]), .B(n53), .CI(carry[50]), .CO(carry[51]), .S(
        DIFF[50]) );
  FA_X1 U2_49 ( .A(A[49]), .B(n52), .CI(carry[49]), .CO(carry[50]), .S(
        DIFF[49]) );
  FA_X1 U2_48 ( .A(A[48]), .B(n51), .CI(carry[48]), .CO(carry[49]), .S(
        DIFF[48]) );
  FA_X1 U2_47 ( .A(A[47]), .B(n50), .CI(carry[47]), .CO(carry[48]), .S(
        DIFF[47]) );
  FA_X1 U2_46 ( .A(A[46]), .B(n49), .CI(carry[46]), .CO(carry[47]), .S(
        DIFF[46]) );
  FA_X1 U2_45 ( .A(A[45]), .B(n48), .CI(carry[45]), .CO(carry[46]), .S(
        DIFF[45]) );
  FA_X1 U2_44 ( .A(A[44]), .B(n47), .CI(carry[44]), .CO(carry[45]), .S(
        DIFF[44]) );
  FA_X1 U2_43 ( .A(A[43]), .B(n46), .CI(carry[43]), .CO(carry[44]), .S(
        DIFF[43]) );
  FA_X1 U2_42 ( .A(A[42]), .B(n45), .CI(carry[42]), .CO(carry[43]), .S(
        DIFF[42]) );
  FA_X1 U2_41 ( .A(A[41]), .B(n44), .CI(carry[41]), .CO(carry[42]), .S(
        DIFF[41]) );
  FA_X1 U2_40 ( .A(A[40]), .B(n43), .CI(carry[40]), .CO(carry[41]), .S(
        DIFF[40]) );
  FA_X1 U2_39 ( .A(A[39]), .B(n42), .CI(carry[39]), .CO(carry[40]), .S(
        DIFF[39]) );
  FA_X1 U2_38 ( .A(A[38]), .B(n41), .CI(carry[38]), .CO(carry[39]), .S(
        DIFF[38]) );
  FA_X1 U2_37 ( .A(A[37]), .B(n40), .CI(carry[37]), .CO(carry[38]), .S(
        DIFF[37]) );
  FA_X1 U2_36 ( .A(A[36]), .B(n39), .CI(carry[36]), .CO(carry[37]), .S(
        DIFF[36]) );
  FA_X1 U2_35 ( .A(A[35]), .B(n38), .CI(carry[35]), .CO(carry[36]), .S(
        DIFF[35]) );
  FA_X1 U2_34 ( .A(A[34]), .B(n37), .CI(carry[34]), .CO(carry[35]), .S(
        DIFF[34]) );
  FA_X1 U2_33 ( .A(A[33]), .B(n36), .CI(carry[33]), .CO(carry[34]), .S(
        DIFF[33]) );
  FA_X1 U2_32 ( .A(A[32]), .B(n35), .CI(carry[32]), .CO(carry[33]), .S(
        DIFF[32]) );
  FA_X1 U2_31 ( .A(A[31]), .B(n34), .CI(carry[31]), .CO(carry[32]), .S(
        DIFF[31]) );
  FA_X1 U2_30 ( .A(A[30]), .B(n33), .CI(carry[30]), .CO(carry[31]), .S(
        DIFF[30]) );
  FA_X1 U2_29 ( .A(A[29]), .B(n32), .CI(carry[29]), .CO(carry[30]), .S(
        DIFF[29]) );
  FA_X1 U2_28 ( .A(A[28]), .B(n31), .CI(carry[28]), .CO(carry[29]), .S(
        DIFF[28]) );
  FA_X1 U2_27 ( .A(A[27]), .B(n30), .CI(carry[27]), .CO(carry[28]), .S(
        DIFF[27]) );
  FA_X1 U2_26 ( .A(A[26]), .B(n29), .CI(carry[26]), .CO(carry[27]), .S(
        DIFF[26]) );
  FA_X1 U2_25 ( .A(A[25]), .B(n28), .CI(carry[25]), .CO(carry[26]), .S(
        DIFF[25]) );
  FA_X1 U2_24 ( .A(A[24]), .B(n27), .CI(carry[24]), .CO(carry[25]), .S(
        DIFF[24]) );
  FA_X1 U2_23 ( .A(A[23]), .B(n26), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  FA_X1 U2_22 ( .A(A[22]), .B(n25), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FA_X1 U2_21 ( .A(A[21]), .B(n24), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FA_X1 U2_20 ( .A(A[20]), .B(n23), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FA_X1 U2_19 ( .A(A[19]), .B(n22), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FA_X1 U2_18 ( .A(A[18]), .B(n21), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FA_X1 U2_17 ( .A(A[17]), .B(n20), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FA_X1 U2_16 ( .A(A[16]), .B(n19), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FA_X1 U2_15 ( .A(A[15]), .B(n18), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FA_X1 U2_14 ( .A(A[14]), .B(n17), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FA_X1 U2_13 ( .A(A[13]), .B(n16), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FA_X1 U2_12 ( .A(A[12]), .B(n15), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FA_X1 U2_11 ( .A(A[11]), .B(n14), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FA_X1 U2_10 ( .A(A[10]), .B(n13), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FA_X1 U2_9 ( .A(A[9]), .B(n12), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FA_X1 U2_8 ( .A(A[8]), .B(n11), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FA_X1 U2_7 ( .A(A[7]), .B(n10), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FA_X1 U2_6 ( .A(A[6]), .B(n9), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA_X1 U2_5 ( .A(A[5]), .B(n8), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n7), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_3 ( .A(A[3]), .B(n6), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA_X1 U2_2 ( .A(A[2]), .B(n5), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA_X1 U2_1 ( .A(A[1]), .B(n4), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  NAND2_X2 U1 ( .A1(B[0]), .A2(n1), .ZN(carry[1]) );
  XNOR2_X2 U2 ( .A(n3), .B(A[0]), .ZN(DIFF[0]) );
  INV_X4 U3 ( .A(A[0]), .ZN(n1) );
  INV_X4 U4 ( .A(carry[56]), .ZN(DIFF[56]) );
  INV_X4 U5 ( .A(B[0]), .ZN(n3) );
  INV_X4 U6 ( .A(B[1]), .ZN(n4) );
  INV_X4 U7 ( .A(B[2]), .ZN(n5) );
  INV_X4 U8 ( .A(B[3]), .ZN(n6) );
  INV_X4 U9 ( .A(B[4]), .ZN(n7) );
  INV_X4 U10 ( .A(B[5]), .ZN(n8) );
  INV_X4 U11 ( .A(B[6]), .ZN(n9) );
  INV_X4 U12 ( .A(B[7]), .ZN(n10) );
  INV_X4 U13 ( .A(B[8]), .ZN(n11) );
  INV_X4 U14 ( .A(B[9]), .ZN(n12) );
  INV_X4 U15 ( .A(B[10]), .ZN(n13) );
  INV_X4 U16 ( .A(B[11]), .ZN(n14) );
  INV_X4 U17 ( .A(B[12]), .ZN(n15) );
  INV_X4 U18 ( .A(B[13]), .ZN(n16) );
  INV_X4 U19 ( .A(B[14]), .ZN(n17) );
  INV_X4 U20 ( .A(B[15]), .ZN(n18) );
  INV_X4 U21 ( .A(B[16]), .ZN(n19) );
  INV_X4 U22 ( .A(B[17]), .ZN(n20) );
  INV_X4 U23 ( .A(B[18]), .ZN(n21) );
  INV_X4 U24 ( .A(B[19]), .ZN(n22) );
  INV_X4 U25 ( .A(B[20]), .ZN(n23) );
  INV_X4 U26 ( .A(B[21]), .ZN(n24) );
  INV_X4 U27 ( .A(B[22]), .ZN(n25) );
  INV_X4 U28 ( .A(B[23]), .ZN(n26) );
  INV_X4 U29 ( .A(B[24]), .ZN(n27) );
  INV_X4 U30 ( .A(B[25]), .ZN(n28) );
  INV_X4 U31 ( .A(B[26]), .ZN(n29) );
  INV_X4 U32 ( .A(B[27]), .ZN(n30) );
  INV_X4 U33 ( .A(B[28]), .ZN(n31) );
  INV_X4 U34 ( .A(B[29]), .ZN(n32) );
  INV_X4 U35 ( .A(B[30]), .ZN(n33) );
  INV_X4 U36 ( .A(B[31]), .ZN(n34) );
  INV_X4 U37 ( .A(B[32]), .ZN(n35) );
  INV_X4 U38 ( .A(B[33]), .ZN(n36) );
  INV_X4 U39 ( .A(B[34]), .ZN(n37) );
  INV_X4 U40 ( .A(B[35]), .ZN(n38) );
  INV_X4 U41 ( .A(B[36]), .ZN(n39) );
  INV_X4 U42 ( .A(B[37]), .ZN(n40) );
  INV_X4 U43 ( .A(B[38]), .ZN(n41) );
  INV_X4 U44 ( .A(B[39]), .ZN(n42) );
  INV_X4 U45 ( .A(B[40]), .ZN(n43) );
  INV_X4 U46 ( .A(B[41]), .ZN(n44) );
  INV_X4 U47 ( .A(B[42]), .ZN(n45) );
  INV_X4 U48 ( .A(B[43]), .ZN(n46) );
  INV_X4 U49 ( .A(B[44]), .ZN(n47) );
  INV_X4 U50 ( .A(B[45]), .ZN(n48) );
  INV_X4 U51 ( .A(B[46]), .ZN(n49) );
  INV_X4 U52 ( .A(B[47]), .ZN(n50) );
  INV_X4 U53 ( .A(B[48]), .ZN(n51) );
  INV_X4 U54 ( .A(B[49]), .ZN(n52) );
  INV_X4 U55 ( .A(B[50]), .ZN(n53) );
  INV_X4 U56 ( .A(B[51]), .ZN(n54) );
  INV_X4 U57 ( .A(B[52]), .ZN(n55) );
  INV_X4 U58 ( .A(B[53]), .ZN(n56) );
  INV_X4 U59 ( .A(B[54]), .ZN(n57) );
  INV_X4 U60 ( .A(B[55]), .ZN(n58) );
endmodule


module fpu_DW01_add_4 ( A, B, CI, SUM, CO );
  input [56:0] A;
  input [56:0] B;
  output [56:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [55:2] carry;

  FA_X1 U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(SUM[56]), .S(SUM[55]) );
  FA_X1 U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  FA_X1 U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  FA_X1 U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  FA_X1 U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  FA_X1 U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  FA_X1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FA_X1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FA_X1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FA_X1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FA_X1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FA_X1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FA_X1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FA_X1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FA_X1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FA_X1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FA_X1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FA_X1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FA_X1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FA_X1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FA_X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FA_X1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FA_X1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FA_X1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X2 U1 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X4 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
endmodule


module fpu_DW01_inc_3 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HA_X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV_X4 U1 ( .A(A[0]), .ZN(SUM[0]) );
  XOR2_X1 U2 ( .A(carry[10]), .B(A[10]), .Z(SUM[10]) );
endmodule


module fpu_DW01_inc_4 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HA_X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV_X4 U1 ( .A(A[0]), .ZN(SUM[0]) );
  XOR2_X1 U2 ( .A(carry[10]), .B(A[10]), .Z(SUM[10]) );
endmodule


module fpu_DW01_add_6 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [10:2] carry;

  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(SUM[11]), .S(SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X2 U1 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X4 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
endmodule


module fpu_DW01_sub_12 ( A, B, CI, DIFF, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] DIFF;
  input CI;
  output CO;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;
  wire   [11:1] carry;

  FA_X1 U2_10 ( .A(A[10]), .B(n3), .CI(carry[10]), .CO(carry[11]), .S(DIFF[10]) );
  FA_X1 U2_9 ( .A(A[9]), .B(n4), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9]) );
  FA_X1 U2_8 ( .A(A[8]), .B(n5), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FA_X1 U2_7 ( .A(A[7]), .B(n6), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FA_X1 U2_6 ( .A(A[6]), .B(n7), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA_X1 U2_5 ( .A(A[5]), .B(n8), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n9), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_3 ( .A(A[3]), .B(n10), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA_X1 U2_2 ( .A(A[2]), .B(n11), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA_X1 U2_1 ( .A(A[1]), .B(n12), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  NAND2_X2 U1 ( .A1(B[0]), .A2(n1), .ZN(carry[1]) );
  XNOR2_X2 U2 ( .A(n13), .B(A[0]), .ZN(DIFF[0]) );
  INV_X4 U3 ( .A(A[0]), .ZN(n1) );
  INV_X4 U4 ( .A(carry[11]), .ZN(DIFF[11]) );
  INV_X4 U5 ( .A(B[10]), .ZN(n3) );
  INV_X4 U6 ( .A(B[9]), .ZN(n4) );
  INV_X4 U7 ( .A(B[8]), .ZN(n5) );
  INV_X4 U8 ( .A(B[7]), .ZN(n6) );
  INV_X4 U9 ( .A(B[6]), .ZN(n7) );
  INV_X4 U10 ( .A(B[5]), .ZN(n8) );
  INV_X4 U11 ( .A(B[4]), .ZN(n9) );
  INV_X4 U12 ( .A(B[3]), .ZN(n10) );
  INV_X4 U13 ( .A(B[2]), .ZN(n11) );
  INV_X4 U14 ( .A(B[1]), .ZN(n12) );
  INV_X4 U15 ( .A(B[0]), .ZN(n13) );
endmodule


module fpu_DW01_cmp2_13 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [55:0] A;
  input [55:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167;

  INV_X4 U1 ( .A(B[9]), .ZN(n1) );
  INV_X4 U2 ( .A(B[8]), .ZN(n2) );
  INV_X4 U3 ( .A(B[7]), .ZN(n3) );
  INV_X4 U4 ( .A(B[6]), .ZN(n4) );
  INV_X4 U5 ( .A(B[5]), .ZN(n5) );
  INV_X4 U6 ( .A(B[55]), .ZN(n6) );
  INV_X4 U7 ( .A(B[54]), .ZN(n7) );
  INV_X4 U8 ( .A(B[53]), .ZN(n8) );
  INV_X4 U9 ( .A(B[52]), .ZN(n9) );
  INV_X4 U10 ( .A(B[51]), .ZN(n10) );
  INV_X4 U11 ( .A(B[50]), .ZN(n11) );
  INV_X4 U12 ( .A(B[4]), .ZN(n12) );
  INV_X4 U13 ( .A(B[49]), .ZN(n13) );
  INV_X4 U14 ( .A(B[48]), .ZN(n14) );
  INV_X4 U15 ( .A(B[47]), .ZN(n15) );
  INV_X4 U16 ( .A(B[46]), .ZN(n16) );
  INV_X4 U17 ( .A(B[45]), .ZN(n17) );
  INV_X4 U18 ( .A(B[44]), .ZN(n18) );
  INV_X4 U19 ( .A(B[43]), .ZN(n19) );
  INV_X4 U20 ( .A(B[42]), .ZN(n20) );
  INV_X4 U21 ( .A(B[41]), .ZN(n21) );
  INV_X4 U22 ( .A(B[40]), .ZN(n22) );
  INV_X4 U23 ( .A(B[3]), .ZN(n23) );
  INV_X4 U24 ( .A(B[39]), .ZN(n24) );
  INV_X4 U25 ( .A(B[38]), .ZN(n25) );
  INV_X4 U26 ( .A(B[37]), .ZN(n26) );
  INV_X4 U27 ( .A(B[36]), .ZN(n27) );
  INV_X4 U28 ( .A(B[35]), .ZN(n28) );
  INV_X4 U29 ( .A(B[34]), .ZN(n29) );
  INV_X4 U30 ( .A(B[33]), .ZN(n30) );
  INV_X4 U31 ( .A(B[32]), .ZN(n31) );
  INV_X4 U32 ( .A(B[31]), .ZN(n32) );
  INV_X4 U33 ( .A(B[30]), .ZN(n33) );
  INV_X4 U34 ( .A(B[29]), .ZN(n34) );
  INV_X4 U35 ( .A(B[28]), .ZN(n35) );
  INV_X4 U36 ( .A(B[27]), .ZN(n36) );
  INV_X4 U37 ( .A(B[26]), .ZN(n37) );
  INV_X4 U38 ( .A(B[25]), .ZN(n38) );
  INV_X4 U39 ( .A(B[24]), .ZN(n39) );
  INV_X4 U40 ( .A(B[23]), .ZN(n40) );
  INV_X4 U41 ( .A(B[22]), .ZN(n41) );
  INV_X4 U42 ( .A(B[21]), .ZN(n42) );
  INV_X4 U43 ( .A(B[20]), .ZN(n43) );
  INV_X4 U44 ( .A(B[19]), .ZN(n44) );
  INV_X4 U45 ( .A(B[18]), .ZN(n45) );
  INV_X4 U46 ( .A(B[17]), .ZN(n46) );
  INV_X4 U47 ( .A(B[16]), .ZN(n47) );
  INV_X4 U48 ( .A(B[15]), .ZN(n48) );
  INV_X4 U49 ( .A(B[14]), .ZN(n49) );
  INV_X4 U50 ( .A(B[13]), .ZN(n50) );
  INV_X4 U51 ( .A(B[12]), .ZN(n51) );
  INV_X4 U52 ( .A(B[11]), .ZN(n52) );
  INV_X4 U53 ( .A(B[10]), .ZN(n53) );
  INV_X4 U54 ( .A(A[9]), .ZN(n54) );
  INV_X4 U55 ( .A(A[8]), .ZN(n55) );
  INV_X4 U56 ( .A(A[7]), .ZN(n56) );
  INV_X4 U57 ( .A(A[6]), .ZN(n57) );
  INV_X4 U58 ( .A(A[5]), .ZN(n58) );
  INV_X4 U59 ( .A(A[55]), .ZN(n59) );
  INV_X4 U60 ( .A(A[53]), .ZN(n60) );
  INV_X4 U61 ( .A(A[52]), .ZN(n61) );
  INV_X4 U62 ( .A(A[51]), .ZN(n62) );
  INV_X4 U63 ( .A(A[50]), .ZN(n63) );
  INV_X4 U64 ( .A(A[4]), .ZN(n64) );
  INV_X4 U65 ( .A(A[49]), .ZN(n65) );
  INV_X4 U66 ( .A(A[48]), .ZN(n66) );
  INV_X4 U67 ( .A(A[47]), .ZN(n67) );
  INV_X4 U68 ( .A(A[46]), .ZN(n68) );
  INV_X4 U69 ( .A(A[45]), .ZN(n69) );
  INV_X4 U70 ( .A(A[44]), .ZN(n70) );
  INV_X4 U71 ( .A(A[43]), .ZN(n71) );
  INV_X4 U72 ( .A(A[42]), .ZN(n72) );
  INV_X4 U73 ( .A(A[41]), .ZN(n73) );
  INV_X4 U74 ( .A(A[40]), .ZN(n74) );
  INV_X4 U75 ( .A(A[3]), .ZN(n75) );
  INV_X4 U76 ( .A(A[39]), .ZN(n76) );
  INV_X4 U77 ( .A(A[38]), .ZN(n77) );
  INV_X4 U78 ( .A(A[37]), .ZN(n78) );
  INV_X4 U79 ( .A(A[36]), .ZN(n79) );
  INV_X4 U80 ( .A(A[35]), .ZN(n80) );
  INV_X4 U81 ( .A(A[34]), .ZN(n81) );
  INV_X4 U82 ( .A(A[33]), .ZN(n82) );
  INV_X4 U83 ( .A(A[32]), .ZN(n83) );
  INV_X4 U84 ( .A(A[31]), .ZN(n84) );
  INV_X4 U85 ( .A(A[30]), .ZN(n85) );
  INV_X4 U86 ( .A(A[2]), .ZN(n86) );
  INV_X4 U87 ( .A(A[29]), .ZN(n87) );
  INV_X4 U88 ( .A(A[28]), .ZN(n88) );
  INV_X4 U89 ( .A(A[27]), .ZN(n89) );
  INV_X4 U90 ( .A(A[26]), .ZN(n90) );
  INV_X4 U91 ( .A(A[25]), .ZN(n91) );
  INV_X4 U92 ( .A(A[24]), .ZN(n92) );
  INV_X4 U93 ( .A(A[23]), .ZN(n93) );
  INV_X4 U94 ( .A(A[22]), .ZN(n94) );
  INV_X4 U95 ( .A(A[21]), .ZN(n95) );
  INV_X4 U96 ( .A(A[20]), .ZN(n96) );
  INV_X4 U97 ( .A(A[1]), .ZN(n97) );
  INV_X4 U98 ( .A(A[19]), .ZN(n98) );
  INV_X4 U99 ( .A(A[18]), .ZN(n99) );
  INV_X4 U100 ( .A(A[17]), .ZN(n100) );
  INV_X4 U101 ( .A(A[16]), .ZN(n101) );
  INV_X4 U102 ( .A(A[15]), .ZN(n102) );
  INV_X4 U103 ( .A(A[14]), .ZN(n103) );
  INV_X4 U104 ( .A(A[13]), .ZN(n104) );
  INV_X4 U105 ( .A(A[12]), .ZN(n105) );
  INV_X4 U106 ( .A(A[11]), .ZN(n106) );
  INV_X4 U107 ( .A(A[10]), .ZN(n107) );
  INV_X4 U108 ( .A(n167), .ZN(n108) );
  INV_X4 U109 ( .A(B[0]), .ZN(n109) );
  INV_X4 U110 ( .A(B[2]), .ZN(n110) );
  OAI21_X1 U111 ( .B1(A[55]), .B2(n6), .A(n111), .ZN(LT_LE) );
  OAI22_X1 U112 ( .A1(n112), .A2(n113), .B1(B[55]), .B2(n59), .ZN(n111) );
  AOI221_X1 U113 ( .B1(A[54]), .B2(n7), .C1(A[53]), .C2(n8), .A(n114), .ZN(
        n113) );
  AOI221_X1 U114 ( .B1(B[53]), .B2(n60), .C1(B[52]), .C2(n61), .A(n115), .ZN(
        n114) );
  AOI221_X1 U115 ( .B1(A[52]), .B2(n9), .C1(A[51]), .C2(n10), .A(n116), .ZN(
        n115) );
  AOI221_X1 U116 ( .B1(B[51]), .B2(n62), .C1(B[50]), .C2(n63), .A(n117), .ZN(
        n116) );
  AOI221_X1 U117 ( .B1(A[50]), .B2(n11), .C1(A[49]), .C2(n13), .A(n118), .ZN(
        n117) );
  AOI221_X1 U118 ( .B1(B[49]), .B2(n65), .C1(B[48]), .C2(n66), .A(n119), .ZN(
        n118) );
  AOI221_X1 U119 ( .B1(A[48]), .B2(n14), .C1(A[47]), .C2(n15), .A(n120), .ZN(
        n119) );
  AOI221_X1 U120 ( .B1(B[47]), .B2(n67), .C1(B[46]), .C2(n68), .A(n121), .ZN(
        n120) );
  AOI221_X1 U121 ( .B1(A[46]), .B2(n16), .C1(A[45]), .C2(n17), .A(n122), .ZN(
        n121) );
  AOI221_X1 U122 ( .B1(B[45]), .B2(n69), .C1(B[44]), .C2(n70), .A(n123), .ZN(
        n122) );
  AOI221_X1 U123 ( .B1(A[44]), .B2(n18), .C1(A[43]), .C2(n19), .A(n124), .ZN(
        n123) );
  AOI221_X1 U124 ( .B1(B[43]), .B2(n71), .C1(B[42]), .C2(n72), .A(n125), .ZN(
        n124) );
  AOI221_X1 U125 ( .B1(A[42]), .B2(n20), .C1(A[41]), .C2(n21), .A(n126), .ZN(
        n125) );
  AOI221_X1 U126 ( .B1(B[41]), .B2(n73), .C1(B[40]), .C2(n74), .A(n127), .ZN(
        n126) );
  AOI221_X1 U127 ( .B1(A[40]), .B2(n22), .C1(A[39]), .C2(n24), .A(n128), .ZN(
        n127) );
  AOI221_X1 U128 ( .B1(B[39]), .B2(n76), .C1(B[38]), .C2(n77), .A(n129), .ZN(
        n128) );
  AOI221_X1 U129 ( .B1(A[38]), .B2(n25), .C1(A[37]), .C2(n26), .A(n130), .ZN(
        n129) );
  AOI221_X1 U130 ( .B1(B[37]), .B2(n78), .C1(B[36]), .C2(n79), .A(n131), .ZN(
        n130) );
  AOI221_X1 U131 ( .B1(A[36]), .B2(n27), .C1(A[35]), .C2(n28), .A(n132), .ZN(
        n131) );
  AOI221_X1 U132 ( .B1(B[35]), .B2(n80), .C1(B[34]), .C2(n81), .A(n133), .ZN(
        n132) );
  AOI221_X1 U133 ( .B1(A[34]), .B2(n29), .C1(A[33]), .C2(n30), .A(n134), .ZN(
        n133) );
  AOI221_X1 U134 ( .B1(B[33]), .B2(n82), .C1(B[32]), .C2(n83), .A(n135), .ZN(
        n134) );
  AOI221_X1 U135 ( .B1(A[32]), .B2(n31), .C1(A[31]), .C2(n32), .A(n136), .ZN(
        n135) );
  AOI221_X1 U136 ( .B1(B[31]), .B2(n84), .C1(B[30]), .C2(n85), .A(n137), .ZN(
        n136) );
  AOI221_X1 U137 ( .B1(A[30]), .B2(n33), .C1(A[29]), .C2(n34), .A(n138), .ZN(
        n137) );
  AOI221_X1 U138 ( .B1(B[29]), .B2(n87), .C1(B[28]), .C2(n88), .A(n139), .ZN(
        n138) );
  AOI221_X1 U139 ( .B1(A[28]), .B2(n35), .C1(A[27]), .C2(n36), .A(n140), .ZN(
        n139) );
  AOI221_X1 U140 ( .B1(B[27]), .B2(n89), .C1(B[26]), .C2(n90), .A(n141), .ZN(
        n140) );
  AOI221_X1 U141 ( .B1(A[26]), .B2(n37), .C1(A[25]), .C2(n38), .A(n142), .ZN(
        n141) );
  AOI221_X1 U142 ( .B1(B[25]), .B2(n91), .C1(B[24]), .C2(n92), .A(n143), .ZN(
        n142) );
  AOI221_X1 U143 ( .B1(A[24]), .B2(n39), .C1(A[23]), .C2(n40), .A(n144), .ZN(
        n143) );
  AOI221_X1 U144 ( .B1(B[23]), .B2(n93), .C1(B[22]), .C2(n94), .A(n145), .ZN(
        n144) );
  AOI221_X1 U145 ( .B1(A[22]), .B2(n41), .C1(A[21]), .C2(n42), .A(n146), .ZN(
        n145) );
  AOI221_X1 U146 ( .B1(B[21]), .B2(n95), .C1(B[20]), .C2(n96), .A(n147), .ZN(
        n146) );
  AOI221_X1 U147 ( .B1(A[20]), .B2(n43), .C1(A[19]), .C2(n44), .A(n148), .ZN(
        n147) );
  AOI221_X1 U148 ( .B1(B[19]), .B2(n98), .C1(B[18]), .C2(n99), .A(n149), .ZN(
        n148) );
  AOI221_X1 U149 ( .B1(A[18]), .B2(n45), .C1(A[17]), .C2(n46), .A(n150), .ZN(
        n149) );
  AOI221_X1 U150 ( .B1(B[17]), .B2(n100), .C1(B[16]), .C2(n101), .A(n151), 
        .ZN(n150) );
  AOI221_X1 U151 ( .B1(A[16]), .B2(n47), .C1(A[15]), .C2(n48), .A(n152), .ZN(
        n151) );
  AOI221_X1 U152 ( .B1(B[15]), .B2(n102), .C1(B[14]), .C2(n103), .A(n153), 
        .ZN(n152) );
  AOI221_X1 U153 ( .B1(A[14]), .B2(n49), .C1(A[13]), .C2(n50), .A(n154), .ZN(
        n153) );
  AOI221_X1 U154 ( .B1(B[13]), .B2(n104), .C1(B[12]), .C2(n105), .A(n155), 
        .ZN(n154) );
  AOI221_X1 U155 ( .B1(A[12]), .B2(n51), .C1(A[11]), .C2(n52), .A(n156), .ZN(
        n155) );
  AOI221_X1 U156 ( .B1(B[11]), .B2(n106), .C1(B[10]), .C2(n107), .A(n157), 
        .ZN(n156) );
  AOI221_X1 U157 ( .B1(A[9]), .B2(n1), .C1(A[10]), .C2(n53), .A(n158), .ZN(
        n157) );
  AOI221_X1 U158 ( .B1(B[9]), .B2(n54), .C1(B[8]), .C2(n55), .A(n159), .ZN(
        n158) );
  AOI221_X1 U159 ( .B1(A[8]), .B2(n2), .C1(A[7]), .C2(n3), .A(n160), .ZN(n159)
         );
  AOI221_X1 U160 ( .B1(B[7]), .B2(n56), .C1(B[6]), .C2(n57), .A(n161), .ZN(
        n160) );
  AOI221_X1 U161 ( .B1(A[6]), .B2(n4), .C1(A[5]), .C2(n5), .A(n162), .ZN(n161)
         );
  AOI221_X1 U162 ( .B1(B[5]), .B2(n58), .C1(B[4]), .C2(n64), .A(n163), .ZN(
        n162) );
  AOI221_X1 U163 ( .B1(A[4]), .B2(n12), .C1(A[3]), .C2(n23), .A(n164), .ZN(
        n163) );
  AOI221_X1 U164 ( .B1(B[3]), .B2(n75), .C1(B[2]), .C2(n86), .A(n165), .ZN(
        n164) );
  AOI221_X1 U165 ( .B1(A[2]), .B2(n110), .C1(A[1]), .C2(n108), .A(n166), .ZN(
        n165) );
  AOI21_X1 U166 ( .B1(n167), .B2(n97), .A(B[1]), .ZN(n166) );
  NOR2_X1 U167 ( .A1(n109), .A2(A[0]), .ZN(n167) );
  NOR2_X1 U168 ( .A1(A[54]), .A2(n7), .ZN(n112) );
endmodule


module fpu_DW_rash_1 ( A, DATA_TC, SH, SH_TC, B );
  input [55:0] A;
  input [5:0] SH;
  output [55:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360;

  NOR2_X2 U3 ( .A1(n94), .A2(n59), .ZN(n237) );
  NOR2_X2 U4 ( .A1(n19), .A2(n8), .ZN(n146) );
  INV_X4 U5 ( .A(n237), .ZN(n58) );
  NOR2_X2 U6 ( .A1(n5), .A2(n8), .ZN(n143) );
  NOR2_X2 U7 ( .A1(n8), .A2(n58), .ZN(n141) );
  NOR2_X2 U8 ( .A1(n98), .A2(SH[4]), .ZN(n145) );
  OR2_X4 U9 ( .A1(n59), .A2(SH[3]), .ZN(n1) );
  NOR2_X2 U10 ( .A1(SH[2]), .A2(SH[3]), .ZN(n2) );
  NAND2_X2 U11 ( .A1(SH[1]), .A2(n93), .ZN(n3) );
  AND2_X4 U12 ( .A1(n97), .A2(n98), .ZN(n4) );
  NOR2_X2 U13 ( .A1(n93), .A2(SH[1]), .ZN(n224) );
  INV_X4 U14 ( .A(n19), .ZN(n18) );
  INV_X4 U15 ( .A(n3), .ZN(n13) );
  INV_X4 U16 ( .A(n198), .ZN(n14) );
  NOR2_X2 U17 ( .A1(n94), .A2(SH[2]), .ZN(n196) );
  INV_X4 U18 ( .A(n2), .ZN(n19) );
  INV_X4 U19 ( .A(n4), .ZN(n8) );
  INV_X4 U20 ( .A(n199), .ZN(n17) );
  INV_X4 U21 ( .A(n1), .ZN(n10) );
  INV_X4 U22 ( .A(n1), .ZN(n11) );
  INV_X4 U23 ( .A(n224), .ZN(n7) );
  INV_X4 U24 ( .A(n163), .ZN(n96) );
  NOR2_X2 U25 ( .A1(n1), .A2(n9), .ZN(n139) );
  INV_X4 U26 ( .A(n196), .ZN(n5) );
  INV_X4 U27 ( .A(n17), .ZN(n16) );
  INV_X4 U28 ( .A(n13), .ZN(n12) );
  INV_X4 U29 ( .A(n14), .ZN(n15) );
  INV_X4 U30 ( .A(n224), .ZN(n6) );
  INV_X4 U31 ( .A(n4), .ZN(n9) );
  INV_X4 U32 ( .A(n289), .ZN(n20) );
  INV_X4 U33 ( .A(n356), .ZN(n21) );
  INV_X4 U34 ( .A(n215), .ZN(n22) );
  INV_X4 U35 ( .A(n343), .ZN(n23) );
  INV_X4 U36 ( .A(n272), .ZN(n24) );
  INV_X4 U37 ( .A(n146), .ZN(n25) );
  INV_X4 U38 ( .A(n230), .ZN(n26) );
  INV_X4 U39 ( .A(n217), .ZN(n27) );
  INV_X4 U40 ( .A(n191), .ZN(n28) );
  INV_X4 U41 ( .A(n190), .ZN(n29) );
  INV_X4 U42 ( .A(n189), .ZN(n30) );
  INV_X4 U43 ( .A(n188), .ZN(n31) );
  INV_X4 U44 ( .A(n214), .ZN(n32) );
  INV_X4 U45 ( .A(n277), .ZN(n33) );
  INV_X4 U46 ( .A(n213), .ZN(n34) );
  INV_X4 U47 ( .A(n226), .ZN(n35) );
  INV_X4 U48 ( .A(n202), .ZN(n36) );
  INV_X4 U49 ( .A(n201), .ZN(n37) );
  INV_X4 U50 ( .A(n210), .ZN(n38) );
  INV_X4 U51 ( .A(n185), .ZN(n39) );
  INV_X4 U52 ( .A(n208), .ZN(n40) );
  INV_X4 U53 ( .A(n175), .ZN(n41) );
  INV_X4 U54 ( .A(n206), .ZN(n42) );
  INV_X4 U55 ( .A(n171), .ZN(n43) );
  INV_X4 U56 ( .A(n203), .ZN(n44) );
  INV_X4 U57 ( .A(n164), .ZN(n45) );
  INV_X4 U58 ( .A(n156), .ZN(n46) );
  INV_X4 U59 ( .A(n148), .ZN(n47) );
  INV_X4 U60 ( .A(n337), .ZN(n48) );
  INV_X4 U61 ( .A(n311), .ZN(n49) );
  INV_X4 U62 ( .A(n295), .ZN(n50) );
  INV_X4 U63 ( .A(n287), .ZN(n51) );
  INV_X4 U64 ( .A(n284), .ZN(n52) );
  INV_X4 U65 ( .A(n268), .ZN(n53) );
  INV_X4 U66 ( .A(n264), .ZN(n54) );
  INV_X4 U67 ( .A(n257), .ZN(n55) );
  INV_X4 U68 ( .A(n244), .ZN(n56) );
  INV_X4 U69 ( .A(n236), .ZN(n57) );
  INV_X4 U70 ( .A(SH[2]), .ZN(n59) );
  INV_X4 U71 ( .A(n270), .ZN(n60) );
  INV_X4 U72 ( .A(n352), .ZN(n61) );
  INV_X4 U73 ( .A(n312), .ZN(n62) );
  INV_X4 U74 ( .A(n351), .ZN(n63) );
  INV_X4 U75 ( .A(n241), .ZN(n64) );
  INV_X4 U76 ( .A(n349), .ZN(n65) );
  INV_X4 U77 ( .A(n179), .ZN(n66) );
  INV_X4 U78 ( .A(n348), .ZN(n67) );
  INV_X4 U79 ( .A(n263), .ZN(n68) );
  INV_X4 U80 ( .A(n336), .ZN(n69) );
  INV_X4 U81 ( .A(n286), .ZN(n70) );
  INV_X4 U82 ( .A(n335), .ZN(n71) );
  INV_X4 U83 ( .A(n177), .ZN(n72) );
  INV_X4 U84 ( .A(n262), .ZN(n73) );
  INV_X4 U85 ( .A(n334), .ZN(n74) );
  INV_X4 U86 ( .A(n279), .ZN(n75) );
  INV_X4 U87 ( .A(n248), .ZN(n76) );
  INV_X4 U88 ( .A(n283), .ZN(n77) );
  INV_X4 U89 ( .A(n324), .ZN(n78) );
  INV_X4 U90 ( .A(n281), .ZN(n79) );
  INV_X4 U91 ( .A(n254), .ZN(n80) );
  INV_X4 U92 ( .A(n321), .ZN(n81) );
  INV_X4 U93 ( .A(n320), .ZN(n82) );
  INV_X4 U94 ( .A(n319), .ZN(n83) );
  INV_X4 U95 ( .A(n161), .ZN(n84) );
  INV_X4 U96 ( .A(n267), .ZN(n85) );
  INV_X4 U97 ( .A(n306), .ZN(n86) );
  INV_X4 U98 ( .A(n238), .ZN(n87) );
  INV_X4 U99 ( .A(n233), .ZN(n88) );
  INV_X4 U100 ( .A(n303), .ZN(n89) );
  INV_X4 U101 ( .A(n178), .ZN(n90) );
  INV_X4 U102 ( .A(n266), .ZN(n91) );
  INV_X4 U103 ( .A(n302), .ZN(n92) );
  INV_X4 U104 ( .A(SH[0]), .ZN(n93) );
  INV_X4 U105 ( .A(SH[3]), .ZN(n94) );
  INV_X4 U106 ( .A(n145), .ZN(n95) );
  INV_X4 U107 ( .A(SH[4]), .ZN(n97) );
  INV_X4 U108 ( .A(SH[5]), .ZN(n98) );
  INV_X4 U109 ( .A(A[12]), .ZN(n99) );
  INV_X4 U110 ( .A(A[11]), .ZN(n100) );
  INV_X4 U111 ( .A(A[10]), .ZN(n101) );
  INV_X4 U112 ( .A(A[9]), .ZN(n102) );
  INV_X4 U113 ( .A(A[8]), .ZN(n103) );
  INV_X4 U114 ( .A(A[7]), .ZN(n104) );
  INV_X4 U115 ( .A(A[6]), .ZN(n105) );
  INV_X4 U116 ( .A(A[40]), .ZN(n106) );
  INV_X4 U117 ( .A(A[39]), .ZN(n107) );
  INV_X4 U118 ( .A(A[38]), .ZN(n108) );
  INV_X4 U119 ( .A(A[37]), .ZN(n109) );
  INV_X4 U120 ( .A(A[36]), .ZN(n110) );
  INV_X4 U121 ( .A(A[35]), .ZN(n111) );
  INV_X4 U122 ( .A(A[34]), .ZN(n112) );
  INV_X4 U123 ( .A(A[33]), .ZN(n113) );
  INV_X4 U124 ( .A(A[5]), .ZN(n114) );
  INV_X4 U125 ( .A(A[32]), .ZN(n115) );
  INV_X4 U126 ( .A(A[31]), .ZN(n116) );
  INV_X4 U127 ( .A(A[30]), .ZN(n117) );
  INV_X4 U128 ( .A(A[29]), .ZN(n118) );
  INV_X4 U129 ( .A(A[28]), .ZN(n119) );
  INV_X4 U130 ( .A(A[27]), .ZN(n120) );
  INV_X4 U131 ( .A(A[26]), .ZN(n121) );
  INV_X4 U132 ( .A(A[25]), .ZN(n122) );
  INV_X4 U133 ( .A(A[24]), .ZN(n123) );
  INV_X4 U134 ( .A(A[23]), .ZN(n124) );
  INV_X4 U135 ( .A(A[4]), .ZN(n125) );
  INV_X4 U136 ( .A(A[22]), .ZN(n126) );
  INV_X4 U137 ( .A(A[21]), .ZN(n127) );
  INV_X4 U138 ( .A(A[20]), .ZN(n128) );
  INV_X4 U139 ( .A(A[19]), .ZN(n129) );
  INV_X4 U140 ( .A(A[18]), .ZN(n130) );
  INV_X4 U141 ( .A(A[17]), .ZN(n131) );
  INV_X4 U142 ( .A(A[16]), .ZN(n132) );
  INV_X4 U143 ( .A(A[15]), .ZN(n133) );
  INV_X4 U144 ( .A(A[14]), .ZN(n134) );
  INV_X4 U145 ( .A(A[13]), .ZN(n135) );
  OAI211_X1 U146 ( .C1(n136), .C2(n96), .A(n137), .B(n138), .ZN(B[9]) );
  AOI222_X1 U147 ( .A1(n139), .A2(n140), .B1(n141), .B2(n142), .C1(n143), .C2(
        n144), .ZN(n138) );
  AOI22_X1 U148 ( .A1(n145), .A2(n47), .B1(n146), .B2(n147), .ZN(n137) );
  OAI211_X1 U149 ( .C1(n149), .C2(n96), .A(n150), .B(n151), .ZN(B[8]) );
  AOI222_X1 U150 ( .A1(n139), .A2(n152), .B1(n141), .B2(n153), .C1(n143), .C2(
        n154), .ZN(n151) );
  AOI22_X1 U151 ( .A1(n145), .A2(n46), .B1(n146), .B2(n155), .ZN(n150) );
  OAI211_X1 U152 ( .C1(n44), .C2(n98), .A(n157), .B(n158), .ZN(B[7]) );
  AOI222_X1 U153 ( .A1(n139), .A2(n159), .B1(n141), .B2(n160), .C1(n143), .C2(
        n161), .ZN(n158) );
  AOI22_X1 U154 ( .A1(n146), .A2(n162), .B1(n163), .B2(n45), .ZN(n157) );
  OAI211_X1 U155 ( .C1(n42), .C2(n98), .A(n165), .B(n166), .ZN(B[6]) );
  AOI222_X1 U156 ( .A1(n139), .A2(n167), .B1(n141), .B2(n168), .C1(n143), .C2(
        n169), .ZN(n166) );
  AOI22_X1 U157 ( .A1(n146), .A2(n170), .B1(n163), .B2(n43), .ZN(n165) );
  OAI211_X1 U158 ( .C1(n40), .C2(n98), .A(n172), .B(n173), .ZN(B[5]) );
  AOI222_X1 U159 ( .A1(n139), .A2(n147), .B1(n141), .B2(n144), .C1(n143), .C2(
        n140), .ZN(n173) );
  AOI22_X1 U160 ( .A1(n146), .A2(n174), .B1(n163), .B2(n41), .ZN(n172) );
  NOR2_X1 U161 ( .A1(n25), .A2(n176), .ZN(B[55]) );
  NOR2_X1 U162 ( .A1(n177), .A2(n25), .ZN(B[54]) );
  NOR2_X1 U163 ( .A1(n178), .A2(n25), .ZN(B[53]) );
  NOR2_X1 U164 ( .A1(n179), .A2(n25), .ZN(B[52]) );
  NOR2_X1 U165 ( .A1(n8), .A2(n180), .ZN(B[51]) );
  NOR2_X1 U166 ( .A1(n181), .A2(n8), .ZN(B[50]) );
  OAI211_X1 U167 ( .C1(n38), .C2(n98), .A(n182), .B(n183), .ZN(B[4]) );
  AOI222_X1 U168 ( .A1(n139), .A2(n155), .B1(n141), .B2(n154), .C1(n143), .C2(
        n152), .ZN(n183) );
  AOI22_X1 U169 ( .A1(n146), .A2(n184), .B1(n163), .B2(n39), .ZN(n182) );
  NOR2_X1 U170 ( .A1(n186), .A2(n8), .ZN(B[49]) );
  NOR2_X1 U171 ( .A1(n187), .A2(n8), .ZN(B[48]) );
  NOR2_X1 U172 ( .A1(n27), .A2(n8), .ZN(B[47]) );
  NOR2_X1 U173 ( .A1(n188), .A2(n8), .ZN(B[46]) );
  NOR2_X1 U174 ( .A1(n189), .A2(n8), .ZN(B[45]) );
  NOR2_X1 U175 ( .A1(n190), .A2(n8), .ZN(B[44]) );
  NOR2_X1 U176 ( .A1(n26), .A2(n8), .ZN(B[43]) );
  NOR2_X1 U177 ( .A1(n191), .A2(n8), .ZN(B[42]) );
  NOR2_X1 U178 ( .A1(n148), .A2(n8), .ZN(B[41]) );
  NOR2_X1 U179 ( .A1(n156), .A2(n8), .ZN(B[40]) );
  MUX2_X1 U180 ( .A(n36), .B(n192), .S(n98), .Z(B[3]) );
  MUX2_X1 U181 ( .A(n37), .B(n193), .S(n97), .Z(n192) );
  OAI221_X1 U182 ( .B1(n194), .B2(n19), .C1(n84), .C2(n58), .A(n195), .ZN(n193) );
  AOI22_X1 U183 ( .A1(n196), .A2(n159), .B1(n11), .B2(n162), .ZN(n195) );
  OAI221_X1 U184 ( .B1(n6), .B2(n103), .C1(n12), .C2(n102), .A(n197), .ZN(n162) );
  AOI22_X1 U185 ( .A1(A[10]), .A2(n198), .B1(A[7]), .B2(n16), .ZN(n197) );
  AOI221_X1 U186 ( .B1(A[6]), .B2(n15), .C1(A[3]), .C2(n199), .A(n200), .ZN(
        n194) );
  OAI22_X1 U187 ( .A1(n3), .A2(n114), .B1(n6), .B2(n125), .ZN(n200) );
  NOR2_X1 U188 ( .A1(SH[5]), .A2(n44), .ZN(B[39]) );
  OAI22_X1 U189 ( .A1(SH[4]), .A2(n204), .B1(n205), .B2(n176), .ZN(n203) );
  NOR2_X1 U190 ( .A1(SH[5]), .A2(n42), .ZN(B[38]) );
  OAI22_X1 U191 ( .A1(SH[4]), .A2(n207), .B1(n177), .B2(n205), .ZN(n206) );
  NOR2_X1 U192 ( .A1(SH[5]), .A2(n40), .ZN(B[37]) );
  OAI22_X1 U193 ( .A1(SH[4]), .A2(n209), .B1(n178), .B2(n205), .ZN(n208) );
  NOR2_X1 U194 ( .A1(SH[5]), .A2(n38), .ZN(B[36]) );
  OAI22_X1 U195 ( .A1(SH[4]), .A2(n211), .B1(n179), .B2(n205), .ZN(n210) );
  NAND2_X1 U196 ( .A1(SH[4]), .A2(n2), .ZN(n205) );
  NOR2_X1 U197 ( .A1(SH[5]), .A2(n202), .ZN(B[35]) );
  MUX2_X1 U198 ( .A(n180), .B(n212), .S(n97), .Z(n202) );
  OAI22_X1 U199 ( .A1(n213), .A2(n9), .B1(n181), .B2(n96), .ZN(B[34]) );
  OAI22_X1 U200 ( .A1(n214), .A2(n9), .B1(n186), .B2(n96), .ZN(B[33]) );
  OAI22_X1 U201 ( .A1(n215), .A2(n8), .B1(n187), .B2(n96), .ZN(B[32]) );
  OAI22_X1 U202 ( .A1(n216), .A2(n9), .B1(n27), .B2(n96), .ZN(B[31]) );
  OAI22_X1 U203 ( .A1(n218), .A2(n8), .B1(n188), .B2(n96), .ZN(B[30]) );
  NAND2_X1 U204 ( .A1(n219), .A2(n220), .ZN(B[2]) );
  AOI221_X1 U205 ( .B1(n141), .B2(n169), .C1(n143), .C2(n167), .A(n221), .ZN(
        n220) );
  OAI22_X1 U206 ( .A1(n222), .A2(n25), .B1(n181), .B2(n223), .ZN(n221) );
  AOI222_X1 U207 ( .A1(A[5]), .A2(n15), .B1(A[3]), .B2(n224), .C1(A[4]), .C2(
        n13), .ZN(n222) );
  AOI222_X1 U208 ( .A1(n163), .A2(n35), .B1(n139), .B2(n170), .C1(n145), .C2(
        n34), .ZN(n219) );
  OAI221_X1 U209 ( .B1(n6), .B2(n104), .C1(n3), .C2(n103), .A(n225), .ZN(n170)
         );
  AOI22_X1 U210 ( .A1(A[9]), .A2(n15), .B1(A[6]), .B2(n199), .ZN(n225) );
  OAI22_X1 U211 ( .A1(n227), .A2(n8), .B1(n189), .B2(n96), .ZN(B[29]) );
  OAI22_X1 U212 ( .A1(n228), .A2(n8), .B1(n190), .B2(n96), .ZN(B[28]) );
  OAI22_X1 U213 ( .A1(n229), .A2(n8), .B1(n26), .B2(n96), .ZN(B[27]) );
  OAI22_X1 U214 ( .A1(n231), .A2(n8), .B1(n191), .B2(n96), .ZN(B[26]) );
  OAI22_X1 U215 ( .A1(n136), .A2(n8), .B1(n148), .B2(n96), .ZN(B[25]) );
  AOI221_X1 U216 ( .B1(n91), .B2(n10), .C1(n85), .C2(n2), .A(n232), .ZN(n148)
         );
  OAI22_X1 U217 ( .A1(n58), .A2(n178), .B1(n5), .B2(n233), .ZN(n232) );
  AOI221_X1 U218 ( .B1(n234), .B2(n10), .C1(n235), .C2(n2), .A(n57), .ZN(n136)
         );
  AOI22_X1 U219 ( .A1(n237), .A2(n238), .B1(n196), .B2(n239), .ZN(n236) );
  OAI22_X1 U220 ( .A1(n149), .A2(n8), .B1(n156), .B2(n96), .ZN(B[24]) );
  AOI221_X1 U221 ( .B1(n60), .B2(n10), .C1(n62), .C2(n2), .A(n240), .ZN(n156)
         );
  OAI22_X1 U222 ( .A1(n58), .A2(n179), .B1(n5), .B2(n241), .ZN(n240) );
  AOI221_X1 U223 ( .B1(n242), .B2(n10), .C1(n243), .C2(n2), .A(n56), .ZN(n149)
         );
  AOI22_X1 U224 ( .A1(n237), .A2(n245), .B1(n196), .B2(n246), .ZN(n244) );
  OAI222_X1 U225 ( .A1(n204), .A2(n96), .B1(n176), .B2(n247), .C1(n164), .C2(
        n9), .ZN(B[23]) );
  AOI221_X1 U226 ( .B1(n248), .B2(n10), .C1(n249), .C2(n2), .A(n250), .ZN(n164) );
  OAI22_X1 U227 ( .A1(n58), .A2(n79), .B1(n5), .B2(n75), .ZN(n250) );
  AOI221_X1 U228 ( .B1(n80), .B2(n10), .C1(n77), .C2(n2), .A(n251), .ZN(n204)
         );
  OAI22_X1 U229 ( .A1(n58), .A2(n252), .B1(n5), .B2(n253), .ZN(n251) );
  OAI222_X1 U230 ( .A1(n207), .A2(n96), .B1(n177), .B2(n247), .C1(n171), .C2(
        n9), .ZN(B[22]) );
  AOI221_X1 U231 ( .B1(n255), .B2(n10), .C1(n256), .C2(n2), .A(n55), .ZN(n171)
         );
  AOI22_X1 U232 ( .A1(n237), .A2(n258), .B1(n196), .B2(n259), .ZN(n257) );
  AOI221_X1 U233 ( .B1(n70), .B2(n10), .C1(n260), .C2(n18), .A(n261), .ZN(n207) );
  OAI22_X1 U234 ( .A1(n58), .A2(n262), .B1(n5), .B2(n263), .ZN(n261) );
  OAI222_X1 U235 ( .A1(n209), .A2(n96), .B1(n178), .B2(n247), .C1(n175), .C2(
        n9), .ZN(B[21]) );
  AOI221_X1 U236 ( .B1(n235), .B2(n10), .C1(n142), .C2(n2), .A(n54), .ZN(n175)
         );
  AOI22_X1 U237 ( .A1(n237), .A2(n239), .B1(n196), .B2(n234), .ZN(n264) );
  AOI221_X1 U238 ( .B1(n85), .B2(n11), .C1(n238), .C2(n18), .A(n265), .ZN(n209) );
  OAI22_X1 U239 ( .A1(n58), .A2(n233), .B1(n5), .B2(n266), .ZN(n265) );
  OAI222_X1 U240 ( .A1(n211), .A2(n96), .B1(n179), .B2(n247), .C1(n185), .C2(
        n9), .ZN(B[20]) );
  AOI221_X1 U241 ( .B1(n243), .B2(n10), .C1(n153), .C2(n18), .A(n53), .ZN(n185) );
  AOI22_X1 U242 ( .A1(n237), .A2(n246), .B1(n196), .B2(n242), .ZN(n268) );
  NAND2_X1 U243 ( .A1(n145), .A2(n2), .ZN(n247) );
  AOI221_X1 U244 ( .B1(n62), .B2(n11), .C1(n245), .C2(n18), .A(n269), .ZN(n211) );
  OAI22_X1 U245 ( .A1(n58), .A2(n241), .B1(n5), .B2(n270), .ZN(n269) );
  NAND2_X1 U246 ( .A1(n271), .A2(n24), .ZN(B[1]) );
  OAI221_X1 U247 ( .B1(n25), .B2(n273), .C1(n223), .C2(n186), .A(n274), .ZN(
        n272) );
  AOI22_X1 U248 ( .A1(n147), .A2(n143), .B1(n140), .B2(n141), .ZN(n274) );
  OAI221_X1 U249 ( .B1(n6), .B2(n101), .C1(n3), .C2(n100), .A(n275), .ZN(n147)
         );
  AOI22_X1 U250 ( .A1(A[12]), .A2(n15), .B1(A[9]), .B2(n199), .ZN(n275) );
  AOI22_X1 U251 ( .A1(n15), .A2(A[4]), .B1(n13), .B2(A[3]), .ZN(n273) );
  AOI222_X1 U252 ( .A1(n163), .A2(n33), .B1(n139), .B2(n174), .C1(n145), .C2(
        n32), .ZN(n271) );
  OAI221_X1 U253 ( .B1(n6), .B2(n105), .C1(n3), .C2(n104), .A(n276), .ZN(n174)
         );
  AOI22_X1 U254 ( .A1(A[8]), .A2(n15), .B1(A[5]), .B2(n199), .ZN(n276) );
  OAI222_X1 U255 ( .A1(n212), .A2(n96), .B1(n95), .B2(n180), .C1(n201), .C2(n9), .ZN(B[19]) );
  AOI221_X1 U256 ( .B1(n249), .B2(n10), .C1(n160), .C2(n18), .A(n278), .ZN(
        n201) );
  OAI22_X1 U257 ( .A1(n58), .A2(n75), .B1(n5), .B2(n76), .ZN(n278) );
  OR2_X1 U258 ( .A1(n280), .A2(SH[3]), .ZN(n180) );
  AOI221_X1 U259 ( .B1(n77), .B2(n11), .C1(n281), .C2(n18), .A(n282), .ZN(n212) );
  OAI22_X1 U260 ( .A1(n58), .A2(n253), .B1(n5), .B2(n254), .ZN(n282) );
  OAI222_X1 U261 ( .A1(n213), .A2(n96), .B1(n181), .B2(n95), .C1(n226), .C2(n9), .ZN(B[18]) );
  AOI221_X1 U262 ( .B1(n256), .B2(n10), .C1(n168), .C2(n18), .A(n52), .ZN(n226) );
  AOI22_X1 U263 ( .A1(n237), .A2(n259), .B1(n196), .B2(n255), .ZN(n284) );
  AOI22_X1 U264 ( .A1(n73), .A2(n18), .B1(n72), .B2(n11), .ZN(n181) );
  AOI221_X1 U265 ( .B1(n260), .B2(n10), .C1(n258), .C2(n18), .A(n285), .ZN(
        n213) );
  OAI22_X1 U266 ( .A1(n58), .A2(n263), .B1(n5), .B2(n286), .ZN(n285) );
  OAI222_X1 U267 ( .A1(n214), .A2(n96), .B1(n186), .B2(n95), .C1(n277), .C2(n9), .ZN(B[17]) );
  AOI221_X1 U268 ( .B1(n142), .B2(n10), .C1(n144), .C2(n18), .A(n51), .ZN(n277) );
  AOI22_X1 U269 ( .A1(n237), .A2(n234), .B1(n196), .B2(n235), .ZN(n287) );
  AOI22_X1 U270 ( .A1(n88), .A2(n2), .B1(n90), .B2(n11), .ZN(n186) );
  AOI221_X1 U271 ( .B1(n238), .B2(n11), .C1(n239), .C2(n18), .A(n288), .ZN(
        n214) );
  OAI22_X1 U272 ( .A1(n58), .A2(n266), .B1(n5), .B2(n267), .ZN(n288) );
  OAI222_X1 U273 ( .A1(n215), .A2(n96), .B1(n187), .B2(n95), .C1(n289), .C2(n9), .ZN(B[16]) );
  OAI211_X1 U274 ( .C1(n216), .C2(n96), .A(n290), .B(n291), .ZN(B[15]) );
  AOI222_X1 U275 ( .A1(n139), .A2(n160), .B1(n141), .B2(n248), .C1(n143), .C2(
        n249), .ZN(n291) );
  AOI22_X1 U276 ( .A1(n145), .A2(n217), .B1(n146), .B2(n161), .ZN(n290) );
  OAI222_X1 U277 ( .A1(n252), .A2(n1), .B1(n5), .B2(n176), .C1(n253), .C2(n19), 
        .ZN(n217) );
  AOI221_X1 U278 ( .B1(n281), .B2(n11), .C1(n279), .C2(n2), .A(n292), .ZN(n216) );
  OAI22_X1 U279 ( .A1(n58), .A2(n254), .B1(n5), .B2(n283), .ZN(n292) );
  OAI211_X1 U280 ( .C1(n218), .C2(n96), .A(n293), .B(n294), .ZN(B[14]) );
  AOI222_X1 U281 ( .A1(n139), .A2(n168), .B1(n141), .B2(n255), .C1(n143), .C2(
        n256), .ZN(n294) );
  AOI22_X1 U282 ( .A1(n145), .A2(n31), .B1(n146), .B2(n169), .ZN(n293) );
  AOI222_X1 U283 ( .A1(n73), .A2(n10), .B1(n72), .B2(n196), .C1(n68), .C2(n2), 
        .ZN(n188) );
  AOI221_X1 U284 ( .B1(n258), .B2(n10), .C1(n259), .C2(n18), .A(n50), .ZN(n218) );
  AOI22_X1 U285 ( .A1(n237), .A2(n70), .B1(n196), .B2(n260), .ZN(n295) );
  OAI211_X1 U286 ( .C1(n227), .C2(n96), .A(n296), .B(n297), .ZN(B[13]) );
  AOI222_X1 U287 ( .A1(n139), .A2(n144), .B1(n141), .B2(n235), .C1(n143), .C2(
        n142), .ZN(n297) );
  OAI221_X1 U288 ( .B1(n6), .B2(n126), .C1(n3), .C2(n124), .A(n298), .ZN(n142)
         );
  AOI22_X1 U289 ( .A1(A[24]), .A2(n15), .B1(A[21]), .B2(n16), .ZN(n298) );
  OAI221_X1 U290 ( .B1(n6), .B2(n121), .C1(n3), .C2(n120), .A(n299), .ZN(n235)
         );
  AOI22_X1 U291 ( .A1(A[28]), .A2(n15), .B1(A[25]), .B2(n16), .ZN(n299) );
  OAI221_X1 U292 ( .B1(n6), .B2(n130), .C1(n3), .C2(n129), .A(n300), .ZN(n144)
         );
  AOI22_X1 U293 ( .A1(A[20]), .A2(n15), .B1(A[17]), .B2(n199), .ZN(n300) );
  AOI22_X1 U294 ( .A1(n145), .A2(n30), .B1(n146), .B2(n140), .ZN(n296) );
  OAI221_X1 U295 ( .B1(n6), .B2(n134), .C1(n3), .C2(n133), .A(n301), .ZN(n140)
         );
  AOI22_X1 U296 ( .A1(A[16]), .A2(n15), .B1(A[13]), .B2(n199), .ZN(n301) );
  AOI222_X1 U297 ( .A1(n88), .A2(n10), .B1(n90), .B2(n196), .C1(n91), .C2(n2), 
        .ZN(n189) );
  AOI221_X1 U298 ( .B1(n224), .B2(A[46]), .C1(n13), .C2(A[47]), .A(n92), .ZN(
        n266) );
  AOI22_X1 U299 ( .A1(A[48]), .A2(n15), .B1(A[45]), .B2(n16), .ZN(n302) );
  AOI222_X1 U300 ( .A1(n13), .A2(A[55]), .B1(n224), .B2(A[54]), .C1(n16), .C2(
        A[53]), .ZN(n178) );
  AOI221_X1 U301 ( .B1(n224), .B2(A[50]), .C1(n13), .C2(A[51]), .A(n89), .ZN(
        n233) );
  AOI22_X1 U302 ( .A1(A[52]), .A2(n15), .B1(A[49]), .B2(n16), .ZN(n303) );
  AOI221_X1 U303 ( .B1(n239), .B2(n11), .C1(n234), .C2(n2), .A(n304), .ZN(n227) );
  OAI22_X1 U304 ( .A1(n58), .A2(n267), .B1(n5), .B2(n87), .ZN(n304) );
  OAI221_X1 U305 ( .B1(n6), .B2(n108), .C1(n3), .C2(n107), .A(n305), .ZN(n238)
         );
  AOI22_X1 U306 ( .A1(A[40]), .A2(n15), .B1(A[37]), .B2(n16), .ZN(n305) );
  AOI221_X1 U307 ( .B1(n224), .B2(A[42]), .C1(n13), .C2(A[43]), .A(n86), .ZN(
        n267) );
  AOI22_X1 U308 ( .A1(A[44]), .A2(n15), .B1(A[41]), .B2(n16), .ZN(n306) );
  OAI221_X1 U309 ( .B1(n6), .B2(n117), .C1(n3), .C2(n116), .A(n307), .ZN(n234)
         );
  AOI22_X1 U310 ( .A1(A[32]), .A2(n15), .B1(A[29]), .B2(n16), .ZN(n307) );
  OAI221_X1 U311 ( .B1(n6), .B2(n112), .C1(n12), .C2(n111), .A(n308), .ZN(n239) );
  AOI22_X1 U312 ( .A1(A[36]), .A2(n15), .B1(A[33]), .B2(n16), .ZN(n308) );
  OAI211_X1 U313 ( .C1(n228), .C2(n96), .A(n309), .B(n310), .ZN(B[12]) );
  AOI222_X1 U314 ( .A1(n139), .A2(n154), .B1(n141), .B2(n243), .C1(n143), .C2(
        n153), .ZN(n310) );
  AOI22_X1 U315 ( .A1(n145), .A2(n29), .B1(n146), .B2(n152), .ZN(n309) );
  AOI222_X1 U316 ( .A1(n64), .A2(n10), .B1(n66), .B2(n196), .C1(n60), .C2(n2), 
        .ZN(n190) );
  AOI221_X1 U317 ( .B1(n246), .B2(n11), .C1(n242), .C2(n2), .A(n49), .ZN(n228)
         );
  AOI22_X1 U318 ( .A1(n237), .A2(n62), .B1(n196), .B2(n245), .ZN(n311) );
  OAI211_X1 U319 ( .C1(n229), .C2(n96), .A(n313), .B(n314), .ZN(B[11]) );
  AOI222_X1 U320 ( .A1(n139), .A2(n161), .B1(n141), .B2(n249), .C1(n143), .C2(
        n160), .ZN(n314) );
  OAI221_X1 U321 ( .B1(n6), .B2(n128), .C1(n12), .C2(n127), .A(n315), .ZN(n160) );
  AOI22_X1 U322 ( .A1(n15), .A2(A[22]), .B1(A[19]), .B2(n16), .ZN(n315) );
  OAI221_X1 U323 ( .B1(n6), .B2(n123), .C1(n12), .C2(n122), .A(n316), .ZN(n249) );
  AOI22_X1 U324 ( .A1(A[26]), .A2(n15), .B1(n199), .B2(A[23]), .ZN(n316) );
  OAI221_X1 U325 ( .B1(n6), .B2(n132), .C1(n12), .C2(n131), .A(n317), .ZN(n161) );
  AOI22_X1 U326 ( .A1(A[18]), .A2(n15), .B1(A[15]), .B2(n16), .ZN(n317) );
  AOI22_X1 U327 ( .A1(n145), .A2(n230), .B1(n146), .B2(n159), .ZN(n313) );
  OAI221_X1 U328 ( .B1(n6), .B2(n99), .C1(n12), .C2(n135), .A(n318), .ZN(n159)
         );
  AOI22_X1 U329 ( .A1(A[14]), .A2(n15), .B1(A[11]), .B2(n16), .ZN(n318) );
  OAI222_X1 U330 ( .A1(n254), .A2(n19), .B1(n253), .B2(n1), .C1(n280), .C2(n94), .ZN(n230) );
  MUX2_X1 U331 ( .A(n176), .B(n252), .S(n59), .Z(n280) );
  AOI221_X1 U332 ( .B1(n224), .B2(A[52]), .C1(n13), .C2(A[53]), .A(n83), .ZN(
        n252) );
  AOI22_X1 U333 ( .A1(A[54]), .A2(n15), .B1(A[51]), .B2(n16), .ZN(n319) );
  NAND2_X1 U334 ( .A1(A[55]), .A2(n199), .ZN(n176) );
  AOI221_X1 U335 ( .B1(n224), .B2(A[48]), .C1(n13), .C2(A[49]), .A(n82), .ZN(
        n253) );
  AOI22_X1 U336 ( .A1(A[50]), .A2(n15), .B1(A[47]), .B2(n16), .ZN(n320) );
  AOI221_X1 U337 ( .B1(n224), .B2(A[44]), .C1(n13), .C2(A[45]), .A(n81), .ZN(
        n254) );
  AOI22_X1 U338 ( .A1(A[46]), .A2(n15), .B1(A[43]), .B2(n16), .ZN(n321) );
  AOI221_X1 U339 ( .B1(n279), .B2(n11), .C1(n248), .C2(n2), .A(n322), .ZN(n229) );
  OAI22_X1 U340 ( .A1(n58), .A2(n283), .B1(n5), .B2(n79), .ZN(n322) );
  OAI221_X1 U341 ( .B1(n6), .B2(n110), .C1(n12), .C2(n109), .A(n323), .ZN(n281) );
  AOI22_X1 U342 ( .A1(A[38]), .A2(n198), .B1(A[35]), .B2(n16), .ZN(n323) );
  AOI221_X1 U343 ( .B1(n224), .B2(A[40]), .C1(n13), .C2(A[41]), .A(n78), .ZN(
        n283) );
  AOI22_X1 U344 ( .A1(A[42]), .A2(n15), .B1(A[39]), .B2(n16), .ZN(n324) );
  OAI221_X1 U345 ( .B1(n6), .B2(n119), .C1(n12), .C2(n118), .A(n325), .ZN(n248) );
  AOI22_X1 U346 ( .A1(A[30]), .A2(n15), .B1(A[27]), .B2(n16), .ZN(n325) );
  OAI221_X1 U347 ( .B1(n6), .B2(n115), .C1(n12), .C2(n113), .A(n326), .ZN(n279) );
  AOI22_X1 U348 ( .A1(A[34]), .A2(n198), .B1(A[31]), .B2(n16), .ZN(n326) );
  OAI211_X1 U349 ( .C1(n231), .C2(n96), .A(n327), .B(n328), .ZN(B[10]) );
  AOI222_X1 U350 ( .A1(n139), .A2(n169), .B1(n141), .B2(n256), .C1(n143), .C2(
        n168), .ZN(n328) );
  OAI221_X1 U351 ( .B1(n6), .B2(n129), .C1(n12), .C2(n128), .A(n329), .ZN(n168) );
  AOI22_X1 U352 ( .A1(A[21]), .A2(n198), .B1(A[18]), .B2(n16), .ZN(n329) );
  OAI221_X1 U353 ( .B1(n6), .B2(n124), .C1(n12), .C2(n123), .A(n330), .ZN(n256) );
  AOI22_X1 U354 ( .A1(A[25]), .A2(n198), .B1(n199), .B2(A[22]), .ZN(n330) );
  OAI221_X1 U355 ( .B1(n6), .B2(n133), .C1(n12), .C2(n132), .A(n331), .ZN(n169) );
  AOI22_X1 U356 ( .A1(A[17]), .A2(n198), .B1(A[14]), .B2(n16), .ZN(n331) );
  AOI22_X1 U357 ( .A1(n145), .A2(n28), .B1(n146), .B2(n167), .ZN(n327) );
  OAI221_X1 U358 ( .B1(n7), .B2(n100), .C1(n12), .C2(n99), .A(n332), .ZN(n167)
         );
  AOI22_X1 U359 ( .A1(A[13]), .A2(n198), .B1(A[10]), .B2(n16), .ZN(n332) );
  AOI221_X1 U360 ( .B1(n68), .B2(n11), .C1(n70), .C2(n2), .A(n333), .ZN(n191)
         );
  OAI22_X1 U361 ( .A1(n58), .A2(n177), .B1(n5), .B2(n262), .ZN(n333) );
  AOI221_X1 U362 ( .B1(n224), .B2(A[51]), .C1(n13), .C2(A[52]), .A(n74), .ZN(
        n262) );
  AOI22_X1 U363 ( .A1(A[53]), .A2(n15), .B1(A[50]), .B2(n16), .ZN(n334) );
  AOI22_X1 U364 ( .A1(n16), .A2(A[54]), .B1(n224), .B2(A[55]), .ZN(n177) );
  AOI221_X1 U365 ( .B1(n224), .B2(A[43]), .C1(n13), .C2(A[44]), .A(n71), .ZN(
        n286) );
  AOI22_X1 U366 ( .A1(A[45]), .A2(n15), .B1(A[42]), .B2(n16), .ZN(n335) );
  AOI221_X1 U367 ( .B1(n224), .B2(A[47]), .C1(n13), .C2(A[48]), .A(n69), .ZN(
        n263) );
  AOI22_X1 U368 ( .A1(A[49]), .A2(n15), .B1(A[46]), .B2(n16), .ZN(n336) );
  AOI221_X1 U369 ( .B1(n259), .B2(n11), .C1(n255), .C2(n2), .A(n48), .ZN(n231)
         );
  AOI22_X1 U370 ( .A1(n237), .A2(n260), .B1(n196), .B2(n258), .ZN(n337) );
  OAI221_X1 U371 ( .B1(n7), .B2(n111), .C1(n12), .C2(n110), .A(n338), .ZN(n258) );
  AOI22_X1 U372 ( .A1(A[37]), .A2(n198), .B1(A[34]), .B2(n16), .ZN(n338) );
  OAI221_X1 U373 ( .B1(n7), .B2(n107), .C1(n12), .C2(n106), .A(n339), .ZN(n260) );
  AOI22_X1 U374 ( .A1(A[41]), .A2(n15), .B1(A[38]), .B2(n16), .ZN(n339) );
  OAI221_X1 U375 ( .B1(n7), .B2(n120), .C1(n12), .C2(n119), .A(n340), .ZN(n255) );
  AOI22_X1 U376 ( .A1(A[29]), .A2(n15), .B1(A[26]), .B2(n16), .ZN(n340) );
  OAI221_X1 U377 ( .B1(n7), .B2(n116), .C1(n12), .C2(n115), .A(n341), .ZN(n259) );
  AOI22_X1 U378 ( .A1(A[33]), .A2(n15), .B1(A[30]), .B2(n16), .ZN(n341) );
  NAND2_X1 U379 ( .A1(n342), .A2(n23), .ZN(B[0]) );
  OAI211_X1 U380 ( .C1(n223), .C2(n187), .A(n344), .B(n345), .ZN(n343) );
  NAND3_X1 U381 ( .A1(A[3]), .A2(n15), .A3(n146), .ZN(n345) );
  AOI22_X1 U382 ( .A1(n155), .A2(n143), .B1(n152), .B2(n141), .ZN(n344) );
  OAI221_X1 U383 ( .B1(n7), .B2(n135), .C1(n12), .C2(n134), .A(n346), .ZN(n152) );
  AOI22_X1 U384 ( .A1(A[15]), .A2(n198), .B1(A[12]), .B2(n16), .ZN(n346) );
  OAI221_X1 U385 ( .B1(n7), .B2(n102), .C1(n12), .C2(n101), .A(n347), .ZN(n155) );
  AOI22_X1 U386 ( .A1(A[11]), .A2(n198), .B1(A[8]), .B2(n16), .ZN(n347) );
  AOI22_X1 U387 ( .A1(n64), .A2(n18), .B1(n66), .B2(n11), .ZN(n187) );
  AOI221_X1 U388 ( .B1(n224), .B2(A[53]), .C1(n13), .C2(A[54]), .A(n67), .ZN(
        n179) );
  AOI22_X1 U389 ( .A1(A[55]), .A2(n15), .B1(A[52]), .B2(n16), .ZN(n348) );
  AOI221_X1 U390 ( .B1(n224), .B2(A[49]), .C1(n13), .C2(A[50]), .A(n65), .ZN(
        n241) );
  AOI22_X1 U391 ( .A1(A[51]), .A2(n15), .B1(A[48]), .B2(n16), .ZN(n349) );
  NAND2_X1 U392 ( .A1(SH[4]), .A2(SH[5]), .ZN(n223) );
  AOI222_X1 U393 ( .A1(n163), .A2(n20), .B1(n139), .B2(n184), .C1(n145), .C2(
        n22), .ZN(n342) );
  AOI221_X1 U394 ( .B1(n245), .B2(n11), .C1(n246), .C2(n18), .A(n350), .ZN(
        n215) );
  OAI22_X1 U395 ( .A1(n58), .A2(n270), .B1(n5), .B2(n312), .ZN(n350) );
  AOI221_X1 U396 ( .B1(n224), .B2(A[41]), .C1(n13), .C2(A[42]), .A(n63), .ZN(
        n312) );
  AOI22_X1 U397 ( .A1(A[43]), .A2(n198), .B1(A[40]), .B2(n199), .ZN(n351) );
  AOI221_X1 U398 ( .B1(n224), .B2(A[45]), .C1(n13), .C2(A[46]), .A(n61), .ZN(
        n270) );
  AOI22_X1 U399 ( .A1(A[47]), .A2(n198), .B1(A[44]), .B2(n199), .ZN(n352) );
  OAI221_X1 U400 ( .B1(n7), .B2(n113), .C1(n12), .C2(n112), .A(n353), .ZN(n246) );
  AOI22_X1 U401 ( .A1(A[35]), .A2(n15), .B1(A[32]), .B2(n16), .ZN(n353) );
  OAI221_X1 U402 ( .B1(n7), .B2(n109), .C1(n12), .C2(n108), .A(n354), .ZN(n245) );
  AOI22_X1 U403 ( .A1(A[39]), .A2(n15), .B1(A[36]), .B2(n16), .ZN(n354) );
  OAI221_X1 U404 ( .B1(n7), .B2(n114), .C1(n12), .C2(n105), .A(n355), .ZN(n184) );
  AOI22_X1 U405 ( .A1(A[7]), .A2(n15), .B1(A[4]), .B2(n16), .ZN(n355) );
  AOI221_X1 U406 ( .B1(n242), .B2(n237), .C1(n243), .C2(n196), .A(n21), .ZN(
        n289) );
  AOI22_X1 U407 ( .A1(n10), .A2(n153), .B1(n2), .B2(n154), .ZN(n356) );
  OAI221_X1 U408 ( .B1(n7), .B2(n131), .C1(n3), .C2(n130), .A(n357), .ZN(n154)
         );
  AOI22_X1 U409 ( .A1(A[19]), .A2(n15), .B1(A[16]), .B2(n16), .ZN(n357) );
  OAI221_X1 U410 ( .B1(n7), .B2(n127), .C1(n126), .C2(n3), .A(n358), .ZN(n153)
         );
  AOI22_X1 U411 ( .A1(n15), .A2(A[23]), .B1(A[20]), .B2(n16), .ZN(n358) );
  OAI221_X1 U412 ( .B1(n6), .B2(n122), .C1(n3), .C2(n121), .A(n359), .ZN(n243)
         );
  AOI22_X1 U413 ( .A1(A[27]), .A2(n15), .B1(n16), .B2(A[24]), .ZN(n359) );
  OAI221_X1 U414 ( .B1(n6), .B2(n118), .C1(n12), .C2(n117), .A(n360), .ZN(n242) );
  AOI22_X1 U415 ( .A1(A[31]), .A2(n15), .B1(A[28]), .B2(n16), .ZN(n360) );
  NOR2_X1 U416 ( .A1(SH[0]), .A2(SH[1]), .ZN(n199) );
  AND2_X1 U417 ( .A1(SH[1]), .A2(SH[0]), .ZN(n198) );
  NOR2_X1 U418 ( .A1(n97), .A2(SH[5]), .ZN(n163) );
endmodule


module fpu_DW01_sub_13 ( A, B, CI, DIFF, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
  wire   [10:1] carry;

  FA_X1 U2_10 ( .A(A[10]), .B(n10), .CI(carry[10]), .S(DIFF[10]) );
  FA_X1 U2_9 ( .A(A[9]), .B(n1), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9]) );
  FA_X1 U2_8 ( .A(A[8]), .B(n2), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FA_X1 U2_7 ( .A(A[7]), .B(n3), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FA_X1 U2_6 ( .A(A[6]), .B(n4), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA_X1 U2_5 ( .A(A[5]), .B(n5), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n6), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_3 ( .A(A[3]), .B(n7), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA_X1 U2_2 ( .A(A[2]), .B(n8), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA_X1 U2_1 ( .A(A[1]), .B(n9), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  FA_X1 U2_0 ( .A(A[0]), .B(n11), .CI(n12), .CO(carry[1]), .S(DIFF[0]) );
  INV_X4 U1 ( .A(B[9]), .ZN(n1) );
  INV_X4 U2 ( .A(B[8]), .ZN(n2) );
  INV_X4 U3 ( .A(B[7]), .ZN(n3) );
  INV_X4 U4 ( .A(B[6]), .ZN(n4) );
  INV_X4 U5 ( .A(B[5]), .ZN(n5) );
  INV_X4 U6 ( .A(B[4]), .ZN(n6) );
  INV_X4 U7 ( .A(B[3]), .ZN(n7) );
  INV_X4 U8 ( .A(B[2]), .ZN(n8) );
  INV_X4 U9 ( .A(B[1]), .ZN(n9) );
  INV_X4 U10 ( .A(B[10]), .ZN(n10) );
  INV_X4 U11 ( .A(B[0]), .ZN(n11) );
  INV_X4 U12 ( .A(CI), .ZN(n12) );
endmodule


module fpu_DW01_sub_14 ( A, B, CI, DIFF, CO );
  input [105:0] A;
  input [105:0] B;
  output [105:0] DIFF;
  input CI;
  output CO;
  wire   n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n97, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171;

  XOR2_X2 U1 ( .A(n116), .B(n95), .Z(DIFF[103]) );
  XOR2_X2 U2 ( .A(n115), .B(n46), .Z(DIFF[104]) );
  XOR2_X2 U3 ( .A(n114), .B(n97), .Z(DIFF[105]) );
  XOR2_X2 U4 ( .A(n140), .B(n48), .Z(DIFF[79]) );
  XOR2_X2 U5 ( .A(n139), .B(n85), .Z(DIFF[80]) );
  AND2_X4 U6 ( .A1(n165), .A2(n39), .ZN(n6) );
  AND2_X4 U7 ( .A1(n167), .A2(n40), .ZN(n7) );
  AND2_X4 U8 ( .A1(n169), .A2(n41), .ZN(n8) );
  AND2_X4 U9 ( .A1(n120), .A2(n42), .ZN(n9) );
  AND2_X4 U10 ( .A1(n125), .A2(n78), .ZN(n10) );
  AND2_X4 U11 ( .A1(n127), .A2(n79), .ZN(n11) );
  AND2_X4 U12 ( .A1(n129), .A2(n80), .ZN(n12) );
  AND2_X4 U13 ( .A1(n131), .A2(n81), .ZN(n13) );
  AND2_X4 U14 ( .A1(n133), .A2(n82), .ZN(n14) );
  AND2_X4 U15 ( .A1(n135), .A2(n83), .ZN(n15) );
  AND2_X4 U16 ( .A1(n137), .A2(n84), .ZN(n16) );
  AND2_X4 U17 ( .A1(n151), .A2(n91), .ZN(n17) );
  AND2_X4 U18 ( .A1(n153), .A2(n92), .ZN(n18) );
  AND2_X4 U19 ( .A1(n155), .A2(n93), .ZN(n19) );
  AND2_X4 U20 ( .A1(n157), .A2(n94), .ZN(n20) );
  AND2_X4 U21 ( .A1(n161), .A2(n37), .ZN(n21) );
  AND2_X4 U22 ( .A1(n163), .A2(n38), .ZN(n22) );
  AND2_X4 U23 ( .A1(n139), .A2(n85), .ZN(n23) );
  XOR2_X2 U24 ( .A(n122), .B(n47), .Z(DIFF[97]) );
  XOR2_X2 U25 ( .A(n123), .B(n77), .Z(DIFF[96]) );
  XOR2_X2 U26 ( .A(n121), .B(n76), .Z(DIFF[98]) );
  XOR2_X2 U27 ( .A(n142), .B(n49), .Z(DIFF[77]) );
  XOR2_X2 U28 ( .A(n141), .B(n86), .Z(DIFF[78]) );
  XOR2_X2 U29 ( .A(n147), .B(n89), .Z(DIFF[72]) );
  XOR2_X2 U30 ( .A(n143), .B(n87), .Z(DIFF[76]) );
  XOR2_X2 U31 ( .A(n149), .B(n90), .Z(DIFF[70]) );
  XOR2_X2 U32 ( .A(n148), .B(n52), .Z(DIFF[71]) );
  XOR2_X2 U33 ( .A(n146), .B(n51), .Z(DIFF[73]) );
  XOR2_X2 U34 ( .A(n145), .B(n88), .Z(DIFF[74]) );
  XOR2_X2 U35 ( .A(n144), .B(n50), .Z(DIFF[75]) );
  AND2_X4 U36 ( .A1(n160), .A2(n21), .ZN(n36) );
  AND2_X4 U37 ( .A1(n162), .A2(n22), .ZN(n37) );
  AND2_X4 U38 ( .A1(n164), .A2(n6), .ZN(n38) );
  AND2_X4 U39 ( .A1(n166), .A2(n7), .ZN(n39) );
  AND2_X4 U40 ( .A1(n168), .A2(n8), .ZN(n40) );
  AND2_X4 U41 ( .A1(n170), .A2(n171), .ZN(n41) );
  AND2_X4 U42 ( .A1(n121), .A2(n76), .ZN(n42) );
  AND2_X4 U43 ( .A1(n119), .A2(n9), .ZN(n43) );
  AND2_X4 U44 ( .A1(n159), .A2(n36), .ZN(n44) );
  AND2_X4 U45 ( .A1(n118), .A2(n43), .ZN(n45) );
  AND2_X4 U46 ( .A1(n116), .A2(n95), .ZN(n46) );
  AND2_X4 U47 ( .A1(n123), .A2(n77), .ZN(n47) );
  AND2_X4 U48 ( .A1(n141), .A2(n86), .ZN(n48) );
  AND2_X4 U49 ( .A1(n143), .A2(n87), .ZN(n49) );
  AND2_X4 U50 ( .A1(n145), .A2(n88), .ZN(n50) );
  AND2_X4 U51 ( .A1(n147), .A2(n89), .ZN(n51) );
  AND2_X4 U52 ( .A1(n149), .A2(n90), .ZN(n52) );
  XOR2_X2 U53 ( .A(n137), .B(n84), .Z(DIFF[82]) );
  XOR2_X2 U54 ( .A(n136), .B(n16), .Z(DIFF[83]) );
  XOR2_X2 U55 ( .A(n131), .B(n81), .Z(DIFF[88]) );
  XOR2_X2 U56 ( .A(n129), .B(n80), .Z(DIFF[90]) );
  XOR2_X2 U57 ( .A(n138), .B(n23), .Z(DIFF[81]) );
  XOR2_X2 U58 ( .A(n135), .B(n83), .Z(DIFF[84]) );
  XOR2_X2 U59 ( .A(n134), .B(n15), .Z(DIFF[85]) );
  XOR2_X2 U60 ( .A(n133), .B(n82), .Z(DIFF[86]) );
  XOR2_X2 U61 ( .A(n132), .B(n14), .Z(DIFF[87]) );
  XOR2_X2 U62 ( .A(n130), .B(n13), .Z(DIFF[89]) );
  XOR2_X2 U63 ( .A(n128), .B(n12), .Z(DIFF[91]) );
  XOR2_X2 U64 ( .A(n127), .B(n79), .Z(DIFF[92]) );
  XOR2_X2 U65 ( .A(n126), .B(n11), .Z(DIFF[93]) );
  XOR2_X2 U66 ( .A(n125), .B(n78), .Z(DIFF[94]) );
  XOR2_X2 U67 ( .A(n124), .B(n10), .Z(DIFF[95]) );
  XOR2_X2 U68 ( .A(n155), .B(n93), .Z(DIFF[64]) );
  XOR2_X2 U69 ( .A(n154), .B(n19), .Z(DIFF[65]) );
  XOR2_X2 U70 ( .A(n153), .B(n92), .Z(DIFF[66]) );
  XOR2_X2 U71 ( .A(n152), .B(n18), .Z(DIFF[67]) );
  XOR2_X2 U72 ( .A(n157), .B(n94), .Z(DIFF[62]) );
  XOR2_X2 U73 ( .A(n156), .B(n20), .Z(DIFF[63]) );
  XOR2_X2 U74 ( .A(n151), .B(n91), .Z(DIFF[68]) );
  XOR2_X2 U75 ( .A(n150), .B(n17), .Z(DIFF[69]) );
  AND2_X4 U76 ( .A1(n122), .A2(n47), .ZN(n76) );
  AND2_X4 U77 ( .A1(n124), .A2(n10), .ZN(n77) );
  AND2_X4 U78 ( .A1(n126), .A2(n11), .ZN(n78) );
  AND2_X4 U79 ( .A1(n128), .A2(n12), .ZN(n79) );
  AND2_X4 U80 ( .A1(n130), .A2(n13), .ZN(n80) );
  AND2_X4 U81 ( .A1(n132), .A2(n14), .ZN(n81) );
  AND2_X4 U82 ( .A1(n134), .A2(n15), .ZN(n82) );
  AND2_X4 U83 ( .A1(n136), .A2(n16), .ZN(n83) );
  AND2_X4 U84 ( .A1(n138), .A2(n23), .ZN(n84) );
  AND2_X4 U85 ( .A1(n140), .A2(n48), .ZN(n85) );
  AND2_X4 U86 ( .A1(n142), .A2(n49), .ZN(n86) );
  AND2_X4 U87 ( .A1(n144), .A2(n50), .ZN(n87) );
  AND2_X4 U88 ( .A1(n146), .A2(n51), .ZN(n88) );
  AND2_X4 U89 ( .A1(n148), .A2(n52), .ZN(n89) );
  AND2_X4 U90 ( .A1(n150), .A2(n17), .ZN(n90) );
  AND2_X4 U91 ( .A1(n152), .A2(n18), .ZN(n91) );
  AND2_X4 U92 ( .A1(n154), .A2(n19), .ZN(n92) );
  AND2_X4 U93 ( .A1(n156), .A2(n20), .ZN(n93) );
  AND2_X4 U94 ( .A1(n158), .A2(n44), .ZN(n94) );
  AND2_X4 U95 ( .A1(n117), .A2(n45), .ZN(n95) );
  XOR2_X2 U96 ( .A(n120), .B(n42), .Z(DIFF[99]) );
  AND2_X4 U97 ( .A1(n115), .A2(n46), .ZN(n97) );
  XOR2_X2 U98 ( .A(n119), .B(n9), .Z(DIFF[100]) );
  XOR2_X2 U99 ( .A(n118), .B(n43), .Z(DIFF[101]) );
  XOR2_X2 U100 ( .A(n117), .B(n45), .Z(DIFF[102]) );
  XOR2_X2 U101 ( .A(n170), .B(n171), .Z(DIFF[49]) );
  XOR2_X2 U102 ( .A(n167), .B(n40), .Z(DIFF[52]) );
  XOR2_X2 U103 ( .A(n166), .B(n7), .Z(DIFF[53]) );
  XOR2_X2 U104 ( .A(n165), .B(n39), .Z(DIFF[54]) );
  XOR2_X2 U105 ( .A(n163), .B(n38), .Z(DIFF[56]) );
  XOR2_X2 U106 ( .A(n169), .B(n41), .Z(DIFF[50]) );
  XOR2_X2 U107 ( .A(n168), .B(n8), .Z(DIFF[51]) );
  XOR2_X2 U108 ( .A(n164), .B(n6), .Z(DIFF[55]) );
  XOR2_X2 U109 ( .A(n162), .B(n22), .Z(DIFF[57]) );
  XOR2_X2 U110 ( .A(n161), .B(n37), .Z(DIFF[58]) );
  XOR2_X2 U111 ( .A(n160), .B(n21), .Z(DIFF[59]) );
  XOR2_X2 U112 ( .A(n159), .B(n36), .Z(DIFF[60]) );
  XOR2_X2 U113 ( .A(n158), .B(n44), .Z(DIFF[61]) );
  INV_X4 U114 ( .A(B[105]), .ZN(n114) );
  INV_X4 U115 ( .A(B[104]), .ZN(n115) );
  INV_X4 U116 ( .A(B[103]), .ZN(n116) );
  INV_X4 U117 ( .A(B[102]), .ZN(n117) );
  INV_X4 U118 ( .A(B[101]), .ZN(n118) );
  INV_X4 U119 ( .A(B[100]), .ZN(n119) );
  INV_X4 U120 ( .A(B[99]), .ZN(n120) );
  INV_X4 U121 ( .A(B[98]), .ZN(n121) );
  INV_X4 U122 ( .A(B[97]), .ZN(n122) );
  INV_X4 U123 ( .A(B[96]), .ZN(n123) );
  INV_X4 U124 ( .A(B[95]), .ZN(n124) );
  INV_X4 U125 ( .A(B[94]), .ZN(n125) );
  INV_X4 U126 ( .A(B[93]), .ZN(n126) );
  INV_X4 U127 ( .A(B[92]), .ZN(n127) );
  INV_X4 U128 ( .A(B[91]), .ZN(n128) );
  INV_X4 U129 ( .A(B[90]), .ZN(n129) );
  INV_X4 U130 ( .A(B[89]), .ZN(n130) );
  INV_X4 U131 ( .A(B[88]), .ZN(n131) );
  INV_X4 U132 ( .A(B[87]), .ZN(n132) );
  INV_X4 U133 ( .A(B[86]), .ZN(n133) );
  INV_X4 U134 ( .A(B[85]), .ZN(n134) );
  INV_X4 U135 ( .A(B[84]), .ZN(n135) );
  INV_X4 U136 ( .A(B[83]), .ZN(n136) );
  INV_X4 U137 ( .A(B[82]), .ZN(n137) );
  INV_X4 U138 ( .A(B[81]), .ZN(n138) );
  INV_X4 U139 ( .A(B[80]), .ZN(n139) );
  INV_X4 U140 ( .A(B[79]), .ZN(n140) );
  INV_X4 U141 ( .A(B[78]), .ZN(n141) );
  INV_X4 U142 ( .A(B[77]), .ZN(n142) );
  INV_X4 U143 ( .A(B[76]), .ZN(n143) );
  INV_X4 U144 ( .A(B[75]), .ZN(n144) );
  INV_X4 U145 ( .A(B[74]), .ZN(n145) );
  INV_X4 U146 ( .A(B[73]), .ZN(n146) );
  INV_X4 U147 ( .A(B[72]), .ZN(n147) );
  INV_X4 U148 ( .A(B[71]), .ZN(n148) );
  INV_X4 U149 ( .A(B[70]), .ZN(n149) );
  INV_X4 U150 ( .A(B[69]), .ZN(n150) );
  INV_X4 U151 ( .A(B[68]), .ZN(n151) );
  INV_X4 U152 ( .A(B[67]), .ZN(n152) );
  INV_X4 U153 ( .A(B[66]), .ZN(n153) );
  INV_X4 U154 ( .A(B[65]), .ZN(n154) );
  INV_X4 U155 ( .A(B[64]), .ZN(n155) );
  INV_X4 U156 ( .A(B[63]), .ZN(n156) );
  INV_X4 U157 ( .A(B[62]), .ZN(n157) );
  INV_X4 U158 ( .A(B[61]), .ZN(n158) );
  INV_X4 U159 ( .A(B[60]), .ZN(n159) );
  INV_X4 U160 ( .A(B[59]), .ZN(n160) );
  INV_X4 U161 ( .A(B[58]), .ZN(n161) );
  INV_X4 U162 ( .A(B[57]), .ZN(n162) );
  INV_X4 U163 ( .A(B[56]), .ZN(n163) );
  INV_X4 U164 ( .A(B[55]), .ZN(n164) );
  INV_X4 U165 ( .A(B[54]), .ZN(n165) );
  INV_X4 U166 ( .A(B[53]), .ZN(n166) );
  INV_X4 U167 ( .A(B[52]), .ZN(n167) );
  INV_X4 U168 ( .A(B[51]), .ZN(n168) );
  INV_X4 U169 ( .A(B[50]), .ZN(n169) );
  INV_X4 U170 ( .A(B[49]), .ZN(n170) );
  INV_X4 U171 ( .A(B[48]), .ZN(n171) );
endmodule


module fpu_DW01_sub_15 ( A, B, CI, DIFF, CO );
  input [53:0] A;
  input [53:0] B;
  output [53:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n1, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  AND2_X4 U1 ( .A1(n106), .A2(n10), .ZN(n1) );
  XOR2_X2 U2 ( .A(n113), .B(n47), .Z(DIFF[44]) );
  XOR2_X2 U3 ( .A(n120), .B(n29), .Z(DIFF[37]) );
  XOR2_X2 U4 ( .A(n119), .B(n50), .Z(DIFF[38]) );
  XOR2_X2 U5 ( .A(n118), .B(n34), .Z(DIFF[39]) );
  XOR2_X2 U6 ( .A(n117), .B(n49), .Z(DIFF[40]) );
  XOR2_X2 U7 ( .A(n116), .B(n33), .Z(DIFF[41]) );
  XOR2_X2 U8 ( .A(n115), .B(n48), .Z(DIFF[42]) );
  XOR2_X2 U9 ( .A(n114), .B(n32), .Z(DIFF[43]) );
  AND2_X4 U10 ( .A1(n107), .A2(n44), .ZN(n10) );
  AND2_X4 U11 ( .A1(n143), .A2(n62), .ZN(n11) );
  AND2_X4 U12 ( .A1(n145), .A2(n63), .ZN(n12) );
  AND2_X4 U13 ( .A1(n147), .A2(n64), .ZN(n13) );
  AND2_X4 U14 ( .A1(n149), .A2(n65), .ZN(n14) );
  AND2_X4 U15 ( .A1(n151), .A2(n66), .ZN(n15) );
  AND2_X4 U16 ( .A1(n111), .A2(n46), .ZN(n16) );
  AND2_X4 U17 ( .A1(n123), .A2(n52), .ZN(n17) );
  AND2_X4 U18 ( .A1(n125), .A2(n53), .ZN(n18) );
  AND2_X4 U19 ( .A1(n127), .A2(n54), .ZN(n19) );
  AND2_X4 U20 ( .A1(n129), .A2(n55), .ZN(n20) );
  AND2_X4 U21 ( .A1(n131), .A2(n56), .ZN(n21) );
  AND2_X4 U22 ( .A1(n133), .A2(n57), .ZN(n22) );
  AND2_X4 U23 ( .A1(n135), .A2(n58), .ZN(n23) );
  AND2_X4 U24 ( .A1(n137), .A2(n59), .ZN(n24) );
  AND2_X4 U25 ( .A1(n139), .A2(n60), .ZN(n25) );
  AND2_X4 U26 ( .A1(n141), .A2(n61), .ZN(n26) );
  AND2_X4 U27 ( .A1(n109), .A2(n45), .ZN(n27) );
  AND2_X4 U28 ( .A1(n153), .A2(n67), .ZN(n28) );
  AND2_X4 U29 ( .A1(n121), .A2(n51), .ZN(n29) );
  AND2_X4 U30 ( .A1(n155), .A2(n68), .ZN(n30) );
  AND2_X4 U31 ( .A1(n113), .A2(n47), .ZN(n31) );
  AND2_X4 U32 ( .A1(n115), .A2(n48), .ZN(n32) );
  AND2_X4 U33 ( .A1(n117), .A2(n49), .ZN(n33) );
  AND2_X4 U34 ( .A1(n119), .A2(n50), .ZN(n34) );
  XOR2_X2 U35 ( .A(n107), .B(n44), .Z(DIFF[50]) );
  XOR2_X2 U36 ( .A(n112), .B(n31), .Z(DIFF[45]) );
  XOR2_X2 U37 ( .A(n109), .B(n45), .Z(DIFF[48]) );
  XOR2_X2 U38 ( .A(n156), .B(n157), .Z(DIFF[1]) );
  XOR2_X2 U39 ( .A(n155), .B(n68), .Z(DIFF[2]) );
  XOR2_X2 U40 ( .A(n154), .B(n30), .Z(DIFF[3]) );
  XOR2_X2 U41 ( .A(n153), .B(n67), .Z(DIFF[4]) );
  XOR2_X2 U42 ( .A(n152), .B(n28), .Z(DIFF[5]) );
  XOR2_X2 U43 ( .A(n151), .B(n66), .Z(DIFF[6]) );
  AND2_X4 U44 ( .A1(n108), .A2(n27), .ZN(n44) );
  AND2_X4 U45 ( .A1(n110), .A2(n16), .ZN(n45) );
  AND2_X4 U46 ( .A1(n112), .A2(n31), .ZN(n46) );
  AND2_X4 U47 ( .A1(n114), .A2(n32), .ZN(n47) );
  AND2_X4 U48 ( .A1(n116), .A2(n33), .ZN(n48) );
  AND2_X4 U49 ( .A1(n118), .A2(n34), .ZN(n49) );
  AND2_X4 U50 ( .A1(n120), .A2(n29), .ZN(n50) );
  AND2_X4 U51 ( .A1(n122), .A2(n17), .ZN(n51) );
  AND2_X4 U52 ( .A1(n124), .A2(n18), .ZN(n52) );
  AND2_X4 U53 ( .A1(n126), .A2(n19), .ZN(n53) );
  AND2_X4 U54 ( .A1(n128), .A2(n20), .ZN(n54) );
  AND2_X4 U55 ( .A1(n130), .A2(n21), .ZN(n55) );
  AND2_X4 U56 ( .A1(n132), .A2(n22), .ZN(n56) );
  AND2_X4 U57 ( .A1(n134), .A2(n23), .ZN(n57) );
  AND2_X4 U58 ( .A1(n136), .A2(n24), .ZN(n58) );
  AND2_X4 U59 ( .A1(n138), .A2(n25), .ZN(n59) );
  AND2_X4 U60 ( .A1(n140), .A2(n26), .ZN(n60) );
  AND2_X4 U61 ( .A1(n142), .A2(n11), .ZN(n61) );
  AND2_X4 U62 ( .A1(n144), .A2(n12), .ZN(n62) );
  AND2_X4 U63 ( .A1(n146), .A2(n13), .ZN(n63) );
  AND2_X4 U64 ( .A1(n148), .A2(n14), .ZN(n64) );
  AND2_X4 U65 ( .A1(n150), .A2(n15), .ZN(n65) );
  AND2_X4 U66 ( .A1(n152), .A2(n28), .ZN(n66) );
  AND2_X4 U67 ( .A1(n154), .A2(n30), .ZN(n67) );
  AND2_X4 U68 ( .A1(n156), .A2(n157), .ZN(n68) );
  XOR2_X2 U69 ( .A(n121), .B(n51), .Z(DIFF[36]) );
  XOR2_X2 U70 ( .A(n111), .B(n46), .Z(DIFF[46]) );
  XOR2_X2 U71 ( .A(n110), .B(n16), .Z(DIFF[47]) );
  XOR2_X2 U72 ( .A(n108), .B(n27), .Z(DIFF[49]) );
  XOR2_X2 U73 ( .A(n106), .B(n10), .Z(DIFF[51]) );
  XOR2_X2 U74 ( .A(n105), .B(n1), .Z(DIFF[52]) );
  XOR2_X2 U75 ( .A(n143), .B(n62), .Z(DIFF[14]) );
  XOR2_X2 U76 ( .A(n142), .B(n11), .Z(DIFF[15]) );
  XOR2_X2 U77 ( .A(n141), .B(n61), .Z(DIFF[16]) );
  XOR2_X2 U78 ( .A(n140), .B(n26), .Z(DIFF[17]) );
  XOR2_X2 U79 ( .A(n139), .B(n60), .Z(DIFF[18]) );
  XOR2_X2 U80 ( .A(n138), .B(n25), .Z(DIFF[19]) );
  XOR2_X2 U81 ( .A(n137), .B(n59), .Z(DIFF[20]) );
  XOR2_X2 U82 ( .A(n136), .B(n24), .Z(DIFF[21]) );
  XOR2_X2 U83 ( .A(n135), .B(n58), .Z(DIFF[22]) );
  XOR2_X2 U84 ( .A(n134), .B(n23), .Z(DIFF[23]) );
  XOR2_X2 U85 ( .A(n133), .B(n57), .Z(DIFF[24]) );
  XOR2_X2 U86 ( .A(n132), .B(n22), .Z(DIFF[25]) );
  XOR2_X2 U87 ( .A(n131), .B(n56), .Z(DIFF[26]) );
  XOR2_X2 U88 ( .A(n130), .B(n21), .Z(DIFF[27]) );
  XOR2_X2 U89 ( .A(n129), .B(n55), .Z(DIFF[28]) );
  XOR2_X2 U90 ( .A(n128), .B(n20), .Z(DIFF[29]) );
  XOR2_X2 U91 ( .A(n127), .B(n54), .Z(DIFF[30]) );
  XOR2_X2 U92 ( .A(n126), .B(n19), .Z(DIFF[31]) );
  XOR2_X2 U93 ( .A(n125), .B(n53), .Z(DIFF[32]) );
  XOR2_X2 U94 ( .A(n124), .B(n18), .Z(DIFF[33]) );
  XOR2_X2 U95 ( .A(n123), .B(n52), .Z(DIFF[34]) );
  XOR2_X2 U96 ( .A(n122), .B(n17), .Z(DIFF[35]) );
  XOR2_X2 U97 ( .A(n150), .B(n15), .Z(DIFF[7]) );
  XOR2_X2 U98 ( .A(n149), .B(n65), .Z(DIFF[8]) );
  XOR2_X2 U99 ( .A(n148), .B(n14), .Z(DIFF[9]) );
  XOR2_X2 U100 ( .A(n147), .B(n64), .Z(DIFF[10]) );
  XOR2_X2 U101 ( .A(n146), .B(n13), .Z(DIFF[11]) );
  XOR2_X2 U102 ( .A(n145), .B(n63), .Z(DIFF[12]) );
  XOR2_X2 U103 ( .A(n144), .B(n12), .Z(DIFF[13]) );
  NAND2_X2 U104 ( .A1(n105), .A2(n1), .ZN(DIFF[53]) );
  INV_X4 U105 ( .A(B[52]), .ZN(n105) );
  INV_X4 U106 ( .A(B[51]), .ZN(n106) );
  INV_X4 U107 ( .A(B[50]), .ZN(n107) );
  INV_X4 U108 ( .A(B[49]), .ZN(n108) );
  INV_X4 U109 ( .A(B[48]), .ZN(n109) );
  INV_X4 U110 ( .A(B[47]), .ZN(n110) );
  INV_X4 U111 ( .A(B[46]), .ZN(n111) );
  INV_X4 U112 ( .A(B[45]), .ZN(n112) );
  INV_X4 U113 ( .A(B[44]), .ZN(n113) );
  INV_X4 U114 ( .A(B[43]), .ZN(n114) );
  INV_X4 U115 ( .A(B[42]), .ZN(n115) );
  INV_X4 U116 ( .A(B[41]), .ZN(n116) );
  INV_X4 U117 ( .A(B[40]), .ZN(n117) );
  INV_X4 U118 ( .A(B[39]), .ZN(n118) );
  INV_X4 U119 ( .A(B[38]), .ZN(n119) );
  INV_X4 U120 ( .A(B[37]), .ZN(n120) );
  INV_X4 U121 ( .A(B[36]), .ZN(n121) );
  INV_X4 U122 ( .A(B[35]), .ZN(n122) );
  INV_X4 U123 ( .A(B[34]), .ZN(n123) );
  INV_X4 U124 ( .A(B[33]), .ZN(n124) );
  INV_X4 U125 ( .A(B[32]), .ZN(n125) );
  INV_X4 U126 ( .A(B[31]), .ZN(n126) );
  INV_X4 U127 ( .A(B[30]), .ZN(n127) );
  INV_X4 U128 ( .A(B[29]), .ZN(n128) );
  INV_X4 U129 ( .A(B[28]), .ZN(n129) );
  INV_X4 U130 ( .A(B[27]), .ZN(n130) );
  INV_X4 U131 ( .A(B[26]), .ZN(n131) );
  INV_X4 U132 ( .A(B[25]), .ZN(n132) );
  INV_X4 U133 ( .A(B[24]), .ZN(n133) );
  INV_X4 U134 ( .A(B[23]), .ZN(n134) );
  INV_X4 U135 ( .A(B[22]), .ZN(n135) );
  INV_X4 U136 ( .A(B[21]), .ZN(n136) );
  INV_X4 U137 ( .A(B[20]), .ZN(n137) );
  INV_X4 U138 ( .A(B[19]), .ZN(n138) );
  INV_X4 U139 ( .A(B[18]), .ZN(n139) );
  INV_X4 U140 ( .A(B[17]), .ZN(n140) );
  INV_X4 U141 ( .A(B[16]), .ZN(n141) );
  INV_X4 U142 ( .A(B[15]), .ZN(n142) );
  INV_X4 U143 ( .A(B[14]), .ZN(n143) );
  INV_X4 U144 ( .A(B[13]), .ZN(n144) );
  INV_X4 U145 ( .A(B[12]), .ZN(n145) );
  INV_X4 U146 ( .A(B[11]), .ZN(n146) );
  INV_X4 U147 ( .A(B[10]), .ZN(n147) );
  INV_X4 U148 ( .A(B[9]), .ZN(n148) );
  INV_X4 U149 ( .A(B[8]), .ZN(n149) );
  INV_X4 U150 ( .A(B[7]), .ZN(n150) );
  INV_X4 U151 ( .A(B[6]), .ZN(n151) );
  INV_X4 U152 ( .A(B[5]), .ZN(n152) );
  INV_X4 U153 ( .A(B[4]), .ZN(n153) );
  INV_X4 U154 ( .A(B[3]), .ZN(n154) );
  INV_X4 U155 ( .A(B[2]), .ZN(n155) );
  INV_X4 U156 ( .A(B[1]), .ZN(n156) );
  INV_X4 U157 ( .A(\B[0] ), .ZN(n157) );
endmodule


module fpu_DW01_ash_2 ( A, DATA_TC, SH, SH_TC, B );
  input [52:0] A;
  input [4:0] SH;
  output [52:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][52] , \ML_int[1][51] , \ML_int[1][50] , \ML_int[1][49] ,
         \ML_int[1][48] , \ML_int[1][47] , \ML_int[1][46] , \ML_int[1][45] ,
         \ML_int[1][44] , \ML_int[1][43] , \ML_int[1][42] , \ML_int[1][41] ,
         \ML_int[1][40] , \ML_int[1][39] , \ML_int[1][38] , \ML_int[1][37] ,
         \ML_int[1][36] , \ML_int[1][35] , \ML_int[1][34] , \ML_int[1][33] ,
         \ML_int[1][32] , \ML_int[1][31] , \ML_int[1][30] , \ML_int[1][29] ,
         \ML_int[1][28] , \ML_int[1][27] , \ML_int[1][26] , \ML_int[1][25] ,
         \ML_int[1][24] , \ML_int[1][23] , \ML_int[1][22] , \ML_int[1][21] ,
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
         \ML_int[1][20] , \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] ,
         \ML_int[1][16] , \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] ,
         \ML_int[1][12] , \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] ,
         \ML_int[1][8] , \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] ,
         \ML_int[1][4] , \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] ,
<<<<<<< HEAD
         \ML_int[1][0] , \ML_int[2][27] , \ML_int[2][26] , \ML_int[2][25] ,
         \ML_int[2][24] , \ML_int[2][23] , \ML_int[2][22] , \ML_int[2][21] ,
         \ML_int[2][20] , \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] ,
         \ML_int[2][16] , \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] ,
         \ML_int[2][12] , \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] ,
         \ML_int[2][8] , \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] ,
         \ML_int[2][4] , \ML_int[2][3] , \ML_int[2][2] , \ML_int[3][27] ,
         \ML_int[3][26] , \ML_int[3][25] , \ML_int[3][24] , \ML_int[3][23] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] ,
         \ML_int[3][8] , \ML_int[3][7] , \ML_int[3][3] , \ML_int[3][2] ,
         \ML_int[3][1] , \ML_int[3][0] , \ML_int[4][27] , \ML_int[4][26] ,
         \ML_int[4][25] , \ML_int[4][24] , \ML_int[4][23] , \ML_int[4][11] ,
         \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] , \ML_int[4][7] ,
         \ML_int[5][27] , \ML_int[5][26] , \ML_int[5][25] , \ML_int[5][24] ,
         \ML_int[5][23] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36;
=======
         \ML_int[1][0] , \ML_int[2][52] , \ML_int[2][51] , \ML_int[2][50] ,
         \ML_int[2][49] , \ML_int[2][48] , \ML_int[2][47] , \ML_int[2][46] ,
         \ML_int[2][45] , \ML_int[2][44] , \ML_int[2][43] , \ML_int[2][42] ,
         \ML_int[2][41] , \ML_int[2][40] , \ML_int[2][39] , \ML_int[2][38] ,
         \ML_int[2][37] , \ML_int[2][36] , \ML_int[2][35] , \ML_int[2][34] ,
         \ML_int[2][33] , \ML_int[2][32] , \ML_int[2][31] , \ML_int[2][30] ,
         \ML_int[2][29] , \ML_int[2][28] , \ML_int[2][27] , \ML_int[2][26] ,
         \ML_int[2][25] , \ML_int[2][24] , \ML_int[2][23] , \ML_int[2][22] ,
         \ML_int[2][21] , \ML_int[2][20] , \ML_int[2][19] , \ML_int[2][18] ,
         \ML_int[2][17] , \ML_int[2][16] , \ML_int[2][15] , \ML_int[2][14] ,
         \ML_int[2][13] , \ML_int[2][12] , \ML_int[2][11] , \ML_int[2][10] ,
         \ML_int[2][9] , \ML_int[2][8] , \ML_int[2][7] , \ML_int[2][6] ,
         \ML_int[2][5] , \ML_int[2][4] , \ML_int[2][3] , \ML_int[2][2] ,
         \ML_int[2][1] , \ML_int[2][0] , \ML_int[3][52] , \ML_int[3][51] ,
         \ML_int[3][50] , \ML_int[3][49] , \ML_int[3][48] , \ML_int[3][47] ,
         \ML_int[3][46] , \ML_int[3][45] , \ML_int[3][44] , \ML_int[3][43] ,
         \ML_int[3][42] , \ML_int[3][41] , \ML_int[3][40] , \ML_int[3][39] ,
         \ML_int[3][38] , \ML_int[3][37] , \ML_int[3][36] , \ML_int[3][35] ,
         \ML_int[3][34] , \ML_int[3][33] , \ML_int[3][32] , \ML_int[3][31] ,
         \ML_int[3][30] , \ML_int[3][29] , \ML_int[3][28] , \ML_int[3][27] ,
         \ML_int[3][26] , \ML_int[3][25] , \ML_int[3][24] , \ML_int[3][23] ,
         \ML_int[3][22] , \ML_int[3][21] , \ML_int[3][20] , \ML_int[3][19] ,
         \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] , \ML_int[3][15] ,
         \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] , \ML_int[3][11] ,
         \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] , \ML_int[3][7] ,
         \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] , \ML_int[3][3] ,
         \ML_int[3][2] , \ML_int[3][1] , \ML_int[3][0] , \ML_int[4][52] ,
         \ML_int[4][51] , \ML_int[4][50] , \ML_int[4][49] , \ML_int[4][48] ,
         \ML_int[4][47] , \ML_int[4][46] , \ML_int[4][45] , \ML_int[4][44] ,
         \ML_int[4][43] , \ML_int[4][42] , \ML_int[4][41] , \ML_int[4][40] ,
         \ML_int[4][39] , \ML_int[4][38] , \ML_int[4][37] , \ML_int[4][36] ,
         \ML_int[4][35] , \ML_int[4][34] , \ML_int[4][33] , \ML_int[4][32] ,
         \ML_int[4][31] , \ML_int[4][30] , \ML_int[4][29] , \ML_int[4][28] ,
         \ML_int[4][27] , \ML_int[4][26] , \ML_int[4][25] , \ML_int[4][24] ,
         \ML_int[4][23] , \ML_int[4][22] , \ML_int[4][21] , \ML_int[4][20] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][16] ,
         \ML_int[4][15] , \ML_int[4][14] , \ML_int[4][13] , \ML_int[4][12] ,
         \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] ,
         \ML_int[5][52] , \ML_int[5][51] , \ML_int[5][50] , \ML_int[5][49] ,
         \ML_int[5][48] , \ML_int[5][47] , \ML_int[5][46] , \ML_int[5][45] ,
         \ML_int[5][44] , \ML_int[5][43] , \ML_int[5][42] , \ML_int[5][41] ,
         \ML_int[5][40] , \ML_int[5][39] , \ML_int[5][38] , \ML_int[5][37] ,
         \ML_int[5][36] , \ML_int[5][35] , \ML_int[5][34] , \ML_int[5][33] ,
         \ML_int[5][32] , \ML_int[5][31] , \ML_int[5][30] , \ML_int[5][29] ,
         \ML_int[5][28] , \ML_int[5][27] , \ML_int[5][26] , \ML_int[5][25] ,
         \ML_int[5][24] , \ML_int[5][23] , \ML_int[5][22] , \ML_int[5][21] ,
         \ML_int[5][20] , \ML_int[5][19] , \ML_int[5][18] , \ML_int[5][17] ,
         \ML_int[5][16] , \ML_int[5][15] , \ML_int[5][14] , \ML_int[5][13] ,
         \ML_int[5][12] , \ML_int[5][11] , \ML_int[5][10] , \ML_int[5][9] ,
         \ML_int[5][8] , \ML_int[5][7] , \ML_int[5][6] , \ML_int[5][5] ,
         \ML_int[5][4] , \ML_int[5][3] , \ML_int[5][2] , \ML_int[5][1] ,
         \ML_int[5][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30;
  assign B[52] = \ML_int[5][52] ;
  assign B[51] = \ML_int[5][51] ;
  assign B[50] = \ML_int[5][50] ;
  assign B[49] = \ML_int[5][49] ;
  assign B[48] = \ML_int[5][48] ;
  assign B[47] = \ML_int[5][47] ;
  assign B[46] = \ML_int[5][46] ;
  assign B[45] = \ML_int[5][45] ;
  assign B[44] = \ML_int[5][44] ;
  assign B[43] = \ML_int[5][43] ;
  assign B[42] = \ML_int[5][42] ;
  assign B[41] = \ML_int[5][41] ;
  assign B[40] = \ML_int[5][40] ;
  assign B[39] = \ML_int[5][39] ;
  assign B[38] = \ML_int[5][38] ;
  assign B[37] = \ML_int[5][37] ;
  assign B[36] = \ML_int[5][36] ;
  assign B[35] = \ML_int[5][35] ;
  assign B[34] = \ML_int[5][34] ;
  assign B[33] = \ML_int[5][33] ;
  assign B[32] = \ML_int[5][32] ;
  assign B[31] = \ML_int[5][31] ;
  assign B[30] = \ML_int[5][30] ;
  assign B[29] = \ML_int[5][29] ;
  assign B[28] = \ML_int[5][28] ;
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  assign B[27] = \ML_int[5][27] ;
  assign B[26] = \ML_int[5][26] ;
  assign B[25] = \ML_int[5][25] ;
  assign B[24] = \ML_int[5][24] ;
  assign B[23] = \ML_int[5][23] ;
<<<<<<< HEAD

  MUX2_X2 M1_4_27 ( .A(\ML_int[4][27] ), .B(\ML_int[4][11] ), .S(SH[4]), .Z(
        \ML_int[5][27] ) );
  MUX2_X2 M1_4_26 ( .A(\ML_int[4][26] ), .B(\ML_int[4][10] ), .S(SH[4]), .Z(
        \ML_int[5][26] ) );
  MUX2_X2 M1_4_23 ( .A(\ML_int[4][23] ), .B(\ML_int[4][7] ), .S(SH[4]), .Z(
        \ML_int[5][23] ) );
=======
  assign B[22] = \ML_int[5][22] ;
  assign B[21] = \ML_int[5][21] ;
  assign B[20] = \ML_int[5][20] ;
  assign B[19] = \ML_int[5][19] ;
  assign B[18] = \ML_int[5][18] ;
  assign B[17] = \ML_int[5][17] ;
  assign B[16] = \ML_int[5][16] ;
  assign B[15] = \ML_int[5][15] ;
  assign B[14] = \ML_int[5][14] ;
  assign B[13] = \ML_int[5][13] ;
  assign B[12] = \ML_int[5][12] ;
  assign B[11] = \ML_int[5][11] ;
  assign B[10] = \ML_int[5][10] ;
  assign B[9] = \ML_int[5][9] ;
  assign B[8] = \ML_int[5][8] ;
  assign B[7] = \ML_int[5][7] ;
  assign B[6] = \ML_int[5][6] ;
  assign B[5] = \ML_int[5][5] ;
  assign B[4] = \ML_int[5][4] ;
  assign B[3] = \ML_int[5][3] ;
  assign B[2] = \ML_int[5][2] ;
  assign B[1] = \ML_int[5][1] ;
  assign B[0] = \ML_int[5][0] ;

  MUX2_X2 M1_4_52 ( .A(\ML_int[4][52] ), .B(\ML_int[4][36] ), .S(n11), .Z(
        \ML_int[5][52] ) );
  MUX2_X2 M1_4_51 ( .A(\ML_int[4][51] ), .B(\ML_int[4][35] ), .S(SH[4]), .Z(
        \ML_int[5][51] ) );
  MUX2_X2 M1_4_50 ( .A(\ML_int[4][50] ), .B(\ML_int[4][34] ), .S(SH[4]), .Z(
        \ML_int[5][50] ) );
  MUX2_X2 M1_4_49 ( .A(\ML_int[4][49] ), .B(\ML_int[4][33] ), .S(SH[4]), .Z(
        \ML_int[5][49] ) );
  MUX2_X2 M1_4_48 ( .A(\ML_int[4][48] ), .B(\ML_int[4][32] ), .S(SH[4]), .Z(
        \ML_int[5][48] ) );
  MUX2_X2 M1_4_47 ( .A(\ML_int[4][47] ), .B(\ML_int[4][31] ), .S(n11), .Z(
        \ML_int[5][47] ) );
  MUX2_X2 M1_4_46 ( .A(\ML_int[4][46] ), .B(\ML_int[4][30] ), .S(SH[4]), .Z(
        \ML_int[5][46] ) );
  MUX2_X2 M1_4_45 ( .A(\ML_int[4][45] ), .B(\ML_int[4][29] ), .S(SH[4]), .Z(
        \ML_int[5][45] ) );
  MUX2_X2 M1_4_44 ( .A(\ML_int[4][44] ), .B(\ML_int[4][28] ), .S(SH[4]), .Z(
        \ML_int[5][44] ) );
  MUX2_X2 M1_4_43 ( .A(\ML_int[4][43] ), .B(\ML_int[4][27] ), .S(SH[4]), .Z(
        \ML_int[5][43] ) );
  MUX2_X2 M1_4_42 ( .A(\ML_int[4][42] ), .B(\ML_int[4][26] ), .S(SH[4]), .Z(
        \ML_int[5][42] ) );
  MUX2_X2 M1_4_41 ( .A(\ML_int[4][41] ), .B(\ML_int[4][25] ), .S(n13), .Z(
        \ML_int[5][41] ) );
  MUX2_X2 M1_4_40 ( .A(\ML_int[4][40] ), .B(\ML_int[4][24] ), .S(n13), .Z(
        \ML_int[5][40] ) );
  MUX2_X2 M1_4_39 ( .A(\ML_int[4][39] ), .B(\ML_int[4][23] ), .S(n13), .Z(
        \ML_int[5][39] ) );
  MUX2_X2 M1_4_38 ( .A(\ML_int[4][38] ), .B(\ML_int[4][22] ), .S(n13), .Z(
        \ML_int[5][38] ) );
  MUX2_X2 M1_4_37 ( .A(\ML_int[4][37] ), .B(\ML_int[4][21] ), .S(n13), .Z(
        \ML_int[5][37] ) );
  MUX2_X2 M1_4_36 ( .A(\ML_int[4][36] ), .B(\ML_int[4][20] ), .S(n13), .Z(
        \ML_int[5][36] ) );
  MUX2_X2 M1_4_35 ( .A(\ML_int[4][35] ), .B(\ML_int[4][19] ), .S(n13), .Z(
        \ML_int[5][35] ) );
  MUX2_X2 M1_4_34 ( .A(\ML_int[4][34] ), .B(\ML_int[4][18] ), .S(n13), .Z(
        \ML_int[5][34] ) );
  MUX2_X2 M1_4_33 ( .A(\ML_int[4][33] ), .B(\ML_int[4][17] ), .S(n13), .Z(
        \ML_int[5][33] ) );
  MUX2_X2 M1_4_32 ( .A(\ML_int[4][32] ), .B(\ML_int[4][16] ), .S(n13), .Z(
        \ML_int[5][32] ) );
  MUX2_X2 M1_4_31 ( .A(\ML_int[4][31] ), .B(\ML_int[4][15] ), .S(n13), .Z(
        \ML_int[5][31] ) );
  MUX2_X2 M1_4_30 ( .A(\ML_int[4][30] ), .B(\ML_int[4][14] ), .S(n14), .Z(
        \ML_int[5][30] ) );
  MUX2_X2 M1_4_29 ( .A(\ML_int[4][29] ), .B(\ML_int[4][13] ), .S(n14), .Z(
        \ML_int[5][29] ) );
  MUX2_X2 M1_4_28 ( .A(\ML_int[4][28] ), .B(\ML_int[4][12] ), .S(n14), .Z(
        \ML_int[5][28] ) );
  MUX2_X2 M1_4_27 ( .A(\ML_int[4][27] ), .B(\ML_int[4][11] ), .S(n14), .Z(
        \ML_int[5][27] ) );
  MUX2_X2 M1_4_26 ( .A(\ML_int[4][26] ), .B(\ML_int[4][10] ), .S(n14), .Z(
        \ML_int[5][26] ) );
  MUX2_X2 M1_4_25 ( .A(\ML_int[4][25] ), .B(\ML_int[4][9] ), .S(n14), .Z(
        \ML_int[5][25] ) );
  MUX2_X2 M1_4_24 ( .A(\ML_int[4][24] ), .B(\ML_int[4][8] ), .S(n14), .Z(
        \ML_int[5][24] ) );
  MUX2_X2 M1_4_23 ( .A(\ML_int[4][23] ), .B(n22), .S(n14), .Z(\ML_int[5][23] )
         );
  MUX2_X2 M1_4_22 ( .A(\ML_int[4][22] ), .B(n21), .S(n14), .Z(\ML_int[5][22] )
         );
  MUX2_X2 M1_4_21 ( .A(\ML_int[4][21] ), .B(n20), .S(n14), .Z(\ML_int[5][21] )
         );
  MUX2_X2 M1_4_20 ( .A(\ML_int[4][20] ), .B(n19), .S(n14), .Z(\ML_int[5][20] )
         );
  MUX2_X2 M1_4_19 ( .A(\ML_int[4][19] ), .B(n15), .S(n11), .Z(\ML_int[5][19] )
         );
  MUX2_X2 M1_4_18 ( .A(\ML_int[4][18] ), .B(n16), .S(n13), .Z(\ML_int[5][18] )
         );
  MUX2_X2 M1_4_17 ( .A(\ML_int[4][17] ), .B(n17), .S(n14), .Z(\ML_int[5][17] )
         );
  MUX2_X2 M1_4_16 ( .A(\ML_int[4][16] ), .B(n18), .S(n11), .Z(\ML_int[5][16] )
         );
  MUX2_X2 M1_3_52 ( .A(\ML_int[3][52] ), .B(\ML_int[3][44] ), .S(n9), .Z(
        \ML_int[4][52] ) );
  MUX2_X2 M1_3_51 ( .A(\ML_int[3][51] ), .B(\ML_int[3][43] ), .S(n9), .Z(
        \ML_int[4][51] ) );
  MUX2_X2 M1_3_50 ( .A(\ML_int[3][50] ), .B(\ML_int[3][42] ), .S(n9), .Z(
        \ML_int[4][50] ) );
  MUX2_X2 M1_3_49 ( .A(\ML_int[3][49] ), .B(\ML_int[3][41] ), .S(n9), .Z(
        \ML_int[4][49] ) );
  MUX2_X2 M1_3_48 ( .A(\ML_int[3][48] ), .B(\ML_int[3][40] ), .S(n9), .Z(
        \ML_int[4][48] ) );
  MUX2_X2 M1_3_47 ( .A(\ML_int[3][47] ), .B(\ML_int[3][39] ), .S(n9), .Z(
        \ML_int[4][47] ) );
  MUX2_X2 M1_3_46 ( .A(\ML_int[3][46] ), .B(\ML_int[3][38] ), .S(n9), .Z(
        \ML_int[4][46] ) );
  MUX2_X2 M1_3_45 ( .A(\ML_int[3][45] ), .B(\ML_int[3][37] ), .S(n9), .Z(
        \ML_int[4][45] ) );
  MUX2_X2 M1_3_44 ( .A(\ML_int[3][44] ), .B(\ML_int[3][36] ), .S(n9), .Z(
        \ML_int[4][44] ) );
  MUX2_X2 M1_3_43 ( .A(\ML_int[3][43] ), .B(\ML_int[3][35] ), .S(n9), .Z(
        \ML_int[4][43] ) );
  MUX2_X2 M1_3_42 ( .A(\ML_int[3][42] ), .B(\ML_int[3][34] ), .S(n9), .Z(
        \ML_int[4][42] ) );
  MUX2_X2 M1_3_41 ( .A(\ML_int[3][41] ), .B(\ML_int[3][33] ), .S(n9), .Z(
        \ML_int[4][41] ) );
  MUX2_X2 M1_3_40 ( .A(\ML_int[3][40] ), .B(\ML_int[3][32] ), .S(n9), .Z(
        \ML_int[4][40] ) );
  MUX2_X2 M1_3_39 ( .A(\ML_int[3][39] ), .B(\ML_int[3][31] ), .S(n9), .Z(
        \ML_int[4][39] ) );
  MUX2_X2 M1_3_38 ( .A(\ML_int[3][38] ), .B(\ML_int[3][30] ), .S(n9), .Z(
        \ML_int[4][38] ) );
  MUX2_X2 M1_3_37 ( .A(\ML_int[3][37] ), .B(\ML_int[3][29] ), .S(n9), .Z(
        \ML_int[4][37] ) );
  MUX2_X2 M1_3_36 ( .A(\ML_int[3][36] ), .B(\ML_int[3][28] ), .S(n9), .Z(
        \ML_int[4][36] ) );
  MUX2_X2 M1_3_35 ( .A(\ML_int[3][35] ), .B(\ML_int[3][27] ), .S(n9), .Z(
        \ML_int[4][35] ) );
  MUX2_X2 M1_3_34 ( .A(\ML_int[3][34] ), .B(\ML_int[3][26] ), .S(n9), .Z(
        \ML_int[4][34] ) );
  MUX2_X2 M1_3_33 ( .A(\ML_int[3][33] ), .B(\ML_int[3][25] ), .S(n9), .Z(
        \ML_int[4][33] ) );
  MUX2_X2 M1_3_32 ( .A(\ML_int[3][32] ), .B(\ML_int[3][24] ), .S(n9), .Z(
        \ML_int[4][32] ) );
  MUX2_X2 M1_3_31 ( .A(\ML_int[3][31] ), .B(\ML_int[3][23] ), .S(n9), .Z(
        \ML_int[4][31] ) );
  MUX2_X2 M1_3_30 ( .A(\ML_int[3][30] ), .B(\ML_int[3][22] ), .S(n9), .Z(
        \ML_int[4][30] ) );
  MUX2_X2 M1_3_29 ( .A(\ML_int[3][29] ), .B(\ML_int[3][21] ), .S(SH[3]), .Z(
        \ML_int[4][29] ) );
  MUX2_X2 M1_3_28 ( .A(\ML_int[3][28] ), .B(\ML_int[3][20] ), .S(SH[3]), .Z(
        \ML_int[4][28] ) );
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  MUX2_X2 M1_3_27 ( .A(\ML_int[3][27] ), .B(\ML_int[3][19] ), .S(SH[3]), .Z(
        \ML_int[4][27] ) );
  MUX2_X2 M1_3_26 ( .A(\ML_int[3][26] ), .B(\ML_int[3][18] ), .S(SH[3]), .Z(
        \ML_int[4][26] ) );
<<<<<<< HEAD
  MUX2_X2 M1_3_23 ( .A(\ML_int[3][23] ), .B(\ML_int[3][15] ), .S(SH[3]), .Z(
        \ML_int[4][23] ) );
=======
  MUX2_X2 M1_3_25 ( .A(\ML_int[3][25] ), .B(\ML_int[3][17] ), .S(SH[3]), .Z(
        \ML_int[4][25] ) );
  MUX2_X2 M1_3_24 ( .A(\ML_int[3][24] ), .B(\ML_int[3][16] ), .S(SH[3]), .Z(
        \ML_int[4][24] ) );
  MUX2_X2 M1_3_23 ( .A(\ML_int[3][23] ), .B(\ML_int[3][15] ), .S(SH[3]), .Z(
        \ML_int[4][23] ) );
  MUX2_X2 M1_3_22 ( .A(\ML_int[3][22] ), .B(\ML_int[3][14] ), .S(SH[3]), .Z(
        \ML_int[4][22] ) );
  MUX2_X2 M1_3_21 ( .A(\ML_int[3][21] ), .B(\ML_int[3][13] ), .S(SH[3]), .Z(
        \ML_int[4][21] ) );
  MUX2_X2 M1_3_20 ( .A(\ML_int[3][20] ), .B(\ML_int[3][12] ), .S(SH[3]), .Z(
        \ML_int[4][20] ) );
  MUX2_X2 M1_3_19 ( .A(\ML_int[3][19] ), .B(\ML_int[3][11] ), .S(SH[3]), .Z(
        \ML_int[4][19] ) );
  MUX2_X2 M1_3_18 ( .A(\ML_int[3][18] ), .B(\ML_int[3][10] ), .S(n9), .Z(
        \ML_int[4][18] ) );
  MUX2_X2 M1_3_17 ( .A(\ML_int[3][17] ), .B(\ML_int[3][9] ), .S(SH[3]), .Z(
        \ML_int[4][17] ) );
  MUX2_X2 M1_3_16 ( .A(\ML_int[3][16] ), .B(\ML_int[3][8] ), .S(SH[3]), .Z(
        \ML_int[4][16] ) );
  MUX2_X2 M1_3_15 ( .A(\ML_int[3][15] ), .B(\ML_int[3][7] ), .S(SH[3]), .Z(
        \ML_int[4][15] ) );
  MUX2_X2 M1_3_14 ( .A(\ML_int[3][14] ), .B(\ML_int[3][6] ), .S(SH[3]), .Z(
        \ML_int[4][14] ) );
  MUX2_X2 M1_3_13 ( .A(\ML_int[3][13] ), .B(\ML_int[3][5] ), .S(SH[3]), .Z(
        \ML_int[4][13] ) );
  MUX2_X2 M1_3_12 ( .A(\ML_int[3][12] ), .B(\ML_int[3][4] ), .S(SH[3]), .Z(
        \ML_int[4][12] ) );
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  MUX2_X2 M1_3_11 ( .A(\ML_int[3][11] ), .B(\ML_int[3][3] ), .S(SH[3]), .Z(
        \ML_int[4][11] ) );
  MUX2_X2 M1_3_10 ( .A(\ML_int[3][10] ), .B(\ML_int[3][2] ), .S(SH[3]), .Z(
        \ML_int[4][10] ) );
  MUX2_X2 M1_3_9 ( .A(\ML_int[3][9] ), .B(\ML_int[3][1] ), .S(SH[3]), .Z(
        \ML_int[4][9] ) );
<<<<<<< HEAD
  MUX2_X2 M1_2_27 ( .A(\ML_int[2][27] ), .B(\ML_int[2][23] ), .S(n28), .Z(
        \ML_int[3][27] ) );
  MUX2_X2 M1_2_26 ( .A(\ML_int[2][26] ), .B(\ML_int[2][22] ), .S(n28), .Z(
        \ML_int[3][26] ) );
  MUX2_X2 M1_2_25 ( .A(\ML_int[2][25] ), .B(\ML_int[2][21] ), .S(n28), .Z(
        \ML_int[3][25] ) );
  MUX2_X2 M1_2_24 ( .A(\ML_int[2][24] ), .B(\ML_int[2][20] ), .S(n28), .Z(
        \ML_int[3][24] ) );
  MUX2_X2 M1_2_23 ( .A(\ML_int[2][23] ), .B(\ML_int[2][19] ), .S(n28), .Z(
        \ML_int[3][23] ) );
  MUX2_X2 M1_2_19 ( .A(\ML_int[2][19] ), .B(\ML_int[2][15] ), .S(n28), .Z(
        \ML_int[3][19] ) );
  MUX2_X2 M1_2_18 ( .A(\ML_int[2][18] ), .B(\ML_int[2][14] ), .S(n28), .Z(
        \ML_int[3][18] ) );
  MUX2_X2 M1_2_15 ( .A(\ML_int[2][15] ), .B(\ML_int[2][11] ), .S(n28), .Z(
        \ML_int[3][15] ) );
  MUX2_X2 M1_2_11 ( .A(\ML_int[2][11] ), .B(\ML_int[2][7] ), .S(n28), .Z(
        \ML_int[3][11] ) );
  MUX2_X2 M1_2_10 ( .A(\ML_int[2][10] ), .B(\ML_int[2][6] ), .S(n28), .Z(
        \ML_int[3][10] ) );
  MUX2_X2 M1_2_9 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S(n28), .Z(
        \ML_int[3][9] ) );
  MUX2_X2 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(n28), .Z(
        \ML_int[3][8] ) );
  MUX2_X2 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(n28), .Z(
        \ML_int[3][7] ) );
  MUX2_X2 M1_1_27 ( .A(\ML_int[1][27] ), .B(\ML_int[1][27] ), .S(n32), .Z(
        \ML_int[2][27] ) );
  MUX2_X2 M1_1_26 ( .A(\ML_int[1][27] ), .B(\ML_int[1][24] ), .S(n32), .Z(
        \ML_int[2][26] ) );
  MUX2_X2 M1_1_23 ( .A(\ML_int[1][27] ), .B(\ML_int[1][21] ), .S(n32), .Z(
        \ML_int[2][23] ) );
  MUX2_X2 M1_1_22 ( .A(\ML_int[1][22] ), .B(\ML_int[1][20] ), .S(n32), .Z(
        \ML_int[2][22] ) );
  MUX2_X2 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S(n32), .Z(
        \ML_int[2][21] ) );
  MUX2_X2 M1_1_19 ( .A(\ML_int[1][19] ), .B(\ML_int[1][17] ), .S(n32), .Z(
        \ML_int[2][19] ) );
  MUX2_X2 M1_1_18 ( .A(\ML_int[1][18] ), .B(\ML_int[1][16] ), .S(n32), .Z(
        \ML_int[2][18] ) );
  MUX2_X2 M1_1_17 ( .A(\ML_int[1][17] ), .B(\ML_int[1][15] ), .S(n32), .Z(
        \ML_int[2][17] ) );
  MUX2_X2 M1_1_16 ( .A(\ML_int[1][16] ), .B(\ML_int[1][14] ), .S(n33), .Z(
        \ML_int[2][16] ) );
  MUX2_X2 M1_1_15 ( .A(\ML_int[1][15] ), .B(\ML_int[1][13] ), .S(n33), .Z(
        \ML_int[2][15] ) );
  MUX2_X2 M1_1_14 ( .A(\ML_int[1][14] ), .B(\ML_int[1][12] ), .S(n33), .Z(
        \ML_int[2][14] ) );
  MUX2_X2 M1_1_11 ( .A(\ML_int[1][11] ), .B(\ML_int[1][9] ), .S(n33), .Z(
        \ML_int[2][11] ) );
  MUX2_X2 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S(n33), .Z(
        \ML_int[2][10] ) );
  MUX2_X2 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S(n33), .Z(
        \ML_int[2][9] ) );
  MUX2_X2 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S(n33), .Z(
        \ML_int[2][8] ) );
  MUX2_X2 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S(n33), .Z(
        \ML_int[2][7] ) );
  MUX2_X2 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(n34), .Z(
        \ML_int[2][3] ) );
  MUX2_X2 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S(n34), .Z(
        \ML_int[2][2] ) );
  MUX2_X2 M1_0_24 ( .A(A[24]), .B(A[23]), .S(n30), .Z(\ML_int[1][24] ) );
  MUX2_X2 M1_0_22 ( .A(A[22]), .B(A[21]), .S(n30), .Z(\ML_int[1][22] ) );
  MUX2_X2 M1_0_21 ( .A(A[21]), .B(A[20]), .S(n30), .Z(\ML_int[1][21] ) );
  MUX2_X2 M1_0_20 ( .A(A[20]), .B(A[19]), .S(n30), .Z(\ML_int[1][20] ) );
  MUX2_X2 M1_0_19 ( .A(A[19]), .B(A[18]), .S(n30), .Z(\ML_int[1][19] ) );
  MUX2_X2 M1_0_18 ( .A(A[18]), .B(A[17]), .S(n30), .Z(\ML_int[1][18] ) );
  MUX2_X2 M1_0_17 ( .A(A[17]), .B(A[16]), .S(n30), .Z(\ML_int[1][17] ) );
  MUX2_X2 M1_0_16 ( .A(A[16]), .B(A[15]), .S(n30), .Z(\ML_int[1][16] ) );
  MUX2_X2 M1_0_15 ( .A(A[15]), .B(A[14]), .S(n30), .Z(\ML_int[1][15] ) );
  MUX2_X2 M1_0_14 ( .A(A[14]), .B(A[13]), .S(n30), .Z(\ML_int[1][14] ) );
  MUX2_X2 M1_0_13 ( .A(A[13]), .B(A[12]), .S(n30), .Z(\ML_int[1][13] ) );
  MUX2_X2 M1_0_12 ( .A(A[12]), .B(A[11]), .S(n30), .Z(\ML_int[1][12] ) );
  MUX2_X2 M1_0_11 ( .A(A[11]), .B(A[10]), .S(n29), .Z(\ML_int[1][11] ) );
  MUX2_X2 M1_0_10 ( .A(A[10]), .B(A[9]), .S(n29), .Z(\ML_int[1][10] ) );
  MUX2_X2 M1_0_9 ( .A(A[9]), .B(A[8]), .S(n29), .Z(\ML_int[1][9] ) );
  MUX2_X2 M1_0_8 ( .A(A[8]), .B(A[7]), .S(n29), .Z(\ML_int[1][8] ) );
  MUX2_X2 M1_0_7 ( .A(A[7]), .B(A[6]), .S(n29), .Z(\ML_int[1][7] ) );
  MUX2_X2 M1_0_6 ( .A(A[6]), .B(A[5]), .S(n29), .Z(\ML_int[1][6] ) );
  MUX2_X2 M1_0_4 ( .A(A[4]), .B(A[3]), .S(n29), .Z(\ML_int[1][4] ) );
  MUX2_X2 M1_0_3 ( .A(A[3]), .B(A[2]), .S(n29), .Z(\ML_int[1][3] ) );
  MUX2_X2 M1_0_2 ( .A(A[2]), .B(A[1]), .S(n29), .Z(\ML_int[1][2] ) );
  MUX2_X2 M1_0_1 ( .A(A[1]), .B(A[0]), .S(n29), .Z(\ML_int[1][1] ) );
  MUX2_X1 M1_2_16 ( .A(\ML_int[2][16] ), .B(\ML_int[2][12] ), .S(n28), .Z(
        \ML_int[3][16] ) );
  MUX2_X1 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S(n33), .Z(
        \ML_int[2][6] ) );
  MUX2_X2 M1_2_17 ( .A(\ML_int[2][17] ), .B(\ML_int[2][13] ), .S(n28), .Z(
        \ML_int[3][17] ) );
  MUX2_X2 M1_0_27 ( .A(A[27]), .B(A[26]), .S(n30), .Z(\ML_int[1][27] ) );
  NAND2_X1 U3 ( .A1(A[5]), .A2(n4), .ZN(n5) );
  NAND2_X4 U4 ( .A1(n25), .A2(n26), .ZN(\ML_int[5][25] ) );
  NAND2_X1 U5 ( .A1(\ML_int[1][3] ), .A2(n1), .ZN(n2) );
  NAND2_X2 U6 ( .A1(\ML_int[1][5] ), .A2(n35), .ZN(n3) );
  NAND2_X2 U7 ( .A1(n2), .A2(n3), .ZN(\ML_int[2][5] ) );
  INV_X1 U8 ( .A(n35), .ZN(n1) );
  NAND2_X1 U9 ( .A1(A[4]), .A2(n29), .ZN(n6) );
  NAND2_X2 U10 ( .A1(n5), .A2(n6), .ZN(\ML_int[1][5] ) );
  INV_X1 U11 ( .A(n29), .ZN(n4) );
  INV_X16 U12 ( .A(n31), .ZN(n30) );
  INV_X16 U13 ( .A(n31), .ZN(n29) );
  INV_X4 U14 ( .A(SH[0]), .ZN(n31) );
  INV_X4 U15 ( .A(n33), .ZN(n21) );
  INV_X4 U16 ( .A(SH[4]), .ZN(n24) );
  INV_X8 U17 ( .A(n27), .ZN(n28) );
  INV_X4 U18 ( .A(SH[2]), .ZN(n27) );
  NAND2_X4 U19 ( .A1(\ML_int[4][25] ), .A2(n24), .ZN(n25) );
  MUX2_X2 U20 ( .A(\ML_int[1][22] ), .B(\ML_int[1][24] ), .S(n21), .Z(
        \ML_int[2][24] ) );
  INV_X8 U21 ( .A(n35), .ZN(n32) );
  OAI21_X2 U22 ( .B1(n7), .B2(SH[3]), .A(n10), .ZN(\ML_int[4][25] ) );
  INV_X4 U23 ( .A(\ML_int[3][25] ), .ZN(n7) );
  NAND2_X2 U24 ( .A1(\ML_int[3][8] ), .A2(n16), .ZN(n8) );
  NAND2_X2 U25 ( .A1(\ML_int[3][0] ), .A2(SH[3]), .ZN(n9) );
  NAND2_X2 U26 ( .A1(n8), .A2(n9), .ZN(\ML_int[4][8] ) );
  NAND2_X4 U27 ( .A1(n17), .A2(n18), .ZN(\ML_int[4][24] ) );
  NAND2_X2 U28 ( .A1(\ML_int[3][16] ), .A2(SH[3]), .ZN(n18) );
  NAND2_X4 U29 ( .A1(\ML_int[4][8] ), .A2(SH[4]), .ZN(n20) );
  NAND2_X4 U30 ( .A1(n19), .A2(n20), .ZN(\ML_int[5][24] ) );
  NAND2_X4 U31 ( .A1(\ML_int[3][24] ), .A2(n16), .ZN(n17) );
  INV_X4 U32 ( .A(n35), .ZN(n34) );
  NAND2_X2 U33 ( .A1(\ML_int[4][9] ), .A2(SH[4]), .ZN(n26) );
  NAND2_X2 U34 ( .A1(\ML_int[3][17] ), .A2(SH[3]), .ZN(n10) );
  NAND2_X1 U35 ( .A1(\ML_int[1][13] ), .A2(n21), .ZN(n11) );
  NAND2_X1 U36 ( .A1(\ML_int[1][11] ), .A2(n33), .ZN(n12) );
  NAND2_X2 U37 ( .A1(n11), .A2(n12), .ZN(\ML_int[2][13] ) );
  NAND2_X1 U38 ( .A1(\ML_int[1][27] ), .A2(n13), .ZN(n14) );
  NAND2_X1 U39 ( .A1(\ML_int[1][27] ), .A2(n32), .ZN(n15) );
  NAND2_X2 U40 ( .A1(n14), .A2(n15), .ZN(\ML_int[2][25] ) );
  INV_X1 U41 ( .A(n32), .ZN(n13) );
  INV_X1 U42 ( .A(SH[3]), .ZN(n16) );
  NAND2_X4 U43 ( .A1(\ML_int[4][24] ), .A2(n24), .ZN(n19) );
  MUX2_X2 U44 ( .A(\ML_int[1][2] ), .B(\ML_int[1][4] ), .S(n35), .Z(
        \ML_int[2][4] ) );
  NAND2_X1 U45 ( .A1(\ML_int[1][12] ), .A2(n21), .ZN(n22) );
  NAND2_X1 U46 ( .A1(\ML_int[1][10] ), .A2(n33), .ZN(n23) );
  NAND2_X2 U47 ( .A1(n22), .A2(n23), .ZN(\ML_int[2][12] ) );
  MUX2_X2 U48 ( .A(\ML_int[1][18] ), .B(\ML_int[1][20] ), .S(n13), .Z(
        \ML_int[2][20] ) );
  INV_X32 U49 ( .A(n35), .ZN(n33) );
  INV_X32 U50 ( .A(SH[1]), .ZN(n35) );
  AND2_X1 U51 ( .A1(\ML_int[3][7] ), .A2(n16), .ZN(\ML_int[4][7] ) );
  AND2_X1 U52 ( .A1(\ML_int[2][3] ), .A2(n27), .ZN(\ML_int[3][3] ) );
  AND2_X1 U53 ( .A1(\ML_int[2][2] ), .A2(n27), .ZN(\ML_int[3][2] ) );
  AND2_X1 U54 ( .A1(\ML_int[1][1] ), .A2(n36), .ZN(\ML_int[3][1] ) );
  AND2_X1 U55 ( .A1(n36), .A2(\ML_int[1][0] ), .ZN(\ML_int[3][0] ) );
  NOR2_X1 U56 ( .A1(n32), .A2(n28), .ZN(n36) );
  AND2_X1 U57 ( .A1(A[0]), .A2(n31), .ZN(\ML_int[1][0] ) );
endmodule


module fpu_DW01_sub_7 ( A, B, CI, DIFF, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;
  wire   [14:1] carry;

  FA_X1 U2_13 ( .A(A[13]), .B(n18), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FA_X1 U2_12 ( .A(A[12]), .B(n17), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FA_X1 U2_11 ( .A(A[11]), .B(n16), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FA_X1 U2_10 ( .A(A[10]), .B(n15), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FA_X1 U2_9 ( .A(A[9]), .B(n14), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FA_X1 U2_8 ( .A(A[8]), .B(n13), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FA_X1 U2_7 ( .A(A[7]), .B(n12), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FA_X1 U2_6 ( .A(A[6]), .B(n11), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA_X1 U2_5 ( .A(A[5]), .B(n10), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n9), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_3 ( .A(A[3]), .B(n8), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA_X1 U2_2 ( .A(A[2]), .B(n7), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA_X1 U2_1 ( .A(A[1]), .B(n6), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  INV_X1 U1 ( .A(n3), .ZN(n1) );
  NAND2_X4 U2 ( .A1(n2), .A2(n3), .ZN(carry[1]) );
  XNOR2_X2 U3 ( .A(n5), .B(n1), .ZN(DIFF[0]) );
  INV_X4 U4 ( .A(n5), .ZN(n2) );
  INV_X4 U5 ( .A(A[0]), .ZN(n3) );
  INV_X4 U6 ( .A(carry[14]), .ZN(DIFF[14]) );
  INV_X4 U7 ( .A(B[0]), .ZN(n5) );
  INV_X4 U8 ( .A(B[1]), .ZN(n6) );
  INV_X4 U9 ( .A(B[2]), .ZN(n7) );
  INV_X4 U10 ( .A(B[3]), .ZN(n8) );
  INV_X4 U11 ( .A(B[4]), .ZN(n9) );
  INV_X4 U12 ( .A(B[5]), .ZN(n10) );
  INV_X4 U13 ( .A(B[6]), .ZN(n11) );
  INV_X4 U14 ( .A(B[7]), .ZN(n12) );
  INV_X4 U15 ( .A(B[8]), .ZN(n13) );
  INV_X4 U16 ( .A(B[9]), .ZN(n14) );
  INV_X4 U17 ( .A(B[10]), .ZN(n15) );
  INV_X4 U18 ( .A(B[11]), .ZN(n16) );
  INV_X4 U19 ( .A(B[12]), .ZN(n17) );
  INV_X4 U20 ( .A(B[13]), .ZN(n18) );
endmodule


module fpu_DW01_add_5 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n4;
  wire   [13:1] carry;

  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(SUM[14]), .S(SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
=======
  MUX2_X2 M1_3_8 ( .A(\ML_int[3][8] ), .B(\ML_int[3][0] ), .S(SH[3]), .Z(
        \ML_int[4][8] ) );
  MUX2_X2 M1_2_52 ( .A(\ML_int[2][52] ), .B(\ML_int[2][48] ), .S(n7), .Z(
        \ML_int[3][52] ) );
  MUX2_X2 M1_2_51 ( .A(\ML_int[2][51] ), .B(\ML_int[2][47] ), .S(n7), .Z(
        \ML_int[3][51] ) );
  MUX2_X2 M1_2_50 ( .A(\ML_int[2][50] ), .B(\ML_int[2][46] ), .S(n7), .Z(
        \ML_int[3][50] ) );
  MUX2_X2 M1_2_49 ( .A(\ML_int[2][49] ), .B(\ML_int[2][45] ), .S(n7), .Z(
        \ML_int[3][49] ) );
  MUX2_X2 M1_2_48 ( .A(\ML_int[2][48] ), .B(\ML_int[2][44] ), .S(n7), .Z(
        \ML_int[3][48] ) );
  MUX2_X2 M1_2_47 ( .A(\ML_int[2][47] ), .B(\ML_int[2][43] ), .S(n7), .Z(
        \ML_int[3][47] ) );
  MUX2_X2 M1_2_46 ( .A(\ML_int[2][46] ), .B(\ML_int[2][42] ), .S(n7), .Z(
        \ML_int[3][46] ) );
  MUX2_X2 M1_2_45 ( .A(\ML_int[2][45] ), .B(\ML_int[2][41] ), .S(n7), .Z(
        \ML_int[3][45] ) );
  MUX2_X2 M1_2_44 ( .A(\ML_int[2][44] ), .B(\ML_int[2][40] ), .S(n7), .Z(
        \ML_int[3][44] ) );
  MUX2_X2 M1_2_43 ( .A(\ML_int[2][43] ), .B(\ML_int[2][39] ), .S(n7), .Z(
        \ML_int[3][43] ) );
  MUX2_X2 M1_2_42 ( .A(\ML_int[2][42] ), .B(\ML_int[2][38] ), .S(n7), .Z(
        \ML_int[3][42] ) );
  MUX2_X2 M1_2_41 ( .A(\ML_int[2][41] ), .B(\ML_int[2][37] ), .S(n7), .Z(
        \ML_int[3][41] ) );
  MUX2_X2 M1_2_40 ( .A(\ML_int[2][40] ), .B(\ML_int[2][36] ), .S(n7), .Z(
        \ML_int[3][40] ) );
  MUX2_X2 M1_2_39 ( .A(\ML_int[2][39] ), .B(\ML_int[2][35] ), .S(n7), .Z(
        \ML_int[3][39] ) );
  MUX2_X2 M1_2_38 ( .A(\ML_int[2][38] ), .B(\ML_int[2][34] ), .S(n7), .Z(
        \ML_int[3][38] ) );
  MUX2_X2 M1_2_37 ( .A(\ML_int[2][37] ), .B(\ML_int[2][33] ), .S(n7), .Z(
        \ML_int[3][37] ) );
  MUX2_X2 M1_2_36 ( .A(\ML_int[2][36] ), .B(\ML_int[2][32] ), .S(n7), .Z(
        \ML_int[3][36] ) );
  MUX2_X2 M1_2_35 ( .A(\ML_int[2][35] ), .B(\ML_int[2][31] ), .S(n7), .Z(
        \ML_int[3][35] ) );
  MUX2_X2 M1_2_34 ( .A(\ML_int[2][34] ), .B(\ML_int[2][30] ), .S(n7), .Z(
        \ML_int[3][34] ) );
  MUX2_X2 M1_2_33 ( .A(\ML_int[2][33] ), .B(\ML_int[2][29] ), .S(n7), .Z(
        \ML_int[3][33] ) );
  MUX2_X2 M1_2_32 ( .A(\ML_int[2][32] ), .B(\ML_int[2][28] ), .S(n7), .Z(
        \ML_int[3][32] ) );
  MUX2_X2 M1_2_31 ( .A(\ML_int[2][31] ), .B(\ML_int[2][27] ), .S(n7), .Z(
        \ML_int[3][31] ) );
  MUX2_X2 M1_2_30 ( .A(\ML_int[2][30] ), .B(\ML_int[2][26] ), .S(n7), .Z(
        \ML_int[3][30] ) );
  MUX2_X2 M1_2_29 ( .A(\ML_int[2][29] ), .B(\ML_int[2][25] ), .S(n7), .Z(
        \ML_int[3][29] ) );
  MUX2_X2 M1_2_28 ( .A(\ML_int[2][28] ), .B(\ML_int[2][24] ), .S(n7), .Z(
        \ML_int[3][28] ) );
  MUX2_X2 M1_2_27 ( .A(\ML_int[2][27] ), .B(\ML_int[2][23] ), .S(n7), .Z(
        \ML_int[3][27] ) );
  MUX2_X2 M1_2_26 ( .A(\ML_int[2][26] ), .B(\ML_int[2][22] ), .S(n7), .Z(
        \ML_int[3][26] ) );
  MUX2_X2 M1_2_25 ( .A(\ML_int[2][25] ), .B(\ML_int[2][21] ), .S(SH[2]), .Z(
        \ML_int[3][25] ) );
  MUX2_X2 M1_2_24 ( .A(\ML_int[2][24] ), .B(\ML_int[2][20] ), .S(SH[2]), .Z(
        \ML_int[3][24] ) );
  MUX2_X2 M1_2_23 ( .A(\ML_int[2][23] ), .B(\ML_int[2][19] ), .S(SH[2]), .Z(
        \ML_int[3][23] ) );
  MUX2_X2 M1_2_22 ( .A(\ML_int[2][22] ), .B(\ML_int[2][18] ), .S(SH[2]), .Z(
        \ML_int[3][22] ) );
  MUX2_X2 M1_2_21 ( .A(\ML_int[2][21] ), .B(\ML_int[2][17] ), .S(SH[2]), .Z(
        \ML_int[3][21] ) );
  MUX2_X2 M1_2_20 ( .A(\ML_int[2][20] ), .B(\ML_int[2][16] ), .S(SH[2]), .Z(
        \ML_int[3][20] ) );
  MUX2_X2 M1_2_19 ( .A(\ML_int[2][19] ), .B(\ML_int[2][15] ), .S(SH[2]), .Z(
        \ML_int[3][19] ) );
  MUX2_X2 M1_2_18 ( .A(\ML_int[2][18] ), .B(\ML_int[2][14] ), .S(SH[2]), .Z(
        \ML_int[3][18] ) );
  MUX2_X2 M1_2_17 ( .A(\ML_int[2][17] ), .B(\ML_int[2][13] ), .S(SH[2]), .Z(
        \ML_int[3][17] ) );
  MUX2_X2 M1_2_16 ( .A(\ML_int[2][16] ), .B(\ML_int[2][12] ), .S(SH[2]), .Z(
        \ML_int[3][16] ) );
  MUX2_X2 M1_2_15 ( .A(\ML_int[2][15] ), .B(\ML_int[2][11] ), .S(SH[2]), .Z(
        \ML_int[3][15] ) );
  MUX2_X2 M1_2_14 ( .A(\ML_int[2][14] ), .B(\ML_int[2][10] ), .S(SH[2]), .Z(
        \ML_int[3][14] ) );
  MUX2_X2 M1_2_13 ( .A(\ML_int[2][13] ), .B(\ML_int[2][9] ), .S(SH[2]), .Z(
        \ML_int[3][13] ) );
  MUX2_X2 M1_2_12 ( .A(\ML_int[2][12] ), .B(\ML_int[2][8] ), .S(SH[2]), .Z(
        \ML_int[3][12] ) );
  MUX2_X2 M1_2_11 ( .A(\ML_int[2][11] ), .B(\ML_int[2][7] ), .S(SH[2]), .Z(
        \ML_int[3][11] ) );
  MUX2_X2 M1_2_10 ( .A(\ML_int[2][10] ), .B(\ML_int[2][6] ), .S(SH[2]), .Z(
        \ML_int[3][10] ) );
  MUX2_X2 M1_2_9 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S(SH[2]), .Z(
        \ML_int[3][9] ) );
  MUX2_X2 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(SH[2]), .Z(
        \ML_int[3][8] ) );
  MUX2_X2 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(SH[2]), .Z(
        \ML_int[3][7] ) );
  MUX2_X2 M1_2_6 ( .A(\ML_int[2][6] ), .B(\ML_int[2][2] ), .S(SH[2]), .Z(
        \ML_int[3][6] ) );
  MUX2_X2 M1_2_5 ( .A(\ML_int[2][5] ), .B(\ML_int[2][1] ), .S(SH[2]), .Z(
        \ML_int[3][5] ) );
  MUX2_X2 M1_2_4 ( .A(\ML_int[2][4] ), .B(\ML_int[2][0] ), .S(SH[2]), .Z(
        \ML_int[3][4] ) );
  MUX2_X2 M1_1_52 ( .A(\ML_int[1][52] ), .B(\ML_int[1][50] ), .S(n4), .Z(
        \ML_int[2][52] ) );
  MUX2_X2 M1_1_51 ( .A(\ML_int[1][51] ), .B(\ML_int[1][49] ), .S(n4), .Z(
        \ML_int[2][51] ) );
  MUX2_X2 M1_1_50 ( .A(\ML_int[1][50] ), .B(\ML_int[1][48] ), .S(n4), .Z(
        \ML_int[2][50] ) );
  MUX2_X2 M1_1_49 ( .A(\ML_int[1][49] ), .B(\ML_int[1][47] ), .S(n4), .Z(
        \ML_int[2][49] ) );
  MUX2_X2 M1_1_48 ( .A(\ML_int[1][48] ), .B(\ML_int[1][46] ), .S(SH[1]), .Z(
        \ML_int[2][48] ) );
  MUX2_X2 M1_1_47 ( .A(\ML_int[1][47] ), .B(\ML_int[1][45] ), .S(SH[1]), .Z(
        \ML_int[2][47] ) );
  MUX2_X2 M1_1_46 ( .A(\ML_int[1][46] ), .B(\ML_int[1][44] ), .S(SH[1]), .Z(
        \ML_int[2][46] ) );
  MUX2_X2 M1_1_45 ( .A(\ML_int[1][45] ), .B(\ML_int[1][43] ), .S(SH[1]), .Z(
        \ML_int[2][45] ) );
  MUX2_X2 M1_1_44 ( .A(\ML_int[1][44] ), .B(\ML_int[1][42] ), .S(SH[1]), .Z(
        \ML_int[2][44] ) );
  MUX2_X2 M1_1_43 ( .A(\ML_int[1][43] ), .B(\ML_int[1][41] ), .S(SH[1]), .Z(
        \ML_int[2][43] ) );
  MUX2_X2 M1_1_42 ( .A(\ML_int[1][42] ), .B(\ML_int[1][40] ), .S(SH[1]), .Z(
        \ML_int[2][42] ) );
  MUX2_X2 M1_1_41 ( .A(\ML_int[1][41] ), .B(\ML_int[1][39] ), .S(SH[1]), .Z(
        \ML_int[2][41] ) );
  MUX2_X2 M1_1_40 ( .A(\ML_int[1][40] ), .B(\ML_int[1][38] ), .S(SH[1]), .Z(
        \ML_int[2][40] ) );
  MUX2_X2 M1_1_39 ( .A(\ML_int[1][39] ), .B(\ML_int[1][37] ), .S(SH[1]), .Z(
        \ML_int[2][39] ) );
  MUX2_X2 M1_1_38 ( .A(\ML_int[1][38] ), .B(\ML_int[1][36] ), .S(SH[1]), .Z(
        \ML_int[2][38] ) );
  MUX2_X2 M1_1_37 ( .A(\ML_int[1][37] ), .B(\ML_int[1][35] ), .S(SH[1]), .Z(
        \ML_int[2][37] ) );
  MUX2_X2 M1_1_36 ( .A(\ML_int[1][36] ), .B(\ML_int[1][34] ), .S(SH[1]), .Z(
        \ML_int[2][36] ) );
  MUX2_X2 M1_1_35 ( .A(\ML_int[1][35] ), .B(\ML_int[1][33] ), .S(SH[1]), .Z(
        \ML_int[2][35] ) );
  MUX2_X2 M1_1_34 ( .A(\ML_int[1][34] ), .B(\ML_int[1][32] ), .S(SH[1]), .Z(
        \ML_int[2][34] ) );
  MUX2_X2 M1_1_33 ( .A(\ML_int[1][33] ), .B(\ML_int[1][31] ), .S(SH[1]), .Z(
        \ML_int[2][33] ) );
  MUX2_X2 M1_1_32 ( .A(\ML_int[1][32] ), .B(\ML_int[1][30] ), .S(SH[1]), .Z(
        \ML_int[2][32] ) );
  MUX2_X2 M1_1_31 ( .A(\ML_int[1][31] ), .B(\ML_int[1][29] ), .S(SH[1]), .Z(
        \ML_int[2][31] ) );
  MUX2_X2 M1_1_30 ( .A(\ML_int[1][30] ), .B(\ML_int[1][28] ), .S(SH[1]), .Z(
        \ML_int[2][30] ) );
  MUX2_X2 M1_1_29 ( .A(\ML_int[1][29] ), .B(\ML_int[1][27] ), .S(SH[1]), .Z(
        \ML_int[2][29] ) );
  MUX2_X2 M1_1_28 ( .A(\ML_int[1][28] ), .B(\ML_int[1][26] ), .S(n4), .Z(
        \ML_int[2][28] ) );
  MUX2_X2 M1_1_27 ( .A(\ML_int[1][27] ), .B(\ML_int[1][25] ), .S(n4), .Z(
        \ML_int[2][27] ) );
  MUX2_X2 M1_1_26 ( .A(\ML_int[1][26] ), .B(\ML_int[1][24] ), .S(SH[1]), .Z(
        \ML_int[2][26] ) );
  MUX2_X2 M1_1_25 ( .A(\ML_int[1][25] ), .B(\ML_int[1][23] ), .S(SH[1]), .Z(
        \ML_int[2][25] ) );
  MUX2_X2 M1_1_24 ( .A(\ML_int[1][24] ), .B(\ML_int[1][22] ), .S(SH[1]), .Z(
        \ML_int[2][24] ) );
  MUX2_X2 M1_1_23 ( .A(\ML_int[1][23] ), .B(\ML_int[1][21] ), .S(n6), .Z(
        \ML_int[2][23] ) );
  MUX2_X2 M1_1_22 ( .A(\ML_int[1][22] ), .B(\ML_int[1][20] ), .S(n6), .Z(
        \ML_int[2][22] ) );
  MUX2_X2 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S(n6), .Z(
        \ML_int[2][21] ) );
  MUX2_X2 M1_1_20 ( .A(\ML_int[1][20] ), .B(\ML_int[1][18] ), .S(n6), .Z(
        \ML_int[2][20] ) );
  MUX2_X2 M1_1_19 ( .A(\ML_int[1][19] ), .B(\ML_int[1][17] ), .S(n6), .Z(
        \ML_int[2][19] ) );
  MUX2_X2 M1_1_18 ( .A(\ML_int[1][18] ), .B(\ML_int[1][16] ), .S(n6), .Z(
        \ML_int[2][18] ) );
  MUX2_X2 M1_1_17 ( .A(\ML_int[1][17] ), .B(\ML_int[1][15] ), .S(n6), .Z(
        \ML_int[2][17] ) );
  MUX2_X2 M1_1_16 ( .A(\ML_int[1][16] ), .B(\ML_int[1][14] ), .S(n6), .Z(
        \ML_int[2][16] ) );
  MUX2_X2 M1_1_15 ( .A(\ML_int[1][15] ), .B(\ML_int[1][13] ), .S(n6), .Z(
        \ML_int[2][15] ) );
  MUX2_X2 M1_1_14 ( .A(\ML_int[1][14] ), .B(\ML_int[1][12] ), .S(n6), .Z(
        \ML_int[2][14] ) );
  MUX2_X2 M1_1_13 ( .A(\ML_int[1][13] ), .B(\ML_int[1][11] ), .S(n6), .Z(
        \ML_int[2][13] ) );
  MUX2_X2 M1_1_12 ( .A(\ML_int[1][12] ), .B(\ML_int[1][10] ), .S(n6), .Z(
        \ML_int[2][12] ) );
  MUX2_X2 M1_1_11 ( .A(\ML_int[1][11] ), .B(\ML_int[1][9] ), .S(n6), .Z(
        \ML_int[2][11] ) );
  MUX2_X2 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S(n6), .Z(
        \ML_int[2][10] ) );
  MUX2_X2 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S(n6), .Z(
        \ML_int[2][9] ) );
  MUX2_X2 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S(n6), .Z(
        \ML_int[2][8] ) );
  MUX2_X2 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S(n6), .Z(
        \ML_int[2][7] ) );
  MUX2_X2 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S(n6), .Z(
        \ML_int[2][6] ) );
  MUX2_X2 M1_1_5 ( .A(\ML_int[1][5] ), .B(\ML_int[1][3] ), .S(n6), .Z(
        \ML_int[2][5] ) );
  MUX2_X2 M1_1_4 ( .A(\ML_int[1][4] ), .B(\ML_int[1][2] ), .S(n6), .Z(
        \ML_int[2][4] ) );
  MUX2_X2 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(n6), .Z(
        \ML_int[2][3] ) );
  MUX2_X2 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S(n6), .Z(
        \ML_int[2][2] ) );
  MUX2_X2 M1_0_52 ( .A(A[52]), .B(A[51]), .S(n1), .Z(\ML_int[1][52] ) );
  MUX2_X2 M1_0_51 ( .A(A[51]), .B(A[50]), .S(n1), .Z(\ML_int[1][51] ) );
  MUX2_X2 M1_0_50 ( .A(A[50]), .B(A[49]), .S(n1), .Z(\ML_int[1][50] ) );
  MUX2_X2 M1_0_49 ( .A(A[49]), .B(A[48]), .S(n1), .Z(\ML_int[1][49] ) );
  MUX2_X2 M1_0_48 ( .A(A[48]), .B(A[47]), .S(n1), .Z(\ML_int[1][48] ) );
  MUX2_X2 M1_0_47 ( .A(A[47]), .B(A[46]), .S(SH[0]), .Z(\ML_int[1][47] ) );
  MUX2_X2 M1_0_46 ( .A(A[46]), .B(A[45]), .S(SH[0]), .Z(\ML_int[1][46] ) );
  MUX2_X2 M1_0_45 ( .A(A[45]), .B(A[44]), .S(SH[0]), .Z(\ML_int[1][45] ) );
  MUX2_X2 M1_0_44 ( .A(A[44]), .B(A[43]), .S(SH[0]), .Z(\ML_int[1][44] ) );
  MUX2_X2 M1_0_43 ( .A(A[43]), .B(A[42]), .S(SH[0]), .Z(\ML_int[1][43] ) );
  MUX2_X2 M1_0_42 ( .A(A[42]), .B(A[41]), .S(SH[0]), .Z(\ML_int[1][42] ) );
  MUX2_X2 M1_0_41 ( .A(A[41]), .B(A[40]), .S(SH[0]), .Z(\ML_int[1][41] ) );
  MUX2_X2 M1_0_40 ( .A(A[40]), .B(A[39]), .S(SH[0]), .Z(\ML_int[1][40] ) );
  MUX2_X2 M1_0_39 ( .A(A[39]), .B(A[38]), .S(SH[0]), .Z(\ML_int[1][39] ) );
  MUX2_X2 M1_0_38 ( .A(A[38]), .B(A[37]), .S(SH[0]), .Z(\ML_int[1][38] ) );
  MUX2_X2 M1_0_37 ( .A(A[37]), .B(A[36]), .S(SH[0]), .Z(\ML_int[1][37] ) );
  MUX2_X2 M1_0_36 ( .A(A[36]), .B(A[35]), .S(SH[0]), .Z(\ML_int[1][36] ) );
  MUX2_X2 M1_0_35 ( .A(A[35]), .B(A[34]), .S(SH[0]), .Z(\ML_int[1][35] ) );
  MUX2_X2 M1_0_34 ( .A(A[34]), .B(A[33]), .S(SH[0]), .Z(\ML_int[1][34] ) );
  MUX2_X2 M1_0_33 ( .A(A[33]), .B(A[32]), .S(SH[0]), .Z(\ML_int[1][33] ) );
  MUX2_X2 M1_0_32 ( .A(A[32]), .B(A[31]), .S(SH[0]), .Z(\ML_int[1][32] ) );
  MUX2_X2 M1_0_31 ( .A(A[31]), .B(A[30]), .S(SH[0]), .Z(\ML_int[1][31] ) );
  MUX2_X2 M1_0_30 ( .A(A[30]), .B(A[29]), .S(SH[0]), .Z(\ML_int[1][30] ) );
  MUX2_X2 M1_0_29 ( .A(A[29]), .B(A[28]), .S(SH[0]), .Z(\ML_int[1][29] ) );
  MUX2_X2 M1_0_28 ( .A(A[28]), .B(A[27]), .S(SH[0]), .Z(\ML_int[1][28] ) );
  MUX2_X2 M1_0_27 ( .A(A[27]), .B(A[26]), .S(SH[0]), .Z(\ML_int[1][27] ) );
  MUX2_X2 M1_0_26 ( .A(A[26]), .B(A[25]), .S(n1), .Z(\ML_int[1][26] ) );
  MUX2_X2 M1_0_25 ( .A(A[25]), .B(A[24]), .S(n1), .Z(\ML_int[1][25] ) );
  MUX2_X2 M1_0_24 ( .A(A[24]), .B(A[23]), .S(SH[0]), .Z(\ML_int[1][24] ) );
  MUX2_X2 M1_0_23 ( .A(A[23]), .B(A[22]), .S(SH[0]), .Z(\ML_int[1][23] ) );
  MUX2_X2 M1_0_22 ( .A(A[22]), .B(A[21]), .S(n3), .Z(\ML_int[1][22] ) );
  MUX2_X2 M1_0_21 ( .A(A[21]), .B(A[20]), .S(n3), .Z(\ML_int[1][21] ) );
  MUX2_X2 M1_0_20 ( .A(A[20]), .B(A[19]), .S(n3), .Z(\ML_int[1][20] ) );
  MUX2_X2 M1_0_19 ( .A(A[19]), .B(A[18]), .S(n3), .Z(\ML_int[1][19] ) );
  MUX2_X2 M1_0_18 ( .A(A[18]), .B(A[17]), .S(n3), .Z(\ML_int[1][18] ) );
  MUX2_X2 M1_0_17 ( .A(A[17]), .B(A[16]), .S(n3), .Z(\ML_int[1][17] ) );
  MUX2_X2 M1_0_16 ( .A(A[16]), .B(A[15]), .S(n3), .Z(\ML_int[1][16] ) );
  MUX2_X2 M1_0_15 ( .A(A[15]), .B(A[14]), .S(n3), .Z(\ML_int[1][15] ) );
  MUX2_X2 M1_0_14 ( .A(A[14]), .B(A[13]), .S(n3), .Z(\ML_int[1][14] ) );
  MUX2_X2 M1_0_13 ( .A(A[13]), .B(A[12]), .S(n3), .Z(\ML_int[1][13] ) );
  MUX2_X2 M1_0_12 ( .A(A[12]), .B(A[11]), .S(n3), .Z(\ML_int[1][12] ) );
  MUX2_X2 M1_0_11 ( .A(A[11]), .B(A[10]), .S(n3), .Z(\ML_int[1][11] ) );
  MUX2_X2 M1_0_10 ( .A(A[10]), .B(A[9]), .S(n3), .Z(\ML_int[1][10] ) );
  MUX2_X2 M1_0_9 ( .A(A[9]), .B(A[8]), .S(n3), .Z(\ML_int[1][9] ) );
  MUX2_X2 M1_0_8 ( .A(A[8]), .B(A[7]), .S(n3), .Z(\ML_int[1][8] ) );
  MUX2_X2 M1_0_7 ( .A(A[7]), .B(A[6]), .S(n3), .Z(\ML_int[1][7] ) );
  MUX2_X2 M1_0_6 ( .A(A[6]), .B(A[5]), .S(n3), .Z(\ML_int[1][6] ) );
  MUX2_X2 M1_0_5 ( .A(A[5]), .B(A[4]), .S(n3), .Z(\ML_int[1][5] ) );
  MUX2_X2 M1_0_4 ( .A(A[4]), .B(A[3]), .S(n3), .Z(\ML_int[1][4] ) );
  MUX2_X2 M1_0_3 ( .A(A[3]), .B(A[2]), .S(n3), .Z(\ML_int[1][3] ) );
  MUX2_X2 M1_0_2 ( .A(A[2]), .B(A[1]), .S(n3), .Z(\ML_int[1][2] ) );
  MUX2_X2 M1_0_1 ( .A(A[1]), .B(A[0]), .S(n3), .Z(\ML_int[1][1] ) );
  INV_X4 U3 ( .A(SH[3]), .ZN(n10) );
  INV_X4 U4 ( .A(SH[2]), .ZN(n8) );
  INV_X4 U5 ( .A(n5), .ZN(n6) );
  INV_X4 U6 ( .A(n2), .ZN(n3) );
  INV_X4 U7 ( .A(SH[4]), .ZN(n12) );
  INV_X4 U8 ( .A(n2), .ZN(n1) );
  INV_X4 U9 ( .A(SH[0]), .ZN(n2) );
  INV_X4 U10 ( .A(n5), .ZN(n4) );
  INV_X4 U11 ( .A(SH[1]), .ZN(n5) );
  INV_X4 U12 ( .A(n8), .ZN(n7) );
  INV_X4 U13 ( .A(n12), .ZN(n11) );
  INV_X4 U14 ( .A(n12), .ZN(n14) );
  INV_X4 U15 ( .A(n12), .ZN(n13) );
  INV_X4 U16 ( .A(n10), .ZN(n9) );
  INV_X4 U17 ( .A(n27), .ZN(n15) );
  INV_X4 U18 ( .A(n28), .ZN(n16) );
  INV_X4 U19 ( .A(n29), .ZN(n17) );
  INV_X4 U20 ( .A(n30), .ZN(n18) );
  INV_X4 U21 ( .A(n26), .ZN(n19) );
  INV_X4 U22 ( .A(n25), .ZN(n20) );
  INV_X4 U23 ( .A(n24), .ZN(n21) );
  INV_X4 U24 ( .A(n23), .ZN(n22) );
  AND2_X1 U25 ( .A1(\ML_int[4][9] ), .A2(n12), .ZN(\ML_int[5][9] ) );
  AND2_X1 U26 ( .A1(\ML_int[4][8] ), .A2(n12), .ZN(\ML_int[5][8] ) );
  NOR2_X1 U27 ( .A1(n11), .A2(n23), .ZN(\ML_int[5][7] ) );
  NOR2_X1 U28 ( .A1(n11), .A2(n24), .ZN(\ML_int[5][6] ) );
  NOR2_X1 U29 ( .A1(n11), .A2(n25), .ZN(\ML_int[5][5] ) );
  NOR2_X1 U30 ( .A1(n11), .A2(n26), .ZN(\ML_int[5][4] ) );
  NOR2_X1 U31 ( .A1(n11), .A2(n27), .ZN(\ML_int[5][3] ) );
  NOR2_X1 U32 ( .A1(n14), .A2(n28), .ZN(\ML_int[5][2] ) );
  NOR2_X1 U33 ( .A1(n13), .A2(n29), .ZN(\ML_int[5][1] ) );
  AND2_X1 U34 ( .A1(\ML_int[4][15] ), .A2(n12), .ZN(\ML_int[5][15] ) );
  AND2_X1 U35 ( .A1(\ML_int[4][14] ), .A2(n12), .ZN(\ML_int[5][14] ) );
  AND2_X1 U36 ( .A1(\ML_int[4][13] ), .A2(n12), .ZN(\ML_int[5][13] ) );
  AND2_X1 U37 ( .A1(\ML_int[4][12] ), .A2(n12), .ZN(\ML_int[5][12] ) );
  AND2_X1 U38 ( .A1(\ML_int[4][11] ), .A2(n12), .ZN(\ML_int[5][11] ) );
  AND2_X1 U39 ( .A1(\ML_int[4][10] ), .A2(n12), .ZN(\ML_int[5][10] ) );
  NOR2_X1 U40 ( .A1(SH[4]), .A2(n30), .ZN(\ML_int[5][0] ) );
  NAND2_X1 U41 ( .A1(\ML_int[3][7] ), .A2(n10), .ZN(n23) );
  NAND2_X1 U42 ( .A1(\ML_int[3][6] ), .A2(n10), .ZN(n24) );
  NAND2_X1 U43 ( .A1(\ML_int[3][5] ), .A2(n10), .ZN(n25) );
  NAND2_X1 U44 ( .A1(\ML_int[3][4] ), .A2(n10), .ZN(n26) );
  NAND2_X1 U45 ( .A1(\ML_int[3][3] ), .A2(n10), .ZN(n27) );
  NAND2_X1 U46 ( .A1(\ML_int[3][2] ), .A2(n10), .ZN(n28) );
  NAND2_X1 U47 ( .A1(\ML_int[3][1] ), .A2(n10), .ZN(n29) );
  NAND2_X1 U48 ( .A1(\ML_int[3][0] ), .A2(n10), .ZN(n30) );
  AND2_X1 U49 ( .A1(\ML_int[2][3] ), .A2(n8), .ZN(\ML_int[3][3] ) );
  AND2_X1 U50 ( .A1(\ML_int[2][2] ), .A2(n8), .ZN(\ML_int[3][2] ) );
  AND2_X1 U51 ( .A1(\ML_int[2][1] ), .A2(n8), .ZN(\ML_int[3][1] ) );
  AND2_X1 U52 ( .A1(\ML_int[2][0] ), .A2(n8), .ZN(\ML_int[3][0] ) );
  AND2_X1 U53 ( .A1(\ML_int[1][1] ), .A2(n5), .ZN(\ML_int[2][1] ) );
  AND2_X1 U54 ( .A1(\ML_int[1][0] ), .A2(n5), .ZN(\ML_int[2][0] ) );
  AND2_X1 U55 ( .A1(A[0]), .A2(n2), .ZN(\ML_int[1][0] ) );
endmodule


module fpu_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [51:0] A;
  input [51:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178;

  INV_X4 U1 ( .A(A[50]), .ZN(n1) );
  INV_X4 U2 ( .A(n87), .ZN(n2) );
  INV_X4 U3 ( .A(n88), .ZN(n3) );
  INV_X4 U4 ( .A(A[1]), .ZN(n4) );
  INV_X4 U5 ( .A(n165), .ZN(n5) );
  INV_X4 U6 ( .A(B[51]), .ZN(n6) );
  INV_X4 U7 ( .A(B[49]), .ZN(n7) );
  INV_X4 U8 ( .A(B[48]), .ZN(n8) );
  INV_X4 U9 ( .A(B[47]), .ZN(n9) );
  INV_X4 U10 ( .A(B[46]), .ZN(n10) );
  INV_X4 U11 ( .A(B[45]), .ZN(n11) );
  INV_X4 U12 ( .A(B[44]), .ZN(n12) );
  INV_X4 U13 ( .A(B[43]), .ZN(n13) );
  INV_X4 U14 ( .A(B[42]), .ZN(n14) );
  INV_X4 U15 ( .A(B[41]), .ZN(n15) );
  INV_X4 U16 ( .A(B[40]), .ZN(n16) );
  INV_X4 U17 ( .A(B[39]), .ZN(n17) );
  INV_X4 U18 ( .A(B[38]), .ZN(n18) );
  INV_X4 U19 ( .A(B[37]), .ZN(n19) );
  INV_X4 U20 ( .A(B[36]), .ZN(n20) );
  INV_X4 U21 ( .A(B[35]), .ZN(n21) );
  INV_X4 U22 ( .A(B[34]), .ZN(n22) );
  INV_X4 U23 ( .A(B[33]), .ZN(n23) );
  INV_X4 U24 ( .A(B[32]), .ZN(n24) );
  INV_X4 U25 ( .A(B[31]), .ZN(n25) );
  INV_X4 U26 ( .A(B[30]), .ZN(n26) );
  INV_X4 U27 ( .A(B[29]), .ZN(n27) );
  INV_X4 U28 ( .A(B[28]), .ZN(n28) );
  INV_X4 U29 ( .A(B[27]), .ZN(n29) );
  INV_X4 U30 ( .A(B[26]), .ZN(n30) );
  INV_X4 U31 ( .A(B[25]), .ZN(n31) );
  INV_X4 U32 ( .A(B[24]), .ZN(n32) );
  INV_X4 U33 ( .A(B[23]), .ZN(n33) );
  INV_X4 U34 ( .A(B[22]), .ZN(n34) );
  INV_X4 U35 ( .A(B[21]), .ZN(n35) );
  INV_X4 U36 ( .A(B[20]), .ZN(n36) );
  INV_X4 U37 ( .A(B[19]), .ZN(n37) );
  INV_X4 U38 ( .A(B[18]), .ZN(n38) );
  INV_X4 U39 ( .A(B[17]), .ZN(n39) );
  INV_X4 U40 ( .A(B[16]), .ZN(n40) );
  INV_X4 U41 ( .A(B[15]), .ZN(n41) );
  INV_X4 U42 ( .A(B[14]), .ZN(n42) );
  INV_X4 U43 ( .A(B[13]), .ZN(n43) );
  INV_X4 U44 ( .A(B[12]), .ZN(n44) );
  INV_X4 U45 ( .A(B[11]), .ZN(n45) );
  INV_X4 U46 ( .A(B[10]), .ZN(n46) );
  INV_X4 U47 ( .A(B[9]), .ZN(n47) );
  INV_X4 U48 ( .A(B[8]), .ZN(n48) );
  INV_X4 U49 ( .A(B[7]), .ZN(n49) );
  INV_X4 U50 ( .A(B[6]), .ZN(n50) );
  INV_X4 U51 ( .A(B[5]), .ZN(n51) );
  INV_X4 U52 ( .A(B[4]), .ZN(n52) );
  INV_X4 U53 ( .A(B[3]), .ZN(n53) );
  INV_X4 U54 ( .A(B[2]), .ZN(n54) );
  INV_X4 U55 ( .A(B[1]), .ZN(n55) );
  INV_X4 U56 ( .A(B[0]), .ZN(n56) );
  NOR4_X1 U57 ( .A1(n57), .A2(n58), .A3(n59), .A4(n60), .ZN(EQ) );
  NAND4_X1 U58 ( .A1(n61), .A2(n62), .A3(n63), .A4(n64), .ZN(n60) );
  AND3_X1 U59 ( .A1(n65), .A2(n66), .A3(n67), .ZN(n64) );
  NAND4_X1 U60 ( .A1(n68), .A2(n69), .A3(n70), .A4(n71), .ZN(n59) );
  AND4_X1 U61 ( .A1(n72), .A2(n73), .A3(n74), .A4(n75), .ZN(n71) );
  NAND3_X1 U62 ( .A1(n76), .A2(n77), .A3(n78), .ZN(n58) );
  AND4_X1 U63 ( .A1(n79), .A2(n80), .A3(n81), .A4(n82), .ZN(n78) );
  AND3_X1 U64 ( .A1(n83), .A2(n84), .A3(n85), .ZN(n79) );
  NOR4_X1 U65 ( .A1(LT), .A2(n86), .A3(n3), .A4(n2), .ZN(n77) );
  OAI22_X1 U66 ( .A1(A[51]), .A2(n6), .B1(n86), .B2(n89), .ZN(LT) );
  AOI22_X1 U67 ( .A1(B[50]), .A2(n1), .B1(n90), .B2(n91), .ZN(n89) );
  OAI221_X1 U68 ( .B1(A[48]), .B2(n8), .C1(A[49]), .C2(n7), .A(n92), .ZN(n91)
         );
  NAND3_X1 U69 ( .A1(n93), .A2(n94), .A3(n95), .ZN(n92) );
  OAI221_X1 U70 ( .B1(A[46]), .B2(n10), .C1(A[47]), .C2(n9), .A(n96), .ZN(n95)
         );
  NAND3_X1 U71 ( .A1(n97), .A2(n98), .A3(n99), .ZN(n96) );
  OAI221_X1 U72 ( .B1(A[44]), .B2(n12), .C1(A[45]), .C2(n11), .A(n100), .ZN(
        n99) );
  NAND3_X1 U73 ( .A1(n101), .A2(n102), .A3(n103), .ZN(n100) );
  OAI221_X1 U74 ( .B1(A[42]), .B2(n14), .C1(A[43]), .C2(n13), .A(n104), .ZN(
        n103) );
  NAND3_X1 U75 ( .A1(n105), .A2(n106), .A3(n107), .ZN(n104) );
  OAI221_X1 U76 ( .B1(A[40]), .B2(n16), .C1(A[41]), .C2(n15), .A(n108), .ZN(
        n107) );
  NAND3_X1 U77 ( .A1(n109), .A2(n110), .A3(n111), .ZN(n108) );
  OAI221_X1 U78 ( .B1(A[38]), .B2(n18), .C1(A[39]), .C2(n17), .A(n112), .ZN(
        n111) );
  NAND3_X1 U79 ( .A1(n113), .A2(n114), .A3(n115), .ZN(n112) );
  OAI221_X1 U80 ( .B1(A[36]), .B2(n20), .C1(A[37]), .C2(n19), .A(n116), .ZN(
        n115) );
  NAND3_X1 U81 ( .A1(n117), .A2(n118), .A3(n119), .ZN(n116) );
  OAI221_X1 U82 ( .B1(A[34]), .B2(n22), .C1(A[35]), .C2(n21), .A(n120), .ZN(
        n119) );
  NAND3_X1 U83 ( .A1(n121), .A2(n122), .A3(n123), .ZN(n120) );
  OAI221_X1 U84 ( .B1(A[32]), .B2(n24), .C1(A[33]), .C2(n23), .A(n124), .ZN(
        n123) );
  NAND3_X1 U85 ( .A1(n125), .A2(n126), .A3(n127), .ZN(n124) );
  OAI221_X1 U86 ( .B1(A[30]), .B2(n26), .C1(A[31]), .C2(n25), .A(n128), .ZN(
        n127) );
  NAND3_X1 U87 ( .A1(n129), .A2(n130), .A3(n131), .ZN(n128) );
  OAI221_X1 U88 ( .B1(A[28]), .B2(n28), .C1(A[29]), .C2(n27), .A(n132), .ZN(
        n131) );
  NAND3_X1 U89 ( .A1(n133), .A2(n134), .A3(n135), .ZN(n132) );
  OAI221_X1 U90 ( .B1(A[26]), .B2(n30), .C1(A[27]), .C2(n29), .A(n136), .ZN(
        n135) );
  NAND3_X1 U91 ( .A1(n137), .A2(n63), .A3(n138), .ZN(n136) );
  OAI221_X1 U92 ( .B1(A[24]), .B2(n32), .C1(A[25]), .C2(n31), .A(n139), .ZN(
        n138) );
  NAND3_X1 U93 ( .A1(n61), .A2(n62), .A3(n140), .ZN(n139) );
  OAI221_X1 U94 ( .B1(A[22]), .B2(n34), .C1(A[23]), .C2(n33), .A(n141), .ZN(
        n140) );
  NAND3_X1 U95 ( .A1(n65), .A2(n67), .A3(n142), .ZN(n141) );
  OAI221_X1 U96 ( .B1(A[20]), .B2(n36), .C1(A[21]), .C2(n35), .A(n143), .ZN(
        n142) );
  NAND3_X1 U97 ( .A1(n66), .A2(n70), .A3(n144), .ZN(n143) );
  OAI221_X1 U98 ( .B1(A[18]), .B2(n38), .C1(A[19]), .C2(n37), .A(n145), .ZN(
        n144) );
  NAND3_X1 U99 ( .A1(n68), .A2(n69), .A3(n146), .ZN(n145) );
  OAI221_X1 U100 ( .B1(A[16]), .B2(n40), .C1(A[17]), .C2(n39), .A(n147), .ZN(
        n146) );
  NAND3_X1 U101 ( .A1(n75), .A2(n74), .A3(n148), .ZN(n147) );
  OAI221_X1 U102 ( .B1(A[14]), .B2(n42), .C1(A[15]), .C2(n41), .A(n149), .ZN(
        n148) );
  NAND3_X1 U103 ( .A1(n73), .A2(n72), .A3(n150), .ZN(n149) );
  OAI221_X1 U104 ( .B1(A[12]), .B2(n44), .C1(A[13]), .C2(n43), .A(n151), .ZN(
        n150) );
  NAND3_X1 U105 ( .A1(n80), .A2(n82), .A3(n152), .ZN(n151) );
  OAI221_X1 U106 ( .B1(A[10]), .B2(n46), .C1(A[11]), .C2(n45), .A(n153), .ZN(
        n152) );
  NAND3_X1 U107 ( .A1(n81), .A2(n85), .A3(n154), .ZN(n153) );
  OAI221_X1 U108 ( .B1(A[8]), .B2(n48), .C1(A[9]), .C2(n47), .A(n155), .ZN(
        n154) );
  NAND3_X1 U109 ( .A1(n83), .A2(n84), .A3(n156), .ZN(n155) );
  OAI221_X1 U110 ( .B1(A[6]), .B2(n50), .C1(A[7]), .C2(n49), .A(n157), .ZN(
        n156) );
  NAND3_X1 U111 ( .A1(n158), .A2(n159), .A3(n160), .ZN(n157) );
  OAI221_X1 U112 ( .B1(A[4]), .B2(n52), .C1(A[5]), .C2(n51), .A(n161), .ZN(
        n160) );
  NAND3_X1 U113 ( .A1(n162), .A2(n87), .A3(n163), .ZN(n161) );
  OAI221_X1 U114 ( .B1(A[2]), .B2(n54), .C1(A[3]), .C2(n53), .A(n164), .ZN(
        n163) );
  OAI211_X1 U115 ( .C1(n165), .C2(n4), .A(n166), .B(n88), .ZN(n164) );
  NAND2_X1 U116 ( .A1(A[2]), .A2(n54), .ZN(n88) );
  OAI21_X1 U117 ( .B1(A[1]), .B2(n5), .A(n55), .ZN(n166) );
  NOR2_X1 U118 ( .A1(n56), .A2(A[0]), .ZN(n165) );
  NAND2_X1 U119 ( .A1(A[3]), .A2(n53), .ZN(n87) );
  NAND2_X1 U120 ( .A1(A[7]), .A2(n49), .ZN(n84) );
  NAND2_X1 U121 ( .A1(A[8]), .A2(n48), .ZN(n83) );
  NAND2_X1 U122 ( .A1(A[9]), .A2(n47), .ZN(n85) );
  NAND2_X1 U123 ( .A1(A[10]), .A2(n46), .ZN(n81) );
  NAND2_X1 U124 ( .A1(A[11]), .A2(n45), .ZN(n82) );
  NAND2_X1 U125 ( .A1(A[12]), .A2(n44), .ZN(n80) );
  NAND2_X1 U126 ( .A1(A[13]), .A2(n43), .ZN(n72) );
  NAND2_X1 U127 ( .A1(A[14]), .A2(n42), .ZN(n73) );
  NAND2_X1 U128 ( .A1(A[15]), .A2(n41), .ZN(n74) );
  NAND2_X1 U129 ( .A1(A[16]), .A2(n40), .ZN(n75) );
  NAND2_X1 U130 ( .A1(A[17]), .A2(n39), .ZN(n69) );
  NAND2_X1 U131 ( .A1(A[18]), .A2(n38), .ZN(n68) );
  NAND2_X1 U132 ( .A1(A[19]), .A2(n37), .ZN(n70) );
  NAND2_X1 U133 ( .A1(A[20]), .A2(n36), .ZN(n66) );
  NAND2_X1 U134 ( .A1(A[21]), .A2(n35), .ZN(n67) );
  NAND2_X1 U135 ( .A1(A[22]), .A2(n34), .ZN(n65) );
  NAND2_X1 U136 ( .A1(A[23]), .A2(n33), .ZN(n62) );
  NAND2_X1 U137 ( .A1(A[24]), .A2(n32), .ZN(n61) );
  NAND2_X1 U138 ( .A1(A[25]), .A2(n31), .ZN(n63) );
  AND2_X1 U139 ( .A1(n167), .A2(n168), .ZN(n90) );
  AND2_X1 U140 ( .A1(A[51]), .A2(n6), .ZN(n86) );
  AND3_X1 U141 ( .A1(n158), .A2(n162), .A3(n159), .ZN(n76) );
  NAND2_X1 U142 ( .A1(A[5]), .A2(n51), .ZN(n159) );
  NAND2_X1 U143 ( .A1(A[4]), .A2(n52), .ZN(n162) );
  NAND2_X1 U144 ( .A1(A[6]), .A2(n50), .ZN(n158) );
  NAND4_X1 U145 ( .A1(n169), .A2(n170), .A3(n171), .A4(n172), .ZN(n57) );
  AND4_X1 U146 ( .A1(n173), .A2(n125), .A3(n129), .A4(n126), .ZN(n172) );
  NAND2_X1 U147 ( .A1(A[31]), .A2(n25), .ZN(n126) );
  NAND2_X1 U148 ( .A1(A[30]), .A2(n26), .ZN(n129) );
  NAND2_X1 U149 ( .A1(A[32]), .A2(n24), .ZN(n125) );
  AND4_X1 U150 ( .A1(n130), .A2(n133), .A3(n134), .A4(n137), .ZN(n173) );
  NAND2_X1 U151 ( .A1(A[26]), .A2(n30), .ZN(n137) );
  NAND2_X1 U152 ( .A1(A[27]), .A2(n29), .ZN(n134) );
  NAND2_X1 U153 ( .A1(A[28]), .A2(n28), .ZN(n133) );
  NAND2_X1 U154 ( .A1(A[29]), .A2(n27), .ZN(n130) );
  AND4_X1 U155 ( .A1(n174), .A2(n113), .A3(n117), .A4(n114), .ZN(n171) );
  NAND2_X1 U156 ( .A1(A[37]), .A2(n19), .ZN(n114) );
  NAND2_X1 U157 ( .A1(A[36]), .A2(n20), .ZN(n117) );
  NAND2_X1 U158 ( .A1(A[38]), .A2(n18), .ZN(n113) );
  AND3_X1 U159 ( .A1(n121), .A2(n122), .A3(n118), .ZN(n174) );
  NAND2_X1 U160 ( .A1(A[35]), .A2(n21), .ZN(n118) );
  NAND2_X1 U161 ( .A1(A[33]), .A2(n23), .ZN(n122) );
  NAND2_X1 U162 ( .A1(A[34]), .A2(n22), .ZN(n121) );
  AND4_X1 U163 ( .A1(n175), .A2(n98), .A3(n102), .A4(n101), .ZN(n170) );
  NAND2_X1 U164 ( .A1(A[44]), .A2(n12), .ZN(n101) );
  NAND2_X1 U165 ( .A1(A[43]), .A2(n13), .ZN(n102) );
  NAND2_X1 U166 ( .A1(A[45]), .A2(n11), .ZN(n98) );
  AND4_X1 U167 ( .A1(n105), .A2(n106), .A3(n109), .A4(n110), .ZN(n175) );
  NAND2_X1 U168 ( .A1(A[39]), .A2(n17), .ZN(n110) );
  NAND2_X1 U169 ( .A1(A[40]), .A2(n16), .ZN(n109) );
  NAND2_X1 U170 ( .A1(A[41]), .A2(n15), .ZN(n106) );
  NAND2_X1 U171 ( .A1(A[42]), .A2(n14), .ZN(n105) );
  AND4_X1 U172 ( .A1(n176), .A2(n93), .A3(n97), .A4(n94), .ZN(n169) );
  NAND2_X1 U173 ( .A1(A[47]), .A2(n9), .ZN(n94) );
  NAND2_X1 U174 ( .A1(A[46]), .A2(n10), .ZN(n97) );
  NAND2_X1 U175 ( .A1(A[48]), .A2(n8), .ZN(n93) );
  AND3_X1 U176 ( .A1(n168), .A2(n167), .A3(n177), .ZN(n176) );
  OAI22_X1 U177 ( .A1(A[1]), .A2(n178), .B1(n178), .B2(n55), .ZN(n177) );
  AND2_X1 U178 ( .A1(A[0]), .A2(n56), .ZN(n178) );
  OR2_X1 U179 ( .A1(n1), .A2(B[50]), .ZN(n167) );
  NAND2_X1 U180 ( .A1(A[49]), .A2(n7), .ZN(n168) );
endmodule


module fpu_DW01_add_9 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4;
  wire   [8:2] carry;

>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
<<<<<<< HEAD
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  BUF_X32 U1 ( .A(A[0]), .Z(n1) );
  BUF_X32 U2 ( .A(B[0]), .Z(n2) );
  XOR2_X1 U3 ( .A(n2), .B(n1), .Z(SUM[0]) );
  NAND2_X2 U4 ( .A1(B[0]), .A2(A[0]), .ZN(n4) );
  INV_X4 U5 ( .A(n4), .ZN(carry[1]) );
endmodule


module fpu_DW01_ash_2 ( A, DATA_TC, SH, SH_TC, B );
  input [10:0] A;
  input [3:0] SH;
  output [10:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] , \ML_int[1][7] ,
         \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] , \ML_int[1][3] ,
         \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] , \ML_int[2][10] ,
         \ML_int[2][9] , \ML_int[2][8] , \ML_int[2][7] , \ML_int[2][6] ,
         \ML_int[2][5] , \ML_int[2][4] , \ML_int[2][3] , \ML_int[2][2] ,
         \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] , \ML_int[3][7] ,
         \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] , \ML_int[3][2] ,
         \ML_int[3][1] , \ML_int[3][0] , \ML_int[4][10] , \ML_int[4][9] ,
         \ML_int[4][8] , \ML_int[4][7] , \ML_int[4][6] , \ML_int[4][5] ,
         \ML_int[4][4] , \ML_int[4][3] , \ML_int[4][2] , \ML_int[4][1] ,
         \ML_int[4][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;
  assign B[10] = \ML_int[4][10] ;
  assign B[9] = \ML_int[4][9] ;
  assign B[8] = \ML_int[4][8] ;
  assign B[7] = \ML_int[4][7] ;
  assign B[6] = \ML_int[4][6] ;
  assign B[5] = \ML_int[4][5] ;
  assign B[4] = \ML_int[4][4] ;
  assign B[3] = \ML_int[4][3] ;
  assign B[2] = \ML_int[4][2] ;
  assign B[1] = \ML_int[4][1] ;
  assign B[0] = \ML_int[4][0] ;

  MUX2_X2 M1_3_10 ( .A(\ML_int[3][10] ), .B(\ML_int[3][2] ), .S(SH[3]), .Z(
        \ML_int[4][10] ) );
  MUX2_X2 M1_3_9 ( .A(\ML_int[3][9] ), .B(\ML_int[3][1] ), .S(SH[3]), .Z(
        \ML_int[4][9] ) );
  MUX2_X2 M1_3_8 ( .A(\ML_int[3][8] ), .B(\ML_int[3][0] ), .S(SH[3]), .Z(
        \ML_int[4][8] ) );
  MUX2_X2 M1_2_10 ( .A(\ML_int[2][10] ), .B(\ML_int[2][6] ), .S(SH[2]), .Z(
        \ML_int[3][10] ) );
  MUX2_X2 M1_2_9 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S(SH[2]), .Z(
        \ML_int[3][9] ) );
  MUX2_X2 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(SH[2]), .Z(
        \ML_int[3][8] ) );
  MUX2_X2 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(SH[2]), .Z(
        \ML_int[3][7] ) );
  MUX2_X2 M1_2_6 ( .A(\ML_int[2][6] ), .B(\ML_int[2][2] ), .S(SH[2]), .Z(
        \ML_int[3][6] ) );
  MUX2_X2 M1_2_5 ( .A(\ML_int[2][5] ), .B(n4), .S(SH[2]), .Z(\ML_int[3][5] )
         );
  MUX2_X2 M1_2_4 ( .A(\ML_int[2][4] ), .B(n2), .S(SH[2]), .Z(\ML_int[3][4] )
         );
  MUX2_X2 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S(SH[1]), .Z(
        \ML_int[2][10] ) );
  MUX2_X2 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S(SH[1]), .Z(
        \ML_int[2][9] ) );
  MUX2_X2 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S(SH[1]), .Z(
        \ML_int[2][8] ) );
  MUX2_X2 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S(SH[1]), .Z(
        \ML_int[2][7] ) );
  MUX2_X2 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S(SH[1]), .Z(
        \ML_int[2][6] ) );
  MUX2_X2 M1_1_5 ( .A(\ML_int[1][5] ), .B(\ML_int[1][3] ), .S(SH[1]), .Z(
        \ML_int[2][5] ) );
  MUX2_X2 M1_1_4 ( .A(\ML_int[1][4] ), .B(\ML_int[1][2] ), .S(SH[1]), .Z(
        \ML_int[2][4] ) );
  MUX2_X2 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(SH[1]), .Z(
        \ML_int[2][3] ) );
  MUX2_X2 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S(SH[1]), .Z(
        \ML_int[2][2] ) );
  MUX2_X2 M1_0_10 ( .A(A[10]), .B(A[9]), .S(SH[0]), .Z(\ML_int[1][10] ) );
  MUX2_X2 M1_0_9 ( .A(A[9]), .B(A[8]), .S(SH[0]), .Z(\ML_int[1][9] ) );
  MUX2_X2 M1_0_8 ( .A(A[8]), .B(A[7]), .S(SH[0]), .Z(\ML_int[1][8] ) );
  MUX2_X2 M1_0_7 ( .A(A[7]), .B(A[6]), .S(SH[0]), .Z(\ML_int[1][7] ) );
  MUX2_X2 M1_0_6 ( .A(A[6]), .B(A[5]), .S(SH[0]), .Z(\ML_int[1][6] ) );
  MUX2_X2 M1_0_5 ( .A(A[5]), .B(A[4]), .S(SH[0]), .Z(\ML_int[1][5] ) );
  MUX2_X2 M1_0_4 ( .A(A[4]), .B(A[3]), .S(SH[0]), .Z(\ML_int[1][4] ) );
  MUX2_X2 M1_0_3 ( .A(A[3]), .B(A[2]), .S(SH[0]), .Z(\ML_int[1][3] ) );
  MUX2_X2 M1_0_2 ( .A(A[2]), .B(A[1]), .S(SH[0]), .Z(\ML_int[1][2] ) );
  MUX2_X2 M1_0_1 ( .A(A[1]), .B(A[0]), .S(SH[0]), .Z(\ML_int[1][1] ) );
  AND2_X2 U3 ( .A1(A[0]), .A2(n1), .ZN(\ML_int[1][0] ) );
  INV_X4 U4 ( .A(SH[0]), .ZN(n1) );
  INV_X4 U5 ( .A(n11), .ZN(n2) );
  INV_X4 U6 ( .A(\ML_int[2][2] ), .ZN(n3) );
  INV_X4 U7 ( .A(n10), .ZN(n4) );
  INV_X4 U8 ( .A(\ML_int[2][3] ), .ZN(n5) );
  INV_X4 U9 ( .A(SH[3]), .ZN(n6) );
  INV_X4 U10 ( .A(SH[2]), .ZN(n7) );
  INV_X4 U11 ( .A(SH[1]), .ZN(n8) );
  AND2_X1 U12 ( .A1(\ML_int[3][7] ), .A2(n6), .ZN(\ML_int[4][7] ) );
  AND2_X1 U13 ( .A1(\ML_int[3][6] ), .A2(n6), .ZN(\ML_int[4][6] ) );
  AND2_X1 U14 ( .A1(\ML_int[3][5] ), .A2(n6), .ZN(\ML_int[4][5] ) );
  AND2_X1 U15 ( .A1(\ML_int[3][4] ), .A2(n6), .ZN(\ML_int[4][4] ) );
  NOR2_X1 U16 ( .A1(n5), .A2(n9), .ZN(\ML_int[4][3] ) );
  NOR2_X1 U17 ( .A1(n9), .A2(n3), .ZN(\ML_int[4][2] ) );
  NOR2_X1 U18 ( .A1(n9), .A2(n10), .ZN(\ML_int[4][1] ) );
  NOR2_X1 U19 ( .A1(n9), .A2(n11), .ZN(\ML_int[4][0] ) );
  NAND2_X1 U20 ( .A1(n7), .A2(n6), .ZN(n9) );
  NOR2_X1 U21 ( .A1(SH[2]), .A2(n3), .ZN(\ML_int[3][2] ) );
  NOR2_X1 U22 ( .A1(SH[2]), .A2(n10), .ZN(\ML_int[3][1] ) );
  NOR2_X1 U23 ( .A1(SH[2]), .A2(n11), .ZN(\ML_int[3][0] ) );
  NAND2_X1 U24 ( .A1(\ML_int[1][1] ), .A2(n8), .ZN(n10) );
  NAND2_X1 U25 ( .A1(\ML_int[1][0] ), .A2(n8), .ZN(n11) );
endmodule


module fpu_DW01_add_11 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   \A[9] , \A[8] , \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] ,
         \A[1] , \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83;
=======
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X2 U1 ( .A(A[8]), .B(carry[8]), .Z(SUM[8]) );
  AND2_X4 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
  AND2_X4 U3 ( .A1(A[8]), .A2(carry[8]), .ZN(n3) );
  AND2_X4 U4 ( .A1(A[9]), .A2(n3), .ZN(n4) );
  XOR2_X2 U5 ( .A(A[9]), .B(n3), .Z(SUM[9]) );
  XOR2_X2 U6 ( .A(A[10]), .B(n4), .Z(SUM[10]) );
  XOR2_X2 U7 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module fpu_DW01_add_8 ( A, B, CI, SUM, CO );
  input [103:0] A;
  input [103:0] B;
  output [103:0] SUM;
  input CI;
  output CO;
  wire   \A[50] , \A[49] , \A[48] , \A[47] , \A[46] , \A[45] , \A[44] ,
         \A[43] , \A[42] , \A[41] , \A[40] , \A[39] , \A[38] , \A[37] ,
         \A[36] , \A[35] , \A[34] , \A[33] , \A[32] , \A[31] , \A[30] ,
         \A[29] , \A[28] , \A[27] , \A[26] , \A[25] , \A[24] , \A[23] ,
         \A[22] , \A[21] , \A[20] , \A[19] , \A[18] , \A[17] , \A[16] ,
         \A[15] , \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] ,
         \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n1,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305;
  assign SUM[51] = A[51];
  assign SUM[50] = \A[50] ;
  assign \A[50]  = A[50];
  assign SUM[49] = \A[49] ;
  assign \A[49]  = A[49];
  assign SUM[48] = \A[48] ;
  assign \A[48]  = A[48];
  assign SUM[47] = \A[47] ;
  assign \A[47]  = A[47];
  assign SUM[46] = \A[46] ;
  assign \A[46]  = A[46];
  assign SUM[45] = \A[45] ;
  assign \A[45]  = A[45];
  assign SUM[44] = \A[44] ;
  assign \A[44]  = A[44];
  assign SUM[43] = \A[43] ;
  assign \A[43]  = A[43];
  assign SUM[42] = \A[42] ;
  assign \A[42]  = A[42];
  assign SUM[41] = \A[41] ;
  assign \A[41]  = A[41];
  assign SUM[40] = \A[40] ;
  assign \A[40]  = A[40];
  assign SUM[39] = \A[39] ;
  assign \A[39]  = A[39];
  assign SUM[38] = \A[38] ;
  assign \A[38]  = A[38];
  assign SUM[37] = \A[37] ;
  assign \A[37]  = A[37];
  assign SUM[36] = \A[36] ;
  assign \A[36]  = A[36];
  assign SUM[35] = \A[35] ;
  assign \A[35]  = A[35];
  assign SUM[34] = \A[34] ;
  assign \A[34]  = A[34];
  assign SUM[33] = \A[33] ;
  assign \A[33]  = A[33];
  assign SUM[32] = \A[32] ;
  assign \A[32]  = A[32];
  assign SUM[31] = \A[31] ;
  assign \A[31]  = A[31];
  assign SUM[30] = \A[30] ;
  assign \A[30]  = A[30];
  assign SUM[29] = \A[29] ;
  assign \A[29]  = A[29];
  assign SUM[28] = \A[28] ;
  assign \A[28]  = A[28];
  assign SUM[27] = \A[27] ;
  assign \A[27]  = A[27];
  assign SUM[26] = \A[26] ;
  assign \A[26]  = A[26];
  assign SUM[25] = \A[25] ;
  assign \A[25]  = A[25];
  assign SUM[24] = \A[24] ;
  assign \A[24]  = A[24];
  assign SUM[23] = \A[23] ;
  assign \A[23]  = A[23];
  assign SUM[22] = \A[22] ;
  assign \A[22]  = A[22];
  assign SUM[21] = \A[21] ;
  assign \A[21]  = A[21];
  assign SUM[20] = \A[20] ;
  assign \A[20]  = A[20];
  assign SUM[19] = \A[19] ;
  assign \A[19]  = A[19];
  assign SUM[18] = \A[18] ;
  assign \A[18]  = A[18];
  assign SUM[17] = \A[17] ;
  assign \A[17]  = A[17];
  assign SUM[16] = \A[16] ;
  assign \A[16]  = A[16];
  assign SUM[15] = \A[15] ;
  assign \A[15]  = A[15];
  assign SUM[14] = \A[14] ;
  assign \A[14]  = A[14];
  assign SUM[13] = \A[13] ;
  assign \A[13]  = A[13];
  assign SUM[12] = \A[12] ;
  assign \A[12]  = A[12];
  assign SUM[11] = \A[11] ;
  assign \A[11]  = A[11];
  assign SUM[10] = \A[10] ;
  assign \A[10]  = A[10];
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign SUM[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign SUM[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign SUM[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

<<<<<<< HEAD
  AND2_X2 U2 ( .A1(A[10]), .A2(B[10]), .ZN(n1) );
  NAND4_X2 U3 ( .A1(n46), .A2(n39), .A3(n78), .A4(n53), .ZN(n52) );
  INV_X4 U4 ( .A(A[11]), .ZN(n83) );
  INV_X4 U5 ( .A(n71), .ZN(n53) );
  AOI21_X2 U6 ( .B1(n23), .B2(n18), .A(n24), .ZN(n22) );
  AOI21_X2 U7 ( .B1(n62), .B2(n46), .A(n63), .ZN(n56) );
  INV_X4 U8 ( .A(n45), .ZN(n78) );
  OR2_X2 U9 ( .A1(n45), .A2(n71), .ZN(n2) );
  OR2_X2 U10 ( .A1(n25), .A2(n26), .ZN(n3) );
  OR2_X1 U11 ( .A1(n80), .A2(n71), .ZN(n4) );
  NOR2_X2 U12 ( .A1(n1), .A2(n48), .ZN(SUM[10]) );
  NOR2_X1 U13 ( .A1(A[10]), .A2(B[10]), .ZN(n48) );
  NAND2_X4 U14 ( .A1(n50), .A2(n51), .ZN(n72) );
  NAND2_X4 U15 ( .A1(n47), .A2(n49), .ZN(n35) );
  NAND2_X4 U16 ( .A1(n50), .A2(n51), .ZN(n49) );
  NAND2_X4 U17 ( .A1(n35), .A2(n36), .ZN(n31) );
  XNOR2_X1 U18 ( .A(n31), .B(n34), .ZN(SUM[16]) );
  INV_X8 U19 ( .A(n31), .ZN(n7) );
  NAND2_X4 U20 ( .A1(n82), .A2(n83), .ZN(n79) );
  NAND2_X1 U21 ( .A1(n51), .A2(n79), .ZN(n81) );
  NOR3_X2 U22 ( .A1(n44), .A2(n40), .A3(n45), .ZN(n37) );
  NOR2_X2 U23 ( .A1(n45), .A2(n69), .ZN(n68) );
  NAND2_X4 U24 ( .A1(n73), .A2(n74), .ZN(n46) );
  INV_X4 U25 ( .A(B[19]), .ZN(n5) );
  XNOR2_X2 U26 ( .A(n6), .B(n5), .ZN(SUM[19]) );
  OAI21_X4 U27 ( .B1(n7), .B2(n8), .A(n9), .ZN(n6) );
  AOI21_X4 U28 ( .B1(n10), .B2(n11), .A(n12), .ZN(n9) );
  INV_X4 U29 ( .A(n13), .ZN(n12) );
  NAND2_X2 U30 ( .A1(n14), .A2(n15), .ZN(n11) );
  NAND2_X2 U31 ( .A1(n10), .A2(n16), .ZN(n8) );
  INV_X4 U32 ( .A(n17), .ZN(n10) );
  NAND2_X2 U33 ( .A1(n18), .A2(n19), .ZN(n17) );
  XNOR2_X2 U34 ( .A(n21), .B(n20), .ZN(SUM[18]) );
  OAI21_X4 U35 ( .B1(n7), .B2(n3), .A(n22), .ZN(n21) );
  INV_X4 U36 ( .A(n14), .ZN(n24) );
  INV_X4 U37 ( .A(n15), .ZN(n23) );
  INV_X4 U38 ( .A(n18), .ZN(n25) );
  NAND2_X2 U39 ( .A1(n19), .A2(n13), .ZN(n20) );
  NAND2_X2 U40 ( .A1(B[18]), .A2(A[18]), .ZN(n13) );
  NAND2_X2 U41 ( .A1(n27), .A2(n28), .ZN(n19) );
  INV_X4 U42 ( .A(A[18]), .ZN(n28) );
  INV_X4 U43 ( .A(B[18]), .ZN(n27) );
  XNOR2_X2 U44 ( .A(n30), .B(n29), .ZN(SUM[17]) );
  OAI21_X4 U45 ( .B1(n7), .B2(n26), .A(n15), .ZN(n30) );
  INV_X4 U46 ( .A(n16), .ZN(n26) );
  NAND2_X2 U47 ( .A1(n14), .A2(n18), .ZN(n29) );
  NAND2_X2 U48 ( .A1(n32), .A2(n33), .ZN(n18) );
  INV_X4 U49 ( .A(A[17]), .ZN(n33) );
  INV_X4 U50 ( .A(B[17]), .ZN(n32) );
  NAND2_X2 U51 ( .A1(B[17]), .A2(A[17]), .ZN(n14) );
  OAI21_X4 U52 ( .B1(n37), .B2(n38), .A(n39), .ZN(n36) );
  OAI211_X2 U53 ( .C1(n40), .C2(n41), .A(n42), .B(n43), .ZN(n38) );
  NAND2_X2 U54 ( .A1(A[13]), .A2(B[13]), .ZN(n41) );
  INV_X4 U55 ( .A(n46), .ZN(n40) );
  NAND2_X2 U56 ( .A1(B[12]), .A2(A[12]), .ZN(n44) );
  INV_X4 U57 ( .A(n52), .ZN(n47) );
  NAND2_X2 U58 ( .A1(n16), .A2(n15), .ZN(n34) );
  NAND2_X2 U59 ( .A1(B[16]), .A2(A[16]), .ZN(n15) );
  NAND2_X2 U60 ( .A1(n54), .A2(n55), .ZN(n16) );
  INV_X4 U61 ( .A(A[16]), .ZN(n55) );
  INV_X4 U62 ( .A(B[16]), .ZN(n54) );
  XNOR2_X2 U63 ( .A(n56), .B(n57), .ZN(SUM[15]) );
  NOR2_X4 U64 ( .A1(n58), .A2(n59), .ZN(n57) );
  INV_X4 U65 ( .A(n42), .ZN(n59) );
  NAND2_X2 U66 ( .A1(B[15]), .A2(A[15]), .ZN(n42) );
  INV_X4 U67 ( .A(n39), .ZN(n58) );
  NAND2_X2 U68 ( .A1(n60), .A2(n61), .ZN(n39) );
  INV_X4 U69 ( .A(A[15]), .ZN(n61) );
  INV_X4 U70 ( .A(B[15]), .ZN(n60) );
  INV_X4 U71 ( .A(n43), .ZN(n63) );
  XNOR2_X2 U72 ( .A(n62), .B(n64), .ZN(SUM[14]) );
  OAI21_X4 U73 ( .B1(n65), .B2(n2), .A(n66), .ZN(n62) );
  NOR2_X4 U74 ( .A1(n67), .A2(n68), .ZN(n66) );
  INV_X4 U75 ( .A(n70), .ZN(n67) );
  INV_X4 U76 ( .A(n72), .ZN(n65) );
  NAND2_X2 U77 ( .A1(n46), .A2(n43), .ZN(n64) );
  NAND2_X2 U78 ( .A1(B[14]), .A2(A[14]), .ZN(n43) );
  INV_X4 U79 ( .A(A[14]), .ZN(n74) );
  INV_X4 U80 ( .A(B[14]), .ZN(n73) );
  XNOR2_X2 U81 ( .A(n76), .B(n75), .ZN(SUM[13]) );
  NAND2_X2 U82 ( .A1(n77), .A2(n69), .ZN(n76) );
  NAND2_X2 U83 ( .A1(n72), .A2(n53), .ZN(n77) );
  NAND2_X2 U84 ( .A1(n78), .A2(n70), .ZN(n75) );
  NAND2_X2 U85 ( .A1(B[13]), .A2(A[13]), .ZN(n70) );
  NOR2_X4 U86 ( .A1(A[13]), .A2(B[13]), .ZN(n45) );
  XNOR2_X2 U87 ( .A(n72), .B(n4), .ZN(SUM[12]) );
  NAND3_X4 U88 ( .A1(n79), .A2(B[10]), .A3(A[10]), .ZN(n50) );
  NOR2_X4 U89 ( .A1(A[12]), .A2(B[12]), .ZN(n71) );
  INV_X4 U90 ( .A(n69), .ZN(n80) );
  NAND2_X2 U91 ( .A1(B[12]), .A2(A[12]), .ZN(n69) );
  XNOR2_X2 U92 ( .A(n1), .B(n81), .ZN(SUM[11]) );
  NAND2_X2 U93 ( .A1(A[11]), .A2(B[11]), .ZN(n51) );
  INV_X4 U94 ( .A(B[11]), .ZN(n82) );
=======
  OR2_X4 U2 ( .A1(B[52]), .A2(A[52]), .ZN(n1) );
  AND2_X4 U3 ( .A1(n1), .A2(n264), .ZN(SUM[52]) );
  INV_X4 U4 ( .A(n266), .ZN(n3) );
  INV_X4 U5 ( .A(n272), .ZN(n4) );
  INV_X4 U6 ( .A(n274), .ZN(n5) );
  INV_X4 U7 ( .A(n72), .ZN(n6) );
  INV_X4 U8 ( .A(n76), .ZN(n7) );
  INV_X4 U9 ( .A(n80), .ZN(n8) );
  INV_X4 U10 ( .A(n84), .ZN(n9) );
  INV_X4 U11 ( .A(n82), .ZN(n10) );
  INV_X4 U12 ( .A(n90), .ZN(n11) );
  INV_X4 U13 ( .A(n92), .ZN(n12) );
  INV_X4 U14 ( .A(n93), .ZN(n13) );
  INV_X4 U15 ( .A(n100), .ZN(n14) );
  INV_X4 U16 ( .A(n283), .ZN(n15) );
  INV_X4 U17 ( .A(n106), .ZN(n16) );
  INV_X4 U18 ( .A(n109), .ZN(n17) );
  INV_X4 U19 ( .A(n107), .ZN(n18) );
  INV_X4 U20 ( .A(n114), .ZN(n19) );
  INV_X4 U21 ( .A(n112), .ZN(n20) );
  INV_X4 U22 ( .A(n115), .ZN(n21) );
  INV_X4 U23 ( .A(n126), .ZN(n22) );
  INV_X4 U24 ( .A(n128), .ZN(n23) );
  INV_X4 U25 ( .A(n129), .ZN(n24) );
  INV_X4 U26 ( .A(n135), .ZN(n25) );
  INV_X4 U27 ( .A(n133), .ZN(n26) );
  INV_X4 U28 ( .A(n289), .ZN(n27) );
  INV_X4 U29 ( .A(n146), .ZN(n28) );
  INV_X4 U30 ( .A(n144), .ZN(n29) );
  INV_X4 U31 ( .A(n148), .ZN(n30) );
  INV_X4 U32 ( .A(n151), .ZN(n31) );
  INV_X4 U33 ( .A(n156), .ZN(n32) );
  INV_X4 U34 ( .A(n157), .ZN(n33) );
  INV_X4 U35 ( .A(n164), .ZN(n34) );
  INV_X4 U36 ( .A(n165), .ZN(n35) );
  INV_X4 U37 ( .A(n177), .ZN(n36) );
  INV_X4 U38 ( .A(n179), .ZN(n37) );
  INV_X4 U39 ( .A(n180), .ZN(n38) );
  INV_X4 U40 ( .A(n186), .ZN(n39) );
  INV_X4 U41 ( .A(n184), .ZN(n40) );
  INV_X4 U42 ( .A(n297), .ZN(n41) );
  INV_X4 U43 ( .A(n298), .ZN(n42) );
  INV_X4 U44 ( .A(n198), .ZN(n43) );
  INV_X4 U45 ( .A(n195), .ZN(n44) );
  INV_X4 U46 ( .A(n197), .ZN(n45) );
  INV_X4 U47 ( .A(n200), .ZN(n46) );
  INV_X4 U48 ( .A(n203), .ZN(n47) );
  INV_X4 U49 ( .A(n208), .ZN(n48) );
  INV_X4 U50 ( .A(n204), .ZN(n49) );
  INV_X4 U51 ( .A(n211), .ZN(n50) );
  INV_X4 U52 ( .A(n209), .ZN(n51) );
  INV_X4 U53 ( .A(n216), .ZN(n52) );
  INV_X4 U54 ( .A(n214), .ZN(n53) );
  INV_X4 U55 ( .A(n218), .ZN(n54) );
  INV_X4 U56 ( .A(n224), .ZN(n55) );
  INV_X4 U57 ( .A(n228), .ZN(n56) );
  INV_X4 U58 ( .A(n232), .ZN(n57) );
  INV_X4 U59 ( .A(n236), .ZN(n58) );
  INV_X4 U60 ( .A(n234), .ZN(n59) );
  INV_X4 U61 ( .A(n240), .ZN(n60) );
  INV_X4 U62 ( .A(n244), .ZN(n61) );
  INV_X4 U63 ( .A(n248), .ZN(n62) );
  INV_X4 U64 ( .A(n252), .ZN(n63) );
  INV_X4 U65 ( .A(n256), .ZN(n64) );
  INV_X4 U66 ( .A(n253), .ZN(n65) );
  INV_X4 U67 ( .A(n260), .ZN(n66) );
  INV_X4 U68 ( .A(n263), .ZN(n67) );
  INV_X4 U69 ( .A(n264), .ZN(n68) );
  XOR2_X1 U70 ( .A(n69), .B(n70), .Z(SUM[99]) );
  NOR2_X1 U71 ( .A1(n71), .A2(n72), .ZN(n70) );
  XOR2_X1 U72 ( .A(n73), .B(n74), .Z(SUM[98]) );
  NAND2_X1 U73 ( .A1(n7), .A2(n75), .ZN(n73) );
  XOR2_X1 U74 ( .A(n77), .B(n78), .Z(SUM[97]) );
  NOR2_X1 U75 ( .A1(n79), .A2(n80), .ZN(n78) );
  XNOR2_X1 U76 ( .A(n81), .B(n82), .ZN(SUM[96]) );
  NAND2_X1 U77 ( .A1(n9), .A2(n83), .ZN(n81) );
  XOR2_X1 U78 ( .A(n85), .B(n86), .Z(SUM[95]) );
  AOI21_X1 U79 ( .B1(n87), .B2(n12), .A(n88), .ZN(n86) );
  NAND2_X1 U80 ( .A1(n11), .A2(n89), .ZN(n85) );
  XOR2_X1 U81 ( .A(n87), .B(n91), .Z(SUM[94]) );
  NOR2_X1 U82 ( .A1(n88), .A2(n92), .ZN(n91) );
  OAI21_X1 U83 ( .B1(n93), .B2(n94), .A(n95), .ZN(n87) );
  XOR2_X1 U84 ( .A(n96), .B(n94), .Z(SUM[93]) );
  AOI21_X1 U85 ( .B1(n14), .B2(n97), .A(n98), .ZN(n94) );
  NAND2_X1 U86 ( .A1(n13), .A2(n95), .ZN(n96) );
  XOR2_X1 U87 ( .A(n97), .B(n99), .Z(SUM[92]) );
  NOR2_X1 U88 ( .A1(n98), .A2(n100), .ZN(n99) );
  OAI21_X1 U89 ( .B1(n101), .B2(n102), .A(n15), .ZN(n97) );
  XOR2_X1 U90 ( .A(n103), .B(n104), .Z(SUM[91]) );
  NOR2_X1 U91 ( .A1(n16), .A2(n105), .ZN(n104) );
  OAI21_X1 U92 ( .B1(n107), .B2(n108), .A(n109), .ZN(n103) );
  XOR2_X1 U93 ( .A(n110), .B(n108), .Z(SUM[90]) );
  AOI21_X1 U94 ( .B1(n20), .B2(n111), .A(n19), .ZN(n108) );
  NAND2_X1 U95 ( .A1(n18), .A2(n109), .ZN(n110) );
  XOR2_X1 U96 ( .A(n111), .B(n113), .Z(SUM[89]) );
  NOR2_X1 U97 ( .A1(n19), .A2(n112), .ZN(n113) );
  OAI21_X1 U98 ( .B1(n115), .B2(n101), .A(n116), .ZN(n111) );
  XOR2_X1 U99 ( .A(n117), .B(n101), .Z(SUM[88]) );
  AOI21_X1 U100 ( .B1(n118), .B2(n119), .A(n120), .ZN(n101) );
  NAND2_X1 U101 ( .A1(n21), .A2(n116), .ZN(n117) );
  XOR2_X1 U102 ( .A(n121), .B(n122), .Z(SUM[87]) );
  AOI21_X1 U103 ( .B1(n123), .B2(n23), .A(n124), .ZN(n122) );
  NAND2_X1 U104 ( .A1(n22), .A2(n125), .ZN(n121) );
  XOR2_X1 U105 ( .A(n123), .B(n127), .Z(SUM[86]) );
  NOR2_X1 U106 ( .A1(n124), .A2(n128), .ZN(n127) );
  OAI21_X1 U107 ( .B1(n129), .B2(n130), .A(n131), .ZN(n123) );
  XOR2_X1 U108 ( .A(n132), .B(n130), .Z(SUM[85]) );
  AOI21_X1 U109 ( .B1(n26), .B2(n118), .A(n25), .ZN(n130) );
  NAND2_X1 U110 ( .A1(n24), .A2(n131), .ZN(n132) );
  XOR2_X1 U111 ( .A(n118), .B(n134), .Z(SUM[84]) );
  NOR2_X1 U112 ( .A1(n25), .A2(n133), .ZN(n134) );
  OR2_X1 U113 ( .A1(n136), .A2(n137), .ZN(n118) );
  XOR2_X1 U114 ( .A(n138), .B(n139), .Z(SUM[83]) );
  AOI21_X1 U115 ( .B1(n140), .B2(n141), .A(n28), .ZN(n139) );
  NAND2_X1 U116 ( .A1(n27), .A2(n142), .ZN(n138) );
  XNOR2_X1 U117 ( .A(n143), .B(n140), .ZN(SUM[82]) );
  OAI21_X1 U118 ( .B1(n144), .B2(n30), .A(n145), .ZN(n140) );
  NAND2_X1 U119 ( .A1(n141), .A2(n146), .ZN(n143) );
  XOR2_X1 U120 ( .A(n147), .B(n30), .Z(SUM[81]) );
  OAI21_X1 U121 ( .B1(n149), .B2(n150), .A(n151), .ZN(n148) );
  NAND2_X1 U122 ( .A1(n29), .A2(n145), .ZN(n147) );
  XNOR2_X1 U123 ( .A(n149), .B(n152), .ZN(SUM[80]) );
  NOR2_X1 U124 ( .A1(n31), .A2(n150), .ZN(n152) );
  XOR2_X1 U125 ( .A(n153), .B(n154), .Z(SUM[79]) );
  NOR2_X1 U126 ( .A1(n155), .A2(n156), .ZN(n154) );
  OAI21_X1 U127 ( .B1(n157), .B2(n158), .A(n159), .ZN(n153) );
  XOR2_X1 U128 ( .A(n160), .B(n158), .Z(SUM[78]) );
  AOI21_X1 U129 ( .B1(n34), .B2(n161), .A(n162), .ZN(n158) );
  NAND2_X1 U130 ( .A1(n33), .A2(n159), .ZN(n160) );
  XOR2_X1 U131 ( .A(n161), .B(n163), .Z(SUM[77]) );
  NOR2_X1 U132 ( .A1(n162), .A2(n164), .ZN(n163) );
  OAI21_X1 U133 ( .B1(n165), .B2(n166), .A(n167), .ZN(n161) );
  XOR2_X1 U134 ( .A(n168), .B(n166), .Z(SUM[76]) );
  AOI21_X1 U135 ( .B1(n169), .B2(n170), .A(n171), .ZN(n166) );
  NAND2_X1 U136 ( .A1(n35), .A2(n167), .ZN(n168) );
  XOR2_X1 U137 ( .A(n172), .B(n173), .Z(SUM[75]) );
  AOI21_X1 U138 ( .B1(n174), .B2(n37), .A(n175), .ZN(n173) );
  NAND2_X1 U139 ( .A1(n36), .A2(n176), .ZN(n172) );
  XOR2_X1 U140 ( .A(n174), .B(n178), .Z(SUM[74]) );
  NOR2_X1 U141 ( .A1(n175), .A2(n179), .ZN(n178) );
  OAI21_X1 U142 ( .B1(n180), .B2(n181), .A(n182), .ZN(n174) );
  XOR2_X1 U143 ( .A(n183), .B(n181), .Z(SUM[73]) );
  AOI21_X1 U144 ( .B1(n40), .B2(n169), .A(n39), .ZN(n181) );
  NAND2_X1 U145 ( .A1(n38), .A2(n182), .ZN(n183) );
  XOR2_X1 U146 ( .A(n169), .B(n185), .Z(SUM[72]) );
  NOR2_X1 U147 ( .A1(n39), .A2(n184), .ZN(n185) );
  OAI21_X1 U148 ( .B1(n187), .B2(n188), .A(n41), .ZN(n169) );
  XOR2_X1 U149 ( .A(n189), .B(n190), .Z(SUM[71]) );
  AOI21_X1 U150 ( .B1(n191), .B2(n192), .A(n43), .ZN(n190) );
  NAND2_X1 U151 ( .A1(n42), .A2(n193), .ZN(n189) );
  XNOR2_X1 U152 ( .A(n194), .B(n191), .ZN(SUM[70]) );
  OAI21_X1 U153 ( .B1(n195), .B2(n45), .A(n196), .ZN(n191) );
  NAND2_X1 U154 ( .A1(n192), .A2(n198), .ZN(n194) );
  XNOR2_X1 U155 ( .A(n199), .B(n197), .ZN(SUM[69]) );
  OAI21_X1 U156 ( .B1(n200), .B2(n187), .A(n201), .ZN(n197) );
  NAND2_X1 U157 ( .A1(n44), .A2(n196), .ZN(n199) );
  XOR2_X1 U158 ( .A(n202), .B(n187), .Z(SUM[68]) );
  NOR2_X1 U159 ( .A1(n203), .A2(n204), .ZN(n187) );
  NAND2_X1 U160 ( .A1(n46), .A2(n201), .ZN(n202) );
  XOR2_X1 U161 ( .A(n205), .B(n206), .Z(SUM[67]) );
  NOR2_X1 U162 ( .A1(n48), .A2(n207), .ZN(n206) );
  OAI21_X1 U163 ( .B1(n209), .B2(n210), .A(n211), .ZN(n205) );
  XOR2_X1 U164 ( .A(n212), .B(n210), .Z(SUM[66]) );
  AOI21_X1 U165 ( .B1(n53), .B2(n213), .A(n52), .ZN(n210) );
  NAND2_X1 U166 ( .A1(n51), .A2(n211), .ZN(n212) );
  XOR2_X1 U167 ( .A(n213), .B(n215), .Z(SUM[65]) );
  NOR2_X1 U168 ( .A1(n52), .A2(n214), .ZN(n215) );
  OAI21_X1 U169 ( .B1(n217), .B2(n218), .A(n219), .ZN(n213) );
  XOR2_X1 U170 ( .A(n220), .B(n217), .Z(SUM[64]) );
  NAND2_X1 U171 ( .A1(n54), .A2(n219), .ZN(n220) );
  XOR2_X1 U172 ( .A(n221), .B(n222), .Z(SUM[63]) );
  NOR2_X1 U173 ( .A1(n223), .A2(n224), .ZN(n222) );
  XOR2_X1 U174 ( .A(n225), .B(n226), .Z(SUM[62]) );
  NAND2_X1 U175 ( .A1(n56), .A2(n227), .ZN(n225) );
  XOR2_X1 U176 ( .A(n229), .B(n230), .Z(SUM[61]) );
  NOR2_X1 U177 ( .A1(n231), .A2(n232), .ZN(n230) );
  XNOR2_X1 U178 ( .A(n233), .B(n234), .ZN(SUM[60]) );
  NAND2_X1 U179 ( .A1(n58), .A2(n235), .ZN(n233) );
  XNOR2_X1 U180 ( .A(n237), .B(n238), .ZN(SUM[59]) );
  NOR2_X1 U181 ( .A1(n60), .A2(n239), .ZN(n238) );
  XNOR2_X1 U182 ( .A(n241), .B(n242), .ZN(SUM[58]) );
  NAND2_X1 U183 ( .A1(n243), .A2(n244), .ZN(n241) );
  XNOR2_X1 U184 ( .A(n245), .B(n246), .ZN(SUM[57]) );
  NOR2_X1 U185 ( .A1(n62), .A2(n247), .ZN(n246) );
  XNOR2_X1 U186 ( .A(n249), .B(n250), .ZN(SUM[56]) );
  NAND2_X1 U187 ( .A1(n251), .A2(n252), .ZN(n249) );
  XOR2_X1 U188 ( .A(n253), .B(n254), .Z(SUM[55]) );
  NOR2_X1 U189 ( .A1(n64), .A2(n255), .ZN(n254) );
  XOR2_X1 U190 ( .A(n257), .B(n258), .Z(SUM[54]) );
  NAND2_X1 U191 ( .A1(n66), .A2(n259), .ZN(n257) );
  XOR2_X1 U192 ( .A(n68), .B(n261), .Z(SUM[53]) );
  NOR2_X1 U193 ( .A1(n262), .A2(n263), .ZN(n261) );
  XOR2_X1 U194 ( .A(n265), .B(B[103]), .Z(SUM[103]) );
  OAI21_X1 U195 ( .B1(n266), .B2(n267), .A(n268), .ZN(n265) );
  XOR2_X1 U196 ( .A(n269), .B(n267), .Z(SUM[102]) );
  AOI21_X1 U197 ( .B1(n4), .B2(n270), .A(n271), .ZN(n267) );
  NAND2_X1 U198 ( .A1(n3), .A2(n268), .ZN(n269) );
  NAND2_X1 U199 ( .A1(B[102]), .A2(A[102]), .ZN(n268) );
  NOR2_X1 U200 ( .A1(B[102]), .A2(A[102]), .ZN(n266) );
  XOR2_X1 U201 ( .A(n270), .B(n273), .Z(SUM[101]) );
  NOR2_X1 U202 ( .A1(n271), .A2(n272), .ZN(n273) );
  NOR2_X1 U203 ( .A1(B[101]), .A2(A[101]), .ZN(n272) );
  AND2_X1 U204 ( .A1(B[101]), .A2(A[101]), .ZN(n271) );
  OAI21_X1 U205 ( .B1(n274), .B2(n275), .A(n276), .ZN(n270) );
  XOR2_X1 U206 ( .A(n277), .B(n275), .Z(SUM[100]) );
  AOI21_X1 U207 ( .B1(n69), .B2(n6), .A(n71), .ZN(n275) );
  AND2_X1 U208 ( .A1(B[99]), .A2(A[99]), .ZN(n71) );
  NOR2_X1 U209 ( .A1(B[99]), .A2(A[99]), .ZN(n72) );
  OAI21_X1 U210 ( .B1(n76), .B2(n74), .A(n75), .ZN(n69) );
  NAND2_X1 U211 ( .A1(B[98]), .A2(A[98]), .ZN(n75) );
  AOI21_X1 U212 ( .B1(n8), .B2(n77), .A(n79), .ZN(n74) );
  AND2_X1 U213 ( .A1(B[97]), .A2(A[97]), .ZN(n79) );
  OAI21_X1 U214 ( .B1(n10), .B2(n84), .A(n83), .ZN(n77) );
  NAND2_X1 U215 ( .A1(B[96]), .A2(A[96]), .ZN(n83) );
  NOR2_X1 U216 ( .A1(B[96]), .A2(A[96]), .ZN(n84) );
  OAI21_X1 U217 ( .B1(n90), .B2(n278), .A(n89), .ZN(n82) );
  NAND2_X1 U218 ( .A1(B[95]), .A2(A[95]), .ZN(n89) );
  AOI21_X1 U219 ( .B1(n279), .B2(n12), .A(n88), .ZN(n278) );
  AND2_X1 U220 ( .A1(B[94]), .A2(A[94]), .ZN(n88) );
  NOR2_X1 U221 ( .A1(B[94]), .A2(A[94]), .ZN(n92) );
  OAI21_X1 U222 ( .B1(n93), .B2(n280), .A(n95), .ZN(n279) );
  NAND2_X1 U223 ( .A1(B[93]), .A2(A[93]), .ZN(n95) );
  AOI21_X1 U224 ( .B1(n281), .B2(n14), .A(n98), .ZN(n280) );
  AND2_X1 U225 ( .A1(B[92]), .A2(A[92]), .ZN(n98) );
  NOR2_X1 U226 ( .A1(B[92]), .A2(A[92]), .ZN(n100) );
  OAI21_X1 U227 ( .B1(n282), .B2(n102), .A(n15), .ZN(n281) );
  OAI21_X1 U228 ( .B1(n105), .B2(n284), .A(n106), .ZN(n283) );
  NAND2_X1 U229 ( .A1(B[91]), .A2(A[91]), .ZN(n106) );
  AOI21_X1 U230 ( .B1(n285), .B2(n18), .A(n17), .ZN(n284) );
  NAND2_X1 U231 ( .A1(B[90]), .A2(A[90]), .ZN(n109) );
  OAI21_X1 U232 ( .B1(n112), .B2(n116), .A(n114), .ZN(n285) );
  NAND2_X1 U233 ( .A1(B[89]), .A2(A[89]), .ZN(n114) );
  NAND2_X1 U234 ( .A1(B[88]), .A2(A[88]), .ZN(n116) );
  OR4_X1 U235 ( .A1(n105), .A2(n107), .A3(n112), .A4(n115), .ZN(n102) );
  NOR2_X1 U236 ( .A1(B[88]), .A2(A[88]), .ZN(n115) );
  NOR2_X1 U237 ( .A1(B[89]), .A2(A[89]), .ZN(n112) );
  NOR2_X1 U238 ( .A1(B[90]), .A2(A[90]), .ZN(n107) );
  NOR2_X1 U239 ( .A1(B[91]), .A2(A[91]), .ZN(n105) );
  AOI221_X1 U240 ( .B1(n119), .B2(n136), .C1(n137), .C2(n119), .A(n120), .ZN(
        n282) );
  OAI21_X1 U241 ( .B1(n126), .B2(n286), .A(n125), .ZN(n120) );
  NAND2_X1 U242 ( .A1(B[87]), .A2(A[87]), .ZN(n125) );
  AOI21_X1 U243 ( .B1(n287), .B2(n23), .A(n124), .ZN(n286) );
  AND2_X1 U244 ( .A1(B[86]), .A2(A[86]), .ZN(n124) );
  OAI21_X1 U245 ( .B1(n129), .B2(n135), .A(n131), .ZN(n287) );
  NAND2_X1 U246 ( .A1(B[85]), .A2(A[85]), .ZN(n131) );
  NAND2_X1 U247 ( .A1(B[84]), .A2(A[84]), .ZN(n135) );
  NOR4_X1 U248 ( .A1(n150), .A2(n149), .A3(n144), .A4(n288), .ZN(n137) );
  NAND2_X1 U249 ( .A1(n141), .A2(n27), .ZN(n288) );
  AOI21_X1 U250 ( .B1(n32), .B2(n290), .A(n155), .ZN(n149) );
  AND2_X1 U251 ( .A1(B[79]), .A2(A[79]), .ZN(n155) );
  OAI21_X1 U252 ( .B1(n291), .B2(n157), .A(n159), .ZN(n290) );
  NAND2_X1 U253 ( .A1(B[78]), .A2(A[78]), .ZN(n159) );
  NOR2_X1 U254 ( .A1(B[78]), .A2(A[78]), .ZN(n157) );
  AOI21_X1 U255 ( .B1(n34), .B2(n292), .A(n162), .ZN(n291) );
  AND2_X1 U256 ( .A1(B[77]), .A2(A[77]), .ZN(n162) );
  OAI21_X1 U257 ( .B1(n293), .B2(n165), .A(n167), .ZN(n292) );
  NAND2_X1 U258 ( .A1(B[76]), .A2(A[76]), .ZN(n167) );
  NOR2_X1 U259 ( .A1(B[76]), .A2(A[76]), .ZN(n165) );
  AOI21_X1 U260 ( .B1(n294), .B2(n170), .A(n171), .ZN(n293) );
  OAI21_X1 U261 ( .B1(n177), .B2(n295), .A(n176), .ZN(n171) );
  NAND2_X1 U262 ( .A1(B[75]), .A2(A[75]), .ZN(n176) );
  AOI21_X1 U263 ( .B1(n296), .B2(n37), .A(n175), .ZN(n295) );
  AND2_X1 U264 ( .A1(B[74]), .A2(A[74]), .ZN(n175) );
  OAI21_X1 U265 ( .B1(n180), .B2(n186), .A(n182), .ZN(n296) );
  NAND2_X1 U266 ( .A1(B[73]), .A2(A[73]), .ZN(n182) );
  NAND2_X1 U267 ( .A1(B[72]), .A2(A[72]), .ZN(n186) );
  NOR4_X1 U268 ( .A1(n177), .A2(n179), .A3(n180), .A4(n184), .ZN(n170) );
  NOR2_X1 U269 ( .A1(B[72]), .A2(A[72]), .ZN(n184) );
  NOR2_X1 U270 ( .A1(B[73]), .A2(A[73]), .ZN(n180) );
  NOR2_X1 U271 ( .A1(B[74]), .A2(A[74]), .ZN(n179) );
  NOR2_X1 U272 ( .A1(B[75]), .A2(A[75]), .ZN(n177) );
  OAI221_X1 U273 ( .B1(n188), .B2(n47), .C1(n49), .C2(n188), .A(n41), .ZN(n294) );
  OAI21_X1 U274 ( .B1(n298), .B2(n299), .A(n193), .ZN(n297) );
  NAND2_X1 U275 ( .A1(B[71]), .A2(A[71]), .ZN(n193) );
  AOI21_X1 U276 ( .B1(n300), .B2(n192), .A(n43), .ZN(n299) );
  NAND2_X1 U277 ( .A1(B[70]), .A2(A[70]), .ZN(n198) );
  OAI21_X1 U278 ( .B1(n195), .B2(n201), .A(n196), .ZN(n300) );
  NAND2_X1 U279 ( .A1(B[69]), .A2(A[69]), .ZN(n196) );
  NAND2_X1 U280 ( .A1(B[68]), .A2(A[68]), .ZN(n201) );
  NOR4_X1 U281 ( .A1(n207), .A2(n209), .A3(n301), .A4(n214), .ZN(n204) );
  OR2_X1 U282 ( .A1(n217), .A2(n218), .ZN(n301) );
  NOR2_X1 U283 ( .A1(B[64]), .A2(A[64]), .ZN(n218) );
  AOI21_X1 U284 ( .B1(n55), .B2(n221), .A(n223), .ZN(n217) );
  AND2_X1 U285 ( .A1(B[63]), .A2(A[63]), .ZN(n223) );
  OAI21_X1 U286 ( .B1(n228), .B2(n226), .A(n227), .ZN(n221) );
  NAND2_X1 U287 ( .A1(B[62]), .A2(A[62]), .ZN(n227) );
  AOI21_X1 U288 ( .B1(n57), .B2(n229), .A(n231), .ZN(n226) );
  AND2_X1 U289 ( .A1(B[61]), .A2(A[61]), .ZN(n231) );
  OAI21_X1 U290 ( .B1(n236), .B2(n59), .A(n235), .ZN(n229) );
  NAND2_X1 U291 ( .A1(B[60]), .A2(A[60]), .ZN(n235) );
  OAI21_X1 U292 ( .B1(n239), .B2(n237), .A(n240), .ZN(n234) );
  NAND2_X1 U293 ( .A1(B[59]), .A2(A[59]), .ZN(n240) );
  AOI21_X1 U294 ( .B1(n243), .B2(n242), .A(n61), .ZN(n237) );
  NAND2_X1 U295 ( .A1(B[58]), .A2(A[58]), .ZN(n244) );
  OAI21_X1 U296 ( .B1(n247), .B2(n245), .A(n248), .ZN(n242) );
  NAND2_X1 U297 ( .A1(B[57]), .A2(A[57]), .ZN(n248) );
  AOI21_X1 U298 ( .B1(n251), .B2(n250), .A(n63), .ZN(n245) );
  NAND2_X1 U299 ( .A1(B[56]), .A2(A[56]), .ZN(n252) );
  OAI21_X1 U300 ( .B1(n255), .B2(n65), .A(n256), .ZN(n250) );
  NAND2_X1 U301 ( .A1(B[55]), .A2(A[55]), .ZN(n256) );
  OAI21_X1 U302 ( .B1(n260), .B2(n258), .A(n259), .ZN(n253) );
  NAND2_X1 U303 ( .A1(B[54]), .A2(A[54]), .ZN(n259) );
  AOI21_X1 U304 ( .B1(n67), .B2(n68), .A(n262), .ZN(n258) );
  AND2_X1 U305 ( .A1(B[53]), .A2(A[53]), .ZN(n262) );
  NAND2_X1 U306 ( .A1(B[52]), .A2(A[52]), .ZN(n264) );
  NOR2_X1 U307 ( .A1(B[53]), .A2(A[53]), .ZN(n263) );
  NOR2_X1 U308 ( .A1(B[54]), .A2(A[54]), .ZN(n260) );
  NOR2_X1 U309 ( .A1(B[55]), .A2(A[55]), .ZN(n255) );
  OR2_X1 U310 ( .A1(B[56]), .A2(A[56]), .ZN(n251) );
  NOR2_X1 U311 ( .A1(B[57]), .A2(A[57]), .ZN(n247) );
  OR2_X1 U312 ( .A1(B[58]), .A2(A[58]), .ZN(n243) );
  NOR2_X1 U313 ( .A1(B[59]), .A2(A[59]), .ZN(n239) );
  NOR2_X1 U314 ( .A1(B[60]), .A2(A[60]), .ZN(n236) );
  NOR2_X1 U315 ( .A1(B[61]), .A2(A[61]), .ZN(n232) );
  NOR2_X1 U316 ( .A1(B[62]), .A2(A[62]), .ZN(n228) );
  NOR2_X1 U317 ( .A1(B[63]), .A2(A[63]), .ZN(n224) );
  OAI21_X1 U318 ( .B1(n207), .B2(n302), .A(n208), .ZN(n203) );
  NAND2_X1 U319 ( .A1(B[67]), .A2(A[67]), .ZN(n208) );
  AOI21_X1 U320 ( .B1(n303), .B2(n51), .A(n50), .ZN(n302) );
  NAND2_X1 U321 ( .A1(B[66]), .A2(A[66]), .ZN(n211) );
  NOR2_X1 U322 ( .A1(B[66]), .A2(A[66]), .ZN(n209) );
  OAI21_X1 U323 ( .B1(n214), .B2(n219), .A(n216), .ZN(n303) );
  NAND2_X1 U324 ( .A1(B[65]), .A2(A[65]), .ZN(n216) );
  NAND2_X1 U325 ( .A1(B[64]), .A2(A[64]), .ZN(n219) );
  NOR2_X1 U326 ( .A1(B[65]), .A2(A[65]), .ZN(n214) );
  NOR2_X1 U327 ( .A1(B[67]), .A2(A[67]), .ZN(n207) );
  NAND4_X1 U328 ( .A1(n42), .A2(n192), .A3(n44), .A4(n46), .ZN(n188) );
  NOR2_X1 U329 ( .A1(B[68]), .A2(A[68]), .ZN(n200) );
  NOR2_X1 U330 ( .A1(B[69]), .A2(A[69]), .ZN(n195) );
  OR2_X1 U331 ( .A1(B[70]), .A2(A[70]), .ZN(n192) );
  NOR2_X1 U332 ( .A1(B[71]), .A2(A[71]), .ZN(n298) );
  NOR2_X1 U333 ( .A1(B[77]), .A2(A[77]), .ZN(n164) );
  NOR2_X1 U334 ( .A1(B[79]), .A2(A[79]), .ZN(n156) );
  NOR2_X1 U335 ( .A1(B[80]), .A2(A[80]), .ZN(n150) );
  OAI21_X1 U336 ( .B1(n289), .B2(n304), .A(n142), .ZN(n136) );
  NAND2_X1 U337 ( .A1(B[83]), .A2(A[83]), .ZN(n142) );
  AOI21_X1 U338 ( .B1(n305), .B2(n141), .A(n28), .ZN(n304) );
  NAND2_X1 U339 ( .A1(B[82]), .A2(A[82]), .ZN(n146) );
  OR2_X1 U340 ( .A1(B[82]), .A2(A[82]), .ZN(n141) );
  OAI21_X1 U341 ( .B1(n144), .B2(n151), .A(n145), .ZN(n305) );
  NAND2_X1 U342 ( .A1(B[81]), .A2(A[81]), .ZN(n145) );
  NAND2_X1 U343 ( .A1(B[80]), .A2(A[80]), .ZN(n151) );
  NOR2_X1 U344 ( .A1(B[81]), .A2(A[81]), .ZN(n144) );
  NOR2_X1 U345 ( .A1(B[83]), .A2(A[83]), .ZN(n289) );
  NOR4_X1 U346 ( .A1(n126), .A2(n128), .A3(n129), .A4(n133), .ZN(n119) );
  NOR2_X1 U347 ( .A1(B[84]), .A2(A[84]), .ZN(n133) );
  NOR2_X1 U348 ( .A1(B[85]), .A2(A[85]), .ZN(n129) );
  NOR2_X1 U349 ( .A1(B[86]), .A2(A[86]), .ZN(n128) );
  NOR2_X1 U350 ( .A1(B[87]), .A2(A[87]), .ZN(n126) );
  NOR2_X1 U351 ( .A1(B[93]), .A2(A[93]), .ZN(n93) );
  NOR2_X1 U352 ( .A1(B[95]), .A2(A[95]), .ZN(n90) );
  NOR2_X1 U353 ( .A1(B[97]), .A2(A[97]), .ZN(n80) );
  NOR2_X1 U354 ( .A1(B[98]), .A2(A[98]), .ZN(n76) );
  NAND2_X1 U355 ( .A1(n5), .A2(n276), .ZN(n277) );
  NAND2_X1 U356 ( .A1(B[100]), .A2(A[100]), .ZN(n276) );
  NOR2_X1 U357 ( .A1(B[100]), .A2(A[100]), .ZN(n274) );
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
endmodule


module fpu_DW02_mult_0 ( A, B, TC, PRODUCT );
<<<<<<< HEAD
  input [10:0] A;
  input [10:0] B;
  output [21:0] PRODUCT;
  input TC;
  wire   \ab[10][10] , \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] ,
         \ab[10][5] , \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] ,
         \ab[10][0] , \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] ,
         \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] ,
         \ab[9][1] , \ab[9][0] , \ab[8][10] , \ab[8][9] , \ab[8][8] ,
         \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] , \ab[8][3] ,
         \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][10] , \ab[7][9] ,
         \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] , \ab[7][4] ,
         \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] , \ab[6][10] ,
         \ab[6][9] , \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] ,
         \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] ,
         \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] ,
         \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] ,
         \ab[5][0] , \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] ,
         \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] ,
         \ab[4][1] , \ab[4][0] , \ab[3][10] , \ab[3][9] , \ab[3][8] ,
         \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][10] , \ab[2][9] ,
         \ab[2][8] , \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] ,
         \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] , \ab[1][10] ,
         \ab[1][9] , \ab[1][8] , \ab[1][7] , \ab[1][6] , \ab[1][5] ,
         \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[1][0] ,
         \ab[0][9] , \ab[0][8] , \ab[0][7] , \ab[0][6] , \ab[0][5] ,
         \ab[0][4] , \ab[0][3] , \ab[0][2] , \ab[0][1] , \CARRYB[10][9] ,
         \CARRYB[10][8] , \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] ,
         \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] ,
         \CARRYB[10][0] , \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] ,
         \CARRYB[9][6] , \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] ,
         \CARRYB[9][2] , \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][9] ,
         \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] ,
         \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] ,
         \CARRYB[8][0] , \CARRYB[7][9] , \CARRYB[7][8] , \CARRYB[7][7] ,
         \CARRYB[7][6] , \CARRYB[7][5] , \CARRYB[7][4] , \CARRYB[7][3] ,
         \CARRYB[7][2] , \CARRYB[7][1] , \CARRYB[7][0] , \CARRYB[6][9] ,
         \CARRYB[6][8] , \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] ,
         \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] ,
         \CARRYB[6][0] , \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] ,
         \CARRYB[5][6] , \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] ,
         \CARRYB[5][2] , \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][9] ,
         \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] ,
         \CARRYB[4][0] , \CARRYB[3][9] , \CARRYB[3][8] , \CARRYB[3][7] ,
         \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][4] , \CARRYB[3][3] ,
         \CARRYB[3][2] , \CARRYB[3][1] , \CARRYB[3][0] , \CARRYB[2][9] ,
         \CARRYB[2][8] , \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \CARRYB[1][9] , \CARRYB[1][8] , \CARRYB[1][7] ,
         \CARRYB[1][6] , \CARRYB[1][5] , \CARRYB[1][4] , \CARRYB[1][3] ,
         \CARRYB[1][2] , \CARRYB[1][1] , \CARRYB[1][0] , \SUMB[10][9] ,
         \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] , \SUMB[10][5] ,
         \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] , \SUMB[10][1] ,
         \SUMB[10][0] , \SUMB[9][9] , \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] ,
         \SUMB[9][5] , \SUMB[9][4] , \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] ,
         \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] ,
         \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][9] ,
         \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] , \SUMB[7][4] ,
         \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][9] , \SUMB[6][8] ,
         \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] , \SUMB[6][4] , \SUMB[6][3] ,
         \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] ,
         \SUMB[5][6] , \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] ,
         \SUMB[5][1] , \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][9] ,
         \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] ,
         \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][9] , \SUMB[1][8] ,
         \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] ,
         \SUMB[1][2] , \SUMB[1][1] , n3, n4, n5, n6, n7, n8, n9, n10, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69;
  wire   [19:16] CLA_CARRY;
  wire   [19:2] CLA_SUM;

  FA_X1 S4_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\SUMB[10][0] ) );
  FA_X1 S4_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA_X1 S4_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA_X1 S4_3 ( .A(\CARRYB[9][3] ), .B(\ab[10][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA_X1 S4_4 ( .A(\CARRYB[9][4] ), .B(\ab[10][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA_X1 S4_5 ( .A(\CARRYB[9][5] ), .B(\ab[10][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA_X1 S4_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA_X1 S4_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA_X1 S4_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA_X1 S5_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\ab[9][10] ), .CO(
        \CARRYB[10][9] ), .S(\SUMB[10][9] ) );
=======
  input [52:0] A;
  input [52:0] B;
  output [105:0] PRODUCT;
  input TC;
  wire   \ab[52][52] , \ab[52][51] , \ab[52][50] , \ab[52][49] , \ab[52][48] ,
         \ab[52][47] , \ab[52][46] , \ab[52][45] , \ab[52][44] , \ab[52][43] ,
         \ab[52][42] , \ab[52][41] , \ab[52][40] , \ab[52][39] , \ab[52][38] ,
         \ab[52][37] , \ab[52][36] , \ab[52][35] , \ab[52][34] , \ab[52][33] ,
         \ab[52][32] , \ab[52][31] , \ab[52][30] , \ab[52][29] , \ab[52][28] ,
         \ab[52][27] , \ab[52][26] , \ab[52][25] , \ab[52][24] , \ab[52][23] ,
         \ab[52][22] , \ab[52][21] , \ab[52][20] , \ab[52][19] , \ab[52][18] ,
         \ab[52][17] , \ab[52][16] , \ab[52][15] , \ab[52][14] , \ab[52][13] ,
         \ab[52][12] , \ab[52][11] , \ab[52][10] , \ab[52][9] , \ab[52][8] ,
         \ab[52][7] , \ab[52][6] , \ab[52][5] , \ab[52][4] , \ab[52][3] ,
         \ab[52][2] , \ab[52][1] , \ab[52][0] , \ab[51][52] , \ab[51][51] ,
         \ab[51][50] , \ab[51][49] , \ab[51][48] , \ab[51][47] , \ab[51][46] ,
         \ab[51][45] , \ab[51][44] , \ab[51][43] , \ab[51][42] , \ab[51][41] ,
         \ab[51][40] , \ab[51][39] , \ab[51][38] , \ab[51][37] , \ab[51][36] ,
         \ab[51][35] , \ab[51][34] , \ab[51][33] , \ab[51][32] , \ab[51][31] ,
         \ab[51][30] , \ab[51][29] , \ab[51][28] , \ab[51][27] , \ab[51][26] ,
         \ab[51][25] , \ab[51][24] , \ab[51][23] , \ab[51][22] , \ab[51][21] ,
         \ab[51][20] , \ab[51][19] , \ab[51][18] , \ab[51][17] , \ab[51][16] ,
         \ab[51][15] , \ab[51][14] , \ab[51][13] , \ab[51][12] , \ab[51][11] ,
         \ab[51][10] , \ab[51][9] , \ab[51][8] , \ab[51][7] , \ab[51][6] ,
         \ab[51][5] , \ab[51][4] , \ab[51][3] , \ab[51][2] , \ab[51][1] ,
         \ab[51][0] , \ab[50][52] , \ab[50][51] , \ab[50][50] , \ab[50][49] ,
         \ab[50][48] , \ab[50][47] , \ab[50][46] , \ab[50][45] , \ab[50][44] ,
         \ab[50][43] , \ab[50][42] , \ab[50][41] , \ab[50][40] , \ab[50][39] ,
         \ab[50][38] , \ab[50][37] , \ab[50][36] , \ab[50][35] , \ab[50][34] ,
         \ab[50][33] , \ab[50][32] , \ab[50][31] , \ab[50][30] , \ab[50][29] ,
         \ab[50][28] , \ab[50][27] , \ab[50][26] , \ab[50][25] , \ab[50][24] ,
         \ab[50][23] , \ab[50][22] , \ab[50][21] , \ab[50][20] , \ab[50][19] ,
         \ab[50][18] , \ab[50][17] , \ab[50][16] , \ab[50][15] , \ab[50][14] ,
         \ab[50][13] , \ab[50][12] , \ab[50][11] , \ab[50][10] , \ab[50][9] ,
         \ab[50][8] , \ab[50][7] , \ab[50][6] , \ab[50][5] , \ab[50][4] ,
         \ab[50][3] , \ab[50][2] , \ab[50][1] , \ab[50][0] , \ab[49][52] ,
         \ab[49][51] , \ab[49][50] , \ab[49][49] , \ab[49][48] , \ab[49][47] ,
         \ab[49][46] , \ab[49][45] , \ab[49][44] , \ab[49][43] , \ab[49][42] ,
         \ab[49][41] , \ab[49][40] , \ab[49][39] , \ab[49][38] , \ab[49][37] ,
         \ab[49][36] , \ab[49][35] , \ab[49][34] , \ab[49][33] , \ab[49][32] ,
         \ab[49][31] , \ab[49][30] , \ab[49][29] , \ab[49][28] , \ab[49][27] ,
         \ab[49][26] , \ab[49][25] , \ab[49][24] , \ab[49][23] , \ab[49][22] ,
         \ab[49][21] , \ab[49][20] , \ab[49][19] , \ab[49][18] , \ab[49][17] ,
         \ab[49][16] , \ab[49][15] , \ab[49][14] , \ab[49][13] , \ab[49][12] ,
         \ab[49][11] , \ab[49][10] , \ab[49][9] , \ab[49][8] , \ab[49][7] ,
         \ab[49][6] , \ab[49][5] , \ab[49][4] , \ab[49][3] , \ab[49][2] ,
         \ab[49][1] , \ab[49][0] , \ab[48][52] , \ab[48][51] , \ab[48][50] ,
         \ab[48][49] , \ab[48][48] , \ab[48][47] , \ab[48][46] , \ab[48][45] ,
         \ab[48][44] , \ab[48][43] , \ab[48][42] , \ab[48][41] , \ab[48][40] ,
         \ab[48][39] , \ab[48][38] , \ab[48][37] , \ab[48][36] , \ab[48][35] ,
         \ab[48][34] , \ab[48][33] , \ab[48][32] , \ab[48][31] , \ab[48][30] ,
         \ab[48][29] , \ab[48][28] , \ab[48][27] , \ab[48][26] , \ab[48][25] ,
         \ab[48][24] , \ab[48][23] , \ab[48][22] , \ab[48][21] , \ab[48][20] ,
         \ab[48][19] , \ab[48][18] , \ab[48][17] , \ab[48][16] , \ab[48][15] ,
         \ab[48][14] , \ab[48][13] , \ab[48][12] , \ab[48][11] , \ab[48][10] ,
         \ab[48][9] , \ab[48][8] , \ab[48][7] , \ab[48][6] , \ab[48][5] ,
         \ab[48][4] , \ab[48][3] , \ab[48][2] , \ab[48][1] , \ab[48][0] ,
         \ab[47][52] , \ab[47][51] , \ab[47][50] , \ab[47][49] , \ab[47][48] ,
         \ab[47][47] , \ab[47][46] , \ab[47][45] , \ab[47][44] , \ab[47][43] ,
         \ab[47][42] , \ab[47][41] , \ab[47][40] , \ab[47][39] , \ab[47][38] ,
         \ab[47][37] , \ab[47][36] , \ab[47][35] , \ab[47][34] , \ab[47][33] ,
         \ab[47][32] , \ab[47][31] , \ab[47][30] , \ab[47][29] , \ab[47][28] ,
         \ab[47][27] , \ab[47][26] , \ab[47][25] , \ab[47][24] , \ab[47][23] ,
         \ab[47][22] , \ab[47][21] , \ab[47][20] , \ab[47][19] , \ab[47][18] ,
         \ab[47][17] , \ab[47][16] , \ab[47][15] , \ab[47][14] , \ab[47][13] ,
         \ab[47][12] , \ab[47][11] , \ab[47][10] , \ab[47][9] , \ab[47][8] ,
         \ab[47][7] , \ab[47][6] , \ab[47][5] , \ab[47][4] , \ab[47][3] ,
         \ab[47][2] , \ab[47][1] , \ab[47][0] , \ab[46][52] , \ab[46][51] ,
         \ab[46][50] , \ab[46][49] , \ab[46][48] , \ab[46][47] , \ab[46][46] ,
         \ab[46][45] , \ab[46][44] , \ab[46][43] , \ab[46][42] , \ab[46][41] ,
         \ab[46][40] , \ab[46][39] , \ab[46][38] , \ab[46][37] , \ab[46][36] ,
         \ab[46][35] , \ab[46][34] , \ab[46][33] , \ab[46][32] , \ab[46][31] ,
         \ab[46][30] , \ab[46][29] , \ab[46][28] , \ab[46][27] , \ab[46][26] ,
         \ab[46][25] , \ab[46][24] , \ab[46][23] , \ab[46][22] , \ab[46][21] ,
         \ab[46][20] , \ab[46][19] , \ab[46][18] , \ab[46][17] , \ab[46][16] ,
         \ab[46][15] , \ab[46][14] , \ab[46][13] , \ab[46][12] , \ab[46][11] ,
         \ab[46][10] , \ab[46][9] , \ab[46][8] , \ab[46][7] , \ab[46][6] ,
         \ab[46][5] , \ab[46][4] , \ab[46][3] , \ab[46][2] , \ab[46][1] ,
         \ab[46][0] , \ab[45][52] , \ab[45][51] , \ab[45][50] , \ab[45][49] ,
         \ab[45][48] , \ab[45][47] , \ab[45][46] , \ab[45][45] , \ab[45][44] ,
         \ab[45][43] , \ab[45][42] , \ab[45][41] , \ab[45][40] , \ab[45][39] ,
         \ab[45][38] , \ab[45][37] , \ab[45][36] , \ab[45][35] , \ab[45][34] ,
         \ab[45][33] , \ab[45][32] , \ab[45][31] , \ab[45][30] , \ab[45][29] ,
         \ab[45][28] , \ab[45][27] , \ab[45][26] , \ab[45][25] , \ab[45][24] ,
         \ab[45][23] , \ab[45][22] , \ab[45][21] , \ab[45][20] , \ab[45][19] ,
         \ab[45][18] , \ab[45][17] , \ab[45][16] , \ab[45][15] , \ab[45][14] ,
         \ab[45][13] , \ab[45][12] , \ab[45][11] , \ab[45][10] , \ab[45][9] ,
         \ab[45][8] , \ab[45][7] , \ab[45][6] , \ab[45][5] , \ab[45][4] ,
         \ab[45][3] , \ab[45][2] , \ab[45][1] , \ab[45][0] , \ab[44][52] ,
         \ab[44][51] , \ab[44][50] , \ab[44][49] , \ab[44][48] , \ab[44][47] ,
         \ab[44][46] , \ab[44][45] , \ab[44][44] , \ab[44][43] , \ab[44][42] ,
         \ab[44][41] , \ab[44][40] , \ab[44][39] , \ab[44][38] , \ab[44][37] ,
         \ab[44][36] , \ab[44][35] , \ab[44][34] , \ab[44][33] , \ab[44][32] ,
         \ab[44][31] , \ab[44][30] , \ab[44][29] , \ab[44][28] , \ab[44][27] ,
         \ab[44][26] , \ab[44][25] , \ab[44][24] , \ab[44][23] , \ab[44][22] ,
         \ab[44][21] , \ab[44][20] , \ab[44][19] , \ab[44][18] , \ab[44][17] ,
         \ab[44][16] , \ab[44][15] , \ab[44][14] , \ab[44][13] , \ab[44][12] ,
         \ab[44][11] , \ab[44][10] , \ab[44][9] , \ab[44][8] , \ab[44][7] ,
         \ab[44][6] , \ab[44][5] , \ab[44][4] , \ab[44][3] , \ab[44][2] ,
         \ab[44][1] , \ab[44][0] , \ab[43][52] , \ab[43][51] , \ab[43][50] ,
         \ab[43][49] , \ab[43][48] , \ab[43][47] , \ab[43][46] , \ab[43][45] ,
         \ab[43][44] , \ab[43][43] , \ab[43][42] , \ab[43][41] , \ab[43][40] ,
         \ab[43][39] , \ab[43][38] , \ab[43][37] , \ab[43][36] , \ab[43][35] ,
         \ab[43][34] , \ab[43][33] , \ab[43][32] , \ab[43][31] , \ab[43][30] ,
         \ab[43][29] , \ab[43][28] , \ab[43][27] , \ab[43][26] , \ab[43][25] ,
         \ab[43][24] , \ab[43][23] , \ab[43][22] , \ab[43][21] , \ab[43][20] ,
         \ab[43][19] , \ab[43][18] , \ab[43][17] , \ab[43][16] , \ab[43][15] ,
         \ab[43][14] , \ab[43][13] , \ab[43][12] , \ab[43][11] , \ab[43][10] ,
         \ab[43][9] , \ab[43][8] , \ab[43][7] , \ab[43][6] , \ab[43][5] ,
         \ab[43][4] , \ab[43][3] , \ab[43][2] , \ab[43][1] , \ab[43][0] ,
         \ab[42][52] , \ab[42][51] , \ab[42][50] , \ab[42][49] , \ab[42][48] ,
         \ab[42][47] , \ab[42][46] , \ab[42][45] , \ab[42][44] , \ab[42][43] ,
         \ab[42][42] , \ab[42][41] , \ab[42][40] , \ab[42][39] , \ab[42][38] ,
         \ab[42][37] , \ab[42][36] , \ab[42][35] , \ab[42][34] , \ab[42][33] ,
         \ab[42][32] , \ab[42][31] , \ab[42][30] , \ab[42][29] , \ab[42][28] ,
         \ab[42][27] , \ab[42][26] , \ab[42][25] , \ab[42][24] , \ab[42][23] ,
         \ab[42][22] , \ab[42][21] , \ab[42][20] , \ab[42][19] , \ab[42][18] ,
         \ab[42][17] , \ab[42][16] , \ab[42][15] , \ab[42][14] , \ab[42][13] ,
         \ab[42][12] , \ab[42][11] , \ab[42][10] , \ab[42][9] , \ab[42][8] ,
         \ab[42][7] , \ab[42][6] , \ab[42][5] , \ab[42][4] , \ab[42][3] ,
         \ab[42][2] , \ab[42][1] , \ab[42][0] , \ab[41][52] , \ab[41][51] ,
         \ab[41][50] , \ab[41][49] , \ab[41][48] , \ab[41][47] , \ab[41][46] ,
         \ab[41][45] , \ab[41][44] , \ab[41][43] , \ab[41][42] , \ab[41][41] ,
         \ab[41][40] , \ab[41][39] , \ab[41][38] , \ab[41][37] , \ab[41][36] ,
         \ab[41][35] , \ab[41][34] , \ab[41][33] , \ab[41][32] , \ab[41][31] ,
         \ab[41][30] , \ab[41][29] , \ab[41][28] , \ab[41][27] , \ab[41][26] ,
         \ab[41][25] , \ab[41][24] , \ab[41][23] , \ab[41][22] , \ab[41][21] ,
         \ab[41][20] , \ab[41][19] , \ab[41][18] , \ab[41][17] , \ab[41][16] ,
         \ab[41][15] , \ab[41][14] , \ab[41][13] , \ab[41][12] , \ab[41][11] ,
         \ab[41][10] , \ab[41][9] , \ab[41][8] , \ab[41][7] , \ab[41][6] ,
         \ab[41][5] , \ab[41][4] , \ab[41][3] , \ab[41][2] , \ab[41][1] ,
         \ab[41][0] , \ab[40][52] , \ab[40][51] , \ab[40][50] , \ab[40][49] ,
         \ab[40][48] , \ab[40][47] , \ab[40][46] , \ab[40][45] , \ab[40][44] ,
         \ab[40][43] , \ab[40][42] , \ab[40][41] , \ab[40][40] , \ab[40][39] ,
         \ab[40][38] , \ab[40][37] , \ab[40][36] , \ab[40][35] , \ab[40][34] ,
         \ab[40][33] , \ab[40][32] , \ab[40][31] , \ab[40][30] , \ab[40][29] ,
         \ab[40][28] , \ab[40][27] , \ab[40][26] , \ab[40][25] , \ab[40][24] ,
         \ab[40][23] , \ab[40][22] , \ab[40][21] , \ab[40][20] , \ab[40][19] ,
         \ab[40][18] , \ab[40][17] , \ab[40][16] , \ab[40][15] , \ab[40][14] ,
         \ab[40][13] , \ab[40][12] , \ab[40][11] , \ab[40][10] , \ab[40][9] ,
         \ab[40][8] , \ab[40][7] , \ab[40][6] , \ab[40][5] , \ab[40][4] ,
         \ab[40][3] , \ab[40][2] , \ab[40][1] , \ab[40][0] , \ab[39][52] ,
         \ab[39][51] , \ab[39][50] , \ab[39][49] , \ab[39][48] , \ab[39][47] ,
         \ab[39][46] , \ab[39][45] , \ab[39][44] , \ab[39][43] , \ab[39][42] ,
         \ab[39][41] , \ab[39][40] , \ab[39][39] , \ab[39][38] , \ab[39][37] ,
         \ab[39][36] , \ab[39][35] , \ab[39][34] , \ab[39][33] , \ab[39][32] ,
         \ab[39][31] , \ab[39][30] , \ab[39][29] , \ab[39][28] , \ab[39][27] ,
         \ab[39][26] , \ab[39][25] , \ab[39][24] , \ab[39][23] , \ab[39][22] ,
         \ab[39][21] , \ab[39][20] , \ab[39][19] , \ab[39][18] , \ab[39][17] ,
         \ab[39][16] , \ab[39][15] , \ab[39][14] , \ab[39][13] , \ab[39][12] ,
         \ab[39][11] , \ab[39][10] , \ab[39][9] , \ab[39][8] , \ab[39][7] ,
         \ab[39][6] , \ab[39][5] , \ab[39][4] , \ab[39][3] , \ab[39][2] ,
         \ab[39][1] , \ab[39][0] , \ab[38][52] , \ab[38][51] , \ab[38][50] ,
         \ab[38][49] , \ab[38][48] , \ab[38][47] , \ab[38][46] , \ab[38][45] ,
         \ab[38][44] , \ab[38][43] , \ab[38][42] , \ab[38][41] , \ab[38][40] ,
         \ab[38][39] , \ab[38][38] , \ab[38][37] , \ab[38][36] , \ab[38][35] ,
         \ab[38][34] , \ab[38][33] , \ab[38][32] , \ab[38][31] , \ab[38][30] ,
         \ab[38][29] , \ab[38][28] , \ab[38][27] , \ab[38][26] , \ab[38][25] ,
         \ab[38][24] , \ab[38][23] , \ab[38][22] , \ab[38][21] , \ab[38][20] ,
         \ab[38][19] , \ab[38][18] , \ab[38][17] , \ab[38][16] , \ab[38][15] ,
         \ab[38][14] , \ab[38][13] , \ab[38][12] , \ab[38][11] , \ab[38][10] ,
         \ab[38][9] , \ab[38][8] , \ab[38][7] , \ab[38][6] , \ab[38][5] ,
         \ab[38][4] , \ab[38][3] , \ab[38][2] , \ab[38][1] , \ab[38][0] ,
         \ab[37][52] , \ab[37][51] , \ab[37][50] , \ab[37][49] , \ab[37][48] ,
         \ab[37][47] , \ab[37][46] , \ab[37][45] , \ab[37][44] , \ab[37][43] ,
         \ab[37][42] , \ab[37][41] , \ab[37][40] , \ab[37][39] , \ab[37][38] ,
         \ab[37][37] , \ab[37][36] , \ab[37][35] , \ab[37][34] , \ab[37][33] ,
         \ab[37][32] , \ab[37][31] , \ab[37][30] , \ab[37][29] , \ab[37][28] ,
         \ab[37][27] , \ab[37][26] , \ab[37][25] , \ab[37][24] , \ab[37][23] ,
         \ab[37][22] , \ab[37][21] , \ab[37][20] , \ab[37][19] , \ab[37][18] ,
         \ab[37][17] , \ab[37][16] , \ab[37][15] , \ab[37][14] , \ab[37][13] ,
         \ab[37][12] , \ab[37][11] , \ab[37][10] , \ab[37][9] , \ab[37][8] ,
         \ab[37][7] , \ab[37][6] , \ab[37][5] , \ab[37][4] , \ab[37][3] ,
         \ab[37][2] , \ab[37][1] , \ab[37][0] , \ab[36][52] , \ab[36][51] ,
         \ab[36][50] , \ab[36][49] , \ab[36][48] , \ab[36][47] , \ab[36][46] ,
         \ab[36][45] , \ab[36][44] , \ab[36][43] , \ab[36][42] , \ab[36][41] ,
         \ab[36][40] , \ab[36][39] , \ab[36][38] , \ab[36][37] , \ab[36][36] ,
         \ab[36][35] , \ab[36][34] , \ab[36][33] , \ab[36][32] , \ab[36][31] ,
         \ab[36][30] , \ab[36][29] , \ab[36][28] , \ab[36][27] , \ab[36][26] ,
         \ab[36][25] , \ab[36][24] , \ab[36][23] , \ab[36][22] , \ab[36][21] ,
         \ab[36][20] , \ab[36][19] , \ab[36][18] , \ab[36][17] , \ab[36][16] ,
         \ab[36][15] , \ab[36][14] , \ab[36][13] , \ab[36][12] , \ab[36][11] ,
         \ab[36][10] , \ab[36][9] , \ab[36][8] , \ab[36][7] , \ab[36][6] ,
         \ab[36][5] , \ab[36][4] , \ab[36][3] , \ab[36][2] , \ab[36][1] ,
         \ab[36][0] , \ab[35][52] , \ab[35][51] , \ab[35][50] , \ab[35][49] ,
         \ab[35][48] , \ab[35][47] , \ab[35][46] , \ab[35][45] , \ab[35][44] ,
         \ab[35][43] , \ab[35][42] , \ab[35][41] , \ab[35][40] , \ab[35][39] ,
         \ab[35][38] , \ab[35][37] , \ab[35][36] , \ab[35][35] , \ab[35][34] ,
         \ab[35][33] , \ab[35][32] , \ab[35][31] , \ab[35][30] , \ab[35][29] ,
         \ab[35][28] , \ab[35][27] , \ab[35][26] , \ab[35][25] , \ab[35][24] ,
         \ab[35][23] , \ab[35][22] , \ab[35][21] , \ab[35][20] , \ab[35][19] ,
         \ab[35][18] , \ab[35][17] , \ab[35][16] , \ab[35][15] , \ab[35][14] ,
         \ab[35][13] , \ab[35][12] , \ab[35][11] , \ab[35][10] , \ab[35][9] ,
         \ab[35][8] , \ab[35][7] , \ab[35][6] , \ab[35][5] , \ab[35][4] ,
         \ab[35][3] , \ab[35][2] , \ab[35][1] , \ab[35][0] , \ab[34][52] ,
         \ab[34][51] , \ab[34][50] , \ab[34][49] , \ab[34][48] , \ab[34][47] ,
         \ab[34][46] , \ab[34][45] , \ab[34][44] , \ab[34][43] , \ab[34][42] ,
         \ab[34][41] , \ab[34][40] , \ab[34][39] , \ab[34][38] , \ab[34][37] ,
         \ab[34][36] , \ab[34][35] , \ab[34][34] , \ab[34][33] , \ab[34][32] ,
         \ab[34][31] , \ab[34][30] , \ab[34][29] , \ab[34][28] , \ab[34][27] ,
         \ab[34][26] , \ab[34][25] , \ab[34][24] , \ab[34][23] , \ab[34][22] ,
         \ab[34][21] , \ab[34][20] , \ab[34][19] , \ab[34][18] , \ab[34][17] ,
         \ab[34][16] , \ab[34][15] , \ab[34][14] , \ab[34][13] , \ab[34][12] ,
         \ab[34][11] , \ab[34][10] , \ab[34][9] , \ab[34][8] , \ab[34][7] ,
         \ab[34][6] , \ab[34][5] , \ab[34][4] , \ab[34][3] , \ab[34][2] ,
         \ab[34][1] , \ab[34][0] , \ab[33][52] , \ab[33][51] , \ab[33][50] ,
         \ab[33][49] , \ab[33][48] , \ab[33][47] , \ab[33][46] , \ab[33][45] ,
         \ab[33][44] , \ab[33][43] , \ab[33][42] , \ab[33][41] , \ab[33][40] ,
         \ab[33][39] , \ab[33][38] , \ab[33][37] , \ab[33][36] , \ab[33][35] ,
         \ab[33][34] , \ab[33][33] , \ab[33][32] , \ab[33][31] , \ab[33][30] ,
         \ab[33][29] , \ab[33][28] , \ab[33][27] , \ab[33][26] , \ab[33][25] ,
         \ab[33][24] , \ab[33][23] , \ab[33][22] , \ab[33][21] , \ab[33][20] ,
         \ab[33][19] , \ab[33][18] , \ab[33][17] , \ab[33][16] , \ab[33][15] ,
         \ab[33][14] , \ab[33][13] , \ab[33][12] , \ab[33][11] , \ab[33][10] ,
         \ab[33][9] , \ab[33][8] , \ab[33][7] , \ab[33][6] , \ab[33][5] ,
         \ab[33][4] , \ab[33][3] , \ab[33][2] , \ab[33][1] , \ab[33][0] ,
         \ab[32][52] , \ab[32][51] , \ab[32][50] , \ab[32][49] , \ab[32][48] ,
         \ab[32][47] , \ab[32][46] , \ab[32][45] , \ab[32][44] , \ab[32][43] ,
         \ab[32][42] , \ab[32][41] , \ab[32][40] , \ab[32][39] , \ab[32][38] ,
         \ab[32][37] , \ab[32][36] , \ab[32][35] , \ab[32][34] , \ab[32][33] ,
         \ab[32][32] , \ab[32][31] , \ab[32][30] , \ab[32][29] , \ab[32][28] ,
         \ab[32][27] , \ab[32][26] , \ab[32][25] , \ab[32][24] , \ab[32][23] ,
         \ab[32][22] , \ab[32][21] , \ab[32][20] , \ab[32][19] , \ab[32][18] ,
         \ab[32][17] , \ab[32][16] , \ab[32][15] , \ab[32][14] , \ab[32][13] ,
         \ab[32][12] , \ab[32][11] , \ab[32][10] , \ab[32][9] , \ab[32][8] ,
         \ab[32][7] , \ab[32][6] , \ab[32][5] , \ab[32][4] , \ab[32][3] ,
         \ab[32][2] , \ab[32][1] , \ab[32][0] , \ab[31][52] , \ab[31][51] ,
         \ab[31][50] , \ab[31][49] , \ab[31][48] , \ab[31][47] , \ab[31][46] ,
         \ab[31][45] , \ab[31][44] , \ab[31][43] , \ab[31][42] , \ab[31][41] ,
         \ab[31][40] , \ab[31][39] , \ab[31][38] , \ab[31][37] , \ab[31][36] ,
         \ab[31][35] , \ab[31][34] , \ab[31][33] , \ab[31][32] , \ab[31][31] ,
         \ab[31][30] , \ab[31][29] , \ab[31][28] , \ab[31][27] , \ab[31][26] ,
         \ab[31][25] , \ab[31][24] , \ab[31][23] , \ab[31][22] , \ab[31][21] ,
         \ab[31][20] , \ab[31][19] , \ab[31][18] , \ab[31][17] , \ab[31][16] ,
         \ab[31][15] , \ab[31][14] , \ab[31][13] , \ab[31][12] , \ab[31][11] ,
         \ab[31][10] , \ab[31][9] , \ab[31][8] , \ab[31][7] , \ab[31][6] ,
         \ab[31][5] , \ab[31][4] , \ab[31][3] , \ab[31][2] , \ab[31][1] ,
         \ab[31][0] , \ab[30][52] , \ab[30][51] , \ab[30][50] , \ab[30][49] ,
         \ab[30][48] , \ab[30][47] , \ab[30][46] , \ab[30][45] , \ab[30][44] ,
         \ab[30][43] , \ab[30][42] , \ab[30][41] , \ab[30][40] , \ab[30][39] ,
         \ab[30][38] , \ab[30][37] , \ab[30][36] , \ab[30][35] , \ab[30][34] ,
         \ab[30][33] , \ab[30][32] , \ab[30][31] , \ab[30][30] , \ab[30][29] ,
         \ab[30][28] , \ab[30][27] , \ab[30][26] , \ab[30][25] , \ab[30][24] ,
         \ab[30][23] , \ab[30][22] , \ab[30][21] , \ab[30][20] , \ab[30][19] ,
         \ab[30][18] , \ab[30][17] , \ab[30][16] , \ab[30][15] , \ab[30][14] ,
         \ab[30][13] , \ab[30][12] , \ab[30][11] , \ab[30][10] , \ab[30][9] ,
         \ab[30][8] , \ab[30][7] , \ab[30][6] , \ab[30][5] , \ab[30][4] ,
         \ab[30][3] , \ab[30][2] , \ab[30][1] , \ab[30][0] , \ab[29][52] ,
         \ab[29][51] , \ab[29][50] , \ab[29][49] , \ab[29][48] , \ab[29][47] ,
         \ab[29][46] , \ab[29][45] , \ab[29][44] , \ab[29][43] , \ab[29][42] ,
         \ab[29][41] , \ab[29][40] , \ab[29][39] , \ab[29][38] , \ab[29][37] ,
         \ab[29][36] , \ab[29][35] , \ab[29][34] , \ab[29][33] , \ab[29][32] ,
         \ab[29][31] , \ab[29][30] , \ab[29][29] , \ab[29][28] , \ab[29][27] ,
         \ab[29][26] , \ab[29][25] , \ab[29][24] , \ab[29][23] , \ab[29][22] ,
         \ab[29][21] , \ab[29][20] , \ab[29][19] , \ab[29][18] , \ab[29][17] ,
         \ab[29][16] , \ab[29][15] , \ab[29][14] , \ab[29][13] , \ab[29][12] ,
         \ab[29][11] , \ab[29][10] , \ab[29][9] , \ab[29][8] , \ab[29][7] ,
         \ab[29][6] , \ab[29][5] , \ab[29][4] , \ab[29][3] , \ab[29][2] ,
         \ab[29][1] , \ab[29][0] , \ab[28][52] , \ab[28][51] , \ab[28][50] ,
         \ab[28][49] , \ab[28][48] , \ab[28][47] , \ab[28][46] , \ab[28][45] ,
         \ab[28][44] , \ab[28][43] , \ab[28][42] , \ab[28][41] , \ab[28][40] ,
         \ab[28][39] , \ab[28][38] , \ab[28][37] , \ab[28][36] , \ab[28][35] ,
         \ab[28][34] , \ab[28][33] , \ab[28][32] , \ab[28][31] , \ab[28][30] ,
         \ab[28][29] , \ab[28][28] , \ab[28][27] , \ab[28][26] , \ab[28][25] ,
         \ab[28][24] , \ab[28][23] , \ab[28][22] , \ab[28][21] , \ab[28][20] ,
         \ab[28][19] , \ab[28][18] , \ab[28][17] , \ab[28][16] , \ab[28][15] ,
         \ab[28][14] , \ab[28][13] , \ab[28][12] , \ab[28][11] , \ab[28][10] ,
         \ab[28][9] , \ab[28][8] , \ab[28][7] , \ab[28][6] , \ab[28][5] ,
         \ab[28][4] , \ab[28][3] , \ab[28][2] , \ab[28][1] , \ab[28][0] ,
         \ab[27][52] , \ab[27][51] , \ab[27][50] , \ab[27][49] , \ab[27][48] ,
         \ab[27][47] , \ab[27][46] , \ab[27][45] , \ab[27][44] , \ab[27][43] ,
         \ab[27][42] , \ab[27][41] , \ab[27][40] , \ab[27][39] , \ab[27][38] ,
         \ab[27][37] , \ab[27][36] , \ab[27][35] , \ab[27][34] , \ab[27][33] ,
         \ab[27][32] , \ab[27][31] , \ab[27][30] , \ab[27][29] , \ab[27][28] ,
         \ab[27][27] , \ab[27][26] , \ab[27][25] , \ab[27][24] , \ab[27][23] ,
         \ab[27][22] , \ab[27][21] , \ab[27][20] , \ab[27][19] , \ab[27][18] ,
         \ab[27][17] , \ab[27][16] , \ab[27][15] , \ab[27][14] , \ab[27][13] ,
         \ab[27][12] , \ab[27][11] , \ab[27][10] , \ab[27][9] , \ab[27][8] ,
         \ab[27][7] , \ab[27][6] , \ab[27][5] , \ab[27][4] , \ab[27][3] ,
         \ab[27][2] , \ab[27][1] , \ab[27][0] , \ab[26][52] , \ab[26][51] ,
         \ab[26][50] , \ab[26][49] , \ab[26][48] , \ab[26][47] , \ab[26][46] ,
         \ab[26][45] , \ab[26][44] , \ab[26][43] , \ab[26][42] , \ab[26][41] ,
         \ab[26][40] , \ab[26][39] , \ab[26][38] , \ab[26][37] , \ab[26][36] ,
         \ab[26][35] , \ab[26][34] , \ab[26][33] , \ab[26][32] , \ab[26][31] ,
         \ab[26][30] , \ab[26][29] , \ab[26][28] , \ab[26][27] , \ab[26][26] ,
         \ab[26][25] , \ab[26][24] , \ab[26][23] , \ab[26][22] , \ab[26][21] ,
         \ab[26][20] , \ab[26][19] , \ab[26][18] , \ab[26][17] , \ab[26][16] ,
         \ab[26][15] , \ab[26][14] , \ab[26][13] , \ab[26][12] , \ab[26][11] ,
         \ab[26][10] , \ab[26][9] , \ab[26][8] , \ab[26][7] , \ab[26][6] ,
         \ab[26][5] , \ab[26][4] , \ab[26][3] , \ab[26][2] , \ab[26][1] ,
         \ab[26][0] , \ab[25][52] , \ab[25][51] , \ab[25][50] , \ab[25][49] ,
         \ab[25][48] , \ab[25][47] , \ab[25][46] , \ab[25][45] , \ab[25][44] ,
         \ab[25][43] , \ab[25][42] , \ab[25][41] , \ab[25][40] , \ab[25][39] ,
         \ab[25][38] , \ab[25][37] , \ab[25][36] , \ab[25][35] , \ab[25][34] ,
         \ab[25][33] , \ab[25][32] , \ab[25][31] , \ab[25][30] , \ab[25][29] ,
         \ab[25][28] , \ab[25][27] , \ab[25][26] , \ab[25][25] , \ab[25][24] ,
         \ab[25][23] , \ab[25][22] , \ab[25][21] , \ab[25][20] , \ab[25][19] ,
         \ab[25][18] , \ab[25][17] , \ab[25][16] , \ab[25][15] , \ab[25][14] ,
         \ab[25][13] , \ab[25][12] , \ab[25][11] , \ab[25][10] , \ab[25][9] ,
         \ab[25][8] , \ab[25][7] , \ab[25][6] , \ab[25][5] , \ab[25][4] ,
         \ab[25][3] , \ab[25][2] , \ab[25][1] , \ab[25][0] , \ab[24][52] ,
         \ab[24][51] , \ab[24][50] , \ab[24][49] , \ab[24][48] , \ab[24][47] ,
         \ab[24][46] , \ab[24][45] , \ab[24][44] , \ab[24][43] , \ab[24][42] ,
         \ab[24][41] , \ab[24][40] , \ab[24][39] , \ab[24][38] , \ab[24][37] ,
         \ab[24][36] , \ab[24][35] , \ab[24][34] , \ab[24][33] , \ab[24][32] ,
         \ab[24][31] , \ab[24][30] , \ab[24][29] , \ab[24][28] , \ab[24][27] ,
         \ab[24][26] , \ab[24][25] , \ab[24][24] , \ab[24][23] , \ab[24][22] ,
         \ab[24][21] , \ab[24][20] , \ab[24][19] , \ab[24][18] , \ab[24][17] ,
         \ab[24][16] , \ab[24][15] , \ab[24][14] , \ab[24][13] , \ab[24][12] ,
         \ab[24][11] , \ab[24][10] , \ab[24][9] , \ab[24][8] , \ab[24][7] ,
         \ab[24][6] , \ab[24][5] , \ab[24][4] , \ab[24][3] , \ab[24][2] ,
         \ab[24][1] , \ab[24][0] , \ab[23][52] , \ab[23][51] , \ab[23][50] ,
         \ab[23][49] , \ab[23][48] , \ab[23][47] , \ab[23][46] , \ab[23][45] ,
         \ab[23][44] , \ab[23][43] , \ab[23][42] , \ab[23][41] , \ab[23][40] ,
         \ab[23][39] , \ab[23][38] , \ab[23][37] , \ab[23][36] , \ab[23][35] ,
         \ab[23][34] , \ab[23][33] , \ab[23][32] , \ab[23][31] , \ab[23][30] ,
         \ab[23][29] , \ab[23][28] , \ab[23][27] , \ab[23][26] , \ab[23][25] ,
         \ab[23][24] , \ab[23][23] , \ab[23][22] , \ab[23][21] , \ab[23][20] ,
         \ab[23][19] , \ab[23][18] , \ab[23][17] , \ab[23][16] , \ab[23][15] ,
         \ab[23][14] , \ab[23][13] , \ab[23][12] , \ab[23][11] , \ab[23][10] ,
         \ab[23][9] , \ab[23][8] , \ab[23][7] , \ab[23][6] , \ab[23][5] ,
         \ab[23][4] , \ab[23][3] , \ab[23][2] , \ab[23][1] , \ab[23][0] ,
         \ab[22][52] , \ab[22][51] , \ab[22][50] , \ab[22][49] , \ab[22][48] ,
         \ab[22][47] , \ab[22][46] , \ab[22][45] , \ab[22][44] , \ab[22][43] ,
         \ab[22][42] , \ab[22][41] , \ab[22][40] , \ab[22][39] , \ab[22][38] ,
         \ab[22][37] , \ab[22][36] , \ab[22][35] , \ab[22][34] , \ab[22][33] ,
         \ab[22][32] , \ab[22][31] , \ab[22][30] , \ab[22][29] , \ab[22][28] ,
         \ab[22][27] , \ab[22][26] , \ab[22][25] , \ab[22][24] , \ab[22][23] ,
         \ab[22][22] , \ab[22][21] , \ab[22][20] , \ab[22][19] , \ab[22][18] ,
         \ab[22][17] , \ab[22][16] , \ab[22][15] , \ab[22][14] , \ab[22][13] ,
         \ab[22][12] , \ab[22][11] , \ab[22][10] , \ab[22][9] , \ab[22][8] ,
         \ab[22][7] , \ab[22][6] , \ab[22][5] , \ab[22][4] , \ab[22][3] ,
         \ab[22][2] , \ab[22][1] , \ab[22][0] , \ab[21][52] , \ab[21][51] ,
         \ab[21][50] , \ab[21][49] , \ab[21][48] , \ab[21][47] , \ab[21][46] ,
         \ab[21][45] , \ab[21][44] , \ab[21][43] , \ab[21][42] , \ab[21][41] ,
         \ab[21][40] , \ab[21][39] , \ab[21][38] , \ab[21][37] , \ab[21][36] ,
         \ab[21][35] , \ab[21][34] , \ab[21][33] , \ab[21][32] , \ab[21][31] ,
         \ab[21][30] , \ab[21][29] , \ab[21][28] , \ab[21][27] , \ab[21][26] ,
         \ab[21][25] , \ab[21][24] , \ab[21][23] , \ab[21][22] , \ab[21][21] ,
         \ab[21][20] , \ab[21][19] , \ab[21][18] , \ab[21][17] , \ab[21][16] ,
         \ab[21][15] , \ab[21][14] , \ab[21][13] , \ab[21][12] , \ab[21][11] ,
         \ab[21][10] , \ab[21][9] , \ab[21][8] , \ab[21][7] , \ab[21][6] ,
         \ab[21][5] , \ab[21][4] , \ab[21][3] , \ab[21][2] , \ab[21][1] ,
         \ab[21][0] , \ab[20][52] , \ab[20][51] , \ab[20][50] , \ab[20][49] ,
         \ab[20][48] , \ab[20][47] , \ab[20][46] , \ab[20][45] , \ab[20][44] ,
         \ab[20][43] , \ab[20][42] , \ab[20][41] , \ab[20][40] , \ab[20][39] ,
         \ab[20][38] , \ab[20][37] , \ab[20][36] , \ab[20][35] , \ab[20][34] ,
         \ab[20][33] , \ab[20][32] , \ab[20][31] , \ab[20][30] , \ab[20][29] ,
         \ab[20][28] , \ab[20][27] , \ab[20][26] , \ab[20][25] , \ab[20][24] ,
         \ab[20][23] , \ab[20][22] , \ab[20][21] , \ab[20][20] , \ab[20][19] ,
         \ab[20][18] , \ab[20][17] , \ab[20][16] , \ab[20][15] , \ab[20][14] ,
         \ab[20][13] , \ab[20][12] , \ab[20][11] , \ab[20][10] , \ab[20][9] ,
         \ab[20][8] , \ab[20][7] , \ab[20][6] , \ab[20][5] , \ab[20][4] ,
         \ab[20][3] , \ab[20][2] , \ab[20][1] , \ab[20][0] , \ab[19][52] ,
         \ab[19][51] , \ab[19][50] , \ab[19][49] , \ab[19][48] , \ab[19][47] ,
         \ab[19][46] , \ab[19][45] , \ab[19][44] , \ab[19][43] , \ab[19][42] ,
         \ab[19][41] , \ab[19][40] , \ab[19][39] , \ab[19][38] , \ab[19][37] ,
         \ab[19][36] , \ab[19][35] , \ab[19][34] , \ab[19][33] , \ab[19][32] ,
         \ab[19][31] , \ab[19][30] , \ab[19][29] , \ab[19][28] , \ab[19][27] ,
         \ab[19][26] , \ab[19][25] , \ab[19][24] , \ab[19][23] , \ab[19][22] ,
         \ab[19][21] , \ab[19][20] , \ab[19][19] , \ab[19][18] , \ab[19][17] ,
         \ab[19][16] , \ab[19][15] , \ab[19][14] , \ab[19][13] , \ab[19][12] ,
         \ab[19][11] , \ab[19][10] , \ab[19][9] , \ab[19][8] , \ab[19][7] ,
         \ab[19][6] , \ab[19][5] , \ab[19][4] , \ab[19][3] , \ab[19][2] ,
         \ab[19][1] , \ab[19][0] , \ab[18][52] , \ab[18][51] , \ab[18][50] ,
         \ab[18][49] , \ab[18][48] , \ab[18][47] , \ab[18][46] , \ab[18][45] ,
         \ab[18][44] , \ab[18][43] , \ab[18][42] , \ab[18][41] , \ab[18][40] ,
         \ab[18][39] , \ab[18][38] , \ab[18][37] , \ab[18][36] , \ab[18][35] ,
         \ab[18][34] , \ab[18][33] , \ab[18][32] , \ab[18][31] , \ab[18][30] ,
         \ab[18][29] , \ab[18][28] , \ab[18][27] , \ab[18][26] , \ab[18][25] ,
         \ab[18][24] , \ab[18][23] , \ab[18][22] , \ab[18][21] , \ab[18][20] ,
         \ab[18][19] , \ab[18][18] , \ab[18][17] , \ab[18][16] , \ab[18][15] ,
         \ab[18][14] , \ab[18][13] , \ab[18][12] , \ab[18][11] , \ab[18][10] ,
         \ab[18][9] , \ab[18][8] , \ab[18][7] , \ab[18][6] , \ab[18][5] ,
         \ab[18][4] , \ab[18][3] , \ab[18][2] , \ab[18][1] , \ab[18][0] ,
         \ab[17][52] , \ab[17][51] , \ab[17][50] , \ab[17][49] , \ab[17][48] ,
         \ab[17][47] , \ab[17][46] , \ab[17][45] , \ab[17][44] , \ab[17][43] ,
         \ab[17][42] , \ab[17][41] , \ab[17][40] , \ab[17][39] , \ab[17][38] ,
         \ab[17][37] , \ab[17][36] , \ab[17][35] , \ab[17][34] , \ab[17][33] ,
         \ab[17][32] , \ab[17][31] , \ab[17][30] , \ab[17][29] , \ab[17][28] ,
         \ab[17][27] , \ab[17][26] , \ab[17][25] , \ab[17][24] , \ab[17][23] ,
         \ab[17][22] , \ab[17][21] , \ab[17][20] , \ab[17][19] , \ab[17][18] ,
         \ab[17][17] , \ab[17][16] , \ab[17][15] , \ab[17][14] , \ab[17][13] ,
         \ab[17][12] , \ab[17][11] , \ab[17][10] , \ab[17][9] , \ab[17][8] ,
         \ab[17][7] , \ab[17][6] , \ab[17][5] , \ab[17][4] , \ab[17][3] ,
         \ab[17][2] , \ab[17][1] , \ab[17][0] , \ab[16][52] , \ab[16][51] ,
         \ab[16][50] , \ab[16][49] , \ab[16][48] , \ab[16][47] , \ab[16][46] ,
         \ab[16][45] , \ab[16][44] , \ab[16][43] , \ab[16][42] , \ab[16][41] ,
         \ab[16][40] , \ab[16][39] , \ab[16][38] , \ab[16][37] , \ab[16][36] ,
         \ab[16][35] , \ab[16][34] , \ab[16][33] , \ab[16][32] , \ab[16][31] ,
         \ab[16][30] , \ab[16][29] , \ab[16][28] , \ab[16][27] , \ab[16][26] ,
         \ab[16][25] , \ab[16][24] , \ab[16][23] , \ab[16][22] , \ab[16][21] ,
         \ab[16][20] , \ab[16][19] , \ab[16][18] , \ab[16][17] , \ab[16][16] ,
         \ab[16][15] , \ab[16][14] , \ab[16][13] , \ab[16][12] , \ab[16][11] ,
         \ab[16][10] , \ab[16][9] , \ab[16][8] , \ab[16][7] , \ab[16][6] ,
         \ab[16][5] , \ab[16][4] , \ab[16][3] , \ab[16][2] , \ab[16][1] ,
         \ab[16][0] , \ab[15][52] , \ab[15][51] , \ab[15][50] , \ab[15][49] ,
         \ab[15][48] , \ab[15][47] , \ab[15][46] , \ab[15][45] , \ab[15][44] ,
         \ab[15][43] , \ab[15][42] , \ab[15][41] , \ab[15][40] , \ab[15][39] ,
         \ab[15][38] , \ab[15][37] , \ab[15][36] , \ab[15][35] , \ab[15][34] ,
         \ab[15][33] , \ab[15][32] , \ab[15][31] , \ab[15][30] , \ab[15][29] ,
         \ab[15][28] , \ab[15][27] , \ab[15][26] , \ab[15][25] , \ab[15][24] ,
         \ab[15][23] , \ab[15][22] , \ab[15][21] , \ab[15][20] , \ab[15][19] ,
         \ab[15][18] , \ab[15][17] , \ab[15][16] , \ab[15][15] , \ab[15][14] ,
         \ab[15][13] , \ab[15][12] , \ab[15][11] , \ab[15][10] , \ab[15][9] ,
         \ab[15][8] , \ab[15][7] , \ab[15][6] , \ab[15][5] , \ab[15][4] ,
         \ab[15][3] , \ab[15][2] , \ab[15][1] , \ab[15][0] , \ab[14][52] ,
         \ab[14][51] , \ab[14][50] , \ab[14][49] , \ab[14][48] , \ab[14][47] ,
         \ab[14][46] , \ab[14][45] , \ab[14][44] , \ab[14][43] , \ab[14][42] ,
         \ab[14][41] , \ab[14][40] , \ab[14][39] , \ab[14][38] , \ab[14][37] ,
         \ab[14][36] , \ab[14][35] , \ab[14][34] , \ab[14][33] , \ab[14][32] ,
         \ab[14][31] , \ab[14][30] , \ab[14][29] , \ab[14][28] , \ab[14][27] ,
         \ab[14][26] , \ab[14][25] , \ab[14][24] , \ab[14][23] , \ab[14][22] ,
         \ab[14][21] , \ab[14][20] , \ab[14][19] , \ab[14][18] , \ab[14][17] ,
         \ab[14][16] , \ab[14][15] , \ab[14][14] , \ab[14][13] , \ab[14][12] ,
         \ab[14][11] , \ab[14][10] , \ab[14][9] , \ab[14][8] , \ab[14][7] ,
         \ab[14][6] , \ab[14][5] , \ab[14][4] , \ab[14][3] , \ab[14][2] ,
         \ab[14][1] , \ab[14][0] , \ab[13][52] , \ab[13][51] , \ab[13][50] ,
         \ab[13][49] , \ab[13][48] , \ab[13][47] , \ab[13][46] , \ab[13][45] ,
         \ab[13][44] , \ab[13][43] , \ab[13][42] , \ab[13][41] , \ab[13][40] ,
         \ab[13][39] , \ab[13][38] , \ab[13][37] , \ab[13][36] , \ab[13][35] ,
         \ab[13][34] , \ab[13][33] , \ab[13][32] , \ab[13][31] , \ab[13][30] ,
         \ab[13][29] , \ab[13][28] , \ab[13][27] , \ab[13][26] , \ab[13][25] ,
         \ab[13][24] , \ab[13][23] , \ab[13][22] , \ab[13][21] , \ab[13][20] ,
         \ab[13][19] , \ab[13][18] , \ab[13][17] , \ab[13][16] , \ab[13][15] ,
         \ab[13][14] , \ab[13][13] , \ab[13][12] , \ab[13][11] , \ab[13][10] ,
         \ab[13][9] , \ab[13][8] , \ab[13][7] , \ab[13][6] , \ab[13][5] ,
         \ab[13][4] , \ab[13][3] , \ab[13][2] , \ab[13][1] , \ab[13][0] ,
         \ab[12][52] , \ab[12][51] , \ab[12][50] , \ab[12][49] , \ab[12][48] ,
         \ab[12][47] , \ab[12][46] , \ab[12][45] , \ab[12][44] , \ab[12][43] ,
         \ab[12][42] , \ab[12][41] , \ab[12][40] , \ab[12][39] , \ab[12][38] ,
         \ab[12][37] , \ab[12][36] , \ab[12][35] , \ab[12][34] , \ab[12][33] ,
         \ab[12][32] , \ab[12][31] , \ab[12][30] , \ab[12][29] , \ab[12][28] ,
         \ab[12][27] , \ab[12][26] , \ab[12][25] , \ab[12][24] , \ab[12][23] ,
         \ab[12][22] , \ab[12][21] , \ab[12][20] , \ab[12][19] , \ab[12][18] ,
         \ab[12][17] , \ab[12][16] , \ab[12][15] , \ab[12][14] , \ab[12][13] ,
         \ab[12][12] , \ab[12][11] , \ab[12][10] , \ab[12][9] , \ab[12][8] ,
         \ab[12][7] , \ab[12][6] , \ab[12][5] , \ab[12][4] , \ab[12][3] ,
         \ab[12][2] , \ab[12][1] , \ab[12][0] , \ab[11][52] , \ab[11][51] ,
         \ab[11][50] , \ab[11][49] , \ab[11][48] , \ab[11][47] , \ab[11][46] ,
         \ab[11][45] , \ab[11][44] , \ab[11][43] , \ab[11][42] , \ab[11][41] ,
         \ab[11][40] , \ab[11][39] , \ab[11][38] , \ab[11][37] , \ab[11][36] ,
         \ab[11][35] , \ab[11][34] , \ab[11][33] , \ab[11][32] , \ab[11][31] ,
         \ab[11][30] , \ab[11][29] , \ab[11][28] , \ab[11][27] , \ab[11][26] ,
         \ab[11][25] , \ab[11][24] , \ab[11][23] , \ab[11][22] , \ab[11][21] ,
         \ab[11][20] , \ab[11][19] , \ab[11][18] , \ab[11][17] , \ab[11][16] ,
         \ab[11][15] , \ab[11][14] , \ab[11][13] , \ab[11][12] , \ab[11][11] ,
         \ab[11][10] , \ab[11][9] , \ab[11][8] , \ab[11][7] , \ab[11][6] ,
         \ab[11][5] , \ab[11][4] , \ab[11][3] , \ab[11][2] , \ab[11][1] ,
         \ab[11][0] , \ab[10][52] , \ab[10][51] , \ab[10][50] , \ab[10][49] ,
         \ab[10][48] , \ab[10][47] , \ab[10][46] , \ab[10][45] , \ab[10][44] ,
         \ab[10][43] , \ab[10][42] , \ab[10][41] , \ab[10][40] , \ab[10][39] ,
         \ab[10][38] , \ab[10][37] , \ab[10][36] , \ab[10][35] , \ab[10][34] ,
         \ab[10][33] , \ab[10][32] , \ab[10][31] , \ab[10][30] , \ab[10][29] ,
         \ab[10][28] , \ab[10][27] , \ab[10][26] , \ab[10][25] , \ab[10][24] ,
         \ab[10][23] , \ab[10][22] , \ab[10][21] , \ab[10][20] , \ab[10][19] ,
         \ab[10][18] , \ab[10][17] , \ab[10][16] , \ab[10][15] , \ab[10][14] ,
         \ab[10][13] , \ab[10][12] , \ab[10][11] , \ab[10][10] , \ab[10][9] ,
         \ab[10][8] , \ab[10][7] , \ab[10][6] , \ab[10][5] , \ab[10][4] ,
         \ab[10][3] , \ab[10][2] , \ab[10][1] , \ab[10][0] , \ab[9][52] ,
         \ab[9][51] , \ab[9][50] , \ab[9][49] , \ab[9][48] , \ab[9][47] ,
         \ab[9][46] , \ab[9][45] , \ab[9][44] , \ab[9][43] , \ab[9][42] ,
         \ab[9][41] , \ab[9][40] , \ab[9][39] , \ab[9][38] , \ab[9][37] ,
         \ab[9][36] , \ab[9][35] , \ab[9][34] , \ab[9][33] , \ab[9][32] ,
         \ab[9][31] , \ab[9][30] , \ab[9][29] , \ab[9][28] , \ab[9][27] ,
         \ab[9][26] , \ab[9][25] , \ab[9][24] , \ab[9][23] , \ab[9][22] ,
         \ab[9][21] , \ab[9][20] , \ab[9][19] , \ab[9][18] , \ab[9][17] ,
         \ab[9][16] , \ab[9][15] , \ab[9][14] , \ab[9][13] , \ab[9][12] ,
         \ab[9][11] , \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] ,
         \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] ,
         \ab[9][1] , \ab[9][0] , \ab[8][52] , \ab[8][51] , \ab[8][50] ,
         \ab[8][49] , \ab[8][48] , \ab[8][47] , \ab[8][46] , \ab[8][45] ,
         \ab[8][44] , \ab[8][43] , \ab[8][42] , \ab[8][41] , \ab[8][40] ,
         \ab[8][39] , \ab[8][38] , \ab[8][37] , \ab[8][36] , \ab[8][35] ,
         \ab[8][34] , \ab[8][33] , \ab[8][32] , \ab[8][31] , \ab[8][30] ,
         \ab[8][29] , \ab[8][28] , \ab[8][27] , \ab[8][26] , \ab[8][25] ,
         \ab[8][24] , \ab[8][23] , \ab[8][22] , \ab[8][21] , \ab[8][20] ,
         \ab[8][19] , \ab[8][18] , \ab[8][17] , \ab[8][16] , \ab[8][15] ,
         \ab[8][14] , \ab[8][13] , \ab[8][12] , \ab[8][11] , \ab[8][10] ,
         \ab[8][9] , \ab[8][8] , \ab[8][7] , \ab[8][6] , \ab[8][5] ,
         \ab[8][4] , \ab[8][3] , \ab[8][2] , \ab[8][1] , \ab[8][0] ,
         \ab[7][52] , \ab[7][51] , \ab[7][50] , \ab[7][49] , \ab[7][48] ,
         \ab[7][47] , \ab[7][46] , \ab[7][45] , \ab[7][44] , \ab[7][43] ,
         \ab[7][42] , \ab[7][41] , \ab[7][40] , \ab[7][39] , \ab[7][38] ,
         \ab[7][37] , \ab[7][36] , \ab[7][35] , \ab[7][34] , \ab[7][33] ,
         \ab[7][32] , \ab[7][31] , \ab[7][30] , \ab[7][29] , \ab[7][28] ,
         \ab[7][27] , \ab[7][26] , \ab[7][25] , \ab[7][24] , \ab[7][23] ,
         \ab[7][22] , \ab[7][21] , \ab[7][20] , \ab[7][19] , \ab[7][18] ,
         \ab[7][17] , \ab[7][16] , \ab[7][15] , \ab[7][14] , \ab[7][13] ,
         \ab[7][12] , \ab[7][11] , \ab[7][10] , \ab[7][9] , \ab[7][8] ,
         \ab[7][7] , \ab[7][6] , \ab[7][5] , \ab[7][4] , \ab[7][3] ,
         \ab[7][2] , \ab[7][1] , \ab[7][0] , \ab[6][52] , \ab[6][51] ,
         \ab[6][50] , \ab[6][49] , \ab[6][48] , \ab[6][47] , \ab[6][46] ,
         \ab[6][45] , \ab[6][44] , \ab[6][43] , \ab[6][42] , \ab[6][41] ,
         \ab[6][40] , \ab[6][39] , \ab[6][38] , \ab[6][37] , \ab[6][36] ,
         \ab[6][35] , \ab[6][34] , \ab[6][33] , \ab[6][32] , \ab[6][31] ,
         \ab[6][30] , \ab[6][29] , \ab[6][28] , \ab[6][27] , \ab[6][26] ,
         \ab[6][25] , \ab[6][24] , \ab[6][23] , \ab[6][22] , \ab[6][21] ,
         \ab[6][20] , \ab[6][19] , \ab[6][18] , \ab[6][17] , \ab[6][16] ,
         \ab[6][15] , \ab[6][14] , \ab[6][13] , \ab[6][12] , \ab[6][11] ,
         \ab[6][10] , \ab[6][9] , \ab[6][8] , \ab[6][7] , \ab[6][6] ,
         \ab[6][5] , \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] ,
         \ab[6][0] , \ab[5][52] , \ab[5][51] , \ab[5][50] , \ab[5][49] ,
         \ab[5][48] , \ab[5][47] , \ab[5][46] , \ab[5][45] , \ab[5][44] ,
         \ab[5][43] , \ab[5][42] , \ab[5][41] , \ab[5][40] , \ab[5][39] ,
         \ab[5][38] , \ab[5][37] , \ab[5][36] , \ab[5][35] , \ab[5][34] ,
         \ab[5][33] , \ab[5][32] , \ab[5][31] , \ab[5][30] , \ab[5][29] ,
         \ab[5][28] , \ab[5][27] , \ab[5][26] , \ab[5][25] , \ab[5][24] ,
         \ab[5][23] , \ab[5][22] , \ab[5][21] , \ab[5][20] , \ab[5][19] ,
         \ab[5][18] , \ab[5][17] , \ab[5][16] , \ab[5][15] , \ab[5][14] ,
         \ab[5][13] , \ab[5][12] , \ab[5][11] , \ab[5][10] , \ab[5][9] ,
         \ab[5][8] , \ab[5][7] , \ab[5][6] , \ab[5][5] , \ab[5][4] ,
         \ab[5][3] , \ab[5][2] , \ab[5][1] , \ab[5][0] , \ab[4][52] ,
         \ab[4][51] , \ab[4][50] , \ab[4][49] , \ab[4][48] , \ab[4][47] ,
         \ab[4][46] , \ab[4][45] , \ab[4][44] , \ab[4][43] , \ab[4][42] ,
         \ab[4][41] , \ab[4][40] , \ab[4][39] , \ab[4][38] , \ab[4][37] ,
         \ab[4][36] , \ab[4][35] , \ab[4][34] , \ab[4][33] , \ab[4][32] ,
         \ab[4][31] , \ab[4][30] , \ab[4][29] , \ab[4][28] , \ab[4][27] ,
         \ab[4][26] , \ab[4][25] , \ab[4][24] , \ab[4][23] , \ab[4][22] ,
         \ab[4][21] , \ab[4][20] , \ab[4][19] , \ab[4][18] , \ab[4][17] ,
         \ab[4][16] , \ab[4][15] , \ab[4][14] , \ab[4][13] , \ab[4][12] ,
         \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] ,
         \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] ,
         \ab[4][1] , \ab[4][0] , \ab[3][52] , \ab[3][51] , \ab[3][50] ,
         \ab[3][49] , \ab[3][48] , \ab[3][47] , \ab[3][46] , \ab[3][45] ,
         \ab[3][44] , \ab[3][43] , \ab[3][42] , \ab[3][41] , \ab[3][40] ,
         \ab[3][39] , \ab[3][38] , \ab[3][37] , \ab[3][36] , \ab[3][35] ,
         \ab[3][34] , \ab[3][33] , \ab[3][32] , \ab[3][31] , \ab[3][30] ,
         \ab[3][29] , \ab[3][28] , \ab[3][27] , \ab[3][26] , \ab[3][25] ,
         \ab[3][24] , \ab[3][23] , \ab[3][22] , \ab[3][21] , \ab[3][20] ,
         \ab[3][19] , \ab[3][18] , \ab[3][17] , \ab[3][16] , \ab[3][15] ,
         \ab[3][14] , \ab[3][13] , \ab[3][12] , \ab[3][11] , \ab[3][10] ,
         \ab[3][9] , \ab[3][8] , \ab[3][7] , \ab[3][6] , \ab[3][5] ,
         \ab[3][4] , \ab[3][3] , \ab[3][2] , \ab[3][1] , \ab[3][0] ,
         \ab[2][52] , \ab[2][51] , \ab[2][50] , \ab[2][49] , \ab[2][48] ,
         \ab[2][47] , \ab[2][46] , \ab[2][45] , \ab[2][44] , \ab[2][43] ,
         \ab[2][42] , \ab[2][41] , \ab[2][40] , \ab[2][39] , \ab[2][38] ,
         \ab[2][37] , \ab[2][36] , \ab[2][35] , \ab[2][34] , \ab[2][33] ,
         \ab[2][32] , \ab[2][31] , \ab[2][30] , \ab[2][29] , \ab[2][28] ,
         \ab[2][27] , \ab[2][26] , \ab[2][25] , \ab[2][24] , \ab[2][23] ,
         \ab[2][22] , \ab[2][21] , \ab[2][20] , \ab[2][19] , \ab[2][18] ,
         \ab[2][17] , \ab[2][16] , \ab[2][15] , \ab[2][14] , \ab[2][13] ,
         \ab[2][12] , \ab[2][11] , \ab[2][10] , \ab[2][9] , \ab[2][8] ,
         \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] ,
         \ab[2][2] , \ab[2][1] , \ab[2][0] , \ab[1][52] , \ab[1][51] ,
         \ab[1][50] , \ab[1][49] , \ab[1][48] , \ab[1][47] , \ab[1][46] ,
         \ab[1][45] , \ab[1][44] , \ab[1][43] , \ab[1][42] , \ab[1][41] ,
         \ab[1][40] , \ab[1][39] , \ab[1][38] , \ab[1][37] , \ab[1][36] ,
         \ab[1][35] , \ab[1][34] , \ab[1][33] , \ab[1][32] , \ab[1][31] ,
         \ab[1][30] , \ab[1][29] , \ab[1][28] , \ab[1][27] , \ab[1][26] ,
         \ab[1][25] , \ab[1][24] , \ab[1][23] , \ab[1][22] , \ab[1][21] ,
         \ab[1][20] , \ab[1][19] , \ab[1][18] , \ab[1][17] , \ab[1][16] ,
         \ab[1][15] , \ab[1][14] , \ab[1][13] , \ab[1][12] , \ab[1][11] ,
         \ab[1][10] , \ab[1][9] , \ab[1][8] , \ab[1][7] , \ab[1][6] ,
         \ab[1][5] , \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] ,
         \ab[1][0] , \ab[0][52] , \ab[0][51] , \ab[0][50] , \ab[0][49] ,
         \ab[0][48] , \ab[0][47] , \ab[0][46] , \ab[0][45] , \ab[0][44] ,
         \ab[0][43] , \ab[0][42] , \ab[0][41] , \ab[0][40] , \ab[0][39] ,
         \ab[0][38] , \ab[0][37] , \ab[0][36] , \ab[0][35] , \ab[0][34] ,
         \ab[0][33] , \ab[0][32] , \ab[0][31] , \ab[0][30] , \ab[0][29] ,
         \ab[0][28] , \ab[0][27] , \ab[0][26] , \ab[0][25] , \ab[0][24] ,
         \ab[0][23] , \ab[0][22] , \ab[0][21] , \ab[0][20] , \ab[0][19] ,
         \ab[0][18] , \ab[0][17] , \ab[0][16] , \ab[0][15] , \ab[0][14] ,
         \ab[0][13] , \ab[0][12] , \ab[0][11] , \ab[0][10] , \ab[0][9] ,
         \ab[0][8] , \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] ,
         \ab[0][3] , \ab[0][2] , \ab[0][1] , \CARRYB[4][36] , \CARRYB[4][35] ,
         \CARRYB[4][34] , \CARRYB[4][33] , \CARRYB[4][32] , \CARRYB[4][31] ,
         \CARRYB[4][30] , \CARRYB[4][29] , \CARRYB[4][28] , \CARRYB[4][27] ,
         \CARRYB[4][26] , \CARRYB[4][25] , \CARRYB[4][24] , \CARRYB[4][23] ,
         \CARRYB[4][22] , \CARRYB[4][21] , \CARRYB[4][20] , \CARRYB[4][19] ,
         \CARRYB[4][18] , \CARRYB[4][17] , \CARRYB[4][16] , \CARRYB[4][15] ,
         \CARRYB[4][14] , \CARRYB[4][13] , \CARRYB[4][12] , \CARRYB[4][11] ,
         \CARRYB[4][10] , \CARRYB[4][9] , \CARRYB[4][8] , \CARRYB[4][7] ,
         \CARRYB[4][6] , \CARRYB[4][5] , \CARRYB[4][4] , \CARRYB[4][3] ,
         \CARRYB[4][2] , \CARRYB[4][1] , \CARRYB[4][0] , \CARRYB[3][51] ,
         \CARRYB[3][50] , \CARRYB[3][49] , \CARRYB[3][48] , \CARRYB[3][47] ,
         \CARRYB[3][46] , \CARRYB[3][45] , \CARRYB[3][44] , \CARRYB[3][43] ,
         \CARRYB[3][42] , \CARRYB[3][41] , \CARRYB[3][40] , \CARRYB[3][39] ,
         \CARRYB[3][38] , \CARRYB[3][37] , \CARRYB[3][36] , \CARRYB[3][35] ,
         \CARRYB[3][34] , \CARRYB[3][33] , \CARRYB[3][32] , \CARRYB[3][31] ,
         \CARRYB[3][30] , \CARRYB[3][29] , \CARRYB[3][28] , \CARRYB[3][27] ,
         \CARRYB[3][26] , \CARRYB[3][25] , \CARRYB[3][24] , \CARRYB[3][23] ,
         \CARRYB[3][22] , \CARRYB[3][21] , \CARRYB[3][20] , \CARRYB[3][19] ,
         \CARRYB[3][18] , \CARRYB[3][17] , \CARRYB[3][16] , \CARRYB[3][15] ,
         \CARRYB[3][14] , \CARRYB[3][13] , \CARRYB[3][12] , \CARRYB[3][11] ,
         \CARRYB[3][10] , \CARRYB[3][9] , \CARRYB[3][8] , \CARRYB[3][7] ,
         \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][4] , \CARRYB[3][3] ,
         \CARRYB[3][2] , \CARRYB[3][1] , \CARRYB[3][0] , \CARRYB[2][51] ,
         \CARRYB[2][50] , \CARRYB[2][49] , \CARRYB[2][48] , \CARRYB[2][47] ,
         \CARRYB[2][46] , \CARRYB[2][45] , \CARRYB[2][44] , \CARRYB[2][43] ,
         \CARRYB[2][42] , \CARRYB[2][41] , \CARRYB[2][40] , \CARRYB[2][39] ,
         \CARRYB[2][38] , \CARRYB[2][37] , \CARRYB[2][36] , \CARRYB[2][35] ,
         \CARRYB[2][34] , \CARRYB[2][33] , \CARRYB[2][32] , \CARRYB[2][31] ,
         \CARRYB[2][30] , \CARRYB[2][29] , \CARRYB[2][28] , \CARRYB[2][27] ,
         \CARRYB[2][26] , \CARRYB[2][25] , \CARRYB[2][24] , \CARRYB[2][23] ,
         \CARRYB[2][22] , \CARRYB[2][21] , \CARRYB[2][20] , \CARRYB[2][19] ,
         \CARRYB[2][18] , \CARRYB[2][17] , \CARRYB[2][16] , \CARRYB[2][15] ,
         \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] , \CARRYB[2][11] ,
         \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][7] ,
         \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] ,
         \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] , \SUMB[4][36] ,
         \SUMB[4][35] , \SUMB[4][34] , \SUMB[4][33] , \SUMB[4][32] ,
         \SUMB[4][31] , \SUMB[4][30] , \SUMB[4][29] , \SUMB[4][28] ,
         \SUMB[4][27] , \SUMB[4][26] , \SUMB[4][25] , \SUMB[4][24] ,
         \SUMB[4][23] , \SUMB[4][22] , \SUMB[4][21] , \SUMB[4][20] ,
         \SUMB[4][19] , \SUMB[4][18] , \SUMB[4][17] , \SUMB[4][16] ,
         \SUMB[4][15] , \SUMB[4][14] , \SUMB[4][13] , \SUMB[4][12] ,
         \SUMB[4][11] , \SUMB[4][10] , \SUMB[4][9] , \SUMB[4][8] ,
         \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] ,
         \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][51] , \SUMB[3][50] ,
         \SUMB[3][49] , \SUMB[3][48] , \SUMB[3][47] , \SUMB[3][46] ,
         \SUMB[3][45] , \SUMB[3][44] , \SUMB[3][43] , \SUMB[3][42] ,
         \SUMB[3][41] , \SUMB[3][40] , \SUMB[3][39] , \SUMB[3][38] ,
         \SUMB[3][37] , \SUMB[3][36] , \SUMB[3][35] , \SUMB[3][34] ,
         \SUMB[3][33] , \SUMB[3][32] , \SUMB[3][31] , \SUMB[3][30] ,
         \SUMB[3][29] , \SUMB[3][28] , \SUMB[3][27] , \SUMB[3][26] ,
         \SUMB[3][25] , \SUMB[3][24] , \SUMB[3][23] , \SUMB[3][22] ,
         \SUMB[3][21] , \SUMB[3][20] , \SUMB[3][19] , \SUMB[3][18] ,
         \SUMB[3][17] , \SUMB[3][16] , \SUMB[3][15] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][51] ,
         \SUMB[2][50] , \SUMB[2][49] , \SUMB[2][48] , \SUMB[2][47] ,
         \SUMB[2][46] , \SUMB[2][45] , \SUMB[2][44] , \SUMB[2][43] ,
         \SUMB[2][42] , \SUMB[2][41] , \SUMB[2][40] , \SUMB[2][39] ,
         \SUMB[2][38] , \SUMB[2][37] , \SUMB[2][36] , \SUMB[2][35] ,
         \SUMB[2][34] , \SUMB[2][33] , \SUMB[2][32] , \SUMB[2][31] ,
         \SUMB[2][30] , \SUMB[2][29] , \SUMB[2][28] , \SUMB[2][27] ,
         \SUMB[2][26] , \SUMB[2][25] , \SUMB[2][24] , \SUMB[2][23] ,
         \SUMB[2][22] , \SUMB[2][21] , \SUMB[2][20] , \SUMB[2][19] ,
         \SUMB[2][18] , \SUMB[2][17] , \SUMB[2][16] , \SUMB[2][15] ,
         \SUMB[2][14] , \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] ,
         \SUMB[2][10] , \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] ,
         \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] ,
         \CARRYB[14][18] , \CARRYB[14][17] , \CARRYB[14][16] ,
         \CARRYB[14][15] , \CARRYB[14][14] , \CARRYB[14][13] ,
         \CARRYB[14][12] , \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] ,
         \CARRYB[14][8] , \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] ,
         \CARRYB[14][4] , \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] ,
         \CARRYB[14][0] , \CARRYB[13][51] , \CARRYB[13][50] , \CARRYB[13][49] ,
         \CARRYB[13][48] , \CARRYB[13][47] , \CARRYB[13][46] ,
         \CARRYB[13][45] , \CARRYB[13][44] , \CARRYB[13][43] ,
         \CARRYB[13][42] , \CARRYB[13][41] , \CARRYB[13][40] ,
         \CARRYB[13][39] , \CARRYB[13][38] , \CARRYB[13][37] ,
         \CARRYB[13][36] , \CARRYB[13][35] , \CARRYB[13][34] ,
         \CARRYB[13][33] , \CARRYB[13][32] , \CARRYB[13][31] ,
         \CARRYB[13][30] , \CARRYB[13][29] , \CARRYB[13][28] ,
         \CARRYB[13][27] , \CARRYB[13][26] , \CARRYB[13][25] ,
         \CARRYB[13][24] , \CARRYB[13][23] , \CARRYB[13][22] ,
         \CARRYB[13][21] , \CARRYB[13][20] , \CARRYB[13][19] ,
         \CARRYB[13][18] , \CARRYB[13][17] , \CARRYB[13][16] ,
         \CARRYB[13][15] , \CARRYB[13][14] , \CARRYB[13][13] ,
         \CARRYB[13][12] , \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] ,
         \CARRYB[13][8] , \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] ,
         \CARRYB[13][4] , \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] ,
         \CARRYB[13][0] , \CARRYB[12][51] , \CARRYB[12][50] , \CARRYB[12][49] ,
         \CARRYB[12][48] , \CARRYB[12][47] , \CARRYB[12][46] ,
         \CARRYB[12][45] , \CARRYB[12][44] , \CARRYB[12][43] ,
         \CARRYB[12][42] , \CARRYB[12][41] , \CARRYB[12][40] ,
         \CARRYB[12][39] , \CARRYB[12][38] , \CARRYB[12][37] ,
         \CARRYB[12][36] , \CARRYB[12][35] , \CARRYB[12][34] ,
         \CARRYB[12][33] , \CARRYB[12][32] , \CARRYB[12][31] ,
         \CARRYB[12][30] , \CARRYB[12][29] , \CARRYB[12][28] ,
         \CARRYB[12][27] , \CARRYB[12][26] , \CARRYB[12][25] ,
         \CARRYB[12][24] , \CARRYB[12][23] , \CARRYB[12][22] ,
         \CARRYB[12][21] , \CARRYB[12][20] , \CARRYB[12][19] ,
         \CARRYB[12][18] , \CARRYB[12][17] , \CARRYB[12][16] ,
         \CARRYB[12][15] , \CARRYB[12][14] , \CARRYB[12][13] ,
         \CARRYB[12][12] , \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] ,
         \CARRYB[12][8] , \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] ,
         \CARRYB[12][4] , \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] ,
         \CARRYB[12][0] , \CARRYB[11][51] , \CARRYB[11][50] , \CARRYB[11][49] ,
         \CARRYB[11][48] , \CARRYB[11][47] , \CARRYB[11][46] ,
         \CARRYB[11][45] , \CARRYB[11][44] , \CARRYB[11][43] ,
         \CARRYB[11][42] , \CARRYB[11][41] , \CARRYB[11][40] ,
         \CARRYB[11][39] , \CARRYB[11][38] , \CARRYB[11][37] ,
         \CARRYB[11][36] , \CARRYB[11][35] , \CARRYB[11][34] ,
         \CARRYB[11][33] , \CARRYB[11][32] , \CARRYB[11][31] ,
         \CARRYB[11][30] , \CARRYB[11][29] , \CARRYB[11][28] ,
         \CARRYB[11][27] , \CARRYB[11][26] , \CARRYB[11][25] ,
         \CARRYB[11][24] , \CARRYB[11][23] , \CARRYB[11][22] ,
         \CARRYB[11][21] , \CARRYB[11][20] , \CARRYB[11][19] ,
         \CARRYB[11][18] , \CARRYB[11][17] , \CARRYB[11][16] ,
         \CARRYB[11][15] , \CARRYB[11][14] , \CARRYB[11][13] ,
         \CARRYB[11][12] , \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] ,
         \CARRYB[11][8] , \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] ,
         \CARRYB[11][4] , \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] ,
         \CARRYB[11][0] , \CARRYB[10][51] , \CARRYB[10][50] , \CARRYB[10][49] ,
         \CARRYB[10][48] , \CARRYB[10][47] , \CARRYB[10][46] ,
         \CARRYB[10][45] , \CARRYB[10][44] , \CARRYB[10][43] ,
         \CARRYB[10][42] , \CARRYB[10][41] , \CARRYB[10][40] ,
         \CARRYB[10][39] , \CARRYB[10][38] , \CARRYB[10][37] ,
         \CARRYB[10][36] , \CARRYB[10][35] , \CARRYB[10][34] ,
         \CARRYB[10][33] , \CARRYB[10][32] , \CARRYB[10][31] ,
         \CARRYB[10][30] , \CARRYB[10][29] , \CARRYB[10][28] ,
         \CARRYB[10][27] , \CARRYB[10][26] , \CARRYB[10][25] ,
         \CARRYB[10][24] , \CARRYB[10][23] , \CARRYB[10][22] ,
         \CARRYB[10][21] , \CARRYB[10][20] , \CARRYB[10][19] ,
         \CARRYB[10][18] , \CARRYB[10][17] , \CARRYB[10][16] ,
         \CARRYB[10][15] , \CARRYB[10][14] , \CARRYB[10][13] ,
         \CARRYB[10][12] , \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] ,
         \CARRYB[10][8] , \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] ,
         \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] ,
         \CARRYB[10][0] , \CARRYB[9][51] , \CARRYB[9][50] , \CARRYB[9][49] ,
         \CARRYB[9][48] , \CARRYB[9][47] , \CARRYB[9][46] , \CARRYB[9][45] ,
         \CARRYB[9][44] , \CARRYB[9][43] , \CARRYB[9][42] , \CARRYB[9][41] ,
         \CARRYB[9][40] , \CARRYB[9][39] , \CARRYB[9][38] , \CARRYB[9][37] ,
         \CARRYB[9][36] , \CARRYB[9][35] , \CARRYB[9][34] , \CARRYB[9][33] ,
         \CARRYB[9][32] , \CARRYB[9][31] , \CARRYB[9][30] , \CARRYB[9][29] ,
         \CARRYB[9][28] , \CARRYB[9][27] , \CARRYB[9][26] , \CARRYB[9][25] ,
         \CARRYB[9][24] , \CARRYB[9][23] , \CARRYB[9][22] , \CARRYB[9][21] ,
         \CARRYB[9][20] , \CARRYB[9][19] , \CARRYB[9][18] , \CARRYB[9][17] ,
         \CARRYB[9][16] , \CARRYB[9][15] , \CARRYB[9][14] , \CARRYB[9][13] ,
         \CARRYB[9][12] , \CARRYB[9][11] , \CARRYB[9][10] , \CARRYB[9][9] ,
         \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] , \CARRYB[9][5] ,
         \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] , \CARRYB[9][1] ,
         \CARRYB[9][0] , \CARRYB[8][51] , \CARRYB[8][50] , \CARRYB[8][49] ,
         \CARRYB[8][48] , \CARRYB[8][47] , \CARRYB[8][46] , \CARRYB[8][45] ,
         \CARRYB[8][44] , \CARRYB[8][43] , \CARRYB[8][42] , \CARRYB[8][41] ,
         \CARRYB[8][40] , \CARRYB[8][39] , \CARRYB[8][38] , \CARRYB[8][37] ,
         \CARRYB[8][36] , \CARRYB[8][35] , \CARRYB[8][34] , \CARRYB[8][33] ,
         \CARRYB[8][32] , \CARRYB[8][31] , \CARRYB[8][30] , \CARRYB[8][29] ,
         \CARRYB[8][28] , \CARRYB[8][27] , \CARRYB[8][26] , \CARRYB[8][25] ,
         \CARRYB[8][24] , \CARRYB[8][23] , \CARRYB[8][22] , \CARRYB[8][21] ,
         \CARRYB[8][20] , \CARRYB[8][19] , \CARRYB[8][18] , \CARRYB[8][17] ,
         \CARRYB[8][16] , \CARRYB[8][15] , \CARRYB[8][14] , \CARRYB[8][13] ,
         \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] , \CARRYB[8][9] ,
         \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] ,
         \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] ,
         \CARRYB[8][0] , \CARRYB[7][51] , \CARRYB[7][50] , \CARRYB[7][49] ,
         \CARRYB[7][48] , \CARRYB[7][47] , \CARRYB[7][46] , \CARRYB[7][45] ,
         \CARRYB[7][44] , \CARRYB[7][43] , \CARRYB[7][42] , \CARRYB[7][41] ,
         \CARRYB[7][40] , \CARRYB[7][39] , \CARRYB[7][38] , \CARRYB[7][37] ,
         \CARRYB[7][36] , \CARRYB[7][35] , \CARRYB[7][34] , \CARRYB[7][33] ,
         \CARRYB[7][32] , \CARRYB[7][31] , \CARRYB[7][30] , \CARRYB[7][29] ,
         \CARRYB[7][28] , \CARRYB[7][27] , \CARRYB[7][26] , \CARRYB[7][25] ,
         \CARRYB[7][24] , \CARRYB[7][23] , \CARRYB[7][22] , \CARRYB[7][21] ,
         \CARRYB[7][20] , \CARRYB[7][19] , \CARRYB[7][18] , \CARRYB[7][17] ,
         \CARRYB[7][16] , \CARRYB[7][15] , \CARRYB[7][14] , \CARRYB[7][13] ,
         \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] ,
         \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] ,
         \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] ,
         \CARRYB[7][0] , \CARRYB[6][51] , \CARRYB[6][50] , \CARRYB[6][49] ,
         \CARRYB[6][48] , \CARRYB[6][47] , \CARRYB[6][46] , \CARRYB[6][45] ,
         \CARRYB[6][44] , \CARRYB[6][43] , \CARRYB[6][42] , \CARRYB[6][41] ,
         \CARRYB[6][40] , \CARRYB[6][39] , \CARRYB[6][38] , \CARRYB[6][37] ,
         \CARRYB[6][36] , \CARRYB[6][35] , \CARRYB[6][34] , \CARRYB[6][33] ,
         \CARRYB[6][32] , \CARRYB[6][31] , \CARRYB[6][30] , \CARRYB[6][29] ,
         \CARRYB[6][28] , \CARRYB[6][27] , \CARRYB[6][26] , \CARRYB[6][25] ,
         \CARRYB[6][24] , \CARRYB[6][23] , \CARRYB[6][22] , \CARRYB[6][21] ,
         \CARRYB[6][20] , \CARRYB[6][19] , \CARRYB[6][18] , \CARRYB[6][17] ,
         \CARRYB[6][16] , \CARRYB[6][15] , \CARRYB[6][14] , \CARRYB[6][13] ,
         \CARRYB[6][12] , \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] ,
         \CARRYB[6][8] , \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] ,
         \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] ,
         \CARRYB[6][0] , \CARRYB[5][51] , \CARRYB[5][50] , \CARRYB[5][49] ,
         \CARRYB[5][48] , \CARRYB[5][47] , \CARRYB[5][46] , \CARRYB[5][45] ,
         \CARRYB[5][44] , \CARRYB[5][43] , \CARRYB[5][42] , \CARRYB[5][41] ,
         \CARRYB[5][40] , \CARRYB[5][39] , \CARRYB[5][38] , \CARRYB[5][37] ,
         \CARRYB[5][36] , \CARRYB[5][35] , \CARRYB[5][34] , \CARRYB[5][33] ,
         \CARRYB[5][32] , \CARRYB[5][31] , \CARRYB[5][30] , \CARRYB[5][29] ,
         \CARRYB[5][28] , \CARRYB[5][27] , \CARRYB[5][26] , \CARRYB[5][25] ,
         \CARRYB[5][24] , \CARRYB[5][23] , \CARRYB[5][22] , \CARRYB[5][21] ,
         \CARRYB[5][20] , \CARRYB[5][19] , \CARRYB[5][18] , \CARRYB[5][17] ,
         \CARRYB[5][16] , \CARRYB[5][15] , \CARRYB[5][14] , \CARRYB[5][13] ,
         \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] , \CARRYB[5][9] ,
         \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] , \CARRYB[5][5] ,
         \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] , \CARRYB[5][1] ,
         \CARRYB[5][0] , \CARRYB[4][51] , \CARRYB[4][50] , \CARRYB[4][49] ,
         \CARRYB[4][48] , \CARRYB[4][47] , \CARRYB[4][46] , \CARRYB[4][45] ,
         \CARRYB[4][44] , \CARRYB[4][43] , \CARRYB[4][42] , \CARRYB[4][41] ,
         \CARRYB[4][40] , \CARRYB[4][39] , \CARRYB[4][38] , \CARRYB[4][37] ,
         \SUMB[14][18] , \SUMB[14][17] , \SUMB[14][16] , \SUMB[14][15] ,
         \SUMB[14][14] , \SUMB[14][13] , \SUMB[14][12] , \SUMB[14][11] ,
         \SUMB[14][10] , \SUMB[14][9] , \SUMB[14][8] , \SUMB[14][7] ,
         \SUMB[14][6] , \SUMB[14][5] , \SUMB[14][4] , \SUMB[14][3] ,
         \SUMB[14][2] , \SUMB[14][1] , \SUMB[13][51] , \SUMB[13][50] ,
         \SUMB[13][49] , \SUMB[13][48] , \SUMB[13][47] , \SUMB[13][46] ,
         \SUMB[13][45] , \SUMB[13][44] , \SUMB[13][43] , \SUMB[13][42] ,
         \SUMB[13][41] , \SUMB[13][40] , \SUMB[13][39] , \SUMB[13][38] ,
         \SUMB[13][37] , \SUMB[13][36] , \SUMB[13][35] , \SUMB[13][34] ,
         \SUMB[13][33] , \SUMB[13][32] , \SUMB[13][31] , \SUMB[13][30] ,
         \SUMB[13][29] , \SUMB[13][28] , \SUMB[13][27] , \SUMB[13][26] ,
         \SUMB[13][25] , \SUMB[13][24] , \SUMB[13][23] , \SUMB[13][22] ,
         \SUMB[13][21] , \SUMB[13][20] , \SUMB[13][19] , \SUMB[13][18] ,
         \SUMB[13][17] , \SUMB[13][16] , \SUMB[13][15] , \SUMB[13][14] ,
         \SUMB[13][13] , \SUMB[13][12] , \SUMB[13][11] , \SUMB[13][10] ,
         \SUMB[13][9] , \SUMB[13][8] , \SUMB[13][7] , \SUMB[13][6] ,
         \SUMB[13][5] , \SUMB[13][4] , \SUMB[13][3] , \SUMB[13][2] ,
         \SUMB[13][1] , \SUMB[12][51] , \SUMB[12][50] , \SUMB[12][49] ,
         \SUMB[12][48] , \SUMB[12][47] , \SUMB[12][46] , \SUMB[12][45] ,
         \SUMB[12][44] , \SUMB[12][43] , \SUMB[12][42] , \SUMB[12][41] ,
         \SUMB[12][40] , \SUMB[12][39] , \SUMB[12][38] , \SUMB[12][37] ,
         \SUMB[12][36] , \SUMB[12][35] , \SUMB[12][34] , \SUMB[12][33] ,
         \SUMB[12][32] , \SUMB[12][31] , \SUMB[12][30] , \SUMB[12][29] ,
         \SUMB[12][28] , \SUMB[12][27] , \SUMB[12][26] , \SUMB[12][25] ,
         \SUMB[12][24] , \SUMB[12][23] , \SUMB[12][22] , \SUMB[12][21] ,
         \SUMB[12][20] , \SUMB[12][19] , \SUMB[12][18] , \SUMB[12][17] ,
         \SUMB[12][16] , \SUMB[12][15] , \SUMB[12][14] , \SUMB[12][13] ,
         \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][10] , \SUMB[12][9] ,
         \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] , \SUMB[12][5] ,
         \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] , \SUMB[12][1] ,
         \SUMB[11][51] , \SUMB[11][50] , \SUMB[11][49] , \SUMB[11][48] ,
         \SUMB[11][47] , \SUMB[11][46] , \SUMB[11][45] , \SUMB[11][44] ,
         \SUMB[11][43] , \SUMB[11][42] , \SUMB[11][41] , \SUMB[11][40] ,
         \SUMB[11][39] , \SUMB[11][38] , \SUMB[11][37] , \SUMB[11][36] ,
         \SUMB[11][35] , \SUMB[11][34] , \SUMB[11][33] , \SUMB[11][32] ,
         \SUMB[11][31] , \SUMB[11][30] , \SUMB[11][29] , \SUMB[11][28] ,
         \SUMB[11][27] , \SUMB[11][26] , \SUMB[11][25] , \SUMB[11][24] ,
         \SUMB[11][23] , \SUMB[11][22] , \SUMB[11][21] , \SUMB[11][20] ,
         \SUMB[11][19] , \SUMB[11][18] , \SUMB[11][17] , \SUMB[11][16] ,
         \SUMB[11][15] , \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] ,
         \SUMB[11][11] , \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] ,
         \SUMB[11][7] , \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] ,
         \SUMB[11][3] , \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][51] ,
         \SUMB[10][50] , \SUMB[10][49] , \SUMB[10][48] , \SUMB[10][47] ,
         \SUMB[10][46] , \SUMB[10][45] , \SUMB[10][44] , \SUMB[10][43] ,
         \SUMB[10][42] , \SUMB[10][41] , \SUMB[10][40] , \SUMB[10][39] ,
         \SUMB[10][38] , \SUMB[10][37] , \SUMB[10][36] , \SUMB[10][35] ,
         \SUMB[10][34] , \SUMB[10][33] , \SUMB[10][32] , \SUMB[10][31] ,
         \SUMB[10][30] , \SUMB[10][29] , \SUMB[10][28] , \SUMB[10][27] ,
         \SUMB[10][26] , \SUMB[10][25] , \SUMB[10][24] , \SUMB[10][23] ,
         \SUMB[10][22] , \SUMB[10][21] , \SUMB[10][20] , \SUMB[10][19] ,
         \SUMB[10][18] , \SUMB[10][17] , \SUMB[10][16] , \SUMB[10][15] ,
         \SUMB[10][14] , \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] ,
         \SUMB[10][10] , \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] ,
         \SUMB[10][6] , \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] ,
         \SUMB[10][2] , \SUMB[10][1] , \SUMB[9][51] , \SUMB[9][50] ,
         \SUMB[9][49] , \SUMB[9][48] , \SUMB[9][47] , \SUMB[9][46] ,
         \SUMB[9][45] , \SUMB[9][44] , \SUMB[9][43] , \SUMB[9][42] ,
         \SUMB[9][41] , \SUMB[9][40] , \SUMB[9][39] , \SUMB[9][38] ,
         \SUMB[9][37] , \SUMB[9][36] , \SUMB[9][35] , \SUMB[9][34] ,
         \SUMB[9][33] , \SUMB[9][32] , \SUMB[9][31] , \SUMB[9][30] ,
         \SUMB[9][29] , \SUMB[9][28] , \SUMB[9][27] , \SUMB[9][26] ,
         \SUMB[9][25] , \SUMB[9][24] , \SUMB[9][23] , \SUMB[9][22] ,
         \SUMB[9][21] , \SUMB[9][20] , \SUMB[9][19] , \SUMB[9][18] ,
         \SUMB[9][17] , \SUMB[9][16] , \SUMB[9][15] , \SUMB[9][14] ,
         \SUMB[9][13] , \SUMB[9][12] , \SUMB[9][11] , \SUMB[9][10] ,
         \SUMB[9][9] , \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] ,
         \SUMB[9][4] , \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][51] ,
         \SUMB[8][50] , \SUMB[8][49] , \SUMB[8][48] , \SUMB[8][47] ,
         \SUMB[8][46] , \SUMB[8][45] , \SUMB[8][44] , \SUMB[8][43] ,
         \SUMB[8][42] , \SUMB[8][41] , \SUMB[8][40] , \SUMB[8][39] ,
         \SUMB[8][38] , \SUMB[8][37] , \SUMB[8][36] , \SUMB[8][35] ,
         \SUMB[8][34] , \SUMB[8][33] , \SUMB[8][32] , \SUMB[8][31] ,
         \SUMB[8][30] , \SUMB[8][29] , \SUMB[8][28] , \SUMB[8][27] ,
         \SUMB[8][26] , \SUMB[8][25] , \SUMB[8][24] , \SUMB[8][23] ,
         \SUMB[8][22] , \SUMB[8][21] , \SUMB[8][20] , \SUMB[8][19] ,
         \SUMB[8][18] , \SUMB[8][17] , \SUMB[8][16] , \SUMB[8][15] ,
         \SUMB[8][14] , \SUMB[8][13] , \SUMB[8][12] , \SUMB[8][11] ,
         \SUMB[8][10] , \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] ,
         \SUMB[8][5] , \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] ,
         \SUMB[7][51] , \SUMB[7][50] , \SUMB[7][49] , \SUMB[7][48] ,
         \SUMB[7][47] , \SUMB[7][46] , \SUMB[7][45] , \SUMB[7][44] ,
         \SUMB[7][43] , \SUMB[7][42] , \SUMB[7][41] , \SUMB[7][40] ,
         \SUMB[7][39] , \SUMB[7][38] , \SUMB[7][37] , \SUMB[7][36] ,
         \SUMB[7][35] , \SUMB[7][34] , \SUMB[7][33] , \SUMB[7][32] ,
         \SUMB[7][31] , \SUMB[7][30] , \SUMB[7][29] , \SUMB[7][28] ,
         \SUMB[7][27] , \SUMB[7][26] , \SUMB[7][25] , \SUMB[7][24] ,
         \SUMB[7][23] , \SUMB[7][22] , \SUMB[7][21] , \SUMB[7][20] ,
         \SUMB[7][19] , \SUMB[7][18] , \SUMB[7][17] , \SUMB[7][16] ,
         \SUMB[7][15] , \SUMB[7][14] , \SUMB[7][13] , \SUMB[7][12] ,
         \SUMB[7][11] , \SUMB[7][10] , \SUMB[7][9] , \SUMB[7][8] ,
         \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] ,
         \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][51] , \SUMB[6][50] ,
         \SUMB[6][49] , \SUMB[6][48] , \SUMB[6][47] , \SUMB[6][46] ,
         \SUMB[6][45] , \SUMB[6][44] , \SUMB[6][43] , \SUMB[6][42] ,
         \SUMB[6][41] , \SUMB[6][40] , \SUMB[6][39] , \SUMB[6][38] ,
         \SUMB[6][37] , \SUMB[6][36] , \SUMB[6][35] , \SUMB[6][34] ,
         \SUMB[6][33] , \SUMB[6][32] , \SUMB[6][31] , \SUMB[6][30] ,
         \SUMB[6][29] , \SUMB[6][28] , \SUMB[6][27] , \SUMB[6][26] ,
         \SUMB[6][25] , \SUMB[6][24] , \SUMB[6][23] , \SUMB[6][22] ,
         \SUMB[6][21] , \SUMB[6][20] , \SUMB[6][19] , \SUMB[6][18] ,
         \SUMB[6][17] , \SUMB[6][16] , \SUMB[6][15] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][51] ,
         \SUMB[5][50] , \SUMB[5][49] , \SUMB[5][48] , \SUMB[5][47] ,
         \SUMB[5][46] , \SUMB[5][45] , \SUMB[5][44] , \SUMB[5][43] ,
         \SUMB[5][42] , \SUMB[5][41] , \SUMB[5][40] , \SUMB[5][39] ,
         \SUMB[5][38] , \SUMB[5][37] , \SUMB[5][36] , \SUMB[5][35] ,
         \SUMB[5][34] , \SUMB[5][33] , \SUMB[5][32] , \SUMB[5][31] ,
         \SUMB[5][30] , \SUMB[5][29] , \SUMB[5][28] , \SUMB[5][27] ,
         \SUMB[5][26] , \SUMB[5][25] , \SUMB[5][24] , \SUMB[5][23] ,
         \SUMB[5][22] , \SUMB[5][21] , \SUMB[5][20] , \SUMB[5][19] ,
         \SUMB[5][18] , \SUMB[5][17] , \SUMB[5][16] , \SUMB[5][15] ,
         \SUMB[5][14] , \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] ,
         \SUMB[5][10] , \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][51] , \SUMB[4][50] , \SUMB[4][49] , \SUMB[4][48] ,
         \SUMB[4][47] , \SUMB[4][46] , \SUMB[4][45] , \SUMB[4][44] ,
         \SUMB[4][43] , \SUMB[4][42] , \SUMB[4][41] , \SUMB[4][40] ,
         \SUMB[4][39] , \SUMB[4][38] , \SUMB[4][37] , \CARRYB[24][0] ,
         \CARRYB[23][51] , \CARRYB[23][50] , \CARRYB[23][49] ,
         \CARRYB[23][48] , \CARRYB[23][47] , \CARRYB[23][46] ,
         \CARRYB[23][45] , \CARRYB[23][44] , \CARRYB[23][43] ,
         \CARRYB[23][42] , \CARRYB[23][41] , \CARRYB[23][40] ,
         \CARRYB[23][39] , \CARRYB[23][38] , \CARRYB[23][37] ,
         \CARRYB[23][36] , \CARRYB[23][35] , \CARRYB[23][34] ,
         \CARRYB[23][33] , \CARRYB[23][32] , \CARRYB[23][31] ,
         \CARRYB[23][30] , \CARRYB[23][29] , \CARRYB[23][28] ,
         \CARRYB[23][27] , \CARRYB[23][26] , \CARRYB[23][25] ,
         \CARRYB[23][24] , \CARRYB[23][23] , \CARRYB[23][22] ,
         \CARRYB[23][21] , \CARRYB[23][20] , \CARRYB[23][19] ,
         \CARRYB[23][18] , \CARRYB[23][17] , \CARRYB[23][16] ,
         \CARRYB[23][15] , \CARRYB[23][14] , \CARRYB[23][13] ,
         \CARRYB[23][12] , \CARRYB[23][11] , \CARRYB[23][10] , \CARRYB[23][9] ,
         \CARRYB[23][8] , \CARRYB[23][7] , \CARRYB[23][6] , \CARRYB[23][5] ,
         \CARRYB[23][4] , \CARRYB[23][3] , \CARRYB[23][2] , \CARRYB[23][1] ,
         \CARRYB[23][0] , \CARRYB[22][51] , \CARRYB[22][50] , \CARRYB[22][49] ,
         \CARRYB[22][48] , \CARRYB[22][47] , \CARRYB[22][46] ,
         \CARRYB[22][45] , \CARRYB[22][44] , \CARRYB[22][43] ,
         \CARRYB[22][42] , \CARRYB[22][41] , \CARRYB[22][40] ,
         \CARRYB[22][39] , \CARRYB[22][38] , \CARRYB[22][37] ,
         \CARRYB[22][36] , \CARRYB[22][35] , \CARRYB[22][34] ,
         \CARRYB[22][33] , \CARRYB[22][32] , \CARRYB[22][31] ,
         \CARRYB[22][30] , \CARRYB[22][29] , \CARRYB[22][28] ,
         \CARRYB[22][27] , \CARRYB[22][26] , \CARRYB[22][25] ,
         \CARRYB[22][24] , \CARRYB[22][23] , \CARRYB[22][22] ,
         \CARRYB[22][21] , \CARRYB[22][20] , \CARRYB[22][19] ,
         \CARRYB[22][18] , \CARRYB[22][17] , \CARRYB[22][16] ,
         \CARRYB[22][15] , \CARRYB[22][14] , \CARRYB[22][13] ,
         \CARRYB[22][12] , \CARRYB[22][11] , \CARRYB[22][10] , \CARRYB[22][9] ,
         \CARRYB[22][8] , \CARRYB[22][7] , \CARRYB[22][6] , \CARRYB[22][5] ,
         \CARRYB[22][4] , \CARRYB[22][3] , \CARRYB[22][2] , \CARRYB[22][1] ,
         \CARRYB[22][0] , \CARRYB[21][51] , \CARRYB[21][50] , \CARRYB[21][49] ,
         \CARRYB[21][48] , \CARRYB[21][47] , \CARRYB[21][46] ,
         \CARRYB[21][45] , \CARRYB[21][44] , \CARRYB[21][43] ,
         \CARRYB[21][42] , \CARRYB[21][41] , \CARRYB[21][40] ,
         \CARRYB[21][39] , \CARRYB[21][38] , \CARRYB[21][37] ,
         \CARRYB[21][36] , \CARRYB[21][35] , \CARRYB[21][34] ,
         \CARRYB[21][33] , \CARRYB[21][32] , \CARRYB[21][31] ,
         \CARRYB[21][30] , \CARRYB[21][29] , \CARRYB[21][28] ,
         \CARRYB[21][27] , \CARRYB[21][26] , \CARRYB[21][25] ,
         \CARRYB[21][24] , \CARRYB[21][23] , \CARRYB[21][22] ,
         \CARRYB[21][21] , \CARRYB[21][20] , \CARRYB[21][19] ,
         \CARRYB[21][18] , \CARRYB[21][17] , \CARRYB[21][16] ,
         \CARRYB[21][15] , \CARRYB[21][14] , \CARRYB[21][13] ,
         \CARRYB[21][12] , \CARRYB[21][11] , \CARRYB[21][10] , \CARRYB[21][9] ,
         \CARRYB[21][8] , \CARRYB[21][7] , \CARRYB[21][6] , \CARRYB[21][5] ,
         \CARRYB[21][4] , \CARRYB[21][3] , \CARRYB[21][2] , \CARRYB[21][1] ,
         \CARRYB[21][0] , \CARRYB[20][51] , \CARRYB[20][50] , \CARRYB[20][49] ,
         \CARRYB[20][48] , \CARRYB[20][47] , \CARRYB[20][46] ,
         \CARRYB[20][45] , \CARRYB[20][44] , \CARRYB[20][43] ,
         \CARRYB[20][42] , \CARRYB[20][41] , \CARRYB[20][40] ,
         \CARRYB[20][39] , \CARRYB[20][38] , \CARRYB[20][37] ,
         \CARRYB[20][36] , \CARRYB[20][35] , \CARRYB[20][34] ,
         \CARRYB[20][33] , \CARRYB[20][32] , \CARRYB[20][31] ,
         \CARRYB[20][30] , \CARRYB[20][29] , \CARRYB[20][28] ,
         \CARRYB[20][27] , \CARRYB[20][26] , \CARRYB[20][25] ,
         \CARRYB[20][24] , \CARRYB[20][23] , \CARRYB[20][22] ,
         \CARRYB[20][21] , \CARRYB[20][20] , \CARRYB[20][19] ,
         \CARRYB[20][18] , \CARRYB[20][17] , \CARRYB[20][16] ,
         \CARRYB[20][15] , \CARRYB[20][14] , \CARRYB[20][13] ,
         \CARRYB[20][12] , \CARRYB[20][11] , \CARRYB[20][10] , \CARRYB[20][9] ,
         \CARRYB[20][8] , \CARRYB[20][7] , \CARRYB[20][6] , \CARRYB[20][5] ,
         \CARRYB[20][4] , \CARRYB[20][3] , \CARRYB[20][2] , \CARRYB[20][1] ,
         \CARRYB[20][0] , \CARRYB[19][51] , \CARRYB[19][50] , \CARRYB[19][49] ,
         \CARRYB[19][48] , \CARRYB[19][47] , \CARRYB[19][46] ,
         \CARRYB[19][45] , \CARRYB[19][44] , \CARRYB[19][43] ,
         \CARRYB[19][42] , \CARRYB[19][41] , \CARRYB[19][40] ,
         \CARRYB[19][39] , \CARRYB[19][38] , \CARRYB[19][37] ,
         \CARRYB[19][36] , \CARRYB[19][35] , \CARRYB[19][34] ,
         \CARRYB[19][33] , \CARRYB[19][32] , \CARRYB[19][31] ,
         \CARRYB[19][30] , \CARRYB[19][29] , \CARRYB[19][28] ,
         \CARRYB[19][27] , \CARRYB[19][26] , \CARRYB[19][25] ,
         \CARRYB[19][24] , \CARRYB[19][23] , \CARRYB[19][22] ,
         \CARRYB[19][21] , \CARRYB[19][20] , \CARRYB[19][19] ,
         \CARRYB[19][18] , \CARRYB[19][17] , \CARRYB[19][16] ,
         \CARRYB[19][15] , \CARRYB[19][14] , \CARRYB[19][13] ,
         \CARRYB[19][12] , \CARRYB[19][11] , \CARRYB[19][10] , \CARRYB[19][9] ,
         \CARRYB[19][8] , \CARRYB[19][7] , \CARRYB[19][6] , \CARRYB[19][5] ,
         \CARRYB[19][4] , \CARRYB[19][3] , \CARRYB[19][2] , \CARRYB[19][1] ,
         \CARRYB[19][0] , \CARRYB[18][51] , \CARRYB[18][50] , \CARRYB[18][49] ,
         \CARRYB[18][48] , \CARRYB[18][47] , \CARRYB[18][46] ,
         \CARRYB[18][45] , \CARRYB[18][44] , \CARRYB[18][43] ,
         \CARRYB[18][42] , \CARRYB[18][41] , \CARRYB[18][40] ,
         \CARRYB[18][39] , \CARRYB[18][38] , \CARRYB[18][37] ,
         \CARRYB[18][36] , \CARRYB[18][35] , \CARRYB[18][34] ,
         \CARRYB[18][33] , \CARRYB[18][32] , \CARRYB[18][31] ,
         \CARRYB[18][30] , \CARRYB[18][29] , \CARRYB[18][28] ,
         \CARRYB[18][27] , \CARRYB[18][26] , \CARRYB[18][25] ,
         \CARRYB[18][24] , \CARRYB[18][23] , \CARRYB[18][22] ,
         \CARRYB[18][21] , \CARRYB[18][20] , \CARRYB[18][19] ,
         \CARRYB[18][18] , \CARRYB[18][17] , \CARRYB[18][16] ,
         \CARRYB[18][15] , \CARRYB[18][14] , \CARRYB[18][13] ,
         \CARRYB[18][12] , \CARRYB[18][11] , \CARRYB[18][10] , \CARRYB[18][9] ,
         \CARRYB[18][8] , \CARRYB[18][7] , \CARRYB[18][6] , \CARRYB[18][5] ,
         \CARRYB[18][4] , \CARRYB[18][3] , \CARRYB[18][2] , \CARRYB[18][1] ,
         \CARRYB[18][0] , \CARRYB[17][51] , \CARRYB[17][50] , \CARRYB[17][49] ,
         \CARRYB[17][48] , \CARRYB[17][47] , \CARRYB[17][46] ,
         \CARRYB[17][45] , \CARRYB[17][44] , \CARRYB[17][43] ,
         \CARRYB[17][42] , \CARRYB[17][41] , \CARRYB[17][40] ,
         \CARRYB[17][39] , \CARRYB[17][38] , \CARRYB[17][37] ,
         \CARRYB[17][36] , \CARRYB[17][35] , \CARRYB[17][34] ,
         \CARRYB[17][33] , \CARRYB[17][32] , \CARRYB[17][31] ,
         \CARRYB[17][30] , \CARRYB[17][29] , \CARRYB[17][28] ,
         \CARRYB[17][27] , \CARRYB[17][26] , \CARRYB[17][25] ,
         \CARRYB[17][24] , \CARRYB[17][23] , \CARRYB[17][22] ,
         \CARRYB[17][21] , \CARRYB[17][20] , \CARRYB[17][19] ,
         \CARRYB[17][18] , \CARRYB[17][17] , \CARRYB[17][16] ,
         \CARRYB[17][15] , \CARRYB[17][14] , \CARRYB[17][13] ,
         \CARRYB[17][12] , \CARRYB[17][11] , \CARRYB[17][10] , \CARRYB[17][9] ,
         \CARRYB[17][8] , \CARRYB[17][7] , \CARRYB[17][6] , \CARRYB[17][5] ,
         \CARRYB[17][4] , \CARRYB[17][3] , \CARRYB[17][2] , \CARRYB[17][1] ,
         \CARRYB[17][0] , \CARRYB[16][51] , \CARRYB[16][50] , \CARRYB[16][49] ,
         \CARRYB[16][48] , \CARRYB[16][47] , \CARRYB[16][46] ,
         \CARRYB[16][45] , \CARRYB[16][44] , \CARRYB[16][43] ,
         \CARRYB[16][42] , \CARRYB[16][41] , \CARRYB[16][40] ,
         \CARRYB[16][39] , \CARRYB[16][38] , \CARRYB[16][37] ,
         \CARRYB[16][36] , \CARRYB[16][35] , \CARRYB[16][34] ,
         \CARRYB[16][33] , \CARRYB[16][32] , \CARRYB[16][31] ,
         \CARRYB[16][30] , \CARRYB[16][29] , \CARRYB[16][28] ,
         \CARRYB[16][27] , \CARRYB[16][26] , \CARRYB[16][25] ,
         \CARRYB[16][24] , \CARRYB[16][23] , \CARRYB[16][22] ,
         \CARRYB[16][21] , \CARRYB[16][20] , \CARRYB[16][19] ,
         \CARRYB[16][18] , \CARRYB[16][17] , \CARRYB[16][16] ,
         \CARRYB[16][15] , \CARRYB[16][14] , \CARRYB[16][13] ,
         \CARRYB[16][12] , \CARRYB[16][11] , \CARRYB[16][10] , \CARRYB[16][9] ,
         \CARRYB[16][8] , \CARRYB[16][7] , \CARRYB[16][6] , \CARRYB[16][5] ,
         \CARRYB[16][4] , \CARRYB[16][3] , \CARRYB[16][2] , \CARRYB[16][1] ,
         \CARRYB[16][0] , \CARRYB[15][51] , \CARRYB[15][50] , \CARRYB[15][49] ,
         \CARRYB[15][48] , \CARRYB[15][47] , \CARRYB[15][46] ,
         \CARRYB[15][45] , \CARRYB[15][44] , \CARRYB[15][43] ,
         \CARRYB[15][42] , \CARRYB[15][41] , \CARRYB[15][40] ,
         \CARRYB[15][39] , \CARRYB[15][38] , \CARRYB[15][37] ,
         \CARRYB[15][36] , \CARRYB[15][35] , \CARRYB[15][34] ,
         \CARRYB[15][33] , \CARRYB[15][32] , \CARRYB[15][31] ,
         \CARRYB[15][30] , \CARRYB[15][29] , \CARRYB[15][28] ,
         \CARRYB[15][27] , \CARRYB[15][26] , \CARRYB[15][25] ,
         \CARRYB[15][24] , \CARRYB[15][23] , \CARRYB[15][22] ,
         \CARRYB[15][21] , \CARRYB[15][20] , \CARRYB[15][19] ,
         \CARRYB[15][18] , \CARRYB[15][17] , \CARRYB[15][16] ,
         \CARRYB[15][15] , \CARRYB[15][14] , \CARRYB[15][13] ,
         \CARRYB[15][12] , \CARRYB[15][11] , \CARRYB[15][10] , \CARRYB[15][9] ,
         \CARRYB[15][8] , \CARRYB[15][7] , \CARRYB[15][6] , \CARRYB[15][5] ,
         \CARRYB[15][4] , \CARRYB[15][3] , \CARRYB[15][2] , \CARRYB[15][1] ,
         \CARRYB[15][0] , \CARRYB[14][51] , \CARRYB[14][50] , \CARRYB[14][49] ,
         \CARRYB[14][48] , \CARRYB[14][47] , \CARRYB[14][46] ,
         \CARRYB[14][45] , \CARRYB[14][44] , \CARRYB[14][43] ,
         \CARRYB[14][42] , \CARRYB[14][41] , \CARRYB[14][40] ,
         \CARRYB[14][39] , \CARRYB[14][38] , \CARRYB[14][37] ,
         \CARRYB[14][36] , \CARRYB[14][35] , \CARRYB[14][34] ,
         \CARRYB[14][33] , \CARRYB[14][32] , \CARRYB[14][31] ,
         \CARRYB[14][30] , \CARRYB[14][29] , \CARRYB[14][28] ,
         \CARRYB[14][27] , \CARRYB[14][26] , \CARRYB[14][25] ,
         \CARRYB[14][24] , \CARRYB[14][23] , \CARRYB[14][22] ,
         \CARRYB[14][21] , \CARRYB[14][20] , \CARRYB[14][19] , \SUMB[23][51] ,
         \SUMB[23][50] , \SUMB[23][49] , \SUMB[23][48] , \SUMB[23][47] ,
         \SUMB[23][46] , \SUMB[23][45] , \SUMB[23][44] , \SUMB[23][43] ,
         \SUMB[23][42] , \SUMB[23][41] , \SUMB[23][40] , \SUMB[23][39] ,
         \SUMB[23][38] , \SUMB[23][37] , \SUMB[23][36] , \SUMB[23][35] ,
         \SUMB[23][34] , \SUMB[23][33] , \SUMB[23][32] , \SUMB[23][31] ,
         \SUMB[23][30] , \SUMB[23][29] , \SUMB[23][28] , \SUMB[23][27] ,
         \SUMB[23][26] , \SUMB[23][25] , \SUMB[23][24] , \SUMB[23][23] ,
         \SUMB[23][22] , \SUMB[23][21] , \SUMB[23][20] , \SUMB[23][19] ,
         \SUMB[23][18] , \SUMB[23][17] , \SUMB[23][16] , \SUMB[23][15] ,
         \SUMB[23][14] , \SUMB[23][13] , \SUMB[23][12] , \SUMB[23][11] ,
         \SUMB[23][10] , \SUMB[23][9] , \SUMB[23][8] , \SUMB[23][7] ,
         \SUMB[23][6] , \SUMB[23][5] , \SUMB[23][4] , \SUMB[23][3] ,
         \SUMB[23][2] , \SUMB[23][1] , \SUMB[22][51] , \SUMB[22][50] ,
         \SUMB[22][49] , \SUMB[22][48] , \SUMB[22][47] , \SUMB[22][46] ,
         \SUMB[22][45] , \SUMB[22][44] , \SUMB[22][43] , \SUMB[22][42] ,
         \SUMB[22][41] , \SUMB[22][40] , \SUMB[22][39] , \SUMB[22][38] ,
         \SUMB[22][37] , \SUMB[22][36] , \SUMB[22][35] , \SUMB[22][34] ,
         \SUMB[22][33] , \SUMB[22][32] , \SUMB[22][31] , \SUMB[22][30] ,
         \SUMB[22][29] , \SUMB[22][28] , \SUMB[22][27] , \SUMB[22][26] ,
         \SUMB[22][25] , \SUMB[22][24] , \SUMB[22][23] , \SUMB[22][22] ,
         \SUMB[22][21] , \SUMB[22][20] , \SUMB[22][19] , \SUMB[22][18] ,
         \SUMB[22][17] , \SUMB[22][16] , \SUMB[22][15] , \SUMB[22][14] ,
         \SUMB[22][13] , \SUMB[22][12] , \SUMB[22][11] , \SUMB[22][10] ,
         \SUMB[22][9] , \SUMB[22][8] , \SUMB[22][7] , \SUMB[22][6] ,
         \SUMB[22][5] , \SUMB[22][4] , \SUMB[22][3] , \SUMB[22][2] ,
         \SUMB[22][1] , \SUMB[21][51] , \SUMB[21][50] , \SUMB[21][49] ,
         \SUMB[21][48] , \SUMB[21][47] , \SUMB[21][46] , \SUMB[21][45] ,
         \SUMB[21][44] , \SUMB[21][43] , \SUMB[21][42] , \SUMB[21][41] ,
         \SUMB[21][40] , \SUMB[21][39] , \SUMB[21][38] , \SUMB[21][37] ,
         \SUMB[21][36] , \SUMB[21][35] , \SUMB[21][34] , \SUMB[21][33] ,
         \SUMB[21][32] , \SUMB[21][31] , \SUMB[21][30] , \SUMB[21][29] ,
         \SUMB[21][28] , \SUMB[21][27] , \SUMB[21][26] , \SUMB[21][25] ,
         \SUMB[21][24] , \SUMB[21][23] , \SUMB[21][22] , \SUMB[21][21] ,
         \SUMB[21][20] , \SUMB[21][19] , \SUMB[21][18] , \SUMB[21][17] ,
         \SUMB[21][16] , \SUMB[21][15] , \SUMB[21][14] , \SUMB[21][13] ,
         \SUMB[21][12] , \SUMB[21][11] , \SUMB[21][10] , \SUMB[21][9] ,
         \SUMB[21][8] , \SUMB[21][7] , \SUMB[21][6] , \SUMB[21][5] ,
         \SUMB[21][4] , \SUMB[21][3] , \SUMB[21][2] , \SUMB[21][1] ,
         \SUMB[20][51] , \SUMB[20][50] , \SUMB[20][49] , \SUMB[20][48] ,
         \SUMB[20][47] , \SUMB[20][46] , \SUMB[20][45] , \SUMB[20][44] ,
         \SUMB[20][43] , \SUMB[20][42] , \SUMB[20][41] , \SUMB[20][40] ,
         \SUMB[20][39] , \SUMB[20][38] , \SUMB[20][37] , \SUMB[20][36] ,
         \SUMB[20][35] , \SUMB[20][34] , \SUMB[20][33] , \SUMB[20][32] ,
         \SUMB[20][31] , \SUMB[20][30] , \SUMB[20][29] , \SUMB[20][28] ,
         \SUMB[20][27] , \SUMB[20][26] , \SUMB[20][25] , \SUMB[20][24] ,
         \SUMB[20][23] , \SUMB[20][22] , \SUMB[20][21] , \SUMB[20][20] ,
         \SUMB[20][19] , \SUMB[20][18] , \SUMB[20][17] , \SUMB[20][16] ,
         \SUMB[20][15] , \SUMB[20][14] , \SUMB[20][13] , \SUMB[20][12] ,
         \SUMB[20][11] , \SUMB[20][10] , \SUMB[20][9] , \SUMB[20][8] ,
         \SUMB[20][7] , \SUMB[20][6] , \SUMB[20][5] , \SUMB[20][4] ,
         \SUMB[20][3] , \SUMB[20][2] , \SUMB[20][1] , \SUMB[19][51] ,
         \SUMB[19][50] , \SUMB[19][49] , \SUMB[19][48] , \SUMB[19][47] ,
         \SUMB[19][46] , \SUMB[19][45] , \SUMB[19][44] , \SUMB[19][43] ,
         \SUMB[19][42] , \SUMB[19][41] , \SUMB[19][40] , \SUMB[19][39] ,
         \SUMB[19][38] , \SUMB[19][37] , \SUMB[19][36] , \SUMB[19][35] ,
         \SUMB[19][34] , \SUMB[19][33] , \SUMB[19][32] , \SUMB[19][31] ,
         \SUMB[19][30] , \SUMB[19][29] , \SUMB[19][28] , \SUMB[19][27] ,
         \SUMB[19][26] , \SUMB[19][25] , \SUMB[19][24] , \SUMB[19][23] ,
         \SUMB[19][22] , \SUMB[19][21] , \SUMB[19][20] , \SUMB[19][19] ,
         \SUMB[19][18] , \SUMB[19][17] , \SUMB[19][16] , \SUMB[19][15] ,
         \SUMB[19][14] , \SUMB[19][13] , \SUMB[19][12] , \SUMB[19][11] ,
         \SUMB[19][10] , \SUMB[19][9] , \SUMB[19][8] , \SUMB[19][7] ,
         \SUMB[19][6] , \SUMB[19][5] , \SUMB[19][4] , \SUMB[19][3] ,
         \SUMB[19][2] , \SUMB[19][1] , \SUMB[18][51] , \SUMB[18][50] ,
         \SUMB[18][49] , \SUMB[18][48] , \SUMB[18][47] , \SUMB[18][46] ,
         \SUMB[18][45] , \SUMB[18][44] , \SUMB[18][43] , \SUMB[18][42] ,
         \SUMB[18][41] , \SUMB[18][40] , \SUMB[18][39] , \SUMB[18][38] ,
         \SUMB[18][37] , \SUMB[18][36] , \SUMB[18][35] , \SUMB[18][34] ,
         \SUMB[18][33] , \SUMB[18][32] , \SUMB[18][31] , \SUMB[18][30] ,
         \SUMB[18][29] , \SUMB[18][28] , \SUMB[18][27] , \SUMB[18][26] ,
         \SUMB[18][25] , \SUMB[18][24] , \SUMB[18][23] , \SUMB[18][22] ,
         \SUMB[18][21] , \SUMB[18][20] , \SUMB[18][19] , \SUMB[18][18] ,
         \SUMB[18][17] , \SUMB[18][16] , \SUMB[18][15] , \SUMB[18][14] ,
         \SUMB[18][13] , \SUMB[18][12] , \SUMB[18][11] , \SUMB[18][10] ,
         \SUMB[18][9] , \SUMB[18][8] , \SUMB[18][7] , \SUMB[18][6] ,
         \SUMB[18][5] , \SUMB[18][4] , \SUMB[18][3] , \SUMB[18][2] ,
         \SUMB[18][1] , \SUMB[17][51] , \SUMB[17][50] , \SUMB[17][49] ,
         \SUMB[17][48] , \SUMB[17][47] , \SUMB[17][46] , \SUMB[17][45] ,
         \SUMB[17][44] , \SUMB[17][43] , \SUMB[17][42] , \SUMB[17][41] ,
         \SUMB[17][40] , \SUMB[17][39] , \SUMB[17][38] , \SUMB[17][37] ,
         \SUMB[17][36] , \SUMB[17][35] , \SUMB[17][34] , \SUMB[17][33] ,
         \SUMB[17][32] , \SUMB[17][31] , \SUMB[17][30] , \SUMB[17][29] ,
         \SUMB[17][28] , \SUMB[17][27] , \SUMB[17][26] , \SUMB[17][25] ,
         \SUMB[17][24] , \SUMB[17][23] , \SUMB[17][22] , \SUMB[17][21] ,
         \SUMB[17][20] , \SUMB[17][19] , \SUMB[17][18] , \SUMB[17][17] ,
         \SUMB[17][16] , \SUMB[17][15] , \SUMB[17][14] , \SUMB[17][13] ,
         \SUMB[17][12] , \SUMB[17][11] , \SUMB[17][10] , \SUMB[17][9] ,
         \SUMB[17][8] , \SUMB[17][7] , \SUMB[17][6] , \SUMB[17][5] ,
         \SUMB[17][4] , \SUMB[17][3] , \SUMB[17][2] , \SUMB[17][1] ,
         \SUMB[16][51] , \SUMB[16][50] , \SUMB[16][49] , \SUMB[16][48] ,
         \SUMB[16][47] , \SUMB[16][46] , \SUMB[16][45] , \SUMB[16][44] ,
         \SUMB[16][43] , \SUMB[16][42] , \SUMB[16][41] , \SUMB[16][40] ,
         \SUMB[16][39] , \SUMB[16][38] , \SUMB[16][37] , \SUMB[16][36] ,
         \SUMB[16][35] , \SUMB[16][34] , \SUMB[16][33] , \SUMB[16][32] ,
         \SUMB[16][31] , \SUMB[16][30] , \SUMB[16][29] , \SUMB[16][28] ,
         \SUMB[16][27] , \SUMB[16][26] , \SUMB[16][25] , \SUMB[16][24] ,
         \SUMB[16][23] , \SUMB[16][22] , \SUMB[16][21] , \SUMB[16][20] ,
         \SUMB[16][19] , \SUMB[16][18] , \SUMB[16][17] , \SUMB[16][16] ,
         \SUMB[16][15] , \SUMB[16][14] , \SUMB[16][13] , \SUMB[16][12] ,
         \SUMB[16][11] , \SUMB[16][10] , \SUMB[16][9] , \SUMB[16][8] ,
         \SUMB[16][7] , \SUMB[16][6] , \SUMB[16][5] , \SUMB[16][4] ,
         \SUMB[16][3] , \SUMB[16][2] , \SUMB[16][1] , \SUMB[15][51] ,
         \SUMB[15][50] , \SUMB[15][49] , \SUMB[15][48] , \SUMB[15][47] ,
         \SUMB[15][46] , \SUMB[15][45] , \SUMB[15][44] , \SUMB[15][43] ,
         \SUMB[15][42] , \SUMB[15][41] , \SUMB[15][40] , \SUMB[15][39] ,
         \SUMB[15][38] , \SUMB[15][37] , \SUMB[15][36] , \SUMB[15][35] ,
         \SUMB[15][34] , \SUMB[15][33] , \SUMB[15][32] , \SUMB[15][31] ,
         \SUMB[15][30] , \SUMB[15][29] , \SUMB[15][28] , \SUMB[15][27] ,
         \SUMB[15][26] , \SUMB[15][25] , \SUMB[15][24] , \SUMB[15][23] ,
         \SUMB[15][22] , \SUMB[15][21] , \SUMB[15][20] , \SUMB[15][19] ,
         \SUMB[15][18] , \SUMB[15][17] , \SUMB[15][16] , \SUMB[15][15] ,
         \SUMB[15][14] , \SUMB[15][13] , \SUMB[15][12] , \SUMB[15][11] ,
         \SUMB[15][10] , \SUMB[15][9] , \SUMB[15][8] , \SUMB[15][7] ,
         \SUMB[15][6] , \SUMB[15][5] , \SUMB[15][4] , \SUMB[15][3] ,
         \SUMB[15][2] , \SUMB[15][1] , \SUMB[14][51] , \SUMB[14][50] ,
         \SUMB[14][49] , \SUMB[14][48] , \SUMB[14][47] , \SUMB[14][46] ,
         \SUMB[14][45] , \SUMB[14][44] , \SUMB[14][43] , \SUMB[14][42] ,
         \SUMB[14][41] , \SUMB[14][40] , \SUMB[14][39] , \SUMB[14][38] ,
         \SUMB[14][37] , \SUMB[14][36] , \SUMB[14][35] , \SUMB[14][34] ,
         \SUMB[14][33] , \SUMB[14][32] , \SUMB[14][31] , \SUMB[14][30] ,
         \SUMB[14][29] , \SUMB[14][28] , \SUMB[14][27] , \SUMB[14][26] ,
         \SUMB[14][25] , \SUMB[14][24] , \SUMB[14][23] , \SUMB[14][22] ,
         \SUMB[14][21] , \SUMB[14][20] , \SUMB[14][19] , \CARRYB[33][35] ,
         \CARRYB[33][34] , \CARRYB[33][33] , \CARRYB[33][32] ,
         \CARRYB[33][31] , \CARRYB[33][30] , \CARRYB[33][29] ,
         \CARRYB[33][28] , \CARRYB[33][27] , \CARRYB[33][26] ,
         \CARRYB[33][25] , \CARRYB[33][24] , \CARRYB[33][23] ,
         \CARRYB[33][22] , \CARRYB[33][21] , \CARRYB[33][20] ,
         \CARRYB[33][19] , \CARRYB[33][18] , \CARRYB[33][17] ,
         \CARRYB[33][16] , \CARRYB[33][15] , \CARRYB[33][14] ,
         \CARRYB[33][13] , \CARRYB[33][12] , \CARRYB[33][11] ,
         \CARRYB[33][10] , \CARRYB[33][9] , \CARRYB[33][8] , \CARRYB[33][7] ,
         \CARRYB[33][6] , \CARRYB[33][5] , \CARRYB[33][4] , \CARRYB[33][3] ,
         \CARRYB[33][2] , \CARRYB[33][1] , \CARRYB[33][0] , \CARRYB[32][51] ,
         \CARRYB[32][50] , \CARRYB[32][49] , \CARRYB[32][48] ,
         \CARRYB[32][47] , \CARRYB[32][46] , \CARRYB[32][45] ,
         \CARRYB[32][44] , \CARRYB[32][43] , \CARRYB[32][42] ,
         \CARRYB[32][41] , \CARRYB[32][40] , \CARRYB[32][39] ,
         \CARRYB[32][38] , \CARRYB[32][37] , \CARRYB[32][36] ,
         \CARRYB[32][35] , \CARRYB[32][34] , \CARRYB[32][33] ,
         \CARRYB[32][32] , \CARRYB[32][31] , \CARRYB[32][30] ,
         \CARRYB[32][29] , \CARRYB[32][28] , \CARRYB[32][27] ,
         \CARRYB[32][26] , \CARRYB[32][25] , \CARRYB[32][24] ,
         \CARRYB[32][23] , \CARRYB[32][22] , \CARRYB[32][21] ,
         \CARRYB[32][20] , \CARRYB[32][19] , \CARRYB[32][18] ,
         \CARRYB[32][17] , \CARRYB[32][16] , \CARRYB[32][15] ,
         \CARRYB[32][14] , \CARRYB[32][13] , \CARRYB[32][12] ,
         \CARRYB[32][11] , \CARRYB[32][10] , \CARRYB[32][9] , \CARRYB[32][8] ,
         \CARRYB[32][7] , \CARRYB[32][6] , \CARRYB[32][5] , \CARRYB[32][4] ,
         \CARRYB[32][3] , \CARRYB[32][2] , \CARRYB[32][1] , \CARRYB[32][0] ,
         \CARRYB[31][51] , \CARRYB[31][50] , \CARRYB[31][49] ,
         \CARRYB[31][48] , \CARRYB[31][47] , \CARRYB[31][46] ,
         \CARRYB[31][45] , \CARRYB[31][44] , \CARRYB[31][43] ,
         \CARRYB[31][42] , \CARRYB[31][41] , \CARRYB[31][40] ,
         \CARRYB[31][39] , \CARRYB[31][38] , \CARRYB[31][37] ,
         \CARRYB[31][36] , \CARRYB[31][35] , \CARRYB[31][34] ,
         \CARRYB[31][33] , \CARRYB[31][32] , \CARRYB[31][31] ,
         \CARRYB[31][30] , \CARRYB[31][29] , \CARRYB[31][28] ,
         \CARRYB[31][27] , \CARRYB[31][26] , \CARRYB[31][25] ,
         \CARRYB[31][24] , \CARRYB[31][23] , \CARRYB[31][22] ,
         \CARRYB[31][21] , \CARRYB[31][20] , \CARRYB[31][19] ,
         \CARRYB[31][18] , \CARRYB[31][17] , \CARRYB[31][16] ,
         \CARRYB[31][15] , \CARRYB[31][14] , \CARRYB[31][13] ,
         \CARRYB[31][12] , \CARRYB[31][11] , \CARRYB[31][10] , \CARRYB[31][9] ,
         \CARRYB[31][8] , \CARRYB[31][7] , \CARRYB[31][6] , \CARRYB[31][5] ,
         \CARRYB[31][4] , \CARRYB[31][3] , \CARRYB[31][2] , \CARRYB[31][1] ,
         \CARRYB[31][0] , \CARRYB[30][51] , \CARRYB[30][50] , \CARRYB[30][49] ,
         \CARRYB[30][48] , \CARRYB[30][47] , \CARRYB[30][46] ,
         \CARRYB[30][45] , \CARRYB[30][44] , \CARRYB[30][43] ,
         \CARRYB[30][42] , \CARRYB[30][41] , \CARRYB[30][40] ,
         \CARRYB[30][39] , \CARRYB[30][38] , \CARRYB[30][37] ,
         \CARRYB[30][36] , \CARRYB[30][35] , \CARRYB[30][34] ,
         \CARRYB[30][33] , \CARRYB[30][32] , \CARRYB[30][31] ,
         \CARRYB[30][30] , \CARRYB[30][29] , \CARRYB[30][28] ,
         \CARRYB[30][27] , \CARRYB[30][26] , \CARRYB[30][25] ,
         \CARRYB[30][24] , \CARRYB[30][23] , \CARRYB[30][22] ,
         \CARRYB[30][21] , \CARRYB[30][20] , \CARRYB[30][19] ,
         \CARRYB[30][18] , \CARRYB[30][17] , \CARRYB[30][16] ,
         \CARRYB[30][15] , \CARRYB[30][14] , \CARRYB[30][13] ,
         \CARRYB[30][12] , \CARRYB[30][11] , \CARRYB[30][10] , \CARRYB[30][9] ,
         \CARRYB[30][8] , \CARRYB[30][7] , \CARRYB[30][6] , \CARRYB[30][5] ,
         \CARRYB[30][4] , \CARRYB[30][3] , \CARRYB[30][2] , \CARRYB[30][1] ,
         \CARRYB[30][0] , \CARRYB[29][51] , \CARRYB[29][50] , \CARRYB[29][49] ,
         \CARRYB[29][48] , \CARRYB[29][47] , \CARRYB[29][46] ,
         \CARRYB[29][45] , \CARRYB[29][44] , \CARRYB[29][43] ,
         \CARRYB[29][42] , \CARRYB[29][41] , \CARRYB[29][40] ,
         \CARRYB[29][39] , \CARRYB[29][38] , \CARRYB[29][37] ,
         \CARRYB[29][36] , \CARRYB[29][35] , \CARRYB[29][34] ,
         \CARRYB[29][33] , \CARRYB[29][32] , \CARRYB[29][31] ,
         \CARRYB[29][30] , \CARRYB[29][29] , \CARRYB[29][28] ,
         \CARRYB[29][27] , \CARRYB[29][26] , \CARRYB[29][25] ,
         \CARRYB[29][24] , \CARRYB[29][23] , \CARRYB[29][22] ,
         \CARRYB[29][21] , \CARRYB[29][20] , \CARRYB[29][19] ,
         \CARRYB[29][18] , \CARRYB[29][17] , \CARRYB[29][16] ,
         \CARRYB[29][15] , \CARRYB[29][14] , \CARRYB[29][13] ,
         \CARRYB[29][12] , \CARRYB[29][11] , \CARRYB[29][10] , \CARRYB[29][9] ,
         \CARRYB[29][8] , \CARRYB[29][7] , \CARRYB[29][6] , \CARRYB[29][5] ,
         \CARRYB[29][4] , \CARRYB[29][3] , \CARRYB[29][2] , \CARRYB[29][1] ,
         \CARRYB[29][0] , \CARRYB[28][51] , \CARRYB[28][50] , \CARRYB[28][49] ,
         \CARRYB[28][48] , \CARRYB[28][47] , \CARRYB[28][46] ,
         \CARRYB[28][45] , \CARRYB[28][44] , \CARRYB[28][43] ,
         \CARRYB[28][42] , \CARRYB[28][41] , \CARRYB[28][40] ,
         \CARRYB[28][39] , \CARRYB[28][38] , \CARRYB[28][37] ,
         \CARRYB[28][36] , \CARRYB[28][35] , \CARRYB[28][34] ,
         \CARRYB[28][33] , \CARRYB[28][32] , \CARRYB[28][31] ,
         \CARRYB[28][30] , \CARRYB[28][29] , \CARRYB[28][28] ,
         \CARRYB[28][27] , \CARRYB[28][26] , \CARRYB[28][25] ,
         \CARRYB[28][24] , \CARRYB[28][23] , \CARRYB[28][22] ,
         \CARRYB[28][21] , \CARRYB[28][20] , \CARRYB[28][19] ,
         \CARRYB[28][18] , \CARRYB[28][17] , \CARRYB[28][16] ,
         \CARRYB[28][15] , \CARRYB[28][14] , \CARRYB[28][13] ,
         \CARRYB[28][12] , \CARRYB[28][11] , \CARRYB[28][10] , \CARRYB[28][9] ,
         \CARRYB[28][8] , \CARRYB[28][7] , \CARRYB[28][6] , \CARRYB[28][5] ,
         \CARRYB[28][4] , \CARRYB[28][3] , \CARRYB[28][2] , \CARRYB[28][1] ,
         \CARRYB[28][0] , \CARRYB[27][51] , \CARRYB[27][50] , \CARRYB[27][49] ,
         \CARRYB[27][48] , \CARRYB[27][47] , \CARRYB[27][46] ,
         \CARRYB[27][45] , \CARRYB[27][44] , \CARRYB[27][43] ,
         \CARRYB[27][42] , \CARRYB[27][41] , \CARRYB[27][40] ,
         \CARRYB[27][39] , \CARRYB[27][38] , \CARRYB[27][37] ,
         \CARRYB[27][36] , \CARRYB[27][35] , \CARRYB[27][34] ,
         \CARRYB[27][33] , \CARRYB[27][32] , \CARRYB[27][31] ,
         \CARRYB[27][30] , \CARRYB[27][29] , \CARRYB[27][28] ,
         \CARRYB[27][27] , \CARRYB[27][26] , \CARRYB[27][25] ,
         \CARRYB[27][24] , \CARRYB[27][23] , \CARRYB[27][22] ,
         \CARRYB[27][21] , \CARRYB[27][20] , \CARRYB[27][19] ,
         \CARRYB[27][18] , \CARRYB[27][17] , \CARRYB[27][16] ,
         \CARRYB[27][15] , \CARRYB[27][14] , \CARRYB[27][13] ,
         \CARRYB[27][12] , \CARRYB[27][11] , \CARRYB[27][10] , \CARRYB[27][9] ,
         \CARRYB[27][8] , \CARRYB[27][7] , \CARRYB[27][6] , \CARRYB[27][5] ,
         \CARRYB[27][4] , \CARRYB[27][3] , \CARRYB[27][2] , \CARRYB[27][1] ,
         \CARRYB[27][0] , \CARRYB[26][51] , \CARRYB[26][50] , \CARRYB[26][49] ,
         \CARRYB[26][48] , \CARRYB[26][47] , \CARRYB[26][46] ,
         \CARRYB[26][45] , \CARRYB[26][44] , \CARRYB[26][43] ,
         \CARRYB[26][42] , \CARRYB[26][41] , \CARRYB[26][40] ,
         \CARRYB[26][39] , \CARRYB[26][38] , \CARRYB[26][37] ,
         \CARRYB[26][36] , \CARRYB[26][35] , \CARRYB[26][34] ,
         \CARRYB[26][33] , \CARRYB[26][32] , \CARRYB[26][31] ,
         \CARRYB[26][30] , \CARRYB[26][29] , \CARRYB[26][28] ,
         \CARRYB[26][27] , \CARRYB[26][26] , \CARRYB[26][25] ,
         \CARRYB[26][24] , \CARRYB[26][23] , \CARRYB[26][22] ,
         \CARRYB[26][21] , \CARRYB[26][20] , \CARRYB[26][19] ,
         \CARRYB[26][18] , \CARRYB[26][17] , \CARRYB[26][16] ,
         \CARRYB[26][15] , \CARRYB[26][14] , \CARRYB[26][13] ,
         \CARRYB[26][12] , \CARRYB[26][11] , \CARRYB[26][10] , \CARRYB[26][9] ,
         \CARRYB[26][8] , \CARRYB[26][7] , \CARRYB[26][6] , \CARRYB[26][5] ,
         \CARRYB[26][4] , \CARRYB[26][3] , \CARRYB[26][2] , \CARRYB[26][1] ,
         \CARRYB[26][0] , \CARRYB[25][51] , \CARRYB[25][50] , \CARRYB[25][49] ,
         \CARRYB[25][48] , \CARRYB[25][47] , \CARRYB[25][46] ,
         \CARRYB[25][45] , \CARRYB[25][44] , \CARRYB[25][43] ,
         \CARRYB[25][42] , \CARRYB[25][41] , \CARRYB[25][40] ,
         \CARRYB[25][39] , \CARRYB[25][38] , \CARRYB[25][37] ,
         \CARRYB[25][36] , \CARRYB[25][35] , \CARRYB[25][34] ,
         \CARRYB[25][33] , \CARRYB[25][32] , \CARRYB[25][31] ,
         \CARRYB[25][30] , \CARRYB[25][29] , \CARRYB[25][28] ,
         \CARRYB[25][27] , \CARRYB[25][26] , \CARRYB[25][25] ,
         \CARRYB[25][24] , \CARRYB[25][23] , \CARRYB[25][22] ,
         \CARRYB[25][21] , \CARRYB[25][20] , \CARRYB[25][19] ,
         \CARRYB[25][18] , \CARRYB[25][17] , \CARRYB[25][16] ,
         \CARRYB[25][15] , \CARRYB[25][14] , \CARRYB[25][13] ,
         \CARRYB[25][12] , \CARRYB[25][11] , \CARRYB[25][10] , \CARRYB[25][9] ,
         \CARRYB[25][8] , \CARRYB[25][7] , \CARRYB[25][6] , \CARRYB[25][5] ,
         \CARRYB[25][4] , \CARRYB[25][3] , \CARRYB[25][2] , \CARRYB[25][1] ,
         \CARRYB[25][0] , \CARRYB[24][51] , \CARRYB[24][50] , \CARRYB[24][49] ,
         \CARRYB[24][48] , \CARRYB[24][47] , \CARRYB[24][46] ,
         \CARRYB[24][45] , \CARRYB[24][44] , \CARRYB[24][43] ,
         \CARRYB[24][42] , \CARRYB[24][41] , \CARRYB[24][40] ,
         \CARRYB[24][39] , \CARRYB[24][38] , \CARRYB[24][37] ,
         \CARRYB[24][36] , \CARRYB[24][35] , \CARRYB[24][34] ,
         \CARRYB[24][33] , \CARRYB[24][32] , \CARRYB[24][31] ,
         \CARRYB[24][30] , \CARRYB[24][29] , \CARRYB[24][28] ,
         \CARRYB[24][27] , \CARRYB[24][26] , \CARRYB[24][25] ,
         \CARRYB[24][24] , \CARRYB[24][23] , \CARRYB[24][22] ,
         \CARRYB[24][21] , \CARRYB[24][20] , \CARRYB[24][19] ,
         \CARRYB[24][18] , \CARRYB[24][17] , \CARRYB[24][16] ,
         \CARRYB[24][15] , \CARRYB[24][14] , \CARRYB[24][13] ,
         \CARRYB[24][12] , \CARRYB[24][11] , \CARRYB[24][10] , \CARRYB[24][9] ,
         \CARRYB[24][8] , \CARRYB[24][7] , \CARRYB[24][6] , \CARRYB[24][5] ,
         \CARRYB[24][4] , \CARRYB[24][3] , \CARRYB[24][2] , \CARRYB[24][1] ,
         \SUMB[33][35] , \SUMB[33][34] , \SUMB[33][33] , \SUMB[33][32] ,
         \SUMB[33][31] , \SUMB[33][30] , \SUMB[33][29] , \SUMB[33][28] ,
         \SUMB[33][27] , \SUMB[33][26] , \SUMB[33][25] , \SUMB[33][24] ,
         \SUMB[33][23] , \SUMB[33][22] , \SUMB[33][21] , \SUMB[33][20] ,
         \SUMB[33][19] , \SUMB[33][18] , \SUMB[33][17] , \SUMB[33][16] ,
         \SUMB[33][15] , \SUMB[33][14] , \SUMB[33][13] , \SUMB[33][12] ,
         \SUMB[33][11] , \SUMB[33][10] , \SUMB[33][9] , \SUMB[33][8] ,
         \SUMB[33][7] , \SUMB[33][6] , \SUMB[33][5] , \SUMB[33][4] ,
         \SUMB[33][3] , \SUMB[33][2] , \SUMB[33][1] , \SUMB[32][51] ,
         \SUMB[32][50] , \SUMB[32][49] , \SUMB[32][48] , \SUMB[32][47] ,
         \SUMB[32][46] , \SUMB[32][45] , \SUMB[32][44] , \SUMB[32][43] ,
         \SUMB[32][42] , \SUMB[32][41] , \SUMB[32][40] , \SUMB[32][39] ,
         \SUMB[32][38] , \SUMB[32][37] , \SUMB[32][36] , \SUMB[32][35] ,
         \SUMB[32][34] , \SUMB[32][33] , \SUMB[32][32] , \SUMB[32][31] ,
         \SUMB[32][30] , \SUMB[32][29] , \SUMB[32][28] , \SUMB[32][27] ,
         \SUMB[32][26] , \SUMB[32][25] , \SUMB[32][24] , \SUMB[32][23] ,
         \SUMB[32][22] , \SUMB[32][21] , \SUMB[32][20] , \SUMB[32][19] ,
         \SUMB[32][18] , \SUMB[32][17] , \SUMB[32][16] , \SUMB[32][15] ,
         \SUMB[32][14] , \SUMB[32][13] , \SUMB[32][12] , \SUMB[32][11] ,
         \SUMB[32][10] , \SUMB[32][9] , \SUMB[32][8] , \SUMB[32][7] ,
         \SUMB[32][6] , \SUMB[32][5] , \SUMB[32][4] , \SUMB[32][3] ,
         \SUMB[32][2] , \SUMB[32][1] , \SUMB[31][51] , \SUMB[31][50] ,
         \SUMB[31][49] , \SUMB[31][48] , \SUMB[31][47] , \SUMB[31][46] ,
         \SUMB[31][45] , \SUMB[31][44] , \SUMB[31][43] , \SUMB[31][42] ,
         \SUMB[31][41] , \SUMB[31][40] , \SUMB[31][39] , \SUMB[31][38] ,
         \SUMB[31][37] , \SUMB[31][36] , \SUMB[31][35] , \SUMB[31][34] ,
         \SUMB[31][33] , \SUMB[31][32] , \SUMB[31][31] , \SUMB[31][30] ,
         \SUMB[31][29] , \SUMB[31][28] , \SUMB[31][27] , \SUMB[31][26] ,
         \SUMB[31][25] , \SUMB[31][24] , \SUMB[31][23] , \SUMB[31][22] ,
         \SUMB[31][21] , \SUMB[31][20] , \SUMB[31][19] , \SUMB[31][18] ,
         \SUMB[31][17] , \SUMB[31][16] , \SUMB[31][15] , \SUMB[31][14] ,
         \SUMB[31][13] , \SUMB[31][12] , \SUMB[31][11] , \SUMB[31][10] ,
         \SUMB[31][9] , \SUMB[31][8] , \SUMB[31][7] , \SUMB[31][6] ,
         \SUMB[31][5] , \SUMB[31][4] , \SUMB[31][3] , \SUMB[31][2] ,
         \SUMB[31][1] , \SUMB[30][51] , \SUMB[30][50] , \SUMB[30][49] ,
         \SUMB[30][48] , \SUMB[30][47] , \SUMB[30][46] , \SUMB[30][45] ,
         \SUMB[30][44] , \SUMB[30][43] , \SUMB[30][42] , \SUMB[30][41] ,
         \SUMB[30][40] , \SUMB[30][39] , \SUMB[30][38] , \SUMB[30][37] ,
         \SUMB[30][36] , \SUMB[30][35] , \SUMB[30][34] , \SUMB[30][33] ,
         \SUMB[30][32] , \SUMB[30][31] , \SUMB[30][30] , \SUMB[30][29] ,
         \SUMB[30][28] , \SUMB[30][27] , \SUMB[30][26] , \SUMB[30][25] ,
         \SUMB[30][24] , \SUMB[30][23] , \SUMB[30][22] , \SUMB[30][21] ,
         \SUMB[30][20] , \SUMB[30][19] , \SUMB[30][18] , \SUMB[30][17] ,
         \SUMB[30][16] , \SUMB[30][15] , \SUMB[30][14] , \SUMB[30][13] ,
         \SUMB[30][12] , \SUMB[30][11] , \SUMB[30][10] , \SUMB[30][9] ,
         \SUMB[30][8] , \SUMB[30][7] , \SUMB[30][6] , \SUMB[30][5] ,
         \SUMB[30][4] , \SUMB[30][3] , \SUMB[30][2] , \SUMB[30][1] ,
         \SUMB[29][51] , \SUMB[29][50] , \SUMB[29][49] , \SUMB[29][48] ,
         \SUMB[29][47] , \SUMB[29][46] , \SUMB[29][45] , \SUMB[29][44] ,
         \SUMB[29][43] , \SUMB[29][42] , \SUMB[29][41] , \SUMB[29][40] ,
         \SUMB[29][39] , \SUMB[29][38] , \SUMB[29][37] , \SUMB[29][36] ,
         \SUMB[29][35] , \SUMB[29][34] , \SUMB[29][33] , \SUMB[29][32] ,
         \SUMB[29][31] , \SUMB[29][30] , \SUMB[29][29] , \SUMB[29][28] ,
         \SUMB[29][27] , \SUMB[29][26] , \SUMB[29][25] , \SUMB[29][24] ,
         \SUMB[29][23] , \SUMB[29][22] , \SUMB[29][21] , \SUMB[29][20] ,
         \SUMB[29][19] , \SUMB[29][18] , \SUMB[29][17] , \SUMB[29][16] ,
         \SUMB[29][15] , \SUMB[29][14] , \SUMB[29][13] , \SUMB[29][12] ,
         \SUMB[29][11] , \SUMB[29][10] , \SUMB[29][9] , \SUMB[29][8] ,
         \SUMB[29][7] , \SUMB[29][6] , \SUMB[29][5] , \SUMB[29][4] ,
         \SUMB[29][3] , \SUMB[29][2] , \SUMB[29][1] , \SUMB[28][51] ,
         \SUMB[28][50] , \SUMB[28][49] , \SUMB[28][48] , \SUMB[28][47] ,
         \SUMB[28][46] , \SUMB[28][45] , \SUMB[28][44] , \SUMB[28][43] ,
         \SUMB[28][42] , \SUMB[28][41] , \SUMB[28][40] , \SUMB[28][39] ,
         \SUMB[28][38] , \SUMB[28][37] , \SUMB[28][36] , \SUMB[28][35] ,
         \SUMB[28][34] , \SUMB[28][33] , \SUMB[28][32] , \SUMB[28][31] ,
         \SUMB[28][30] , \SUMB[28][29] , \SUMB[28][28] , \SUMB[28][27] ,
         \SUMB[28][26] , \SUMB[28][25] , \SUMB[28][24] , \SUMB[28][23] ,
         \SUMB[28][22] , \SUMB[28][21] , \SUMB[28][20] , \SUMB[28][19] ,
         \SUMB[28][18] , \SUMB[28][17] , \SUMB[28][16] , \SUMB[28][15] ,
         \SUMB[28][14] , \SUMB[28][13] , \SUMB[28][12] , \SUMB[28][11] ,
         \SUMB[28][10] , \SUMB[28][9] , \SUMB[28][8] , \SUMB[28][7] ,
         \SUMB[28][6] , \SUMB[28][5] , \SUMB[28][4] , \SUMB[28][3] ,
         \SUMB[28][2] , \SUMB[28][1] , \SUMB[27][51] , \SUMB[27][50] ,
         \SUMB[27][49] , \SUMB[27][48] , \SUMB[27][47] , \SUMB[27][46] ,
         \SUMB[27][45] , \SUMB[27][44] , \SUMB[27][43] , \SUMB[27][42] ,
         \SUMB[27][41] , \SUMB[27][40] , \SUMB[27][39] , \SUMB[27][38] ,
         \SUMB[27][37] , \SUMB[27][36] , \SUMB[27][35] , \SUMB[27][34] ,
         \SUMB[27][33] , \SUMB[27][32] , \SUMB[27][31] , \SUMB[27][30] ,
         \SUMB[27][29] , \SUMB[27][28] , \SUMB[27][27] , \SUMB[27][26] ,
         \SUMB[27][25] , \SUMB[27][24] , \SUMB[27][23] , \SUMB[27][22] ,
         \SUMB[27][21] , \SUMB[27][20] , \SUMB[27][19] , \SUMB[27][18] ,
         \SUMB[27][17] , \SUMB[27][16] , \SUMB[27][15] , \SUMB[27][14] ,
         \SUMB[27][13] , \SUMB[27][12] , \SUMB[27][11] , \SUMB[27][10] ,
         \SUMB[27][9] , \SUMB[27][8] , \SUMB[27][7] , \SUMB[27][6] ,
         \SUMB[27][5] , \SUMB[27][4] , \SUMB[27][3] , \SUMB[27][2] ,
         \SUMB[27][1] , \SUMB[26][51] , \SUMB[26][50] , \SUMB[26][49] ,
         \SUMB[26][48] , \SUMB[26][47] , \SUMB[26][46] , \SUMB[26][45] ,
         \SUMB[26][44] , \SUMB[26][43] , \SUMB[26][42] , \SUMB[26][41] ,
         \SUMB[26][40] , \SUMB[26][39] , \SUMB[26][38] , \SUMB[26][37] ,
         \SUMB[26][36] , \SUMB[26][35] , \SUMB[26][34] , \SUMB[26][33] ,
         \SUMB[26][32] , \SUMB[26][31] , \SUMB[26][30] , \SUMB[26][29] ,
         \SUMB[26][28] , \SUMB[26][27] , \SUMB[26][26] , \SUMB[26][25] ,
         \SUMB[26][24] , \SUMB[26][23] , \SUMB[26][22] , \SUMB[26][21] ,
         \SUMB[26][20] , \SUMB[26][19] , \SUMB[26][18] , \SUMB[26][17] ,
         \SUMB[26][16] , \SUMB[26][15] , \SUMB[26][14] , \SUMB[26][13] ,
         \SUMB[26][12] , \SUMB[26][11] , \SUMB[26][10] , \SUMB[26][9] ,
         \SUMB[26][8] , \SUMB[26][7] , \SUMB[26][6] , \SUMB[26][5] ,
         \SUMB[26][4] , \SUMB[26][3] , \SUMB[26][2] , \SUMB[26][1] ,
         \SUMB[25][51] , \SUMB[25][50] , \SUMB[25][49] , \SUMB[25][48] ,
         \SUMB[25][47] , \SUMB[25][46] , \SUMB[25][45] , \SUMB[25][44] ,
         \SUMB[25][43] , \SUMB[25][42] , \SUMB[25][41] , \SUMB[25][40] ,
         \SUMB[25][39] , \SUMB[25][38] , \SUMB[25][37] , \SUMB[25][36] ,
         \SUMB[25][35] , \SUMB[25][34] , \SUMB[25][33] , \SUMB[25][32] ,
         \SUMB[25][31] , \SUMB[25][30] , \SUMB[25][29] , \SUMB[25][28] ,
         \SUMB[25][27] , \SUMB[25][26] , \SUMB[25][25] , \SUMB[25][24] ,
         \SUMB[25][23] , \SUMB[25][22] , \SUMB[25][21] , \SUMB[25][20] ,
         \SUMB[25][19] , \SUMB[25][18] , \SUMB[25][17] , \SUMB[25][16] ,
         \SUMB[25][15] , \SUMB[25][14] , \SUMB[25][13] , \SUMB[25][12] ,
         \SUMB[25][11] , \SUMB[25][10] , \SUMB[25][9] , \SUMB[25][8] ,
         \SUMB[25][7] , \SUMB[25][6] , \SUMB[25][5] , \SUMB[25][4] ,
         \SUMB[25][3] , \SUMB[25][2] , \SUMB[25][1] , \SUMB[24][51] ,
         \SUMB[24][50] , \SUMB[24][49] , \SUMB[24][48] , \SUMB[24][47] ,
         \SUMB[24][46] , \SUMB[24][45] , \SUMB[24][44] , \SUMB[24][43] ,
         \SUMB[24][42] , \SUMB[24][41] , \SUMB[24][40] , \SUMB[24][39] ,
         \SUMB[24][38] , \SUMB[24][37] , \SUMB[24][36] , \SUMB[24][35] ,
         \SUMB[24][34] , \SUMB[24][33] , \SUMB[24][32] , \SUMB[24][31] ,
         \SUMB[24][30] , \SUMB[24][29] , \SUMB[24][28] , \SUMB[24][27] ,
         \SUMB[24][26] , \SUMB[24][25] , \SUMB[24][24] , \SUMB[24][23] ,
         \SUMB[24][22] , \SUMB[24][21] , \SUMB[24][20] , \SUMB[24][19] ,
         \SUMB[24][18] , \SUMB[24][17] , \SUMB[24][16] , \SUMB[24][15] ,
         \SUMB[24][14] , \SUMB[24][13] , \SUMB[24][12] , \SUMB[24][11] ,
         \SUMB[24][10] , \SUMB[24][9] , \SUMB[24][8] , \SUMB[24][7] ,
         \SUMB[24][6] , \SUMB[24][5] , \SUMB[24][4] , \SUMB[24][3] ,
         \SUMB[24][2] , \SUMB[24][1] , \CARRYB[43][17] , \CARRYB[43][16] ,
         \CARRYB[43][15] , \CARRYB[43][14] , \CARRYB[43][13] ,
         \CARRYB[43][12] , \CARRYB[43][11] , \CARRYB[43][10] , \CARRYB[43][9] ,
         \CARRYB[43][8] , \CARRYB[43][7] , \CARRYB[43][6] , \CARRYB[43][5] ,
         \CARRYB[43][4] , \CARRYB[43][3] , \CARRYB[43][2] , \CARRYB[43][1] ,
         \CARRYB[43][0] , \CARRYB[42][51] , \CARRYB[42][50] , \CARRYB[42][49] ,
         \CARRYB[42][48] , \CARRYB[42][47] , \CARRYB[42][46] ,
         \CARRYB[42][45] , \CARRYB[42][44] , \CARRYB[42][43] ,
         \CARRYB[42][42] , \CARRYB[42][41] , \CARRYB[42][40] ,
         \CARRYB[42][39] , \CARRYB[42][38] , \CARRYB[42][37] ,
         \CARRYB[42][36] , \CARRYB[42][35] , \CARRYB[42][34] ,
         \CARRYB[42][33] , \CARRYB[42][32] , \CARRYB[42][31] ,
         \CARRYB[42][30] , \CARRYB[42][29] , \CARRYB[42][28] ,
         \CARRYB[42][27] , \CARRYB[42][26] , \CARRYB[42][25] ,
         \CARRYB[42][24] , \CARRYB[42][23] , \CARRYB[42][22] ,
         \CARRYB[42][21] , \CARRYB[42][20] , \CARRYB[42][19] ,
         \CARRYB[42][18] , \CARRYB[42][17] , \CARRYB[42][16] ,
         \CARRYB[42][15] , \CARRYB[42][14] , \CARRYB[42][13] ,
         \CARRYB[42][12] , \CARRYB[42][11] , \CARRYB[42][10] , \CARRYB[42][9] ,
         \CARRYB[42][8] , \CARRYB[42][7] , \CARRYB[42][6] , \CARRYB[42][5] ,
         \CARRYB[42][4] , \CARRYB[42][3] , \CARRYB[42][2] , \CARRYB[42][1] ,
         \CARRYB[42][0] , \CARRYB[41][51] , \CARRYB[41][50] , \CARRYB[41][49] ,
         \CARRYB[41][48] , \CARRYB[41][47] , \CARRYB[41][46] ,
         \CARRYB[41][45] , \CARRYB[41][44] , \CARRYB[41][43] ,
         \CARRYB[41][42] , \CARRYB[41][41] , \CARRYB[41][40] ,
         \CARRYB[41][39] , \CARRYB[41][38] , \CARRYB[41][37] ,
         \CARRYB[41][36] , \CARRYB[41][35] , \CARRYB[41][34] ,
         \CARRYB[41][33] , \CARRYB[41][32] , \CARRYB[41][31] ,
         \CARRYB[41][30] , \CARRYB[41][29] , \CARRYB[41][28] ,
         \CARRYB[41][27] , \CARRYB[41][26] , \CARRYB[41][25] ,
         \CARRYB[41][24] , \CARRYB[41][23] , \CARRYB[41][22] ,
         \CARRYB[41][21] , \CARRYB[41][20] , \CARRYB[41][19] ,
         \CARRYB[41][18] , \CARRYB[41][17] , \CARRYB[41][16] ,
         \CARRYB[41][15] , \CARRYB[41][14] , \CARRYB[41][13] ,
         \CARRYB[41][12] , \CARRYB[41][11] , \CARRYB[41][10] , \CARRYB[41][9] ,
         \CARRYB[41][8] , \CARRYB[41][7] , \CARRYB[41][6] , \CARRYB[41][5] ,
         \CARRYB[41][4] , \CARRYB[41][3] , \CARRYB[41][2] , \CARRYB[41][1] ,
         \CARRYB[41][0] , \CARRYB[40][51] , \CARRYB[40][50] , \CARRYB[40][49] ,
         \CARRYB[40][48] , \CARRYB[40][47] , \CARRYB[40][46] ,
         \CARRYB[40][45] , \CARRYB[40][44] , \CARRYB[40][43] ,
         \CARRYB[40][42] , \CARRYB[40][41] , \CARRYB[40][40] ,
         \CARRYB[40][39] , \CARRYB[40][38] , \CARRYB[40][37] ,
         \CARRYB[40][36] , \CARRYB[40][35] , \CARRYB[40][34] ,
         \CARRYB[40][33] , \CARRYB[40][32] , \CARRYB[40][31] ,
         \CARRYB[40][30] , \CARRYB[40][29] , \CARRYB[40][28] ,
         \CARRYB[40][27] , \CARRYB[40][26] , \CARRYB[40][25] ,
         \CARRYB[40][24] , \CARRYB[40][23] , \CARRYB[40][22] ,
         \CARRYB[40][21] , \CARRYB[40][20] , \CARRYB[40][19] ,
         \CARRYB[40][18] , \CARRYB[40][17] , \CARRYB[40][16] ,
         \CARRYB[40][15] , \CARRYB[40][14] , \CARRYB[40][13] ,
         \CARRYB[40][12] , \CARRYB[40][11] , \CARRYB[40][10] , \CARRYB[40][9] ,
         \CARRYB[40][8] , \CARRYB[40][7] , \CARRYB[40][6] , \CARRYB[40][5] ,
         \CARRYB[40][4] , \CARRYB[40][3] , \CARRYB[40][2] , \CARRYB[40][1] ,
         \CARRYB[40][0] , \CARRYB[39][51] , \CARRYB[39][50] , \CARRYB[39][49] ,
         \CARRYB[39][48] , \CARRYB[39][47] , \CARRYB[39][46] ,
         \CARRYB[39][45] , \CARRYB[39][44] , \CARRYB[39][43] ,
         \CARRYB[39][42] , \CARRYB[39][41] , \CARRYB[39][40] ,
         \CARRYB[39][39] , \CARRYB[39][38] , \CARRYB[39][37] ,
         \CARRYB[39][36] , \CARRYB[39][35] , \CARRYB[39][34] ,
         \CARRYB[39][33] , \CARRYB[39][32] , \CARRYB[39][31] ,
         \CARRYB[39][30] , \CARRYB[39][29] , \CARRYB[39][28] ,
         \CARRYB[39][27] , \CARRYB[39][26] , \CARRYB[39][25] ,
         \CARRYB[39][24] , \CARRYB[39][23] , \CARRYB[39][22] ,
         \CARRYB[39][21] , \CARRYB[39][20] , \CARRYB[39][19] ,
         \CARRYB[39][18] , \CARRYB[39][17] , \CARRYB[39][16] ,
         \CARRYB[39][15] , \CARRYB[39][14] , \CARRYB[39][13] ,
         \CARRYB[39][12] , \CARRYB[39][11] , \CARRYB[39][10] , \CARRYB[39][9] ,
         \CARRYB[39][8] , \CARRYB[39][7] , \CARRYB[39][6] , \CARRYB[39][5] ,
         \CARRYB[39][4] , \CARRYB[39][3] , \CARRYB[39][2] , \CARRYB[39][1] ,
         \CARRYB[39][0] , \CARRYB[38][51] , \CARRYB[38][50] , \CARRYB[38][49] ,
         \CARRYB[38][48] , \CARRYB[38][47] , \CARRYB[38][46] ,
         \CARRYB[38][45] , \CARRYB[38][44] , \CARRYB[38][43] ,
         \CARRYB[38][42] , \CARRYB[38][41] , \CARRYB[38][40] ,
         \CARRYB[38][39] , \CARRYB[38][38] , \CARRYB[38][37] ,
         \CARRYB[38][36] , \CARRYB[38][35] , \CARRYB[38][34] ,
         \CARRYB[38][33] , \CARRYB[38][32] , \CARRYB[38][31] ,
         \CARRYB[38][30] , \CARRYB[38][29] , \CARRYB[38][28] ,
         \CARRYB[38][27] , \CARRYB[38][26] , \CARRYB[38][25] ,
         \CARRYB[38][24] , \CARRYB[38][23] , \CARRYB[38][22] ,
         \CARRYB[38][21] , \CARRYB[38][20] , \CARRYB[38][19] ,
         \CARRYB[38][18] , \CARRYB[38][17] , \CARRYB[38][16] ,
         \CARRYB[38][15] , \CARRYB[38][14] , \CARRYB[38][13] ,
         \CARRYB[38][12] , \CARRYB[38][11] , \CARRYB[38][10] , \CARRYB[38][9] ,
         \CARRYB[38][8] , \CARRYB[38][7] , \CARRYB[38][6] , \CARRYB[38][5] ,
         \CARRYB[38][4] , \CARRYB[38][3] , \CARRYB[38][2] , \CARRYB[38][1] ,
         \CARRYB[38][0] , \CARRYB[37][51] , \CARRYB[37][50] , \CARRYB[37][49] ,
         \CARRYB[37][48] , \CARRYB[37][47] , \CARRYB[37][46] ,
         \CARRYB[37][45] , \CARRYB[37][44] , \CARRYB[37][43] ,
         \CARRYB[37][42] , \CARRYB[37][41] , \CARRYB[37][40] ,
         \CARRYB[37][39] , \CARRYB[37][38] , \CARRYB[37][37] ,
         \CARRYB[37][36] , \CARRYB[37][35] , \CARRYB[37][34] ,
         \CARRYB[37][33] , \CARRYB[37][32] , \CARRYB[37][31] ,
         \CARRYB[37][30] , \CARRYB[37][29] , \CARRYB[37][28] ,
         \CARRYB[37][27] , \CARRYB[37][26] , \CARRYB[37][25] ,
         \CARRYB[37][24] , \CARRYB[37][23] , \CARRYB[37][22] ,
         \CARRYB[37][21] , \CARRYB[37][20] , \CARRYB[37][19] ,
         \CARRYB[37][18] , \CARRYB[37][17] , \CARRYB[37][16] ,
         \CARRYB[37][15] , \CARRYB[37][14] , \CARRYB[37][13] ,
         \CARRYB[37][12] , \CARRYB[37][11] , \CARRYB[37][10] , \CARRYB[37][9] ,
         \CARRYB[37][8] , \CARRYB[37][7] , \CARRYB[37][6] , \CARRYB[37][5] ,
         \CARRYB[37][4] , \CARRYB[37][3] , \CARRYB[37][2] , \CARRYB[37][1] ,
         \CARRYB[37][0] , \CARRYB[36][51] , \CARRYB[36][50] , \CARRYB[36][49] ,
         \CARRYB[36][48] , \CARRYB[36][47] , \CARRYB[36][46] ,
         \CARRYB[36][45] , \CARRYB[36][44] , \CARRYB[36][43] ,
         \CARRYB[36][42] , \CARRYB[36][41] , \CARRYB[36][40] ,
         \CARRYB[36][39] , \CARRYB[36][38] , \CARRYB[36][37] ,
         \CARRYB[36][36] , \CARRYB[36][35] , \CARRYB[36][34] ,
         \CARRYB[36][33] , \CARRYB[36][32] , \CARRYB[36][31] ,
         \CARRYB[36][30] , \CARRYB[36][29] , \CARRYB[36][28] ,
         \CARRYB[36][27] , \CARRYB[36][26] , \CARRYB[36][25] ,
         \CARRYB[36][24] , \CARRYB[36][23] , \CARRYB[36][22] ,
         \CARRYB[36][21] , \CARRYB[36][20] , \CARRYB[36][19] ,
         \CARRYB[36][18] , \CARRYB[36][17] , \CARRYB[36][16] ,
         \CARRYB[36][15] , \CARRYB[36][14] , \CARRYB[36][13] ,
         \CARRYB[36][12] , \CARRYB[36][11] , \CARRYB[36][10] , \CARRYB[36][9] ,
         \CARRYB[36][8] , \CARRYB[36][7] , \CARRYB[36][6] , \CARRYB[36][5] ,
         \CARRYB[36][4] , \CARRYB[36][3] , \CARRYB[36][2] , \CARRYB[36][1] ,
         \CARRYB[36][0] , \CARRYB[35][51] , \CARRYB[35][50] , \CARRYB[35][49] ,
         \CARRYB[35][48] , \CARRYB[35][47] , \CARRYB[35][46] ,
         \CARRYB[35][45] , \CARRYB[35][44] , \CARRYB[35][43] ,
         \CARRYB[35][42] , \CARRYB[35][41] , \CARRYB[35][40] ,
         \CARRYB[35][39] , \CARRYB[35][38] , \CARRYB[35][37] ,
         \CARRYB[35][36] , \CARRYB[35][35] , \CARRYB[35][34] ,
         \CARRYB[35][33] , \CARRYB[35][32] , \CARRYB[35][31] ,
         \CARRYB[35][30] , \CARRYB[35][29] , \CARRYB[35][28] ,
         \CARRYB[35][27] , \CARRYB[35][26] , \CARRYB[35][25] ,
         \CARRYB[35][24] , \CARRYB[35][23] , \CARRYB[35][22] ,
         \CARRYB[35][21] , \CARRYB[35][20] , \CARRYB[35][19] ,
         \CARRYB[35][18] , \CARRYB[35][17] , \CARRYB[35][16] ,
         \CARRYB[35][15] , \CARRYB[35][14] , \CARRYB[35][13] ,
         \CARRYB[35][12] , \CARRYB[35][11] , \CARRYB[35][10] , \CARRYB[35][9] ,
         \CARRYB[35][8] , \CARRYB[35][7] , \CARRYB[35][6] , \CARRYB[35][5] ,
         \CARRYB[35][4] , \CARRYB[35][3] , \CARRYB[35][2] , \CARRYB[35][1] ,
         \CARRYB[35][0] , \CARRYB[34][51] , \CARRYB[34][50] , \CARRYB[34][49] ,
         \CARRYB[34][48] , \CARRYB[34][47] , \CARRYB[34][46] ,
         \CARRYB[34][45] , \CARRYB[34][44] , \CARRYB[34][43] ,
         \CARRYB[34][42] , \CARRYB[34][41] , \CARRYB[34][40] ,
         \CARRYB[34][39] , \CARRYB[34][38] , \CARRYB[34][37] ,
         \CARRYB[34][36] , \CARRYB[34][35] , \CARRYB[34][34] ,
         \CARRYB[34][33] , \CARRYB[34][32] , \CARRYB[34][31] ,
         \CARRYB[34][30] , \CARRYB[34][29] , \CARRYB[34][28] ,
         \CARRYB[34][27] , \CARRYB[34][26] , \CARRYB[34][25] ,
         \CARRYB[34][24] , \CARRYB[34][23] , \CARRYB[34][22] ,
         \CARRYB[34][21] , \CARRYB[34][20] , \CARRYB[34][19] ,
         \CARRYB[34][18] , \CARRYB[34][17] , \CARRYB[34][16] ,
         \CARRYB[34][15] , \CARRYB[34][14] , \CARRYB[34][13] ,
         \CARRYB[34][12] , \CARRYB[34][11] , \CARRYB[34][10] , \CARRYB[34][9] ,
         \CARRYB[34][8] , \CARRYB[34][7] , \CARRYB[34][6] , \CARRYB[34][5] ,
         \CARRYB[34][4] , \CARRYB[34][3] , \CARRYB[34][2] , \CARRYB[34][1] ,
         \CARRYB[34][0] , \CARRYB[33][51] , \CARRYB[33][50] , \CARRYB[33][49] ,
         \CARRYB[33][48] , \CARRYB[33][47] , \CARRYB[33][46] ,
         \CARRYB[33][45] , \CARRYB[33][44] , \CARRYB[33][43] ,
         \CARRYB[33][42] , \CARRYB[33][41] , \CARRYB[33][40] ,
         \CARRYB[33][39] , \CARRYB[33][38] , \CARRYB[33][37] ,
         \CARRYB[33][36] , \SUMB[43][17] , \SUMB[43][16] , \SUMB[43][15] ,
         \SUMB[43][14] , \SUMB[43][13] , \SUMB[43][12] , \SUMB[43][11] ,
         \SUMB[43][10] , \SUMB[43][9] , \SUMB[43][8] , \SUMB[43][7] ,
         \SUMB[43][6] , \SUMB[43][5] , \SUMB[43][4] , \SUMB[43][3] ,
         \SUMB[43][2] , \SUMB[43][1] , \SUMB[42][51] , \SUMB[42][50] ,
         \SUMB[42][49] , \SUMB[42][48] , \SUMB[42][47] , \SUMB[42][46] ,
         \SUMB[42][45] , \SUMB[42][44] , \SUMB[42][43] , \SUMB[42][42] ,
         \SUMB[42][41] , \SUMB[42][40] , \SUMB[42][39] , \SUMB[42][38] ,
         \SUMB[42][37] , \SUMB[42][36] , \SUMB[42][35] , \SUMB[42][34] ,
         \SUMB[42][33] , \SUMB[42][32] , \SUMB[42][31] , \SUMB[42][30] ,
         \SUMB[42][29] , \SUMB[42][28] , \SUMB[42][27] , \SUMB[42][26] ,
         \SUMB[42][25] , \SUMB[42][24] , \SUMB[42][23] , \SUMB[42][22] ,
         \SUMB[42][21] , \SUMB[42][20] , \SUMB[42][19] , \SUMB[42][18] ,
         \SUMB[42][17] , \SUMB[42][16] , \SUMB[42][15] , \SUMB[42][14] ,
         \SUMB[42][13] , \SUMB[42][12] , \SUMB[42][11] , \SUMB[42][10] ,
         \SUMB[42][9] , \SUMB[42][8] , \SUMB[42][7] , \SUMB[42][6] ,
         \SUMB[42][5] , \SUMB[42][4] , \SUMB[42][3] , \SUMB[42][2] ,
         \SUMB[42][1] , \SUMB[41][51] , \SUMB[41][50] , \SUMB[41][49] ,
         \SUMB[41][48] , \SUMB[41][47] , \SUMB[41][46] , \SUMB[41][45] ,
         \SUMB[41][44] , \SUMB[41][43] , \SUMB[41][42] , \SUMB[41][41] ,
         \SUMB[41][40] , \SUMB[41][39] , \SUMB[41][38] , \SUMB[41][37] ,
         \SUMB[41][36] , \SUMB[41][35] , \SUMB[41][34] , \SUMB[41][33] ,
         \SUMB[41][32] , \SUMB[41][31] , \SUMB[41][30] , \SUMB[41][29] ,
         \SUMB[41][28] , \SUMB[41][27] , \SUMB[41][26] , \SUMB[41][25] ,
         \SUMB[41][24] , \SUMB[41][23] , \SUMB[41][22] , \SUMB[41][21] ,
         \SUMB[41][20] , \SUMB[41][19] , \SUMB[41][18] , \SUMB[41][17] ,
         \SUMB[41][16] , \SUMB[41][15] , \SUMB[41][14] , \SUMB[41][13] ,
         \SUMB[41][12] , \SUMB[41][11] , \SUMB[41][10] , \SUMB[41][9] ,
         \SUMB[41][8] , \SUMB[41][7] , \SUMB[41][6] , \SUMB[41][5] ,
         \SUMB[41][4] , \SUMB[41][3] , \SUMB[41][2] , \SUMB[41][1] ,
         \SUMB[40][51] , \SUMB[40][50] , \SUMB[40][49] , \SUMB[40][48] ,
         \SUMB[40][47] , \SUMB[40][46] , \SUMB[40][45] , \SUMB[40][44] ,
         \SUMB[40][43] , \SUMB[40][42] , \SUMB[40][41] , \SUMB[40][40] ,
         \SUMB[40][39] , \SUMB[40][38] , \SUMB[40][37] , \SUMB[40][36] ,
         \SUMB[40][35] , \SUMB[40][34] , \SUMB[40][33] , \SUMB[40][32] ,
         \SUMB[40][31] , \SUMB[40][30] , \SUMB[40][29] , \SUMB[40][28] ,
         \SUMB[40][27] , \SUMB[40][26] , \SUMB[40][25] , \SUMB[40][24] ,
         \SUMB[40][23] , \SUMB[40][22] , \SUMB[40][21] , \SUMB[40][20] ,
         \SUMB[40][19] , \SUMB[40][18] , \SUMB[40][17] , \SUMB[40][16] ,
         \SUMB[40][15] , \SUMB[40][14] , \SUMB[40][13] , \SUMB[40][12] ,
         \SUMB[40][11] , \SUMB[40][10] , \SUMB[40][9] , \SUMB[40][8] ,
         \SUMB[40][7] , \SUMB[40][6] , \SUMB[40][5] , \SUMB[40][4] ,
         \SUMB[40][3] , \SUMB[40][2] , \SUMB[40][1] , \SUMB[39][51] ,
         \SUMB[39][50] , \SUMB[39][49] , \SUMB[39][48] , \SUMB[39][47] ,
         \SUMB[39][46] , \SUMB[39][45] , \SUMB[39][44] , \SUMB[39][43] ,
         \SUMB[39][42] , \SUMB[39][41] , \SUMB[39][40] , \SUMB[39][39] ,
         \SUMB[39][38] , \SUMB[39][37] , \SUMB[39][36] , \SUMB[39][35] ,
         \SUMB[39][34] , \SUMB[39][33] , \SUMB[39][32] , \SUMB[39][31] ,
         \SUMB[39][30] , \SUMB[39][29] , \SUMB[39][28] , \SUMB[39][27] ,
         \SUMB[39][26] , \SUMB[39][25] , \SUMB[39][24] , \SUMB[39][23] ,
         \SUMB[39][22] , \SUMB[39][21] , \SUMB[39][20] , \SUMB[39][19] ,
         \SUMB[39][18] , \SUMB[39][17] , \SUMB[39][16] , \SUMB[39][15] ,
         \SUMB[39][14] , \SUMB[39][13] , \SUMB[39][12] , \SUMB[39][11] ,
         \SUMB[39][10] , \SUMB[39][9] , \SUMB[39][8] , \SUMB[39][7] ,
         \SUMB[39][6] , \SUMB[39][5] , \SUMB[39][4] , \SUMB[39][3] ,
         \SUMB[39][2] , \SUMB[39][1] , \SUMB[38][51] , \SUMB[38][50] ,
         \SUMB[38][49] , \SUMB[38][48] , \SUMB[38][47] , \SUMB[38][46] ,
         \SUMB[38][45] , \SUMB[38][44] , \SUMB[38][43] , \SUMB[38][42] ,
         \SUMB[38][41] , \SUMB[38][40] , \SUMB[38][39] , \SUMB[38][38] ,
         \SUMB[38][37] , \SUMB[38][36] , \SUMB[38][35] , \SUMB[38][34] ,
         \SUMB[38][33] , \SUMB[38][32] , \SUMB[38][31] , \SUMB[38][30] ,
         \SUMB[38][29] , \SUMB[38][28] , \SUMB[38][27] , \SUMB[38][26] ,
         \SUMB[38][25] , \SUMB[38][24] , \SUMB[38][23] , \SUMB[38][22] ,
         \SUMB[38][21] , \SUMB[38][20] , \SUMB[38][19] , \SUMB[38][18] ,
         \SUMB[38][17] , \SUMB[38][16] , \SUMB[38][15] , \SUMB[38][14] ,
         \SUMB[38][13] , \SUMB[38][12] , \SUMB[38][11] , \SUMB[38][10] ,
         \SUMB[38][9] , \SUMB[38][8] , \SUMB[38][7] , \SUMB[38][6] ,
         \SUMB[38][5] , \SUMB[38][4] , \SUMB[38][3] , \SUMB[38][2] ,
         \SUMB[38][1] , \SUMB[37][51] , \SUMB[37][50] , \SUMB[37][49] ,
         \SUMB[37][48] , \SUMB[37][47] , \SUMB[37][46] , \SUMB[37][45] ,
         \SUMB[37][44] , \SUMB[37][43] , \SUMB[37][42] , \SUMB[37][41] ,
         \SUMB[37][40] , \SUMB[37][39] , \SUMB[37][38] , \SUMB[37][37] ,
         \SUMB[37][36] , \SUMB[37][35] , \SUMB[37][34] , \SUMB[37][33] ,
         \SUMB[37][32] , \SUMB[37][31] , \SUMB[37][30] , \SUMB[37][29] ,
         \SUMB[37][28] , \SUMB[37][27] , \SUMB[37][26] , \SUMB[37][25] ,
         \SUMB[37][24] , \SUMB[37][23] , \SUMB[37][22] , \SUMB[37][21] ,
         \SUMB[37][20] , \SUMB[37][19] , \SUMB[37][18] , \SUMB[37][17] ,
         \SUMB[37][16] , \SUMB[37][15] , \SUMB[37][14] , \SUMB[37][13] ,
         \SUMB[37][12] , \SUMB[37][11] , \SUMB[37][10] , \SUMB[37][9] ,
         \SUMB[37][8] , \SUMB[37][7] , \SUMB[37][6] , \SUMB[37][5] ,
         \SUMB[37][4] , \SUMB[37][3] , \SUMB[37][2] , \SUMB[37][1] ,
         \SUMB[36][51] , \SUMB[36][50] , \SUMB[36][49] , \SUMB[36][48] ,
         \SUMB[36][47] , \SUMB[36][46] , \SUMB[36][45] , \SUMB[36][44] ,
         \SUMB[36][43] , \SUMB[36][42] , \SUMB[36][41] , \SUMB[36][40] ,
         \SUMB[36][39] , \SUMB[36][38] , \SUMB[36][37] , \SUMB[36][36] ,
         \SUMB[36][35] , \SUMB[36][34] , \SUMB[36][33] , \SUMB[36][32] ,
         \SUMB[36][31] , \SUMB[36][30] , \SUMB[36][29] , \SUMB[36][28] ,
         \SUMB[36][27] , \SUMB[36][26] , \SUMB[36][25] , \SUMB[36][24] ,
         \SUMB[36][23] , \SUMB[36][22] , \SUMB[36][21] , \SUMB[36][20] ,
         \SUMB[36][19] , \SUMB[36][18] , \SUMB[36][17] , \SUMB[36][16] ,
         \SUMB[36][15] , \SUMB[36][14] , \SUMB[36][13] , \SUMB[36][12] ,
         \SUMB[36][11] , \SUMB[36][10] , \SUMB[36][9] , \SUMB[36][8] ,
         \SUMB[36][7] , \SUMB[36][6] , \SUMB[36][5] , \SUMB[36][4] ,
         \SUMB[36][3] , \SUMB[36][2] , \SUMB[36][1] , \SUMB[35][51] ,
         \SUMB[35][50] , \SUMB[35][49] , \SUMB[35][48] , \SUMB[35][47] ,
         \SUMB[35][46] , \SUMB[35][45] , \SUMB[35][44] , \SUMB[35][43] ,
         \SUMB[35][42] , \SUMB[35][41] , \SUMB[35][40] , \SUMB[35][39] ,
         \SUMB[35][38] , \SUMB[35][37] , \SUMB[35][36] , \SUMB[35][35] ,
         \SUMB[35][34] , \SUMB[35][33] , \SUMB[35][32] , \SUMB[35][31] ,
         \SUMB[35][30] , \SUMB[35][29] , \SUMB[35][28] , \SUMB[35][27] ,
         \SUMB[35][26] , \SUMB[35][25] , \SUMB[35][24] , \SUMB[35][23] ,
         \SUMB[35][22] , \SUMB[35][21] , \SUMB[35][20] , \SUMB[35][19] ,
         \SUMB[35][18] , \SUMB[35][17] , \SUMB[35][16] , \SUMB[35][15] ,
         \SUMB[35][14] , \SUMB[35][13] , \SUMB[35][12] , \SUMB[35][11] ,
         \SUMB[35][10] , \SUMB[35][9] , \SUMB[35][8] , \SUMB[35][7] ,
         \SUMB[35][6] , \SUMB[35][5] , \SUMB[35][4] , \SUMB[35][3] ,
         \SUMB[35][2] , \SUMB[35][1] , \SUMB[34][51] , \SUMB[34][50] ,
         \SUMB[34][49] , \SUMB[34][48] , \SUMB[34][47] , \SUMB[34][46] ,
         \SUMB[34][45] , \SUMB[34][44] , \SUMB[34][43] , \SUMB[34][42] ,
         \SUMB[34][41] , \SUMB[34][40] , \SUMB[34][39] , \SUMB[34][38] ,
         \SUMB[34][37] , \SUMB[34][36] , \SUMB[34][35] , \SUMB[34][34] ,
         \SUMB[34][33] , \SUMB[34][32] , \SUMB[34][31] , \SUMB[34][30] ,
         \SUMB[34][29] , \SUMB[34][28] , \SUMB[34][27] , \SUMB[34][26] ,
         \SUMB[34][25] , \SUMB[34][24] , \SUMB[34][23] , \SUMB[34][22] ,
         \SUMB[34][21] , \SUMB[34][20] , \SUMB[34][19] , \SUMB[34][18] ,
         \SUMB[34][17] , \SUMB[34][16] , \SUMB[34][15] , \SUMB[34][14] ,
         \SUMB[34][13] , \SUMB[34][12] , \SUMB[34][11] , \SUMB[34][10] ,
         \SUMB[34][9] , \SUMB[34][8] , \SUMB[34][7] , \SUMB[34][6] ,
         \SUMB[34][5] , \SUMB[34][4] , \SUMB[34][3] , \SUMB[34][2] ,
         \SUMB[34][1] , \SUMB[33][51] , \SUMB[33][50] , \SUMB[33][49] ,
         \SUMB[33][48] , \SUMB[33][47] , \SUMB[33][46] , \SUMB[33][45] ,
         \SUMB[33][44] , \SUMB[33][43] , \SUMB[33][42] , \SUMB[33][41] ,
         \SUMB[33][40] , \SUMB[33][39] , \SUMB[33][38] , \SUMB[33][37] ,
         \SUMB[33][36] , \CARRYB[52][51] , \CARRYB[52][50] , \CARRYB[52][49] ,
         \CARRYB[52][48] , \CARRYB[52][47] , \CARRYB[52][46] ,
         \CARRYB[52][45] , \CARRYB[52][44] , \CARRYB[52][43] ,
         \CARRYB[52][42] , \CARRYB[52][41] , \CARRYB[52][40] ,
         \CARRYB[52][39] , \CARRYB[52][38] , \CARRYB[52][37] ,
         \CARRYB[52][36] , \CARRYB[52][35] , \CARRYB[52][34] ,
         \CARRYB[52][33] , \CARRYB[52][32] , \CARRYB[52][31] ,
         \CARRYB[52][30] , \CARRYB[52][29] , \CARRYB[52][28] ,
         \CARRYB[52][27] , \CARRYB[52][26] , \CARRYB[52][25] ,
         \CARRYB[52][24] , \CARRYB[52][23] , \CARRYB[52][22] ,
         \CARRYB[52][21] , \CARRYB[52][20] , \CARRYB[52][19] ,
         \CARRYB[52][18] , \CARRYB[52][17] , \CARRYB[52][16] ,
         \CARRYB[52][15] , \CARRYB[52][14] , \CARRYB[52][13] ,
         \CARRYB[52][12] , \CARRYB[52][11] , \CARRYB[52][10] , \CARRYB[52][9] ,
         \CARRYB[52][8] , \CARRYB[52][7] , \CARRYB[52][6] , \CARRYB[52][5] ,
         \CARRYB[52][4] , \CARRYB[52][3] , \CARRYB[52][2] , \CARRYB[52][1] ,
         \CARRYB[52][0] , \CARRYB[51][51] , \CARRYB[51][50] , \CARRYB[51][49] ,
         \CARRYB[51][48] , \CARRYB[51][47] , \CARRYB[51][46] ,
         \CARRYB[51][45] , \CARRYB[51][44] , \CARRYB[51][43] ,
         \CARRYB[51][42] , \CARRYB[51][41] , \CARRYB[51][40] ,
         \CARRYB[51][39] , \CARRYB[51][38] , \CARRYB[51][37] ,
         \CARRYB[51][36] , \CARRYB[51][35] , \CARRYB[51][34] ,
         \CARRYB[51][33] , \CARRYB[51][32] , \CARRYB[51][31] ,
         \CARRYB[51][30] , \CARRYB[51][29] , \CARRYB[51][28] ,
         \CARRYB[51][27] , \CARRYB[51][26] , \CARRYB[51][25] ,
         \CARRYB[51][24] , \CARRYB[51][23] , \CARRYB[51][22] ,
         \CARRYB[51][21] , \CARRYB[51][20] , \CARRYB[51][19] ,
         \CARRYB[51][18] , \CARRYB[51][17] , \CARRYB[51][16] ,
         \CARRYB[51][15] , \CARRYB[51][14] , \CARRYB[51][13] ,
         \CARRYB[51][12] , \CARRYB[51][11] , \CARRYB[51][10] , \CARRYB[51][9] ,
         \CARRYB[51][8] , \CARRYB[51][7] , \CARRYB[51][6] , \CARRYB[51][5] ,
         \CARRYB[51][4] , \CARRYB[51][3] , \CARRYB[51][2] , \CARRYB[51][1] ,
         \CARRYB[51][0] , \CARRYB[50][51] , \CARRYB[50][50] , \CARRYB[50][49] ,
         \CARRYB[50][48] , \CARRYB[50][47] , \CARRYB[50][46] ,
         \CARRYB[50][45] , \CARRYB[50][44] , \CARRYB[50][43] ,
         \CARRYB[50][42] , \CARRYB[50][41] , \CARRYB[50][40] ,
         \CARRYB[50][39] , \CARRYB[50][38] , \CARRYB[50][37] ,
         \CARRYB[50][36] , \CARRYB[50][35] , \CARRYB[50][34] ,
         \CARRYB[50][33] , \CARRYB[50][32] , \CARRYB[50][31] ,
         \CARRYB[50][30] , \CARRYB[50][29] , \CARRYB[50][28] ,
         \CARRYB[50][27] , \CARRYB[50][26] , \CARRYB[50][25] ,
         \CARRYB[50][24] , \CARRYB[50][23] , \CARRYB[50][22] ,
         \CARRYB[50][21] , \CARRYB[50][20] , \CARRYB[50][19] ,
         \CARRYB[50][18] , \CARRYB[50][17] , \CARRYB[50][16] ,
         \CARRYB[50][15] , \CARRYB[50][14] , \CARRYB[50][13] ,
         \CARRYB[50][12] , \CARRYB[50][11] , \CARRYB[50][10] , \CARRYB[50][9] ,
         \CARRYB[50][8] , \CARRYB[50][7] , \CARRYB[50][6] , \CARRYB[50][5] ,
         \CARRYB[50][4] , \CARRYB[50][3] , \CARRYB[50][2] , \CARRYB[50][1] ,
         \CARRYB[50][0] , \CARRYB[49][51] , \CARRYB[49][50] , \CARRYB[49][49] ,
         \CARRYB[49][48] , \CARRYB[49][47] , \CARRYB[49][46] ,
         \CARRYB[49][45] , \CARRYB[49][44] , \CARRYB[49][43] ,
         \CARRYB[49][42] , \CARRYB[49][41] , \CARRYB[49][40] ,
         \CARRYB[49][39] , \CARRYB[49][38] , \CARRYB[49][37] ,
         \CARRYB[49][36] , \CARRYB[49][35] , \CARRYB[49][34] ,
         \CARRYB[49][33] , \CARRYB[49][32] , \CARRYB[49][31] ,
         \CARRYB[49][30] , \CARRYB[49][29] , \CARRYB[49][28] ,
         \CARRYB[49][27] , \CARRYB[49][26] , \CARRYB[49][25] ,
         \CARRYB[49][24] , \CARRYB[49][23] , \CARRYB[49][22] ,
         \CARRYB[49][21] , \CARRYB[49][20] , \CARRYB[49][19] ,
         \CARRYB[49][18] , \CARRYB[49][17] , \CARRYB[49][16] ,
         \CARRYB[49][15] , \CARRYB[49][14] , \CARRYB[49][13] ,
         \CARRYB[49][12] , \CARRYB[49][11] , \CARRYB[49][10] , \CARRYB[49][9] ,
         \CARRYB[49][8] , \CARRYB[49][7] , \CARRYB[49][6] , \CARRYB[49][5] ,
         \CARRYB[49][4] , \CARRYB[49][3] , \CARRYB[49][2] , \CARRYB[49][1] ,
         \CARRYB[49][0] , \CARRYB[48][51] , \CARRYB[48][50] , \CARRYB[48][49] ,
         \CARRYB[48][48] , \CARRYB[48][47] , \CARRYB[48][46] ,
         \CARRYB[48][45] , \CARRYB[48][44] , \CARRYB[48][43] ,
         \CARRYB[48][42] , \CARRYB[48][41] , \CARRYB[48][40] ,
         \CARRYB[48][39] , \CARRYB[48][38] , \CARRYB[48][37] ,
         \CARRYB[48][36] , \CARRYB[48][35] , \CARRYB[48][34] ,
         \CARRYB[48][33] , \CARRYB[48][32] , \CARRYB[48][31] ,
         \CARRYB[48][30] , \CARRYB[48][29] , \CARRYB[48][28] ,
         \CARRYB[48][27] , \CARRYB[48][26] , \CARRYB[48][25] ,
         \CARRYB[48][24] , \CARRYB[48][23] , \CARRYB[48][22] ,
         \CARRYB[48][21] , \CARRYB[48][20] , \CARRYB[48][19] ,
         \CARRYB[48][18] , \CARRYB[48][17] , \CARRYB[48][16] ,
         \CARRYB[48][15] , \CARRYB[48][14] , \CARRYB[48][13] ,
         \CARRYB[48][12] , \CARRYB[48][11] , \CARRYB[48][10] , \CARRYB[48][9] ,
         \CARRYB[48][8] , \CARRYB[48][7] , \CARRYB[48][6] , \CARRYB[48][5] ,
         \CARRYB[48][4] , \CARRYB[48][3] , \CARRYB[48][2] , \CARRYB[48][1] ,
         \CARRYB[48][0] , \CARRYB[47][51] , \CARRYB[47][50] , \CARRYB[47][49] ,
         \CARRYB[47][48] , \CARRYB[47][47] , \CARRYB[47][46] ,
         \CARRYB[47][45] , \CARRYB[47][44] , \CARRYB[47][43] ,
         \CARRYB[47][42] , \CARRYB[47][41] , \CARRYB[47][40] ,
         \CARRYB[47][39] , \CARRYB[47][38] , \CARRYB[47][37] ,
         \CARRYB[47][36] , \CARRYB[47][35] , \CARRYB[47][34] ,
         \CARRYB[47][33] , \CARRYB[47][32] , \CARRYB[47][31] ,
         \CARRYB[47][30] , \CARRYB[47][29] , \CARRYB[47][28] ,
         \CARRYB[47][27] , \CARRYB[47][26] , \CARRYB[47][25] ,
         \CARRYB[47][24] , \CARRYB[47][23] , \CARRYB[47][22] ,
         \CARRYB[47][21] , \CARRYB[47][20] , \CARRYB[47][19] ,
         \CARRYB[47][18] , \CARRYB[47][17] , \CARRYB[47][16] ,
         \CARRYB[47][15] , \CARRYB[47][14] , \CARRYB[47][13] ,
         \CARRYB[47][12] , \CARRYB[47][11] , \CARRYB[47][10] , \CARRYB[47][9] ,
         \CARRYB[47][8] , \CARRYB[47][7] , \CARRYB[47][6] , \CARRYB[47][5] ,
         \CARRYB[47][4] , \CARRYB[47][3] , \CARRYB[47][2] , \CARRYB[47][1] ,
         \CARRYB[47][0] , \CARRYB[46][51] , \CARRYB[46][50] , \CARRYB[46][49] ,
         \CARRYB[46][48] , \CARRYB[46][47] , \CARRYB[46][46] ,
         \CARRYB[46][45] , \CARRYB[46][44] , \CARRYB[46][43] ,
         \CARRYB[46][42] , \CARRYB[46][41] , \CARRYB[46][40] ,
         \CARRYB[46][39] , \CARRYB[46][38] , \CARRYB[46][37] ,
         \CARRYB[46][36] , \CARRYB[46][35] , \CARRYB[46][34] ,
         \CARRYB[46][33] , \CARRYB[46][32] , \CARRYB[46][31] ,
         \CARRYB[46][30] , \CARRYB[46][29] , \CARRYB[46][28] ,
         \CARRYB[46][27] , \CARRYB[46][26] , \CARRYB[46][25] ,
         \CARRYB[46][24] , \CARRYB[46][23] , \CARRYB[46][22] ,
         \CARRYB[46][21] , \CARRYB[46][20] , \CARRYB[46][19] ,
         \CARRYB[46][18] , \CARRYB[46][17] , \CARRYB[46][16] ,
         \CARRYB[46][15] , \CARRYB[46][14] , \CARRYB[46][13] ,
         \CARRYB[46][12] , \CARRYB[46][11] , \CARRYB[46][10] , \CARRYB[46][9] ,
         \CARRYB[46][8] , \CARRYB[46][7] , \CARRYB[46][6] , \CARRYB[46][5] ,
         \CARRYB[46][4] , \CARRYB[46][3] , \CARRYB[46][2] , \CARRYB[46][1] ,
         \CARRYB[46][0] , \CARRYB[45][51] , \CARRYB[45][50] , \CARRYB[45][49] ,
         \CARRYB[45][48] , \CARRYB[45][47] , \CARRYB[45][46] ,
         \CARRYB[45][45] , \CARRYB[45][44] , \CARRYB[45][43] ,
         \CARRYB[45][42] , \CARRYB[45][41] , \CARRYB[45][40] ,
         \CARRYB[45][39] , \CARRYB[45][38] , \CARRYB[45][37] ,
         \CARRYB[45][36] , \CARRYB[45][35] , \CARRYB[45][34] ,
         \CARRYB[45][33] , \CARRYB[45][32] , \CARRYB[45][31] ,
         \CARRYB[45][30] , \CARRYB[45][29] , \CARRYB[45][28] ,
         \CARRYB[45][27] , \CARRYB[45][26] , \CARRYB[45][25] ,
         \CARRYB[45][24] , \CARRYB[45][23] , \CARRYB[45][22] ,
         \CARRYB[45][21] , \CARRYB[45][20] , \CARRYB[45][19] ,
         \CARRYB[45][18] , \CARRYB[45][17] , \CARRYB[45][16] ,
         \CARRYB[45][15] , \CARRYB[45][14] , \CARRYB[45][13] ,
         \CARRYB[45][12] , \CARRYB[45][11] , \CARRYB[45][10] , \CARRYB[45][9] ,
         \CARRYB[45][8] , \CARRYB[45][7] , \CARRYB[45][6] , \CARRYB[45][5] ,
         \CARRYB[45][4] , \CARRYB[45][3] , \CARRYB[45][2] , \CARRYB[45][1] ,
         \CARRYB[45][0] , \CARRYB[44][51] , \CARRYB[44][50] , \CARRYB[44][49] ,
         \CARRYB[44][48] , \CARRYB[44][47] , \CARRYB[44][46] ,
         \CARRYB[44][45] , \CARRYB[44][44] , \CARRYB[44][43] ,
         \CARRYB[44][42] , \CARRYB[44][41] , \CARRYB[44][40] ,
         \CARRYB[44][39] , \CARRYB[44][38] , \CARRYB[44][37] ,
         \CARRYB[44][36] , \CARRYB[44][35] , \CARRYB[44][34] ,
         \CARRYB[44][33] , \CARRYB[44][32] , \CARRYB[44][31] ,
         \CARRYB[44][30] , \CARRYB[44][29] , \CARRYB[44][28] ,
         \CARRYB[44][27] , \CARRYB[44][26] , \CARRYB[44][25] ,
         \CARRYB[44][24] , \CARRYB[44][23] , \CARRYB[44][22] ,
         \CARRYB[44][21] , \CARRYB[44][20] , \CARRYB[44][19] ,
         \CARRYB[44][18] , \CARRYB[44][17] , \CARRYB[44][16] ,
         \CARRYB[44][15] , \CARRYB[44][14] , \CARRYB[44][13] ,
         \CARRYB[44][12] , \CARRYB[44][11] , \CARRYB[44][10] , \CARRYB[44][9] ,
         \CARRYB[44][8] , \CARRYB[44][7] , \CARRYB[44][6] , \CARRYB[44][5] ,
         \CARRYB[44][4] , \CARRYB[44][3] , \CARRYB[44][2] , \CARRYB[44][1] ,
         \CARRYB[44][0] , \CARRYB[43][51] , \CARRYB[43][50] , \CARRYB[43][49] ,
         \CARRYB[43][48] , \CARRYB[43][47] , \CARRYB[43][46] ,
         \CARRYB[43][45] , \CARRYB[43][44] , \CARRYB[43][43] ,
         \CARRYB[43][42] , \CARRYB[43][41] , \CARRYB[43][40] ,
         \CARRYB[43][39] , \CARRYB[43][38] , \CARRYB[43][37] ,
         \CARRYB[43][36] , \CARRYB[43][35] , \CARRYB[43][34] ,
         \CARRYB[43][33] , \CARRYB[43][32] , \CARRYB[43][31] ,
         \CARRYB[43][30] , \CARRYB[43][29] , \CARRYB[43][28] ,
         \CARRYB[43][27] , \CARRYB[43][26] , \CARRYB[43][25] ,
         \CARRYB[43][24] , \CARRYB[43][23] , \CARRYB[43][22] ,
         \CARRYB[43][21] , \CARRYB[43][20] , \CARRYB[43][19] ,
         \CARRYB[43][18] , \SUMB[52][51] , \SUMB[52][50] , \SUMB[52][49] ,
         \SUMB[52][48] , \SUMB[52][47] , \SUMB[52][46] , \SUMB[52][45] ,
         \SUMB[52][44] , \SUMB[52][43] , \SUMB[52][42] , \SUMB[52][41] ,
         \SUMB[52][40] , \SUMB[52][39] , \SUMB[52][38] , \SUMB[52][37] ,
         \SUMB[52][36] , \SUMB[52][35] , \SUMB[52][34] , \SUMB[52][33] ,
         \SUMB[52][32] , \SUMB[52][31] , \SUMB[52][30] , \SUMB[52][29] ,
         \SUMB[52][28] , \SUMB[52][27] , \SUMB[52][26] , \SUMB[52][25] ,
         \SUMB[52][24] , \SUMB[52][23] , \SUMB[52][22] , \SUMB[52][21] ,
         \SUMB[52][20] , \SUMB[52][19] , \SUMB[52][18] , \SUMB[52][17] ,
         \SUMB[52][16] , \SUMB[52][15] , \SUMB[52][14] , \SUMB[52][13] ,
         \SUMB[52][12] , \SUMB[52][11] , \SUMB[52][10] , \SUMB[52][9] ,
         \SUMB[52][8] , \SUMB[52][7] , \SUMB[52][6] , \SUMB[52][5] ,
         \SUMB[52][4] , \SUMB[52][3] , \SUMB[52][2] , \SUMB[52][1] ,
         \SUMB[52][0] , \SUMB[51][51] , \SUMB[51][50] , \SUMB[51][49] ,
         \SUMB[51][48] , \SUMB[51][47] , \SUMB[51][46] , \SUMB[51][45] ,
         \SUMB[51][44] , \SUMB[51][43] , \SUMB[51][42] , \SUMB[51][41] ,
         \SUMB[51][40] , \SUMB[51][39] , \SUMB[51][38] , \SUMB[51][37] ,
         \SUMB[51][36] , \SUMB[51][35] , \SUMB[51][34] , \SUMB[51][33] ,
         \SUMB[51][32] , \SUMB[51][31] , \SUMB[51][30] , \SUMB[51][29] ,
         \SUMB[51][28] , \SUMB[51][27] , \SUMB[51][26] , \SUMB[51][25] ,
         \SUMB[51][24] , \SUMB[51][23] , \SUMB[51][22] , \SUMB[51][21] ,
         \SUMB[51][20] , \SUMB[51][19] , \SUMB[51][18] , \SUMB[51][17] ,
         \SUMB[51][16] , \SUMB[51][15] , \SUMB[51][14] , \SUMB[51][13] ,
         \SUMB[51][12] , \SUMB[51][11] , \SUMB[51][10] , \SUMB[51][9] ,
         \SUMB[51][8] , \SUMB[51][7] , \SUMB[51][6] , \SUMB[51][5] ,
         \SUMB[51][4] , \SUMB[51][3] , \SUMB[51][2] , \SUMB[51][1] ,
         \SUMB[50][51] , \SUMB[50][50] , \SUMB[50][49] , \SUMB[50][48] ,
         \SUMB[50][47] , \SUMB[50][46] , \SUMB[50][45] , \SUMB[50][44] ,
         \SUMB[50][43] , \SUMB[50][42] , \SUMB[50][41] , \SUMB[50][40] ,
         \SUMB[50][39] , \SUMB[50][38] , \SUMB[50][37] , \SUMB[50][36] ,
         \SUMB[50][35] , \SUMB[50][34] , \SUMB[50][33] , \SUMB[50][32] ,
         \SUMB[50][31] , \SUMB[50][30] , \SUMB[50][29] , \SUMB[50][28] ,
         \SUMB[50][27] , \SUMB[50][26] , \SUMB[50][25] , \SUMB[50][24] ,
         \SUMB[50][23] , \SUMB[50][22] , \SUMB[50][21] , \SUMB[50][20] ,
         \SUMB[50][19] , \SUMB[50][18] , \SUMB[50][17] , \SUMB[50][16] ,
         \SUMB[50][15] , \SUMB[50][14] , \SUMB[50][13] , \SUMB[50][12] ,
         \SUMB[50][11] , \SUMB[50][10] , \SUMB[50][9] , \SUMB[50][8] ,
         \SUMB[50][7] , \SUMB[50][6] , \SUMB[50][5] , \SUMB[50][4] ,
         \SUMB[50][3] , \SUMB[50][2] , \SUMB[50][1] , \SUMB[49][51] ,
         \SUMB[49][50] , \SUMB[49][49] , \SUMB[49][48] , \SUMB[49][47] ,
         \SUMB[49][46] , \SUMB[49][45] , \SUMB[49][44] , \SUMB[49][43] ,
         \SUMB[49][42] , \SUMB[49][41] , \SUMB[49][40] , \SUMB[49][39] ,
         \SUMB[49][38] , \SUMB[49][37] , \SUMB[49][36] , \SUMB[49][35] ,
         \SUMB[49][34] , \SUMB[49][33] , \SUMB[49][32] , \SUMB[49][31] ,
         \SUMB[49][30] , \SUMB[49][29] , \SUMB[49][28] , \SUMB[49][27] ,
         \SUMB[49][26] , \SUMB[49][25] , \SUMB[49][24] , \SUMB[49][23] ,
         \SUMB[49][22] , \SUMB[49][21] , \SUMB[49][20] , \SUMB[49][19] ,
         \SUMB[49][18] , \SUMB[49][17] , \SUMB[49][16] , \SUMB[49][15] ,
         \SUMB[49][14] , \SUMB[49][13] , \SUMB[49][12] , \SUMB[49][11] ,
         \SUMB[49][10] , \SUMB[49][9] , \SUMB[49][8] , \SUMB[49][7] ,
         \SUMB[49][6] , \SUMB[49][5] , \SUMB[49][4] , \SUMB[49][3] ,
         \SUMB[49][2] , \SUMB[49][1] , \SUMB[48][51] , \SUMB[48][50] ,
         \SUMB[48][49] , \SUMB[48][48] , \SUMB[48][47] , \SUMB[48][46] ,
         \SUMB[48][45] , \SUMB[48][44] , \SUMB[48][43] , \SUMB[48][42] ,
         \SUMB[48][41] , \SUMB[48][40] , \SUMB[48][39] , \SUMB[48][38] ,
         \SUMB[48][37] , \SUMB[48][36] , \SUMB[48][35] , \SUMB[48][34] ,
         \SUMB[48][33] , \SUMB[48][32] , \SUMB[48][31] , \SUMB[48][30] ,
         \SUMB[48][29] , \SUMB[48][28] , \SUMB[48][27] , \SUMB[48][26] ,
         \SUMB[48][25] , \SUMB[48][24] , \SUMB[48][23] , \SUMB[48][22] ,
         \SUMB[48][21] , \SUMB[48][20] , \SUMB[48][19] , \SUMB[48][18] ,
         \SUMB[48][17] , \SUMB[48][16] , \SUMB[48][15] , \SUMB[48][14] ,
         \SUMB[48][13] , \SUMB[48][12] , \SUMB[48][11] , \SUMB[48][10] ,
         \SUMB[48][9] , \SUMB[48][8] , \SUMB[48][7] , \SUMB[48][6] ,
         \SUMB[48][5] , \SUMB[48][4] , \SUMB[48][3] , \SUMB[48][2] ,
         \SUMB[48][1] , \SUMB[47][51] , \SUMB[47][50] , \SUMB[47][49] ,
         \SUMB[47][48] , \SUMB[47][47] , \SUMB[47][46] , \SUMB[47][45] ,
         \SUMB[47][44] , \SUMB[47][43] , \SUMB[47][42] , \SUMB[47][41] ,
         \SUMB[47][40] , \SUMB[47][39] , \SUMB[47][38] , \SUMB[47][37] ,
         \SUMB[47][36] , \SUMB[47][35] , \SUMB[47][34] , \SUMB[47][33] ,
         \SUMB[47][32] , \SUMB[47][31] , \SUMB[47][30] , \SUMB[47][29] ,
         \SUMB[47][28] , \SUMB[47][27] , \SUMB[47][26] , \SUMB[47][25] ,
         \SUMB[47][24] , \SUMB[47][23] , \SUMB[47][22] , \SUMB[47][21] ,
         \SUMB[47][20] , \SUMB[47][19] , \SUMB[47][18] , \SUMB[47][17] ,
         \SUMB[47][16] , \SUMB[47][15] , \SUMB[47][14] , \SUMB[47][13] ,
         \SUMB[47][12] , \SUMB[47][11] , \SUMB[47][10] , \SUMB[47][9] ,
         \SUMB[47][8] , \SUMB[47][7] , \SUMB[47][6] , \SUMB[47][5] ,
         \SUMB[47][4] , \SUMB[47][3] , \SUMB[47][2] , \SUMB[47][1] ,
         \SUMB[46][51] , \SUMB[46][50] , \SUMB[46][49] , \SUMB[46][48] ,
         \SUMB[46][47] , \SUMB[46][46] , \SUMB[46][45] , \SUMB[46][44] ,
         \SUMB[46][43] , \SUMB[46][42] , \SUMB[46][41] , \SUMB[46][40] ,
         \SUMB[46][39] , \SUMB[46][38] , \SUMB[46][37] , \SUMB[46][36] ,
         \SUMB[46][35] , \SUMB[46][34] , \SUMB[46][33] , \SUMB[46][32] ,
         \SUMB[46][31] , \SUMB[46][30] , \SUMB[46][29] , \SUMB[46][28] ,
         \SUMB[46][27] , \SUMB[46][26] , \SUMB[46][25] , \SUMB[46][24] ,
         \SUMB[46][23] , \SUMB[46][22] , \SUMB[46][21] , \SUMB[46][20] ,
         \SUMB[46][19] , \SUMB[46][18] , \SUMB[46][17] , \SUMB[46][16] ,
         \SUMB[46][15] , \SUMB[46][14] , \SUMB[46][13] , \SUMB[46][12] ,
         \SUMB[46][11] , \SUMB[46][10] , \SUMB[46][9] , \SUMB[46][8] ,
         \SUMB[46][7] , \SUMB[46][6] , \SUMB[46][5] , \SUMB[46][4] ,
         \SUMB[46][3] , \SUMB[46][2] , \SUMB[46][1] , \SUMB[45][51] ,
         \SUMB[45][50] , \SUMB[45][49] , \SUMB[45][48] , \SUMB[45][47] ,
         \SUMB[45][46] , \SUMB[45][45] , \SUMB[45][44] , \SUMB[45][43] ,
         \SUMB[45][42] , \SUMB[45][41] , \SUMB[45][40] , \SUMB[45][39] ,
         \SUMB[45][38] , \SUMB[45][37] , \SUMB[45][36] , \SUMB[45][35] ,
         \SUMB[45][34] , \SUMB[45][33] , \SUMB[45][32] , \SUMB[45][31] ,
         \SUMB[45][30] , \SUMB[45][29] , \SUMB[45][28] , \SUMB[45][27] ,
         \SUMB[45][26] , \SUMB[45][25] , \SUMB[45][24] , \SUMB[45][23] ,
         \SUMB[45][22] , \SUMB[45][21] , \SUMB[45][20] , \SUMB[45][19] ,
         \SUMB[45][18] , \SUMB[45][17] , \SUMB[45][16] , \SUMB[45][15] ,
         \SUMB[45][14] , \SUMB[45][13] , \SUMB[45][12] , \SUMB[45][11] ,
         \SUMB[45][10] , \SUMB[45][9] , \SUMB[45][8] , \SUMB[45][7] ,
         \SUMB[45][6] , \SUMB[45][5] , \SUMB[45][4] , \SUMB[45][3] ,
         \SUMB[45][2] , \SUMB[45][1] , \SUMB[44][51] , \SUMB[44][50] ,
         \SUMB[44][49] , \SUMB[44][48] , \SUMB[44][47] , \SUMB[44][46] ,
         \SUMB[44][45] , \SUMB[44][44] , \SUMB[44][43] , \SUMB[44][42] ,
         \SUMB[44][41] , \SUMB[44][40] , \SUMB[44][39] , \SUMB[44][38] ,
         \SUMB[44][37] , \SUMB[44][36] , \SUMB[44][35] , \SUMB[44][34] ,
         \SUMB[44][33] , \SUMB[44][32] , \SUMB[44][31] , \SUMB[44][30] ,
         \SUMB[44][29] , \SUMB[44][28] , \SUMB[44][27] , \SUMB[44][26] ,
         \SUMB[44][25] , \SUMB[44][24] , \SUMB[44][23] , \SUMB[44][22] ,
         \SUMB[44][21] , \SUMB[44][20] , \SUMB[44][19] , \SUMB[44][18] ,
         \SUMB[44][17] , \SUMB[44][16] , \SUMB[44][15] , \SUMB[44][14] ,
         \SUMB[44][13] , \SUMB[44][12] , \SUMB[44][11] , \SUMB[44][10] ,
         \SUMB[44][9] , \SUMB[44][8] , \SUMB[44][7] , \SUMB[44][6] ,
         \SUMB[44][5] , \SUMB[44][4] , \SUMB[44][3] , \SUMB[44][2] ,
         \SUMB[44][1] , \SUMB[43][51] , \SUMB[43][50] , \SUMB[43][49] ,
         \SUMB[43][48] , \SUMB[43][47] , \SUMB[43][46] , \SUMB[43][45] ,
         \SUMB[43][44] , \SUMB[43][43] , \SUMB[43][42] , \SUMB[43][41] ,
         \SUMB[43][40] , \SUMB[43][39] , \SUMB[43][38] , \SUMB[43][37] ,
         \SUMB[43][36] , \SUMB[43][35] , \SUMB[43][34] , \SUMB[43][33] ,
         \SUMB[43][32] , \SUMB[43][31] , \SUMB[43][30] , \SUMB[43][29] ,
         \SUMB[43][28] , \SUMB[43][27] , \SUMB[43][26] , \SUMB[43][25] ,
         \SUMB[43][24] , \SUMB[43][23] , \SUMB[43][22] , \SUMB[43][21] ,
         \SUMB[43][20] , \SUMB[43][19] , \SUMB[43][18] , n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480;
  wire   [51:2] CLA_SUM;

  FA_X1 S4_0 ( .A(\ab[52][0] ), .B(\CARRYB[51][0] ), .CI(\SUMB[51][1] ), .CO(
        \CARRYB[52][0] ), .S(\SUMB[52][0] ) );
  FA_X1 S4_1 ( .A(\ab[52][1] ), .B(\CARRYB[51][1] ), .CI(\SUMB[51][2] ), .CO(
        \CARRYB[52][1] ), .S(\SUMB[52][1] ) );
  FA_X1 S4_2 ( .A(\ab[52][2] ), .B(\CARRYB[51][2] ), .CI(\SUMB[51][3] ), .CO(
        \CARRYB[52][2] ), .S(\SUMB[52][2] ) );
  FA_X1 S4_3 ( .A(\ab[52][3] ), .B(\CARRYB[51][3] ), .CI(\SUMB[51][4] ), .CO(
        \CARRYB[52][3] ), .S(\SUMB[52][3] ) );
  FA_X1 S4_4 ( .A(\ab[52][4] ), .B(\CARRYB[51][4] ), .CI(\SUMB[51][5] ), .CO(
        \CARRYB[52][4] ), .S(\SUMB[52][4] ) );
  FA_X1 S4_5 ( .A(\ab[52][5] ), .B(\CARRYB[51][5] ), .CI(\SUMB[51][6] ), .CO(
        \CARRYB[52][5] ), .S(\SUMB[52][5] ) );
  FA_X1 S4_6 ( .A(\ab[52][6] ), .B(\CARRYB[51][6] ), .CI(\SUMB[51][7] ), .CO(
        \CARRYB[52][6] ), .S(\SUMB[52][6] ) );
  FA_X1 S4_7 ( .A(\ab[52][7] ), .B(\CARRYB[51][7] ), .CI(\SUMB[51][8] ), .CO(
        \CARRYB[52][7] ), .S(\SUMB[52][7] ) );
  FA_X1 S4_8 ( .A(\ab[52][8] ), .B(\CARRYB[51][8] ), .CI(\SUMB[51][9] ), .CO(
        \CARRYB[52][8] ), .S(\SUMB[52][8] ) );
  FA_X1 S4_9 ( .A(\ab[52][9] ), .B(\CARRYB[51][9] ), .CI(\SUMB[51][10] ), .CO(
        \CARRYB[52][9] ), .S(\SUMB[52][9] ) );
  FA_X1 S4_10 ( .A(\ab[52][10] ), .B(\CARRYB[51][10] ), .CI(\SUMB[51][11] ), 
        .CO(\CARRYB[52][10] ), .S(\SUMB[52][10] ) );
  FA_X1 S4_11 ( .A(\ab[52][11] ), .B(\CARRYB[51][11] ), .CI(\SUMB[51][12] ), 
        .CO(\CARRYB[52][11] ), .S(\SUMB[52][11] ) );
  FA_X1 S4_12 ( .A(\ab[52][12] ), .B(\CARRYB[51][12] ), .CI(\SUMB[51][13] ), 
        .CO(\CARRYB[52][12] ), .S(\SUMB[52][12] ) );
  FA_X1 S4_13 ( .A(\ab[52][13] ), .B(\CARRYB[51][13] ), .CI(\SUMB[51][14] ), 
        .CO(\CARRYB[52][13] ), .S(\SUMB[52][13] ) );
  FA_X1 S4_14 ( .A(\ab[52][14] ), .B(\CARRYB[51][14] ), .CI(\SUMB[51][15] ), 
        .CO(\CARRYB[52][14] ), .S(\SUMB[52][14] ) );
  FA_X1 S4_15 ( .A(\ab[52][15] ), .B(\CARRYB[51][15] ), .CI(\SUMB[51][16] ), 
        .CO(\CARRYB[52][15] ), .S(\SUMB[52][15] ) );
  FA_X1 S4_16 ( .A(\ab[52][16] ), .B(\CARRYB[51][16] ), .CI(\SUMB[51][17] ), 
        .CO(\CARRYB[52][16] ), .S(\SUMB[52][16] ) );
  FA_X1 S4_17 ( .A(\ab[52][17] ), .B(\CARRYB[51][17] ), .CI(\SUMB[51][18] ), 
        .CO(\CARRYB[52][17] ), .S(\SUMB[52][17] ) );
  FA_X1 S4_18 ( .A(\ab[52][18] ), .B(\CARRYB[51][18] ), .CI(\SUMB[51][19] ), 
        .CO(\CARRYB[52][18] ), .S(\SUMB[52][18] ) );
  FA_X1 S4_19 ( .A(\ab[52][19] ), .B(\CARRYB[51][19] ), .CI(\SUMB[51][20] ), 
        .CO(\CARRYB[52][19] ), .S(\SUMB[52][19] ) );
  FA_X1 S4_20 ( .A(\ab[52][20] ), .B(\CARRYB[51][20] ), .CI(\SUMB[51][21] ), 
        .CO(\CARRYB[52][20] ), .S(\SUMB[52][20] ) );
  FA_X1 S4_21 ( .A(\ab[52][21] ), .B(\CARRYB[51][21] ), .CI(\SUMB[51][22] ), 
        .CO(\CARRYB[52][21] ), .S(\SUMB[52][21] ) );
  FA_X1 S4_22 ( .A(\ab[52][22] ), .B(\CARRYB[51][22] ), .CI(\SUMB[51][23] ), 
        .CO(\CARRYB[52][22] ), .S(\SUMB[52][22] ) );
  FA_X1 S4_23 ( .A(\ab[52][23] ), .B(\CARRYB[51][23] ), .CI(\SUMB[51][24] ), 
        .CO(\CARRYB[52][23] ), .S(\SUMB[52][23] ) );
  FA_X1 S4_24 ( .A(\ab[52][24] ), .B(\CARRYB[51][24] ), .CI(\SUMB[51][25] ), 
        .CO(\CARRYB[52][24] ), .S(\SUMB[52][24] ) );
  FA_X1 S4_25 ( .A(\ab[52][25] ), .B(\CARRYB[51][25] ), .CI(\SUMB[51][26] ), 
        .CO(\CARRYB[52][25] ), .S(\SUMB[52][25] ) );
  FA_X1 S4_26 ( .A(\ab[52][26] ), .B(\CARRYB[51][26] ), .CI(\SUMB[51][27] ), 
        .CO(\CARRYB[52][26] ), .S(\SUMB[52][26] ) );
  FA_X1 S4_27 ( .A(\ab[52][27] ), .B(\CARRYB[51][27] ), .CI(\SUMB[51][28] ), 
        .CO(\CARRYB[52][27] ), .S(\SUMB[52][27] ) );
  FA_X1 S4_28 ( .A(\ab[52][28] ), .B(\CARRYB[51][28] ), .CI(\SUMB[51][29] ), 
        .CO(\CARRYB[52][28] ), .S(\SUMB[52][28] ) );
  FA_X1 S4_29 ( .A(\ab[52][29] ), .B(\CARRYB[51][29] ), .CI(\SUMB[51][30] ), 
        .CO(\CARRYB[52][29] ), .S(\SUMB[52][29] ) );
  FA_X1 S4_30 ( .A(\ab[52][30] ), .B(\CARRYB[51][30] ), .CI(\SUMB[51][31] ), 
        .CO(\CARRYB[52][30] ), .S(\SUMB[52][30] ) );
  FA_X1 S4_31 ( .A(\ab[52][31] ), .B(\CARRYB[51][31] ), .CI(\SUMB[51][32] ), 
        .CO(\CARRYB[52][31] ), .S(\SUMB[52][31] ) );
  FA_X1 S4_32 ( .A(\ab[52][32] ), .B(\CARRYB[51][32] ), .CI(\SUMB[51][33] ), 
        .CO(\CARRYB[52][32] ), .S(\SUMB[52][32] ) );
  FA_X1 S4_33 ( .A(\ab[52][33] ), .B(\CARRYB[51][33] ), .CI(\SUMB[51][34] ), 
        .CO(\CARRYB[52][33] ), .S(\SUMB[52][33] ) );
  FA_X1 S4_34 ( .A(\ab[52][34] ), .B(\CARRYB[51][34] ), .CI(\SUMB[51][35] ), 
        .CO(\CARRYB[52][34] ), .S(\SUMB[52][34] ) );
  FA_X1 S4_35 ( .A(\ab[52][35] ), .B(\CARRYB[51][35] ), .CI(\SUMB[51][36] ), 
        .CO(\CARRYB[52][35] ), .S(\SUMB[52][35] ) );
  FA_X1 S4_36 ( .A(\ab[52][36] ), .B(\CARRYB[51][36] ), .CI(\SUMB[51][37] ), 
        .CO(\CARRYB[52][36] ), .S(\SUMB[52][36] ) );
  FA_X1 S4_37 ( .A(\ab[52][37] ), .B(\CARRYB[51][37] ), .CI(\SUMB[51][38] ), 
        .CO(\CARRYB[52][37] ), .S(\SUMB[52][37] ) );
  FA_X1 S4_38 ( .A(\ab[52][38] ), .B(\CARRYB[51][38] ), .CI(\SUMB[51][39] ), 
        .CO(\CARRYB[52][38] ), .S(\SUMB[52][38] ) );
  FA_X1 S4_39 ( .A(\ab[52][39] ), .B(\CARRYB[51][39] ), .CI(\SUMB[51][40] ), 
        .CO(\CARRYB[52][39] ), .S(\SUMB[52][39] ) );
  FA_X1 S4_40 ( .A(\ab[52][40] ), .B(\CARRYB[51][40] ), .CI(\SUMB[51][41] ), 
        .CO(\CARRYB[52][40] ), .S(\SUMB[52][40] ) );
  FA_X1 S4_41 ( .A(\ab[52][41] ), .B(\CARRYB[51][41] ), .CI(\SUMB[51][42] ), 
        .CO(\CARRYB[52][41] ), .S(\SUMB[52][41] ) );
  FA_X1 S4_42 ( .A(\ab[52][42] ), .B(\CARRYB[51][42] ), .CI(\SUMB[51][43] ), 
        .CO(\CARRYB[52][42] ), .S(\SUMB[52][42] ) );
  FA_X1 S4_43 ( .A(\ab[52][43] ), .B(\CARRYB[51][43] ), .CI(\SUMB[51][44] ), 
        .CO(\CARRYB[52][43] ), .S(\SUMB[52][43] ) );
  FA_X1 S4_44 ( .A(\ab[52][44] ), .B(\CARRYB[51][44] ), .CI(\SUMB[51][45] ), 
        .CO(\CARRYB[52][44] ), .S(\SUMB[52][44] ) );
  FA_X1 S4_45 ( .A(\ab[52][45] ), .B(\CARRYB[51][45] ), .CI(\SUMB[51][46] ), 
        .CO(\CARRYB[52][45] ), .S(\SUMB[52][45] ) );
  FA_X1 S4_46 ( .A(\ab[52][46] ), .B(\CARRYB[51][46] ), .CI(\SUMB[51][47] ), 
        .CO(\CARRYB[52][46] ), .S(\SUMB[52][46] ) );
  FA_X1 S4_47 ( .A(\ab[52][47] ), .B(\CARRYB[51][47] ), .CI(\SUMB[51][48] ), 
        .CO(\CARRYB[52][47] ), .S(\SUMB[52][47] ) );
  FA_X1 S4_48 ( .A(\ab[52][48] ), .B(\CARRYB[51][48] ), .CI(\SUMB[51][49] ), 
        .CO(\CARRYB[52][48] ), .S(\SUMB[52][48] ) );
  FA_X1 S4_49 ( .A(\ab[52][49] ), .B(\CARRYB[51][49] ), .CI(\SUMB[51][50] ), 
        .CO(\CARRYB[52][49] ), .S(\SUMB[52][49] ) );
  FA_X1 S4_50 ( .A(\ab[52][50] ), .B(\CARRYB[51][50] ), .CI(\SUMB[51][51] ), 
        .CO(\CARRYB[52][50] ), .S(\SUMB[52][50] ) );
  FA_X1 S5_51 ( .A(\ab[52][51] ), .B(\CARRYB[51][51] ), .CI(\ab[51][52] ), 
        .CO(\CARRYB[52][51] ), .S(\SUMB[52][51] ) );
  FA_X1 S1_51_0 ( .A(\ab[51][0] ), .B(\CARRYB[50][0] ), .CI(\SUMB[50][1] ), 
        .CO(\CARRYB[51][0] ), .S(CLA_SUM[51]) );
  FA_X1 S2_51_1 ( .A(\ab[51][1] ), .B(\CARRYB[50][1] ), .CI(\SUMB[50][2] ), 
        .CO(\CARRYB[51][1] ), .S(\SUMB[51][1] ) );
  FA_X1 S2_51_2 ( .A(\ab[51][2] ), .B(\CARRYB[50][2] ), .CI(\SUMB[50][3] ), 
        .CO(\CARRYB[51][2] ), .S(\SUMB[51][2] ) );
  FA_X1 S2_51_3 ( .A(\ab[51][3] ), .B(\CARRYB[50][3] ), .CI(\SUMB[50][4] ), 
        .CO(\CARRYB[51][3] ), .S(\SUMB[51][3] ) );
  FA_X1 S2_51_4 ( .A(\ab[51][4] ), .B(\CARRYB[50][4] ), .CI(\SUMB[50][5] ), 
        .CO(\CARRYB[51][4] ), .S(\SUMB[51][4] ) );
  FA_X1 S2_51_5 ( .A(\ab[51][5] ), .B(\CARRYB[50][5] ), .CI(\SUMB[50][6] ), 
        .CO(\CARRYB[51][5] ), .S(\SUMB[51][5] ) );
  FA_X1 S2_51_6 ( .A(\ab[51][6] ), .B(\CARRYB[50][6] ), .CI(\SUMB[50][7] ), 
        .CO(\CARRYB[51][6] ), .S(\SUMB[51][6] ) );
  FA_X1 S2_51_7 ( .A(\ab[51][7] ), .B(\CARRYB[50][7] ), .CI(\SUMB[50][8] ), 
        .CO(\CARRYB[51][7] ), .S(\SUMB[51][7] ) );
  FA_X1 S2_51_8 ( .A(\ab[51][8] ), .B(\CARRYB[50][8] ), .CI(\SUMB[50][9] ), 
        .CO(\CARRYB[51][8] ), .S(\SUMB[51][8] ) );
  FA_X1 S2_51_9 ( .A(\ab[51][9] ), .B(\CARRYB[50][9] ), .CI(\SUMB[50][10] ), 
        .CO(\CARRYB[51][9] ), .S(\SUMB[51][9] ) );
  FA_X1 S2_51_10 ( .A(\ab[51][10] ), .B(\CARRYB[50][10] ), .CI(\SUMB[50][11] ), 
        .CO(\CARRYB[51][10] ), .S(\SUMB[51][10] ) );
  FA_X1 S2_51_11 ( .A(\ab[51][11] ), .B(\CARRYB[50][11] ), .CI(\SUMB[50][12] ), 
        .CO(\CARRYB[51][11] ), .S(\SUMB[51][11] ) );
  FA_X1 S2_51_12 ( .A(\ab[51][12] ), .B(\CARRYB[50][12] ), .CI(\SUMB[50][13] ), 
        .CO(\CARRYB[51][12] ), .S(\SUMB[51][12] ) );
  FA_X1 S2_51_13 ( .A(\ab[51][13] ), .B(\CARRYB[50][13] ), .CI(\SUMB[50][14] ), 
        .CO(\CARRYB[51][13] ), .S(\SUMB[51][13] ) );
  FA_X1 S2_51_14 ( .A(\ab[51][14] ), .B(\CARRYB[50][14] ), .CI(\SUMB[50][15] ), 
        .CO(\CARRYB[51][14] ), .S(\SUMB[51][14] ) );
  FA_X1 S2_51_15 ( .A(\ab[51][15] ), .B(\CARRYB[50][15] ), .CI(\SUMB[50][16] ), 
        .CO(\CARRYB[51][15] ), .S(\SUMB[51][15] ) );
  FA_X1 S2_51_16 ( .A(\ab[51][16] ), .B(\CARRYB[50][16] ), .CI(\SUMB[50][17] ), 
        .CO(\CARRYB[51][16] ), .S(\SUMB[51][16] ) );
  FA_X1 S2_51_17 ( .A(\ab[51][17] ), .B(\CARRYB[50][17] ), .CI(\SUMB[50][18] ), 
        .CO(\CARRYB[51][17] ), .S(\SUMB[51][17] ) );
  FA_X1 S2_51_18 ( .A(\ab[51][18] ), .B(\CARRYB[50][18] ), .CI(\SUMB[50][19] ), 
        .CO(\CARRYB[51][18] ), .S(\SUMB[51][18] ) );
  FA_X1 S2_51_19 ( .A(\ab[51][19] ), .B(\CARRYB[50][19] ), .CI(\SUMB[50][20] ), 
        .CO(\CARRYB[51][19] ), .S(\SUMB[51][19] ) );
  FA_X1 S2_51_20 ( .A(\ab[51][20] ), .B(\CARRYB[50][20] ), .CI(\SUMB[50][21] ), 
        .CO(\CARRYB[51][20] ), .S(\SUMB[51][20] ) );
  FA_X1 S2_51_21 ( .A(\ab[51][21] ), .B(\CARRYB[50][21] ), .CI(\SUMB[50][22] ), 
        .CO(\CARRYB[51][21] ), .S(\SUMB[51][21] ) );
  FA_X1 S2_51_22 ( .A(\ab[51][22] ), .B(\CARRYB[50][22] ), .CI(\SUMB[50][23] ), 
        .CO(\CARRYB[51][22] ), .S(\SUMB[51][22] ) );
  FA_X1 S2_51_23 ( .A(\ab[51][23] ), .B(\CARRYB[50][23] ), .CI(\SUMB[50][24] ), 
        .CO(\CARRYB[51][23] ), .S(\SUMB[51][23] ) );
  FA_X1 S2_51_24 ( .A(\ab[51][24] ), .B(\CARRYB[50][24] ), .CI(\SUMB[50][25] ), 
        .CO(\CARRYB[51][24] ), .S(\SUMB[51][24] ) );
  FA_X1 S2_51_25 ( .A(\ab[51][25] ), .B(\CARRYB[50][25] ), .CI(\SUMB[50][26] ), 
        .CO(\CARRYB[51][25] ), .S(\SUMB[51][25] ) );
  FA_X1 S2_51_26 ( .A(\ab[51][26] ), .B(\CARRYB[50][26] ), .CI(\SUMB[50][27] ), 
        .CO(\CARRYB[51][26] ), .S(\SUMB[51][26] ) );
  FA_X1 S2_51_27 ( .A(\ab[51][27] ), .B(\CARRYB[50][27] ), .CI(\SUMB[50][28] ), 
        .CO(\CARRYB[51][27] ), .S(\SUMB[51][27] ) );
  FA_X1 S2_51_28 ( .A(\ab[51][28] ), .B(\CARRYB[50][28] ), .CI(\SUMB[50][29] ), 
        .CO(\CARRYB[51][28] ), .S(\SUMB[51][28] ) );
  FA_X1 S2_51_29 ( .A(\ab[51][29] ), .B(\CARRYB[50][29] ), .CI(\SUMB[50][30] ), 
        .CO(\CARRYB[51][29] ), .S(\SUMB[51][29] ) );
  FA_X1 S2_51_30 ( .A(\ab[51][30] ), .B(\CARRYB[50][30] ), .CI(\SUMB[50][31] ), 
        .CO(\CARRYB[51][30] ), .S(\SUMB[51][30] ) );
  FA_X1 S2_51_31 ( .A(\ab[51][31] ), .B(\CARRYB[50][31] ), .CI(\SUMB[50][32] ), 
        .CO(\CARRYB[51][31] ), .S(\SUMB[51][31] ) );
  FA_X1 S2_51_32 ( .A(\ab[51][32] ), .B(\CARRYB[50][32] ), .CI(\SUMB[50][33] ), 
        .CO(\CARRYB[51][32] ), .S(\SUMB[51][32] ) );
  FA_X1 S2_51_33 ( .A(\ab[51][33] ), .B(\CARRYB[50][33] ), .CI(\SUMB[50][34] ), 
        .CO(\CARRYB[51][33] ), .S(\SUMB[51][33] ) );
  FA_X1 S2_51_34 ( .A(\ab[51][34] ), .B(\CARRYB[50][34] ), .CI(\SUMB[50][35] ), 
        .CO(\CARRYB[51][34] ), .S(\SUMB[51][34] ) );
  FA_X1 S2_51_35 ( .A(\ab[51][35] ), .B(\CARRYB[50][35] ), .CI(\SUMB[50][36] ), 
        .CO(\CARRYB[51][35] ), .S(\SUMB[51][35] ) );
  FA_X1 S2_51_36 ( .A(\ab[51][36] ), .B(\CARRYB[50][36] ), .CI(\SUMB[50][37] ), 
        .CO(\CARRYB[51][36] ), .S(\SUMB[51][36] ) );
  FA_X1 S2_51_37 ( .A(\ab[51][37] ), .B(\CARRYB[50][37] ), .CI(\SUMB[50][38] ), 
        .CO(\CARRYB[51][37] ), .S(\SUMB[51][37] ) );
  FA_X1 S2_51_38 ( .A(\ab[51][38] ), .B(\CARRYB[50][38] ), .CI(\SUMB[50][39] ), 
        .CO(\CARRYB[51][38] ), .S(\SUMB[51][38] ) );
  FA_X1 S2_51_39 ( .A(\ab[51][39] ), .B(\CARRYB[50][39] ), .CI(\SUMB[50][40] ), 
        .CO(\CARRYB[51][39] ), .S(\SUMB[51][39] ) );
  FA_X1 S2_51_40 ( .A(\ab[51][40] ), .B(\CARRYB[50][40] ), .CI(\SUMB[50][41] ), 
        .CO(\CARRYB[51][40] ), .S(\SUMB[51][40] ) );
  FA_X1 S2_51_41 ( .A(\ab[51][41] ), .B(\CARRYB[50][41] ), .CI(\SUMB[50][42] ), 
        .CO(\CARRYB[51][41] ), .S(\SUMB[51][41] ) );
  FA_X1 S2_51_42 ( .A(\ab[51][42] ), .B(\CARRYB[50][42] ), .CI(\SUMB[50][43] ), 
        .CO(\CARRYB[51][42] ), .S(\SUMB[51][42] ) );
  FA_X1 S2_51_43 ( .A(\ab[51][43] ), .B(\CARRYB[50][43] ), .CI(\SUMB[50][44] ), 
        .CO(\CARRYB[51][43] ), .S(\SUMB[51][43] ) );
  FA_X1 S2_51_44 ( .A(\ab[51][44] ), .B(\CARRYB[50][44] ), .CI(\SUMB[50][45] ), 
        .CO(\CARRYB[51][44] ), .S(\SUMB[51][44] ) );
  FA_X1 S2_51_45 ( .A(\ab[51][45] ), .B(\CARRYB[50][45] ), .CI(\SUMB[50][46] ), 
        .CO(\CARRYB[51][45] ), .S(\SUMB[51][45] ) );
  FA_X1 S2_51_46 ( .A(\ab[51][46] ), .B(\CARRYB[50][46] ), .CI(\SUMB[50][47] ), 
        .CO(\CARRYB[51][46] ), .S(\SUMB[51][46] ) );
  FA_X1 S2_51_47 ( .A(\ab[51][47] ), .B(\CARRYB[50][47] ), .CI(\SUMB[50][48] ), 
        .CO(\CARRYB[51][47] ), .S(\SUMB[51][47] ) );
  FA_X1 S2_51_48 ( .A(\ab[51][48] ), .B(\CARRYB[50][48] ), .CI(\SUMB[50][49] ), 
        .CO(\CARRYB[51][48] ), .S(\SUMB[51][48] ) );
  FA_X1 S2_51_49 ( .A(\ab[51][49] ), .B(\CARRYB[50][49] ), .CI(\SUMB[50][50] ), 
        .CO(\CARRYB[51][49] ), .S(\SUMB[51][49] ) );
  FA_X1 S2_51_50 ( .A(\ab[51][50] ), .B(\CARRYB[50][50] ), .CI(\SUMB[50][51] ), 
        .CO(\CARRYB[51][50] ), .S(\SUMB[51][50] ) );
  FA_X1 S3_51_51 ( .A(\ab[51][51] ), .B(\CARRYB[50][51] ), .CI(\ab[50][52] ), 
        .CO(\CARRYB[51][51] ), .S(\SUMB[51][51] ) );
  FA_X1 S1_50_0 ( .A(\ab[50][0] ), .B(\CARRYB[49][0] ), .CI(\SUMB[49][1] ), 
        .CO(\CARRYB[50][0] ), .S(CLA_SUM[50]) );
  FA_X1 S2_50_1 ( .A(\ab[50][1] ), .B(\CARRYB[49][1] ), .CI(\SUMB[49][2] ), 
        .CO(\CARRYB[50][1] ), .S(\SUMB[50][1] ) );
  FA_X1 S2_50_2 ( .A(\ab[50][2] ), .B(\CARRYB[49][2] ), .CI(\SUMB[49][3] ), 
        .CO(\CARRYB[50][2] ), .S(\SUMB[50][2] ) );
  FA_X1 S2_50_3 ( .A(\ab[50][3] ), .B(\CARRYB[49][3] ), .CI(\SUMB[49][4] ), 
        .CO(\CARRYB[50][3] ), .S(\SUMB[50][3] ) );
  FA_X1 S2_50_4 ( .A(\ab[50][4] ), .B(\CARRYB[49][4] ), .CI(\SUMB[49][5] ), 
        .CO(\CARRYB[50][4] ), .S(\SUMB[50][4] ) );
  FA_X1 S2_50_5 ( .A(\ab[50][5] ), .B(\CARRYB[49][5] ), .CI(\SUMB[49][6] ), 
        .CO(\CARRYB[50][5] ), .S(\SUMB[50][5] ) );
  FA_X1 S2_50_6 ( .A(\ab[50][6] ), .B(\CARRYB[49][6] ), .CI(\SUMB[49][7] ), 
        .CO(\CARRYB[50][6] ), .S(\SUMB[50][6] ) );
  FA_X1 S2_50_7 ( .A(\ab[50][7] ), .B(\CARRYB[49][7] ), .CI(\SUMB[49][8] ), 
        .CO(\CARRYB[50][7] ), .S(\SUMB[50][7] ) );
  FA_X1 S2_50_8 ( .A(\ab[50][8] ), .B(\CARRYB[49][8] ), .CI(\SUMB[49][9] ), 
        .CO(\CARRYB[50][8] ), .S(\SUMB[50][8] ) );
  FA_X1 S2_50_9 ( .A(\ab[50][9] ), .B(\CARRYB[49][9] ), .CI(\SUMB[49][10] ), 
        .CO(\CARRYB[50][9] ), .S(\SUMB[50][9] ) );
  FA_X1 S2_50_10 ( .A(\ab[50][10] ), .B(\CARRYB[49][10] ), .CI(\SUMB[49][11] ), 
        .CO(\CARRYB[50][10] ), .S(\SUMB[50][10] ) );
  FA_X1 S2_50_11 ( .A(\ab[50][11] ), .B(\CARRYB[49][11] ), .CI(\SUMB[49][12] ), 
        .CO(\CARRYB[50][11] ), .S(\SUMB[50][11] ) );
  FA_X1 S2_50_12 ( .A(\ab[50][12] ), .B(\CARRYB[49][12] ), .CI(\SUMB[49][13] ), 
        .CO(\CARRYB[50][12] ), .S(\SUMB[50][12] ) );
  FA_X1 S2_50_13 ( .A(\ab[50][13] ), .B(\CARRYB[49][13] ), .CI(\SUMB[49][14] ), 
        .CO(\CARRYB[50][13] ), .S(\SUMB[50][13] ) );
  FA_X1 S2_50_14 ( .A(\ab[50][14] ), .B(\CARRYB[49][14] ), .CI(\SUMB[49][15] ), 
        .CO(\CARRYB[50][14] ), .S(\SUMB[50][14] ) );
  FA_X1 S2_50_15 ( .A(\ab[50][15] ), .B(\CARRYB[49][15] ), .CI(\SUMB[49][16] ), 
        .CO(\CARRYB[50][15] ), .S(\SUMB[50][15] ) );
  FA_X1 S2_50_16 ( .A(\ab[50][16] ), .B(\CARRYB[49][16] ), .CI(\SUMB[49][17] ), 
        .CO(\CARRYB[50][16] ), .S(\SUMB[50][16] ) );
  FA_X1 S2_50_17 ( .A(\ab[50][17] ), .B(\CARRYB[49][17] ), .CI(\SUMB[49][18] ), 
        .CO(\CARRYB[50][17] ), .S(\SUMB[50][17] ) );
  FA_X1 S2_50_18 ( .A(\ab[50][18] ), .B(\CARRYB[49][18] ), .CI(\SUMB[49][19] ), 
        .CO(\CARRYB[50][18] ), .S(\SUMB[50][18] ) );
  FA_X1 S2_50_19 ( .A(\ab[50][19] ), .B(\CARRYB[49][19] ), .CI(\SUMB[49][20] ), 
        .CO(\CARRYB[50][19] ), .S(\SUMB[50][19] ) );
  FA_X1 S2_50_20 ( .A(\ab[50][20] ), .B(\CARRYB[49][20] ), .CI(\SUMB[49][21] ), 
        .CO(\CARRYB[50][20] ), .S(\SUMB[50][20] ) );
  FA_X1 S2_50_21 ( .A(\ab[50][21] ), .B(\CARRYB[49][21] ), .CI(\SUMB[49][22] ), 
        .CO(\CARRYB[50][21] ), .S(\SUMB[50][21] ) );
  FA_X1 S2_50_22 ( .A(\ab[50][22] ), .B(\CARRYB[49][22] ), .CI(\SUMB[49][23] ), 
        .CO(\CARRYB[50][22] ), .S(\SUMB[50][22] ) );
  FA_X1 S2_50_23 ( .A(\ab[50][23] ), .B(\CARRYB[49][23] ), .CI(\SUMB[49][24] ), 
        .CO(\CARRYB[50][23] ), .S(\SUMB[50][23] ) );
  FA_X1 S2_50_24 ( .A(\ab[50][24] ), .B(\CARRYB[49][24] ), .CI(\SUMB[49][25] ), 
        .CO(\CARRYB[50][24] ), .S(\SUMB[50][24] ) );
  FA_X1 S2_50_25 ( .A(\ab[50][25] ), .B(\CARRYB[49][25] ), .CI(\SUMB[49][26] ), 
        .CO(\CARRYB[50][25] ), .S(\SUMB[50][25] ) );
  FA_X1 S2_50_26 ( .A(\ab[50][26] ), .B(\CARRYB[49][26] ), .CI(\SUMB[49][27] ), 
        .CO(\CARRYB[50][26] ), .S(\SUMB[50][26] ) );
  FA_X1 S2_50_27 ( .A(\ab[50][27] ), .B(\CARRYB[49][27] ), .CI(\SUMB[49][28] ), 
        .CO(\CARRYB[50][27] ), .S(\SUMB[50][27] ) );
  FA_X1 S2_50_28 ( .A(\ab[50][28] ), .B(\CARRYB[49][28] ), .CI(\SUMB[49][29] ), 
        .CO(\CARRYB[50][28] ), .S(\SUMB[50][28] ) );
  FA_X1 S2_50_29 ( .A(\ab[50][29] ), .B(\CARRYB[49][29] ), .CI(\SUMB[49][30] ), 
        .CO(\CARRYB[50][29] ), .S(\SUMB[50][29] ) );
  FA_X1 S2_50_30 ( .A(\ab[50][30] ), .B(\CARRYB[49][30] ), .CI(\SUMB[49][31] ), 
        .CO(\CARRYB[50][30] ), .S(\SUMB[50][30] ) );
  FA_X1 S2_50_31 ( .A(\ab[50][31] ), .B(\CARRYB[49][31] ), .CI(\SUMB[49][32] ), 
        .CO(\CARRYB[50][31] ), .S(\SUMB[50][31] ) );
  FA_X1 S2_50_32 ( .A(\ab[50][32] ), .B(\CARRYB[49][32] ), .CI(\SUMB[49][33] ), 
        .CO(\CARRYB[50][32] ), .S(\SUMB[50][32] ) );
  FA_X1 S2_50_33 ( .A(\ab[50][33] ), .B(\CARRYB[49][33] ), .CI(\SUMB[49][34] ), 
        .CO(\CARRYB[50][33] ), .S(\SUMB[50][33] ) );
  FA_X1 S2_50_34 ( .A(\ab[50][34] ), .B(\CARRYB[49][34] ), .CI(\SUMB[49][35] ), 
        .CO(\CARRYB[50][34] ), .S(\SUMB[50][34] ) );
  FA_X1 S2_50_35 ( .A(\ab[50][35] ), .B(\CARRYB[49][35] ), .CI(\SUMB[49][36] ), 
        .CO(\CARRYB[50][35] ), .S(\SUMB[50][35] ) );
  FA_X1 S2_50_36 ( .A(\ab[50][36] ), .B(\CARRYB[49][36] ), .CI(\SUMB[49][37] ), 
        .CO(\CARRYB[50][36] ), .S(\SUMB[50][36] ) );
  FA_X1 S2_50_37 ( .A(\ab[50][37] ), .B(\CARRYB[49][37] ), .CI(\SUMB[49][38] ), 
        .CO(\CARRYB[50][37] ), .S(\SUMB[50][37] ) );
  FA_X1 S2_50_38 ( .A(\ab[50][38] ), .B(\CARRYB[49][38] ), .CI(\SUMB[49][39] ), 
        .CO(\CARRYB[50][38] ), .S(\SUMB[50][38] ) );
  FA_X1 S2_50_39 ( .A(\ab[50][39] ), .B(\CARRYB[49][39] ), .CI(\SUMB[49][40] ), 
        .CO(\CARRYB[50][39] ), .S(\SUMB[50][39] ) );
  FA_X1 S2_50_40 ( .A(\ab[50][40] ), .B(\CARRYB[49][40] ), .CI(\SUMB[49][41] ), 
        .CO(\CARRYB[50][40] ), .S(\SUMB[50][40] ) );
  FA_X1 S2_50_41 ( .A(\ab[50][41] ), .B(\CARRYB[49][41] ), .CI(\SUMB[49][42] ), 
        .CO(\CARRYB[50][41] ), .S(\SUMB[50][41] ) );
  FA_X1 S2_50_42 ( .A(\ab[50][42] ), .B(\CARRYB[49][42] ), .CI(\SUMB[49][43] ), 
        .CO(\CARRYB[50][42] ), .S(\SUMB[50][42] ) );
  FA_X1 S2_50_43 ( .A(\ab[50][43] ), .B(\CARRYB[49][43] ), .CI(\SUMB[49][44] ), 
        .CO(\CARRYB[50][43] ), .S(\SUMB[50][43] ) );
  FA_X1 S2_50_44 ( .A(\ab[50][44] ), .B(\CARRYB[49][44] ), .CI(\SUMB[49][45] ), 
        .CO(\CARRYB[50][44] ), .S(\SUMB[50][44] ) );
  FA_X1 S2_50_45 ( .A(\ab[50][45] ), .B(\CARRYB[49][45] ), .CI(\SUMB[49][46] ), 
        .CO(\CARRYB[50][45] ), .S(\SUMB[50][45] ) );
  FA_X1 S2_50_46 ( .A(\ab[50][46] ), .B(\CARRYB[49][46] ), .CI(\SUMB[49][47] ), 
        .CO(\CARRYB[50][46] ), .S(\SUMB[50][46] ) );
  FA_X1 S2_50_47 ( .A(\ab[50][47] ), .B(\CARRYB[49][47] ), .CI(\SUMB[49][48] ), 
        .CO(\CARRYB[50][47] ), .S(\SUMB[50][47] ) );
  FA_X1 S2_50_48 ( .A(\ab[50][48] ), .B(\CARRYB[49][48] ), .CI(\SUMB[49][49] ), 
        .CO(\CARRYB[50][48] ), .S(\SUMB[50][48] ) );
  FA_X1 S2_50_49 ( .A(\ab[50][49] ), .B(\CARRYB[49][49] ), .CI(\SUMB[49][50] ), 
        .CO(\CARRYB[50][49] ), .S(\SUMB[50][49] ) );
  FA_X1 S2_50_50 ( .A(\ab[50][50] ), .B(\CARRYB[49][50] ), .CI(\SUMB[49][51] ), 
        .CO(\CARRYB[50][50] ), .S(\SUMB[50][50] ) );
  FA_X1 S3_50_51 ( .A(\ab[50][51] ), .B(\CARRYB[49][51] ), .CI(\ab[49][52] ), 
        .CO(\CARRYB[50][51] ), .S(\SUMB[50][51] ) );
  FA_X1 S1_49_0 ( .A(\ab[49][0] ), .B(\CARRYB[48][0] ), .CI(\SUMB[48][1] ), 
        .CO(\CARRYB[49][0] ), .S(CLA_SUM[49]) );
  FA_X1 S2_49_1 ( .A(\ab[49][1] ), .B(\CARRYB[48][1] ), .CI(\SUMB[48][2] ), 
        .CO(\CARRYB[49][1] ), .S(\SUMB[49][1] ) );
  FA_X1 S2_49_2 ( .A(\ab[49][2] ), .B(\CARRYB[48][2] ), .CI(\SUMB[48][3] ), 
        .CO(\CARRYB[49][2] ), .S(\SUMB[49][2] ) );
  FA_X1 S2_49_3 ( .A(\ab[49][3] ), .B(\CARRYB[48][3] ), .CI(\SUMB[48][4] ), 
        .CO(\CARRYB[49][3] ), .S(\SUMB[49][3] ) );
  FA_X1 S2_49_4 ( .A(\ab[49][4] ), .B(\CARRYB[48][4] ), .CI(\SUMB[48][5] ), 
        .CO(\CARRYB[49][4] ), .S(\SUMB[49][4] ) );
  FA_X1 S2_49_5 ( .A(\ab[49][5] ), .B(\CARRYB[48][5] ), .CI(\SUMB[48][6] ), 
        .CO(\CARRYB[49][5] ), .S(\SUMB[49][5] ) );
  FA_X1 S2_49_6 ( .A(\ab[49][6] ), .B(\CARRYB[48][6] ), .CI(\SUMB[48][7] ), 
        .CO(\CARRYB[49][6] ), .S(\SUMB[49][6] ) );
  FA_X1 S2_49_7 ( .A(\ab[49][7] ), .B(\CARRYB[48][7] ), .CI(\SUMB[48][8] ), 
        .CO(\CARRYB[49][7] ), .S(\SUMB[49][7] ) );
  FA_X1 S2_49_8 ( .A(\ab[49][8] ), .B(\CARRYB[48][8] ), .CI(\SUMB[48][9] ), 
        .CO(\CARRYB[49][8] ), .S(\SUMB[49][8] ) );
  FA_X1 S2_49_9 ( .A(\ab[49][9] ), .B(\CARRYB[48][9] ), .CI(\SUMB[48][10] ), 
        .CO(\CARRYB[49][9] ), .S(\SUMB[49][9] ) );
  FA_X1 S2_49_10 ( .A(\ab[49][10] ), .B(\CARRYB[48][10] ), .CI(\SUMB[48][11] ), 
        .CO(\CARRYB[49][10] ), .S(\SUMB[49][10] ) );
  FA_X1 S2_49_11 ( .A(\ab[49][11] ), .B(\CARRYB[48][11] ), .CI(\SUMB[48][12] ), 
        .CO(\CARRYB[49][11] ), .S(\SUMB[49][11] ) );
  FA_X1 S2_49_12 ( .A(\ab[49][12] ), .B(\CARRYB[48][12] ), .CI(\SUMB[48][13] ), 
        .CO(\CARRYB[49][12] ), .S(\SUMB[49][12] ) );
  FA_X1 S2_49_13 ( .A(\ab[49][13] ), .B(\CARRYB[48][13] ), .CI(\SUMB[48][14] ), 
        .CO(\CARRYB[49][13] ), .S(\SUMB[49][13] ) );
  FA_X1 S2_49_14 ( .A(\ab[49][14] ), .B(\CARRYB[48][14] ), .CI(\SUMB[48][15] ), 
        .CO(\CARRYB[49][14] ), .S(\SUMB[49][14] ) );
  FA_X1 S2_49_15 ( .A(\ab[49][15] ), .B(\CARRYB[48][15] ), .CI(\SUMB[48][16] ), 
        .CO(\CARRYB[49][15] ), .S(\SUMB[49][15] ) );
  FA_X1 S2_49_16 ( .A(\ab[49][16] ), .B(\CARRYB[48][16] ), .CI(\SUMB[48][17] ), 
        .CO(\CARRYB[49][16] ), .S(\SUMB[49][16] ) );
  FA_X1 S2_49_17 ( .A(\ab[49][17] ), .B(\CARRYB[48][17] ), .CI(\SUMB[48][18] ), 
        .CO(\CARRYB[49][17] ), .S(\SUMB[49][17] ) );
  FA_X1 S2_49_18 ( .A(\ab[49][18] ), .B(\CARRYB[48][18] ), .CI(\SUMB[48][19] ), 
        .CO(\CARRYB[49][18] ), .S(\SUMB[49][18] ) );
  FA_X1 S2_49_19 ( .A(\ab[49][19] ), .B(\CARRYB[48][19] ), .CI(\SUMB[48][20] ), 
        .CO(\CARRYB[49][19] ), .S(\SUMB[49][19] ) );
  FA_X1 S2_49_20 ( .A(\ab[49][20] ), .B(\CARRYB[48][20] ), .CI(\SUMB[48][21] ), 
        .CO(\CARRYB[49][20] ), .S(\SUMB[49][20] ) );
  FA_X1 S2_49_21 ( .A(\ab[49][21] ), .B(\CARRYB[48][21] ), .CI(\SUMB[48][22] ), 
        .CO(\CARRYB[49][21] ), .S(\SUMB[49][21] ) );
  FA_X1 S2_49_22 ( .A(\ab[49][22] ), .B(\CARRYB[48][22] ), .CI(\SUMB[48][23] ), 
        .CO(\CARRYB[49][22] ), .S(\SUMB[49][22] ) );
  FA_X1 S2_49_23 ( .A(\ab[49][23] ), .B(\CARRYB[48][23] ), .CI(\SUMB[48][24] ), 
        .CO(\CARRYB[49][23] ), .S(\SUMB[49][23] ) );
  FA_X1 S2_49_24 ( .A(\ab[49][24] ), .B(\CARRYB[48][24] ), .CI(\SUMB[48][25] ), 
        .CO(\CARRYB[49][24] ), .S(\SUMB[49][24] ) );
  FA_X1 S2_49_25 ( .A(\ab[49][25] ), .B(\CARRYB[48][25] ), .CI(\SUMB[48][26] ), 
        .CO(\CARRYB[49][25] ), .S(\SUMB[49][25] ) );
  FA_X1 S2_49_26 ( .A(\ab[49][26] ), .B(\CARRYB[48][26] ), .CI(\SUMB[48][27] ), 
        .CO(\CARRYB[49][26] ), .S(\SUMB[49][26] ) );
  FA_X1 S2_49_27 ( .A(\ab[49][27] ), .B(\CARRYB[48][27] ), .CI(\SUMB[48][28] ), 
        .CO(\CARRYB[49][27] ), .S(\SUMB[49][27] ) );
  FA_X1 S2_49_28 ( .A(\ab[49][28] ), .B(\CARRYB[48][28] ), .CI(\SUMB[48][29] ), 
        .CO(\CARRYB[49][28] ), .S(\SUMB[49][28] ) );
  FA_X1 S2_49_29 ( .A(\ab[49][29] ), .B(\CARRYB[48][29] ), .CI(\SUMB[48][30] ), 
        .CO(\CARRYB[49][29] ), .S(\SUMB[49][29] ) );
  FA_X1 S2_49_30 ( .A(\ab[49][30] ), .B(\CARRYB[48][30] ), .CI(\SUMB[48][31] ), 
        .CO(\CARRYB[49][30] ), .S(\SUMB[49][30] ) );
  FA_X1 S2_49_31 ( .A(\ab[49][31] ), .B(\CARRYB[48][31] ), .CI(\SUMB[48][32] ), 
        .CO(\CARRYB[49][31] ), .S(\SUMB[49][31] ) );
  FA_X1 S2_49_32 ( .A(\ab[49][32] ), .B(\CARRYB[48][32] ), .CI(\SUMB[48][33] ), 
        .CO(\CARRYB[49][32] ), .S(\SUMB[49][32] ) );
  FA_X1 S2_49_33 ( .A(\ab[49][33] ), .B(\CARRYB[48][33] ), .CI(\SUMB[48][34] ), 
        .CO(\CARRYB[49][33] ), .S(\SUMB[49][33] ) );
  FA_X1 S2_49_34 ( .A(\ab[49][34] ), .B(\CARRYB[48][34] ), .CI(\SUMB[48][35] ), 
        .CO(\CARRYB[49][34] ), .S(\SUMB[49][34] ) );
  FA_X1 S2_49_35 ( .A(\ab[49][35] ), .B(\CARRYB[48][35] ), .CI(\SUMB[48][36] ), 
        .CO(\CARRYB[49][35] ), .S(\SUMB[49][35] ) );
  FA_X1 S2_49_36 ( .A(\ab[49][36] ), .B(\CARRYB[48][36] ), .CI(\SUMB[48][37] ), 
        .CO(\CARRYB[49][36] ), .S(\SUMB[49][36] ) );
  FA_X1 S2_49_37 ( .A(\ab[49][37] ), .B(\CARRYB[48][37] ), .CI(\SUMB[48][38] ), 
        .CO(\CARRYB[49][37] ), .S(\SUMB[49][37] ) );
  FA_X1 S2_49_38 ( .A(\ab[49][38] ), .B(\CARRYB[48][38] ), .CI(\SUMB[48][39] ), 
        .CO(\CARRYB[49][38] ), .S(\SUMB[49][38] ) );
  FA_X1 S2_49_39 ( .A(\ab[49][39] ), .B(\CARRYB[48][39] ), .CI(\SUMB[48][40] ), 
        .CO(\CARRYB[49][39] ), .S(\SUMB[49][39] ) );
  FA_X1 S2_49_40 ( .A(\ab[49][40] ), .B(\CARRYB[48][40] ), .CI(\SUMB[48][41] ), 
        .CO(\CARRYB[49][40] ), .S(\SUMB[49][40] ) );
  FA_X1 S2_49_41 ( .A(\ab[49][41] ), .B(\CARRYB[48][41] ), .CI(\SUMB[48][42] ), 
        .CO(\CARRYB[49][41] ), .S(\SUMB[49][41] ) );
  FA_X1 S2_49_42 ( .A(\ab[49][42] ), .B(\CARRYB[48][42] ), .CI(\SUMB[48][43] ), 
        .CO(\CARRYB[49][42] ), .S(\SUMB[49][42] ) );
  FA_X1 S2_49_43 ( .A(\ab[49][43] ), .B(\CARRYB[48][43] ), .CI(\SUMB[48][44] ), 
        .CO(\CARRYB[49][43] ), .S(\SUMB[49][43] ) );
  FA_X1 S2_49_44 ( .A(\ab[49][44] ), .B(\CARRYB[48][44] ), .CI(\SUMB[48][45] ), 
        .CO(\CARRYB[49][44] ), .S(\SUMB[49][44] ) );
  FA_X1 S2_49_45 ( .A(\ab[49][45] ), .B(\CARRYB[48][45] ), .CI(\SUMB[48][46] ), 
        .CO(\CARRYB[49][45] ), .S(\SUMB[49][45] ) );
  FA_X1 S2_49_46 ( .A(\ab[49][46] ), .B(\CARRYB[48][46] ), .CI(\SUMB[48][47] ), 
        .CO(\CARRYB[49][46] ), .S(\SUMB[49][46] ) );
  FA_X1 S2_49_47 ( .A(\ab[49][47] ), .B(\CARRYB[48][47] ), .CI(\SUMB[48][48] ), 
        .CO(\CARRYB[49][47] ), .S(\SUMB[49][47] ) );
  FA_X1 S2_49_48 ( .A(\ab[49][48] ), .B(\CARRYB[48][48] ), .CI(\SUMB[48][49] ), 
        .CO(\CARRYB[49][48] ), .S(\SUMB[49][48] ) );
  FA_X1 S2_49_49 ( .A(\ab[49][49] ), .B(\CARRYB[48][49] ), .CI(\SUMB[48][50] ), 
        .CO(\CARRYB[49][49] ), .S(\SUMB[49][49] ) );
  FA_X1 S2_49_50 ( .A(\ab[49][50] ), .B(\CARRYB[48][50] ), .CI(\SUMB[48][51] ), 
        .CO(\CARRYB[49][50] ), .S(\SUMB[49][50] ) );
  FA_X1 S3_49_51 ( .A(\ab[49][51] ), .B(\CARRYB[48][51] ), .CI(\ab[48][52] ), 
        .CO(\CARRYB[49][51] ), .S(\SUMB[49][51] ) );
  FA_X1 S1_48_0 ( .A(\ab[48][0] ), .B(\CARRYB[47][0] ), .CI(\SUMB[47][1] ), 
        .CO(\CARRYB[48][0] ), .S(CLA_SUM[48]) );
  FA_X1 S2_48_1 ( .A(\ab[48][1] ), .B(\CARRYB[47][1] ), .CI(\SUMB[47][2] ), 
        .CO(\CARRYB[48][1] ), .S(\SUMB[48][1] ) );
  FA_X1 S2_48_2 ( .A(\ab[48][2] ), .B(\CARRYB[47][2] ), .CI(\SUMB[47][3] ), 
        .CO(\CARRYB[48][2] ), .S(\SUMB[48][2] ) );
  FA_X1 S2_48_3 ( .A(\ab[48][3] ), .B(\CARRYB[47][3] ), .CI(\SUMB[47][4] ), 
        .CO(\CARRYB[48][3] ), .S(\SUMB[48][3] ) );
  FA_X1 S2_48_4 ( .A(\ab[48][4] ), .B(\CARRYB[47][4] ), .CI(\SUMB[47][5] ), 
        .CO(\CARRYB[48][4] ), .S(\SUMB[48][4] ) );
  FA_X1 S2_48_5 ( .A(\ab[48][5] ), .B(\CARRYB[47][5] ), .CI(\SUMB[47][6] ), 
        .CO(\CARRYB[48][5] ), .S(\SUMB[48][5] ) );
  FA_X1 S2_48_6 ( .A(\ab[48][6] ), .B(\CARRYB[47][6] ), .CI(\SUMB[47][7] ), 
        .CO(\CARRYB[48][6] ), .S(\SUMB[48][6] ) );
  FA_X1 S2_48_7 ( .A(\ab[48][7] ), .B(\CARRYB[47][7] ), .CI(\SUMB[47][8] ), 
        .CO(\CARRYB[48][7] ), .S(\SUMB[48][7] ) );
  FA_X1 S2_48_8 ( .A(\ab[48][8] ), .B(\CARRYB[47][8] ), .CI(\SUMB[47][9] ), 
        .CO(\CARRYB[48][8] ), .S(\SUMB[48][8] ) );
  FA_X1 S2_48_9 ( .A(\ab[48][9] ), .B(\CARRYB[47][9] ), .CI(\SUMB[47][10] ), 
        .CO(\CARRYB[48][9] ), .S(\SUMB[48][9] ) );
  FA_X1 S2_48_10 ( .A(\ab[48][10] ), .B(\CARRYB[47][10] ), .CI(\SUMB[47][11] ), 
        .CO(\CARRYB[48][10] ), .S(\SUMB[48][10] ) );
  FA_X1 S2_48_11 ( .A(\ab[48][11] ), .B(\CARRYB[47][11] ), .CI(\SUMB[47][12] ), 
        .CO(\CARRYB[48][11] ), .S(\SUMB[48][11] ) );
  FA_X1 S2_48_12 ( .A(\ab[48][12] ), .B(\CARRYB[47][12] ), .CI(\SUMB[47][13] ), 
        .CO(\CARRYB[48][12] ), .S(\SUMB[48][12] ) );
  FA_X1 S2_48_13 ( .A(\ab[48][13] ), .B(\CARRYB[47][13] ), .CI(\SUMB[47][14] ), 
        .CO(\CARRYB[48][13] ), .S(\SUMB[48][13] ) );
  FA_X1 S2_48_14 ( .A(\ab[48][14] ), .B(\CARRYB[47][14] ), .CI(\SUMB[47][15] ), 
        .CO(\CARRYB[48][14] ), .S(\SUMB[48][14] ) );
  FA_X1 S2_48_15 ( .A(\ab[48][15] ), .B(\CARRYB[47][15] ), .CI(\SUMB[47][16] ), 
        .CO(\CARRYB[48][15] ), .S(\SUMB[48][15] ) );
  FA_X1 S2_48_16 ( .A(\ab[48][16] ), .B(\CARRYB[47][16] ), .CI(\SUMB[47][17] ), 
        .CO(\CARRYB[48][16] ), .S(\SUMB[48][16] ) );
  FA_X1 S2_48_17 ( .A(\ab[48][17] ), .B(\CARRYB[47][17] ), .CI(\SUMB[47][18] ), 
        .CO(\CARRYB[48][17] ), .S(\SUMB[48][17] ) );
  FA_X1 S2_48_18 ( .A(\ab[48][18] ), .B(\CARRYB[47][18] ), .CI(\SUMB[47][19] ), 
        .CO(\CARRYB[48][18] ), .S(\SUMB[48][18] ) );
  FA_X1 S2_48_19 ( .A(\ab[48][19] ), .B(\CARRYB[47][19] ), .CI(\SUMB[47][20] ), 
        .CO(\CARRYB[48][19] ), .S(\SUMB[48][19] ) );
  FA_X1 S2_48_20 ( .A(\ab[48][20] ), .B(\CARRYB[47][20] ), .CI(\SUMB[47][21] ), 
        .CO(\CARRYB[48][20] ), .S(\SUMB[48][20] ) );
  FA_X1 S2_48_21 ( .A(\ab[48][21] ), .B(\CARRYB[47][21] ), .CI(\SUMB[47][22] ), 
        .CO(\CARRYB[48][21] ), .S(\SUMB[48][21] ) );
  FA_X1 S2_48_22 ( .A(\ab[48][22] ), .B(\CARRYB[47][22] ), .CI(\SUMB[47][23] ), 
        .CO(\CARRYB[48][22] ), .S(\SUMB[48][22] ) );
  FA_X1 S2_48_23 ( .A(\ab[48][23] ), .B(\CARRYB[47][23] ), .CI(\SUMB[47][24] ), 
        .CO(\CARRYB[48][23] ), .S(\SUMB[48][23] ) );
  FA_X1 S2_48_24 ( .A(\ab[48][24] ), .B(\CARRYB[47][24] ), .CI(\SUMB[47][25] ), 
        .CO(\CARRYB[48][24] ), .S(\SUMB[48][24] ) );
  FA_X1 S2_48_25 ( .A(\ab[48][25] ), .B(\CARRYB[47][25] ), .CI(\SUMB[47][26] ), 
        .CO(\CARRYB[48][25] ), .S(\SUMB[48][25] ) );
  FA_X1 S2_48_26 ( .A(\ab[48][26] ), .B(\CARRYB[47][26] ), .CI(\SUMB[47][27] ), 
        .CO(\CARRYB[48][26] ), .S(\SUMB[48][26] ) );
  FA_X1 S2_48_27 ( .A(\ab[48][27] ), .B(\CARRYB[47][27] ), .CI(\SUMB[47][28] ), 
        .CO(\CARRYB[48][27] ), .S(\SUMB[48][27] ) );
  FA_X1 S2_48_28 ( .A(\ab[48][28] ), .B(\CARRYB[47][28] ), .CI(\SUMB[47][29] ), 
        .CO(\CARRYB[48][28] ), .S(\SUMB[48][28] ) );
  FA_X1 S2_48_29 ( .A(\ab[48][29] ), .B(\CARRYB[47][29] ), .CI(\SUMB[47][30] ), 
        .CO(\CARRYB[48][29] ), .S(\SUMB[48][29] ) );
  FA_X1 S2_48_30 ( .A(\ab[48][30] ), .B(\CARRYB[47][30] ), .CI(\SUMB[47][31] ), 
        .CO(\CARRYB[48][30] ), .S(\SUMB[48][30] ) );
  FA_X1 S2_48_31 ( .A(\ab[48][31] ), .B(\CARRYB[47][31] ), .CI(\SUMB[47][32] ), 
        .CO(\CARRYB[48][31] ), .S(\SUMB[48][31] ) );
  FA_X1 S2_48_32 ( .A(\ab[48][32] ), .B(\CARRYB[47][32] ), .CI(\SUMB[47][33] ), 
        .CO(\CARRYB[48][32] ), .S(\SUMB[48][32] ) );
  FA_X1 S2_48_33 ( .A(\ab[48][33] ), .B(\CARRYB[47][33] ), .CI(\SUMB[47][34] ), 
        .CO(\CARRYB[48][33] ), .S(\SUMB[48][33] ) );
  FA_X1 S2_48_34 ( .A(\ab[48][34] ), .B(\CARRYB[47][34] ), .CI(\SUMB[47][35] ), 
        .CO(\CARRYB[48][34] ), .S(\SUMB[48][34] ) );
  FA_X1 S2_48_35 ( .A(\ab[48][35] ), .B(\CARRYB[47][35] ), .CI(\SUMB[47][36] ), 
        .CO(\CARRYB[48][35] ), .S(\SUMB[48][35] ) );
  FA_X1 S2_48_36 ( .A(\ab[48][36] ), .B(\CARRYB[47][36] ), .CI(\SUMB[47][37] ), 
        .CO(\CARRYB[48][36] ), .S(\SUMB[48][36] ) );
  FA_X1 S2_48_37 ( .A(\ab[48][37] ), .B(\CARRYB[47][37] ), .CI(\SUMB[47][38] ), 
        .CO(\CARRYB[48][37] ), .S(\SUMB[48][37] ) );
  FA_X1 S2_48_38 ( .A(\ab[48][38] ), .B(\CARRYB[47][38] ), .CI(\SUMB[47][39] ), 
        .CO(\CARRYB[48][38] ), .S(\SUMB[48][38] ) );
  FA_X1 S2_48_39 ( .A(\ab[48][39] ), .B(\CARRYB[47][39] ), .CI(\SUMB[47][40] ), 
        .CO(\CARRYB[48][39] ), .S(\SUMB[48][39] ) );
  FA_X1 S2_48_40 ( .A(\ab[48][40] ), .B(\CARRYB[47][40] ), .CI(\SUMB[47][41] ), 
        .CO(\CARRYB[48][40] ), .S(\SUMB[48][40] ) );
  FA_X1 S2_48_41 ( .A(\ab[48][41] ), .B(\CARRYB[47][41] ), .CI(\SUMB[47][42] ), 
        .CO(\CARRYB[48][41] ), .S(\SUMB[48][41] ) );
  FA_X1 S2_48_42 ( .A(\ab[48][42] ), .B(\CARRYB[47][42] ), .CI(\SUMB[47][43] ), 
        .CO(\CARRYB[48][42] ), .S(\SUMB[48][42] ) );
  FA_X1 S2_48_43 ( .A(\ab[48][43] ), .B(\CARRYB[47][43] ), .CI(\SUMB[47][44] ), 
        .CO(\CARRYB[48][43] ), .S(\SUMB[48][43] ) );
  FA_X1 S2_48_44 ( .A(\ab[48][44] ), .B(\CARRYB[47][44] ), .CI(\SUMB[47][45] ), 
        .CO(\CARRYB[48][44] ), .S(\SUMB[48][44] ) );
  FA_X1 S2_48_45 ( .A(\ab[48][45] ), .B(\CARRYB[47][45] ), .CI(\SUMB[47][46] ), 
        .CO(\CARRYB[48][45] ), .S(\SUMB[48][45] ) );
  FA_X1 S2_48_46 ( .A(\ab[48][46] ), .B(\CARRYB[47][46] ), .CI(\SUMB[47][47] ), 
        .CO(\CARRYB[48][46] ), .S(\SUMB[48][46] ) );
  FA_X1 S2_48_47 ( .A(\ab[48][47] ), .B(\CARRYB[47][47] ), .CI(\SUMB[47][48] ), 
        .CO(\CARRYB[48][47] ), .S(\SUMB[48][47] ) );
  FA_X1 S2_48_48 ( .A(\ab[48][48] ), .B(\CARRYB[47][48] ), .CI(\SUMB[47][49] ), 
        .CO(\CARRYB[48][48] ), .S(\SUMB[48][48] ) );
  FA_X1 S2_48_49 ( .A(\ab[48][49] ), .B(\CARRYB[47][49] ), .CI(\SUMB[47][50] ), 
        .CO(\CARRYB[48][49] ), .S(\SUMB[48][49] ) );
  FA_X1 S2_48_50 ( .A(\ab[48][50] ), .B(\CARRYB[47][50] ), .CI(\SUMB[47][51] ), 
        .CO(\CARRYB[48][50] ), .S(\SUMB[48][50] ) );
  FA_X1 S3_48_51 ( .A(\ab[48][51] ), .B(\CARRYB[47][51] ), .CI(\ab[47][52] ), 
        .CO(\CARRYB[48][51] ), .S(\SUMB[48][51] ) );
  FA_X1 S1_47_0 ( .A(\ab[47][0] ), .B(\CARRYB[46][0] ), .CI(\SUMB[46][1] ), 
        .CO(\CARRYB[47][0] ), .S(CLA_SUM[47]) );
  FA_X1 S2_47_1 ( .A(\ab[47][1] ), .B(\CARRYB[46][1] ), .CI(\SUMB[46][2] ), 
        .CO(\CARRYB[47][1] ), .S(\SUMB[47][1] ) );
  FA_X1 S2_47_2 ( .A(\ab[47][2] ), .B(\CARRYB[46][2] ), .CI(\SUMB[46][3] ), 
        .CO(\CARRYB[47][2] ), .S(\SUMB[47][2] ) );
  FA_X1 S2_47_3 ( .A(\ab[47][3] ), .B(\CARRYB[46][3] ), .CI(\SUMB[46][4] ), 
        .CO(\CARRYB[47][3] ), .S(\SUMB[47][3] ) );
  FA_X1 S2_47_4 ( .A(\ab[47][4] ), .B(\CARRYB[46][4] ), .CI(\SUMB[46][5] ), 
        .CO(\CARRYB[47][4] ), .S(\SUMB[47][4] ) );
  FA_X1 S2_47_5 ( .A(\ab[47][5] ), .B(\CARRYB[46][5] ), .CI(\SUMB[46][6] ), 
        .CO(\CARRYB[47][5] ), .S(\SUMB[47][5] ) );
  FA_X1 S2_47_6 ( .A(\ab[47][6] ), .B(\CARRYB[46][6] ), .CI(\SUMB[46][7] ), 
        .CO(\CARRYB[47][6] ), .S(\SUMB[47][6] ) );
  FA_X1 S2_47_7 ( .A(\ab[47][7] ), .B(\CARRYB[46][7] ), .CI(\SUMB[46][8] ), 
        .CO(\CARRYB[47][7] ), .S(\SUMB[47][7] ) );
  FA_X1 S2_47_8 ( .A(\ab[47][8] ), .B(\CARRYB[46][8] ), .CI(\SUMB[46][9] ), 
        .CO(\CARRYB[47][8] ), .S(\SUMB[47][8] ) );
  FA_X1 S2_47_9 ( .A(\ab[47][9] ), .B(\CARRYB[46][9] ), .CI(\SUMB[46][10] ), 
        .CO(\CARRYB[47][9] ), .S(\SUMB[47][9] ) );
  FA_X1 S2_47_10 ( .A(\ab[47][10] ), .B(\CARRYB[46][10] ), .CI(\SUMB[46][11] ), 
        .CO(\CARRYB[47][10] ), .S(\SUMB[47][10] ) );
  FA_X1 S2_47_11 ( .A(\ab[47][11] ), .B(\CARRYB[46][11] ), .CI(\SUMB[46][12] ), 
        .CO(\CARRYB[47][11] ), .S(\SUMB[47][11] ) );
  FA_X1 S2_47_12 ( .A(\ab[47][12] ), .B(\CARRYB[46][12] ), .CI(\SUMB[46][13] ), 
        .CO(\CARRYB[47][12] ), .S(\SUMB[47][12] ) );
  FA_X1 S2_47_13 ( .A(\ab[47][13] ), .B(\CARRYB[46][13] ), .CI(\SUMB[46][14] ), 
        .CO(\CARRYB[47][13] ), .S(\SUMB[47][13] ) );
  FA_X1 S2_47_14 ( .A(\ab[47][14] ), .B(\CARRYB[46][14] ), .CI(\SUMB[46][15] ), 
        .CO(\CARRYB[47][14] ), .S(\SUMB[47][14] ) );
  FA_X1 S2_47_15 ( .A(\ab[47][15] ), .B(\CARRYB[46][15] ), .CI(\SUMB[46][16] ), 
        .CO(\CARRYB[47][15] ), .S(\SUMB[47][15] ) );
  FA_X1 S2_47_16 ( .A(\ab[47][16] ), .B(\CARRYB[46][16] ), .CI(\SUMB[46][17] ), 
        .CO(\CARRYB[47][16] ), .S(\SUMB[47][16] ) );
  FA_X1 S2_47_17 ( .A(\ab[47][17] ), .B(\CARRYB[46][17] ), .CI(\SUMB[46][18] ), 
        .CO(\CARRYB[47][17] ), .S(\SUMB[47][17] ) );
  FA_X1 S2_47_18 ( .A(\ab[47][18] ), .B(\CARRYB[46][18] ), .CI(\SUMB[46][19] ), 
        .CO(\CARRYB[47][18] ), .S(\SUMB[47][18] ) );
  FA_X1 S2_47_19 ( .A(\ab[47][19] ), .B(\CARRYB[46][19] ), .CI(\SUMB[46][20] ), 
        .CO(\CARRYB[47][19] ), .S(\SUMB[47][19] ) );
  FA_X1 S2_47_20 ( .A(\ab[47][20] ), .B(\CARRYB[46][20] ), .CI(\SUMB[46][21] ), 
        .CO(\CARRYB[47][20] ), .S(\SUMB[47][20] ) );
  FA_X1 S2_47_21 ( .A(\ab[47][21] ), .B(\CARRYB[46][21] ), .CI(\SUMB[46][22] ), 
        .CO(\CARRYB[47][21] ), .S(\SUMB[47][21] ) );
  FA_X1 S2_47_22 ( .A(\ab[47][22] ), .B(\CARRYB[46][22] ), .CI(\SUMB[46][23] ), 
        .CO(\CARRYB[47][22] ), .S(\SUMB[47][22] ) );
  FA_X1 S2_47_23 ( .A(\ab[47][23] ), .B(\CARRYB[46][23] ), .CI(\SUMB[46][24] ), 
        .CO(\CARRYB[47][23] ), .S(\SUMB[47][23] ) );
  FA_X1 S2_47_24 ( .A(\ab[47][24] ), .B(\CARRYB[46][24] ), .CI(\SUMB[46][25] ), 
        .CO(\CARRYB[47][24] ), .S(\SUMB[47][24] ) );
  FA_X1 S2_47_25 ( .A(\ab[47][25] ), .B(\CARRYB[46][25] ), .CI(\SUMB[46][26] ), 
        .CO(\CARRYB[47][25] ), .S(\SUMB[47][25] ) );
  FA_X1 S2_47_26 ( .A(\ab[47][26] ), .B(\CARRYB[46][26] ), .CI(\SUMB[46][27] ), 
        .CO(\CARRYB[47][26] ), .S(\SUMB[47][26] ) );
  FA_X1 S2_47_27 ( .A(\ab[47][27] ), .B(\CARRYB[46][27] ), .CI(\SUMB[46][28] ), 
        .CO(\CARRYB[47][27] ), .S(\SUMB[47][27] ) );
  FA_X1 S2_47_28 ( .A(\ab[47][28] ), .B(\CARRYB[46][28] ), .CI(\SUMB[46][29] ), 
        .CO(\CARRYB[47][28] ), .S(\SUMB[47][28] ) );
  FA_X1 S2_47_29 ( .A(\ab[47][29] ), .B(\CARRYB[46][29] ), .CI(\SUMB[46][30] ), 
        .CO(\CARRYB[47][29] ), .S(\SUMB[47][29] ) );
  FA_X1 S2_47_30 ( .A(\ab[47][30] ), .B(\CARRYB[46][30] ), .CI(\SUMB[46][31] ), 
        .CO(\CARRYB[47][30] ), .S(\SUMB[47][30] ) );
  FA_X1 S2_47_31 ( .A(\ab[47][31] ), .B(\CARRYB[46][31] ), .CI(\SUMB[46][32] ), 
        .CO(\CARRYB[47][31] ), .S(\SUMB[47][31] ) );
  FA_X1 S2_47_32 ( .A(\ab[47][32] ), .B(\CARRYB[46][32] ), .CI(\SUMB[46][33] ), 
        .CO(\CARRYB[47][32] ), .S(\SUMB[47][32] ) );
  FA_X1 S2_47_33 ( .A(\ab[47][33] ), .B(\CARRYB[46][33] ), .CI(\SUMB[46][34] ), 
        .CO(\CARRYB[47][33] ), .S(\SUMB[47][33] ) );
  FA_X1 S2_47_34 ( .A(\ab[47][34] ), .B(\CARRYB[46][34] ), .CI(\SUMB[46][35] ), 
        .CO(\CARRYB[47][34] ), .S(\SUMB[47][34] ) );
  FA_X1 S2_47_35 ( .A(\ab[47][35] ), .B(\CARRYB[46][35] ), .CI(\SUMB[46][36] ), 
        .CO(\CARRYB[47][35] ), .S(\SUMB[47][35] ) );
  FA_X1 S2_47_36 ( .A(\ab[47][36] ), .B(\CARRYB[46][36] ), .CI(\SUMB[46][37] ), 
        .CO(\CARRYB[47][36] ), .S(\SUMB[47][36] ) );
  FA_X1 S2_47_37 ( .A(\ab[47][37] ), .B(\CARRYB[46][37] ), .CI(\SUMB[46][38] ), 
        .CO(\CARRYB[47][37] ), .S(\SUMB[47][37] ) );
  FA_X1 S2_47_38 ( .A(\ab[47][38] ), .B(\CARRYB[46][38] ), .CI(\SUMB[46][39] ), 
        .CO(\CARRYB[47][38] ), .S(\SUMB[47][38] ) );
  FA_X1 S2_47_39 ( .A(\ab[47][39] ), .B(\CARRYB[46][39] ), .CI(\SUMB[46][40] ), 
        .CO(\CARRYB[47][39] ), .S(\SUMB[47][39] ) );
  FA_X1 S2_47_40 ( .A(\ab[47][40] ), .B(\CARRYB[46][40] ), .CI(\SUMB[46][41] ), 
        .CO(\CARRYB[47][40] ), .S(\SUMB[47][40] ) );
  FA_X1 S2_47_41 ( .A(\ab[47][41] ), .B(\CARRYB[46][41] ), .CI(\SUMB[46][42] ), 
        .CO(\CARRYB[47][41] ), .S(\SUMB[47][41] ) );
  FA_X1 S2_47_42 ( .A(\ab[47][42] ), .B(\CARRYB[46][42] ), .CI(\SUMB[46][43] ), 
        .CO(\CARRYB[47][42] ), .S(\SUMB[47][42] ) );
  FA_X1 S2_47_43 ( .A(\ab[47][43] ), .B(\CARRYB[46][43] ), .CI(\SUMB[46][44] ), 
        .CO(\CARRYB[47][43] ), .S(\SUMB[47][43] ) );
  FA_X1 S2_47_44 ( .A(\ab[47][44] ), .B(\CARRYB[46][44] ), .CI(\SUMB[46][45] ), 
        .CO(\CARRYB[47][44] ), .S(\SUMB[47][44] ) );
  FA_X1 S2_47_45 ( .A(\ab[47][45] ), .B(\CARRYB[46][45] ), .CI(\SUMB[46][46] ), 
        .CO(\CARRYB[47][45] ), .S(\SUMB[47][45] ) );
  FA_X1 S2_47_46 ( .A(\ab[47][46] ), .B(\CARRYB[46][46] ), .CI(\SUMB[46][47] ), 
        .CO(\CARRYB[47][46] ), .S(\SUMB[47][46] ) );
  FA_X1 S2_47_47 ( .A(\ab[47][47] ), .B(\CARRYB[46][47] ), .CI(\SUMB[46][48] ), 
        .CO(\CARRYB[47][47] ), .S(\SUMB[47][47] ) );
  FA_X1 S2_47_48 ( .A(\ab[47][48] ), .B(\CARRYB[46][48] ), .CI(\SUMB[46][49] ), 
        .CO(\CARRYB[47][48] ), .S(\SUMB[47][48] ) );
  FA_X1 S2_47_49 ( .A(\ab[47][49] ), .B(\CARRYB[46][49] ), .CI(\SUMB[46][50] ), 
        .CO(\CARRYB[47][49] ), .S(\SUMB[47][49] ) );
  FA_X1 S2_47_50 ( .A(\ab[47][50] ), .B(\CARRYB[46][50] ), .CI(\SUMB[46][51] ), 
        .CO(\CARRYB[47][50] ), .S(\SUMB[47][50] ) );
  FA_X1 S3_47_51 ( .A(\ab[47][51] ), .B(\CARRYB[46][51] ), .CI(\ab[46][52] ), 
        .CO(\CARRYB[47][51] ), .S(\SUMB[47][51] ) );
  FA_X1 S1_46_0 ( .A(\ab[46][0] ), .B(\CARRYB[45][0] ), .CI(\SUMB[45][1] ), 
        .CO(\CARRYB[46][0] ), .S(CLA_SUM[46]) );
  FA_X1 S2_46_1 ( .A(\ab[46][1] ), .B(\CARRYB[45][1] ), .CI(\SUMB[45][2] ), 
        .CO(\CARRYB[46][1] ), .S(\SUMB[46][1] ) );
  FA_X1 S2_46_2 ( .A(\ab[46][2] ), .B(\CARRYB[45][2] ), .CI(\SUMB[45][3] ), 
        .CO(\CARRYB[46][2] ), .S(\SUMB[46][2] ) );
  FA_X1 S2_46_3 ( .A(\ab[46][3] ), .B(\CARRYB[45][3] ), .CI(\SUMB[45][4] ), 
        .CO(\CARRYB[46][3] ), .S(\SUMB[46][3] ) );
  FA_X1 S2_46_4 ( .A(\ab[46][4] ), .B(\CARRYB[45][4] ), .CI(\SUMB[45][5] ), 
        .CO(\CARRYB[46][4] ), .S(\SUMB[46][4] ) );
  FA_X1 S2_46_5 ( .A(\ab[46][5] ), .B(\CARRYB[45][5] ), .CI(\SUMB[45][6] ), 
        .CO(\CARRYB[46][5] ), .S(\SUMB[46][5] ) );
  FA_X1 S2_46_6 ( .A(\ab[46][6] ), .B(\CARRYB[45][6] ), .CI(\SUMB[45][7] ), 
        .CO(\CARRYB[46][6] ), .S(\SUMB[46][6] ) );
  FA_X1 S2_46_7 ( .A(\ab[46][7] ), .B(\CARRYB[45][7] ), .CI(\SUMB[45][8] ), 
        .CO(\CARRYB[46][7] ), .S(\SUMB[46][7] ) );
  FA_X1 S2_46_8 ( .A(\ab[46][8] ), .B(\CARRYB[45][8] ), .CI(\SUMB[45][9] ), 
        .CO(\CARRYB[46][8] ), .S(\SUMB[46][8] ) );
  FA_X1 S2_46_9 ( .A(\ab[46][9] ), .B(\CARRYB[45][9] ), .CI(\SUMB[45][10] ), 
        .CO(\CARRYB[46][9] ), .S(\SUMB[46][9] ) );
  FA_X1 S2_46_10 ( .A(\ab[46][10] ), .B(\CARRYB[45][10] ), .CI(\SUMB[45][11] ), 
        .CO(\CARRYB[46][10] ), .S(\SUMB[46][10] ) );
  FA_X1 S2_46_11 ( .A(\ab[46][11] ), .B(\CARRYB[45][11] ), .CI(\SUMB[45][12] ), 
        .CO(\CARRYB[46][11] ), .S(\SUMB[46][11] ) );
  FA_X1 S2_46_12 ( .A(\ab[46][12] ), .B(\CARRYB[45][12] ), .CI(\SUMB[45][13] ), 
        .CO(\CARRYB[46][12] ), .S(\SUMB[46][12] ) );
  FA_X1 S2_46_13 ( .A(\ab[46][13] ), .B(\CARRYB[45][13] ), .CI(\SUMB[45][14] ), 
        .CO(\CARRYB[46][13] ), .S(\SUMB[46][13] ) );
  FA_X1 S2_46_14 ( .A(\ab[46][14] ), .B(\CARRYB[45][14] ), .CI(\SUMB[45][15] ), 
        .CO(\CARRYB[46][14] ), .S(\SUMB[46][14] ) );
  FA_X1 S2_46_15 ( .A(\ab[46][15] ), .B(\CARRYB[45][15] ), .CI(\SUMB[45][16] ), 
        .CO(\CARRYB[46][15] ), .S(\SUMB[46][15] ) );
  FA_X1 S2_46_16 ( .A(\ab[46][16] ), .B(\CARRYB[45][16] ), .CI(\SUMB[45][17] ), 
        .CO(\CARRYB[46][16] ), .S(\SUMB[46][16] ) );
  FA_X1 S2_46_17 ( .A(\ab[46][17] ), .B(\CARRYB[45][17] ), .CI(\SUMB[45][18] ), 
        .CO(\CARRYB[46][17] ), .S(\SUMB[46][17] ) );
  FA_X1 S2_46_18 ( .A(\ab[46][18] ), .B(\CARRYB[45][18] ), .CI(\SUMB[45][19] ), 
        .CO(\CARRYB[46][18] ), .S(\SUMB[46][18] ) );
  FA_X1 S2_46_19 ( .A(\ab[46][19] ), .B(\CARRYB[45][19] ), .CI(\SUMB[45][20] ), 
        .CO(\CARRYB[46][19] ), .S(\SUMB[46][19] ) );
  FA_X1 S2_46_20 ( .A(\ab[46][20] ), .B(\CARRYB[45][20] ), .CI(\SUMB[45][21] ), 
        .CO(\CARRYB[46][20] ), .S(\SUMB[46][20] ) );
  FA_X1 S2_46_21 ( .A(\ab[46][21] ), .B(\CARRYB[45][21] ), .CI(\SUMB[45][22] ), 
        .CO(\CARRYB[46][21] ), .S(\SUMB[46][21] ) );
  FA_X1 S2_46_22 ( .A(\ab[46][22] ), .B(\CARRYB[45][22] ), .CI(\SUMB[45][23] ), 
        .CO(\CARRYB[46][22] ), .S(\SUMB[46][22] ) );
  FA_X1 S2_46_23 ( .A(\ab[46][23] ), .B(\CARRYB[45][23] ), .CI(\SUMB[45][24] ), 
        .CO(\CARRYB[46][23] ), .S(\SUMB[46][23] ) );
  FA_X1 S2_46_24 ( .A(\ab[46][24] ), .B(\CARRYB[45][24] ), .CI(\SUMB[45][25] ), 
        .CO(\CARRYB[46][24] ), .S(\SUMB[46][24] ) );
  FA_X1 S2_46_25 ( .A(\ab[46][25] ), .B(\CARRYB[45][25] ), .CI(\SUMB[45][26] ), 
        .CO(\CARRYB[46][25] ), .S(\SUMB[46][25] ) );
  FA_X1 S2_46_26 ( .A(\ab[46][26] ), .B(\CARRYB[45][26] ), .CI(\SUMB[45][27] ), 
        .CO(\CARRYB[46][26] ), .S(\SUMB[46][26] ) );
  FA_X1 S2_46_27 ( .A(\ab[46][27] ), .B(\CARRYB[45][27] ), .CI(\SUMB[45][28] ), 
        .CO(\CARRYB[46][27] ), .S(\SUMB[46][27] ) );
  FA_X1 S2_46_28 ( .A(\ab[46][28] ), .B(\CARRYB[45][28] ), .CI(\SUMB[45][29] ), 
        .CO(\CARRYB[46][28] ), .S(\SUMB[46][28] ) );
  FA_X1 S2_46_29 ( .A(\ab[46][29] ), .B(\CARRYB[45][29] ), .CI(\SUMB[45][30] ), 
        .CO(\CARRYB[46][29] ), .S(\SUMB[46][29] ) );
  FA_X1 S2_46_30 ( .A(\ab[46][30] ), .B(\CARRYB[45][30] ), .CI(\SUMB[45][31] ), 
        .CO(\CARRYB[46][30] ), .S(\SUMB[46][30] ) );
  FA_X1 S2_46_31 ( .A(\ab[46][31] ), .B(\CARRYB[45][31] ), .CI(\SUMB[45][32] ), 
        .CO(\CARRYB[46][31] ), .S(\SUMB[46][31] ) );
  FA_X1 S2_46_32 ( .A(\ab[46][32] ), .B(\CARRYB[45][32] ), .CI(\SUMB[45][33] ), 
        .CO(\CARRYB[46][32] ), .S(\SUMB[46][32] ) );
  FA_X1 S2_46_33 ( .A(\ab[46][33] ), .B(\CARRYB[45][33] ), .CI(\SUMB[45][34] ), 
        .CO(\CARRYB[46][33] ), .S(\SUMB[46][33] ) );
  FA_X1 S2_46_34 ( .A(\ab[46][34] ), .B(\CARRYB[45][34] ), .CI(\SUMB[45][35] ), 
        .CO(\CARRYB[46][34] ), .S(\SUMB[46][34] ) );
  FA_X1 S2_46_35 ( .A(\ab[46][35] ), .B(\CARRYB[45][35] ), .CI(\SUMB[45][36] ), 
        .CO(\CARRYB[46][35] ), .S(\SUMB[46][35] ) );
  FA_X1 S2_46_36 ( .A(\ab[46][36] ), .B(\CARRYB[45][36] ), .CI(\SUMB[45][37] ), 
        .CO(\CARRYB[46][36] ), .S(\SUMB[46][36] ) );
  FA_X1 S2_46_37 ( .A(\ab[46][37] ), .B(\CARRYB[45][37] ), .CI(\SUMB[45][38] ), 
        .CO(\CARRYB[46][37] ), .S(\SUMB[46][37] ) );
  FA_X1 S2_46_38 ( .A(\ab[46][38] ), .B(\CARRYB[45][38] ), .CI(\SUMB[45][39] ), 
        .CO(\CARRYB[46][38] ), .S(\SUMB[46][38] ) );
  FA_X1 S2_46_39 ( .A(\ab[46][39] ), .B(\CARRYB[45][39] ), .CI(\SUMB[45][40] ), 
        .CO(\CARRYB[46][39] ), .S(\SUMB[46][39] ) );
  FA_X1 S2_46_40 ( .A(\ab[46][40] ), .B(\CARRYB[45][40] ), .CI(\SUMB[45][41] ), 
        .CO(\CARRYB[46][40] ), .S(\SUMB[46][40] ) );
  FA_X1 S2_46_41 ( .A(\ab[46][41] ), .B(\CARRYB[45][41] ), .CI(\SUMB[45][42] ), 
        .CO(\CARRYB[46][41] ), .S(\SUMB[46][41] ) );
  FA_X1 S2_46_42 ( .A(\ab[46][42] ), .B(\CARRYB[45][42] ), .CI(\SUMB[45][43] ), 
        .CO(\CARRYB[46][42] ), .S(\SUMB[46][42] ) );
  FA_X1 S2_46_43 ( .A(\ab[46][43] ), .B(\CARRYB[45][43] ), .CI(\SUMB[45][44] ), 
        .CO(\CARRYB[46][43] ), .S(\SUMB[46][43] ) );
  FA_X1 S2_46_44 ( .A(\ab[46][44] ), .B(\CARRYB[45][44] ), .CI(\SUMB[45][45] ), 
        .CO(\CARRYB[46][44] ), .S(\SUMB[46][44] ) );
  FA_X1 S2_46_45 ( .A(\ab[46][45] ), .B(\CARRYB[45][45] ), .CI(\SUMB[45][46] ), 
        .CO(\CARRYB[46][45] ), .S(\SUMB[46][45] ) );
  FA_X1 S2_46_46 ( .A(\ab[46][46] ), .B(\CARRYB[45][46] ), .CI(\SUMB[45][47] ), 
        .CO(\CARRYB[46][46] ), .S(\SUMB[46][46] ) );
  FA_X1 S2_46_47 ( .A(\ab[46][47] ), .B(\CARRYB[45][47] ), .CI(\SUMB[45][48] ), 
        .CO(\CARRYB[46][47] ), .S(\SUMB[46][47] ) );
  FA_X1 S2_46_48 ( .A(\ab[46][48] ), .B(\CARRYB[45][48] ), .CI(\SUMB[45][49] ), 
        .CO(\CARRYB[46][48] ), .S(\SUMB[46][48] ) );
  FA_X1 S2_46_49 ( .A(\ab[46][49] ), .B(\CARRYB[45][49] ), .CI(\SUMB[45][50] ), 
        .CO(\CARRYB[46][49] ), .S(\SUMB[46][49] ) );
  FA_X1 S2_46_50 ( .A(\ab[46][50] ), .B(\CARRYB[45][50] ), .CI(\SUMB[45][51] ), 
        .CO(\CARRYB[46][50] ), .S(\SUMB[46][50] ) );
  FA_X1 S3_46_51 ( .A(\ab[46][51] ), .B(\CARRYB[45][51] ), .CI(\ab[45][52] ), 
        .CO(\CARRYB[46][51] ), .S(\SUMB[46][51] ) );
  FA_X1 S1_45_0 ( .A(\ab[45][0] ), .B(\CARRYB[44][0] ), .CI(\SUMB[44][1] ), 
        .CO(\CARRYB[45][0] ), .S(CLA_SUM[45]) );
  FA_X1 S2_45_1 ( .A(\ab[45][1] ), .B(\CARRYB[44][1] ), .CI(\SUMB[44][2] ), 
        .CO(\CARRYB[45][1] ), .S(\SUMB[45][1] ) );
  FA_X1 S2_45_2 ( .A(\ab[45][2] ), .B(\CARRYB[44][2] ), .CI(\SUMB[44][3] ), 
        .CO(\CARRYB[45][2] ), .S(\SUMB[45][2] ) );
  FA_X1 S2_45_3 ( .A(\ab[45][3] ), .B(\CARRYB[44][3] ), .CI(\SUMB[44][4] ), 
        .CO(\CARRYB[45][3] ), .S(\SUMB[45][3] ) );
  FA_X1 S2_45_4 ( .A(\ab[45][4] ), .B(\CARRYB[44][4] ), .CI(\SUMB[44][5] ), 
        .CO(\CARRYB[45][4] ), .S(\SUMB[45][4] ) );
  FA_X1 S2_45_5 ( .A(\ab[45][5] ), .B(\CARRYB[44][5] ), .CI(\SUMB[44][6] ), 
        .CO(\CARRYB[45][5] ), .S(\SUMB[45][5] ) );
  FA_X1 S2_45_6 ( .A(\ab[45][6] ), .B(\CARRYB[44][6] ), .CI(\SUMB[44][7] ), 
        .CO(\CARRYB[45][6] ), .S(\SUMB[45][6] ) );
  FA_X1 S2_45_7 ( .A(\ab[45][7] ), .B(\CARRYB[44][7] ), .CI(\SUMB[44][8] ), 
        .CO(\CARRYB[45][7] ), .S(\SUMB[45][7] ) );
  FA_X1 S2_45_8 ( .A(\ab[45][8] ), .B(\CARRYB[44][8] ), .CI(\SUMB[44][9] ), 
        .CO(\CARRYB[45][8] ), .S(\SUMB[45][8] ) );
  FA_X1 S2_45_9 ( .A(\ab[45][9] ), .B(\CARRYB[44][9] ), .CI(\SUMB[44][10] ), 
        .CO(\CARRYB[45][9] ), .S(\SUMB[45][9] ) );
  FA_X1 S2_45_10 ( .A(\ab[45][10] ), .B(\CARRYB[44][10] ), .CI(\SUMB[44][11] ), 
        .CO(\CARRYB[45][10] ), .S(\SUMB[45][10] ) );
  FA_X1 S2_45_11 ( .A(\ab[45][11] ), .B(\CARRYB[44][11] ), .CI(\SUMB[44][12] ), 
        .CO(\CARRYB[45][11] ), .S(\SUMB[45][11] ) );
  FA_X1 S2_45_12 ( .A(\ab[45][12] ), .B(\CARRYB[44][12] ), .CI(\SUMB[44][13] ), 
        .CO(\CARRYB[45][12] ), .S(\SUMB[45][12] ) );
  FA_X1 S2_45_13 ( .A(\ab[45][13] ), .B(\CARRYB[44][13] ), .CI(\SUMB[44][14] ), 
        .CO(\CARRYB[45][13] ), .S(\SUMB[45][13] ) );
  FA_X1 S2_45_14 ( .A(\ab[45][14] ), .B(\CARRYB[44][14] ), .CI(\SUMB[44][15] ), 
        .CO(\CARRYB[45][14] ), .S(\SUMB[45][14] ) );
  FA_X1 S2_45_15 ( .A(\ab[45][15] ), .B(\CARRYB[44][15] ), .CI(\SUMB[44][16] ), 
        .CO(\CARRYB[45][15] ), .S(\SUMB[45][15] ) );
  FA_X1 S2_45_16 ( .A(\ab[45][16] ), .B(\CARRYB[44][16] ), .CI(\SUMB[44][17] ), 
        .CO(\CARRYB[45][16] ), .S(\SUMB[45][16] ) );
  FA_X1 S2_45_17 ( .A(\ab[45][17] ), .B(\CARRYB[44][17] ), .CI(\SUMB[44][18] ), 
        .CO(\CARRYB[45][17] ), .S(\SUMB[45][17] ) );
  FA_X1 S2_45_18 ( .A(\ab[45][18] ), .B(\CARRYB[44][18] ), .CI(\SUMB[44][19] ), 
        .CO(\CARRYB[45][18] ), .S(\SUMB[45][18] ) );
  FA_X1 S2_45_19 ( .A(\ab[45][19] ), .B(\CARRYB[44][19] ), .CI(\SUMB[44][20] ), 
        .CO(\CARRYB[45][19] ), .S(\SUMB[45][19] ) );
  FA_X1 S2_45_20 ( .A(\ab[45][20] ), .B(\CARRYB[44][20] ), .CI(\SUMB[44][21] ), 
        .CO(\CARRYB[45][20] ), .S(\SUMB[45][20] ) );
  FA_X1 S2_45_21 ( .A(\ab[45][21] ), .B(\CARRYB[44][21] ), .CI(\SUMB[44][22] ), 
        .CO(\CARRYB[45][21] ), .S(\SUMB[45][21] ) );
  FA_X1 S2_45_22 ( .A(\ab[45][22] ), .B(\CARRYB[44][22] ), .CI(\SUMB[44][23] ), 
        .CO(\CARRYB[45][22] ), .S(\SUMB[45][22] ) );
  FA_X1 S2_45_23 ( .A(\ab[45][23] ), .B(\CARRYB[44][23] ), .CI(\SUMB[44][24] ), 
        .CO(\CARRYB[45][23] ), .S(\SUMB[45][23] ) );
  FA_X1 S2_45_24 ( .A(\ab[45][24] ), .B(\CARRYB[44][24] ), .CI(\SUMB[44][25] ), 
        .CO(\CARRYB[45][24] ), .S(\SUMB[45][24] ) );
  FA_X1 S2_45_25 ( .A(\ab[45][25] ), .B(\CARRYB[44][25] ), .CI(\SUMB[44][26] ), 
        .CO(\CARRYB[45][25] ), .S(\SUMB[45][25] ) );
  FA_X1 S2_45_26 ( .A(\ab[45][26] ), .B(\CARRYB[44][26] ), .CI(\SUMB[44][27] ), 
        .CO(\CARRYB[45][26] ), .S(\SUMB[45][26] ) );
  FA_X1 S2_45_27 ( .A(\ab[45][27] ), .B(\CARRYB[44][27] ), .CI(\SUMB[44][28] ), 
        .CO(\CARRYB[45][27] ), .S(\SUMB[45][27] ) );
  FA_X1 S2_45_28 ( .A(\ab[45][28] ), .B(\CARRYB[44][28] ), .CI(\SUMB[44][29] ), 
        .CO(\CARRYB[45][28] ), .S(\SUMB[45][28] ) );
  FA_X1 S2_45_29 ( .A(\ab[45][29] ), .B(\CARRYB[44][29] ), .CI(\SUMB[44][30] ), 
        .CO(\CARRYB[45][29] ), .S(\SUMB[45][29] ) );
  FA_X1 S2_45_30 ( .A(\ab[45][30] ), .B(\CARRYB[44][30] ), .CI(\SUMB[44][31] ), 
        .CO(\CARRYB[45][30] ), .S(\SUMB[45][30] ) );
  FA_X1 S2_45_31 ( .A(\ab[45][31] ), .B(\CARRYB[44][31] ), .CI(\SUMB[44][32] ), 
        .CO(\CARRYB[45][31] ), .S(\SUMB[45][31] ) );
  FA_X1 S2_45_32 ( .A(\ab[45][32] ), .B(\CARRYB[44][32] ), .CI(\SUMB[44][33] ), 
        .CO(\CARRYB[45][32] ), .S(\SUMB[45][32] ) );
  FA_X1 S2_45_33 ( .A(\ab[45][33] ), .B(\CARRYB[44][33] ), .CI(\SUMB[44][34] ), 
        .CO(\CARRYB[45][33] ), .S(\SUMB[45][33] ) );
  FA_X1 S2_45_34 ( .A(\ab[45][34] ), .B(\CARRYB[44][34] ), .CI(\SUMB[44][35] ), 
        .CO(\CARRYB[45][34] ), .S(\SUMB[45][34] ) );
  FA_X1 S2_45_35 ( .A(\ab[45][35] ), .B(\CARRYB[44][35] ), .CI(\SUMB[44][36] ), 
        .CO(\CARRYB[45][35] ), .S(\SUMB[45][35] ) );
  FA_X1 S2_45_36 ( .A(\ab[45][36] ), .B(\CARRYB[44][36] ), .CI(\SUMB[44][37] ), 
        .CO(\CARRYB[45][36] ), .S(\SUMB[45][36] ) );
  FA_X1 S2_45_37 ( .A(\ab[45][37] ), .B(\CARRYB[44][37] ), .CI(\SUMB[44][38] ), 
        .CO(\CARRYB[45][37] ), .S(\SUMB[45][37] ) );
  FA_X1 S2_45_38 ( .A(\ab[45][38] ), .B(\CARRYB[44][38] ), .CI(\SUMB[44][39] ), 
        .CO(\CARRYB[45][38] ), .S(\SUMB[45][38] ) );
  FA_X1 S2_45_39 ( .A(\ab[45][39] ), .B(\CARRYB[44][39] ), .CI(\SUMB[44][40] ), 
        .CO(\CARRYB[45][39] ), .S(\SUMB[45][39] ) );
  FA_X1 S2_45_40 ( .A(\ab[45][40] ), .B(\CARRYB[44][40] ), .CI(\SUMB[44][41] ), 
        .CO(\CARRYB[45][40] ), .S(\SUMB[45][40] ) );
  FA_X1 S2_45_41 ( .A(\ab[45][41] ), .B(\CARRYB[44][41] ), .CI(\SUMB[44][42] ), 
        .CO(\CARRYB[45][41] ), .S(\SUMB[45][41] ) );
  FA_X1 S2_45_42 ( .A(\ab[45][42] ), .B(\CARRYB[44][42] ), .CI(\SUMB[44][43] ), 
        .CO(\CARRYB[45][42] ), .S(\SUMB[45][42] ) );
  FA_X1 S2_45_43 ( .A(\ab[45][43] ), .B(\CARRYB[44][43] ), .CI(\SUMB[44][44] ), 
        .CO(\CARRYB[45][43] ), .S(\SUMB[45][43] ) );
  FA_X1 S2_45_44 ( .A(\ab[45][44] ), .B(\CARRYB[44][44] ), .CI(\SUMB[44][45] ), 
        .CO(\CARRYB[45][44] ), .S(\SUMB[45][44] ) );
  FA_X1 S2_45_45 ( .A(\ab[45][45] ), .B(\CARRYB[44][45] ), .CI(\SUMB[44][46] ), 
        .CO(\CARRYB[45][45] ), .S(\SUMB[45][45] ) );
  FA_X1 S2_45_46 ( .A(\ab[45][46] ), .B(\CARRYB[44][46] ), .CI(\SUMB[44][47] ), 
        .CO(\CARRYB[45][46] ), .S(\SUMB[45][46] ) );
  FA_X1 S2_45_47 ( .A(\ab[45][47] ), .B(\CARRYB[44][47] ), .CI(\SUMB[44][48] ), 
        .CO(\CARRYB[45][47] ), .S(\SUMB[45][47] ) );
  FA_X1 S2_45_48 ( .A(\ab[45][48] ), .B(\CARRYB[44][48] ), .CI(\SUMB[44][49] ), 
        .CO(\CARRYB[45][48] ), .S(\SUMB[45][48] ) );
  FA_X1 S2_45_49 ( .A(\ab[45][49] ), .B(\CARRYB[44][49] ), .CI(\SUMB[44][50] ), 
        .CO(\CARRYB[45][49] ), .S(\SUMB[45][49] ) );
  FA_X1 S2_45_50 ( .A(\ab[45][50] ), .B(\CARRYB[44][50] ), .CI(\SUMB[44][51] ), 
        .CO(\CARRYB[45][50] ), .S(\SUMB[45][50] ) );
  FA_X1 S3_45_51 ( .A(\ab[45][51] ), .B(\CARRYB[44][51] ), .CI(\ab[44][52] ), 
        .CO(\CARRYB[45][51] ), .S(\SUMB[45][51] ) );
  FA_X1 S1_44_0 ( .A(\ab[44][0] ), .B(\CARRYB[43][0] ), .CI(\SUMB[43][1] ), 
        .CO(\CARRYB[44][0] ), .S(CLA_SUM[44]) );
  FA_X1 S2_44_1 ( .A(\ab[44][1] ), .B(\CARRYB[43][1] ), .CI(\SUMB[43][2] ), 
        .CO(\CARRYB[44][1] ), .S(\SUMB[44][1] ) );
  FA_X1 S2_44_2 ( .A(\ab[44][2] ), .B(\CARRYB[43][2] ), .CI(\SUMB[43][3] ), 
        .CO(\CARRYB[44][2] ), .S(\SUMB[44][2] ) );
  FA_X1 S2_44_3 ( .A(\ab[44][3] ), .B(\CARRYB[43][3] ), .CI(\SUMB[43][4] ), 
        .CO(\CARRYB[44][3] ), .S(\SUMB[44][3] ) );
  FA_X1 S2_44_4 ( .A(\ab[44][4] ), .B(\CARRYB[43][4] ), .CI(\SUMB[43][5] ), 
        .CO(\CARRYB[44][4] ), .S(\SUMB[44][4] ) );
  FA_X1 S2_44_5 ( .A(\ab[44][5] ), .B(\CARRYB[43][5] ), .CI(\SUMB[43][6] ), 
        .CO(\CARRYB[44][5] ), .S(\SUMB[44][5] ) );
  FA_X1 S2_44_6 ( .A(\ab[44][6] ), .B(\CARRYB[43][6] ), .CI(\SUMB[43][7] ), 
        .CO(\CARRYB[44][6] ), .S(\SUMB[44][6] ) );
  FA_X1 S2_44_7 ( .A(\ab[44][7] ), .B(\CARRYB[43][7] ), .CI(\SUMB[43][8] ), 
        .CO(\CARRYB[44][7] ), .S(\SUMB[44][7] ) );
  FA_X1 S2_44_8 ( .A(\ab[44][8] ), .B(\CARRYB[43][8] ), .CI(\SUMB[43][9] ), 
        .CO(\CARRYB[44][8] ), .S(\SUMB[44][8] ) );
  FA_X1 S2_44_9 ( .A(\ab[44][9] ), .B(\CARRYB[43][9] ), .CI(\SUMB[43][10] ), 
        .CO(\CARRYB[44][9] ), .S(\SUMB[44][9] ) );
  FA_X1 S2_44_10 ( .A(\ab[44][10] ), .B(\CARRYB[43][10] ), .CI(\SUMB[43][11] ), 
        .CO(\CARRYB[44][10] ), .S(\SUMB[44][10] ) );
  FA_X1 S2_44_11 ( .A(\ab[44][11] ), .B(\CARRYB[43][11] ), .CI(\SUMB[43][12] ), 
        .CO(\CARRYB[44][11] ), .S(\SUMB[44][11] ) );
  FA_X1 S2_44_12 ( .A(\ab[44][12] ), .B(\CARRYB[43][12] ), .CI(\SUMB[43][13] ), 
        .CO(\CARRYB[44][12] ), .S(\SUMB[44][12] ) );
  FA_X1 S2_44_13 ( .A(\ab[44][13] ), .B(\CARRYB[43][13] ), .CI(\SUMB[43][14] ), 
        .CO(\CARRYB[44][13] ), .S(\SUMB[44][13] ) );
  FA_X1 S2_44_14 ( .A(\ab[44][14] ), .B(\CARRYB[43][14] ), .CI(\SUMB[43][15] ), 
        .CO(\CARRYB[44][14] ), .S(\SUMB[44][14] ) );
  FA_X1 S2_44_15 ( .A(\ab[44][15] ), .B(\CARRYB[43][15] ), .CI(\SUMB[43][16] ), 
        .CO(\CARRYB[44][15] ), .S(\SUMB[44][15] ) );
  FA_X1 S2_44_16 ( .A(\ab[44][16] ), .B(\CARRYB[43][16] ), .CI(\SUMB[43][17] ), 
        .CO(\CARRYB[44][16] ), .S(\SUMB[44][16] ) );
  FA_X1 S2_44_17 ( .A(\ab[44][17] ), .B(\CARRYB[43][17] ), .CI(\SUMB[43][18] ), 
        .CO(\CARRYB[44][17] ), .S(\SUMB[44][17] ) );
  FA_X1 S2_44_18 ( .A(\ab[44][18] ), .B(\CARRYB[43][18] ), .CI(\SUMB[43][19] ), 
        .CO(\CARRYB[44][18] ), .S(\SUMB[44][18] ) );
  FA_X1 S2_44_19 ( .A(\ab[44][19] ), .B(\CARRYB[43][19] ), .CI(\SUMB[43][20] ), 
        .CO(\CARRYB[44][19] ), .S(\SUMB[44][19] ) );
  FA_X1 S2_44_20 ( .A(\ab[44][20] ), .B(\CARRYB[43][20] ), .CI(\SUMB[43][21] ), 
        .CO(\CARRYB[44][20] ), .S(\SUMB[44][20] ) );
  FA_X1 S2_44_21 ( .A(\ab[44][21] ), .B(\CARRYB[43][21] ), .CI(\SUMB[43][22] ), 
        .CO(\CARRYB[44][21] ), .S(\SUMB[44][21] ) );
  FA_X1 S2_44_22 ( .A(\ab[44][22] ), .B(\CARRYB[43][22] ), .CI(\SUMB[43][23] ), 
        .CO(\CARRYB[44][22] ), .S(\SUMB[44][22] ) );
  FA_X1 S2_44_23 ( .A(\ab[44][23] ), .B(\CARRYB[43][23] ), .CI(\SUMB[43][24] ), 
        .CO(\CARRYB[44][23] ), .S(\SUMB[44][23] ) );
  FA_X1 S2_44_24 ( .A(\ab[44][24] ), .B(\CARRYB[43][24] ), .CI(\SUMB[43][25] ), 
        .CO(\CARRYB[44][24] ), .S(\SUMB[44][24] ) );
  FA_X1 S2_44_25 ( .A(\ab[44][25] ), .B(\CARRYB[43][25] ), .CI(\SUMB[43][26] ), 
        .CO(\CARRYB[44][25] ), .S(\SUMB[44][25] ) );
  FA_X1 S2_44_26 ( .A(\ab[44][26] ), .B(\CARRYB[43][26] ), .CI(\SUMB[43][27] ), 
        .CO(\CARRYB[44][26] ), .S(\SUMB[44][26] ) );
  FA_X1 S2_44_27 ( .A(\ab[44][27] ), .B(\CARRYB[43][27] ), .CI(\SUMB[43][28] ), 
        .CO(\CARRYB[44][27] ), .S(\SUMB[44][27] ) );
  FA_X1 S2_44_28 ( .A(\ab[44][28] ), .B(\CARRYB[43][28] ), .CI(\SUMB[43][29] ), 
        .CO(\CARRYB[44][28] ), .S(\SUMB[44][28] ) );
  FA_X1 S2_44_29 ( .A(\ab[44][29] ), .B(\CARRYB[43][29] ), .CI(\SUMB[43][30] ), 
        .CO(\CARRYB[44][29] ), .S(\SUMB[44][29] ) );
  FA_X1 S2_44_30 ( .A(\ab[44][30] ), .B(\CARRYB[43][30] ), .CI(\SUMB[43][31] ), 
        .CO(\CARRYB[44][30] ), .S(\SUMB[44][30] ) );
  FA_X1 S2_44_31 ( .A(\ab[44][31] ), .B(\CARRYB[43][31] ), .CI(\SUMB[43][32] ), 
        .CO(\CARRYB[44][31] ), .S(\SUMB[44][31] ) );
  FA_X1 S2_44_32 ( .A(\ab[44][32] ), .B(\CARRYB[43][32] ), .CI(\SUMB[43][33] ), 
        .CO(\CARRYB[44][32] ), .S(\SUMB[44][32] ) );
  FA_X1 S2_44_33 ( .A(\ab[44][33] ), .B(\CARRYB[43][33] ), .CI(\SUMB[43][34] ), 
        .CO(\CARRYB[44][33] ), .S(\SUMB[44][33] ) );
  FA_X1 S2_44_34 ( .A(\ab[44][34] ), .B(\CARRYB[43][34] ), .CI(\SUMB[43][35] ), 
        .CO(\CARRYB[44][34] ), .S(\SUMB[44][34] ) );
  FA_X1 S2_44_35 ( .A(\ab[44][35] ), .B(\CARRYB[43][35] ), .CI(\SUMB[43][36] ), 
        .CO(\CARRYB[44][35] ), .S(\SUMB[44][35] ) );
  FA_X1 S2_44_36 ( .A(\ab[44][36] ), .B(\CARRYB[43][36] ), .CI(\SUMB[43][37] ), 
        .CO(\CARRYB[44][36] ), .S(\SUMB[44][36] ) );
  FA_X1 S2_44_37 ( .A(\ab[44][37] ), .B(\CARRYB[43][37] ), .CI(\SUMB[43][38] ), 
        .CO(\CARRYB[44][37] ), .S(\SUMB[44][37] ) );
  FA_X1 S2_44_38 ( .A(\ab[44][38] ), .B(\CARRYB[43][38] ), .CI(\SUMB[43][39] ), 
        .CO(\CARRYB[44][38] ), .S(\SUMB[44][38] ) );
  FA_X1 S2_44_39 ( .A(\ab[44][39] ), .B(\CARRYB[43][39] ), .CI(\SUMB[43][40] ), 
        .CO(\CARRYB[44][39] ), .S(\SUMB[44][39] ) );
  FA_X1 S2_44_40 ( .A(\ab[44][40] ), .B(\CARRYB[43][40] ), .CI(\SUMB[43][41] ), 
        .CO(\CARRYB[44][40] ), .S(\SUMB[44][40] ) );
  FA_X1 S2_44_41 ( .A(\ab[44][41] ), .B(\CARRYB[43][41] ), .CI(\SUMB[43][42] ), 
        .CO(\CARRYB[44][41] ), .S(\SUMB[44][41] ) );
  FA_X1 S2_44_42 ( .A(\ab[44][42] ), .B(\CARRYB[43][42] ), .CI(\SUMB[43][43] ), 
        .CO(\CARRYB[44][42] ), .S(\SUMB[44][42] ) );
  FA_X1 S2_44_43 ( .A(\ab[44][43] ), .B(\CARRYB[43][43] ), .CI(\SUMB[43][44] ), 
        .CO(\CARRYB[44][43] ), .S(\SUMB[44][43] ) );
  FA_X1 S2_44_44 ( .A(\ab[44][44] ), .B(\CARRYB[43][44] ), .CI(\SUMB[43][45] ), 
        .CO(\CARRYB[44][44] ), .S(\SUMB[44][44] ) );
  FA_X1 S2_44_45 ( .A(\ab[44][45] ), .B(\CARRYB[43][45] ), .CI(\SUMB[43][46] ), 
        .CO(\CARRYB[44][45] ), .S(\SUMB[44][45] ) );
  FA_X1 S2_44_46 ( .A(\ab[44][46] ), .B(\CARRYB[43][46] ), .CI(\SUMB[43][47] ), 
        .CO(\CARRYB[44][46] ), .S(\SUMB[44][46] ) );
  FA_X1 S2_44_47 ( .A(\ab[44][47] ), .B(\CARRYB[43][47] ), .CI(\SUMB[43][48] ), 
        .CO(\CARRYB[44][47] ), .S(\SUMB[44][47] ) );
  FA_X1 S2_44_48 ( .A(\ab[44][48] ), .B(\CARRYB[43][48] ), .CI(\SUMB[43][49] ), 
        .CO(\CARRYB[44][48] ), .S(\SUMB[44][48] ) );
  FA_X1 S2_44_49 ( .A(\ab[44][49] ), .B(\CARRYB[43][49] ), .CI(\SUMB[43][50] ), 
        .CO(\CARRYB[44][49] ), .S(\SUMB[44][49] ) );
  FA_X1 S2_44_50 ( .A(\ab[44][50] ), .B(\CARRYB[43][50] ), .CI(\SUMB[43][51] ), 
        .CO(\CARRYB[44][50] ), .S(\SUMB[44][50] ) );
  FA_X1 S3_44_51 ( .A(\ab[44][51] ), .B(\CARRYB[43][51] ), .CI(\ab[43][52] ), 
        .CO(\CARRYB[44][51] ), .S(\SUMB[44][51] ) );
  FA_X1 S1_43_0 ( .A(\ab[43][0] ), .B(\CARRYB[42][0] ), .CI(\SUMB[42][1] ), 
        .CO(\CARRYB[43][0] ), .S(CLA_SUM[43]) );
  FA_X1 S2_43_1 ( .A(\ab[43][1] ), .B(\CARRYB[42][1] ), .CI(\SUMB[42][2] ), 
        .CO(\CARRYB[43][1] ), .S(\SUMB[43][1] ) );
  FA_X1 S2_43_2 ( .A(\ab[43][2] ), .B(\CARRYB[42][2] ), .CI(\SUMB[42][3] ), 
        .CO(\CARRYB[43][2] ), .S(\SUMB[43][2] ) );
  FA_X1 S2_43_3 ( .A(\ab[43][3] ), .B(\CARRYB[42][3] ), .CI(\SUMB[42][4] ), 
        .CO(\CARRYB[43][3] ), .S(\SUMB[43][3] ) );
  FA_X1 S2_43_4 ( .A(\ab[43][4] ), .B(\CARRYB[42][4] ), .CI(\SUMB[42][5] ), 
        .CO(\CARRYB[43][4] ), .S(\SUMB[43][4] ) );
  FA_X1 S2_43_5 ( .A(\ab[43][5] ), .B(\CARRYB[42][5] ), .CI(\SUMB[42][6] ), 
        .CO(\CARRYB[43][5] ), .S(\SUMB[43][5] ) );
  FA_X1 S2_43_6 ( .A(\ab[43][6] ), .B(\CARRYB[42][6] ), .CI(\SUMB[42][7] ), 
        .CO(\CARRYB[43][6] ), .S(\SUMB[43][6] ) );
  FA_X1 S2_43_7 ( .A(\ab[43][7] ), .B(\CARRYB[42][7] ), .CI(\SUMB[42][8] ), 
        .CO(\CARRYB[43][7] ), .S(\SUMB[43][7] ) );
  FA_X1 S2_43_8 ( .A(\ab[43][8] ), .B(\CARRYB[42][8] ), .CI(\SUMB[42][9] ), 
        .CO(\CARRYB[43][8] ), .S(\SUMB[43][8] ) );
  FA_X1 S2_43_9 ( .A(\ab[43][9] ), .B(\CARRYB[42][9] ), .CI(\SUMB[42][10] ), 
        .CO(\CARRYB[43][9] ), .S(\SUMB[43][9] ) );
  FA_X1 S2_43_10 ( .A(\ab[43][10] ), .B(\CARRYB[42][10] ), .CI(\SUMB[42][11] ), 
        .CO(\CARRYB[43][10] ), .S(\SUMB[43][10] ) );
  FA_X1 S2_43_11 ( .A(\ab[43][11] ), .B(\CARRYB[42][11] ), .CI(\SUMB[42][12] ), 
        .CO(\CARRYB[43][11] ), .S(\SUMB[43][11] ) );
  FA_X1 S2_43_12 ( .A(\ab[43][12] ), .B(\CARRYB[42][12] ), .CI(\SUMB[42][13] ), 
        .CO(\CARRYB[43][12] ), .S(\SUMB[43][12] ) );
  FA_X1 S2_43_13 ( .A(\ab[43][13] ), .B(\CARRYB[42][13] ), .CI(\SUMB[42][14] ), 
        .CO(\CARRYB[43][13] ), .S(\SUMB[43][13] ) );
  FA_X1 S2_43_14 ( .A(\ab[43][14] ), .B(\CARRYB[42][14] ), .CI(\SUMB[42][15] ), 
        .CO(\CARRYB[43][14] ), .S(\SUMB[43][14] ) );
  FA_X1 S2_43_15 ( .A(\ab[43][15] ), .B(\CARRYB[42][15] ), .CI(\SUMB[42][16] ), 
        .CO(\CARRYB[43][15] ), .S(\SUMB[43][15] ) );
  FA_X1 S2_43_16 ( .A(\ab[43][16] ), .B(\CARRYB[42][16] ), .CI(\SUMB[42][17] ), 
        .CO(\CARRYB[43][16] ), .S(\SUMB[43][16] ) );
  FA_X1 S2_43_17 ( .A(\ab[43][17] ), .B(\CARRYB[42][17] ), .CI(\SUMB[42][18] ), 
        .CO(\CARRYB[43][17] ), .S(\SUMB[43][17] ) );
  FA_X1 S2_43_18 ( .A(\ab[43][18] ), .B(\CARRYB[42][18] ), .CI(\SUMB[42][19] ), 
        .CO(\CARRYB[43][18] ), .S(\SUMB[43][18] ) );
  FA_X1 S2_43_19 ( .A(\ab[43][19] ), .B(\CARRYB[42][19] ), .CI(\SUMB[42][20] ), 
        .CO(\CARRYB[43][19] ), .S(\SUMB[43][19] ) );
  FA_X1 S2_43_20 ( .A(\ab[43][20] ), .B(\CARRYB[42][20] ), .CI(\SUMB[42][21] ), 
        .CO(\CARRYB[43][20] ), .S(\SUMB[43][20] ) );
  FA_X1 S2_43_21 ( .A(\ab[43][21] ), .B(\CARRYB[42][21] ), .CI(\SUMB[42][22] ), 
        .CO(\CARRYB[43][21] ), .S(\SUMB[43][21] ) );
  FA_X1 S2_43_22 ( .A(\ab[43][22] ), .B(\CARRYB[42][22] ), .CI(\SUMB[42][23] ), 
        .CO(\CARRYB[43][22] ), .S(\SUMB[43][22] ) );
  FA_X1 S2_43_23 ( .A(\ab[43][23] ), .B(\CARRYB[42][23] ), .CI(\SUMB[42][24] ), 
        .CO(\CARRYB[43][23] ), .S(\SUMB[43][23] ) );
  FA_X1 S2_43_24 ( .A(\ab[43][24] ), .B(\CARRYB[42][24] ), .CI(\SUMB[42][25] ), 
        .CO(\CARRYB[43][24] ), .S(\SUMB[43][24] ) );
  FA_X1 S2_43_25 ( .A(\ab[43][25] ), .B(\CARRYB[42][25] ), .CI(\SUMB[42][26] ), 
        .CO(\CARRYB[43][25] ), .S(\SUMB[43][25] ) );
  FA_X1 S2_43_26 ( .A(\ab[43][26] ), .B(\CARRYB[42][26] ), .CI(\SUMB[42][27] ), 
        .CO(\CARRYB[43][26] ), .S(\SUMB[43][26] ) );
  FA_X1 S2_43_27 ( .A(\ab[43][27] ), .B(\CARRYB[42][27] ), .CI(\SUMB[42][28] ), 
        .CO(\CARRYB[43][27] ), .S(\SUMB[43][27] ) );
  FA_X1 S2_43_28 ( .A(\ab[43][28] ), .B(\CARRYB[42][28] ), .CI(\SUMB[42][29] ), 
        .CO(\CARRYB[43][28] ), .S(\SUMB[43][28] ) );
  FA_X1 S2_43_29 ( .A(\ab[43][29] ), .B(\CARRYB[42][29] ), .CI(\SUMB[42][30] ), 
        .CO(\CARRYB[43][29] ), .S(\SUMB[43][29] ) );
  FA_X1 S2_43_30 ( .A(\ab[43][30] ), .B(\CARRYB[42][30] ), .CI(\SUMB[42][31] ), 
        .CO(\CARRYB[43][30] ), .S(\SUMB[43][30] ) );
  FA_X1 S2_43_31 ( .A(\ab[43][31] ), .B(\CARRYB[42][31] ), .CI(\SUMB[42][32] ), 
        .CO(\CARRYB[43][31] ), .S(\SUMB[43][31] ) );
  FA_X1 S2_43_32 ( .A(\ab[43][32] ), .B(\CARRYB[42][32] ), .CI(\SUMB[42][33] ), 
        .CO(\CARRYB[43][32] ), .S(\SUMB[43][32] ) );
  FA_X1 S2_43_33 ( .A(\ab[43][33] ), .B(\CARRYB[42][33] ), .CI(\SUMB[42][34] ), 
        .CO(\CARRYB[43][33] ), .S(\SUMB[43][33] ) );
  FA_X1 S2_43_34 ( .A(\ab[43][34] ), .B(\CARRYB[42][34] ), .CI(\SUMB[42][35] ), 
        .CO(\CARRYB[43][34] ), .S(\SUMB[43][34] ) );
  FA_X1 S2_43_35 ( .A(\ab[43][35] ), .B(\CARRYB[42][35] ), .CI(\SUMB[42][36] ), 
        .CO(\CARRYB[43][35] ), .S(\SUMB[43][35] ) );
  FA_X1 S2_43_36 ( .A(\ab[43][36] ), .B(\CARRYB[42][36] ), .CI(\SUMB[42][37] ), 
        .CO(\CARRYB[43][36] ), .S(\SUMB[43][36] ) );
  FA_X1 S2_43_37 ( .A(\ab[43][37] ), .B(\CARRYB[42][37] ), .CI(\SUMB[42][38] ), 
        .CO(\CARRYB[43][37] ), .S(\SUMB[43][37] ) );
  FA_X1 S2_43_38 ( .A(\ab[43][38] ), .B(\CARRYB[42][38] ), .CI(\SUMB[42][39] ), 
        .CO(\CARRYB[43][38] ), .S(\SUMB[43][38] ) );
  FA_X1 S2_43_39 ( .A(\ab[43][39] ), .B(\CARRYB[42][39] ), .CI(\SUMB[42][40] ), 
        .CO(\CARRYB[43][39] ), .S(\SUMB[43][39] ) );
  FA_X1 S2_43_40 ( .A(\ab[43][40] ), .B(\CARRYB[42][40] ), .CI(\SUMB[42][41] ), 
        .CO(\CARRYB[43][40] ), .S(\SUMB[43][40] ) );
  FA_X1 S2_43_41 ( .A(\ab[43][41] ), .B(\CARRYB[42][41] ), .CI(\SUMB[42][42] ), 
        .CO(\CARRYB[43][41] ), .S(\SUMB[43][41] ) );
  FA_X1 S2_43_42 ( .A(\ab[43][42] ), .B(\CARRYB[42][42] ), .CI(\SUMB[42][43] ), 
        .CO(\CARRYB[43][42] ), .S(\SUMB[43][42] ) );
  FA_X1 S2_43_43 ( .A(\ab[43][43] ), .B(\CARRYB[42][43] ), .CI(\SUMB[42][44] ), 
        .CO(\CARRYB[43][43] ), .S(\SUMB[43][43] ) );
  FA_X1 S2_43_44 ( .A(\ab[43][44] ), .B(\CARRYB[42][44] ), .CI(\SUMB[42][45] ), 
        .CO(\CARRYB[43][44] ), .S(\SUMB[43][44] ) );
  FA_X1 S2_43_45 ( .A(\ab[43][45] ), .B(\CARRYB[42][45] ), .CI(\SUMB[42][46] ), 
        .CO(\CARRYB[43][45] ), .S(\SUMB[43][45] ) );
  FA_X1 S2_43_46 ( .A(\ab[43][46] ), .B(\CARRYB[42][46] ), .CI(\SUMB[42][47] ), 
        .CO(\CARRYB[43][46] ), .S(\SUMB[43][46] ) );
  FA_X1 S2_43_47 ( .A(\ab[43][47] ), .B(\CARRYB[42][47] ), .CI(\SUMB[42][48] ), 
        .CO(\CARRYB[43][47] ), .S(\SUMB[43][47] ) );
  FA_X1 S2_43_48 ( .A(\ab[43][48] ), .B(\CARRYB[42][48] ), .CI(\SUMB[42][49] ), 
        .CO(\CARRYB[43][48] ), .S(\SUMB[43][48] ) );
  FA_X1 S2_43_49 ( .A(\ab[43][49] ), .B(\CARRYB[42][49] ), .CI(\SUMB[42][50] ), 
        .CO(\CARRYB[43][49] ), .S(\SUMB[43][49] ) );
  FA_X1 S2_43_50 ( .A(\ab[43][50] ), .B(\CARRYB[42][50] ), .CI(\SUMB[42][51] ), 
        .CO(\CARRYB[43][50] ), .S(\SUMB[43][50] ) );
  FA_X1 S3_43_51 ( .A(\ab[43][51] ), .B(\CARRYB[42][51] ), .CI(\ab[42][52] ), 
        .CO(\CARRYB[43][51] ), .S(\SUMB[43][51] ) );
  FA_X1 S1_42_0 ( .A(\ab[42][0] ), .B(\CARRYB[41][0] ), .CI(\SUMB[41][1] ), 
        .CO(\CARRYB[42][0] ), .S(CLA_SUM[42]) );
  FA_X1 S2_42_1 ( .A(\ab[42][1] ), .B(\CARRYB[41][1] ), .CI(\SUMB[41][2] ), 
        .CO(\CARRYB[42][1] ), .S(\SUMB[42][1] ) );
  FA_X1 S2_42_2 ( .A(\ab[42][2] ), .B(\CARRYB[41][2] ), .CI(\SUMB[41][3] ), 
        .CO(\CARRYB[42][2] ), .S(\SUMB[42][2] ) );
  FA_X1 S2_42_3 ( .A(\ab[42][3] ), .B(\CARRYB[41][3] ), .CI(\SUMB[41][4] ), 
        .CO(\CARRYB[42][3] ), .S(\SUMB[42][3] ) );
  FA_X1 S2_42_4 ( .A(\ab[42][4] ), .B(\CARRYB[41][4] ), .CI(\SUMB[41][5] ), 
        .CO(\CARRYB[42][4] ), .S(\SUMB[42][4] ) );
  FA_X1 S2_42_5 ( .A(\ab[42][5] ), .B(\CARRYB[41][5] ), .CI(\SUMB[41][6] ), 
        .CO(\CARRYB[42][5] ), .S(\SUMB[42][5] ) );
  FA_X1 S2_42_6 ( .A(\ab[42][6] ), .B(\CARRYB[41][6] ), .CI(\SUMB[41][7] ), 
        .CO(\CARRYB[42][6] ), .S(\SUMB[42][6] ) );
  FA_X1 S2_42_7 ( .A(\ab[42][7] ), .B(\CARRYB[41][7] ), .CI(\SUMB[41][8] ), 
        .CO(\CARRYB[42][7] ), .S(\SUMB[42][7] ) );
  FA_X1 S2_42_8 ( .A(\ab[42][8] ), .B(\CARRYB[41][8] ), .CI(\SUMB[41][9] ), 
        .CO(\CARRYB[42][8] ), .S(\SUMB[42][8] ) );
  FA_X1 S2_42_9 ( .A(\ab[42][9] ), .B(\CARRYB[41][9] ), .CI(\SUMB[41][10] ), 
        .CO(\CARRYB[42][9] ), .S(\SUMB[42][9] ) );
  FA_X1 S2_42_10 ( .A(\ab[42][10] ), .B(\CARRYB[41][10] ), .CI(\SUMB[41][11] ), 
        .CO(\CARRYB[42][10] ), .S(\SUMB[42][10] ) );
  FA_X1 S2_42_11 ( .A(\ab[42][11] ), .B(\CARRYB[41][11] ), .CI(\SUMB[41][12] ), 
        .CO(\CARRYB[42][11] ), .S(\SUMB[42][11] ) );
  FA_X1 S2_42_12 ( .A(\ab[42][12] ), .B(\CARRYB[41][12] ), .CI(\SUMB[41][13] ), 
        .CO(\CARRYB[42][12] ), .S(\SUMB[42][12] ) );
  FA_X1 S2_42_13 ( .A(\ab[42][13] ), .B(\CARRYB[41][13] ), .CI(\SUMB[41][14] ), 
        .CO(\CARRYB[42][13] ), .S(\SUMB[42][13] ) );
  FA_X1 S2_42_14 ( .A(\ab[42][14] ), .B(\CARRYB[41][14] ), .CI(\SUMB[41][15] ), 
        .CO(\CARRYB[42][14] ), .S(\SUMB[42][14] ) );
  FA_X1 S2_42_15 ( .A(\ab[42][15] ), .B(\CARRYB[41][15] ), .CI(\SUMB[41][16] ), 
        .CO(\CARRYB[42][15] ), .S(\SUMB[42][15] ) );
  FA_X1 S2_42_16 ( .A(\ab[42][16] ), .B(\CARRYB[41][16] ), .CI(\SUMB[41][17] ), 
        .CO(\CARRYB[42][16] ), .S(\SUMB[42][16] ) );
  FA_X1 S2_42_17 ( .A(\ab[42][17] ), .B(\CARRYB[41][17] ), .CI(\SUMB[41][18] ), 
        .CO(\CARRYB[42][17] ), .S(\SUMB[42][17] ) );
  FA_X1 S2_42_18 ( .A(\ab[42][18] ), .B(\CARRYB[41][18] ), .CI(\SUMB[41][19] ), 
        .CO(\CARRYB[42][18] ), .S(\SUMB[42][18] ) );
  FA_X1 S2_42_19 ( .A(\ab[42][19] ), .B(\CARRYB[41][19] ), .CI(\SUMB[41][20] ), 
        .CO(\CARRYB[42][19] ), .S(\SUMB[42][19] ) );
  FA_X1 S2_42_20 ( .A(\ab[42][20] ), .B(\CARRYB[41][20] ), .CI(\SUMB[41][21] ), 
        .CO(\CARRYB[42][20] ), .S(\SUMB[42][20] ) );
  FA_X1 S2_42_21 ( .A(\ab[42][21] ), .B(\CARRYB[41][21] ), .CI(\SUMB[41][22] ), 
        .CO(\CARRYB[42][21] ), .S(\SUMB[42][21] ) );
  FA_X1 S2_42_22 ( .A(\ab[42][22] ), .B(\CARRYB[41][22] ), .CI(\SUMB[41][23] ), 
        .CO(\CARRYB[42][22] ), .S(\SUMB[42][22] ) );
  FA_X1 S2_42_23 ( .A(\ab[42][23] ), .B(\CARRYB[41][23] ), .CI(\SUMB[41][24] ), 
        .CO(\CARRYB[42][23] ), .S(\SUMB[42][23] ) );
  FA_X1 S2_42_24 ( .A(\ab[42][24] ), .B(\CARRYB[41][24] ), .CI(\SUMB[41][25] ), 
        .CO(\CARRYB[42][24] ), .S(\SUMB[42][24] ) );
  FA_X1 S2_42_25 ( .A(\ab[42][25] ), .B(\CARRYB[41][25] ), .CI(\SUMB[41][26] ), 
        .CO(\CARRYB[42][25] ), .S(\SUMB[42][25] ) );
  FA_X1 S2_42_26 ( .A(\ab[42][26] ), .B(\CARRYB[41][26] ), .CI(\SUMB[41][27] ), 
        .CO(\CARRYB[42][26] ), .S(\SUMB[42][26] ) );
  FA_X1 S2_42_27 ( .A(\ab[42][27] ), .B(\CARRYB[41][27] ), .CI(\SUMB[41][28] ), 
        .CO(\CARRYB[42][27] ), .S(\SUMB[42][27] ) );
  FA_X1 S2_42_28 ( .A(\ab[42][28] ), .B(\CARRYB[41][28] ), .CI(\SUMB[41][29] ), 
        .CO(\CARRYB[42][28] ), .S(\SUMB[42][28] ) );
  FA_X1 S2_42_29 ( .A(\ab[42][29] ), .B(\CARRYB[41][29] ), .CI(\SUMB[41][30] ), 
        .CO(\CARRYB[42][29] ), .S(\SUMB[42][29] ) );
  FA_X1 S2_42_30 ( .A(\ab[42][30] ), .B(\CARRYB[41][30] ), .CI(\SUMB[41][31] ), 
        .CO(\CARRYB[42][30] ), .S(\SUMB[42][30] ) );
  FA_X1 S2_42_31 ( .A(\ab[42][31] ), .B(\CARRYB[41][31] ), .CI(\SUMB[41][32] ), 
        .CO(\CARRYB[42][31] ), .S(\SUMB[42][31] ) );
  FA_X1 S2_42_32 ( .A(\ab[42][32] ), .B(\CARRYB[41][32] ), .CI(\SUMB[41][33] ), 
        .CO(\CARRYB[42][32] ), .S(\SUMB[42][32] ) );
  FA_X1 S2_42_33 ( .A(\ab[42][33] ), .B(\CARRYB[41][33] ), .CI(\SUMB[41][34] ), 
        .CO(\CARRYB[42][33] ), .S(\SUMB[42][33] ) );
  FA_X1 S2_42_34 ( .A(\ab[42][34] ), .B(\CARRYB[41][34] ), .CI(\SUMB[41][35] ), 
        .CO(\CARRYB[42][34] ), .S(\SUMB[42][34] ) );
  FA_X1 S2_42_35 ( .A(\ab[42][35] ), .B(\CARRYB[41][35] ), .CI(\SUMB[41][36] ), 
        .CO(\CARRYB[42][35] ), .S(\SUMB[42][35] ) );
  FA_X1 S2_42_36 ( .A(\ab[42][36] ), .B(\CARRYB[41][36] ), .CI(\SUMB[41][37] ), 
        .CO(\CARRYB[42][36] ), .S(\SUMB[42][36] ) );
  FA_X1 S2_42_37 ( .A(\ab[42][37] ), .B(\CARRYB[41][37] ), .CI(\SUMB[41][38] ), 
        .CO(\CARRYB[42][37] ), .S(\SUMB[42][37] ) );
  FA_X1 S2_42_38 ( .A(\ab[42][38] ), .B(\CARRYB[41][38] ), .CI(\SUMB[41][39] ), 
        .CO(\CARRYB[42][38] ), .S(\SUMB[42][38] ) );
  FA_X1 S2_42_39 ( .A(\ab[42][39] ), .B(\CARRYB[41][39] ), .CI(\SUMB[41][40] ), 
        .CO(\CARRYB[42][39] ), .S(\SUMB[42][39] ) );
  FA_X1 S2_42_40 ( .A(\ab[42][40] ), .B(\CARRYB[41][40] ), .CI(\SUMB[41][41] ), 
        .CO(\CARRYB[42][40] ), .S(\SUMB[42][40] ) );
  FA_X1 S2_42_41 ( .A(\ab[42][41] ), .B(\CARRYB[41][41] ), .CI(\SUMB[41][42] ), 
        .CO(\CARRYB[42][41] ), .S(\SUMB[42][41] ) );
  FA_X1 S2_42_42 ( .A(\ab[42][42] ), .B(\CARRYB[41][42] ), .CI(\SUMB[41][43] ), 
        .CO(\CARRYB[42][42] ), .S(\SUMB[42][42] ) );
  FA_X1 S2_42_43 ( .A(\ab[42][43] ), .B(\CARRYB[41][43] ), .CI(\SUMB[41][44] ), 
        .CO(\CARRYB[42][43] ), .S(\SUMB[42][43] ) );
  FA_X1 S2_42_44 ( .A(\ab[42][44] ), .B(\CARRYB[41][44] ), .CI(\SUMB[41][45] ), 
        .CO(\CARRYB[42][44] ), .S(\SUMB[42][44] ) );
  FA_X1 S2_42_45 ( .A(\ab[42][45] ), .B(\CARRYB[41][45] ), .CI(\SUMB[41][46] ), 
        .CO(\CARRYB[42][45] ), .S(\SUMB[42][45] ) );
  FA_X1 S2_42_46 ( .A(\ab[42][46] ), .B(\CARRYB[41][46] ), .CI(\SUMB[41][47] ), 
        .CO(\CARRYB[42][46] ), .S(\SUMB[42][46] ) );
  FA_X1 S2_42_47 ( .A(\ab[42][47] ), .B(\CARRYB[41][47] ), .CI(\SUMB[41][48] ), 
        .CO(\CARRYB[42][47] ), .S(\SUMB[42][47] ) );
  FA_X1 S2_42_48 ( .A(\ab[42][48] ), .B(\CARRYB[41][48] ), .CI(\SUMB[41][49] ), 
        .CO(\CARRYB[42][48] ), .S(\SUMB[42][48] ) );
  FA_X1 S2_42_49 ( .A(\ab[42][49] ), .B(\CARRYB[41][49] ), .CI(\SUMB[41][50] ), 
        .CO(\CARRYB[42][49] ), .S(\SUMB[42][49] ) );
  FA_X1 S2_42_50 ( .A(\ab[42][50] ), .B(\CARRYB[41][50] ), .CI(\SUMB[41][51] ), 
        .CO(\CARRYB[42][50] ), .S(\SUMB[42][50] ) );
  FA_X1 S3_42_51 ( .A(\ab[42][51] ), .B(\CARRYB[41][51] ), .CI(\ab[41][52] ), 
        .CO(\CARRYB[42][51] ), .S(\SUMB[42][51] ) );
  FA_X1 S1_41_0 ( .A(\ab[41][0] ), .B(\CARRYB[40][0] ), .CI(\SUMB[40][1] ), 
        .CO(\CARRYB[41][0] ), .S(CLA_SUM[41]) );
  FA_X1 S2_41_1 ( .A(\ab[41][1] ), .B(\CARRYB[40][1] ), .CI(\SUMB[40][2] ), 
        .CO(\CARRYB[41][1] ), .S(\SUMB[41][1] ) );
  FA_X1 S2_41_2 ( .A(\ab[41][2] ), .B(\CARRYB[40][2] ), .CI(\SUMB[40][3] ), 
        .CO(\CARRYB[41][2] ), .S(\SUMB[41][2] ) );
  FA_X1 S2_41_3 ( .A(\ab[41][3] ), .B(\CARRYB[40][3] ), .CI(\SUMB[40][4] ), 
        .CO(\CARRYB[41][3] ), .S(\SUMB[41][3] ) );
  FA_X1 S2_41_4 ( .A(\ab[41][4] ), .B(\CARRYB[40][4] ), .CI(\SUMB[40][5] ), 
        .CO(\CARRYB[41][4] ), .S(\SUMB[41][4] ) );
  FA_X1 S2_41_5 ( .A(\ab[41][5] ), .B(\CARRYB[40][5] ), .CI(\SUMB[40][6] ), 
        .CO(\CARRYB[41][5] ), .S(\SUMB[41][5] ) );
  FA_X1 S2_41_6 ( .A(\ab[41][6] ), .B(\CARRYB[40][6] ), .CI(\SUMB[40][7] ), 
        .CO(\CARRYB[41][6] ), .S(\SUMB[41][6] ) );
  FA_X1 S2_41_7 ( .A(\ab[41][7] ), .B(\CARRYB[40][7] ), .CI(\SUMB[40][8] ), 
        .CO(\CARRYB[41][7] ), .S(\SUMB[41][7] ) );
  FA_X1 S2_41_8 ( .A(\ab[41][8] ), .B(\CARRYB[40][8] ), .CI(\SUMB[40][9] ), 
        .CO(\CARRYB[41][8] ), .S(\SUMB[41][8] ) );
  FA_X1 S2_41_9 ( .A(\ab[41][9] ), .B(\CARRYB[40][9] ), .CI(\SUMB[40][10] ), 
        .CO(\CARRYB[41][9] ), .S(\SUMB[41][9] ) );
  FA_X1 S2_41_10 ( .A(\ab[41][10] ), .B(\CARRYB[40][10] ), .CI(\SUMB[40][11] ), 
        .CO(\CARRYB[41][10] ), .S(\SUMB[41][10] ) );
  FA_X1 S2_41_11 ( .A(\ab[41][11] ), .B(\CARRYB[40][11] ), .CI(\SUMB[40][12] ), 
        .CO(\CARRYB[41][11] ), .S(\SUMB[41][11] ) );
  FA_X1 S2_41_12 ( .A(\ab[41][12] ), .B(\CARRYB[40][12] ), .CI(\SUMB[40][13] ), 
        .CO(\CARRYB[41][12] ), .S(\SUMB[41][12] ) );
  FA_X1 S2_41_13 ( .A(\ab[41][13] ), .B(\CARRYB[40][13] ), .CI(\SUMB[40][14] ), 
        .CO(\CARRYB[41][13] ), .S(\SUMB[41][13] ) );
  FA_X1 S2_41_14 ( .A(\ab[41][14] ), .B(\CARRYB[40][14] ), .CI(\SUMB[40][15] ), 
        .CO(\CARRYB[41][14] ), .S(\SUMB[41][14] ) );
  FA_X1 S2_41_15 ( .A(\ab[41][15] ), .B(\CARRYB[40][15] ), .CI(\SUMB[40][16] ), 
        .CO(\CARRYB[41][15] ), .S(\SUMB[41][15] ) );
  FA_X1 S2_41_16 ( .A(\ab[41][16] ), .B(\CARRYB[40][16] ), .CI(\SUMB[40][17] ), 
        .CO(\CARRYB[41][16] ), .S(\SUMB[41][16] ) );
  FA_X1 S2_41_17 ( .A(\ab[41][17] ), .B(\CARRYB[40][17] ), .CI(\SUMB[40][18] ), 
        .CO(\CARRYB[41][17] ), .S(\SUMB[41][17] ) );
  FA_X1 S2_41_18 ( .A(\ab[41][18] ), .B(\CARRYB[40][18] ), .CI(\SUMB[40][19] ), 
        .CO(\CARRYB[41][18] ), .S(\SUMB[41][18] ) );
  FA_X1 S2_41_19 ( .A(\ab[41][19] ), .B(\CARRYB[40][19] ), .CI(\SUMB[40][20] ), 
        .CO(\CARRYB[41][19] ), .S(\SUMB[41][19] ) );
  FA_X1 S2_41_20 ( .A(\ab[41][20] ), .B(\CARRYB[40][20] ), .CI(\SUMB[40][21] ), 
        .CO(\CARRYB[41][20] ), .S(\SUMB[41][20] ) );
  FA_X1 S2_41_21 ( .A(\ab[41][21] ), .B(\CARRYB[40][21] ), .CI(\SUMB[40][22] ), 
        .CO(\CARRYB[41][21] ), .S(\SUMB[41][21] ) );
  FA_X1 S2_41_22 ( .A(\ab[41][22] ), .B(\CARRYB[40][22] ), .CI(\SUMB[40][23] ), 
        .CO(\CARRYB[41][22] ), .S(\SUMB[41][22] ) );
  FA_X1 S2_41_23 ( .A(\ab[41][23] ), .B(\CARRYB[40][23] ), .CI(\SUMB[40][24] ), 
        .CO(\CARRYB[41][23] ), .S(\SUMB[41][23] ) );
  FA_X1 S2_41_24 ( .A(\ab[41][24] ), .B(\CARRYB[40][24] ), .CI(\SUMB[40][25] ), 
        .CO(\CARRYB[41][24] ), .S(\SUMB[41][24] ) );
  FA_X1 S2_41_25 ( .A(\ab[41][25] ), .B(\CARRYB[40][25] ), .CI(\SUMB[40][26] ), 
        .CO(\CARRYB[41][25] ), .S(\SUMB[41][25] ) );
  FA_X1 S2_41_26 ( .A(\ab[41][26] ), .B(\CARRYB[40][26] ), .CI(\SUMB[40][27] ), 
        .CO(\CARRYB[41][26] ), .S(\SUMB[41][26] ) );
  FA_X1 S2_41_27 ( .A(\ab[41][27] ), .B(\CARRYB[40][27] ), .CI(\SUMB[40][28] ), 
        .CO(\CARRYB[41][27] ), .S(\SUMB[41][27] ) );
  FA_X1 S2_41_28 ( .A(\ab[41][28] ), .B(\CARRYB[40][28] ), .CI(\SUMB[40][29] ), 
        .CO(\CARRYB[41][28] ), .S(\SUMB[41][28] ) );
  FA_X1 S2_41_29 ( .A(\ab[41][29] ), .B(\CARRYB[40][29] ), .CI(\SUMB[40][30] ), 
        .CO(\CARRYB[41][29] ), .S(\SUMB[41][29] ) );
  FA_X1 S2_41_30 ( .A(\ab[41][30] ), .B(\CARRYB[40][30] ), .CI(\SUMB[40][31] ), 
        .CO(\CARRYB[41][30] ), .S(\SUMB[41][30] ) );
  FA_X1 S2_41_31 ( .A(\ab[41][31] ), .B(\CARRYB[40][31] ), .CI(\SUMB[40][32] ), 
        .CO(\CARRYB[41][31] ), .S(\SUMB[41][31] ) );
  FA_X1 S2_41_32 ( .A(\ab[41][32] ), .B(\CARRYB[40][32] ), .CI(\SUMB[40][33] ), 
        .CO(\CARRYB[41][32] ), .S(\SUMB[41][32] ) );
  FA_X1 S2_41_33 ( .A(\ab[41][33] ), .B(\CARRYB[40][33] ), .CI(\SUMB[40][34] ), 
        .CO(\CARRYB[41][33] ), .S(\SUMB[41][33] ) );
  FA_X1 S2_41_34 ( .A(\ab[41][34] ), .B(\CARRYB[40][34] ), .CI(\SUMB[40][35] ), 
        .CO(\CARRYB[41][34] ), .S(\SUMB[41][34] ) );
  FA_X1 S2_41_35 ( .A(\ab[41][35] ), .B(\CARRYB[40][35] ), .CI(\SUMB[40][36] ), 
        .CO(\CARRYB[41][35] ), .S(\SUMB[41][35] ) );
  FA_X1 S2_41_36 ( .A(\ab[41][36] ), .B(\CARRYB[40][36] ), .CI(\SUMB[40][37] ), 
        .CO(\CARRYB[41][36] ), .S(\SUMB[41][36] ) );
  FA_X1 S2_41_37 ( .A(\ab[41][37] ), .B(\CARRYB[40][37] ), .CI(\SUMB[40][38] ), 
        .CO(\CARRYB[41][37] ), .S(\SUMB[41][37] ) );
  FA_X1 S2_41_38 ( .A(\ab[41][38] ), .B(\CARRYB[40][38] ), .CI(\SUMB[40][39] ), 
        .CO(\CARRYB[41][38] ), .S(\SUMB[41][38] ) );
  FA_X1 S2_41_39 ( .A(\ab[41][39] ), .B(\CARRYB[40][39] ), .CI(\SUMB[40][40] ), 
        .CO(\CARRYB[41][39] ), .S(\SUMB[41][39] ) );
  FA_X1 S2_41_40 ( .A(\ab[41][40] ), .B(\CARRYB[40][40] ), .CI(\SUMB[40][41] ), 
        .CO(\CARRYB[41][40] ), .S(\SUMB[41][40] ) );
  FA_X1 S2_41_41 ( .A(\ab[41][41] ), .B(\CARRYB[40][41] ), .CI(\SUMB[40][42] ), 
        .CO(\CARRYB[41][41] ), .S(\SUMB[41][41] ) );
  FA_X1 S2_41_42 ( .A(\ab[41][42] ), .B(\CARRYB[40][42] ), .CI(\SUMB[40][43] ), 
        .CO(\CARRYB[41][42] ), .S(\SUMB[41][42] ) );
  FA_X1 S2_41_43 ( .A(\ab[41][43] ), .B(\CARRYB[40][43] ), .CI(\SUMB[40][44] ), 
        .CO(\CARRYB[41][43] ), .S(\SUMB[41][43] ) );
  FA_X1 S2_41_44 ( .A(\ab[41][44] ), .B(\CARRYB[40][44] ), .CI(\SUMB[40][45] ), 
        .CO(\CARRYB[41][44] ), .S(\SUMB[41][44] ) );
  FA_X1 S2_41_45 ( .A(\ab[41][45] ), .B(\CARRYB[40][45] ), .CI(\SUMB[40][46] ), 
        .CO(\CARRYB[41][45] ), .S(\SUMB[41][45] ) );
  FA_X1 S2_41_46 ( .A(\ab[41][46] ), .B(\CARRYB[40][46] ), .CI(\SUMB[40][47] ), 
        .CO(\CARRYB[41][46] ), .S(\SUMB[41][46] ) );
  FA_X1 S2_41_47 ( .A(\ab[41][47] ), .B(\CARRYB[40][47] ), .CI(\SUMB[40][48] ), 
        .CO(\CARRYB[41][47] ), .S(\SUMB[41][47] ) );
  FA_X1 S2_41_48 ( .A(\ab[41][48] ), .B(\CARRYB[40][48] ), .CI(\SUMB[40][49] ), 
        .CO(\CARRYB[41][48] ), .S(\SUMB[41][48] ) );
  FA_X1 S2_41_49 ( .A(\ab[41][49] ), .B(\CARRYB[40][49] ), .CI(\SUMB[40][50] ), 
        .CO(\CARRYB[41][49] ), .S(\SUMB[41][49] ) );
  FA_X1 S2_41_50 ( .A(\ab[41][50] ), .B(\CARRYB[40][50] ), .CI(\SUMB[40][51] ), 
        .CO(\CARRYB[41][50] ), .S(\SUMB[41][50] ) );
  FA_X1 S3_41_51 ( .A(\ab[41][51] ), .B(\CARRYB[40][51] ), .CI(\ab[40][52] ), 
        .CO(\CARRYB[41][51] ), .S(\SUMB[41][51] ) );
  FA_X1 S1_40_0 ( .A(\ab[40][0] ), .B(\CARRYB[39][0] ), .CI(\SUMB[39][1] ), 
        .CO(\CARRYB[40][0] ), .S(CLA_SUM[40]) );
  FA_X1 S2_40_1 ( .A(\ab[40][1] ), .B(\CARRYB[39][1] ), .CI(\SUMB[39][2] ), 
        .CO(\CARRYB[40][1] ), .S(\SUMB[40][1] ) );
  FA_X1 S2_40_2 ( .A(\ab[40][2] ), .B(\CARRYB[39][2] ), .CI(\SUMB[39][3] ), 
        .CO(\CARRYB[40][2] ), .S(\SUMB[40][2] ) );
  FA_X1 S2_40_3 ( .A(\ab[40][3] ), .B(\CARRYB[39][3] ), .CI(\SUMB[39][4] ), 
        .CO(\CARRYB[40][3] ), .S(\SUMB[40][3] ) );
  FA_X1 S2_40_4 ( .A(\ab[40][4] ), .B(\CARRYB[39][4] ), .CI(\SUMB[39][5] ), 
        .CO(\CARRYB[40][4] ), .S(\SUMB[40][4] ) );
  FA_X1 S2_40_5 ( .A(\ab[40][5] ), .B(\CARRYB[39][5] ), .CI(\SUMB[39][6] ), 
        .CO(\CARRYB[40][5] ), .S(\SUMB[40][5] ) );
  FA_X1 S2_40_6 ( .A(\ab[40][6] ), .B(\CARRYB[39][6] ), .CI(\SUMB[39][7] ), 
        .CO(\CARRYB[40][6] ), .S(\SUMB[40][6] ) );
  FA_X1 S2_40_7 ( .A(\ab[40][7] ), .B(\CARRYB[39][7] ), .CI(\SUMB[39][8] ), 
        .CO(\CARRYB[40][7] ), .S(\SUMB[40][7] ) );
  FA_X1 S2_40_8 ( .A(\ab[40][8] ), .B(\CARRYB[39][8] ), .CI(\SUMB[39][9] ), 
        .CO(\CARRYB[40][8] ), .S(\SUMB[40][8] ) );
  FA_X1 S2_40_9 ( .A(\ab[40][9] ), .B(\CARRYB[39][9] ), .CI(\SUMB[39][10] ), 
        .CO(\CARRYB[40][9] ), .S(\SUMB[40][9] ) );
  FA_X1 S2_40_10 ( .A(\ab[40][10] ), .B(\CARRYB[39][10] ), .CI(\SUMB[39][11] ), 
        .CO(\CARRYB[40][10] ), .S(\SUMB[40][10] ) );
  FA_X1 S2_40_11 ( .A(\ab[40][11] ), .B(\CARRYB[39][11] ), .CI(\SUMB[39][12] ), 
        .CO(\CARRYB[40][11] ), .S(\SUMB[40][11] ) );
  FA_X1 S2_40_12 ( .A(\ab[40][12] ), .B(\CARRYB[39][12] ), .CI(\SUMB[39][13] ), 
        .CO(\CARRYB[40][12] ), .S(\SUMB[40][12] ) );
  FA_X1 S2_40_13 ( .A(\ab[40][13] ), .B(\CARRYB[39][13] ), .CI(\SUMB[39][14] ), 
        .CO(\CARRYB[40][13] ), .S(\SUMB[40][13] ) );
  FA_X1 S2_40_14 ( .A(\ab[40][14] ), .B(\CARRYB[39][14] ), .CI(\SUMB[39][15] ), 
        .CO(\CARRYB[40][14] ), .S(\SUMB[40][14] ) );
  FA_X1 S2_40_15 ( .A(\ab[40][15] ), .B(\CARRYB[39][15] ), .CI(\SUMB[39][16] ), 
        .CO(\CARRYB[40][15] ), .S(\SUMB[40][15] ) );
  FA_X1 S2_40_16 ( .A(\ab[40][16] ), .B(\CARRYB[39][16] ), .CI(\SUMB[39][17] ), 
        .CO(\CARRYB[40][16] ), .S(\SUMB[40][16] ) );
  FA_X1 S2_40_17 ( .A(\ab[40][17] ), .B(\CARRYB[39][17] ), .CI(\SUMB[39][18] ), 
        .CO(\CARRYB[40][17] ), .S(\SUMB[40][17] ) );
  FA_X1 S2_40_18 ( .A(\ab[40][18] ), .B(\CARRYB[39][18] ), .CI(\SUMB[39][19] ), 
        .CO(\CARRYB[40][18] ), .S(\SUMB[40][18] ) );
  FA_X1 S2_40_19 ( .A(\ab[40][19] ), .B(\CARRYB[39][19] ), .CI(\SUMB[39][20] ), 
        .CO(\CARRYB[40][19] ), .S(\SUMB[40][19] ) );
  FA_X1 S2_40_20 ( .A(\ab[40][20] ), .B(\CARRYB[39][20] ), .CI(\SUMB[39][21] ), 
        .CO(\CARRYB[40][20] ), .S(\SUMB[40][20] ) );
  FA_X1 S2_40_21 ( .A(\ab[40][21] ), .B(\CARRYB[39][21] ), .CI(\SUMB[39][22] ), 
        .CO(\CARRYB[40][21] ), .S(\SUMB[40][21] ) );
  FA_X1 S2_40_22 ( .A(\ab[40][22] ), .B(\CARRYB[39][22] ), .CI(\SUMB[39][23] ), 
        .CO(\CARRYB[40][22] ), .S(\SUMB[40][22] ) );
  FA_X1 S2_40_23 ( .A(\ab[40][23] ), .B(\CARRYB[39][23] ), .CI(\SUMB[39][24] ), 
        .CO(\CARRYB[40][23] ), .S(\SUMB[40][23] ) );
  FA_X1 S2_40_24 ( .A(\ab[40][24] ), .B(\CARRYB[39][24] ), .CI(\SUMB[39][25] ), 
        .CO(\CARRYB[40][24] ), .S(\SUMB[40][24] ) );
  FA_X1 S2_40_25 ( .A(\ab[40][25] ), .B(\CARRYB[39][25] ), .CI(\SUMB[39][26] ), 
        .CO(\CARRYB[40][25] ), .S(\SUMB[40][25] ) );
  FA_X1 S2_40_26 ( .A(\ab[40][26] ), .B(\CARRYB[39][26] ), .CI(\SUMB[39][27] ), 
        .CO(\CARRYB[40][26] ), .S(\SUMB[40][26] ) );
  FA_X1 S2_40_27 ( .A(\ab[40][27] ), .B(\CARRYB[39][27] ), .CI(\SUMB[39][28] ), 
        .CO(\CARRYB[40][27] ), .S(\SUMB[40][27] ) );
  FA_X1 S2_40_28 ( .A(\ab[40][28] ), .B(\CARRYB[39][28] ), .CI(\SUMB[39][29] ), 
        .CO(\CARRYB[40][28] ), .S(\SUMB[40][28] ) );
  FA_X1 S2_40_29 ( .A(\ab[40][29] ), .B(\CARRYB[39][29] ), .CI(\SUMB[39][30] ), 
        .CO(\CARRYB[40][29] ), .S(\SUMB[40][29] ) );
  FA_X1 S2_40_30 ( .A(\ab[40][30] ), .B(\CARRYB[39][30] ), .CI(\SUMB[39][31] ), 
        .CO(\CARRYB[40][30] ), .S(\SUMB[40][30] ) );
  FA_X1 S2_40_31 ( .A(\ab[40][31] ), .B(\CARRYB[39][31] ), .CI(\SUMB[39][32] ), 
        .CO(\CARRYB[40][31] ), .S(\SUMB[40][31] ) );
  FA_X1 S2_40_32 ( .A(\ab[40][32] ), .B(\CARRYB[39][32] ), .CI(\SUMB[39][33] ), 
        .CO(\CARRYB[40][32] ), .S(\SUMB[40][32] ) );
  FA_X1 S2_40_33 ( .A(\ab[40][33] ), .B(\CARRYB[39][33] ), .CI(\SUMB[39][34] ), 
        .CO(\CARRYB[40][33] ), .S(\SUMB[40][33] ) );
  FA_X1 S2_40_34 ( .A(\ab[40][34] ), .B(\CARRYB[39][34] ), .CI(\SUMB[39][35] ), 
        .CO(\CARRYB[40][34] ), .S(\SUMB[40][34] ) );
  FA_X1 S2_40_35 ( .A(\ab[40][35] ), .B(\CARRYB[39][35] ), .CI(\SUMB[39][36] ), 
        .CO(\CARRYB[40][35] ), .S(\SUMB[40][35] ) );
  FA_X1 S2_40_36 ( .A(\ab[40][36] ), .B(\CARRYB[39][36] ), .CI(\SUMB[39][37] ), 
        .CO(\CARRYB[40][36] ), .S(\SUMB[40][36] ) );
  FA_X1 S2_40_37 ( .A(\ab[40][37] ), .B(\CARRYB[39][37] ), .CI(\SUMB[39][38] ), 
        .CO(\CARRYB[40][37] ), .S(\SUMB[40][37] ) );
  FA_X1 S2_40_38 ( .A(\ab[40][38] ), .B(\CARRYB[39][38] ), .CI(\SUMB[39][39] ), 
        .CO(\CARRYB[40][38] ), .S(\SUMB[40][38] ) );
  FA_X1 S2_40_39 ( .A(\ab[40][39] ), .B(\CARRYB[39][39] ), .CI(\SUMB[39][40] ), 
        .CO(\CARRYB[40][39] ), .S(\SUMB[40][39] ) );
  FA_X1 S2_40_40 ( .A(\ab[40][40] ), .B(\CARRYB[39][40] ), .CI(\SUMB[39][41] ), 
        .CO(\CARRYB[40][40] ), .S(\SUMB[40][40] ) );
  FA_X1 S2_40_41 ( .A(\ab[40][41] ), .B(\CARRYB[39][41] ), .CI(\SUMB[39][42] ), 
        .CO(\CARRYB[40][41] ), .S(\SUMB[40][41] ) );
  FA_X1 S2_40_42 ( .A(\ab[40][42] ), .B(\CARRYB[39][42] ), .CI(\SUMB[39][43] ), 
        .CO(\CARRYB[40][42] ), .S(\SUMB[40][42] ) );
  FA_X1 S2_40_43 ( .A(\ab[40][43] ), .B(\CARRYB[39][43] ), .CI(\SUMB[39][44] ), 
        .CO(\CARRYB[40][43] ), .S(\SUMB[40][43] ) );
  FA_X1 S2_40_44 ( .A(\ab[40][44] ), .B(\CARRYB[39][44] ), .CI(\SUMB[39][45] ), 
        .CO(\CARRYB[40][44] ), .S(\SUMB[40][44] ) );
  FA_X1 S2_40_45 ( .A(\ab[40][45] ), .B(\CARRYB[39][45] ), .CI(\SUMB[39][46] ), 
        .CO(\CARRYB[40][45] ), .S(\SUMB[40][45] ) );
  FA_X1 S2_40_46 ( .A(\ab[40][46] ), .B(\CARRYB[39][46] ), .CI(\SUMB[39][47] ), 
        .CO(\CARRYB[40][46] ), .S(\SUMB[40][46] ) );
  FA_X1 S2_40_47 ( .A(\ab[40][47] ), .B(\CARRYB[39][47] ), .CI(\SUMB[39][48] ), 
        .CO(\CARRYB[40][47] ), .S(\SUMB[40][47] ) );
  FA_X1 S2_40_48 ( .A(\ab[40][48] ), .B(\CARRYB[39][48] ), .CI(\SUMB[39][49] ), 
        .CO(\CARRYB[40][48] ), .S(\SUMB[40][48] ) );
  FA_X1 S2_40_49 ( .A(\ab[40][49] ), .B(\CARRYB[39][49] ), .CI(\SUMB[39][50] ), 
        .CO(\CARRYB[40][49] ), .S(\SUMB[40][49] ) );
  FA_X1 S2_40_50 ( .A(\ab[40][50] ), .B(\CARRYB[39][50] ), .CI(\SUMB[39][51] ), 
        .CO(\CARRYB[40][50] ), .S(\SUMB[40][50] ) );
  FA_X1 S3_40_51 ( .A(\ab[40][51] ), .B(\CARRYB[39][51] ), .CI(\ab[39][52] ), 
        .CO(\CARRYB[40][51] ), .S(\SUMB[40][51] ) );
  FA_X1 S1_39_0 ( .A(\ab[39][0] ), .B(\CARRYB[38][0] ), .CI(\SUMB[38][1] ), 
        .CO(\CARRYB[39][0] ), .S(CLA_SUM[39]) );
  FA_X1 S2_39_1 ( .A(\ab[39][1] ), .B(\CARRYB[38][1] ), .CI(\SUMB[38][2] ), 
        .CO(\CARRYB[39][1] ), .S(\SUMB[39][1] ) );
  FA_X1 S2_39_2 ( .A(\ab[39][2] ), .B(\CARRYB[38][2] ), .CI(\SUMB[38][3] ), 
        .CO(\CARRYB[39][2] ), .S(\SUMB[39][2] ) );
  FA_X1 S2_39_3 ( .A(\ab[39][3] ), .B(\CARRYB[38][3] ), .CI(\SUMB[38][4] ), 
        .CO(\CARRYB[39][3] ), .S(\SUMB[39][3] ) );
  FA_X1 S2_39_4 ( .A(\ab[39][4] ), .B(\CARRYB[38][4] ), .CI(\SUMB[38][5] ), 
        .CO(\CARRYB[39][4] ), .S(\SUMB[39][4] ) );
  FA_X1 S2_39_5 ( .A(\ab[39][5] ), .B(\CARRYB[38][5] ), .CI(\SUMB[38][6] ), 
        .CO(\CARRYB[39][5] ), .S(\SUMB[39][5] ) );
  FA_X1 S2_39_6 ( .A(\ab[39][6] ), .B(\CARRYB[38][6] ), .CI(\SUMB[38][7] ), 
        .CO(\CARRYB[39][6] ), .S(\SUMB[39][6] ) );
  FA_X1 S2_39_7 ( .A(\ab[39][7] ), .B(\CARRYB[38][7] ), .CI(\SUMB[38][8] ), 
        .CO(\CARRYB[39][7] ), .S(\SUMB[39][7] ) );
  FA_X1 S2_39_8 ( .A(\ab[39][8] ), .B(\CARRYB[38][8] ), .CI(\SUMB[38][9] ), 
        .CO(\CARRYB[39][8] ), .S(\SUMB[39][8] ) );
  FA_X1 S2_39_9 ( .A(\ab[39][9] ), .B(\CARRYB[38][9] ), .CI(\SUMB[38][10] ), 
        .CO(\CARRYB[39][9] ), .S(\SUMB[39][9] ) );
  FA_X1 S2_39_10 ( .A(\ab[39][10] ), .B(\CARRYB[38][10] ), .CI(\SUMB[38][11] ), 
        .CO(\CARRYB[39][10] ), .S(\SUMB[39][10] ) );
  FA_X1 S2_39_11 ( .A(\ab[39][11] ), .B(\CARRYB[38][11] ), .CI(\SUMB[38][12] ), 
        .CO(\CARRYB[39][11] ), .S(\SUMB[39][11] ) );
  FA_X1 S2_39_12 ( .A(\ab[39][12] ), .B(\CARRYB[38][12] ), .CI(\SUMB[38][13] ), 
        .CO(\CARRYB[39][12] ), .S(\SUMB[39][12] ) );
  FA_X1 S2_39_13 ( .A(\ab[39][13] ), .B(\CARRYB[38][13] ), .CI(\SUMB[38][14] ), 
        .CO(\CARRYB[39][13] ), .S(\SUMB[39][13] ) );
  FA_X1 S2_39_14 ( .A(\ab[39][14] ), .B(\CARRYB[38][14] ), .CI(\SUMB[38][15] ), 
        .CO(\CARRYB[39][14] ), .S(\SUMB[39][14] ) );
  FA_X1 S2_39_15 ( .A(\ab[39][15] ), .B(\CARRYB[38][15] ), .CI(\SUMB[38][16] ), 
        .CO(\CARRYB[39][15] ), .S(\SUMB[39][15] ) );
  FA_X1 S2_39_16 ( .A(\ab[39][16] ), .B(\CARRYB[38][16] ), .CI(\SUMB[38][17] ), 
        .CO(\CARRYB[39][16] ), .S(\SUMB[39][16] ) );
  FA_X1 S2_39_17 ( .A(\ab[39][17] ), .B(\CARRYB[38][17] ), .CI(\SUMB[38][18] ), 
        .CO(\CARRYB[39][17] ), .S(\SUMB[39][17] ) );
  FA_X1 S2_39_18 ( .A(\ab[39][18] ), .B(\CARRYB[38][18] ), .CI(\SUMB[38][19] ), 
        .CO(\CARRYB[39][18] ), .S(\SUMB[39][18] ) );
  FA_X1 S2_39_19 ( .A(\ab[39][19] ), .B(\CARRYB[38][19] ), .CI(\SUMB[38][20] ), 
        .CO(\CARRYB[39][19] ), .S(\SUMB[39][19] ) );
  FA_X1 S2_39_20 ( .A(\ab[39][20] ), .B(\CARRYB[38][20] ), .CI(\SUMB[38][21] ), 
        .CO(\CARRYB[39][20] ), .S(\SUMB[39][20] ) );
  FA_X1 S2_39_21 ( .A(\ab[39][21] ), .B(\CARRYB[38][21] ), .CI(\SUMB[38][22] ), 
        .CO(\CARRYB[39][21] ), .S(\SUMB[39][21] ) );
  FA_X1 S2_39_22 ( .A(\ab[39][22] ), .B(\CARRYB[38][22] ), .CI(\SUMB[38][23] ), 
        .CO(\CARRYB[39][22] ), .S(\SUMB[39][22] ) );
  FA_X1 S2_39_23 ( .A(\ab[39][23] ), .B(\CARRYB[38][23] ), .CI(\SUMB[38][24] ), 
        .CO(\CARRYB[39][23] ), .S(\SUMB[39][23] ) );
  FA_X1 S2_39_24 ( .A(\ab[39][24] ), .B(\CARRYB[38][24] ), .CI(\SUMB[38][25] ), 
        .CO(\CARRYB[39][24] ), .S(\SUMB[39][24] ) );
  FA_X1 S2_39_25 ( .A(\ab[39][25] ), .B(\CARRYB[38][25] ), .CI(\SUMB[38][26] ), 
        .CO(\CARRYB[39][25] ), .S(\SUMB[39][25] ) );
  FA_X1 S2_39_26 ( .A(\ab[39][26] ), .B(\CARRYB[38][26] ), .CI(\SUMB[38][27] ), 
        .CO(\CARRYB[39][26] ), .S(\SUMB[39][26] ) );
  FA_X1 S2_39_27 ( .A(\ab[39][27] ), .B(\CARRYB[38][27] ), .CI(\SUMB[38][28] ), 
        .CO(\CARRYB[39][27] ), .S(\SUMB[39][27] ) );
  FA_X1 S2_39_28 ( .A(\ab[39][28] ), .B(\CARRYB[38][28] ), .CI(\SUMB[38][29] ), 
        .CO(\CARRYB[39][28] ), .S(\SUMB[39][28] ) );
  FA_X1 S2_39_29 ( .A(\ab[39][29] ), .B(\CARRYB[38][29] ), .CI(\SUMB[38][30] ), 
        .CO(\CARRYB[39][29] ), .S(\SUMB[39][29] ) );
  FA_X1 S2_39_30 ( .A(\ab[39][30] ), .B(\CARRYB[38][30] ), .CI(\SUMB[38][31] ), 
        .CO(\CARRYB[39][30] ), .S(\SUMB[39][30] ) );
  FA_X1 S2_39_31 ( .A(\ab[39][31] ), .B(\CARRYB[38][31] ), .CI(\SUMB[38][32] ), 
        .CO(\CARRYB[39][31] ), .S(\SUMB[39][31] ) );
  FA_X1 S2_39_32 ( .A(\ab[39][32] ), .B(\CARRYB[38][32] ), .CI(\SUMB[38][33] ), 
        .CO(\CARRYB[39][32] ), .S(\SUMB[39][32] ) );
  FA_X1 S2_39_33 ( .A(\ab[39][33] ), .B(\CARRYB[38][33] ), .CI(\SUMB[38][34] ), 
        .CO(\CARRYB[39][33] ), .S(\SUMB[39][33] ) );
  FA_X1 S2_39_34 ( .A(\ab[39][34] ), .B(\CARRYB[38][34] ), .CI(\SUMB[38][35] ), 
        .CO(\CARRYB[39][34] ), .S(\SUMB[39][34] ) );
  FA_X1 S2_39_35 ( .A(\ab[39][35] ), .B(\CARRYB[38][35] ), .CI(\SUMB[38][36] ), 
        .CO(\CARRYB[39][35] ), .S(\SUMB[39][35] ) );
  FA_X1 S2_39_36 ( .A(\ab[39][36] ), .B(\CARRYB[38][36] ), .CI(\SUMB[38][37] ), 
        .CO(\CARRYB[39][36] ), .S(\SUMB[39][36] ) );
  FA_X1 S2_39_37 ( .A(\ab[39][37] ), .B(\CARRYB[38][37] ), .CI(\SUMB[38][38] ), 
        .CO(\CARRYB[39][37] ), .S(\SUMB[39][37] ) );
  FA_X1 S2_39_38 ( .A(\ab[39][38] ), .B(\CARRYB[38][38] ), .CI(\SUMB[38][39] ), 
        .CO(\CARRYB[39][38] ), .S(\SUMB[39][38] ) );
  FA_X1 S2_39_39 ( .A(\ab[39][39] ), .B(\CARRYB[38][39] ), .CI(\SUMB[38][40] ), 
        .CO(\CARRYB[39][39] ), .S(\SUMB[39][39] ) );
  FA_X1 S2_39_40 ( .A(\ab[39][40] ), .B(\CARRYB[38][40] ), .CI(\SUMB[38][41] ), 
        .CO(\CARRYB[39][40] ), .S(\SUMB[39][40] ) );
  FA_X1 S2_39_41 ( .A(\ab[39][41] ), .B(\CARRYB[38][41] ), .CI(\SUMB[38][42] ), 
        .CO(\CARRYB[39][41] ), .S(\SUMB[39][41] ) );
  FA_X1 S2_39_42 ( .A(\ab[39][42] ), .B(\CARRYB[38][42] ), .CI(\SUMB[38][43] ), 
        .CO(\CARRYB[39][42] ), .S(\SUMB[39][42] ) );
  FA_X1 S2_39_43 ( .A(\ab[39][43] ), .B(\CARRYB[38][43] ), .CI(\SUMB[38][44] ), 
        .CO(\CARRYB[39][43] ), .S(\SUMB[39][43] ) );
  FA_X1 S2_39_44 ( .A(\ab[39][44] ), .B(\CARRYB[38][44] ), .CI(\SUMB[38][45] ), 
        .CO(\CARRYB[39][44] ), .S(\SUMB[39][44] ) );
  FA_X1 S2_39_45 ( .A(\ab[39][45] ), .B(\CARRYB[38][45] ), .CI(\SUMB[38][46] ), 
        .CO(\CARRYB[39][45] ), .S(\SUMB[39][45] ) );
  FA_X1 S2_39_46 ( .A(\ab[39][46] ), .B(\CARRYB[38][46] ), .CI(\SUMB[38][47] ), 
        .CO(\CARRYB[39][46] ), .S(\SUMB[39][46] ) );
  FA_X1 S2_39_47 ( .A(\ab[39][47] ), .B(\CARRYB[38][47] ), .CI(\SUMB[38][48] ), 
        .CO(\CARRYB[39][47] ), .S(\SUMB[39][47] ) );
  FA_X1 S2_39_48 ( .A(\ab[39][48] ), .B(\CARRYB[38][48] ), .CI(\SUMB[38][49] ), 
        .CO(\CARRYB[39][48] ), .S(\SUMB[39][48] ) );
  FA_X1 S2_39_49 ( .A(\ab[39][49] ), .B(\CARRYB[38][49] ), .CI(\SUMB[38][50] ), 
        .CO(\CARRYB[39][49] ), .S(\SUMB[39][49] ) );
  FA_X1 S2_39_50 ( .A(\ab[39][50] ), .B(\CARRYB[38][50] ), .CI(\SUMB[38][51] ), 
        .CO(\CARRYB[39][50] ), .S(\SUMB[39][50] ) );
  FA_X1 S3_39_51 ( .A(\ab[39][51] ), .B(\CARRYB[38][51] ), .CI(\ab[38][52] ), 
        .CO(\CARRYB[39][51] ), .S(\SUMB[39][51] ) );
  FA_X1 S1_38_0 ( .A(\ab[38][0] ), .B(\CARRYB[37][0] ), .CI(\SUMB[37][1] ), 
        .CO(\CARRYB[38][0] ), .S(CLA_SUM[38]) );
  FA_X1 S2_38_1 ( .A(\ab[38][1] ), .B(\CARRYB[37][1] ), .CI(\SUMB[37][2] ), 
        .CO(\CARRYB[38][1] ), .S(\SUMB[38][1] ) );
  FA_X1 S2_38_2 ( .A(\ab[38][2] ), .B(\CARRYB[37][2] ), .CI(\SUMB[37][3] ), 
        .CO(\CARRYB[38][2] ), .S(\SUMB[38][2] ) );
  FA_X1 S2_38_3 ( .A(\ab[38][3] ), .B(\CARRYB[37][3] ), .CI(\SUMB[37][4] ), 
        .CO(\CARRYB[38][3] ), .S(\SUMB[38][3] ) );
  FA_X1 S2_38_4 ( .A(\ab[38][4] ), .B(\CARRYB[37][4] ), .CI(\SUMB[37][5] ), 
        .CO(\CARRYB[38][4] ), .S(\SUMB[38][4] ) );
  FA_X1 S2_38_5 ( .A(\ab[38][5] ), .B(\CARRYB[37][5] ), .CI(\SUMB[37][6] ), 
        .CO(\CARRYB[38][5] ), .S(\SUMB[38][5] ) );
  FA_X1 S2_38_6 ( .A(\ab[38][6] ), .B(\CARRYB[37][6] ), .CI(\SUMB[37][7] ), 
        .CO(\CARRYB[38][6] ), .S(\SUMB[38][6] ) );
  FA_X1 S2_38_7 ( .A(\ab[38][7] ), .B(\CARRYB[37][7] ), .CI(\SUMB[37][8] ), 
        .CO(\CARRYB[38][7] ), .S(\SUMB[38][7] ) );
  FA_X1 S2_38_8 ( .A(\ab[38][8] ), .B(\CARRYB[37][8] ), .CI(\SUMB[37][9] ), 
        .CO(\CARRYB[38][8] ), .S(\SUMB[38][8] ) );
  FA_X1 S2_38_9 ( .A(\ab[38][9] ), .B(\CARRYB[37][9] ), .CI(\SUMB[37][10] ), 
        .CO(\CARRYB[38][9] ), .S(\SUMB[38][9] ) );
  FA_X1 S2_38_10 ( .A(\ab[38][10] ), .B(\CARRYB[37][10] ), .CI(\SUMB[37][11] ), 
        .CO(\CARRYB[38][10] ), .S(\SUMB[38][10] ) );
  FA_X1 S2_38_11 ( .A(\ab[38][11] ), .B(\CARRYB[37][11] ), .CI(\SUMB[37][12] ), 
        .CO(\CARRYB[38][11] ), .S(\SUMB[38][11] ) );
  FA_X1 S2_38_12 ( .A(\ab[38][12] ), .B(\CARRYB[37][12] ), .CI(\SUMB[37][13] ), 
        .CO(\CARRYB[38][12] ), .S(\SUMB[38][12] ) );
  FA_X1 S2_38_13 ( .A(\ab[38][13] ), .B(\CARRYB[37][13] ), .CI(\SUMB[37][14] ), 
        .CO(\CARRYB[38][13] ), .S(\SUMB[38][13] ) );
  FA_X1 S2_38_14 ( .A(\ab[38][14] ), .B(\CARRYB[37][14] ), .CI(\SUMB[37][15] ), 
        .CO(\CARRYB[38][14] ), .S(\SUMB[38][14] ) );
  FA_X1 S2_38_15 ( .A(\ab[38][15] ), .B(\CARRYB[37][15] ), .CI(\SUMB[37][16] ), 
        .CO(\CARRYB[38][15] ), .S(\SUMB[38][15] ) );
  FA_X1 S2_38_16 ( .A(\ab[38][16] ), .B(\CARRYB[37][16] ), .CI(\SUMB[37][17] ), 
        .CO(\CARRYB[38][16] ), .S(\SUMB[38][16] ) );
  FA_X1 S2_38_17 ( .A(\ab[38][17] ), .B(\CARRYB[37][17] ), .CI(\SUMB[37][18] ), 
        .CO(\CARRYB[38][17] ), .S(\SUMB[38][17] ) );
  FA_X1 S2_38_18 ( .A(\ab[38][18] ), .B(\CARRYB[37][18] ), .CI(\SUMB[37][19] ), 
        .CO(\CARRYB[38][18] ), .S(\SUMB[38][18] ) );
  FA_X1 S2_38_19 ( .A(\ab[38][19] ), .B(\CARRYB[37][19] ), .CI(\SUMB[37][20] ), 
        .CO(\CARRYB[38][19] ), .S(\SUMB[38][19] ) );
  FA_X1 S2_38_20 ( .A(\ab[38][20] ), .B(\CARRYB[37][20] ), .CI(\SUMB[37][21] ), 
        .CO(\CARRYB[38][20] ), .S(\SUMB[38][20] ) );
  FA_X1 S2_38_21 ( .A(\ab[38][21] ), .B(\CARRYB[37][21] ), .CI(\SUMB[37][22] ), 
        .CO(\CARRYB[38][21] ), .S(\SUMB[38][21] ) );
  FA_X1 S2_38_22 ( .A(\ab[38][22] ), .B(\CARRYB[37][22] ), .CI(\SUMB[37][23] ), 
        .CO(\CARRYB[38][22] ), .S(\SUMB[38][22] ) );
  FA_X1 S2_38_23 ( .A(\ab[38][23] ), .B(\CARRYB[37][23] ), .CI(\SUMB[37][24] ), 
        .CO(\CARRYB[38][23] ), .S(\SUMB[38][23] ) );
  FA_X1 S2_38_24 ( .A(\ab[38][24] ), .B(\CARRYB[37][24] ), .CI(\SUMB[37][25] ), 
        .CO(\CARRYB[38][24] ), .S(\SUMB[38][24] ) );
  FA_X1 S2_38_25 ( .A(\ab[38][25] ), .B(\CARRYB[37][25] ), .CI(\SUMB[37][26] ), 
        .CO(\CARRYB[38][25] ), .S(\SUMB[38][25] ) );
  FA_X1 S2_38_26 ( .A(\ab[38][26] ), .B(\CARRYB[37][26] ), .CI(\SUMB[37][27] ), 
        .CO(\CARRYB[38][26] ), .S(\SUMB[38][26] ) );
  FA_X1 S2_38_27 ( .A(\ab[38][27] ), .B(\CARRYB[37][27] ), .CI(\SUMB[37][28] ), 
        .CO(\CARRYB[38][27] ), .S(\SUMB[38][27] ) );
  FA_X1 S2_38_28 ( .A(\ab[38][28] ), .B(\CARRYB[37][28] ), .CI(\SUMB[37][29] ), 
        .CO(\CARRYB[38][28] ), .S(\SUMB[38][28] ) );
  FA_X1 S2_38_29 ( .A(\ab[38][29] ), .B(\CARRYB[37][29] ), .CI(\SUMB[37][30] ), 
        .CO(\CARRYB[38][29] ), .S(\SUMB[38][29] ) );
  FA_X1 S2_38_30 ( .A(\ab[38][30] ), .B(\CARRYB[37][30] ), .CI(\SUMB[37][31] ), 
        .CO(\CARRYB[38][30] ), .S(\SUMB[38][30] ) );
  FA_X1 S2_38_31 ( .A(\ab[38][31] ), .B(\CARRYB[37][31] ), .CI(\SUMB[37][32] ), 
        .CO(\CARRYB[38][31] ), .S(\SUMB[38][31] ) );
  FA_X1 S2_38_32 ( .A(\ab[38][32] ), .B(\CARRYB[37][32] ), .CI(\SUMB[37][33] ), 
        .CO(\CARRYB[38][32] ), .S(\SUMB[38][32] ) );
  FA_X1 S2_38_33 ( .A(\ab[38][33] ), .B(\CARRYB[37][33] ), .CI(\SUMB[37][34] ), 
        .CO(\CARRYB[38][33] ), .S(\SUMB[38][33] ) );
  FA_X1 S2_38_34 ( .A(\ab[38][34] ), .B(\CARRYB[37][34] ), .CI(\SUMB[37][35] ), 
        .CO(\CARRYB[38][34] ), .S(\SUMB[38][34] ) );
  FA_X1 S2_38_35 ( .A(\ab[38][35] ), .B(\CARRYB[37][35] ), .CI(\SUMB[37][36] ), 
        .CO(\CARRYB[38][35] ), .S(\SUMB[38][35] ) );
  FA_X1 S2_38_36 ( .A(\ab[38][36] ), .B(\CARRYB[37][36] ), .CI(\SUMB[37][37] ), 
        .CO(\CARRYB[38][36] ), .S(\SUMB[38][36] ) );
  FA_X1 S2_38_37 ( .A(\ab[38][37] ), .B(\CARRYB[37][37] ), .CI(\SUMB[37][38] ), 
        .CO(\CARRYB[38][37] ), .S(\SUMB[38][37] ) );
  FA_X1 S2_38_38 ( .A(\ab[38][38] ), .B(\CARRYB[37][38] ), .CI(\SUMB[37][39] ), 
        .CO(\CARRYB[38][38] ), .S(\SUMB[38][38] ) );
  FA_X1 S2_38_39 ( .A(\ab[38][39] ), .B(\CARRYB[37][39] ), .CI(\SUMB[37][40] ), 
        .CO(\CARRYB[38][39] ), .S(\SUMB[38][39] ) );
  FA_X1 S2_38_40 ( .A(\ab[38][40] ), .B(\CARRYB[37][40] ), .CI(\SUMB[37][41] ), 
        .CO(\CARRYB[38][40] ), .S(\SUMB[38][40] ) );
  FA_X1 S2_38_41 ( .A(\ab[38][41] ), .B(\CARRYB[37][41] ), .CI(\SUMB[37][42] ), 
        .CO(\CARRYB[38][41] ), .S(\SUMB[38][41] ) );
  FA_X1 S2_38_42 ( .A(\ab[38][42] ), .B(\CARRYB[37][42] ), .CI(\SUMB[37][43] ), 
        .CO(\CARRYB[38][42] ), .S(\SUMB[38][42] ) );
  FA_X1 S2_38_43 ( .A(\ab[38][43] ), .B(\CARRYB[37][43] ), .CI(\SUMB[37][44] ), 
        .CO(\CARRYB[38][43] ), .S(\SUMB[38][43] ) );
  FA_X1 S2_38_44 ( .A(\ab[38][44] ), .B(\CARRYB[37][44] ), .CI(\SUMB[37][45] ), 
        .CO(\CARRYB[38][44] ), .S(\SUMB[38][44] ) );
  FA_X1 S2_38_45 ( .A(\ab[38][45] ), .B(\CARRYB[37][45] ), .CI(\SUMB[37][46] ), 
        .CO(\CARRYB[38][45] ), .S(\SUMB[38][45] ) );
  FA_X1 S2_38_46 ( .A(\ab[38][46] ), .B(\CARRYB[37][46] ), .CI(\SUMB[37][47] ), 
        .CO(\CARRYB[38][46] ), .S(\SUMB[38][46] ) );
  FA_X1 S2_38_47 ( .A(\ab[38][47] ), .B(\CARRYB[37][47] ), .CI(\SUMB[37][48] ), 
        .CO(\CARRYB[38][47] ), .S(\SUMB[38][47] ) );
  FA_X1 S2_38_48 ( .A(\ab[38][48] ), .B(\CARRYB[37][48] ), .CI(\SUMB[37][49] ), 
        .CO(\CARRYB[38][48] ), .S(\SUMB[38][48] ) );
  FA_X1 S2_38_49 ( .A(\ab[38][49] ), .B(\CARRYB[37][49] ), .CI(\SUMB[37][50] ), 
        .CO(\CARRYB[38][49] ), .S(\SUMB[38][49] ) );
  FA_X1 S2_38_50 ( .A(\ab[38][50] ), .B(\CARRYB[37][50] ), .CI(\SUMB[37][51] ), 
        .CO(\CARRYB[38][50] ), .S(\SUMB[38][50] ) );
  FA_X1 S3_38_51 ( .A(\ab[38][51] ), .B(\CARRYB[37][51] ), .CI(\ab[37][52] ), 
        .CO(\CARRYB[38][51] ), .S(\SUMB[38][51] ) );
  FA_X1 S1_37_0 ( .A(\ab[37][0] ), .B(\CARRYB[36][0] ), .CI(\SUMB[36][1] ), 
        .CO(\CARRYB[37][0] ), .S(CLA_SUM[37]) );
  FA_X1 S2_37_1 ( .A(\ab[37][1] ), .B(\CARRYB[36][1] ), .CI(\SUMB[36][2] ), 
        .CO(\CARRYB[37][1] ), .S(\SUMB[37][1] ) );
  FA_X1 S2_37_2 ( .A(\ab[37][2] ), .B(\CARRYB[36][2] ), .CI(\SUMB[36][3] ), 
        .CO(\CARRYB[37][2] ), .S(\SUMB[37][2] ) );
  FA_X1 S2_37_3 ( .A(\ab[37][3] ), .B(\CARRYB[36][3] ), .CI(\SUMB[36][4] ), 
        .CO(\CARRYB[37][3] ), .S(\SUMB[37][3] ) );
  FA_X1 S2_37_4 ( .A(\ab[37][4] ), .B(\CARRYB[36][4] ), .CI(\SUMB[36][5] ), 
        .CO(\CARRYB[37][4] ), .S(\SUMB[37][4] ) );
  FA_X1 S2_37_5 ( .A(\ab[37][5] ), .B(\CARRYB[36][5] ), .CI(\SUMB[36][6] ), 
        .CO(\CARRYB[37][5] ), .S(\SUMB[37][5] ) );
  FA_X1 S2_37_6 ( .A(\ab[37][6] ), .B(\CARRYB[36][6] ), .CI(\SUMB[36][7] ), 
        .CO(\CARRYB[37][6] ), .S(\SUMB[37][6] ) );
  FA_X1 S2_37_7 ( .A(\ab[37][7] ), .B(\CARRYB[36][7] ), .CI(\SUMB[36][8] ), 
        .CO(\CARRYB[37][7] ), .S(\SUMB[37][7] ) );
  FA_X1 S2_37_8 ( .A(\ab[37][8] ), .B(\CARRYB[36][8] ), .CI(\SUMB[36][9] ), 
        .CO(\CARRYB[37][8] ), .S(\SUMB[37][8] ) );
  FA_X1 S2_37_9 ( .A(\ab[37][9] ), .B(\CARRYB[36][9] ), .CI(\SUMB[36][10] ), 
        .CO(\CARRYB[37][9] ), .S(\SUMB[37][9] ) );
  FA_X1 S2_37_10 ( .A(\ab[37][10] ), .B(\CARRYB[36][10] ), .CI(\SUMB[36][11] ), 
        .CO(\CARRYB[37][10] ), .S(\SUMB[37][10] ) );
  FA_X1 S2_37_11 ( .A(\ab[37][11] ), .B(\CARRYB[36][11] ), .CI(\SUMB[36][12] ), 
        .CO(\CARRYB[37][11] ), .S(\SUMB[37][11] ) );
  FA_X1 S2_37_12 ( .A(\ab[37][12] ), .B(\CARRYB[36][12] ), .CI(\SUMB[36][13] ), 
        .CO(\CARRYB[37][12] ), .S(\SUMB[37][12] ) );
  FA_X1 S2_37_13 ( .A(\ab[37][13] ), .B(\CARRYB[36][13] ), .CI(\SUMB[36][14] ), 
        .CO(\CARRYB[37][13] ), .S(\SUMB[37][13] ) );
  FA_X1 S2_37_14 ( .A(\ab[37][14] ), .B(\CARRYB[36][14] ), .CI(\SUMB[36][15] ), 
        .CO(\CARRYB[37][14] ), .S(\SUMB[37][14] ) );
  FA_X1 S2_37_15 ( .A(\ab[37][15] ), .B(\CARRYB[36][15] ), .CI(\SUMB[36][16] ), 
        .CO(\CARRYB[37][15] ), .S(\SUMB[37][15] ) );
  FA_X1 S2_37_16 ( .A(\ab[37][16] ), .B(\CARRYB[36][16] ), .CI(\SUMB[36][17] ), 
        .CO(\CARRYB[37][16] ), .S(\SUMB[37][16] ) );
  FA_X1 S2_37_17 ( .A(\ab[37][17] ), .B(\CARRYB[36][17] ), .CI(\SUMB[36][18] ), 
        .CO(\CARRYB[37][17] ), .S(\SUMB[37][17] ) );
  FA_X1 S2_37_18 ( .A(\ab[37][18] ), .B(\CARRYB[36][18] ), .CI(\SUMB[36][19] ), 
        .CO(\CARRYB[37][18] ), .S(\SUMB[37][18] ) );
  FA_X1 S2_37_19 ( .A(\ab[37][19] ), .B(\CARRYB[36][19] ), .CI(\SUMB[36][20] ), 
        .CO(\CARRYB[37][19] ), .S(\SUMB[37][19] ) );
  FA_X1 S2_37_20 ( .A(\ab[37][20] ), .B(\CARRYB[36][20] ), .CI(\SUMB[36][21] ), 
        .CO(\CARRYB[37][20] ), .S(\SUMB[37][20] ) );
  FA_X1 S2_37_21 ( .A(\ab[37][21] ), .B(\CARRYB[36][21] ), .CI(\SUMB[36][22] ), 
        .CO(\CARRYB[37][21] ), .S(\SUMB[37][21] ) );
  FA_X1 S2_37_22 ( .A(\ab[37][22] ), .B(\CARRYB[36][22] ), .CI(\SUMB[36][23] ), 
        .CO(\CARRYB[37][22] ), .S(\SUMB[37][22] ) );
  FA_X1 S2_37_23 ( .A(\ab[37][23] ), .B(\CARRYB[36][23] ), .CI(\SUMB[36][24] ), 
        .CO(\CARRYB[37][23] ), .S(\SUMB[37][23] ) );
  FA_X1 S2_37_24 ( .A(\ab[37][24] ), .B(\CARRYB[36][24] ), .CI(\SUMB[36][25] ), 
        .CO(\CARRYB[37][24] ), .S(\SUMB[37][24] ) );
  FA_X1 S2_37_25 ( .A(\ab[37][25] ), .B(\CARRYB[36][25] ), .CI(\SUMB[36][26] ), 
        .CO(\CARRYB[37][25] ), .S(\SUMB[37][25] ) );
  FA_X1 S2_37_26 ( .A(\ab[37][26] ), .B(\CARRYB[36][26] ), .CI(\SUMB[36][27] ), 
        .CO(\CARRYB[37][26] ), .S(\SUMB[37][26] ) );
  FA_X1 S2_37_27 ( .A(\ab[37][27] ), .B(\CARRYB[36][27] ), .CI(\SUMB[36][28] ), 
        .CO(\CARRYB[37][27] ), .S(\SUMB[37][27] ) );
  FA_X1 S2_37_28 ( .A(\ab[37][28] ), .B(\CARRYB[36][28] ), .CI(\SUMB[36][29] ), 
        .CO(\CARRYB[37][28] ), .S(\SUMB[37][28] ) );
  FA_X1 S2_37_29 ( .A(\ab[37][29] ), .B(\CARRYB[36][29] ), .CI(\SUMB[36][30] ), 
        .CO(\CARRYB[37][29] ), .S(\SUMB[37][29] ) );
  FA_X1 S2_37_30 ( .A(\ab[37][30] ), .B(\CARRYB[36][30] ), .CI(\SUMB[36][31] ), 
        .CO(\CARRYB[37][30] ), .S(\SUMB[37][30] ) );
  FA_X1 S2_37_31 ( .A(\ab[37][31] ), .B(\CARRYB[36][31] ), .CI(\SUMB[36][32] ), 
        .CO(\CARRYB[37][31] ), .S(\SUMB[37][31] ) );
  FA_X1 S2_37_32 ( .A(\ab[37][32] ), .B(\CARRYB[36][32] ), .CI(\SUMB[36][33] ), 
        .CO(\CARRYB[37][32] ), .S(\SUMB[37][32] ) );
  FA_X1 S2_37_33 ( .A(\ab[37][33] ), .B(\CARRYB[36][33] ), .CI(\SUMB[36][34] ), 
        .CO(\CARRYB[37][33] ), .S(\SUMB[37][33] ) );
  FA_X1 S2_37_34 ( .A(\ab[37][34] ), .B(\CARRYB[36][34] ), .CI(\SUMB[36][35] ), 
        .CO(\CARRYB[37][34] ), .S(\SUMB[37][34] ) );
  FA_X1 S2_37_35 ( .A(\ab[37][35] ), .B(\CARRYB[36][35] ), .CI(\SUMB[36][36] ), 
        .CO(\CARRYB[37][35] ), .S(\SUMB[37][35] ) );
  FA_X1 S2_37_36 ( .A(\ab[37][36] ), .B(\CARRYB[36][36] ), .CI(\SUMB[36][37] ), 
        .CO(\CARRYB[37][36] ), .S(\SUMB[37][36] ) );
  FA_X1 S2_37_37 ( .A(\ab[37][37] ), .B(\CARRYB[36][37] ), .CI(\SUMB[36][38] ), 
        .CO(\CARRYB[37][37] ), .S(\SUMB[37][37] ) );
  FA_X1 S2_37_38 ( .A(\ab[37][38] ), .B(\CARRYB[36][38] ), .CI(\SUMB[36][39] ), 
        .CO(\CARRYB[37][38] ), .S(\SUMB[37][38] ) );
  FA_X1 S2_37_39 ( .A(\ab[37][39] ), .B(\CARRYB[36][39] ), .CI(\SUMB[36][40] ), 
        .CO(\CARRYB[37][39] ), .S(\SUMB[37][39] ) );
  FA_X1 S2_37_40 ( .A(\ab[37][40] ), .B(\CARRYB[36][40] ), .CI(\SUMB[36][41] ), 
        .CO(\CARRYB[37][40] ), .S(\SUMB[37][40] ) );
  FA_X1 S2_37_41 ( .A(\ab[37][41] ), .B(\CARRYB[36][41] ), .CI(\SUMB[36][42] ), 
        .CO(\CARRYB[37][41] ), .S(\SUMB[37][41] ) );
  FA_X1 S2_37_42 ( .A(\ab[37][42] ), .B(\CARRYB[36][42] ), .CI(\SUMB[36][43] ), 
        .CO(\CARRYB[37][42] ), .S(\SUMB[37][42] ) );
  FA_X1 S2_37_43 ( .A(\ab[37][43] ), .B(\CARRYB[36][43] ), .CI(\SUMB[36][44] ), 
        .CO(\CARRYB[37][43] ), .S(\SUMB[37][43] ) );
  FA_X1 S2_37_44 ( .A(\ab[37][44] ), .B(\CARRYB[36][44] ), .CI(\SUMB[36][45] ), 
        .CO(\CARRYB[37][44] ), .S(\SUMB[37][44] ) );
  FA_X1 S2_37_45 ( .A(\ab[37][45] ), .B(\CARRYB[36][45] ), .CI(\SUMB[36][46] ), 
        .CO(\CARRYB[37][45] ), .S(\SUMB[37][45] ) );
  FA_X1 S2_37_46 ( .A(\ab[37][46] ), .B(\CARRYB[36][46] ), .CI(\SUMB[36][47] ), 
        .CO(\CARRYB[37][46] ), .S(\SUMB[37][46] ) );
  FA_X1 S2_37_47 ( .A(\ab[37][47] ), .B(\CARRYB[36][47] ), .CI(\SUMB[36][48] ), 
        .CO(\CARRYB[37][47] ), .S(\SUMB[37][47] ) );
  FA_X1 S2_37_48 ( .A(\ab[37][48] ), .B(\CARRYB[36][48] ), .CI(\SUMB[36][49] ), 
        .CO(\CARRYB[37][48] ), .S(\SUMB[37][48] ) );
  FA_X1 S2_37_49 ( .A(\ab[37][49] ), .B(\CARRYB[36][49] ), .CI(\SUMB[36][50] ), 
        .CO(\CARRYB[37][49] ), .S(\SUMB[37][49] ) );
  FA_X1 S2_37_50 ( .A(\ab[37][50] ), .B(\CARRYB[36][50] ), .CI(\SUMB[36][51] ), 
        .CO(\CARRYB[37][50] ), .S(\SUMB[37][50] ) );
  FA_X1 S3_37_51 ( .A(\ab[37][51] ), .B(\CARRYB[36][51] ), .CI(\ab[36][52] ), 
        .CO(\CARRYB[37][51] ), .S(\SUMB[37][51] ) );
  FA_X1 S1_36_0 ( .A(\ab[36][0] ), .B(\CARRYB[35][0] ), .CI(\SUMB[35][1] ), 
        .CO(\CARRYB[36][0] ), .S(CLA_SUM[36]) );
  FA_X1 S2_36_1 ( .A(\ab[36][1] ), .B(\CARRYB[35][1] ), .CI(\SUMB[35][2] ), 
        .CO(\CARRYB[36][1] ), .S(\SUMB[36][1] ) );
  FA_X1 S2_36_2 ( .A(\ab[36][2] ), .B(\CARRYB[35][2] ), .CI(\SUMB[35][3] ), 
        .CO(\CARRYB[36][2] ), .S(\SUMB[36][2] ) );
  FA_X1 S2_36_3 ( .A(\ab[36][3] ), .B(\CARRYB[35][3] ), .CI(\SUMB[35][4] ), 
        .CO(\CARRYB[36][3] ), .S(\SUMB[36][3] ) );
  FA_X1 S2_36_4 ( .A(\ab[36][4] ), .B(\CARRYB[35][4] ), .CI(\SUMB[35][5] ), 
        .CO(\CARRYB[36][4] ), .S(\SUMB[36][4] ) );
  FA_X1 S2_36_5 ( .A(\ab[36][5] ), .B(\CARRYB[35][5] ), .CI(\SUMB[35][6] ), 
        .CO(\CARRYB[36][5] ), .S(\SUMB[36][5] ) );
  FA_X1 S2_36_6 ( .A(\ab[36][6] ), .B(\CARRYB[35][6] ), .CI(\SUMB[35][7] ), 
        .CO(\CARRYB[36][6] ), .S(\SUMB[36][6] ) );
  FA_X1 S2_36_7 ( .A(\ab[36][7] ), .B(\CARRYB[35][7] ), .CI(\SUMB[35][8] ), 
        .CO(\CARRYB[36][7] ), .S(\SUMB[36][7] ) );
  FA_X1 S2_36_8 ( .A(\ab[36][8] ), .B(\CARRYB[35][8] ), .CI(\SUMB[35][9] ), 
        .CO(\CARRYB[36][8] ), .S(\SUMB[36][8] ) );
  FA_X1 S2_36_9 ( .A(\ab[36][9] ), .B(\CARRYB[35][9] ), .CI(\SUMB[35][10] ), 
        .CO(\CARRYB[36][9] ), .S(\SUMB[36][9] ) );
  FA_X1 S2_36_10 ( .A(\ab[36][10] ), .B(\CARRYB[35][10] ), .CI(\SUMB[35][11] ), 
        .CO(\CARRYB[36][10] ), .S(\SUMB[36][10] ) );
  FA_X1 S2_36_11 ( .A(\ab[36][11] ), .B(\CARRYB[35][11] ), .CI(\SUMB[35][12] ), 
        .CO(\CARRYB[36][11] ), .S(\SUMB[36][11] ) );
  FA_X1 S2_36_12 ( .A(\ab[36][12] ), .B(\CARRYB[35][12] ), .CI(\SUMB[35][13] ), 
        .CO(\CARRYB[36][12] ), .S(\SUMB[36][12] ) );
  FA_X1 S2_36_13 ( .A(\ab[36][13] ), .B(\CARRYB[35][13] ), .CI(\SUMB[35][14] ), 
        .CO(\CARRYB[36][13] ), .S(\SUMB[36][13] ) );
  FA_X1 S2_36_14 ( .A(\ab[36][14] ), .B(\CARRYB[35][14] ), .CI(\SUMB[35][15] ), 
        .CO(\CARRYB[36][14] ), .S(\SUMB[36][14] ) );
  FA_X1 S2_36_15 ( .A(\ab[36][15] ), .B(\CARRYB[35][15] ), .CI(\SUMB[35][16] ), 
        .CO(\CARRYB[36][15] ), .S(\SUMB[36][15] ) );
  FA_X1 S2_36_16 ( .A(\ab[36][16] ), .B(\CARRYB[35][16] ), .CI(\SUMB[35][17] ), 
        .CO(\CARRYB[36][16] ), .S(\SUMB[36][16] ) );
  FA_X1 S2_36_17 ( .A(\ab[36][17] ), .B(\CARRYB[35][17] ), .CI(\SUMB[35][18] ), 
        .CO(\CARRYB[36][17] ), .S(\SUMB[36][17] ) );
  FA_X1 S2_36_18 ( .A(\ab[36][18] ), .B(\CARRYB[35][18] ), .CI(\SUMB[35][19] ), 
        .CO(\CARRYB[36][18] ), .S(\SUMB[36][18] ) );
  FA_X1 S2_36_19 ( .A(\ab[36][19] ), .B(\CARRYB[35][19] ), .CI(\SUMB[35][20] ), 
        .CO(\CARRYB[36][19] ), .S(\SUMB[36][19] ) );
  FA_X1 S2_36_20 ( .A(\ab[36][20] ), .B(\CARRYB[35][20] ), .CI(\SUMB[35][21] ), 
        .CO(\CARRYB[36][20] ), .S(\SUMB[36][20] ) );
  FA_X1 S2_36_21 ( .A(\ab[36][21] ), .B(\CARRYB[35][21] ), .CI(\SUMB[35][22] ), 
        .CO(\CARRYB[36][21] ), .S(\SUMB[36][21] ) );
  FA_X1 S2_36_22 ( .A(\ab[36][22] ), .B(\CARRYB[35][22] ), .CI(\SUMB[35][23] ), 
        .CO(\CARRYB[36][22] ), .S(\SUMB[36][22] ) );
  FA_X1 S2_36_23 ( .A(\ab[36][23] ), .B(\CARRYB[35][23] ), .CI(\SUMB[35][24] ), 
        .CO(\CARRYB[36][23] ), .S(\SUMB[36][23] ) );
  FA_X1 S2_36_24 ( .A(\ab[36][24] ), .B(\CARRYB[35][24] ), .CI(\SUMB[35][25] ), 
        .CO(\CARRYB[36][24] ), .S(\SUMB[36][24] ) );
  FA_X1 S2_36_25 ( .A(\ab[36][25] ), .B(\CARRYB[35][25] ), .CI(\SUMB[35][26] ), 
        .CO(\CARRYB[36][25] ), .S(\SUMB[36][25] ) );
  FA_X1 S2_36_26 ( .A(\ab[36][26] ), .B(\CARRYB[35][26] ), .CI(\SUMB[35][27] ), 
        .CO(\CARRYB[36][26] ), .S(\SUMB[36][26] ) );
  FA_X1 S2_36_27 ( .A(\ab[36][27] ), .B(\CARRYB[35][27] ), .CI(\SUMB[35][28] ), 
        .CO(\CARRYB[36][27] ), .S(\SUMB[36][27] ) );
  FA_X1 S2_36_28 ( .A(\ab[36][28] ), .B(\CARRYB[35][28] ), .CI(\SUMB[35][29] ), 
        .CO(\CARRYB[36][28] ), .S(\SUMB[36][28] ) );
  FA_X1 S2_36_29 ( .A(\ab[36][29] ), .B(\CARRYB[35][29] ), .CI(\SUMB[35][30] ), 
        .CO(\CARRYB[36][29] ), .S(\SUMB[36][29] ) );
  FA_X1 S2_36_30 ( .A(\ab[36][30] ), .B(\CARRYB[35][30] ), .CI(\SUMB[35][31] ), 
        .CO(\CARRYB[36][30] ), .S(\SUMB[36][30] ) );
  FA_X1 S2_36_31 ( .A(\ab[36][31] ), .B(\CARRYB[35][31] ), .CI(\SUMB[35][32] ), 
        .CO(\CARRYB[36][31] ), .S(\SUMB[36][31] ) );
  FA_X1 S2_36_32 ( .A(\ab[36][32] ), .B(\CARRYB[35][32] ), .CI(\SUMB[35][33] ), 
        .CO(\CARRYB[36][32] ), .S(\SUMB[36][32] ) );
  FA_X1 S2_36_33 ( .A(\ab[36][33] ), .B(\CARRYB[35][33] ), .CI(\SUMB[35][34] ), 
        .CO(\CARRYB[36][33] ), .S(\SUMB[36][33] ) );
  FA_X1 S2_36_34 ( .A(\ab[36][34] ), .B(\CARRYB[35][34] ), .CI(\SUMB[35][35] ), 
        .CO(\CARRYB[36][34] ), .S(\SUMB[36][34] ) );
  FA_X1 S2_36_35 ( .A(\ab[36][35] ), .B(\CARRYB[35][35] ), .CI(\SUMB[35][36] ), 
        .CO(\CARRYB[36][35] ), .S(\SUMB[36][35] ) );
  FA_X1 S2_36_36 ( .A(\ab[36][36] ), .B(\CARRYB[35][36] ), .CI(\SUMB[35][37] ), 
        .CO(\CARRYB[36][36] ), .S(\SUMB[36][36] ) );
  FA_X1 S2_36_37 ( .A(\ab[36][37] ), .B(\CARRYB[35][37] ), .CI(\SUMB[35][38] ), 
        .CO(\CARRYB[36][37] ), .S(\SUMB[36][37] ) );
  FA_X1 S2_36_38 ( .A(\ab[36][38] ), .B(\CARRYB[35][38] ), .CI(\SUMB[35][39] ), 
        .CO(\CARRYB[36][38] ), .S(\SUMB[36][38] ) );
  FA_X1 S2_36_39 ( .A(\ab[36][39] ), .B(\CARRYB[35][39] ), .CI(\SUMB[35][40] ), 
        .CO(\CARRYB[36][39] ), .S(\SUMB[36][39] ) );
  FA_X1 S2_36_40 ( .A(\ab[36][40] ), .B(\CARRYB[35][40] ), .CI(\SUMB[35][41] ), 
        .CO(\CARRYB[36][40] ), .S(\SUMB[36][40] ) );
  FA_X1 S2_36_41 ( .A(\ab[36][41] ), .B(\CARRYB[35][41] ), .CI(\SUMB[35][42] ), 
        .CO(\CARRYB[36][41] ), .S(\SUMB[36][41] ) );
  FA_X1 S2_36_42 ( .A(\ab[36][42] ), .B(\CARRYB[35][42] ), .CI(\SUMB[35][43] ), 
        .CO(\CARRYB[36][42] ), .S(\SUMB[36][42] ) );
  FA_X1 S2_36_43 ( .A(\ab[36][43] ), .B(\CARRYB[35][43] ), .CI(\SUMB[35][44] ), 
        .CO(\CARRYB[36][43] ), .S(\SUMB[36][43] ) );
  FA_X1 S2_36_44 ( .A(\ab[36][44] ), .B(\CARRYB[35][44] ), .CI(\SUMB[35][45] ), 
        .CO(\CARRYB[36][44] ), .S(\SUMB[36][44] ) );
  FA_X1 S2_36_45 ( .A(\ab[36][45] ), .B(\CARRYB[35][45] ), .CI(\SUMB[35][46] ), 
        .CO(\CARRYB[36][45] ), .S(\SUMB[36][45] ) );
  FA_X1 S2_36_46 ( .A(\ab[36][46] ), .B(\CARRYB[35][46] ), .CI(\SUMB[35][47] ), 
        .CO(\CARRYB[36][46] ), .S(\SUMB[36][46] ) );
  FA_X1 S2_36_47 ( .A(\ab[36][47] ), .B(\CARRYB[35][47] ), .CI(\SUMB[35][48] ), 
        .CO(\CARRYB[36][47] ), .S(\SUMB[36][47] ) );
  FA_X1 S2_36_48 ( .A(\ab[36][48] ), .B(\CARRYB[35][48] ), .CI(\SUMB[35][49] ), 
        .CO(\CARRYB[36][48] ), .S(\SUMB[36][48] ) );
  FA_X1 S2_36_49 ( .A(\ab[36][49] ), .B(\CARRYB[35][49] ), .CI(\SUMB[35][50] ), 
        .CO(\CARRYB[36][49] ), .S(\SUMB[36][49] ) );
  FA_X1 S2_36_50 ( .A(\ab[36][50] ), .B(\CARRYB[35][50] ), .CI(\SUMB[35][51] ), 
        .CO(\CARRYB[36][50] ), .S(\SUMB[36][50] ) );
  FA_X1 S3_36_51 ( .A(\ab[36][51] ), .B(\CARRYB[35][51] ), .CI(\ab[35][52] ), 
        .CO(\CARRYB[36][51] ), .S(\SUMB[36][51] ) );
  FA_X1 S1_35_0 ( .A(\ab[35][0] ), .B(\CARRYB[34][0] ), .CI(\SUMB[34][1] ), 
        .CO(\CARRYB[35][0] ), .S(CLA_SUM[35]) );
  FA_X1 S2_35_1 ( .A(\ab[35][1] ), .B(\CARRYB[34][1] ), .CI(\SUMB[34][2] ), 
        .CO(\CARRYB[35][1] ), .S(\SUMB[35][1] ) );
  FA_X1 S2_35_2 ( .A(\ab[35][2] ), .B(\CARRYB[34][2] ), .CI(\SUMB[34][3] ), 
        .CO(\CARRYB[35][2] ), .S(\SUMB[35][2] ) );
  FA_X1 S2_35_3 ( .A(\ab[35][3] ), .B(\CARRYB[34][3] ), .CI(\SUMB[34][4] ), 
        .CO(\CARRYB[35][3] ), .S(\SUMB[35][3] ) );
  FA_X1 S2_35_4 ( .A(\ab[35][4] ), .B(\CARRYB[34][4] ), .CI(\SUMB[34][5] ), 
        .CO(\CARRYB[35][4] ), .S(\SUMB[35][4] ) );
  FA_X1 S2_35_5 ( .A(\ab[35][5] ), .B(\CARRYB[34][5] ), .CI(\SUMB[34][6] ), 
        .CO(\CARRYB[35][5] ), .S(\SUMB[35][5] ) );
  FA_X1 S2_35_6 ( .A(\ab[35][6] ), .B(\CARRYB[34][6] ), .CI(\SUMB[34][7] ), 
        .CO(\CARRYB[35][6] ), .S(\SUMB[35][6] ) );
  FA_X1 S2_35_7 ( .A(\ab[35][7] ), .B(\CARRYB[34][7] ), .CI(\SUMB[34][8] ), 
        .CO(\CARRYB[35][7] ), .S(\SUMB[35][7] ) );
  FA_X1 S2_35_8 ( .A(\ab[35][8] ), .B(\CARRYB[34][8] ), .CI(\SUMB[34][9] ), 
        .CO(\CARRYB[35][8] ), .S(\SUMB[35][8] ) );
  FA_X1 S2_35_9 ( .A(\ab[35][9] ), .B(\CARRYB[34][9] ), .CI(\SUMB[34][10] ), 
        .CO(\CARRYB[35][9] ), .S(\SUMB[35][9] ) );
  FA_X1 S2_35_10 ( .A(\ab[35][10] ), .B(\CARRYB[34][10] ), .CI(\SUMB[34][11] ), 
        .CO(\CARRYB[35][10] ), .S(\SUMB[35][10] ) );
  FA_X1 S2_35_11 ( .A(\ab[35][11] ), .B(\CARRYB[34][11] ), .CI(\SUMB[34][12] ), 
        .CO(\CARRYB[35][11] ), .S(\SUMB[35][11] ) );
  FA_X1 S2_35_12 ( .A(\ab[35][12] ), .B(\CARRYB[34][12] ), .CI(\SUMB[34][13] ), 
        .CO(\CARRYB[35][12] ), .S(\SUMB[35][12] ) );
  FA_X1 S2_35_13 ( .A(\ab[35][13] ), .B(\CARRYB[34][13] ), .CI(\SUMB[34][14] ), 
        .CO(\CARRYB[35][13] ), .S(\SUMB[35][13] ) );
  FA_X1 S2_35_14 ( .A(\ab[35][14] ), .B(\CARRYB[34][14] ), .CI(\SUMB[34][15] ), 
        .CO(\CARRYB[35][14] ), .S(\SUMB[35][14] ) );
  FA_X1 S2_35_15 ( .A(\ab[35][15] ), .B(\CARRYB[34][15] ), .CI(\SUMB[34][16] ), 
        .CO(\CARRYB[35][15] ), .S(\SUMB[35][15] ) );
  FA_X1 S2_35_16 ( .A(\ab[35][16] ), .B(\CARRYB[34][16] ), .CI(\SUMB[34][17] ), 
        .CO(\CARRYB[35][16] ), .S(\SUMB[35][16] ) );
  FA_X1 S2_35_17 ( .A(\ab[35][17] ), .B(\CARRYB[34][17] ), .CI(\SUMB[34][18] ), 
        .CO(\CARRYB[35][17] ), .S(\SUMB[35][17] ) );
  FA_X1 S2_35_18 ( .A(\ab[35][18] ), .B(\CARRYB[34][18] ), .CI(\SUMB[34][19] ), 
        .CO(\CARRYB[35][18] ), .S(\SUMB[35][18] ) );
  FA_X1 S2_35_19 ( .A(\ab[35][19] ), .B(\CARRYB[34][19] ), .CI(\SUMB[34][20] ), 
        .CO(\CARRYB[35][19] ), .S(\SUMB[35][19] ) );
  FA_X1 S2_35_20 ( .A(\ab[35][20] ), .B(\CARRYB[34][20] ), .CI(\SUMB[34][21] ), 
        .CO(\CARRYB[35][20] ), .S(\SUMB[35][20] ) );
  FA_X1 S2_35_21 ( .A(\ab[35][21] ), .B(\CARRYB[34][21] ), .CI(\SUMB[34][22] ), 
        .CO(\CARRYB[35][21] ), .S(\SUMB[35][21] ) );
  FA_X1 S2_35_22 ( .A(\ab[35][22] ), .B(\CARRYB[34][22] ), .CI(\SUMB[34][23] ), 
        .CO(\CARRYB[35][22] ), .S(\SUMB[35][22] ) );
  FA_X1 S2_35_23 ( .A(\ab[35][23] ), .B(\CARRYB[34][23] ), .CI(\SUMB[34][24] ), 
        .CO(\CARRYB[35][23] ), .S(\SUMB[35][23] ) );
  FA_X1 S2_35_24 ( .A(\ab[35][24] ), .B(\CARRYB[34][24] ), .CI(\SUMB[34][25] ), 
        .CO(\CARRYB[35][24] ), .S(\SUMB[35][24] ) );
  FA_X1 S2_35_25 ( .A(\ab[35][25] ), .B(\CARRYB[34][25] ), .CI(\SUMB[34][26] ), 
        .CO(\CARRYB[35][25] ), .S(\SUMB[35][25] ) );
  FA_X1 S2_35_26 ( .A(\ab[35][26] ), .B(\CARRYB[34][26] ), .CI(\SUMB[34][27] ), 
        .CO(\CARRYB[35][26] ), .S(\SUMB[35][26] ) );
  FA_X1 S2_35_27 ( .A(\ab[35][27] ), .B(\CARRYB[34][27] ), .CI(\SUMB[34][28] ), 
        .CO(\CARRYB[35][27] ), .S(\SUMB[35][27] ) );
  FA_X1 S2_35_28 ( .A(\ab[35][28] ), .B(\CARRYB[34][28] ), .CI(\SUMB[34][29] ), 
        .CO(\CARRYB[35][28] ), .S(\SUMB[35][28] ) );
  FA_X1 S2_35_29 ( .A(\ab[35][29] ), .B(\CARRYB[34][29] ), .CI(\SUMB[34][30] ), 
        .CO(\CARRYB[35][29] ), .S(\SUMB[35][29] ) );
  FA_X1 S2_35_30 ( .A(\ab[35][30] ), .B(\CARRYB[34][30] ), .CI(\SUMB[34][31] ), 
        .CO(\CARRYB[35][30] ), .S(\SUMB[35][30] ) );
  FA_X1 S2_35_31 ( .A(\ab[35][31] ), .B(\CARRYB[34][31] ), .CI(\SUMB[34][32] ), 
        .CO(\CARRYB[35][31] ), .S(\SUMB[35][31] ) );
  FA_X1 S2_35_32 ( .A(\ab[35][32] ), .B(\CARRYB[34][32] ), .CI(\SUMB[34][33] ), 
        .CO(\CARRYB[35][32] ), .S(\SUMB[35][32] ) );
  FA_X1 S2_35_33 ( .A(\ab[35][33] ), .B(\CARRYB[34][33] ), .CI(\SUMB[34][34] ), 
        .CO(\CARRYB[35][33] ), .S(\SUMB[35][33] ) );
  FA_X1 S2_35_34 ( .A(\ab[35][34] ), .B(\CARRYB[34][34] ), .CI(\SUMB[34][35] ), 
        .CO(\CARRYB[35][34] ), .S(\SUMB[35][34] ) );
  FA_X1 S2_35_35 ( .A(\ab[35][35] ), .B(\CARRYB[34][35] ), .CI(\SUMB[34][36] ), 
        .CO(\CARRYB[35][35] ), .S(\SUMB[35][35] ) );
  FA_X1 S2_35_36 ( .A(\ab[35][36] ), .B(\CARRYB[34][36] ), .CI(\SUMB[34][37] ), 
        .CO(\CARRYB[35][36] ), .S(\SUMB[35][36] ) );
  FA_X1 S2_35_37 ( .A(\ab[35][37] ), .B(\CARRYB[34][37] ), .CI(\SUMB[34][38] ), 
        .CO(\CARRYB[35][37] ), .S(\SUMB[35][37] ) );
  FA_X1 S2_35_38 ( .A(\ab[35][38] ), .B(\CARRYB[34][38] ), .CI(\SUMB[34][39] ), 
        .CO(\CARRYB[35][38] ), .S(\SUMB[35][38] ) );
  FA_X1 S2_35_39 ( .A(\ab[35][39] ), .B(\CARRYB[34][39] ), .CI(\SUMB[34][40] ), 
        .CO(\CARRYB[35][39] ), .S(\SUMB[35][39] ) );
  FA_X1 S2_35_40 ( .A(\ab[35][40] ), .B(\CARRYB[34][40] ), .CI(\SUMB[34][41] ), 
        .CO(\CARRYB[35][40] ), .S(\SUMB[35][40] ) );
  FA_X1 S2_35_41 ( .A(\ab[35][41] ), .B(\CARRYB[34][41] ), .CI(\SUMB[34][42] ), 
        .CO(\CARRYB[35][41] ), .S(\SUMB[35][41] ) );
  FA_X1 S2_35_42 ( .A(\ab[35][42] ), .B(\CARRYB[34][42] ), .CI(\SUMB[34][43] ), 
        .CO(\CARRYB[35][42] ), .S(\SUMB[35][42] ) );
  FA_X1 S2_35_43 ( .A(\ab[35][43] ), .B(\CARRYB[34][43] ), .CI(\SUMB[34][44] ), 
        .CO(\CARRYB[35][43] ), .S(\SUMB[35][43] ) );
  FA_X1 S2_35_44 ( .A(\ab[35][44] ), .B(\CARRYB[34][44] ), .CI(\SUMB[34][45] ), 
        .CO(\CARRYB[35][44] ), .S(\SUMB[35][44] ) );
  FA_X1 S2_35_45 ( .A(\ab[35][45] ), .B(\CARRYB[34][45] ), .CI(\SUMB[34][46] ), 
        .CO(\CARRYB[35][45] ), .S(\SUMB[35][45] ) );
  FA_X1 S2_35_46 ( .A(\ab[35][46] ), .B(\CARRYB[34][46] ), .CI(\SUMB[34][47] ), 
        .CO(\CARRYB[35][46] ), .S(\SUMB[35][46] ) );
  FA_X1 S2_35_47 ( .A(\ab[35][47] ), .B(\CARRYB[34][47] ), .CI(\SUMB[34][48] ), 
        .CO(\CARRYB[35][47] ), .S(\SUMB[35][47] ) );
  FA_X1 S2_35_48 ( .A(\ab[35][48] ), .B(\CARRYB[34][48] ), .CI(\SUMB[34][49] ), 
        .CO(\CARRYB[35][48] ), .S(\SUMB[35][48] ) );
  FA_X1 S2_35_49 ( .A(\ab[35][49] ), .B(\CARRYB[34][49] ), .CI(\SUMB[34][50] ), 
        .CO(\CARRYB[35][49] ), .S(\SUMB[35][49] ) );
  FA_X1 S2_35_50 ( .A(\ab[35][50] ), .B(\CARRYB[34][50] ), .CI(\SUMB[34][51] ), 
        .CO(\CARRYB[35][50] ), .S(\SUMB[35][50] ) );
  FA_X1 S3_35_51 ( .A(\ab[35][51] ), .B(\CARRYB[34][51] ), .CI(\ab[34][52] ), 
        .CO(\CARRYB[35][51] ), .S(\SUMB[35][51] ) );
  FA_X1 S1_34_0 ( .A(\ab[34][0] ), .B(\CARRYB[33][0] ), .CI(\SUMB[33][1] ), 
        .CO(\CARRYB[34][0] ), .S(CLA_SUM[34]) );
  FA_X1 S2_34_1 ( .A(\ab[34][1] ), .B(\CARRYB[33][1] ), .CI(\SUMB[33][2] ), 
        .CO(\CARRYB[34][1] ), .S(\SUMB[34][1] ) );
  FA_X1 S2_34_2 ( .A(\ab[34][2] ), .B(\CARRYB[33][2] ), .CI(\SUMB[33][3] ), 
        .CO(\CARRYB[34][2] ), .S(\SUMB[34][2] ) );
  FA_X1 S2_34_3 ( .A(\ab[34][3] ), .B(\CARRYB[33][3] ), .CI(\SUMB[33][4] ), 
        .CO(\CARRYB[34][3] ), .S(\SUMB[34][3] ) );
  FA_X1 S2_34_4 ( .A(\ab[34][4] ), .B(\CARRYB[33][4] ), .CI(\SUMB[33][5] ), 
        .CO(\CARRYB[34][4] ), .S(\SUMB[34][4] ) );
  FA_X1 S2_34_5 ( .A(\ab[34][5] ), .B(\CARRYB[33][5] ), .CI(\SUMB[33][6] ), 
        .CO(\CARRYB[34][5] ), .S(\SUMB[34][5] ) );
  FA_X1 S2_34_6 ( .A(\ab[34][6] ), .B(\CARRYB[33][6] ), .CI(\SUMB[33][7] ), 
        .CO(\CARRYB[34][6] ), .S(\SUMB[34][6] ) );
  FA_X1 S2_34_7 ( .A(\ab[34][7] ), .B(\CARRYB[33][7] ), .CI(\SUMB[33][8] ), 
        .CO(\CARRYB[34][7] ), .S(\SUMB[34][7] ) );
  FA_X1 S2_34_8 ( .A(\ab[34][8] ), .B(\CARRYB[33][8] ), .CI(\SUMB[33][9] ), 
        .CO(\CARRYB[34][8] ), .S(\SUMB[34][8] ) );
  FA_X1 S2_34_9 ( .A(\ab[34][9] ), .B(\CARRYB[33][9] ), .CI(\SUMB[33][10] ), 
        .CO(\CARRYB[34][9] ), .S(\SUMB[34][9] ) );
  FA_X1 S2_34_10 ( .A(\ab[34][10] ), .B(\CARRYB[33][10] ), .CI(\SUMB[33][11] ), 
        .CO(\CARRYB[34][10] ), .S(\SUMB[34][10] ) );
  FA_X1 S2_34_11 ( .A(\ab[34][11] ), .B(\CARRYB[33][11] ), .CI(\SUMB[33][12] ), 
        .CO(\CARRYB[34][11] ), .S(\SUMB[34][11] ) );
  FA_X1 S2_34_12 ( .A(\ab[34][12] ), .B(\CARRYB[33][12] ), .CI(\SUMB[33][13] ), 
        .CO(\CARRYB[34][12] ), .S(\SUMB[34][12] ) );
  FA_X1 S2_34_13 ( .A(\ab[34][13] ), .B(\CARRYB[33][13] ), .CI(\SUMB[33][14] ), 
        .CO(\CARRYB[34][13] ), .S(\SUMB[34][13] ) );
  FA_X1 S2_34_14 ( .A(\ab[34][14] ), .B(\CARRYB[33][14] ), .CI(\SUMB[33][15] ), 
        .CO(\CARRYB[34][14] ), .S(\SUMB[34][14] ) );
  FA_X1 S2_34_15 ( .A(\ab[34][15] ), .B(\CARRYB[33][15] ), .CI(\SUMB[33][16] ), 
        .CO(\CARRYB[34][15] ), .S(\SUMB[34][15] ) );
  FA_X1 S2_34_16 ( .A(\ab[34][16] ), .B(\CARRYB[33][16] ), .CI(\SUMB[33][17] ), 
        .CO(\CARRYB[34][16] ), .S(\SUMB[34][16] ) );
  FA_X1 S2_34_17 ( .A(\ab[34][17] ), .B(\CARRYB[33][17] ), .CI(\SUMB[33][18] ), 
        .CO(\CARRYB[34][17] ), .S(\SUMB[34][17] ) );
  FA_X1 S2_34_18 ( .A(\ab[34][18] ), .B(\CARRYB[33][18] ), .CI(\SUMB[33][19] ), 
        .CO(\CARRYB[34][18] ), .S(\SUMB[34][18] ) );
  FA_X1 S2_34_19 ( .A(\ab[34][19] ), .B(\CARRYB[33][19] ), .CI(\SUMB[33][20] ), 
        .CO(\CARRYB[34][19] ), .S(\SUMB[34][19] ) );
  FA_X1 S2_34_20 ( .A(\ab[34][20] ), .B(\CARRYB[33][20] ), .CI(\SUMB[33][21] ), 
        .CO(\CARRYB[34][20] ), .S(\SUMB[34][20] ) );
  FA_X1 S2_34_21 ( .A(\ab[34][21] ), .B(\CARRYB[33][21] ), .CI(\SUMB[33][22] ), 
        .CO(\CARRYB[34][21] ), .S(\SUMB[34][21] ) );
  FA_X1 S2_34_22 ( .A(\ab[34][22] ), .B(\CARRYB[33][22] ), .CI(\SUMB[33][23] ), 
        .CO(\CARRYB[34][22] ), .S(\SUMB[34][22] ) );
  FA_X1 S2_34_23 ( .A(\ab[34][23] ), .B(\CARRYB[33][23] ), .CI(\SUMB[33][24] ), 
        .CO(\CARRYB[34][23] ), .S(\SUMB[34][23] ) );
  FA_X1 S2_34_24 ( .A(\ab[34][24] ), .B(\CARRYB[33][24] ), .CI(\SUMB[33][25] ), 
        .CO(\CARRYB[34][24] ), .S(\SUMB[34][24] ) );
  FA_X1 S2_34_25 ( .A(\ab[34][25] ), .B(\CARRYB[33][25] ), .CI(\SUMB[33][26] ), 
        .CO(\CARRYB[34][25] ), .S(\SUMB[34][25] ) );
  FA_X1 S2_34_26 ( .A(\ab[34][26] ), .B(\CARRYB[33][26] ), .CI(\SUMB[33][27] ), 
        .CO(\CARRYB[34][26] ), .S(\SUMB[34][26] ) );
  FA_X1 S2_34_27 ( .A(\ab[34][27] ), .B(\CARRYB[33][27] ), .CI(\SUMB[33][28] ), 
        .CO(\CARRYB[34][27] ), .S(\SUMB[34][27] ) );
  FA_X1 S2_34_28 ( .A(\ab[34][28] ), .B(\CARRYB[33][28] ), .CI(\SUMB[33][29] ), 
        .CO(\CARRYB[34][28] ), .S(\SUMB[34][28] ) );
  FA_X1 S2_34_29 ( .A(\ab[34][29] ), .B(\CARRYB[33][29] ), .CI(\SUMB[33][30] ), 
        .CO(\CARRYB[34][29] ), .S(\SUMB[34][29] ) );
  FA_X1 S2_34_30 ( .A(\ab[34][30] ), .B(\CARRYB[33][30] ), .CI(\SUMB[33][31] ), 
        .CO(\CARRYB[34][30] ), .S(\SUMB[34][30] ) );
  FA_X1 S2_34_31 ( .A(\ab[34][31] ), .B(\CARRYB[33][31] ), .CI(\SUMB[33][32] ), 
        .CO(\CARRYB[34][31] ), .S(\SUMB[34][31] ) );
  FA_X1 S2_34_32 ( .A(\ab[34][32] ), .B(\CARRYB[33][32] ), .CI(\SUMB[33][33] ), 
        .CO(\CARRYB[34][32] ), .S(\SUMB[34][32] ) );
  FA_X1 S2_34_33 ( .A(\ab[34][33] ), .B(\CARRYB[33][33] ), .CI(\SUMB[33][34] ), 
        .CO(\CARRYB[34][33] ), .S(\SUMB[34][33] ) );
  FA_X1 S2_34_34 ( .A(\ab[34][34] ), .B(\CARRYB[33][34] ), .CI(\SUMB[33][35] ), 
        .CO(\CARRYB[34][34] ), .S(\SUMB[34][34] ) );
  FA_X1 S2_34_35 ( .A(\ab[34][35] ), .B(\CARRYB[33][35] ), .CI(\SUMB[33][36] ), 
        .CO(\CARRYB[34][35] ), .S(\SUMB[34][35] ) );
  FA_X1 S2_34_36 ( .A(\ab[34][36] ), .B(\CARRYB[33][36] ), .CI(\SUMB[33][37] ), 
        .CO(\CARRYB[34][36] ), .S(\SUMB[34][36] ) );
  FA_X1 S2_34_37 ( .A(\ab[34][37] ), .B(\CARRYB[33][37] ), .CI(\SUMB[33][38] ), 
        .CO(\CARRYB[34][37] ), .S(\SUMB[34][37] ) );
  FA_X1 S2_34_38 ( .A(\ab[34][38] ), .B(\CARRYB[33][38] ), .CI(\SUMB[33][39] ), 
        .CO(\CARRYB[34][38] ), .S(\SUMB[34][38] ) );
  FA_X1 S2_34_39 ( .A(\ab[34][39] ), .B(\CARRYB[33][39] ), .CI(\SUMB[33][40] ), 
        .CO(\CARRYB[34][39] ), .S(\SUMB[34][39] ) );
  FA_X1 S2_34_40 ( .A(\ab[34][40] ), .B(\CARRYB[33][40] ), .CI(\SUMB[33][41] ), 
        .CO(\CARRYB[34][40] ), .S(\SUMB[34][40] ) );
  FA_X1 S2_34_41 ( .A(\ab[34][41] ), .B(\CARRYB[33][41] ), .CI(\SUMB[33][42] ), 
        .CO(\CARRYB[34][41] ), .S(\SUMB[34][41] ) );
  FA_X1 S2_34_42 ( .A(\ab[34][42] ), .B(\CARRYB[33][42] ), .CI(\SUMB[33][43] ), 
        .CO(\CARRYB[34][42] ), .S(\SUMB[34][42] ) );
  FA_X1 S2_34_43 ( .A(\ab[34][43] ), .B(\CARRYB[33][43] ), .CI(\SUMB[33][44] ), 
        .CO(\CARRYB[34][43] ), .S(\SUMB[34][43] ) );
  FA_X1 S2_34_44 ( .A(\ab[34][44] ), .B(\CARRYB[33][44] ), .CI(\SUMB[33][45] ), 
        .CO(\CARRYB[34][44] ), .S(\SUMB[34][44] ) );
  FA_X1 S2_34_45 ( .A(\ab[34][45] ), .B(\CARRYB[33][45] ), .CI(\SUMB[33][46] ), 
        .CO(\CARRYB[34][45] ), .S(\SUMB[34][45] ) );
  FA_X1 S2_34_46 ( .A(\ab[34][46] ), .B(\CARRYB[33][46] ), .CI(\SUMB[33][47] ), 
        .CO(\CARRYB[34][46] ), .S(\SUMB[34][46] ) );
  FA_X1 S2_34_47 ( .A(\ab[34][47] ), .B(\CARRYB[33][47] ), .CI(\SUMB[33][48] ), 
        .CO(\CARRYB[34][47] ), .S(\SUMB[34][47] ) );
  FA_X1 S2_34_48 ( .A(\ab[34][48] ), .B(\CARRYB[33][48] ), .CI(\SUMB[33][49] ), 
        .CO(\CARRYB[34][48] ), .S(\SUMB[34][48] ) );
  FA_X1 S2_34_49 ( .A(\ab[34][49] ), .B(\CARRYB[33][49] ), .CI(\SUMB[33][50] ), 
        .CO(\CARRYB[34][49] ), .S(\SUMB[34][49] ) );
  FA_X1 S2_34_50 ( .A(\ab[34][50] ), .B(\CARRYB[33][50] ), .CI(\SUMB[33][51] ), 
        .CO(\CARRYB[34][50] ), .S(\SUMB[34][50] ) );
  FA_X1 S3_34_51 ( .A(\ab[34][51] ), .B(\CARRYB[33][51] ), .CI(\ab[33][52] ), 
        .CO(\CARRYB[34][51] ), .S(\SUMB[34][51] ) );
  FA_X1 S1_33_0 ( .A(\ab[33][0] ), .B(\CARRYB[32][0] ), .CI(\SUMB[32][1] ), 
        .CO(\CARRYB[33][0] ), .S(CLA_SUM[33]) );
  FA_X1 S2_33_1 ( .A(\ab[33][1] ), .B(\CARRYB[32][1] ), .CI(\SUMB[32][2] ), 
        .CO(\CARRYB[33][1] ), .S(\SUMB[33][1] ) );
  FA_X1 S2_33_2 ( .A(\ab[33][2] ), .B(\CARRYB[32][2] ), .CI(\SUMB[32][3] ), 
        .CO(\CARRYB[33][2] ), .S(\SUMB[33][2] ) );
  FA_X1 S2_33_3 ( .A(\ab[33][3] ), .B(\CARRYB[32][3] ), .CI(\SUMB[32][4] ), 
        .CO(\CARRYB[33][3] ), .S(\SUMB[33][3] ) );
  FA_X1 S2_33_4 ( .A(\ab[33][4] ), .B(\CARRYB[32][4] ), .CI(\SUMB[32][5] ), 
        .CO(\CARRYB[33][4] ), .S(\SUMB[33][4] ) );
  FA_X1 S2_33_5 ( .A(\ab[33][5] ), .B(\CARRYB[32][5] ), .CI(\SUMB[32][6] ), 
        .CO(\CARRYB[33][5] ), .S(\SUMB[33][5] ) );
  FA_X1 S2_33_6 ( .A(\ab[33][6] ), .B(\CARRYB[32][6] ), .CI(\SUMB[32][7] ), 
        .CO(\CARRYB[33][6] ), .S(\SUMB[33][6] ) );
  FA_X1 S2_33_7 ( .A(\ab[33][7] ), .B(\CARRYB[32][7] ), .CI(\SUMB[32][8] ), 
        .CO(\CARRYB[33][7] ), .S(\SUMB[33][7] ) );
  FA_X1 S2_33_8 ( .A(\ab[33][8] ), .B(\CARRYB[32][8] ), .CI(\SUMB[32][9] ), 
        .CO(\CARRYB[33][8] ), .S(\SUMB[33][8] ) );
  FA_X1 S2_33_9 ( .A(\ab[33][9] ), .B(\CARRYB[32][9] ), .CI(\SUMB[32][10] ), 
        .CO(\CARRYB[33][9] ), .S(\SUMB[33][9] ) );
  FA_X1 S2_33_10 ( .A(\ab[33][10] ), .B(\CARRYB[32][10] ), .CI(\SUMB[32][11] ), 
        .CO(\CARRYB[33][10] ), .S(\SUMB[33][10] ) );
  FA_X1 S2_33_11 ( .A(\ab[33][11] ), .B(\CARRYB[32][11] ), .CI(\SUMB[32][12] ), 
        .CO(\CARRYB[33][11] ), .S(\SUMB[33][11] ) );
  FA_X1 S2_33_12 ( .A(\ab[33][12] ), .B(\CARRYB[32][12] ), .CI(\SUMB[32][13] ), 
        .CO(\CARRYB[33][12] ), .S(\SUMB[33][12] ) );
  FA_X1 S2_33_13 ( .A(\ab[33][13] ), .B(\CARRYB[32][13] ), .CI(\SUMB[32][14] ), 
        .CO(\CARRYB[33][13] ), .S(\SUMB[33][13] ) );
  FA_X1 S2_33_14 ( .A(\ab[33][14] ), .B(\CARRYB[32][14] ), .CI(\SUMB[32][15] ), 
        .CO(\CARRYB[33][14] ), .S(\SUMB[33][14] ) );
  FA_X1 S2_33_15 ( .A(\ab[33][15] ), .B(\CARRYB[32][15] ), .CI(\SUMB[32][16] ), 
        .CO(\CARRYB[33][15] ), .S(\SUMB[33][15] ) );
  FA_X1 S2_33_16 ( .A(\ab[33][16] ), .B(\CARRYB[32][16] ), .CI(\SUMB[32][17] ), 
        .CO(\CARRYB[33][16] ), .S(\SUMB[33][16] ) );
  FA_X1 S2_33_17 ( .A(\ab[33][17] ), .B(\CARRYB[32][17] ), .CI(\SUMB[32][18] ), 
        .CO(\CARRYB[33][17] ), .S(\SUMB[33][17] ) );
  FA_X1 S2_33_18 ( .A(\ab[33][18] ), .B(\CARRYB[32][18] ), .CI(\SUMB[32][19] ), 
        .CO(\CARRYB[33][18] ), .S(\SUMB[33][18] ) );
  FA_X1 S2_33_19 ( .A(\ab[33][19] ), .B(\CARRYB[32][19] ), .CI(\SUMB[32][20] ), 
        .CO(\CARRYB[33][19] ), .S(\SUMB[33][19] ) );
  FA_X1 S2_33_20 ( .A(\ab[33][20] ), .B(\CARRYB[32][20] ), .CI(\SUMB[32][21] ), 
        .CO(\CARRYB[33][20] ), .S(\SUMB[33][20] ) );
  FA_X1 S2_33_21 ( .A(\ab[33][21] ), .B(\CARRYB[32][21] ), .CI(\SUMB[32][22] ), 
        .CO(\CARRYB[33][21] ), .S(\SUMB[33][21] ) );
  FA_X1 S2_33_22 ( .A(\ab[33][22] ), .B(\CARRYB[32][22] ), .CI(\SUMB[32][23] ), 
        .CO(\CARRYB[33][22] ), .S(\SUMB[33][22] ) );
  FA_X1 S2_33_23 ( .A(\ab[33][23] ), .B(\CARRYB[32][23] ), .CI(\SUMB[32][24] ), 
        .CO(\CARRYB[33][23] ), .S(\SUMB[33][23] ) );
  FA_X1 S2_33_24 ( .A(\ab[33][24] ), .B(\CARRYB[32][24] ), .CI(\SUMB[32][25] ), 
        .CO(\CARRYB[33][24] ), .S(\SUMB[33][24] ) );
  FA_X1 S2_33_25 ( .A(\ab[33][25] ), .B(\CARRYB[32][25] ), .CI(\SUMB[32][26] ), 
        .CO(\CARRYB[33][25] ), .S(\SUMB[33][25] ) );
  FA_X1 S2_33_26 ( .A(\ab[33][26] ), .B(\CARRYB[32][26] ), .CI(\SUMB[32][27] ), 
        .CO(\CARRYB[33][26] ), .S(\SUMB[33][26] ) );
  FA_X1 S2_33_27 ( .A(\ab[33][27] ), .B(\CARRYB[32][27] ), .CI(\SUMB[32][28] ), 
        .CO(\CARRYB[33][27] ), .S(\SUMB[33][27] ) );
  FA_X1 S2_33_28 ( .A(\ab[33][28] ), .B(\CARRYB[32][28] ), .CI(\SUMB[32][29] ), 
        .CO(\CARRYB[33][28] ), .S(\SUMB[33][28] ) );
  FA_X1 S2_33_29 ( .A(\ab[33][29] ), .B(\CARRYB[32][29] ), .CI(\SUMB[32][30] ), 
        .CO(\CARRYB[33][29] ), .S(\SUMB[33][29] ) );
  FA_X1 S2_33_30 ( .A(\ab[33][30] ), .B(\CARRYB[32][30] ), .CI(\SUMB[32][31] ), 
        .CO(\CARRYB[33][30] ), .S(\SUMB[33][30] ) );
  FA_X1 S2_33_31 ( .A(\ab[33][31] ), .B(\CARRYB[32][31] ), .CI(\SUMB[32][32] ), 
        .CO(\CARRYB[33][31] ), .S(\SUMB[33][31] ) );
  FA_X1 S2_33_32 ( .A(\ab[33][32] ), .B(\CARRYB[32][32] ), .CI(\SUMB[32][33] ), 
        .CO(\CARRYB[33][32] ), .S(\SUMB[33][32] ) );
  FA_X1 S2_33_33 ( .A(\ab[33][33] ), .B(\CARRYB[32][33] ), .CI(\SUMB[32][34] ), 
        .CO(\CARRYB[33][33] ), .S(\SUMB[33][33] ) );
  FA_X1 S2_33_34 ( .A(\ab[33][34] ), .B(\CARRYB[32][34] ), .CI(\SUMB[32][35] ), 
        .CO(\CARRYB[33][34] ), .S(\SUMB[33][34] ) );
  FA_X1 S2_33_35 ( .A(\ab[33][35] ), .B(\CARRYB[32][35] ), .CI(\SUMB[32][36] ), 
        .CO(\CARRYB[33][35] ), .S(\SUMB[33][35] ) );
  FA_X1 S2_33_36 ( .A(\ab[33][36] ), .B(\CARRYB[32][36] ), .CI(\SUMB[32][37] ), 
        .CO(\CARRYB[33][36] ), .S(\SUMB[33][36] ) );
  FA_X1 S2_33_37 ( .A(\ab[33][37] ), .B(\CARRYB[32][37] ), .CI(\SUMB[32][38] ), 
        .CO(\CARRYB[33][37] ), .S(\SUMB[33][37] ) );
  FA_X1 S2_33_38 ( .A(\ab[33][38] ), .B(\CARRYB[32][38] ), .CI(\SUMB[32][39] ), 
        .CO(\CARRYB[33][38] ), .S(\SUMB[33][38] ) );
  FA_X1 S2_33_39 ( .A(\ab[33][39] ), .B(\CARRYB[32][39] ), .CI(\SUMB[32][40] ), 
        .CO(\CARRYB[33][39] ), .S(\SUMB[33][39] ) );
  FA_X1 S2_33_40 ( .A(\ab[33][40] ), .B(\CARRYB[32][40] ), .CI(\SUMB[32][41] ), 
        .CO(\CARRYB[33][40] ), .S(\SUMB[33][40] ) );
  FA_X1 S2_33_41 ( .A(\ab[33][41] ), .B(\CARRYB[32][41] ), .CI(\SUMB[32][42] ), 
        .CO(\CARRYB[33][41] ), .S(\SUMB[33][41] ) );
  FA_X1 S2_33_42 ( .A(\ab[33][42] ), .B(\CARRYB[32][42] ), .CI(\SUMB[32][43] ), 
        .CO(\CARRYB[33][42] ), .S(\SUMB[33][42] ) );
  FA_X1 S2_33_43 ( .A(\ab[33][43] ), .B(\CARRYB[32][43] ), .CI(\SUMB[32][44] ), 
        .CO(\CARRYB[33][43] ), .S(\SUMB[33][43] ) );
  FA_X1 S2_33_44 ( .A(\ab[33][44] ), .B(\CARRYB[32][44] ), .CI(\SUMB[32][45] ), 
        .CO(\CARRYB[33][44] ), .S(\SUMB[33][44] ) );
  FA_X1 S2_33_45 ( .A(\ab[33][45] ), .B(\CARRYB[32][45] ), .CI(\SUMB[32][46] ), 
        .CO(\CARRYB[33][45] ), .S(\SUMB[33][45] ) );
  FA_X1 S2_33_46 ( .A(\ab[33][46] ), .B(\CARRYB[32][46] ), .CI(\SUMB[32][47] ), 
        .CO(\CARRYB[33][46] ), .S(\SUMB[33][46] ) );
  FA_X1 S2_33_47 ( .A(\ab[33][47] ), .B(\CARRYB[32][47] ), .CI(\SUMB[32][48] ), 
        .CO(\CARRYB[33][47] ), .S(\SUMB[33][47] ) );
  FA_X1 S2_33_48 ( .A(\ab[33][48] ), .B(\CARRYB[32][48] ), .CI(\SUMB[32][49] ), 
        .CO(\CARRYB[33][48] ), .S(\SUMB[33][48] ) );
  FA_X1 S2_33_49 ( .A(\ab[33][49] ), .B(\CARRYB[32][49] ), .CI(\SUMB[32][50] ), 
        .CO(\CARRYB[33][49] ), .S(\SUMB[33][49] ) );
  FA_X1 S2_33_50 ( .A(\ab[33][50] ), .B(\CARRYB[32][50] ), .CI(\SUMB[32][51] ), 
        .CO(\CARRYB[33][50] ), .S(\SUMB[33][50] ) );
  FA_X1 S3_33_51 ( .A(\ab[33][51] ), .B(\CARRYB[32][51] ), .CI(\ab[32][52] ), 
        .CO(\CARRYB[33][51] ), .S(\SUMB[33][51] ) );
  FA_X1 S1_32_0 ( .A(\ab[32][0] ), .B(\CARRYB[31][0] ), .CI(\SUMB[31][1] ), 
        .CO(\CARRYB[32][0] ), .S(CLA_SUM[32]) );
  FA_X1 S2_32_1 ( .A(\ab[32][1] ), .B(\CARRYB[31][1] ), .CI(\SUMB[31][2] ), 
        .CO(\CARRYB[32][1] ), .S(\SUMB[32][1] ) );
  FA_X1 S2_32_2 ( .A(\ab[32][2] ), .B(\CARRYB[31][2] ), .CI(\SUMB[31][3] ), 
        .CO(\CARRYB[32][2] ), .S(\SUMB[32][2] ) );
  FA_X1 S2_32_3 ( .A(\ab[32][3] ), .B(\CARRYB[31][3] ), .CI(\SUMB[31][4] ), 
        .CO(\CARRYB[32][3] ), .S(\SUMB[32][3] ) );
  FA_X1 S2_32_4 ( .A(\ab[32][4] ), .B(\CARRYB[31][4] ), .CI(\SUMB[31][5] ), 
        .CO(\CARRYB[32][4] ), .S(\SUMB[32][4] ) );
  FA_X1 S2_32_5 ( .A(\ab[32][5] ), .B(\CARRYB[31][5] ), .CI(\SUMB[31][6] ), 
        .CO(\CARRYB[32][5] ), .S(\SUMB[32][5] ) );
  FA_X1 S2_32_6 ( .A(\ab[32][6] ), .B(\CARRYB[31][6] ), .CI(\SUMB[31][7] ), 
        .CO(\CARRYB[32][6] ), .S(\SUMB[32][6] ) );
  FA_X1 S2_32_7 ( .A(\ab[32][7] ), .B(\CARRYB[31][7] ), .CI(\SUMB[31][8] ), 
        .CO(\CARRYB[32][7] ), .S(\SUMB[32][7] ) );
  FA_X1 S2_32_8 ( .A(\ab[32][8] ), .B(\CARRYB[31][8] ), .CI(\SUMB[31][9] ), 
        .CO(\CARRYB[32][8] ), .S(\SUMB[32][8] ) );
  FA_X1 S2_32_9 ( .A(\ab[32][9] ), .B(\CARRYB[31][9] ), .CI(\SUMB[31][10] ), 
        .CO(\CARRYB[32][9] ), .S(\SUMB[32][9] ) );
  FA_X1 S2_32_10 ( .A(\ab[32][10] ), .B(\CARRYB[31][10] ), .CI(\SUMB[31][11] ), 
        .CO(\CARRYB[32][10] ), .S(\SUMB[32][10] ) );
  FA_X1 S2_32_11 ( .A(\ab[32][11] ), .B(\CARRYB[31][11] ), .CI(\SUMB[31][12] ), 
        .CO(\CARRYB[32][11] ), .S(\SUMB[32][11] ) );
  FA_X1 S2_32_12 ( .A(\ab[32][12] ), .B(\CARRYB[31][12] ), .CI(\SUMB[31][13] ), 
        .CO(\CARRYB[32][12] ), .S(\SUMB[32][12] ) );
  FA_X1 S2_32_13 ( .A(\ab[32][13] ), .B(\CARRYB[31][13] ), .CI(\SUMB[31][14] ), 
        .CO(\CARRYB[32][13] ), .S(\SUMB[32][13] ) );
  FA_X1 S2_32_14 ( .A(\ab[32][14] ), .B(\CARRYB[31][14] ), .CI(\SUMB[31][15] ), 
        .CO(\CARRYB[32][14] ), .S(\SUMB[32][14] ) );
  FA_X1 S2_32_15 ( .A(\ab[32][15] ), .B(\CARRYB[31][15] ), .CI(\SUMB[31][16] ), 
        .CO(\CARRYB[32][15] ), .S(\SUMB[32][15] ) );
  FA_X1 S2_32_16 ( .A(\ab[32][16] ), .B(\CARRYB[31][16] ), .CI(\SUMB[31][17] ), 
        .CO(\CARRYB[32][16] ), .S(\SUMB[32][16] ) );
  FA_X1 S2_32_17 ( .A(\ab[32][17] ), .B(\CARRYB[31][17] ), .CI(\SUMB[31][18] ), 
        .CO(\CARRYB[32][17] ), .S(\SUMB[32][17] ) );
  FA_X1 S2_32_18 ( .A(\ab[32][18] ), .B(\CARRYB[31][18] ), .CI(\SUMB[31][19] ), 
        .CO(\CARRYB[32][18] ), .S(\SUMB[32][18] ) );
  FA_X1 S2_32_19 ( .A(\ab[32][19] ), .B(\CARRYB[31][19] ), .CI(\SUMB[31][20] ), 
        .CO(\CARRYB[32][19] ), .S(\SUMB[32][19] ) );
  FA_X1 S2_32_20 ( .A(\ab[32][20] ), .B(\CARRYB[31][20] ), .CI(\SUMB[31][21] ), 
        .CO(\CARRYB[32][20] ), .S(\SUMB[32][20] ) );
  FA_X1 S2_32_21 ( .A(\ab[32][21] ), .B(\CARRYB[31][21] ), .CI(\SUMB[31][22] ), 
        .CO(\CARRYB[32][21] ), .S(\SUMB[32][21] ) );
  FA_X1 S2_32_22 ( .A(\ab[32][22] ), .B(\CARRYB[31][22] ), .CI(\SUMB[31][23] ), 
        .CO(\CARRYB[32][22] ), .S(\SUMB[32][22] ) );
  FA_X1 S2_32_23 ( .A(\ab[32][23] ), .B(\CARRYB[31][23] ), .CI(\SUMB[31][24] ), 
        .CO(\CARRYB[32][23] ), .S(\SUMB[32][23] ) );
  FA_X1 S2_32_24 ( .A(\ab[32][24] ), .B(\CARRYB[31][24] ), .CI(\SUMB[31][25] ), 
        .CO(\CARRYB[32][24] ), .S(\SUMB[32][24] ) );
  FA_X1 S2_32_25 ( .A(\ab[32][25] ), .B(\CARRYB[31][25] ), .CI(\SUMB[31][26] ), 
        .CO(\CARRYB[32][25] ), .S(\SUMB[32][25] ) );
  FA_X1 S2_32_26 ( .A(\ab[32][26] ), .B(\CARRYB[31][26] ), .CI(\SUMB[31][27] ), 
        .CO(\CARRYB[32][26] ), .S(\SUMB[32][26] ) );
  FA_X1 S2_32_27 ( .A(\ab[32][27] ), .B(\CARRYB[31][27] ), .CI(\SUMB[31][28] ), 
        .CO(\CARRYB[32][27] ), .S(\SUMB[32][27] ) );
  FA_X1 S2_32_28 ( .A(\ab[32][28] ), .B(\CARRYB[31][28] ), .CI(\SUMB[31][29] ), 
        .CO(\CARRYB[32][28] ), .S(\SUMB[32][28] ) );
  FA_X1 S2_32_29 ( .A(\ab[32][29] ), .B(\CARRYB[31][29] ), .CI(\SUMB[31][30] ), 
        .CO(\CARRYB[32][29] ), .S(\SUMB[32][29] ) );
  FA_X1 S2_32_30 ( .A(\ab[32][30] ), .B(\CARRYB[31][30] ), .CI(\SUMB[31][31] ), 
        .CO(\CARRYB[32][30] ), .S(\SUMB[32][30] ) );
  FA_X1 S2_32_31 ( .A(\ab[32][31] ), .B(\CARRYB[31][31] ), .CI(\SUMB[31][32] ), 
        .CO(\CARRYB[32][31] ), .S(\SUMB[32][31] ) );
  FA_X1 S2_32_32 ( .A(\ab[32][32] ), .B(\CARRYB[31][32] ), .CI(\SUMB[31][33] ), 
        .CO(\CARRYB[32][32] ), .S(\SUMB[32][32] ) );
  FA_X1 S2_32_33 ( .A(\ab[32][33] ), .B(\CARRYB[31][33] ), .CI(\SUMB[31][34] ), 
        .CO(\CARRYB[32][33] ), .S(\SUMB[32][33] ) );
  FA_X1 S2_32_34 ( .A(\ab[32][34] ), .B(\CARRYB[31][34] ), .CI(\SUMB[31][35] ), 
        .CO(\CARRYB[32][34] ), .S(\SUMB[32][34] ) );
  FA_X1 S2_32_35 ( .A(\ab[32][35] ), .B(\CARRYB[31][35] ), .CI(\SUMB[31][36] ), 
        .CO(\CARRYB[32][35] ), .S(\SUMB[32][35] ) );
  FA_X1 S2_32_36 ( .A(\ab[32][36] ), .B(\CARRYB[31][36] ), .CI(\SUMB[31][37] ), 
        .CO(\CARRYB[32][36] ), .S(\SUMB[32][36] ) );
  FA_X1 S2_32_37 ( .A(\ab[32][37] ), .B(\CARRYB[31][37] ), .CI(\SUMB[31][38] ), 
        .CO(\CARRYB[32][37] ), .S(\SUMB[32][37] ) );
  FA_X1 S2_32_38 ( .A(\ab[32][38] ), .B(\CARRYB[31][38] ), .CI(\SUMB[31][39] ), 
        .CO(\CARRYB[32][38] ), .S(\SUMB[32][38] ) );
  FA_X1 S2_32_39 ( .A(\ab[32][39] ), .B(\CARRYB[31][39] ), .CI(\SUMB[31][40] ), 
        .CO(\CARRYB[32][39] ), .S(\SUMB[32][39] ) );
  FA_X1 S2_32_40 ( .A(\ab[32][40] ), .B(\CARRYB[31][40] ), .CI(\SUMB[31][41] ), 
        .CO(\CARRYB[32][40] ), .S(\SUMB[32][40] ) );
  FA_X1 S2_32_41 ( .A(\ab[32][41] ), .B(\CARRYB[31][41] ), .CI(\SUMB[31][42] ), 
        .CO(\CARRYB[32][41] ), .S(\SUMB[32][41] ) );
  FA_X1 S2_32_42 ( .A(\ab[32][42] ), .B(\CARRYB[31][42] ), .CI(\SUMB[31][43] ), 
        .CO(\CARRYB[32][42] ), .S(\SUMB[32][42] ) );
  FA_X1 S2_32_43 ( .A(\ab[32][43] ), .B(\CARRYB[31][43] ), .CI(\SUMB[31][44] ), 
        .CO(\CARRYB[32][43] ), .S(\SUMB[32][43] ) );
  FA_X1 S2_32_44 ( .A(\ab[32][44] ), .B(\CARRYB[31][44] ), .CI(\SUMB[31][45] ), 
        .CO(\CARRYB[32][44] ), .S(\SUMB[32][44] ) );
  FA_X1 S2_32_45 ( .A(\ab[32][45] ), .B(\CARRYB[31][45] ), .CI(\SUMB[31][46] ), 
        .CO(\CARRYB[32][45] ), .S(\SUMB[32][45] ) );
  FA_X1 S2_32_46 ( .A(\ab[32][46] ), .B(\CARRYB[31][46] ), .CI(\SUMB[31][47] ), 
        .CO(\CARRYB[32][46] ), .S(\SUMB[32][46] ) );
  FA_X1 S2_32_47 ( .A(\ab[32][47] ), .B(\CARRYB[31][47] ), .CI(\SUMB[31][48] ), 
        .CO(\CARRYB[32][47] ), .S(\SUMB[32][47] ) );
  FA_X1 S2_32_48 ( .A(\ab[32][48] ), .B(\CARRYB[31][48] ), .CI(\SUMB[31][49] ), 
        .CO(\CARRYB[32][48] ), .S(\SUMB[32][48] ) );
  FA_X1 S2_32_49 ( .A(\ab[32][49] ), .B(\CARRYB[31][49] ), .CI(\SUMB[31][50] ), 
        .CO(\CARRYB[32][49] ), .S(\SUMB[32][49] ) );
  FA_X1 S2_32_50 ( .A(\ab[32][50] ), .B(\CARRYB[31][50] ), .CI(\SUMB[31][51] ), 
        .CO(\CARRYB[32][50] ), .S(\SUMB[32][50] ) );
  FA_X1 S3_32_51 ( .A(\ab[32][51] ), .B(\CARRYB[31][51] ), .CI(\ab[31][52] ), 
        .CO(\CARRYB[32][51] ), .S(\SUMB[32][51] ) );
  FA_X1 S1_31_0 ( .A(\ab[31][0] ), .B(\CARRYB[30][0] ), .CI(\SUMB[30][1] ), 
        .CO(\CARRYB[31][0] ), .S(CLA_SUM[31]) );
  FA_X1 S2_31_1 ( .A(\ab[31][1] ), .B(\CARRYB[30][1] ), .CI(\SUMB[30][2] ), 
        .CO(\CARRYB[31][1] ), .S(\SUMB[31][1] ) );
  FA_X1 S2_31_2 ( .A(\ab[31][2] ), .B(\CARRYB[30][2] ), .CI(\SUMB[30][3] ), 
        .CO(\CARRYB[31][2] ), .S(\SUMB[31][2] ) );
  FA_X1 S2_31_3 ( .A(\ab[31][3] ), .B(\CARRYB[30][3] ), .CI(\SUMB[30][4] ), 
        .CO(\CARRYB[31][3] ), .S(\SUMB[31][3] ) );
  FA_X1 S2_31_4 ( .A(\ab[31][4] ), .B(\CARRYB[30][4] ), .CI(\SUMB[30][5] ), 
        .CO(\CARRYB[31][4] ), .S(\SUMB[31][4] ) );
  FA_X1 S2_31_5 ( .A(\ab[31][5] ), .B(\CARRYB[30][5] ), .CI(\SUMB[30][6] ), 
        .CO(\CARRYB[31][5] ), .S(\SUMB[31][5] ) );
  FA_X1 S2_31_6 ( .A(\ab[31][6] ), .B(\CARRYB[30][6] ), .CI(\SUMB[30][7] ), 
        .CO(\CARRYB[31][6] ), .S(\SUMB[31][6] ) );
  FA_X1 S2_31_7 ( .A(\ab[31][7] ), .B(\CARRYB[30][7] ), .CI(\SUMB[30][8] ), 
        .CO(\CARRYB[31][7] ), .S(\SUMB[31][7] ) );
  FA_X1 S2_31_8 ( .A(\ab[31][8] ), .B(\CARRYB[30][8] ), .CI(\SUMB[30][9] ), 
        .CO(\CARRYB[31][8] ), .S(\SUMB[31][8] ) );
  FA_X1 S2_31_9 ( .A(\ab[31][9] ), .B(\CARRYB[30][9] ), .CI(\SUMB[30][10] ), 
        .CO(\CARRYB[31][9] ), .S(\SUMB[31][9] ) );
  FA_X1 S2_31_10 ( .A(\ab[31][10] ), .B(\CARRYB[30][10] ), .CI(\SUMB[30][11] ), 
        .CO(\CARRYB[31][10] ), .S(\SUMB[31][10] ) );
  FA_X1 S2_31_11 ( .A(\ab[31][11] ), .B(\CARRYB[30][11] ), .CI(\SUMB[30][12] ), 
        .CO(\CARRYB[31][11] ), .S(\SUMB[31][11] ) );
  FA_X1 S2_31_12 ( .A(\ab[31][12] ), .B(\CARRYB[30][12] ), .CI(\SUMB[30][13] ), 
        .CO(\CARRYB[31][12] ), .S(\SUMB[31][12] ) );
  FA_X1 S2_31_13 ( .A(\ab[31][13] ), .B(\CARRYB[30][13] ), .CI(\SUMB[30][14] ), 
        .CO(\CARRYB[31][13] ), .S(\SUMB[31][13] ) );
  FA_X1 S2_31_14 ( .A(\ab[31][14] ), .B(\CARRYB[30][14] ), .CI(\SUMB[30][15] ), 
        .CO(\CARRYB[31][14] ), .S(\SUMB[31][14] ) );
  FA_X1 S2_31_15 ( .A(\ab[31][15] ), .B(\CARRYB[30][15] ), .CI(\SUMB[30][16] ), 
        .CO(\CARRYB[31][15] ), .S(\SUMB[31][15] ) );
  FA_X1 S2_31_16 ( .A(\ab[31][16] ), .B(\CARRYB[30][16] ), .CI(\SUMB[30][17] ), 
        .CO(\CARRYB[31][16] ), .S(\SUMB[31][16] ) );
  FA_X1 S2_31_17 ( .A(\ab[31][17] ), .B(\CARRYB[30][17] ), .CI(\SUMB[30][18] ), 
        .CO(\CARRYB[31][17] ), .S(\SUMB[31][17] ) );
  FA_X1 S2_31_18 ( .A(\ab[31][18] ), .B(\CARRYB[30][18] ), .CI(\SUMB[30][19] ), 
        .CO(\CARRYB[31][18] ), .S(\SUMB[31][18] ) );
  FA_X1 S2_31_19 ( .A(\ab[31][19] ), .B(\CARRYB[30][19] ), .CI(\SUMB[30][20] ), 
        .CO(\CARRYB[31][19] ), .S(\SUMB[31][19] ) );
  FA_X1 S2_31_20 ( .A(\ab[31][20] ), .B(\CARRYB[30][20] ), .CI(\SUMB[30][21] ), 
        .CO(\CARRYB[31][20] ), .S(\SUMB[31][20] ) );
  FA_X1 S2_31_21 ( .A(\ab[31][21] ), .B(\CARRYB[30][21] ), .CI(\SUMB[30][22] ), 
        .CO(\CARRYB[31][21] ), .S(\SUMB[31][21] ) );
  FA_X1 S2_31_22 ( .A(\ab[31][22] ), .B(\CARRYB[30][22] ), .CI(\SUMB[30][23] ), 
        .CO(\CARRYB[31][22] ), .S(\SUMB[31][22] ) );
  FA_X1 S2_31_23 ( .A(\ab[31][23] ), .B(\CARRYB[30][23] ), .CI(\SUMB[30][24] ), 
        .CO(\CARRYB[31][23] ), .S(\SUMB[31][23] ) );
  FA_X1 S2_31_24 ( .A(\ab[31][24] ), .B(\CARRYB[30][24] ), .CI(\SUMB[30][25] ), 
        .CO(\CARRYB[31][24] ), .S(\SUMB[31][24] ) );
  FA_X1 S2_31_25 ( .A(\ab[31][25] ), .B(\CARRYB[30][25] ), .CI(\SUMB[30][26] ), 
        .CO(\CARRYB[31][25] ), .S(\SUMB[31][25] ) );
  FA_X1 S2_31_26 ( .A(\ab[31][26] ), .B(\CARRYB[30][26] ), .CI(\SUMB[30][27] ), 
        .CO(\CARRYB[31][26] ), .S(\SUMB[31][26] ) );
  FA_X1 S2_31_27 ( .A(\ab[31][27] ), .B(\CARRYB[30][27] ), .CI(\SUMB[30][28] ), 
        .CO(\CARRYB[31][27] ), .S(\SUMB[31][27] ) );
  FA_X1 S2_31_28 ( .A(\ab[31][28] ), .B(\CARRYB[30][28] ), .CI(\SUMB[30][29] ), 
        .CO(\CARRYB[31][28] ), .S(\SUMB[31][28] ) );
  FA_X1 S2_31_29 ( .A(\ab[31][29] ), .B(\CARRYB[30][29] ), .CI(\SUMB[30][30] ), 
        .CO(\CARRYB[31][29] ), .S(\SUMB[31][29] ) );
  FA_X1 S2_31_30 ( .A(\ab[31][30] ), .B(\CARRYB[30][30] ), .CI(\SUMB[30][31] ), 
        .CO(\CARRYB[31][30] ), .S(\SUMB[31][30] ) );
  FA_X1 S2_31_31 ( .A(\ab[31][31] ), .B(\CARRYB[30][31] ), .CI(\SUMB[30][32] ), 
        .CO(\CARRYB[31][31] ), .S(\SUMB[31][31] ) );
  FA_X1 S2_31_32 ( .A(\ab[31][32] ), .B(\CARRYB[30][32] ), .CI(\SUMB[30][33] ), 
        .CO(\CARRYB[31][32] ), .S(\SUMB[31][32] ) );
  FA_X1 S2_31_33 ( .A(\ab[31][33] ), .B(\CARRYB[30][33] ), .CI(\SUMB[30][34] ), 
        .CO(\CARRYB[31][33] ), .S(\SUMB[31][33] ) );
  FA_X1 S2_31_34 ( .A(\ab[31][34] ), .B(\CARRYB[30][34] ), .CI(\SUMB[30][35] ), 
        .CO(\CARRYB[31][34] ), .S(\SUMB[31][34] ) );
  FA_X1 S2_31_35 ( .A(\ab[31][35] ), .B(\CARRYB[30][35] ), .CI(\SUMB[30][36] ), 
        .CO(\CARRYB[31][35] ), .S(\SUMB[31][35] ) );
  FA_X1 S2_31_36 ( .A(\ab[31][36] ), .B(\CARRYB[30][36] ), .CI(\SUMB[30][37] ), 
        .CO(\CARRYB[31][36] ), .S(\SUMB[31][36] ) );
  FA_X1 S2_31_37 ( .A(\ab[31][37] ), .B(\CARRYB[30][37] ), .CI(\SUMB[30][38] ), 
        .CO(\CARRYB[31][37] ), .S(\SUMB[31][37] ) );
  FA_X1 S2_31_38 ( .A(\ab[31][38] ), .B(\CARRYB[30][38] ), .CI(\SUMB[30][39] ), 
        .CO(\CARRYB[31][38] ), .S(\SUMB[31][38] ) );
  FA_X1 S2_31_39 ( .A(\ab[31][39] ), .B(\CARRYB[30][39] ), .CI(\SUMB[30][40] ), 
        .CO(\CARRYB[31][39] ), .S(\SUMB[31][39] ) );
  FA_X1 S2_31_40 ( .A(\ab[31][40] ), .B(\CARRYB[30][40] ), .CI(\SUMB[30][41] ), 
        .CO(\CARRYB[31][40] ), .S(\SUMB[31][40] ) );
  FA_X1 S2_31_41 ( .A(\ab[31][41] ), .B(\CARRYB[30][41] ), .CI(\SUMB[30][42] ), 
        .CO(\CARRYB[31][41] ), .S(\SUMB[31][41] ) );
  FA_X1 S2_31_42 ( .A(\ab[31][42] ), .B(\CARRYB[30][42] ), .CI(\SUMB[30][43] ), 
        .CO(\CARRYB[31][42] ), .S(\SUMB[31][42] ) );
  FA_X1 S2_31_43 ( .A(\ab[31][43] ), .B(\CARRYB[30][43] ), .CI(\SUMB[30][44] ), 
        .CO(\CARRYB[31][43] ), .S(\SUMB[31][43] ) );
  FA_X1 S2_31_44 ( .A(\ab[31][44] ), .B(\CARRYB[30][44] ), .CI(\SUMB[30][45] ), 
        .CO(\CARRYB[31][44] ), .S(\SUMB[31][44] ) );
  FA_X1 S2_31_45 ( .A(\ab[31][45] ), .B(\CARRYB[30][45] ), .CI(\SUMB[30][46] ), 
        .CO(\CARRYB[31][45] ), .S(\SUMB[31][45] ) );
  FA_X1 S2_31_46 ( .A(\ab[31][46] ), .B(\CARRYB[30][46] ), .CI(\SUMB[30][47] ), 
        .CO(\CARRYB[31][46] ), .S(\SUMB[31][46] ) );
  FA_X1 S2_31_47 ( .A(\ab[31][47] ), .B(\CARRYB[30][47] ), .CI(\SUMB[30][48] ), 
        .CO(\CARRYB[31][47] ), .S(\SUMB[31][47] ) );
  FA_X1 S2_31_48 ( .A(\ab[31][48] ), .B(\CARRYB[30][48] ), .CI(\SUMB[30][49] ), 
        .CO(\CARRYB[31][48] ), .S(\SUMB[31][48] ) );
  FA_X1 S2_31_49 ( .A(\ab[31][49] ), .B(\CARRYB[30][49] ), .CI(\SUMB[30][50] ), 
        .CO(\CARRYB[31][49] ), .S(\SUMB[31][49] ) );
  FA_X1 S2_31_50 ( .A(\ab[31][50] ), .B(\CARRYB[30][50] ), .CI(\SUMB[30][51] ), 
        .CO(\CARRYB[31][50] ), .S(\SUMB[31][50] ) );
  FA_X1 S3_31_51 ( .A(\ab[31][51] ), .B(\CARRYB[30][51] ), .CI(\ab[30][52] ), 
        .CO(\CARRYB[31][51] ), .S(\SUMB[31][51] ) );
  FA_X1 S1_30_0 ( .A(\ab[30][0] ), .B(\CARRYB[29][0] ), .CI(\SUMB[29][1] ), 
        .CO(\CARRYB[30][0] ), .S(CLA_SUM[30]) );
  FA_X1 S2_30_1 ( .A(\ab[30][1] ), .B(\CARRYB[29][1] ), .CI(\SUMB[29][2] ), 
        .CO(\CARRYB[30][1] ), .S(\SUMB[30][1] ) );
  FA_X1 S2_30_2 ( .A(\ab[30][2] ), .B(\CARRYB[29][2] ), .CI(\SUMB[29][3] ), 
        .CO(\CARRYB[30][2] ), .S(\SUMB[30][2] ) );
  FA_X1 S2_30_3 ( .A(\ab[30][3] ), .B(\CARRYB[29][3] ), .CI(\SUMB[29][4] ), 
        .CO(\CARRYB[30][3] ), .S(\SUMB[30][3] ) );
  FA_X1 S2_30_4 ( .A(\ab[30][4] ), .B(\CARRYB[29][4] ), .CI(\SUMB[29][5] ), 
        .CO(\CARRYB[30][4] ), .S(\SUMB[30][4] ) );
  FA_X1 S2_30_5 ( .A(\ab[30][5] ), .B(\CARRYB[29][5] ), .CI(\SUMB[29][6] ), 
        .CO(\CARRYB[30][5] ), .S(\SUMB[30][5] ) );
  FA_X1 S2_30_6 ( .A(\ab[30][6] ), .B(\CARRYB[29][6] ), .CI(\SUMB[29][7] ), 
        .CO(\CARRYB[30][6] ), .S(\SUMB[30][6] ) );
  FA_X1 S2_30_7 ( .A(\ab[30][7] ), .B(\CARRYB[29][7] ), .CI(\SUMB[29][8] ), 
        .CO(\CARRYB[30][7] ), .S(\SUMB[30][7] ) );
  FA_X1 S2_30_8 ( .A(\ab[30][8] ), .B(\CARRYB[29][8] ), .CI(\SUMB[29][9] ), 
        .CO(\CARRYB[30][8] ), .S(\SUMB[30][8] ) );
  FA_X1 S2_30_9 ( .A(\ab[30][9] ), .B(\CARRYB[29][9] ), .CI(\SUMB[29][10] ), 
        .CO(\CARRYB[30][9] ), .S(\SUMB[30][9] ) );
  FA_X1 S2_30_10 ( .A(\ab[30][10] ), .B(\CARRYB[29][10] ), .CI(\SUMB[29][11] ), 
        .CO(\CARRYB[30][10] ), .S(\SUMB[30][10] ) );
  FA_X1 S2_30_11 ( .A(\ab[30][11] ), .B(\CARRYB[29][11] ), .CI(\SUMB[29][12] ), 
        .CO(\CARRYB[30][11] ), .S(\SUMB[30][11] ) );
  FA_X1 S2_30_12 ( .A(\ab[30][12] ), .B(\CARRYB[29][12] ), .CI(\SUMB[29][13] ), 
        .CO(\CARRYB[30][12] ), .S(\SUMB[30][12] ) );
  FA_X1 S2_30_13 ( .A(\ab[30][13] ), .B(\CARRYB[29][13] ), .CI(\SUMB[29][14] ), 
        .CO(\CARRYB[30][13] ), .S(\SUMB[30][13] ) );
  FA_X1 S2_30_14 ( .A(\ab[30][14] ), .B(\CARRYB[29][14] ), .CI(\SUMB[29][15] ), 
        .CO(\CARRYB[30][14] ), .S(\SUMB[30][14] ) );
  FA_X1 S2_30_15 ( .A(\ab[30][15] ), .B(\CARRYB[29][15] ), .CI(\SUMB[29][16] ), 
        .CO(\CARRYB[30][15] ), .S(\SUMB[30][15] ) );
  FA_X1 S2_30_16 ( .A(\ab[30][16] ), .B(\CARRYB[29][16] ), .CI(\SUMB[29][17] ), 
        .CO(\CARRYB[30][16] ), .S(\SUMB[30][16] ) );
  FA_X1 S2_30_17 ( .A(\ab[30][17] ), .B(\CARRYB[29][17] ), .CI(\SUMB[29][18] ), 
        .CO(\CARRYB[30][17] ), .S(\SUMB[30][17] ) );
  FA_X1 S2_30_18 ( .A(\ab[30][18] ), .B(\CARRYB[29][18] ), .CI(\SUMB[29][19] ), 
        .CO(\CARRYB[30][18] ), .S(\SUMB[30][18] ) );
  FA_X1 S2_30_19 ( .A(\ab[30][19] ), .B(\CARRYB[29][19] ), .CI(\SUMB[29][20] ), 
        .CO(\CARRYB[30][19] ), .S(\SUMB[30][19] ) );
  FA_X1 S2_30_20 ( .A(\ab[30][20] ), .B(\CARRYB[29][20] ), .CI(\SUMB[29][21] ), 
        .CO(\CARRYB[30][20] ), .S(\SUMB[30][20] ) );
  FA_X1 S2_30_21 ( .A(\ab[30][21] ), .B(\CARRYB[29][21] ), .CI(\SUMB[29][22] ), 
        .CO(\CARRYB[30][21] ), .S(\SUMB[30][21] ) );
  FA_X1 S2_30_22 ( .A(\ab[30][22] ), .B(\CARRYB[29][22] ), .CI(\SUMB[29][23] ), 
        .CO(\CARRYB[30][22] ), .S(\SUMB[30][22] ) );
  FA_X1 S2_30_23 ( .A(\ab[30][23] ), .B(\CARRYB[29][23] ), .CI(\SUMB[29][24] ), 
        .CO(\CARRYB[30][23] ), .S(\SUMB[30][23] ) );
  FA_X1 S2_30_24 ( .A(\ab[30][24] ), .B(\CARRYB[29][24] ), .CI(\SUMB[29][25] ), 
        .CO(\CARRYB[30][24] ), .S(\SUMB[30][24] ) );
  FA_X1 S2_30_25 ( .A(\ab[30][25] ), .B(\CARRYB[29][25] ), .CI(\SUMB[29][26] ), 
        .CO(\CARRYB[30][25] ), .S(\SUMB[30][25] ) );
  FA_X1 S2_30_26 ( .A(\ab[30][26] ), .B(\CARRYB[29][26] ), .CI(\SUMB[29][27] ), 
        .CO(\CARRYB[30][26] ), .S(\SUMB[30][26] ) );
  FA_X1 S2_30_27 ( .A(\ab[30][27] ), .B(\CARRYB[29][27] ), .CI(\SUMB[29][28] ), 
        .CO(\CARRYB[30][27] ), .S(\SUMB[30][27] ) );
  FA_X1 S2_30_28 ( .A(\ab[30][28] ), .B(\CARRYB[29][28] ), .CI(\SUMB[29][29] ), 
        .CO(\CARRYB[30][28] ), .S(\SUMB[30][28] ) );
  FA_X1 S2_30_29 ( .A(\ab[30][29] ), .B(\CARRYB[29][29] ), .CI(\SUMB[29][30] ), 
        .CO(\CARRYB[30][29] ), .S(\SUMB[30][29] ) );
  FA_X1 S2_30_30 ( .A(\ab[30][30] ), .B(\CARRYB[29][30] ), .CI(\SUMB[29][31] ), 
        .CO(\CARRYB[30][30] ), .S(\SUMB[30][30] ) );
  FA_X1 S2_30_31 ( .A(\ab[30][31] ), .B(\CARRYB[29][31] ), .CI(\SUMB[29][32] ), 
        .CO(\CARRYB[30][31] ), .S(\SUMB[30][31] ) );
  FA_X1 S2_30_32 ( .A(\ab[30][32] ), .B(\CARRYB[29][32] ), .CI(\SUMB[29][33] ), 
        .CO(\CARRYB[30][32] ), .S(\SUMB[30][32] ) );
  FA_X1 S2_30_33 ( .A(\ab[30][33] ), .B(\CARRYB[29][33] ), .CI(\SUMB[29][34] ), 
        .CO(\CARRYB[30][33] ), .S(\SUMB[30][33] ) );
  FA_X1 S2_30_34 ( .A(\ab[30][34] ), .B(\CARRYB[29][34] ), .CI(\SUMB[29][35] ), 
        .CO(\CARRYB[30][34] ), .S(\SUMB[30][34] ) );
  FA_X1 S2_30_35 ( .A(\ab[30][35] ), .B(\CARRYB[29][35] ), .CI(\SUMB[29][36] ), 
        .CO(\CARRYB[30][35] ), .S(\SUMB[30][35] ) );
  FA_X1 S2_30_36 ( .A(\ab[30][36] ), .B(\CARRYB[29][36] ), .CI(\SUMB[29][37] ), 
        .CO(\CARRYB[30][36] ), .S(\SUMB[30][36] ) );
  FA_X1 S2_30_37 ( .A(\ab[30][37] ), .B(\CARRYB[29][37] ), .CI(\SUMB[29][38] ), 
        .CO(\CARRYB[30][37] ), .S(\SUMB[30][37] ) );
  FA_X1 S2_30_38 ( .A(\ab[30][38] ), .B(\CARRYB[29][38] ), .CI(\SUMB[29][39] ), 
        .CO(\CARRYB[30][38] ), .S(\SUMB[30][38] ) );
  FA_X1 S2_30_39 ( .A(\ab[30][39] ), .B(\CARRYB[29][39] ), .CI(\SUMB[29][40] ), 
        .CO(\CARRYB[30][39] ), .S(\SUMB[30][39] ) );
  FA_X1 S2_30_40 ( .A(\ab[30][40] ), .B(\CARRYB[29][40] ), .CI(\SUMB[29][41] ), 
        .CO(\CARRYB[30][40] ), .S(\SUMB[30][40] ) );
  FA_X1 S2_30_41 ( .A(\ab[30][41] ), .B(\CARRYB[29][41] ), .CI(\SUMB[29][42] ), 
        .CO(\CARRYB[30][41] ), .S(\SUMB[30][41] ) );
  FA_X1 S2_30_42 ( .A(\ab[30][42] ), .B(\CARRYB[29][42] ), .CI(\SUMB[29][43] ), 
        .CO(\CARRYB[30][42] ), .S(\SUMB[30][42] ) );
  FA_X1 S2_30_43 ( .A(\ab[30][43] ), .B(\CARRYB[29][43] ), .CI(\SUMB[29][44] ), 
        .CO(\CARRYB[30][43] ), .S(\SUMB[30][43] ) );
  FA_X1 S2_30_44 ( .A(\ab[30][44] ), .B(\CARRYB[29][44] ), .CI(\SUMB[29][45] ), 
        .CO(\CARRYB[30][44] ), .S(\SUMB[30][44] ) );
  FA_X1 S2_30_45 ( .A(\ab[30][45] ), .B(\CARRYB[29][45] ), .CI(\SUMB[29][46] ), 
        .CO(\CARRYB[30][45] ), .S(\SUMB[30][45] ) );
  FA_X1 S2_30_46 ( .A(\ab[30][46] ), .B(\CARRYB[29][46] ), .CI(\SUMB[29][47] ), 
        .CO(\CARRYB[30][46] ), .S(\SUMB[30][46] ) );
  FA_X1 S2_30_47 ( .A(\ab[30][47] ), .B(\CARRYB[29][47] ), .CI(\SUMB[29][48] ), 
        .CO(\CARRYB[30][47] ), .S(\SUMB[30][47] ) );
  FA_X1 S2_30_48 ( .A(\ab[30][48] ), .B(\CARRYB[29][48] ), .CI(\SUMB[29][49] ), 
        .CO(\CARRYB[30][48] ), .S(\SUMB[30][48] ) );
  FA_X1 S2_30_49 ( .A(\ab[30][49] ), .B(\CARRYB[29][49] ), .CI(\SUMB[29][50] ), 
        .CO(\CARRYB[30][49] ), .S(\SUMB[30][49] ) );
  FA_X1 S2_30_50 ( .A(\ab[30][50] ), .B(\CARRYB[29][50] ), .CI(\SUMB[29][51] ), 
        .CO(\CARRYB[30][50] ), .S(\SUMB[30][50] ) );
  FA_X1 S3_30_51 ( .A(\ab[30][51] ), .B(\CARRYB[29][51] ), .CI(\ab[29][52] ), 
        .CO(\CARRYB[30][51] ), .S(\SUMB[30][51] ) );
  FA_X1 S1_29_0 ( .A(\ab[29][0] ), .B(\CARRYB[28][0] ), .CI(\SUMB[28][1] ), 
        .CO(\CARRYB[29][0] ), .S(CLA_SUM[29]) );
  FA_X1 S2_29_1 ( .A(\ab[29][1] ), .B(\CARRYB[28][1] ), .CI(\SUMB[28][2] ), 
        .CO(\CARRYB[29][1] ), .S(\SUMB[29][1] ) );
  FA_X1 S2_29_2 ( .A(\ab[29][2] ), .B(\CARRYB[28][2] ), .CI(\SUMB[28][3] ), 
        .CO(\CARRYB[29][2] ), .S(\SUMB[29][2] ) );
  FA_X1 S2_29_3 ( .A(\ab[29][3] ), .B(\CARRYB[28][3] ), .CI(\SUMB[28][4] ), 
        .CO(\CARRYB[29][3] ), .S(\SUMB[29][3] ) );
  FA_X1 S2_29_4 ( .A(\ab[29][4] ), .B(\CARRYB[28][4] ), .CI(\SUMB[28][5] ), 
        .CO(\CARRYB[29][4] ), .S(\SUMB[29][4] ) );
  FA_X1 S2_29_5 ( .A(\ab[29][5] ), .B(\CARRYB[28][5] ), .CI(\SUMB[28][6] ), 
        .CO(\CARRYB[29][5] ), .S(\SUMB[29][5] ) );
  FA_X1 S2_29_6 ( .A(\ab[29][6] ), .B(\CARRYB[28][6] ), .CI(\SUMB[28][7] ), 
        .CO(\CARRYB[29][6] ), .S(\SUMB[29][6] ) );
  FA_X1 S2_29_7 ( .A(\ab[29][7] ), .B(\CARRYB[28][7] ), .CI(\SUMB[28][8] ), 
        .CO(\CARRYB[29][7] ), .S(\SUMB[29][7] ) );
  FA_X1 S2_29_8 ( .A(\ab[29][8] ), .B(\CARRYB[28][8] ), .CI(\SUMB[28][9] ), 
        .CO(\CARRYB[29][8] ), .S(\SUMB[29][8] ) );
  FA_X1 S2_29_9 ( .A(\ab[29][9] ), .B(\CARRYB[28][9] ), .CI(\SUMB[28][10] ), 
        .CO(\CARRYB[29][9] ), .S(\SUMB[29][9] ) );
  FA_X1 S2_29_10 ( .A(\ab[29][10] ), .B(\CARRYB[28][10] ), .CI(\SUMB[28][11] ), 
        .CO(\CARRYB[29][10] ), .S(\SUMB[29][10] ) );
  FA_X1 S2_29_11 ( .A(\ab[29][11] ), .B(\CARRYB[28][11] ), .CI(\SUMB[28][12] ), 
        .CO(\CARRYB[29][11] ), .S(\SUMB[29][11] ) );
  FA_X1 S2_29_12 ( .A(\ab[29][12] ), .B(\CARRYB[28][12] ), .CI(\SUMB[28][13] ), 
        .CO(\CARRYB[29][12] ), .S(\SUMB[29][12] ) );
  FA_X1 S2_29_13 ( .A(\ab[29][13] ), .B(\CARRYB[28][13] ), .CI(\SUMB[28][14] ), 
        .CO(\CARRYB[29][13] ), .S(\SUMB[29][13] ) );
  FA_X1 S2_29_14 ( .A(\ab[29][14] ), .B(\CARRYB[28][14] ), .CI(\SUMB[28][15] ), 
        .CO(\CARRYB[29][14] ), .S(\SUMB[29][14] ) );
  FA_X1 S2_29_15 ( .A(\ab[29][15] ), .B(\CARRYB[28][15] ), .CI(\SUMB[28][16] ), 
        .CO(\CARRYB[29][15] ), .S(\SUMB[29][15] ) );
  FA_X1 S2_29_16 ( .A(\ab[29][16] ), .B(\CARRYB[28][16] ), .CI(\SUMB[28][17] ), 
        .CO(\CARRYB[29][16] ), .S(\SUMB[29][16] ) );
  FA_X1 S2_29_17 ( .A(\ab[29][17] ), .B(\CARRYB[28][17] ), .CI(\SUMB[28][18] ), 
        .CO(\CARRYB[29][17] ), .S(\SUMB[29][17] ) );
  FA_X1 S2_29_18 ( .A(\ab[29][18] ), .B(\CARRYB[28][18] ), .CI(\SUMB[28][19] ), 
        .CO(\CARRYB[29][18] ), .S(\SUMB[29][18] ) );
  FA_X1 S2_29_19 ( .A(\ab[29][19] ), .B(\CARRYB[28][19] ), .CI(\SUMB[28][20] ), 
        .CO(\CARRYB[29][19] ), .S(\SUMB[29][19] ) );
  FA_X1 S2_29_20 ( .A(\ab[29][20] ), .B(\CARRYB[28][20] ), .CI(\SUMB[28][21] ), 
        .CO(\CARRYB[29][20] ), .S(\SUMB[29][20] ) );
  FA_X1 S2_29_21 ( .A(\ab[29][21] ), .B(\CARRYB[28][21] ), .CI(\SUMB[28][22] ), 
        .CO(\CARRYB[29][21] ), .S(\SUMB[29][21] ) );
  FA_X1 S2_29_22 ( .A(\ab[29][22] ), .B(\CARRYB[28][22] ), .CI(\SUMB[28][23] ), 
        .CO(\CARRYB[29][22] ), .S(\SUMB[29][22] ) );
  FA_X1 S2_29_23 ( .A(\ab[29][23] ), .B(\CARRYB[28][23] ), .CI(\SUMB[28][24] ), 
        .CO(\CARRYB[29][23] ), .S(\SUMB[29][23] ) );
  FA_X1 S2_29_24 ( .A(\ab[29][24] ), .B(\CARRYB[28][24] ), .CI(\SUMB[28][25] ), 
        .CO(\CARRYB[29][24] ), .S(\SUMB[29][24] ) );
  FA_X1 S2_29_25 ( .A(\ab[29][25] ), .B(\CARRYB[28][25] ), .CI(\SUMB[28][26] ), 
        .CO(\CARRYB[29][25] ), .S(\SUMB[29][25] ) );
  FA_X1 S2_29_26 ( .A(\ab[29][26] ), .B(\CARRYB[28][26] ), .CI(\SUMB[28][27] ), 
        .CO(\CARRYB[29][26] ), .S(\SUMB[29][26] ) );
  FA_X1 S2_29_27 ( .A(\ab[29][27] ), .B(\CARRYB[28][27] ), .CI(\SUMB[28][28] ), 
        .CO(\CARRYB[29][27] ), .S(\SUMB[29][27] ) );
  FA_X1 S2_29_28 ( .A(\ab[29][28] ), .B(\CARRYB[28][28] ), .CI(\SUMB[28][29] ), 
        .CO(\CARRYB[29][28] ), .S(\SUMB[29][28] ) );
  FA_X1 S2_29_29 ( .A(\ab[29][29] ), .B(\CARRYB[28][29] ), .CI(\SUMB[28][30] ), 
        .CO(\CARRYB[29][29] ), .S(\SUMB[29][29] ) );
  FA_X1 S2_29_30 ( .A(\ab[29][30] ), .B(\CARRYB[28][30] ), .CI(\SUMB[28][31] ), 
        .CO(\CARRYB[29][30] ), .S(\SUMB[29][30] ) );
  FA_X1 S2_29_31 ( .A(\ab[29][31] ), .B(\CARRYB[28][31] ), .CI(\SUMB[28][32] ), 
        .CO(\CARRYB[29][31] ), .S(\SUMB[29][31] ) );
  FA_X1 S2_29_32 ( .A(\ab[29][32] ), .B(\CARRYB[28][32] ), .CI(\SUMB[28][33] ), 
        .CO(\CARRYB[29][32] ), .S(\SUMB[29][32] ) );
  FA_X1 S2_29_33 ( .A(\ab[29][33] ), .B(\CARRYB[28][33] ), .CI(\SUMB[28][34] ), 
        .CO(\CARRYB[29][33] ), .S(\SUMB[29][33] ) );
  FA_X1 S2_29_34 ( .A(\ab[29][34] ), .B(\CARRYB[28][34] ), .CI(\SUMB[28][35] ), 
        .CO(\CARRYB[29][34] ), .S(\SUMB[29][34] ) );
  FA_X1 S2_29_35 ( .A(\ab[29][35] ), .B(\CARRYB[28][35] ), .CI(\SUMB[28][36] ), 
        .CO(\CARRYB[29][35] ), .S(\SUMB[29][35] ) );
  FA_X1 S2_29_36 ( .A(\ab[29][36] ), .B(\CARRYB[28][36] ), .CI(\SUMB[28][37] ), 
        .CO(\CARRYB[29][36] ), .S(\SUMB[29][36] ) );
  FA_X1 S2_29_37 ( .A(\ab[29][37] ), .B(\CARRYB[28][37] ), .CI(\SUMB[28][38] ), 
        .CO(\CARRYB[29][37] ), .S(\SUMB[29][37] ) );
  FA_X1 S2_29_38 ( .A(\ab[29][38] ), .B(\CARRYB[28][38] ), .CI(\SUMB[28][39] ), 
        .CO(\CARRYB[29][38] ), .S(\SUMB[29][38] ) );
  FA_X1 S2_29_39 ( .A(\ab[29][39] ), .B(\CARRYB[28][39] ), .CI(\SUMB[28][40] ), 
        .CO(\CARRYB[29][39] ), .S(\SUMB[29][39] ) );
  FA_X1 S2_29_40 ( .A(\ab[29][40] ), .B(\CARRYB[28][40] ), .CI(\SUMB[28][41] ), 
        .CO(\CARRYB[29][40] ), .S(\SUMB[29][40] ) );
  FA_X1 S2_29_41 ( .A(\ab[29][41] ), .B(\CARRYB[28][41] ), .CI(\SUMB[28][42] ), 
        .CO(\CARRYB[29][41] ), .S(\SUMB[29][41] ) );
  FA_X1 S2_29_42 ( .A(\ab[29][42] ), .B(\CARRYB[28][42] ), .CI(\SUMB[28][43] ), 
        .CO(\CARRYB[29][42] ), .S(\SUMB[29][42] ) );
  FA_X1 S2_29_43 ( .A(\ab[29][43] ), .B(\CARRYB[28][43] ), .CI(\SUMB[28][44] ), 
        .CO(\CARRYB[29][43] ), .S(\SUMB[29][43] ) );
  FA_X1 S2_29_44 ( .A(\ab[29][44] ), .B(\CARRYB[28][44] ), .CI(\SUMB[28][45] ), 
        .CO(\CARRYB[29][44] ), .S(\SUMB[29][44] ) );
  FA_X1 S2_29_45 ( .A(\ab[29][45] ), .B(\CARRYB[28][45] ), .CI(\SUMB[28][46] ), 
        .CO(\CARRYB[29][45] ), .S(\SUMB[29][45] ) );
  FA_X1 S2_29_46 ( .A(\ab[29][46] ), .B(\CARRYB[28][46] ), .CI(\SUMB[28][47] ), 
        .CO(\CARRYB[29][46] ), .S(\SUMB[29][46] ) );
  FA_X1 S2_29_47 ( .A(\ab[29][47] ), .B(\CARRYB[28][47] ), .CI(\SUMB[28][48] ), 
        .CO(\CARRYB[29][47] ), .S(\SUMB[29][47] ) );
  FA_X1 S2_29_48 ( .A(\ab[29][48] ), .B(\CARRYB[28][48] ), .CI(\SUMB[28][49] ), 
        .CO(\CARRYB[29][48] ), .S(\SUMB[29][48] ) );
  FA_X1 S2_29_49 ( .A(\ab[29][49] ), .B(\CARRYB[28][49] ), .CI(\SUMB[28][50] ), 
        .CO(\CARRYB[29][49] ), .S(\SUMB[29][49] ) );
  FA_X1 S2_29_50 ( .A(\ab[29][50] ), .B(\CARRYB[28][50] ), .CI(\SUMB[28][51] ), 
        .CO(\CARRYB[29][50] ), .S(\SUMB[29][50] ) );
  FA_X1 S3_29_51 ( .A(\ab[29][51] ), .B(\CARRYB[28][51] ), .CI(\ab[28][52] ), 
        .CO(\CARRYB[29][51] ), .S(\SUMB[29][51] ) );
  FA_X1 S1_28_0 ( .A(\ab[28][0] ), .B(\CARRYB[27][0] ), .CI(\SUMB[27][1] ), 
        .CO(\CARRYB[28][0] ), .S(CLA_SUM[28]) );
  FA_X1 S2_28_1 ( .A(\ab[28][1] ), .B(\CARRYB[27][1] ), .CI(\SUMB[27][2] ), 
        .CO(\CARRYB[28][1] ), .S(\SUMB[28][1] ) );
  FA_X1 S2_28_2 ( .A(\ab[28][2] ), .B(\CARRYB[27][2] ), .CI(\SUMB[27][3] ), 
        .CO(\CARRYB[28][2] ), .S(\SUMB[28][2] ) );
  FA_X1 S2_28_3 ( .A(\ab[28][3] ), .B(\CARRYB[27][3] ), .CI(\SUMB[27][4] ), 
        .CO(\CARRYB[28][3] ), .S(\SUMB[28][3] ) );
  FA_X1 S2_28_4 ( .A(\ab[28][4] ), .B(\CARRYB[27][4] ), .CI(\SUMB[27][5] ), 
        .CO(\CARRYB[28][4] ), .S(\SUMB[28][4] ) );
  FA_X1 S2_28_5 ( .A(\ab[28][5] ), .B(\CARRYB[27][5] ), .CI(\SUMB[27][6] ), 
        .CO(\CARRYB[28][5] ), .S(\SUMB[28][5] ) );
  FA_X1 S2_28_6 ( .A(\ab[28][6] ), .B(\CARRYB[27][6] ), .CI(\SUMB[27][7] ), 
        .CO(\CARRYB[28][6] ), .S(\SUMB[28][6] ) );
  FA_X1 S2_28_7 ( .A(\ab[28][7] ), .B(\CARRYB[27][7] ), .CI(\SUMB[27][8] ), 
        .CO(\CARRYB[28][7] ), .S(\SUMB[28][7] ) );
  FA_X1 S2_28_8 ( .A(\ab[28][8] ), .B(\CARRYB[27][8] ), .CI(\SUMB[27][9] ), 
        .CO(\CARRYB[28][8] ), .S(\SUMB[28][8] ) );
  FA_X1 S2_28_9 ( .A(\ab[28][9] ), .B(\CARRYB[27][9] ), .CI(\SUMB[27][10] ), 
        .CO(\CARRYB[28][9] ), .S(\SUMB[28][9] ) );
  FA_X1 S2_28_10 ( .A(\ab[28][10] ), .B(\CARRYB[27][10] ), .CI(\SUMB[27][11] ), 
        .CO(\CARRYB[28][10] ), .S(\SUMB[28][10] ) );
  FA_X1 S2_28_11 ( .A(\ab[28][11] ), .B(\CARRYB[27][11] ), .CI(\SUMB[27][12] ), 
        .CO(\CARRYB[28][11] ), .S(\SUMB[28][11] ) );
  FA_X1 S2_28_12 ( .A(\ab[28][12] ), .B(\CARRYB[27][12] ), .CI(\SUMB[27][13] ), 
        .CO(\CARRYB[28][12] ), .S(\SUMB[28][12] ) );
  FA_X1 S2_28_13 ( .A(\ab[28][13] ), .B(\CARRYB[27][13] ), .CI(\SUMB[27][14] ), 
        .CO(\CARRYB[28][13] ), .S(\SUMB[28][13] ) );
  FA_X1 S2_28_14 ( .A(\ab[28][14] ), .B(\CARRYB[27][14] ), .CI(\SUMB[27][15] ), 
        .CO(\CARRYB[28][14] ), .S(\SUMB[28][14] ) );
  FA_X1 S2_28_15 ( .A(\ab[28][15] ), .B(\CARRYB[27][15] ), .CI(\SUMB[27][16] ), 
        .CO(\CARRYB[28][15] ), .S(\SUMB[28][15] ) );
  FA_X1 S2_28_16 ( .A(\ab[28][16] ), .B(\CARRYB[27][16] ), .CI(\SUMB[27][17] ), 
        .CO(\CARRYB[28][16] ), .S(\SUMB[28][16] ) );
  FA_X1 S2_28_17 ( .A(\ab[28][17] ), .B(\CARRYB[27][17] ), .CI(\SUMB[27][18] ), 
        .CO(\CARRYB[28][17] ), .S(\SUMB[28][17] ) );
  FA_X1 S2_28_18 ( .A(\ab[28][18] ), .B(\CARRYB[27][18] ), .CI(\SUMB[27][19] ), 
        .CO(\CARRYB[28][18] ), .S(\SUMB[28][18] ) );
  FA_X1 S2_28_19 ( .A(\ab[28][19] ), .B(\CARRYB[27][19] ), .CI(\SUMB[27][20] ), 
        .CO(\CARRYB[28][19] ), .S(\SUMB[28][19] ) );
  FA_X1 S2_28_20 ( .A(\ab[28][20] ), .B(\CARRYB[27][20] ), .CI(\SUMB[27][21] ), 
        .CO(\CARRYB[28][20] ), .S(\SUMB[28][20] ) );
  FA_X1 S2_28_21 ( .A(\ab[28][21] ), .B(\CARRYB[27][21] ), .CI(\SUMB[27][22] ), 
        .CO(\CARRYB[28][21] ), .S(\SUMB[28][21] ) );
  FA_X1 S2_28_22 ( .A(\ab[28][22] ), .B(\CARRYB[27][22] ), .CI(\SUMB[27][23] ), 
        .CO(\CARRYB[28][22] ), .S(\SUMB[28][22] ) );
  FA_X1 S2_28_23 ( .A(\ab[28][23] ), .B(\CARRYB[27][23] ), .CI(\SUMB[27][24] ), 
        .CO(\CARRYB[28][23] ), .S(\SUMB[28][23] ) );
  FA_X1 S2_28_24 ( .A(\ab[28][24] ), .B(\CARRYB[27][24] ), .CI(\SUMB[27][25] ), 
        .CO(\CARRYB[28][24] ), .S(\SUMB[28][24] ) );
  FA_X1 S2_28_25 ( .A(\ab[28][25] ), .B(\CARRYB[27][25] ), .CI(\SUMB[27][26] ), 
        .CO(\CARRYB[28][25] ), .S(\SUMB[28][25] ) );
  FA_X1 S2_28_26 ( .A(\ab[28][26] ), .B(\CARRYB[27][26] ), .CI(\SUMB[27][27] ), 
        .CO(\CARRYB[28][26] ), .S(\SUMB[28][26] ) );
  FA_X1 S2_28_27 ( .A(\ab[28][27] ), .B(\CARRYB[27][27] ), .CI(\SUMB[27][28] ), 
        .CO(\CARRYB[28][27] ), .S(\SUMB[28][27] ) );
  FA_X1 S2_28_28 ( .A(\ab[28][28] ), .B(\CARRYB[27][28] ), .CI(\SUMB[27][29] ), 
        .CO(\CARRYB[28][28] ), .S(\SUMB[28][28] ) );
  FA_X1 S2_28_29 ( .A(\ab[28][29] ), .B(\CARRYB[27][29] ), .CI(\SUMB[27][30] ), 
        .CO(\CARRYB[28][29] ), .S(\SUMB[28][29] ) );
  FA_X1 S2_28_30 ( .A(\ab[28][30] ), .B(\CARRYB[27][30] ), .CI(\SUMB[27][31] ), 
        .CO(\CARRYB[28][30] ), .S(\SUMB[28][30] ) );
  FA_X1 S2_28_31 ( .A(\ab[28][31] ), .B(\CARRYB[27][31] ), .CI(\SUMB[27][32] ), 
        .CO(\CARRYB[28][31] ), .S(\SUMB[28][31] ) );
  FA_X1 S2_28_32 ( .A(\ab[28][32] ), .B(\CARRYB[27][32] ), .CI(\SUMB[27][33] ), 
        .CO(\CARRYB[28][32] ), .S(\SUMB[28][32] ) );
  FA_X1 S2_28_33 ( .A(\ab[28][33] ), .B(\CARRYB[27][33] ), .CI(\SUMB[27][34] ), 
        .CO(\CARRYB[28][33] ), .S(\SUMB[28][33] ) );
  FA_X1 S2_28_34 ( .A(\ab[28][34] ), .B(\CARRYB[27][34] ), .CI(\SUMB[27][35] ), 
        .CO(\CARRYB[28][34] ), .S(\SUMB[28][34] ) );
  FA_X1 S2_28_35 ( .A(\ab[28][35] ), .B(\CARRYB[27][35] ), .CI(\SUMB[27][36] ), 
        .CO(\CARRYB[28][35] ), .S(\SUMB[28][35] ) );
  FA_X1 S2_28_36 ( .A(\ab[28][36] ), .B(\CARRYB[27][36] ), .CI(\SUMB[27][37] ), 
        .CO(\CARRYB[28][36] ), .S(\SUMB[28][36] ) );
  FA_X1 S2_28_37 ( .A(\ab[28][37] ), .B(\CARRYB[27][37] ), .CI(\SUMB[27][38] ), 
        .CO(\CARRYB[28][37] ), .S(\SUMB[28][37] ) );
  FA_X1 S2_28_38 ( .A(\ab[28][38] ), .B(\CARRYB[27][38] ), .CI(\SUMB[27][39] ), 
        .CO(\CARRYB[28][38] ), .S(\SUMB[28][38] ) );
  FA_X1 S2_28_39 ( .A(\ab[28][39] ), .B(\CARRYB[27][39] ), .CI(\SUMB[27][40] ), 
        .CO(\CARRYB[28][39] ), .S(\SUMB[28][39] ) );
  FA_X1 S2_28_40 ( .A(\ab[28][40] ), .B(\CARRYB[27][40] ), .CI(\SUMB[27][41] ), 
        .CO(\CARRYB[28][40] ), .S(\SUMB[28][40] ) );
  FA_X1 S2_28_41 ( .A(\ab[28][41] ), .B(\CARRYB[27][41] ), .CI(\SUMB[27][42] ), 
        .CO(\CARRYB[28][41] ), .S(\SUMB[28][41] ) );
  FA_X1 S2_28_42 ( .A(\ab[28][42] ), .B(\CARRYB[27][42] ), .CI(\SUMB[27][43] ), 
        .CO(\CARRYB[28][42] ), .S(\SUMB[28][42] ) );
  FA_X1 S2_28_43 ( .A(\ab[28][43] ), .B(\CARRYB[27][43] ), .CI(\SUMB[27][44] ), 
        .CO(\CARRYB[28][43] ), .S(\SUMB[28][43] ) );
  FA_X1 S2_28_44 ( .A(\ab[28][44] ), .B(\CARRYB[27][44] ), .CI(\SUMB[27][45] ), 
        .CO(\CARRYB[28][44] ), .S(\SUMB[28][44] ) );
  FA_X1 S2_28_45 ( .A(\ab[28][45] ), .B(\CARRYB[27][45] ), .CI(\SUMB[27][46] ), 
        .CO(\CARRYB[28][45] ), .S(\SUMB[28][45] ) );
  FA_X1 S2_28_46 ( .A(\ab[28][46] ), .B(\CARRYB[27][46] ), .CI(\SUMB[27][47] ), 
        .CO(\CARRYB[28][46] ), .S(\SUMB[28][46] ) );
  FA_X1 S2_28_47 ( .A(\ab[28][47] ), .B(\CARRYB[27][47] ), .CI(\SUMB[27][48] ), 
        .CO(\CARRYB[28][47] ), .S(\SUMB[28][47] ) );
  FA_X1 S2_28_48 ( .A(\ab[28][48] ), .B(\CARRYB[27][48] ), .CI(\SUMB[27][49] ), 
        .CO(\CARRYB[28][48] ), .S(\SUMB[28][48] ) );
  FA_X1 S2_28_49 ( .A(\ab[28][49] ), .B(\CARRYB[27][49] ), .CI(\SUMB[27][50] ), 
        .CO(\CARRYB[28][49] ), .S(\SUMB[28][49] ) );
  FA_X1 S2_28_50 ( .A(\ab[28][50] ), .B(\CARRYB[27][50] ), .CI(\SUMB[27][51] ), 
        .CO(\CARRYB[28][50] ), .S(\SUMB[28][50] ) );
  FA_X1 S3_28_51 ( .A(\ab[28][51] ), .B(\CARRYB[27][51] ), .CI(\ab[27][52] ), 
        .CO(\CARRYB[28][51] ), .S(\SUMB[28][51] ) );
  FA_X1 S1_27_0 ( .A(\ab[27][0] ), .B(\CARRYB[26][0] ), .CI(\SUMB[26][1] ), 
        .CO(\CARRYB[27][0] ), .S(CLA_SUM[27]) );
  FA_X1 S2_27_1 ( .A(\ab[27][1] ), .B(\CARRYB[26][1] ), .CI(\SUMB[26][2] ), 
        .CO(\CARRYB[27][1] ), .S(\SUMB[27][1] ) );
  FA_X1 S2_27_2 ( .A(\ab[27][2] ), .B(\CARRYB[26][2] ), .CI(\SUMB[26][3] ), 
        .CO(\CARRYB[27][2] ), .S(\SUMB[27][2] ) );
  FA_X1 S2_27_3 ( .A(\ab[27][3] ), .B(\CARRYB[26][3] ), .CI(\SUMB[26][4] ), 
        .CO(\CARRYB[27][3] ), .S(\SUMB[27][3] ) );
  FA_X1 S2_27_4 ( .A(\ab[27][4] ), .B(\CARRYB[26][4] ), .CI(\SUMB[26][5] ), 
        .CO(\CARRYB[27][4] ), .S(\SUMB[27][4] ) );
  FA_X1 S2_27_5 ( .A(\ab[27][5] ), .B(\CARRYB[26][5] ), .CI(\SUMB[26][6] ), 
        .CO(\CARRYB[27][5] ), .S(\SUMB[27][5] ) );
  FA_X1 S2_27_6 ( .A(\ab[27][6] ), .B(\CARRYB[26][6] ), .CI(\SUMB[26][7] ), 
        .CO(\CARRYB[27][6] ), .S(\SUMB[27][6] ) );
  FA_X1 S2_27_7 ( .A(\ab[27][7] ), .B(\CARRYB[26][7] ), .CI(\SUMB[26][8] ), 
        .CO(\CARRYB[27][7] ), .S(\SUMB[27][7] ) );
  FA_X1 S2_27_8 ( .A(\ab[27][8] ), .B(\CARRYB[26][8] ), .CI(\SUMB[26][9] ), 
        .CO(\CARRYB[27][8] ), .S(\SUMB[27][8] ) );
  FA_X1 S2_27_9 ( .A(\ab[27][9] ), .B(\CARRYB[26][9] ), .CI(\SUMB[26][10] ), 
        .CO(\CARRYB[27][9] ), .S(\SUMB[27][9] ) );
  FA_X1 S2_27_10 ( .A(\ab[27][10] ), .B(\CARRYB[26][10] ), .CI(\SUMB[26][11] ), 
        .CO(\CARRYB[27][10] ), .S(\SUMB[27][10] ) );
  FA_X1 S2_27_11 ( .A(\ab[27][11] ), .B(\CARRYB[26][11] ), .CI(\SUMB[26][12] ), 
        .CO(\CARRYB[27][11] ), .S(\SUMB[27][11] ) );
  FA_X1 S2_27_12 ( .A(\ab[27][12] ), .B(\CARRYB[26][12] ), .CI(\SUMB[26][13] ), 
        .CO(\CARRYB[27][12] ), .S(\SUMB[27][12] ) );
  FA_X1 S2_27_13 ( .A(\ab[27][13] ), .B(\CARRYB[26][13] ), .CI(\SUMB[26][14] ), 
        .CO(\CARRYB[27][13] ), .S(\SUMB[27][13] ) );
  FA_X1 S2_27_14 ( .A(\ab[27][14] ), .B(\CARRYB[26][14] ), .CI(\SUMB[26][15] ), 
        .CO(\CARRYB[27][14] ), .S(\SUMB[27][14] ) );
  FA_X1 S2_27_15 ( .A(\ab[27][15] ), .B(\CARRYB[26][15] ), .CI(\SUMB[26][16] ), 
        .CO(\CARRYB[27][15] ), .S(\SUMB[27][15] ) );
  FA_X1 S2_27_16 ( .A(\ab[27][16] ), .B(\CARRYB[26][16] ), .CI(\SUMB[26][17] ), 
        .CO(\CARRYB[27][16] ), .S(\SUMB[27][16] ) );
  FA_X1 S2_27_17 ( .A(\ab[27][17] ), .B(\CARRYB[26][17] ), .CI(\SUMB[26][18] ), 
        .CO(\CARRYB[27][17] ), .S(\SUMB[27][17] ) );
  FA_X1 S2_27_18 ( .A(\ab[27][18] ), .B(\CARRYB[26][18] ), .CI(\SUMB[26][19] ), 
        .CO(\CARRYB[27][18] ), .S(\SUMB[27][18] ) );
  FA_X1 S2_27_19 ( .A(\ab[27][19] ), .B(\CARRYB[26][19] ), .CI(\SUMB[26][20] ), 
        .CO(\CARRYB[27][19] ), .S(\SUMB[27][19] ) );
  FA_X1 S2_27_20 ( .A(\ab[27][20] ), .B(\CARRYB[26][20] ), .CI(\SUMB[26][21] ), 
        .CO(\CARRYB[27][20] ), .S(\SUMB[27][20] ) );
  FA_X1 S2_27_21 ( .A(\ab[27][21] ), .B(\CARRYB[26][21] ), .CI(\SUMB[26][22] ), 
        .CO(\CARRYB[27][21] ), .S(\SUMB[27][21] ) );
  FA_X1 S2_27_22 ( .A(\ab[27][22] ), .B(\CARRYB[26][22] ), .CI(\SUMB[26][23] ), 
        .CO(\CARRYB[27][22] ), .S(\SUMB[27][22] ) );
  FA_X1 S2_27_23 ( .A(\ab[27][23] ), .B(\CARRYB[26][23] ), .CI(\SUMB[26][24] ), 
        .CO(\CARRYB[27][23] ), .S(\SUMB[27][23] ) );
  FA_X1 S2_27_24 ( .A(\ab[27][24] ), .B(\CARRYB[26][24] ), .CI(\SUMB[26][25] ), 
        .CO(\CARRYB[27][24] ), .S(\SUMB[27][24] ) );
  FA_X1 S2_27_25 ( .A(\ab[27][25] ), .B(\CARRYB[26][25] ), .CI(\SUMB[26][26] ), 
        .CO(\CARRYB[27][25] ), .S(\SUMB[27][25] ) );
  FA_X1 S2_27_26 ( .A(\ab[27][26] ), .B(\CARRYB[26][26] ), .CI(\SUMB[26][27] ), 
        .CO(\CARRYB[27][26] ), .S(\SUMB[27][26] ) );
  FA_X1 S2_27_27 ( .A(\ab[27][27] ), .B(\CARRYB[26][27] ), .CI(\SUMB[26][28] ), 
        .CO(\CARRYB[27][27] ), .S(\SUMB[27][27] ) );
  FA_X1 S2_27_28 ( .A(\ab[27][28] ), .B(\CARRYB[26][28] ), .CI(\SUMB[26][29] ), 
        .CO(\CARRYB[27][28] ), .S(\SUMB[27][28] ) );
  FA_X1 S2_27_29 ( .A(\ab[27][29] ), .B(\CARRYB[26][29] ), .CI(\SUMB[26][30] ), 
        .CO(\CARRYB[27][29] ), .S(\SUMB[27][29] ) );
  FA_X1 S2_27_30 ( .A(\ab[27][30] ), .B(\CARRYB[26][30] ), .CI(\SUMB[26][31] ), 
        .CO(\CARRYB[27][30] ), .S(\SUMB[27][30] ) );
  FA_X1 S2_27_31 ( .A(\ab[27][31] ), .B(\CARRYB[26][31] ), .CI(\SUMB[26][32] ), 
        .CO(\CARRYB[27][31] ), .S(\SUMB[27][31] ) );
  FA_X1 S2_27_32 ( .A(\ab[27][32] ), .B(\CARRYB[26][32] ), .CI(\SUMB[26][33] ), 
        .CO(\CARRYB[27][32] ), .S(\SUMB[27][32] ) );
  FA_X1 S2_27_33 ( .A(\ab[27][33] ), .B(\CARRYB[26][33] ), .CI(\SUMB[26][34] ), 
        .CO(\CARRYB[27][33] ), .S(\SUMB[27][33] ) );
  FA_X1 S2_27_34 ( .A(\ab[27][34] ), .B(\CARRYB[26][34] ), .CI(\SUMB[26][35] ), 
        .CO(\CARRYB[27][34] ), .S(\SUMB[27][34] ) );
  FA_X1 S2_27_35 ( .A(\ab[27][35] ), .B(\CARRYB[26][35] ), .CI(\SUMB[26][36] ), 
        .CO(\CARRYB[27][35] ), .S(\SUMB[27][35] ) );
  FA_X1 S2_27_36 ( .A(\ab[27][36] ), .B(\CARRYB[26][36] ), .CI(\SUMB[26][37] ), 
        .CO(\CARRYB[27][36] ), .S(\SUMB[27][36] ) );
  FA_X1 S2_27_37 ( .A(\ab[27][37] ), .B(\CARRYB[26][37] ), .CI(\SUMB[26][38] ), 
        .CO(\CARRYB[27][37] ), .S(\SUMB[27][37] ) );
  FA_X1 S2_27_38 ( .A(\ab[27][38] ), .B(\CARRYB[26][38] ), .CI(\SUMB[26][39] ), 
        .CO(\CARRYB[27][38] ), .S(\SUMB[27][38] ) );
  FA_X1 S2_27_39 ( .A(\ab[27][39] ), .B(\CARRYB[26][39] ), .CI(\SUMB[26][40] ), 
        .CO(\CARRYB[27][39] ), .S(\SUMB[27][39] ) );
  FA_X1 S2_27_40 ( .A(\ab[27][40] ), .B(\CARRYB[26][40] ), .CI(\SUMB[26][41] ), 
        .CO(\CARRYB[27][40] ), .S(\SUMB[27][40] ) );
  FA_X1 S2_27_41 ( .A(\ab[27][41] ), .B(\CARRYB[26][41] ), .CI(\SUMB[26][42] ), 
        .CO(\CARRYB[27][41] ), .S(\SUMB[27][41] ) );
  FA_X1 S2_27_42 ( .A(\ab[27][42] ), .B(\CARRYB[26][42] ), .CI(\SUMB[26][43] ), 
        .CO(\CARRYB[27][42] ), .S(\SUMB[27][42] ) );
  FA_X1 S2_27_43 ( .A(\ab[27][43] ), .B(\CARRYB[26][43] ), .CI(\SUMB[26][44] ), 
        .CO(\CARRYB[27][43] ), .S(\SUMB[27][43] ) );
  FA_X1 S2_27_44 ( .A(\ab[27][44] ), .B(\CARRYB[26][44] ), .CI(\SUMB[26][45] ), 
        .CO(\CARRYB[27][44] ), .S(\SUMB[27][44] ) );
  FA_X1 S2_27_45 ( .A(\ab[27][45] ), .B(\CARRYB[26][45] ), .CI(\SUMB[26][46] ), 
        .CO(\CARRYB[27][45] ), .S(\SUMB[27][45] ) );
  FA_X1 S2_27_46 ( .A(\ab[27][46] ), .B(\CARRYB[26][46] ), .CI(\SUMB[26][47] ), 
        .CO(\CARRYB[27][46] ), .S(\SUMB[27][46] ) );
  FA_X1 S2_27_47 ( .A(\ab[27][47] ), .B(\CARRYB[26][47] ), .CI(\SUMB[26][48] ), 
        .CO(\CARRYB[27][47] ), .S(\SUMB[27][47] ) );
  FA_X1 S2_27_48 ( .A(\ab[27][48] ), .B(\CARRYB[26][48] ), .CI(\SUMB[26][49] ), 
        .CO(\CARRYB[27][48] ), .S(\SUMB[27][48] ) );
  FA_X1 S2_27_49 ( .A(\ab[27][49] ), .B(\CARRYB[26][49] ), .CI(\SUMB[26][50] ), 
        .CO(\CARRYB[27][49] ), .S(\SUMB[27][49] ) );
  FA_X1 S2_27_50 ( .A(\ab[27][50] ), .B(\CARRYB[26][50] ), .CI(\SUMB[26][51] ), 
        .CO(\CARRYB[27][50] ), .S(\SUMB[27][50] ) );
  FA_X1 S3_27_51 ( .A(\ab[27][51] ), .B(\CARRYB[26][51] ), .CI(\ab[26][52] ), 
        .CO(\CARRYB[27][51] ), .S(\SUMB[27][51] ) );
  FA_X1 S1_26_0 ( .A(\ab[26][0] ), .B(\CARRYB[25][0] ), .CI(\SUMB[25][1] ), 
        .CO(\CARRYB[26][0] ), .S(CLA_SUM[26]) );
  FA_X1 S2_26_1 ( .A(\ab[26][1] ), .B(\CARRYB[25][1] ), .CI(\SUMB[25][2] ), 
        .CO(\CARRYB[26][1] ), .S(\SUMB[26][1] ) );
  FA_X1 S2_26_2 ( .A(\ab[26][2] ), .B(\CARRYB[25][2] ), .CI(\SUMB[25][3] ), 
        .CO(\CARRYB[26][2] ), .S(\SUMB[26][2] ) );
  FA_X1 S2_26_3 ( .A(\ab[26][3] ), .B(\CARRYB[25][3] ), .CI(\SUMB[25][4] ), 
        .CO(\CARRYB[26][3] ), .S(\SUMB[26][3] ) );
  FA_X1 S2_26_4 ( .A(\ab[26][4] ), .B(\CARRYB[25][4] ), .CI(\SUMB[25][5] ), 
        .CO(\CARRYB[26][4] ), .S(\SUMB[26][4] ) );
  FA_X1 S2_26_5 ( .A(\ab[26][5] ), .B(\CARRYB[25][5] ), .CI(\SUMB[25][6] ), 
        .CO(\CARRYB[26][5] ), .S(\SUMB[26][5] ) );
  FA_X1 S2_26_6 ( .A(\ab[26][6] ), .B(\CARRYB[25][6] ), .CI(\SUMB[25][7] ), 
        .CO(\CARRYB[26][6] ), .S(\SUMB[26][6] ) );
  FA_X1 S2_26_7 ( .A(\ab[26][7] ), .B(\CARRYB[25][7] ), .CI(\SUMB[25][8] ), 
        .CO(\CARRYB[26][7] ), .S(\SUMB[26][7] ) );
  FA_X1 S2_26_8 ( .A(\ab[26][8] ), .B(\CARRYB[25][8] ), .CI(\SUMB[25][9] ), 
        .CO(\CARRYB[26][8] ), .S(\SUMB[26][8] ) );
  FA_X1 S2_26_9 ( .A(\ab[26][9] ), .B(\CARRYB[25][9] ), .CI(\SUMB[25][10] ), 
        .CO(\CARRYB[26][9] ), .S(\SUMB[26][9] ) );
  FA_X1 S2_26_10 ( .A(\ab[26][10] ), .B(\CARRYB[25][10] ), .CI(\SUMB[25][11] ), 
        .CO(\CARRYB[26][10] ), .S(\SUMB[26][10] ) );
  FA_X1 S2_26_11 ( .A(\ab[26][11] ), .B(\CARRYB[25][11] ), .CI(\SUMB[25][12] ), 
        .CO(\CARRYB[26][11] ), .S(\SUMB[26][11] ) );
  FA_X1 S2_26_12 ( .A(\ab[26][12] ), .B(\CARRYB[25][12] ), .CI(\SUMB[25][13] ), 
        .CO(\CARRYB[26][12] ), .S(\SUMB[26][12] ) );
  FA_X1 S2_26_13 ( .A(\ab[26][13] ), .B(\CARRYB[25][13] ), .CI(\SUMB[25][14] ), 
        .CO(\CARRYB[26][13] ), .S(\SUMB[26][13] ) );
  FA_X1 S2_26_14 ( .A(\ab[26][14] ), .B(\CARRYB[25][14] ), .CI(\SUMB[25][15] ), 
        .CO(\CARRYB[26][14] ), .S(\SUMB[26][14] ) );
  FA_X1 S2_26_15 ( .A(\ab[26][15] ), .B(\CARRYB[25][15] ), .CI(\SUMB[25][16] ), 
        .CO(\CARRYB[26][15] ), .S(\SUMB[26][15] ) );
  FA_X1 S2_26_16 ( .A(\ab[26][16] ), .B(\CARRYB[25][16] ), .CI(\SUMB[25][17] ), 
        .CO(\CARRYB[26][16] ), .S(\SUMB[26][16] ) );
  FA_X1 S2_26_17 ( .A(\ab[26][17] ), .B(\CARRYB[25][17] ), .CI(\SUMB[25][18] ), 
        .CO(\CARRYB[26][17] ), .S(\SUMB[26][17] ) );
  FA_X1 S2_26_18 ( .A(\ab[26][18] ), .B(\CARRYB[25][18] ), .CI(\SUMB[25][19] ), 
        .CO(\CARRYB[26][18] ), .S(\SUMB[26][18] ) );
  FA_X1 S2_26_19 ( .A(\ab[26][19] ), .B(\CARRYB[25][19] ), .CI(\SUMB[25][20] ), 
        .CO(\CARRYB[26][19] ), .S(\SUMB[26][19] ) );
  FA_X1 S2_26_20 ( .A(\ab[26][20] ), .B(\CARRYB[25][20] ), .CI(\SUMB[25][21] ), 
        .CO(\CARRYB[26][20] ), .S(\SUMB[26][20] ) );
  FA_X1 S2_26_21 ( .A(\ab[26][21] ), .B(\CARRYB[25][21] ), .CI(\SUMB[25][22] ), 
        .CO(\CARRYB[26][21] ), .S(\SUMB[26][21] ) );
  FA_X1 S2_26_22 ( .A(\ab[26][22] ), .B(\CARRYB[25][22] ), .CI(\SUMB[25][23] ), 
        .CO(\CARRYB[26][22] ), .S(\SUMB[26][22] ) );
  FA_X1 S2_26_23 ( .A(\ab[26][23] ), .B(\CARRYB[25][23] ), .CI(\SUMB[25][24] ), 
        .CO(\CARRYB[26][23] ), .S(\SUMB[26][23] ) );
  FA_X1 S2_26_24 ( .A(\ab[26][24] ), .B(\CARRYB[25][24] ), .CI(\SUMB[25][25] ), 
        .CO(\CARRYB[26][24] ), .S(\SUMB[26][24] ) );
  FA_X1 S2_26_25 ( .A(\ab[26][25] ), .B(\CARRYB[25][25] ), .CI(\SUMB[25][26] ), 
        .CO(\CARRYB[26][25] ), .S(\SUMB[26][25] ) );
  FA_X1 S2_26_26 ( .A(\ab[26][26] ), .B(\CARRYB[25][26] ), .CI(\SUMB[25][27] ), 
        .CO(\CARRYB[26][26] ), .S(\SUMB[26][26] ) );
  FA_X1 S2_26_27 ( .A(\ab[26][27] ), .B(\CARRYB[25][27] ), .CI(\SUMB[25][28] ), 
        .CO(\CARRYB[26][27] ), .S(\SUMB[26][27] ) );
  FA_X1 S2_26_28 ( .A(\ab[26][28] ), .B(\CARRYB[25][28] ), .CI(\SUMB[25][29] ), 
        .CO(\CARRYB[26][28] ), .S(\SUMB[26][28] ) );
  FA_X1 S2_26_29 ( .A(\ab[26][29] ), .B(\CARRYB[25][29] ), .CI(\SUMB[25][30] ), 
        .CO(\CARRYB[26][29] ), .S(\SUMB[26][29] ) );
  FA_X1 S2_26_30 ( .A(\ab[26][30] ), .B(\CARRYB[25][30] ), .CI(\SUMB[25][31] ), 
        .CO(\CARRYB[26][30] ), .S(\SUMB[26][30] ) );
  FA_X1 S2_26_31 ( .A(\ab[26][31] ), .B(\CARRYB[25][31] ), .CI(\SUMB[25][32] ), 
        .CO(\CARRYB[26][31] ), .S(\SUMB[26][31] ) );
  FA_X1 S2_26_32 ( .A(\ab[26][32] ), .B(\CARRYB[25][32] ), .CI(\SUMB[25][33] ), 
        .CO(\CARRYB[26][32] ), .S(\SUMB[26][32] ) );
  FA_X1 S2_26_33 ( .A(\ab[26][33] ), .B(\CARRYB[25][33] ), .CI(\SUMB[25][34] ), 
        .CO(\CARRYB[26][33] ), .S(\SUMB[26][33] ) );
  FA_X1 S2_26_34 ( .A(\ab[26][34] ), .B(\CARRYB[25][34] ), .CI(\SUMB[25][35] ), 
        .CO(\CARRYB[26][34] ), .S(\SUMB[26][34] ) );
  FA_X1 S2_26_35 ( .A(\ab[26][35] ), .B(\CARRYB[25][35] ), .CI(\SUMB[25][36] ), 
        .CO(\CARRYB[26][35] ), .S(\SUMB[26][35] ) );
  FA_X1 S2_26_36 ( .A(\ab[26][36] ), .B(\CARRYB[25][36] ), .CI(\SUMB[25][37] ), 
        .CO(\CARRYB[26][36] ), .S(\SUMB[26][36] ) );
  FA_X1 S2_26_37 ( .A(\ab[26][37] ), .B(\CARRYB[25][37] ), .CI(\SUMB[25][38] ), 
        .CO(\CARRYB[26][37] ), .S(\SUMB[26][37] ) );
  FA_X1 S2_26_38 ( .A(\ab[26][38] ), .B(\CARRYB[25][38] ), .CI(\SUMB[25][39] ), 
        .CO(\CARRYB[26][38] ), .S(\SUMB[26][38] ) );
  FA_X1 S2_26_39 ( .A(\ab[26][39] ), .B(\CARRYB[25][39] ), .CI(\SUMB[25][40] ), 
        .CO(\CARRYB[26][39] ), .S(\SUMB[26][39] ) );
  FA_X1 S2_26_40 ( .A(\ab[26][40] ), .B(\CARRYB[25][40] ), .CI(\SUMB[25][41] ), 
        .CO(\CARRYB[26][40] ), .S(\SUMB[26][40] ) );
  FA_X1 S2_26_41 ( .A(\ab[26][41] ), .B(\CARRYB[25][41] ), .CI(\SUMB[25][42] ), 
        .CO(\CARRYB[26][41] ), .S(\SUMB[26][41] ) );
  FA_X1 S2_26_42 ( .A(\ab[26][42] ), .B(\CARRYB[25][42] ), .CI(\SUMB[25][43] ), 
        .CO(\CARRYB[26][42] ), .S(\SUMB[26][42] ) );
  FA_X1 S2_26_43 ( .A(\ab[26][43] ), .B(\CARRYB[25][43] ), .CI(\SUMB[25][44] ), 
        .CO(\CARRYB[26][43] ), .S(\SUMB[26][43] ) );
  FA_X1 S2_26_44 ( .A(\ab[26][44] ), .B(\CARRYB[25][44] ), .CI(\SUMB[25][45] ), 
        .CO(\CARRYB[26][44] ), .S(\SUMB[26][44] ) );
  FA_X1 S2_26_45 ( .A(\ab[26][45] ), .B(\CARRYB[25][45] ), .CI(\SUMB[25][46] ), 
        .CO(\CARRYB[26][45] ), .S(\SUMB[26][45] ) );
  FA_X1 S2_26_46 ( .A(\ab[26][46] ), .B(\CARRYB[25][46] ), .CI(\SUMB[25][47] ), 
        .CO(\CARRYB[26][46] ), .S(\SUMB[26][46] ) );
  FA_X1 S2_26_47 ( .A(\ab[26][47] ), .B(\CARRYB[25][47] ), .CI(\SUMB[25][48] ), 
        .CO(\CARRYB[26][47] ), .S(\SUMB[26][47] ) );
  FA_X1 S2_26_48 ( .A(\ab[26][48] ), .B(\CARRYB[25][48] ), .CI(\SUMB[25][49] ), 
        .CO(\CARRYB[26][48] ), .S(\SUMB[26][48] ) );
  FA_X1 S2_26_49 ( .A(\ab[26][49] ), .B(\CARRYB[25][49] ), .CI(\SUMB[25][50] ), 
        .CO(\CARRYB[26][49] ), .S(\SUMB[26][49] ) );
  FA_X1 S2_26_50 ( .A(\ab[26][50] ), .B(\CARRYB[25][50] ), .CI(\SUMB[25][51] ), 
        .CO(\CARRYB[26][50] ), .S(\SUMB[26][50] ) );
  FA_X1 S3_26_51 ( .A(\ab[26][51] ), .B(\CARRYB[25][51] ), .CI(\ab[25][52] ), 
        .CO(\CARRYB[26][51] ), .S(\SUMB[26][51] ) );
  FA_X1 S1_25_0 ( .A(\ab[25][0] ), .B(\CARRYB[24][0] ), .CI(\SUMB[24][1] ), 
        .CO(\CARRYB[25][0] ), .S(CLA_SUM[25]) );
  FA_X1 S2_25_1 ( .A(\ab[25][1] ), .B(\CARRYB[24][1] ), .CI(\SUMB[24][2] ), 
        .CO(\CARRYB[25][1] ), .S(\SUMB[25][1] ) );
  FA_X1 S2_25_2 ( .A(\ab[25][2] ), .B(\CARRYB[24][2] ), .CI(\SUMB[24][3] ), 
        .CO(\CARRYB[25][2] ), .S(\SUMB[25][2] ) );
  FA_X1 S2_25_3 ( .A(\ab[25][3] ), .B(\CARRYB[24][3] ), .CI(\SUMB[24][4] ), 
        .CO(\CARRYB[25][3] ), .S(\SUMB[25][3] ) );
  FA_X1 S2_25_4 ( .A(\ab[25][4] ), .B(\CARRYB[24][4] ), .CI(\SUMB[24][5] ), 
        .CO(\CARRYB[25][4] ), .S(\SUMB[25][4] ) );
  FA_X1 S2_25_5 ( .A(\ab[25][5] ), .B(\CARRYB[24][5] ), .CI(\SUMB[24][6] ), 
        .CO(\CARRYB[25][5] ), .S(\SUMB[25][5] ) );
  FA_X1 S2_25_6 ( .A(\ab[25][6] ), .B(\CARRYB[24][6] ), .CI(\SUMB[24][7] ), 
        .CO(\CARRYB[25][6] ), .S(\SUMB[25][6] ) );
  FA_X1 S2_25_7 ( .A(\ab[25][7] ), .B(\CARRYB[24][7] ), .CI(\SUMB[24][8] ), 
        .CO(\CARRYB[25][7] ), .S(\SUMB[25][7] ) );
  FA_X1 S2_25_8 ( .A(\ab[25][8] ), .B(\CARRYB[24][8] ), .CI(\SUMB[24][9] ), 
        .CO(\CARRYB[25][8] ), .S(\SUMB[25][8] ) );
  FA_X1 S2_25_9 ( .A(\ab[25][9] ), .B(\CARRYB[24][9] ), .CI(\SUMB[24][10] ), 
        .CO(\CARRYB[25][9] ), .S(\SUMB[25][9] ) );
  FA_X1 S2_25_10 ( .A(\ab[25][10] ), .B(\CARRYB[24][10] ), .CI(\SUMB[24][11] ), 
        .CO(\CARRYB[25][10] ), .S(\SUMB[25][10] ) );
  FA_X1 S2_25_11 ( .A(\ab[25][11] ), .B(\CARRYB[24][11] ), .CI(\SUMB[24][12] ), 
        .CO(\CARRYB[25][11] ), .S(\SUMB[25][11] ) );
  FA_X1 S2_25_12 ( .A(\ab[25][12] ), .B(\CARRYB[24][12] ), .CI(\SUMB[24][13] ), 
        .CO(\CARRYB[25][12] ), .S(\SUMB[25][12] ) );
  FA_X1 S2_25_13 ( .A(\ab[25][13] ), .B(\CARRYB[24][13] ), .CI(\SUMB[24][14] ), 
        .CO(\CARRYB[25][13] ), .S(\SUMB[25][13] ) );
  FA_X1 S2_25_14 ( .A(\ab[25][14] ), .B(\CARRYB[24][14] ), .CI(\SUMB[24][15] ), 
        .CO(\CARRYB[25][14] ), .S(\SUMB[25][14] ) );
  FA_X1 S2_25_15 ( .A(\ab[25][15] ), .B(\CARRYB[24][15] ), .CI(\SUMB[24][16] ), 
        .CO(\CARRYB[25][15] ), .S(\SUMB[25][15] ) );
  FA_X1 S2_25_16 ( .A(\ab[25][16] ), .B(\CARRYB[24][16] ), .CI(\SUMB[24][17] ), 
        .CO(\CARRYB[25][16] ), .S(\SUMB[25][16] ) );
  FA_X1 S2_25_17 ( .A(\ab[25][17] ), .B(\CARRYB[24][17] ), .CI(\SUMB[24][18] ), 
        .CO(\CARRYB[25][17] ), .S(\SUMB[25][17] ) );
  FA_X1 S2_25_18 ( .A(\ab[25][18] ), .B(\CARRYB[24][18] ), .CI(\SUMB[24][19] ), 
        .CO(\CARRYB[25][18] ), .S(\SUMB[25][18] ) );
  FA_X1 S2_25_19 ( .A(\ab[25][19] ), .B(\CARRYB[24][19] ), .CI(\SUMB[24][20] ), 
        .CO(\CARRYB[25][19] ), .S(\SUMB[25][19] ) );
  FA_X1 S2_25_20 ( .A(\ab[25][20] ), .B(\CARRYB[24][20] ), .CI(\SUMB[24][21] ), 
        .CO(\CARRYB[25][20] ), .S(\SUMB[25][20] ) );
  FA_X1 S2_25_21 ( .A(\ab[25][21] ), .B(\CARRYB[24][21] ), .CI(\SUMB[24][22] ), 
        .CO(\CARRYB[25][21] ), .S(\SUMB[25][21] ) );
  FA_X1 S2_25_22 ( .A(\ab[25][22] ), .B(\CARRYB[24][22] ), .CI(\SUMB[24][23] ), 
        .CO(\CARRYB[25][22] ), .S(\SUMB[25][22] ) );
  FA_X1 S2_25_23 ( .A(\ab[25][23] ), .B(\CARRYB[24][23] ), .CI(\SUMB[24][24] ), 
        .CO(\CARRYB[25][23] ), .S(\SUMB[25][23] ) );
  FA_X1 S2_25_24 ( .A(\ab[25][24] ), .B(\CARRYB[24][24] ), .CI(\SUMB[24][25] ), 
        .CO(\CARRYB[25][24] ), .S(\SUMB[25][24] ) );
  FA_X1 S2_25_25 ( .A(\ab[25][25] ), .B(\CARRYB[24][25] ), .CI(\SUMB[24][26] ), 
        .CO(\CARRYB[25][25] ), .S(\SUMB[25][25] ) );
  FA_X1 S2_25_26 ( .A(\ab[25][26] ), .B(\CARRYB[24][26] ), .CI(\SUMB[24][27] ), 
        .CO(\CARRYB[25][26] ), .S(\SUMB[25][26] ) );
  FA_X1 S2_25_27 ( .A(\ab[25][27] ), .B(\CARRYB[24][27] ), .CI(\SUMB[24][28] ), 
        .CO(\CARRYB[25][27] ), .S(\SUMB[25][27] ) );
  FA_X1 S2_25_28 ( .A(\ab[25][28] ), .B(\CARRYB[24][28] ), .CI(\SUMB[24][29] ), 
        .CO(\CARRYB[25][28] ), .S(\SUMB[25][28] ) );
  FA_X1 S2_25_29 ( .A(\ab[25][29] ), .B(\CARRYB[24][29] ), .CI(\SUMB[24][30] ), 
        .CO(\CARRYB[25][29] ), .S(\SUMB[25][29] ) );
  FA_X1 S2_25_30 ( .A(\ab[25][30] ), .B(\CARRYB[24][30] ), .CI(\SUMB[24][31] ), 
        .CO(\CARRYB[25][30] ), .S(\SUMB[25][30] ) );
  FA_X1 S2_25_31 ( .A(\ab[25][31] ), .B(\CARRYB[24][31] ), .CI(\SUMB[24][32] ), 
        .CO(\CARRYB[25][31] ), .S(\SUMB[25][31] ) );
  FA_X1 S2_25_32 ( .A(\ab[25][32] ), .B(\CARRYB[24][32] ), .CI(\SUMB[24][33] ), 
        .CO(\CARRYB[25][32] ), .S(\SUMB[25][32] ) );
  FA_X1 S2_25_33 ( .A(\ab[25][33] ), .B(\CARRYB[24][33] ), .CI(\SUMB[24][34] ), 
        .CO(\CARRYB[25][33] ), .S(\SUMB[25][33] ) );
  FA_X1 S2_25_34 ( .A(\ab[25][34] ), .B(\CARRYB[24][34] ), .CI(\SUMB[24][35] ), 
        .CO(\CARRYB[25][34] ), .S(\SUMB[25][34] ) );
  FA_X1 S2_25_35 ( .A(\ab[25][35] ), .B(\CARRYB[24][35] ), .CI(\SUMB[24][36] ), 
        .CO(\CARRYB[25][35] ), .S(\SUMB[25][35] ) );
  FA_X1 S2_25_36 ( .A(\ab[25][36] ), .B(\CARRYB[24][36] ), .CI(\SUMB[24][37] ), 
        .CO(\CARRYB[25][36] ), .S(\SUMB[25][36] ) );
  FA_X1 S2_25_37 ( .A(\ab[25][37] ), .B(\CARRYB[24][37] ), .CI(\SUMB[24][38] ), 
        .CO(\CARRYB[25][37] ), .S(\SUMB[25][37] ) );
  FA_X1 S2_25_38 ( .A(\ab[25][38] ), .B(\CARRYB[24][38] ), .CI(\SUMB[24][39] ), 
        .CO(\CARRYB[25][38] ), .S(\SUMB[25][38] ) );
  FA_X1 S2_25_39 ( .A(\ab[25][39] ), .B(\CARRYB[24][39] ), .CI(\SUMB[24][40] ), 
        .CO(\CARRYB[25][39] ), .S(\SUMB[25][39] ) );
  FA_X1 S2_25_40 ( .A(\ab[25][40] ), .B(\CARRYB[24][40] ), .CI(\SUMB[24][41] ), 
        .CO(\CARRYB[25][40] ), .S(\SUMB[25][40] ) );
  FA_X1 S2_25_41 ( .A(\ab[25][41] ), .B(\CARRYB[24][41] ), .CI(\SUMB[24][42] ), 
        .CO(\CARRYB[25][41] ), .S(\SUMB[25][41] ) );
  FA_X1 S2_25_42 ( .A(\ab[25][42] ), .B(\CARRYB[24][42] ), .CI(\SUMB[24][43] ), 
        .CO(\CARRYB[25][42] ), .S(\SUMB[25][42] ) );
  FA_X1 S2_25_43 ( .A(\ab[25][43] ), .B(\CARRYB[24][43] ), .CI(\SUMB[24][44] ), 
        .CO(\CARRYB[25][43] ), .S(\SUMB[25][43] ) );
  FA_X1 S2_25_44 ( .A(\ab[25][44] ), .B(\CARRYB[24][44] ), .CI(\SUMB[24][45] ), 
        .CO(\CARRYB[25][44] ), .S(\SUMB[25][44] ) );
  FA_X1 S2_25_45 ( .A(\ab[25][45] ), .B(\CARRYB[24][45] ), .CI(\SUMB[24][46] ), 
        .CO(\CARRYB[25][45] ), .S(\SUMB[25][45] ) );
  FA_X1 S2_25_46 ( .A(\ab[25][46] ), .B(\CARRYB[24][46] ), .CI(\SUMB[24][47] ), 
        .CO(\CARRYB[25][46] ), .S(\SUMB[25][46] ) );
  FA_X1 S2_25_47 ( .A(\ab[25][47] ), .B(\CARRYB[24][47] ), .CI(\SUMB[24][48] ), 
        .CO(\CARRYB[25][47] ), .S(\SUMB[25][47] ) );
  FA_X1 S2_25_48 ( .A(\ab[25][48] ), .B(\CARRYB[24][48] ), .CI(\SUMB[24][49] ), 
        .CO(\CARRYB[25][48] ), .S(\SUMB[25][48] ) );
  FA_X1 S2_25_49 ( .A(\ab[25][49] ), .B(\CARRYB[24][49] ), .CI(\SUMB[24][50] ), 
        .CO(\CARRYB[25][49] ), .S(\SUMB[25][49] ) );
  FA_X1 S2_25_50 ( .A(\ab[25][50] ), .B(\CARRYB[24][50] ), .CI(\SUMB[24][51] ), 
        .CO(\CARRYB[25][50] ), .S(\SUMB[25][50] ) );
  FA_X1 S3_25_51 ( .A(\ab[25][51] ), .B(\CARRYB[24][51] ), .CI(\ab[24][52] ), 
        .CO(\CARRYB[25][51] ), .S(\SUMB[25][51] ) );
  FA_X1 S1_24_0 ( .A(\ab[24][0] ), .B(\CARRYB[23][0] ), .CI(\SUMB[23][1] ), 
        .CO(\CARRYB[24][0] ), .S(CLA_SUM[24]) );
  FA_X1 S2_24_1 ( .A(\ab[24][1] ), .B(\CARRYB[23][1] ), .CI(\SUMB[23][2] ), 
        .CO(\CARRYB[24][1] ), .S(\SUMB[24][1] ) );
  FA_X1 S2_24_2 ( .A(\ab[24][2] ), .B(\CARRYB[23][2] ), .CI(\SUMB[23][3] ), 
        .CO(\CARRYB[24][2] ), .S(\SUMB[24][2] ) );
  FA_X1 S2_24_3 ( .A(\ab[24][3] ), .B(\CARRYB[23][3] ), .CI(\SUMB[23][4] ), 
        .CO(\CARRYB[24][3] ), .S(\SUMB[24][3] ) );
  FA_X1 S2_24_4 ( .A(\ab[24][4] ), .B(\CARRYB[23][4] ), .CI(\SUMB[23][5] ), 
        .CO(\CARRYB[24][4] ), .S(\SUMB[24][4] ) );
  FA_X1 S2_24_5 ( .A(\ab[24][5] ), .B(\CARRYB[23][5] ), .CI(\SUMB[23][6] ), 
        .CO(\CARRYB[24][5] ), .S(\SUMB[24][5] ) );
  FA_X1 S2_24_6 ( .A(\ab[24][6] ), .B(\CARRYB[23][6] ), .CI(\SUMB[23][7] ), 
        .CO(\CARRYB[24][6] ), .S(\SUMB[24][6] ) );
  FA_X1 S2_24_7 ( .A(\ab[24][7] ), .B(\CARRYB[23][7] ), .CI(\SUMB[23][8] ), 
        .CO(\CARRYB[24][7] ), .S(\SUMB[24][7] ) );
  FA_X1 S2_24_8 ( .A(\ab[24][8] ), .B(\CARRYB[23][8] ), .CI(\SUMB[23][9] ), 
        .CO(\CARRYB[24][8] ), .S(\SUMB[24][8] ) );
  FA_X1 S2_24_9 ( .A(\ab[24][9] ), .B(\CARRYB[23][9] ), .CI(\SUMB[23][10] ), 
        .CO(\CARRYB[24][9] ), .S(\SUMB[24][9] ) );
  FA_X1 S2_24_10 ( .A(\ab[24][10] ), .B(\CARRYB[23][10] ), .CI(\SUMB[23][11] ), 
        .CO(\CARRYB[24][10] ), .S(\SUMB[24][10] ) );
  FA_X1 S2_24_11 ( .A(\ab[24][11] ), .B(\CARRYB[23][11] ), .CI(\SUMB[23][12] ), 
        .CO(\CARRYB[24][11] ), .S(\SUMB[24][11] ) );
  FA_X1 S2_24_12 ( .A(\ab[24][12] ), .B(\CARRYB[23][12] ), .CI(\SUMB[23][13] ), 
        .CO(\CARRYB[24][12] ), .S(\SUMB[24][12] ) );
  FA_X1 S2_24_13 ( .A(\ab[24][13] ), .B(\CARRYB[23][13] ), .CI(\SUMB[23][14] ), 
        .CO(\CARRYB[24][13] ), .S(\SUMB[24][13] ) );
  FA_X1 S2_24_14 ( .A(\ab[24][14] ), .B(\CARRYB[23][14] ), .CI(\SUMB[23][15] ), 
        .CO(\CARRYB[24][14] ), .S(\SUMB[24][14] ) );
  FA_X1 S2_24_15 ( .A(\ab[24][15] ), .B(\CARRYB[23][15] ), .CI(\SUMB[23][16] ), 
        .CO(\CARRYB[24][15] ), .S(\SUMB[24][15] ) );
  FA_X1 S2_24_16 ( .A(\ab[24][16] ), .B(\CARRYB[23][16] ), .CI(\SUMB[23][17] ), 
        .CO(\CARRYB[24][16] ), .S(\SUMB[24][16] ) );
  FA_X1 S2_24_17 ( .A(\ab[24][17] ), .B(\CARRYB[23][17] ), .CI(\SUMB[23][18] ), 
        .CO(\CARRYB[24][17] ), .S(\SUMB[24][17] ) );
  FA_X1 S2_24_18 ( .A(\ab[24][18] ), .B(\CARRYB[23][18] ), .CI(\SUMB[23][19] ), 
        .CO(\CARRYB[24][18] ), .S(\SUMB[24][18] ) );
  FA_X1 S2_24_19 ( .A(\ab[24][19] ), .B(\CARRYB[23][19] ), .CI(\SUMB[23][20] ), 
        .CO(\CARRYB[24][19] ), .S(\SUMB[24][19] ) );
  FA_X1 S2_24_20 ( .A(\ab[24][20] ), .B(\CARRYB[23][20] ), .CI(\SUMB[23][21] ), 
        .CO(\CARRYB[24][20] ), .S(\SUMB[24][20] ) );
  FA_X1 S2_24_21 ( .A(\ab[24][21] ), .B(\CARRYB[23][21] ), .CI(\SUMB[23][22] ), 
        .CO(\CARRYB[24][21] ), .S(\SUMB[24][21] ) );
  FA_X1 S2_24_22 ( .A(\ab[24][22] ), .B(\CARRYB[23][22] ), .CI(\SUMB[23][23] ), 
        .CO(\CARRYB[24][22] ), .S(\SUMB[24][22] ) );
  FA_X1 S2_24_23 ( .A(\ab[24][23] ), .B(\CARRYB[23][23] ), .CI(\SUMB[23][24] ), 
        .CO(\CARRYB[24][23] ), .S(\SUMB[24][23] ) );
  FA_X1 S2_24_24 ( .A(\ab[24][24] ), .B(\CARRYB[23][24] ), .CI(\SUMB[23][25] ), 
        .CO(\CARRYB[24][24] ), .S(\SUMB[24][24] ) );
  FA_X1 S2_24_25 ( .A(\ab[24][25] ), .B(\CARRYB[23][25] ), .CI(\SUMB[23][26] ), 
        .CO(\CARRYB[24][25] ), .S(\SUMB[24][25] ) );
  FA_X1 S2_24_26 ( .A(\ab[24][26] ), .B(\CARRYB[23][26] ), .CI(\SUMB[23][27] ), 
        .CO(\CARRYB[24][26] ), .S(\SUMB[24][26] ) );
  FA_X1 S2_24_27 ( .A(\ab[24][27] ), .B(\CARRYB[23][27] ), .CI(\SUMB[23][28] ), 
        .CO(\CARRYB[24][27] ), .S(\SUMB[24][27] ) );
  FA_X1 S2_24_28 ( .A(\ab[24][28] ), .B(\CARRYB[23][28] ), .CI(\SUMB[23][29] ), 
        .CO(\CARRYB[24][28] ), .S(\SUMB[24][28] ) );
  FA_X1 S2_24_29 ( .A(\ab[24][29] ), .B(\CARRYB[23][29] ), .CI(\SUMB[23][30] ), 
        .CO(\CARRYB[24][29] ), .S(\SUMB[24][29] ) );
  FA_X1 S2_24_30 ( .A(\ab[24][30] ), .B(\CARRYB[23][30] ), .CI(\SUMB[23][31] ), 
        .CO(\CARRYB[24][30] ), .S(\SUMB[24][30] ) );
  FA_X1 S2_24_31 ( .A(\ab[24][31] ), .B(\CARRYB[23][31] ), .CI(\SUMB[23][32] ), 
        .CO(\CARRYB[24][31] ), .S(\SUMB[24][31] ) );
  FA_X1 S2_24_32 ( .A(\ab[24][32] ), .B(\CARRYB[23][32] ), .CI(\SUMB[23][33] ), 
        .CO(\CARRYB[24][32] ), .S(\SUMB[24][32] ) );
  FA_X1 S2_24_33 ( .A(\ab[24][33] ), .B(\CARRYB[23][33] ), .CI(\SUMB[23][34] ), 
        .CO(\CARRYB[24][33] ), .S(\SUMB[24][33] ) );
  FA_X1 S2_24_34 ( .A(\ab[24][34] ), .B(\CARRYB[23][34] ), .CI(\SUMB[23][35] ), 
        .CO(\CARRYB[24][34] ), .S(\SUMB[24][34] ) );
  FA_X1 S2_24_35 ( .A(\ab[24][35] ), .B(\CARRYB[23][35] ), .CI(\SUMB[23][36] ), 
        .CO(\CARRYB[24][35] ), .S(\SUMB[24][35] ) );
  FA_X1 S2_24_36 ( .A(\ab[24][36] ), .B(\CARRYB[23][36] ), .CI(\SUMB[23][37] ), 
        .CO(\CARRYB[24][36] ), .S(\SUMB[24][36] ) );
  FA_X1 S2_24_37 ( .A(\ab[24][37] ), .B(\CARRYB[23][37] ), .CI(\SUMB[23][38] ), 
        .CO(\CARRYB[24][37] ), .S(\SUMB[24][37] ) );
  FA_X1 S2_24_38 ( .A(\ab[24][38] ), .B(\CARRYB[23][38] ), .CI(\SUMB[23][39] ), 
        .CO(\CARRYB[24][38] ), .S(\SUMB[24][38] ) );
  FA_X1 S2_24_39 ( .A(\ab[24][39] ), .B(\CARRYB[23][39] ), .CI(\SUMB[23][40] ), 
        .CO(\CARRYB[24][39] ), .S(\SUMB[24][39] ) );
  FA_X1 S2_24_40 ( .A(\ab[24][40] ), .B(\CARRYB[23][40] ), .CI(\SUMB[23][41] ), 
        .CO(\CARRYB[24][40] ), .S(\SUMB[24][40] ) );
  FA_X1 S2_24_41 ( .A(\ab[24][41] ), .B(\CARRYB[23][41] ), .CI(\SUMB[23][42] ), 
        .CO(\CARRYB[24][41] ), .S(\SUMB[24][41] ) );
  FA_X1 S2_24_42 ( .A(\ab[24][42] ), .B(\CARRYB[23][42] ), .CI(\SUMB[23][43] ), 
        .CO(\CARRYB[24][42] ), .S(\SUMB[24][42] ) );
  FA_X1 S2_24_43 ( .A(\ab[24][43] ), .B(\CARRYB[23][43] ), .CI(\SUMB[23][44] ), 
        .CO(\CARRYB[24][43] ), .S(\SUMB[24][43] ) );
  FA_X1 S2_24_44 ( .A(\ab[24][44] ), .B(\CARRYB[23][44] ), .CI(\SUMB[23][45] ), 
        .CO(\CARRYB[24][44] ), .S(\SUMB[24][44] ) );
  FA_X1 S2_24_45 ( .A(\ab[24][45] ), .B(\CARRYB[23][45] ), .CI(\SUMB[23][46] ), 
        .CO(\CARRYB[24][45] ), .S(\SUMB[24][45] ) );
  FA_X1 S2_24_46 ( .A(\ab[24][46] ), .B(\CARRYB[23][46] ), .CI(\SUMB[23][47] ), 
        .CO(\CARRYB[24][46] ), .S(\SUMB[24][46] ) );
  FA_X1 S2_24_47 ( .A(\ab[24][47] ), .B(\CARRYB[23][47] ), .CI(\SUMB[23][48] ), 
        .CO(\CARRYB[24][47] ), .S(\SUMB[24][47] ) );
  FA_X1 S2_24_48 ( .A(\ab[24][48] ), .B(\CARRYB[23][48] ), .CI(\SUMB[23][49] ), 
        .CO(\CARRYB[24][48] ), .S(\SUMB[24][48] ) );
  FA_X1 S2_24_49 ( .A(\ab[24][49] ), .B(\CARRYB[23][49] ), .CI(\SUMB[23][50] ), 
        .CO(\CARRYB[24][49] ), .S(\SUMB[24][49] ) );
  FA_X1 S2_24_50 ( .A(\ab[24][50] ), .B(\CARRYB[23][50] ), .CI(\SUMB[23][51] ), 
        .CO(\CARRYB[24][50] ), .S(\SUMB[24][50] ) );
  FA_X1 S3_24_51 ( .A(\ab[24][51] ), .B(\CARRYB[23][51] ), .CI(\ab[23][52] ), 
        .CO(\CARRYB[24][51] ), .S(\SUMB[24][51] ) );
  FA_X1 S1_23_0 ( .A(\ab[23][0] ), .B(\CARRYB[22][0] ), .CI(\SUMB[22][1] ), 
        .CO(\CARRYB[23][0] ), .S(CLA_SUM[23]) );
  FA_X1 S2_23_1 ( .A(\ab[23][1] ), .B(\CARRYB[22][1] ), .CI(\SUMB[22][2] ), 
        .CO(\CARRYB[23][1] ), .S(\SUMB[23][1] ) );
  FA_X1 S2_23_2 ( .A(\ab[23][2] ), .B(\CARRYB[22][2] ), .CI(\SUMB[22][3] ), 
        .CO(\CARRYB[23][2] ), .S(\SUMB[23][2] ) );
  FA_X1 S2_23_3 ( .A(\ab[23][3] ), .B(\CARRYB[22][3] ), .CI(\SUMB[22][4] ), 
        .CO(\CARRYB[23][3] ), .S(\SUMB[23][3] ) );
  FA_X1 S2_23_4 ( .A(\ab[23][4] ), .B(\CARRYB[22][4] ), .CI(\SUMB[22][5] ), 
        .CO(\CARRYB[23][4] ), .S(\SUMB[23][4] ) );
  FA_X1 S2_23_5 ( .A(\ab[23][5] ), .B(\CARRYB[22][5] ), .CI(\SUMB[22][6] ), 
        .CO(\CARRYB[23][5] ), .S(\SUMB[23][5] ) );
  FA_X1 S2_23_6 ( .A(\ab[23][6] ), .B(\CARRYB[22][6] ), .CI(\SUMB[22][7] ), 
        .CO(\CARRYB[23][6] ), .S(\SUMB[23][6] ) );
  FA_X1 S2_23_7 ( .A(\ab[23][7] ), .B(\CARRYB[22][7] ), .CI(\SUMB[22][8] ), 
        .CO(\CARRYB[23][7] ), .S(\SUMB[23][7] ) );
  FA_X1 S2_23_8 ( .A(\ab[23][8] ), .B(\CARRYB[22][8] ), .CI(\SUMB[22][9] ), 
        .CO(\CARRYB[23][8] ), .S(\SUMB[23][8] ) );
  FA_X1 S2_23_9 ( .A(\ab[23][9] ), .B(\CARRYB[22][9] ), .CI(\SUMB[22][10] ), 
        .CO(\CARRYB[23][9] ), .S(\SUMB[23][9] ) );
  FA_X1 S2_23_10 ( .A(\ab[23][10] ), .B(\CARRYB[22][10] ), .CI(\SUMB[22][11] ), 
        .CO(\CARRYB[23][10] ), .S(\SUMB[23][10] ) );
  FA_X1 S2_23_11 ( .A(\ab[23][11] ), .B(\CARRYB[22][11] ), .CI(\SUMB[22][12] ), 
        .CO(\CARRYB[23][11] ), .S(\SUMB[23][11] ) );
  FA_X1 S2_23_12 ( .A(\ab[23][12] ), .B(\CARRYB[22][12] ), .CI(\SUMB[22][13] ), 
        .CO(\CARRYB[23][12] ), .S(\SUMB[23][12] ) );
  FA_X1 S2_23_13 ( .A(\ab[23][13] ), .B(\CARRYB[22][13] ), .CI(\SUMB[22][14] ), 
        .CO(\CARRYB[23][13] ), .S(\SUMB[23][13] ) );
  FA_X1 S2_23_14 ( .A(\ab[23][14] ), .B(\CARRYB[22][14] ), .CI(\SUMB[22][15] ), 
        .CO(\CARRYB[23][14] ), .S(\SUMB[23][14] ) );
  FA_X1 S2_23_15 ( .A(\ab[23][15] ), .B(\CARRYB[22][15] ), .CI(\SUMB[22][16] ), 
        .CO(\CARRYB[23][15] ), .S(\SUMB[23][15] ) );
  FA_X1 S2_23_16 ( .A(\ab[23][16] ), .B(\CARRYB[22][16] ), .CI(\SUMB[22][17] ), 
        .CO(\CARRYB[23][16] ), .S(\SUMB[23][16] ) );
  FA_X1 S2_23_17 ( .A(\ab[23][17] ), .B(\CARRYB[22][17] ), .CI(\SUMB[22][18] ), 
        .CO(\CARRYB[23][17] ), .S(\SUMB[23][17] ) );
  FA_X1 S2_23_18 ( .A(\ab[23][18] ), .B(\CARRYB[22][18] ), .CI(\SUMB[22][19] ), 
        .CO(\CARRYB[23][18] ), .S(\SUMB[23][18] ) );
  FA_X1 S2_23_19 ( .A(\ab[23][19] ), .B(\CARRYB[22][19] ), .CI(\SUMB[22][20] ), 
        .CO(\CARRYB[23][19] ), .S(\SUMB[23][19] ) );
  FA_X1 S2_23_20 ( .A(\ab[23][20] ), .B(\CARRYB[22][20] ), .CI(\SUMB[22][21] ), 
        .CO(\CARRYB[23][20] ), .S(\SUMB[23][20] ) );
  FA_X1 S2_23_21 ( .A(\ab[23][21] ), .B(\CARRYB[22][21] ), .CI(\SUMB[22][22] ), 
        .CO(\CARRYB[23][21] ), .S(\SUMB[23][21] ) );
  FA_X1 S2_23_22 ( .A(\ab[23][22] ), .B(\CARRYB[22][22] ), .CI(\SUMB[22][23] ), 
        .CO(\CARRYB[23][22] ), .S(\SUMB[23][22] ) );
  FA_X1 S2_23_23 ( .A(\ab[23][23] ), .B(\CARRYB[22][23] ), .CI(\SUMB[22][24] ), 
        .CO(\CARRYB[23][23] ), .S(\SUMB[23][23] ) );
  FA_X1 S2_23_24 ( .A(\ab[23][24] ), .B(\CARRYB[22][24] ), .CI(\SUMB[22][25] ), 
        .CO(\CARRYB[23][24] ), .S(\SUMB[23][24] ) );
  FA_X1 S2_23_25 ( .A(\ab[23][25] ), .B(\CARRYB[22][25] ), .CI(\SUMB[22][26] ), 
        .CO(\CARRYB[23][25] ), .S(\SUMB[23][25] ) );
  FA_X1 S2_23_26 ( .A(\ab[23][26] ), .B(\CARRYB[22][26] ), .CI(\SUMB[22][27] ), 
        .CO(\CARRYB[23][26] ), .S(\SUMB[23][26] ) );
  FA_X1 S2_23_27 ( .A(\ab[23][27] ), .B(\CARRYB[22][27] ), .CI(\SUMB[22][28] ), 
        .CO(\CARRYB[23][27] ), .S(\SUMB[23][27] ) );
  FA_X1 S2_23_28 ( .A(\ab[23][28] ), .B(\CARRYB[22][28] ), .CI(\SUMB[22][29] ), 
        .CO(\CARRYB[23][28] ), .S(\SUMB[23][28] ) );
  FA_X1 S2_23_29 ( .A(\ab[23][29] ), .B(\CARRYB[22][29] ), .CI(\SUMB[22][30] ), 
        .CO(\CARRYB[23][29] ), .S(\SUMB[23][29] ) );
  FA_X1 S2_23_30 ( .A(\ab[23][30] ), .B(\CARRYB[22][30] ), .CI(\SUMB[22][31] ), 
        .CO(\CARRYB[23][30] ), .S(\SUMB[23][30] ) );
  FA_X1 S2_23_31 ( .A(\ab[23][31] ), .B(\CARRYB[22][31] ), .CI(\SUMB[22][32] ), 
        .CO(\CARRYB[23][31] ), .S(\SUMB[23][31] ) );
  FA_X1 S2_23_32 ( .A(\ab[23][32] ), .B(\CARRYB[22][32] ), .CI(\SUMB[22][33] ), 
        .CO(\CARRYB[23][32] ), .S(\SUMB[23][32] ) );
  FA_X1 S2_23_33 ( .A(\ab[23][33] ), .B(\CARRYB[22][33] ), .CI(\SUMB[22][34] ), 
        .CO(\CARRYB[23][33] ), .S(\SUMB[23][33] ) );
  FA_X1 S2_23_34 ( .A(\ab[23][34] ), .B(\CARRYB[22][34] ), .CI(\SUMB[22][35] ), 
        .CO(\CARRYB[23][34] ), .S(\SUMB[23][34] ) );
  FA_X1 S2_23_35 ( .A(\ab[23][35] ), .B(\CARRYB[22][35] ), .CI(\SUMB[22][36] ), 
        .CO(\CARRYB[23][35] ), .S(\SUMB[23][35] ) );
  FA_X1 S2_23_36 ( .A(\ab[23][36] ), .B(\CARRYB[22][36] ), .CI(\SUMB[22][37] ), 
        .CO(\CARRYB[23][36] ), .S(\SUMB[23][36] ) );
  FA_X1 S2_23_37 ( .A(\ab[23][37] ), .B(\CARRYB[22][37] ), .CI(\SUMB[22][38] ), 
        .CO(\CARRYB[23][37] ), .S(\SUMB[23][37] ) );
  FA_X1 S2_23_38 ( .A(\ab[23][38] ), .B(\CARRYB[22][38] ), .CI(\SUMB[22][39] ), 
        .CO(\CARRYB[23][38] ), .S(\SUMB[23][38] ) );
  FA_X1 S2_23_39 ( .A(\ab[23][39] ), .B(\CARRYB[22][39] ), .CI(\SUMB[22][40] ), 
        .CO(\CARRYB[23][39] ), .S(\SUMB[23][39] ) );
  FA_X1 S2_23_40 ( .A(\ab[23][40] ), .B(\CARRYB[22][40] ), .CI(\SUMB[22][41] ), 
        .CO(\CARRYB[23][40] ), .S(\SUMB[23][40] ) );
  FA_X1 S2_23_41 ( .A(\ab[23][41] ), .B(\CARRYB[22][41] ), .CI(\SUMB[22][42] ), 
        .CO(\CARRYB[23][41] ), .S(\SUMB[23][41] ) );
  FA_X1 S2_23_42 ( .A(\ab[23][42] ), .B(\CARRYB[22][42] ), .CI(\SUMB[22][43] ), 
        .CO(\CARRYB[23][42] ), .S(\SUMB[23][42] ) );
  FA_X1 S2_23_43 ( .A(\ab[23][43] ), .B(\CARRYB[22][43] ), .CI(\SUMB[22][44] ), 
        .CO(\CARRYB[23][43] ), .S(\SUMB[23][43] ) );
  FA_X1 S2_23_44 ( .A(\ab[23][44] ), .B(\CARRYB[22][44] ), .CI(\SUMB[22][45] ), 
        .CO(\CARRYB[23][44] ), .S(\SUMB[23][44] ) );
  FA_X1 S2_23_45 ( .A(\ab[23][45] ), .B(\CARRYB[22][45] ), .CI(\SUMB[22][46] ), 
        .CO(\CARRYB[23][45] ), .S(\SUMB[23][45] ) );
  FA_X1 S2_23_46 ( .A(\ab[23][46] ), .B(\CARRYB[22][46] ), .CI(\SUMB[22][47] ), 
        .CO(\CARRYB[23][46] ), .S(\SUMB[23][46] ) );
  FA_X1 S2_23_47 ( .A(\ab[23][47] ), .B(\CARRYB[22][47] ), .CI(\SUMB[22][48] ), 
        .CO(\CARRYB[23][47] ), .S(\SUMB[23][47] ) );
  FA_X1 S2_23_48 ( .A(\ab[23][48] ), .B(\CARRYB[22][48] ), .CI(\SUMB[22][49] ), 
        .CO(\CARRYB[23][48] ), .S(\SUMB[23][48] ) );
  FA_X1 S2_23_49 ( .A(\ab[23][49] ), .B(\CARRYB[22][49] ), .CI(\SUMB[22][50] ), 
        .CO(\CARRYB[23][49] ), .S(\SUMB[23][49] ) );
  FA_X1 S2_23_50 ( .A(\ab[23][50] ), .B(\CARRYB[22][50] ), .CI(\SUMB[22][51] ), 
        .CO(\CARRYB[23][50] ), .S(\SUMB[23][50] ) );
  FA_X1 S3_23_51 ( .A(\ab[23][51] ), .B(\CARRYB[22][51] ), .CI(\ab[22][52] ), 
        .CO(\CARRYB[23][51] ), .S(\SUMB[23][51] ) );
  FA_X1 S1_22_0 ( .A(\ab[22][0] ), .B(\CARRYB[21][0] ), .CI(\SUMB[21][1] ), 
        .CO(\CARRYB[22][0] ), .S(CLA_SUM[22]) );
  FA_X1 S2_22_1 ( .A(\ab[22][1] ), .B(\CARRYB[21][1] ), .CI(\SUMB[21][2] ), 
        .CO(\CARRYB[22][1] ), .S(\SUMB[22][1] ) );
  FA_X1 S2_22_2 ( .A(\ab[22][2] ), .B(\CARRYB[21][2] ), .CI(\SUMB[21][3] ), 
        .CO(\CARRYB[22][2] ), .S(\SUMB[22][2] ) );
  FA_X1 S2_22_3 ( .A(\ab[22][3] ), .B(\CARRYB[21][3] ), .CI(\SUMB[21][4] ), 
        .CO(\CARRYB[22][3] ), .S(\SUMB[22][3] ) );
  FA_X1 S2_22_4 ( .A(\ab[22][4] ), .B(\CARRYB[21][4] ), .CI(\SUMB[21][5] ), 
        .CO(\CARRYB[22][4] ), .S(\SUMB[22][4] ) );
  FA_X1 S2_22_5 ( .A(\ab[22][5] ), .B(\CARRYB[21][5] ), .CI(\SUMB[21][6] ), 
        .CO(\CARRYB[22][5] ), .S(\SUMB[22][5] ) );
  FA_X1 S2_22_6 ( .A(\ab[22][6] ), .B(\CARRYB[21][6] ), .CI(\SUMB[21][7] ), 
        .CO(\CARRYB[22][6] ), .S(\SUMB[22][6] ) );
  FA_X1 S2_22_7 ( .A(\ab[22][7] ), .B(\CARRYB[21][7] ), .CI(\SUMB[21][8] ), 
        .CO(\CARRYB[22][7] ), .S(\SUMB[22][7] ) );
  FA_X1 S2_22_8 ( .A(\ab[22][8] ), .B(\CARRYB[21][8] ), .CI(\SUMB[21][9] ), 
        .CO(\CARRYB[22][8] ), .S(\SUMB[22][8] ) );
  FA_X1 S2_22_9 ( .A(\ab[22][9] ), .B(\CARRYB[21][9] ), .CI(\SUMB[21][10] ), 
        .CO(\CARRYB[22][9] ), .S(\SUMB[22][9] ) );
  FA_X1 S2_22_10 ( .A(\ab[22][10] ), .B(\CARRYB[21][10] ), .CI(\SUMB[21][11] ), 
        .CO(\CARRYB[22][10] ), .S(\SUMB[22][10] ) );
  FA_X1 S2_22_11 ( .A(\ab[22][11] ), .B(\CARRYB[21][11] ), .CI(\SUMB[21][12] ), 
        .CO(\CARRYB[22][11] ), .S(\SUMB[22][11] ) );
  FA_X1 S2_22_12 ( .A(\ab[22][12] ), .B(\CARRYB[21][12] ), .CI(\SUMB[21][13] ), 
        .CO(\CARRYB[22][12] ), .S(\SUMB[22][12] ) );
  FA_X1 S2_22_13 ( .A(\ab[22][13] ), .B(\CARRYB[21][13] ), .CI(\SUMB[21][14] ), 
        .CO(\CARRYB[22][13] ), .S(\SUMB[22][13] ) );
  FA_X1 S2_22_14 ( .A(\ab[22][14] ), .B(\CARRYB[21][14] ), .CI(\SUMB[21][15] ), 
        .CO(\CARRYB[22][14] ), .S(\SUMB[22][14] ) );
  FA_X1 S2_22_15 ( .A(\ab[22][15] ), .B(\CARRYB[21][15] ), .CI(\SUMB[21][16] ), 
        .CO(\CARRYB[22][15] ), .S(\SUMB[22][15] ) );
  FA_X1 S2_22_16 ( .A(\ab[22][16] ), .B(\CARRYB[21][16] ), .CI(\SUMB[21][17] ), 
        .CO(\CARRYB[22][16] ), .S(\SUMB[22][16] ) );
  FA_X1 S2_22_17 ( .A(\ab[22][17] ), .B(\CARRYB[21][17] ), .CI(\SUMB[21][18] ), 
        .CO(\CARRYB[22][17] ), .S(\SUMB[22][17] ) );
  FA_X1 S2_22_18 ( .A(\ab[22][18] ), .B(\CARRYB[21][18] ), .CI(\SUMB[21][19] ), 
        .CO(\CARRYB[22][18] ), .S(\SUMB[22][18] ) );
  FA_X1 S2_22_19 ( .A(\ab[22][19] ), .B(\CARRYB[21][19] ), .CI(\SUMB[21][20] ), 
        .CO(\CARRYB[22][19] ), .S(\SUMB[22][19] ) );
  FA_X1 S2_22_20 ( .A(\ab[22][20] ), .B(\CARRYB[21][20] ), .CI(\SUMB[21][21] ), 
        .CO(\CARRYB[22][20] ), .S(\SUMB[22][20] ) );
  FA_X1 S2_22_21 ( .A(\ab[22][21] ), .B(\CARRYB[21][21] ), .CI(\SUMB[21][22] ), 
        .CO(\CARRYB[22][21] ), .S(\SUMB[22][21] ) );
  FA_X1 S2_22_22 ( .A(\ab[22][22] ), .B(\CARRYB[21][22] ), .CI(\SUMB[21][23] ), 
        .CO(\CARRYB[22][22] ), .S(\SUMB[22][22] ) );
  FA_X1 S2_22_23 ( .A(\ab[22][23] ), .B(\CARRYB[21][23] ), .CI(\SUMB[21][24] ), 
        .CO(\CARRYB[22][23] ), .S(\SUMB[22][23] ) );
  FA_X1 S2_22_24 ( .A(\ab[22][24] ), .B(\CARRYB[21][24] ), .CI(\SUMB[21][25] ), 
        .CO(\CARRYB[22][24] ), .S(\SUMB[22][24] ) );
  FA_X1 S2_22_25 ( .A(\ab[22][25] ), .B(\CARRYB[21][25] ), .CI(\SUMB[21][26] ), 
        .CO(\CARRYB[22][25] ), .S(\SUMB[22][25] ) );
  FA_X1 S2_22_26 ( .A(\ab[22][26] ), .B(\CARRYB[21][26] ), .CI(\SUMB[21][27] ), 
        .CO(\CARRYB[22][26] ), .S(\SUMB[22][26] ) );
  FA_X1 S2_22_27 ( .A(\ab[22][27] ), .B(\CARRYB[21][27] ), .CI(\SUMB[21][28] ), 
        .CO(\CARRYB[22][27] ), .S(\SUMB[22][27] ) );
  FA_X1 S2_22_28 ( .A(\ab[22][28] ), .B(\CARRYB[21][28] ), .CI(\SUMB[21][29] ), 
        .CO(\CARRYB[22][28] ), .S(\SUMB[22][28] ) );
  FA_X1 S2_22_29 ( .A(\ab[22][29] ), .B(\CARRYB[21][29] ), .CI(\SUMB[21][30] ), 
        .CO(\CARRYB[22][29] ), .S(\SUMB[22][29] ) );
  FA_X1 S2_22_30 ( .A(\ab[22][30] ), .B(\CARRYB[21][30] ), .CI(\SUMB[21][31] ), 
        .CO(\CARRYB[22][30] ), .S(\SUMB[22][30] ) );
  FA_X1 S2_22_31 ( .A(\ab[22][31] ), .B(\CARRYB[21][31] ), .CI(\SUMB[21][32] ), 
        .CO(\CARRYB[22][31] ), .S(\SUMB[22][31] ) );
  FA_X1 S2_22_32 ( .A(\ab[22][32] ), .B(\CARRYB[21][32] ), .CI(\SUMB[21][33] ), 
        .CO(\CARRYB[22][32] ), .S(\SUMB[22][32] ) );
  FA_X1 S2_22_33 ( .A(\ab[22][33] ), .B(\CARRYB[21][33] ), .CI(\SUMB[21][34] ), 
        .CO(\CARRYB[22][33] ), .S(\SUMB[22][33] ) );
  FA_X1 S2_22_34 ( .A(\ab[22][34] ), .B(\CARRYB[21][34] ), .CI(\SUMB[21][35] ), 
        .CO(\CARRYB[22][34] ), .S(\SUMB[22][34] ) );
  FA_X1 S2_22_35 ( .A(\ab[22][35] ), .B(\CARRYB[21][35] ), .CI(\SUMB[21][36] ), 
        .CO(\CARRYB[22][35] ), .S(\SUMB[22][35] ) );
  FA_X1 S2_22_36 ( .A(\ab[22][36] ), .B(\CARRYB[21][36] ), .CI(\SUMB[21][37] ), 
        .CO(\CARRYB[22][36] ), .S(\SUMB[22][36] ) );
  FA_X1 S2_22_37 ( .A(\ab[22][37] ), .B(\CARRYB[21][37] ), .CI(\SUMB[21][38] ), 
        .CO(\CARRYB[22][37] ), .S(\SUMB[22][37] ) );
  FA_X1 S2_22_38 ( .A(\ab[22][38] ), .B(\CARRYB[21][38] ), .CI(\SUMB[21][39] ), 
        .CO(\CARRYB[22][38] ), .S(\SUMB[22][38] ) );
  FA_X1 S2_22_39 ( .A(\ab[22][39] ), .B(\CARRYB[21][39] ), .CI(\SUMB[21][40] ), 
        .CO(\CARRYB[22][39] ), .S(\SUMB[22][39] ) );
  FA_X1 S2_22_40 ( .A(\ab[22][40] ), .B(\CARRYB[21][40] ), .CI(\SUMB[21][41] ), 
        .CO(\CARRYB[22][40] ), .S(\SUMB[22][40] ) );
  FA_X1 S2_22_41 ( .A(\ab[22][41] ), .B(\CARRYB[21][41] ), .CI(\SUMB[21][42] ), 
        .CO(\CARRYB[22][41] ), .S(\SUMB[22][41] ) );
  FA_X1 S2_22_42 ( .A(\ab[22][42] ), .B(\CARRYB[21][42] ), .CI(\SUMB[21][43] ), 
        .CO(\CARRYB[22][42] ), .S(\SUMB[22][42] ) );
  FA_X1 S2_22_43 ( .A(\ab[22][43] ), .B(\CARRYB[21][43] ), .CI(\SUMB[21][44] ), 
        .CO(\CARRYB[22][43] ), .S(\SUMB[22][43] ) );
  FA_X1 S2_22_44 ( .A(\ab[22][44] ), .B(\CARRYB[21][44] ), .CI(\SUMB[21][45] ), 
        .CO(\CARRYB[22][44] ), .S(\SUMB[22][44] ) );
  FA_X1 S2_22_45 ( .A(\ab[22][45] ), .B(\CARRYB[21][45] ), .CI(\SUMB[21][46] ), 
        .CO(\CARRYB[22][45] ), .S(\SUMB[22][45] ) );
  FA_X1 S2_22_46 ( .A(\ab[22][46] ), .B(\CARRYB[21][46] ), .CI(\SUMB[21][47] ), 
        .CO(\CARRYB[22][46] ), .S(\SUMB[22][46] ) );
  FA_X1 S2_22_47 ( .A(\ab[22][47] ), .B(\CARRYB[21][47] ), .CI(\SUMB[21][48] ), 
        .CO(\CARRYB[22][47] ), .S(\SUMB[22][47] ) );
  FA_X1 S2_22_48 ( .A(\ab[22][48] ), .B(\CARRYB[21][48] ), .CI(\SUMB[21][49] ), 
        .CO(\CARRYB[22][48] ), .S(\SUMB[22][48] ) );
  FA_X1 S2_22_49 ( .A(\ab[22][49] ), .B(\CARRYB[21][49] ), .CI(\SUMB[21][50] ), 
        .CO(\CARRYB[22][49] ), .S(\SUMB[22][49] ) );
  FA_X1 S2_22_50 ( .A(\ab[22][50] ), .B(\CARRYB[21][50] ), .CI(\SUMB[21][51] ), 
        .CO(\CARRYB[22][50] ), .S(\SUMB[22][50] ) );
  FA_X1 S3_22_51 ( .A(\ab[22][51] ), .B(\CARRYB[21][51] ), .CI(\ab[21][52] ), 
        .CO(\CARRYB[22][51] ), .S(\SUMB[22][51] ) );
  FA_X1 S1_21_0 ( .A(\ab[21][0] ), .B(\CARRYB[20][0] ), .CI(\SUMB[20][1] ), 
        .CO(\CARRYB[21][0] ), .S(CLA_SUM[21]) );
  FA_X1 S2_21_1 ( .A(\ab[21][1] ), .B(\CARRYB[20][1] ), .CI(\SUMB[20][2] ), 
        .CO(\CARRYB[21][1] ), .S(\SUMB[21][1] ) );
  FA_X1 S2_21_2 ( .A(\ab[21][2] ), .B(\CARRYB[20][2] ), .CI(\SUMB[20][3] ), 
        .CO(\CARRYB[21][2] ), .S(\SUMB[21][2] ) );
  FA_X1 S2_21_3 ( .A(\ab[21][3] ), .B(\CARRYB[20][3] ), .CI(\SUMB[20][4] ), 
        .CO(\CARRYB[21][3] ), .S(\SUMB[21][3] ) );
  FA_X1 S2_21_4 ( .A(\ab[21][4] ), .B(\CARRYB[20][4] ), .CI(\SUMB[20][5] ), 
        .CO(\CARRYB[21][4] ), .S(\SUMB[21][4] ) );
  FA_X1 S2_21_5 ( .A(\ab[21][5] ), .B(\CARRYB[20][5] ), .CI(\SUMB[20][6] ), 
        .CO(\CARRYB[21][5] ), .S(\SUMB[21][5] ) );
  FA_X1 S2_21_6 ( .A(\ab[21][6] ), .B(\CARRYB[20][6] ), .CI(\SUMB[20][7] ), 
        .CO(\CARRYB[21][6] ), .S(\SUMB[21][6] ) );
  FA_X1 S2_21_7 ( .A(\ab[21][7] ), .B(\CARRYB[20][7] ), .CI(\SUMB[20][8] ), 
        .CO(\CARRYB[21][7] ), .S(\SUMB[21][7] ) );
  FA_X1 S2_21_8 ( .A(\ab[21][8] ), .B(\CARRYB[20][8] ), .CI(\SUMB[20][9] ), 
        .CO(\CARRYB[21][8] ), .S(\SUMB[21][8] ) );
  FA_X1 S2_21_9 ( .A(\ab[21][9] ), .B(\CARRYB[20][9] ), .CI(\SUMB[20][10] ), 
        .CO(\CARRYB[21][9] ), .S(\SUMB[21][9] ) );
  FA_X1 S2_21_10 ( .A(\ab[21][10] ), .B(\CARRYB[20][10] ), .CI(\SUMB[20][11] ), 
        .CO(\CARRYB[21][10] ), .S(\SUMB[21][10] ) );
  FA_X1 S2_21_11 ( .A(\ab[21][11] ), .B(\CARRYB[20][11] ), .CI(\SUMB[20][12] ), 
        .CO(\CARRYB[21][11] ), .S(\SUMB[21][11] ) );
  FA_X1 S2_21_12 ( .A(\ab[21][12] ), .B(\CARRYB[20][12] ), .CI(\SUMB[20][13] ), 
        .CO(\CARRYB[21][12] ), .S(\SUMB[21][12] ) );
  FA_X1 S2_21_13 ( .A(\ab[21][13] ), .B(\CARRYB[20][13] ), .CI(\SUMB[20][14] ), 
        .CO(\CARRYB[21][13] ), .S(\SUMB[21][13] ) );
  FA_X1 S2_21_14 ( .A(\ab[21][14] ), .B(\CARRYB[20][14] ), .CI(\SUMB[20][15] ), 
        .CO(\CARRYB[21][14] ), .S(\SUMB[21][14] ) );
  FA_X1 S2_21_15 ( .A(\ab[21][15] ), .B(\CARRYB[20][15] ), .CI(\SUMB[20][16] ), 
        .CO(\CARRYB[21][15] ), .S(\SUMB[21][15] ) );
  FA_X1 S2_21_16 ( .A(\ab[21][16] ), .B(\CARRYB[20][16] ), .CI(\SUMB[20][17] ), 
        .CO(\CARRYB[21][16] ), .S(\SUMB[21][16] ) );
  FA_X1 S2_21_17 ( .A(\ab[21][17] ), .B(\CARRYB[20][17] ), .CI(\SUMB[20][18] ), 
        .CO(\CARRYB[21][17] ), .S(\SUMB[21][17] ) );
  FA_X1 S2_21_18 ( .A(\ab[21][18] ), .B(\CARRYB[20][18] ), .CI(\SUMB[20][19] ), 
        .CO(\CARRYB[21][18] ), .S(\SUMB[21][18] ) );
  FA_X1 S2_21_19 ( .A(\ab[21][19] ), .B(\CARRYB[20][19] ), .CI(\SUMB[20][20] ), 
        .CO(\CARRYB[21][19] ), .S(\SUMB[21][19] ) );
  FA_X1 S2_21_20 ( .A(\ab[21][20] ), .B(\CARRYB[20][20] ), .CI(\SUMB[20][21] ), 
        .CO(\CARRYB[21][20] ), .S(\SUMB[21][20] ) );
  FA_X1 S2_21_21 ( .A(\ab[21][21] ), .B(\CARRYB[20][21] ), .CI(\SUMB[20][22] ), 
        .CO(\CARRYB[21][21] ), .S(\SUMB[21][21] ) );
  FA_X1 S2_21_22 ( .A(\ab[21][22] ), .B(\CARRYB[20][22] ), .CI(\SUMB[20][23] ), 
        .CO(\CARRYB[21][22] ), .S(\SUMB[21][22] ) );
  FA_X1 S2_21_23 ( .A(\ab[21][23] ), .B(\CARRYB[20][23] ), .CI(\SUMB[20][24] ), 
        .CO(\CARRYB[21][23] ), .S(\SUMB[21][23] ) );
  FA_X1 S2_21_24 ( .A(\ab[21][24] ), .B(\CARRYB[20][24] ), .CI(\SUMB[20][25] ), 
        .CO(\CARRYB[21][24] ), .S(\SUMB[21][24] ) );
  FA_X1 S2_21_25 ( .A(\ab[21][25] ), .B(\CARRYB[20][25] ), .CI(\SUMB[20][26] ), 
        .CO(\CARRYB[21][25] ), .S(\SUMB[21][25] ) );
  FA_X1 S2_21_26 ( .A(\ab[21][26] ), .B(\CARRYB[20][26] ), .CI(\SUMB[20][27] ), 
        .CO(\CARRYB[21][26] ), .S(\SUMB[21][26] ) );
  FA_X1 S2_21_27 ( .A(\ab[21][27] ), .B(\CARRYB[20][27] ), .CI(\SUMB[20][28] ), 
        .CO(\CARRYB[21][27] ), .S(\SUMB[21][27] ) );
  FA_X1 S2_21_28 ( .A(\ab[21][28] ), .B(\CARRYB[20][28] ), .CI(\SUMB[20][29] ), 
        .CO(\CARRYB[21][28] ), .S(\SUMB[21][28] ) );
  FA_X1 S2_21_29 ( .A(\ab[21][29] ), .B(\CARRYB[20][29] ), .CI(\SUMB[20][30] ), 
        .CO(\CARRYB[21][29] ), .S(\SUMB[21][29] ) );
  FA_X1 S2_21_30 ( .A(\ab[21][30] ), .B(\CARRYB[20][30] ), .CI(\SUMB[20][31] ), 
        .CO(\CARRYB[21][30] ), .S(\SUMB[21][30] ) );
  FA_X1 S2_21_31 ( .A(\ab[21][31] ), .B(\CARRYB[20][31] ), .CI(\SUMB[20][32] ), 
        .CO(\CARRYB[21][31] ), .S(\SUMB[21][31] ) );
  FA_X1 S2_21_32 ( .A(\ab[21][32] ), .B(\CARRYB[20][32] ), .CI(\SUMB[20][33] ), 
        .CO(\CARRYB[21][32] ), .S(\SUMB[21][32] ) );
  FA_X1 S2_21_33 ( .A(\ab[21][33] ), .B(\CARRYB[20][33] ), .CI(\SUMB[20][34] ), 
        .CO(\CARRYB[21][33] ), .S(\SUMB[21][33] ) );
  FA_X1 S2_21_34 ( .A(\ab[21][34] ), .B(\CARRYB[20][34] ), .CI(\SUMB[20][35] ), 
        .CO(\CARRYB[21][34] ), .S(\SUMB[21][34] ) );
  FA_X1 S2_21_35 ( .A(\ab[21][35] ), .B(\CARRYB[20][35] ), .CI(\SUMB[20][36] ), 
        .CO(\CARRYB[21][35] ), .S(\SUMB[21][35] ) );
  FA_X1 S2_21_36 ( .A(\ab[21][36] ), .B(\CARRYB[20][36] ), .CI(\SUMB[20][37] ), 
        .CO(\CARRYB[21][36] ), .S(\SUMB[21][36] ) );
  FA_X1 S2_21_37 ( .A(\ab[21][37] ), .B(\CARRYB[20][37] ), .CI(\SUMB[20][38] ), 
        .CO(\CARRYB[21][37] ), .S(\SUMB[21][37] ) );
  FA_X1 S2_21_38 ( .A(\ab[21][38] ), .B(\CARRYB[20][38] ), .CI(\SUMB[20][39] ), 
        .CO(\CARRYB[21][38] ), .S(\SUMB[21][38] ) );
  FA_X1 S2_21_39 ( .A(\ab[21][39] ), .B(\CARRYB[20][39] ), .CI(\SUMB[20][40] ), 
        .CO(\CARRYB[21][39] ), .S(\SUMB[21][39] ) );
  FA_X1 S2_21_40 ( .A(\ab[21][40] ), .B(\CARRYB[20][40] ), .CI(\SUMB[20][41] ), 
        .CO(\CARRYB[21][40] ), .S(\SUMB[21][40] ) );
  FA_X1 S2_21_41 ( .A(\ab[21][41] ), .B(\CARRYB[20][41] ), .CI(\SUMB[20][42] ), 
        .CO(\CARRYB[21][41] ), .S(\SUMB[21][41] ) );
  FA_X1 S2_21_42 ( .A(\ab[21][42] ), .B(\CARRYB[20][42] ), .CI(\SUMB[20][43] ), 
        .CO(\CARRYB[21][42] ), .S(\SUMB[21][42] ) );
  FA_X1 S2_21_43 ( .A(\ab[21][43] ), .B(\CARRYB[20][43] ), .CI(\SUMB[20][44] ), 
        .CO(\CARRYB[21][43] ), .S(\SUMB[21][43] ) );
  FA_X1 S2_21_44 ( .A(\ab[21][44] ), .B(\CARRYB[20][44] ), .CI(\SUMB[20][45] ), 
        .CO(\CARRYB[21][44] ), .S(\SUMB[21][44] ) );
  FA_X1 S2_21_45 ( .A(\ab[21][45] ), .B(\CARRYB[20][45] ), .CI(\SUMB[20][46] ), 
        .CO(\CARRYB[21][45] ), .S(\SUMB[21][45] ) );
  FA_X1 S2_21_46 ( .A(\ab[21][46] ), .B(\CARRYB[20][46] ), .CI(\SUMB[20][47] ), 
        .CO(\CARRYB[21][46] ), .S(\SUMB[21][46] ) );
  FA_X1 S2_21_47 ( .A(\ab[21][47] ), .B(\CARRYB[20][47] ), .CI(\SUMB[20][48] ), 
        .CO(\CARRYB[21][47] ), .S(\SUMB[21][47] ) );
  FA_X1 S2_21_48 ( .A(\ab[21][48] ), .B(\CARRYB[20][48] ), .CI(\SUMB[20][49] ), 
        .CO(\CARRYB[21][48] ), .S(\SUMB[21][48] ) );
  FA_X1 S2_21_49 ( .A(\ab[21][49] ), .B(\CARRYB[20][49] ), .CI(\SUMB[20][50] ), 
        .CO(\CARRYB[21][49] ), .S(\SUMB[21][49] ) );
  FA_X1 S2_21_50 ( .A(\ab[21][50] ), .B(\CARRYB[20][50] ), .CI(\SUMB[20][51] ), 
        .CO(\CARRYB[21][50] ), .S(\SUMB[21][50] ) );
  FA_X1 S3_21_51 ( .A(\ab[21][51] ), .B(\CARRYB[20][51] ), .CI(\ab[20][52] ), 
        .CO(\CARRYB[21][51] ), .S(\SUMB[21][51] ) );
  FA_X1 S1_20_0 ( .A(\ab[20][0] ), .B(\CARRYB[19][0] ), .CI(\SUMB[19][1] ), 
        .CO(\CARRYB[20][0] ), .S(CLA_SUM[20]) );
  FA_X1 S2_20_1 ( .A(\ab[20][1] ), .B(\CARRYB[19][1] ), .CI(\SUMB[19][2] ), 
        .CO(\CARRYB[20][1] ), .S(\SUMB[20][1] ) );
  FA_X1 S2_20_2 ( .A(\ab[20][2] ), .B(\CARRYB[19][2] ), .CI(\SUMB[19][3] ), 
        .CO(\CARRYB[20][2] ), .S(\SUMB[20][2] ) );
  FA_X1 S2_20_3 ( .A(\ab[20][3] ), .B(\CARRYB[19][3] ), .CI(\SUMB[19][4] ), 
        .CO(\CARRYB[20][3] ), .S(\SUMB[20][3] ) );
  FA_X1 S2_20_4 ( .A(\ab[20][4] ), .B(\CARRYB[19][4] ), .CI(\SUMB[19][5] ), 
        .CO(\CARRYB[20][4] ), .S(\SUMB[20][4] ) );
  FA_X1 S2_20_5 ( .A(\ab[20][5] ), .B(\CARRYB[19][5] ), .CI(\SUMB[19][6] ), 
        .CO(\CARRYB[20][5] ), .S(\SUMB[20][5] ) );
  FA_X1 S2_20_6 ( .A(\ab[20][6] ), .B(\CARRYB[19][6] ), .CI(\SUMB[19][7] ), 
        .CO(\CARRYB[20][6] ), .S(\SUMB[20][6] ) );
  FA_X1 S2_20_7 ( .A(\ab[20][7] ), .B(\CARRYB[19][7] ), .CI(\SUMB[19][8] ), 
        .CO(\CARRYB[20][7] ), .S(\SUMB[20][7] ) );
  FA_X1 S2_20_8 ( .A(\ab[20][8] ), .B(\CARRYB[19][8] ), .CI(\SUMB[19][9] ), 
        .CO(\CARRYB[20][8] ), .S(\SUMB[20][8] ) );
  FA_X1 S2_20_9 ( .A(\ab[20][9] ), .B(\CARRYB[19][9] ), .CI(\SUMB[19][10] ), 
        .CO(\CARRYB[20][9] ), .S(\SUMB[20][9] ) );
  FA_X1 S2_20_10 ( .A(\ab[20][10] ), .B(\CARRYB[19][10] ), .CI(\SUMB[19][11] ), 
        .CO(\CARRYB[20][10] ), .S(\SUMB[20][10] ) );
  FA_X1 S2_20_11 ( .A(\ab[20][11] ), .B(\CARRYB[19][11] ), .CI(\SUMB[19][12] ), 
        .CO(\CARRYB[20][11] ), .S(\SUMB[20][11] ) );
  FA_X1 S2_20_12 ( .A(\ab[20][12] ), .B(\CARRYB[19][12] ), .CI(\SUMB[19][13] ), 
        .CO(\CARRYB[20][12] ), .S(\SUMB[20][12] ) );
  FA_X1 S2_20_13 ( .A(\ab[20][13] ), .B(\CARRYB[19][13] ), .CI(\SUMB[19][14] ), 
        .CO(\CARRYB[20][13] ), .S(\SUMB[20][13] ) );
  FA_X1 S2_20_14 ( .A(\ab[20][14] ), .B(\CARRYB[19][14] ), .CI(\SUMB[19][15] ), 
        .CO(\CARRYB[20][14] ), .S(\SUMB[20][14] ) );
  FA_X1 S2_20_15 ( .A(\ab[20][15] ), .B(\CARRYB[19][15] ), .CI(\SUMB[19][16] ), 
        .CO(\CARRYB[20][15] ), .S(\SUMB[20][15] ) );
  FA_X1 S2_20_16 ( .A(\ab[20][16] ), .B(\CARRYB[19][16] ), .CI(\SUMB[19][17] ), 
        .CO(\CARRYB[20][16] ), .S(\SUMB[20][16] ) );
  FA_X1 S2_20_17 ( .A(\ab[20][17] ), .B(\CARRYB[19][17] ), .CI(\SUMB[19][18] ), 
        .CO(\CARRYB[20][17] ), .S(\SUMB[20][17] ) );
  FA_X1 S2_20_18 ( .A(\ab[20][18] ), .B(\CARRYB[19][18] ), .CI(\SUMB[19][19] ), 
        .CO(\CARRYB[20][18] ), .S(\SUMB[20][18] ) );
  FA_X1 S2_20_19 ( .A(\ab[20][19] ), .B(\CARRYB[19][19] ), .CI(\SUMB[19][20] ), 
        .CO(\CARRYB[20][19] ), .S(\SUMB[20][19] ) );
  FA_X1 S2_20_20 ( .A(\ab[20][20] ), .B(\CARRYB[19][20] ), .CI(\SUMB[19][21] ), 
        .CO(\CARRYB[20][20] ), .S(\SUMB[20][20] ) );
  FA_X1 S2_20_21 ( .A(\ab[20][21] ), .B(\CARRYB[19][21] ), .CI(\SUMB[19][22] ), 
        .CO(\CARRYB[20][21] ), .S(\SUMB[20][21] ) );
  FA_X1 S2_20_22 ( .A(\ab[20][22] ), .B(\CARRYB[19][22] ), .CI(\SUMB[19][23] ), 
        .CO(\CARRYB[20][22] ), .S(\SUMB[20][22] ) );
  FA_X1 S2_20_23 ( .A(\ab[20][23] ), .B(\CARRYB[19][23] ), .CI(\SUMB[19][24] ), 
        .CO(\CARRYB[20][23] ), .S(\SUMB[20][23] ) );
  FA_X1 S2_20_24 ( .A(\ab[20][24] ), .B(\CARRYB[19][24] ), .CI(\SUMB[19][25] ), 
        .CO(\CARRYB[20][24] ), .S(\SUMB[20][24] ) );
  FA_X1 S2_20_25 ( .A(\ab[20][25] ), .B(\CARRYB[19][25] ), .CI(\SUMB[19][26] ), 
        .CO(\CARRYB[20][25] ), .S(\SUMB[20][25] ) );
  FA_X1 S2_20_26 ( .A(\ab[20][26] ), .B(\CARRYB[19][26] ), .CI(\SUMB[19][27] ), 
        .CO(\CARRYB[20][26] ), .S(\SUMB[20][26] ) );
  FA_X1 S2_20_27 ( .A(\ab[20][27] ), .B(\CARRYB[19][27] ), .CI(\SUMB[19][28] ), 
        .CO(\CARRYB[20][27] ), .S(\SUMB[20][27] ) );
  FA_X1 S2_20_28 ( .A(\ab[20][28] ), .B(\CARRYB[19][28] ), .CI(\SUMB[19][29] ), 
        .CO(\CARRYB[20][28] ), .S(\SUMB[20][28] ) );
  FA_X1 S2_20_29 ( .A(\ab[20][29] ), .B(\CARRYB[19][29] ), .CI(\SUMB[19][30] ), 
        .CO(\CARRYB[20][29] ), .S(\SUMB[20][29] ) );
  FA_X1 S2_20_30 ( .A(\ab[20][30] ), .B(\CARRYB[19][30] ), .CI(\SUMB[19][31] ), 
        .CO(\CARRYB[20][30] ), .S(\SUMB[20][30] ) );
  FA_X1 S2_20_31 ( .A(\ab[20][31] ), .B(\CARRYB[19][31] ), .CI(\SUMB[19][32] ), 
        .CO(\CARRYB[20][31] ), .S(\SUMB[20][31] ) );
  FA_X1 S2_20_32 ( .A(\ab[20][32] ), .B(\CARRYB[19][32] ), .CI(\SUMB[19][33] ), 
        .CO(\CARRYB[20][32] ), .S(\SUMB[20][32] ) );
  FA_X1 S2_20_33 ( .A(\ab[20][33] ), .B(\CARRYB[19][33] ), .CI(\SUMB[19][34] ), 
        .CO(\CARRYB[20][33] ), .S(\SUMB[20][33] ) );
  FA_X1 S2_20_34 ( .A(\ab[20][34] ), .B(\CARRYB[19][34] ), .CI(\SUMB[19][35] ), 
        .CO(\CARRYB[20][34] ), .S(\SUMB[20][34] ) );
  FA_X1 S2_20_35 ( .A(\ab[20][35] ), .B(\CARRYB[19][35] ), .CI(\SUMB[19][36] ), 
        .CO(\CARRYB[20][35] ), .S(\SUMB[20][35] ) );
  FA_X1 S2_20_36 ( .A(\ab[20][36] ), .B(\CARRYB[19][36] ), .CI(\SUMB[19][37] ), 
        .CO(\CARRYB[20][36] ), .S(\SUMB[20][36] ) );
  FA_X1 S2_20_37 ( .A(\ab[20][37] ), .B(\CARRYB[19][37] ), .CI(\SUMB[19][38] ), 
        .CO(\CARRYB[20][37] ), .S(\SUMB[20][37] ) );
  FA_X1 S2_20_38 ( .A(\ab[20][38] ), .B(\CARRYB[19][38] ), .CI(\SUMB[19][39] ), 
        .CO(\CARRYB[20][38] ), .S(\SUMB[20][38] ) );
  FA_X1 S2_20_39 ( .A(\ab[20][39] ), .B(\CARRYB[19][39] ), .CI(\SUMB[19][40] ), 
        .CO(\CARRYB[20][39] ), .S(\SUMB[20][39] ) );
  FA_X1 S2_20_40 ( .A(\ab[20][40] ), .B(\CARRYB[19][40] ), .CI(\SUMB[19][41] ), 
        .CO(\CARRYB[20][40] ), .S(\SUMB[20][40] ) );
  FA_X1 S2_20_41 ( .A(\ab[20][41] ), .B(\CARRYB[19][41] ), .CI(\SUMB[19][42] ), 
        .CO(\CARRYB[20][41] ), .S(\SUMB[20][41] ) );
  FA_X1 S2_20_42 ( .A(\ab[20][42] ), .B(\CARRYB[19][42] ), .CI(\SUMB[19][43] ), 
        .CO(\CARRYB[20][42] ), .S(\SUMB[20][42] ) );
  FA_X1 S2_20_43 ( .A(\ab[20][43] ), .B(\CARRYB[19][43] ), .CI(\SUMB[19][44] ), 
        .CO(\CARRYB[20][43] ), .S(\SUMB[20][43] ) );
  FA_X1 S2_20_44 ( .A(\ab[20][44] ), .B(\CARRYB[19][44] ), .CI(\SUMB[19][45] ), 
        .CO(\CARRYB[20][44] ), .S(\SUMB[20][44] ) );
  FA_X1 S2_20_45 ( .A(\ab[20][45] ), .B(\CARRYB[19][45] ), .CI(\SUMB[19][46] ), 
        .CO(\CARRYB[20][45] ), .S(\SUMB[20][45] ) );
  FA_X1 S2_20_46 ( .A(\ab[20][46] ), .B(\CARRYB[19][46] ), .CI(\SUMB[19][47] ), 
        .CO(\CARRYB[20][46] ), .S(\SUMB[20][46] ) );
  FA_X1 S2_20_47 ( .A(\ab[20][47] ), .B(\CARRYB[19][47] ), .CI(\SUMB[19][48] ), 
        .CO(\CARRYB[20][47] ), .S(\SUMB[20][47] ) );
  FA_X1 S2_20_48 ( .A(\ab[20][48] ), .B(\CARRYB[19][48] ), .CI(\SUMB[19][49] ), 
        .CO(\CARRYB[20][48] ), .S(\SUMB[20][48] ) );
  FA_X1 S2_20_49 ( .A(\ab[20][49] ), .B(\CARRYB[19][49] ), .CI(\SUMB[19][50] ), 
        .CO(\CARRYB[20][49] ), .S(\SUMB[20][49] ) );
  FA_X1 S2_20_50 ( .A(\ab[20][50] ), .B(\CARRYB[19][50] ), .CI(\SUMB[19][51] ), 
        .CO(\CARRYB[20][50] ), .S(\SUMB[20][50] ) );
  FA_X1 S3_20_51 ( .A(\ab[20][51] ), .B(\CARRYB[19][51] ), .CI(\ab[19][52] ), 
        .CO(\CARRYB[20][51] ), .S(\SUMB[20][51] ) );
  FA_X1 S1_19_0 ( .A(\ab[19][0] ), .B(\CARRYB[18][0] ), .CI(\SUMB[18][1] ), 
        .CO(\CARRYB[19][0] ), .S(CLA_SUM[19]) );
  FA_X1 S2_19_1 ( .A(\ab[19][1] ), .B(\CARRYB[18][1] ), .CI(\SUMB[18][2] ), 
        .CO(\CARRYB[19][1] ), .S(\SUMB[19][1] ) );
  FA_X1 S2_19_2 ( .A(\ab[19][2] ), .B(\CARRYB[18][2] ), .CI(\SUMB[18][3] ), 
        .CO(\CARRYB[19][2] ), .S(\SUMB[19][2] ) );
  FA_X1 S2_19_3 ( .A(\ab[19][3] ), .B(\CARRYB[18][3] ), .CI(\SUMB[18][4] ), 
        .CO(\CARRYB[19][3] ), .S(\SUMB[19][3] ) );
  FA_X1 S2_19_4 ( .A(\ab[19][4] ), .B(\CARRYB[18][4] ), .CI(\SUMB[18][5] ), 
        .CO(\CARRYB[19][4] ), .S(\SUMB[19][4] ) );
  FA_X1 S2_19_5 ( .A(\ab[19][5] ), .B(\CARRYB[18][5] ), .CI(\SUMB[18][6] ), 
        .CO(\CARRYB[19][5] ), .S(\SUMB[19][5] ) );
  FA_X1 S2_19_6 ( .A(\ab[19][6] ), .B(\CARRYB[18][6] ), .CI(\SUMB[18][7] ), 
        .CO(\CARRYB[19][6] ), .S(\SUMB[19][6] ) );
  FA_X1 S2_19_7 ( .A(\ab[19][7] ), .B(\CARRYB[18][7] ), .CI(\SUMB[18][8] ), 
        .CO(\CARRYB[19][7] ), .S(\SUMB[19][7] ) );
  FA_X1 S2_19_8 ( .A(\ab[19][8] ), .B(\CARRYB[18][8] ), .CI(\SUMB[18][9] ), 
        .CO(\CARRYB[19][8] ), .S(\SUMB[19][8] ) );
  FA_X1 S2_19_9 ( .A(\ab[19][9] ), .B(\CARRYB[18][9] ), .CI(\SUMB[18][10] ), 
        .CO(\CARRYB[19][9] ), .S(\SUMB[19][9] ) );
  FA_X1 S2_19_10 ( .A(\ab[19][10] ), .B(\CARRYB[18][10] ), .CI(\SUMB[18][11] ), 
        .CO(\CARRYB[19][10] ), .S(\SUMB[19][10] ) );
  FA_X1 S2_19_11 ( .A(\ab[19][11] ), .B(\CARRYB[18][11] ), .CI(\SUMB[18][12] ), 
        .CO(\CARRYB[19][11] ), .S(\SUMB[19][11] ) );
  FA_X1 S2_19_12 ( .A(\ab[19][12] ), .B(\CARRYB[18][12] ), .CI(\SUMB[18][13] ), 
        .CO(\CARRYB[19][12] ), .S(\SUMB[19][12] ) );
  FA_X1 S2_19_13 ( .A(\ab[19][13] ), .B(\CARRYB[18][13] ), .CI(\SUMB[18][14] ), 
        .CO(\CARRYB[19][13] ), .S(\SUMB[19][13] ) );
  FA_X1 S2_19_14 ( .A(\ab[19][14] ), .B(\CARRYB[18][14] ), .CI(\SUMB[18][15] ), 
        .CO(\CARRYB[19][14] ), .S(\SUMB[19][14] ) );
  FA_X1 S2_19_15 ( .A(\ab[19][15] ), .B(\CARRYB[18][15] ), .CI(\SUMB[18][16] ), 
        .CO(\CARRYB[19][15] ), .S(\SUMB[19][15] ) );
  FA_X1 S2_19_16 ( .A(\ab[19][16] ), .B(\CARRYB[18][16] ), .CI(\SUMB[18][17] ), 
        .CO(\CARRYB[19][16] ), .S(\SUMB[19][16] ) );
  FA_X1 S2_19_17 ( .A(\ab[19][17] ), .B(\CARRYB[18][17] ), .CI(\SUMB[18][18] ), 
        .CO(\CARRYB[19][17] ), .S(\SUMB[19][17] ) );
  FA_X1 S2_19_18 ( .A(\ab[19][18] ), .B(\CARRYB[18][18] ), .CI(\SUMB[18][19] ), 
        .CO(\CARRYB[19][18] ), .S(\SUMB[19][18] ) );
  FA_X1 S2_19_19 ( .A(\ab[19][19] ), .B(\CARRYB[18][19] ), .CI(\SUMB[18][20] ), 
        .CO(\CARRYB[19][19] ), .S(\SUMB[19][19] ) );
  FA_X1 S2_19_20 ( .A(\ab[19][20] ), .B(\CARRYB[18][20] ), .CI(\SUMB[18][21] ), 
        .CO(\CARRYB[19][20] ), .S(\SUMB[19][20] ) );
  FA_X1 S2_19_21 ( .A(\ab[19][21] ), .B(\CARRYB[18][21] ), .CI(\SUMB[18][22] ), 
        .CO(\CARRYB[19][21] ), .S(\SUMB[19][21] ) );
  FA_X1 S2_19_22 ( .A(\ab[19][22] ), .B(\CARRYB[18][22] ), .CI(\SUMB[18][23] ), 
        .CO(\CARRYB[19][22] ), .S(\SUMB[19][22] ) );
  FA_X1 S2_19_23 ( .A(\ab[19][23] ), .B(\CARRYB[18][23] ), .CI(\SUMB[18][24] ), 
        .CO(\CARRYB[19][23] ), .S(\SUMB[19][23] ) );
  FA_X1 S2_19_24 ( .A(\ab[19][24] ), .B(\CARRYB[18][24] ), .CI(\SUMB[18][25] ), 
        .CO(\CARRYB[19][24] ), .S(\SUMB[19][24] ) );
  FA_X1 S2_19_25 ( .A(\ab[19][25] ), .B(\CARRYB[18][25] ), .CI(\SUMB[18][26] ), 
        .CO(\CARRYB[19][25] ), .S(\SUMB[19][25] ) );
  FA_X1 S2_19_26 ( .A(\ab[19][26] ), .B(\CARRYB[18][26] ), .CI(\SUMB[18][27] ), 
        .CO(\CARRYB[19][26] ), .S(\SUMB[19][26] ) );
  FA_X1 S2_19_27 ( .A(\ab[19][27] ), .B(\CARRYB[18][27] ), .CI(\SUMB[18][28] ), 
        .CO(\CARRYB[19][27] ), .S(\SUMB[19][27] ) );
  FA_X1 S2_19_28 ( .A(\ab[19][28] ), .B(\CARRYB[18][28] ), .CI(\SUMB[18][29] ), 
        .CO(\CARRYB[19][28] ), .S(\SUMB[19][28] ) );
  FA_X1 S2_19_29 ( .A(\ab[19][29] ), .B(\CARRYB[18][29] ), .CI(\SUMB[18][30] ), 
        .CO(\CARRYB[19][29] ), .S(\SUMB[19][29] ) );
  FA_X1 S2_19_30 ( .A(\ab[19][30] ), .B(\CARRYB[18][30] ), .CI(\SUMB[18][31] ), 
        .CO(\CARRYB[19][30] ), .S(\SUMB[19][30] ) );
  FA_X1 S2_19_31 ( .A(\ab[19][31] ), .B(\CARRYB[18][31] ), .CI(\SUMB[18][32] ), 
        .CO(\CARRYB[19][31] ), .S(\SUMB[19][31] ) );
  FA_X1 S2_19_32 ( .A(\ab[19][32] ), .B(\CARRYB[18][32] ), .CI(\SUMB[18][33] ), 
        .CO(\CARRYB[19][32] ), .S(\SUMB[19][32] ) );
  FA_X1 S2_19_33 ( .A(\ab[19][33] ), .B(\CARRYB[18][33] ), .CI(\SUMB[18][34] ), 
        .CO(\CARRYB[19][33] ), .S(\SUMB[19][33] ) );
  FA_X1 S2_19_34 ( .A(\ab[19][34] ), .B(\CARRYB[18][34] ), .CI(\SUMB[18][35] ), 
        .CO(\CARRYB[19][34] ), .S(\SUMB[19][34] ) );
  FA_X1 S2_19_35 ( .A(\ab[19][35] ), .B(\CARRYB[18][35] ), .CI(\SUMB[18][36] ), 
        .CO(\CARRYB[19][35] ), .S(\SUMB[19][35] ) );
  FA_X1 S2_19_36 ( .A(\ab[19][36] ), .B(\CARRYB[18][36] ), .CI(\SUMB[18][37] ), 
        .CO(\CARRYB[19][36] ), .S(\SUMB[19][36] ) );
  FA_X1 S2_19_37 ( .A(\ab[19][37] ), .B(\CARRYB[18][37] ), .CI(\SUMB[18][38] ), 
        .CO(\CARRYB[19][37] ), .S(\SUMB[19][37] ) );
  FA_X1 S2_19_38 ( .A(\ab[19][38] ), .B(\CARRYB[18][38] ), .CI(\SUMB[18][39] ), 
        .CO(\CARRYB[19][38] ), .S(\SUMB[19][38] ) );
  FA_X1 S2_19_39 ( .A(\ab[19][39] ), .B(\CARRYB[18][39] ), .CI(\SUMB[18][40] ), 
        .CO(\CARRYB[19][39] ), .S(\SUMB[19][39] ) );
  FA_X1 S2_19_40 ( .A(\ab[19][40] ), .B(\CARRYB[18][40] ), .CI(\SUMB[18][41] ), 
        .CO(\CARRYB[19][40] ), .S(\SUMB[19][40] ) );
  FA_X1 S2_19_41 ( .A(\ab[19][41] ), .B(\CARRYB[18][41] ), .CI(\SUMB[18][42] ), 
        .CO(\CARRYB[19][41] ), .S(\SUMB[19][41] ) );
  FA_X1 S2_19_42 ( .A(\ab[19][42] ), .B(\CARRYB[18][42] ), .CI(\SUMB[18][43] ), 
        .CO(\CARRYB[19][42] ), .S(\SUMB[19][42] ) );
  FA_X1 S2_19_43 ( .A(\ab[19][43] ), .B(\CARRYB[18][43] ), .CI(\SUMB[18][44] ), 
        .CO(\CARRYB[19][43] ), .S(\SUMB[19][43] ) );
  FA_X1 S2_19_44 ( .A(\ab[19][44] ), .B(\CARRYB[18][44] ), .CI(\SUMB[18][45] ), 
        .CO(\CARRYB[19][44] ), .S(\SUMB[19][44] ) );
  FA_X1 S2_19_45 ( .A(\ab[19][45] ), .B(\CARRYB[18][45] ), .CI(\SUMB[18][46] ), 
        .CO(\CARRYB[19][45] ), .S(\SUMB[19][45] ) );
  FA_X1 S2_19_46 ( .A(\ab[19][46] ), .B(\CARRYB[18][46] ), .CI(\SUMB[18][47] ), 
        .CO(\CARRYB[19][46] ), .S(\SUMB[19][46] ) );
  FA_X1 S2_19_47 ( .A(\ab[19][47] ), .B(\CARRYB[18][47] ), .CI(\SUMB[18][48] ), 
        .CO(\CARRYB[19][47] ), .S(\SUMB[19][47] ) );
  FA_X1 S2_19_48 ( .A(\ab[19][48] ), .B(\CARRYB[18][48] ), .CI(\SUMB[18][49] ), 
        .CO(\CARRYB[19][48] ), .S(\SUMB[19][48] ) );
  FA_X1 S2_19_49 ( .A(\ab[19][49] ), .B(\CARRYB[18][49] ), .CI(\SUMB[18][50] ), 
        .CO(\CARRYB[19][49] ), .S(\SUMB[19][49] ) );
  FA_X1 S2_19_50 ( .A(\ab[19][50] ), .B(\CARRYB[18][50] ), .CI(\SUMB[18][51] ), 
        .CO(\CARRYB[19][50] ), .S(\SUMB[19][50] ) );
  FA_X1 S3_19_51 ( .A(\ab[19][51] ), .B(\CARRYB[18][51] ), .CI(\ab[18][52] ), 
        .CO(\CARRYB[19][51] ), .S(\SUMB[19][51] ) );
  FA_X1 S1_18_0 ( .A(\ab[18][0] ), .B(\CARRYB[17][0] ), .CI(\SUMB[17][1] ), 
        .CO(\CARRYB[18][0] ), .S(CLA_SUM[18]) );
  FA_X1 S2_18_1 ( .A(\ab[18][1] ), .B(\CARRYB[17][1] ), .CI(\SUMB[17][2] ), 
        .CO(\CARRYB[18][1] ), .S(\SUMB[18][1] ) );
  FA_X1 S2_18_2 ( .A(\ab[18][2] ), .B(\CARRYB[17][2] ), .CI(\SUMB[17][3] ), 
        .CO(\CARRYB[18][2] ), .S(\SUMB[18][2] ) );
  FA_X1 S2_18_3 ( .A(\ab[18][3] ), .B(\CARRYB[17][3] ), .CI(\SUMB[17][4] ), 
        .CO(\CARRYB[18][3] ), .S(\SUMB[18][3] ) );
  FA_X1 S2_18_4 ( .A(\ab[18][4] ), .B(\CARRYB[17][4] ), .CI(\SUMB[17][5] ), 
        .CO(\CARRYB[18][4] ), .S(\SUMB[18][4] ) );
  FA_X1 S2_18_5 ( .A(\ab[18][5] ), .B(\CARRYB[17][5] ), .CI(\SUMB[17][6] ), 
        .CO(\CARRYB[18][5] ), .S(\SUMB[18][5] ) );
  FA_X1 S2_18_6 ( .A(\ab[18][6] ), .B(\CARRYB[17][6] ), .CI(\SUMB[17][7] ), 
        .CO(\CARRYB[18][6] ), .S(\SUMB[18][6] ) );
  FA_X1 S2_18_7 ( .A(\ab[18][7] ), .B(\CARRYB[17][7] ), .CI(\SUMB[17][8] ), 
        .CO(\CARRYB[18][7] ), .S(\SUMB[18][7] ) );
  FA_X1 S2_18_8 ( .A(\ab[18][8] ), .B(\CARRYB[17][8] ), .CI(\SUMB[17][9] ), 
        .CO(\CARRYB[18][8] ), .S(\SUMB[18][8] ) );
  FA_X1 S2_18_9 ( .A(\ab[18][9] ), .B(\CARRYB[17][9] ), .CI(\SUMB[17][10] ), 
        .CO(\CARRYB[18][9] ), .S(\SUMB[18][9] ) );
  FA_X1 S2_18_10 ( .A(\ab[18][10] ), .B(\CARRYB[17][10] ), .CI(\SUMB[17][11] ), 
        .CO(\CARRYB[18][10] ), .S(\SUMB[18][10] ) );
  FA_X1 S2_18_11 ( .A(\ab[18][11] ), .B(\CARRYB[17][11] ), .CI(\SUMB[17][12] ), 
        .CO(\CARRYB[18][11] ), .S(\SUMB[18][11] ) );
  FA_X1 S2_18_12 ( .A(\ab[18][12] ), .B(\CARRYB[17][12] ), .CI(\SUMB[17][13] ), 
        .CO(\CARRYB[18][12] ), .S(\SUMB[18][12] ) );
  FA_X1 S2_18_13 ( .A(\ab[18][13] ), .B(\CARRYB[17][13] ), .CI(\SUMB[17][14] ), 
        .CO(\CARRYB[18][13] ), .S(\SUMB[18][13] ) );
  FA_X1 S2_18_14 ( .A(\ab[18][14] ), .B(\CARRYB[17][14] ), .CI(\SUMB[17][15] ), 
        .CO(\CARRYB[18][14] ), .S(\SUMB[18][14] ) );
  FA_X1 S2_18_15 ( .A(\ab[18][15] ), .B(\CARRYB[17][15] ), .CI(\SUMB[17][16] ), 
        .CO(\CARRYB[18][15] ), .S(\SUMB[18][15] ) );
  FA_X1 S2_18_16 ( .A(\ab[18][16] ), .B(\CARRYB[17][16] ), .CI(\SUMB[17][17] ), 
        .CO(\CARRYB[18][16] ), .S(\SUMB[18][16] ) );
  FA_X1 S2_18_17 ( .A(\ab[18][17] ), .B(\CARRYB[17][17] ), .CI(\SUMB[17][18] ), 
        .CO(\CARRYB[18][17] ), .S(\SUMB[18][17] ) );
  FA_X1 S2_18_18 ( .A(\ab[18][18] ), .B(\CARRYB[17][18] ), .CI(\SUMB[17][19] ), 
        .CO(\CARRYB[18][18] ), .S(\SUMB[18][18] ) );
  FA_X1 S2_18_19 ( .A(\ab[18][19] ), .B(\CARRYB[17][19] ), .CI(\SUMB[17][20] ), 
        .CO(\CARRYB[18][19] ), .S(\SUMB[18][19] ) );
  FA_X1 S2_18_20 ( .A(\ab[18][20] ), .B(\CARRYB[17][20] ), .CI(\SUMB[17][21] ), 
        .CO(\CARRYB[18][20] ), .S(\SUMB[18][20] ) );
  FA_X1 S2_18_21 ( .A(\ab[18][21] ), .B(\CARRYB[17][21] ), .CI(\SUMB[17][22] ), 
        .CO(\CARRYB[18][21] ), .S(\SUMB[18][21] ) );
  FA_X1 S2_18_22 ( .A(\ab[18][22] ), .B(\CARRYB[17][22] ), .CI(\SUMB[17][23] ), 
        .CO(\CARRYB[18][22] ), .S(\SUMB[18][22] ) );
  FA_X1 S2_18_23 ( .A(\ab[18][23] ), .B(\CARRYB[17][23] ), .CI(\SUMB[17][24] ), 
        .CO(\CARRYB[18][23] ), .S(\SUMB[18][23] ) );
  FA_X1 S2_18_24 ( .A(\ab[18][24] ), .B(\CARRYB[17][24] ), .CI(\SUMB[17][25] ), 
        .CO(\CARRYB[18][24] ), .S(\SUMB[18][24] ) );
  FA_X1 S2_18_25 ( .A(\ab[18][25] ), .B(\CARRYB[17][25] ), .CI(\SUMB[17][26] ), 
        .CO(\CARRYB[18][25] ), .S(\SUMB[18][25] ) );
  FA_X1 S2_18_26 ( .A(\ab[18][26] ), .B(\CARRYB[17][26] ), .CI(\SUMB[17][27] ), 
        .CO(\CARRYB[18][26] ), .S(\SUMB[18][26] ) );
  FA_X1 S2_18_27 ( .A(\ab[18][27] ), .B(\CARRYB[17][27] ), .CI(\SUMB[17][28] ), 
        .CO(\CARRYB[18][27] ), .S(\SUMB[18][27] ) );
  FA_X1 S2_18_28 ( .A(\ab[18][28] ), .B(\CARRYB[17][28] ), .CI(\SUMB[17][29] ), 
        .CO(\CARRYB[18][28] ), .S(\SUMB[18][28] ) );
  FA_X1 S2_18_29 ( .A(\ab[18][29] ), .B(\CARRYB[17][29] ), .CI(\SUMB[17][30] ), 
        .CO(\CARRYB[18][29] ), .S(\SUMB[18][29] ) );
  FA_X1 S2_18_30 ( .A(\ab[18][30] ), .B(\CARRYB[17][30] ), .CI(\SUMB[17][31] ), 
        .CO(\CARRYB[18][30] ), .S(\SUMB[18][30] ) );
  FA_X1 S2_18_31 ( .A(\ab[18][31] ), .B(\CARRYB[17][31] ), .CI(\SUMB[17][32] ), 
        .CO(\CARRYB[18][31] ), .S(\SUMB[18][31] ) );
  FA_X1 S2_18_32 ( .A(\ab[18][32] ), .B(\CARRYB[17][32] ), .CI(\SUMB[17][33] ), 
        .CO(\CARRYB[18][32] ), .S(\SUMB[18][32] ) );
  FA_X1 S2_18_33 ( .A(\ab[18][33] ), .B(\CARRYB[17][33] ), .CI(\SUMB[17][34] ), 
        .CO(\CARRYB[18][33] ), .S(\SUMB[18][33] ) );
  FA_X1 S2_18_34 ( .A(\ab[18][34] ), .B(\CARRYB[17][34] ), .CI(\SUMB[17][35] ), 
        .CO(\CARRYB[18][34] ), .S(\SUMB[18][34] ) );
  FA_X1 S2_18_35 ( .A(\ab[18][35] ), .B(\CARRYB[17][35] ), .CI(\SUMB[17][36] ), 
        .CO(\CARRYB[18][35] ), .S(\SUMB[18][35] ) );
  FA_X1 S2_18_36 ( .A(\ab[18][36] ), .B(\CARRYB[17][36] ), .CI(\SUMB[17][37] ), 
        .CO(\CARRYB[18][36] ), .S(\SUMB[18][36] ) );
  FA_X1 S2_18_37 ( .A(\ab[18][37] ), .B(\CARRYB[17][37] ), .CI(\SUMB[17][38] ), 
        .CO(\CARRYB[18][37] ), .S(\SUMB[18][37] ) );
  FA_X1 S2_18_38 ( .A(\ab[18][38] ), .B(\CARRYB[17][38] ), .CI(\SUMB[17][39] ), 
        .CO(\CARRYB[18][38] ), .S(\SUMB[18][38] ) );
  FA_X1 S2_18_39 ( .A(\ab[18][39] ), .B(\CARRYB[17][39] ), .CI(\SUMB[17][40] ), 
        .CO(\CARRYB[18][39] ), .S(\SUMB[18][39] ) );
  FA_X1 S2_18_40 ( .A(\ab[18][40] ), .B(\CARRYB[17][40] ), .CI(\SUMB[17][41] ), 
        .CO(\CARRYB[18][40] ), .S(\SUMB[18][40] ) );
  FA_X1 S2_18_41 ( .A(\ab[18][41] ), .B(\CARRYB[17][41] ), .CI(\SUMB[17][42] ), 
        .CO(\CARRYB[18][41] ), .S(\SUMB[18][41] ) );
  FA_X1 S2_18_42 ( .A(\ab[18][42] ), .B(\CARRYB[17][42] ), .CI(\SUMB[17][43] ), 
        .CO(\CARRYB[18][42] ), .S(\SUMB[18][42] ) );
  FA_X1 S2_18_43 ( .A(\ab[18][43] ), .B(\CARRYB[17][43] ), .CI(\SUMB[17][44] ), 
        .CO(\CARRYB[18][43] ), .S(\SUMB[18][43] ) );
  FA_X1 S2_18_44 ( .A(\ab[18][44] ), .B(\CARRYB[17][44] ), .CI(\SUMB[17][45] ), 
        .CO(\CARRYB[18][44] ), .S(\SUMB[18][44] ) );
  FA_X1 S2_18_45 ( .A(\ab[18][45] ), .B(\CARRYB[17][45] ), .CI(\SUMB[17][46] ), 
        .CO(\CARRYB[18][45] ), .S(\SUMB[18][45] ) );
  FA_X1 S2_18_46 ( .A(\ab[18][46] ), .B(\CARRYB[17][46] ), .CI(\SUMB[17][47] ), 
        .CO(\CARRYB[18][46] ), .S(\SUMB[18][46] ) );
  FA_X1 S2_18_47 ( .A(\ab[18][47] ), .B(\CARRYB[17][47] ), .CI(\SUMB[17][48] ), 
        .CO(\CARRYB[18][47] ), .S(\SUMB[18][47] ) );
  FA_X1 S2_18_48 ( .A(\ab[18][48] ), .B(\CARRYB[17][48] ), .CI(\SUMB[17][49] ), 
        .CO(\CARRYB[18][48] ), .S(\SUMB[18][48] ) );
  FA_X1 S2_18_49 ( .A(\ab[18][49] ), .B(\CARRYB[17][49] ), .CI(\SUMB[17][50] ), 
        .CO(\CARRYB[18][49] ), .S(\SUMB[18][49] ) );
  FA_X1 S2_18_50 ( .A(\ab[18][50] ), .B(\CARRYB[17][50] ), .CI(\SUMB[17][51] ), 
        .CO(\CARRYB[18][50] ), .S(\SUMB[18][50] ) );
  FA_X1 S3_18_51 ( .A(\ab[18][51] ), .B(\CARRYB[17][51] ), .CI(\ab[17][52] ), 
        .CO(\CARRYB[18][51] ), .S(\SUMB[18][51] ) );
  FA_X1 S1_17_0 ( .A(\ab[17][0] ), .B(\CARRYB[16][0] ), .CI(\SUMB[16][1] ), 
        .CO(\CARRYB[17][0] ), .S(CLA_SUM[17]) );
  FA_X1 S2_17_1 ( .A(\ab[17][1] ), .B(\CARRYB[16][1] ), .CI(\SUMB[16][2] ), 
        .CO(\CARRYB[17][1] ), .S(\SUMB[17][1] ) );
  FA_X1 S2_17_2 ( .A(\ab[17][2] ), .B(\CARRYB[16][2] ), .CI(\SUMB[16][3] ), 
        .CO(\CARRYB[17][2] ), .S(\SUMB[17][2] ) );
  FA_X1 S2_17_3 ( .A(\ab[17][3] ), .B(\CARRYB[16][3] ), .CI(\SUMB[16][4] ), 
        .CO(\CARRYB[17][3] ), .S(\SUMB[17][3] ) );
  FA_X1 S2_17_4 ( .A(\ab[17][4] ), .B(\CARRYB[16][4] ), .CI(\SUMB[16][5] ), 
        .CO(\CARRYB[17][4] ), .S(\SUMB[17][4] ) );
  FA_X1 S2_17_5 ( .A(\ab[17][5] ), .B(\CARRYB[16][5] ), .CI(\SUMB[16][6] ), 
        .CO(\CARRYB[17][5] ), .S(\SUMB[17][5] ) );
  FA_X1 S2_17_6 ( .A(\ab[17][6] ), .B(\CARRYB[16][6] ), .CI(\SUMB[16][7] ), 
        .CO(\CARRYB[17][6] ), .S(\SUMB[17][6] ) );
  FA_X1 S2_17_7 ( .A(\ab[17][7] ), .B(\CARRYB[16][7] ), .CI(\SUMB[16][8] ), 
        .CO(\CARRYB[17][7] ), .S(\SUMB[17][7] ) );
  FA_X1 S2_17_8 ( .A(\ab[17][8] ), .B(\CARRYB[16][8] ), .CI(\SUMB[16][9] ), 
        .CO(\CARRYB[17][8] ), .S(\SUMB[17][8] ) );
  FA_X1 S2_17_9 ( .A(\ab[17][9] ), .B(\CARRYB[16][9] ), .CI(\SUMB[16][10] ), 
        .CO(\CARRYB[17][9] ), .S(\SUMB[17][9] ) );
  FA_X1 S2_17_10 ( .A(\ab[17][10] ), .B(\CARRYB[16][10] ), .CI(\SUMB[16][11] ), 
        .CO(\CARRYB[17][10] ), .S(\SUMB[17][10] ) );
  FA_X1 S2_17_11 ( .A(\ab[17][11] ), .B(\CARRYB[16][11] ), .CI(\SUMB[16][12] ), 
        .CO(\CARRYB[17][11] ), .S(\SUMB[17][11] ) );
  FA_X1 S2_17_12 ( .A(\ab[17][12] ), .B(\CARRYB[16][12] ), .CI(\SUMB[16][13] ), 
        .CO(\CARRYB[17][12] ), .S(\SUMB[17][12] ) );
  FA_X1 S2_17_13 ( .A(\ab[17][13] ), .B(\CARRYB[16][13] ), .CI(\SUMB[16][14] ), 
        .CO(\CARRYB[17][13] ), .S(\SUMB[17][13] ) );
  FA_X1 S2_17_14 ( .A(\ab[17][14] ), .B(\CARRYB[16][14] ), .CI(\SUMB[16][15] ), 
        .CO(\CARRYB[17][14] ), .S(\SUMB[17][14] ) );
  FA_X1 S2_17_15 ( .A(\ab[17][15] ), .B(\CARRYB[16][15] ), .CI(\SUMB[16][16] ), 
        .CO(\CARRYB[17][15] ), .S(\SUMB[17][15] ) );
  FA_X1 S2_17_16 ( .A(\ab[17][16] ), .B(\CARRYB[16][16] ), .CI(\SUMB[16][17] ), 
        .CO(\CARRYB[17][16] ), .S(\SUMB[17][16] ) );
  FA_X1 S2_17_17 ( .A(\ab[17][17] ), .B(\CARRYB[16][17] ), .CI(\SUMB[16][18] ), 
        .CO(\CARRYB[17][17] ), .S(\SUMB[17][17] ) );
  FA_X1 S2_17_18 ( .A(\ab[17][18] ), .B(\CARRYB[16][18] ), .CI(\SUMB[16][19] ), 
        .CO(\CARRYB[17][18] ), .S(\SUMB[17][18] ) );
  FA_X1 S2_17_19 ( .A(\ab[17][19] ), .B(\CARRYB[16][19] ), .CI(\SUMB[16][20] ), 
        .CO(\CARRYB[17][19] ), .S(\SUMB[17][19] ) );
  FA_X1 S2_17_20 ( .A(\ab[17][20] ), .B(\CARRYB[16][20] ), .CI(\SUMB[16][21] ), 
        .CO(\CARRYB[17][20] ), .S(\SUMB[17][20] ) );
  FA_X1 S2_17_21 ( .A(\ab[17][21] ), .B(\CARRYB[16][21] ), .CI(\SUMB[16][22] ), 
        .CO(\CARRYB[17][21] ), .S(\SUMB[17][21] ) );
  FA_X1 S2_17_22 ( .A(\ab[17][22] ), .B(\CARRYB[16][22] ), .CI(\SUMB[16][23] ), 
        .CO(\CARRYB[17][22] ), .S(\SUMB[17][22] ) );
  FA_X1 S2_17_23 ( .A(\ab[17][23] ), .B(\CARRYB[16][23] ), .CI(\SUMB[16][24] ), 
        .CO(\CARRYB[17][23] ), .S(\SUMB[17][23] ) );
  FA_X1 S2_17_24 ( .A(\ab[17][24] ), .B(\CARRYB[16][24] ), .CI(\SUMB[16][25] ), 
        .CO(\CARRYB[17][24] ), .S(\SUMB[17][24] ) );
  FA_X1 S2_17_25 ( .A(\ab[17][25] ), .B(\CARRYB[16][25] ), .CI(\SUMB[16][26] ), 
        .CO(\CARRYB[17][25] ), .S(\SUMB[17][25] ) );
  FA_X1 S2_17_26 ( .A(\ab[17][26] ), .B(\CARRYB[16][26] ), .CI(\SUMB[16][27] ), 
        .CO(\CARRYB[17][26] ), .S(\SUMB[17][26] ) );
  FA_X1 S2_17_27 ( .A(\ab[17][27] ), .B(\CARRYB[16][27] ), .CI(\SUMB[16][28] ), 
        .CO(\CARRYB[17][27] ), .S(\SUMB[17][27] ) );
  FA_X1 S2_17_28 ( .A(\ab[17][28] ), .B(\CARRYB[16][28] ), .CI(\SUMB[16][29] ), 
        .CO(\CARRYB[17][28] ), .S(\SUMB[17][28] ) );
  FA_X1 S2_17_29 ( .A(\ab[17][29] ), .B(\CARRYB[16][29] ), .CI(\SUMB[16][30] ), 
        .CO(\CARRYB[17][29] ), .S(\SUMB[17][29] ) );
  FA_X1 S2_17_30 ( .A(\ab[17][30] ), .B(\CARRYB[16][30] ), .CI(\SUMB[16][31] ), 
        .CO(\CARRYB[17][30] ), .S(\SUMB[17][30] ) );
  FA_X1 S2_17_31 ( .A(\ab[17][31] ), .B(\CARRYB[16][31] ), .CI(\SUMB[16][32] ), 
        .CO(\CARRYB[17][31] ), .S(\SUMB[17][31] ) );
  FA_X1 S2_17_32 ( .A(\ab[17][32] ), .B(\CARRYB[16][32] ), .CI(\SUMB[16][33] ), 
        .CO(\CARRYB[17][32] ), .S(\SUMB[17][32] ) );
  FA_X1 S2_17_33 ( .A(\ab[17][33] ), .B(\CARRYB[16][33] ), .CI(\SUMB[16][34] ), 
        .CO(\CARRYB[17][33] ), .S(\SUMB[17][33] ) );
  FA_X1 S2_17_34 ( .A(\ab[17][34] ), .B(\CARRYB[16][34] ), .CI(\SUMB[16][35] ), 
        .CO(\CARRYB[17][34] ), .S(\SUMB[17][34] ) );
  FA_X1 S2_17_35 ( .A(\ab[17][35] ), .B(\CARRYB[16][35] ), .CI(\SUMB[16][36] ), 
        .CO(\CARRYB[17][35] ), .S(\SUMB[17][35] ) );
  FA_X1 S2_17_36 ( .A(\ab[17][36] ), .B(\CARRYB[16][36] ), .CI(\SUMB[16][37] ), 
        .CO(\CARRYB[17][36] ), .S(\SUMB[17][36] ) );
  FA_X1 S2_17_37 ( .A(\ab[17][37] ), .B(\CARRYB[16][37] ), .CI(\SUMB[16][38] ), 
        .CO(\CARRYB[17][37] ), .S(\SUMB[17][37] ) );
  FA_X1 S2_17_38 ( .A(\ab[17][38] ), .B(\CARRYB[16][38] ), .CI(\SUMB[16][39] ), 
        .CO(\CARRYB[17][38] ), .S(\SUMB[17][38] ) );
  FA_X1 S2_17_39 ( .A(\ab[17][39] ), .B(\CARRYB[16][39] ), .CI(\SUMB[16][40] ), 
        .CO(\CARRYB[17][39] ), .S(\SUMB[17][39] ) );
  FA_X1 S2_17_40 ( .A(\ab[17][40] ), .B(\CARRYB[16][40] ), .CI(\SUMB[16][41] ), 
        .CO(\CARRYB[17][40] ), .S(\SUMB[17][40] ) );
  FA_X1 S2_17_41 ( .A(\ab[17][41] ), .B(\CARRYB[16][41] ), .CI(\SUMB[16][42] ), 
        .CO(\CARRYB[17][41] ), .S(\SUMB[17][41] ) );
  FA_X1 S2_17_42 ( .A(\ab[17][42] ), .B(\CARRYB[16][42] ), .CI(\SUMB[16][43] ), 
        .CO(\CARRYB[17][42] ), .S(\SUMB[17][42] ) );
  FA_X1 S2_17_43 ( .A(\ab[17][43] ), .B(\CARRYB[16][43] ), .CI(\SUMB[16][44] ), 
        .CO(\CARRYB[17][43] ), .S(\SUMB[17][43] ) );
  FA_X1 S2_17_44 ( .A(\ab[17][44] ), .B(\CARRYB[16][44] ), .CI(\SUMB[16][45] ), 
        .CO(\CARRYB[17][44] ), .S(\SUMB[17][44] ) );
  FA_X1 S2_17_45 ( .A(\ab[17][45] ), .B(\CARRYB[16][45] ), .CI(\SUMB[16][46] ), 
        .CO(\CARRYB[17][45] ), .S(\SUMB[17][45] ) );
  FA_X1 S2_17_46 ( .A(\ab[17][46] ), .B(\CARRYB[16][46] ), .CI(\SUMB[16][47] ), 
        .CO(\CARRYB[17][46] ), .S(\SUMB[17][46] ) );
  FA_X1 S2_17_47 ( .A(\ab[17][47] ), .B(\CARRYB[16][47] ), .CI(\SUMB[16][48] ), 
        .CO(\CARRYB[17][47] ), .S(\SUMB[17][47] ) );
  FA_X1 S2_17_48 ( .A(\ab[17][48] ), .B(\CARRYB[16][48] ), .CI(\SUMB[16][49] ), 
        .CO(\CARRYB[17][48] ), .S(\SUMB[17][48] ) );
  FA_X1 S2_17_49 ( .A(\ab[17][49] ), .B(\CARRYB[16][49] ), .CI(\SUMB[16][50] ), 
        .CO(\CARRYB[17][49] ), .S(\SUMB[17][49] ) );
  FA_X1 S2_17_50 ( .A(\ab[17][50] ), .B(\CARRYB[16][50] ), .CI(\SUMB[16][51] ), 
        .CO(\CARRYB[17][50] ), .S(\SUMB[17][50] ) );
  FA_X1 S3_17_51 ( .A(\ab[17][51] ), .B(\CARRYB[16][51] ), .CI(\ab[16][52] ), 
        .CO(\CARRYB[17][51] ), .S(\SUMB[17][51] ) );
  FA_X1 S1_16_0 ( .A(\ab[16][0] ), .B(\CARRYB[15][0] ), .CI(\SUMB[15][1] ), 
        .CO(\CARRYB[16][0] ), .S(CLA_SUM[16]) );
  FA_X1 S2_16_1 ( .A(\ab[16][1] ), .B(\CARRYB[15][1] ), .CI(\SUMB[15][2] ), 
        .CO(\CARRYB[16][1] ), .S(\SUMB[16][1] ) );
  FA_X1 S2_16_2 ( .A(\ab[16][2] ), .B(\CARRYB[15][2] ), .CI(\SUMB[15][3] ), 
        .CO(\CARRYB[16][2] ), .S(\SUMB[16][2] ) );
  FA_X1 S2_16_3 ( .A(\ab[16][3] ), .B(\CARRYB[15][3] ), .CI(\SUMB[15][4] ), 
        .CO(\CARRYB[16][3] ), .S(\SUMB[16][3] ) );
  FA_X1 S2_16_4 ( .A(\ab[16][4] ), .B(\CARRYB[15][4] ), .CI(\SUMB[15][5] ), 
        .CO(\CARRYB[16][4] ), .S(\SUMB[16][4] ) );
  FA_X1 S2_16_5 ( .A(\ab[16][5] ), .B(\CARRYB[15][5] ), .CI(\SUMB[15][6] ), 
        .CO(\CARRYB[16][5] ), .S(\SUMB[16][5] ) );
  FA_X1 S2_16_6 ( .A(\ab[16][6] ), .B(\CARRYB[15][6] ), .CI(\SUMB[15][7] ), 
        .CO(\CARRYB[16][6] ), .S(\SUMB[16][6] ) );
  FA_X1 S2_16_7 ( .A(\ab[16][7] ), .B(\CARRYB[15][7] ), .CI(\SUMB[15][8] ), 
        .CO(\CARRYB[16][7] ), .S(\SUMB[16][7] ) );
  FA_X1 S2_16_8 ( .A(\ab[16][8] ), .B(\CARRYB[15][8] ), .CI(\SUMB[15][9] ), 
        .CO(\CARRYB[16][8] ), .S(\SUMB[16][8] ) );
  FA_X1 S2_16_9 ( .A(\ab[16][9] ), .B(\CARRYB[15][9] ), .CI(\SUMB[15][10] ), 
        .CO(\CARRYB[16][9] ), .S(\SUMB[16][9] ) );
  FA_X1 S2_16_10 ( .A(\ab[16][10] ), .B(\CARRYB[15][10] ), .CI(\SUMB[15][11] ), 
        .CO(\CARRYB[16][10] ), .S(\SUMB[16][10] ) );
  FA_X1 S2_16_11 ( .A(\ab[16][11] ), .B(\CARRYB[15][11] ), .CI(\SUMB[15][12] ), 
        .CO(\CARRYB[16][11] ), .S(\SUMB[16][11] ) );
  FA_X1 S2_16_12 ( .A(\ab[16][12] ), .B(\CARRYB[15][12] ), .CI(\SUMB[15][13] ), 
        .CO(\CARRYB[16][12] ), .S(\SUMB[16][12] ) );
  FA_X1 S2_16_13 ( .A(\ab[16][13] ), .B(\CARRYB[15][13] ), .CI(\SUMB[15][14] ), 
        .CO(\CARRYB[16][13] ), .S(\SUMB[16][13] ) );
  FA_X1 S2_16_14 ( .A(\ab[16][14] ), .B(\CARRYB[15][14] ), .CI(\SUMB[15][15] ), 
        .CO(\CARRYB[16][14] ), .S(\SUMB[16][14] ) );
  FA_X1 S2_16_15 ( .A(\ab[16][15] ), .B(\CARRYB[15][15] ), .CI(\SUMB[15][16] ), 
        .CO(\CARRYB[16][15] ), .S(\SUMB[16][15] ) );
  FA_X1 S2_16_16 ( .A(\ab[16][16] ), .B(\CARRYB[15][16] ), .CI(\SUMB[15][17] ), 
        .CO(\CARRYB[16][16] ), .S(\SUMB[16][16] ) );
  FA_X1 S2_16_17 ( .A(\ab[16][17] ), .B(\CARRYB[15][17] ), .CI(\SUMB[15][18] ), 
        .CO(\CARRYB[16][17] ), .S(\SUMB[16][17] ) );
  FA_X1 S2_16_18 ( .A(\ab[16][18] ), .B(\CARRYB[15][18] ), .CI(\SUMB[15][19] ), 
        .CO(\CARRYB[16][18] ), .S(\SUMB[16][18] ) );
  FA_X1 S2_16_19 ( .A(\ab[16][19] ), .B(\CARRYB[15][19] ), .CI(\SUMB[15][20] ), 
        .CO(\CARRYB[16][19] ), .S(\SUMB[16][19] ) );
  FA_X1 S2_16_20 ( .A(\ab[16][20] ), .B(\CARRYB[15][20] ), .CI(\SUMB[15][21] ), 
        .CO(\CARRYB[16][20] ), .S(\SUMB[16][20] ) );
  FA_X1 S2_16_21 ( .A(\ab[16][21] ), .B(\CARRYB[15][21] ), .CI(\SUMB[15][22] ), 
        .CO(\CARRYB[16][21] ), .S(\SUMB[16][21] ) );
  FA_X1 S2_16_22 ( .A(\ab[16][22] ), .B(\CARRYB[15][22] ), .CI(\SUMB[15][23] ), 
        .CO(\CARRYB[16][22] ), .S(\SUMB[16][22] ) );
  FA_X1 S2_16_23 ( .A(\ab[16][23] ), .B(\CARRYB[15][23] ), .CI(\SUMB[15][24] ), 
        .CO(\CARRYB[16][23] ), .S(\SUMB[16][23] ) );
  FA_X1 S2_16_24 ( .A(\ab[16][24] ), .B(\CARRYB[15][24] ), .CI(\SUMB[15][25] ), 
        .CO(\CARRYB[16][24] ), .S(\SUMB[16][24] ) );
  FA_X1 S2_16_25 ( .A(\ab[16][25] ), .B(\CARRYB[15][25] ), .CI(\SUMB[15][26] ), 
        .CO(\CARRYB[16][25] ), .S(\SUMB[16][25] ) );
  FA_X1 S2_16_26 ( .A(\ab[16][26] ), .B(\CARRYB[15][26] ), .CI(\SUMB[15][27] ), 
        .CO(\CARRYB[16][26] ), .S(\SUMB[16][26] ) );
  FA_X1 S2_16_27 ( .A(\ab[16][27] ), .B(\CARRYB[15][27] ), .CI(\SUMB[15][28] ), 
        .CO(\CARRYB[16][27] ), .S(\SUMB[16][27] ) );
  FA_X1 S2_16_28 ( .A(\ab[16][28] ), .B(\CARRYB[15][28] ), .CI(\SUMB[15][29] ), 
        .CO(\CARRYB[16][28] ), .S(\SUMB[16][28] ) );
  FA_X1 S2_16_29 ( .A(\ab[16][29] ), .B(\CARRYB[15][29] ), .CI(\SUMB[15][30] ), 
        .CO(\CARRYB[16][29] ), .S(\SUMB[16][29] ) );
  FA_X1 S2_16_30 ( .A(\ab[16][30] ), .B(\CARRYB[15][30] ), .CI(\SUMB[15][31] ), 
        .CO(\CARRYB[16][30] ), .S(\SUMB[16][30] ) );
  FA_X1 S2_16_31 ( .A(\ab[16][31] ), .B(\CARRYB[15][31] ), .CI(\SUMB[15][32] ), 
        .CO(\CARRYB[16][31] ), .S(\SUMB[16][31] ) );
  FA_X1 S2_16_32 ( .A(\ab[16][32] ), .B(\CARRYB[15][32] ), .CI(\SUMB[15][33] ), 
        .CO(\CARRYB[16][32] ), .S(\SUMB[16][32] ) );
  FA_X1 S2_16_33 ( .A(\ab[16][33] ), .B(\CARRYB[15][33] ), .CI(\SUMB[15][34] ), 
        .CO(\CARRYB[16][33] ), .S(\SUMB[16][33] ) );
  FA_X1 S2_16_34 ( .A(\ab[16][34] ), .B(\CARRYB[15][34] ), .CI(\SUMB[15][35] ), 
        .CO(\CARRYB[16][34] ), .S(\SUMB[16][34] ) );
  FA_X1 S2_16_35 ( .A(\ab[16][35] ), .B(\CARRYB[15][35] ), .CI(\SUMB[15][36] ), 
        .CO(\CARRYB[16][35] ), .S(\SUMB[16][35] ) );
  FA_X1 S2_16_36 ( .A(\ab[16][36] ), .B(\CARRYB[15][36] ), .CI(\SUMB[15][37] ), 
        .CO(\CARRYB[16][36] ), .S(\SUMB[16][36] ) );
  FA_X1 S2_16_37 ( .A(\ab[16][37] ), .B(\CARRYB[15][37] ), .CI(\SUMB[15][38] ), 
        .CO(\CARRYB[16][37] ), .S(\SUMB[16][37] ) );
  FA_X1 S2_16_38 ( .A(\ab[16][38] ), .B(\CARRYB[15][38] ), .CI(\SUMB[15][39] ), 
        .CO(\CARRYB[16][38] ), .S(\SUMB[16][38] ) );
  FA_X1 S2_16_39 ( .A(\ab[16][39] ), .B(\CARRYB[15][39] ), .CI(\SUMB[15][40] ), 
        .CO(\CARRYB[16][39] ), .S(\SUMB[16][39] ) );
  FA_X1 S2_16_40 ( .A(\ab[16][40] ), .B(\CARRYB[15][40] ), .CI(\SUMB[15][41] ), 
        .CO(\CARRYB[16][40] ), .S(\SUMB[16][40] ) );
  FA_X1 S2_16_41 ( .A(\ab[16][41] ), .B(\CARRYB[15][41] ), .CI(\SUMB[15][42] ), 
        .CO(\CARRYB[16][41] ), .S(\SUMB[16][41] ) );
  FA_X1 S2_16_42 ( .A(\ab[16][42] ), .B(\CARRYB[15][42] ), .CI(\SUMB[15][43] ), 
        .CO(\CARRYB[16][42] ), .S(\SUMB[16][42] ) );
  FA_X1 S2_16_43 ( .A(\ab[16][43] ), .B(\CARRYB[15][43] ), .CI(\SUMB[15][44] ), 
        .CO(\CARRYB[16][43] ), .S(\SUMB[16][43] ) );
  FA_X1 S2_16_44 ( .A(\ab[16][44] ), .B(\CARRYB[15][44] ), .CI(\SUMB[15][45] ), 
        .CO(\CARRYB[16][44] ), .S(\SUMB[16][44] ) );
  FA_X1 S2_16_45 ( .A(\ab[16][45] ), .B(\CARRYB[15][45] ), .CI(\SUMB[15][46] ), 
        .CO(\CARRYB[16][45] ), .S(\SUMB[16][45] ) );
  FA_X1 S2_16_46 ( .A(\ab[16][46] ), .B(\CARRYB[15][46] ), .CI(\SUMB[15][47] ), 
        .CO(\CARRYB[16][46] ), .S(\SUMB[16][46] ) );
  FA_X1 S2_16_47 ( .A(\ab[16][47] ), .B(\CARRYB[15][47] ), .CI(\SUMB[15][48] ), 
        .CO(\CARRYB[16][47] ), .S(\SUMB[16][47] ) );
  FA_X1 S2_16_48 ( .A(\ab[16][48] ), .B(\CARRYB[15][48] ), .CI(\SUMB[15][49] ), 
        .CO(\CARRYB[16][48] ), .S(\SUMB[16][48] ) );
  FA_X1 S2_16_49 ( .A(\ab[16][49] ), .B(\CARRYB[15][49] ), .CI(\SUMB[15][50] ), 
        .CO(\CARRYB[16][49] ), .S(\SUMB[16][49] ) );
  FA_X1 S2_16_50 ( .A(\ab[16][50] ), .B(\CARRYB[15][50] ), .CI(\SUMB[15][51] ), 
        .CO(\CARRYB[16][50] ), .S(\SUMB[16][50] ) );
  FA_X1 S3_16_51 ( .A(\ab[16][51] ), .B(\CARRYB[15][51] ), .CI(\ab[15][52] ), 
        .CO(\CARRYB[16][51] ), .S(\SUMB[16][51] ) );
  FA_X1 S1_15_0 ( .A(\ab[15][0] ), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), 
        .CO(\CARRYB[15][0] ), .S(CLA_SUM[15]) );
  FA_X1 S2_15_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), 
        .CO(\CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FA_X1 S2_15_2 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), 
        .CO(\CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FA_X1 S2_15_3 ( .A(\ab[15][3] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), 
        .CO(\CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FA_X1 S2_15_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), 
        .CO(\CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FA_X1 S2_15_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), 
        .CO(\CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FA_X1 S2_15_6 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), 
        .CO(\CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FA_X1 S2_15_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), 
        .CO(\CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FA_X1 S2_15_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), 
        .CO(\CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FA_X1 S2_15_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), 
        .CO(\CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FA_X1 S2_15_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .CI(\SUMB[14][11] ), 
        .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FA_X1 S2_15_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .CI(\SUMB[14][12] ), 
        .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FA_X1 S2_15_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .CI(\SUMB[14][13] ), 
        .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FA_X1 S2_15_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), 
        .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FA_X1 S2_15_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(\SUMB[14][15] ), 
        .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FA_X1 S2_15_15 ( .A(\ab[15][15] ), .B(\CARRYB[14][15] ), .CI(\SUMB[14][16] ), 
        .CO(\CARRYB[15][15] ), .S(\SUMB[15][15] ) );
  FA_X1 S2_15_16 ( .A(\ab[15][16] ), .B(\CARRYB[14][16] ), .CI(\SUMB[14][17] ), 
        .CO(\CARRYB[15][16] ), .S(\SUMB[15][16] ) );
  FA_X1 S2_15_17 ( .A(\ab[15][17] ), .B(\CARRYB[14][17] ), .CI(\SUMB[14][18] ), 
        .CO(\CARRYB[15][17] ), .S(\SUMB[15][17] ) );
  FA_X1 S2_15_18 ( .A(\ab[15][18] ), .B(\CARRYB[14][18] ), .CI(\SUMB[14][19] ), 
        .CO(\CARRYB[15][18] ), .S(\SUMB[15][18] ) );
  FA_X1 S2_15_19 ( .A(\ab[15][19] ), .B(\CARRYB[14][19] ), .CI(\SUMB[14][20] ), 
        .CO(\CARRYB[15][19] ), .S(\SUMB[15][19] ) );
  FA_X1 S2_15_20 ( .A(\ab[15][20] ), .B(\CARRYB[14][20] ), .CI(\SUMB[14][21] ), 
        .CO(\CARRYB[15][20] ), .S(\SUMB[15][20] ) );
  FA_X1 S2_15_21 ( .A(\ab[15][21] ), .B(\CARRYB[14][21] ), .CI(\SUMB[14][22] ), 
        .CO(\CARRYB[15][21] ), .S(\SUMB[15][21] ) );
  FA_X1 S2_15_22 ( .A(\ab[15][22] ), .B(\CARRYB[14][22] ), .CI(\SUMB[14][23] ), 
        .CO(\CARRYB[15][22] ), .S(\SUMB[15][22] ) );
  FA_X1 S2_15_23 ( .A(\ab[15][23] ), .B(\CARRYB[14][23] ), .CI(\SUMB[14][24] ), 
        .CO(\CARRYB[15][23] ), .S(\SUMB[15][23] ) );
  FA_X1 S2_15_24 ( .A(\ab[15][24] ), .B(\CARRYB[14][24] ), .CI(\SUMB[14][25] ), 
        .CO(\CARRYB[15][24] ), .S(\SUMB[15][24] ) );
  FA_X1 S2_15_25 ( .A(\ab[15][25] ), .B(\CARRYB[14][25] ), .CI(\SUMB[14][26] ), 
        .CO(\CARRYB[15][25] ), .S(\SUMB[15][25] ) );
  FA_X1 S2_15_26 ( .A(\ab[15][26] ), .B(\CARRYB[14][26] ), .CI(\SUMB[14][27] ), 
        .CO(\CARRYB[15][26] ), .S(\SUMB[15][26] ) );
  FA_X1 S2_15_27 ( .A(\ab[15][27] ), .B(\CARRYB[14][27] ), .CI(\SUMB[14][28] ), 
        .CO(\CARRYB[15][27] ), .S(\SUMB[15][27] ) );
  FA_X1 S2_15_28 ( .A(\ab[15][28] ), .B(\CARRYB[14][28] ), .CI(\SUMB[14][29] ), 
        .CO(\CARRYB[15][28] ), .S(\SUMB[15][28] ) );
  FA_X1 S2_15_29 ( .A(\ab[15][29] ), .B(\CARRYB[14][29] ), .CI(\SUMB[14][30] ), 
        .CO(\CARRYB[15][29] ), .S(\SUMB[15][29] ) );
  FA_X1 S2_15_30 ( .A(\ab[15][30] ), .B(\CARRYB[14][30] ), .CI(\SUMB[14][31] ), 
        .CO(\CARRYB[15][30] ), .S(\SUMB[15][30] ) );
  FA_X1 S2_15_31 ( .A(\ab[15][31] ), .B(\CARRYB[14][31] ), .CI(\SUMB[14][32] ), 
        .CO(\CARRYB[15][31] ), .S(\SUMB[15][31] ) );
  FA_X1 S2_15_32 ( .A(\ab[15][32] ), .B(\CARRYB[14][32] ), .CI(\SUMB[14][33] ), 
        .CO(\CARRYB[15][32] ), .S(\SUMB[15][32] ) );
  FA_X1 S2_15_33 ( .A(\ab[15][33] ), .B(\CARRYB[14][33] ), .CI(\SUMB[14][34] ), 
        .CO(\CARRYB[15][33] ), .S(\SUMB[15][33] ) );
  FA_X1 S2_15_34 ( .A(\ab[15][34] ), .B(\CARRYB[14][34] ), .CI(\SUMB[14][35] ), 
        .CO(\CARRYB[15][34] ), .S(\SUMB[15][34] ) );
  FA_X1 S2_15_35 ( .A(\ab[15][35] ), .B(\CARRYB[14][35] ), .CI(\SUMB[14][36] ), 
        .CO(\CARRYB[15][35] ), .S(\SUMB[15][35] ) );
  FA_X1 S2_15_36 ( .A(\ab[15][36] ), .B(\CARRYB[14][36] ), .CI(\SUMB[14][37] ), 
        .CO(\CARRYB[15][36] ), .S(\SUMB[15][36] ) );
  FA_X1 S2_15_37 ( .A(\ab[15][37] ), .B(\CARRYB[14][37] ), .CI(\SUMB[14][38] ), 
        .CO(\CARRYB[15][37] ), .S(\SUMB[15][37] ) );
  FA_X1 S2_15_38 ( .A(\ab[15][38] ), .B(\CARRYB[14][38] ), .CI(\SUMB[14][39] ), 
        .CO(\CARRYB[15][38] ), .S(\SUMB[15][38] ) );
  FA_X1 S2_15_39 ( .A(\ab[15][39] ), .B(\CARRYB[14][39] ), .CI(\SUMB[14][40] ), 
        .CO(\CARRYB[15][39] ), .S(\SUMB[15][39] ) );
  FA_X1 S2_15_40 ( .A(\ab[15][40] ), .B(\CARRYB[14][40] ), .CI(\SUMB[14][41] ), 
        .CO(\CARRYB[15][40] ), .S(\SUMB[15][40] ) );
  FA_X1 S2_15_41 ( .A(\ab[15][41] ), .B(\CARRYB[14][41] ), .CI(\SUMB[14][42] ), 
        .CO(\CARRYB[15][41] ), .S(\SUMB[15][41] ) );
  FA_X1 S2_15_42 ( .A(\ab[15][42] ), .B(\CARRYB[14][42] ), .CI(\SUMB[14][43] ), 
        .CO(\CARRYB[15][42] ), .S(\SUMB[15][42] ) );
  FA_X1 S2_15_43 ( .A(\ab[15][43] ), .B(\CARRYB[14][43] ), .CI(\SUMB[14][44] ), 
        .CO(\CARRYB[15][43] ), .S(\SUMB[15][43] ) );
  FA_X1 S2_15_44 ( .A(\ab[15][44] ), .B(\CARRYB[14][44] ), .CI(\SUMB[14][45] ), 
        .CO(\CARRYB[15][44] ), .S(\SUMB[15][44] ) );
  FA_X1 S2_15_45 ( .A(\ab[15][45] ), .B(\CARRYB[14][45] ), .CI(\SUMB[14][46] ), 
        .CO(\CARRYB[15][45] ), .S(\SUMB[15][45] ) );
  FA_X1 S2_15_46 ( .A(\ab[15][46] ), .B(\CARRYB[14][46] ), .CI(\SUMB[14][47] ), 
        .CO(\CARRYB[15][46] ), .S(\SUMB[15][46] ) );
  FA_X1 S2_15_47 ( .A(\ab[15][47] ), .B(\CARRYB[14][47] ), .CI(\SUMB[14][48] ), 
        .CO(\CARRYB[15][47] ), .S(\SUMB[15][47] ) );
  FA_X1 S2_15_48 ( .A(\ab[15][48] ), .B(\CARRYB[14][48] ), .CI(\SUMB[14][49] ), 
        .CO(\CARRYB[15][48] ), .S(\SUMB[15][48] ) );
  FA_X1 S2_15_49 ( .A(\ab[15][49] ), .B(\CARRYB[14][49] ), .CI(\SUMB[14][50] ), 
        .CO(\CARRYB[15][49] ), .S(\SUMB[15][49] ) );
  FA_X1 S2_15_50 ( .A(\ab[15][50] ), .B(\CARRYB[14][50] ), .CI(\SUMB[14][51] ), 
        .CO(\CARRYB[15][50] ), .S(\SUMB[15][50] ) );
  FA_X1 S3_15_51 ( .A(\ab[15][51] ), .B(\CARRYB[14][51] ), .CI(\ab[14][52] ), 
        .CO(\CARRYB[15][51] ), .S(\SUMB[15][51] ) );
  FA_X1 S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), 
        .CO(\CARRYB[14][0] ), .S(CLA_SUM[14]) );
  FA_X1 S2_14_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), 
        .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA_X1 S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), 
        .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA_X1 S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), 
        .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FA_X1 S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA_X1 S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), 
        .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA_X1 S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), 
        .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FA_X1 S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), 
        .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA_X1 S2_14_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA_X1 S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), 
        .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA_X1 S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA_X1 S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), 
        .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA_X1 S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), 
        .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA_X1 S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), 
        .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FA_X1 S2_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\SUMB[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA_X1 S2_14_15 ( .A(\ab[14][15] ), .B(\CARRYB[13][15] ), .CI(\SUMB[13][16] ), 
        .CO(\CARRYB[14][15] ), .S(\SUMB[14][15] ) );
  FA_X1 S2_14_16 ( .A(\ab[14][16] ), .B(\CARRYB[13][16] ), .CI(\SUMB[13][17] ), 
        .CO(\CARRYB[14][16] ), .S(\SUMB[14][16] ) );
  FA_X1 S2_14_17 ( .A(\ab[14][17] ), .B(\CARRYB[13][17] ), .CI(\SUMB[13][18] ), 
        .CO(\CARRYB[14][17] ), .S(\SUMB[14][17] ) );
  FA_X1 S2_14_18 ( .A(\ab[14][18] ), .B(\CARRYB[13][18] ), .CI(\SUMB[13][19] ), 
        .CO(\CARRYB[14][18] ), .S(\SUMB[14][18] ) );
  FA_X1 S2_14_19 ( .A(\ab[14][19] ), .B(\CARRYB[13][19] ), .CI(\SUMB[13][20] ), 
        .CO(\CARRYB[14][19] ), .S(\SUMB[14][19] ) );
  FA_X1 S2_14_20 ( .A(\ab[14][20] ), .B(\CARRYB[13][20] ), .CI(\SUMB[13][21] ), 
        .CO(\CARRYB[14][20] ), .S(\SUMB[14][20] ) );
  FA_X1 S2_14_21 ( .A(\ab[14][21] ), .B(\CARRYB[13][21] ), .CI(\SUMB[13][22] ), 
        .CO(\CARRYB[14][21] ), .S(\SUMB[14][21] ) );
  FA_X1 S2_14_22 ( .A(\ab[14][22] ), .B(\CARRYB[13][22] ), .CI(\SUMB[13][23] ), 
        .CO(\CARRYB[14][22] ), .S(\SUMB[14][22] ) );
  FA_X1 S2_14_23 ( .A(\ab[14][23] ), .B(\CARRYB[13][23] ), .CI(\SUMB[13][24] ), 
        .CO(\CARRYB[14][23] ), .S(\SUMB[14][23] ) );
  FA_X1 S2_14_24 ( .A(\ab[14][24] ), .B(\CARRYB[13][24] ), .CI(\SUMB[13][25] ), 
        .CO(\CARRYB[14][24] ), .S(\SUMB[14][24] ) );
  FA_X1 S2_14_25 ( .A(\ab[14][25] ), .B(\CARRYB[13][25] ), .CI(\SUMB[13][26] ), 
        .CO(\CARRYB[14][25] ), .S(\SUMB[14][25] ) );
  FA_X1 S2_14_26 ( .A(\ab[14][26] ), .B(\CARRYB[13][26] ), .CI(\SUMB[13][27] ), 
        .CO(\CARRYB[14][26] ), .S(\SUMB[14][26] ) );
  FA_X1 S2_14_27 ( .A(\ab[14][27] ), .B(\CARRYB[13][27] ), .CI(\SUMB[13][28] ), 
        .CO(\CARRYB[14][27] ), .S(\SUMB[14][27] ) );
  FA_X1 S2_14_28 ( .A(\ab[14][28] ), .B(\CARRYB[13][28] ), .CI(\SUMB[13][29] ), 
        .CO(\CARRYB[14][28] ), .S(\SUMB[14][28] ) );
  FA_X1 S2_14_29 ( .A(\ab[14][29] ), .B(\CARRYB[13][29] ), .CI(\SUMB[13][30] ), 
        .CO(\CARRYB[14][29] ), .S(\SUMB[14][29] ) );
  FA_X1 S2_14_30 ( .A(\ab[14][30] ), .B(\CARRYB[13][30] ), .CI(\SUMB[13][31] ), 
        .CO(\CARRYB[14][30] ), .S(\SUMB[14][30] ) );
  FA_X1 S2_14_31 ( .A(\ab[14][31] ), .B(\CARRYB[13][31] ), .CI(\SUMB[13][32] ), 
        .CO(\CARRYB[14][31] ), .S(\SUMB[14][31] ) );
  FA_X1 S2_14_32 ( .A(\ab[14][32] ), .B(\CARRYB[13][32] ), .CI(\SUMB[13][33] ), 
        .CO(\CARRYB[14][32] ), .S(\SUMB[14][32] ) );
  FA_X1 S2_14_33 ( .A(\ab[14][33] ), .B(\CARRYB[13][33] ), .CI(\SUMB[13][34] ), 
        .CO(\CARRYB[14][33] ), .S(\SUMB[14][33] ) );
  FA_X1 S2_14_34 ( .A(\ab[14][34] ), .B(\CARRYB[13][34] ), .CI(\SUMB[13][35] ), 
        .CO(\CARRYB[14][34] ), .S(\SUMB[14][34] ) );
  FA_X1 S2_14_35 ( .A(\ab[14][35] ), .B(\CARRYB[13][35] ), .CI(\SUMB[13][36] ), 
        .CO(\CARRYB[14][35] ), .S(\SUMB[14][35] ) );
  FA_X1 S2_14_36 ( .A(\ab[14][36] ), .B(\CARRYB[13][36] ), .CI(\SUMB[13][37] ), 
        .CO(\CARRYB[14][36] ), .S(\SUMB[14][36] ) );
  FA_X1 S2_14_37 ( .A(\ab[14][37] ), .B(\CARRYB[13][37] ), .CI(\SUMB[13][38] ), 
        .CO(\CARRYB[14][37] ), .S(\SUMB[14][37] ) );
  FA_X1 S2_14_38 ( .A(\ab[14][38] ), .B(\CARRYB[13][38] ), .CI(\SUMB[13][39] ), 
        .CO(\CARRYB[14][38] ), .S(\SUMB[14][38] ) );
  FA_X1 S2_14_39 ( .A(\ab[14][39] ), .B(\CARRYB[13][39] ), .CI(\SUMB[13][40] ), 
        .CO(\CARRYB[14][39] ), .S(\SUMB[14][39] ) );
  FA_X1 S2_14_40 ( .A(\ab[14][40] ), .B(\CARRYB[13][40] ), .CI(\SUMB[13][41] ), 
        .CO(\CARRYB[14][40] ), .S(\SUMB[14][40] ) );
  FA_X1 S2_14_41 ( .A(\ab[14][41] ), .B(\CARRYB[13][41] ), .CI(\SUMB[13][42] ), 
        .CO(\CARRYB[14][41] ), .S(\SUMB[14][41] ) );
  FA_X1 S2_14_42 ( .A(\ab[14][42] ), .B(\CARRYB[13][42] ), .CI(\SUMB[13][43] ), 
        .CO(\CARRYB[14][42] ), .S(\SUMB[14][42] ) );
  FA_X1 S2_14_43 ( .A(\ab[14][43] ), .B(\CARRYB[13][43] ), .CI(\SUMB[13][44] ), 
        .CO(\CARRYB[14][43] ), .S(\SUMB[14][43] ) );
  FA_X1 S2_14_44 ( .A(\ab[14][44] ), .B(\CARRYB[13][44] ), .CI(\SUMB[13][45] ), 
        .CO(\CARRYB[14][44] ), .S(\SUMB[14][44] ) );
  FA_X1 S2_14_45 ( .A(\ab[14][45] ), .B(\CARRYB[13][45] ), .CI(\SUMB[13][46] ), 
        .CO(\CARRYB[14][45] ), .S(\SUMB[14][45] ) );
  FA_X1 S2_14_46 ( .A(\ab[14][46] ), .B(\CARRYB[13][46] ), .CI(\SUMB[13][47] ), 
        .CO(\CARRYB[14][46] ), .S(\SUMB[14][46] ) );
  FA_X1 S2_14_47 ( .A(\ab[14][47] ), .B(\CARRYB[13][47] ), .CI(\SUMB[13][48] ), 
        .CO(\CARRYB[14][47] ), .S(\SUMB[14][47] ) );
  FA_X1 S2_14_48 ( .A(\ab[14][48] ), .B(\CARRYB[13][48] ), .CI(\SUMB[13][49] ), 
        .CO(\CARRYB[14][48] ), .S(\SUMB[14][48] ) );
  FA_X1 S2_14_49 ( .A(\ab[14][49] ), .B(\CARRYB[13][49] ), .CI(\SUMB[13][50] ), 
        .CO(\CARRYB[14][49] ), .S(\SUMB[14][49] ) );
  FA_X1 S2_14_50 ( .A(\ab[14][50] ), .B(\CARRYB[13][50] ), .CI(\SUMB[13][51] ), 
        .CO(\CARRYB[14][50] ), .S(\SUMB[14][50] ) );
  FA_X1 S3_14_51 ( .A(\ab[14][51] ), .B(\CARRYB[13][51] ), .CI(\ab[13][52] ), 
        .CO(\CARRYB[14][51] ), .S(\SUMB[14][51] ) );
  FA_X1 S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(CLA_SUM[13]) );
  FA_X1 S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA_X1 S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA_X1 S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA_X1 S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA_X1 S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA_X1 S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA_X1 S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA_X1 S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA_X1 S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA_X1 S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA_X1 S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), 
        .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FA_X1 S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), 
        .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FA_X1 S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), 
        .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA_X1 S2_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\SUMB[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA_X1 S2_13_15 ( .A(\ab[13][15] ), .B(\CARRYB[12][15] ), .CI(\SUMB[12][16] ), 
        .CO(\CARRYB[13][15] ), .S(\SUMB[13][15] ) );
  FA_X1 S2_13_16 ( .A(\ab[13][16] ), .B(\CARRYB[12][16] ), .CI(\SUMB[12][17] ), 
        .CO(\CARRYB[13][16] ), .S(\SUMB[13][16] ) );
  FA_X1 S2_13_17 ( .A(\ab[13][17] ), .B(\CARRYB[12][17] ), .CI(\SUMB[12][18] ), 
        .CO(\CARRYB[13][17] ), .S(\SUMB[13][17] ) );
  FA_X1 S2_13_18 ( .A(\ab[13][18] ), .B(\CARRYB[12][18] ), .CI(\SUMB[12][19] ), 
        .CO(\CARRYB[13][18] ), .S(\SUMB[13][18] ) );
  FA_X1 S2_13_19 ( .A(\ab[13][19] ), .B(\CARRYB[12][19] ), .CI(\SUMB[12][20] ), 
        .CO(\CARRYB[13][19] ), .S(\SUMB[13][19] ) );
  FA_X1 S2_13_20 ( .A(\ab[13][20] ), .B(\CARRYB[12][20] ), .CI(\SUMB[12][21] ), 
        .CO(\CARRYB[13][20] ), .S(\SUMB[13][20] ) );
  FA_X1 S2_13_21 ( .A(\ab[13][21] ), .B(\CARRYB[12][21] ), .CI(\SUMB[12][22] ), 
        .CO(\CARRYB[13][21] ), .S(\SUMB[13][21] ) );
  FA_X1 S2_13_22 ( .A(\ab[13][22] ), .B(\CARRYB[12][22] ), .CI(\SUMB[12][23] ), 
        .CO(\CARRYB[13][22] ), .S(\SUMB[13][22] ) );
  FA_X1 S2_13_23 ( .A(\ab[13][23] ), .B(\CARRYB[12][23] ), .CI(\SUMB[12][24] ), 
        .CO(\CARRYB[13][23] ), .S(\SUMB[13][23] ) );
  FA_X1 S2_13_24 ( .A(\ab[13][24] ), .B(\CARRYB[12][24] ), .CI(\SUMB[12][25] ), 
        .CO(\CARRYB[13][24] ), .S(\SUMB[13][24] ) );
  FA_X1 S2_13_25 ( .A(\ab[13][25] ), .B(\CARRYB[12][25] ), .CI(\SUMB[12][26] ), 
        .CO(\CARRYB[13][25] ), .S(\SUMB[13][25] ) );
  FA_X1 S2_13_26 ( .A(\ab[13][26] ), .B(\CARRYB[12][26] ), .CI(\SUMB[12][27] ), 
        .CO(\CARRYB[13][26] ), .S(\SUMB[13][26] ) );
  FA_X1 S2_13_27 ( .A(\ab[13][27] ), .B(\CARRYB[12][27] ), .CI(\SUMB[12][28] ), 
        .CO(\CARRYB[13][27] ), .S(\SUMB[13][27] ) );
  FA_X1 S2_13_28 ( .A(\ab[13][28] ), .B(\CARRYB[12][28] ), .CI(\SUMB[12][29] ), 
        .CO(\CARRYB[13][28] ), .S(\SUMB[13][28] ) );
  FA_X1 S2_13_29 ( .A(\ab[13][29] ), .B(\CARRYB[12][29] ), .CI(\SUMB[12][30] ), 
        .CO(\CARRYB[13][29] ), .S(\SUMB[13][29] ) );
  FA_X1 S2_13_30 ( .A(\ab[13][30] ), .B(\CARRYB[12][30] ), .CI(\SUMB[12][31] ), 
        .CO(\CARRYB[13][30] ), .S(\SUMB[13][30] ) );
  FA_X1 S2_13_31 ( .A(\ab[13][31] ), .B(\CARRYB[12][31] ), .CI(\SUMB[12][32] ), 
        .CO(\CARRYB[13][31] ), .S(\SUMB[13][31] ) );
  FA_X1 S2_13_32 ( .A(\ab[13][32] ), .B(\CARRYB[12][32] ), .CI(\SUMB[12][33] ), 
        .CO(\CARRYB[13][32] ), .S(\SUMB[13][32] ) );
  FA_X1 S2_13_33 ( .A(\ab[13][33] ), .B(\CARRYB[12][33] ), .CI(\SUMB[12][34] ), 
        .CO(\CARRYB[13][33] ), .S(\SUMB[13][33] ) );
  FA_X1 S2_13_34 ( .A(\ab[13][34] ), .B(\CARRYB[12][34] ), .CI(\SUMB[12][35] ), 
        .CO(\CARRYB[13][34] ), .S(\SUMB[13][34] ) );
  FA_X1 S2_13_35 ( .A(\ab[13][35] ), .B(\CARRYB[12][35] ), .CI(\SUMB[12][36] ), 
        .CO(\CARRYB[13][35] ), .S(\SUMB[13][35] ) );
  FA_X1 S2_13_36 ( .A(\ab[13][36] ), .B(\CARRYB[12][36] ), .CI(\SUMB[12][37] ), 
        .CO(\CARRYB[13][36] ), .S(\SUMB[13][36] ) );
  FA_X1 S2_13_37 ( .A(\ab[13][37] ), .B(\CARRYB[12][37] ), .CI(\SUMB[12][38] ), 
        .CO(\CARRYB[13][37] ), .S(\SUMB[13][37] ) );
  FA_X1 S2_13_38 ( .A(\ab[13][38] ), .B(\CARRYB[12][38] ), .CI(\SUMB[12][39] ), 
        .CO(\CARRYB[13][38] ), .S(\SUMB[13][38] ) );
  FA_X1 S2_13_39 ( .A(\ab[13][39] ), .B(\CARRYB[12][39] ), .CI(\SUMB[12][40] ), 
        .CO(\CARRYB[13][39] ), .S(\SUMB[13][39] ) );
  FA_X1 S2_13_40 ( .A(\ab[13][40] ), .B(\CARRYB[12][40] ), .CI(\SUMB[12][41] ), 
        .CO(\CARRYB[13][40] ), .S(\SUMB[13][40] ) );
  FA_X1 S2_13_41 ( .A(\ab[13][41] ), .B(\CARRYB[12][41] ), .CI(\SUMB[12][42] ), 
        .CO(\CARRYB[13][41] ), .S(\SUMB[13][41] ) );
  FA_X1 S2_13_42 ( .A(\ab[13][42] ), .B(\CARRYB[12][42] ), .CI(\SUMB[12][43] ), 
        .CO(\CARRYB[13][42] ), .S(\SUMB[13][42] ) );
  FA_X1 S2_13_43 ( .A(\ab[13][43] ), .B(\CARRYB[12][43] ), .CI(\SUMB[12][44] ), 
        .CO(\CARRYB[13][43] ), .S(\SUMB[13][43] ) );
  FA_X1 S2_13_44 ( .A(\ab[13][44] ), .B(\CARRYB[12][44] ), .CI(\SUMB[12][45] ), 
        .CO(\CARRYB[13][44] ), .S(\SUMB[13][44] ) );
  FA_X1 S2_13_45 ( .A(\ab[13][45] ), .B(\CARRYB[12][45] ), .CI(\SUMB[12][46] ), 
        .CO(\CARRYB[13][45] ), .S(\SUMB[13][45] ) );
  FA_X1 S2_13_46 ( .A(\ab[13][46] ), .B(\CARRYB[12][46] ), .CI(\SUMB[12][47] ), 
        .CO(\CARRYB[13][46] ), .S(\SUMB[13][46] ) );
  FA_X1 S2_13_47 ( .A(\ab[13][47] ), .B(\CARRYB[12][47] ), .CI(\SUMB[12][48] ), 
        .CO(\CARRYB[13][47] ), .S(\SUMB[13][47] ) );
  FA_X1 S2_13_48 ( .A(\ab[13][48] ), .B(\CARRYB[12][48] ), .CI(\SUMB[12][49] ), 
        .CO(\CARRYB[13][48] ), .S(\SUMB[13][48] ) );
  FA_X1 S2_13_49 ( .A(\ab[13][49] ), .B(\CARRYB[12][49] ), .CI(\SUMB[12][50] ), 
        .CO(\CARRYB[13][49] ), .S(\SUMB[13][49] ) );
  FA_X1 S2_13_50 ( .A(\ab[13][50] ), .B(\CARRYB[12][50] ), .CI(\SUMB[12][51] ), 
        .CO(\CARRYB[13][50] ), .S(\SUMB[13][50] ) );
  FA_X1 S3_13_51 ( .A(\ab[13][51] ), .B(\CARRYB[12][51] ), .CI(\ab[12][52] ), 
        .CO(\CARRYB[13][51] ), .S(\SUMB[13][51] ) );
  FA_X1 S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(CLA_SUM[12]) );
  FA_X1 S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA_X1 S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA_X1 S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FA_X1 S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA_X1 S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA_X1 S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA_X1 S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA_X1 S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA_X1 S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA_X1 S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA_X1 S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), 
        .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA_X1 S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), 
        .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FA_X1 S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), 
        .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA_X1 S2_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\SUMB[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FA_X1 S2_12_15 ( .A(\ab[12][15] ), .B(\CARRYB[11][15] ), .CI(\SUMB[11][16] ), 
        .CO(\CARRYB[12][15] ), .S(\SUMB[12][15] ) );
  FA_X1 S2_12_16 ( .A(\ab[12][16] ), .B(\CARRYB[11][16] ), .CI(\SUMB[11][17] ), 
        .CO(\CARRYB[12][16] ), .S(\SUMB[12][16] ) );
  FA_X1 S2_12_17 ( .A(\ab[12][17] ), .B(\CARRYB[11][17] ), .CI(\SUMB[11][18] ), 
        .CO(\CARRYB[12][17] ), .S(\SUMB[12][17] ) );
  FA_X1 S2_12_18 ( .A(\ab[12][18] ), .B(\CARRYB[11][18] ), .CI(\SUMB[11][19] ), 
        .CO(\CARRYB[12][18] ), .S(\SUMB[12][18] ) );
  FA_X1 S2_12_19 ( .A(\ab[12][19] ), .B(\CARRYB[11][19] ), .CI(\SUMB[11][20] ), 
        .CO(\CARRYB[12][19] ), .S(\SUMB[12][19] ) );
  FA_X1 S2_12_20 ( .A(\ab[12][20] ), .B(\CARRYB[11][20] ), .CI(\SUMB[11][21] ), 
        .CO(\CARRYB[12][20] ), .S(\SUMB[12][20] ) );
  FA_X1 S2_12_21 ( .A(\ab[12][21] ), .B(\CARRYB[11][21] ), .CI(\SUMB[11][22] ), 
        .CO(\CARRYB[12][21] ), .S(\SUMB[12][21] ) );
  FA_X1 S2_12_22 ( .A(\ab[12][22] ), .B(\CARRYB[11][22] ), .CI(\SUMB[11][23] ), 
        .CO(\CARRYB[12][22] ), .S(\SUMB[12][22] ) );
  FA_X1 S2_12_23 ( .A(\ab[12][23] ), .B(\CARRYB[11][23] ), .CI(\SUMB[11][24] ), 
        .CO(\CARRYB[12][23] ), .S(\SUMB[12][23] ) );
  FA_X1 S2_12_24 ( .A(\ab[12][24] ), .B(\CARRYB[11][24] ), .CI(\SUMB[11][25] ), 
        .CO(\CARRYB[12][24] ), .S(\SUMB[12][24] ) );
  FA_X1 S2_12_25 ( .A(\ab[12][25] ), .B(\CARRYB[11][25] ), .CI(\SUMB[11][26] ), 
        .CO(\CARRYB[12][25] ), .S(\SUMB[12][25] ) );
  FA_X1 S2_12_26 ( .A(\ab[12][26] ), .B(\CARRYB[11][26] ), .CI(\SUMB[11][27] ), 
        .CO(\CARRYB[12][26] ), .S(\SUMB[12][26] ) );
  FA_X1 S2_12_27 ( .A(\ab[12][27] ), .B(\CARRYB[11][27] ), .CI(\SUMB[11][28] ), 
        .CO(\CARRYB[12][27] ), .S(\SUMB[12][27] ) );
  FA_X1 S2_12_28 ( .A(\ab[12][28] ), .B(\CARRYB[11][28] ), .CI(\SUMB[11][29] ), 
        .CO(\CARRYB[12][28] ), .S(\SUMB[12][28] ) );
  FA_X1 S2_12_29 ( .A(\ab[12][29] ), .B(\CARRYB[11][29] ), .CI(\SUMB[11][30] ), 
        .CO(\CARRYB[12][29] ), .S(\SUMB[12][29] ) );
  FA_X1 S2_12_30 ( .A(\ab[12][30] ), .B(\CARRYB[11][30] ), .CI(\SUMB[11][31] ), 
        .CO(\CARRYB[12][30] ), .S(\SUMB[12][30] ) );
  FA_X1 S2_12_31 ( .A(\ab[12][31] ), .B(\CARRYB[11][31] ), .CI(\SUMB[11][32] ), 
        .CO(\CARRYB[12][31] ), .S(\SUMB[12][31] ) );
  FA_X1 S2_12_32 ( .A(\ab[12][32] ), .B(\CARRYB[11][32] ), .CI(\SUMB[11][33] ), 
        .CO(\CARRYB[12][32] ), .S(\SUMB[12][32] ) );
  FA_X1 S2_12_33 ( .A(\ab[12][33] ), .B(\CARRYB[11][33] ), .CI(\SUMB[11][34] ), 
        .CO(\CARRYB[12][33] ), .S(\SUMB[12][33] ) );
  FA_X1 S2_12_34 ( .A(\ab[12][34] ), .B(\CARRYB[11][34] ), .CI(\SUMB[11][35] ), 
        .CO(\CARRYB[12][34] ), .S(\SUMB[12][34] ) );
  FA_X1 S2_12_35 ( .A(\ab[12][35] ), .B(\CARRYB[11][35] ), .CI(\SUMB[11][36] ), 
        .CO(\CARRYB[12][35] ), .S(\SUMB[12][35] ) );
  FA_X1 S2_12_36 ( .A(\ab[12][36] ), .B(\CARRYB[11][36] ), .CI(\SUMB[11][37] ), 
        .CO(\CARRYB[12][36] ), .S(\SUMB[12][36] ) );
  FA_X1 S2_12_37 ( .A(\ab[12][37] ), .B(\CARRYB[11][37] ), .CI(\SUMB[11][38] ), 
        .CO(\CARRYB[12][37] ), .S(\SUMB[12][37] ) );
  FA_X1 S2_12_38 ( .A(\ab[12][38] ), .B(\CARRYB[11][38] ), .CI(\SUMB[11][39] ), 
        .CO(\CARRYB[12][38] ), .S(\SUMB[12][38] ) );
  FA_X1 S2_12_39 ( .A(\ab[12][39] ), .B(\CARRYB[11][39] ), .CI(\SUMB[11][40] ), 
        .CO(\CARRYB[12][39] ), .S(\SUMB[12][39] ) );
  FA_X1 S2_12_40 ( .A(\ab[12][40] ), .B(\CARRYB[11][40] ), .CI(\SUMB[11][41] ), 
        .CO(\CARRYB[12][40] ), .S(\SUMB[12][40] ) );
  FA_X1 S2_12_41 ( .A(\ab[12][41] ), .B(\CARRYB[11][41] ), .CI(\SUMB[11][42] ), 
        .CO(\CARRYB[12][41] ), .S(\SUMB[12][41] ) );
  FA_X1 S2_12_42 ( .A(\ab[12][42] ), .B(\CARRYB[11][42] ), .CI(\SUMB[11][43] ), 
        .CO(\CARRYB[12][42] ), .S(\SUMB[12][42] ) );
  FA_X1 S2_12_43 ( .A(\ab[12][43] ), .B(\CARRYB[11][43] ), .CI(\SUMB[11][44] ), 
        .CO(\CARRYB[12][43] ), .S(\SUMB[12][43] ) );
  FA_X1 S2_12_44 ( .A(\ab[12][44] ), .B(\CARRYB[11][44] ), .CI(\SUMB[11][45] ), 
        .CO(\CARRYB[12][44] ), .S(\SUMB[12][44] ) );
  FA_X1 S2_12_45 ( .A(\ab[12][45] ), .B(\CARRYB[11][45] ), .CI(\SUMB[11][46] ), 
        .CO(\CARRYB[12][45] ), .S(\SUMB[12][45] ) );
  FA_X1 S2_12_46 ( .A(\ab[12][46] ), .B(\CARRYB[11][46] ), .CI(\SUMB[11][47] ), 
        .CO(\CARRYB[12][46] ), .S(\SUMB[12][46] ) );
  FA_X1 S2_12_47 ( .A(\ab[12][47] ), .B(\CARRYB[11][47] ), .CI(\SUMB[11][48] ), 
        .CO(\CARRYB[12][47] ), .S(\SUMB[12][47] ) );
  FA_X1 S2_12_48 ( .A(\ab[12][48] ), .B(\CARRYB[11][48] ), .CI(\SUMB[11][49] ), 
        .CO(\CARRYB[12][48] ), .S(\SUMB[12][48] ) );
  FA_X1 S2_12_49 ( .A(\ab[12][49] ), .B(\CARRYB[11][49] ), .CI(\SUMB[11][50] ), 
        .CO(\CARRYB[12][49] ), .S(\SUMB[12][49] ) );
  FA_X1 S2_12_50 ( .A(\ab[12][50] ), .B(\CARRYB[11][50] ), .CI(\SUMB[11][51] ), 
        .CO(\CARRYB[12][50] ), .S(\SUMB[12][50] ) );
  FA_X1 S3_12_51 ( .A(\ab[12][51] ), .B(\CARRYB[11][51] ), .CI(\ab[11][52] ), 
        .CO(\CARRYB[12][51] ), .S(\SUMB[12][51] ) );
  FA_X1 S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(CLA_SUM[11]) );
  FA_X1 S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA_X1 S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA_X1 S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA_X1 S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA_X1 S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA_X1 S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA_X1 S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA_X1 S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA_X1 S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA_X1 S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA_X1 S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA_X1 S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA_X1 S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA_X1 S2_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\SUMB[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA_X1 S2_11_15 ( .A(\ab[11][15] ), .B(\CARRYB[10][15] ), .CI(\SUMB[10][16] ), 
        .CO(\CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FA_X1 S2_11_16 ( .A(\ab[11][16] ), .B(\CARRYB[10][16] ), .CI(\SUMB[10][17] ), 
        .CO(\CARRYB[11][16] ), .S(\SUMB[11][16] ) );
  FA_X1 S2_11_17 ( .A(\ab[11][17] ), .B(\CARRYB[10][17] ), .CI(\SUMB[10][18] ), 
        .CO(\CARRYB[11][17] ), .S(\SUMB[11][17] ) );
  FA_X1 S2_11_18 ( .A(\ab[11][18] ), .B(\CARRYB[10][18] ), .CI(\SUMB[10][19] ), 
        .CO(\CARRYB[11][18] ), .S(\SUMB[11][18] ) );
  FA_X1 S2_11_19 ( .A(\ab[11][19] ), .B(\CARRYB[10][19] ), .CI(\SUMB[10][20] ), 
        .CO(\CARRYB[11][19] ), .S(\SUMB[11][19] ) );
  FA_X1 S2_11_20 ( .A(\ab[11][20] ), .B(\CARRYB[10][20] ), .CI(\SUMB[10][21] ), 
        .CO(\CARRYB[11][20] ), .S(\SUMB[11][20] ) );
  FA_X1 S2_11_21 ( .A(\ab[11][21] ), .B(\CARRYB[10][21] ), .CI(\SUMB[10][22] ), 
        .CO(\CARRYB[11][21] ), .S(\SUMB[11][21] ) );
  FA_X1 S2_11_22 ( .A(\ab[11][22] ), .B(\CARRYB[10][22] ), .CI(\SUMB[10][23] ), 
        .CO(\CARRYB[11][22] ), .S(\SUMB[11][22] ) );
  FA_X1 S2_11_23 ( .A(\ab[11][23] ), .B(\CARRYB[10][23] ), .CI(\SUMB[10][24] ), 
        .CO(\CARRYB[11][23] ), .S(\SUMB[11][23] ) );
  FA_X1 S2_11_24 ( .A(\ab[11][24] ), .B(\CARRYB[10][24] ), .CI(\SUMB[10][25] ), 
        .CO(\CARRYB[11][24] ), .S(\SUMB[11][24] ) );
  FA_X1 S2_11_25 ( .A(\ab[11][25] ), .B(\CARRYB[10][25] ), .CI(\SUMB[10][26] ), 
        .CO(\CARRYB[11][25] ), .S(\SUMB[11][25] ) );
  FA_X1 S2_11_26 ( .A(\ab[11][26] ), .B(\CARRYB[10][26] ), .CI(\SUMB[10][27] ), 
        .CO(\CARRYB[11][26] ), .S(\SUMB[11][26] ) );
  FA_X1 S2_11_27 ( .A(\ab[11][27] ), .B(\CARRYB[10][27] ), .CI(\SUMB[10][28] ), 
        .CO(\CARRYB[11][27] ), .S(\SUMB[11][27] ) );
  FA_X1 S2_11_28 ( .A(\ab[11][28] ), .B(\CARRYB[10][28] ), .CI(\SUMB[10][29] ), 
        .CO(\CARRYB[11][28] ), .S(\SUMB[11][28] ) );
  FA_X1 S2_11_29 ( .A(\ab[11][29] ), .B(\CARRYB[10][29] ), .CI(\SUMB[10][30] ), 
        .CO(\CARRYB[11][29] ), .S(\SUMB[11][29] ) );
  FA_X1 S2_11_30 ( .A(\ab[11][30] ), .B(\CARRYB[10][30] ), .CI(\SUMB[10][31] ), 
        .CO(\CARRYB[11][30] ), .S(\SUMB[11][30] ) );
  FA_X1 S2_11_31 ( .A(\ab[11][31] ), .B(\CARRYB[10][31] ), .CI(\SUMB[10][32] ), 
        .CO(\CARRYB[11][31] ), .S(\SUMB[11][31] ) );
  FA_X1 S2_11_32 ( .A(\ab[11][32] ), .B(\CARRYB[10][32] ), .CI(\SUMB[10][33] ), 
        .CO(\CARRYB[11][32] ), .S(\SUMB[11][32] ) );
  FA_X1 S2_11_33 ( .A(\ab[11][33] ), .B(\CARRYB[10][33] ), .CI(\SUMB[10][34] ), 
        .CO(\CARRYB[11][33] ), .S(\SUMB[11][33] ) );
  FA_X1 S2_11_34 ( .A(\ab[11][34] ), .B(\CARRYB[10][34] ), .CI(\SUMB[10][35] ), 
        .CO(\CARRYB[11][34] ), .S(\SUMB[11][34] ) );
  FA_X1 S2_11_35 ( .A(\ab[11][35] ), .B(\CARRYB[10][35] ), .CI(\SUMB[10][36] ), 
        .CO(\CARRYB[11][35] ), .S(\SUMB[11][35] ) );
  FA_X1 S2_11_36 ( .A(\ab[11][36] ), .B(\CARRYB[10][36] ), .CI(\SUMB[10][37] ), 
        .CO(\CARRYB[11][36] ), .S(\SUMB[11][36] ) );
  FA_X1 S2_11_37 ( .A(\ab[11][37] ), .B(\CARRYB[10][37] ), .CI(\SUMB[10][38] ), 
        .CO(\CARRYB[11][37] ), .S(\SUMB[11][37] ) );
  FA_X1 S2_11_38 ( .A(\ab[11][38] ), .B(\CARRYB[10][38] ), .CI(\SUMB[10][39] ), 
        .CO(\CARRYB[11][38] ), .S(\SUMB[11][38] ) );
  FA_X1 S2_11_39 ( .A(\ab[11][39] ), .B(\CARRYB[10][39] ), .CI(\SUMB[10][40] ), 
        .CO(\CARRYB[11][39] ), .S(\SUMB[11][39] ) );
  FA_X1 S2_11_40 ( .A(\ab[11][40] ), .B(\CARRYB[10][40] ), .CI(\SUMB[10][41] ), 
        .CO(\CARRYB[11][40] ), .S(\SUMB[11][40] ) );
  FA_X1 S2_11_41 ( .A(\ab[11][41] ), .B(\CARRYB[10][41] ), .CI(\SUMB[10][42] ), 
        .CO(\CARRYB[11][41] ), .S(\SUMB[11][41] ) );
  FA_X1 S2_11_42 ( .A(\ab[11][42] ), .B(\CARRYB[10][42] ), .CI(\SUMB[10][43] ), 
        .CO(\CARRYB[11][42] ), .S(\SUMB[11][42] ) );
  FA_X1 S2_11_43 ( .A(\ab[11][43] ), .B(\CARRYB[10][43] ), .CI(\SUMB[10][44] ), 
        .CO(\CARRYB[11][43] ), .S(\SUMB[11][43] ) );
  FA_X1 S2_11_44 ( .A(\ab[11][44] ), .B(\CARRYB[10][44] ), .CI(\SUMB[10][45] ), 
        .CO(\CARRYB[11][44] ), .S(\SUMB[11][44] ) );
  FA_X1 S2_11_45 ( .A(\ab[11][45] ), .B(\CARRYB[10][45] ), .CI(\SUMB[10][46] ), 
        .CO(\CARRYB[11][45] ), .S(\SUMB[11][45] ) );
  FA_X1 S2_11_46 ( .A(\ab[11][46] ), .B(\CARRYB[10][46] ), .CI(\SUMB[10][47] ), 
        .CO(\CARRYB[11][46] ), .S(\SUMB[11][46] ) );
  FA_X1 S2_11_47 ( .A(\ab[11][47] ), .B(\CARRYB[10][47] ), .CI(\SUMB[10][48] ), 
        .CO(\CARRYB[11][47] ), .S(\SUMB[11][47] ) );
  FA_X1 S2_11_48 ( .A(\ab[11][48] ), .B(\CARRYB[10][48] ), .CI(\SUMB[10][49] ), 
        .CO(\CARRYB[11][48] ), .S(\SUMB[11][48] ) );
  FA_X1 S2_11_49 ( .A(\ab[11][49] ), .B(\CARRYB[10][49] ), .CI(\SUMB[10][50] ), 
        .CO(\CARRYB[11][49] ), .S(\SUMB[11][49] ) );
  FA_X1 S2_11_50 ( .A(\ab[11][50] ), .B(\CARRYB[10][50] ), .CI(\SUMB[10][51] ), 
        .CO(\CARRYB[11][50] ), .S(\SUMB[11][50] ) );
  FA_X1 S3_11_51 ( .A(\ab[11][51] ), .B(\CARRYB[10][51] ), .CI(\ab[10][52] ), 
        .CO(\CARRYB[11][51] ), .S(\SUMB[11][51] ) );
  FA_X1 S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(CLA_SUM[10]) );
  FA_X1 S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA_X1 S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA_X1 S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA_X1 S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA_X1 S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA_X1 S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA_X1 S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA_X1 S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA_X1 S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), 
        .CO(\CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA_X1 S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA_X1 S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA_X1 S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA_X1 S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA_X1 S2_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\SUMB[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA_X1 S2_10_15 ( .A(\ab[10][15] ), .B(\CARRYB[9][15] ), .CI(\SUMB[9][16] ), 
        .CO(\CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FA_X1 S2_10_16 ( .A(\ab[10][16] ), .B(\CARRYB[9][16] ), .CI(\SUMB[9][17] ), 
        .CO(\CARRYB[10][16] ), .S(\SUMB[10][16] ) );
  FA_X1 S2_10_17 ( .A(\ab[10][17] ), .B(\CARRYB[9][17] ), .CI(\SUMB[9][18] ), 
        .CO(\CARRYB[10][17] ), .S(\SUMB[10][17] ) );
  FA_X1 S2_10_18 ( .A(\ab[10][18] ), .B(\CARRYB[9][18] ), .CI(\SUMB[9][19] ), 
        .CO(\CARRYB[10][18] ), .S(\SUMB[10][18] ) );
  FA_X1 S2_10_19 ( .A(\ab[10][19] ), .B(\CARRYB[9][19] ), .CI(\SUMB[9][20] ), 
        .CO(\CARRYB[10][19] ), .S(\SUMB[10][19] ) );
  FA_X1 S2_10_20 ( .A(\ab[10][20] ), .B(\CARRYB[9][20] ), .CI(\SUMB[9][21] ), 
        .CO(\CARRYB[10][20] ), .S(\SUMB[10][20] ) );
  FA_X1 S2_10_21 ( .A(\ab[10][21] ), .B(\CARRYB[9][21] ), .CI(\SUMB[9][22] ), 
        .CO(\CARRYB[10][21] ), .S(\SUMB[10][21] ) );
  FA_X1 S2_10_22 ( .A(\ab[10][22] ), .B(\CARRYB[9][22] ), .CI(\SUMB[9][23] ), 
        .CO(\CARRYB[10][22] ), .S(\SUMB[10][22] ) );
  FA_X1 S2_10_23 ( .A(\ab[10][23] ), .B(\CARRYB[9][23] ), .CI(\SUMB[9][24] ), 
        .CO(\CARRYB[10][23] ), .S(\SUMB[10][23] ) );
  FA_X1 S2_10_24 ( .A(\ab[10][24] ), .B(\CARRYB[9][24] ), .CI(\SUMB[9][25] ), 
        .CO(\CARRYB[10][24] ), .S(\SUMB[10][24] ) );
  FA_X1 S2_10_25 ( .A(\ab[10][25] ), .B(\CARRYB[9][25] ), .CI(\SUMB[9][26] ), 
        .CO(\CARRYB[10][25] ), .S(\SUMB[10][25] ) );
  FA_X1 S2_10_26 ( .A(\ab[10][26] ), .B(\CARRYB[9][26] ), .CI(\SUMB[9][27] ), 
        .CO(\CARRYB[10][26] ), .S(\SUMB[10][26] ) );
  FA_X1 S2_10_27 ( .A(\ab[10][27] ), .B(\CARRYB[9][27] ), .CI(\SUMB[9][28] ), 
        .CO(\CARRYB[10][27] ), .S(\SUMB[10][27] ) );
  FA_X1 S2_10_28 ( .A(\ab[10][28] ), .B(\CARRYB[9][28] ), .CI(\SUMB[9][29] ), 
        .CO(\CARRYB[10][28] ), .S(\SUMB[10][28] ) );
  FA_X1 S2_10_29 ( .A(\ab[10][29] ), .B(\CARRYB[9][29] ), .CI(\SUMB[9][30] ), 
        .CO(\CARRYB[10][29] ), .S(\SUMB[10][29] ) );
  FA_X1 S2_10_30 ( .A(\ab[10][30] ), .B(\CARRYB[9][30] ), .CI(\SUMB[9][31] ), 
        .CO(\CARRYB[10][30] ), .S(\SUMB[10][30] ) );
  FA_X1 S2_10_31 ( .A(\ab[10][31] ), .B(\CARRYB[9][31] ), .CI(\SUMB[9][32] ), 
        .CO(\CARRYB[10][31] ), .S(\SUMB[10][31] ) );
  FA_X1 S2_10_32 ( .A(\ab[10][32] ), .B(\CARRYB[9][32] ), .CI(\SUMB[9][33] ), 
        .CO(\CARRYB[10][32] ), .S(\SUMB[10][32] ) );
  FA_X1 S2_10_33 ( .A(\ab[10][33] ), .B(\CARRYB[9][33] ), .CI(\SUMB[9][34] ), 
        .CO(\CARRYB[10][33] ), .S(\SUMB[10][33] ) );
  FA_X1 S2_10_34 ( .A(\ab[10][34] ), .B(\CARRYB[9][34] ), .CI(\SUMB[9][35] ), 
        .CO(\CARRYB[10][34] ), .S(\SUMB[10][34] ) );
  FA_X1 S2_10_35 ( .A(\ab[10][35] ), .B(\CARRYB[9][35] ), .CI(\SUMB[9][36] ), 
        .CO(\CARRYB[10][35] ), .S(\SUMB[10][35] ) );
  FA_X1 S2_10_36 ( .A(\ab[10][36] ), .B(\CARRYB[9][36] ), .CI(\SUMB[9][37] ), 
        .CO(\CARRYB[10][36] ), .S(\SUMB[10][36] ) );
  FA_X1 S2_10_37 ( .A(\ab[10][37] ), .B(\CARRYB[9][37] ), .CI(\SUMB[9][38] ), 
        .CO(\CARRYB[10][37] ), .S(\SUMB[10][37] ) );
  FA_X1 S2_10_38 ( .A(\ab[10][38] ), .B(\CARRYB[9][38] ), .CI(\SUMB[9][39] ), 
        .CO(\CARRYB[10][38] ), .S(\SUMB[10][38] ) );
  FA_X1 S2_10_39 ( .A(\ab[10][39] ), .B(\CARRYB[9][39] ), .CI(\SUMB[9][40] ), 
        .CO(\CARRYB[10][39] ), .S(\SUMB[10][39] ) );
  FA_X1 S2_10_40 ( .A(\ab[10][40] ), .B(\CARRYB[9][40] ), .CI(\SUMB[9][41] ), 
        .CO(\CARRYB[10][40] ), .S(\SUMB[10][40] ) );
  FA_X1 S2_10_41 ( .A(\ab[10][41] ), .B(\CARRYB[9][41] ), .CI(\SUMB[9][42] ), 
        .CO(\CARRYB[10][41] ), .S(\SUMB[10][41] ) );
  FA_X1 S2_10_42 ( .A(\ab[10][42] ), .B(\CARRYB[9][42] ), .CI(\SUMB[9][43] ), 
        .CO(\CARRYB[10][42] ), .S(\SUMB[10][42] ) );
  FA_X1 S2_10_43 ( .A(\ab[10][43] ), .B(\CARRYB[9][43] ), .CI(\SUMB[9][44] ), 
        .CO(\CARRYB[10][43] ), .S(\SUMB[10][43] ) );
  FA_X1 S2_10_44 ( .A(\ab[10][44] ), .B(\CARRYB[9][44] ), .CI(\SUMB[9][45] ), 
        .CO(\CARRYB[10][44] ), .S(\SUMB[10][44] ) );
  FA_X1 S2_10_45 ( .A(\ab[10][45] ), .B(\CARRYB[9][45] ), .CI(\SUMB[9][46] ), 
        .CO(\CARRYB[10][45] ), .S(\SUMB[10][45] ) );
  FA_X1 S2_10_46 ( .A(\ab[10][46] ), .B(\CARRYB[9][46] ), .CI(\SUMB[9][47] ), 
        .CO(\CARRYB[10][46] ), .S(\SUMB[10][46] ) );
  FA_X1 S2_10_47 ( .A(\ab[10][47] ), .B(\CARRYB[9][47] ), .CI(\SUMB[9][48] ), 
        .CO(\CARRYB[10][47] ), .S(\SUMB[10][47] ) );
  FA_X1 S2_10_48 ( .A(\ab[10][48] ), .B(\CARRYB[9][48] ), .CI(\SUMB[9][49] ), 
        .CO(\CARRYB[10][48] ), .S(\SUMB[10][48] ) );
  FA_X1 S2_10_49 ( .A(\ab[10][49] ), .B(\CARRYB[9][49] ), .CI(\SUMB[9][50] ), 
        .CO(\CARRYB[10][49] ), .S(\SUMB[10][49] ) );
  FA_X1 S2_10_50 ( .A(\ab[10][50] ), .B(\CARRYB[9][50] ), .CI(\SUMB[9][51] ), 
        .CO(\CARRYB[10][50] ), .S(\SUMB[10][50] ) );
  FA_X1 S3_10_51 ( .A(\ab[10][51] ), .B(\CARRYB[9][51] ), .CI(\ab[9][52] ), 
        .CO(\CARRYB[10][51] ), .S(\SUMB[10][51] ) );
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  FA_X1 S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(CLA_SUM[9]) );
  FA_X1 S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA_X1 S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
<<<<<<< HEAD
  FA_X1 S2_9_3 ( .A(\CARRYB[8][3] ), .B(\ab[9][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA_X1 S2_9_4 ( .A(\CARRYB[8][4] ), .B(\ab[9][4] ), .CI(\SUMB[8][5] ), .CO(
=======
  FA_X1 S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA_X1 S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA_X1 S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA_X1 S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA_X1 S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA_X1 S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
<<<<<<< HEAD
  FA_X1 S3_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\ab[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
=======
  FA_X1 S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA_X1 S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA_X1 S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA_X1 S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA_X1 S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA_X1 S2_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\SUMB[8][15] ), 
        .CO(\CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA_X1 S2_9_15 ( .A(\ab[9][15] ), .B(\CARRYB[8][15] ), .CI(\SUMB[8][16] ), 
        .CO(\CARRYB[9][15] ), .S(\SUMB[9][15] ) );
  FA_X1 S2_9_16 ( .A(\ab[9][16] ), .B(\CARRYB[8][16] ), .CI(\SUMB[8][17] ), 
        .CO(\CARRYB[9][16] ), .S(\SUMB[9][16] ) );
  FA_X1 S2_9_17 ( .A(\ab[9][17] ), .B(\CARRYB[8][17] ), .CI(\SUMB[8][18] ), 
        .CO(\CARRYB[9][17] ), .S(\SUMB[9][17] ) );
  FA_X1 S2_9_18 ( .A(\ab[9][18] ), .B(\CARRYB[8][18] ), .CI(\SUMB[8][19] ), 
        .CO(\CARRYB[9][18] ), .S(\SUMB[9][18] ) );
  FA_X1 S2_9_19 ( .A(\ab[9][19] ), .B(\CARRYB[8][19] ), .CI(\SUMB[8][20] ), 
        .CO(\CARRYB[9][19] ), .S(\SUMB[9][19] ) );
  FA_X1 S2_9_20 ( .A(\ab[9][20] ), .B(\CARRYB[8][20] ), .CI(\SUMB[8][21] ), 
        .CO(\CARRYB[9][20] ), .S(\SUMB[9][20] ) );
  FA_X1 S2_9_21 ( .A(\ab[9][21] ), .B(\CARRYB[8][21] ), .CI(\SUMB[8][22] ), 
        .CO(\CARRYB[9][21] ), .S(\SUMB[9][21] ) );
  FA_X1 S2_9_22 ( .A(\ab[9][22] ), .B(\CARRYB[8][22] ), .CI(\SUMB[8][23] ), 
        .CO(\CARRYB[9][22] ), .S(\SUMB[9][22] ) );
  FA_X1 S2_9_23 ( .A(\ab[9][23] ), .B(\CARRYB[8][23] ), .CI(\SUMB[8][24] ), 
        .CO(\CARRYB[9][23] ), .S(\SUMB[9][23] ) );
  FA_X1 S2_9_24 ( .A(\ab[9][24] ), .B(\CARRYB[8][24] ), .CI(\SUMB[8][25] ), 
        .CO(\CARRYB[9][24] ), .S(\SUMB[9][24] ) );
  FA_X1 S2_9_25 ( .A(\ab[9][25] ), .B(\CARRYB[8][25] ), .CI(\SUMB[8][26] ), 
        .CO(\CARRYB[9][25] ), .S(\SUMB[9][25] ) );
  FA_X1 S2_9_26 ( .A(\ab[9][26] ), .B(\CARRYB[8][26] ), .CI(\SUMB[8][27] ), 
        .CO(\CARRYB[9][26] ), .S(\SUMB[9][26] ) );
  FA_X1 S2_9_27 ( .A(\ab[9][27] ), .B(\CARRYB[8][27] ), .CI(\SUMB[8][28] ), 
        .CO(\CARRYB[9][27] ), .S(\SUMB[9][27] ) );
  FA_X1 S2_9_28 ( .A(\ab[9][28] ), .B(\CARRYB[8][28] ), .CI(\SUMB[8][29] ), 
        .CO(\CARRYB[9][28] ), .S(\SUMB[9][28] ) );
  FA_X1 S2_9_29 ( .A(\ab[9][29] ), .B(\CARRYB[8][29] ), .CI(\SUMB[8][30] ), 
        .CO(\CARRYB[9][29] ), .S(\SUMB[9][29] ) );
  FA_X1 S2_9_30 ( .A(\ab[9][30] ), .B(\CARRYB[8][30] ), .CI(\SUMB[8][31] ), 
        .CO(\CARRYB[9][30] ), .S(\SUMB[9][30] ) );
  FA_X1 S2_9_31 ( .A(\ab[9][31] ), .B(\CARRYB[8][31] ), .CI(\SUMB[8][32] ), 
        .CO(\CARRYB[9][31] ), .S(\SUMB[9][31] ) );
  FA_X1 S2_9_32 ( .A(\ab[9][32] ), .B(\CARRYB[8][32] ), .CI(\SUMB[8][33] ), 
        .CO(\CARRYB[9][32] ), .S(\SUMB[9][32] ) );
  FA_X1 S2_9_33 ( .A(\ab[9][33] ), .B(\CARRYB[8][33] ), .CI(\SUMB[8][34] ), 
        .CO(\CARRYB[9][33] ), .S(\SUMB[9][33] ) );
  FA_X1 S2_9_34 ( .A(\ab[9][34] ), .B(\CARRYB[8][34] ), .CI(\SUMB[8][35] ), 
        .CO(\CARRYB[9][34] ), .S(\SUMB[9][34] ) );
  FA_X1 S2_9_35 ( .A(\ab[9][35] ), .B(\CARRYB[8][35] ), .CI(\SUMB[8][36] ), 
        .CO(\CARRYB[9][35] ), .S(\SUMB[9][35] ) );
  FA_X1 S2_9_36 ( .A(\ab[9][36] ), .B(\CARRYB[8][36] ), .CI(\SUMB[8][37] ), 
        .CO(\CARRYB[9][36] ), .S(\SUMB[9][36] ) );
  FA_X1 S2_9_37 ( .A(\ab[9][37] ), .B(\CARRYB[8][37] ), .CI(\SUMB[8][38] ), 
        .CO(\CARRYB[9][37] ), .S(\SUMB[9][37] ) );
  FA_X1 S2_9_38 ( .A(\ab[9][38] ), .B(\CARRYB[8][38] ), .CI(\SUMB[8][39] ), 
        .CO(\CARRYB[9][38] ), .S(\SUMB[9][38] ) );
  FA_X1 S2_9_39 ( .A(\ab[9][39] ), .B(\CARRYB[8][39] ), .CI(\SUMB[8][40] ), 
        .CO(\CARRYB[9][39] ), .S(\SUMB[9][39] ) );
  FA_X1 S2_9_40 ( .A(\ab[9][40] ), .B(\CARRYB[8][40] ), .CI(\SUMB[8][41] ), 
        .CO(\CARRYB[9][40] ), .S(\SUMB[9][40] ) );
  FA_X1 S2_9_41 ( .A(\ab[9][41] ), .B(\CARRYB[8][41] ), .CI(\SUMB[8][42] ), 
        .CO(\CARRYB[9][41] ), .S(\SUMB[9][41] ) );
  FA_X1 S2_9_42 ( .A(\ab[9][42] ), .B(\CARRYB[8][42] ), .CI(\SUMB[8][43] ), 
        .CO(\CARRYB[9][42] ), .S(\SUMB[9][42] ) );
  FA_X1 S2_9_43 ( .A(\ab[9][43] ), .B(\CARRYB[8][43] ), .CI(\SUMB[8][44] ), 
        .CO(\CARRYB[9][43] ), .S(\SUMB[9][43] ) );
  FA_X1 S2_9_44 ( .A(\ab[9][44] ), .B(\CARRYB[8][44] ), .CI(\SUMB[8][45] ), 
        .CO(\CARRYB[9][44] ), .S(\SUMB[9][44] ) );
  FA_X1 S2_9_45 ( .A(\ab[9][45] ), .B(\CARRYB[8][45] ), .CI(\SUMB[8][46] ), 
        .CO(\CARRYB[9][45] ), .S(\SUMB[9][45] ) );
  FA_X1 S2_9_46 ( .A(\ab[9][46] ), .B(\CARRYB[8][46] ), .CI(\SUMB[8][47] ), 
        .CO(\CARRYB[9][46] ), .S(\SUMB[9][46] ) );
  FA_X1 S2_9_47 ( .A(\ab[9][47] ), .B(\CARRYB[8][47] ), .CI(\SUMB[8][48] ), 
        .CO(\CARRYB[9][47] ), .S(\SUMB[9][47] ) );
  FA_X1 S2_9_48 ( .A(\ab[9][48] ), .B(\CARRYB[8][48] ), .CI(\SUMB[8][49] ), 
        .CO(\CARRYB[9][48] ), .S(\SUMB[9][48] ) );
  FA_X1 S2_9_49 ( .A(\ab[9][49] ), .B(\CARRYB[8][49] ), .CI(\SUMB[8][50] ), 
        .CO(\CARRYB[9][49] ), .S(\SUMB[9][49] ) );
  FA_X1 S2_9_50 ( .A(\ab[9][50] ), .B(\CARRYB[8][50] ), .CI(\SUMB[8][51] ), 
        .CO(\CARRYB[9][50] ), .S(\SUMB[9][50] ) );
  FA_X1 S3_9_51 ( .A(\ab[9][51] ), .B(\CARRYB[8][51] ), .CI(\ab[8][52] ), .CO(
        \CARRYB[9][51] ), .S(\SUMB[9][51] ) );
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  FA_X1 S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(CLA_SUM[8]) );
  FA_X1 S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA_X1 S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
<<<<<<< HEAD
  FA_X1 S2_8_3 ( .A(\CARRYB[7][3] ), .B(\ab[8][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA_X1 S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA_X1 S2_8_5 ( .A(\CARRYB[7][5] ), .B(\ab[8][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA_X1 S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA_X1 S2_8_7 ( .A(\ab[8][7] ), .B(\SUMB[7][8] ), .CI(\CARRYB[7][7] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA_X1 S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA_X1 S3_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\ab[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
=======
  FA_X1 S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA_X1 S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA_X1 S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA_X1 S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA_X1 S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA_X1 S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA_X1 S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA_X1 S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA_X1 S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA_X1 S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA_X1 S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA_X1 S2_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\SUMB[7][15] ), 
        .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA_X1 S2_8_15 ( .A(\ab[8][15] ), .B(\CARRYB[7][15] ), .CI(\SUMB[7][16] ), 
        .CO(\CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FA_X1 S2_8_16 ( .A(\ab[8][16] ), .B(\CARRYB[7][16] ), .CI(\SUMB[7][17] ), 
        .CO(\CARRYB[8][16] ), .S(\SUMB[8][16] ) );
  FA_X1 S2_8_17 ( .A(\ab[8][17] ), .B(\CARRYB[7][17] ), .CI(\SUMB[7][18] ), 
        .CO(\CARRYB[8][17] ), .S(\SUMB[8][17] ) );
  FA_X1 S2_8_18 ( .A(\ab[8][18] ), .B(\CARRYB[7][18] ), .CI(\SUMB[7][19] ), 
        .CO(\CARRYB[8][18] ), .S(\SUMB[8][18] ) );
  FA_X1 S2_8_19 ( .A(\ab[8][19] ), .B(\CARRYB[7][19] ), .CI(\SUMB[7][20] ), 
        .CO(\CARRYB[8][19] ), .S(\SUMB[8][19] ) );
  FA_X1 S2_8_20 ( .A(\ab[8][20] ), .B(\CARRYB[7][20] ), .CI(\SUMB[7][21] ), 
        .CO(\CARRYB[8][20] ), .S(\SUMB[8][20] ) );
  FA_X1 S2_8_21 ( .A(\ab[8][21] ), .B(\CARRYB[7][21] ), .CI(\SUMB[7][22] ), 
        .CO(\CARRYB[8][21] ), .S(\SUMB[8][21] ) );
  FA_X1 S2_8_22 ( .A(\ab[8][22] ), .B(\CARRYB[7][22] ), .CI(\SUMB[7][23] ), 
        .CO(\CARRYB[8][22] ), .S(\SUMB[8][22] ) );
  FA_X1 S2_8_23 ( .A(\ab[8][23] ), .B(\CARRYB[7][23] ), .CI(\SUMB[7][24] ), 
        .CO(\CARRYB[8][23] ), .S(\SUMB[8][23] ) );
  FA_X1 S2_8_24 ( .A(\ab[8][24] ), .B(\CARRYB[7][24] ), .CI(\SUMB[7][25] ), 
        .CO(\CARRYB[8][24] ), .S(\SUMB[8][24] ) );
  FA_X1 S2_8_25 ( .A(\ab[8][25] ), .B(\CARRYB[7][25] ), .CI(\SUMB[7][26] ), 
        .CO(\CARRYB[8][25] ), .S(\SUMB[8][25] ) );
  FA_X1 S2_8_26 ( .A(\ab[8][26] ), .B(\CARRYB[7][26] ), .CI(\SUMB[7][27] ), 
        .CO(\CARRYB[8][26] ), .S(\SUMB[8][26] ) );
  FA_X1 S2_8_27 ( .A(\ab[8][27] ), .B(\CARRYB[7][27] ), .CI(\SUMB[7][28] ), 
        .CO(\CARRYB[8][27] ), .S(\SUMB[8][27] ) );
  FA_X1 S2_8_28 ( .A(\ab[8][28] ), .B(\CARRYB[7][28] ), .CI(\SUMB[7][29] ), 
        .CO(\CARRYB[8][28] ), .S(\SUMB[8][28] ) );
  FA_X1 S2_8_29 ( .A(\ab[8][29] ), .B(\CARRYB[7][29] ), .CI(\SUMB[7][30] ), 
        .CO(\CARRYB[8][29] ), .S(\SUMB[8][29] ) );
  FA_X1 S2_8_30 ( .A(\ab[8][30] ), .B(\CARRYB[7][30] ), .CI(\SUMB[7][31] ), 
        .CO(\CARRYB[8][30] ), .S(\SUMB[8][30] ) );
  FA_X1 S2_8_31 ( .A(\ab[8][31] ), .B(\CARRYB[7][31] ), .CI(\SUMB[7][32] ), 
        .CO(\CARRYB[8][31] ), .S(\SUMB[8][31] ) );
  FA_X1 S2_8_32 ( .A(\ab[8][32] ), .B(\CARRYB[7][32] ), .CI(\SUMB[7][33] ), 
        .CO(\CARRYB[8][32] ), .S(\SUMB[8][32] ) );
  FA_X1 S2_8_33 ( .A(\ab[8][33] ), .B(\CARRYB[7][33] ), .CI(\SUMB[7][34] ), 
        .CO(\CARRYB[8][33] ), .S(\SUMB[8][33] ) );
  FA_X1 S2_8_34 ( .A(\ab[8][34] ), .B(\CARRYB[7][34] ), .CI(\SUMB[7][35] ), 
        .CO(\CARRYB[8][34] ), .S(\SUMB[8][34] ) );
  FA_X1 S2_8_35 ( .A(\ab[8][35] ), .B(\CARRYB[7][35] ), .CI(\SUMB[7][36] ), 
        .CO(\CARRYB[8][35] ), .S(\SUMB[8][35] ) );
  FA_X1 S2_8_36 ( .A(\ab[8][36] ), .B(\CARRYB[7][36] ), .CI(\SUMB[7][37] ), 
        .CO(\CARRYB[8][36] ), .S(\SUMB[8][36] ) );
  FA_X1 S2_8_37 ( .A(\ab[8][37] ), .B(\CARRYB[7][37] ), .CI(\SUMB[7][38] ), 
        .CO(\CARRYB[8][37] ), .S(\SUMB[8][37] ) );
  FA_X1 S2_8_38 ( .A(\ab[8][38] ), .B(\CARRYB[7][38] ), .CI(\SUMB[7][39] ), 
        .CO(\CARRYB[8][38] ), .S(\SUMB[8][38] ) );
  FA_X1 S2_8_39 ( .A(\ab[8][39] ), .B(\CARRYB[7][39] ), .CI(\SUMB[7][40] ), 
        .CO(\CARRYB[8][39] ), .S(\SUMB[8][39] ) );
  FA_X1 S2_8_40 ( .A(\ab[8][40] ), .B(\CARRYB[7][40] ), .CI(\SUMB[7][41] ), 
        .CO(\CARRYB[8][40] ), .S(\SUMB[8][40] ) );
  FA_X1 S2_8_41 ( .A(\ab[8][41] ), .B(\CARRYB[7][41] ), .CI(\SUMB[7][42] ), 
        .CO(\CARRYB[8][41] ), .S(\SUMB[8][41] ) );
  FA_X1 S2_8_42 ( .A(\ab[8][42] ), .B(\CARRYB[7][42] ), .CI(\SUMB[7][43] ), 
        .CO(\CARRYB[8][42] ), .S(\SUMB[8][42] ) );
  FA_X1 S2_8_43 ( .A(\ab[8][43] ), .B(\CARRYB[7][43] ), .CI(\SUMB[7][44] ), 
        .CO(\CARRYB[8][43] ), .S(\SUMB[8][43] ) );
  FA_X1 S2_8_44 ( .A(\ab[8][44] ), .B(\CARRYB[7][44] ), .CI(\SUMB[7][45] ), 
        .CO(\CARRYB[8][44] ), .S(\SUMB[8][44] ) );
  FA_X1 S2_8_45 ( .A(\ab[8][45] ), .B(\CARRYB[7][45] ), .CI(\SUMB[7][46] ), 
        .CO(\CARRYB[8][45] ), .S(\SUMB[8][45] ) );
  FA_X1 S2_8_46 ( .A(\ab[8][46] ), .B(\CARRYB[7][46] ), .CI(\SUMB[7][47] ), 
        .CO(\CARRYB[8][46] ), .S(\SUMB[8][46] ) );
  FA_X1 S2_8_47 ( .A(\ab[8][47] ), .B(\CARRYB[7][47] ), .CI(\SUMB[7][48] ), 
        .CO(\CARRYB[8][47] ), .S(\SUMB[8][47] ) );
  FA_X1 S2_8_48 ( .A(\ab[8][48] ), .B(\CARRYB[7][48] ), .CI(\SUMB[7][49] ), 
        .CO(\CARRYB[8][48] ), .S(\SUMB[8][48] ) );
  FA_X1 S2_8_49 ( .A(\ab[8][49] ), .B(\CARRYB[7][49] ), .CI(\SUMB[7][50] ), 
        .CO(\CARRYB[8][49] ), .S(\SUMB[8][49] ) );
  FA_X1 S2_8_50 ( .A(\ab[8][50] ), .B(\CARRYB[7][50] ), .CI(\SUMB[7][51] ), 
        .CO(\CARRYB[8][50] ), .S(\SUMB[8][50] ) );
  FA_X1 S3_8_51 ( .A(\ab[8][51] ), .B(\CARRYB[7][51] ), .CI(\ab[7][52] ), .CO(
        \CARRYB[8][51] ), .S(\SUMB[8][51] ) );
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  FA_X1 S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(CLA_SUM[7]) );
  FA_X1 S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA_X1 S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA_X1 S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA_X1 S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
<<<<<<< HEAD
  FA_X1 S2_7_5 ( .A(\CARRYB[6][5] ), .B(\ab[7][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA_X1 S2_7_6 ( .A(\CARRYB[6][6] ), .B(\ab[7][6] ), .CI(\SUMB[6][7] ), .CO(
=======
  FA_X1 S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA_X1 S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA_X1 S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA_X1 S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
<<<<<<< HEAD
  FA_X1 S3_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\ab[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
=======
  FA_X1 S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA_X1 S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA_X1 S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA_X1 S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA_X1 S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA_X1 S2_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\SUMB[6][15] ), 
        .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA_X1 S2_7_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .CI(\SUMB[6][16] ), 
        .CO(\CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FA_X1 S2_7_16 ( .A(\ab[7][16] ), .B(\CARRYB[6][16] ), .CI(\SUMB[6][17] ), 
        .CO(\CARRYB[7][16] ), .S(\SUMB[7][16] ) );
  FA_X1 S2_7_17 ( .A(\ab[7][17] ), .B(\CARRYB[6][17] ), .CI(\SUMB[6][18] ), 
        .CO(\CARRYB[7][17] ), .S(\SUMB[7][17] ) );
  FA_X1 S2_7_18 ( .A(\ab[7][18] ), .B(\CARRYB[6][18] ), .CI(\SUMB[6][19] ), 
        .CO(\CARRYB[7][18] ), .S(\SUMB[7][18] ) );
  FA_X1 S2_7_19 ( .A(\ab[7][19] ), .B(\CARRYB[6][19] ), .CI(\SUMB[6][20] ), 
        .CO(\CARRYB[7][19] ), .S(\SUMB[7][19] ) );
  FA_X1 S2_7_20 ( .A(\ab[7][20] ), .B(\CARRYB[6][20] ), .CI(\SUMB[6][21] ), 
        .CO(\CARRYB[7][20] ), .S(\SUMB[7][20] ) );
  FA_X1 S2_7_21 ( .A(\ab[7][21] ), .B(\CARRYB[6][21] ), .CI(\SUMB[6][22] ), 
        .CO(\CARRYB[7][21] ), .S(\SUMB[7][21] ) );
  FA_X1 S2_7_22 ( .A(\ab[7][22] ), .B(\CARRYB[6][22] ), .CI(\SUMB[6][23] ), 
        .CO(\CARRYB[7][22] ), .S(\SUMB[7][22] ) );
  FA_X1 S2_7_23 ( .A(\ab[7][23] ), .B(\CARRYB[6][23] ), .CI(\SUMB[6][24] ), 
        .CO(\CARRYB[7][23] ), .S(\SUMB[7][23] ) );
  FA_X1 S2_7_24 ( .A(\ab[7][24] ), .B(\CARRYB[6][24] ), .CI(\SUMB[6][25] ), 
        .CO(\CARRYB[7][24] ), .S(\SUMB[7][24] ) );
  FA_X1 S2_7_25 ( .A(\ab[7][25] ), .B(\CARRYB[6][25] ), .CI(\SUMB[6][26] ), 
        .CO(\CARRYB[7][25] ), .S(\SUMB[7][25] ) );
  FA_X1 S2_7_26 ( .A(\ab[7][26] ), .B(\CARRYB[6][26] ), .CI(\SUMB[6][27] ), 
        .CO(\CARRYB[7][26] ), .S(\SUMB[7][26] ) );
  FA_X1 S2_7_27 ( .A(\ab[7][27] ), .B(\CARRYB[6][27] ), .CI(\SUMB[6][28] ), 
        .CO(\CARRYB[7][27] ), .S(\SUMB[7][27] ) );
  FA_X1 S2_7_28 ( .A(\ab[7][28] ), .B(\CARRYB[6][28] ), .CI(\SUMB[6][29] ), 
        .CO(\CARRYB[7][28] ), .S(\SUMB[7][28] ) );
  FA_X1 S2_7_29 ( .A(\ab[7][29] ), .B(\CARRYB[6][29] ), .CI(\SUMB[6][30] ), 
        .CO(\CARRYB[7][29] ), .S(\SUMB[7][29] ) );
  FA_X1 S2_7_30 ( .A(\ab[7][30] ), .B(\CARRYB[6][30] ), .CI(\SUMB[6][31] ), 
        .CO(\CARRYB[7][30] ), .S(\SUMB[7][30] ) );
  FA_X1 S2_7_31 ( .A(\ab[7][31] ), .B(\CARRYB[6][31] ), .CI(\SUMB[6][32] ), 
        .CO(\CARRYB[7][31] ), .S(\SUMB[7][31] ) );
  FA_X1 S2_7_32 ( .A(\ab[7][32] ), .B(\CARRYB[6][32] ), .CI(\SUMB[6][33] ), 
        .CO(\CARRYB[7][32] ), .S(\SUMB[7][32] ) );
  FA_X1 S2_7_33 ( .A(\ab[7][33] ), .B(\CARRYB[6][33] ), .CI(\SUMB[6][34] ), 
        .CO(\CARRYB[7][33] ), .S(\SUMB[7][33] ) );
  FA_X1 S2_7_34 ( .A(\ab[7][34] ), .B(\CARRYB[6][34] ), .CI(\SUMB[6][35] ), 
        .CO(\CARRYB[7][34] ), .S(\SUMB[7][34] ) );
  FA_X1 S2_7_35 ( .A(\ab[7][35] ), .B(\CARRYB[6][35] ), .CI(\SUMB[6][36] ), 
        .CO(\CARRYB[7][35] ), .S(\SUMB[7][35] ) );
  FA_X1 S2_7_36 ( .A(\ab[7][36] ), .B(\CARRYB[6][36] ), .CI(\SUMB[6][37] ), 
        .CO(\CARRYB[7][36] ), .S(\SUMB[7][36] ) );
  FA_X1 S2_7_37 ( .A(\ab[7][37] ), .B(\CARRYB[6][37] ), .CI(\SUMB[6][38] ), 
        .CO(\CARRYB[7][37] ), .S(\SUMB[7][37] ) );
  FA_X1 S2_7_38 ( .A(\ab[7][38] ), .B(\CARRYB[6][38] ), .CI(\SUMB[6][39] ), 
        .CO(\CARRYB[7][38] ), .S(\SUMB[7][38] ) );
  FA_X1 S2_7_39 ( .A(\ab[7][39] ), .B(\CARRYB[6][39] ), .CI(\SUMB[6][40] ), 
        .CO(\CARRYB[7][39] ), .S(\SUMB[7][39] ) );
  FA_X1 S2_7_40 ( .A(\ab[7][40] ), .B(\CARRYB[6][40] ), .CI(\SUMB[6][41] ), 
        .CO(\CARRYB[7][40] ), .S(\SUMB[7][40] ) );
  FA_X1 S2_7_41 ( .A(\ab[7][41] ), .B(\CARRYB[6][41] ), .CI(\SUMB[6][42] ), 
        .CO(\CARRYB[7][41] ), .S(\SUMB[7][41] ) );
  FA_X1 S2_7_42 ( .A(\ab[7][42] ), .B(\CARRYB[6][42] ), .CI(\SUMB[6][43] ), 
        .CO(\CARRYB[7][42] ), .S(\SUMB[7][42] ) );
  FA_X1 S2_7_43 ( .A(\ab[7][43] ), .B(\CARRYB[6][43] ), .CI(\SUMB[6][44] ), 
        .CO(\CARRYB[7][43] ), .S(\SUMB[7][43] ) );
  FA_X1 S2_7_44 ( .A(\ab[7][44] ), .B(\CARRYB[6][44] ), .CI(\SUMB[6][45] ), 
        .CO(\CARRYB[7][44] ), .S(\SUMB[7][44] ) );
  FA_X1 S2_7_45 ( .A(\ab[7][45] ), .B(\CARRYB[6][45] ), .CI(\SUMB[6][46] ), 
        .CO(\CARRYB[7][45] ), .S(\SUMB[7][45] ) );
  FA_X1 S2_7_46 ( .A(\ab[7][46] ), .B(\CARRYB[6][46] ), .CI(\SUMB[6][47] ), 
        .CO(\CARRYB[7][46] ), .S(\SUMB[7][46] ) );
  FA_X1 S2_7_47 ( .A(\ab[7][47] ), .B(\CARRYB[6][47] ), .CI(\SUMB[6][48] ), 
        .CO(\CARRYB[7][47] ), .S(\SUMB[7][47] ) );
  FA_X1 S2_7_48 ( .A(\ab[7][48] ), .B(\CARRYB[6][48] ), .CI(\SUMB[6][49] ), 
        .CO(\CARRYB[7][48] ), .S(\SUMB[7][48] ) );
  FA_X1 S2_7_49 ( .A(\ab[7][49] ), .B(\CARRYB[6][49] ), .CI(\SUMB[6][50] ), 
        .CO(\CARRYB[7][49] ), .S(\SUMB[7][49] ) );
  FA_X1 S2_7_50 ( .A(\ab[7][50] ), .B(\CARRYB[6][50] ), .CI(\SUMB[6][51] ), 
        .CO(\CARRYB[7][50] ), .S(\SUMB[7][50] ) );
  FA_X1 S3_7_51 ( .A(\ab[7][51] ), .B(\CARRYB[6][51] ), .CI(\ab[6][52] ), .CO(
        \CARRYB[7][51] ), .S(\SUMB[7][51] ) );
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  FA_X1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(CLA_SUM[6]) );
  FA_X1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA_X1 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA_X1 S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA_X1 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
<<<<<<< HEAD
  FA_X1 S2_6_5 ( .A(\CARRYB[5][5] ), .B(\ab[6][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA_X1 S2_6_6 ( .A(\CARRYB[5][6] ), .B(\ab[6][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA_X1 S2_6_7 ( .A(\ab[6][7] ), .B(\SUMB[5][8] ), .CI(\CARRYB[5][7] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA_X1 S2_6_8 ( .A(\CARRYB[5][8] ), .B(\ab[6][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA_X1 S3_6_9 ( .A(\ab[6][9] ), .B(\ab[5][10] ), .CI(\CARRYB[5][9] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
=======
  FA_X1 S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA_X1 S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA_X1 S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA_X1 S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA_X1 S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA_X1 S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA_X1 S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA_X1 S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA_X1 S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA_X1 S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\SUMB[5][15] ), 
        .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA_X1 S2_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .CI(\SUMB[5][16] ), 
        .CO(\CARRYB[6][15] ), .S(\SUMB[6][15] ) );
  FA_X1 S2_6_16 ( .A(\ab[6][16] ), .B(\CARRYB[5][16] ), .CI(\SUMB[5][17] ), 
        .CO(\CARRYB[6][16] ), .S(\SUMB[6][16] ) );
  FA_X1 S2_6_17 ( .A(\ab[6][17] ), .B(\CARRYB[5][17] ), .CI(\SUMB[5][18] ), 
        .CO(\CARRYB[6][17] ), .S(\SUMB[6][17] ) );
  FA_X1 S2_6_18 ( .A(\ab[6][18] ), .B(\CARRYB[5][18] ), .CI(\SUMB[5][19] ), 
        .CO(\CARRYB[6][18] ), .S(\SUMB[6][18] ) );
  FA_X1 S2_6_19 ( .A(\ab[6][19] ), .B(\CARRYB[5][19] ), .CI(\SUMB[5][20] ), 
        .CO(\CARRYB[6][19] ), .S(\SUMB[6][19] ) );
  FA_X1 S2_6_20 ( .A(\ab[6][20] ), .B(\CARRYB[5][20] ), .CI(\SUMB[5][21] ), 
        .CO(\CARRYB[6][20] ), .S(\SUMB[6][20] ) );
  FA_X1 S2_6_21 ( .A(\ab[6][21] ), .B(\CARRYB[5][21] ), .CI(\SUMB[5][22] ), 
        .CO(\CARRYB[6][21] ), .S(\SUMB[6][21] ) );
  FA_X1 S2_6_22 ( .A(\ab[6][22] ), .B(\CARRYB[5][22] ), .CI(\SUMB[5][23] ), 
        .CO(\CARRYB[6][22] ), .S(\SUMB[6][22] ) );
  FA_X1 S2_6_23 ( .A(\ab[6][23] ), .B(\CARRYB[5][23] ), .CI(\SUMB[5][24] ), 
        .CO(\CARRYB[6][23] ), .S(\SUMB[6][23] ) );
  FA_X1 S2_6_24 ( .A(\ab[6][24] ), .B(\CARRYB[5][24] ), .CI(\SUMB[5][25] ), 
        .CO(\CARRYB[6][24] ), .S(\SUMB[6][24] ) );
  FA_X1 S2_6_25 ( .A(\ab[6][25] ), .B(\CARRYB[5][25] ), .CI(\SUMB[5][26] ), 
        .CO(\CARRYB[6][25] ), .S(\SUMB[6][25] ) );
  FA_X1 S2_6_26 ( .A(\ab[6][26] ), .B(\CARRYB[5][26] ), .CI(\SUMB[5][27] ), 
        .CO(\CARRYB[6][26] ), .S(\SUMB[6][26] ) );
  FA_X1 S2_6_27 ( .A(\ab[6][27] ), .B(\CARRYB[5][27] ), .CI(\SUMB[5][28] ), 
        .CO(\CARRYB[6][27] ), .S(\SUMB[6][27] ) );
  FA_X1 S2_6_28 ( .A(\ab[6][28] ), .B(\CARRYB[5][28] ), .CI(\SUMB[5][29] ), 
        .CO(\CARRYB[6][28] ), .S(\SUMB[6][28] ) );
  FA_X1 S2_6_29 ( .A(\ab[6][29] ), .B(\CARRYB[5][29] ), .CI(\SUMB[5][30] ), 
        .CO(\CARRYB[6][29] ), .S(\SUMB[6][29] ) );
  FA_X1 S2_6_30 ( .A(\ab[6][30] ), .B(\CARRYB[5][30] ), .CI(\SUMB[5][31] ), 
        .CO(\CARRYB[6][30] ), .S(\SUMB[6][30] ) );
  FA_X1 S2_6_31 ( .A(\ab[6][31] ), .B(\CARRYB[5][31] ), .CI(\SUMB[5][32] ), 
        .CO(\CARRYB[6][31] ), .S(\SUMB[6][31] ) );
  FA_X1 S2_6_32 ( .A(\ab[6][32] ), .B(\CARRYB[5][32] ), .CI(\SUMB[5][33] ), 
        .CO(\CARRYB[6][32] ), .S(\SUMB[6][32] ) );
  FA_X1 S2_6_33 ( .A(\ab[6][33] ), .B(\CARRYB[5][33] ), .CI(\SUMB[5][34] ), 
        .CO(\CARRYB[6][33] ), .S(\SUMB[6][33] ) );
  FA_X1 S2_6_34 ( .A(\ab[6][34] ), .B(\CARRYB[5][34] ), .CI(\SUMB[5][35] ), 
        .CO(\CARRYB[6][34] ), .S(\SUMB[6][34] ) );
  FA_X1 S2_6_35 ( .A(\ab[6][35] ), .B(\CARRYB[5][35] ), .CI(\SUMB[5][36] ), 
        .CO(\CARRYB[6][35] ), .S(\SUMB[6][35] ) );
  FA_X1 S2_6_36 ( .A(\ab[6][36] ), .B(\CARRYB[5][36] ), .CI(\SUMB[5][37] ), 
        .CO(\CARRYB[6][36] ), .S(\SUMB[6][36] ) );
  FA_X1 S2_6_37 ( .A(\ab[6][37] ), .B(\CARRYB[5][37] ), .CI(\SUMB[5][38] ), 
        .CO(\CARRYB[6][37] ), .S(\SUMB[6][37] ) );
  FA_X1 S2_6_38 ( .A(\ab[6][38] ), .B(\CARRYB[5][38] ), .CI(\SUMB[5][39] ), 
        .CO(\CARRYB[6][38] ), .S(\SUMB[6][38] ) );
  FA_X1 S2_6_39 ( .A(\ab[6][39] ), .B(\CARRYB[5][39] ), .CI(\SUMB[5][40] ), 
        .CO(\CARRYB[6][39] ), .S(\SUMB[6][39] ) );
  FA_X1 S2_6_40 ( .A(\ab[6][40] ), .B(\CARRYB[5][40] ), .CI(\SUMB[5][41] ), 
        .CO(\CARRYB[6][40] ), .S(\SUMB[6][40] ) );
  FA_X1 S2_6_41 ( .A(\ab[6][41] ), .B(\CARRYB[5][41] ), .CI(\SUMB[5][42] ), 
        .CO(\CARRYB[6][41] ), .S(\SUMB[6][41] ) );
  FA_X1 S2_6_42 ( .A(\ab[6][42] ), .B(\CARRYB[5][42] ), .CI(\SUMB[5][43] ), 
        .CO(\CARRYB[6][42] ), .S(\SUMB[6][42] ) );
  FA_X1 S2_6_43 ( .A(\ab[6][43] ), .B(\CARRYB[5][43] ), .CI(\SUMB[5][44] ), 
        .CO(\CARRYB[6][43] ), .S(\SUMB[6][43] ) );
  FA_X1 S2_6_44 ( .A(\ab[6][44] ), .B(\CARRYB[5][44] ), .CI(\SUMB[5][45] ), 
        .CO(\CARRYB[6][44] ), .S(\SUMB[6][44] ) );
  FA_X1 S2_6_45 ( .A(\ab[6][45] ), .B(\CARRYB[5][45] ), .CI(\SUMB[5][46] ), 
        .CO(\CARRYB[6][45] ), .S(\SUMB[6][45] ) );
  FA_X1 S2_6_46 ( .A(\ab[6][46] ), .B(\CARRYB[5][46] ), .CI(\SUMB[5][47] ), 
        .CO(\CARRYB[6][46] ), .S(\SUMB[6][46] ) );
  FA_X1 S2_6_47 ( .A(\ab[6][47] ), .B(\CARRYB[5][47] ), .CI(\SUMB[5][48] ), 
        .CO(\CARRYB[6][47] ), .S(\SUMB[6][47] ) );
  FA_X1 S2_6_48 ( .A(\ab[6][48] ), .B(\CARRYB[5][48] ), .CI(\SUMB[5][49] ), 
        .CO(\CARRYB[6][48] ), .S(\SUMB[6][48] ) );
  FA_X1 S2_6_49 ( .A(\ab[6][49] ), .B(\CARRYB[5][49] ), .CI(\SUMB[5][50] ), 
        .CO(\CARRYB[6][49] ), .S(\SUMB[6][49] ) );
  FA_X1 S2_6_50 ( .A(\ab[6][50] ), .B(\CARRYB[5][50] ), .CI(\SUMB[5][51] ), 
        .CO(\CARRYB[6][50] ), .S(\SUMB[6][50] ) );
  FA_X1 S3_6_51 ( .A(\ab[6][51] ), .B(\CARRYB[5][51] ), .CI(\ab[5][52] ), .CO(
        \CARRYB[6][51] ), .S(\SUMB[6][51] ) );
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  FA_X1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(CLA_SUM[5]) );
  FA_X1 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA_X1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA_X1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA_X1 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA_X1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
<<<<<<< HEAD
  FA_X1 S2_5_6 ( .A(\CARRYB[4][6] ), .B(\ab[5][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA_X1 S2_5_7 ( .A(\CARRYB[4][7] ), .B(\ab[5][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA_X1 S2_5_8 ( .A(\CARRYB[4][8] ), .B(\ab[5][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA_X1 S3_5_9 ( .A(\ab[5][9] ), .B(\ab[4][10] ), .CI(\CARRYB[4][9] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
=======
  FA_X1 S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA_X1 S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA_X1 S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA_X1 S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA_X1 S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA_X1 S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA_X1 S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA_X1 S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA_X1 S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\SUMB[4][15] ), 
        .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA_X1 S2_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .CI(\SUMB[4][16] ), 
        .CO(\CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FA_X1 S2_5_16 ( .A(\ab[5][16] ), .B(\CARRYB[4][16] ), .CI(\SUMB[4][17] ), 
        .CO(\CARRYB[5][16] ), .S(\SUMB[5][16] ) );
  FA_X1 S2_5_17 ( .A(\ab[5][17] ), .B(\CARRYB[4][17] ), .CI(\SUMB[4][18] ), 
        .CO(\CARRYB[5][17] ), .S(\SUMB[5][17] ) );
  FA_X1 S2_5_18 ( .A(\ab[5][18] ), .B(\CARRYB[4][18] ), .CI(\SUMB[4][19] ), 
        .CO(\CARRYB[5][18] ), .S(\SUMB[5][18] ) );
  FA_X1 S2_5_19 ( .A(\ab[5][19] ), .B(\CARRYB[4][19] ), .CI(\SUMB[4][20] ), 
        .CO(\CARRYB[5][19] ), .S(\SUMB[5][19] ) );
  FA_X1 S2_5_20 ( .A(\ab[5][20] ), .B(\CARRYB[4][20] ), .CI(\SUMB[4][21] ), 
        .CO(\CARRYB[5][20] ), .S(\SUMB[5][20] ) );
  FA_X1 S2_5_21 ( .A(\ab[5][21] ), .B(\CARRYB[4][21] ), .CI(\SUMB[4][22] ), 
        .CO(\CARRYB[5][21] ), .S(\SUMB[5][21] ) );
  FA_X1 S2_5_22 ( .A(\ab[5][22] ), .B(\CARRYB[4][22] ), .CI(\SUMB[4][23] ), 
        .CO(\CARRYB[5][22] ), .S(\SUMB[5][22] ) );
  FA_X1 S2_5_23 ( .A(\ab[5][23] ), .B(\CARRYB[4][23] ), .CI(\SUMB[4][24] ), 
        .CO(\CARRYB[5][23] ), .S(\SUMB[5][23] ) );
  FA_X1 S2_5_24 ( .A(\ab[5][24] ), .B(\CARRYB[4][24] ), .CI(\SUMB[4][25] ), 
        .CO(\CARRYB[5][24] ), .S(\SUMB[5][24] ) );
  FA_X1 S2_5_25 ( .A(\ab[5][25] ), .B(\CARRYB[4][25] ), .CI(\SUMB[4][26] ), 
        .CO(\CARRYB[5][25] ), .S(\SUMB[5][25] ) );
  FA_X1 S2_5_26 ( .A(\ab[5][26] ), .B(\CARRYB[4][26] ), .CI(\SUMB[4][27] ), 
        .CO(\CARRYB[5][26] ), .S(\SUMB[5][26] ) );
  FA_X1 S2_5_27 ( .A(\ab[5][27] ), .B(\CARRYB[4][27] ), .CI(\SUMB[4][28] ), 
        .CO(\CARRYB[5][27] ), .S(\SUMB[5][27] ) );
  FA_X1 S2_5_28 ( .A(\ab[5][28] ), .B(\CARRYB[4][28] ), .CI(\SUMB[4][29] ), 
        .CO(\CARRYB[5][28] ), .S(\SUMB[5][28] ) );
  FA_X1 S2_5_29 ( .A(\ab[5][29] ), .B(\CARRYB[4][29] ), .CI(\SUMB[4][30] ), 
        .CO(\CARRYB[5][29] ), .S(\SUMB[5][29] ) );
  FA_X1 S2_5_30 ( .A(\ab[5][30] ), .B(\CARRYB[4][30] ), .CI(\SUMB[4][31] ), 
        .CO(\CARRYB[5][30] ), .S(\SUMB[5][30] ) );
  FA_X1 S2_5_31 ( .A(\ab[5][31] ), .B(\CARRYB[4][31] ), .CI(\SUMB[4][32] ), 
        .CO(\CARRYB[5][31] ), .S(\SUMB[5][31] ) );
  FA_X1 S2_5_32 ( .A(\ab[5][32] ), .B(\CARRYB[4][32] ), .CI(\SUMB[4][33] ), 
        .CO(\CARRYB[5][32] ), .S(\SUMB[5][32] ) );
  FA_X1 S2_5_33 ( .A(\ab[5][33] ), .B(\CARRYB[4][33] ), .CI(\SUMB[4][34] ), 
        .CO(\CARRYB[5][33] ), .S(\SUMB[5][33] ) );
  FA_X1 S2_5_34 ( .A(\ab[5][34] ), .B(\CARRYB[4][34] ), .CI(\SUMB[4][35] ), 
        .CO(\CARRYB[5][34] ), .S(\SUMB[5][34] ) );
  FA_X1 S2_5_35 ( .A(\ab[5][35] ), .B(\CARRYB[4][35] ), .CI(\SUMB[4][36] ), 
        .CO(\CARRYB[5][35] ), .S(\SUMB[5][35] ) );
  FA_X1 S2_5_36 ( .A(\ab[5][36] ), .B(\CARRYB[4][36] ), .CI(\SUMB[4][37] ), 
        .CO(\CARRYB[5][36] ), .S(\SUMB[5][36] ) );
  FA_X1 S2_5_37 ( .A(\ab[5][37] ), .B(\CARRYB[4][37] ), .CI(\SUMB[4][38] ), 
        .CO(\CARRYB[5][37] ), .S(\SUMB[5][37] ) );
  FA_X1 S2_5_38 ( .A(\ab[5][38] ), .B(\CARRYB[4][38] ), .CI(\SUMB[4][39] ), 
        .CO(\CARRYB[5][38] ), .S(\SUMB[5][38] ) );
  FA_X1 S2_5_39 ( .A(\ab[5][39] ), .B(\CARRYB[4][39] ), .CI(\SUMB[4][40] ), 
        .CO(\CARRYB[5][39] ), .S(\SUMB[5][39] ) );
  FA_X1 S2_5_40 ( .A(\ab[5][40] ), .B(\CARRYB[4][40] ), .CI(\SUMB[4][41] ), 
        .CO(\CARRYB[5][40] ), .S(\SUMB[5][40] ) );
  FA_X1 S2_5_41 ( .A(\ab[5][41] ), .B(\CARRYB[4][41] ), .CI(\SUMB[4][42] ), 
        .CO(\CARRYB[5][41] ), .S(\SUMB[5][41] ) );
  FA_X1 S2_5_42 ( .A(\ab[5][42] ), .B(\CARRYB[4][42] ), .CI(\SUMB[4][43] ), 
        .CO(\CARRYB[5][42] ), .S(\SUMB[5][42] ) );
  FA_X1 S2_5_43 ( .A(\ab[5][43] ), .B(\CARRYB[4][43] ), .CI(\SUMB[4][44] ), 
        .CO(\CARRYB[5][43] ), .S(\SUMB[5][43] ) );
  FA_X1 S2_5_44 ( .A(\ab[5][44] ), .B(\CARRYB[4][44] ), .CI(\SUMB[4][45] ), 
        .CO(\CARRYB[5][44] ), .S(\SUMB[5][44] ) );
  FA_X1 S2_5_45 ( .A(\ab[5][45] ), .B(\CARRYB[4][45] ), .CI(\SUMB[4][46] ), 
        .CO(\CARRYB[5][45] ), .S(\SUMB[5][45] ) );
  FA_X1 S2_5_46 ( .A(\ab[5][46] ), .B(\CARRYB[4][46] ), .CI(\SUMB[4][47] ), 
        .CO(\CARRYB[5][46] ), .S(\SUMB[5][46] ) );
  FA_X1 S2_5_47 ( .A(\ab[5][47] ), .B(\CARRYB[4][47] ), .CI(\SUMB[4][48] ), 
        .CO(\CARRYB[5][47] ), .S(\SUMB[5][47] ) );
  FA_X1 S2_5_48 ( .A(\ab[5][48] ), .B(\CARRYB[4][48] ), .CI(\SUMB[4][49] ), 
        .CO(\CARRYB[5][48] ), .S(\SUMB[5][48] ) );
  FA_X1 S2_5_49 ( .A(\ab[5][49] ), .B(\CARRYB[4][49] ), .CI(\SUMB[4][50] ), 
        .CO(\CARRYB[5][49] ), .S(\SUMB[5][49] ) );
  FA_X1 S2_5_50 ( .A(\ab[5][50] ), .B(\CARRYB[4][50] ), .CI(\SUMB[4][51] ), 
        .CO(\CARRYB[5][50] ), .S(\SUMB[5][50] ) );
  FA_X1 S3_5_51 ( .A(\ab[5][51] ), .B(\CARRYB[4][51] ), .CI(\ab[4][52] ), .CO(
        \CARRYB[5][51] ), .S(\SUMB[5][51] ) );
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  FA_X1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(CLA_SUM[4]) );
  FA_X1 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA_X1 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA_X1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA_X1 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA_X1 S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA_X1 S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA_X1 S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
<<<<<<< HEAD
  FA_X1 S2_4_8 ( .A(\SUMB[3][9] ), .B(\ab[4][8] ), .CI(\CARRYB[3][8] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA_X1 S3_4_9 ( .A(\ab[4][9] ), .B(\ab[3][10] ), .CI(\CARRYB[3][9] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
=======
  FA_X1 S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA_X1 S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA_X1 S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA_X1 S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA_X1 S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA_X1 S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA_X1 S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), 
        .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA_X1 S2_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .CI(\SUMB[3][16] ), 
        .CO(\CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FA_X1 S2_4_16 ( .A(\ab[4][16] ), .B(\CARRYB[3][16] ), .CI(\SUMB[3][17] ), 
        .CO(\CARRYB[4][16] ), .S(\SUMB[4][16] ) );
  FA_X1 S2_4_17 ( .A(\ab[4][17] ), .B(\CARRYB[3][17] ), .CI(\SUMB[3][18] ), 
        .CO(\CARRYB[4][17] ), .S(\SUMB[4][17] ) );
  FA_X1 S2_4_18 ( .A(\ab[4][18] ), .B(\CARRYB[3][18] ), .CI(\SUMB[3][19] ), 
        .CO(\CARRYB[4][18] ), .S(\SUMB[4][18] ) );
  FA_X1 S2_4_19 ( .A(\ab[4][19] ), .B(\CARRYB[3][19] ), .CI(\SUMB[3][20] ), 
        .CO(\CARRYB[4][19] ), .S(\SUMB[4][19] ) );
  FA_X1 S2_4_20 ( .A(\ab[4][20] ), .B(\CARRYB[3][20] ), .CI(\SUMB[3][21] ), 
        .CO(\CARRYB[4][20] ), .S(\SUMB[4][20] ) );
  FA_X1 S2_4_21 ( .A(\ab[4][21] ), .B(\CARRYB[3][21] ), .CI(\SUMB[3][22] ), 
        .CO(\CARRYB[4][21] ), .S(\SUMB[4][21] ) );
  FA_X1 S2_4_22 ( .A(\ab[4][22] ), .B(\CARRYB[3][22] ), .CI(\SUMB[3][23] ), 
        .CO(\CARRYB[4][22] ), .S(\SUMB[4][22] ) );
  FA_X1 S2_4_23 ( .A(\ab[4][23] ), .B(\CARRYB[3][23] ), .CI(\SUMB[3][24] ), 
        .CO(\CARRYB[4][23] ), .S(\SUMB[4][23] ) );
  FA_X1 S2_4_24 ( .A(\ab[4][24] ), .B(\CARRYB[3][24] ), .CI(\SUMB[3][25] ), 
        .CO(\CARRYB[4][24] ), .S(\SUMB[4][24] ) );
  FA_X1 S2_4_25 ( .A(\ab[4][25] ), .B(\CARRYB[3][25] ), .CI(\SUMB[3][26] ), 
        .CO(\CARRYB[4][25] ), .S(\SUMB[4][25] ) );
  FA_X1 S2_4_26 ( .A(\ab[4][26] ), .B(\CARRYB[3][26] ), .CI(\SUMB[3][27] ), 
        .CO(\CARRYB[4][26] ), .S(\SUMB[4][26] ) );
  FA_X1 S2_4_27 ( .A(\ab[4][27] ), .B(\CARRYB[3][27] ), .CI(\SUMB[3][28] ), 
        .CO(\CARRYB[4][27] ), .S(\SUMB[4][27] ) );
  FA_X1 S2_4_28 ( .A(\ab[4][28] ), .B(\CARRYB[3][28] ), .CI(\SUMB[3][29] ), 
        .CO(\CARRYB[4][28] ), .S(\SUMB[4][28] ) );
  FA_X1 S2_4_29 ( .A(\ab[4][29] ), .B(\CARRYB[3][29] ), .CI(\SUMB[3][30] ), 
        .CO(\CARRYB[4][29] ), .S(\SUMB[4][29] ) );
  FA_X1 S2_4_30 ( .A(\ab[4][30] ), .B(\CARRYB[3][30] ), .CI(\SUMB[3][31] ), 
        .CO(\CARRYB[4][30] ), .S(\SUMB[4][30] ) );
  FA_X1 S2_4_31 ( .A(\ab[4][31] ), .B(\CARRYB[3][31] ), .CI(\SUMB[3][32] ), 
        .CO(\CARRYB[4][31] ), .S(\SUMB[4][31] ) );
  FA_X1 S2_4_32 ( .A(\ab[4][32] ), .B(\CARRYB[3][32] ), .CI(\SUMB[3][33] ), 
        .CO(\CARRYB[4][32] ), .S(\SUMB[4][32] ) );
  FA_X1 S2_4_33 ( .A(\ab[4][33] ), .B(\CARRYB[3][33] ), .CI(\SUMB[3][34] ), 
        .CO(\CARRYB[4][33] ), .S(\SUMB[4][33] ) );
  FA_X1 S2_4_34 ( .A(\ab[4][34] ), .B(\CARRYB[3][34] ), .CI(\SUMB[3][35] ), 
        .CO(\CARRYB[4][34] ), .S(\SUMB[4][34] ) );
  FA_X1 S2_4_35 ( .A(\ab[4][35] ), .B(\CARRYB[3][35] ), .CI(\SUMB[3][36] ), 
        .CO(\CARRYB[4][35] ), .S(\SUMB[4][35] ) );
  FA_X1 S2_4_36 ( .A(\ab[4][36] ), .B(\CARRYB[3][36] ), .CI(\SUMB[3][37] ), 
        .CO(\CARRYB[4][36] ), .S(\SUMB[4][36] ) );
  FA_X1 S2_4_37 ( .A(\ab[4][37] ), .B(\CARRYB[3][37] ), .CI(\SUMB[3][38] ), 
        .CO(\CARRYB[4][37] ), .S(\SUMB[4][37] ) );
  FA_X1 S2_4_38 ( .A(\ab[4][38] ), .B(\CARRYB[3][38] ), .CI(\SUMB[3][39] ), 
        .CO(\CARRYB[4][38] ), .S(\SUMB[4][38] ) );
  FA_X1 S2_4_39 ( .A(\ab[4][39] ), .B(\CARRYB[3][39] ), .CI(\SUMB[3][40] ), 
        .CO(\CARRYB[4][39] ), .S(\SUMB[4][39] ) );
  FA_X1 S2_4_40 ( .A(\ab[4][40] ), .B(\CARRYB[3][40] ), .CI(\SUMB[3][41] ), 
        .CO(\CARRYB[4][40] ), .S(\SUMB[4][40] ) );
  FA_X1 S2_4_41 ( .A(\ab[4][41] ), .B(\CARRYB[3][41] ), .CI(\SUMB[3][42] ), 
        .CO(\CARRYB[4][41] ), .S(\SUMB[4][41] ) );
  FA_X1 S2_4_42 ( .A(\ab[4][42] ), .B(\CARRYB[3][42] ), .CI(\SUMB[3][43] ), 
        .CO(\CARRYB[4][42] ), .S(\SUMB[4][42] ) );
  FA_X1 S2_4_43 ( .A(\ab[4][43] ), .B(\CARRYB[3][43] ), .CI(\SUMB[3][44] ), 
        .CO(\CARRYB[4][43] ), .S(\SUMB[4][43] ) );
  FA_X1 S2_4_44 ( .A(\ab[4][44] ), .B(\CARRYB[3][44] ), .CI(\SUMB[3][45] ), 
        .CO(\CARRYB[4][44] ), .S(\SUMB[4][44] ) );
  FA_X1 S2_4_45 ( .A(\ab[4][45] ), .B(\CARRYB[3][45] ), .CI(\SUMB[3][46] ), 
        .CO(\CARRYB[4][45] ), .S(\SUMB[4][45] ) );
  FA_X1 S2_4_46 ( .A(\ab[4][46] ), .B(\CARRYB[3][46] ), .CI(\SUMB[3][47] ), 
        .CO(\CARRYB[4][46] ), .S(\SUMB[4][46] ) );
  FA_X1 S2_4_47 ( .A(\ab[4][47] ), .B(\CARRYB[3][47] ), .CI(\SUMB[3][48] ), 
        .CO(\CARRYB[4][47] ), .S(\SUMB[4][47] ) );
  FA_X1 S2_4_48 ( .A(\ab[4][48] ), .B(\CARRYB[3][48] ), .CI(\SUMB[3][49] ), 
        .CO(\CARRYB[4][48] ), .S(\SUMB[4][48] ) );
  FA_X1 S2_4_49 ( .A(\ab[4][49] ), .B(\CARRYB[3][49] ), .CI(\SUMB[3][50] ), 
        .CO(\CARRYB[4][49] ), .S(\SUMB[4][49] ) );
  FA_X1 S2_4_50 ( .A(\ab[4][50] ), .B(\CARRYB[3][50] ), .CI(\SUMB[3][51] ), 
        .CO(\CARRYB[4][50] ), .S(\SUMB[4][50] ) );
  FA_X1 S3_4_51 ( .A(\ab[4][51] ), .B(\CARRYB[3][51] ), .CI(\ab[3][52] ), .CO(
        \CARRYB[4][51] ), .S(\SUMB[4][51] ) );
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  FA_X1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(CLA_SUM[3]) );
  FA_X1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA_X1 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA_X1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA_X1 S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA_X1 S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA_X1 S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA_X1 S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
<<<<<<< HEAD
  FA_X1 S2_3_8 ( .A(\CARRYB[2][8] ), .B(\ab[3][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA_X1 S3_3_9 ( .A(\ab[3][9] ), .B(\ab[2][10] ), .CI(\CARRYB[2][9] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA_X1 S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(CLA_SUM[2]) );
  FA_X1 S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FA_X1 S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FA_X1 S2_2_3 ( .A(\ab[2][3] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FA_X1 S2_2_4 ( .A(\ab[2][4] ), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FA_X1 S2_2_5 ( .A(\ab[2][5] ), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FA_X1 S2_2_6 ( .A(\ab[2][6] ), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FA_X1 S2_2_7 ( .A(\ab[2][7] ), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FA_X1 S2_2_8 ( .A(\ab[2][8] ), .B(\CARRYB[1][8] ), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FA_X1 S3_2_9 ( .A(\CARRYB[1][9] ), .B(\ab[2][9] ), .CI(\ab[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  fpu_DW01_add_11 FS_1 ( .A({1'b0, n8, CLA_SUM[19:11], \SUMB[10][0] , 
        CLA_SUM[9:2]}), .B({n12, CLA_CARRY, n9, n5, n6, n10, n7, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM(
        PRODUCT[21:2]) );
  INV_X1 U2 ( .A(n56), .ZN(n3) );
  INV_X4 U3 ( .A(n3), .ZN(n4) );
  INV_X8 U4 ( .A(B[8]), .ZN(n56) );
  NOR2_X2 U5 ( .A1(n55), .A2(n53), .ZN(\ab[6][9] ) );
  INV_X16 U6 ( .A(B[9]), .ZN(n55) );
  NAND2_X4 U7 ( .A1(\ab[0][9] ), .A2(\ab[1][8] ), .ZN(n44) );
  NOR2_X1 U8 ( .A1(n61), .A2(n54), .ZN(\ab[7][3] ) );
  INV_X8 U9 ( .A(B[2]), .ZN(n62) );
  NOR2_X1 U10 ( .A1(n63), .A2(n54), .ZN(\ab[7][1] ) );
  INV_X8 U11 ( .A(B[0]), .ZN(n65) );
  NOR2_X1 U12 ( .A1(n59), .A2(n50), .ZN(\ab[3][5] ) );
  INV_X8 U13 ( .A(B[4]), .ZN(n60) );
  NOR2_X1 U14 ( .A1(n61), .A2(n52), .ZN(\ab[5][3] ) );
  NOR2_X1 U15 ( .A1(n69), .A2(n61), .ZN(\ab[8][3] ) );
  NOR2_X1 U16 ( .A1(n69), .A2(n62), .ZN(\ab[8][2] ) );
  INV_X8 U17 ( .A(B[1]), .ZN(n63) );
  NOR2_X1 U18 ( .A1(n69), .A2(n65), .ZN(\ab[8][0] ) );
  NOR2_X2 U19 ( .A1(n57), .A2(n52), .ZN(\ab[5][7] ) );
  NOR2_X2 U20 ( .A1(n58), .A2(n52), .ZN(\ab[5][6] ) );
  NOR2_X2 U21 ( .A1(n59), .A2(n52), .ZN(\ab[5][5] ) );
  NOR2_X1 U22 ( .A1(n69), .A2(n4), .ZN(\ab[8][8] ) );
  NOR2_X2 U23 ( .A1(n69), .A2(n57), .ZN(\ab[8][7] ) );
  NOR2_X2 U24 ( .A1(n69), .A2(n58), .ZN(\ab[8][6] ) );
  NOR2_X2 U25 ( .A1(n69), .A2(n59), .ZN(\ab[8][5] ) );
  NOR2_X1 U26 ( .A1(n60), .A2(n51), .ZN(\ab[4][4] ) );
  INV_X8 U27 ( .A(B[7]), .ZN(n57) );
  INV_X8 U28 ( .A(B[6]), .ZN(n58) );
  INV_X8 U29 ( .A(B[5]), .ZN(n59) );
  NOR2_X1 U30 ( .A1(n69), .A2(n60), .ZN(\ab[8][4] ) );
  NOR2_X1 U31 ( .A1(n61), .A2(n51), .ZN(\ab[4][3] ) );
  NOR2_X1 U32 ( .A1(n68), .A2(n62), .ZN(\ab[9][2] ) );
  NOR2_X1 U33 ( .A1(n62), .A2(n51), .ZN(\ab[4][2] ) );
  NOR2_X1 U34 ( .A1(n69), .A2(n63), .ZN(\ab[8][1] ) );
  NOR2_X1 U35 ( .A1(n63), .A2(n51), .ZN(\ab[4][1] ) );
  NOR2_X1 U36 ( .A1(n65), .A2(n54), .ZN(\ab[7][0] ) );
  NOR2_X1 U37 ( .A1(n65), .A2(n51), .ZN(\ab[4][0] ) );
  NOR2_X1 U38 ( .A1(n57), .A2(n50), .ZN(\ab[3][7] ) );
  NOR2_X1 U39 ( .A1(n57), .A2(n53), .ZN(\ab[6][7] ) );
  NOR2_X1 U40 ( .A1(n58), .A2(n53), .ZN(\ab[6][6] ) );
  NOR2_X1 U41 ( .A1(n58), .A2(n50), .ZN(\ab[3][6] ) );
  NOR2_X1 U42 ( .A1(n59), .A2(n53), .ZN(\ab[6][5] ) );
  NOR2_X1 U43 ( .A1(n68), .A2(n4), .ZN(\ab[9][8] ) );
  NOR2_X1 U44 ( .A1(n68), .A2(n57), .ZN(\ab[9][7] ) );
  NOR2_X1 U45 ( .A1(n68), .A2(n58), .ZN(\ab[9][6] ) );
  NOR2_X1 U46 ( .A1(n68), .A2(n59), .ZN(\ab[9][5] ) );
  NOR2_X1 U47 ( .A1(n68), .A2(n60), .ZN(\ab[9][4] ) );
  NOR2_X1 U48 ( .A1(n60), .A2(n52), .ZN(\ab[5][4] ) );
  NOR2_X1 U49 ( .A1(n68), .A2(n61), .ZN(\ab[9][3] ) );
  NOR2_X1 U50 ( .A1(n61), .A2(n50), .ZN(\ab[3][3] ) );
  NOR2_X1 U51 ( .A1(n62), .A2(n54), .ZN(\ab[7][2] ) );
  NOR2_X1 U52 ( .A1(n62), .A2(n50), .ZN(\ab[3][2] ) );
  NOR2_X1 U53 ( .A1(n67), .A2(n63), .ZN(\ab[10][1] ) );
  INV_X4 U54 ( .A(A[9]), .ZN(n68) );
  NOR2_X1 U55 ( .A1(n63), .A2(n53), .ZN(\ab[6][1] ) );
  NOR2_X1 U56 ( .A1(n63), .A2(n50), .ZN(\ab[3][1] ) );
  INV_X8 U57 ( .A(A[2]), .ZN(n49) );
  NOR2_X1 U58 ( .A1(n67), .A2(n65), .ZN(\ab[10][0] ) );
  NOR2_X1 U59 ( .A1(n65), .A2(n53), .ZN(\ab[6][0] ) );
  NOR2_X1 U60 ( .A1(n65), .A2(n50), .ZN(\ab[3][0] ) );
  NOR2_X1 U61 ( .A1(n57), .A2(n51), .ZN(\ab[4][7] ) );
  NOR2_X1 U62 ( .A1(n58), .A2(n51), .ZN(\ab[4][6] ) );
  NOR2_X1 U63 ( .A1(n57), .A2(n54), .ZN(\ab[7][7] ) );
  NOR2_X1 U64 ( .A1(n58), .A2(n54), .ZN(\ab[7][6] ) );
  NOR2_X1 U65 ( .A1(n59), .A2(n54), .ZN(\ab[7][5] ) );
  NOR2_X1 U66 ( .A1(n59), .A2(n51), .ZN(\ab[4][5] ) );
  NOR2_X1 U67 ( .A1(n60), .A2(n54), .ZN(\ab[7][4] ) );
  NOR2_X1 U68 ( .A1(n60), .A2(n50), .ZN(\ab[3][4] ) );
  INV_X4 U69 ( .A(B[10]), .ZN(n64) );
  NOR2_X1 U70 ( .A1(n67), .A2(n4), .ZN(\ab[10][8] ) );
  NOR2_X1 U71 ( .A1(n67), .A2(n57), .ZN(\ab[10][7] ) );
  NOR2_X1 U72 ( .A1(n67), .A2(n58), .ZN(\ab[10][6] ) );
  NOR2_X1 U73 ( .A1(n67), .A2(n59), .ZN(\ab[10][5] ) );
  NOR2_X1 U74 ( .A1(n67), .A2(n60), .ZN(\ab[10][4] ) );
  NOR2_X1 U75 ( .A1(n67), .A2(n61), .ZN(\ab[10][3] ) );
  NOR2_X1 U76 ( .A1(n61), .A2(n53), .ZN(\ab[6][3] ) );
  NOR2_X1 U77 ( .A1(n67), .A2(n62), .ZN(\ab[10][2] ) );
  NOR2_X1 U78 ( .A1(n62), .A2(n52), .ZN(\ab[5][2] ) );
  INV_X4 U79 ( .A(A[8]), .ZN(n69) );
  INV_X1 U80 ( .A(A[10]), .ZN(n67) );
  NOR2_X1 U81 ( .A1(n68), .A2(n63), .ZN(\ab[9][1] ) );
  INV_X8 U82 ( .A(A[7]), .ZN(n54) );
  NOR2_X1 U83 ( .A1(n63), .A2(n52), .ZN(\ab[5][1] ) );
  NOR2_X1 U84 ( .A1(n68), .A2(n65), .ZN(\ab[9][0] ) );
  NOR2_X1 U85 ( .A1(n65), .A2(n52), .ZN(\ab[5][0] ) );
  NOR2_X1 U86 ( .A1(n65), .A2(n49), .ZN(\ab[2][0] ) );
  AND2_X4 U87 ( .A1(\SUMB[10][4] ), .A2(\CARRYB[10][3] ), .ZN(n5) );
  AND2_X4 U88 ( .A1(\CARRYB[10][2] ), .A2(\SUMB[10][3] ), .ZN(n6) );
  AND2_X4 U89 ( .A1(\SUMB[10][1] ), .A2(\CARRYB[10][0] ), .ZN(n7) );
  XOR2_X2 U90 ( .A(\CARRYB[10][9] ), .B(\ab[10][10] ), .Z(n8) );
  AND2_X4 U91 ( .A1(\SUMB[10][5] ), .A2(\CARRYB[10][4] ), .ZN(n9) );
  AND2_X4 U92 ( .A1(\SUMB[10][2] ), .A2(\CARRYB[10][1] ), .ZN(n10) );
  XOR2_X1 U93 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Z(PRODUCT[1]) );
  AND2_X2 U94 ( .A1(\ab[10][10] ), .A2(\CARRYB[10][9] ), .ZN(n12) );
  NOR2_X2 U95 ( .A1(n58), .A2(n48), .ZN(\ab[1][6] ) );
  NOR2_X1 U96 ( .A1(n66), .A2(n65), .ZN(PRODUCT[0]) );
  NOR2_X2 U97 ( .A1(n55), .A2(n51), .ZN(\ab[4][9] ) );
  NOR2_X2 U98 ( .A1(n55), .A2(n52), .ZN(\ab[5][9] ) );
  NOR2_X2 U99 ( .A1(n66), .A2(n56), .ZN(\ab[0][8] ) );
  NOR2_X2 U100 ( .A1(n66), .A2(n58), .ZN(\ab[0][6] ) );
  NOR2_X2 U101 ( .A1(n57), .A2(n48), .ZN(\ab[1][7] ) );
  NOR2_X2 U102 ( .A1(n57), .A2(n49), .ZN(\ab[2][7] ) );
  NOR2_X2 U103 ( .A1(n14), .A2(n49), .ZN(\ab[2][10] ) );
  NOR2_X2 U104 ( .A1(n58), .A2(n49), .ZN(\ab[2][6] ) );
  NOR2_X2 U105 ( .A1(n59), .A2(n49), .ZN(\ab[2][5] ) );
  NOR2_X2 U106 ( .A1(n60), .A2(n49), .ZN(\ab[2][4] ) );
  NOR2_X2 U107 ( .A1(n61), .A2(n49), .ZN(\ab[2][3] ) );
  NOR2_X2 U108 ( .A1(n62), .A2(n49), .ZN(\ab[2][2] ) );
  NOR2_X2 U109 ( .A1(n63), .A2(n49), .ZN(\ab[2][1] ) );
  INV_X2 U110 ( .A(n16), .ZN(CLA_SUM[11]) );
  NOR2_X4 U111 ( .A1(n14), .A2(n48), .ZN(\ab[1][10] ) );
  NOR2_X1 U112 ( .A1(n67), .A2(n55), .ZN(\ab[10][9] ) );
  NOR2_X1 U113 ( .A1(n55), .A2(n50), .ZN(\ab[3][9] ) );
  NOR2_X1 U114 ( .A1(n55), .A2(n49), .ZN(\ab[2][9] ) );
  NOR2_X2 U115 ( .A1(n66), .A2(n57), .ZN(\ab[0][7] ) );
  NOR2_X2 U116 ( .A1(n66), .A2(n60), .ZN(\ab[0][4] ) );
  NOR2_X2 U117 ( .A1(n66), .A2(n59), .ZN(\ab[0][5] ) );
  NOR2_X2 U118 ( .A1(n66), .A2(n61), .ZN(\ab[0][3] ) );
  NOR2_X2 U119 ( .A1(n66), .A2(n62), .ZN(\ab[0][2] ) );
  NOR2_X2 U120 ( .A1(n66), .A2(n63), .ZN(\ab[0][1] ) );
  NOR2_X2 U121 ( .A1(n56), .A2(n49), .ZN(\ab[2][8] ) );
  NOR2_X2 U122 ( .A1(n56), .A2(n50), .ZN(\ab[3][8] ) );
  NOR2_X2 U123 ( .A1(n56), .A2(n51), .ZN(\ab[4][8] ) );
  NOR2_X2 U124 ( .A1(n56), .A2(n52), .ZN(\ab[5][8] ) );
  NOR2_X2 U125 ( .A1(n56), .A2(n53), .ZN(\ab[6][8] ) );
  NOR2_X1 U126 ( .A1(n4), .A2(n54), .ZN(\ab[7][8] ) );
  INV_X8 U127 ( .A(n13), .ZN(n14) );
  INV_X2 U128 ( .A(n64), .ZN(n13) );
  NOR2_X1 U129 ( .A1(n55), .A2(n54), .ZN(\ab[7][9] ) );
  NOR2_X1 U130 ( .A1(n69), .A2(n55), .ZN(\ab[8][9] ) );
  NOR2_X1 U131 ( .A1(n68), .A2(n55), .ZN(\ab[9][9] ) );
  NOR2_X1 U132 ( .A1(n65), .A2(n48), .ZN(\ab[1][0] ) );
  NOR2_X1 U133 ( .A1(n63), .A2(n48), .ZN(\ab[1][1] ) );
  NOR2_X1 U134 ( .A1(n62), .A2(n48), .ZN(\ab[1][2] ) );
  NOR2_X1 U135 ( .A1(n61), .A2(n48), .ZN(\ab[1][3] ) );
  NOR2_X1 U136 ( .A1(n60), .A2(n48), .ZN(\ab[1][4] ) );
  NOR2_X1 U137 ( .A1(n59), .A2(n48), .ZN(\ab[1][5] ) );
  NOR2_X1 U138 ( .A1(n67), .A2(n14), .ZN(\ab[10][10] ) );
  NOR2_X1 U139 ( .A1(n68), .A2(n14), .ZN(\ab[9][10] ) );
  NOR2_X1 U140 ( .A1(n69), .A2(n14), .ZN(\ab[8][10] ) );
  NOR2_X1 U141 ( .A1(n14), .A2(n54), .ZN(\ab[7][10] ) );
  NOR2_X1 U142 ( .A1(n14), .A2(n53), .ZN(\ab[6][10] ) );
  NOR2_X1 U143 ( .A1(n14), .A2(n52), .ZN(\ab[5][10] ) );
  NOR2_X1 U144 ( .A1(n14), .A2(n51), .ZN(\ab[4][10] ) );
  NOR2_X1 U145 ( .A1(n14), .A2(n50), .ZN(\ab[3][10] ) );
  NOR2_X4 U146 ( .A1(n64), .A2(n66), .ZN(n15) );
  XNOR2_X1 U147 ( .A(\SUMB[10][1] ), .B(\CARRYB[10][0] ), .ZN(n16) );
  INV_X8 U148 ( .A(n17), .ZN(CLA_SUM[12]) );
  XNOR2_X2 U149 ( .A(\SUMB[10][3] ), .B(\CARRYB[10][2] ), .ZN(n18) );
  XNOR2_X2 U150 ( .A(\SUMB[10][2] ), .B(\CARRYB[10][1] ), .ZN(n17) );
  INV_X4 U151 ( .A(n18), .ZN(CLA_SUM[13]) );
  XNOR2_X2 U152 ( .A(\SUMB[10][4] ), .B(\CARRYB[10][3] ), .ZN(n19) );
  INV_X4 U153 ( .A(n19), .ZN(CLA_SUM[14]) );
  XNOR2_X2 U154 ( .A(\SUMB[10][5] ), .B(\CARRYB[10][4] ), .ZN(n20) );
  INV_X4 U155 ( .A(n20), .ZN(CLA_SUM[15]) );
  NAND2_X2 U156 ( .A1(\SUMB[10][6] ), .A2(\CARRYB[10][5] ), .ZN(n21) );
  INV_X4 U157 ( .A(n21), .ZN(CLA_CARRY[16]) );
  XNOR2_X2 U158 ( .A(\CARRYB[10][5] ), .B(\SUMB[10][6] ), .ZN(n22) );
  INV_X4 U159 ( .A(n22), .ZN(CLA_SUM[16]) );
  NAND2_X2 U160 ( .A1(\SUMB[10][7] ), .A2(\CARRYB[10][6] ), .ZN(n23) );
  INV_X4 U161 ( .A(n23), .ZN(CLA_CARRY[17]) );
  XNOR2_X2 U162 ( .A(\CARRYB[10][6] ), .B(\SUMB[10][7] ), .ZN(n24) );
  INV_X4 U163 ( .A(n24), .ZN(CLA_SUM[17]) );
  NAND2_X2 U164 ( .A1(\SUMB[10][8] ), .A2(\CARRYB[10][7] ), .ZN(n25) );
  INV_X4 U165 ( .A(n25), .ZN(CLA_CARRY[18]) );
  XNOR2_X2 U166 ( .A(\CARRYB[10][7] ), .B(\SUMB[10][8] ), .ZN(n26) );
  INV_X4 U167 ( .A(n26), .ZN(CLA_SUM[18]) );
  NAND2_X2 U168 ( .A1(\SUMB[10][9] ), .A2(\CARRYB[10][8] ), .ZN(n27) );
  INV_X4 U169 ( .A(n27), .ZN(CLA_CARRY[19]) );
  XNOR2_X2 U170 ( .A(\CARRYB[10][8] ), .B(\SUMB[10][9] ), .ZN(n28) );
  INV_X4 U171 ( .A(n28), .ZN(CLA_SUM[19]) );
  NAND2_X2 U172 ( .A1(\ab[0][1] ), .A2(\ab[1][0] ), .ZN(n29) );
  INV_X4 U173 ( .A(n29), .ZN(\CARRYB[1][0] ) );
  NAND2_X2 U174 ( .A1(\ab[0][2] ), .A2(\ab[1][1] ), .ZN(n30) );
  INV_X4 U175 ( .A(n30), .ZN(\CARRYB[1][1] ) );
  XNOR2_X2 U176 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .ZN(n31) );
  INV_X4 U177 ( .A(n31), .ZN(\SUMB[1][1] ) );
  NAND2_X2 U178 ( .A1(\ab[0][3] ), .A2(\ab[1][2] ), .ZN(n32) );
  INV_X4 U179 ( .A(n32), .ZN(\CARRYB[1][2] ) );
  XNOR2_X2 U180 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .ZN(n33) );
  INV_X4 U181 ( .A(n33), .ZN(\SUMB[1][2] ) );
  NAND2_X2 U182 ( .A1(\ab[0][4] ), .A2(\ab[1][3] ), .ZN(n34) );
  INV_X4 U183 ( .A(n34), .ZN(\CARRYB[1][3] ) );
  XNOR2_X2 U184 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .ZN(n35) );
  INV_X4 U185 ( .A(n35), .ZN(\SUMB[1][3] ) );
  NAND2_X2 U186 ( .A1(\ab[0][5] ), .A2(\ab[1][4] ), .ZN(n36) );
  INV_X4 U187 ( .A(n36), .ZN(\CARRYB[1][4] ) );
  XNOR2_X2 U188 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .ZN(n37) );
  INV_X4 U189 ( .A(n37), .ZN(\SUMB[1][4] ) );
  NAND2_X2 U190 ( .A1(\ab[0][6] ), .A2(\ab[1][5] ), .ZN(n38) );
  INV_X4 U191 ( .A(n38), .ZN(\CARRYB[1][5] ) );
  XNOR2_X2 U192 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .ZN(n39) );
  INV_X4 U193 ( .A(n39), .ZN(\SUMB[1][5] ) );
  NAND2_X2 U194 ( .A1(\ab[0][7] ), .A2(\ab[1][6] ), .ZN(n40) );
  INV_X4 U195 ( .A(n40), .ZN(\CARRYB[1][6] ) );
  XNOR2_X2 U196 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .ZN(n41) );
  INV_X4 U197 ( .A(n41), .ZN(\SUMB[1][6] ) );
  NAND2_X2 U198 ( .A1(\ab[0][8] ), .A2(\ab[1][7] ), .ZN(n42) );
  INV_X4 U199 ( .A(n42), .ZN(\CARRYB[1][7] ) );
  XNOR2_X2 U200 ( .A(\ab[0][8] ), .B(\ab[1][7] ), .ZN(n43) );
  INV_X4 U201 ( .A(n43), .ZN(\SUMB[1][7] ) );
  INV_X4 U202 ( .A(n44), .ZN(\CARRYB[1][8] ) );
  XNOR2_X2 U203 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .ZN(n45) );
  INV_X4 U204 ( .A(n45), .ZN(\SUMB[1][8] ) );
  NAND2_X2 U205 ( .A1(n15), .A2(\ab[1][9] ), .ZN(n46) );
  INV_X4 U206 ( .A(n46), .ZN(\CARRYB[1][9] ) );
  XNOR2_X2 U207 ( .A(n15), .B(\ab[1][9] ), .ZN(n47) );
  INV_X4 U208 ( .A(n47), .ZN(\SUMB[1][9] ) );
  INV_X16 U209 ( .A(A[0]), .ZN(n66) );
  INV_X16 U210 ( .A(A[1]), .ZN(n48) );
  INV_X16 U211 ( .A(B[3]), .ZN(n61) );
  INV_X16 U212 ( .A(A[3]), .ZN(n50) );
  INV_X16 U213 ( .A(A[4]), .ZN(n51) );
  INV_X16 U214 ( .A(A[5]), .ZN(n52) );
  INV_X16 U215 ( .A(A[6]), .ZN(n53) );
  NOR2_X4 U216 ( .A1(n55), .A2(n48), .ZN(\ab[1][9] ) );
  NOR2_X4 U217 ( .A1(n66), .A2(n55), .ZN(\ab[0][9] ) );
  NOR2_X4 U218 ( .A1(n56), .A2(n48), .ZN(\ab[1][8] ) );
  NOR2_X4 U219 ( .A1(n60), .A2(n53), .ZN(\ab[6][4] ) );
  NOR2_X4 U220 ( .A1(n62), .A2(n53), .ZN(\ab[6][2] ) );
endmodule


module fpu_DW01_inc_5 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  XOR2_X1 U2 ( .A(n4), .B(A[1]), .Z(SUM[1]) );
  NAND3_X4 U3 ( .A1(A[8]), .A2(A[7]), .A3(A[9]), .ZN(n30) );
  AND3_X4 U4 ( .A1(A[4]), .A2(A[5]), .A3(n11), .ZN(n2) );
  INV_X1 U5 ( .A(A[0]), .ZN(n3) );
  INV_X4 U6 ( .A(n3), .ZN(n4) );
  NAND4_X1 U7 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(n19) );
  INV_X4 U8 ( .A(n4), .ZN(SUM[0]) );
  NAND2_X4 U9 ( .A1(A[4]), .A2(A[3]), .ZN(n29) );
  INV_X2 U10 ( .A(A[3]), .ZN(n22) );
  NAND2_X1 U11 ( .A1(n2), .A2(A[6]), .ZN(n15) );
  INV_X1 U12 ( .A(A[6]), .ZN(n16) );
  NAND2_X4 U13 ( .A1(n26), .A2(n27), .ZN(n25) );
  NOR2_X4 U14 ( .A1(n28), .A2(n29), .ZN(n27) );
  INV_X8 U15 ( .A(n25), .ZN(SUM[10]) );
  CLKBUF_X2 U16 ( .A(A[2]), .Z(n5) );
  INV_X2 U17 ( .A(A[4]), .ZN(n20) );
  INV_X1 U18 ( .A(A[9]), .ZN(n7) );
  XNOR2_X1 U19 ( .A(A[7]), .B(n15), .ZN(SUM[7]) );
  NOR2_X2 U20 ( .A1(n23), .A2(n24), .ZN(n21) );
  INV_X1 U21 ( .A(A[8]), .ZN(n9) );
  NAND3_X2 U22 ( .A1(A[0]), .A2(A[2]), .A3(A[1]), .ZN(n28) );
  NOR2_X2 U23 ( .A1(n13), .A2(n14), .ZN(n12) );
  NOR2_X2 U24 ( .A1(n8), .A2(n9), .ZN(n6) );
  INV_X1 U25 ( .A(A[5]), .ZN(n18) );
  NAND2_X1 U26 ( .A1(A[6]), .A2(A[5]), .ZN(n31) );
  NAND2_X1 U27 ( .A1(A[7]), .A2(A[6]), .ZN(n13) );
  NOR2_X1 U28 ( .A1(n19), .A2(n20), .ZN(n17) );
  NAND2_X1 U29 ( .A1(A[4]), .A2(A[5]), .ZN(n14) );
  NAND2_X1 U30 ( .A1(A[1]), .A2(n4), .ZN(n24) );
  NOR2_X2 U31 ( .A1(n30), .A2(n31), .ZN(n26) );
  XNOR2_X2 U32 ( .A(n6), .B(n7), .ZN(SUM[9]) );
  XNOR2_X2 U33 ( .A(n10), .B(n9), .ZN(SUM[8]) );
  INV_X4 U34 ( .A(n8), .ZN(n10) );
  NAND2_X2 U35 ( .A1(n11), .A2(n12), .ZN(n8) );
  XNOR2_X2 U36 ( .A(n2), .B(n16), .ZN(SUM[6]) );
  XNOR2_X2 U37 ( .A(n17), .B(n18), .ZN(SUM[5]) );
  XNOR2_X2 U38 ( .A(n11), .B(n20), .ZN(SUM[4]) );
  INV_X4 U39 ( .A(n19), .ZN(n11) );
  XNOR2_X2 U40 ( .A(n21), .B(n22), .ZN(SUM[3]) );
  INV_X4 U41 ( .A(A[2]), .ZN(n23) );
  XNOR2_X2 U42 ( .A(n5), .B(n24), .ZN(SUM[2]) );
endmodule


module fpu_DW_rash_2 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [2:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   n2, n3, n4, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170;

  OAI211_X2 U3 ( .C1(SH[2]), .C2(n152), .A(1'b1), .B(n153), .ZN(B[10]) );
  OAI211_X2 U4 ( .C1(SH[2]), .C2(n138), .A(1'b1), .B(n139), .ZN(B[11]) );
  OAI211_X2 U5 ( .C1(n132), .C2(SH[2]), .A(1'b1), .B(n133), .ZN(B[12]) );
  NAND2_X2 U6 ( .A1(n118), .A2(n119), .ZN(B[13]) );
  OAI21_X4 U7 ( .B1(n94), .B2(n112), .A(n113), .ZN(B[14]) );
  OAI211_X2 U8 ( .C1(n94), .C2(n106), .A(1'b1), .B(n107), .ZN(B[15]) );
  OAI211_X2 U9 ( .C1(SH[2]), .C2(n96), .A(1'b1), .B(n97), .ZN(B[16]) );
  OAI211_X2 U10 ( .C1(n74), .C2(n94), .A(1'b1), .B(n95), .ZN(B[17]) );
  NAND2_X2 U11 ( .A1(n79), .A2(n80), .ZN(B[1]) );
  INV_X4 U12 ( .A(n76), .ZN(B[20]) );
  INV_X4 U13 ( .A(n72), .ZN(B[21]) );
  NAND2_X2 U14 ( .A1(n65), .A2(n66), .ZN(B[2]) );
  NAND2_X2 U15 ( .A1(n55), .A2(n56), .ZN(B[3]) );
  AOI21_X1 U16 ( .B1(A[19]), .B2(n20), .A(n105), .ZN(n135) );
  AOI21_X1 U17 ( .B1(A[15]), .B2(n20), .A(n2), .ZN(n100) );
  AND2_X2 U18 ( .A1(n92), .A2(n25), .ZN(B[18]) );
  INV_X4 U19 ( .A(SH[1]), .ZN(n19) );
  INV_X4 U20 ( .A(SH[0]), .ZN(n22) );
  INV_X4 U21 ( .A(n17), .ZN(n16) );
  AND2_X2 U22 ( .A1(A[14]), .A2(n22), .ZN(n2) );
  AND2_X2 U23 ( .A1(A[16]), .A2(n54), .ZN(n3) );
  AND2_X2 U24 ( .A1(A[10]), .A2(n22), .ZN(n4) );
  AND2_X2 U25 ( .A1(n90), .A2(n25), .ZN(B[19]) );
  NAND2_X1 U26 ( .A1(A[7]), .A2(n84), .ZN(n159) );
  NAND2_X1 U27 ( .A1(A[7]), .A2(n15), .ZN(n146) );
  INV_X1 U28 ( .A(A[4]), .ZN(n71) );
  NAND2_X1 U29 ( .A1(A[4]), .A2(n14), .ZN(n169) );
  NAND2_X1 U30 ( .A1(A[14]), .A2(n54), .ZN(n156) );
  NAND2_X1 U31 ( .A1(A[14]), .A2(n84), .ZN(n121) );
  NAND2_X1 U32 ( .A1(A[18]), .A2(n14), .ZN(n116) );
  NAND2_X1 U33 ( .A1(A[18]), .A2(n84), .ZN(n125) );
  NAND2_X1 U34 ( .A1(A[18]), .A2(n22), .ZN(n136) );
  INV_X4 U35 ( .A(SH[2]), .ZN(n94) );
  NAND2_X2 U36 ( .A1(n49), .A2(n50), .ZN(B[4]) );
  NAND2_X2 U37 ( .A1(n46), .A2(n47), .ZN(B[5]) );
  NAND2_X2 U38 ( .A1(n41), .A2(n42), .ZN(B[6]) );
  NAND2_X2 U39 ( .A1(n36), .A2(n37), .ZN(B[7]) );
  NAND2_X2 U40 ( .A1(n30), .A2(n31), .ZN(B[8]) );
  NAND2_X2 U41 ( .A1(n23), .A2(n24), .ZN(B[9]) );
  NAND2_X2 U42 ( .A1(n98), .A2(n99), .ZN(n77) );
  NAND2_X2 U49 ( .A1(n54), .A2(n12), .ZN(n74) );
  INV_X4 U50 ( .A(n17), .ZN(n12) );
  NOR2_X4 U51 ( .A1(n21), .A2(n13), .ZN(n111) );
  INV_X4 U52 ( .A(n16), .ZN(n13) );
  NAND2_X1 U53 ( .A1(A[19]), .A2(n84), .ZN(n115) );
  NAND2_X1 U54 ( .A1(A[19]), .A2(n15), .ZN(n110) );
  NAND2_X1 U55 ( .A1(A[6]), .A2(n15), .ZN(n160) );
  NAND2_X1 U56 ( .A1(A[6]), .A2(n84), .ZN(n82) );
  INV_X1 U57 ( .A(A[6]), .ZN(n64) );
  NAND2_X1 U58 ( .A1(A[10]), .A2(n84), .ZN(n129) );
  NAND2_X1 U59 ( .A1(n15), .A2(A[10]), .ZN(n164) );
  NAND2_X1 U60 ( .A1(A[20]), .A2(n15), .ZN(n99) );
  NAND2_X1 U61 ( .A1(A[17]), .A2(n15), .ZN(n126) );
  NAND2_X1 U62 ( .A1(A[17]), .A2(n84), .ZN(n103) );
  NAND2_X1 U63 ( .A1(A[5]), .A2(n84), .ZN(n168) );
  NAND2_X1 U64 ( .A1(A[5]), .A2(n54), .ZN(n83) );
  NAND2_X1 U65 ( .A1(A[20]), .A2(n84), .ZN(n109) );
  INV_X2 U66 ( .A(A[21]), .ZN(n17) );
  OAI21_X2 U67 ( .B1(n135), .B2(n19), .A(n103), .ZN(n134) );
  AOI21_X1 U68 ( .B1(A[11]), .B2(n20), .A(n4), .ZN(n51) );
  NAND2_X1 U69 ( .A1(A[11]), .A2(n14), .ZN(n150) );
  NAND2_X1 U70 ( .A1(A[11]), .A2(n84), .ZN(n163) );
  NAND2_X1 U71 ( .A1(A[9]), .A2(n84), .ZN(n52) );
  NAND2_X1 U72 ( .A1(A[9]), .A2(n14), .ZN(n130) );
  NAND2_X1 U73 ( .A1(A[8]), .A2(n14), .ZN(n53) );
  NAND2_X1 U74 ( .A1(A[8]), .A2(n84), .ZN(n145) );
  INV_X16 U75 ( .A(SH[2]), .ZN(n25) );
  NOR2_X4 U76 ( .A1(n18), .A2(n20), .ZN(n14) );
  NOR2_X4 U77 ( .A1(n18), .A2(n20), .ZN(n15) );
  INV_X8 U78 ( .A(n58), .ZN(n84) );
  INV_X8 U79 ( .A(n94), .ZN(n27) );
  INV_X32 U80 ( .A(n19), .ZN(n18) );
  INV_X32 U81 ( .A(n22), .ZN(n20) );
  INV_X32 U82 ( .A(n22), .ZN(n21) );
  NAND2_X2 U83 ( .A1(n25), .A2(n26), .ZN(n24) );
  NAND2_X2 U84 ( .A1(n27), .A2(n28), .ZN(n23) );
  NAND2_X2 U85 ( .A1(n32), .A2(n25), .ZN(n31) );
  NAND2_X2 U86 ( .A1(n27), .A2(n33), .ZN(n30) );
  NAND2_X2 U87 ( .A1(n38), .A2(n25), .ZN(n37) );
  NAND2_X2 U88 ( .A1(n27), .A2(n39), .ZN(n36) );
  NAND2_X2 U89 ( .A1(n43), .A2(n25), .ZN(n42) );
  NAND2_X2 U90 ( .A1(n27), .A2(n44), .ZN(n41) );
  NAND2_X2 U91 ( .A1(n25), .A2(n29), .ZN(n47) );
  NAND2_X2 U92 ( .A1(n27), .A2(n26), .ZN(n46) );
  NAND2_X2 U93 ( .A1(n27), .A2(n32), .ZN(n50) );
  OAI211_X2 U94 ( .C1(n51), .C2(n19), .A(n52), .B(n53), .ZN(n32) );
  NAND2_X2 U95 ( .A1(n34), .A2(n25), .ZN(n49) );
  NAND2_X2 U96 ( .A1(n27), .A2(n38), .ZN(n56) );
  NAND2_X2 U97 ( .A1(n60), .A2(n25), .ZN(n55) );
  INV_X4 U98 ( .A(n35), .ZN(n60) );
  MUX2_X2 U99 ( .A(n61), .B(n62), .S(n18), .Z(n35) );
  MUX2_X2 U100 ( .A(n63), .B(n64), .S(n20), .Z(n62) );
  NAND2_X2 U101 ( .A1(n68), .A2(n25), .ZN(n66) );
  INV_X4 U102 ( .A(n40), .ZN(n68) );
  MUX2_X2 U103 ( .A(n69), .B(n70), .S(n18), .Z(n40) );
  MUX2_X2 U104 ( .A(n71), .B(n63), .S(n21), .Z(n70) );
  INV_X4 U105 ( .A(A[5]), .ZN(n63) );
  NAND2_X2 U106 ( .A1(n27), .A2(n43), .ZN(n65) );
  NAND2_X2 U107 ( .A1(n73), .A2(n25), .ZN(n72) );
  INV_X4 U108 ( .A(n74), .ZN(n73) );
  NAND2_X2 U109 ( .A1(n77), .A2(n25), .ZN(n76) );
  NAND2_X2 U110 ( .A1(n27), .A2(n29), .ZN(n80) );
  NAND3_X2 U111 ( .A1(n81), .A2(n82), .A3(n83), .ZN(n29) );
  NAND2_X2 U112 ( .A1(n85), .A2(n18), .ZN(n81) );
  MUX2_X2 U113 ( .A(A[7]), .B(A[8]), .S(n21), .Z(n85) );
  NAND2_X2 U114 ( .A1(n86), .A2(n25), .ZN(n79) );
  INV_X4 U115 ( .A(n45), .ZN(n86) );
  MUX2_X2 U116 ( .A(n57), .B(n61), .S(n18), .Z(n45) );
  MUX2_X2 U117 ( .A(n87), .B(n71), .S(n21), .Z(n61) );
  MUX2_X2 U118 ( .A(n88), .B(n89), .S(n21), .Z(n57) );
  NAND2_X2 U119 ( .A1(n75), .A2(n25), .ZN(n95) );
  NAND2_X2 U120 ( .A1(n27), .A2(n77), .ZN(n97) );
  NAND2_X2 U121 ( .A1(n16), .A2(n84), .ZN(n98) );
  OAI211_X2 U122 ( .C1(n100), .C2(n19), .A(n101), .B(n102), .ZN(n33) );
  NAND2_X2 U123 ( .A1(A[12]), .A2(n14), .ZN(n102) );
  INV_X4 U124 ( .A(n78), .ZN(n96) );
  OAI211_X2 U125 ( .C1(n135), .C2(n19), .A(n103), .B(n104), .ZN(n78) );
  NAND2_X2 U126 ( .A1(A[16]), .A2(n54), .ZN(n104) );
  NAND2_X2 U127 ( .A1(n91), .A2(n25), .ZN(n107) );
  INV_X4 U128 ( .A(n90), .ZN(n106) );
  NAND3_X2 U129 ( .A1(n108), .A2(n109), .A3(n110), .ZN(n90) );
  NAND2_X2 U130 ( .A1(n111), .A2(n18), .ZN(n108) );
  NAND2_X2 U131 ( .A1(n93), .A2(n25), .ZN(n113) );
  INV_X4 U132 ( .A(n92), .ZN(n112) );
  NAND3_X2 U133 ( .A1(n114), .A2(n115), .A3(n116), .ZN(n92) );
  NAND2_X2 U134 ( .A1(n117), .A2(n18), .ZN(n114) );
  MUX2_X2 U135 ( .A(A[20]), .B(n16), .S(n21), .Z(n117) );
  NAND2_X2 U136 ( .A1(n25), .A2(n28), .ZN(n119) );
  NAND3_X2 U137 ( .A1(n120), .A2(n121), .A3(n122), .ZN(n28) );
  NAND2_X2 U138 ( .A1(A[13]), .A2(n54), .ZN(n122) );
  NAND2_X2 U139 ( .A1(n123), .A2(n18), .ZN(n120) );
  MUX2_X2 U140 ( .A(A[15]), .B(A[16]), .S(n21), .Z(n123) );
  NAND2_X2 U141 ( .A1(n27), .A2(n75), .ZN(n118) );
  NAND3_X2 U142 ( .A1(n124), .A2(n125), .A3(n126), .ZN(n75) );
  NAND2_X2 U143 ( .A1(n127), .A2(n18), .ZN(n124) );
  MUX2_X2 U144 ( .A(A[19]), .B(A[20]), .S(n21), .Z(n127) );
  NAND3_X2 U145 ( .A1(n128), .A2(n129), .A3(n130), .ZN(n26) );
  NAND2_X2 U146 ( .A1(n131), .A2(n18), .ZN(n128) );
  MUX2_X2 U147 ( .A(A[11]), .B(A[12]), .S(n21), .Z(n131) );
  OAI21_X4 U148 ( .B1(n134), .B2(n3), .A(n27), .ZN(n133) );
  INV_X4 U149 ( .A(n136), .ZN(n105) );
  INV_X4 U150 ( .A(n137), .ZN(n132) );
  OAI211_X2 U151 ( .C1(n100), .C2(n19), .A(n101), .B(n102), .ZN(n137) );
  NAND2_X2 U152 ( .A1(A[13]), .A2(n84), .ZN(n101) );
  NAND2_X2 U153 ( .A1(n27), .A2(n91), .ZN(n139) );
  NAND3_X2 U154 ( .A1(n140), .A2(n141), .A3(n142), .ZN(n91) );
  NAND2_X2 U155 ( .A1(A[15]), .A2(n54), .ZN(n142) );
  NAND2_X2 U156 ( .A1(A[16]), .A2(n84), .ZN(n141) );
  NAND2_X2 U157 ( .A1(n143), .A2(n18), .ZN(n140) );
  MUX2_X2 U158 ( .A(A[17]), .B(A[18]), .S(n20), .Z(n143) );
  NAND3_X2 U159 ( .A1(n144), .A2(n145), .A3(n146), .ZN(n38) );
  NAND2_X2 U160 ( .A1(n147), .A2(n18), .ZN(n144) );
  MUX2_X2 U161 ( .A(A[9]), .B(A[10]), .S(n21), .Z(n147) );
  INV_X4 U162 ( .A(n39), .ZN(n138) );
  NAND3_X2 U163 ( .A1(n148), .A2(n149), .A3(n150), .ZN(n39) );
  NAND2_X2 U164 ( .A1(A[12]), .A2(n84), .ZN(n149) );
  NAND2_X2 U165 ( .A1(n151), .A2(n18), .ZN(n148) );
  MUX2_X2 U166 ( .A(A[13]), .B(A[14]), .S(n20), .Z(n151) );
  NAND2_X2 U167 ( .A1(n27), .A2(n93), .ZN(n153) );
  NAND3_X2 U168 ( .A1(n154), .A2(n155), .A3(n156), .ZN(n93) );
  NAND2_X2 U169 ( .A1(A[15]), .A2(n84), .ZN(n155) );
  NAND2_X2 U170 ( .A1(n157), .A2(n18), .ZN(n154) );
  MUX2_X2 U171 ( .A(A[16]), .B(A[17]), .S(n21), .Z(n157) );
  NAND3_X2 U172 ( .A1(n158), .A2(n159), .A3(n160), .ZN(n43) );
  NAND2_X2 U173 ( .A1(n161), .A2(n18), .ZN(n158) );
  MUX2_X2 U174 ( .A(A[8]), .B(A[9]), .S(n20), .Z(n161) );
  INV_X4 U175 ( .A(n44), .ZN(n152) );
  NAND3_X2 U176 ( .A1(n162), .A2(n163), .A3(n164), .ZN(n44) );
  NAND2_X2 U177 ( .A1(n165), .A2(n18), .ZN(n162) );
  MUX2_X2 U178 ( .A(A[12]), .B(A[13]), .S(n20), .Z(n165) );
  OAI21_X4 U179 ( .B1(SH[2]), .B2(n48), .A(n166), .ZN(B[0]) );
  NAND2_X2 U180 ( .A1(n27), .A2(n34), .ZN(n166) );
  NAND3_X2 U181 ( .A1(n167), .A2(n168), .A3(n169), .ZN(n34) );
  NOR2_X4 U182 ( .A1(n18), .A2(n20), .ZN(n54) );
  NAND2_X2 U183 ( .A1(n21), .A2(n19), .ZN(n58) );
  NAND2_X2 U184 ( .A1(n170), .A2(n18), .ZN(n167) );
  MUX2_X2 U185 ( .A(A[6]), .B(A[7]), .S(n20), .Z(n170) );
  MUX2_X2 U186 ( .A(n67), .B(n69), .S(n18), .Z(n48) );
  MUX2_X2 U187 ( .A(n89), .B(n87), .S(n20), .Z(n69) );
  INV_X4 U188 ( .A(A[3]), .ZN(n87) );
  INV_X4 U189 ( .A(A[2]), .ZN(n89) );
  MUX2_X2 U190 ( .A(n59), .B(n88), .S(n21), .Z(n67) );
  INV_X4 U191 ( .A(A[1]), .ZN(n88) );
  INV_X4 U192 ( .A(A[0]), .ZN(n59) );
endmodule


module fpu_DW01_ash_4 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [2:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][20] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][0] , \ML_int[2][20] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][16] , \ML_int[2][15] ,
         \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][11] , \ML_int[2][9] ,
         \ML_int[2][8] , \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] ,
         \ML_int[2][4] , \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] ,
         \ML_int[2][0] , net85895, net85899, net85903, net88351, net88458,
         net88600, net88672, net88766, net88778, net88783, net88852, net88861,
         net88908, net88921, net88980, net88998, net89007, net89012, net89040,
         net89046, net89052, net89050, net89170, net89236, net89240, net89257,
         net89339, net89358, net89354, net89420, net89441, net89694, net89773,
         net90992, net91003, net91001, net91017, net91147, net91155, net91202,
         net91269, net91311, net91388, net91392, net91526, net99829, net99836,
         net99835, \ML_int[1][15] , net99764, net89357, net88995, net88994,
         net88993, net88992, net88991, net88990, net85898, net85894,
         \ML_int[2][21] , \ML_int[2][17] , \ML_int[1][21] , \ML_int[1][19] ,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100
;

  MUX2_X2 M1_2_10 ( .A(n16), .B(\ML_int[2][6] ), .S(net85895), .Z(B[10]) );
  MUX2_X2 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(net85895), .Z(
        B[8]) );
  MUX2_X2 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(net85895), .Z(
        B[7]) );
  MUX2_X2 M1_2_5 ( .A(\ML_int[2][5] ), .B(\ML_int[2][1] ), .S(net85895), .Z(
        B[5]) );
  MUX2_X2 M1_0_20 ( .A(A[20]), .B(A[19]), .S(net88600), .Z(\ML_int[1][20] ) );
  MUX2_X2 M1_0_11 ( .A(A[11]), .B(A[10]), .S(net85903), .Z(\ML_int[1][11] ) );
  MUX2_X2 M1_0_9 ( .A(A[9]), .B(A[8]), .S(net88672), .Z(\ML_int[1][9] ) );
  MUX2_X2 M1_0_14 ( .A(A[14]), .B(A[13]), .S(net88672), .Z(\ML_int[1][14] ) );
  MUX2_X2 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S(net85899), 
        .Z(\ML_int[2][21] ) );
  MUX2_X2 M0_0_0 ( .A(A[0]), .B(1'b0), .S(net88672), .Z(\ML_int[1][0] ) );
  NAND2_X2 U3 ( .A1(net99764), .A2(net88990), .ZN(net88991) );
  NAND2_X2 U4 ( .A1(A[19]), .A2(net89357), .ZN(n10) );
  NAND2_X2 U5 ( .A1(\ML_int[1][5] ), .A2(net88766), .ZN(n18) );
  NAND2_X4 U6 ( .A1(n77), .A2(n78), .ZN(n1) );
  NAND2_X1 U7 ( .A1(n77), .A2(n78), .ZN(n16) );
  NAND2_X1 U8 ( .A1(\ML_int[2][11] ), .A2(net89236), .ZN(n53) );
  NAND2_X2 U9 ( .A1(n63), .A2(n64), .ZN(n2) );
  NAND2_X2 U10 ( .A1(A[11]), .A2(n4), .ZN(n64) );
  NAND2_X2 U11 ( .A1(\ML_int[1][7] ), .A2(net89012), .ZN(n27) );
  NAND2_X1 U12 ( .A1(A[21]), .A2(net89257), .ZN(n11) );
  NAND2_X1 U13 ( .A1(\ML_int[1][20] ), .A2(net91392), .ZN(n83) );
  NAND2_X2 U14 ( .A1(\ML_int[1][6] ), .A2(net89046), .ZN(n61) );
  NAND2_X2 U15 ( .A1(n24), .A2(n25), .ZN(\ML_int[2][14] ) );
  INV_X4 U16 ( .A(net88600), .ZN(n3) );
  INV_X4 U17 ( .A(n3), .ZN(n4) );
  NAND2_X2 U18 ( .A1(A[3]), .A2(net85903), .ZN(n62) );
  INV_X1 U19 ( .A(n76), .ZN(n5) );
  INV_X4 U20 ( .A(net85895), .ZN(net88351) );
  INV_X4 U21 ( .A(net88351), .ZN(net88861) );
  NAND2_X4 U22 ( .A1(net88458), .A2(n2), .ZN(n96) );
  NOR2_X2 U23 ( .A1(n40), .A2(net85898), .ZN(n8) );
  INV_X1 U24 ( .A(A[9]), .ZN(n46) );
  NAND2_X2 U25 ( .A1(\ML_int[1][10] ), .A2(net85899), .ZN(n97) );
  NAND2_X2 U26 ( .A1(\ML_int[1][6] ), .A2(net85899), .ZN(n57) );
  NAND2_X2 U27 ( .A1(n33), .A2(n34), .ZN(\ML_int[2][13] ) );
  NAND2_X2 U28 ( .A1(n22), .A2(n23), .ZN(\ML_int[2][9] ) );
  INV_X1 U29 ( .A(A[0]), .ZN(n42) );
  INV_X1 U30 ( .A(A[1]), .ZN(n41) );
  INV_X8 U31 ( .A(net85895), .ZN(net91311) );
  NAND2_X2 U32 ( .A1(n60), .A2(n61), .ZN(\ML_int[2][6] ) );
  NAND2_X2 U33 ( .A1(\ML_int[1][4] ), .A2(net89354), .ZN(n60) );
  NAND2_X2 U34 ( .A1(\ML_int[2][8] ), .A2(net88861), .ZN(n87) );
  NAND2_X2 U35 ( .A1(net88351), .A2(n17), .ZN(n88) );
  NAND2_X2 U36 ( .A1(\ML_int[2][7] ), .A2(net88861), .ZN(n52) );
  NAND2_X2 U37 ( .A1(n70), .A2(n69), .ZN(B[13]) );
  NAND2_X2 U38 ( .A1(net88600), .A2(A[18]), .ZN(net89773) );
  INV_X8 U39 ( .A(net88600), .ZN(net89257) );
  INV_X8 U40 ( .A(n13), .ZN(net85903) );
  NAND2_X2 U41 ( .A1(n31), .A2(n32), .ZN(\ML_int[2][18] ) );
  NAND2_X4 U42 ( .A1(n48), .A2(n49), .ZN(B[15]) );
  NAND2_X4 U43 ( .A1(\ML_int[1][3] ), .A2(net89007), .ZN(n75) );
  NAND2_X2 U44 ( .A1(\ML_int[1][3] ), .A2(net85899), .ZN(n19) );
  NAND2_X1 U45 ( .A1(A[20]), .A2(net85903), .ZN(n12) );
  NAND2_X4 U46 ( .A1(n36), .A2(n37), .ZN(B[19]) );
  NAND2_X2 U47 ( .A1(\ML_int[2][15] ), .A2(net85895), .ZN(n37) );
  NAND2_X2 U48 ( .A1(\ML_int[1][8] ), .A2(net89441), .ZN(n56) );
  NAND2_X4 U49 ( .A1(n73), .A2(net89040), .ZN(B[17]) );
  NAND2_X4 U50 ( .A1(\ML_int[2][17] ), .A2(net88778), .ZN(net89040) );
  NAND2_X4 U51 ( .A1(n95), .A2(n94), .ZN(\ML_int[2][16] ) );
  MUX2_X2 U52 ( .A(A[18]), .B(A[17]), .S(net88600), .Z(n6) );
  NAND2_X4 U53 ( .A1(n47), .A2(net88908), .ZN(n82) );
  NAND2_X2 U54 ( .A1(\ML_int[1][15] ), .A2(net85899), .ZN(net88992) );
  NAND2_X2 U55 ( .A1(\ML_int[1][15] ), .A2(net88766), .ZN(net88783) );
  NAND2_X2 U56 ( .A1(net99836), .A2(net89050), .ZN(n72) );
  INV_X4 U57 ( .A(net99835), .ZN(net99836) );
  NAND2_X4 U58 ( .A1(n17), .A2(net85895), .ZN(n29) );
  NAND2_X4 U59 ( .A1(n97), .A2(n96), .ZN(n17) );
  NOR2_X4 U60 ( .A1(n100), .A2(net85899), .ZN(\ML_int[2][0] ) );
  INV_X4 U61 ( .A(\ML_int[1][0] ), .ZN(n100) );
  INV_X2 U62 ( .A(net85899), .ZN(net89046) );
  OAI21_X1 U63 ( .B1(n5), .B2(n9), .A(net85894), .ZN(n7) );
  INV_X2 U64 ( .A(n7), .ZN(B[3]) );
  INV_X4 U65 ( .A(n8), .ZN(n76) );
  INV_X1 U66 ( .A(n75), .ZN(n9) );
  AND2_X2 U67 ( .A1(\ML_int[2][1] ), .A2(net85894), .ZN(B[1]) );
  NAND2_X4 U68 ( .A1(net88994), .A2(net88995), .ZN(B[21]) );
  NAND2_X4 U69 ( .A1(\ML_int[2][17] ), .A2(net85895), .ZN(net88995) );
  INV_X32 U70 ( .A(net85894), .ZN(net85895) );
  INV_X8 U71 ( .A(SH[2]), .ZN(net85894) );
  NAND2_X4 U72 ( .A1(\ML_int[2][21] ), .A2(net88993), .ZN(net88994) );
  INV_X1 U73 ( .A(net85895), .ZN(net88993) );
  INV_X32 U74 ( .A(net85898), .ZN(net85899) );
  INV_X8 U75 ( .A(SH[1]), .ZN(net85898) );
  NAND2_X2 U76 ( .A1(n12), .A2(n11), .ZN(\ML_int[1][21] ) );
  INV_X2 U77 ( .A(net89257), .ZN(net91526) );
  NAND2_X1 U78 ( .A1(A[13]), .A2(net89257), .ZN(net91001) );
  INV_X16 U79 ( .A(n13), .ZN(net88600) );
  INV_X16 U80 ( .A(SH[0]), .ZN(n13) );
  INV_X16 U81 ( .A(n13), .ZN(net88672) );
  NAND2_X4 U82 ( .A1(net88991), .A2(net88992), .ZN(\ML_int[2][17] ) );
  INV_X1 U83 ( .A(net85899), .ZN(net88990) );
  NAND2_X4 U84 ( .A1(net89773), .A2(n10), .ZN(\ML_int[1][19] ) );
  INV_X1 U85 ( .A(\ML_int[1][19] ), .ZN(net99835) );
  INV_X4 U86 ( .A(net85903), .ZN(net89357) );
  NAND2_X1 U87 ( .A1(A[2]), .A2(net89357), .ZN(net91147) );
  NAND2_X1 U88 ( .A1(A[4]), .A2(net89357), .ZN(net89358) );
  MUX2_X2 U89 ( .A(A[17]), .B(A[16]), .S(net88672), .Z(net99764) );
  NAND2_X2 U90 ( .A1(net85899), .A2(net99764), .ZN(net89052) );
  MUX2_X2 U91 ( .A(A[16]), .B(A[15]), .S(net88600), .Z(net99829) );
  NAND2_X4 U92 ( .A1(n14), .A2(n15), .ZN(\ML_int[1][15] ) );
  NAND2_X1 U93 ( .A1(A[14]), .A2(net88600), .ZN(n15) );
  NAND2_X2 U94 ( .A1(A[15]), .A2(net89257), .ZN(n14) );
  NAND2_X1 U95 ( .A1(A[3]), .A2(net89257), .ZN(net89170) );
  NAND2_X4 U96 ( .A1(\ML_int[2][13] ), .A2(net88980), .ZN(n73) );
  NAND2_X2 U97 ( .A1(\ML_int[2][14] ), .A2(net89420), .ZN(n58) );
  INV_X1 U98 ( .A(net85899), .ZN(net88908) );
  NAND2_X4 U99 ( .A1(\ML_int[2][14] ), .A2(net88980), .ZN(n79) );
  NAND2_X4 U100 ( .A1(n1), .A2(net85895), .ZN(n59) );
  NAND2_X4 U101 ( .A1(\ML_int[2][11] ), .A2(net88980), .ZN(n48) );
  NAND2_X4 U102 ( .A1(n81), .A2(n82), .ZN(\ML_int[2][11] ) );
  INV_X4 U103 ( .A(net85895), .ZN(net88778) );
  NAND2_X4 U104 ( .A1(n59), .A2(n58), .ZN(B[14]) );
  INV_X1 U105 ( .A(A[10]), .ZN(n45) );
  NAND2_X2 U106 ( .A1(net85899), .A2(net99829), .ZN(n32) );
  NAND2_X2 U107 ( .A1(n85), .A2(n86), .ZN(\ML_int[1][6] ) );
  NAND2_X1 U108 ( .A1(A[8]), .A2(net89257), .ZN(n54) );
  NAND2_X2 U109 ( .A1(n62), .A2(net89358), .ZN(\ML_int[1][4] ) );
  NAND2_X1 U110 ( .A1(A[2]), .A2(net85903), .ZN(n71) );
  NAND2_X2 U111 ( .A1(n54), .A2(n55), .ZN(\ML_int[1][8] ) );
  NAND2_X2 U112 ( .A1(n18), .A2(n19), .ZN(\ML_int[2][5] ) );
  NAND2_X2 U113 ( .A1(\ML_int[2][5] ), .A2(net85895), .ZN(n51) );
  NAND2_X1 U114 ( .A1(A[4]), .A2(net88600), .ZN(n68) );
  INV_X2 U115 ( .A(net88908), .ZN(net88921) );
  INV_X2 U116 ( .A(net89046), .ZN(net89354) );
  INV_X2 U117 ( .A(net89012), .ZN(net91202) );
  NAND2_X4 U118 ( .A1(\ML_int[2][19] ), .A2(net91003), .ZN(n36) );
  NAND2_X2 U119 ( .A1(\ML_int[2][15] ), .A2(net88351), .ZN(n49) );
  NAND2_X4 U120 ( .A1(n91), .A2(net88783), .ZN(\ML_int[2][15] ) );
  NAND2_X2 U121 ( .A1(\ML_int[1][11] ), .A2(net85899), .ZN(n34) );
  NAND2_X2 U122 ( .A1(\ML_int[1][9] ), .A2(net88921), .ZN(n81) );
  NAND2_X2 U123 ( .A1(n74), .A2(net91392), .ZN(n20) );
  NAND2_X1 U124 ( .A1(\ML_int[1][0] ), .A2(net85899), .ZN(n21) );
  NAND2_X2 U125 ( .A1(n20), .A2(n21), .ZN(\ML_int[2][2] ) );
  INV_X1 U126 ( .A(net85899), .ZN(net91392) );
  NOR2_X1 U127 ( .A1(net85895), .A2(n99), .ZN(B[0]) );
  NOR2_X1 U128 ( .A1(n98), .A2(net85895), .ZN(B[2]) );
  NAND2_X2 U129 ( .A1(\ML_int[1][9] ), .A2(net91388), .ZN(n22) );
  NAND2_X2 U130 ( .A1(\ML_int[1][7] ), .A2(net85899), .ZN(n23) );
  INV_X1 U131 ( .A(net85899), .ZN(net91388) );
  NAND2_X2 U132 ( .A1(\ML_int[2][9] ), .A2(net85895), .ZN(n70) );
  NAND2_X2 U133 ( .A1(\ML_int[2][9] ), .A2(net89694), .ZN(n50) );
  NAND2_X1 U134 ( .A1(A[6]), .A2(n4), .ZN(n93) );
  NAND2_X1 U135 ( .A1(\ML_int[1][12] ), .A2(net85899), .ZN(n25) );
  NAND2_X2 U136 ( .A1(\ML_int[1][14] ), .A2(net91269), .ZN(n24) );
  NAND2_X2 U137 ( .A1(n6), .A2(net91017), .ZN(n31) );
  NAND2_X2 U138 ( .A1(\ML_int[1][14] ), .A2(net91202), .ZN(n94) );
  MUX2_X2 U139 ( .A(\ML_int[2][0] ), .B(\ML_int[2][4] ), .S(net91311), .Z(B[4]) );
  NAND2_X4 U140 ( .A1(\ML_int[2][16] ), .A2(net91155), .ZN(n28) );
  NAND2_X1 U141 ( .A1(A[7]), .A2(net89257), .ZN(n92) );
  INV_X1 U142 ( .A(net85899), .ZN(net91269) );
  NAND2_X2 U143 ( .A1(\ML_int[2][16] ), .A2(net85895), .ZN(n39) );
  NAND2_X4 U144 ( .A1(\ML_int[2][18] ), .A2(net88778), .ZN(n80) );
  NAND2_X4 U145 ( .A1(n80), .A2(n79), .ZN(B[18]) );
  NAND2_X1 U146 ( .A1(\ML_int[1][5] ), .A2(net91202), .ZN(n26) );
  NAND2_X2 U147 ( .A1(n26), .A2(n27), .ZN(\ML_int[2][7] ) );
  NAND2_X2 U148 ( .A1(n92), .A2(n93), .ZN(\ML_int[1][7] ) );
  INV_X1 U149 ( .A(net85899), .ZN(net89012) );
  NAND2_X4 U150 ( .A1(n29), .A2(n28), .ZN(B[16]) );
  INV_X1 U151 ( .A(net85895), .ZN(net91155) );
  NAND2_X1 U152 ( .A1(A[1]), .A2(net88600), .ZN(n30) );
  NAND2_X2 U153 ( .A1(net91147), .A2(n30), .ZN(\ML_int[1][2] ) );
  NAND2_X2 U154 ( .A1(net99829), .A2(net91388), .ZN(n95) );
  NAND2_X1 U155 ( .A1(A[5]), .A2(net88600), .ZN(n86) );
  INV_X1 U156 ( .A(net85899), .ZN(net91017) );
  NAND2_X2 U157 ( .A1(n43), .A2(net91269), .ZN(n33) );
  NAND2_X2 U158 ( .A1(\ML_int[2][13] ), .A2(net89240), .ZN(n69) );
  NAND2_X1 U159 ( .A1(A[12]), .A2(net91526), .ZN(n35) );
  NAND2_X2 U160 ( .A1(net91001), .A2(n35), .ZN(\ML_int[1][13] ) );
  INV_X1 U161 ( .A(net85895), .ZN(net91003) );
  NAND2_X2 U162 ( .A1(\ML_int[1][13] ), .A2(net88921), .ZN(n91) );
  NAND2_X2 U163 ( .A1(\ML_int[2][20] ), .A2(net90992), .ZN(n38) );
  NAND2_X2 U164 ( .A1(n38), .A2(n39), .ZN(B[20]) );
  INV_X1 U165 ( .A(net85895), .ZN(net90992) );
  NAND2_X2 U166 ( .A1(\ML_int[1][2] ), .A2(net85899), .ZN(n66) );
  MUX2_X2 U167 ( .A(n41), .B(n42), .S(net88600), .Z(n40) );
  MUX2_X2 U168 ( .A(A[13]), .B(A[12]), .S(net88600), .Z(n43) );
  MUX2_X2 U169 ( .A(n45), .B(n46), .S(net88672), .Z(n44) );
  INV_X4 U170 ( .A(n44), .ZN(\ML_int[1][10] ) );
  INV_X1 U171 ( .A(\ML_int[2][0] ), .ZN(n99) );
  MUX2_X2 U172 ( .A(A[11]), .B(A[10]), .S(net85903), .Z(n47) );
  NAND2_X2 U173 ( .A1(n75), .A2(n76), .ZN(\ML_int[2][3] ) );
  NAND2_X2 U174 ( .A1(n50), .A2(n51), .ZN(B[9]) );
  INV_X1 U175 ( .A(net85895), .ZN(net89694) );
  NAND2_X1 U176 ( .A1(\ML_int[2][6] ), .A2(net88852), .ZN(n89) );
  NAND2_X2 U177 ( .A1(\ML_int[2][2] ), .A2(net85895), .ZN(n90) );
  NAND2_X4 U178 ( .A1(n52), .A2(n53), .ZN(B[11]) );
  INV_X1 U179 ( .A(net85895), .ZN(net89236) );
  NAND2_X1 U180 ( .A1(A[7]), .A2(net85903), .ZN(n55) );
  NAND2_X4 U181 ( .A1(n56), .A2(n57), .ZN(\ML_int[2][8] ) );
  INV_X1 U182 ( .A(net85899), .ZN(net89441) );
  NAND2_X2 U183 ( .A1(\ML_int[1][8] ), .A2(net85899), .ZN(n78) );
  INV_X1 U184 ( .A(net85895), .ZN(net89420) );
  INV_X2 U185 ( .A(\ML_int[2][2] ), .ZN(n98) );
  NAND2_X4 U186 ( .A1(\ML_int[1][4] ), .A2(net89339), .ZN(n65) );
  NAND2_X2 U187 ( .A1(n6), .A2(net85899), .ZN(n84) );
  NAND2_X2 U188 ( .A1(A[12]), .A2(net89357), .ZN(n63) );
  NAND2_X2 U189 ( .A1(n63), .A2(n64), .ZN(\ML_int[1][12] ) );
  NAND2_X2 U190 ( .A1(n65), .A2(n66), .ZN(\ML_int[2][4] ) );
  INV_X1 U191 ( .A(net85899), .ZN(net89339) );
  NAND2_X1 U192 ( .A1(A[5]), .A2(net89257), .ZN(n67) );
  NAND2_X2 U193 ( .A1(n67), .A2(n68), .ZN(\ML_int[1][5] ) );
  NOR2_X2 U194 ( .A1(net85899), .A2(n40), .ZN(\ML_int[2][1] ) );
  INV_X1 U195 ( .A(net85895), .ZN(net89240) );
  NAND2_X2 U196 ( .A1(net89170), .A2(n71), .ZN(\ML_int[1][3] ) );
  NAND2_X2 U197 ( .A1(n72), .A2(net89052), .ZN(\ML_int[2][19] ) );
  INV_X1 U198 ( .A(net85899), .ZN(net89050) );
  MUX2_X2 U199 ( .A(A[2]), .B(A[1]), .S(net85903), .Z(n74) );
  INV_X1 U200 ( .A(net85899), .ZN(net89007) );
  NAND2_X2 U201 ( .A1(\ML_int[1][10] ), .A2(net88998), .ZN(n77) );
  INV_X1 U202 ( .A(net85899), .ZN(net88998) );
  INV_X4 U203 ( .A(net88778), .ZN(net88980) );
  NAND2_X2 U204 ( .A1(n83), .A2(n84), .ZN(\ML_int[2][20] ) );
  NAND2_X1 U205 ( .A1(A[6]), .A2(net89257), .ZN(n85) );
  NAND2_X4 U206 ( .A1(n87), .A2(n88), .ZN(B[12]) );
  NAND2_X2 U207 ( .A1(n90), .A2(n89), .ZN(B[6]) );
  INV_X1 U208 ( .A(net85895), .ZN(net88852) );
  INV_X1 U209 ( .A(net85899), .ZN(net88766) );
  INV_X1 U210 ( .A(net85899), .ZN(net88458) );
endmodule


module fpu_DW01_sub_23 ( A, B, CI, DIFF, CO );
  input [6:0] A;
  input [6:0] B;
  output [6:0] DIFF;
  input CI;
  output CO;
  wire   net64864, net64862, net64843, net64841, net64840, net85706, net89571,
         net89670, net89739, net64871, net90964, net90963, net90960, net90954,
         net90950, net90938, net90300, net64870, net64847, net64863, net64848,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;
  assign net85706 = A[1];

  OAI21_X2 U3 ( .B1(net64840), .B2(net64841), .A(net64864), .ZN(n17) );
  INV_X4 U4 ( .A(n23), .ZN(n19) );
  NAND2_X2 U5 ( .A1(net89739), .A2(net64843), .ZN(net64864) );
  NAND2_X1 U6 ( .A1(n1), .A2(n4), .ZN(net90938) );
  INV_X1 U7 ( .A(n9), .ZN(net89739) );
  INV_X8 U8 ( .A(A[2]), .ZN(net64843) );
  NAND2_X1 U9 ( .A1(net89571), .A2(n8), .ZN(net64841) );
  INV_X4 U10 ( .A(net85706), .ZN(n1) );
  NOR2_X4 U11 ( .A1(n2), .A2(n1), .ZN(n3) );
  AOI21_X4 U12 ( .B1(net64863), .B2(net90300), .A(n3), .ZN(net64870) );
  NAND2_X2 U13 ( .A1(n2), .A2(n1), .ZN(net64863) );
  INV_X8 U14 ( .A(net64848), .ZN(n2) );
  BUF_X32 U15 ( .A(n2), .Z(n4) );
  INV_X8 U16 ( .A(B[1]), .ZN(net64848) );
  NAND2_X1 U17 ( .A1(net85706), .A2(net64848), .ZN(net89571) );
  NOR2_X1 U18 ( .A1(net85706), .A2(net64848), .ZN(net64847) );
  XNOR2_X2 U19 ( .A(B[1]), .B(net85706), .ZN(net90964) );
  XNOR2_X2 U20 ( .A(net64870), .B(net64871), .ZN(DIFF[2]) );
  INV_X8 U21 ( .A(net90954), .ZN(net90300) );
  NAND3_X1 U22 ( .A1(net90938), .A2(net90300), .A3(net64864), .ZN(net64862) );
  INV_X4 U23 ( .A(net90950), .ZN(net90954) );
  NOR2_X2 U24 ( .A1(net64847), .A2(net90954), .ZN(net64840) );
  XNOR2_X2 U25 ( .A(net90954), .B(net90964), .ZN(DIFF[1]) );
  NAND2_X4 U26 ( .A1(B[0]), .A2(n5), .ZN(net90950) );
  NAND2_X2 U27 ( .A1(net90950), .A2(net90963), .ZN(DIFF[0]) );
  INV_X4 U28 ( .A(A[0]), .ZN(n5) );
  INV_X4 U29 ( .A(B[0]), .ZN(net90960) );
  NAND2_X2 U30 ( .A1(A[0]), .A2(net90960), .ZN(net90963) );
  NOR2_X4 U31 ( .A1(n7), .A2(n6), .ZN(net64871) );
  NOR2_X4 U32 ( .A1(n9), .A2(A[2]), .ZN(n6) );
  INV_X8 U33 ( .A(B[2]), .ZN(n9) );
  NAND2_X4 U34 ( .A1(n9), .A2(A[2]), .ZN(n8) );
  INV_X8 U35 ( .A(n8), .ZN(n7) );
  NOR2_X2 U36 ( .A1(n22), .A2(B[4]), .ZN(n10) );
  INV_X4 U37 ( .A(n10), .ZN(n21) );
  NAND2_X4 U38 ( .A1(n24), .A2(n25), .ZN(n16) );
  INV_X4 U39 ( .A(n15), .ZN(n11) );
  NAND2_X1 U40 ( .A1(n22), .A2(B[4]), .ZN(n25) );
  INV_X4 U41 ( .A(B[3]), .ZN(n35) );
  NAND2_X1 U42 ( .A1(n29), .A2(n24), .ZN(n28) );
  INV_X1 U43 ( .A(net89571), .ZN(net89670) );
  NAND2_X2 U44 ( .A1(n15), .A2(A[5]), .ZN(n13) );
  NAND2_X4 U45 ( .A1(n11), .A2(n12), .ZN(n14) );
  NAND2_X4 U46 ( .A1(n14), .A2(n13), .ZN(DIFF[5]) );
  INV_X4 U47 ( .A(A[5]), .ZN(n12) );
  AOI21_X1 U48 ( .B1(n34), .B2(net89670), .A(n7), .ZN(n33) );
  NAND2_X1 U49 ( .A1(n25), .A2(n21), .ZN(n26) );
  NAND2_X4 U50 ( .A1(n35), .A2(A[3]), .ZN(n23) );
  NAND2_X2 U51 ( .A1(B[4]), .A2(n22), .ZN(n20) );
  NAND2_X1 U52 ( .A1(n24), .A2(n23), .ZN(n31) );
  NAND2_X1 U53 ( .A1(n28), .A2(n23), .ZN(n27) );
  NAND2_X1 U54 ( .A1(net64843), .A2(net89739), .ZN(n34) );
  OAI21_X4 U55 ( .B1(n17), .B2(n16), .A(n18), .ZN(n15) );
  AOI21_X4 U56 ( .B1(n19), .B2(n20), .A(n10), .ZN(n18) );
  XNOR2_X2 U57 ( .A(n26), .B(n27), .ZN(DIFF[4]) );
  INV_X4 U58 ( .A(A[4]), .ZN(n22) );
  INV_X4 U59 ( .A(n30), .ZN(DIFF[3]) );
  XNOR2_X2 U60 ( .A(n31), .B(n32), .ZN(n30) );
  INV_X4 U61 ( .A(n29), .ZN(n32) );
  NAND2_X2 U62 ( .A1(n33), .A2(net64862), .ZN(n29) );
  NAND2_X2 U63 ( .A1(n36), .A2(B[3]), .ZN(n24) );
  INV_X4 U64 ( .A(A[3]), .ZN(n36) );
endmodule


module fpu_DW_rash_11 ( A, DATA_TC, SH, SH_TC, B );
  input [13:0] A;
  input [3:0] SH;
  output [13:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140;

  NAND2_X2 U3 ( .A1(A[9]), .A2(n130), .ZN(n129) );
  NAND2_X2 U4 ( .A1(A[8]), .A2(n130), .ZN(n103) );
  NAND2_X2 U5 ( .A1(n130), .A2(A[4]), .ZN(n99) );
  NAND2_X2 U6 ( .A1(A[11]), .A2(n130), .ZN(n112) );
  NAND2_X2 U7 ( .A1(A[7]), .A2(n130), .ZN(n118) );
  INV_X8 U8 ( .A(n131), .ZN(n130) );
  NAND2_X4 U9 ( .A1(A[10]), .A2(n69), .ZN(n89) );
  NAND2_X4 U10 ( .A1(n34), .A2(n35), .ZN(B[5]) );
  NOR2_X2 U11 ( .A1(n73), .A2(n74), .ZN(n63) );
  NOR2_X1 U12 ( .A1(n32), .A2(n14), .ZN(n53) );
  NOR2_X1 U13 ( .A1(n15), .A2(n12), .ZN(n132) );
  NAND2_X2 U14 ( .A1(A[5]), .A2(n130), .ZN(n137) );
  NOR2_X2 U15 ( .A1(n21), .A2(n12), .ZN(n41) );
  NOR2_X1 U16 ( .A1(n20), .A2(n14), .ZN(n17) );
  NOR2_X1 U17 ( .A1(n19), .A2(n12), .ZN(n18) );
  NOR3_X2 U18 ( .A1(n59), .A2(SH[2]), .A3(n2), .ZN(n58) );
  NOR2_X2 U19 ( .A1(n9), .A2(n10), .ZN(n6) );
  NOR2_X1 U20 ( .A1(n13), .A2(n14), .ZN(n9) );
  NOR2_X1 U21 ( .A1(n13), .A2(n12), .ZN(n72) );
  NOR2_X1 U22 ( .A1(n5), .A2(n12), .ZN(n54) );
  NOR2_X2 U23 ( .A1(n132), .A2(n133), .ZN(n123) );
  INV_X4 U24 ( .A(SH[3]), .ZN(n134) );
  AND2_X2 U25 ( .A1(SH[0]), .A2(SH[1]), .ZN(n1) );
  AND2_X2 U26 ( .A1(n27), .A2(n8), .ZN(n2) );
  OR2_X4 U27 ( .A1(n19), .A2(n14), .ZN(n3) );
  AND2_X2 U28 ( .A1(A[7]), .A2(n69), .ZN(n4) );
  AND3_X4 U29 ( .A1(n121), .A2(n122), .A3(n120), .ZN(n5) );
  NOR2_X2 U30 ( .A1(n20), .A2(n12), .ZN(B[12]) );
  NOR2_X1 U31 ( .A1(n33), .A2(n12), .ZN(B[10]) );
  NAND2_X4 U32 ( .A1(n36), .A2(n64), .ZN(n35) );
  OAI21_X2 U33 ( .B1(n7), .B2(SH[3]), .A(n37), .ZN(n36) );
  NOR2_X2 U34 ( .A1(n11), .A2(n44), .ZN(n59) );
  NOR2_X1 U35 ( .A1(n11), .A2(n14), .ZN(n38) );
  NOR2_X1 U36 ( .A1(n11), .A2(n12), .ZN(n10) );
  AND4_X4 U37 ( .A1(n75), .A2(n76), .A3(n77), .A4(n78), .ZN(n11) );
  NAND2_X1 U38 ( .A1(n27), .A2(n28), .ZN(n22) );
  NAND3_X2 U39 ( .A1(n45), .A2(n46), .A3(n47), .ZN(B[3]) );
  INV_X1 U40 ( .A(SH[0]), .ZN(n140) );
  NAND3_X2 U41 ( .A1(n89), .A2(n90), .A3(n91), .ZN(n88) );
  NAND3_X2 U42 ( .A1(n107), .A2(n108), .A3(n106), .ZN(n26) );
  NAND2_X2 U43 ( .A1(A[6]), .A2(n130), .ZN(n84) );
  NOR2_X4 U44 ( .A1(SH[1]), .A2(SH[0]), .ZN(n24) );
  NAND2_X2 U45 ( .A1(A[5]), .A2(n24), .ZN(n82) );
  NAND2_X2 U46 ( .A1(A[12]), .A2(n24), .ZN(n87) );
  NOR2_X2 U47 ( .A1(SH[2]), .A2(SH[3]), .ZN(n27) );
  NOR2_X1 U48 ( .A1(n21), .A2(n14), .ZN(n133) );
  AND4_X4 U49 ( .A1(n135), .A2(n136), .A3(n137), .A4(n138), .ZN(n21) );
  NAND2_X1 U50 ( .A1(n130), .A2(A[3]), .ZN(n121) );
  INV_X2 U51 ( .A(SH[1]), .ZN(n70) );
  NAND2_X1 U52 ( .A1(n87), .A2(n86), .ZN(n127) );
  NOR2_X2 U53 ( .A1(n7), .A2(SH[3]), .ZN(n65) );
  INV_X1 U54 ( .A(n24), .ZN(n73) );
  NAND2_X2 U55 ( .A1(SH[0]), .A2(n70), .ZN(n131) );
  NAND2_X1 U56 ( .A1(A[6]), .A2(n24), .ZN(n116) );
  NAND2_X1 U57 ( .A1(A[10]), .A2(n24), .ZN(n110) );
  NAND2_X1 U58 ( .A1(A[3]), .A2(n24), .ZN(n97) );
  NAND2_X1 U59 ( .A1(A[7]), .A2(n24), .ZN(n101) );
  NAND2_X1 U60 ( .A1(A[9]), .A2(n24), .ZN(n75) );
  NAND2_X1 U61 ( .A1(A[4]), .A2(n24), .ZN(n135) );
  NAND2_X4 U62 ( .A1(A[8]), .A2(n24), .ZN(n95) );
  NAND3_X1 U63 ( .A1(SH[1]), .A2(SH[0]), .A3(A[8]), .ZN(n83) );
  NAND3_X1 U64 ( .A1(A[13]), .A2(n70), .A3(SH[0]), .ZN(n86) );
  INV_X4 U65 ( .A(n6), .ZN(B[9]) );
  NAND2_X2 U66 ( .A1(n66), .A2(n67), .ZN(n8) );
  NAND2_X2 U67 ( .A1(n86), .A2(n87), .ZN(n43) );
  INV_X4 U68 ( .A(n96), .ZN(B[11]) );
  NAND2_X2 U69 ( .A1(n51), .A2(n52), .ZN(B[2]) );
  NAND3_X4 U70 ( .A1(n3), .A2(n40), .A3(n39), .ZN(B[4]) );
  NAND2_X2 U71 ( .A1(n22), .A2(n23), .ZN(B[7]) );
  INV_X4 U72 ( .A(n29), .ZN(B[6]) );
  INV_X4 U73 ( .A(n16), .ZN(B[8]) );
  INV_X4 U74 ( .A(n37), .ZN(n60) );
  NAND2_X2 U75 ( .A1(n1), .A2(A[3]), .ZN(n15) );
  INV_X4 U76 ( .A(n72), .ZN(n71) );
  INV_X4 U77 ( .A(n48), .ZN(n47) );
  NAND2_X4 U78 ( .A1(SH[2]), .A2(n134), .ZN(n14) );
  INV_X8 U79 ( .A(n139), .ZN(n69) );
  NAND2_X4 U80 ( .A1(SH[1]), .A2(SH[0]), .ZN(n68) );
  INV_X8 U81 ( .A(n27), .ZN(n12) );
  NOR2_X4 U82 ( .A1(n17), .A2(n18), .ZN(n16) );
  NAND2_X2 U83 ( .A1(n25), .A2(n26), .ZN(n23) );
  INV_X4 U84 ( .A(n14), .ZN(n25) );
  NOR2_X4 U85 ( .A1(n30), .A2(n31), .ZN(n29) );
  NOR2_X4 U86 ( .A1(n32), .A2(n12), .ZN(n31) );
  NOR2_X4 U87 ( .A1(n33), .A2(n14), .ZN(n30) );
  INV_X4 U88 ( .A(n38), .ZN(n34) );
  INV_X4 U89 ( .A(n41), .ZN(n40) );
  NAND2_X2 U90 ( .A1(n42), .A2(n43), .ZN(n39) );
  INV_X4 U91 ( .A(n44), .ZN(n42) );
  NOR2_X4 U92 ( .A1(n49), .A2(n44), .ZN(n48) );
  INV_X4 U93 ( .A(n26), .ZN(n49) );
  NAND2_X2 U94 ( .A1(n25), .A2(n28), .ZN(n46) );
  NAND2_X2 U95 ( .A1(n27), .A2(n50), .ZN(n45) );
  NOR2_X4 U96 ( .A1(n53), .A2(n54), .ZN(n52) );
  NAND2_X2 U97 ( .A1(n42), .A2(n55), .ZN(n51) );
  AOI21_X4 U98 ( .B1(n56), .B2(n57), .A(n58), .ZN(B[1]) );
  NOR2_X4 U99 ( .A1(n59), .A2(n60), .ZN(n57) );
  NAND2_X2 U100 ( .A1(n62), .A2(n63), .ZN(n37) );
  NAND2_X2 U101 ( .A1(n62), .A2(n64), .ZN(n44) );
  NOR2_X4 U102 ( .A1(n2), .A2(n65), .ZN(n56) );
  NAND2_X2 U103 ( .A1(A[4]), .A2(n61), .ZN(n67) );
  INV_X4 U104 ( .A(n68), .ZN(n61) );
  NAND2_X2 U105 ( .A1(A[3]), .A2(n69), .ZN(n66) );
  INV_X4 U106 ( .A(n71), .ZN(B[13]) );
  INV_X4 U107 ( .A(n63), .ZN(n13) );
  INV_X4 U108 ( .A(A[13]), .ZN(n74) );
  NAND2_X2 U109 ( .A1(A[11]), .A2(n69), .ZN(n78) );
  NAND2_X2 U110 ( .A1(A[10]), .A2(n130), .ZN(n77) );
  NAND2_X2 U111 ( .A1(A[12]), .A2(n79), .ZN(n76) );
  INV_X4 U112 ( .A(n68), .ZN(n79) );
  NOR3_X4 U113 ( .A1(n4), .A2(n80), .A3(n81), .ZN(n7) );
  NAND2_X2 U114 ( .A1(n82), .A2(n83), .ZN(n81) );
  INV_X4 U115 ( .A(n84), .ZN(n80) );
  INV_X4 U116 ( .A(n43), .ZN(n20) );
  INV_X4 U117 ( .A(n88), .ZN(n19) );
  NOR2_X4 U118 ( .A1(n92), .A2(n93), .ZN(n91) );
  NOR2_X4 U119 ( .A1(n68), .A2(n94), .ZN(n93) );
  INV_X4 U120 ( .A(A[11]), .ZN(n94) );
  INV_X4 U121 ( .A(n95), .ZN(n92) );
  NAND2_X2 U122 ( .A1(A[9]), .A2(n130), .ZN(n90) );
  NAND4_X2 U123 ( .A1(n97), .A2(n98), .A3(n99), .A4(n100), .ZN(n50) );
  NAND2_X2 U124 ( .A1(A[5]), .A2(n69), .ZN(n100) );
  NAND2_X2 U125 ( .A1(A[6]), .A2(n61), .ZN(n98) );
  NAND4_X2 U126 ( .A1(n101), .A2(n102), .A3(n103), .A4(n104), .ZN(n28) );
  NAND2_X2 U127 ( .A1(A[9]), .A2(n69), .ZN(n104) );
  NAND2_X2 U128 ( .A1(A[10]), .A2(n105), .ZN(n102) );
  INV_X4 U129 ( .A(n68), .ZN(n105) );
  NAND2_X2 U130 ( .A1(n27), .A2(n26), .ZN(n96) );
  NAND2_X2 U131 ( .A1(A[13]), .A2(n69), .ZN(n108) );
  NAND2_X2 U132 ( .A1(A[12]), .A2(n130), .ZN(n107) );
  NAND2_X2 U133 ( .A1(A[11]), .A2(n24), .ZN(n106) );
  INV_X4 U134 ( .A(n55), .ZN(n33) );
  NAND4_X2 U135 ( .A1(n110), .A2(n111), .A3(n112), .A4(n113), .ZN(n55) );
  NAND2_X2 U136 ( .A1(A[12]), .A2(n69), .ZN(n113) );
  NAND2_X2 U137 ( .A1(A[13]), .A2(n114), .ZN(n111) );
  INV_X4 U138 ( .A(n68), .ZN(n114) );
  INV_X4 U139 ( .A(n115), .ZN(n32) );
  NAND4_X2 U140 ( .A1(n116), .A2(n117), .A3(n118), .A4(n119), .ZN(n115) );
  NAND2_X2 U141 ( .A1(A[8]), .A2(n69), .ZN(n119) );
  NAND2_X2 U142 ( .A1(A[9]), .A2(n61), .ZN(n117) );
  INV_X4 U143 ( .A(SH[2]), .ZN(n64) );
  NAND2_X2 U144 ( .A1(A[4]), .A2(n69), .ZN(n122) );
  NAND2_X2 U145 ( .A1(A[5]), .A2(n114), .ZN(n120) );
  NAND2_X2 U146 ( .A1(n123), .A2(n124), .ZN(B[0]) );
  NAND2_X2 U147 ( .A1(n125), .A2(n62), .ZN(n124) );
  INV_X4 U148 ( .A(n134), .ZN(n62) );
  MUX2_X2 U149 ( .A(n126), .B(n127), .S(SH[2]), .Z(n125) );
  NAND4_X2 U150 ( .A1(n128), .A2(n129), .A3(n89), .A4(n95), .ZN(n126) );
  NAND2_X2 U151 ( .A1(A[11]), .A2(n105), .ZN(n128) );
  NAND2_X2 U152 ( .A1(A[6]), .A2(n69), .ZN(n138) );
  NAND2_X2 U153 ( .A1(SH[1]), .A2(n140), .ZN(n139) );
  NAND2_X2 U154 ( .A1(A[7]), .A2(n79), .ZN(n136) );
=======
  FA_X1 S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA_X1 S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA_X1 S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA_X1 S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA_X1 S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA_X1 S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA_X1 S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), 
        .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA_X1 S2_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .CI(\SUMB[2][16] ), 
        .CO(\CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FA_X1 S2_3_16 ( .A(\ab[3][16] ), .B(\CARRYB[2][16] ), .CI(\SUMB[2][17] ), 
        .CO(\CARRYB[3][16] ), .S(\SUMB[3][16] ) );
  FA_X1 S2_3_17 ( .A(\ab[3][17] ), .B(\CARRYB[2][17] ), .CI(\SUMB[2][18] ), 
        .CO(\CARRYB[3][17] ), .S(\SUMB[3][17] ) );
  FA_X1 S2_3_18 ( .A(\ab[3][18] ), .B(\CARRYB[2][18] ), .CI(\SUMB[2][19] ), 
        .CO(\CARRYB[3][18] ), .S(\SUMB[3][18] ) );
  FA_X1 S2_3_19 ( .A(\ab[3][19] ), .B(\CARRYB[2][19] ), .CI(\SUMB[2][20] ), 
        .CO(\CARRYB[3][19] ), .S(\SUMB[3][19] ) );
  FA_X1 S2_3_20 ( .A(\ab[3][20] ), .B(\CARRYB[2][20] ), .CI(\SUMB[2][21] ), 
        .CO(\CARRYB[3][20] ), .S(\SUMB[3][20] ) );
  FA_X1 S2_3_21 ( .A(\ab[3][21] ), .B(\CARRYB[2][21] ), .CI(\SUMB[2][22] ), 
        .CO(\CARRYB[3][21] ), .S(\SUMB[3][21] ) );
  FA_X1 S2_3_22 ( .A(\ab[3][22] ), .B(\CARRYB[2][22] ), .CI(\SUMB[2][23] ), 
        .CO(\CARRYB[3][22] ), .S(\SUMB[3][22] ) );
  FA_X1 S2_3_23 ( .A(\ab[3][23] ), .B(\CARRYB[2][23] ), .CI(\SUMB[2][24] ), 
        .CO(\CARRYB[3][23] ), .S(\SUMB[3][23] ) );
  FA_X1 S2_3_24 ( .A(\ab[3][24] ), .B(\CARRYB[2][24] ), .CI(\SUMB[2][25] ), 
        .CO(\CARRYB[3][24] ), .S(\SUMB[3][24] ) );
  FA_X1 S2_3_25 ( .A(\ab[3][25] ), .B(\CARRYB[2][25] ), .CI(\SUMB[2][26] ), 
        .CO(\CARRYB[3][25] ), .S(\SUMB[3][25] ) );
  FA_X1 S2_3_26 ( .A(\ab[3][26] ), .B(\CARRYB[2][26] ), .CI(\SUMB[2][27] ), 
        .CO(\CARRYB[3][26] ), .S(\SUMB[3][26] ) );
  FA_X1 S2_3_27 ( .A(\ab[3][27] ), .B(\CARRYB[2][27] ), .CI(\SUMB[2][28] ), 
        .CO(\CARRYB[3][27] ), .S(\SUMB[3][27] ) );
  FA_X1 S2_3_28 ( .A(\ab[3][28] ), .B(\CARRYB[2][28] ), .CI(\SUMB[2][29] ), 
        .CO(\CARRYB[3][28] ), .S(\SUMB[3][28] ) );
  FA_X1 S2_3_29 ( .A(\ab[3][29] ), .B(\CARRYB[2][29] ), .CI(\SUMB[2][30] ), 
        .CO(\CARRYB[3][29] ), .S(\SUMB[3][29] ) );
  FA_X1 S2_3_30 ( .A(\ab[3][30] ), .B(\CARRYB[2][30] ), .CI(\SUMB[2][31] ), 
        .CO(\CARRYB[3][30] ), .S(\SUMB[3][30] ) );
  FA_X1 S2_3_31 ( .A(\ab[3][31] ), .B(\CARRYB[2][31] ), .CI(\SUMB[2][32] ), 
        .CO(\CARRYB[3][31] ), .S(\SUMB[3][31] ) );
  FA_X1 S2_3_32 ( .A(\ab[3][32] ), .B(\CARRYB[2][32] ), .CI(\SUMB[2][33] ), 
        .CO(\CARRYB[3][32] ), .S(\SUMB[3][32] ) );
  FA_X1 S2_3_33 ( .A(\ab[3][33] ), .B(\CARRYB[2][33] ), .CI(\SUMB[2][34] ), 
        .CO(\CARRYB[3][33] ), .S(\SUMB[3][33] ) );
  FA_X1 S2_3_34 ( .A(\ab[3][34] ), .B(\CARRYB[2][34] ), .CI(\SUMB[2][35] ), 
        .CO(\CARRYB[3][34] ), .S(\SUMB[3][34] ) );
  FA_X1 S2_3_35 ( .A(\ab[3][35] ), .B(\CARRYB[2][35] ), .CI(\SUMB[2][36] ), 
        .CO(\CARRYB[3][35] ), .S(\SUMB[3][35] ) );
  FA_X1 S2_3_36 ( .A(\ab[3][36] ), .B(\CARRYB[2][36] ), .CI(\SUMB[2][37] ), 
        .CO(\CARRYB[3][36] ), .S(\SUMB[3][36] ) );
  FA_X1 S2_3_37 ( .A(\ab[3][37] ), .B(\CARRYB[2][37] ), .CI(\SUMB[2][38] ), 
        .CO(\CARRYB[3][37] ), .S(\SUMB[3][37] ) );
  FA_X1 S2_3_38 ( .A(\ab[3][38] ), .B(\CARRYB[2][38] ), .CI(\SUMB[2][39] ), 
        .CO(\CARRYB[3][38] ), .S(\SUMB[3][38] ) );
  FA_X1 S2_3_39 ( .A(\ab[3][39] ), .B(\CARRYB[2][39] ), .CI(\SUMB[2][40] ), 
        .CO(\CARRYB[3][39] ), .S(\SUMB[3][39] ) );
  FA_X1 S2_3_40 ( .A(\ab[3][40] ), .B(\CARRYB[2][40] ), .CI(\SUMB[2][41] ), 
        .CO(\CARRYB[3][40] ), .S(\SUMB[3][40] ) );
  FA_X1 S2_3_41 ( .A(\ab[3][41] ), .B(\CARRYB[2][41] ), .CI(\SUMB[2][42] ), 
        .CO(\CARRYB[3][41] ), .S(\SUMB[3][41] ) );
  FA_X1 S2_3_42 ( .A(\ab[3][42] ), .B(\CARRYB[2][42] ), .CI(\SUMB[2][43] ), 
        .CO(\CARRYB[3][42] ), .S(\SUMB[3][42] ) );
  FA_X1 S2_3_43 ( .A(\ab[3][43] ), .B(\CARRYB[2][43] ), .CI(\SUMB[2][44] ), 
        .CO(\CARRYB[3][43] ), .S(\SUMB[3][43] ) );
  FA_X1 S2_3_44 ( .A(\ab[3][44] ), .B(\CARRYB[2][44] ), .CI(\SUMB[2][45] ), 
        .CO(\CARRYB[3][44] ), .S(\SUMB[3][44] ) );
  FA_X1 S2_3_45 ( .A(\ab[3][45] ), .B(\CARRYB[2][45] ), .CI(\SUMB[2][46] ), 
        .CO(\CARRYB[3][45] ), .S(\SUMB[3][45] ) );
  FA_X1 S2_3_46 ( .A(\ab[3][46] ), .B(\CARRYB[2][46] ), .CI(\SUMB[2][47] ), 
        .CO(\CARRYB[3][46] ), .S(\SUMB[3][46] ) );
  FA_X1 S2_3_47 ( .A(\ab[3][47] ), .B(\CARRYB[2][47] ), .CI(\SUMB[2][48] ), 
        .CO(\CARRYB[3][47] ), .S(\SUMB[3][47] ) );
  FA_X1 S2_3_48 ( .A(\ab[3][48] ), .B(\CARRYB[2][48] ), .CI(\SUMB[2][49] ), 
        .CO(\CARRYB[3][48] ), .S(\SUMB[3][48] ) );
  FA_X1 S2_3_49 ( .A(\ab[3][49] ), .B(\CARRYB[2][49] ), .CI(\SUMB[2][50] ), 
        .CO(\CARRYB[3][49] ), .S(\SUMB[3][49] ) );
  FA_X1 S2_3_50 ( .A(\ab[3][50] ), .B(\CARRYB[2][50] ), .CI(\SUMB[2][51] ), 
        .CO(\CARRYB[3][50] ), .S(\SUMB[3][50] ) );
  FA_X1 S3_3_51 ( .A(\ab[3][51] ), .B(\CARRYB[2][51] ), .CI(\ab[2][52] ), .CO(
        \CARRYB[3][51] ), .S(\SUMB[3][51] ) );
  FA_X1 S1_2_0 ( .A(\ab[2][0] ), .B(n72), .CI(n171), .CO(\CARRYB[2][0] ), .S(
        CLA_SUM[2]) );
  FA_X1 S2_2_1 ( .A(\ab[2][1] ), .B(n29), .CI(n158), .CO(\CARRYB[2][1] ), .S(
        \SUMB[2][1] ) );
  FA_X1 S2_2_2 ( .A(\ab[2][2] ), .B(n28), .CI(n157), .CO(\CARRYB[2][2] ), .S(
        \SUMB[2][2] ) );
  FA_X1 S2_2_3 ( .A(\ab[2][3] ), .B(n33), .CI(n156), .CO(\CARRYB[2][3] ), .S(
        \SUMB[2][3] ) );
  FA_X1 S2_2_4 ( .A(\ab[2][4] ), .B(n32), .CI(n155), .CO(\CARRYB[2][4] ), .S(
        \SUMB[2][4] ) );
  FA_X1 S2_2_5 ( .A(\ab[2][5] ), .B(n55), .CI(n154), .CO(\CARRYB[2][5] ), .S(
        \SUMB[2][5] ) );
  FA_X1 S2_2_6 ( .A(\ab[2][6] ), .B(n31), .CI(n153), .CO(\CARRYB[2][6] ), .S(
        \SUMB[2][6] ) );
  FA_X1 S2_2_7 ( .A(\ab[2][7] ), .B(n54), .CI(n152), .CO(\CARRYB[2][7] ), .S(
        \SUMB[2][7] ) );
  FA_X1 S2_2_8 ( .A(\ab[2][8] ), .B(n30), .CI(n151), .CO(\CARRYB[2][8] ), .S(
        \SUMB[2][8] ) );
  FA_X1 S2_2_9 ( .A(\ab[2][9] ), .B(n53), .CI(n150), .CO(\CARRYB[2][9] ), .S(
        \SUMB[2][9] ) );
  FA_X1 S2_2_10 ( .A(\ab[2][10] ), .B(n52), .CI(n149), .CO(\CARRYB[2][10] ), 
        .S(\SUMB[2][10] ) );
  FA_X1 S2_2_11 ( .A(\ab[2][11] ), .B(n51), .CI(n148), .CO(\CARRYB[2][11] ), 
        .S(\SUMB[2][11] ) );
  FA_X1 S2_2_12 ( .A(\ab[2][12] ), .B(n50), .CI(n147), .CO(\CARRYB[2][12] ), 
        .S(\SUMB[2][12] ) );
  FA_X1 S2_2_13 ( .A(\ab[2][13] ), .B(n49), .CI(n146), .CO(\CARRYB[2][13] ), 
        .S(\SUMB[2][13] ) );
  FA_X1 S2_2_14 ( .A(\ab[2][14] ), .B(n48), .CI(n145), .CO(\CARRYB[2][14] ), 
        .S(\SUMB[2][14] ) );
  FA_X1 S2_2_15 ( .A(\ab[2][15] ), .B(n47), .CI(n144), .CO(\CARRYB[2][15] ), 
        .S(\SUMB[2][15] ) );
  FA_X1 S2_2_16 ( .A(\ab[2][16] ), .B(n46), .CI(n143), .CO(\CARRYB[2][16] ), 
        .S(\SUMB[2][16] ) );
  FA_X1 S2_2_17 ( .A(\ab[2][17] ), .B(n45), .CI(n142), .CO(\CARRYB[2][17] ), 
        .S(\SUMB[2][17] ) );
  FA_X1 S2_2_18 ( .A(\ab[2][18] ), .B(n44), .CI(n141), .CO(\CARRYB[2][18] ), 
        .S(\SUMB[2][18] ) );
  FA_X1 S2_2_19 ( .A(\ab[2][19] ), .B(n43), .CI(n140), .CO(\CARRYB[2][19] ), 
        .S(\SUMB[2][19] ) );
  FA_X1 S2_2_20 ( .A(\ab[2][20] ), .B(n42), .CI(n139), .CO(\CARRYB[2][20] ), 
        .S(\SUMB[2][20] ) );
  FA_X1 S2_2_21 ( .A(\ab[2][21] ), .B(n41), .CI(n138), .CO(\CARRYB[2][21] ), 
        .S(\SUMB[2][21] ) );
  FA_X1 S2_2_22 ( .A(\ab[2][22] ), .B(n40), .CI(n137), .CO(\CARRYB[2][22] ), 
        .S(\SUMB[2][22] ) );
  FA_X1 S2_2_23 ( .A(\ab[2][23] ), .B(n39), .CI(n136), .CO(\CARRYB[2][23] ), 
        .S(\SUMB[2][23] ) );
  FA_X1 S2_2_24 ( .A(\ab[2][24] ), .B(n38), .CI(n135), .CO(\CARRYB[2][24] ), 
        .S(\SUMB[2][24] ) );
  FA_X1 S2_2_25 ( .A(\ab[2][25] ), .B(n37), .CI(n134), .CO(\CARRYB[2][25] ), 
        .S(\SUMB[2][25] ) );
  FA_X1 S2_2_26 ( .A(\ab[2][26] ), .B(n36), .CI(n133), .CO(\CARRYB[2][26] ), 
        .S(\SUMB[2][26] ) );
  FA_X1 S2_2_27 ( .A(\ab[2][27] ), .B(n35), .CI(n132), .CO(\CARRYB[2][27] ), 
        .S(\SUMB[2][27] ) );
  FA_X1 S2_2_28 ( .A(\ab[2][28] ), .B(n34), .CI(n131), .CO(\CARRYB[2][28] ), 
        .S(\SUMB[2][28] ) );
  FA_X1 S2_2_29 ( .A(\ab[2][29] ), .B(n27), .CI(n130), .CO(\CARRYB[2][29] ), 
        .S(\SUMB[2][29] ) );
  FA_X1 S2_2_30 ( .A(\ab[2][30] ), .B(n26), .CI(n129), .CO(\CARRYB[2][30] ), 
        .S(\SUMB[2][30] ) );
  FA_X1 S2_2_31 ( .A(\ab[2][31] ), .B(n25), .CI(n128), .CO(\CARRYB[2][31] ), 
        .S(\SUMB[2][31] ) );
  FA_X1 S2_2_32 ( .A(\ab[2][32] ), .B(n24), .CI(n127), .CO(\CARRYB[2][32] ), 
        .S(\SUMB[2][32] ) );
  FA_X1 S2_2_33 ( .A(\ab[2][33] ), .B(n23), .CI(n126), .CO(\CARRYB[2][33] ), 
        .S(\SUMB[2][33] ) );
  FA_X1 S2_2_34 ( .A(\ab[2][34] ), .B(n22), .CI(n125), .CO(\CARRYB[2][34] ), 
        .S(\SUMB[2][34] ) );
  FA_X1 S2_2_35 ( .A(\ab[2][35] ), .B(n21), .CI(n124), .CO(\CARRYB[2][35] ), 
        .S(\SUMB[2][35] ) );
  FA_X1 S2_2_36 ( .A(\ab[2][36] ), .B(n20), .CI(n123), .CO(\CARRYB[2][36] ), 
        .S(\SUMB[2][36] ) );
  FA_X1 S2_2_37 ( .A(\ab[2][37] ), .B(n19), .CI(n122), .CO(\CARRYB[2][37] ), 
        .S(\SUMB[2][37] ) );
  FA_X1 S2_2_38 ( .A(\ab[2][38] ), .B(n18), .CI(n121), .CO(\CARRYB[2][38] ), 
        .S(\SUMB[2][38] ) );
  FA_X1 S2_2_39 ( .A(\ab[2][39] ), .B(n17), .CI(n120), .CO(\CARRYB[2][39] ), 
        .S(\SUMB[2][39] ) );
  FA_X1 S2_2_40 ( .A(\ab[2][40] ), .B(n16), .CI(n119), .CO(\CARRYB[2][40] ), 
        .S(\SUMB[2][40] ) );
  FA_X1 S2_2_41 ( .A(\ab[2][41] ), .B(n15), .CI(n118), .CO(\CARRYB[2][41] ), 
        .S(\SUMB[2][41] ) );
  FA_X1 S2_2_42 ( .A(\ab[2][42] ), .B(n14), .CI(n117), .CO(\CARRYB[2][42] ), 
        .S(\SUMB[2][42] ) );
  FA_X1 S2_2_43 ( .A(\ab[2][43] ), .B(n13), .CI(n116), .CO(\CARRYB[2][43] ), 
        .S(\SUMB[2][43] ) );
  FA_X1 S2_2_44 ( .A(\ab[2][44] ), .B(n12), .CI(n115), .CO(\CARRYB[2][44] ), 
        .S(\SUMB[2][44] ) );
  FA_X1 S2_2_45 ( .A(\ab[2][45] ), .B(n11), .CI(n114), .CO(\CARRYB[2][45] ), 
        .S(\SUMB[2][45] ) );
  FA_X1 S2_2_46 ( .A(\ab[2][46] ), .B(n10), .CI(n113), .CO(\CARRYB[2][46] ), 
        .S(\SUMB[2][46] ) );
  FA_X1 S2_2_47 ( .A(\ab[2][47] ), .B(n9), .CI(n112), .CO(\CARRYB[2][47] ), 
        .S(\SUMB[2][47] ) );
  FA_X1 S2_2_48 ( .A(\ab[2][48] ), .B(n8), .CI(n111), .CO(\CARRYB[2][48] ), 
        .S(\SUMB[2][48] ) );
  FA_X1 S2_2_49 ( .A(\ab[2][49] ), .B(n3), .CI(n110), .CO(\CARRYB[2][49] ), 
        .S(\SUMB[2][49] ) );
  FA_X1 S2_2_50 ( .A(\ab[2][50] ), .B(n109), .CI(n4), .CO(\CARRYB[2][50] ), 
        .S(\SUMB[2][50] ) );
  FA_X1 S3_2_51 ( .A(\ab[2][51] ), .B(n105), .CI(\ab[1][52] ), .CO(
        \CARRYB[2][51] ), .S(\SUMB[2][51] ) );
  fpu_DW01_add_8 FS_1 ( .A({1'b0, n94, n95, n104, n96, n103, n99, n100, n102, 
        n97, n101, n98, n81, n80, n79, n78, n93, n76, n92, n91, n90, n77, n89, 
        n88, n75, n82, n74, n83, n86, n73, n85, n84, n87, n60, n71, n70, n69, 
        n66, n68, n67, n57, n65, n56, n64, n63, n59, n62, n58, n61, n7, n5, n6, 
        n207, \SUMB[52][0] , CLA_SUM}), .B({n208, n209, n196, n206, n197, n205, 
        n200, n201, n204, n198, n203, n199, n202, n180, n179, n178, n195, n177, 
        n194, n193, n192, n173, n191, n190, n176, n181, n175, n182, n185, n174, 
        n184, n183, n189, n172, n188, n187, n186, n168, n170, n169, n162, n167, 
        n161, n166, n165, n160, n164, n159, n163, n108, n106, n107, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM(PRODUCT[105:2]) );
  INV_X4 U2 ( .A(A[9]), .ZN(n311) );
  INV_X4 U3 ( .A(A[13]), .ZN(n305) );
  INV_X4 U4 ( .A(A[12]), .ZN(n307) );
  INV_X4 U5 ( .A(B[20]), .ZN(n403) );
  INV_X4 U6 ( .A(A[15]), .ZN(n302) );
  INV_X4 U7 ( .A(A[16]), .ZN(n300) );
  INV_X4 U8 ( .A(B[52]), .ZN(n336) );
  INV_X4 U9 ( .A(B[25]), .ZN(n393) );
  INV_X4 U10 ( .A(B[23]), .ZN(n397) );
  INV_X4 U11 ( .A(B[29]), .ZN(n385) );
  INV_X4 U12 ( .A(A[6]), .ZN(n317) );
  INV_X4 U13 ( .A(B[6]), .ZN(n434) );
  INV_X4 U14 ( .A(B[4]), .ZN(n438) );
  INV_X4 U15 ( .A(B[9]), .ZN(n428) );
  INV_X4 U16 ( .A(B[7]), .ZN(n432) );
  INV_X4 U17 ( .A(B[26]), .ZN(n391) );
  INV_X4 U18 ( .A(B[24]), .ZN(n395) );
  INV_X4 U19 ( .A(B[27]), .ZN(n389) );
  INV_X4 U20 ( .A(B[17]), .ZN(n408) );
  INV_X4 U21 ( .A(B[11]), .ZN(n425) );
  INV_X4 U22 ( .A(B[22]), .ZN(n399) );
  INV_X4 U23 ( .A(B[21]), .ZN(n401) );
  INV_X4 U24 ( .A(B[5]), .ZN(n436) );
  INV_X4 U25 ( .A(B[28]), .ZN(n387) );
  INV_X4 U26 ( .A(B[0]), .ZN(n446) );
  INV_X4 U27 ( .A(A[14]), .ZN(n303) );
  INV_X4 U28 ( .A(A[25]), .ZN(n282) );
  INV_X4 U29 ( .A(B[8]), .ZN(n430) );
  INV_X4 U30 ( .A(B[51]), .ZN(n338) );
  INV_X4 U31 ( .A(B[18]), .ZN(n406) );
  INV_X4 U32 ( .A(B[39]), .ZN(n365) );
  INV_X4 U33 ( .A(B[33]), .ZN(n377) );
  INV_X4 U34 ( .A(B[45]), .ZN(n351) );
  INV_X4 U35 ( .A(B[40]), .ZN(n363) );
  INV_X4 U36 ( .A(B[31]), .ZN(n381) );
  INV_X4 U37 ( .A(B[46]), .ZN(n349) );
  INV_X4 U38 ( .A(B[41]), .ZN(n361) );
  INV_X4 U39 ( .A(B[30]), .ZN(n383) );
  INV_X4 U40 ( .A(B[47]), .ZN(n347) );
  INV_X4 U41 ( .A(B[48]), .ZN(n345) );
  INV_X4 U42 ( .A(B[35]), .ZN(n373) );
  INV_X4 U43 ( .A(B[13]), .ZN(n419) );
  INV_X4 U44 ( .A(B[14]), .ZN(n416) );
  INV_X4 U45 ( .A(B[12]), .ZN(n422) );
  INV_X4 U46 ( .A(B[44]), .ZN(n353) );
  INV_X4 U47 ( .A(B[42]), .ZN(n358) );
  INV_X4 U48 ( .A(B[37]), .ZN(n370) );
  INV_X4 U49 ( .A(B[32]), .ZN(n380) );
  INV_X4 U50 ( .A(B[16]), .ZN(n410) );
  INV_X4 U51 ( .A(B[15]), .ZN(n413) );
  INV_X4 U52 ( .A(B[10]), .ZN(n427) );
  INV_X4 U53 ( .A(B[3]), .ZN(n440) );
  INV_X4 U54 ( .A(B[4]), .ZN(n439) );
  INV_X4 U55 ( .A(B[6]), .ZN(n435) );
  INV_X4 U56 ( .A(B[5]), .ZN(n437) );
  INV_X4 U57 ( .A(A[7]), .ZN(n315) );
  INV_X4 U58 ( .A(A[19]), .ZN(n293) );
  INV_X4 U59 ( .A(A[20]), .ZN(n292) );
  INV_X4 U60 ( .A(A[23]), .ZN(n286) );
  INV_X4 U61 ( .A(A[24]), .ZN(n284) );
  INV_X4 U62 ( .A(A[22]), .ZN(n288) );
  INV_X4 U63 ( .A(A[21]), .ZN(n290) );
  INV_X4 U64 ( .A(A[29]), .ZN(n274) );
  INV_X4 U65 ( .A(A[1]), .ZN(n330) );
  INV_X4 U66 ( .A(A[5]), .ZN(n319) );
  INV_X4 U67 ( .A(B[51]), .ZN(n340) );
  INV_X4 U68 ( .A(B[51]), .ZN(n339) );
  INV_X4 U69 ( .A(B[49]), .ZN(n343) );
  INV_X4 U70 ( .A(B[43]), .ZN(n356) );
  INV_X4 U71 ( .A(B[34]), .ZN(n375) );
  INV_X4 U72 ( .A(B[52]), .ZN(n337) );
  INV_X4 U73 ( .A(B[50]), .ZN(n341) );
  INV_X4 U74 ( .A(B[19]), .ZN(n404) );
  INV_X4 U75 ( .A(B[36]), .ZN(n372) );
  INV_X4 U76 ( .A(B[32]), .ZN(n379) );
  INV_X4 U77 ( .A(B[17]), .ZN(n409) );
  INV_X4 U78 ( .A(B[11]), .ZN(n426) );
  INV_X4 U79 ( .A(B[38]), .ZN(n369) );
  INV_X4 U80 ( .A(A[6]), .ZN(n316) );
  INV_X4 U81 ( .A(B[8]), .ZN(n431) );
  INV_X4 U82 ( .A(B[9]), .ZN(n429) );
  INV_X4 U83 ( .A(B[7]), .ZN(n433) );
  INV_X4 U84 ( .A(B[2]), .ZN(n442) );
  INV_X4 U85 ( .A(A[18]), .ZN(n296) );
  INV_X4 U86 ( .A(A[26]), .ZN(n281) );
  INV_X4 U87 ( .A(A[28]), .ZN(n277) );
  INV_X4 U88 ( .A(A[31]), .ZN(n269) );
  INV_X4 U89 ( .A(A[35]), .ZN(n261) );
  INV_X4 U90 ( .A(n454), .ZN(n235) );
  INV_X4 U91 ( .A(A[39]), .ZN(n248) );
  INV_X4 U92 ( .A(A[41]), .ZN(n243) );
  INV_X4 U93 ( .A(A[52]), .ZN(n449) );
  INV_X4 U94 ( .A(A[50]), .ZN(n214) );
  INV_X4 U95 ( .A(A[46]), .ZN(n224) );
  AND2_X4 U96 ( .A1(\ab[0][50] ), .A2(\ab[1][49] ), .ZN(n3) );
  XOR2_X2 U97 ( .A(\ab[1][51] ), .B(\ab[0][52] ), .Z(n4) );
  XOR2_X2 U98 ( .A(\CARRYB[52][2] ), .B(\SUMB[52][3] ), .Z(n5) );
  XOR2_X2 U99 ( .A(\CARRYB[52][1] ), .B(\SUMB[52][2] ), .Z(n6) );
  XOR2_X2 U100 ( .A(\CARRYB[52][3] ), .B(\SUMB[52][4] ), .Z(n7) );
  AND2_X4 U101 ( .A1(\ab[0][49] ), .A2(\ab[1][48] ), .ZN(n8) );
  AND2_X4 U102 ( .A1(\ab[0][48] ), .A2(\ab[1][47] ), .ZN(n9) );
  AND2_X4 U103 ( .A1(\ab[0][47] ), .A2(\ab[1][46] ), .ZN(n10) );
  AND2_X4 U104 ( .A1(\ab[0][46] ), .A2(\ab[1][45] ), .ZN(n11) );
  AND2_X4 U105 ( .A1(\ab[0][45] ), .A2(\ab[1][44] ), .ZN(n12) );
  AND2_X4 U106 ( .A1(\ab[0][44] ), .A2(\ab[1][43] ), .ZN(n13) );
  AND2_X4 U107 ( .A1(\ab[0][43] ), .A2(\ab[1][42] ), .ZN(n14) );
  AND2_X4 U108 ( .A1(\ab[0][42] ), .A2(\ab[1][41] ), .ZN(n15) );
  AND2_X4 U109 ( .A1(\ab[0][41] ), .A2(\ab[1][40] ), .ZN(n16) );
  AND2_X4 U110 ( .A1(\ab[0][40] ), .A2(\ab[1][39] ), .ZN(n17) );
  AND2_X4 U111 ( .A1(\ab[0][39] ), .A2(\ab[1][38] ), .ZN(n18) );
  AND2_X4 U112 ( .A1(\ab[0][38] ), .A2(\ab[1][37] ), .ZN(n19) );
  AND2_X4 U113 ( .A1(\ab[0][37] ), .A2(\ab[1][36] ), .ZN(n20) );
  AND2_X4 U114 ( .A1(\ab[0][36] ), .A2(\ab[1][35] ), .ZN(n21) );
  AND2_X4 U115 ( .A1(\ab[0][35] ), .A2(\ab[1][34] ), .ZN(n22) );
  AND2_X4 U116 ( .A1(\ab[0][34] ), .A2(\ab[1][33] ), .ZN(n23) );
  AND2_X4 U117 ( .A1(\ab[0][33] ), .A2(\ab[1][32] ), .ZN(n24) );
  AND2_X4 U118 ( .A1(\ab[0][32] ), .A2(\ab[1][31] ), .ZN(n25) );
  AND2_X4 U119 ( .A1(\ab[0][31] ), .A2(\ab[1][30] ), .ZN(n26) );
  AND2_X4 U120 ( .A1(\ab[0][30] ), .A2(\ab[1][29] ), .ZN(n27) );
  AND2_X4 U121 ( .A1(\ab[0][3] ), .A2(\ab[1][2] ), .ZN(n28) );
  AND2_X4 U122 ( .A1(\ab[0][2] ), .A2(\ab[1][1] ), .ZN(n29) );
  AND2_X4 U123 ( .A1(\ab[0][9] ), .A2(\ab[1][8] ), .ZN(n30) );
  AND2_X4 U124 ( .A1(\ab[0][7] ), .A2(\ab[1][6] ), .ZN(n31) );
  AND2_X4 U125 ( .A1(\ab[0][5] ), .A2(\ab[1][4] ), .ZN(n32) );
  AND2_X4 U126 ( .A1(\ab[0][4] ), .A2(\ab[1][3] ), .ZN(n33) );
  AND2_X4 U127 ( .A1(\ab[0][29] ), .A2(\ab[1][28] ), .ZN(n34) );
  AND2_X4 U128 ( .A1(\ab[0][28] ), .A2(\ab[1][27] ), .ZN(n35) );
  AND2_X4 U129 ( .A1(\ab[0][27] ), .A2(\ab[1][26] ), .ZN(n36) );
  AND2_X4 U130 ( .A1(\ab[0][26] ), .A2(\ab[1][25] ), .ZN(n37) );
  AND2_X4 U131 ( .A1(\ab[0][25] ), .A2(\ab[1][24] ), .ZN(n38) );
  AND2_X4 U132 ( .A1(\ab[0][24] ), .A2(\ab[1][23] ), .ZN(n39) );
  AND2_X4 U133 ( .A1(\ab[0][23] ), .A2(\ab[1][22] ), .ZN(n40) );
  AND2_X4 U134 ( .A1(\ab[0][22] ), .A2(\ab[1][21] ), .ZN(n41) );
  AND2_X4 U135 ( .A1(\ab[0][21] ), .A2(\ab[1][20] ), .ZN(n42) );
  AND2_X4 U136 ( .A1(\ab[0][20] ), .A2(\ab[1][19] ), .ZN(n43) );
  AND2_X4 U137 ( .A1(\ab[0][19] ), .A2(\ab[1][18] ), .ZN(n44) );
  AND2_X4 U138 ( .A1(\ab[0][18] ), .A2(\ab[1][17] ), .ZN(n45) );
  AND2_X4 U139 ( .A1(\ab[0][17] ), .A2(\ab[1][16] ), .ZN(n46) );
  AND2_X4 U140 ( .A1(\ab[0][16] ), .A2(\ab[1][15] ), .ZN(n47) );
  AND2_X4 U141 ( .A1(\ab[0][15] ), .A2(\ab[1][14] ), .ZN(n48) );
  AND2_X4 U142 ( .A1(\ab[0][14] ), .A2(\ab[1][13] ), .ZN(n49) );
  AND2_X4 U143 ( .A1(\ab[0][13] ), .A2(\ab[1][12] ), .ZN(n50) );
  AND2_X4 U144 ( .A1(\ab[0][12] ), .A2(\ab[1][11] ), .ZN(n51) );
  AND2_X4 U145 ( .A1(\ab[0][11] ), .A2(\ab[1][10] ), .ZN(n52) );
  AND2_X4 U146 ( .A1(\ab[0][10] ), .A2(\ab[1][9] ), .ZN(n53) );
  AND2_X4 U147 ( .A1(\ab[0][8] ), .A2(\ab[1][7] ), .ZN(n54) );
  AND2_X4 U148 ( .A1(\ab[0][6] ), .A2(\ab[1][5] ), .ZN(n55) );
  XOR2_X2 U149 ( .A(\CARRYB[52][10] ), .B(\SUMB[52][11] ), .Z(n56) );
  XOR2_X2 U150 ( .A(\CARRYB[52][12] ), .B(\SUMB[52][13] ), .Z(n57) );
  XOR2_X2 U151 ( .A(\CARRYB[52][5] ), .B(\SUMB[52][6] ), .Z(n58) );
  XOR2_X2 U152 ( .A(\CARRYB[52][7] ), .B(\SUMB[52][8] ), .Z(n59) );
  XOR2_X2 U153 ( .A(\CARRYB[52][19] ), .B(\SUMB[52][20] ), .Z(n60) );
  XOR2_X2 U154 ( .A(\CARRYB[52][4] ), .B(\SUMB[52][5] ), .Z(n61) );
  XOR2_X2 U155 ( .A(\CARRYB[52][6] ), .B(\SUMB[52][7] ), .Z(n62) );
  XOR2_X2 U156 ( .A(\CARRYB[52][8] ), .B(\SUMB[52][9] ), .Z(n63) );
  XOR2_X2 U157 ( .A(\CARRYB[52][9] ), .B(\SUMB[52][10] ), .Z(n64) );
  XOR2_X2 U158 ( .A(\CARRYB[52][11] ), .B(\SUMB[52][12] ), .Z(n65) );
  XOR2_X2 U159 ( .A(\CARRYB[52][15] ), .B(\SUMB[52][16] ), .Z(n66) );
  XOR2_X2 U160 ( .A(\CARRYB[52][13] ), .B(\SUMB[52][14] ), .Z(n67) );
  XOR2_X2 U161 ( .A(\CARRYB[52][14] ), .B(\SUMB[52][15] ), .Z(n68) );
  XOR2_X2 U162 ( .A(\CARRYB[52][16] ), .B(\SUMB[52][17] ), .Z(n69) );
  XOR2_X2 U163 ( .A(\CARRYB[52][17] ), .B(\SUMB[52][18] ), .Z(n70) );
  XOR2_X2 U164 ( .A(\CARRYB[52][18] ), .B(\SUMB[52][19] ), .Z(n71) );
  INV_X4 U165 ( .A(A[2]), .ZN(n327) );
  INV_X4 U166 ( .A(B[28]), .ZN(n388) );
  INV_X4 U167 ( .A(B[27]), .ZN(n390) );
  INV_X4 U168 ( .A(B[22]), .ZN(n400) );
  INV_X4 U169 ( .A(B[44]), .ZN(n355) );
  INV_X4 U170 ( .A(B[44]), .ZN(n354) );
  INV_X4 U171 ( .A(B[42]), .ZN(n360) );
  INV_X4 U172 ( .A(B[42]), .ZN(n359) );
  INV_X4 U173 ( .A(B[38]), .ZN(n368) );
  INV_X4 U174 ( .A(B[38]), .ZN(n367) );
  INV_X4 U175 ( .A(B[25]), .ZN(n394) );
  INV_X4 U176 ( .A(B[24]), .ZN(n396) );
  INV_X4 U177 ( .A(B[23]), .ZN(n398) );
  INV_X4 U178 ( .A(B[29]), .ZN(n386) );
  INV_X4 U179 ( .A(B[26]), .ZN(n392) );
  INV_X4 U180 ( .A(B[34]), .ZN(n376) );
  INV_X4 U181 ( .A(B[21]), .ZN(n402) );
  INV_X4 U182 ( .A(B[48]), .ZN(n346) );
  INV_X4 U183 ( .A(B[47]), .ZN(n348) );
  INV_X4 U184 ( .A(B[46]), .ZN(n350) );
  INV_X4 U185 ( .A(B[45]), .ZN(n352) );
  INV_X4 U186 ( .A(B[41]), .ZN(n362) );
  INV_X4 U187 ( .A(B[40]), .ZN(n364) );
  INV_X4 U188 ( .A(B[39]), .ZN(n366) );
  INV_X4 U189 ( .A(B[35]), .ZN(n374) );
  INV_X4 U190 ( .A(B[33]), .ZN(n378) );
  INV_X4 U191 ( .A(B[31]), .ZN(n382) );
  INV_X4 U192 ( .A(B[30]), .ZN(n384) );
  INV_X4 U193 ( .A(B[37]), .ZN(n371) );
  AND2_X4 U194 ( .A1(\ab[0][1] ), .A2(\ab[1][0] ), .ZN(n72) );
  XOR2_X2 U195 ( .A(\CARRYB[52][23] ), .B(\SUMB[52][24] ), .Z(n73) );
  XOR2_X2 U196 ( .A(\CARRYB[52][26] ), .B(\SUMB[52][27] ), .Z(n74) );
  XOR2_X2 U197 ( .A(\CARRYB[52][28] ), .B(\SUMB[52][29] ), .Z(n75) );
  XOR2_X2 U198 ( .A(\CARRYB[52][35] ), .B(\SUMB[52][36] ), .Z(n76) );
  XOR2_X2 U199 ( .A(\CARRYB[52][31] ), .B(\SUMB[52][32] ), .Z(n77) );
  XOR2_X2 U200 ( .A(\CARRYB[52][37] ), .B(\SUMB[52][38] ), .Z(n78) );
  XOR2_X2 U201 ( .A(\CARRYB[52][38] ), .B(\SUMB[52][39] ), .Z(n79) );
  XOR2_X2 U202 ( .A(\CARRYB[52][39] ), .B(\SUMB[52][40] ), .Z(n80) );
  XOR2_X2 U203 ( .A(\CARRYB[52][40] ), .B(\SUMB[52][41] ), .Z(n81) );
  XOR2_X2 U204 ( .A(\CARRYB[52][27] ), .B(\SUMB[52][28] ), .Z(n82) );
  XOR2_X2 U205 ( .A(\CARRYB[52][25] ), .B(\SUMB[52][26] ), .Z(n83) );
  XOR2_X2 U206 ( .A(\CARRYB[52][21] ), .B(\SUMB[52][22] ), .Z(n84) );
  XOR2_X2 U207 ( .A(\CARRYB[52][22] ), .B(\SUMB[52][23] ), .Z(n85) );
  XOR2_X2 U208 ( .A(\CARRYB[52][24] ), .B(\SUMB[52][25] ), .Z(n86) );
  XOR2_X2 U209 ( .A(\CARRYB[52][20] ), .B(\SUMB[52][21] ), .Z(n87) );
  XOR2_X2 U210 ( .A(\CARRYB[52][29] ), .B(\SUMB[52][30] ), .Z(n88) );
  XOR2_X2 U211 ( .A(\CARRYB[52][30] ), .B(\SUMB[52][31] ), .Z(n89) );
  XOR2_X2 U212 ( .A(\CARRYB[52][32] ), .B(\SUMB[52][33] ), .Z(n90) );
  XOR2_X2 U213 ( .A(\CARRYB[52][33] ), .B(\SUMB[52][34] ), .Z(n91) );
  XOR2_X2 U214 ( .A(\CARRYB[52][34] ), .B(\SUMB[52][35] ), .Z(n92) );
  XOR2_X2 U215 ( .A(\CARRYB[52][36] ), .B(\SUMB[52][37] ), .Z(n93) );
  INV_X4 U216 ( .A(B[3]), .ZN(n441) );
  INV_X4 U217 ( .A(B[1]), .ZN(n445) );
  INV_X4 U218 ( .A(B[1]), .ZN(n443) );
  XOR2_X2 U219 ( .A(\CARRYB[52][51] ), .B(\ab[52][52] ), .Z(n94) );
  XOR2_X2 U220 ( .A(\CARRYB[52][50] ), .B(\SUMB[52][51] ), .Z(n95) );
  XOR2_X2 U221 ( .A(\CARRYB[52][48] ), .B(\SUMB[52][49] ), .Z(n96) );
  XOR2_X2 U222 ( .A(\CARRYB[52][43] ), .B(\SUMB[52][44] ), .Z(n97) );
  XOR2_X2 U223 ( .A(\CARRYB[52][41] ), .B(\SUMB[52][42] ), .Z(n98) );
  XOR2_X2 U224 ( .A(\CARRYB[52][46] ), .B(\SUMB[52][47] ), .Z(n99) );
  XOR2_X2 U225 ( .A(\CARRYB[52][45] ), .B(\SUMB[52][46] ), .Z(n100) );
  XOR2_X2 U226 ( .A(\CARRYB[52][42] ), .B(\SUMB[52][43] ), .Z(n101) );
  XOR2_X2 U227 ( .A(\CARRYB[52][44] ), .B(\SUMB[52][45] ), .Z(n102) );
  XOR2_X2 U228 ( .A(\CARRYB[52][47] ), .B(\SUMB[52][48] ), .Z(n103) );
  XOR2_X2 U229 ( .A(\CARRYB[52][49] ), .B(\SUMB[52][50] ), .Z(n104) );
  INV_X4 U230 ( .A(A[13]), .ZN(n304) );
  INV_X4 U231 ( .A(A[17]), .ZN(n298) );
  INV_X4 U232 ( .A(A[26]), .ZN(n280) );
  INV_X4 U233 ( .A(A[28]), .ZN(n275) );
  INV_X4 U234 ( .A(A[32]), .ZN(n267) );
  INV_X4 U235 ( .A(A[27]), .ZN(n278) );
  INV_X4 U236 ( .A(A[29]), .ZN(n272) );
  INV_X4 U237 ( .A(A[29]), .ZN(n273) );
  INV_X4 U238 ( .A(A[30]), .ZN(n271) );
  INV_X4 U239 ( .A(A[30]), .ZN(n270) );
  INV_X4 U240 ( .A(A[25]), .ZN(n283) );
  INV_X4 U241 ( .A(A[36]), .ZN(n258) );
  INV_X4 U242 ( .A(A[35]), .ZN(n260) );
  INV_X4 U243 ( .A(A[35]), .ZN(n259) );
  INV_X4 U244 ( .A(A[38]), .ZN(n252) );
  INV_X4 U245 ( .A(A[39]), .ZN(n247) );
  INV_X4 U246 ( .A(A[41]), .ZN(n242) );
  INV_X4 U247 ( .A(A[41]), .ZN(n241) );
  INV_X4 U248 ( .A(A[41]), .ZN(n240) );
  INV_X4 U249 ( .A(n235), .ZN(n234) );
  INV_X4 U250 ( .A(A[42]), .ZN(n239) );
  INV_X4 U251 ( .A(A[44]), .ZN(n231) );
  INV_X4 U252 ( .A(A[47]), .ZN(n221) );
  INV_X4 U253 ( .A(A[48]), .ZN(n218) );
  INV_X4 U254 ( .A(A[49]), .ZN(n215) );
  INV_X4 U255 ( .A(A[51]), .ZN(n212) );
  INV_X4 U256 ( .A(A[46]), .ZN(n225) );
  INV_X4 U257 ( .A(A[50]), .ZN(n213) );
  INV_X4 U258 ( .A(A[52]), .ZN(n448) );
  AND2_X4 U259 ( .A1(\ab[0][52] ), .A2(\ab[1][51] ), .ZN(n105) );
  AND2_X4 U260 ( .A1(\SUMB[52][2] ), .A2(\CARRYB[52][1] ), .ZN(n106) );
  AND2_X4 U261 ( .A1(\SUMB[52][1] ), .A2(\CARRYB[52][0] ), .ZN(n107) );
  AND2_X4 U262 ( .A1(\SUMB[52][3] ), .A2(\CARRYB[52][2] ), .ZN(n108) );
  AND2_X4 U263 ( .A1(\ab[0][51] ), .A2(\ab[1][50] ), .ZN(n109) );
  XOR2_X2 U264 ( .A(\ab[1][50] ), .B(\ab[0][51] ), .Z(n110) );
  XOR2_X2 U265 ( .A(\ab[1][49] ), .B(\ab[0][50] ), .Z(n111) );
  XOR2_X2 U266 ( .A(\ab[1][48] ), .B(\ab[0][49] ), .Z(n112) );
  XOR2_X2 U267 ( .A(\ab[1][47] ), .B(\ab[0][48] ), .Z(n113) );
  XOR2_X2 U268 ( .A(\ab[1][46] ), .B(\ab[0][47] ), .Z(n114) );
  XOR2_X2 U269 ( .A(\ab[1][45] ), .B(\ab[0][46] ), .Z(n115) );
  XOR2_X2 U270 ( .A(\ab[1][44] ), .B(\ab[0][45] ), .Z(n116) );
  XOR2_X2 U271 ( .A(\ab[1][43] ), .B(\ab[0][44] ), .Z(n117) );
  XOR2_X2 U272 ( .A(\ab[1][42] ), .B(\ab[0][43] ), .Z(n118) );
  XOR2_X2 U273 ( .A(\ab[1][41] ), .B(\ab[0][42] ), .Z(n119) );
  XOR2_X2 U274 ( .A(\ab[1][40] ), .B(\ab[0][41] ), .Z(n120) );
  XOR2_X2 U275 ( .A(\ab[1][39] ), .B(\ab[0][40] ), .Z(n121) );
  XOR2_X2 U276 ( .A(\ab[1][38] ), .B(\ab[0][39] ), .Z(n122) );
  XOR2_X2 U277 ( .A(\ab[1][37] ), .B(\ab[0][38] ), .Z(n123) );
  XOR2_X2 U278 ( .A(\ab[1][36] ), .B(\ab[0][37] ), .Z(n124) );
  XOR2_X2 U279 ( .A(\ab[1][35] ), .B(\ab[0][36] ), .Z(n125) );
  XOR2_X2 U280 ( .A(\ab[1][34] ), .B(\ab[0][35] ), .Z(n126) );
  XOR2_X2 U281 ( .A(\ab[1][33] ), .B(\ab[0][34] ), .Z(n127) );
  XOR2_X2 U282 ( .A(\ab[1][32] ), .B(\ab[0][33] ), .Z(n128) );
  XOR2_X2 U283 ( .A(\ab[1][31] ), .B(\ab[0][32] ), .Z(n129) );
  XOR2_X2 U284 ( .A(\ab[1][30] ), .B(\ab[0][31] ), .Z(n130) );
  XOR2_X2 U285 ( .A(\ab[1][29] ), .B(\ab[0][30] ), .Z(n131) );
  XOR2_X2 U286 ( .A(\ab[1][28] ), .B(\ab[0][29] ), .Z(n132) );
  XOR2_X2 U287 ( .A(\ab[1][27] ), .B(\ab[0][28] ), .Z(n133) );
  XOR2_X2 U288 ( .A(\ab[1][26] ), .B(\ab[0][27] ), .Z(n134) );
  XOR2_X2 U289 ( .A(\ab[1][25] ), .B(\ab[0][26] ), .Z(n135) );
  XOR2_X2 U290 ( .A(\ab[1][24] ), .B(\ab[0][25] ), .Z(n136) );
  XOR2_X2 U291 ( .A(\ab[1][23] ), .B(\ab[0][24] ), .Z(n137) );
  XOR2_X2 U292 ( .A(\ab[1][22] ), .B(\ab[0][23] ), .Z(n138) );
  XOR2_X2 U293 ( .A(\ab[1][21] ), .B(\ab[0][22] ), .Z(n139) );
  XOR2_X2 U294 ( .A(\ab[1][20] ), .B(\ab[0][21] ), .Z(n140) );
  XOR2_X2 U295 ( .A(\ab[1][19] ), .B(\ab[0][20] ), .Z(n141) );
  XOR2_X2 U296 ( .A(\ab[1][18] ), .B(\ab[0][19] ), .Z(n142) );
  XOR2_X2 U297 ( .A(\ab[1][17] ), .B(\ab[0][18] ), .Z(n143) );
  XOR2_X2 U298 ( .A(\ab[1][16] ), .B(\ab[0][17] ), .Z(n144) );
  XOR2_X2 U299 ( .A(\ab[1][15] ), .B(\ab[0][16] ), .Z(n145) );
  XOR2_X2 U300 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Z(n146) );
  XOR2_X2 U301 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Z(n147) );
  XOR2_X2 U302 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(n148) );
  XOR2_X2 U303 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(n149) );
  XOR2_X2 U304 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(n150) );
  XOR2_X2 U305 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(n151) );
  XOR2_X2 U306 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(n152) );
  XOR2_X2 U307 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(n153) );
  XOR2_X2 U308 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(n154) );
  XOR2_X2 U309 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(n155) );
  XOR2_X2 U310 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(n156) );
  XOR2_X2 U311 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(n157) );
  XOR2_X2 U312 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(n158) );
  INV_X4 U313 ( .A(B[50]), .ZN(n342) );
  AND2_X4 U314 ( .A1(\SUMB[52][5] ), .A2(\CARRYB[52][4] ), .ZN(n159) );
  AND2_X4 U315 ( .A1(\SUMB[52][7] ), .A2(\CARRYB[52][6] ), .ZN(n160) );
  AND2_X4 U316 ( .A1(\SUMB[52][10] ), .A2(\CARRYB[52][9] ), .ZN(n161) );
  AND2_X4 U317 ( .A1(\SUMB[52][12] ), .A2(\CARRYB[52][11] ), .ZN(n162) );
  AND2_X4 U318 ( .A1(\SUMB[52][4] ), .A2(\CARRYB[52][3] ), .ZN(n163) );
  AND2_X4 U319 ( .A1(\SUMB[52][6] ), .A2(\CARRYB[52][5] ), .ZN(n164) );
  AND2_X4 U320 ( .A1(\SUMB[52][8] ), .A2(\CARRYB[52][7] ), .ZN(n165) );
  AND2_X4 U321 ( .A1(\SUMB[52][9] ), .A2(\CARRYB[52][8] ), .ZN(n166) );
  AND2_X4 U322 ( .A1(\SUMB[52][11] ), .A2(\CARRYB[52][10] ), .ZN(n167) );
  AND2_X4 U323 ( .A1(\SUMB[52][15] ), .A2(\CARRYB[52][14] ), .ZN(n168) );
  AND2_X4 U324 ( .A1(\SUMB[52][13] ), .A2(\CARRYB[52][12] ), .ZN(n169) );
  AND2_X4 U325 ( .A1(\SUMB[52][14] ), .A2(\CARRYB[52][13] ), .ZN(n170) );
  INV_X4 U326 ( .A(B[14]), .ZN(n418) );
  INV_X4 U327 ( .A(B[14]), .ZN(n417) );
  INV_X4 U328 ( .A(B[13]), .ZN(n421) );
  INV_X4 U329 ( .A(B[13]), .ZN(n420) );
  INV_X4 U330 ( .A(B[12]), .ZN(n424) );
  INV_X4 U331 ( .A(B[12]), .ZN(n423) );
  INV_X4 U332 ( .A(B[16]), .ZN(n412) );
  INV_X4 U333 ( .A(B[16]), .ZN(n411) );
  INV_X4 U334 ( .A(B[15]), .ZN(n415) );
  INV_X4 U335 ( .A(B[15]), .ZN(n414) );
  INV_X4 U336 ( .A(B[19]), .ZN(n405) );
  INV_X4 U337 ( .A(B[49]), .ZN(n344) );
  INV_X4 U338 ( .A(B[43]), .ZN(n357) );
  INV_X4 U339 ( .A(A[2]), .ZN(n329) );
  INV_X4 U340 ( .A(A[2]), .ZN(n328) );
  INV_X4 U341 ( .A(A[5]), .ZN(n322) );
  INV_X4 U342 ( .A(A[5]), .ZN(n321) );
  INV_X4 U343 ( .A(A[5]), .ZN(n320) );
  INV_X4 U344 ( .A(A[1]), .ZN(n332) );
  INV_X4 U345 ( .A(A[1]), .ZN(n331) );
  INV_X4 U346 ( .A(A[4]), .ZN(n324) );
  INV_X4 U347 ( .A(A[4]), .ZN(n323) );
  INV_X4 U348 ( .A(A[3]), .ZN(n326) );
  INV_X4 U349 ( .A(A[3]), .ZN(n325) );
  INV_X4 U350 ( .A(A[0]), .ZN(n335) );
  INV_X4 U351 ( .A(A[0]), .ZN(n334) );
  INV_X4 U352 ( .A(A[0]), .ZN(n333) );
  XOR2_X2 U353 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(n171) );
  INV_X4 U354 ( .A(A[6]), .ZN(n318) );
  AND2_X4 U355 ( .A1(\SUMB[52][19] ), .A2(\CARRYB[52][18] ), .ZN(n172) );
  AND2_X4 U356 ( .A1(\SUMB[52][31] ), .A2(\CARRYB[52][30] ), .ZN(n173) );
  AND2_X4 U357 ( .A1(\SUMB[52][23] ), .A2(\CARRYB[52][22] ), .ZN(n174) );
  AND2_X4 U358 ( .A1(\SUMB[52][26] ), .A2(\CARRYB[52][25] ), .ZN(n175) );
  AND2_X4 U359 ( .A1(\SUMB[52][28] ), .A2(\CARRYB[52][27] ), .ZN(n176) );
  AND2_X4 U360 ( .A1(\SUMB[52][35] ), .A2(\CARRYB[52][34] ), .ZN(n177) );
  AND2_X4 U361 ( .A1(\SUMB[52][37] ), .A2(\CARRYB[52][36] ), .ZN(n178) );
  AND2_X4 U362 ( .A1(\SUMB[52][38] ), .A2(\CARRYB[52][37] ), .ZN(n179) );
  AND2_X4 U363 ( .A1(\SUMB[52][39] ), .A2(\CARRYB[52][38] ), .ZN(n180) );
  AND2_X4 U364 ( .A1(\SUMB[52][27] ), .A2(\CARRYB[52][26] ), .ZN(n181) );
  AND2_X4 U365 ( .A1(\SUMB[52][25] ), .A2(\CARRYB[52][24] ), .ZN(n182) );
  AND2_X4 U366 ( .A1(\SUMB[52][21] ), .A2(\CARRYB[52][20] ), .ZN(n183) );
  AND2_X4 U367 ( .A1(\SUMB[52][22] ), .A2(\CARRYB[52][21] ), .ZN(n184) );
  AND2_X4 U368 ( .A1(\SUMB[52][24] ), .A2(\CARRYB[52][23] ), .ZN(n185) );
  AND2_X4 U369 ( .A1(\SUMB[52][16] ), .A2(\CARRYB[52][15] ), .ZN(n186) );
  AND2_X4 U370 ( .A1(\SUMB[52][17] ), .A2(\CARRYB[52][16] ), .ZN(n187) );
  AND2_X4 U371 ( .A1(\SUMB[52][18] ), .A2(\CARRYB[52][17] ), .ZN(n188) );
  AND2_X4 U372 ( .A1(\SUMB[52][20] ), .A2(\CARRYB[52][19] ), .ZN(n189) );
  AND2_X4 U373 ( .A1(\SUMB[52][29] ), .A2(\CARRYB[52][28] ), .ZN(n190) );
  AND2_X4 U374 ( .A1(\SUMB[52][30] ), .A2(\CARRYB[52][29] ), .ZN(n191) );
  AND2_X4 U375 ( .A1(\SUMB[52][32] ), .A2(\CARRYB[52][31] ), .ZN(n192) );
  AND2_X4 U376 ( .A1(\SUMB[52][33] ), .A2(\CARRYB[52][32] ), .ZN(n193) );
  AND2_X4 U377 ( .A1(\SUMB[52][34] ), .A2(\CARRYB[52][33] ), .ZN(n194) );
  AND2_X4 U378 ( .A1(\SUMB[52][36] ), .A2(\CARRYB[52][35] ), .ZN(n195) );
  INV_X4 U379 ( .A(A[9]), .ZN(n310) );
  INV_X4 U380 ( .A(B[1]), .ZN(n444) );
  INV_X4 U381 ( .A(B[18]), .ZN(n407) );
  INV_X4 U382 ( .A(A[11]), .ZN(n308) );
  INV_X4 U383 ( .A(A[10]), .ZN(n309) );
  INV_X4 U384 ( .A(A[7]), .ZN(n314) );
  INV_X4 U385 ( .A(A[8]), .ZN(n313) );
  INV_X4 U386 ( .A(A[8]), .ZN(n312) );
  AND2_X4 U387 ( .A1(\SUMB[52][50] ), .A2(\CARRYB[52][49] ), .ZN(n196) );
  AND2_X4 U388 ( .A1(\SUMB[52][48] ), .A2(\CARRYB[52][47] ), .ZN(n197) );
  AND2_X4 U389 ( .A1(\SUMB[52][43] ), .A2(\CARRYB[52][42] ), .ZN(n198) );
  AND2_X4 U390 ( .A1(\SUMB[52][41] ), .A2(\CARRYB[52][40] ), .ZN(n199) );
  AND2_X4 U391 ( .A1(\SUMB[52][46] ), .A2(\CARRYB[52][45] ), .ZN(n200) );
  AND2_X4 U392 ( .A1(\SUMB[52][45] ), .A2(\CARRYB[52][44] ), .ZN(n201) );
  AND2_X4 U393 ( .A1(\SUMB[52][40] ), .A2(\CARRYB[52][39] ), .ZN(n202) );
  AND2_X4 U394 ( .A1(\SUMB[52][42] ), .A2(\CARRYB[52][41] ), .ZN(n203) );
  AND2_X4 U395 ( .A1(\SUMB[52][44] ), .A2(\CARRYB[52][43] ), .ZN(n204) );
  AND2_X4 U396 ( .A1(\SUMB[52][47] ), .A2(\CARRYB[52][46] ), .ZN(n205) );
  AND2_X4 U397 ( .A1(\SUMB[52][49] ), .A2(\CARRYB[52][48] ), .ZN(n206) );
  XOR2_X2 U398 ( .A(\CARRYB[52][0] ), .B(\SUMB[52][1] ), .Z(n207) );
  INV_X4 U399 ( .A(A[17]), .ZN(n297) );
  INV_X4 U400 ( .A(A[12]), .ZN(n306) );
  INV_X4 U401 ( .A(A[16]), .ZN(n299) );
  INV_X4 U402 ( .A(A[15]), .ZN(n301) );
  AND2_X4 U403 ( .A1(\ab[52][52] ), .A2(\CARRYB[52][51] ), .ZN(n208) );
  AND2_X4 U404 ( .A1(\SUMB[52][51] ), .A2(\CARRYB[52][50] ), .ZN(n209) );
  INV_X4 U405 ( .A(A[23]), .ZN(n287) );
  INV_X4 U406 ( .A(A[19]), .ZN(n294) );
  INV_X4 U407 ( .A(A[24]), .ZN(n285) );
  INV_X4 U408 ( .A(A[18]), .ZN(n295) );
  INV_X4 U409 ( .A(A[22]), .ZN(n289) );
  INV_X4 U410 ( .A(A[21]), .ZN(n291) );
  INV_X4 U411 ( .A(A[28]), .ZN(n276) );
  INV_X4 U412 ( .A(A[27]), .ZN(n279) );
  INV_X4 U413 ( .A(A[32]), .ZN(n266) );
  INV_X4 U414 ( .A(A[31]), .ZN(n268) );
  INV_X4 U415 ( .A(A[34]), .ZN(n263) );
  INV_X4 U416 ( .A(A[34]), .ZN(n262) );
  INV_X4 U417 ( .A(A[33]), .ZN(n265) );
  INV_X4 U418 ( .A(A[33]), .ZN(n264) );
  INV_X4 U419 ( .A(A[37]), .ZN(n253) );
  INV_X4 U420 ( .A(A[37]), .ZN(n255) );
  INV_X4 U421 ( .A(A[37]), .ZN(n254) );
  INV_X4 U422 ( .A(A[36]), .ZN(n257) );
  INV_X4 U423 ( .A(A[36]), .ZN(n256) );
  INV_X4 U424 ( .A(A[38]), .ZN(n251) );
  INV_X4 U425 ( .A(A[38]), .ZN(n249) );
  INV_X4 U426 ( .A(A[38]), .ZN(n250) );
  INV_X4 U427 ( .A(A[45]), .ZN(n228) );
  INV_X4 U428 ( .A(A[45]), .ZN(n227) );
  INV_X4 U429 ( .A(A[45]), .ZN(n226) );
  INV_X4 U430 ( .A(A[40]), .ZN(n246) );
  INV_X4 U431 ( .A(A[40]), .ZN(n245) );
  INV_X4 U432 ( .A(A[40]), .ZN(n244) );
  INV_X4 U433 ( .A(n235), .ZN(n233) );
  INV_X4 U434 ( .A(n235), .ZN(n232) );
  INV_X4 U435 ( .A(A[42]), .ZN(n238) );
  INV_X4 U436 ( .A(A[42]), .ZN(n237) );
  INV_X4 U437 ( .A(A[42]), .ZN(n236) );
  INV_X4 U438 ( .A(A[44]), .ZN(n230) );
  INV_X4 U439 ( .A(A[44]), .ZN(n229) );
  INV_X4 U440 ( .A(A[52]), .ZN(n447) );
  INV_X4 U441 ( .A(A[51]), .ZN(n211) );
  INV_X4 U442 ( .A(A[47]), .ZN(n223) );
  INV_X4 U443 ( .A(A[47]), .ZN(n222) );
  INV_X4 U444 ( .A(A[48]), .ZN(n220) );
  INV_X4 U445 ( .A(A[48]), .ZN(n219) );
  INV_X4 U446 ( .A(A[49]), .ZN(n217) );
  INV_X4 U447 ( .A(A[49]), .ZN(n216) );
  XOR2_X2 U448 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Z(PRODUCT[1]) );
  INV_X4 U449 ( .A(A[50]), .ZN(n450) );
  INV_X4 U450 ( .A(A[46]), .ZN(n451) );
  INV_X4 U451 ( .A(A[45]), .ZN(n452) );
  INV_X4 U452 ( .A(A[44]), .ZN(n453) );
  INV_X4 U453 ( .A(A[43]), .ZN(n454) );
  INV_X4 U454 ( .A(A[39]), .ZN(n455) );
  INV_X4 U455 ( .A(A[34]), .ZN(n456) );
  INV_X4 U456 ( .A(A[33]), .ZN(n457) );
  INV_X4 U457 ( .A(A[32]), .ZN(n458) );
  INV_X4 U458 ( .A(A[31]), .ZN(n459) );
  INV_X4 U459 ( .A(A[30]), .ZN(n460) );
  INV_X4 U460 ( .A(A[27]), .ZN(n461) );
  INV_X4 U461 ( .A(A[25]), .ZN(n462) );
  INV_X4 U462 ( .A(A[21]), .ZN(n463) );
  INV_X4 U463 ( .A(A[20]), .ZN(n464) );
  INV_X4 U464 ( .A(A[18]), .ZN(n465) );
  INV_X4 U465 ( .A(A[17]), .ZN(n466) );
  INV_X4 U466 ( .A(A[16]), .ZN(n467) );
  INV_X4 U467 ( .A(A[15]), .ZN(n468) );
  INV_X4 U468 ( .A(A[14]), .ZN(n469) );
  INV_X4 U469 ( .A(A[11]), .ZN(n470) );
  INV_X4 U470 ( .A(A[10]), .ZN(n471) );
  INV_X4 U471 ( .A(A[8]), .ZN(n472) );
  INV_X4 U472 ( .A(A[7]), .ZN(n473) );
  INV_X4 U473 ( .A(B[36]), .ZN(n474) );
  INV_X4 U474 ( .A(B[20]), .ZN(n475) );
  INV_X4 U475 ( .A(B[18]), .ZN(n476) );
  INV_X4 U476 ( .A(B[10]), .ZN(n477) );
  INV_X4 U477 ( .A(B[3]), .ZN(n478) );
  INV_X4 U478 ( .A(B[2]), .ZN(n479) );
  INV_X4 U479 ( .A(B[0]), .ZN(n480) );
  NOR2_X1 U481 ( .A1(n310), .A2(n429), .ZN(\ab[9][9] ) );
  NOR2_X1 U482 ( .A1(n310), .A2(n431), .ZN(\ab[9][8] ) );
  NOR2_X1 U483 ( .A1(n310), .A2(n433), .ZN(\ab[9][7] ) );
  NOR2_X1 U484 ( .A1(n310), .A2(n435), .ZN(\ab[9][6] ) );
  NOR2_X1 U485 ( .A1(n310), .A2(n437), .ZN(\ab[9][5] ) );
  NOR2_X1 U486 ( .A1(n310), .A2(n337), .ZN(\ab[9][52] ) );
  NOR2_X1 U487 ( .A1(n310), .A2(n340), .ZN(\ab[9][51] ) );
  NOR2_X1 U488 ( .A1(n310), .A2(n341), .ZN(\ab[9][50] ) );
  NOR2_X1 U489 ( .A1(n310), .A2(n439), .ZN(\ab[9][4] ) );
  NOR2_X1 U490 ( .A1(n311), .A2(n344), .ZN(\ab[9][49] ) );
  NOR2_X1 U491 ( .A1(n311), .A2(n345), .ZN(\ab[9][48] ) );
  NOR2_X1 U492 ( .A1(n311), .A2(n347), .ZN(\ab[9][47] ) );
  NOR2_X1 U493 ( .A1(n311), .A2(n349), .ZN(\ab[9][46] ) );
  NOR2_X1 U494 ( .A1(n311), .A2(n351), .ZN(\ab[9][45] ) );
  NOR2_X1 U495 ( .A1(n311), .A2(n355), .ZN(\ab[9][44] ) );
  NOR2_X1 U496 ( .A1(n311), .A2(n357), .ZN(\ab[9][43] ) );
  NOR2_X1 U497 ( .A1(n311), .A2(n360), .ZN(\ab[9][42] ) );
  NOR2_X1 U498 ( .A1(n311), .A2(n361), .ZN(\ab[9][41] ) );
  NOR2_X1 U499 ( .A1(n311), .A2(n363), .ZN(\ab[9][40] ) );
  NOR2_X1 U500 ( .A1(n311), .A2(n441), .ZN(\ab[9][3] ) );
  NOR2_X1 U501 ( .A1(n310), .A2(n365), .ZN(\ab[9][39] ) );
  NOR2_X1 U502 ( .A1(n311), .A2(n368), .ZN(\ab[9][38] ) );
  NOR2_X1 U503 ( .A1(n311), .A2(n371), .ZN(\ab[9][37] ) );
  NOR2_X1 U504 ( .A1(n311), .A2(n474), .ZN(\ab[9][36] ) );
  NOR2_X1 U505 ( .A1(n311), .A2(n373), .ZN(\ab[9][35] ) );
  NOR2_X1 U506 ( .A1(n311), .A2(n375), .ZN(\ab[9][34] ) );
  NOR2_X1 U507 ( .A1(n310), .A2(n377), .ZN(\ab[9][33] ) );
  NOR2_X1 U508 ( .A1(n311), .A2(n380), .ZN(\ab[9][32] ) );
  NOR2_X1 U509 ( .A1(n311), .A2(n381), .ZN(\ab[9][31] ) );
  NOR2_X1 U510 ( .A1(n310), .A2(n383), .ZN(\ab[9][30] ) );
  NOR2_X1 U511 ( .A1(n310), .A2(n479), .ZN(\ab[9][2] ) );
  NOR2_X1 U512 ( .A1(n310), .A2(n386), .ZN(\ab[9][29] ) );
  NOR2_X1 U513 ( .A1(n310), .A2(n388), .ZN(\ab[9][28] ) );
  NOR2_X1 U514 ( .A1(n310), .A2(n390), .ZN(\ab[9][27] ) );
  NOR2_X1 U515 ( .A1(n310), .A2(n392), .ZN(\ab[9][26] ) );
  NOR2_X1 U516 ( .A1(n310), .A2(n394), .ZN(\ab[9][25] ) );
  NOR2_X1 U517 ( .A1(n310), .A2(n396), .ZN(\ab[9][24] ) );
  NOR2_X1 U518 ( .A1(n310), .A2(n398), .ZN(\ab[9][23] ) );
  NOR2_X1 U519 ( .A1(n310), .A2(n400), .ZN(\ab[9][22] ) );
  NOR2_X1 U520 ( .A1(n310), .A2(n402), .ZN(\ab[9][21] ) );
  NOR2_X1 U521 ( .A1(n310), .A2(n475), .ZN(\ab[9][20] ) );
  NOR2_X1 U522 ( .A1(n310), .A2(n444), .ZN(\ab[9][1] ) );
  NOR2_X1 U523 ( .A1(n310), .A2(n405), .ZN(\ab[9][19] ) );
  NOR2_X1 U524 ( .A1(n310), .A2(n407), .ZN(\ab[9][18] ) );
  NOR2_X1 U525 ( .A1(n310), .A2(n409), .ZN(\ab[9][17] ) );
  NOR2_X1 U526 ( .A1(n310), .A2(n412), .ZN(\ab[9][16] ) );
  NOR2_X1 U527 ( .A1(n310), .A2(n415), .ZN(\ab[9][15] ) );
  NOR2_X1 U528 ( .A1(n310), .A2(n418), .ZN(\ab[9][14] ) );
  NOR2_X1 U529 ( .A1(n310), .A2(n421), .ZN(\ab[9][13] ) );
  NOR2_X1 U530 ( .A1(n310), .A2(n424), .ZN(\ab[9][12] ) );
  NOR2_X1 U531 ( .A1(n310), .A2(n426), .ZN(\ab[9][11] ) );
  NOR2_X1 U532 ( .A1(n310), .A2(n477), .ZN(\ab[9][10] ) );
  NOR2_X1 U533 ( .A1(n310), .A2(n446), .ZN(\ab[9][0] ) );
  NOR2_X1 U534 ( .A1(n429), .A2(n312), .ZN(\ab[8][9] ) );
  NOR2_X1 U535 ( .A1(n431), .A2(n312), .ZN(\ab[8][8] ) );
  NOR2_X1 U536 ( .A1(n433), .A2(n312), .ZN(\ab[8][7] ) );
  NOR2_X1 U537 ( .A1(n435), .A2(n312), .ZN(\ab[8][6] ) );
  NOR2_X1 U538 ( .A1(n437), .A2(n312), .ZN(\ab[8][5] ) );
  NOR2_X1 U539 ( .A1(n337), .A2(n312), .ZN(\ab[8][52] ) );
  NOR2_X1 U540 ( .A1(n340), .A2(n312), .ZN(\ab[8][51] ) );
  NOR2_X1 U541 ( .A1(n341), .A2(n313), .ZN(\ab[8][50] ) );
  NOR2_X1 U542 ( .A1(n439), .A2(n312), .ZN(\ab[8][4] ) );
  NOR2_X1 U543 ( .A1(n344), .A2(n312), .ZN(\ab[8][49] ) );
  NOR2_X1 U544 ( .A1(n346), .A2(n472), .ZN(\ab[8][48] ) );
  NOR2_X1 U545 ( .A1(n348), .A2(n472), .ZN(\ab[8][47] ) );
  NOR2_X1 U546 ( .A1(n350), .A2(n472), .ZN(\ab[8][46] ) );
  NOR2_X1 U547 ( .A1(n352), .A2(n472), .ZN(\ab[8][45] ) );
  NOR2_X1 U548 ( .A1(n355), .A2(n472), .ZN(\ab[8][44] ) );
  NOR2_X1 U549 ( .A1(n357), .A2(n472), .ZN(\ab[8][43] ) );
  NOR2_X1 U550 ( .A1(n360), .A2(n472), .ZN(\ab[8][42] ) );
  NOR2_X1 U551 ( .A1(n362), .A2(n313), .ZN(\ab[8][41] ) );
  NOR2_X1 U552 ( .A1(n364), .A2(n472), .ZN(\ab[8][40] ) );
  NOR2_X1 U553 ( .A1(n441), .A2(n312), .ZN(\ab[8][3] ) );
  NOR2_X1 U554 ( .A1(n366), .A2(n313), .ZN(\ab[8][39] ) );
  NOR2_X1 U555 ( .A1(n368), .A2(n313), .ZN(\ab[8][38] ) );
  NOR2_X1 U556 ( .A1(n371), .A2(n312), .ZN(\ab[8][37] ) );
  NOR2_X1 U557 ( .A1(n372), .A2(n312), .ZN(\ab[8][36] ) );
  NOR2_X1 U558 ( .A1(n374), .A2(n312), .ZN(\ab[8][35] ) );
  NOR2_X1 U559 ( .A1(n376), .A2(n312), .ZN(\ab[8][34] ) );
  NOR2_X1 U560 ( .A1(n378), .A2(n312), .ZN(\ab[8][33] ) );
  NOR2_X1 U561 ( .A1(n379), .A2(n313), .ZN(\ab[8][32] ) );
  NOR2_X1 U562 ( .A1(n382), .A2(n312), .ZN(\ab[8][31] ) );
  NOR2_X1 U563 ( .A1(n384), .A2(n313), .ZN(\ab[8][30] ) );
  NOR2_X1 U564 ( .A1(n479), .A2(n312), .ZN(\ab[8][2] ) );
  NOR2_X1 U565 ( .A1(n385), .A2(n313), .ZN(\ab[8][29] ) );
  NOR2_X1 U566 ( .A1(n388), .A2(n313), .ZN(\ab[8][28] ) );
  NOR2_X1 U567 ( .A1(n389), .A2(n313), .ZN(\ab[8][27] ) );
  NOR2_X1 U568 ( .A1(n391), .A2(n313), .ZN(\ab[8][26] ) );
  NOR2_X1 U569 ( .A1(n393), .A2(n313), .ZN(\ab[8][25] ) );
  NOR2_X1 U570 ( .A1(n395), .A2(n313), .ZN(\ab[8][24] ) );
  NOR2_X1 U571 ( .A1(n397), .A2(n313), .ZN(\ab[8][23] ) );
  NOR2_X1 U572 ( .A1(n399), .A2(n313), .ZN(\ab[8][22] ) );
  NOR2_X1 U573 ( .A1(n401), .A2(n313), .ZN(\ab[8][21] ) );
  NOR2_X1 U574 ( .A1(n475), .A2(n313), .ZN(\ab[8][20] ) );
  NOR2_X1 U575 ( .A1(n444), .A2(n313), .ZN(\ab[8][1] ) );
  NOR2_X1 U576 ( .A1(n405), .A2(n312), .ZN(\ab[8][19] ) );
  NOR2_X1 U577 ( .A1(n407), .A2(n312), .ZN(\ab[8][18] ) );
  NOR2_X1 U578 ( .A1(n408), .A2(n312), .ZN(\ab[8][17] ) );
  NOR2_X1 U579 ( .A1(n412), .A2(n312), .ZN(\ab[8][16] ) );
  NOR2_X1 U580 ( .A1(n415), .A2(n312), .ZN(\ab[8][15] ) );
  NOR2_X1 U581 ( .A1(n418), .A2(n312), .ZN(\ab[8][14] ) );
  NOR2_X1 U582 ( .A1(n421), .A2(n312), .ZN(\ab[8][13] ) );
  NOR2_X1 U583 ( .A1(n424), .A2(n312), .ZN(\ab[8][12] ) );
  NOR2_X1 U584 ( .A1(n425), .A2(n312), .ZN(\ab[8][11] ) );
  NOR2_X1 U585 ( .A1(n427), .A2(n312), .ZN(\ab[8][10] ) );
  NOR2_X1 U586 ( .A1(n480), .A2(n312), .ZN(\ab[8][0] ) );
  NOR2_X1 U587 ( .A1(n429), .A2(n314), .ZN(\ab[7][9] ) );
  NOR2_X1 U588 ( .A1(n431), .A2(n314), .ZN(\ab[7][8] ) );
  NOR2_X1 U589 ( .A1(n433), .A2(n314), .ZN(\ab[7][7] ) );
  NOR2_X1 U590 ( .A1(n435), .A2(n314), .ZN(\ab[7][6] ) );
  NOR2_X1 U591 ( .A1(n437), .A2(n314), .ZN(\ab[7][5] ) );
  NOR2_X1 U592 ( .A1(n337), .A2(n314), .ZN(\ab[7][52] ) );
  NOR2_X1 U593 ( .A1(n340), .A2(n314), .ZN(\ab[7][51] ) );
  NOR2_X1 U594 ( .A1(n341), .A2(n314), .ZN(\ab[7][50] ) );
  NOR2_X1 U595 ( .A1(n439), .A2(n314), .ZN(\ab[7][4] ) );
  NOR2_X1 U596 ( .A1(n344), .A2(n315), .ZN(\ab[7][49] ) );
  NOR2_X1 U597 ( .A1(n346), .A2(n473), .ZN(\ab[7][48] ) );
  NOR2_X1 U598 ( .A1(n348), .A2(n473), .ZN(\ab[7][47] ) );
  NOR2_X1 U599 ( .A1(n350), .A2(n473), .ZN(\ab[7][46] ) );
  NOR2_X1 U600 ( .A1(n352), .A2(n473), .ZN(\ab[7][45] ) );
  NOR2_X1 U601 ( .A1(n355), .A2(n473), .ZN(\ab[7][44] ) );
  NOR2_X1 U602 ( .A1(n357), .A2(n315), .ZN(\ab[7][43] ) );
  NOR2_X1 U603 ( .A1(n360), .A2(n315), .ZN(\ab[7][42] ) );
  NOR2_X1 U604 ( .A1(n362), .A2(n473), .ZN(\ab[7][41] ) );
  NOR2_X1 U605 ( .A1(n364), .A2(n473), .ZN(\ab[7][40] ) );
  NOR2_X1 U606 ( .A1(n441), .A2(n314), .ZN(\ab[7][3] ) );
  NOR2_X1 U607 ( .A1(n366), .A2(n315), .ZN(\ab[7][39] ) );
  NOR2_X1 U608 ( .A1(n368), .A2(n315), .ZN(\ab[7][38] ) );
  NOR2_X1 U609 ( .A1(n371), .A2(n315), .ZN(\ab[7][37] ) );
  NOR2_X1 U610 ( .A1(n474), .A2(n315), .ZN(\ab[7][36] ) );
  NOR2_X1 U611 ( .A1(n374), .A2(n315), .ZN(\ab[7][35] ) );
  NOR2_X1 U612 ( .A1(n376), .A2(n315), .ZN(\ab[7][34] ) );
  NOR2_X1 U613 ( .A1(n378), .A2(n315), .ZN(\ab[7][33] ) );
  NOR2_X1 U614 ( .A1(n380), .A2(n315), .ZN(\ab[7][32] ) );
  NOR2_X1 U615 ( .A1(n382), .A2(n315), .ZN(\ab[7][31] ) );
  NOR2_X1 U616 ( .A1(n384), .A2(n315), .ZN(\ab[7][30] ) );
  NOR2_X1 U617 ( .A1(n479), .A2(n315), .ZN(\ab[7][2] ) );
  NOR2_X1 U618 ( .A1(n386), .A2(n314), .ZN(\ab[7][29] ) );
  NOR2_X1 U619 ( .A1(n388), .A2(n314), .ZN(\ab[7][28] ) );
  NOR2_X1 U620 ( .A1(n390), .A2(n314), .ZN(\ab[7][27] ) );
  NOR2_X1 U621 ( .A1(n392), .A2(n314), .ZN(\ab[7][26] ) );
  NOR2_X1 U622 ( .A1(n394), .A2(n314), .ZN(\ab[7][25] ) );
  NOR2_X1 U623 ( .A1(n396), .A2(n314), .ZN(\ab[7][24] ) );
  NOR2_X1 U624 ( .A1(n398), .A2(n314), .ZN(\ab[7][23] ) );
  NOR2_X1 U625 ( .A1(n400), .A2(n314), .ZN(\ab[7][22] ) );
  NOR2_X1 U626 ( .A1(n402), .A2(n315), .ZN(\ab[7][21] ) );
  NOR2_X1 U627 ( .A1(n403), .A2(n315), .ZN(\ab[7][20] ) );
  NOR2_X1 U628 ( .A1(n444), .A2(n315), .ZN(\ab[7][1] ) );
  NOR2_X1 U629 ( .A1(n405), .A2(n314), .ZN(\ab[7][19] ) );
  NOR2_X1 U630 ( .A1(n407), .A2(n314), .ZN(\ab[7][18] ) );
  NOR2_X1 U631 ( .A1(n409), .A2(n314), .ZN(\ab[7][17] ) );
  NOR2_X1 U632 ( .A1(n412), .A2(n314), .ZN(\ab[7][16] ) );
  NOR2_X1 U633 ( .A1(n415), .A2(n314), .ZN(\ab[7][15] ) );
  NOR2_X1 U634 ( .A1(n418), .A2(n314), .ZN(\ab[7][14] ) );
  NOR2_X1 U635 ( .A1(n421), .A2(n314), .ZN(\ab[7][13] ) );
  NOR2_X1 U636 ( .A1(n424), .A2(n314), .ZN(\ab[7][12] ) );
  NOR2_X1 U637 ( .A1(n426), .A2(n314), .ZN(\ab[7][11] ) );
  NOR2_X1 U638 ( .A1(n477), .A2(n314), .ZN(\ab[7][10] ) );
  NOR2_X1 U639 ( .A1(n480), .A2(n314), .ZN(\ab[7][0] ) );
  NOR2_X1 U640 ( .A1(n429), .A2(n316), .ZN(\ab[6][9] ) );
  NOR2_X1 U641 ( .A1(n431), .A2(n316), .ZN(\ab[6][8] ) );
  NOR2_X1 U642 ( .A1(n433), .A2(n316), .ZN(\ab[6][7] ) );
  NOR2_X1 U643 ( .A1(n435), .A2(n316), .ZN(\ab[6][6] ) );
  NOR2_X1 U644 ( .A1(n437), .A2(n316), .ZN(\ab[6][5] ) );
  NOR2_X1 U645 ( .A1(n337), .A2(n316), .ZN(\ab[6][52] ) );
  NOR2_X1 U646 ( .A1(n340), .A2(n316), .ZN(\ab[6][51] ) );
  NOR2_X1 U647 ( .A1(n341), .A2(n317), .ZN(\ab[6][50] ) );
  NOR2_X1 U648 ( .A1(n439), .A2(n316), .ZN(\ab[6][4] ) );
  NOR2_X1 U649 ( .A1(n344), .A2(n318), .ZN(\ab[6][49] ) );
  NOR2_X1 U650 ( .A1(n346), .A2(n318), .ZN(\ab[6][48] ) );
  NOR2_X1 U651 ( .A1(n348), .A2(n318), .ZN(\ab[6][47] ) );
  NOR2_X1 U652 ( .A1(n350), .A2(n318), .ZN(\ab[6][46] ) );
  NOR2_X1 U653 ( .A1(n352), .A2(n317), .ZN(\ab[6][45] ) );
  NOR2_X1 U654 ( .A1(n355), .A2(n318), .ZN(\ab[6][44] ) );
  NOR2_X1 U655 ( .A1(n357), .A2(n318), .ZN(\ab[6][43] ) );
  NOR2_X1 U656 ( .A1(n360), .A2(n318), .ZN(\ab[6][42] ) );
  NOR2_X1 U657 ( .A1(n362), .A2(n316), .ZN(\ab[6][41] ) );
  NOR2_X1 U658 ( .A1(n364), .A2(n316), .ZN(\ab[6][40] ) );
  NOR2_X1 U659 ( .A1(n441), .A2(n316), .ZN(\ab[6][3] ) );
  NOR2_X1 U660 ( .A1(n366), .A2(n317), .ZN(\ab[6][39] ) );
  NOR2_X1 U661 ( .A1(n368), .A2(n317), .ZN(\ab[6][38] ) );
  NOR2_X1 U662 ( .A1(n371), .A2(n317), .ZN(\ab[6][37] ) );
  NOR2_X1 U663 ( .A1(n474), .A2(n317), .ZN(\ab[6][36] ) );
  NOR2_X1 U664 ( .A1(n374), .A2(n317), .ZN(\ab[6][35] ) );
  NOR2_X1 U665 ( .A1(n376), .A2(n317), .ZN(\ab[6][34] ) );
  NOR2_X1 U666 ( .A1(n378), .A2(n317), .ZN(\ab[6][33] ) );
  NOR2_X1 U667 ( .A1(n380), .A2(n317), .ZN(\ab[6][32] ) );
  NOR2_X1 U668 ( .A1(n382), .A2(n317), .ZN(\ab[6][31] ) );
  NOR2_X1 U669 ( .A1(n384), .A2(n317), .ZN(\ab[6][30] ) );
  NOR2_X1 U670 ( .A1(n479), .A2(n317), .ZN(\ab[6][2] ) );
  NOR2_X1 U671 ( .A1(n385), .A2(n316), .ZN(\ab[6][29] ) );
  NOR2_X1 U672 ( .A1(n388), .A2(n316), .ZN(\ab[6][28] ) );
  NOR2_X1 U673 ( .A1(n389), .A2(n316), .ZN(\ab[6][27] ) );
  NOR2_X1 U674 ( .A1(n391), .A2(n316), .ZN(\ab[6][26] ) );
  NOR2_X1 U675 ( .A1(n393), .A2(n316), .ZN(\ab[6][25] ) );
  NOR2_X1 U676 ( .A1(n395), .A2(n316), .ZN(\ab[6][24] ) );
  NOR2_X1 U677 ( .A1(n397), .A2(n316), .ZN(\ab[6][23] ) );
  NOR2_X1 U678 ( .A1(n399), .A2(n316), .ZN(\ab[6][22] ) );
  NOR2_X1 U679 ( .A1(n401), .A2(n316), .ZN(\ab[6][21] ) );
  NOR2_X1 U680 ( .A1(n475), .A2(n316), .ZN(\ab[6][20] ) );
  NOR2_X1 U681 ( .A1(n444), .A2(n316), .ZN(\ab[6][1] ) );
  NOR2_X1 U682 ( .A1(n405), .A2(n316), .ZN(\ab[6][19] ) );
  NOR2_X1 U683 ( .A1(n407), .A2(n316), .ZN(\ab[6][18] ) );
  NOR2_X1 U684 ( .A1(n408), .A2(n316), .ZN(\ab[6][17] ) );
  NOR2_X1 U685 ( .A1(n412), .A2(n316), .ZN(\ab[6][16] ) );
  NOR2_X1 U686 ( .A1(n415), .A2(n316), .ZN(\ab[6][15] ) );
  NOR2_X1 U687 ( .A1(n418), .A2(n316), .ZN(\ab[6][14] ) );
  NOR2_X1 U688 ( .A1(n421), .A2(n316), .ZN(\ab[6][13] ) );
  NOR2_X1 U689 ( .A1(n424), .A2(n316), .ZN(\ab[6][12] ) );
  NOR2_X1 U690 ( .A1(n425), .A2(n316), .ZN(\ab[6][11] ) );
  NOR2_X1 U691 ( .A1(n477), .A2(n316), .ZN(\ab[6][10] ) );
  NOR2_X1 U692 ( .A1(n480), .A2(n316), .ZN(\ab[6][0] ) );
  NOR2_X1 U693 ( .A1(n429), .A2(n319), .ZN(\ab[5][9] ) );
  NOR2_X1 U694 ( .A1(n431), .A2(n319), .ZN(\ab[5][8] ) );
  NOR2_X1 U695 ( .A1(n433), .A2(n319), .ZN(\ab[5][7] ) );
  NOR2_X1 U696 ( .A1(n435), .A2(n319), .ZN(\ab[5][6] ) );
  NOR2_X1 U697 ( .A1(n437), .A2(n319), .ZN(\ab[5][5] ) );
  NOR2_X1 U698 ( .A1(n337), .A2(n320), .ZN(\ab[5][52] ) );
  NOR2_X1 U699 ( .A1(n340), .A2(n321), .ZN(\ab[5][51] ) );
  NOR2_X1 U700 ( .A1(n341), .A2(n322), .ZN(\ab[5][50] ) );
  NOR2_X1 U701 ( .A1(n439), .A2(n319), .ZN(\ab[5][4] ) );
  NOR2_X1 U702 ( .A1(n344), .A2(n322), .ZN(\ab[5][49] ) );
  NOR2_X1 U703 ( .A1(n346), .A2(n322), .ZN(\ab[5][48] ) );
  NOR2_X1 U704 ( .A1(n348), .A2(n319), .ZN(\ab[5][47] ) );
  NOR2_X1 U705 ( .A1(n350), .A2(n319), .ZN(\ab[5][46] ) );
  NOR2_X1 U706 ( .A1(n352), .A2(n320), .ZN(\ab[5][45] ) );
  NOR2_X1 U707 ( .A1(n355), .A2(n321), .ZN(\ab[5][44] ) );
  NOR2_X1 U708 ( .A1(n357), .A2(n320), .ZN(\ab[5][43] ) );
  NOR2_X1 U709 ( .A1(n360), .A2(n321), .ZN(\ab[5][42] ) );
  NOR2_X1 U710 ( .A1(n362), .A2(n320), .ZN(\ab[5][41] ) );
  NOR2_X1 U711 ( .A1(n364), .A2(n319), .ZN(\ab[5][40] ) );
  NOR2_X1 U712 ( .A1(n441), .A2(n319), .ZN(\ab[5][3] ) );
  NOR2_X1 U713 ( .A1(n366), .A2(n321), .ZN(\ab[5][39] ) );
  NOR2_X1 U714 ( .A1(n368), .A2(n321), .ZN(\ab[5][38] ) );
  NOR2_X1 U715 ( .A1(n371), .A2(n321), .ZN(\ab[5][37] ) );
  NOR2_X1 U716 ( .A1(n474), .A2(n321), .ZN(\ab[5][36] ) );
  NOR2_X1 U717 ( .A1(n374), .A2(n321), .ZN(\ab[5][35] ) );
  NOR2_X1 U718 ( .A1(n376), .A2(n321), .ZN(\ab[5][34] ) );
  NOR2_X1 U719 ( .A1(n378), .A2(n321), .ZN(\ab[5][33] ) );
  NOR2_X1 U720 ( .A1(n380), .A2(n321), .ZN(\ab[5][32] ) );
  NOR2_X1 U721 ( .A1(n382), .A2(n321), .ZN(\ab[5][31] ) );
  NOR2_X1 U722 ( .A1(n384), .A2(n321), .ZN(\ab[5][30] ) );
  NOR2_X1 U723 ( .A1(n479), .A2(n321), .ZN(\ab[5][2] ) );
  NOR2_X1 U724 ( .A1(n386), .A2(n320), .ZN(\ab[5][29] ) );
  NOR2_X1 U725 ( .A1(n388), .A2(n320), .ZN(\ab[5][28] ) );
  NOR2_X1 U726 ( .A1(n390), .A2(n320), .ZN(\ab[5][27] ) );
  NOR2_X1 U727 ( .A1(n392), .A2(n320), .ZN(\ab[5][26] ) );
  NOR2_X1 U728 ( .A1(n394), .A2(n320), .ZN(\ab[5][25] ) );
  NOR2_X1 U729 ( .A1(n396), .A2(n320), .ZN(\ab[5][24] ) );
  NOR2_X1 U730 ( .A1(n398), .A2(n320), .ZN(\ab[5][23] ) );
  NOR2_X1 U731 ( .A1(n400), .A2(n320), .ZN(\ab[5][22] ) );
  NOR2_X1 U732 ( .A1(n402), .A2(n320), .ZN(\ab[5][21] ) );
  NOR2_X1 U733 ( .A1(n475), .A2(n320), .ZN(\ab[5][20] ) );
  NOR2_X1 U734 ( .A1(n444), .A2(n320), .ZN(\ab[5][1] ) );
  NOR2_X1 U735 ( .A1(n405), .A2(n319), .ZN(\ab[5][19] ) );
  NOR2_X1 U736 ( .A1(n407), .A2(n319), .ZN(\ab[5][18] ) );
  NOR2_X1 U737 ( .A1(n409), .A2(n319), .ZN(\ab[5][17] ) );
  NOR2_X1 U738 ( .A1(n412), .A2(n319), .ZN(\ab[5][16] ) );
  NOR2_X1 U739 ( .A1(n415), .A2(n319), .ZN(\ab[5][15] ) );
  NOR2_X1 U740 ( .A1(n418), .A2(n319), .ZN(\ab[5][14] ) );
  NOR2_X1 U741 ( .A1(n421), .A2(n319), .ZN(\ab[5][13] ) );
  NOR2_X1 U742 ( .A1(n424), .A2(n319), .ZN(\ab[5][12] ) );
  NOR2_X1 U743 ( .A1(n426), .A2(n319), .ZN(\ab[5][11] ) );
  NOR2_X1 U744 ( .A1(n477), .A2(n319), .ZN(\ab[5][10] ) );
  NOR2_X1 U745 ( .A1(n480), .A2(n319), .ZN(\ab[5][0] ) );
  NOR2_X1 U746 ( .A1(n429), .A2(n447), .ZN(\ab[52][9] ) );
  NOR2_X1 U747 ( .A1(n431), .A2(n447), .ZN(\ab[52][8] ) );
  NOR2_X1 U748 ( .A1(n433), .A2(n447), .ZN(\ab[52][7] ) );
  NOR2_X1 U749 ( .A1(n435), .A2(n447), .ZN(\ab[52][6] ) );
  NOR2_X1 U750 ( .A1(n437), .A2(n447), .ZN(\ab[52][5] ) );
  NOR2_X1 U751 ( .A1(n337), .A2(n447), .ZN(\ab[52][52] ) );
  NOR2_X1 U752 ( .A1(n340), .A2(n447), .ZN(\ab[52][51] ) );
  NOR2_X1 U753 ( .A1(n341), .A2(n447), .ZN(\ab[52][50] ) );
  NOR2_X1 U754 ( .A1(n439), .A2(n447), .ZN(\ab[52][4] ) );
  NOR2_X1 U755 ( .A1(n344), .A2(n447), .ZN(\ab[52][49] ) );
  NOR2_X1 U756 ( .A1(n346), .A2(n447), .ZN(\ab[52][48] ) );
  NOR2_X1 U757 ( .A1(n348), .A2(n448), .ZN(\ab[52][47] ) );
  NOR2_X1 U758 ( .A1(n350), .A2(n448), .ZN(\ab[52][46] ) );
  NOR2_X1 U759 ( .A1(n352), .A2(n448), .ZN(\ab[52][45] ) );
  NOR2_X1 U760 ( .A1(n355), .A2(n448), .ZN(\ab[52][44] ) );
  NOR2_X1 U761 ( .A1(n357), .A2(n448), .ZN(\ab[52][43] ) );
  NOR2_X1 U762 ( .A1(n360), .A2(n448), .ZN(\ab[52][42] ) );
  NOR2_X1 U763 ( .A1(n362), .A2(n448), .ZN(\ab[52][41] ) );
  NOR2_X1 U764 ( .A1(n364), .A2(n448), .ZN(\ab[52][40] ) );
  NOR2_X1 U765 ( .A1(n441), .A2(n447), .ZN(\ab[52][3] ) );
  NOR2_X1 U766 ( .A1(n366), .A2(n448), .ZN(\ab[52][39] ) );
  NOR2_X1 U767 ( .A1(n368), .A2(n448), .ZN(\ab[52][38] ) );
  NOR2_X1 U768 ( .A1(n371), .A2(n447), .ZN(\ab[52][37] ) );
  NOR2_X1 U769 ( .A1(n372), .A2(n449), .ZN(\ab[52][36] ) );
  NOR2_X1 U770 ( .A1(n374), .A2(n449), .ZN(\ab[52][35] ) );
  NOR2_X1 U771 ( .A1(n376), .A2(n449), .ZN(\ab[52][34] ) );
  NOR2_X1 U772 ( .A1(n378), .A2(n449), .ZN(\ab[52][33] ) );
  NOR2_X1 U773 ( .A1(n379), .A2(n449), .ZN(\ab[52][32] ) );
  NOR2_X1 U774 ( .A1(n382), .A2(n448), .ZN(\ab[52][31] ) );
  NOR2_X1 U775 ( .A1(n384), .A2(n449), .ZN(\ab[52][30] ) );
  NOR2_X1 U776 ( .A1(n479), .A2(n449), .ZN(\ab[52][2] ) );
  NOR2_X1 U777 ( .A1(n385), .A2(n449), .ZN(\ab[52][29] ) );
  NOR2_X1 U778 ( .A1(n388), .A2(n449), .ZN(\ab[52][28] ) );
  NOR2_X1 U779 ( .A1(n389), .A2(n448), .ZN(\ab[52][27] ) );
  NOR2_X1 U780 ( .A1(n391), .A2(n448), .ZN(\ab[52][26] ) );
  NOR2_X1 U781 ( .A1(n393), .A2(n448), .ZN(\ab[52][25] ) );
  NOR2_X1 U782 ( .A1(n395), .A2(n448), .ZN(\ab[52][24] ) );
  NOR2_X1 U783 ( .A1(n397), .A2(n448), .ZN(\ab[52][23] ) );
  NOR2_X1 U784 ( .A1(n399), .A2(n448), .ZN(\ab[52][22] ) );
  NOR2_X1 U785 ( .A1(n401), .A2(n448), .ZN(\ab[52][21] ) );
  NOR2_X1 U786 ( .A1(n403), .A2(n448), .ZN(\ab[52][20] ) );
  NOR2_X1 U787 ( .A1(n444), .A2(n448), .ZN(\ab[52][1] ) );
  NOR2_X1 U788 ( .A1(n405), .A2(n448), .ZN(\ab[52][19] ) );
  NOR2_X1 U789 ( .A1(n407), .A2(n448), .ZN(\ab[52][18] ) );
  NOR2_X1 U790 ( .A1(n408), .A2(n447), .ZN(\ab[52][17] ) );
  NOR2_X1 U791 ( .A1(n412), .A2(n447), .ZN(\ab[52][16] ) );
  NOR2_X1 U792 ( .A1(n415), .A2(n447), .ZN(\ab[52][15] ) );
  NOR2_X1 U793 ( .A1(n418), .A2(n447), .ZN(\ab[52][14] ) );
  NOR2_X1 U794 ( .A1(n421), .A2(n447), .ZN(\ab[52][13] ) );
  NOR2_X1 U795 ( .A1(n424), .A2(n447), .ZN(\ab[52][12] ) );
  NOR2_X1 U796 ( .A1(n425), .A2(n447), .ZN(\ab[52][11] ) );
  NOR2_X1 U797 ( .A1(n477), .A2(n447), .ZN(\ab[52][10] ) );
  NOR2_X1 U798 ( .A1(n480), .A2(n447), .ZN(\ab[52][0] ) );
  NOR2_X1 U799 ( .A1(n429), .A2(n211), .ZN(\ab[51][9] ) );
  NOR2_X1 U800 ( .A1(n431), .A2(n211), .ZN(\ab[51][8] ) );
  NOR2_X1 U801 ( .A1(n433), .A2(n211), .ZN(\ab[51][7] ) );
  NOR2_X1 U802 ( .A1(n435), .A2(n211), .ZN(\ab[51][6] ) );
  NOR2_X1 U803 ( .A1(n437), .A2(n211), .ZN(\ab[51][5] ) );
  NOR2_X1 U804 ( .A1(n337), .A2(n211), .ZN(\ab[51][52] ) );
  NOR2_X1 U805 ( .A1(n340), .A2(n211), .ZN(\ab[51][51] ) );
  NOR2_X1 U806 ( .A1(n341), .A2(n211), .ZN(\ab[51][50] ) );
  NOR2_X1 U807 ( .A1(n439), .A2(n212), .ZN(\ab[51][4] ) );
  NOR2_X1 U808 ( .A1(n344), .A2(n212), .ZN(\ab[51][49] ) );
  NOR2_X1 U809 ( .A1(n345), .A2(n211), .ZN(\ab[51][48] ) );
  NOR2_X1 U810 ( .A1(n347), .A2(n212), .ZN(\ab[51][47] ) );
  NOR2_X1 U811 ( .A1(n349), .A2(n211), .ZN(\ab[51][46] ) );
  NOR2_X1 U812 ( .A1(n351), .A2(n211), .ZN(\ab[51][45] ) );
  NOR2_X1 U813 ( .A1(n355), .A2(n211), .ZN(\ab[51][44] ) );
  NOR2_X1 U814 ( .A1(n357), .A2(n211), .ZN(\ab[51][43] ) );
  NOR2_X1 U815 ( .A1(n360), .A2(n211), .ZN(\ab[51][42] ) );
  NOR2_X1 U816 ( .A1(n361), .A2(n211), .ZN(\ab[51][41] ) );
  NOR2_X1 U817 ( .A1(n363), .A2(n211), .ZN(\ab[51][40] ) );
  NOR2_X1 U818 ( .A1(n441), .A2(n211), .ZN(\ab[51][3] ) );
  NOR2_X1 U819 ( .A1(n365), .A2(n212), .ZN(\ab[51][39] ) );
  NOR2_X1 U820 ( .A1(n368), .A2(n212), .ZN(\ab[51][38] ) );
  NOR2_X1 U821 ( .A1(n371), .A2(n212), .ZN(\ab[51][37] ) );
  NOR2_X1 U822 ( .A1(n474), .A2(n212), .ZN(\ab[51][36] ) );
  NOR2_X1 U823 ( .A1(n373), .A2(n212), .ZN(\ab[51][35] ) );
  NOR2_X1 U824 ( .A1(n375), .A2(n212), .ZN(\ab[51][34] ) );
  NOR2_X1 U825 ( .A1(n377), .A2(n212), .ZN(\ab[51][33] ) );
  NOR2_X1 U826 ( .A1(n380), .A2(n212), .ZN(\ab[51][32] ) );
  NOR2_X1 U827 ( .A1(n381), .A2(n212), .ZN(\ab[51][31] ) );
  NOR2_X1 U828 ( .A1(n383), .A2(n212), .ZN(\ab[51][30] ) );
  NOR2_X1 U829 ( .A1(n479), .A2(n212), .ZN(\ab[51][2] ) );
  NOR2_X1 U830 ( .A1(n386), .A2(n212), .ZN(\ab[51][29] ) );
  NOR2_X1 U831 ( .A1(n388), .A2(n212), .ZN(\ab[51][28] ) );
  NOR2_X1 U832 ( .A1(n390), .A2(n212), .ZN(\ab[51][27] ) );
  NOR2_X1 U833 ( .A1(n392), .A2(n211), .ZN(\ab[51][26] ) );
  NOR2_X1 U834 ( .A1(n394), .A2(n212), .ZN(\ab[51][25] ) );
  NOR2_X1 U835 ( .A1(n396), .A2(n211), .ZN(\ab[51][24] ) );
  NOR2_X1 U836 ( .A1(n398), .A2(n212), .ZN(\ab[51][23] ) );
  NOR2_X1 U837 ( .A1(n400), .A2(n212), .ZN(\ab[51][22] ) );
  NOR2_X1 U838 ( .A1(n402), .A2(n211), .ZN(\ab[51][21] ) );
  NOR2_X1 U839 ( .A1(n475), .A2(n211), .ZN(\ab[51][20] ) );
  NOR2_X1 U840 ( .A1(n444), .A2(n212), .ZN(\ab[51][1] ) );
  NOR2_X1 U841 ( .A1(n405), .A2(n211), .ZN(\ab[51][19] ) );
  NOR2_X1 U842 ( .A1(n407), .A2(n211), .ZN(\ab[51][18] ) );
  NOR2_X1 U843 ( .A1(n409), .A2(n211), .ZN(\ab[51][17] ) );
  NOR2_X1 U844 ( .A1(n412), .A2(n211), .ZN(\ab[51][16] ) );
  NOR2_X1 U845 ( .A1(n415), .A2(n211), .ZN(\ab[51][15] ) );
  NOR2_X1 U846 ( .A1(n418), .A2(n211), .ZN(\ab[51][14] ) );
  NOR2_X1 U847 ( .A1(n421), .A2(n211), .ZN(\ab[51][13] ) );
  NOR2_X1 U848 ( .A1(n424), .A2(n211), .ZN(\ab[51][12] ) );
  NOR2_X1 U849 ( .A1(n426), .A2(n211), .ZN(\ab[51][11] ) );
  NOR2_X1 U850 ( .A1(n427), .A2(n211), .ZN(\ab[51][10] ) );
  NOR2_X1 U851 ( .A1(n446), .A2(n211), .ZN(\ab[51][0] ) );
  NOR2_X1 U852 ( .A1(n429), .A2(n213), .ZN(\ab[50][9] ) );
  NOR2_X1 U853 ( .A1(n431), .A2(n213), .ZN(\ab[50][8] ) );
  NOR2_X1 U854 ( .A1(n433), .A2(n213), .ZN(\ab[50][7] ) );
  NOR2_X1 U855 ( .A1(n435), .A2(n213), .ZN(\ab[50][6] ) );
  NOR2_X1 U856 ( .A1(n437), .A2(n450), .ZN(\ab[50][5] ) );
  NOR2_X1 U857 ( .A1(n337), .A2(n213), .ZN(\ab[50][52] ) );
  NOR2_X1 U858 ( .A1(n340), .A2(n213), .ZN(\ab[50][51] ) );
  NOR2_X1 U859 ( .A1(n341), .A2(n213), .ZN(\ab[50][50] ) );
  NOR2_X1 U860 ( .A1(n439), .A2(n450), .ZN(\ab[50][4] ) );
  NOR2_X1 U861 ( .A1(n344), .A2(n214), .ZN(\ab[50][49] ) );
  NOR2_X1 U862 ( .A1(n346), .A2(n214), .ZN(\ab[50][48] ) );
  NOR2_X1 U863 ( .A1(n348), .A2(n214), .ZN(\ab[50][47] ) );
  NOR2_X1 U864 ( .A1(n350), .A2(n214), .ZN(\ab[50][46] ) );
  NOR2_X1 U865 ( .A1(n352), .A2(n214), .ZN(\ab[50][45] ) );
  NOR2_X1 U866 ( .A1(n355), .A2(n214), .ZN(\ab[50][44] ) );
  NOR2_X1 U867 ( .A1(n357), .A2(n214), .ZN(\ab[50][43] ) );
  NOR2_X1 U868 ( .A1(n360), .A2(n214), .ZN(\ab[50][42] ) );
  NOR2_X1 U869 ( .A1(n362), .A2(n214), .ZN(\ab[50][41] ) );
  NOR2_X1 U870 ( .A1(n364), .A2(n214), .ZN(\ab[50][40] ) );
  NOR2_X1 U871 ( .A1(n441), .A2(n214), .ZN(\ab[50][3] ) );
  NOR2_X1 U872 ( .A1(n366), .A2(n450), .ZN(\ab[50][39] ) );
  NOR2_X1 U873 ( .A1(n368), .A2(n214), .ZN(\ab[50][38] ) );
  NOR2_X1 U874 ( .A1(n371), .A2(n450), .ZN(\ab[50][37] ) );
  NOR2_X1 U875 ( .A1(n372), .A2(n213), .ZN(\ab[50][36] ) );
  NOR2_X1 U876 ( .A1(n374), .A2(n450), .ZN(\ab[50][35] ) );
  NOR2_X1 U877 ( .A1(n376), .A2(n450), .ZN(\ab[50][34] ) );
  NOR2_X1 U878 ( .A1(n378), .A2(n450), .ZN(\ab[50][33] ) );
  NOR2_X1 U879 ( .A1(n379), .A2(n450), .ZN(\ab[50][32] ) );
  NOR2_X1 U880 ( .A1(n382), .A2(n214), .ZN(\ab[50][31] ) );
  NOR2_X1 U881 ( .A1(n384), .A2(n450), .ZN(\ab[50][30] ) );
  NOR2_X1 U882 ( .A1(n479), .A2(n450), .ZN(\ab[50][2] ) );
  NOR2_X1 U883 ( .A1(n385), .A2(n450), .ZN(\ab[50][29] ) );
  NOR2_X1 U884 ( .A1(n388), .A2(n214), .ZN(\ab[50][28] ) );
  NOR2_X1 U885 ( .A1(n389), .A2(n214), .ZN(\ab[50][27] ) );
  NOR2_X1 U886 ( .A1(n391), .A2(n214), .ZN(\ab[50][26] ) );
  NOR2_X1 U887 ( .A1(n393), .A2(n213), .ZN(\ab[50][25] ) );
  NOR2_X1 U888 ( .A1(n396), .A2(n214), .ZN(\ab[50][24] ) );
  NOR2_X1 U889 ( .A1(n397), .A2(n213), .ZN(\ab[50][23] ) );
  NOR2_X1 U890 ( .A1(n399), .A2(n213), .ZN(\ab[50][22] ) );
  NOR2_X1 U891 ( .A1(n401), .A2(n213), .ZN(\ab[50][21] ) );
  NOR2_X1 U892 ( .A1(n403), .A2(n213), .ZN(\ab[50][20] ) );
  NOR2_X1 U893 ( .A1(n444), .A2(n213), .ZN(\ab[50][1] ) );
  NOR2_X1 U894 ( .A1(n405), .A2(n213), .ZN(\ab[50][19] ) );
  NOR2_X1 U895 ( .A1(n407), .A2(n213), .ZN(\ab[50][18] ) );
  NOR2_X1 U896 ( .A1(n408), .A2(n213), .ZN(\ab[50][17] ) );
  NOR2_X1 U897 ( .A1(n412), .A2(n213), .ZN(\ab[50][16] ) );
  NOR2_X1 U898 ( .A1(n415), .A2(n213), .ZN(\ab[50][15] ) );
  NOR2_X1 U899 ( .A1(n418), .A2(n213), .ZN(\ab[50][14] ) );
  NOR2_X1 U900 ( .A1(n421), .A2(n213), .ZN(\ab[50][13] ) );
  NOR2_X1 U901 ( .A1(n424), .A2(n213), .ZN(\ab[50][12] ) );
  NOR2_X1 U902 ( .A1(n425), .A2(n213), .ZN(\ab[50][11] ) );
  NOR2_X1 U903 ( .A1(n477), .A2(n213), .ZN(\ab[50][10] ) );
  NOR2_X1 U904 ( .A1(n480), .A2(n213), .ZN(\ab[50][0] ) );
  NOR2_X1 U905 ( .A1(n429), .A2(n323), .ZN(\ab[4][9] ) );
  NOR2_X1 U906 ( .A1(n431), .A2(n324), .ZN(\ab[4][8] ) );
  NOR2_X1 U907 ( .A1(n433), .A2(n323), .ZN(\ab[4][7] ) );
  NOR2_X1 U908 ( .A1(n435), .A2(n324), .ZN(\ab[4][6] ) );
  NOR2_X1 U909 ( .A1(n437), .A2(n323), .ZN(\ab[4][5] ) );
  NOR2_X1 U910 ( .A1(n337), .A2(n323), .ZN(\ab[4][52] ) );
  NOR2_X1 U911 ( .A1(n340), .A2(n324), .ZN(\ab[4][51] ) );
  NOR2_X1 U912 ( .A1(n341), .A2(n324), .ZN(\ab[4][50] ) );
  NOR2_X1 U913 ( .A1(n439), .A2(n324), .ZN(\ab[4][4] ) );
  NOR2_X1 U914 ( .A1(n344), .A2(n324), .ZN(\ab[4][49] ) );
  NOR2_X1 U915 ( .A1(n346), .A2(n324), .ZN(\ab[4][48] ) );
  NOR2_X1 U916 ( .A1(n348), .A2(n324), .ZN(\ab[4][47] ) );
  NOR2_X1 U917 ( .A1(n350), .A2(n324), .ZN(\ab[4][46] ) );
  NOR2_X1 U918 ( .A1(n352), .A2(n323), .ZN(\ab[4][45] ) );
  NOR2_X1 U919 ( .A1(n355), .A2(n323), .ZN(\ab[4][44] ) );
  NOR2_X1 U920 ( .A1(n357), .A2(n323), .ZN(\ab[4][43] ) );
  NOR2_X1 U921 ( .A1(n360), .A2(n323), .ZN(\ab[4][42] ) );
  NOR2_X1 U922 ( .A1(n362), .A2(n323), .ZN(\ab[4][41] ) );
  NOR2_X1 U923 ( .A1(n364), .A2(n323), .ZN(\ab[4][40] ) );
  NOR2_X1 U924 ( .A1(n441), .A2(n323), .ZN(\ab[4][3] ) );
  NOR2_X1 U925 ( .A1(n366), .A2(n323), .ZN(\ab[4][39] ) );
  NOR2_X1 U926 ( .A1(n368), .A2(n323), .ZN(\ab[4][38] ) );
  NOR2_X1 U927 ( .A1(n371), .A2(n323), .ZN(\ab[4][37] ) );
  NOR2_X1 U928 ( .A1(n474), .A2(n323), .ZN(\ab[4][36] ) );
  NOR2_X1 U929 ( .A1(n374), .A2(n323), .ZN(\ab[4][35] ) );
  NOR2_X1 U930 ( .A1(n376), .A2(n323), .ZN(\ab[4][34] ) );
  NOR2_X1 U931 ( .A1(n378), .A2(n323), .ZN(\ab[4][33] ) );
  NOR2_X1 U932 ( .A1(n380), .A2(n323), .ZN(\ab[4][32] ) );
  NOR2_X1 U933 ( .A1(n382), .A2(n323), .ZN(\ab[4][31] ) );
  NOR2_X1 U934 ( .A1(n384), .A2(n323), .ZN(\ab[4][30] ) );
  NOR2_X1 U935 ( .A1(n479), .A2(n323), .ZN(\ab[4][2] ) );
  NOR2_X1 U936 ( .A1(n386), .A2(n323), .ZN(\ab[4][29] ) );
  NOR2_X1 U937 ( .A1(n388), .A2(n323), .ZN(\ab[4][28] ) );
  NOR2_X1 U938 ( .A1(n390), .A2(n323), .ZN(\ab[4][27] ) );
  NOR2_X1 U939 ( .A1(n392), .A2(n323), .ZN(\ab[4][26] ) );
  NOR2_X1 U940 ( .A1(n394), .A2(n323), .ZN(\ab[4][25] ) );
  NOR2_X1 U941 ( .A1(n396), .A2(n323), .ZN(\ab[4][24] ) );
  NOR2_X1 U942 ( .A1(n398), .A2(n323), .ZN(\ab[4][23] ) );
  NOR2_X1 U943 ( .A1(n400), .A2(n323), .ZN(\ab[4][22] ) );
  NOR2_X1 U944 ( .A1(n402), .A2(n323), .ZN(\ab[4][21] ) );
  NOR2_X1 U945 ( .A1(n475), .A2(n323), .ZN(\ab[4][20] ) );
  NOR2_X1 U946 ( .A1(n444), .A2(n323), .ZN(\ab[4][1] ) );
  NOR2_X1 U947 ( .A1(n405), .A2(n324), .ZN(\ab[4][19] ) );
  NOR2_X1 U948 ( .A1(n407), .A2(n323), .ZN(\ab[4][18] ) );
  NOR2_X1 U949 ( .A1(n409), .A2(n324), .ZN(\ab[4][17] ) );
  NOR2_X1 U950 ( .A1(n412), .A2(n323), .ZN(\ab[4][16] ) );
  NOR2_X1 U951 ( .A1(n415), .A2(n324), .ZN(\ab[4][15] ) );
  NOR2_X1 U952 ( .A1(n418), .A2(n324), .ZN(\ab[4][14] ) );
  NOR2_X1 U953 ( .A1(n421), .A2(n323), .ZN(\ab[4][13] ) );
  NOR2_X1 U954 ( .A1(n424), .A2(n324), .ZN(\ab[4][12] ) );
  NOR2_X1 U955 ( .A1(n426), .A2(n323), .ZN(\ab[4][11] ) );
  NOR2_X1 U956 ( .A1(n477), .A2(n324), .ZN(\ab[4][10] ) );
  NOR2_X1 U957 ( .A1(n480), .A2(n324), .ZN(\ab[4][0] ) );
  NOR2_X1 U958 ( .A1(n429), .A2(n215), .ZN(\ab[49][9] ) );
  NOR2_X1 U959 ( .A1(n431), .A2(n215), .ZN(\ab[49][8] ) );
  NOR2_X1 U960 ( .A1(n433), .A2(n216), .ZN(\ab[49][7] ) );
  NOR2_X1 U961 ( .A1(n435), .A2(n216), .ZN(\ab[49][6] ) );
  NOR2_X1 U962 ( .A1(n437), .A2(n216), .ZN(\ab[49][5] ) );
  NOR2_X1 U963 ( .A1(n337), .A2(n215), .ZN(\ab[49][52] ) );
  NOR2_X1 U964 ( .A1(n339), .A2(n215), .ZN(\ab[49][51] ) );
  NOR2_X1 U965 ( .A1(n341), .A2(n215), .ZN(\ab[49][50] ) );
  NOR2_X1 U966 ( .A1(n439), .A2(n217), .ZN(\ab[49][4] ) );
  NOR2_X1 U967 ( .A1(n344), .A2(n217), .ZN(\ab[49][49] ) );
  NOR2_X1 U968 ( .A1(n345), .A2(n217), .ZN(\ab[49][48] ) );
  NOR2_X1 U969 ( .A1(n347), .A2(n217), .ZN(\ab[49][47] ) );
  NOR2_X1 U970 ( .A1(n349), .A2(n217), .ZN(\ab[49][46] ) );
  NOR2_X1 U971 ( .A1(n351), .A2(n217), .ZN(\ab[49][45] ) );
  NOR2_X1 U972 ( .A1(n354), .A2(n217), .ZN(\ab[49][44] ) );
  NOR2_X1 U973 ( .A1(n357), .A2(n217), .ZN(\ab[49][43] ) );
  NOR2_X1 U974 ( .A1(n359), .A2(n217), .ZN(\ab[49][42] ) );
  NOR2_X1 U975 ( .A1(n361), .A2(n217), .ZN(\ab[49][41] ) );
  NOR2_X1 U976 ( .A1(n363), .A2(n217), .ZN(\ab[49][40] ) );
  NOR2_X1 U977 ( .A1(n478), .A2(n217), .ZN(\ab[49][3] ) );
  NOR2_X1 U978 ( .A1(n365), .A2(n216), .ZN(\ab[49][39] ) );
  NOR2_X1 U979 ( .A1(n367), .A2(n216), .ZN(\ab[49][38] ) );
  NOR2_X1 U980 ( .A1(n371), .A2(n216), .ZN(\ab[49][37] ) );
  NOR2_X1 U981 ( .A1(n474), .A2(n216), .ZN(\ab[49][36] ) );
  NOR2_X1 U982 ( .A1(n373), .A2(n216), .ZN(\ab[49][35] ) );
  NOR2_X1 U983 ( .A1(n375), .A2(n216), .ZN(\ab[49][34] ) );
  NOR2_X1 U984 ( .A1(n377), .A2(n216), .ZN(\ab[49][33] ) );
  NOR2_X1 U985 ( .A1(n380), .A2(n216), .ZN(\ab[49][32] ) );
  NOR2_X1 U986 ( .A1(n381), .A2(n216), .ZN(\ab[49][31] ) );
  NOR2_X1 U987 ( .A1(n383), .A2(n216), .ZN(\ab[49][30] ) );
  NOR2_X1 U988 ( .A1(n479), .A2(n216), .ZN(\ab[49][2] ) );
  NOR2_X1 U989 ( .A1(n386), .A2(n215), .ZN(\ab[49][29] ) );
  NOR2_X1 U990 ( .A1(n388), .A2(n215), .ZN(\ab[49][28] ) );
  NOR2_X1 U991 ( .A1(n390), .A2(n215), .ZN(\ab[49][27] ) );
  NOR2_X1 U992 ( .A1(n392), .A2(n215), .ZN(\ab[49][26] ) );
  NOR2_X1 U993 ( .A1(n394), .A2(n215), .ZN(\ab[49][25] ) );
  NOR2_X1 U994 ( .A1(n395), .A2(n215), .ZN(\ab[49][24] ) );
  NOR2_X1 U995 ( .A1(n398), .A2(n215), .ZN(\ab[49][23] ) );
  NOR2_X1 U996 ( .A1(n400), .A2(n215), .ZN(\ab[49][22] ) );
  NOR2_X1 U997 ( .A1(n402), .A2(n215), .ZN(\ab[49][21] ) );
  NOR2_X1 U998 ( .A1(n475), .A2(n215), .ZN(\ab[49][20] ) );
  NOR2_X1 U999 ( .A1(n444), .A2(n215), .ZN(\ab[49][1] ) );
  NOR2_X1 U1000 ( .A1(n405), .A2(n215), .ZN(\ab[49][19] ) );
  NOR2_X1 U1001 ( .A1(n407), .A2(n215), .ZN(\ab[49][18] ) );
  NOR2_X1 U1002 ( .A1(n409), .A2(n215), .ZN(\ab[49][17] ) );
  NOR2_X1 U1003 ( .A1(n411), .A2(n215), .ZN(\ab[49][16] ) );
  NOR2_X1 U1004 ( .A1(n414), .A2(n215), .ZN(\ab[49][15] ) );
  NOR2_X1 U1005 ( .A1(n417), .A2(n215), .ZN(\ab[49][14] ) );
  NOR2_X1 U1006 ( .A1(n420), .A2(n215), .ZN(\ab[49][13] ) );
  NOR2_X1 U1007 ( .A1(n423), .A2(n215), .ZN(\ab[49][12] ) );
  NOR2_X1 U1008 ( .A1(n426), .A2(n215), .ZN(\ab[49][11] ) );
  NOR2_X1 U1009 ( .A1(n427), .A2(n215), .ZN(\ab[49][10] ) );
  NOR2_X1 U1010 ( .A1(n446), .A2(n215), .ZN(\ab[49][0] ) );
  NOR2_X1 U1011 ( .A1(n429), .A2(n218), .ZN(\ab[48][9] ) );
  NOR2_X1 U1012 ( .A1(n431), .A2(n219), .ZN(\ab[48][8] ) );
  NOR2_X1 U1013 ( .A1(n433), .A2(n219), .ZN(\ab[48][7] ) );
  NOR2_X1 U1014 ( .A1(n435), .A2(n220), .ZN(\ab[48][6] ) );
  NOR2_X1 U1015 ( .A1(n437), .A2(n219), .ZN(\ab[48][5] ) );
  NOR2_X1 U1016 ( .A1(n337), .A2(n218), .ZN(\ab[48][52] ) );
  NOR2_X1 U1017 ( .A1(n339), .A2(n218), .ZN(\ab[48][51] ) );
  NOR2_X1 U1018 ( .A1(n341), .A2(n218), .ZN(\ab[48][50] ) );
  NOR2_X1 U1019 ( .A1(n439), .A2(n220), .ZN(\ab[48][4] ) );
  NOR2_X1 U1020 ( .A1(n344), .A2(n220), .ZN(\ab[48][49] ) );
  NOR2_X1 U1021 ( .A1(n346), .A2(n220), .ZN(\ab[48][48] ) );
  NOR2_X1 U1022 ( .A1(n348), .A2(n220), .ZN(\ab[48][47] ) );
  NOR2_X1 U1023 ( .A1(n350), .A2(n220), .ZN(\ab[48][46] ) );
  NOR2_X1 U1024 ( .A1(n352), .A2(n220), .ZN(\ab[48][45] ) );
  NOR2_X1 U1025 ( .A1(n354), .A2(n220), .ZN(\ab[48][44] ) );
  NOR2_X1 U1026 ( .A1(n357), .A2(n220), .ZN(\ab[48][43] ) );
  NOR2_X1 U1027 ( .A1(n359), .A2(n220), .ZN(\ab[48][42] ) );
  NOR2_X1 U1028 ( .A1(n362), .A2(n220), .ZN(\ab[48][41] ) );
  NOR2_X1 U1029 ( .A1(n364), .A2(n220), .ZN(\ab[48][40] ) );
  NOR2_X1 U1030 ( .A1(n478), .A2(n220), .ZN(\ab[48][3] ) );
  NOR2_X1 U1031 ( .A1(n366), .A2(n219), .ZN(\ab[48][39] ) );
  NOR2_X1 U1032 ( .A1(n367), .A2(n219), .ZN(\ab[48][38] ) );
  NOR2_X1 U1033 ( .A1(n371), .A2(n219), .ZN(\ab[48][37] ) );
  NOR2_X1 U1034 ( .A1(n372), .A2(n219), .ZN(\ab[48][36] ) );
  NOR2_X1 U1035 ( .A1(n374), .A2(n219), .ZN(\ab[48][35] ) );
  NOR2_X1 U1036 ( .A1(n376), .A2(n219), .ZN(\ab[48][34] ) );
  NOR2_X1 U1037 ( .A1(n378), .A2(n219), .ZN(\ab[48][33] ) );
  NOR2_X1 U1038 ( .A1(n379), .A2(n219), .ZN(\ab[48][32] ) );
  NOR2_X1 U1039 ( .A1(n382), .A2(n219), .ZN(\ab[48][31] ) );
  NOR2_X1 U1040 ( .A1(n384), .A2(n219), .ZN(\ab[48][30] ) );
  NOR2_X1 U1041 ( .A1(n479), .A2(n219), .ZN(\ab[48][2] ) );
  NOR2_X1 U1042 ( .A1(n385), .A2(n218), .ZN(\ab[48][29] ) );
  NOR2_X1 U1043 ( .A1(n388), .A2(n218), .ZN(\ab[48][28] ) );
  NOR2_X1 U1044 ( .A1(n389), .A2(n218), .ZN(\ab[48][27] ) );
  NOR2_X1 U1045 ( .A1(n391), .A2(n218), .ZN(\ab[48][26] ) );
  NOR2_X1 U1046 ( .A1(n394), .A2(n218), .ZN(\ab[48][25] ) );
  NOR2_X1 U1047 ( .A1(n396), .A2(n218), .ZN(\ab[48][24] ) );
  NOR2_X1 U1048 ( .A1(n397), .A2(n218), .ZN(\ab[48][23] ) );
  NOR2_X1 U1049 ( .A1(n399), .A2(n218), .ZN(\ab[48][22] ) );
  NOR2_X1 U1050 ( .A1(n401), .A2(n218), .ZN(\ab[48][21] ) );
  NOR2_X1 U1051 ( .A1(n403), .A2(n218), .ZN(\ab[48][20] ) );
  NOR2_X1 U1052 ( .A1(n444), .A2(n218), .ZN(\ab[48][1] ) );
  NOR2_X1 U1053 ( .A1(n405), .A2(n218), .ZN(\ab[48][19] ) );
  NOR2_X1 U1054 ( .A1(n407), .A2(n218), .ZN(\ab[48][18] ) );
  NOR2_X1 U1055 ( .A1(n408), .A2(n218), .ZN(\ab[48][17] ) );
  NOR2_X1 U1056 ( .A1(n411), .A2(n218), .ZN(\ab[48][16] ) );
  NOR2_X1 U1057 ( .A1(n414), .A2(n218), .ZN(\ab[48][15] ) );
  NOR2_X1 U1058 ( .A1(n417), .A2(n218), .ZN(\ab[48][14] ) );
  NOR2_X1 U1059 ( .A1(n420), .A2(n218), .ZN(\ab[48][13] ) );
  NOR2_X1 U1060 ( .A1(n423), .A2(n218), .ZN(\ab[48][12] ) );
  NOR2_X1 U1061 ( .A1(n425), .A2(n218), .ZN(\ab[48][11] ) );
  NOR2_X1 U1062 ( .A1(n477), .A2(n218), .ZN(\ab[48][10] ) );
  NOR2_X1 U1063 ( .A1(n480), .A2(n218), .ZN(\ab[48][0] ) );
  NOR2_X1 U1064 ( .A1(n429), .A2(n221), .ZN(\ab[47][9] ) );
  NOR2_X1 U1065 ( .A1(n431), .A2(n222), .ZN(\ab[47][8] ) );
  NOR2_X1 U1066 ( .A1(n433), .A2(n222), .ZN(\ab[47][7] ) );
  NOR2_X1 U1067 ( .A1(n435), .A2(n223), .ZN(\ab[47][6] ) );
  NOR2_X1 U1068 ( .A1(n437), .A2(n222), .ZN(\ab[47][5] ) );
  NOR2_X1 U1069 ( .A1(n337), .A2(n221), .ZN(\ab[47][52] ) );
  NOR2_X1 U1070 ( .A1(n339), .A2(n221), .ZN(\ab[47][51] ) );
  NOR2_X1 U1071 ( .A1(n341), .A2(n221), .ZN(\ab[47][50] ) );
  NOR2_X1 U1072 ( .A1(n439), .A2(n221), .ZN(\ab[47][4] ) );
  NOR2_X1 U1073 ( .A1(n344), .A2(n223), .ZN(\ab[47][49] ) );
  NOR2_X1 U1074 ( .A1(n345), .A2(n223), .ZN(\ab[47][48] ) );
  NOR2_X1 U1075 ( .A1(n347), .A2(n223), .ZN(\ab[47][47] ) );
  NOR2_X1 U1076 ( .A1(n349), .A2(n223), .ZN(\ab[47][46] ) );
  NOR2_X1 U1077 ( .A1(n351), .A2(n223), .ZN(\ab[47][45] ) );
  NOR2_X1 U1078 ( .A1(n354), .A2(n223), .ZN(\ab[47][44] ) );
  NOR2_X1 U1079 ( .A1(n357), .A2(n223), .ZN(\ab[47][43] ) );
  NOR2_X1 U1080 ( .A1(n359), .A2(n223), .ZN(\ab[47][42] ) );
  NOR2_X1 U1081 ( .A1(n361), .A2(n223), .ZN(\ab[47][41] ) );
  NOR2_X1 U1082 ( .A1(n363), .A2(n223), .ZN(\ab[47][40] ) );
  NOR2_X1 U1083 ( .A1(n478), .A2(n223), .ZN(\ab[47][3] ) );
  NOR2_X1 U1084 ( .A1(n365), .A2(n222), .ZN(\ab[47][39] ) );
  NOR2_X1 U1085 ( .A1(n367), .A2(n222), .ZN(\ab[47][38] ) );
  NOR2_X1 U1086 ( .A1(n371), .A2(n222), .ZN(\ab[47][37] ) );
  NOR2_X1 U1087 ( .A1(n474), .A2(n222), .ZN(\ab[47][36] ) );
  NOR2_X1 U1088 ( .A1(n373), .A2(n222), .ZN(\ab[47][35] ) );
  NOR2_X1 U1089 ( .A1(n375), .A2(n222), .ZN(\ab[47][34] ) );
  NOR2_X1 U1090 ( .A1(n377), .A2(n222), .ZN(\ab[47][33] ) );
  NOR2_X1 U1091 ( .A1(n380), .A2(n222), .ZN(\ab[47][32] ) );
  NOR2_X1 U1092 ( .A1(n381), .A2(n222), .ZN(\ab[47][31] ) );
  NOR2_X1 U1093 ( .A1(n383), .A2(n222), .ZN(\ab[47][30] ) );
  NOR2_X1 U1094 ( .A1(n479), .A2(n222), .ZN(\ab[47][2] ) );
  NOR2_X1 U1095 ( .A1(n386), .A2(n221), .ZN(\ab[47][29] ) );
  NOR2_X1 U1096 ( .A1(n388), .A2(n221), .ZN(\ab[47][28] ) );
  NOR2_X1 U1097 ( .A1(n390), .A2(n221), .ZN(\ab[47][27] ) );
  NOR2_X1 U1098 ( .A1(n392), .A2(n221), .ZN(\ab[47][26] ) );
  NOR2_X1 U1099 ( .A1(n393), .A2(n221), .ZN(\ab[47][25] ) );
  NOR2_X1 U1100 ( .A1(n395), .A2(n221), .ZN(\ab[47][24] ) );
  NOR2_X1 U1101 ( .A1(n398), .A2(n221), .ZN(\ab[47][23] ) );
  NOR2_X1 U1102 ( .A1(n400), .A2(n221), .ZN(\ab[47][22] ) );
  NOR2_X1 U1103 ( .A1(n402), .A2(n221), .ZN(\ab[47][21] ) );
  NOR2_X1 U1104 ( .A1(n475), .A2(n221), .ZN(\ab[47][20] ) );
  NOR2_X1 U1105 ( .A1(n444), .A2(n221), .ZN(\ab[47][1] ) );
  NOR2_X1 U1106 ( .A1(n405), .A2(n221), .ZN(\ab[47][19] ) );
  NOR2_X1 U1107 ( .A1(n407), .A2(n221), .ZN(\ab[47][18] ) );
  NOR2_X1 U1108 ( .A1(n409), .A2(n221), .ZN(\ab[47][17] ) );
  NOR2_X1 U1109 ( .A1(n411), .A2(n221), .ZN(\ab[47][16] ) );
  NOR2_X1 U1110 ( .A1(n414), .A2(n221), .ZN(\ab[47][15] ) );
  NOR2_X1 U1111 ( .A1(n417), .A2(n221), .ZN(\ab[47][14] ) );
  NOR2_X1 U1112 ( .A1(n420), .A2(n221), .ZN(\ab[47][13] ) );
  NOR2_X1 U1113 ( .A1(n423), .A2(n221), .ZN(\ab[47][12] ) );
  NOR2_X1 U1114 ( .A1(n426), .A2(n221), .ZN(\ab[47][11] ) );
  NOR2_X1 U1115 ( .A1(n427), .A2(n221), .ZN(\ab[47][10] ) );
  NOR2_X1 U1116 ( .A1(n446), .A2(n221), .ZN(\ab[47][0] ) );
  NOR2_X1 U1117 ( .A1(n429), .A2(n451), .ZN(\ab[46][9] ) );
  NOR2_X1 U1118 ( .A1(n431), .A2(n451), .ZN(\ab[46][8] ) );
  NOR2_X1 U1119 ( .A1(n433), .A2(n451), .ZN(\ab[46][7] ) );
  NOR2_X1 U1120 ( .A1(n435), .A2(n451), .ZN(\ab[46][6] ) );
  NOR2_X1 U1121 ( .A1(n437), .A2(n225), .ZN(\ab[46][5] ) );
  NOR2_X1 U1122 ( .A1(n337), .A2(n451), .ZN(\ab[46][52] ) );
  NOR2_X1 U1123 ( .A1(n339), .A2(n225), .ZN(\ab[46][51] ) );
  NOR2_X1 U1124 ( .A1(n341), .A2(n225), .ZN(\ab[46][50] ) );
  NOR2_X1 U1125 ( .A1(n439), .A2(n225), .ZN(\ab[46][4] ) );
  NOR2_X1 U1126 ( .A1(n344), .A2(n224), .ZN(\ab[46][49] ) );
  NOR2_X1 U1127 ( .A1(n346), .A2(n224), .ZN(\ab[46][48] ) );
  NOR2_X1 U1128 ( .A1(n348), .A2(n224), .ZN(\ab[46][47] ) );
  NOR2_X1 U1129 ( .A1(n350), .A2(n224), .ZN(\ab[46][46] ) );
  NOR2_X1 U1130 ( .A1(n352), .A2(n224), .ZN(\ab[46][45] ) );
  NOR2_X1 U1131 ( .A1(n354), .A2(n224), .ZN(\ab[46][44] ) );
  NOR2_X1 U1132 ( .A1(n357), .A2(n224), .ZN(\ab[46][43] ) );
  NOR2_X1 U1133 ( .A1(n359), .A2(n224), .ZN(\ab[46][42] ) );
  NOR2_X1 U1134 ( .A1(n362), .A2(n224), .ZN(\ab[46][41] ) );
  NOR2_X1 U1135 ( .A1(n364), .A2(n224), .ZN(\ab[46][40] ) );
  NOR2_X1 U1136 ( .A1(n478), .A2(n224), .ZN(\ab[46][3] ) );
  NOR2_X1 U1137 ( .A1(n366), .A2(n225), .ZN(\ab[46][39] ) );
  NOR2_X1 U1138 ( .A1(n367), .A2(n225), .ZN(\ab[46][38] ) );
  NOR2_X1 U1139 ( .A1(n371), .A2(n225), .ZN(\ab[46][37] ) );
  NOR2_X1 U1140 ( .A1(n372), .A2(n225), .ZN(\ab[46][36] ) );
  NOR2_X1 U1141 ( .A1(n374), .A2(n225), .ZN(\ab[46][35] ) );
  NOR2_X1 U1142 ( .A1(n376), .A2(n225), .ZN(\ab[46][34] ) );
  NOR2_X1 U1143 ( .A1(n378), .A2(n225), .ZN(\ab[46][33] ) );
  NOR2_X1 U1144 ( .A1(n379), .A2(n225), .ZN(\ab[46][32] ) );
  NOR2_X1 U1145 ( .A1(n382), .A2(n225), .ZN(\ab[46][31] ) );
  NOR2_X1 U1146 ( .A1(n384), .A2(n225), .ZN(\ab[46][30] ) );
  NOR2_X1 U1147 ( .A1(n479), .A2(n225), .ZN(\ab[46][2] ) );
  NOR2_X1 U1148 ( .A1(n385), .A2(n225), .ZN(\ab[46][29] ) );
  NOR2_X1 U1149 ( .A1(n388), .A2(n225), .ZN(\ab[46][28] ) );
  NOR2_X1 U1150 ( .A1(n389), .A2(n225), .ZN(\ab[46][27] ) );
  NOR2_X1 U1151 ( .A1(n391), .A2(n225), .ZN(\ab[46][26] ) );
  NOR2_X1 U1152 ( .A1(n394), .A2(n225), .ZN(\ab[46][25] ) );
  NOR2_X1 U1153 ( .A1(n396), .A2(n225), .ZN(\ab[46][24] ) );
  NOR2_X1 U1154 ( .A1(n397), .A2(n225), .ZN(\ab[46][23] ) );
  NOR2_X1 U1155 ( .A1(n399), .A2(n225), .ZN(\ab[46][22] ) );
  NOR2_X1 U1156 ( .A1(n401), .A2(n225), .ZN(\ab[46][21] ) );
  NOR2_X1 U1157 ( .A1(n403), .A2(n225), .ZN(\ab[46][20] ) );
  NOR2_X1 U1158 ( .A1(n444), .A2(n225), .ZN(\ab[46][1] ) );
  NOR2_X1 U1159 ( .A1(n405), .A2(n224), .ZN(\ab[46][19] ) );
  NOR2_X1 U1160 ( .A1(n407), .A2(n224), .ZN(\ab[46][18] ) );
  NOR2_X1 U1161 ( .A1(n408), .A2(n224), .ZN(\ab[46][17] ) );
  NOR2_X1 U1162 ( .A1(n411), .A2(n224), .ZN(\ab[46][16] ) );
  NOR2_X1 U1163 ( .A1(n414), .A2(n224), .ZN(\ab[46][15] ) );
  NOR2_X1 U1164 ( .A1(n417), .A2(n224), .ZN(\ab[46][14] ) );
  NOR2_X1 U1165 ( .A1(n420), .A2(n224), .ZN(\ab[46][13] ) );
  NOR2_X1 U1166 ( .A1(n423), .A2(n224), .ZN(\ab[46][12] ) );
  NOR2_X1 U1167 ( .A1(n425), .A2(n224), .ZN(\ab[46][11] ) );
  NOR2_X1 U1168 ( .A1(n477), .A2(n224), .ZN(\ab[46][10] ) );
  NOR2_X1 U1169 ( .A1(n480), .A2(n224), .ZN(\ab[46][0] ) );
  NOR2_X1 U1170 ( .A1(n429), .A2(n228), .ZN(\ab[45][9] ) );
  NOR2_X1 U1171 ( .A1(n431), .A2(n227), .ZN(\ab[45][8] ) );
  NOR2_X1 U1172 ( .A1(n433), .A2(n226), .ZN(\ab[45][7] ) );
  NOR2_X1 U1173 ( .A1(n435), .A2(n226), .ZN(\ab[45][6] ) );
  NOR2_X1 U1174 ( .A1(n437), .A2(n226), .ZN(\ab[45][5] ) );
  NOR2_X1 U1175 ( .A1(n337), .A2(n226), .ZN(\ab[45][52] ) );
  NOR2_X1 U1176 ( .A1(n339), .A2(n226), .ZN(\ab[45][51] ) );
  NOR2_X1 U1177 ( .A1(n341), .A2(n226), .ZN(\ab[45][50] ) );
  NOR2_X1 U1178 ( .A1(n439), .A2(n226), .ZN(\ab[45][4] ) );
  NOR2_X1 U1179 ( .A1(n344), .A2(n228), .ZN(\ab[45][49] ) );
  NOR2_X1 U1180 ( .A1(n345), .A2(n228), .ZN(\ab[45][48] ) );
  NOR2_X1 U1181 ( .A1(n347), .A2(n228), .ZN(\ab[45][47] ) );
  NOR2_X1 U1182 ( .A1(n349), .A2(n228), .ZN(\ab[45][46] ) );
  NOR2_X1 U1183 ( .A1(n351), .A2(n228), .ZN(\ab[45][45] ) );
  NOR2_X1 U1184 ( .A1(n354), .A2(n228), .ZN(\ab[45][44] ) );
  NOR2_X1 U1185 ( .A1(n357), .A2(n228), .ZN(\ab[45][43] ) );
  NOR2_X1 U1186 ( .A1(n359), .A2(n228), .ZN(\ab[45][42] ) );
  NOR2_X1 U1187 ( .A1(n361), .A2(n228), .ZN(\ab[45][41] ) );
  NOR2_X1 U1188 ( .A1(n363), .A2(n228), .ZN(\ab[45][40] ) );
  NOR2_X1 U1189 ( .A1(n478), .A2(n228), .ZN(\ab[45][3] ) );
  NOR2_X1 U1190 ( .A1(n365), .A2(n227), .ZN(\ab[45][39] ) );
  NOR2_X1 U1191 ( .A1(n367), .A2(n227), .ZN(\ab[45][38] ) );
  NOR2_X1 U1192 ( .A1(n371), .A2(n227), .ZN(\ab[45][37] ) );
  NOR2_X1 U1193 ( .A1(n474), .A2(n227), .ZN(\ab[45][36] ) );
  NOR2_X1 U1194 ( .A1(n373), .A2(n227), .ZN(\ab[45][35] ) );
  NOR2_X1 U1195 ( .A1(n375), .A2(n227), .ZN(\ab[45][34] ) );
  NOR2_X1 U1196 ( .A1(n377), .A2(n227), .ZN(\ab[45][33] ) );
  NOR2_X1 U1197 ( .A1(n380), .A2(n227), .ZN(\ab[45][32] ) );
  NOR2_X1 U1198 ( .A1(n381), .A2(n227), .ZN(\ab[45][31] ) );
  NOR2_X1 U1199 ( .A1(n383), .A2(n227), .ZN(\ab[45][30] ) );
  NOR2_X1 U1200 ( .A1(n479), .A2(n227), .ZN(\ab[45][2] ) );
  NOR2_X1 U1201 ( .A1(n386), .A2(n226), .ZN(\ab[45][29] ) );
  NOR2_X1 U1202 ( .A1(n388), .A2(n226), .ZN(\ab[45][28] ) );
  NOR2_X1 U1203 ( .A1(n390), .A2(n226), .ZN(\ab[45][27] ) );
  NOR2_X1 U1204 ( .A1(n392), .A2(n226), .ZN(\ab[45][26] ) );
  NOR2_X1 U1205 ( .A1(n393), .A2(n226), .ZN(\ab[45][25] ) );
  NOR2_X1 U1206 ( .A1(n395), .A2(n226), .ZN(\ab[45][24] ) );
  NOR2_X1 U1207 ( .A1(n398), .A2(n226), .ZN(\ab[45][23] ) );
  NOR2_X1 U1208 ( .A1(n400), .A2(n226), .ZN(\ab[45][22] ) );
  NOR2_X1 U1209 ( .A1(n402), .A2(n226), .ZN(\ab[45][21] ) );
  NOR2_X1 U1210 ( .A1(n475), .A2(n226), .ZN(\ab[45][20] ) );
  NOR2_X1 U1211 ( .A1(n444), .A2(n226), .ZN(\ab[45][1] ) );
  NOR2_X1 U1212 ( .A1(n405), .A2(n452), .ZN(\ab[45][19] ) );
  NOR2_X1 U1213 ( .A1(n407), .A2(n452), .ZN(\ab[45][18] ) );
  NOR2_X1 U1214 ( .A1(n409), .A2(n452), .ZN(\ab[45][17] ) );
  NOR2_X1 U1215 ( .A1(n411), .A2(n452), .ZN(\ab[45][16] ) );
  NOR2_X1 U1216 ( .A1(n414), .A2(n452), .ZN(\ab[45][15] ) );
  NOR2_X1 U1217 ( .A1(n417), .A2(n452), .ZN(\ab[45][14] ) );
  NOR2_X1 U1218 ( .A1(n420), .A2(n228), .ZN(\ab[45][13] ) );
  NOR2_X1 U1219 ( .A1(n423), .A2(n226), .ZN(\ab[45][12] ) );
  NOR2_X1 U1220 ( .A1(n426), .A2(n226), .ZN(\ab[45][11] ) );
  NOR2_X1 U1221 ( .A1(n427), .A2(n227), .ZN(\ab[45][10] ) );
  NOR2_X1 U1222 ( .A1(n446), .A2(n452), .ZN(\ab[45][0] ) );
  NOR2_X1 U1223 ( .A1(n429), .A2(n453), .ZN(\ab[44][9] ) );
  NOR2_X1 U1224 ( .A1(n431), .A2(n230), .ZN(\ab[44][8] ) );
  NOR2_X1 U1225 ( .A1(n433), .A2(n229), .ZN(\ab[44][7] ) );
  NOR2_X1 U1226 ( .A1(n435), .A2(n229), .ZN(\ab[44][6] ) );
  NOR2_X1 U1227 ( .A1(n437), .A2(n229), .ZN(\ab[44][5] ) );
  NOR2_X1 U1228 ( .A1(n337), .A2(n229), .ZN(\ab[44][52] ) );
  NOR2_X1 U1229 ( .A1(n339), .A2(n229), .ZN(\ab[44][51] ) );
  NOR2_X1 U1230 ( .A1(n341), .A2(n229), .ZN(\ab[44][50] ) );
  NOR2_X1 U1231 ( .A1(n439), .A2(n229), .ZN(\ab[44][4] ) );
  NOR2_X1 U1232 ( .A1(n344), .A2(n453), .ZN(\ab[44][49] ) );
  NOR2_X1 U1233 ( .A1(n346), .A2(n453), .ZN(\ab[44][48] ) );
  NOR2_X1 U1234 ( .A1(n348), .A2(n453), .ZN(\ab[44][47] ) );
  NOR2_X1 U1235 ( .A1(n350), .A2(n453), .ZN(\ab[44][46] ) );
  NOR2_X1 U1236 ( .A1(n352), .A2(n453), .ZN(\ab[44][45] ) );
  NOR2_X1 U1237 ( .A1(n354), .A2(n453), .ZN(\ab[44][44] ) );
  NOR2_X1 U1238 ( .A1(n357), .A2(n453), .ZN(\ab[44][43] ) );
  NOR2_X1 U1239 ( .A1(n359), .A2(n453), .ZN(\ab[44][42] ) );
  NOR2_X1 U1240 ( .A1(n362), .A2(n453), .ZN(\ab[44][41] ) );
  NOR2_X1 U1241 ( .A1(n364), .A2(n453), .ZN(\ab[44][40] ) );
  NOR2_X1 U1242 ( .A1(n478), .A2(n453), .ZN(\ab[44][3] ) );
  NOR2_X1 U1243 ( .A1(n366), .A2(n230), .ZN(\ab[44][39] ) );
  NOR2_X1 U1244 ( .A1(n367), .A2(n230), .ZN(\ab[44][38] ) );
  NOR2_X1 U1245 ( .A1(n371), .A2(n230), .ZN(\ab[44][37] ) );
  NOR2_X1 U1246 ( .A1(n372), .A2(n230), .ZN(\ab[44][36] ) );
  NOR2_X1 U1247 ( .A1(n374), .A2(n230), .ZN(\ab[44][35] ) );
  NOR2_X1 U1248 ( .A1(n376), .A2(n230), .ZN(\ab[44][34] ) );
  NOR2_X1 U1249 ( .A1(n378), .A2(n230), .ZN(\ab[44][33] ) );
  NOR2_X1 U1250 ( .A1(n379), .A2(n230), .ZN(\ab[44][32] ) );
  NOR2_X1 U1251 ( .A1(n382), .A2(n230), .ZN(\ab[44][31] ) );
  NOR2_X1 U1252 ( .A1(n384), .A2(n230), .ZN(\ab[44][30] ) );
  NOR2_X1 U1253 ( .A1(n479), .A2(n230), .ZN(\ab[44][2] ) );
  NOR2_X1 U1254 ( .A1(n385), .A2(n229), .ZN(\ab[44][29] ) );
  NOR2_X1 U1255 ( .A1(n388), .A2(n229), .ZN(\ab[44][28] ) );
  NOR2_X1 U1256 ( .A1(n389), .A2(n229), .ZN(\ab[44][27] ) );
  NOR2_X1 U1257 ( .A1(n391), .A2(n229), .ZN(\ab[44][26] ) );
  NOR2_X1 U1258 ( .A1(n394), .A2(n229), .ZN(\ab[44][25] ) );
  NOR2_X1 U1259 ( .A1(n396), .A2(n229), .ZN(\ab[44][24] ) );
  NOR2_X1 U1260 ( .A1(n398), .A2(n229), .ZN(\ab[44][23] ) );
  NOR2_X1 U1261 ( .A1(n399), .A2(n229), .ZN(\ab[44][22] ) );
  NOR2_X1 U1262 ( .A1(n401), .A2(n229), .ZN(\ab[44][21] ) );
  NOR2_X1 U1263 ( .A1(n403), .A2(n229), .ZN(\ab[44][20] ) );
  NOR2_X1 U1264 ( .A1(n444), .A2(n229), .ZN(\ab[44][1] ) );
  NOR2_X1 U1265 ( .A1(n405), .A2(n453), .ZN(\ab[44][19] ) );
  NOR2_X1 U1266 ( .A1(n407), .A2(n231), .ZN(\ab[44][18] ) );
  NOR2_X1 U1267 ( .A1(n408), .A2(n231), .ZN(\ab[44][17] ) );
  NOR2_X1 U1268 ( .A1(n411), .A2(n231), .ZN(\ab[44][16] ) );
  NOR2_X1 U1269 ( .A1(n414), .A2(n231), .ZN(\ab[44][15] ) );
  NOR2_X1 U1270 ( .A1(n417), .A2(n229), .ZN(\ab[44][14] ) );
  NOR2_X1 U1271 ( .A1(n420), .A2(n230), .ZN(\ab[44][13] ) );
  NOR2_X1 U1272 ( .A1(n423), .A2(n229), .ZN(\ab[44][12] ) );
  NOR2_X1 U1273 ( .A1(n425), .A2(n230), .ZN(\ab[44][11] ) );
  NOR2_X1 U1274 ( .A1(n477), .A2(n231), .ZN(\ab[44][10] ) );
  NOR2_X1 U1275 ( .A1(n480), .A2(n231), .ZN(\ab[44][0] ) );
  NOR2_X1 U1276 ( .A1(n429), .A2(n233), .ZN(\ab[43][9] ) );
  NOR2_X1 U1277 ( .A1(n431), .A2(n233), .ZN(\ab[43][8] ) );
  NOR2_X1 U1278 ( .A1(n433), .A2(n232), .ZN(\ab[43][7] ) );
  NOR2_X1 U1279 ( .A1(n435), .A2(n232), .ZN(\ab[43][6] ) );
  NOR2_X1 U1280 ( .A1(n437), .A2(n232), .ZN(\ab[43][5] ) );
  NOR2_X1 U1281 ( .A1(n337), .A2(n232), .ZN(\ab[43][52] ) );
  NOR2_X1 U1282 ( .A1(n339), .A2(n232), .ZN(\ab[43][51] ) );
  NOR2_X1 U1283 ( .A1(n341), .A2(n232), .ZN(\ab[43][50] ) );
  NOR2_X1 U1284 ( .A1(n439), .A2(n232), .ZN(\ab[43][4] ) );
  NOR2_X1 U1285 ( .A1(n344), .A2(n233), .ZN(\ab[43][49] ) );
  NOR2_X1 U1286 ( .A1(n345), .A2(n233), .ZN(\ab[43][48] ) );
  NOR2_X1 U1287 ( .A1(n347), .A2(n233), .ZN(\ab[43][47] ) );
  NOR2_X1 U1288 ( .A1(n349), .A2(n233), .ZN(\ab[43][46] ) );
  NOR2_X1 U1289 ( .A1(n351), .A2(n233), .ZN(\ab[43][45] ) );
  NOR2_X1 U1290 ( .A1(n354), .A2(n233), .ZN(\ab[43][44] ) );
  NOR2_X1 U1291 ( .A1(n357), .A2(n233), .ZN(\ab[43][43] ) );
  NOR2_X1 U1292 ( .A1(n359), .A2(n233), .ZN(\ab[43][42] ) );
  NOR2_X1 U1293 ( .A1(n361), .A2(n233), .ZN(\ab[43][41] ) );
  NOR2_X1 U1294 ( .A1(n363), .A2(n233), .ZN(\ab[43][40] ) );
  NOR2_X1 U1295 ( .A1(n441), .A2(n233), .ZN(\ab[43][3] ) );
  NOR2_X1 U1296 ( .A1(n365), .A2(n454), .ZN(\ab[43][39] ) );
  NOR2_X1 U1297 ( .A1(n367), .A2(n454), .ZN(\ab[43][38] ) );
  NOR2_X1 U1298 ( .A1(n371), .A2(n454), .ZN(\ab[43][37] ) );
  NOR2_X1 U1299 ( .A1(n474), .A2(n454), .ZN(\ab[43][36] ) );
  NOR2_X1 U1300 ( .A1(n373), .A2(n454), .ZN(\ab[43][35] ) );
  NOR2_X1 U1301 ( .A1(n375), .A2(n454), .ZN(\ab[43][34] ) );
  NOR2_X1 U1302 ( .A1(n377), .A2(n454), .ZN(\ab[43][33] ) );
  NOR2_X1 U1303 ( .A1(n380), .A2(n232), .ZN(\ab[43][32] ) );
  NOR2_X1 U1304 ( .A1(n381), .A2(n233), .ZN(\ab[43][31] ) );
  NOR2_X1 U1305 ( .A1(n383), .A2(n232), .ZN(\ab[43][30] ) );
  NOR2_X1 U1306 ( .A1(n479), .A2(n233), .ZN(\ab[43][2] ) );
  NOR2_X1 U1307 ( .A1(n386), .A2(n232), .ZN(\ab[43][29] ) );
  NOR2_X1 U1308 ( .A1(n388), .A2(n232), .ZN(\ab[43][28] ) );
  NOR2_X1 U1309 ( .A1(n390), .A2(n232), .ZN(\ab[43][27] ) );
  NOR2_X1 U1310 ( .A1(n392), .A2(n232), .ZN(\ab[43][26] ) );
  NOR2_X1 U1311 ( .A1(n393), .A2(n232), .ZN(\ab[43][25] ) );
  NOR2_X1 U1312 ( .A1(n395), .A2(n232), .ZN(\ab[43][24] ) );
  NOR2_X1 U1313 ( .A1(n397), .A2(n232), .ZN(\ab[43][23] ) );
  NOR2_X1 U1314 ( .A1(n400), .A2(n232), .ZN(\ab[43][22] ) );
  NOR2_X1 U1315 ( .A1(n402), .A2(n232), .ZN(\ab[43][21] ) );
  NOR2_X1 U1316 ( .A1(n475), .A2(n232), .ZN(\ab[43][20] ) );
  NOR2_X1 U1317 ( .A1(n444), .A2(n232), .ZN(\ab[43][1] ) );
  NOR2_X1 U1318 ( .A1(n405), .A2(n454), .ZN(\ab[43][19] ) );
  NOR2_X1 U1319 ( .A1(n407), .A2(n454), .ZN(\ab[43][18] ) );
  NOR2_X1 U1320 ( .A1(n409), .A2(n234), .ZN(\ab[43][17] ) );
  NOR2_X1 U1321 ( .A1(n411), .A2(n234), .ZN(\ab[43][16] ) );
  NOR2_X1 U1322 ( .A1(n414), .A2(n234), .ZN(\ab[43][15] ) );
  NOR2_X1 U1323 ( .A1(n417), .A2(n232), .ZN(\ab[43][14] ) );
  NOR2_X1 U1324 ( .A1(n420), .A2(n232), .ZN(\ab[43][13] ) );
  NOR2_X1 U1325 ( .A1(n423), .A2(n234), .ZN(\ab[43][12] ) );
  NOR2_X1 U1326 ( .A1(n426), .A2(n234), .ZN(\ab[43][11] ) );
  NOR2_X1 U1327 ( .A1(n427), .A2(n454), .ZN(\ab[43][10] ) );
  NOR2_X1 U1328 ( .A1(n446), .A2(n234), .ZN(\ab[43][0] ) );
  NOR2_X1 U1329 ( .A1(n429), .A2(n238), .ZN(\ab[42][9] ) );
  NOR2_X1 U1330 ( .A1(n431), .A2(n237), .ZN(\ab[42][8] ) );
  NOR2_X1 U1331 ( .A1(n433), .A2(n236), .ZN(\ab[42][7] ) );
  NOR2_X1 U1332 ( .A1(n435), .A2(n236), .ZN(\ab[42][6] ) );
  NOR2_X1 U1333 ( .A1(n437), .A2(n236), .ZN(\ab[42][5] ) );
  NOR2_X1 U1334 ( .A1(n337), .A2(n236), .ZN(\ab[42][52] ) );
  NOR2_X1 U1335 ( .A1(n339), .A2(n236), .ZN(\ab[42][51] ) );
  NOR2_X1 U1336 ( .A1(n341), .A2(n236), .ZN(\ab[42][50] ) );
  NOR2_X1 U1337 ( .A1(n439), .A2(n236), .ZN(\ab[42][4] ) );
  NOR2_X1 U1338 ( .A1(n344), .A2(n238), .ZN(\ab[42][49] ) );
  NOR2_X1 U1339 ( .A1(n346), .A2(n238), .ZN(\ab[42][48] ) );
  NOR2_X1 U1340 ( .A1(n348), .A2(n238), .ZN(\ab[42][47] ) );
  NOR2_X1 U1341 ( .A1(n350), .A2(n238), .ZN(\ab[42][46] ) );
  NOR2_X1 U1342 ( .A1(n352), .A2(n238), .ZN(\ab[42][45] ) );
  NOR2_X1 U1343 ( .A1(n354), .A2(n238), .ZN(\ab[42][44] ) );
  NOR2_X1 U1344 ( .A1(n357), .A2(n238), .ZN(\ab[42][43] ) );
  NOR2_X1 U1345 ( .A1(n359), .A2(n238), .ZN(\ab[42][42] ) );
  NOR2_X1 U1346 ( .A1(n362), .A2(n238), .ZN(\ab[42][41] ) );
  NOR2_X1 U1347 ( .A1(n364), .A2(n238), .ZN(\ab[42][40] ) );
  NOR2_X1 U1348 ( .A1(n478), .A2(n238), .ZN(\ab[42][3] ) );
  NOR2_X1 U1349 ( .A1(n366), .A2(n237), .ZN(\ab[42][39] ) );
  NOR2_X1 U1350 ( .A1(n367), .A2(n237), .ZN(\ab[42][38] ) );
  NOR2_X1 U1351 ( .A1(n371), .A2(n237), .ZN(\ab[42][37] ) );
  NOR2_X1 U1352 ( .A1(n372), .A2(n237), .ZN(\ab[42][36] ) );
  NOR2_X1 U1353 ( .A1(n374), .A2(n237), .ZN(\ab[42][35] ) );
  NOR2_X1 U1354 ( .A1(n376), .A2(n237), .ZN(\ab[42][34] ) );
  NOR2_X1 U1355 ( .A1(n378), .A2(n237), .ZN(\ab[42][33] ) );
  NOR2_X1 U1356 ( .A1(n379), .A2(n237), .ZN(\ab[42][32] ) );
  NOR2_X1 U1357 ( .A1(n382), .A2(n237), .ZN(\ab[42][31] ) );
  NOR2_X1 U1358 ( .A1(n384), .A2(n237), .ZN(\ab[42][30] ) );
  NOR2_X1 U1359 ( .A1(n479), .A2(n237), .ZN(\ab[42][2] ) );
  NOR2_X1 U1360 ( .A1(n385), .A2(n236), .ZN(\ab[42][29] ) );
  NOR2_X1 U1361 ( .A1(n388), .A2(n236), .ZN(\ab[42][28] ) );
  NOR2_X1 U1362 ( .A1(n389), .A2(n236), .ZN(\ab[42][27] ) );
  NOR2_X1 U1363 ( .A1(n391), .A2(n236), .ZN(\ab[42][26] ) );
  NOR2_X1 U1364 ( .A1(n394), .A2(n236), .ZN(\ab[42][25] ) );
  NOR2_X1 U1365 ( .A1(n396), .A2(n236), .ZN(\ab[42][24] ) );
  NOR2_X1 U1366 ( .A1(n398), .A2(n236), .ZN(\ab[42][23] ) );
  NOR2_X1 U1367 ( .A1(n399), .A2(n236), .ZN(\ab[42][22] ) );
  NOR2_X1 U1368 ( .A1(n401), .A2(n236), .ZN(\ab[42][21] ) );
  NOR2_X1 U1369 ( .A1(n403), .A2(n236), .ZN(\ab[42][20] ) );
  NOR2_X1 U1370 ( .A1(n444), .A2(n236), .ZN(\ab[42][1] ) );
  NOR2_X1 U1371 ( .A1(n405), .A2(n239), .ZN(\ab[42][19] ) );
  NOR2_X1 U1372 ( .A1(n407), .A2(n239), .ZN(\ab[42][18] ) );
  NOR2_X1 U1373 ( .A1(n408), .A2(n239), .ZN(\ab[42][17] ) );
  NOR2_X1 U1374 ( .A1(n411), .A2(n239), .ZN(\ab[42][16] ) );
  NOR2_X1 U1375 ( .A1(n414), .A2(n236), .ZN(\ab[42][15] ) );
  NOR2_X1 U1376 ( .A1(n417), .A2(n236), .ZN(\ab[42][14] ) );
  NOR2_X1 U1377 ( .A1(n420), .A2(n239), .ZN(\ab[42][13] ) );
  NOR2_X1 U1378 ( .A1(n423), .A2(n239), .ZN(\ab[42][12] ) );
  NOR2_X1 U1379 ( .A1(n425), .A2(n239), .ZN(\ab[42][11] ) );
  NOR2_X1 U1380 ( .A1(n477), .A2(n237), .ZN(\ab[42][10] ) );
  NOR2_X1 U1381 ( .A1(n480), .A2(n239), .ZN(\ab[42][0] ) );
  NOR2_X1 U1382 ( .A1(n429), .A2(n242), .ZN(\ab[41][9] ) );
  NOR2_X1 U1383 ( .A1(n431), .A2(n241), .ZN(\ab[41][8] ) );
  NOR2_X1 U1384 ( .A1(n433), .A2(n240), .ZN(\ab[41][7] ) );
  NOR2_X1 U1385 ( .A1(n435), .A2(n240), .ZN(\ab[41][6] ) );
  NOR2_X1 U1386 ( .A1(n437), .A2(n240), .ZN(\ab[41][5] ) );
  NOR2_X1 U1387 ( .A1(n337), .A2(n240), .ZN(\ab[41][52] ) );
  NOR2_X1 U1388 ( .A1(n339), .A2(n240), .ZN(\ab[41][51] ) );
  NOR2_X1 U1389 ( .A1(n341), .A2(n240), .ZN(\ab[41][50] ) );
  NOR2_X1 U1390 ( .A1(n439), .A2(n240), .ZN(\ab[41][4] ) );
  NOR2_X1 U1391 ( .A1(n344), .A2(n242), .ZN(\ab[41][49] ) );
  NOR2_X1 U1392 ( .A1(n345), .A2(n242), .ZN(\ab[41][48] ) );
  NOR2_X1 U1393 ( .A1(n347), .A2(n242), .ZN(\ab[41][47] ) );
  NOR2_X1 U1394 ( .A1(n349), .A2(n242), .ZN(\ab[41][46] ) );
  NOR2_X1 U1395 ( .A1(n351), .A2(n242), .ZN(\ab[41][45] ) );
  NOR2_X1 U1396 ( .A1(n354), .A2(n242), .ZN(\ab[41][44] ) );
  NOR2_X1 U1397 ( .A1(n357), .A2(n242), .ZN(\ab[41][43] ) );
  NOR2_X1 U1398 ( .A1(n359), .A2(n242), .ZN(\ab[41][42] ) );
  NOR2_X1 U1399 ( .A1(n361), .A2(n242), .ZN(\ab[41][41] ) );
  NOR2_X1 U1400 ( .A1(n363), .A2(n242), .ZN(\ab[41][40] ) );
  NOR2_X1 U1401 ( .A1(n478), .A2(n242), .ZN(\ab[41][3] ) );
  NOR2_X1 U1402 ( .A1(n365), .A2(n241), .ZN(\ab[41][39] ) );
  NOR2_X1 U1403 ( .A1(n367), .A2(n241), .ZN(\ab[41][38] ) );
  NOR2_X1 U1404 ( .A1(n371), .A2(n241), .ZN(\ab[41][37] ) );
  NOR2_X1 U1405 ( .A1(n474), .A2(n241), .ZN(\ab[41][36] ) );
  NOR2_X1 U1406 ( .A1(n373), .A2(n241), .ZN(\ab[41][35] ) );
  NOR2_X1 U1407 ( .A1(n375), .A2(n241), .ZN(\ab[41][34] ) );
  NOR2_X1 U1408 ( .A1(n377), .A2(n241), .ZN(\ab[41][33] ) );
  NOR2_X1 U1409 ( .A1(n380), .A2(n241), .ZN(\ab[41][32] ) );
  NOR2_X1 U1410 ( .A1(n381), .A2(n241), .ZN(\ab[41][31] ) );
  NOR2_X1 U1411 ( .A1(n383), .A2(n241), .ZN(\ab[41][30] ) );
  NOR2_X1 U1412 ( .A1(n479), .A2(n241), .ZN(\ab[41][2] ) );
  NOR2_X1 U1413 ( .A1(n386), .A2(n240), .ZN(\ab[41][29] ) );
  NOR2_X1 U1414 ( .A1(n388), .A2(n240), .ZN(\ab[41][28] ) );
  NOR2_X1 U1415 ( .A1(n390), .A2(n240), .ZN(\ab[41][27] ) );
  NOR2_X1 U1416 ( .A1(n392), .A2(n240), .ZN(\ab[41][26] ) );
  NOR2_X1 U1417 ( .A1(n393), .A2(n240), .ZN(\ab[41][25] ) );
  NOR2_X1 U1418 ( .A1(n395), .A2(n240), .ZN(\ab[41][24] ) );
  NOR2_X1 U1419 ( .A1(n397), .A2(n240), .ZN(\ab[41][23] ) );
  NOR2_X1 U1420 ( .A1(n400), .A2(n240), .ZN(\ab[41][22] ) );
  NOR2_X1 U1421 ( .A1(n402), .A2(n240), .ZN(\ab[41][21] ) );
  NOR2_X1 U1422 ( .A1(n475), .A2(n240), .ZN(\ab[41][20] ) );
  NOR2_X1 U1423 ( .A1(n444), .A2(n240), .ZN(\ab[41][1] ) );
  NOR2_X1 U1424 ( .A1(n405), .A2(n241), .ZN(\ab[41][19] ) );
  NOR2_X1 U1425 ( .A1(n407), .A2(n240), .ZN(\ab[41][18] ) );
  NOR2_X1 U1426 ( .A1(n409), .A2(n240), .ZN(\ab[41][17] ) );
  NOR2_X1 U1427 ( .A1(n411), .A2(n240), .ZN(\ab[41][16] ) );
  NOR2_X1 U1428 ( .A1(n414), .A2(n241), .ZN(\ab[41][15] ) );
  NOR2_X1 U1429 ( .A1(n417), .A2(n243), .ZN(\ab[41][14] ) );
  NOR2_X1 U1430 ( .A1(n420), .A2(n243), .ZN(\ab[41][13] ) );
  NOR2_X1 U1431 ( .A1(n423), .A2(n243), .ZN(\ab[41][12] ) );
  NOR2_X1 U1432 ( .A1(n426), .A2(n243), .ZN(\ab[41][11] ) );
  NOR2_X1 U1433 ( .A1(n427), .A2(n243), .ZN(\ab[41][10] ) );
  NOR2_X1 U1434 ( .A1(n446), .A2(n242), .ZN(\ab[41][0] ) );
  NOR2_X1 U1435 ( .A1(n429), .A2(n246), .ZN(\ab[40][9] ) );
  NOR2_X1 U1436 ( .A1(n431), .A2(n245), .ZN(\ab[40][8] ) );
  NOR2_X1 U1437 ( .A1(n433), .A2(n244), .ZN(\ab[40][7] ) );
  NOR2_X1 U1438 ( .A1(n435), .A2(n244), .ZN(\ab[40][6] ) );
  NOR2_X1 U1439 ( .A1(n437), .A2(n244), .ZN(\ab[40][5] ) );
  NOR2_X1 U1440 ( .A1(n337), .A2(n244), .ZN(\ab[40][52] ) );
  NOR2_X1 U1441 ( .A1(n339), .A2(n244), .ZN(\ab[40][51] ) );
  NOR2_X1 U1442 ( .A1(n341), .A2(n244), .ZN(\ab[40][50] ) );
  NOR2_X1 U1443 ( .A1(n439), .A2(n244), .ZN(\ab[40][4] ) );
  NOR2_X1 U1444 ( .A1(n344), .A2(n246), .ZN(\ab[40][49] ) );
  NOR2_X1 U1445 ( .A1(n346), .A2(n246), .ZN(\ab[40][48] ) );
  NOR2_X1 U1446 ( .A1(n348), .A2(n246), .ZN(\ab[40][47] ) );
  NOR2_X1 U1447 ( .A1(n350), .A2(n246), .ZN(\ab[40][46] ) );
  NOR2_X1 U1448 ( .A1(n352), .A2(n246), .ZN(\ab[40][45] ) );
  NOR2_X1 U1449 ( .A1(n354), .A2(n246), .ZN(\ab[40][44] ) );
  NOR2_X1 U1450 ( .A1(n357), .A2(n246), .ZN(\ab[40][43] ) );
  NOR2_X1 U1451 ( .A1(n359), .A2(n246), .ZN(\ab[40][42] ) );
  NOR2_X1 U1452 ( .A1(n362), .A2(n246), .ZN(\ab[40][41] ) );
  NOR2_X1 U1453 ( .A1(n364), .A2(n246), .ZN(\ab[40][40] ) );
  NOR2_X1 U1454 ( .A1(n478), .A2(n246), .ZN(\ab[40][3] ) );
  NOR2_X1 U1455 ( .A1(n366), .A2(n245), .ZN(\ab[40][39] ) );
  NOR2_X1 U1456 ( .A1(n367), .A2(n245), .ZN(\ab[40][38] ) );
  NOR2_X1 U1457 ( .A1(n371), .A2(n245), .ZN(\ab[40][37] ) );
  NOR2_X1 U1458 ( .A1(n372), .A2(n245), .ZN(\ab[40][36] ) );
  NOR2_X1 U1459 ( .A1(n374), .A2(n245), .ZN(\ab[40][35] ) );
  NOR2_X1 U1460 ( .A1(n376), .A2(n245), .ZN(\ab[40][34] ) );
  NOR2_X1 U1461 ( .A1(n378), .A2(n245), .ZN(\ab[40][33] ) );
  NOR2_X1 U1462 ( .A1(n379), .A2(n245), .ZN(\ab[40][32] ) );
  NOR2_X1 U1463 ( .A1(n382), .A2(n245), .ZN(\ab[40][31] ) );
  NOR2_X1 U1464 ( .A1(n384), .A2(n245), .ZN(\ab[40][30] ) );
  NOR2_X1 U1465 ( .A1(n479), .A2(n245), .ZN(\ab[40][2] ) );
  NOR2_X1 U1466 ( .A1(n385), .A2(n244), .ZN(\ab[40][29] ) );
  NOR2_X1 U1467 ( .A1(n388), .A2(n244), .ZN(\ab[40][28] ) );
  NOR2_X1 U1468 ( .A1(n389), .A2(n244), .ZN(\ab[40][27] ) );
  NOR2_X1 U1469 ( .A1(n391), .A2(n244), .ZN(\ab[40][26] ) );
  NOR2_X1 U1470 ( .A1(n394), .A2(n244), .ZN(\ab[40][25] ) );
  NOR2_X1 U1471 ( .A1(n396), .A2(n244), .ZN(\ab[40][24] ) );
  NOR2_X1 U1472 ( .A1(n398), .A2(n244), .ZN(\ab[40][23] ) );
  NOR2_X1 U1473 ( .A1(n399), .A2(n244), .ZN(\ab[40][22] ) );
  NOR2_X1 U1474 ( .A1(n401), .A2(n244), .ZN(\ab[40][21] ) );
  NOR2_X1 U1475 ( .A1(n403), .A2(n244), .ZN(\ab[40][20] ) );
  NOR2_X1 U1476 ( .A1(n444), .A2(n244), .ZN(\ab[40][1] ) );
  NOR2_X1 U1477 ( .A1(n405), .A2(n244), .ZN(\ab[40][19] ) );
  NOR2_X1 U1478 ( .A1(n407), .A2(n244), .ZN(\ab[40][18] ) );
  NOR2_X1 U1479 ( .A1(n408), .A2(n244), .ZN(\ab[40][17] ) );
  NOR2_X1 U1480 ( .A1(n411), .A2(n245), .ZN(\ab[40][16] ) );
  NOR2_X1 U1481 ( .A1(n414), .A2(n246), .ZN(\ab[40][15] ) );
  NOR2_X1 U1482 ( .A1(n417), .A2(n246), .ZN(\ab[40][14] ) );
  NOR2_X1 U1483 ( .A1(n420), .A2(n245), .ZN(\ab[40][13] ) );
  NOR2_X1 U1484 ( .A1(n423), .A2(n245), .ZN(\ab[40][12] ) );
  NOR2_X1 U1485 ( .A1(n425), .A2(n246), .ZN(\ab[40][11] ) );
  NOR2_X1 U1486 ( .A1(n477), .A2(n245), .ZN(\ab[40][10] ) );
  NOR2_X1 U1487 ( .A1(n480), .A2(n244), .ZN(\ab[40][0] ) );
  NOR2_X1 U1488 ( .A1(n429), .A2(n325), .ZN(\ab[3][9] ) );
  NOR2_X1 U1489 ( .A1(n431), .A2(n325), .ZN(\ab[3][8] ) );
  NOR2_X1 U1490 ( .A1(n433), .A2(n325), .ZN(\ab[3][7] ) );
  NOR2_X1 U1491 ( .A1(n435), .A2(n325), .ZN(\ab[3][6] ) );
  NOR2_X1 U1492 ( .A1(n437), .A2(n325), .ZN(\ab[3][5] ) );
  NOR2_X1 U1493 ( .A1(n337), .A2(n326), .ZN(\ab[3][52] ) );
  NOR2_X1 U1494 ( .A1(n339), .A2(n326), .ZN(\ab[3][51] ) );
  NOR2_X1 U1495 ( .A1(n341), .A2(n326), .ZN(\ab[3][50] ) );
  NOR2_X1 U1496 ( .A1(n439), .A2(n325), .ZN(\ab[3][4] ) );
  NOR2_X1 U1497 ( .A1(n344), .A2(n326), .ZN(\ab[3][49] ) );
  NOR2_X1 U1498 ( .A1(n346), .A2(n326), .ZN(\ab[3][48] ) );
  NOR2_X1 U1499 ( .A1(n348), .A2(n326), .ZN(\ab[3][47] ) );
  NOR2_X1 U1500 ( .A1(n350), .A2(n326), .ZN(\ab[3][46] ) );
  NOR2_X1 U1501 ( .A1(n352), .A2(n325), .ZN(\ab[3][45] ) );
  NOR2_X1 U1502 ( .A1(n354), .A2(n325), .ZN(\ab[3][44] ) );
  NOR2_X1 U1503 ( .A1(n357), .A2(n325), .ZN(\ab[3][43] ) );
  NOR2_X1 U1504 ( .A1(n359), .A2(n325), .ZN(\ab[3][42] ) );
  NOR2_X1 U1505 ( .A1(n362), .A2(n325), .ZN(\ab[3][41] ) );
  NOR2_X1 U1506 ( .A1(n364), .A2(n326), .ZN(\ab[3][40] ) );
  NOR2_X1 U1507 ( .A1(n441), .A2(n325), .ZN(\ab[3][3] ) );
  NOR2_X1 U1508 ( .A1(n366), .A2(n326), .ZN(\ab[3][39] ) );
  NOR2_X1 U1509 ( .A1(n367), .A2(n326), .ZN(\ab[3][38] ) );
  NOR2_X1 U1510 ( .A1(n371), .A2(n326), .ZN(\ab[3][37] ) );
  NOR2_X1 U1511 ( .A1(n474), .A2(n326), .ZN(\ab[3][36] ) );
  NOR2_X1 U1512 ( .A1(n374), .A2(n326), .ZN(\ab[3][35] ) );
  NOR2_X1 U1513 ( .A1(n376), .A2(n326), .ZN(\ab[3][34] ) );
  NOR2_X1 U1514 ( .A1(n378), .A2(n326), .ZN(\ab[3][33] ) );
  NOR2_X1 U1515 ( .A1(n380), .A2(n326), .ZN(\ab[3][32] ) );
  NOR2_X1 U1516 ( .A1(n382), .A2(n326), .ZN(\ab[3][31] ) );
  NOR2_X1 U1517 ( .A1(n384), .A2(n326), .ZN(\ab[3][30] ) );
  NOR2_X1 U1518 ( .A1(n442), .A2(n326), .ZN(\ab[3][2] ) );
  NOR2_X1 U1519 ( .A1(n386), .A2(n325), .ZN(\ab[3][29] ) );
  NOR2_X1 U1520 ( .A1(n388), .A2(n325), .ZN(\ab[3][28] ) );
  NOR2_X1 U1521 ( .A1(n390), .A2(n325), .ZN(\ab[3][27] ) );
  NOR2_X1 U1522 ( .A1(n392), .A2(n325), .ZN(\ab[3][26] ) );
  NOR2_X1 U1523 ( .A1(n394), .A2(n325), .ZN(\ab[3][25] ) );
  NOR2_X1 U1524 ( .A1(n396), .A2(n325), .ZN(\ab[3][24] ) );
  NOR2_X1 U1525 ( .A1(n398), .A2(n325), .ZN(\ab[3][23] ) );
  NOR2_X1 U1526 ( .A1(n400), .A2(n325), .ZN(\ab[3][22] ) );
  NOR2_X1 U1527 ( .A1(n402), .A2(n325), .ZN(\ab[3][21] ) );
  NOR2_X1 U1528 ( .A1(n475), .A2(n325), .ZN(\ab[3][20] ) );
  NOR2_X1 U1529 ( .A1(n444), .A2(n325), .ZN(\ab[3][1] ) );
  NOR2_X1 U1530 ( .A1(n405), .A2(n325), .ZN(\ab[3][19] ) );
  NOR2_X1 U1531 ( .A1(n407), .A2(n325), .ZN(\ab[3][18] ) );
  NOR2_X1 U1532 ( .A1(n409), .A2(n325), .ZN(\ab[3][17] ) );
  NOR2_X1 U1533 ( .A1(n411), .A2(n325), .ZN(\ab[3][16] ) );
  NOR2_X1 U1534 ( .A1(n414), .A2(n325), .ZN(\ab[3][15] ) );
  NOR2_X1 U1535 ( .A1(n417), .A2(n325), .ZN(\ab[3][14] ) );
  NOR2_X1 U1536 ( .A1(n420), .A2(n325), .ZN(\ab[3][13] ) );
  NOR2_X1 U1537 ( .A1(n423), .A2(n325), .ZN(\ab[3][12] ) );
  NOR2_X1 U1538 ( .A1(n426), .A2(n325), .ZN(\ab[3][11] ) );
  NOR2_X1 U1539 ( .A1(n477), .A2(n325), .ZN(\ab[3][10] ) );
  NOR2_X1 U1540 ( .A1(n480), .A2(n325), .ZN(\ab[3][0] ) );
  NOR2_X1 U1541 ( .A1(n428), .A2(n248), .ZN(\ab[39][9] ) );
  NOR2_X1 U1542 ( .A1(n430), .A2(n248), .ZN(\ab[39][8] ) );
  NOR2_X1 U1543 ( .A1(n432), .A2(n248), .ZN(\ab[39][7] ) );
  NOR2_X1 U1544 ( .A1(n435), .A2(n248), .ZN(\ab[39][6] ) );
  NOR2_X1 U1545 ( .A1(n437), .A2(n248), .ZN(\ab[39][5] ) );
  NOR2_X1 U1546 ( .A1(n337), .A2(n248), .ZN(\ab[39][52] ) );
  NOR2_X1 U1547 ( .A1(n338), .A2(n248), .ZN(\ab[39][51] ) );
  NOR2_X1 U1548 ( .A1(n342), .A2(n248), .ZN(\ab[39][50] ) );
  NOR2_X1 U1549 ( .A1(n439), .A2(n248), .ZN(\ab[39][4] ) );
  NOR2_X1 U1550 ( .A1(n343), .A2(n247), .ZN(\ab[39][49] ) );
  NOR2_X1 U1551 ( .A1(n345), .A2(n248), .ZN(\ab[39][48] ) );
  NOR2_X1 U1552 ( .A1(n347), .A2(n248), .ZN(\ab[39][47] ) );
  NOR2_X1 U1553 ( .A1(n349), .A2(n248), .ZN(\ab[39][46] ) );
  NOR2_X1 U1554 ( .A1(n351), .A2(n247), .ZN(\ab[39][45] ) );
  NOR2_X1 U1555 ( .A1(n353), .A2(n248), .ZN(\ab[39][44] ) );
  NOR2_X1 U1556 ( .A1(n356), .A2(n248), .ZN(\ab[39][43] ) );
  NOR2_X1 U1557 ( .A1(n358), .A2(n248), .ZN(\ab[39][42] ) );
  NOR2_X1 U1558 ( .A1(n361), .A2(n247), .ZN(\ab[39][41] ) );
  NOR2_X1 U1559 ( .A1(n363), .A2(n247), .ZN(\ab[39][40] ) );
  NOR2_X1 U1560 ( .A1(n478), .A2(n247), .ZN(\ab[39][3] ) );
  NOR2_X1 U1561 ( .A1(n365), .A2(n247), .ZN(\ab[39][39] ) );
  NOR2_X1 U1562 ( .A1(n369), .A2(n247), .ZN(\ab[39][38] ) );
  NOR2_X1 U1563 ( .A1(n370), .A2(n247), .ZN(\ab[39][37] ) );
  NOR2_X1 U1564 ( .A1(n372), .A2(n247), .ZN(\ab[39][36] ) );
  NOR2_X1 U1565 ( .A1(n373), .A2(n247), .ZN(\ab[39][35] ) );
  NOR2_X1 U1566 ( .A1(n375), .A2(n247), .ZN(\ab[39][34] ) );
  NOR2_X1 U1567 ( .A1(n377), .A2(n247), .ZN(\ab[39][33] ) );
  NOR2_X1 U1568 ( .A1(n379), .A2(n247), .ZN(\ab[39][32] ) );
  NOR2_X1 U1569 ( .A1(n381), .A2(n247), .ZN(\ab[39][31] ) );
  NOR2_X1 U1570 ( .A1(n383), .A2(n247), .ZN(\ab[39][30] ) );
  NOR2_X1 U1571 ( .A1(n479), .A2(n247), .ZN(\ab[39][2] ) );
  NOR2_X1 U1572 ( .A1(n385), .A2(n247), .ZN(\ab[39][29] ) );
  NOR2_X1 U1573 ( .A1(n387), .A2(n247), .ZN(\ab[39][28] ) );
  NOR2_X1 U1574 ( .A1(n389), .A2(n247), .ZN(\ab[39][27] ) );
  NOR2_X1 U1575 ( .A1(n391), .A2(n247), .ZN(\ab[39][26] ) );
  NOR2_X1 U1576 ( .A1(n393), .A2(n247), .ZN(\ab[39][25] ) );
  NOR2_X1 U1577 ( .A1(n395), .A2(n247), .ZN(\ab[39][24] ) );
  NOR2_X1 U1578 ( .A1(n397), .A2(n247), .ZN(\ab[39][23] ) );
  NOR2_X1 U1579 ( .A1(n399), .A2(n247), .ZN(\ab[39][22] ) );
  NOR2_X1 U1580 ( .A1(n401), .A2(n247), .ZN(\ab[39][21] ) );
  NOR2_X1 U1581 ( .A1(n403), .A2(n247), .ZN(\ab[39][20] ) );
  NOR2_X1 U1582 ( .A1(n444), .A2(n247), .ZN(\ab[39][1] ) );
  NOR2_X1 U1583 ( .A1(n404), .A2(n247), .ZN(\ab[39][19] ) );
  NOR2_X1 U1584 ( .A1(n406), .A2(n247), .ZN(\ab[39][18] ) );
  NOR2_X1 U1585 ( .A1(n408), .A2(n248), .ZN(\ab[39][17] ) );
  NOR2_X1 U1586 ( .A1(n410), .A2(n455), .ZN(\ab[39][16] ) );
  NOR2_X1 U1587 ( .A1(n413), .A2(n455), .ZN(\ab[39][15] ) );
  NOR2_X1 U1588 ( .A1(n416), .A2(n455), .ZN(\ab[39][14] ) );
  NOR2_X1 U1589 ( .A1(n419), .A2(n455), .ZN(\ab[39][13] ) );
  NOR2_X1 U1590 ( .A1(n422), .A2(n455), .ZN(\ab[39][12] ) );
  NOR2_X1 U1591 ( .A1(n425), .A2(n455), .ZN(\ab[39][11] ) );
  NOR2_X1 U1592 ( .A1(n427), .A2(n248), .ZN(\ab[39][10] ) );
  NOR2_X1 U1593 ( .A1(n446), .A2(n247), .ZN(\ab[39][0] ) );
  NOR2_X1 U1594 ( .A1(n428), .A2(n251), .ZN(\ab[38][9] ) );
  NOR2_X1 U1595 ( .A1(n430), .A2(n249), .ZN(\ab[38][8] ) );
  NOR2_X1 U1596 ( .A1(n432), .A2(n250), .ZN(\ab[38][7] ) );
  NOR2_X1 U1597 ( .A1(n435), .A2(n250), .ZN(\ab[38][6] ) );
  NOR2_X1 U1598 ( .A1(n437), .A2(n250), .ZN(\ab[38][5] ) );
  NOR2_X1 U1599 ( .A1(n337), .A2(n250), .ZN(\ab[38][52] ) );
  NOR2_X1 U1600 ( .A1(n338), .A2(n250), .ZN(\ab[38][51] ) );
  NOR2_X1 U1601 ( .A1(n342), .A2(n250), .ZN(\ab[38][50] ) );
  NOR2_X1 U1602 ( .A1(n439), .A2(n250), .ZN(\ab[38][4] ) );
  NOR2_X1 U1603 ( .A1(n343), .A2(n251), .ZN(\ab[38][49] ) );
  NOR2_X1 U1604 ( .A1(n345), .A2(n251), .ZN(\ab[38][48] ) );
  NOR2_X1 U1605 ( .A1(n347), .A2(n251), .ZN(\ab[38][47] ) );
  NOR2_X1 U1606 ( .A1(n349), .A2(n251), .ZN(\ab[38][46] ) );
  NOR2_X1 U1607 ( .A1(n351), .A2(n251), .ZN(\ab[38][45] ) );
  NOR2_X1 U1608 ( .A1(n353), .A2(n251), .ZN(\ab[38][44] ) );
  NOR2_X1 U1609 ( .A1(n356), .A2(n251), .ZN(\ab[38][43] ) );
  NOR2_X1 U1610 ( .A1(n358), .A2(n251), .ZN(\ab[38][42] ) );
  NOR2_X1 U1611 ( .A1(n361), .A2(n251), .ZN(\ab[38][41] ) );
  NOR2_X1 U1612 ( .A1(n363), .A2(n251), .ZN(\ab[38][40] ) );
  NOR2_X1 U1613 ( .A1(n478), .A2(n251), .ZN(\ab[38][3] ) );
  NOR2_X1 U1614 ( .A1(n365), .A2(n250), .ZN(\ab[38][39] ) );
  NOR2_X1 U1615 ( .A1(n369), .A2(n250), .ZN(\ab[38][38] ) );
  NOR2_X1 U1616 ( .A1(n370), .A2(n250), .ZN(\ab[38][37] ) );
  NOR2_X1 U1617 ( .A1(n372), .A2(n250), .ZN(\ab[38][36] ) );
  NOR2_X1 U1618 ( .A1(n373), .A2(n250), .ZN(\ab[38][35] ) );
  NOR2_X1 U1619 ( .A1(n375), .A2(n250), .ZN(\ab[38][34] ) );
  NOR2_X1 U1620 ( .A1(n377), .A2(n250), .ZN(\ab[38][33] ) );
  NOR2_X1 U1621 ( .A1(n379), .A2(n250), .ZN(\ab[38][32] ) );
  NOR2_X1 U1622 ( .A1(n381), .A2(n250), .ZN(\ab[38][31] ) );
  NOR2_X1 U1623 ( .A1(n383), .A2(n250), .ZN(\ab[38][30] ) );
  NOR2_X1 U1624 ( .A1(n479), .A2(n250), .ZN(\ab[38][2] ) );
  NOR2_X1 U1625 ( .A1(n385), .A2(n249), .ZN(\ab[38][29] ) );
  NOR2_X1 U1626 ( .A1(n387), .A2(n249), .ZN(\ab[38][28] ) );
  NOR2_X1 U1627 ( .A1(n389), .A2(n249), .ZN(\ab[38][27] ) );
  NOR2_X1 U1628 ( .A1(n391), .A2(n249), .ZN(\ab[38][26] ) );
  NOR2_X1 U1629 ( .A1(n393), .A2(n249), .ZN(\ab[38][25] ) );
  NOR2_X1 U1630 ( .A1(n395), .A2(n249), .ZN(\ab[38][24] ) );
  NOR2_X1 U1631 ( .A1(n397), .A2(n249), .ZN(\ab[38][23] ) );
  NOR2_X1 U1632 ( .A1(n399), .A2(n249), .ZN(\ab[38][22] ) );
  NOR2_X1 U1633 ( .A1(n401), .A2(n249), .ZN(\ab[38][21] ) );
  NOR2_X1 U1634 ( .A1(n403), .A2(n249), .ZN(\ab[38][20] ) );
  NOR2_X1 U1635 ( .A1(n444), .A2(n249), .ZN(\ab[38][1] ) );
  NOR2_X1 U1636 ( .A1(n405), .A2(n250), .ZN(\ab[38][19] ) );
  NOR2_X1 U1637 ( .A1(n406), .A2(n249), .ZN(\ab[38][18] ) );
  NOR2_X1 U1638 ( .A1(n408), .A2(n252), .ZN(\ab[38][17] ) );
  NOR2_X1 U1639 ( .A1(n410), .A2(n252), .ZN(\ab[38][16] ) );
  NOR2_X1 U1640 ( .A1(n413), .A2(n252), .ZN(\ab[38][15] ) );
  NOR2_X1 U1641 ( .A1(n416), .A2(n252), .ZN(\ab[38][14] ) );
  NOR2_X1 U1642 ( .A1(n419), .A2(n252), .ZN(\ab[38][13] ) );
  NOR2_X1 U1643 ( .A1(n422), .A2(n249), .ZN(\ab[38][12] ) );
  NOR2_X1 U1644 ( .A1(n425), .A2(n251), .ZN(\ab[38][11] ) );
  NOR2_X1 U1645 ( .A1(n427), .A2(n250), .ZN(\ab[38][10] ) );
  NOR2_X1 U1646 ( .A1(n446), .A2(n250), .ZN(\ab[38][0] ) );
  NOR2_X1 U1647 ( .A1(n428), .A2(n253), .ZN(\ab[37][9] ) );
  NOR2_X1 U1648 ( .A1(n430), .A2(n255), .ZN(\ab[37][8] ) );
  NOR2_X1 U1649 ( .A1(n432), .A2(n254), .ZN(\ab[37][7] ) );
  NOR2_X1 U1650 ( .A1(n435), .A2(n254), .ZN(\ab[37][6] ) );
  NOR2_X1 U1651 ( .A1(n437), .A2(n254), .ZN(\ab[37][5] ) );
  NOR2_X1 U1652 ( .A1(n337), .A2(n254), .ZN(\ab[37][52] ) );
  NOR2_X1 U1653 ( .A1(n338), .A2(n254), .ZN(\ab[37][51] ) );
  NOR2_X1 U1654 ( .A1(n342), .A2(n254), .ZN(\ab[37][50] ) );
  NOR2_X1 U1655 ( .A1(n439), .A2(n254), .ZN(\ab[37][4] ) );
  NOR2_X1 U1656 ( .A1(n343), .A2(n255), .ZN(\ab[37][49] ) );
  NOR2_X1 U1657 ( .A1(n345), .A2(n255), .ZN(\ab[37][48] ) );
  NOR2_X1 U1658 ( .A1(n347), .A2(n255), .ZN(\ab[37][47] ) );
  NOR2_X1 U1659 ( .A1(n349), .A2(n255), .ZN(\ab[37][46] ) );
  NOR2_X1 U1660 ( .A1(n351), .A2(n255), .ZN(\ab[37][45] ) );
  NOR2_X1 U1661 ( .A1(n353), .A2(n255), .ZN(\ab[37][44] ) );
  NOR2_X1 U1662 ( .A1(n356), .A2(n255), .ZN(\ab[37][43] ) );
  NOR2_X1 U1663 ( .A1(n358), .A2(n255), .ZN(\ab[37][42] ) );
  NOR2_X1 U1664 ( .A1(n361), .A2(n255), .ZN(\ab[37][41] ) );
  NOR2_X1 U1665 ( .A1(n363), .A2(n255), .ZN(\ab[37][40] ) );
  NOR2_X1 U1666 ( .A1(n478), .A2(n255), .ZN(\ab[37][3] ) );
  NOR2_X1 U1667 ( .A1(n365), .A2(n254), .ZN(\ab[37][39] ) );
  NOR2_X1 U1668 ( .A1(n368), .A2(n254), .ZN(\ab[37][38] ) );
  NOR2_X1 U1669 ( .A1(n370), .A2(n254), .ZN(\ab[37][37] ) );
  NOR2_X1 U1670 ( .A1(n372), .A2(n254), .ZN(\ab[37][36] ) );
  NOR2_X1 U1671 ( .A1(n373), .A2(n254), .ZN(\ab[37][35] ) );
  NOR2_X1 U1672 ( .A1(n375), .A2(n254), .ZN(\ab[37][34] ) );
  NOR2_X1 U1673 ( .A1(n377), .A2(n254), .ZN(\ab[37][33] ) );
  NOR2_X1 U1674 ( .A1(n379), .A2(n254), .ZN(\ab[37][32] ) );
  NOR2_X1 U1675 ( .A1(n381), .A2(n254), .ZN(\ab[37][31] ) );
  NOR2_X1 U1676 ( .A1(n383), .A2(n254), .ZN(\ab[37][30] ) );
  NOR2_X1 U1677 ( .A1(n479), .A2(n254), .ZN(\ab[37][2] ) );
  NOR2_X1 U1678 ( .A1(n385), .A2(n253), .ZN(\ab[37][29] ) );
  NOR2_X1 U1679 ( .A1(n387), .A2(n253), .ZN(\ab[37][28] ) );
  NOR2_X1 U1680 ( .A1(n389), .A2(n253), .ZN(\ab[37][27] ) );
  NOR2_X1 U1681 ( .A1(n391), .A2(n253), .ZN(\ab[37][26] ) );
  NOR2_X1 U1682 ( .A1(n393), .A2(n253), .ZN(\ab[37][25] ) );
  NOR2_X1 U1683 ( .A1(n395), .A2(n253), .ZN(\ab[37][24] ) );
  NOR2_X1 U1684 ( .A1(n397), .A2(n253), .ZN(\ab[37][23] ) );
  NOR2_X1 U1685 ( .A1(n399), .A2(n253), .ZN(\ab[37][22] ) );
  NOR2_X1 U1686 ( .A1(n401), .A2(n253), .ZN(\ab[37][21] ) );
  NOR2_X1 U1687 ( .A1(n403), .A2(n253), .ZN(\ab[37][20] ) );
  NOR2_X1 U1688 ( .A1(n444), .A2(n253), .ZN(\ab[37][1] ) );
  NOR2_X1 U1689 ( .A1(n404), .A2(n253), .ZN(\ab[37][19] ) );
  NOR2_X1 U1690 ( .A1(n406), .A2(n253), .ZN(\ab[37][18] ) );
  NOR2_X1 U1691 ( .A1(n408), .A2(n255), .ZN(\ab[37][17] ) );
  NOR2_X1 U1692 ( .A1(n410), .A2(n253), .ZN(\ab[37][16] ) );
  NOR2_X1 U1693 ( .A1(n413), .A2(n255), .ZN(\ab[37][15] ) );
  NOR2_X1 U1694 ( .A1(n416), .A2(n253), .ZN(\ab[37][14] ) );
  NOR2_X1 U1695 ( .A1(n419), .A2(n255), .ZN(\ab[37][13] ) );
  NOR2_X1 U1696 ( .A1(n422), .A2(n254), .ZN(\ab[37][12] ) );
  NOR2_X1 U1697 ( .A1(n425), .A2(n254), .ZN(\ab[37][11] ) );
  NOR2_X1 U1698 ( .A1(n427), .A2(n254), .ZN(\ab[37][10] ) );
  NOR2_X1 U1699 ( .A1(n446), .A2(n255), .ZN(\ab[37][0] ) );
  NOR2_X1 U1700 ( .A1(n428), .A2(n257), .ZN(\ab[36][9] ) );
  NOR2_X1 U1701 ( .A1(n430), .A2(n256), .ZN(\ab[36][8] ) );
  NOR2_X1 U1702 ( .A1(n432), .A2(n256), .ZN(\ab[36][7] ) );
  NOR2_X1 U1703 ( .A1(n435), .A2(n256), .ZN(\ab[36][6] ) );
  NOR2_X1 U1704 ( .A1(n437), .A2(n256), .ZN(\ab[36][5] ) );
  NOR2_X1 U1705 ( .A1(n337), .A2(n256), .ZN(\ab[36][52] ) );
  NOR2_X1 U1706 ( .A1(n338), .A2(n256), .ZN(\ab[36][51] ) );
  NOR2_X1 U1707 ( .A1(n342), .A2(n256), .ZN(\ab[36][50] ) );
  NOR2_X1 U1708 ( .A1(n439), .A2(n256), .ZN(\ab[36][4] ) );
  NOR2_X1 U1709 ( .A1(n343), .A2(n257), .ZN(\ab[36][49] ) );
  NOR2_X1 U1710 ( .A1(n345), .A2(n257), .ZN(\ab[36][48] ) );
  NOR2_X1 U1711 ( .A1(n347), .A2(n257), .ZN(\ab[36][47] ) );
  NOR2_X1 U1712 ( .A1(n349), .A2(n257), .ZN(\ab[36][46] ) );
  NOR2_X1 U1713 ( .A1(n351), .A2(n257), .ZN(\ab[36][45] ) );
  NOR2_X1 U1714 ( .A1(n353), .A2(n257), .ZN(\ab[36][44] ) );
  NOR2_X1 U1715 ( .A1(n356), .A2(n257), .ZN(\ab[36][43] ) );
  NOR2_X1 U1716 ( .A1(n358), .A2(n257), .ZN(\ab[36][42] ) );
  NOR2_X1 U1717 ( .A1(n361), .A2(n257), .ZN(\ab[36][41] ) );
  NOR2_X1 U1718 ( .A1(n363), .A2(n257), .ZN(\ab[36][40] ) );
  NOR2_X1 U1719 ( .A1(n441), .A2(n257), .ZN(\ab[36][3] ) );
  NOR2_X1 U1720 ( .A1(n365), .A2(n256), .ZN(\ab[36][39] ) );
  NOR2_X1 U1721 ( .A1(n367), .A2(n256), .ZN(\ab[36][38] ) );
  NOR2_X1 U1722 ( .A1(n370), .A2(n256), .ZN(\ab[36][37] ) );
  NOR2_X1 U1723 ( .A1(n372), .A2(n256), .ZN(\ab[36][36] ) );
  NOR2_X1 U1724 ( .A1(n373), .A2(n256), .ZN(\ab[36][35] ) );
  NOR2_X1 U1725 ( .A1(n375), .A2(n256), .ZN(\ab[36][34] ) );
  NOR2_X1 U1726 ( .A1(n377), .A2(n256), .ZN(\ab[36][33] ) );
  NOR2_X1 U1727 ( .A1(n379), .A2(n256), .ZN(\ab[36][32] ) );
  NOR2_X1 U1728 ( .A1(n381), .A2(n256), .ZN(\ab[36][31] ) );
  NOR2_X1 U1729 ( .A1(n383), .A2(n256), .ZN(\ab[36][30] ) );
  NOR2_X1 U1730 ( .A1(n479), .A2(n256), .ZN(\ab[36][2] ) );
  NOR2_X1 U1731 ( .A1(n385), .A2(n258), .ZN(\ab[36][29] ) );
  NOR2_X1 U1732 ( .A1(n387), .A2(n258), .ZN(\ab[36][28] ) );
  NOR2_X1 U1733 ( .A1(n389), .A2(n258), .ZN(\ab[36][27] ) );
  NOR2_X1 U1734 ( .A1(n391), .A2(n258), .ZN(\ab[36][26] ) );
  NOR2_X1 U1735 ( .A1(n393), .A2(n258), .ZN(\ab[36][25] ) );
  NOR2_X1 U1736 ( .A1(n395), .A2(n258), .ZN(\ab[36][24] ) );
  NOR2_X1 U1737 ( .A1(n397), .A2(n258), .ZN(\ab[36][23] ) );
  NOR2_X1 U1738 ( .A1(n399), .A2(n258), .ZN(\ab[36][22] ) );
  NOR2_X1 U1739 ( .A1(n401), .A2(n258), .ZN(\ab[36][21] ) );
  NOR2_X1 U1740 ( .A1(n403), .A2(n257), .ZN(\ab[36][20] ) );
  NOR2_X1 U1741 ( .A1(n444), .A2(n258), .ZN(\ab[36][1] ) );
  NOR2_X1 U1742 ( .A1(n405), .A2(n258), .ZN(\ab[36][19] ) );
  NOR2_X1 U1743 ( .A1(n406), .A2(n258), .ZN(\ab[36][18] ) );
  NOR2_X1 U1744 ( .A1(n408), .A2(n258), .ZN(\ab[36][17] ) );
  NOR2_X1 U1745 ( .A1(n410), .A2(n258), .ZN(\ab[36][16] ) );
  NOR2_X1 U1746 ( .A1(n413), .A2(n257), .ZN(\ab[36][15] ) );
  NOR2_X1 U1747 ( .A1(n416), .A2(n257), .ZN(\ab[36][14] ) );
  NOR2_X1 U1748 ( .A1(n419), .A2(n257), .ZN(\ab[36][13] ) );
  NOR2_X1 U1749 ( .A1(n422), .A2(n256), .ZN(\ab[36][12] ) );
  NOR2_X1 U1750 ( .A1(n425), .A2(n256), .ZN(\ab[36][11] ) );
  NOR2_X1 U1751 ( .A1(n427), .A2(n256), .ZN(\ab[36][10] ) );
  NOR2_X1 U1752 ( .A1(n446), .A2(n258), .ZN(\ab[36][0] ) );
  NOR2_X1 U1753 ( .A1(n428), .A2(n260), .ZN(\ab[35][9] ) );
  NOR2_X1 U1754 ( .A1(n430), .A2(n259), .ZN(\ab[35][8] ) );
  NOR2_X1 U1755 ( .A1(n432), .A2(n259), .ZN(\ab[35][7] ) );
  NOR2_X1 U1756 ( .A1(n435), .A2(n259), .ZN(\ab[35][6] ) );
  NOR2_X1 U1757 ( .A1(n437), .A2(n259), .ZN(\ab[35][5] ) );
  NOR2_X1 U1758 ( .A1(n337), .A2(n259), .ZN(\ab[35][52] ) );
  NOR2_X1 U1759 ( .A1(n338), .A2(n259), .ZN(\ab[35][51] ) );
  NOR2_X1 U1760 ( .A1(n341), .A2(n259), .ZN(\ab[35][50] ) );
  NOR2_X1 U1761 ( .A1(n439), .A2(n259), .ZN(\ab[35][4] ) );
  NOR2_X1 U1762 ( .A1(n343), .A2(n260), .ZN(\ab[35][49] ) );
  NOR2_X1 U1763 ( .A1(n345), .A2(n260), .ZN(\ab[35][48] ) );
  NOR2_X1 U1764 ( .A1(n347), .A2(n260), .ZN(\ab[35][47] ) );
  NOR2_X1 U1765 ( .A1(n349), .A2(n260), .ZN(\ab[35][46] ) );
  NOR2_X1 U1766 ( .A1(n351), .A2(n260), .ZN(\ab[35][45] ) );
  NOR2_X1 U1767 ( .A1(n353), .A2(n260), .ZN(\ab[35][44] ) );
  NOR2_X1 U1768 ( .A1(n356), .A2(n260), .ZN(\ab[35][43] ) );
  NOR2_X1 U1769 ( .A1(n358), .A2(n260), .ZN(\ab[35][42] ) );
  NOR2_X1 U1770 ( .A1(n361), .A2(n260), .ZN(\ab[35][41] ) );
  NOR2_X1 U1771 ( .A1(n363), .A2(n260), .ZN(\ab[35][40] ) );
  NOR2_X1 U1772 ( .A1(n440), .A2(n260), .ZN(\ab[35][3] ) );
  NOR2_X1 U1773 ( .A1(n365), .A2(n259), .ZN(\ab[35][39] ) );
  NOR2_X1 U1774 ( .A1(n368), .A2(n259), .ZN(\ab[35][38] ) );
  NOR2_X1 U1775 ( .A1(n370), .A2(n259), .ZN(\ab[35][37] ) );
  NOR2_X1 U1776 ( .A1(n372), .A2(n259), .ZN(\ab[35][36] ) );
  NOR2_X1 U1777 ( .A1(n373), .A2(n259), .ZN(\ab[35][35] ) );
  NOR2_X1 U1778 ( .A1(n375), .A2(n259), .ZN(\ab[35][34] ) );
  NOR2_X1 U1779 ( .A1(n377), .A2(n259), .ZN(\ab[35][33] ) );
  NOR2_X1 U1780 ( .A1(n379), .A2(n259), .ZN(\ab[35][32] ) );
  NOR2_X1 U1781 ( .A1(n381), .A2(n259), .ZN(\ab[35][31] ) );
  NOR2_X1 U1782 ( .A1(n383), .A2(n259), .ZN(\ab[35][30] ) );
  NOR2_X1 U1783 ( .A1(n479), .A2(n259), .ZN(\ab[35][2] ) );
  NOR2_X1 U1784 ( .A1(n385), .A2(n261), .ZN(\ab[35][29] ) );
  NOR2_X1 U1785 ( .A1(n387), .A2(n261), .ZN(\ab[35][28] ) );
  NOR2_X1 U1786 ( .A1(n389), .A2(n261), .ZN(\ab[35][27] ) );
  NOR2_X1 U1787 ( .A1(n391), .A2(n261), .ZN(\ab[35][26] ) );
  NOR2_X1 U1788 ( .A1(n393), .A2(n261), .ZN(\ab[35][25] ) );
  NOR2_X1 U1789 ( .A1(n395), .A2(n261), .ZN(\ab[35][24] ) );
  NOR2_X1 U1790 ( .A1(n397), .A2(n260), .ZN(\ab[35][23] ) );
  NOR2_X1 U1791 ( .A1(n399), .A2(n260), .ZN(\ab[35][22] ) );
  NOR2_X1 U1792 ( .A1(n401), .A2(n260), .ZN(\ab[35][21] ) );
  NOR2_X1 U1793 ( .A1(n403), .A2(n261), .ZN(\ab[35][20] ) );
  NOR2_X1 U1794 ( .A1(n444), .A2(n261), .ZN(\ab[35][1] ) );
  NOR2_X1 U1795 ( .A1(n404), .A2(n261), .ZN(\ab[35][19] ) );
  NOR2_X1 U1796 ( .A1(n406), .A2(n261), .ZN(\ab[35][18] ) );
  NOR2_X1 U1797 ( .A1(n408), .A2(n261), .ZN(\ab[35][17] ) );
  NOR2_X1 U1798 ( .A1(n410), .A2(n260), .ZN(\ab[35][16] ) );
  NOR2_X1 U1799 ( .A1(n413), .A2(n259), .ZN(\ab[35][15] ) );
  NOR2_X1 U1800 ( .A1(n416), .A2(n259), .ZN(\ab[35][14] ) );
  NOR2_X1 U1801 ( .A1(n419), .A2(n261), .ZN(\ab[35][13] ) );
  NOR2_X1 U1802 ( .A1(n422), .A2(n261), .ZN(\ab[35][12] ) );
  NOR2_X1 U1803 ( .A1(n425), .A2(n261), .ZN(\ab[35][11] ) );
  NOR2_X1 U1804 ( .A1(n427), .A2(n261), .ZN(\ab[35][10] ) );
  NOR2_X1 U1805 ( .A1(n446), .A2(n261), .ZN(\ab[35][0] ) );
  NOR2_X1 U1806 ( .A1(n428), .A2(n263), .ZN(\ab[34][9] ) );
  NOR2_X1 U1807 ( .A1(n430), .A2(n262), .ZN(\ab[34][8] ) );
  NOR2_X1 U1808 ( .A1(n432), .A2(n262), .ZN(\ab[34][7] ) );
  NOR2_X1 U1809 ( .A1(n435), .A2(n262), .ZN(\ab[34][6] ) );
  NOR2_X1 U1810 ( .A1(n437), .A2(n262), .ZN(\ab[34][5] ) );
  NOR2_X1 U1811 ( .A1(n337), .A2(n262), .ZN(\ab[34][52] ) );
  NOR2_X1 U1812 ( .A1(n338), .A2(n262), .ZN(\ab[34][51] ) );
  NOR2_X1 U1813 ( .A1(n341), .A2(n262), .ZN(\ab[34][50] ) );
  NOR2_X1 U1814 ( .A1(n439), .A2(n262), .ZN(\ab[34][4] ) );
  NOR2_X1 U1815 ( .A1(n343), .A2(n263), .ZN(\ab[34][49] ) );
  NOR2_X1 U1816 ( .A1(n345), .A2(n263), .ZN(\ab[34][48] ) );
  NOR2_X1 U1817 ( .A1(n347), .A2(n263), .ZN(\ab[34][47] ) );
  NOR2_X1 U1818 ( .A1(n349), .A2(n263), .ZN(\ab[34][46] ) );
  NOR2_X1 U1819 ( .A1(n351), .A2(n263), .ZN(\ab[34][45] ) );
  NOR2_X1 U1820 ( .A1(n353), .A2(n263), .ZN(\ab[34][44] ) );
  NOR2_X1 U1821 ( .A1(n356), .A2(n263), .ZN(\ab[34][43] ) );
  NOR2_X1 U1822 ( .A1(n358), .A2(n263), .ZN(\ab[34][42] ) );
  NOR2_X1 U1823 ( .A1(n361), .A2(n263), .ZN(\ab[34][41] ) );
  NOR2_X1 U1824 ( .A1(n363), .A2(n263), .ZN(\ab[34][40] ) );
  NOR2_X1 U1825 ( .A1(n440), .A2(n263), .ZN(\ab[34][3] ) );
  NOR2_X1 U1826 ( .A1(n365), .A2(n262), .ZN(\ab[34][39] ) );
  NOR2_X1 U1827 ( .A1(n367), .A2(n262), .ZN(\ab[34][38] ) );
  NOR2_X1 U1828 ( .A1(n370), .A2(n262), .ZN(\ab[34][37] ) );
  NOR2_X1 U1829 ( .A1(n372), .A2(n262), .ZN(\ab[34][36] ) );
  NOR2_X1 U1830 ( .A1(n373), .A2(n262), .ZN(\ab[34][35] ) );
  NOR2_X1 U1831 ( .A1(n375), .A2(n262), .ZN(\ab[34][34] ) );
  NOR2_X1 U1832 ( .A1(n377), .A2(n262), .ZN(\ab[34][33] ) );
  NOR2_X1 U1833 ( .A1(n379), .A2(n262), .ZN(\ab[34][32] ) );
  NOR2_X1 U1834 ( .A1(n381), .A2(n262), .ZN(\ab[34][31] ) );
  NOR2_X1 U1835 ( .A1(n383), .A2(n262), .ZN(\ab[34][30] ) );
  NOR2_X1 U1836 ( .A1(n479), .A2(n262), .ZN(\ab[34][2] ) );
  NOR2_X1 U1837 ( .A1(n385), .A2(n456), .ZN(\ab[34][29] ) );
  NOR2_X1 U1838 ( .A1(n387), .A2(n456), .ZN(\ab[34][28] ) );
  NOR2_X1 U1839 ( .A1(n389), .A2(n456), .ZN(\ab[34][27] ) );
  NOR2_X1 U1840 ( .A1(n391), .A2(n456), .ZN(\ab[34][26] ) );
  NOR2_X1 U1841 ( .A1(n393), .A2(n456), .ZN(\ab[34][25] ) );
  NOR2_X1 U1842 ( .A1(n395), .A2(n456), .ZN(\ab[34][24] ) );
  NOR2_X1 U1843 ( .A1(n397), .A2(n263), .ZN(\ab[34][23] ) );
  NOR2_X1 U1844 ( .A1(n399), .A2(n263), .ZN(\ab[34][22] ) );
  NOR2_X1 U1845 ( .A1(n401), .A2(n456), .ZN(\ab[34][21] ) );
  NOR2_X1 U1846 ( .A1(n403), .A2(n456), .ZN(\ab[34][20] ) );
  NOR2_X1 U1847 ( .A1(n444), .A2(n456), .ZN(\ab[34][1] ) );
  NOR2_X1 U1848 ( .A1(n405), .A2(n263), .ZN(\ab[34][19] ) );
  NOR2_X1 U1849 ( .A1(n406), .A2(n263), .ZN(\ab[34][18] ) );
  NOR2_X1 U1850 ( .A1(n408), .A2(n456), .ZN(\ab[34][17] ) );
  NOR2_X1 U1851 ( .A1(n410), .A2(n262), .ZN(\ab[34][16] ) );
  NOR2_X1 U1852 ( .A1(n413), .A2(n262), .ZN(\ab[34][15] ) );
  NOR2_X1 U1853 ( .A1(n416), .A2(n262), .ZN(\ab[34][14] ) );
  NOR2_X1 U1854 ( .A1(n419), .A2(n456), .ZN(\ab[34][13] ) );
  NOR2_X1 U1855 ( .A1(n422), .A2(n456), .ZN(\ab[34][12] ) );
  NOR2_X1 U1856 ( .A1(n425), .A2(n456), .ZN(\ab[34][11] ) );
  NOR2_X1 U1857 ( .A1(n427), .A2(n456), .ZN(\ab[34][10] ) );
  NOR2_X1 U1858 ( .A1(n446), .A2(n456), .ZN(\ab[34][0] ) );
  NOR2_X1 U1859 ( .A1(n428), .A2(n265), .ZN(\ab[33][9] ) );
  NOR2_X1 U1860 ( .A1(n430), .A2(n264), .ZN(\ab[33][8] ) );
  NOR2_X1 U1861 ( .A1(n432), .A2(n264), .ZN(\ab[33][7] ) );
  NOR2_X1 U1862 ( .A1(n435), .A2(n264), .ZN(\ab[33][6] ) );
  NOR2_X1 U1863 ( .A1(n437), .A2(n264), .ZN(\ab[33][5] ) );
  NOR2_X1 U1864 ( .A1(n337), .A2(n264), .ZN(\ab[33][52] ) );
  NOR2_X1 U1865 ( .A1(n338), .A2(n264), .ZN(\ab[33][51] ) );
  NOR2_X1 U1866 ( .A1(n341), .A2(n264), .ZN(\ab[33][50] ) );
  NOR2_X1 U1867 ( .A1(n439), .A2(n264), .ZN(\ab[33][4] ) );
  NOR2_X1 U1868 ( .A1(n343), .A2(n265), .ZN(\ab[33][49] ) );
  NOR2_X1 U1869 ( .A1(n345), .A2(n265), .ZN(\ab[33][48] ) );
  NOR2_X1 U1870 ( .A1(n347), .A2(n265), .ZN(\ab[33][47] ) );
  NOR2_X1 U1871 ( .A1(n349), .A2(n265), .ZN(\ab[33][46] ) );
  NOR2_X1 U1872 ( .A1(n351), .A2(n265), .ZN(\ab[33][45] ) );
  NOR2_X1 U1873 ( .A1(n353), .A2(n265), .ZN(\ab[33][44] ) );
  NOR2_X1 U1874 ( .A1(n356), .A2(n265), .ZN(\ab[33][43] ) );
  NOR2_X1 U1875 ( .A1(n358), .A2(n265), .ZN(\ab[33][42] ) );
  NOR2_X1 U1876 ( .A1(n361), .A2(n265), .ZN(\ab[33][41] ) );
  NOR2_X1 U1877 ( .A1(n363), .A2(n265), .ZN(\ab[33][40] ) );
  NOR2_X1 U1878 ( .A1(n440), .A2(n265), .ZN(\ab[33][3] ) );
  NOR2_X1 U1879 ( .A1(n365), .A2(n264), .ZN(\ab[33][39] ) );
  NOR2_X1 U1880 ( .A1(n368), .A2(n264), .ZN(\ab[33][38] ) );
  NOR2_X1 U1881 ( .A1(n370), .A2(n264), .ZN(\ab[33][37] ) );
  NOR2_X1 U1882 ( .A1(n372), .A2(n264), .ZN(\ab[33][36] ) );
  NOR2_X1 U1883 ( .A1(n373), .A2(n264), .ZN(\ab[33][35] ) );
  NOR2_X1 U1884 ( .A1(n375), .A2(n264), .ZN(\ab[33][34] ) );
  NOR2_X1 U1885 ( .A1(n377), .A2(n264), .ZN(\ab[33][33] ) );
  NOR2_X1 U1886 ( .A1(n379), .A2(n264), .ZN(\ab[33][32] ) );
  NOR2_X1 U1887 ( .A1(n381), .A2(n264), .ZN(\ab[33][31] ) );
  NOR2_X1 U1888 ( .A1(n383), .A2(n264), .ZN(\ab[33][30] ) );
  NOR2_X1 U1889 ( .A1(n479), .A2(n264), .ZN(\ab[33][2] ) );
  NOR2_X1 U1890 ( .A1(n385), .A2(n457), .ZN(\ab[33][29] ) );
  NOR2_X1 U1891 ( .A1(n387), .A2(n457), .ZN(\ab[33][28] ) );
  NOR2_X1 U1892 ( .A1(n389), .A2(n457), .ZN(\ab[33][27] ) );
  NOR2_X1 U1893 ( .A1(n391), .A2(n457), .ZN(\ab[33][26] ) );
  NOR2_X1 U1894 ( .A1(n393), .A2(n457), .ZN(\ab[33][25] ) );
  NOR2_X1 U1895 ( .A1(n395), .A2(n457), .ZN(\ab[33][24] ) );
  NOR2_X1 U1896 ( .A1(n397), .A2(n457), .ZN(\ab[33][23] ) );
  NOR2_X1 U1897 ( .A1(n399), .A2(n457), .ZN(\ab[33][22] ) );
  NOR2_X1 U1898 ( .A1(n401), .A2(n457), .ZN(\ab[33][21] ) );
  NOR2_X1 U1899 ( .A1(n403), .A2(n265), .ZN(\ab[33][20] ) );
  NOR2_X1 U1900 ( .A1(n444), .A2(n457), .ZN(\ab[33][1] ) );
  NOR2_X1 U1901 ( .A1(n404), .A2(n265), .ZN(\ab[33][19] ) );
  NOR2_X1 U1902 ( .A1(n406), .A2(n265), .ZN(\ab[33][18] ) );
  NOR2_X1 U1903 ( .A1(n408), .A2(n264), .ZN(\ab[33][17] ) );
  NOR2_X1 U1904 ( .A1(n410), .A2(n264), .ZN(\ab[33][16] ) );
  NOR2_X1 U1905 ( .A1(n413), .A2(n264), .ZN(\ab[33][15] ) );
  NOR2_X1 U1906 ( .A1(n416), .A2(n264), .ZN(\ab[33][14] ) );
  NOR2_X1 U1907 ( .A1(n419), .A2(n264), .ZN(\ab[33][13] ) );
  NOR2_X1 U1908 ( .A1(n422), .A2(n265), .ZN(\ab[33][12] ) );
  NOR2_X1 U1909 ( .A1(n425), .A2(n264), .ZN(\ab[33][11] ) );
  NOR2_X1 U1910 ( .A1(n427), .A2(n265), .ZN(\ab[33][10] ) );
  NOR2_X1 U1911 ( .A1(n446), .A2(n264), .ZN(\ab[33][0] ) );
  NOR2_X1 U1912 ( .A1(n428), .A2(n267), .ZN(\ab[32][9] ) );
  NOR2_X1 U1913 ( .A1(n430), .A2(n267), .ZN(\ab[32][8] ) );
  NOR2_X1 U1914 ( .A1(n432), .A2(n267), .ZN(\ab[32][7] ) );
  NOR2_X1 U1915 ( .A1(n435), .A2(n267), .ZN(\ab[32][6] ) );
  NOR2_X1 U1916 ( .A1(n437), .A2(n267), .ZN(\ab[32][5] ) );
  NOR2_X1 U1917 ( .A1(n337), .A2(n267), .ZN(\ab[32][52] ) );
  NOR2_X1 U1918 ( .A1(n338), .A2(n267), .ZN(\ab[32][51] ) );
  NOR2_X1 U1919 ( .A1(n341), .A2(n267), .ZN(\ab[32][50] ) );
  NOR2_X1 U1920 ( .A1(n439), .A2(n267), .ZN(\ab[32][4] ) );
  NOR2_X1 U1921 ( .A1(n343), .A2(n266), .ZN(\ab[32][49] ) );
  NOR2_X1 U1922 ( .A1(n345), .A2(n266), .ZN(\ab[32][48] ) );
  NOR2_X1 U1923 ( .A1(n347), .A2(n266), .ZN(\ab[32][47] ) );
  NOR2_X1 U1924 ( .A1(n349), .A2(n266), .ZN(\ab[32][46] ) );
  NOR2_X1 U1925 ( .A1(n351), .A2(n266), .ZN(\ab[32][45] ) );
  NOR2_X1 U1926 ( .A1(n353), .A2(n266), .ZN(\ab[32][44] ) );
  NOR2_X1 U1927 ( .A1(n356), .A2(n266), .ZN(\ab[32][43] ) );
  NOR2_X1 U1928 ( .A1(n358), .A2(n266), .ZN(\ab[32][42] ) );
  NOR2_X1 U1929 ( .A1(n361), .A2(n266), .ZN(\ab[32][41] ) );
  NOR2_X1 U1930 ( .A1(n363), .A2(n266), .ZN(\ab[32][40] ) );
  NOR2_X1 U1931 ( .A1(n440), .A2(n266), .ZN(\ab[32][3] ) );
  NOR2_X1 U1932 ( .A1(n365), .A2(n266), .ZN(\ab[32][39] ) );
  NOR2_X1 U1933 ( .A1(n367), .A2(n266), .ZN(\ab[32][38] ) );
  NOR2_X1 U1934 ( .A1(n370), .A2(n266), .ZN(\ab[32][37] ) );
  NOR2_X1 U1935 ( .A1(n372), .A2(n266), .ZN(\ab[32][36] ) );
  NOR2_X1 U1936 ( .A1(n373), .A2(n266), .ZN(\ab[32][35] ) );
  NOR2_X1 U1937 ( .A1(n375), .A2(n266), .ZN(\ab[32][34] ) );
  NOR2_X1 U1938 ( .A1(n377), .A2(n266), .ZN(\ab[32][33] ) );
  NOR2_X1 U1939 ( .A1(n379), .A2(n266), .ZN(\ab[32][32] ) );
  NOR2_X1 U1940 ( .A1(n381), .A2(n266), .ZN(\ab[32][31] ) );
  NOR2_X1 U1941 ( .A1(n383), .A2(n266), .ZN(\ab[32][30] ) );
  NOR2_X1 U1942 ( .A1(n479), .A2(n266), .ZN(\ab[32][2] ) );
  NOR2_X1 U1943 ( .A1(n385), .A2(n458), .ZN(\ab[32][29] ) );
  NOR2_X1 U1944 ( .A1(n387), .A2(n458), .ZN(\ab[32][28] ) );
  NOR2_X1 U1945 ( .A1(n389), .A2(n458), .ZN(\ab[32][27] ) );
  NOR2_X1 U1946 ( .A1(n391), .A2(n458), .ZN(\ab[32][26] ) );
  NOR2_X1 U1947 ( .A1(n393), .A2(n458), .ZN(\ab[32][25] ) );
  NOR2_X1 U1948 ( .A1(n395), .A2(n266), .ZN(\ab[32][24] ) );
  NOR2_X1 U1949 ( .A1(n397), .A2(n458), .ZN(\ab[32][23] ) );
  NOR2_X1 U1950 ( .A1(n399), .A2(n458), .ZN(\ab[32][22] ) );
  NOR2_X1 U1951 ( .A1(n401), .A2(n458), .ZN(\ab[32][21] ) );
  NOR2_X1 U1952 ( .A1(n403), .A2(n458), .ZN(\ab[32][20] ) );
  NOR2_X1 U1953 ( .A1(n444), .A2(n458), .ZN(\ab[32][1] ) );
  NOR2_X1 U1954 ( .A1(n405), .A2(n267), .ZN(\ab[32][19] ) );
  NOR2_X1 U1955 ( .A1(n406), .A2(n267), .ZN(\ab[32][18] ) );
  NOR2_X1 U1956 ( .A1(n408), .A2(n267), .ZN(\ab[32][17] ) );
  NOR2_X1 U1957 ( .A1(n410), .A2(n267), .ZN(\ab[32][16] ) );
  NOR2_X1 U1958 ( .A1(n413), .A2(n266), .ZN(\ab[32][15] ) );
  NOR2_X1 U1959 ( .A1(n416), .A2(n267), .ZN(\ab[32][14] ) );
  NOR2_X1 U1960 ( .A1(n419), .A2(n267), .ZN(\ab[32][13] ) );
  NOR2_X1 U1961 ( .A1(n422), .A2(n266), .ZN(\ab[32][12] ) );
  NOR2_X1 U1962 ( .A1(n425), .A2(n267), .ZN(\ab[32][11] ) );
  NOR2_X1 U1963 ( .A1(n427), .A2(n267), .ZN(\ab[32][10] ) );
  NOR2_X1 U1964 ( .A1(n446), .A2(n267), .ZN(\ab[32][0] ) );
  NOR2_X1 U1965 ( .A1(n428), .A2(n269), .ZN(\ab[31][9] ) );
  NOR2_X1 U1966 ( .A1(n430), .A2(n269), .ZN(\ab[31][8] ) );
  NOR2_X1 U1967 ( .A1(n432), .A2(n269), .ZN(\ab[31][7] ) );
  NOR2_X1 U1968 ( .A1(n435), .A2(n269), .ZN(\ab[31][6] ) );
  NOR2_X1 U1969 ( .A1(n437), .A2(n269), .ZN(\ab[31][5] ) );
  NOR2_X1 U1970 ( .A1(n337), .A2(n269), .ZN(\ab[31][52] ) );
  NOR2_X1 U1971 ( .A1(n338), .A2(n269), .ZN(\ab[31][51] ) );
  NOR2_X1 U1972 ( .A1(n341), .A2(n269), .ZN(\ab[31][50] ) );
  NOR2_X1 U1973 ( .A1(n439), .A2(n269), .ZN(\ab[31][4] ) );
  NOR2_X1 U1974 ( .A1(n343), .A2(n268), .ZN(\ab[31][49] ) );
  NOR2_X1 U1975 ( .A1(n345), .A2(n268), .ZN(\ab[31][48] ) );
  NOR2_X1 U1976 ( .A1(n347), .A2(n268), .ZN(\ab[31][47] ) );
  NOR2_X1 U1977 ( .A1(n349), .A2(n268), .ZN(\ab[31][46] ) );
  NOR2_X1 U1978 ( .A1(n351), .A2(n268), .ZN(\ab[31][45] ) );
  NOR2_X1 U1979 ( .A1(n353), .A2(n268), .ZN(\ab[31][44] ) );
  NOR2_X1 U1980 ( .A1(n356), .A2(n268), .ZN(\ab[31][43] ) );
  NOR2_X1 U1981 ( .A1(n358), .A2(n268), .ZN(\ab[31][42] ) );
  NOR2_X1 U1982 ( .A1(n361), .A2(n268), .ZN(\ab[31][41] ) );
  NOR2_X1 U1983 ( .A1(n363), .A2(n268), .ZN(\ab[31][40] ) );
  NOR2_X1 U1984 ( .A1(n441), .A2(n268), .ZN(\ab[31][3] ) );
  NOR2_X1 U1985 ( .A1(n365), .A2(n268), .ZN(\ab[31][39] ) );
  NOR2_X1 U1986 ( .A1(n368), .A2(n268), .ZN(\ab[31][38] ) );
  NOR2_X1 U1987 ( .A1(n370), .A2(n268), .ZN(\ab[31][37] ) );
  NOR2_X1 U1988 ( .A1(n372), .A2(n268), .ZN(\ab[31][36] ) );
  NOR2_X1 U1989 ( .A1(n373), .A2(n268), .ZN(\ab[31][35] ) );
  NOR2_X1 U1990 ( .A1(n375), .A2(n268), .ZN(\ab[31][34] ) );
  NOR2_X1 U1991 ( .A1(n377), .A2(n268), .ZN(\ab[31][33] ) );
  NOR2_X1 U1992 ( .A1(n379), .A2(n268), .ZN(\ab[31][32] ) );
  NOR2_X1 U1993 ( .A1(n381), .A2(n268), .ZN(\ab[31][31] ) );
  NOR2_X1 U1994 ( .A1(n383), .A2(n268), .ZN(\ab[31][30] ) );
  NOR2_X1 U1995 ( .A1(n479), .A2(n268), .ZN(\ab[31][2] ) );
  NOR2_X1 U1996 ( .A1(n385), .A2(n268), .ZN(\ab[31][29] ) );
  NOR2_X1 U1997 ( .A1(n387), .A2(n268), .ZN(\ab[31][28] ) );
  NOR2_X1 U1998 ( .A1(n389), .A2(n268), .ZN(\ab[31][27] ) );
  NOR2_X1 U1999 ( .A1(n391), .A2(n268), .ZN(\ab[31][26] ) );
  NOR2_X1 U2000 ( .A1(n393), .A2(n459), .ZN(\ab[31][25] ) );
  NOR2_X1 U2001 ( .A1(n395), .A2(n459), .ZN(\ab[31][24] ) );
  NOR2_X1 U2002 ( .A1(n397), .A2(n459), .ZN(\ab[31][23] ) );
  NOR2_X1 U2003 ( .A1(n399), .A2(n459), .ZN(\ab[31][22] ) );
  NOR2_X1 U2004 ( .A1(n401), .A2(n459), .ZN(\ab[31][21] ) );
  NOR2_X1 U2005 ( .A1(n403), .A2(n459), .ZN(\ab[31][20] ) );
  NOR2_X1 U2006 ( .A1(n444), .A2(n268), .ZN(\ab[31][1] ) );
  NOR2_X1 U2007 ( .A1(n404), .A2(n269), .ZN(\ab[31][19] ) );
  NOR2_X1 U2008 ( .A1(n406), .A2(n269), .ZN(\ab[31][18] ) );
  NOR2_X1 U2009 ( .A1(n408), .A2(n269), .ZN(\ab[31][17] ) );
  NOR2_X1 U2010 ( .A1(n410), .A2(n269), .ZN(\ab[31][16] ) );
  NOR2_X1 U2011 ( .A1(n413), .A2(n268), .ZN(\ab[31][15] ) );
  NOR2_X1 U2012 ( .A1(n416), .A2(n269), .ZN(\ab[31][14] ) );
  NOR2_X1 U2013 ( .A1(n419), .A2(n269), .ZN(\ab[31][13] ) );
  NOR2_X1 U2014 ( .A1(n422), .A2(n268), .ZN(\ab[31][12] ) );
  NOR2_X1 U2015 ( .A1(n425), .A2(n269), .ZN(\ab[31][11] ) );
  NOR2_X1 U2016 ( .A1(n427), .A2(n269), .ZN(\ab[31][10] ) );
  NOR2_X1 U2017 ( .A1(n446), .A2(n269), .ZN(\ab[31][0] ) );
  NOR2_X1 U2018 ( .A1(n428), .A2(n271), .ZN(\ab[30][9] ) );
  NOR2_X1 U2019 ( .A1(n430), .A2(n270), .ZN(\ab[30][8] ) );
  NOR2_X1 U2020 ( .A1(n432), .A2(n270), .ZN(\ab[30][7] ) );
  NOR2_X1 U2021 ( .A1(n435), .A2(n270), .ZN(\ab[30][6] ) );
  NOR2_X1 U2022 ( .A1(n437), .A2(n270), .ZN(\ab[30][5] ) );
  NOR2_X1 U2023 ( .A1(n337), .A2(n270), .ZN(\ab[30][52] ) );
  NOR2_X1 U2024 ( .A1(n338), .A2(n270), .ZN(\ab[30][51] ) );
  NOR2_X1 U2025 ( .A1(n341), .A2(n270), .ZN(\ab[30][50] ) );
  NOR2_X1 U2026 ( .A1(n439), .A2(n270), .ZN(\ab[30][4] ) );
  NOR2_X1 U2027 ( .A1(n343), .A2(n271), .ZN(\ab[30][49] ) );
  NOR2_X1 U2028 ( .A1(n345), .A2(n271), .ZN(\ab[30][48] ) );
  NOR2_X1 U2029 ( .A1(n347), .A2(n271), .ZN(\ab[30][47] ) );
  NOR2_X1 U2030 ( .A1(n349), .A2(n271), .ZN(\ab[30][46] ) );
  NOR2_X1 U2031 ( .A1(n351), .A2(n271), .ZN(\ab[30][45] ) );
  NOR2_X1 U2032 ( .A1(n353), .A2(n271), .ZN(\ab[30][44] ) );
  NOR2_X1 U2033 ( .A1(n356), .A2(n271), .ZN(\ab[30][43] ) );
  NOR2_X1 U2034 ( .A1(n358), .A2(n271), .ZN(\ab[30][42] ) );
  NOR2_X1 U2035 ( .A1(n361), .A2(n271), .ZN(\ab[30][41] ) );
  NOR2_X1 U2036 ( .A1(n363), .A2(n271), .ZN(\ab[30][40] ) );
  NOR2_X1 U2037 ( .A1(n441), .A2(n271), .ZN(\ab[30][3] ) );
  NOR2_X1 U2038 ( .A1(n365), .A2(n270), .ZN(\ab[30][39] ) );
  NOR2_X1 U2039 ( .A1(n367), .A2(n270), .ZN(\ab[30][38] ) );
  NOR2_X1 U2040 ( .A1(n370), .A2(n270), .ZN(\ab[30][37] ) );
  NOR2_X1 U2041 ( .A1(n372), .A2(n270), .ZN(\ab[30][36] ) );
  NOR2_X1 U2042 ( .A1(n373), .A2(n270), .ZN(\ab[30][35] ) );
  NOR2_X1 U2043 ( .A1(n375), .A2(n270), .ZN(\ab[30][34] ) );
  NOR2_X1 U2044 ( .A1(n377), .A2(n270), .ZN(\ab[30][33] ) );
  NOR2_X1 U2045 ( .A1(n379), .A2(n270), .ZN(\ab[30][32] ) );
  NOR2_X1 U2046 ( .A1(n381), .A2(n270), .ZN(\ab[30][31] ) );
  NOR2_X1 U2047 ( .A1(n383), .A2(n270), .ZN(\ab[30][30] ) );
  NOR2_X1 U2048 ( .A1(n479), .A2(n270), .ZN(\ab[30][2] ) );
  NOR2_X1 U2049 ( .A1(n385), .A2(n460), .ZN(\ab[30][29] ) );
  NOR2_X1 U2050 ( .A1(n387), .A2(n460), .ZN(\ab[30][28] ) );
  NOR2_X1 U2051 ( .A1(n389), .A2(n460), .ZN(\ab[30][27] ) );
  NOR2_X1 U2052 ( .A1(n391), .A2(n271), .ZN(\ab[30][26] ) );
  NOR2_X1 U2053 ( .A1(n393), .A2(n460), .ZN(\ab[30][25] ) );
  NOR2_X1 U2054 ( .A1(n395), .A2(n460), .ZN(\ab[30][24] ) );
  NOR2_X1 U2055 ( .A1(n397), .A2(n460), .ZN(\ab[30][23] ) );
  NOR2_X1 U2056 ( .A1(n399), .A2(n460), .ZN(\ab[30][22] ) );
  NOR2_X1 U2057 ( .A1(n401), .A2(n460), .ZN(\ab[30][21] ) );
  NOR2_X1 U2058 ( .A1(n403), .A2(n460), .ZN(\ab[30][20] ) );
  NOR2_X1 U2059 ( .A1(n444), .A2(n460), .ZN(\ab[30][1] ) );
  NOR2_X1 U2060 ( .A1(n405), .A2(n271), .ZN(\ab[30][19] ) );
  NOR2_X1 U2061 ( .A1(n406), .A2(n271), .ZN(\ab[30][18] ) );
  NOR2_X1 U2062 ( .A1(n408), .A2(n270), .ZN(\ab[30][17] ) );
  NOR2_X1 U2063 ( .A1(n410), .A2(n270), .ZN(\ab[30][16] ) );
  NOR2_X1 U2064 ( .A1(n413), .A2(n270), .ZN(\ab[30][15] ) );
  NOR2_X1 U2065 ( .A1(n416), .A2(n270), .ZN(\ab[30][14] ) );
  NOR2_X1 U2066 ( .A1(n419), .A2(n270), .ZN(\ab[30][13] ) );
  NOR2_X1 U2067 ( .A1(n422), .A2(n271), .ZN(\ab[30][12] ) );
  NOR2_X1 U2068 ( .A1(n425), .A2(n270), .ZN(\ab[30][11] ) );
  NOR2_X1 U2069 ( .A1(n427), .A2(n271), .ZN(\ab[30][10] ) );
  NOR2_X1 U2070 ( .A1(n446), .A2(n270), .ZN(\ab[30][0] ) );
  NOR2_X1 U2071 ( .A1(n428), .A2(n327), .ZN(\ab[2][9] ) );
  NOR2_X1 U2072 ( .A1(n430), .A2(n327), .ZN(\ab[2][8] ) );
  NOR2_X1 U2073 ( .A1(n432), .A2(n327), .ZN(\ab[2][7] ) );
  NOR2_X1 U2074 ( .A1(n435), .A2(n327), .ZN(\ab[2][6] ) );
  NOR2_X1 U2075 ( .A1(n437), .A2(n327), .ZN(\ab[2][5] ) );
  NOR2_X1 U2076 ( .A1(n337), .A2(n328), .ZN(\ab[2][52] ) );
  NOR2_X1 U2077 ( .A1(n338), .A2(n328), .ZN(\ab[2][51] ) );
  NOR2_X1 U2078 ( .A1(n342), .A2(n329), .ZN(\ab[2][50] ) );
  NOR2_X1 U2079 ( .A1(n439), .A2(n327), .ZN(\ab[2][4] ) );
  NOR2_X1 U2080 ( .A1(n343), .A2(n329), .ZN(\ab[2][49] ) );
  NOR2_X1 U2081 ( .A1(n345), .A2(n329), .ZN(\ab[2][48] ) );
  NOR2_X1 U2082 ( .A1(n347), .A2(n329), .ZN(\ab[2][47] ) );
  NOR2_X1 U2083 ( .A1(n349), .A2(n329), .ZN(\ab[2][46] ) );
  NOR2_X1 U2084 ( .A1(n351), .A2(n329), .ZN(\ab[2][45] ) );
  NOR2_X1 U2085 ( .A1(n353), .A2(n329), .ZN(\ab[2][44] ) );
  NOR2_X1 U2086 ( .A1(n356), .A2(n329), .ZN(\ab[2][43] ) );
  NOR2_X1 U2087 ( .A1(n358), .A2(n329), .ZN(\ab[2][42] ) );
  NOR2_X1 U2088 ( .A1(n361), .A2(n329), .ZN(\ab[2][41] ) );
  NOR2_X1 U2089 ( .A1(n363), .A2(n329), .ZN(\ab[2][40] ) );
  NOR2_X1 U2090 ( .A1(n441), .A2(n329), .ZN(\ab[2][3] ) );
  NOR2_X1 U2091 ( .A1(n365), .A2(n328), .ZN(\ab[2][39] ) );
  NOR2_X1 U2092 ( .A1(n367), .A2(n328), .ZN(\ab[2][38] ) );
  NOR2_X1 U2093 ( .A1(n370), .A2(n328), .ZN(\ab[2][37] ) );
  NOR2_X1 U2094 ( .A1(n372), .A2(n328), .ZN(\ab[2][36] ) );
  NOR2_X1 U2095 ( .A1(n373), .A2(n328), .ZN(\ab[2][35] ) );
  NOR2_X1 U2096 ( .A1(n375), .A2(n328), .ZN(\ab[2][34] ) );
  NOR2_X1 U2097 ( .A1(n377), .A2(n328), .ZN(\ab[2][33] ) );
  NOR2_X1 U2098 ( .A1(n379), .A2(n328), .ZN(\ab[2][32] ) );
  NOR2_X1 U2099 ( .A1(n381), .A2(n328), .ZN(\ab[2][31] ) );
  NOR2_X1 U2100 ( .A1(n383), .A2(n328), .ZN(\ab[2][30] ) );
  NOR2_X1 U2101 ( .A1(n442), .A2(n328), .ZN(\ab[2][2] ) );
  NOR2_X1 U2102 ( .A1(n385), .A2(n327), .ZN(\ab[2][29] ) );
  NOR2_X1 U2103 ( .A1(n387), .A2(n327), .ZN(\ab[2][28] ) );
  NOR2_X1 U2104 ( .A1(n389), .A2(n327), .ZN(\ab[2][27] ) );
  NOR2_X1 U2105 ( .A1(n391), .A2(n327), .ZN(\ab[2][26] ) );
  NOR2_X1 U2106 ( .A1(n393), .A2(n327), .ZN(\ab[2][25] ) );
  NOR2_X1 U2107 ( .A1(n395), .A2(n327), .ZN(\ab[2][24] ) );
  NOR2_X1 U2108 ( .A1(n397), .A2(n327), .ZN(\ab[2][23] ) );
  NOR2_X1 U2109 ( .A1(n399), .A2(n327), .ZN(\ab[2][22] ) );
  NOR2_X1 U2110 ( .A1(n401), .A2(n327), .ZN(\ab[2][21] ) );
  NOR2_X1 U2111 ( .A1(n403), .A2(n327), .ZN(\ab[2][20] ) );
  NOR2_X1 U2112 ( .A1(n445), .A2(n327), .ZN(\ab[2][1] ) );
  NOR2_X1 U2113 ( .A1(n405), .A2(n327), .ZN(\ab[2][19] ) );
  NOR2_X1 U2114 ( .A1(n406), .A2(n327), .ZN(\ab[2][18] ) );
  NOR2_X1 U2115 ( .A1(n408), .A2(n327), .ZN(\ab[2][17] ) );
  NOR2_X1 U2116 ( .A1(n410), .A2(n327), .ZN(\ab[2][16] ) );
  NOR2_X1 U2117 ( .A1(n413), .A2(n327), .ZN(\ab[2][15] ) );
  NOR2_X1 U2118 ( .A1(n416), .A2(n327), .ZN(\ab[2][14] ) );
  NOR2_X1 U2119 ( .A1(n419), .A2(n327), .ZN(\ab[2][13] ) );
  NOR2_X1 U2120 ( .A1(n422), .A2(n327), .ZN(\ab[2][12] ) );
  NOR2_X1 U2121 ( .A1(n425), .A2(n327), .ZN(\ab[2][11] ) );
  NOR2_X1 U2122 ( .A1(n427), .A2(n327), .ZN(\ab[2][10] ) );
  NOR2_X1 U2123 ( .A1(n446), .A2(n327), .ZN(\ab[2][0] ) );
  NOR2_X1 U2124 ( .A1(n429), .A2(n272), .ZN(\ab[29][9] ) );
  NOR2_X1 U2125 ( .A1(n431), .A2(n273), .ZN(\ab[29][8] ) );
  NOR2_X1 U2126 ( .A1(n433), .A2(n273), .ZN(\ab[29][7] ) );
  NOR2_X1 U2127 ( .A1(n434), .A2(n273), .ZN(\ab[29][6] ) );
  NOR2_X1 U2128 ( .A1(n436), .A2(n273), .ZN(\ab[29][5] ) );
  NOR2_X1 U2129 ( .A1(n336), .A2(n273), .ZN(\ab[29][52] ) );
  NOR2_X1 U2130 ( .A1(n339), .A2(n273), .ZN(\ab[29][51] ) );
  NOR2_X1 U2131 ( .A1(n341), .A2(n273), .ZN(\ab[29][50] ) );
  NOR2_X1 U2132 ( .A1(n438), .A2(n273), .ZN(\ab[29][4] ) );
  NOR2_X1 U2133 ( .A1(n344), .A2(n273), .ZN(\ab[29][49] ) );
  NOR2_X1 U2134 ( .A1(n345), .A2(n273), .ZN(\ab[29][48] ) );
  NOR2_X1 U2135 ( .A1(n347), .A2(n273), .ZN(\ab[29][47] ) );
  NOR2_X1 U2136 ( .A1(n349), .A2(n273), .ZN(\ab[29][46] ) );
  NOR2_X1 U2137 ( .A1(n351), .A2(n273), .ZN(\ab[29][45] ) );
  NOR2_X1 U2138 ( .A1(n354), .A2(n273), .ZN(\ab[29][44] ) );
  NOR2_X1 U2139 ( .A1(n357), .A2(n273), .ZN(\ab[29][43] ) );
  NOR2_X1 U2140 ( .A1(n359), .A2(n273), .ZN(\ab[29][42] ) );
  NOR2_X1 U2141 ( .A1(n361), .A2(n273), .ZN(\ab[29][41] ) );
  NOR2_X1 U2142 ( .A1(n363), .A2(n273), .ZN(\ab[29][40] ) );
  NOR2_X1 U2143 ( .A1(n440), .A2(n273), .ZN(\ab[29][3] ) );
  NOR2_X1 U2144 ( .A1(n365), .A2(n272), .ZN(\ab[29][39] ) );
  NOR2_X1 U2145 ( .A1(n369), .A2(n272), .ZN(\ab[29][38] ) );
  NOR2_X1 U2146 ( .A1(n371), .A2(n272), .ZN(\ab[29][37] ) );
  NOR2_X1 U2147 ( .A1(n474), .A2(n272), .ZN(\ab[29][36] ) );
  NOR2_X1 U2148 ( .A1(n373), .A2(n272), .ZN(\ab[29][35] ) );
  NOR2_X1 U2149 ( .A1(n375), .A2(n272), .ZN(\ab[29][34] ) );
  NOR2_X1 U2150 ( .A1(n377), .A2(n272), .ZN(\ab[29][33] ) );
  NOR2_X1 U2151 ( .A1(n380), .A2(n272), .ZN(\ab[29][32] ) );
  NOR2_X1 U2152 ( .A1(n381), .A2(n272), .ZN(\ab[29][31] ) );
  NOR2_X1 U2153 ( .A1(n383), .A2(n272), .ZN(\ab[29][30] ) );
  NOR2_X1 U2154 ( .A1(n442), .A2(n272), .ZN(\ab[29][2] ) );
  NOR2_X1 U2155 ( .A1(n386), .A2(n273), .ZN(\ab[29][29] ) );
  NOR2_X1 U2156 ( .A1(n388), .A2(n273), .ZN(\ab[29][28] ) );
  NOR2_X1 U2157 ( .A1(n390), .A2(n272), .ZN(\ab[29][27] ) );
  NOR2_X1 U2158 ( .A1(n392), .A2(n274), .ZN(\ab[29][26] ) );
  NOR2_X1 U2159 ( .A1(n393), .A2(n274), .ZN(\ab[29][25] ) );
  NOR2_X1 U2160 ( .A1(n395), .A2(n274), .ZN(\ab[29][24] ) );
  NOR2_X1 U2161 ( .A1(n397), .A2(n274), .ZN(\ab[29][23] ) );
  NOR2_X1 U2162 ( .A1(n400), .A2(n274), .ZN(\ab[29][22] ) );
  NOR2_X1 U2163 ( .A1(n402), .A2(n274), .ZN(\ab[29][21] ) );
  NOR2_X1 U2164 ( .A1(n403), .A2(n272), .ZN(\ab[29][20] ) );
  NOR2_X1 U2165 ( .A1(n443), .A2(n273), .ZN(\ab[29][1] ) );
  NOR2_X1 U2166 ( .A1(n404), .A2(n272), .ZN(\ab[29][19] ) );
  NOR2_X1 U2167 ( .A1(n476), .A2(n272), .ZN(\ab[29][18] ) );
  NOR2_X1 U2168 ( .A1(n408), .A2(n273), .ZN(\ab[29][17] ) );
  NOR2_X1 U2169 ( .A1(n411), .A2(n273), .ZN(\ab[29][16] ) );
  NOR2_X1 U2170 ( .A1(n414), .A2(n273), .ZN(\ab[29][15] ) );
  NOR2_X1 U2171 ( .A1(n417), .A2(n273), .ZN(\ab[29][14] ) );
  NOR2_X1 U2172 ( .A1(n420), .A2(n273), .ZN(\ab[29][13] ) );
  NOR2_X1 U2173 ( .A1(n423), .A2(n272), .ZN(\ab[29][12] ) );
  NOR2_X1 U2174 ( .A1(n425), .A2(n273), .ZN(\ab[29][11] ) );
  NOR2_X1 U2175 ( .A1(n427), .A2(n272), .ZN(\ab[29][10] ) );
  NOR2_X1 U2176 ( .A1(n446), .A2(n273), .ZN(\ab[29][0] ) );
  NOR2_X1 U2177 ( .A1(n429), .A2(n276), .ZN(\ab[28][9] ) );
  NOR2_X1 U2178 ( .A1(n431), .A2(n276), .ZN(\ab[28][8] ) );
  NOR2_X1 U2179 ( .A1(n433), .A2(n276), .ZN(\ab[28][7] ) );
  NOR2_X1 U2180 ( .A1(n434), .A2(n276), .ZN(\ab[28][6] ) );
  NOR2_X1 U2181 ( .A1(n436), .A2(n276), .ZN(\ab[28][5] ) );
  NOR2_X1 U2182 ( .A1(n336), .A2(n276), .ZN(\ab[28][52] ) );
  NOR2_X1 U2183 ( .A1(n339), .A2(n276), .ZN(\ab[28][51] ) );
  NOR2_X1 U2184 ( .A1(n341), .A2(n276), .ZN(\ab[28][50] ) );
  NOR2_X1 U2185 ( .A1(n438), .A2(n276), .ZN(\ab[28][4] ) );
  NOR2_X1 U2186 ( .A1(n343), .A2(n276), .ZN(\ab[28][49] ) );
  NOR2_X1 U2187 ( .A1(n345), .A2(n276), .ZN(\ab[28][48] ) );
  NOR2_X1 U2188 ( .A1(n347), .A2(n276), .ZN(\ab[28][47] ) );
  NOR2_X1 U2189 ( .A1(n349), .A2(n276), .ZN(\ab[28][46] ) );
  NOR2_X1 U2190 ( .A1(n351), .A2(n276), .ZN(\ab[28][45] ) );
  NOR2_X1 U2191 ( .A1(n354), .A2(n276), .ZN(\ab[28][44] ) );
  NOR2_X1 U2192 ( .A1(n356), .A2(n276), .ZN(\ab[28][43] ) );
  NOR2_X1 U2193 ( .A1(n359), .A2(n276), .ZN(\ab[28][42] ) );
  NOR2_X1 U2194 ( .A1(n361), .A2(n276), .ZN(\ab[28][41] ) );
  NOR2_X1 U2195 ( .A1(n363), .A2(n276), .ZN(\ab[28][40] ) );
  NOR2_X1 U2196 ( .A1(n440), .A2(n276), .ZN(\ab[28][3] ) );
  NOR2_X1 U2197 ( .A1(n365), .A2(n275), .ZN(\ab[28][39] ) );
  NOR2_X1 U2198 ( .A1(n369), .A2(n275), .ZN(\ab[28][38] ) );
  NOR2_X1 U2199 ( .A1(n370), .A2(n275), .ZN(\ab[28][37] ) );
  NOR2_X1 U2200 ( .A1(n372), .A2(n275), .ZN(\ab[28][36] ) );
  NOR2_X1 U2201 ( .A1(n373), .A2(n275), .ZN(\ab[28][35] ) );
  NOR2_X1 U2202 ( .A1(n375), .A2(n275), .ZN(\ab[28][34] ) );
  NOR2_X1 U2203 ( .A1(n377), .A2(n275), .ZN(\ab[28][33] ) );
  NOR2_X1 U2204 ( .A1(n379), .A2(n275), .ZN(\ab[28][32] ) );
  NOR2_X1 U2205 ( .A1(n381), .A2(n275), .ZN(\ab[28][31] ) );
  NOR2_X1 U2206 ( .A1(n383), .A2(n275), .ZN(\ab[28][30] ) );
  NOR2_X1 U2207 ( .A1(n442), .A2(n275), .ZN(\ab[28][2] ) );
  NOR2_X1 U2208 ( .A1(n385), .A2(n275), .ZN(\ab[28][29] ) );
  NOR2_X1 U2209 ( .A1(n388), .A2(n277), .ZN(\ab[28][28] ) );
  NOR2_X1 U2210 ( .A1(n389), .A2(n277), .ZN(\ab[28][27] ) );
  NOR2_X1 U2211 ( .A1(n391), .A2(n277), .ZN(\ab[28][26] ) );
  NOR2_X1 U2212 ( .A1(n394), .A2(n277), .ZN(\ab[28][25] ) );
  NOR2_X1 U2213 ( .A1(n396), .A2(n277), .ZN(\ab[28][24] ) );
  NOR2_X1 U2214 ( .A1(n398), .A2(n277), .ZN(\ab[28][23] ) );
  NOR2_X1 U2215 ( .A1(n399), .A2(n277), .ZN(\ab[28][22] ) );
  NOR2_X1 U2216 ( .A1(n401), .A2(n275), .ZN(\ab[28][21] ) );
  NOR2_X1 U2217 ( .A1(n403), .A2(n276), .ZN(\ab[28][20] ) );
  NOR2_X1 U2218 ( .A1(n443), .A2(n276), .ZN(\ab[28][1] ) );
  NOR2_X1 U2219 ( .A1(n404), .A2(n275), .ZN(\ab[28][19] ) );
  NOR2_X1 U2220 ( .A1(n476), .A2(n275), .ZN(\ab[28][18] ) );
  NOR2_X1 U2221 ( .A1(n408), .A2(n275), .ZN(\ab[28][17] ) );
  NOR2_X1 U2222 ( .A1(n411), .A2(n276), .ZN(\ab[28][16] ) );
  NOR2_X1 U2223 ( .A1(n414), .A2(n276), .ZN(\ab[28][15] ) );
  NOR2_X1 U2224 ( .A1(n417), .A2(n275), .ZN(\ab[28][14] ) );
  NOR2_X1 U2225 ( .A1(n420), .A2(n275), .ZN(\ab[28][13] ) );
  NOR2_X1 U2226 ( .A1(n423), .A2(n275), .ZN(\ab[28][12] ) );
  NOR2_X1 U2227 ( .A1(n425), .A2(n275), .ZN(\ab[28][11] ) );
  NOR2_X1 U2228 ( .A1(n477), .A2(n275), .ZN(\ab[28][10] ) );
  NOR2_X1 U2229 ( .A1(n446), .A2(n276), .ZN(\ab[28][0] ) );
  NOR2_X1 U2230 ( .A1(n429), .A2(n279), .ZN(\ab[27][9] ) );
  NOR2_X1 U2231 ( .A1(n431), .A2(n279), .ZN(\ab[27][8] ) );
  NOR2_X1 U2232 ( .A1(n433), .A2(n279), .ZN(\ab[27][7] ) );
  NOR2_X1 U2233 ( .A1(n434), .A2(n279), .ZN(\ab[27][6] ) );
  NOR2_X1 U2234 ( .A1(n436), .A2(n279), .ZN(\ab[27][5] ) );
  NOR2_X1 U2235 ( .A1(n336), .A2(n279), .ZN(\ab[27][52] ) );
  NOR2_X1 U2236 ( .A1(n339), .A2(n279), .ZN(\ab[27][51] ) );
  NOR2_X1 U2237 ( .A1(n341), .A2(n279), .ZN(\ab[27][50] ) );
  NOR2_X1 U2238 ( .A1(n438), .A2(n279), .ZN(\ab[27][4] ) );
  NOR2_X1 U2239 ( .A1(n343), .A2(n279), .ZN(\ab[27][49] ) );
  NOR2_X1 U2240 ( .A1(n345), .A2(n279), .ZN(\ab[27][48] ) );
  NOR2_X1 U2241 ( .A1(n347), .A2(n279), .ZN(\ab[27][47] ) );
  NOR2_X1 U2242 ( .A1(n349), .A2(n279), .ZN(\ab[27][46] ) );
  NOR2_X1 U2243 ( .A1(n351), .A2(n279), .ZN(\ab[27][45] ) );
  NOR2_X1 U2244 ( .A1(n354), .A2(n279), .ZN(\ab[27][44] ) );
  NOR2_X1 U2245 ( .A1(n356), .A2(n279), .ZN(\ab[27][43] ) );
  NOR2_X1 U2246 ( .A1(n359), .A2(n279), .ZN(\ab[27][42] ) );
  NOR2_X1 U2247 ( .A1(n361), .A2(n279), .ZN(\ab[27][41] ) );
  NOR2_X1 U2248 ( .A1(n363), .A2(n279), .ZN(\ab[27][40] ) );
  NOR2_X1 U2249 ( .A1(n440), .A2(n279), .ZN(\ab[27][3] ) );
  NOR2_X1 U2250 ( .A1(n365), .A2(n278), .ZN(\ab[27][39] ) );
  NOR2_X1 U2251 ( .A1(n369), .A2(n278), .ZN(\ab[27][38] ) );
  NOR2_X1 U2252 ( .A1(n370), .A2(n278), .ZN(\ab[27][37] ) );
  NOR2_X1 U2253 ( .A1(n474), .A2(n278), .ZN(\ab[27][36] ) );
  NOR2_X1 U2254 ( .A1(n373), .A2(n278), .ZN(\ab[27][35] ) );
  NOR2_X1 U2255 ( .A1(n375), .A2(n278), .ZN(\ab[27][34] ) );
  NOR2_X1 U2256 ( .A1(n377), .A2(n278), .ZN(\ab[27][33] ) );
  NOR2_X1 U2257 ( .A1(n380), .A2(n278), .ZN(\ab[27][32] ) );
  NOR2_X1 U2258 ( .A1(n381), .A2(n278), .ZN(\ab[27][31] ) );
  NOR2_X1 U2259 ( .A1(n383), .A2(n278), .ZN(\ab[27][30] ) );
  NOR2_X1 U2260 ( .A1(n442), .A2(n278), .ZN(\ab[27][2] ) );
  NOR2_X1 U2261 ( .A1(n386), .A2(n461), .ZN(\ab[27][29] ) );
  NOR2_X1 U2262 ( .A1(n388), .A2(n461), .ZN(\ab[27][28] ) );
  NOR2_X1 U2263 ( .A1(n390), .A2(n461), .ZN(\ab[27][27] ) );
  NOR2_X1 U2264 ( .A1(n392), .A2(n461), .ZN(\ab[27][26] ) );
  NOR2_X1 U2265 ( .A1(n393), .A2(n461), .ZN(\ab[27][25] ) );
  NOR2_X1 U2266 ( .A1(n395), .A2(n461), .ZN(\ab[27][24] ) );
  NOR2_X1 U2267 ( .A1(n397), .A2(n461), .ZN(\ab[27][23] ) );
  NOR2_X1 U2268 ( .A1(n400), .A2(n461), .ZN(\ab[27][22] ) );
  NOR2_X1 U2269 ( .A1(n402), .A2(n461), .ZN(\ab[27][21] ) );
  NOR2_X1 U2270 ( .A1(n403), .A2(n278), .ZN(\ab[27][20] ) );
  NOR2_X1 U2271 ( .A1(n443), .A2(n279), .ZN(\ab[27][1] ) );
  NOR2_X1 U2272 ( .A1(n404), .A2(n278), .ZN(\ab[27][19] ) );
  NOR2_X1 U2273 ( .A1(n476), .A2(n278), .ZN(\ab[27][18] ) );
  NOR2_X1 U2274 ( .A1(n409), .A2(n278), .ZN(\ab[27][17] ) );
  NOR2_X1 U2275 ( .A1(n411), .A2(n279), .ZN(\ab[27][16] ) );
  NOR2_X1 U2276 ( .A1(n414), .A2(n279), .ZN(\ab[27][15] ) );
  NOR2_X1 U2277 ( .A1(n417), .A2(n278), .ZN(\ab[27][14] ) );
  NOR2_X1 U2278 ( .A1(n420), .A2(n278), .ZN(\ab[27][13] ) );
  NOR2_X1 U2279 ( .A1(n423), .A2(n278), .ZN(\ab[27][12] ) );
  NOR2_X1 U2280 ( .A1(n426), .A2(n278), .ZN(\ab[27][11] ) );
  NOR2_X1 U2281 ( .A1(n427), .A2(n278), .ZN(\ab[27][10] ) );
  NOR2_X1 U2282 ( .A1(n446), .A2(n279), .ZN(\ab[27][0] ) );
  NOR2_X1 U2283 ( .A1(n429), .A2(n280), .ZN(\ab[26][9] ) );
  NOR2_X1 U2284 ( .A1(n431), .A2(n280), .ZN(\ab[26][8] ) );
  NOR2_X1 U2285 ( .A1(n433), .A2(n280), .ZN(\ab[26][7] ) );
  NOR2_X1 U2286 ( .A1(n434), .A2(n280), .ZN(\ab[26][6] ) );
  NOR2_X1 U2287 ( .A1(n436), .A2(n280), .ZN(\ab[26][5] ) );
  NOR2_X1 U2288 ( .A1(n336), .A2(n280), .ZN(\ab[26][52] ) );
  NOR2_X1 U2289 ( .A1(n339), .A2(n280), .ZN(\ab[26][51] ) );
  NOR2_X1 U2290 ( .A1(n341), .A2(n280), .ZN(\ab[26][50] ) );
  NOR2_X1 U2291 ( .A1(n438), .A2(n280), .ZN(\ab[26][4] ) );
  NOR2_X1 U2292 ( .A1(n343), .A2(n280), .ZN(\ab[26][49] ) );
  NOR2_X1 U2293 ( .A1(n345), .A2(n280), .ZN(\ab[26][48] ) );
  NOR2_X1 U2294 ( .A1(n347), .A2(n280), .ZN(\ab[26][47] ) );
  NOR2_X1 U2295 ( .A1(n349), .A2(n280), .ZN(\ab[26][46] ) );
  NOR2_X1 U2296 ( .A1(n351), .A2(n280), .ZN(\ab[26][45] ) );
  NOR2_X1 U2297 ( .A1(n354), .A2(n280), .ZN(\ab[26][44] ) );
  NOR2_X1 U2298 ( .A1(n356), .A2(n280), .ZN(\ab[26][43] ) );
  NOR2_X1 U2299 ( .A1(n359), .A2(n280), .ZN(\ab[26][42] ) );
  NOR2_X1 U2300 ( .A1(n361), .A2(n280), .ZN(\ab[26][41] ) );
  NOR2_X1 U2301 ( .A1(n363), .A2(n280), .ZN(\ab[26][40] ) );
  NOR2_X1 U2302 ( .A1(n440), .A2(n280), .ZN(\ab[26][3] ) );
  NOR2_X1 U2303 ( .A1(n365), .A2(n281), .ZN(\ab[26][39] ) );
  NOR2_X1 U2304 ( .A1(n369), .A2(n281), .ZN(\ab[26][38] ) );
  NOR2_X1 U2305 ( .A1(n370), .A2(n281), .ZN(\ab[26][37] ) );
  NOR2_X1 U2306 ( .A1(n372), .A2(n281), .ZN(\ab[26][36] ) );
  NOR2_X1 U2307 ( .A1(n373), .A2(n281), .ZN(\ab[26][35] ) );
  NOR2_X1 U2308 ( .A1(n375), .A2(n281), .ZN(\ab[26][34] ) );
  NOR2_X1 U2309 ( .A1(n377), .A2(n281), .ZN(\ab[26][33] ) );
  NOR2_X1 U2310 ( .A1(n379), .A2(n281), .ZN(\ab[26][32] ) );
  NOR2_X1 U2311 ( .A1(n381), .A2(n281), .ZN(\ab[26][31] ) );
  NOR2_X1 U2312 ( .A1(n383), .A2(n281), .ZN(\ab[26][30] ) );
  NOR2_X1 U2313 ( .A1(n442), .A2(n281), .ZN(\ab[26][2] ) );
  NOR2_X1 U2314 ( .A1(n385), .A2(n281), .ZN(\ab[26][29] ) );
  NOR2_X1 U2315 ( .A1(n388), .A2(n281), .ZN(\ab[26][28] ) );
  NOR2_X1 U2316 ( .A1(n389), .A2(n281), .ZN(\ab[26][27] ) );
  NOR2_X1 U2317 ( .A1(n391), .A2(n281), .ZN(\ab[26][26] ) );
  NOR2_X1 U2318 ( .A1(n394), .A2(n281), .ZN(\ab[26][25] ) );
  NOR2_X1 U2319 ( .A1(n396), .A2(n281), .ZN(\ab[26][24] ) );
  NOR2_X1 U2320 ( .A1(n398), .A2(n281), .ZN(\ab[26][23] ) );
  NOR2_X1 U2321 ( .A1(n399), .A2(n281), .ZN(\ab[26][22] ) );
  NOR2_X1 U2322 ( .A1(n401), .A2(n281), .ZN(\ab[26][21] ) );
  NOR2_X1 U2323 ( .A1(n403), .A2(n281), .ZN(\ab[26][20] ) );
  NOR2_X1 U2324 ( .A1(n443), .A2(n281), .ZN(\ab[26][1] ) );
  NOR2_X1 U2325 ( .A1(n404), .A2(n280), .ZN(\ab[26][19] ) );
  NOR2_X1 U2326 ( .A1(n476), .A2(n280), .ZN(\ab[26][18] ) );
  NOR2_X1 U2327 ( .A1(n408), .A2(n280), .ZN(\ab[26][17] ) );
  NOR2_X1 U2328 ( .A1(n411), .A2(n280), .ZN(\ab[26][16] ) );
  NOR2_X1 U2329 ( .A1(n414), .A2(n280), .ZN(\ab[26][15] ) );
  NOR2_X1 U2330 ( .A1(n417), .A2(n280), .ZN(\ab[26][14] ) );
  NOR2_X1 U2331 ( .A1(n420), .A2(n280), .ZN(\ab[26][13] ) );
  NOR2_X1 U2332 ( .A1(n423), .A2(n280), .ZN(\ab[26][12] ) );
  NOR2_X1 U2333 ( .A1(n425), .A2(n280), .ZN(\ab[26][11] ) );
  NOR2_X1 U2334 ( .A1(n477), .A2(n280), .ZN(\ab[26][10] ) );
  NOR2_X1 U2335 ( .A1(n446), .A2(n280), .ZN(\ab[26][0] ) );
  NOR2_X1 U2336 ( .A1(n429), .A2(n283), .ZN(\ab[25][9] ) );
  NOR2_X1 U2337 ( .A1(n431), .A2(n283), .ZN(\ab[25][8] ) );
  NOR2_X1 U2338 ( .A1(n433), .A2(n283), .ZN(\ab[25][7] ) );
  NOR2_X1 U2339 ( .A1(n434), .A2(n283), .ZN(\ab[25][6] ) );
  NOR2_X1 U2340 ( .A1(n436), .A2(n283), .ZN(\ab[25][5] ) );
  NOR2_X1 U2341 ( .A1(n336), .A2(n283), .ZN(\ab[25][52] ) );
  NOR2_X1 U2342 ( .A1(n339), .A2(n283), .ZN(\ab[25][51] ) );
  NOR2_X1 U2343 ( .A1(n341), .A2(n283), .ZN(\ab[25][50] ) );
  NOR2_X1 U2344 ( .A1(n438), .A2(n283), .ZN(\ab[25][4] ) );
  NOR2_X1 U2345 ( .A1(n343), .A2(n283), .ZN(\ab[25][49] ) );
  NOR2_X1 U2346 ( .A1(n345), .A2(n283), .ZN(\ab[25][48] ) );
  NOR2_X1 U2347 ( .A1(n347), .A2(n283), .ZN(\ab[25][47] ) );
  NOR2_X1 U2348 ( .A1(n349), .A2(n283), .ZN(\ab[25][46] ) );
  NOR2_X1 U2349 ( .A1(n351), .A2(n283), .ZN(\ab[25][45] ) );
  NOR2_X1 U2350 ( .A1(n354), .A2(n283), .ZN(\ab[25][44] ) );
  NOR2_X1 U2351 ( .A1(n356), .A2(n283), .ZN(\ab[25][43] ) );
  NOR2_X1 U2352 ( .A1(n359), .A2(n283), .ZN(\ab[25][42] ) );
  NOR2_X1 U2353 ( .A1(n361), .A2(n283), .ZN(\ab[25][41] ) );
  NOR2_X1 U2354 ( .A1(n363), .A2(n283), .ZN(\ab[25][40] ) );
  NOR2_X1 U2355 ( .A1(n440), .A2(n283), .ZN(\ab[25][3] ) );
  NOR2_X1 U2356 ( .A1(n365), .A2(n282), .ZN(\ab[25][39] ) );
  NOR2_X1 U2357 ( .A1(n369), .A2(n282), .ZN(\ab[25][38] ) );
  NOR2_X1 U2358 ( .A1(n370), .A2(n282), .ZN(\ab[25][37] ) );
  NOR2_X1 U2359 ( .A1(n474), .A2(n282), .ZN(\ab[25][36] ) );
  NOR2_X1 U2360 ( .A1(n373), .A2(n282), .ZN(\ab[25][35] ) );
  NOR2_X1 U2361 ( .A1(n375), .A2(n282), .ZN(\ab[25][34] ) );
  NOR2_X1 U2362 ( .A1(n377), .A2(n282), .ZN(\ab[25][33] ) );
  NOR2_X1 U2363 ( .A1(n380), .A2(n282), .ZN(\ab[25][32] ) );
  NOR2_X1 U2364 ( .A1(n381), .A2(n282), .ZN(\ab[25][31] ) );
  NOR2_X1 U2365 ( .A1(n383), .A2(n282), .ZN(\ab[25][30] ) );
  NOR2_X1 U2366 ( .A1(n442), .A2(n282), .ZN(\ab[25][2] ) );
  NOR2_X1 U2367 ( .A1(n386), .A2(n462), .ZN(\ab[25][29] ) );
  NOR2_X1 U2368 ( .A1(n388), .A2(n462), .ZN(\ab[25][28] ) );
  NOR2_X1 U2369 ( .A1(n390), .A2(n282), .ZN(\ab[25][27] ) );
  NOR2_X1 U2370 ( .A1(n392), .A2(n282), .ZN(\ab[25][26] ) );
  NOR2_X1 U2371 ( .A1(n393), .A2(n462), .ZN(\ab[25][25] ) );
  NOR2_X1 U2372 ( .A1(n395), .A2(n462), .ZN(\ab[25][24] ) );
  NOR2_X1 U2373 ( .A1(n397), .A2(n462), .ZN(\ab[25][23] ) );
  NOR2_X1 U2374 ( .A1(n400), .A2(n462), .ZN(\ab[25][22] ) );
  NOR2_X1 U2375 ( .A1(n402), .A2(n283), .ZN(\ab[25][21] ) );
  NOR2_X1 U2376 ( .A1(n403), .A2(n283), .ZN(\ab[25][20] ) );
  NOR2_X1 U2377 ( .A1(n443), .A2(n283), .ZN(\ab[25][1] ) );
  NOR2_X1 U2378 ( .A1(n404), .A2(n283), .ZN(\ab[25][19] ) );
  NOR2_X1 U2379 ( .A1(n407), .A2(n283), .ZN(\ab[25][18] ) );
  NOR2_X1 U2380 ( .A1(n408), .A2(n283), .ZN(\ab[25][17] ) );
  NOR2_X1 U2381 ( .A1(n411), .A2(n283), .ZN(\ab[25][16] ) );
  NOR2_X1 U2382 ( .A1(n414), .A2(n283), .ZN(\ab[25][15] ) );
  NOR2_X1 U2383 ( .A1(n417), .A2(n283), .ZN(\ab[25][14] ) );
  NOR2_X1 U2384 ( .A1(n420), .A2(n283), .ZN(\ab[25][13] ) );
  NOR2_X1 U2385 ( .A1(n423), .A2(n283), .ZN(\ab[25][12] ) );
  NOR2_X1 U2386 ( .A1(n425), .A2(n283), .ZN(\ab[25][11] ) );
  NOR2_X1 U2387 ( .A1(n427), .A2(n283), .ZN(\ab[25][10] ) );
  NOR2_X1 U2388 ( .A1(n446), .A2(n283), .ZN(\ab[25][0] ) );
  NOR2_X1 U2389 ( .A1(n429), .A2(n285), .ZN(\ab[24][9] ) );
  NOR2_X1 U2390 ( .A1(n431), .A2(n285), .ZN(\ab[24][8] ) );
  NOR2_X1 U2391 ( .A1(n433), .A2(n285), .ZN(\ab[24][7] ) );
  NOR2_X1 U2392 ( .A1(n434), .A2(n285), .ZN(\ab[24][6] ) );
  NOR2_X1 U2393 ( .A1(n436), .A2(n285), .ZN(\ab[24][5] ) );
  NOR2_X1 U2394 ( .A1(n336), .A2(n285), .ZN(\ab[24][52] ) );
  NOR2_X1 U2395 ( .A1(n339), .A2(n285), .ZN(\ab[24][51] ) );
  NOR2_X1 U2396 ( .A1(n341), .A2(n285), .ZN(\ab[24][50] ) );
  NOR2_X1 U2397 ( .A1(n438), .A2(n285), .ZN(\ab[24][4] ) );
  NOR2_X1 U2398 ( .A1(n343), .A2(n285), .ZN(\ab[24][49] ) );
  NOR2_X1 U2399 ( .A1(n345), .A2(n285), .ZN(\ab[24][48] ) );
  NOR2_X1 U2400 ( .A1(n347), .A2(n285), .ZN(\ab[24][47] ) );
  NOR2_X1 U2401 ( .A1(n349), .A2(n285), .ZN(\ab[24][46] ) );
  NOR2_X1 U2402 ( .A1(n351), .A2(n285), .ZN(\ab[24][45] ) );
  NOR2_X1 U2403 ( .A1(n354), .A2(n285), .ZN(\ab[24][44] ) );
  NOR2_X1 U2404 ( .A1(n356), .A2(n285), .ZN(\ab[24][43] ) );
  NOR2_X1 U2405 ( .A1(n359), .A2(n285), .ZN(\ab[24][42] ) );
  NOR2_X1 U2406 ( .A1(n361), .A2(n285), .ZN(\ab[24][41] ) );
  NOR2_X1 U2407 ( .A1(n363), .A2(n285), .ZN(\ab[24][40] ) );
  NOR2_X1 U2408 ( .A1(n440), .A2(n285), .ZN(\ab[24][3] ) );
  NOR2_X1 U2409 ( .A1(n365), .A2(n284), .ZN(\ab[24][39] ) );
  NOR2_X1 U2410 ( .A1(n369), .A2(n284), .ZN(\ab[24][38] ) );
  NOR2_X1 U2411 ( .A1(n370), .A2(n284), .ZN(\ab[24][37] ) );
  NOR2_X1 U2412 ( .A1(n372), .A2(n284), .ZN(\ab[24][36] ) );
  NOR2_X1 U2413 ( .A1(n373), .A2(n284), .ZN(\ab[24][35] ) );
  NOR2_X1 U2414 ( .A1(n375), .A2(n284), .ZN(\ab[24][34] ) );
  NOR2_X1 U2415 ( .A1(n377), .A2(n284), .ZN(\ab[24][33] ) );
  NOR2_X1 U2416 ( .A1(n379), .A2(n284), .ZN(\ab[24][32] ) );
  NOR2_X1 U2417 ( .A1(n381), .A2(n284), .ZN(\ab[24][31] ) );
  NOR2_X1 U2418 ( .A1(n383), .A2(n284), .ZN(\ab[24][30] ) );
  NOR2_X1 U2419 ( .A1(n442), .A2(n284), .ZN(\ab[24][2] ) );
  NOR2_X1 U2420 ( .A1(n385), .A2(n284), .ZN(\ab[24][29] ) );
  NOR2_X1 U2421 ( .A1(n388), .A2(n284), .ZN(\ab[24][28] ) );
  NOR2_X1 U2422 ( .A1(n389), .A2(n284), .ZN(\ab[24][27] ) );
  NOR2_X1 U2423 ( .A1(n391), .A2(n284), .ZN(\ab[24][26] ) );
  NOR2_X1 U2424 ( .A1(n393), .A2(n284), .ZN(\ab[24][25] ) );
  NOR2_X1 U2425 ( .A1(n395), .A2(n284), .ZN(\ab[24][24] ) );
  NOR2_X1 U2426 ( .A1(n397), .A2(n285), .ZN(\ab[24][23] ) );
  NOR2_X1 U2427 ( .A1(n399), .A2(n285), .ZN(\ab[24][22] ) );
  NOR2_X1 U2428 ( .A1(n401), .A2(n285), .ZN(\ab[24][21] ) );
  NOR2_X1 U2429 ( .A1(n403), .A2(n285), .ZN(\ab[24][20] ) );
  NOR2_X1 U2430 ( .A1(n443), .A2(n285), .ZN(\ab[24][1] ) );
  NOR2_X1 U2431 ( .A1(n404), .A2(n285), .ZN(\ab[24][19] ) );
  NOR2_X1 U2432 ( .A1(n406), .A2(n285), .ZN(\ab[24][18] ) );
  NOR2_X1 U2433 ( .A1(n408), .A2(n285), .ZN(\ab[24][17] ) );
  NOR2_X1 U2434 ( .A1(n411), .A2(n285), .ZN(\ab[24][16] ) );
  NOR2_X1 U2435 ( .A1(n414), .A2(n285), .ZN(\ab[24][15] ) );
  NOR2_X1 U2436 ( .A1(n417), .A2(n285), .ZN(\ab[24][14] ) );
  NOR2_X1 U2437 ( .A1(n420), .A2(n285), .ZN(\ab[24][13] ) );
  NOR2_X1 U2438 ( .A1(n423), .A2(n285), .ZN(\ab[24][12] ) );
  NOR2_X1 U2439 ( .A1(n425), .A2(n285), .ZN(\ab[24][11] ) );
  NOR2_X1 U2440 ( .A1(n477), .A2(n285), .ZN(\ab[24][10] ) );
  NOR2_X1 U2441 ( .A1(n446), .A2(n285), .ZN(\ab[24][0] ) );
  NOR2_X1 U2442 ( .A1(n429), .A2(n287), .ZN(\ab[23][9] ) );
  NOR2_X1 U2443 ( .A1(n431), .A2(n287), .ZN(\ab[23][8] ) );
  NOR2_X1 U2444 ( .A1(n433), .A2(n287), .ZN(\ab[23][7] ) );
  NOR2_X1 U2445 ( .A1(n434), .A2(n287), .ZN(\ab[23][6] ) );
  NOR2_X1 U2446 ( .A1(n436), .A2(n287), .ZN(\ab[23][5] ) );
  NOR2_X1 U2447 ( .A1(n336), .A2(n287), .ZN(\ab[23][52] ) );
  NOR2_X1 U2448 ( .A1(n339), .A2(n287), .ZN(\ab[23][51] ) );
  NOR2_X1 U2449 ( .A1(n341), .A2(n287), .ZN(\ab[23][50] ) );
  NOR2_X1 U2450 ( .A1(n438), .A2(n287), .ZN(\ab[23][4] ) );
  NOR2_X1 U2451 ( .A1(n343), .A2(n287), .ZN(\ab[23][49] ) );
  NOR2_X1 U2452 ( .A1(n345), .A2(n287), .ZN(\ab[23][48] ) );
  NOR2_X1 U2453 ( .A1(n347), .A2(n287), .ZN(\ab[23][47] ) );
  NOR2_X1 U2454 ( .A1(n349), .A2(n287), .ZN(\ab[23][46] ) );
  NOR2_X1 U2455 ( .A1(n351), .A2(n287), .ZN(\ab[23][45] ) );
  NOR2_X1 U2456 ( .A1(n354), .A2(n287), .ZN(\ab[23][44] ) );
  NOR2_X1 U2457 ( .A1(n356), .A2(n287), .ZN(\ab[23][43] ) );
  NOR2_X1 U2458 ( .A1(n359), .A2(n287), .ZN(\ab[23][42] ) );
  NOR2_X1 U2459 ( .A1(n361), .A2(n287), .ZN(\ab[23][41] ) );
  NOR2_X1 U2460 ( .A1(n363), .A2(n287), .ZN(\ab[23][40] ) );
  NOR2_X1 U2461 ( .A1(n440), .A2(n287), .ZN(\ab[23][3] ) );
  NOR2_X1 U2462 ( .A1(n365), .A2(n286), .ZN(\ab[23][39] ) );
  NOR2_X1 U2463 ( .A1(n369), .A2(n286), .ZN(\ab[23][38] ) );
  NOR2_X1 U2464 ( .A1(n370), .A2(n286), .ZN(\ab[23][37] ) );
  NOR2_X1 U2465 ( .A1(n474), .A2(n286), .ZN(\ab[23][36] ) );
  NOR2_X1 U2466 ( .A1(n373), .A2(n286), .ZN(\ab[23][35] ) );
  NOR2_X1 U2467 ( .A1(n375), .A2(n286), .ZN(\ab[23][34] ) );
  NOR2_X1 U2468 ( .A1(n377), .A2(n286), .ZN(\ab[23][33] ) );
  NOR2_X1 U2469 ( .A1(n380), .A2(n286), .ZN(\ab[23][32] ) );
  NOR2_X1 U2470 ( .A1(n381), .A2(n286), .ZN(\ab[23][31] ) );
  NOR2_X1 U2471 ( .A1(n383), .A2(n286), .ZN(\ab[23][30] ) );
  NOR2_X1 U2472 ( .A1(n442), .A2(n286), .ZN(\ab[23][2] ) );
  NOR2_X1 U2473 ( .A1(n386), .A2(n286), .ZN(\ab[23][29] ) );
  NOR2_X1 U2474 ( .A1(n388), .A2(n286), .ZN(\ab[23][28] ) );
  NOR2_X1 U2475 ( .A1(n390), .A2(n286), .ZN(\ab[23][27] ) );
  NOR2_X1 U2476 ( .A1(n392), .A2(n286), .ZN(\ab[23][26] ) );
  NOR2_X1 U2477 ( .A1(n394), .A2(n287), .ZN(\ab[23][25] ) );
  NOR2_X1 U2478 ( .A1(n396), .A2(n287), .ZN(\ab[23][24] ) );
  NOR2_X1 U2479 ( .A1(n398), .A2(n287), .ZN(\ab[23][23] ) );
  NOR2_X1 U2480 ( .A1(n400), .A2(n286), .ZN(\ab[23][22] ) );
  NOR2_X1 U2481 ( .A1(n402), .A2(n286), .ZN(\ab[23][21] ) );
  NOR2_X1 U2482 ( .A1(n403), .A2(n287), .ZN(\ab[23][20] ) );
  NOR2_X1 U2483 ( .A1(n443), .A2(n286), .ZN(\ab[23][1] ) );
  NOR2_X1 U2484 ( .A1(n404), .A2(n287), .ZN(\ab[23][19] ) );
  NOR2_X1 U2485 ( .A1(n406), .A2(n287), .ZN(\ab[23][18] ) );
  NOR2_X1 U2486 ( .A1(n408), .A2(n287), .ZN(\ab[23][17] ) );
  NOR2_X1 U2487 ( .A1(n411), .A2(n287), .ZN(\ab[23][16] ) );
  NOR2_X1 U2488 ( .A1(n414), .A2(n287), .ZN(\ab[23][15] ) );
  NOR2_X1 U2489 ( .A1(n417), .A2(n287), .ZN(\ab[23][14] ) );
  NOR2_X1 U2490 ( .A1(n420), .A2(n287), .ZN(\ab[23][13] ) );
  NOR2_X1 U2491 ( .A1(n423), .A2(n287), .ZN(\ab[23][12] ) );
  NOR2_X1 U2492 ( .A1(n425), .A2(n287), .ZN(\ab[23][11] ) );
  NOR2_X1 U2493 ( .A1(n427), .A2(n287), .ZN(\ab[23][10] ) );
  NOR2_X1 U2494 ( .A1(n446), .A2(n287), .ZN(\ab[23][0] ) );
  NOR2_X1 U2495 ( .A1(n429), .A2(n289), .ZN(\ab[22][9] ) );
  NOR2_X1 U2496 ( .A1(n431), .A2(n289), .ZN(\ab[22][8] ) );
  NOR2_X1 U2497 ( .A1(n433), .A2(n289), .ZN(\ab[22][7] ) );
  NOR2_X1 U2498 ( .A1(n434), .A2(n289), .ZN(\ab[22][6] ) );
  NOR2_X1 U2499 ( .A1(n436), .A2(n289), .ZN(\ab[22][5] ) );
  NOR2_X1 U2500 ( .A1(n336), .A2(n289), .ZN(\ab[22][52] ) );
  NOR2_X1 U2501 ( .A1(n339), .A2(n289), .ZN(\ab[22][51] ) );
  NOR2_X1 U2502 ( .A1(n341), .A2(n289), .ZN(\ab[22][50] ) );
  NOR2_X1 U2503 ( .A1(n438), .A2(n289), .ZN(\ab[22][4] ) );
  NOR2_X1 U2504 ( .A1(n343), .A2(n289), .ZN(\ab[22][49] ) );
  NOR2_X1 U2505 ( .A1(n345), .A2(n289), .ZN(\ab[22][48] ) );
  NOR2_X1 U2506 ( .A1(n347), .A2(n289), .ZN(\ab[22][47] ) );
  NOR2_X1 U2507 ( .A1(n349), .A2(n289), .ZN(\ab[22][46] ) );
  NOR2_X1 U2508 ( .A1(n351), .A2(n289), .ZN(\ab[22][45] ) );
  NOR2_X1 U2509 ( .A1(n354), .A2(n289), .ZN(\ab[22][44] ) );
  NOR2_X1 U2510 ( .A1(n356), .A2(n289), .ZN(\ab[22][43] ) );
  NOR2_X1 U2511 ( .A1(n359), .A2(n289), .ZN(\ab[22][42] ) );
  NOR2_X1 U2512 ( .A1(n361), .A2(n289), .ZN(\ab[22][41] ) );
  NOR2_X1 U2513 ( .A1(n363), .A2(n289), .ZN(\ab[22][40] ) );
  NOR2_X1 U2514 ( .A1(n440), .A2(n289), .ZN(\ab[22][3] ) );
  NOR2_X1 U2515 ( .A1(n365), .A2(n288), .ZN(\ab[22][39] ) );
  NOR2_X1 U2516 ( .A1(n369), .A2(n288), .ZN(\ab[22][38] ) );
  NOR2_X1 U2517 ( .A1(n370), .A2(n288), .ZN(\ab[22][37] ) );
  NOR2_X1 U2518 ( .A1(n372), .A2(n288), .ZN(\ab[22][36] ) );
  NOR2_X1 U2519 ( .A1(n373), .A2(n288), .ZN(\ab[22][35] ) );
  NOR2_X1 U2520 ( .A1(n375), .A2(n288), .ZN(\ab[22][34] ) );
  NOR2_X1 U2521 ( .A1(n377), .A2(n288), .ZN(\ab[22][33] ) );
  NOR2_X1 U2522 ( .A1(n379), .A2(n288), .ZN(\ab[22][32] ) );
  NOR2_X1 U2523 ( .A1(n381), .A2(n288), .ZN(\ab[22][31] ) );
  NOR2_X1 U2524 ( .A1(n383), .A2(n288), .ZN(\ab[22][30] ) );
  NOR2_X1 U2525 ( .A1(n442), .A2(n288), .ZN(\ab[22][2] ) );
  NOR2_X1 U2526 ( .A1(n386), .A2(n288), .ZN(\ab[22][29] ) );
  NOR2_X1 U2527 ( .A1(n388), .A2(n288), .ZN(\ab[22][28] ) );
  NOR2_X1 U2528 ( .A1(n390), .A2(n288), .ZN(\ab[22][27] ) );
  NOR2_X1 U2529 ( .A1(n392), .A2(n288), .ZN(\ab[22][26] ) );
  NOR2_X1 U2530 ( .A1(n394), .A2(n289), .ZN(\ab[22][25] ) );
  NOR2_X1 U2531 ( .A1(n396), .A2(n289), .ZN(\ab[22][24] ) );
  NOR2_X1 U2532 ( .A1(n398), .A2(n289), .ZN(\ab[22][23] ) );
  NOR2_X1 U2533 ( .A1(n400), .A2(n289), .ZN(\ab[22][22] ) );
  NOR2_X1 U2534 ( .A1(n402), .A2(n289), .ZN(\ab[22][21] ) );
  NOR2_X1 U2535 ( .A1(n475), .A2(n289), .ZN(\ab[22][20] ) );
  NOR2_X1 U2536 ( .A1(n443), .A2(n289), .ZN(\ab[22][1] ) );
  NOR2_X1 U2537 ( .A1(n404), .A2(n289), .ZN(\ab[22][19] ) );
  NOR2_X1 U2538 ( .A1(n406), .A2(n289), .ZN(\ab[22][18] ) );
  NOR2_X1 U2539 ( .A1(n408), .A2(n289), .ZN(\ab[22][17] ) );
  NOR2_X1 U2540 ( .A1(n411), .A2(n289), .ZN(\ab[22][16] ) );
  NOR2_X1 U2541 ( .A1(n414), .A2(n289), .ZN(\ab[22][15] ) );
  NOR2_X1 U2542 ( .A1(n417), .A2(n289), .ZN(\ab[22][14] ) );
  NOR2_X1 U2543 ( .A1(n420), .A2(n289), .ZN(\ab[22][13] ) );
  NOR2_X1 U2544 ( .A1(n423), .A2(n289), .ZN(\ab[22][12] ) );
  NOR2_X1 U2545 ( .A1(n425), .A2(n289), .ZN(\ab[22][11] ) );
  NOR2_X1 U2546 ( .A1(n477), .A2(n289), .ZN(\ab[22][10] ) );
  NOR2_X1 U2547 ( .A1(n446), .A2(n289), .ZN(\ab[22][0] ) );
  NOR2_X1 U2548 ( .A1(n429), .A2(n291), .ZN(\ab[21][9] ) );
  NOR2_X1 U2549 ( .A1(n431), .A2(n291), .ZN(\ab[21][8] ) );
  NOR2_X1 U2550 ( .A1(n433), .A2(n291), .ZN(\ab[21][7] ) );
  NOR2_X1 U2551 ( .A1(n434), .A2(n291), .ZN(\ab[21][6] ) );
  NOR2_X1 U2552 ( .A1(n436), .A2(n291), .ZN(\ab[21][5] ) );
  NOR2_X1 U2553 ( .A1(n336), .A2(n291), .ZN(\ab[21][52] ) );
  NOR2_X1 U2554 ( .A1(n339), .A2(n291), .ZN(\ab[21][51] ) );
  NOR2_X1 U2555 ( .A1(n341), .A2(n291), .ZN(\ab[21][50] ) );
  NOR2_X1 U2556 ( .A1(n438), .A2(n291), .ZN(\ab[21][4] ) );
  NOR2_X1 U2557 ( .A1(n343), .A2(n291), .ZN(\ab[21][49] ) );
  NOR2_X1 U2558 ( .A1(n345), .A2(n291), .ZN(\ab[21][48] ) );
  NOR2_X1 U2559 ( .A1(n347), .A2(n291), .ZN(\ab[21][47] ) );
  NOR2_X1 U2560 ( .A1(n349), .A2(n291), .ZN(\ab[21][46] ) );
  NOR2_X1 U2561 ( .A1(n351), .A2(n291), .ZN(\ab[21][45] ) );
  NOR2_X1 U2562 ( .A1(n354), .A2(n291), .ZN(\ab[21][44] ) );
  NOR2_X1 U2563 ( .A1(n356), .A2(n291), .ZN(\ab[21][43] ) );
  NOR2_X1 U2564 ( .A1(n359), .A2(n291), .ZN(\ab[21][42] ) );
  NOR2_X1 U2565 ( .A1(n361), .A2(n291), .ZN(\ab[21][41] ) );
  NOR2_X1 U2566 ( .A1(n363), .A2(n291), .ZN(\ab[21][40] ) );
  NOR2_X1 U2567 ( .A1(n440), .A2(n291), .ZN(\ab[21][3] ) );
  NOR2_X1 U2568 ( .A1(n365), .A2(n290), .ZN(\ab[21][39] ) );
  NOR2_X1 U2569 ( .A1(n368), .A2(n290), .ZN(\ab[21][38] ) );
  NOR2_X1 U2570 ( .A1(n370), .A2(n290), .ZN(\ab[21][37] ) );
  NOR2_X1 U2571 ( .A1(n474), .A2(n290), .ZN(\ab[21][36] ) );
  NOR2_X1 U2572 ( .A1(n373), .A2(n290), .ZN(\ab[21][35] ) );
  NOR2_X1 U2573 ( .A1(n375), .A2(n290), .ZN(\ab[21][34] ) );
  NOR2_X1 U2574 ( .A1(n377), .A2(n290), .ZN(\ab[21][33] ) );
  NOR2_X1 U2575 ( .A1(n380), .A2(n290), .ZN(\ab[21][32] ) );
  NOR2_X1 U2576 ( .A1(n381), .A2(n290), .ZN(\ab[21][31] ) );
  NOR2_X1 U2577 ( .A1(n383), .A2(n290), .ZN(\ab[21][30] ) );
  NOR2_X1 U2578 ( .A1(n442), .A2(n290), .ZN(\ab[21][2] ) );
  NOR2_X1 U2579 ( .A1(n385), .A2(n290), .ZN(\ab[21][29] ) );
  NOR2_X1 U2580 ( .A1(n388), .A2(n290), .ZN(\ab[21][28] ) );
  NOR2_X1 U2581 ( .A1(n389), .A2(n291), .ZN(\ab[21][27] ) );
  NOR2_X1 U2582 ( .A1(n391), .A2(n290), .ZN(\ab[21][26] ) );
  NOR2_X1 U2583 ( .A1(n393), .A2(n290), .ZN(\ab[21][25] ) );
  NOR2_X1 U2584 ( .A1(n395), .A2(n290), .ZN(\ab[21][24] ) );
  NOR2_X1 U2585 ( .A1(n397), .A2(n290), .ZN(\ab[21][23] ) );
  NOR2_X1 U2586 ( .A1(n399), .A2(n291), .ZN(\ab[21][22] ) );
  NOR2_X1 U2587 ( .A1(n401), .A2(n463), .ZN(\ab[21][21] ) );
  NOR2_X1 U2588 ( .A1(n403), .A2(n463), .ZN(\ab[21][20] ) );
  NOR2_X1 U2589 ( .A1(n443), .A2(n463), .ZN(\ab[21][1] ) );
  NOR2_X1 U2590 ( .A1(n404), .A2(n291), .ZN(\ab[21][19] ) );
  NOR2_X1 U2591 ( .A1(n406), .A2(n291), .ZN(\ab[21][18] ) );
  NOR2_X1 U2592 ( .A1(n408), .A2(n291), .ZN(\ab[21][17] ) );
  NOR2_X1 U2593 ( .A1(n411), .A2(n291), .ZN(\ab[21][16] ) );
  NOR2_X1 U2594 ( .A1(n414), .A2(n291), .ZN(\ab[21][15] ) );
  NOR2_X1 U2595 ( .A1(n417), .A2(n291), .ZN(\ab[21][14] ) );
  NOR2_X1 U2596 ( .A1(n420), .A2(n291), .ZN(\ab[21][13] ) );
  NOR2_X1 U2597 ( .A1(n423), .A2(n291), .ZN(\ab[21][12] ) );
  NOR2_X1 U2598 ( .A1(n425), .A2(n291), .ZN(\ab[21][11] ) );
  NOR2_X1 U2599 ( .A1(n427), .A2(n291), .ZN(\ab[21][10] ) );
  NOR2_X1 U2600 ( .A1(n446), .A2(n291), .ZN(\ab[21][0] ) );
  NOR2_X1 U2601 ( .A1(n429), .A2(n292), .ZN(\ab[20][9] ) );
  NOR2_X1 U2602 ( .A1(n431), .A2(n292), .ZN(\ab[20][8] ) );
  NOR2_X1 U2603 ( .A1(n433), .A2(n292), .ZN(\ab[20][7] ) );
  NOR2_X1 U2604 ( .A1(n434), .A2(n292), .ZN(\ab[20][6] ) );
  NOR2_X1 U2605 ( .A1(n436), .A2(n292), .ZN(\ab[20][5] ) );
  NOR2_X1 U2606 ( .A1(n336), .A2(n292), .ZN(\ab[20][52] ) );
  NOR2_X1 U2607 ( .A1(n339), .A2(n292), .ZN(\ab[20][51] ) );
  NOR2_X1 U2608 ( .A1(n341), .A2(n292), .ZN(\ab[20][50] ) );
  NOR2_X1 U2609 ( .A1(n438), .A2(n292), .ZN(\ab[20][4] ) );
  NOR2_X1 U2610 ( .A1(n343), .A2(n292), .ZN(\ab[20][49] ) );
  NOR2_X1 U2611 ( .A1(n345), .A2(n292), .ZN(\ab[20][48] ) );
  NOR2_X1 U2612 ( .A1(n347), .A2(n292), .ZN(\ab[20][47] ) );
  NOR2_X1 U2613 ( .A1(n349), .A2(n292), .ZN(\ab[20][46] ) );
  NOR2_X1 U2614 ( .A1(n351), .A2(n292), .ZN(\ab[20][45] ) );
  NOR2_X1 U2615 ( .A1(n354), .A2(n292), .ZN(\ab[20][44] ) );
  NOR2_X1 U2616 ( .A1(n356), .A2(n292), .ZN(\ab[20][43] ) );
  NOR2_X1 U2617 ( .A1(n359), .A2(n292), .ZN(\ab[20][42] ) );
  NOR2_X1 U2618 ( .A1(n361), .A2(n292), .ZN(\ab[20][41] ) );
  NOR2_X1 U2619 ( .A1(n363), .A2(n292), .ZN(\ab[20][40] ) );
  NOR2_X1 U2620 ( .A1(n440), .A2(n292), .ZN(\ab[20][3] ) );
  NOR2_X1 U2621 ( .A1(n365), .A2(n464), .ZN(\ab[20][39] ) );
  NOR2_X1 U2622 ( .A1(n368), .A2(n464), .ZN(\ab[20][38] ) );
  NOR2_X1 U2623 ( .A1(n370), .A2(n464), .ZN(\ab[20][37] ) );
  NOR2_X1 U2624 ( .A1(n372), .A2(n464), .ZN(\ab[20][36] ) );
  NOR2_X1 U2625 ( .A1(n373), .A2(n464), .ZN(\ab[20][35] ) );
  NOR2_X1 U2626 ( .A1(n375), .A2(n464), .ZN(\ab[20][34] ) );
  NOR2_X1 U2627 ( .A1(n377), .A2(n464), .ZN(\ab[20][33] ) );
  NOR2_X1 U2628 ( .A1(n379), .A2(n464), .ZN(\ab[20][32] ) );
  NOR2_X1 U2629 ( .A1(n381), .A2(n464), .ZN(\ab[20][31] ) );
  NOR2_X1 U2630 ( .A1(n383), .A2(n464), .ZN(\ab[20][30] ) );
  NOR2_X1 U2631 ( .A1(n442), .A2(n464), .ZN(\ab[20][2] ) );
  NOR2_X1 U2632 ( .A1(n386), .A2(n292), .ZN(\ab[20][29] ) );
  NOR2_X1 U2633 ( .A1(n388), .A2(n292), .ZN(\ab[20][28] ) );
  NOR2_X1 U2634 ( .A1(n390), .A2(n292), .ZN(\ab[20][27] ) );
  NOR2_X1 U2635 ( .A1(n392), .A2(n292), .ZN(\ab[20][26] ) );
  NOR2_X1 U2636 ( .A1(n394), .A2(n292), .ZN(\ab[20][25] ) );
  NOR2_X1 U2637 ( .A1(n396), .A2(n292), .ZN(\ab[20][24] ) );
  NOR2_X1 U2638 ( .A1(n398), .A2(n292), .ZN(\ab[20][23] ) );
  NOR2_X1 U2639 ( .A1(n400), .A2(n292), .ZN(\ab[20][22] ) );
  NOR2_X1 U2640 ( .A1(n402), .A2(n292), .ZN(\ab[20][21] ) );
  NOR2_X1 U2641 ( .A1(n403), .A2(n292), .ZN(\ab[20][20] ) );
  NOR2_X1 U2642 ( .A1(n443), .A2(n292), .ZN(\ab[20][1] ) );
  NOR2_X1 U2643 ( .A1(n404), .A2(n292), .ZN(\ab[20][19] ) );
  NOR2_X1 U2644 ( .A1(n407), .A2(n292), .ZN(\ab[20][18] ) );
  NOR2_X1 U2645 ( .A1(n408), .A2(n292), .ZN(\ab[20][17] ) );
  NOR2_X1 U2646 ( .A1(n411), .A2(n292), .ZN(\ab[20][16] ) );
  NOR2_X1 U2647 ( .A1(n414), .A2(n292), .ZN(\ab[20][15] ) );
  NOR2_X1 U2648 ( .A1(n417), .A2(n292), .ZN(\ab[20][14] ) );
  NOR2_X1 U2649 ( .A1(n420), .A2(n292), .ZN(\ab[20][13] ) );
  NOR2_X1 U2650 ( .A1(n423), .A2(n292), .ZN(\ab[20][12] ) );
  NOR2_X1 U2651 ( .A1(n425), .A2(n292), .ZN(\ab[20][11] ) );
  NOR2_X1 U2652 ( .A1(n477), .A2(n292), .ZN(\ab[20][10] ) );
  NOR2_X1 U2653 ( .A1(n446), .A2(n292), .ZN(\ab[20][0] ) );
  NOR2_X1 U2654 ( .A1(n428), .A2(n330), .ZN(\ab[1][9] ) );
  NOR2_X1 U2655 ( .A1(n430), .A2(n330), .ZN(\ab[1][8] ) );
  NOR2_X1 U2656 ( .A1(n432), .A2(n330), .ZN(\ab[1][7] ) );
  NOR2_X1 U2657 ( .A1(n434), .A2(n330), .ZN(\ab[1][6] ) );
  NOR2_X1 U2658 ( .A1(n436), .A2(n330), .ZN(\ab[1][5] ) );
  NOR2_X1 U2659 ( .A1(n336), .A2(n331), .ZN(\ab[1][52] ) );
  NOR2_X1 U2660 ( .A1(n340), .A2(n331), .ZN(\ab[1][51] ) );
  NOR2_X1 U2661 ( .A1(n342), .A2(n332), .ZN(\ab[1][50] ) );
  NOR2_X1 U2662 ( .A1(n438), .A2(n330), .ZN(\ab[1][4] ) );
  NOR2_X1 U2663 ( .A1(n343), .A2(n332), .ZN(\ab[1][49] ) );
  NOR2_X1 U2664 ( .A1(n346), .A2(n332), .ZN(\ab[1][48] ) );
  NOR2_X1 U2665 ( .A1(n348), .A2(n332), .ZN(\ab[1][47] ) );
  NOR2_X1 U2666 ( .A1(n350), .A2(n332), .ZN(\ab[1][46] ) );
  NOR2_X1 U2667 ( .A1(n352), .A2(n332), .ZN(\ab[1][45] ) );
  NOR2_X1 U2668 ( .A1(n353), .A2(n332), .ZN(\ab[1][44] ) );
  NOR2_X1 U2669 ( .A1(n356), .A2(n332), .ZN(\ab[1][43] ) );
  NOR2_X1 U2670 ( .A1(n358), .A2(n332), .ZN(\ab[1][42] ) );
  NOR2_X1 U2671 ( .A1(n362), .A2(n332), .ZN(\ab[1][41] ) );
  NOR2_X1 U2672 ( .A1(n364), .A2(n332), .ZN(\ab[1][40] ) );
  NOR2_X1 U2673 ( .A1(n440), .A2(n332), .ZN(\ab[1][3] ) );
  NOR2_X1 U2674 ( .A1(n366), .A2(n331), .ZN(\ab[1][39] ) );
  NOR2_X1 U2675 ( .A1(n368), .A2(n331), .ZN(\ab[1][38] ) );
  NOR2_X1 U2676 ( .A1(n370), .A2(n331), .ZN(\ab[1][37] ) );
  NOR2_X1 U2677 ( .A1(n474), .A2(n331), .ZN(\ab[1][36] ) );
  NOR2_X1 U2678 ( .A1(n374), .A2(n331), .ZN(\ab[1][35] ) );
  NOR2_X1 U2679 ( .A1(n376), .A2(n331), .ZN(\ab[1][34] ) );
  NOR2_X1 U2680 ( .A1(n378), .A2(n331), .ZN(\ab[1][33] ) );
  NOR2_X1 U2681 ( .A1(n380), .A2(n331), .ZN(\ab[1][32] ) );
  NOR2_X1 U2682 ( .A1(n382), .A2(n331), .ZN(\ab[1][31] ) );
  NOR2_X1 U2683 ( .A1(n384), .A2(n331), .ZN(\ab[1][30] ) );
  NOR2_X1 U2684 ( .A1(n442), .A2(n331), .ZN(\ab[1][2] ) );
  NOR2_X1 U2685 ( .A1(n386), .A2(n330), .ZN(\ab[1][29] ) );
  NOR2_X1 U2686 ( .A1(n387), .A2(n330), .ZN(\ab[1][28] ) );
  NOR2_X1 U2687 ( .A1(n390), .A2(n330), .ZN(\ab[1][27] ) );
  NOR2_X1 U2688 ( .A1(n392), .A2(n330), .ZN(\ab[1][26] ) );
  NOR2_X1 U2689 ( .A1(n394), .A2(n330), .ZN(\ab[1][25] ) );
  NOR2_X1 U2690 ( .A1(n396), .A2(n330), .ZN(\ab[1][24] ) );
  NOR2_X1 U2691 ( .A1(n398), .A2(n330), .ZN(\ab[1][23] ) );
  NOR2_X1 U2692 ( .A1(n400), .A2(n330), .ZN(\ab[1][22] ) );
  NOR2_X1 U2693 ( .A1(n402), .A2(n330), .ZN(\ab[1][21] ) );
  NOR2_X1 U2694 ( .A1(n475), .A2(n330), .ZN(\ab[1][20] ) );
  NOR2_X1 U2695 ( .A1(n445), .A2(n330), .ZN(\ab[1][1] ) );
  NOR2_X1 U2696 ( .A1(n404), .A2(n330), .ZN(\ab[1][19] ) );
  NOR2_X1 U2697 ( .A1(n476), .A2(n330), .ZN(\ab[1][18] ) );
  NOR2_X1 U2698 ( .A1(n409), .A2(n330), .ZN(\ab[1][17] ) );
  NOR2_X1 U2699 ( .A1(n410), .A2(n330), .ZN(\ab[1][16] ) );
  NOR2_X1 U2700 ( .A1(n413), .A2(n330), .ZN(\ab[1][15] ) );
  NOR2_X1 U2701 ( .A1(n416), .A2(n330), .ZN(\ab[1][14] ) );
  NOR2_X1 U2702 ( .A1(n419), .A2(n330), .ZN(\ab[1][13] ) );
  NOR2_X1 U2703 ( .A1(n422), .A2(n330), .ZN(\ab[1][12] ) );
  NOR2_X1 U2704 ( .A1(n426), .A2(n330), .ZN(\ab[1][11] ) );
  NOR2_X1 U2705 ( .A1(n477), .A2(n330), .ZN(\ab[1][10] ) );
  NOR2_X1 U2706 ( .A1(n480), .A2(n330), .ZN(\ab[1][0] ) );
  NOR2_X1 U2707 ( .A1(n428), .A2(n294), .ZN(\ab[19][9] ) );
  NOR2_X1 U2708 ( .A1(n431), .A2(n294), .ZN(\ab[19][8] ) );
  NOR2_X1 U2709 ( .A1(n432), .A2(n294), .ZN(\ab[19][7] ) );
  NOR2_X1 U2710 ( .A1(n434), .A2(n294), .ZN(\ab[19][6] ) );
  NOR2_X1 U2711 ( .A1(n436), .A2(n294), .ZN(\ab[19][5] ) );
  NOR2_X1 U2712 ( .A1(n336), .A2(n294), .ZN(\ab[19][52] ) );
  NOR2_X1 U2713 ( .A1(n339), .A2(n294), .ZN(\ab[19][51] ) );
  NOR2_X1 U2714 ( .A1(n341), .A2(n294), .ZN(\ab[19][50] ) );
  NOR2_X1 U2715 ( .A1(n438), .A2(n294), .ZN(\ab[19][4] ) );
  NOR2_X1 U2716 ( .A1(n344), .A2(n294), .ZN(\ab[19][49] ) );
  NOR2_X1 U2717 ( .A1(n346), .A2(n294), .ZN(\ab[19][48] ) );
  NOR2_X1 U2718 ( .A1(n348), .A2(n294), .ZN(\ab[19][47] ) );
  NOR2_X1 U2719 ( .A1(n350), .A2(n294), .ZN(\ab[19][46] ) );
  NOR2_X1 U2720 ( .A1(n352), .A2(n294), .ZN(\ab[19][45] ) );
  NOR2_X1 U2721 ( .A1(n354), .A2(n294), .ZN(\ab[19][44] ) );
  NOR2_X1 U2722 ( .A1(n357), .A2(n294), .ZN(\ab[19][43] ) );
  NOR2_X1 U2723 ( .A1(n359), .A2(n294), .ZN(\ab[19][42] ) );
  NOR2_X1 U2724 ( .A1(n362), .A2(n294), .ZN(\ab[19][41] ) );
  NOR2_X1 U2725 ( .A1(n364), .A2(n294), .ZN(\ab[19][40] ) );
  NOR2_X1 U2726 ( .A1(n441), .A2(n294), .ZN(\ab[19][3] ) );
  NOR2_X1 U2727 ( .A1(n366), .A2(n293), .ZN(\ab[19][39] ) );
  NOR2_X1 U2728 ( .A1(n367), .A2(n293), .ZN(\ab[19][38] ) );
  NOR2_X1 U2729 ( .A1(n371), .A2(n293), .ZN(\ab[19][37] ) );
  NOR2_X1 U2730 ( .A1(n474), .A2(n293), .ZN(\ab[19][36] ) );
  NOR2_X1 U2731 ( .A1(n374), .A2(n293), .ZN(\ab[19][35] ) );
  NOR2_X1 U2732 ( .A1(n376), .A2(n293), .ZN(\ab[19][34] ) );
  NOR2_X1 U2733 ( .A1(n378), .A2(n293), .ZN(\ab[19][33] ) );
  NOR2_X1 U2734 ( .A1(n380), .A2(n293), .ZN(\ab[19][32] ) );
  NOR2_X1 U2735 ( .A1(n382), .A2(n293), .ZN(\ab[19][31] ) );
  NOR2_X1 U2736 ( .A1(n384), .A2(n293), .ZN(\ab[19][30] ) );
  NOR2_X1 U2737 ( .A1(n479), .A2(n293), .ZN(\ab[19][2] ) );
  NOR2_X1 U2738 ( .A1(n385), .A2(n294), .ZN(\ab[19][29] ) );
  NOR2_X1 U2739 ( .A1(n388), .A2(n294), .ZN(\ab[19][28] ) );
  NOR2_X1 U2740 ( .A1(n389), .A2(n294), .ZN(\ab[19][27] ) );
  NOR2_X1 U2741 ( .A1(n391), .A2(n294), .ZN(\ab[19][26] ) );
  NOR2_X1 U2742 ( .A1(n393), .A2(n294), .ZN(\ab[19][25] ) );
  NOR2_X1 U2743 ( .A1(n395), .A2(n293), .ZN(\ab[19][24] ) );
  NOR2_X1 U2744 ( .A1(n397), .A2(n293), .ZN(\ab[19][23] ) );
  NOR2_X1 U2745 ( .A1(n399), .A2(n293), .ZN(\ab[19][22] ) );
  NOR2_X1 U2746 ( .A1(n401), .A2(n293), .ZN(\ab[19][21] ) );
  NOR2_X1 U2747 ( .A1(n403), .A2(n293), .ZN(\ab[19][20] ) );
  NOR2_X1 U2748 ( .A1(n443), .A2(n293), .ZN(\ab[19][1] ) );
  NOR2_X1 U2749 ( .A1(n405), .A2(n294), .ZN(\ab[19][19] ) );
  NOR2_X1 U2750 ( .A1(n407), .A2(n294), .ZN(\ab[19][18] ) );
  NOR2_X1 U2751 ( .A1(n409), .A2(n294), .ZN(\ab[19][17] ) );
  NOR2_X1 U2752 ( .A1(n411), .A2(n294), .ZN(\ab[19][16] ) );
  NOR2_X1 U2753 ( .A1(n414), .A2(n294), .ZN(\ab[19][15] ) );
  NOR2_X1 U2754 ( .A1(n417), .A2(n294), .ZN(\ab[19][14] ) );
  NOR2_X1 U2755 ( .A1(n420), .A2(n294), .ZN(\ab[19][13] ) );
  NOR2_X1 U2756 ( .A1(n423), .A2(n294), .ZN(\ab[19][12] ) );
  NOR2_X1 U2757 ( .A1(n426), .A2(n294), .ZN(\ab[19][11] ) );
  NOR2_X1 U2758 ( .A1(n427), .A2(n294), .ZN(\ab[19][10] ) );
  NOR2_X1 U2759 ( .A1(n480), .A2(n294), .ZN(\ab[19][0] ) );
  NOR2_X1 U2760 ( .A1(n428), .A2(n295), .ZN(\ab[18][9] ) );
  NOR2_X1 U2761 ( .A1(n431), .A2(n295), .ZN(\ab[18][8] ) );
  NOR2_X1 U2762 ( .A1(n432), .A2(n295), .ZN(\ab[18][7] ) );
  NOR2_X1 U2763 ( .A1(n434), .A2(n295), .ZN(\ab[18][6] ) );
  NOR2_X1 U2764 ( .A1(n436), .A2(n295), .ZN(\ab[18][5] ) );
  NOR2_X1 U2765 ( .A1(n336), .A2(n295), .ZN(\ab[18][52] ) );
  NOR2_X1 U2766 ( .A1(n339), .A2(n295), .ZN(\ab[18][51] ) );
  NOR2_X1 U2767 ( .A1(n341), .A2(n295), .ZN(\ab[18][50] ) );
  NOR2_X1 U2768 ( .A1(n438), .A2(n295), .ZN(\ab[18][4] ) );
  NOR2_X1 U2769 ( .A1(n344), .A2(n296), .ZN(\ab[18][49] ) );
  NOR2_X1 U2770 ( .A1(n345), .A2(n296), .ZN(\ab[18][48] ) );
  NOR2_X1 U2771 ( .A1(n347), .A2(n296), .ZN(\ab[18][47] ) );
  NOR2_X1 U2772 ( .A1(n349), .A2(n296), .ZN(\ab[18][46] ) );
  NOR2_X1 U2773 ( .A1(n351), .A2(n296), .ZN(\ab[18][45] ) );
  NOR2_X1 U2774 ( .A1(n354), .A2(n296), .ZN(\ab[18][44] ) );
  NOR2_X1 U2775 ( .A1(n357), .A2(n296), .ZN(\ab[18][43] ) );
  NOR2_X1 U2776 ( .A1(n359), .A2(n296), .ZN(\ab[18][42] ) );
  NOR2_X1 U2777 ( .A1(n361), .A2(n296), .ZN(\ab[18][41] ) );
  NOR2_X1 U2778 ( .A1(n363), .A2(n296), .ZN(\ab[18][40] ) );
  NOR2_X1 U2779 ( .A1(n441), .A2(n296), .ZN(\ab[18][3] ) );
  NOR2_X1 U2780 ( .A1(n365), .A2(n295), .ZN(\ab[18][39] ) );
  NOR2_X1 U2781 ( .A1(n367), .A2(n465), .ZN(\ab[18][38] ) );
  NOR2_X1 U2782 ( .A1(n371), .A2(n465), .ZN(\ab[18][37] ) );
  NOR2_X1 U2783 ( .A1(n372), .A2(n465), .ZN(\ab[18][36] ) );
  NOR2_X1 U2784 ( .A1(n373), .A2(n465), .ZN(\ab[18][35] ) );
  NOR2_X1 U2785 ( .A1(n375), .A2(n465), .ZN(\ab[18][34] ) );
  NOR2_X1 U2786 ( .A1(n377), .A2(n465), .ZN(\ab[18][33] ) );
  NOR2_X1 U2787 ( .A1(n379), .A2(n465), .ZN(\ab[18][32] ) );
  NOR2_X1 U2788 ( .A1(n381), .A2(n296), .ZN(\ab[18][31] ) );
  NOR2_X1 U2789 ( .A1(n383), .A2(n296), .ZN(\ab[18][30] ) );
  NOR2_X1 U2790 ( .A1(n479), .A2(n295), .ZN(\ab[18][2] ) );
  NOR2_X1 U2791 ( .A1(n385), .A2(n296), .ZN(\ab[18][29] ) );
  NOR2_X1 U2792 ( .A1(n388), .A2(n296), .ZN(\ab[18][28] ) );
  NOR2_X1 U2793 ( .A1(n389), .A2(n295), .ZN(\ab[18][27] ) );
  NOR2_X1 U2794 ( .A1(n391), .A2(n295), .ZN(\ab[18][26] ) );
  NOR2_X1 U2795 ( .A1(n393), .A2(n295), .ZN(\ab[18][25] ) );
  NOR2_X1 U2796 ( .A1(n395), .A2(n295), .ZN(\ab[18][24] ) );
  NOR2_X1 U2797 ( .A1(n397), .A2(n296), .ZN(\ab[18][23] ) );
  NOR2_X1 U2798 ( .A1(n399), .A2(n296), .ZN(\ab[18][22] ) );
  NOR2_X1 U2799 ( .A1(n401), .A2(n295), .ZN(\ab[18][21] ) );
  NOR2_X1 U2800 ( .A1(n475), .A2(n296), .ZN(\ab[18][20] ) );
  NOR2_X1 U2801 ( .A1(n443), .A2(n296), .ZN(\ab[18][1] ) );
  NOR2_X1 U2802 ( .A1(n405), .A2(n295), .ZN(\ab[18][19] ) );
  NOR2_X1 U2803 ( .A1(n407), .A2(n295), .ZN(\ab[18][18] ) );
  NOR2_X1 U2804 ( .A1(n408), .A2(n295), .ZN(\ab[18][17] ) );
  NOR2_X1 U2805 ( .A1(n411), .A2(n295), .ZN(\ab[18][16] ) );
  NOR2_X1 U2806 ( .A1(n414), .A2(n295), .ZN(\ab[18][15] ) );
  NOR2_X1 U2807 ( .A1(n417), .A2(n295), .ZN(\ab[18][14] ) );
  NOR2_X1 U2808 ( .A1(n420), .A2(n295), .ZN(\ab[18][13] ) );
  NOR2_X1 U2809 ( .A1(n423), .A2(n295), .ZN(\ab[18][12] ) );
  NOR2_X1 U2810 ( .A1(n425), .A2(n295), .ZN(\ab[18][11] ) );
  NOR2_X1 U2811 ( .A1(n477), .A2(n295), .ZN(\ab[18][10] ) );
  NOR2_X1 U2812 ( .A1(n446), .A2(n295), .ZN(\ab[18][0] ) );
  NOR2_X1 U2813 ( .A1(n428), .A2(n297), .ZN(\ab[17][9] ) );
  NOR2_X1 U2814 ( .A1(n431), .A2(n297), .ZN(\ab[17][8] ) );
  NOR2_X1 U2815 ( .A1(n432), .A2(n297), .ZN(\ab[17][7] ) );
  NOR2_X1 U2816 ( .A1(n434), .A2(n297), .ZN(\ab[17][6] ) );
  NOR2_X1 U2817 ( .A1(n436), .A2(n297), .ZN(\ab[17][5] ) );
  NOR2_X1 U2818 ( .A1(n336), .A2(n297), .ZN(\ab[17][52] ) );
  NOR2_X1 U2819 ( .A1(n339), .A2(n297), .ZN(\ab[17][51] ) );
  NOR2_X1 U2820 ( .A1(n341), .A2(n297), .ZN(\ab[17][50] ) );
  NOR2_X1 U2821 ( .A1(n438), .A2(n297), .ZN(\ab[17][4] ) );
  NOR2_X1 U2822 ( .A1(n344), .A2(n298), .ZN(\ab[17][49] ) );
  NOR2_X1 U2823 ( .A1(n346), .A2(n298), .ZN(\ab[17][48] ) );
  NOR2_X1 U2824 ( .A1(n348), .A2(n298), .ZN(\ab[17][47] ) );
  NOR2_X1 U2825 ( .A1(n350), .A2(n298), .ZN(\ab[17][46] ) );
  NOR2_X1 U2826 ( .A1(n352), .A2(n298), .ZN(\ab[17][45] ) );
  NOR2_X1 U2827 ( .A1(n354), .A2(n298), .ZN(\ab[17][44] ) );
  NOR2_X1 U2828 ( .A1(n357), .A2(n298), .ZN(\ab[17][43] ) );
  NOR2_X1 U2829 ( .A1(n359), .A2(n298), .ZN(\ab[17][42] ) );
  NOR2_X1 U2830 ( .A1(n362), .A2(n298), .ZN(\ab[17][41] ) );
  NOR2_X1 U2831 ( .A1(n364), .A2(n298), .ZN(\ab[17][40] ) );
  NOR2_X1 U2832 ( .A1(n441), .A2(n298), .ZN(\ab[17][3] ) );
  NOR2_X1 U2833 ( .A1(n366), .A2(n466), .ZN(\ab[17][39] ) );
  NOR2_X1 U2834 ( .A1(n367), .A2(n466), .ZN(\ab[17][38] ) );
  NOR2_X1 U2835 ( .A1(n371), .A2(n466), .ZN(\ab[17][37] ) );
  NOR2_X1 U2836 ( .A1(n474), .A2(n466), .ZN(\ab[17][36] ) );
  NOR2_X1 U2837 ( .A1(n374), .A2(n466), .ZN(\ab[17][35] ) );
  NOR2_X1 U2838 ( .A1(n376), .A2(n466), .ZN(\ab[17][34] ) );
  NOR2_X1 U2839 ( .A1(n378), .A2(n466), .ZN(\ab[17][33] ) );
  NOR2_X1 U2840 ( .A1(n380), .A2(n466), .ZN(\ab[17][32] ) );
  NOR2_X1 U2841 ( .A1(n382), .A2(n298), .ZN(\ab[17][31] ) );
  NOR2_X1 U2842 ( .A1(n384), .A2(n298), .ZN(\ab[17][30] ) );
  NOR2_X1 U2843 ( .A1(n479), .A2(n297), .ZN(\ab[17][2] ) );
  NOR2_X1 U2844 ( .A1(n385), .A2(n298), .ZN(\ab[17][29] ) );
  NOR2_X1 U2845 ( .A1(n388), .A2(n297), .ZN(\ab[17][28] ) );
  NOR2_X1 U2846 ( .A1(n389), .A2(n297), .ZN(\ab[17][27] ) );
  NOR2_X1 U2847 ( .A1(n391), .A2(n298), .ZN(\ab[17][26] ) );
  NOR2_X1 U2848 ( .A1(n393), .A2(n297), .ZN(\ab[17][25] ) );
  NOR2_X1 U2849 ( .A1(n395), .A2(n298), .ZN(\ab[17][24] ) );
  NOR2_X1 U2850 ( .A1(n397), .A2(n298), .ZN(\ab[17][23] ) );
  NOR2_X1 U2851 ( .A1(n399), .A2(n298), .ZN(\ab[17][22] ) );
  NOR2_X1 U2852 ( .A1(n401), .A2(n298), .ZN(\ab[17][21] ) );
  NOR2_X1 U2853 ( .A1(n403), .A2(n298), .ZN(\ab[17][20] ) );
  NOR2_X1 U2854 ( .A1(n443), .A2(n297), .ZN(\ab[17][1] ) );
  NOR2_X1 U2855 ( .A1(n405), .A2(n297), .ZN(\ab[17][19] ) );
  NOR2_X1 U2856 ( .A1(n407), .A2(n297), .ZN(\ab[17][18] ) );
  NOR2_X1 U2857 ( .A1(n409), .A2(n297), .ZN(\ab[17][17] ) );
  NOR2_X1 U2858 ( .A1(n411), .A2(n297), .ZN(\ab[17][16] ) );
  NOR2_X1 U2859 ( .A1(n414), .A2(n297), .ZN(\ab[17][15] ) );
  NOR2_X1 U2860 ( .A1(n417), .A2(n297), .ZN(\ab[17][14] ) );
  NOR2_X1 U2861 ( .A1(n420), .A2(n297), .ZN(\ab[17][13] ) );
  NOR2_X1 U2862 ( .A1(n423), .A2(n297), .ZN(\ab[17][12] ) );
  NOR2_X1 U2863 ( .A1(n426), .A2(n297), .ZN(\ab[17][11] ) );
  NOR2_X1 U2864 ( .A1(n427), .A2(n297), .ZN(\ab[17][10] ) );
  NOR2_X1 U2865 ( .A1(n480), .A2(n297), .ZN(\ab[17][0] ) );
  NOR2_X1 U2866 ( .A1(n428), .A2(n299), .ZN(\ab[16][9] ) );
  NOR2_X1 U2867 ( .A1(n431), .A2(n299), .ZN(\ab[16][8] ) );
  NOR2_X1 U2868 ( .A1(n432), .A2(n299), .ZN(\ab[16][7] ) );
  NOR2_X1 U2869 ( .A1(n434), .A2(n299), .ZN(\ab[16][6] ) );
  NOR2_X1 U2870 ( .A1(n436), .A2(n299), .ZN(\ab[16][5] ) );
  NOR2_X1 U2871 ( .A1(n336), .A2(n299), .ZN(\ab[16][52] ) );
  NOR2_X1 U2872 ( .A1(n339), .A2(n299), .ZN(\ab[16][51] ) );
  NOR2_X1 U2873 ( .A1(n341), .A2(n299), .ZN(\ab[16][50] ) );
  NOR2_X1 U2874 ( .A1(n438), .A2(n299), .ZN(\ab[16][4] ) );
  NOR2_X1 U2875 ( .A1(n344), .A2(n300), .ZN(\ab[16][49] ) );
  NOR2_X1 U2876 ( .A1(n345), .A2(n300), .ZN(\ab[16][48] ) );
  NOR2_X1 U2877 ( .A1(n347), .A2(n300), .ZN(\ab[16][47] ) );
  NOR2_X1 U2878 ( .A1(n349), .A2(n300), .ZN(\ab[16][46] ) );
  NOR2_X1 U2879 ( .A1(n351), .A2(n300), .ZN(\ab[16][45] ) );
  NOR2_X1 U2880 ( .A1(n354), .A2(n300), .ZN(\ab[16][44] ) );
  NOR2_X1 U2881 ( .A1(n357), .A2(n300), .ZN(\ab[16][43] ) );
  NOR2_X1 U2882 ( .A1(n359), .A2(n300), .ZN(\ab[16][42] ) );
  NOR2_X1 U2883 ( .A1(n361), .A2(n300), .ZN(\ab[16][41] ) );
  NOR2_X1 U2884 ( .A1(n363), .A2(n300), .ZN(\ab[16][40] ) );
  NOR2_X1 U2885 ( .A1(n441), .A2(n300), .ZN(\ab[16][3] ) );
  NOR2_X1 U2886 ( .A1(n365), .A2(n467), .ZN(\ab[16][39] ) );
  NOR2_X1 U2887 ( .A1(n367), .A2(n467), .ZN(\ab[16][38] ) );
  NOR2_X1 U2888 ( .A1(n371), .A2(n467), .ZN(\ab[16][37] ) );
  NOR2_X1 U2889 ( .A1(n372), .A2(n467), .ZN(\ab[16][36] ) );
  NOR2_X1 U2890 ( .A1(n373), .A2(n300), .ZN(\ab[16][35] ) );
  NOR2_X1 U2891 ( .A1(n375), .A2(n300), .ZN(\ab[16][34] ) );
  NOR2_X1 U2892 ( .A1(n377), .A2(n300), .ZN(\ab[16][33] ) );
  NOR2_X1 U2893 ( .A1(n379), .A2(n300), .ZN(\ab[16][32] ) );
  NOR2_X1 U2894 ( .A1(n381), .A2(n300), .ZN(\ab[16][31] ) );
  NOR2_X1 U2895 ( .A1(n383), .A2(n300), .ZN(\ab[16][30] ) );
  NOR2_X1 U2896 ( .A1(n479), .A2(n300), .ZN(\ab[16][2] ) );
  NOR2_X1 U2897 ( .A1(n386), .A2(n299), .ZN(\ab[16][29] ) );
  NOR2_X1 U2898 ( .A1(n388), .A2(n299), .ZN(\ab[16][28] ) );
  NOR2_X1 U2899 ( .A1(n390), .A2(n299), .ZN(\ab[16][27] ) );
  NOR2_X1 U2900 ( .A1(n391), .A2(n299), .ZN(\ab[16][26] ) );
  NOR2_X1 U2901 ( .A1(n394), .A2(n299), .ZN(\ab[16][25] ) );
  NOR2_X1 U2902 ( .A1(n395), .A2(n299), .ZN(\ab[16][24] ) );
  NOR2_X1 U2903 ( .A1(n398), .A2(n299), .ZN(\ab[16][23] ) );
  NOR2_X1 U2904 ( .A1(n400), .A2(n299), .ZN(\ab[16][22] ) );
  NOR2_X1 U2905 ( .A1(n402), .A2(n299), .ZN(\ab[16][21] ) );
  NOR2_X1 U2906 ( .A1(n475), .A2(n299), .ZN(\ab[16][20] ) );
  NOR2_X1 U2907 ( .A1(n443), .A2(n299), .ZN(\ab[16][1] ) );
  NOR2_X1 U2908 ( .A1(n405), .A2(n299), .ZN(\ab[16][19] ) );
  NOR2_X1 U2909 ( .A1(n407), .A2(n299), .ZN(\ab[16][18] ) );
  NOR2_X1 U2910 ( .A1(n408), .A2(n299), .ZN(\ab[16][17] ) );
  NOR2_X1 U2911 ( .A1(n411), .A2(n299), .ZN(\ab[16][16] ) );
  NOR2_X1 U2912 ( .A1(n414), .A2(n299), .ZN(\ab[16][15] ) );
  NOR2_X1 U2913 ( .A1(n417), .A2(n299), .ZN(\ab[16][14] ) );
  NOR2_X1 U2914 ( .A1(n420), .A2(n299), .ZN(\ab[16][13] ) );
  NOR2_X1 U2915 ( .A1(n423), .A2(n299), .ZN(\ab[16][12] ) );
  NOR2_X1 U2916 ( .A1(n425), .A2(n299), .ZN(\ab[16][11] ) );
  NOR2_X1 U2917 ( .A1(n477), .A2(n299), .ZN(\ab[16][10] ) );
  NOR2_X1 U2918 ( .A1(n446), .A2(n299), .ZN(\ab[16][0] ) );
  NOR2_X1 U2919 ( .A1(n429), .A2(n301), .ZN(\ab[15][9] ) );
  NOR2_X1 U2920 ( .A1(n431), .A2(n301), .ZN(\ab[15][8] ) );
  NOR2_X1 U2921 ( .A1(n433), .A2(n301), .ZN(\ab[15][7] ) );
  NOR2_X1 U2922 ( .A1(n434), .A2(n301), .ZN(\ab[15][6] ) );
  NOR2_X1 U2923 ( .A1(n436), .A2(n301), .ZN(\ab[15][5] ) );
  NOR2_X1 U2924 ( .A1(n336), .A2(n301), .ZN(\ab[15][52] ) );
  NOR2_X1 U2925 ( .A1(n339), .A2(n301), .ZN(\ab[15][51] ) );
  NOR2_X1 U2926 ( .A1(n341), .A2(n301), .ZN(\ab[15][50] ) );
  NOR2_X1 U2927 ( .A1(n438), .A2(n301), .ZN(\ab[15][4] ) );
  NOR2_X1 U2928 ( .A1(n344), .A2(n302), .ZN(\ab[15][49] ) );
  NOR2_X1 U2929 ( .A1(n346), .A2(n302), .ZN(\ab[15][48] ) );
  NOR2_X1 U2930 ( .A1(n348), .A2(n302), .ZN(\ab[15][47] ) );
  NOR2_X1 U2931 ( .A1(n350), .A2(n302), .ZN(\ab[15][46] ) );
  NOR2_X1 U2932 ( .A1(n352), .A2(n302), .ZN(\ab[15][45] ) );
  NOR2_X1 U2933 ( .A1(n354), .A2(n302), .ZN(\ab[15][44] ) );
  NOR2_X1 U2934 ( .A1(n357), .A2(n302), .ZN(\ab[15][43] ) );
  NOR2_X1 U2935 ( .A1(n359), .A2(n302), .ZN(\ab[15][42] ) );
  NOR2_X1 U2936 ( .A1(n362), .A2(n302), .ZN(\ab[15][41] ) );
  NOR2_X1 U2937 ( .A1(n364), .A2(n302), .ZN(\ab[15][40] ) );
  NOR2_X1 U2938 ( .A1(n441), .A2(n302), .ZN(\ab[15][3] ) );
  NOR2_X1 U2939 ( .A1(n366), .A2(n468), .ZN(\ab[15][39] ) );
  NOR2_X1 U2940 ( .A1(n367), .A2(n302), .ZN(\ab[15][38] ) );
  NOR2_X1 U2941 ( .A1(n371), .A2(n302), .ZN(\ab[15][37] ) );
  NOR2_X1 U2942 ( .A1(n474), .A2(n302), .ZN(\ab[15][36] ) );
  NOR2_X1 U2943 ( .A1(n374), .A2(n302), .ZN(\ab[15][35] ) );
  NOR2_X1 U2944 ( .A1(n376), .A2(n468), .ZN(\ab[15][34] ) );
  NOR2_X1 U2945 ( .A1(n378), .A2(n468), .ZN(\ab[15][33] ) );
  NOR2_X1 U2946 ( .A1(n380), .A2(n468), .ZN(\ab[15][32] ) );
  NOR2_X1 U2947 ( .A1(n382), .A2(n301), .ZN(\ab[15][31] ) );
  NOR2_X1 U2948 ( .A1(n384), .A2(n301), .ZN(\ab[15][30] ) );
  NOR2_X1 U2949 ( .A1(n479), .A2(n301), .ZN(\ab[15][2] ) );
  NOR2_X1 U2950 ( .A1(n385), .A2(n301), .ZN(\ab[15][29] ) );
  NOR2_X1 U2951 ( .A1(n388), .A2(n301), .ZN(\ab[15][28] ) );
  NOR2_X1 U2952 ( .A1(n389), .A2(n301), .ZN(\ab[15][27] ) );
  NOR2_X1 U2953 ( .A1(n392), .A2(n301), .ZN(\ab[15][26] ) );
  NOR2_X1 U2954 ( .A1(n393), .A2(n301), .ZN(\ab[15][25] ) );
  NOR2_X1 U2955 ( .A1(n396), .A2(n301), .ZN(\ab[15][24] ) );
  NOR2_X1 U2956 ( .A1(n397), .A2(n301), .ZN(\ab[15][23] ) );
  NOR2_X1 U2957 ( .A1(n399), .A2(n301), .ZN(\ab[15][22] ) );
  NOR2_X1 U2958 ( .A1(n401), .A2(n301), .ZN(\ab[15][21] ) );
  NOR2_X1 U2959 ( .A1(n403), .A2(n301), .ZN(\ab[15][20] ) );
  NOR2_X1 U2960 ( .A1(n443), .A2(n301), .ZN(\ab[15][1] ) );
  NOR2_X1 U2961 ( .A1(n405), .A2(n301), .ZN(\ab[15][19] ) );
  NOR2_X1 U2962 ( .A1(n407), .A2(n301), .ZN(\ab[15][18] ) );
  NOR2_X1 U2963 ( .A1(n409), .A2(n301), .ZN(\ab[15][17] ) );
  NOR2_X1 U2964 ( .A1(n411), .A2(n301), .ZN(\ab[15][16] ) );
  NOR2_X1 U2965 ( .A1(n414), .A2(n301), .ZN(\ab[15][15] ) );
  NOR2_X1 U2966 ( .A1(n417), .A2(n301), .ZN(\ab[15][14] ) );
  NOR2_X1 U2967 ( .A1(n420), .A2(n301), .ZN(\ab[15][13] ) );
  NOR2_X1 U2968 ( .A1(n423), .A2(n301), .ZN(\ab[15][12] ) );
  NOR2_X1 U2969 ( .A1(n426), .A2(n301), .ZN(\ab[15][11] ) );
  NOR2_X1 U2970 ( .A1(n427), .A2(n301), .ZN(\ab[15][10] ) );
  NOR2_X1 U2971 ( .A1(n480), .A2(n301), .ZN(\ab[15][0] ) );
  NOR2_X1 U2972 ( .A1(n428), .A2(n303), .ZN(\ab[14][9] ) );
  NOR2_X1 U2973 ( .A1(n431), .A2(n303), .ZN(\ab[14][8] ) );
  NOR2_X1 U2974 ( .A1(n432), .A2(n303), .ZN(\ab[14][7] ) );
  NOR2_X1 U2975 ( .A1(n434), .A2(n303), .ZN(\ab[14][6] ) );
  NOR2_X1 U2976 ( .A1(n436), .A2(n303), .ZN(\ab[14][5] ) );
  NOR2_X1 U2977 ( .A1(n337), .A2(n303), .ZN(\ab[14][52] ) );
  NOR2_X1 U2978 ( .A1(n339), .A2(n303), .ZN(\ab[14][51] ) );
  NOR2_X1 U2979 ( .A1(n341), .A2(n303), .ZN(\ab[14][50] ) );
  NOR2_X1 U2980 ( .A1(n438), .A2(n303), .ZN(\ab[14][4] ) );
  NOR2_X1 U2981 ( .A1(n344), .A2(n469), .ZN(\ab[14][49] ) );
  NOR2_X1 U2982 ( .A1(n345), .A2(n469), .ZN(\ab[14][48] ) );
  NOR2_X1 U2983 ( .A1(n347), .A2(n469), .ZN(\ab[14][47] ) );
  NOR2_X1 U2984 ( .A1(n349), .A2(n469), .ZN(\ab[14][46] ) );
  NOR2_X1 U2985 ( .A1(n351), .A2(n469), .ZN(\ab[14][45] ) );
  NOR2_X1 U2986 ( .A1(n354), .A2(n469), .ZN(\ab[14][44] ) );
  NOR2_X1 U2987 ( .A1(n357), .A2(n469), .ZN(\ab[14][43] ) );
  NOR2_X1 U2988 ( .A1(n359), .A2(n469), .ZN(\ab[14][42] ) );
  NOR2_X1 U2989 ( .A1(n361), .A2(n469), .ZN(\ab[14][41] ) );
  NOR2_X1 U2990 ( .A1(n363), .A2(n303), .ZN(\ab[14][40] ) );
  NOR2_X1 U2991 ( .A1(n441), .A2(n469), .ZN(\ab[14][3] ) );
  NOR2_X1 U2992 ( .A1(n365), .A2(n303), .ZN(\ab[14][39] ) );
  NOR2_X1 U2993 ( .A1(n367), .A2(n303), .ZN(\ab[14][38] ) );
  NOR2_X1 U2994 ( .A1(n371), .A2(n303), .ZN(\ab[14][37] ) );
  NOR2_X1 U2995 ( .A1(n474), .A2(n303), .ZN(\ab[14][36] ) );
  NOR2_X1 U2996 ( .A1(n373), .A2(n303), .ZN(\ab[14][35] ) );
  NOR2_X1 U2997 ( .A1(n375), .A2(n303), .ZN(\ab[14][34] ) );
  NOR2_X1 U2998 ( .A1(n377), .A2(n303), .ZN(\ab[14][33] ) );
  NOR2_X1 U2999 ( .A1(n380), .A2(n303), .ZN(\ab[14][32] ) );
  NOR2_X1 U3000 ( .A1(n381), .A2(n303), .ZN(\ab[14][31] ) );
  NOR2_X1 U3001 ( .A1(n383), .A2(n303), .ZN(\ab[14][30] ) );
  NOR2_X1 U3002 ( .A1(n479), .A2(n303), .ZN(\ab[14][2] ) );
  NOR2_X1 U3003 ( .A1(n385), .A2(n303), .ZN(\ab[14][29] ) );
  NOR2_X1 U3004 ( .A1(n388), .A2(n303), .ZN(\ab[14][28] ) );
  NOR2_X1 U3005 ( .A1(n389), .A2(n303), .ZN(\ab[14][27] ) );
  NOR2_X1 U3006 ( .A1(n391), .A2(n303), .ZN(\ab[14][26] ) );
  NOR2_X1 U3007 ( .A1(n393), .A2(n303), .ZN(\ab[14][25] ) );
  NOR2_X1 U3008 ( .A1(n395), .A2(n303), .ZN(\ab[14][24] ) );
  NOR2_X1 U3009 ( .A1(n397), .A2(n303), .ZN(\ab[14][23] ) );
  NOR2_X1 U3010 ( .A1(n399), .A2(n303), .ZN(\ab[14][22] ) );
  NOR2_X1 U3011 ( .A1(n401), .A2(n303), .ZN(\ab[14][21] ) );
  NOR2_X1 U3012 ( .A1(n475), .A2(n303), .ZN(\ab[14][20] ) );
  NOR2_X1 U3013 ( .A1(n443), .A2(n303), .ZN(\ab[14][1] ) );
  NOR2_X1 U3014 ( .A1(n405), .A2(n303), .ZN(\ab[14][19] ) );
  NOR2_X1 U3015 ( .A1(n407), .A2(n303), .ZN(\ab[14][18] ) );
  NOR2_X1 U3016 ( .A1(n409), .A2(n303), .ZN(\ab[14][17] ) );
  NOR2_X1 U3017 ( .A1(n411), .A2(n303), .ZN(\ab[14][16] ) );
  NOR2_X1 U3018 ( .A1(n414), .A2(n303), .ZN(\ab[14][15] ) );
  NOR2_X1 U3019 ( .A1(n417), .A2(n303), .ZN(\ab[14][14] ) );
  NOR2_X1 U3020 ( .A1(n420), .A2(n303), .ZN(\ab[14][13] ) );
  NOR2_X1 U3021 ( .A1(n423), .A2(n303), .ZN(\ab[14][12] ) );
  NOR2_X1 U3022 ( .A1(n426), .A2(n303), .ZN(\ab[14][11] ) );
  NOR2_X1 U3023 ( .A1(n477), .A2(n303), .ZN(\ab[14][10] ) );
  NOR2_X1 U3024 ( .A1(n446), .A2(n303), .ZN(\ab[14][0] ) );
  NOR2_X1 U3025 ( .A1(n428), .A2(n304), .ZN(\ab[13][9] ) );
  NOR2_X1 U3026 ( .A1(n431), .A2(n304), .ZN(\ab[13][8] ) );
  NOR2_X1 U3027 ( .A1(n432), .A2(n304), .ZN(\ab[13][7] ) );
  NOR2_X1 U3028 ( .A1(n434), .A2(n304), .ZN(\ab[13][6] ) );
  NOR2_X1 U3029 ( .A1(n436), .A2(n304), .ZN(\ab[13][5] ) );
  NOR2_X1 U3030 ( .A1(n336), .A2(n304), .ZN(\ab[13][52] ) );
  NOR2_X1 U3031 ( .A1(n339), .A2(n304), .ZN(\ab[13][51] ) );
  NOR2_X1 U3032 ( .A1(n341), .A2(n304), .ZN(\ab[13][50] ) );
  NOR2_X1 U3033 ( .A1(n438), .A2(n304), .ZN(\ab[13][4] ) );
  NOR2_X1 U3034 ( .A1(n344), .A2(n305), .ZN(\ab[13][49] ) );
  NOR2_X1 U3035 ( .A1(n346), .A2(n305), .ZN(\ab[13][48] ) );
  NOR2_X1 U3036 ( .A1(n348), .A2(n305), .ZN(\ab[13][47] ) );
  NOR2_X1 U3037 ( .A1(n350), .A2(n305), .ZN(\ab[13][46] ) );
  NOR2_X1 U3038 ( .A1(n352), .A2(n305), .ZN(\ab[13][45] ) );
  NOR2_X1 U3039 ( .A1(n354), .A2(n305), .ZN(\ab[13][44] ) );
  NOR2_X1 U3040 ( .A1(n357), .A2(n305), .ZN(\ab[13][43] ) );
  NOR2_X1 U3041 ( .A1(n359), .A2(n305), .ZN(\ab[13][42] ) );
  NOR2_X1 U3042 ( .A1(n362), .A2(n305), .ZN(\ab[13][41] ) );
  NOR2_X1 U3043 ( .A1(n364), .A2(n305), .ZN(\ab[13][40] ) );
  NOR2_X1 U3044 ( .A1(n441), .A2(n305), .ZN(\ab[13][3] ) );
  NOR2_X1 U3045 ( .A1(n366), .A2(n305), .ZN(\ab[13][39] ) );
  NOR2_X1 U3046 ( .A1(n367), .A2(n305), .ZN(\ab[13][38] ) );
  NOR2_X1 U3047 ( .A1(n371), .A2(n305), .ZN(\ab[13][37] ) );
  NOR2_X1 U3048 ( .A1(n372), .A2(n305), .ZN(\ab[13][36] ) );
  NOR2_X1 U3049 ( .A1(n374), .A2(n304), .ZN(\ab[13][35] ) );
  NOR2_X1 U3050 ( .A1(n376), .A2(n304), .ZN(\ab[13][34] ) );
  NOR2_X1 U3051 ( .A1(n378), .A2(n304), .ZN(\ab[13][33] ) );
  NOR2_X1 U3052 ( .A1(n379), .A2(n305), .ZN(\ab[13][32] ) );
  NOR2_X1 U3053 ( .A1(n382), .A2(n305), .ZN(\ab[13][31] ) );
  NOR2_X1 U3054 ( .A1(n384), .A2(n305), .ZN(\ab[13][30] ) );
  NOR2_X1 U3055 ( .A1(n479), .A2(n304), .ZN(\ab[13][2] ) );
  NOR2_X1 U3056 ( .A1(n385), .A2(n304), .ZN(\ab[13][29] ) );
  NOR2_X1 U3057 ( .A1(n388), .A2(n304), .ZN(\ab[13][28] ) );
  NOR2_X1 U3058 ( .A1(n389), .A2(n304), .ZN(\ab[13][27] ) );
  NOR2_X1 U3059 ( .A1(n391), .A2(n304), .ZN(\ab[13][26] ) );
  NOR2_X1 U3060 ( .A1(n393), .A2(n304), .ZN(\ab[13][25] ) );
  NOR2_X1 U3061 ( .A1(n395), .A2(n304), .ZN(\ab[13][24] ) );
  NOR2_X1 U3062 ( .A1(n397), .A2(n304), .ZN(\ab[13][23] ) );
  NOR2_X1 U3063 ( .A1(n399), .A2(n304), .ZN(\ab[13][22] ) );
  NOR2_X1 U3064 ( .A1(n401), .A2(n304), .ZN(\ab[13][21] ) );
  NOR2_X1 U3065 ( .A1(n475), .A2(n304), .ZN(\ab[13][20] ) );
  NOR2_X1 U3066 ( .A1(n443), .A2(n304), .ZN(\ab[13][1] ) );
  NOR2_X1 U3067 ( .A1(n405), .A2(n304), .ZN(\ab[13][19] ) );
  NOR2_X1 U3068 ( .A1(n407), .A2(n304), .ZN(\ab[13][18] ) );
  NOR2_X1 U3069 ( .A1(n408), .A2(n304), .ZN(\ab[13][17] ) );
  NOR2_X1 U3070 ( .A1(n411), .A2(n304), .ZN(\ab[13][16] ) );
  NOR2_X1 U3071 ( .A1(n414), .A2(n304), .ZN(\ab[13][15] ) );
  NOR2_X1 U3072 ( .A1(n417), .A2(n304), .ZN(\ab[13][14] ) );
  NOR2_X1 U3073 ( .A1(n420), .A2(n304), .ZN(\ab[13][13] ) );
  NOR2_X1 U3074 ( .A1(n423), .A2(n304), .ZN(\ab[13][12] ) );
  NOR2_X1 U3075 ( .A1(n425), .A2(n304), .ZN(\ab[13][11] ) );
  NOR2_X1 U3076 ( .A1(n477), .A2(n304), .ZN(\ab[13][10] ) );
  NOR2_X1 U3077 ( .A1(n480), .A2(n304), .ZN(\ab[13][0] ) );
  NOR2_X1 U3078 ( .A1(n428), .A2(n306), .ZN(\ab[12][9] ) );
  NOR2_X1 U3079 ( .A1(n431), .A2(n306), .ZN(\ab[12][8] ) );
  NOR2_X1 U3080 ( .A1(n432), .A2(n306), .ZN(\ab[12][7] ) );
  NOR2_X1 U3081 ( .A1(n434), .A2(n306), .ZN(\ab[12][6] ) );
  NOR2_X1 U3082 ( .A1(n436), .A2(n306), .ZN(\ab[12][5] ) );
  NOR2_X1 U3083 ( .A1(n336), .A2(n306), .ZN(\ab[12][52] ) );
  NOR2_X1 U3084 ( .A1(n339), .A2(n306), .ZN(\ab[12][51] ) );
  NOR2_X1 U3085 ( .A1(n341), .A2(n306), .ZN(\ab[12][50] ) );
  NOR2_X1 U3086 ( .A1(n438), .A2(n306), .ZN(\ab[12][4] ) );
  NOR2_X1 U3087 ( .A1(n344), .A2(n307), .ZN(\ab[12][49] ) );
  NOR2_X1 U3088 ( .A1(n346), .A2(n307), .ZN(\ab[12][48] ) );
  NOR2_X1 U3089 ( .A1(n348), .A2(n307), .ZN(\ab[12][47] ) );
  NOR2_X1 U3090 ( .A1(n350), .A2(n307), .ZN(\ab[12][46] ) );
  NOR2_X1 U3091 ( .A1(n352), .A2(n307), .ZN(\ab[12][45] ) );
  NOR2_X1 U3092 ( .A1(n354), .A2(n307), .ZN(\ab[12][44] ) );
  NOR2_X1 U3093 ( .A1(n357), .A2(n307), .ZN(\ab[12][43] ) );
  NOR2_X1 U3094 ( .A1(n359), .A2(n307), .ZN(\ab[12][42] ) );
  NOR2_X1 U3095 ( .A1(n362), .A2(n307), .ZN(\ab[12][41] ) );
  NOR2_X1 U3096 ( .A1(n364), .A2(n307), .ZN(\ab[12][40] ) );
  NOR2_X1 U3097 ( .A1(n441), .A2(n307), .ZN(\ab[12][3] ) );
  NOR2_X1 U3098 ( .A1(n366), .A2(n307), .ZN(\ab[12][39] ) );
  NOR2_X1 U3099 ( .A1(n367), .A2(n307), .ZN(\ab[12][38] ) );
  NOR2_X1 U3100 ( .A1(n371), .A2(n307), .ZN(\ab[12][37] ) );
  NOR2_X1 U3101 ( .A1(n474), .A2(n307), .ZN(\ab[12][36] ) );
  NOR2_X1 U3102 ( .A1(n374), .A2(n306), .ZN(\ab[12][35] ) );
  NOR2_X1 U3103 ( .A1(n376), .A2(n306), .ZN(\ab[12][34] ) );
  NOR2_X1 U3104 ( .A1(n378), .A2(n306), .ZN(\ab[12][33] ) );
  NOR2_X1 U3105 ( .A1(n380), .A2(n306), .ZN(\ab[12][32] ) );
  NOR2_X1 U3106 ( .A1(n382), .A2(n306), .ZN(\ab[12][31] ) );
  NOR2_X1 U3107 ( .A1(n384), .A2(n306), .ZN(\ab[12][30] ) );
  NOR2_X1 U3108 ( .A1(n479), .A2(n306), .ZN(\ab[12][2] ) );
  NOR2_X1 U3109 ( .A1(n385), .A2(n306), .ZN(\ab[12][29] ) );
  NOR2_X1 U3110 ( .A1(n388), .A2(n306), .ZN(\ab[12][28] ) );
  NOR2_X1 U3111 ( .A1(n389), .A2(n306), .ZN(\ab[12][27] ) );
  NOR2_X1 U3112 ( .A1(n391), .A2(n306), .ZN(\ab[12][26] ) );
  NOR2_X1 U3113 ( .A1(n393), .A2(n306), .ZN(\ab[12][25] ) );
  NOR2_X1 U3114 ( .A1(n395), .A2(n306), .ZN(\ab[12][24] ) );
  NOR2_X1 U3115 ( .A1(n397), .A2(n306), .ZN(\ab[12][23] ) );
  NOR2_X1 U3116 ( .A1(n399), .A2(n306), .ZN(\ab[12][22] ) );
  NOR2_X1 U3117 ( .A1(n401), .A2(n306), .ZN(\ab[12][21] ) );
  NOR2_X1 U3118 ( .A1(n403), .A2(n306), .ZN(\ab[12][20] ) );
  NOR2_X1 U3119 ( .A1(n443), .A2(n306), .ZN(\ab[12][1] ) );
  NOR2_X1 U3120 ( .A1(n405), .A2(n306), .ZN(\ab[12][19] ) );
  NOR2_X1 U3121 ( .A1(n407), .A2(n306), .ZN(\ab[12][18] ) );
  NOR2_X1 U3122 ( .A1(n409), .A2(n306), .ZN(\ab[12][17] ) );
  NOR2_X1 U3123 ( .A1(n411), .A2(n306), .ZN(\ab[12][16] ) );
  NOR2_X1 U3124 ( .A1(n414), .A2(n306), .ZN(\ab[12][15] ) );
  NOR2_X1 U3125 ( .A1(n417), .A2(n306), .ZN(\ab[12][14] ) );
  NOR2_X1 U3126 ( .A1(n420), .A2(n306), .ZN(\ab[12][13] ) );
  NOR2_X1 U3127 ( .A1(n423), .A2(n306), .ZN(\ab[12][12] ) );
  NOR2_X1 U3128 ( .A1(n426), .A2(n306), .ZN(\ab[12][11] ) );
  NOR2_X1 U3129 ( .A1(n427), .A2(n306), .ZN(\ab[12][10] ) );
  NOR2_X1 U3130 ( .A1(n480), .A2(n306), .ZN(\ab[12][0] ) );
  NOR2_X1 U3131 ( .A1(n428), .A2(n308), .ZN(\ab[11][9] ) );
  NOR2_X1 U3132 ( .A1(n431), .A2(n308), .ZN(\ab[11][8] ) );
  NOR2_X1 U3133 ( .A1(n432), .A2(n308), .ZN(\ab[11][7] ) );
  NOR2_X1 U3134 ( .A1(n434), .A2(n308), .ZN(\ab[11][6] ) );
  NOR2_X1 U3135 ( .A1(n436), .A2(n308), .ZN(\ab[11][5] ) );
  NOR2_X1 U3136 ( .A1(n336), .A2(n308), .ZN(\ab[11][52] ) );
  NOR2_X1 U3137 ( .A1(n339), .A2(n308), .ZN(\ab[11][51] ) );
  NOR2_X1 U3138 ( .A1(n341), .A2(n308), .ZN(\ab[11][50] ) );
  NOR2_X1 U3139 ( .A1(n438), .A2(n308), .ZN(\ab[11][4] ) );
  NOR2_X1 U3140 ( .A1(n344), .A2(n308), .ZN(\ab[11][49] ) );
  NOR2_X1 U3141 ( .A1(n345), .A2(n470), .ZN(\ab[11][48] ) );
  NOR2_X1 U3142 ( .A1(n347), .A2(n308), .ZN(\ab[11][47] ) );
  NOR2_X1 U3143 ( .A1(n349), .A2(n308), .ZN(\ab[11][46] ) );
  NOR2_X1 U3144 ( .A1(n351), .A2(n470), .ZN(\ab[11][45] ) );
  NOR2_X1 U3145 ( .A1(n354), .A2(n470), .ZN(\ab[11][44] ) );
  NOR2_X1 U3146 ( .A1(n357), .A2(n470), .ZN(\ab[11][43] ) );
  NOR2_X1 U3147 ( .A1(n359), .A2(n470), .ZN(\ab[11][42] ) );
  NOR2_X1 U3148 ( .A1(n361), .A2(n470), .ZN(\ab[11][41] ) );
  NOR2_X1 U3149 ( .A1(n363), .A2(n470), .ZN(\ab[11][40] ) );
  NOR2_X1 U3150 ( .A1(n441), .A2(n470), .ZN(\ab[11][3] ) );
  NOR2_X1 U3151 ( .A1(n365), .A2(n470), .ZN(\ab[11][39] ) );
  NOR2_X1 U3152 ( .A1(n367), .A2(n470), .ZN(\ab[11][38] ) );
  NOR2_X1 U3153 ( .A1(n371), .A2(n308), .ZN(\ab[11][37] ) );
  NOR2_X1 U3154 ( .A1(n372), .A2(n308), .ZN(\ab[11][36] ) );
  NOR2_X1 U3155 ( .A1(n373), .A2(n308), .ZN(\ab[11][35] ) );
  NOR2_X1 U3156 ( .A1(n375), .A2(n308), .ZN(\ab[11][34] ) );
  NOR2_X1 U3157 ( .A1(n377), .A2(n470), .ZN(\ab[11][33] ) );
  NOR2_X1 U3158 ( .A1(n379), .A2(n308), .ZN(\ab[11][32] ) );
  NOR2_X1 U3159 ( .A1(n381), .A2(n470), .ZN(\ab[11][31] ) );
  NOR2_X1 U3160 ( .A1(n383), .A2(n470), .ZN(\ab[11][30] ) );
  NOR2_X1 U3161 ( .A1(n479), .A2(n470), .ZN(\ab[11][2] ) );
  NOR2_X1 U3162 ( .A1(n385), .A2(n308), .ZN(\ab[11][29] ) );
  NOR2_X1 U3163 ( .A1(n388), .A2(n308), .ZN(\ab[11][28] ) );
  NOR2_X1 U3164 ( .A1(n389), .A2(n308), .ZN(\ab[11][27] ) );
  NOR2_X1 U3165 ( .A1(n391), .A2(n308), .ZN(\ab[11][26] ) );
  NOR2_X1 U3166 ( .A1(n393), .A2(n308), .ZN(\ab[11][25] ) );
  NOR2_X1 U3167 ( .A1(n395), .A2(n308), .ZN(\ab[11][24] ) );
  NOR2_X1 U3168 ( .A1(n397), .A2(n308), .ZN(\ab[11][23] ) );
  NOR2_X1 U3169 ( .A1(n399), .A2(n308), .ZN(\ab[11][22] ) );
  NOR2_X1 U3170 ( .A1(n401), .A2(n308), .ZN(\ab[11][21] ) );
  NOR2_X1 U3171 ( .A1(n475), .A2(n308), .ZN(\ab[11][20] ) );
  NOR2_X1 U3172 ( .A1(n443), .A2(n308), .ZN(\ab[11][1] ) );
  NOR2_X1 U3173 ( .A1(n405), .A2(n308), .ZN(\ab[11][19] ) );
  NOR2_X1 U3174 ( .A1(n407), .A2(n308), .ZN(\ab[11][18] ) );
  NOR2_X1 U3175 ( .A1(n409), .A2(n308), .ZN(\ab[11][17] ) );
  NOR2_X1 U3176 ( .A1(n411), .A2(n308), .ZN(\ab[11][16] ) );
  NOR2_X1 U3177 ( .A1(n414), .A2(n308), .ZN(\ab[11][15] ) );
  NOR2_X1 U3178 ( .A1(n417), .A2(n308), .ZN(\ab[11][14] ) );
  NOR2_X1 U3179 ( .A1(n420), .A2(n308), .ZN(\ab[11][13] ) );
  NOR2_X1 U3180 ( .A1(n423), .A2(n308), .ZN(\ab[11][12] ) );
  NOR2_X1 U3181 ( .A1(n426), .A2(n308), .ZN(\ab[11][11] ) );
  NOR2_X1 U3182 ( .A1(n477), .A2(n308), .ZN(\ab[11][10] ) );
  NOR2_X1 U3183 ( .A1(n446), .A2(n308), .ZN(\ab[11][0] ) );
  NOR2_X1 U3184 ( .A1(n429), .A2(n309), .ZN(\ab[10][9] ) );
  NOR2_X1 U3185 ( .A1(n431), .A2(n309), .ZN(\ab[10][8] ) );
  NOR2_X1 U3186 ( .A1(n433), .A2(n309), .ZN(\ab[10][7] ) );
  NOR2_X1 U3187 ( .A1(n434), .A2(n309), .ZN(\ab[10][6] ) );
  NOR2_X1 U3188 ( .A1(n436), .A2(n309), .ZN(\ab[10][5] ) );
  NOR2_X1 U3189 ( .A1(n336), .A2(n309), .ZN(\ab[10][52] ) );
  NOR2_X1 U3190 ( .A1(n339), .A2(n309), .ZN(\ab[10][51] ) );
  NOR2_X1 U3191 ( .A1(n341), .A2(n309), .ZN(\ab[10][50] ) );
  NOR2_X1 U3192 ( .A1(n438), .A2(n309), .ZN(\ab[10][4] ) );
  NOR2_X1 U3193 ( .A1(n344), .A2(n309), .ZN(\ab[10][49] ) );
  NOR2_X1 U3194 ( .A1(n346), .A2(n471), .ZN(\ab[10][48] ) );
  NOR2_X1 U3195 ( .A1(n348), .A2(n309), .ZN(\ab[10][47] ) );
  NOR2_X1 U3196 ( .A1(n350), .A2(n471), .ZN(\ab[10][46] ) );
  NOR2_X1 U3197 ( .A1(n352), .A2(n471), .ZN(\ab[10][45] ) );
  NOR2_X1 U3198 ( .A1(n354), .A2(n471), .ZN(\ab[10][44] ) );
  NOR2_X1 U3199 ( .A1(n357), .A2(n471), .ZN(\ab[10][43] ) );
  NOR2_X1 U3200 ( .A1(n359), .A2(n471), .ZN(\ab[10][42] ) );
  NOR2_X1 U3201 ( .A1(n362), .A2(n471), .ZN(\ab[10][41] ) );
  NOR2_X1 U3202 ( .A1(n364), .A2(n471), .ZN(\ab[10][40] ) );
  NOR2_X1 U3203 ( .A1(n441), .A2(n471), .ZN(\ab[10][3] ) );
  NOR2_X1 U3204 ( .A1(n366), .A2(n471), .ZN(\ab[10][39] ) );
  NOR2_X1 U3205 ( .A1(n367), .A2(n309), .ZN(\ab[10][38] ) );
  NOR2_X1 U3206 ( .A1(n371), .A2(n309), .ZN(\ab[10][37] ) );
  NOR2_X1 U3207 ( .A1(n474), .A2(n309), .ZN(\ab[10][36] ) );
  NOR2_X1 U3208 ( .A1(n374), .A2(n471), .ZN(\ab[10][35] ) );
  NOR2_X1 U3209 ( .A1(n376), .A2(n309), .ZN(\ab[10][34] ) );
  NOR2_X1 U3210 ( .A1(n378), .A2(n471), .ZN(\ab[10][33] ) );
  NOR2_X1 U3211 ( .A1(n380), .A2(n471), .ZN(\ab[10][32] ) );
  NOR2_X1 U3212 ( .A1(n382), .A2(n309), .ZN(\ab[10][31] ) );
  NOR2_X1 U3213 ( .A1(n384), .A2(n471), .ZN(\ab[10][30] ) );
  NOR2_X1 U3214 ( .A1(n479), .A2(n471), .ZN(\ab[10][2] ) );
  NOR2_X1 U3215 ( .A1(n385), .A2(n309), .ZN(\ab[10][29] ) );
  NOR2_X1 U3216 ( .A1(n388), .A2(n309), .ZN(\ab[10][28] ) );
  NOR2_X1 U3217 ( .A1(n389), .A2(n309), .ZN(\ab[10][27] ) );
  NOR2_X1 U3218 ( .A1(n391), .A2(n309), .ZN(\ab[10][26] ) );
  NOR2_X1 U3219 ( .A1(n393), .A2(n309), .ZN(\ab[10][25] ) );
  NOR2_X1 U3220 ( .A1(n395), .A2(n309), .ZN(\ab[10][24] ) );
  NOR2_X1 U3221 ( .A1(n397), .A2(n309), .ZN(\ab[10][23] ) );
  NOR2_X1 U3222 ( .A1(n399), .A2(n309), .ZN(\ab[10][22] ) );
  NOR2_X1 U3223 ( .A1(n401), .A2(n309), .ZN(\ab[10][21] ) );
  NOR2_X1 U3224 ( .A1(n403), .A2(n309), .ZN(\ab[10][20] ) );
  NOR2_X1 U3225 ( .A1(n443), .A2(n309), .ZN(\ab[10][1] ) );
  NOR2_X1 U3226 ( .A1(n405), .A2(n309), .ZN(\ab[10][19] ) );
  NOR2_X1 U3227 ( .A1(n407), .A2(n309), .ZN(\ab[10][18] ) );
  NOR2_X1 U3228 ( .A1(n408), .A2(n309), .ZN(\ab[10][17] ) );
  NOR2_X1 U3229 ( .A1(n411), .A2(n309), .ZN(\ab[10][16] ) );
  NOR2_X1 U3230 ( .A1(n414), .A2(n309), .ZN(\ab[10][15] ) );
  NOR2_X1 U3231 ( .A1(n417), .A2(n309), .ZN(\ab[10][14] ) );
  NOR2_X1 U3232 ( .A1(n420), .A2(n309), .ZN(\ab[10][13] ) );
  NOR2_X1 U3233 ( .A1(n423), .A2(n309), .ZN(\ab[10][12] ) );
  NOR2_X1 U3234 ( .A1(n425), .A2(n309), .ZN(\ab[10][11] ) );
  NOR2_X1 U3235 ( .A1(n427), .A2(n309), .ZN(\ab[10][10] ) );
  NOR2_X1 U3236 ( .A1(n480), .A2(n309), .ZN(\ab[10][0] ) );
  NOR2_X1 U3237 ( .A1(n428), .A2(n334), .ZN(\ab[0][9] ) );
  NOR2_X1 U3238 ( .A1(n430), .A2(n333), .ZN(\ab[0][8] ) );
  NOR2_X1 U3239 ( .A1(n432), .A2(n335), .ZN(\ab[0][7] ) );
  NOR2_X1 U3240 ( .A1(n434), .A2(n334), .ZN(\ab[0][6] ) );
  NOR2_X1 U3241 ( .A1(n436), .A2(n333), .ZN(\ab[0][5] ) );
  NOR2_X1 U3242 ( .A1(n336), .A2(n335), .ZN(\ab[0][52] ) );
  NOR2_X1 U3243 ( .A1(n338), .A2(n334), .ZN(\ab[0][51] ) );
  NOR2_X1 U3244 ( .A1(n342), .A2(n333), .ZN(\ab[0][50] ) );
  NOR2_X1 U3245 ( .A1(n438), .A2(n335), .ZN(\ab[0][4] ) );
  NOR2_X1 U3246 ( .A1(n343), .A2(n334), .ZN(\ab[0][49] ) );
  NOR2_X1 U3247 ( .A1(n346), .A2(n334), .ZN(\ab[0][48] ) );
  NOR2_X1 U3248 ( .A1(n348), .A2(n334), .ZN(\ab[0][47] ) );
  NOR2_X1 U3249 ( .A1(n350), .A2(n334), .ZN(\ab[0][46] ) );
  NOR2_X1 U3250 ( .A1(n352), .A2(n334), .ZN(\ab[0][45] ) );
  NOR2_X1 U3251 ( .A1(n355), .A2(n334), .ZN(\ab[0][44] ) );
  NOR2_X1 U3252 ( .A1(n356), .A2(n334), .ZN(\ab[0][43] ) );
  NOR2_X1 U3253 ( .A1(n360), .A2(n334), .ZN(\ab[0][42] ) );
  NOR2_X1 U3254 ( .A1(n362), .A2(n334), .ZN(\ab[0][41] ) );
  NOR2_X1 U3255 ( .A1(n364), .A2(n334), .ZN(\ab[0][40] ) );
  NOR2_X1 U3256 ( .A1(n478), .A2(n334), .ZN(\ab[0][3] ) );
  NOR2_X1 U3257 ( .A1(n366), .A2(n333), .ZN(\ab[0][39] ) );
  NOR2_X1 U3258 ( .A1(n368), .A2(n333), .ZN(\ab[0][38] ) );
  NOR2_X1 U3259 ( .A1(n370), .A2(n333), .ZN(\ab[0][37] ) );
  NOR2_X1 U3260 ( .A1(n372), .A2(n333), .ZN(\ab[0][36] ) );
  NOR2_X1 U3261 ( .A1(n374), .A2(n333), .ZN(\ab[0][35] ) );
  NOR2_X1 U3262 ( .A1(n376), .A2(n333), .ZN(\ab[0][34] ) );
  NOR2_X1 U3263 ( .A1(n378), .A2(n333), .ZN(\ab[0][33] ) );
  NOR2_X1 U3264 ( .A1(n379), .A2(n333), .ZN(\ab[0][32] ) );
  NOR2_X1 U3265 ( .A1(n382), .A2(n333), .ZN(\ab[0][31] ) );
  NOR2_X1 U3266 ( .A1(n384), .A2(n333), .ZN(\ab[0][30] ) );
  NOR2_X1 U3267 ( .A1(n442), .A2(n333), .ZN(\ab[0][2] ) );
  NOR2_X1 U3268 ( .A1(n386), .A2(n335), .ZN(\ab[0][29] ) );
  NOR2_X1 U3269 ( .A1(n387), .A2(n335), .ZN(\ab[0][28] ) );
  NOR2_X1 U3270 ( .A1(n390), .A2(n335), .ZN(\ab[0][27] ) );
  NOR2_X1 U3271 ( .A1(n392), .A2(n333), .ZN(\ab[0][26] ) );
  NOR2_X1 U3272 ( .A1(n394), .A2(n335), .ZN(\ab[0][25] ) );
  NOR2_X1 U3273 ( .A1(n396), .A2(n333), .ZN(\ab[0][24] ) );
  NOR2_X1 U3274 ( .A1(n398), .A2(n335), .ZN(\ab[0][23] ) );
  NOR2_X1 U3275 ( .A1(n400), .A2(n335), .ZN(\ab[0][22] ) );
  NOR2_X1 U3276 ( .A1(n402), .A2(n333), .ZN(\ab[0][21] ) );
  NOR2_X1 U3277 ( .A1(n475), .A2(n335), .ZN(\ab[0][20] ) );
  NOR2_X1 U3278 ( .A1(n443), .A2(n334), .ZN(\ab[0][1] ) );
  NOR2_X1 U3279 ( .A1(n404), .A2(n333), .ZN(\ab[0][19] ) );
  NOR2_X1 U3280 ( .A1(n476), .A2(n335), .ZN(\ab[0][18] ) );
  NOR2_X1 U3281 ( .A1(n409), .A2(n333), .ZN(\ab[0][17] ) );
  NOR2_X1 U3282 ( .A1(n412), .A2(n335), .ZN(\ab[0][16] ) );
  NOR2_X1 U3283 ( .A1(n415), .A2(n335), .ZN(\ab[0][15] ) );
  NOR2_X1 U3284 ( .A1(n418), .A2(n333), .ZN(\ab[0][14] ) );
  NOR2_X1 U3285 ( .A1(n421), .A2(n335), .ZN(\ab[0][13] ) );
  NOR2_X1 U3286 ( .A1(n424), .A2(n334), .ZN(\ab[0][12] ) );
  NOR2_X1 U3287 ( .A1(n426), .A2(n333), .ZN(\ab[0][11] ) );
  NOR2_X1 U3288 ( .A1(n427), .A2(n335), .ZN(\ab[0][10] ) );
  NOR2_X1 U3289 ( .A1(n446), .A2(n333), .ZN(PRODUCT[0]) );
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
endmodule


module fpu ( clk, rmode, fpu_op, opa, opb, out, inf, snan, qnan, ine, overflow, 
        underflow, zero, div_by_zero );
  input [1:0] rmode;
  input [2:0] fpu_op;
<<<<<<< HEAD
  input [15:0] opa;
  input [15:0] opb;
  output [15:0] out;
  input clk;
  output inf, snan, qnan, ine, overflow, underflow, zero, div_by_zero;
  wire   snan_d, opa_nan, opb_nan, opa_00, opb_00, opa_inf, opb_inf, opa_dn,
         opb_dn, sign_fasu, nan_sign_d, result_zero_sign_d, fasu_op,
         sign_fasu_r, sign_mul, sign_exe, inf_mul, sign_mul_r, sign_exe_r, N34,
         N44, N56, N65, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77,
         N96, N97, N98, N99, N100, N106, N110, N111, N112, N113, N114, N115,
         N116, \fract_i2f[7] , N138, N139, N140, N141, N150, N151, N179, N180,
         N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191,
         N192, N193, N194, N195, N196, opas_r1, opas_r2, sign, N216,
         fasu_op_r1, N220, N221, N222, N223, N224, N225, N226, N227, N228,
         N229, N230, N231, N232, N233, N234, N254, N278, N281, N283, N285,
         N290, N291, N292, N296, \u0/N17 , \u0/N16 , \u0/expb_00 ,
         \u0/expa_00 , \u0/N11 , \u0/N10 , \u0/N7 , \u0/N6 , \u0/N5 , \u0/N4 ,
         \u0/infb_f_r , \u0/infa_f_r , \u0/expb_ff , \u0/expa_ff , \u1/N133 ,
         \u1/fracta_eq_fractb , \u1/N124 , \u1/fracta_lt_fractb , \u1/N123 ,
         \u1/N122 , \u1/add_r , \u1/signa_r , \u1/sign_d ,
         \u1/adj_op_out_sft[0] , \u1/adj_op_out_sft[1] ,
=======
  input [63:0] opa;
  input [63:0] opb;
  output [63:0] out;
  input clk;
  output inf, snan, qnan, ine, overflow, underflow, zero, div_by_zero;
  wire   inf_d, ind_d, qnan_d, snan_d, opa_nan, opb_nan, opa_00, opb_00,
         opa_inf, opb_inf, opb_dn, sign_fasu, nan_sign_d, result_zero_sign_d,
         fasu_op, sign_fasu_r, sign_mul, sign_exe, inf_mul, sign_mul_r,
         inf_mul_r, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265,
         N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276,
         N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287,
         N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298,
         N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N327,
         N328, N329, N330, N331, N332, N333, N334, N335, N336, N337,
         \fract_div[105] , N340, N343, N344, N345, N346, N347, N348, N349,
         N350, N351, N352, N353, N354, N355, N356, N357, N358, N359, N360,
         N361, N362, N363, N364, N365, N366, N367, N368, N369, N370, N371,
         N372, N373, N374, N375, N376, N377, N378, N379, N380, N381, N382,
         N383, N384, N385, N386, N387, N388, N389, N390, N391, N392, N393,
         N394, N395, N396, N501, N502, N503, N504, N505, N506, N507, N508,
         N509, N510, N511, N512, N513, N514, N515, N516, N517, N518, N519,
         N520, N521, N522, N523, N524, N525, N526, N527, N528, N529, N530,
         N531, N532, N533, N534, N535, N536, N537, N538, N539, N540, N541,
         N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552,
         N553, N554, N555, N556, N557, N710, N711, N712, N713, N714, N715,
         N716, N717, N718, N719, N720, N721, N722, N723, N724, N725, N726,
         N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737,
         N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748,
         N749, N750, N751, N752, N753, N754, N755, N756, N757, N758, N759,
         N760, N761, N762, N763, N764, N765, N766, N767, N768, N769, opas_r1,
         opas_r2, sign, N789, fasu_op_r1, fasu_op_r2, inf_mul2, N793, N794,
         N795, N796, N797, N798, N799, N800, N801, N802, N803, N804, N805,
         N806, N807, N808, N809, N810, N811, N812, N813, N814, N815, N816,
         N817, N818, N819, N820, N821, N822, N823, N824, N825, N826, N827,
         N828, N829, N830, N831, N832, N833, N834, N835, N836, N837, N838,
         N839, N840, N841, N842, N843, N844, N845, N846, N847, N848, N849,
         N850, N851, N852, N853, N854, N855, N875, N889, N899, N902, N904,
         N906, N911, N912, opa_nan_r, N913, N923, \u0/N17 , \u0/N16 ,
         \u0/fractb_00 , \u0/fracta_00 , \u0/expb_00 , \u0/expa_00 , \u0/N11 ,
         \u0/N10 , \u0/N7 , \u0/N6 , \u0/snan_r_b , \u0/N5 , \u0/qnan_r_b ,
         \u0/snan_r_a , \u0/N4 , \u0/qnan_r_a , \u0/infb_f_r , \u0/infa_f_r ,
         \u0/expb_ff , \u0/expa_ff , \u1/N232 , \u1/N229 ,
         \u1/fracta_eq_fractb , \u1/N220 , \u1/fracta_lt_fractb , \u1/N219 ,
         \u1/N218 , \u1/add_r , \u1/signb_r , \u1/signa_r , \u1/sign_d ,
         \u1/fractb_lt_fracta , \u1/adj_op_out_sft[0] , \u1/adj_op_out_sft[1] ,
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
         \u1/adj_op_out_sft[2] , \u1/adj_op_out_sft[3] ,
         \u1/adj_op_out_sft[4] , \u1/adj_op_out_sft[5] ,
         \u1/adj_op_out_sft[6] , \u1/adj_op_out_sft[7] ,
         \u1/adj_op_out_sft[8] , \u1/adj_op_out_sft[9] ,
         \u1/adj_op_out_sft[10] , \u1/adj_op_out_sft[11] ,
         \u1/adj_op_out_sft[12] , \u1/adj_op_out_sft[13] ,
<<<<<<< HEAD
         \u1/exp_diff_sft[0] , \u1/adj_op[9] , \u1/N39 , \u1/N38 , \u1/N37 ,
         \u1/N36 , \u1/N35 , \u2/N73 , \u2/sign_d , \u2/N66 ,
         \u2/exp_ovf_d[0] , \u2/exp_ovf_d[1] , \u2/N44 , \u2/N43 , \u2/N42 ,
         \u2/N41 , \u2/N40 , \u2/N37 , \u2/N34 , \u2/N33 , \u2/N32 , \u2/N31 ,
         \u2/exp_tmp4[0] , \u2/exp_tmp4[1] , \u2/exp_tmp4[2] ,
         \u2/exp_tmp4[3] , \u2/exp_tmp4[4] , \u2/exp_tmp3[1] ,
         \u2/exp_tmp3[2] , \u2/exp_tmp3[3] , \u2/exp_tmp3[4] , \u2/N29 ,
         \u2/N28 , \u2/N27 , \u2/N26 , \u2/N25 , \u2/N23 , \u2/N22 , \u2/N21 ,
         \u2/N20 , \u2/N19 , \u2/N17 , \u2/N16 , \u2/N15 , \u2/N14 , \u2/N13 ,
         \u2/N12 , \u2/N11 , \u2/N10 , \u2/N9 , \u2/N8 , \u2/N7 , \u2/N6 ,
         \u3/N32 , \u3/N31 , \u3/N30 , \u3/N29 , \u3/N28 , \u3/N27 , \u3/N26 ,
         \u3/N25 , \u3/N24 , \u3/N23 , \u3/N22 , \u3/N21 , \u3/N20 , \u3/N19 ,
         \u3/N18 , \u3/N17 , \u3/N16 , \u3/N15 , \u3/N14 , \u3/N13 , \u3/N12 ,
         \u3/N11 , \u3/N10 , \u3/N9 , \u3/N8 , \u3/N7 , \u3/N6 , \u3/N5 ,
         \u3/N4 , \u3/N3 , \u5/N21 , \u5/N20 , \u5/N19 , \u5/N18 , \u5/N17 ,
         \u5/N16 , \u5/N15 , \u5/N14 , \u5/N13 , \u5/N12 , \u5/N11 , \u5/N10 ,
         \u5/N9 , \u5/N8 , \u5/N7 , \u5/N6 , \u5/N5 , \u5/N4 , \u5/N3 ,
         \u5/N2 , \u5/N1 , \u5/N0 , \u6/N23 , \u6/N22 , \u6/N21 , \u6/N20 ,
         \u6/N19 , \u6/N18 , \u6/N17 , \u6/N16 , \u6/N15 , \u6/N14 , \u6/N13 ,
         \u6/N10 , \u6/N9 , \u6/N8 , \u6/N7 , \u6/N6 , \u6/N5 , \u6/N4 ,
         \u6/N3 , \u6/N2 , \u6/N1 , \u6/N0 , \u4/N656 , \u4/N655 , \u4/N653 ,
         \u4/div_exp3[1] , \u4/fi_ldz_mi1[2] , \u4/fi_ldz_mi1[3] , \u4/N433 ,
         \u4/N432 , \u4/N431 , \u4/N430 , \u4/N429 , \u4/N428 , \u4/N427 ,
         \u4/N426 , \u4/N425 , \u4/N424 , \u4/N423 , \u4/N422 , \u4/N421 ,
         \u4/N420 , \u4/N419 , \u4/N418 , \u4/N417 , \u4/N416 , \u4/N415 ,
         \u4/N414 , \u4/N413 , \u4/N412 , \u4/N409 , \u4/N408 , \u4/N407 ,
         \u4/N406 , \u4/N405 , \u4/N404 , \u4/N403 , \u4/N402 , \u4/N401 ,
         \u4/N400 , \u4/N399 , \u4/N398 , \u4/N397 , \u4/N396 , \u4/N395 ,
         \u4/N394 , \u4/N393 , \u4/N392 , \u4/N391 , \u4/N390 , \u4/N389 ,
         \u4/N388 , \u4/N386 , \u4/exp_in_pl1[2] , \u4/exp_in_pl1[3] ,
         \u4/exp_in_pl1[4] , \u4/exp_in_pl1[5] , \u4/f2i_shft[2] ,
         \u4/f2i_shft[3] , \u4/f2i_shft[4] , \u4/div_shft2[0] ,
         \u4/fract_out_pl1[0] , \u4/fract_out_pl1[1] , \u4/fract_out_pl1[2] ,
         \u4/fract_out_pl1[3] , \u4/fract_out_pl1[4] , \u4/fract_out_pl1[5] ,
         \u4/fract_out_pl1[6] , \u4/fract_out_pl1[7] , \u4/fract_out_pl1[8] ,
         \u4/fract_out_pl1[9] , \u4/fract_out_pl1[10] , \u4/exp_next_mi[0] ,
         \u4/exp_next_mi[1] , \u4/exp_next_mi[2] , \u4/exp_next_mi[3] ,
         \u4/exp_next_mi[4] , \u4/exp_next_mi[5] , \u4/fract_out[1] ,
         \u4/fract_out[5] , \u4/exp_out[2] , n845, n851, n872, n888, n1521,
         net10316, \u2/lt_130/A[0] , \u2/lt_130/A[1] , \u2/lt_130/A[2] ,
         \u2/lt_130/A[3] , \u2/gt_140/B[5] , net11677, net11676, net11675,
         net11671, net11670, net11627, net11582, net11576, net11567, net11566,
         net11564, net11562, net11560, net11558, net11555, net11485,
         \u4/sub_409/net10540 , \u2/add_113/A[0] , \u2/add_113/A[1] ,
         \u2/add_113/A[2] , \u2/add_113/A[3] , \u2/add_113/A[4] ,
         \u2/sub_111/carry[2] , \u2/sub_111/carry[3] , \u2/sub_111/carry[4] ,
         \u2/sub_111/carry[5] , \u2/add_111/carry[2] , \u2/add_111/carry[3] ,
         \u2/add_111/carry[4] , \u2/add_111/carry[5] , net15448, net15944,
         net30297, net33278, net60630, net76048, net76254, net76619, net76645,
         net76672, net76926, net77045, net77073, net77161, net77637, net77815,
         net83296, net83361, net83364, net83368, net83402, net83403, net83407,
         net83408, net83414, net83419, net83421, net83423, net83427, net83429,
         net83432, net83438, net83439, net83736, net83747, net83754, net83765,
         net83779, net83780, net83781, net83787, net83791, net83800, net83802,
         net83806, net83807, net83811, net83812, net83820, net83821, net83827,
         net83833, net83836, net83844, net83849, net83853, net83855, net83856,
         net83860, net83861, net83862, net83863, net83864, net83868, net83869,
         net83871, net83874, net83875, net83876, net83878, net83883, net83906,
         net83913, net83925, net83927, net83933, net83934, net83936, net83940,
         net83941, net83942, net83945, net83946, net83950, net83951, net83959,
         net83963, net83967, net83968, net83969, net83971, net83972, net83973,
         net83975, net83987, net83990, net83993, net83994, net83995, net84003,
         net84010, net84012, net84015, net84021, net84024, net84044, net84047,
         net84048, net84050, net84055, net84059, net84060, net84069, net84070,
         net84072, net84073, net84076, net84079, net84080, net84081, net84083,
         net84095, net84096, net84103, net84107, net84115, net84118, net84119,
         net84128, net84133, net84134, net84135, net84136, net84138, net84146,
         net84148, net84149, net84150, net84151, net84157, net84159, net84160,
         net84165, net84166, net84167, net84168, net84169, net84191, net84199,
         net84200, net84211, net84214, net84215, net84216, net84218, net84220,
         net84236, net84249, net84253, net84254, net84263, net84265, net84266,
         net84276, net84277, net84278, net84279, net84280, net84290, net84297,
         net84298, net84299, net84305, net84310, net84312, net84314, net84315,
         net84322, net84326, net84327, net84329, net84332, net84333, net84334,
         net84341, net84343, net84344, net84347, net84352, net84366, net84368,
         net84371, net84373, net84374, net84381, net84398, net84402, net84403,
         net84421, net84445, net84448, net84449, net84450, net84453, net84458,
         net84465, net84468, net84469, net84474, net84475, net84480, net84482,
         net84487, net84488, net84490, net84498, net84500, net84501, net84502,
         net84506, net84511, net84520, net84522, net84523, net84524, net84531,
         net84532, net84548, net84549, net84550, net84551, net84552, net84555,
         net84561, net84564, net84565, net84568, net84571, net84579, net84590,
         net84591, net84595, net84598, net84599, net84600, net84601, net84602,
         net84604, net84605, net84609, net84610, net84611, net84614, net84615,
         net84617, net84619, net84624, net84625, net84626, net84629, net84632,
         net84633, net84637, net84639, net84642, net84643, net84644, net84645,
         net84647, net84648, net84649, net84652, net84655, net84656, net84659,
         net84660, net84661, net84662, net84663, net84664, net84667, net84668,
         net84669, net84672, net84675, net84684, net84702, net84722, net84749,
         net84753, net84754, net84755, net84758, net84761, net84762, net84763,
         net84764, net84765, net84766, net84767, net84768, net84774, net84775,
         net84777, net84778, net84783, net84784, net84810, net84814, net84822,
         net84823, net84839, net84840, net84842, net84847, net84848, net84853,
         net84856, net84858, net84867, net84869, net84870, net84884, net84886,
         net84887, net84890, net84900, net84901, net84906, net84907, net84911,
         net84912, net84915, net84916, net84921, net84953, net84968, net84975,
         net84982, net84983, net84990, net84992, net84995, net84996, net85004,
         net85006, net85010, net85015, net85027, net85030, net85032, net85037,
         net85038, net85039, net85040, net85041, net85043, net85045, net85046,
         net85051, net85059, net85060, net85061, net85067, net85068, net85069,
         net85071, net85076, net85080, net85091, net85093, net85095, net85096,
         net85099, net85103, net85104, net85105, net85111, net85112, net85113,
         net85114, net85115, net85116, net85123, net85124, net85126, net85127,
         net85131, net85136, net85137, net85140, net85141, net85144, net85150,
         net85164, net85168, net85169, net85170, net85171, net85176, net85178,
         net85182, net85191, net85192, net85194, net85195, net85196, net85197,
         net85200, net85203, net85204, net85205, net85206, net85207, net85210,
         net85211, net85212, net85213, net85216, net85220, net85224, net85227,
         net85232, net85234, net85247, net85257, net85263, net85280, net85281,
         net85285, net85292, net85310, net85313, net85316, net85320, net85331,
         net85336, net85351, net85361, net85365, net85369, net85373, net85374,
         net85393, net85676, net85674, net85712, net85710, net85722, net85720,
         net85718, net85716, net85738, net85736, net85732, net85730, net85728,
         net85752, net85748, net85746, net85744, net85778, net85788, net85786,
         net85794, net85790, net85828, net85832, net85842, net85847, net85854,
         net85853, net85974, net85998, net86004, net86006, net86010, net86016,
         net86038, net86037, net86061, net86090, net86096, net86106, net86113,
         net86112, net86125, net86169, net86263, net88287, net88293, net88292,
         net88319, net88421, net88427, net88440, net88500, net88503, net88510,
         net88545, net88566, net88585, net88618, net88695, net88699, net88721,
         net88877, net88896, net88950, net88972, net89029, net89078, net89121,
         net89120, net89129, net89250, net89266, net89314, net89412, net89411,
         net89485, net89537, net89543, net89546, net89624, net89677, net89681,
         net89680, net89679, net89692, net89716, net89741, net89753, net89819,
         net89817, net89863, net89862, net89919, net89924, net89926, net89933,
         net89943, net89948, net89964, net89965, net89975, net89987, net89998,
         net90007, net90026, net90031, net90037, net90047, net90064, net90074,
         net90080, net90115, net90122, net90124, net90126, net90144, net90207,
         net90211, net90210, net90217, net90252, net90268, net90287, net90290,
         net90292, net90299, net90302, net86262, net85081, net91047, net91057,
         net91056, net91059, net91070, net91069, net91075, net91095, net91112,
         net91128, net91159, net91299, net91298, net91325, net91512, net91542,
         net91548, net91555, net83406, net85166, net85160, net85157, net85155,
         net85135, net85125, net85120, net85133, net85107, net84830, net90035,
         net85337, net85335, net85162, net85147, net84910, net91467, net90997,
         net84994, net89447, net89446, net83420, net90072, net85165, net85042,
         net84909, net88895, net84452, net89856, net99868, net99874, net85272,
         net85270, net85265, net85264, net85254, net85253, net85252, net85251,
         net85250, net85189, net85163, net85684, net85261, net85187, net91177,
         net85033, net84984, net84673, net91109, net88551, net85239, net85215,
         net85214, net85177, net85098, net85087, net84503, net85260, net90215,
         net89935, net88605, net86027, net86026, net85290, net85283, net85240,
         net84969, net84960, net84957, net90019, net89300, net88636, net85360,
         net85357, net85159, net85158, net85097, net85089, net85085, net110929,
         net110951, net99862, net85079, net85190, net85188, net85184, net85083,
         net86060, net85317, net76872, net84213, net84071, net83870, net91353,
         net86171, net86015, net84677, net84394, net84393, net84387, net84386,
         net91015, net84882, \u4/fract_out[8] , \u4/fract_out[3] , net84845,
         net84844, net84456, net84110, net85199, net85193, net85185, net85143,
         net85142, net84043, net84033, net84029, net84028, net84026, net85342,
         net86174, net84414, net84075, net85020, net85018, net84974, net85021,
         net84913, net84895, net89073, net84484, net84409, net84401, net84390,
         \u4/fract_out[6] , net84113, net89595, net84553, net84473, net84770,
         net84678, net84573, net84519, net84518, net90110, net88332, net85297,
         net85296, net85186, net85161, net85048, net84030, net84027, net89917,
         net89077, net89076, net86160, net84408, net84385, net84372, net89372,
         net85017, net84967, net84956, net85384, net85248, net85180, net85179,
         net85084, net85082, net85077, net84757, net76352, net84584, net85975,
         net85678, net85387, net85349, net85181, net85174, net85128, net85108,
         net84301, net91511, net91404, net84576, net84575, net84574, net88374,
         net84206, net84204, net84202, net84201, net84085, net84074, net91375,
         net89842, net89224, net89055, net89054, net85831, net84963, net84950,
         net84948, net99831, net84651, net84554, net84483, net89615, net86165,
         net85827, net83974, net83813, net84854, net84846, net84566, net84064,
         net84052, net84051, net84025, net83819, \u4/fract_out[7] ,
         \u4/fract_out[4] , net91150, net84908, net84836, net84829, net84811,
         net84808, net84769, net84586, net84572, net84570, net84569, net89664,
         net89663, net84683, net84679, net84676, net84674, net84472, net84471,
         net84451, net86067, net83394, net83393, net84606, net83395, net89736,
         net89658, net89657, net88646, net83398, \u4/exp_out[4] , net85742,
         net85740, net85726, net85724, net85323, net85028, net84588, net91144,
         net90079, net85846, net85756, net85754, net84658, net84657, net84654,
         net84014, \u4/f2i_shft[1] , net83417, net83416, net83392, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1539, n1541, n1543, n1546, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1718,
         n1719, n1720, n1721, n1722, n1723, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1736, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1969, n1970, n1971, n1972, n1973, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323;
  wire   [15:10] opa_r;
  wire   [15:10] opb_r;
=======
         \u1/adj_op_out_sft[14] , \u1/adj_op_out_sft[15] ,
         \u1/adj_op_out_sft[16] , \u1/adj_op_out_sft[17] ,
         \u1/adj_op_out_sft[18] , \u1/adj_op_out_sft[19] ,
         \u1/adj_op_out_sft[20] , \u1/adj_op_out_sft[21] ,
         \u1/adj_op_out_sft[22] , \u1/adj_op_out_sft[23] ,
         \u1/adj_op_out_sft[24] , \u1/adj_op_out_sft[25] ,
         \u1/adj_op_out_sft[26] , \u1/adj_op_out_sft[27] ,
         \u1/adj_op_out_sft[28] , \u1/adj_op_out_sft[29] ,
         \u1/adj_op_out_sft[30] , \u1/adj_op_out_sft[31] ,
         \u1/adj_op_out_sft[32] , \u1/adj_op_out_sft[33] ,
         \u1/adj_op_out_sft[34] , \u1/adj_op_out_sft[35] ,
         \u1/adj_op_out_sft[36] , \u1/adj_op_out_sft[37] ,
         \u1/adj_op_out_sft[38] , \u1/adj_op_out_sft[39] ,
         \u1/adj_op_out_sft[40] , \u1/adj_op_out_sft[41] ,
         \u1/adj_op_out_sft[42] , \u1/adj_op_out_sft[43] ,
         \u1/adj_op_out_sft[44] , \u1/adj_op_out_sft[45] ,
         \u1/adj_op_out_sft[46] , \u1/adj_op_out_sft[47] ,
         \u1/adj_op_out_sft[48] , \u1/adj_op_out_sft[49] ,
         \u1/adj_op_out_sft[50] , \u1/adj_op_out_sft[51] ,
         \u1/adj_op_out_sft[52] , \u1/adj_op_out_sft[53] ,
         \u1/adj_op_out_sft[54] , \u1/adj_op_out_sft[55] , \u1/exp_lt_27 ,
         \u1/adj_op[0] , \u1/adj_op[3] , \u1/adj_op[10] , \u1/adj_op[11] ,
         \u1/adj_op[15] , \u1/adj_op[16] , \u1/adj_op[17] , \u1/adj_op[20] ,
         \u1/adj_op[21] , \u1/adj_op[22] , \u1/adj_op[27] , \u1/adj_op[28] ,
         \u1/adj_op[32] , \u1/adj_op[36] , \u1/adj_op[37] , \u1/adj_op[38] ,
         \u1/adj_op[42] , \u1/adj_op[44] , \u1/adj_op[51] , \u1/N62 , \u1/N61 ,
         \u1/N60 , \u1/N59 , \u1/N58 , \u1/N57 , \u1/N56 , \u1/N55 , \u1/N54 ,
         \u1/N53 , \u1/N52 , \u1/N49 , \u1/exp_diff[0] , \u1/exp_diff[1] ,
         \u1/exp_diff[2] , \u1/exp_diff[3] , \u1/exp_diff[4] ,
         \u1/exp_diff[5] , \u1/exp_diff[6] , \u1/exp_diff[7] ,
         \u1/exp_diff[8] , \u1/exp_diff[9] , \u1/exp_diff[10] , \u1/N46 ,
         \u1/exp_large[0] , \u1/exp_large[1] , \u1/exp_large[2] ,
         \u1/exp_large[3] , \u1/exp_large[4] , \u1/exp_large[5] ,
         \u1/exp_large[6] , \u1/exp_large[7] , \u1/exp_large[10] ,
         \u1/expa_lt_expb , \u2/N157 , \u2/N121 , \u2/sign_d , \u2/N114 ,
         \u2/N113 , \u2/N111 , \u2/exp_ovf_d[0] , \u2/exp_ovf_d[1] , \u2/N86 ,
         \u2/N85 , \u2/N84 , \u2/N83 , \u2/N82 , \u2/N81 , \u2/N80 , \u2/N79 ,
         \u2/N78 , \u2/N77 , \u2/N76 , \u2/N75 , \u2/N74 , \u2/N73 , \u2/N72 ,
         \u2/N71 , \u2/N70 , \u2/N69 , \u2/N68 , \u2/N67 , \u2/N66 , \u2/N64 ,
         \u2/N63 , \u2/N62 , \u2/N61 , \u2/N60 , \u2/N59 , \u2/N58 , \u2/N57 ,
         \u2/N56 , \u2/N55 , \u2/N54 , \u2/exp_tmp4[1] , \u2/exp_tmp4[2] ,
         \u2/exp_tmp4[3] , \u2/exp_tmp4[4] , \u2/exp_tmp4[10] ,
         \u2/exp_tmp3[0] , \u2/exp_tmp3[1] , \u2/exp_tmp3[2] ,
         \u2/exp_tmp3[3] , \u2/exp_tmp3[4] , \u2/exp_tmp3[5] ,
         \u2/exp_tmp3[6] , \u2/exp_tmp3[7] , \u2/exp_tmp3[8] ,
         \u2/exp_tmp3[9] , \u2/exp_tmp3[10] , \u2/N53 , \u2/N52 , \u2/N51 ,
         \u2/N50 , \u2/N49 , \u2/N48 , \u2/N47 , \u2/N46 , \u2/N45 , \u2/N44 ,
         \u2/N43 , \u2/N41 , \u2/N40 , \u2/N39 , \u2/N38 , \u2/N37 , \u2/N36 ,
         \u2/N35 , \u2/N34 , \u2/N33 , \u2/N32 , \u2/N31 , \u2/exp_tmp1[1] ,
         \u2/exp_tmp1[2] , \u2/exp_tmp1[3] , \u2/exp_tmp1[4] , \u2/N29 ,
         \u2/N28 , \u2/N27 , \u2/N26 , \u2/N25 , \u2/N24 , \u2/N23 , \u2/N22 ,
         \u2/N21 , \u2/N20 , \u2/N19 , \u2/N18 , \u2/N17 , \u2/N16 , \u2/N15 ,
         \u2/N14 , \u2/N13 , \u2/N12 , \u2/N11 , \u2/N10 , \u2/N9 , \u2/N8 ,
         \u2/N7 , \u2/N6 , \u3/N116 , \u3/N115 , \u3/N114 , \u3/N113 ,
         \u3/N112 , \u3/N111 , \u3/N110 , \u3/N109 , \u3/N108 , \u3/N107 ,
         \u3/N106 , \u3/N105 , \u3/N104 , \u3/N103 , \u3/N102 , \u3/N101 ,
         \u3/N100 , \u3/N99 , \u3/N98 , \u3/N97 , \u3/N96 , \u3/N95 , \u3/N94 ,
         \u3/N93 , \u3/N92 , \u3/N91 , \u3/N90 , \u3/N89 , \u3/N88 , \u3/N87 ,
         \u3/N86 , \u3/N85 , \u3/N84 , \u3/N83 , \u3/N82 , \u3/N81 , \u3/N80 ,
         \u3/N79 , \u3/N78 , \u3/N77 , \u3/N76 , \u3/N75 , \u3/N74 , \u3/N73 ,
         \u3/N72 , \u3/N71 , \u3/N70 , \u3/N69 , \u3/N68 , \u3/N67 , \u3/N66 ,
         \u3/N65 , \u3/N64 , \u3/N63 , \u3/N62 , \u3/N61 , \u3/N60 , \u3/N59 ,
         \u3/N58 , \u3/N57 , \u3/N56 , \u3/N55 , \u3/N54 , \u3/N53 , \u3/N52 ,
         \u3/N51 , \u3/N50 , \u3/N49 , \u3/N48 , \u3/N47 , \u3/N46 , \u3/N45 ,
         \u3/N44 , \u3/N43 , \u3/N42 , \u3/N41 , \u3/N40 , \u3/N39 , \u3/N38 ,
         \u3/N37 , \u3/N36 , \u3/N35 , \u3/N34 , \u3/N33 , \u3/N32 , \u3/N31 ,
         \u3/N30 , \u3/N29 , \u3/N28 , \u3/N27 , \u3/N26 , \u3/N25 , \u3/N24 ,
         \u3/N23 , \u3/N22 , \u3/N21 , \u3/N20 , \u3/N19 , \u3/N18 , \u3/N17 ,
         \u3/N16 , \u3/N15 , \u3/N14 , \u3/N13 , \u3/N12 , \u3/N11 , \u3/N10 ,
         \u3/N9 , \u3/N8 , \u3/N7 , \u3/N6 , \u3/N5 , \u3/N4 , \u3/N3 ,
         \u5/N105 , \u5/N104 , \u5/N103 , \u5/N102 , \u5/N101 , \u5/N100 ,
         \u5/N99 , \u5/N98 , \u5/N97 , \u5/N96 , \u5/N95 , \u5/N94 , \u5/N93 ,
         \u5/N92 , \u5/N91 , \u5/N90 , \u5/N89 , \u5/N88 , \u5/N87 , \u5/N86 ,
         \u5/N85 , \u5/N84 , \u5/N83 , \u5/N82 , \u5/N81 , \u5/N80 , \u5/N79 ,
         \u5/N78 , \u5/N77 , \u5/N76 , \u5/N75 , \u5/N74 , \u5/N73 , \u5/N72 ,
         \u5/N71 , \u5/N70 , \u5/N69 , \u5/N68 , \u5/N67 , \u5/N66 , \u5/N65 ,
         \u5/N64 , \u5/N63 , \u5/N62 , \u5/N61 , \u5/N60 , \u5/N59 , \u5/N58 ,
         \u5/N57 , \u5/N56 , \u5/N55 , \u5/N54 , \u5/N53 , \u5/N52 , \u5/N51 ,
         \u5/N50 , \u5/N49 , \u5/N48 , \u5/N47 , \u5/N46 , \u5/N45 , \u5/N44 ,
         \u5/N43 , \u5/N42 , \u5/N41 , \u5/N40 , \u5/N39 , \u5/N38 , \u5/N37 ,
         \u5/N36 , \u5/N35 , \u5/N34 , \u5/N33 , \u5/N32 , \u5/N31 , \u5/N30 ,
         \u5/N29 , \u5/N28 , \u5/N27 , \u5/N26 , \u5/N25 , \u5/N24 , \u5/N23 ,
         \u5/N22 , \u5/N21 , \u5/N20 , \u5/N19 , \u5/N18 , \u5/N17 , \u5/N16 ,
         \u5/N15 , \u5/N14 , \u5/N13 , \u5/N12 , \u5/N11 , \u5/N10 , \u5/N9 ,
         \u5/N8 , \u5/N7 , \u5/N6 , \u5/N5 , \u5/N4 , \u5/N3 , \u5/N2 ,
         \u5/N1 , \u5/N0 , \u6/N107 , \u6/N106 , \u6/N105 , \u6/N104 ,
         \u6/N103 , \u6/N102 , \u6/N101 , \u6/N100 , \u6/N99 , \u6/N98 ,
         \u6/N97 , \u6/N96 , \u6/N95 , \u6/N94 , \u6/N93 , \u6/N92 , \u6/N91 ,
         \u6/N90 , \u6/N89 , \u6/N88 , \u6/N87 , \u6/N86 , \u6/N85 , \u6/N84 ,
         \u6/N83 , \u6/N82 , \u6/N81 , \u6/N80 , \u6/N79 , \u6/N78 , \u6/N77 ,
         \u6/N76 , \u6/N75 , \u6/N74 , \u6/N73 , \u6/N72 , \u6/N71 , \u6/N70 ,
         \u6/N69 , \u6/N68 , \u6/N67 , \u6/N66 , \u6/N65 , \u6/N64 , \u6/N63 ,
         \u6/N62 , \u6/N61 , \u6/N60 , \u6/N59 , \u6/N58 , \u6/N57 , \u6/N56 ,
         \u6/N55 , \u6/N52 , \u6/N51 , \u6/N50 , \u6/N49 , \u6/N48 , \u6/N47 ,
         \u6/N46 , \u6/N45 , \u6/N44 , \u6/N43 , \u6/N42 , \u6/N41 , \u6/N40 ,
         \u6/N39 , \u6/N38 , \u6/N37 , \u6/N36 , \u6/N35 , \u6/N34 , \u6/N33 ,
         \u6/N32 , \u6/N31 , \u6/N30 , \u6/N29 , \u6/N28 , \u6/N27 , \u6/N26 ,
         \u6/N25 , \u6/N24 , \u6/N23 , \u6/N22 , \u6/N21 , \u6/N20 , \u6/N19 ,
         \u6/N18 , \u6/N17 , \u6/N16 , \u6/N15 , \u6/N14 , \u6/N13 , \u6/N12 ,
         \u6/N11 , \u6/N10 , \u6/N9 , \u6/N8 , \u6/N7 , \u6/N6 , \u6/N5 ,
         \u6/N4 , \u6/N3 , \u6/N2 , \u6/N1 , \u6/N0 , \u4/N6917 , \u4/N6916 ,
         \u4/N6915 , \u4/N6463 , \u4/N6462 , \u4/N6461 , \u4/N6460 ,
         \u4/N6459 , \u4/N6458 , \u4/N6457 , \u4/N6456 , \u4/N6455 ,
         \u4/N6454 , \u4/N6410 , \u4/N6286 , \u4/N6284 , \u4/N6283 ,
         \u4/N6280 , \u4/N6279 , \u4/N6278 , \u4/N6251 , \u4/N6249 ,
         \u4/N6203 , \u4/N6194 , \u4/N6172 , \u4/N6171 , \u4/div_exp2[0] ,
         \u4/div_exp2[1] , \u4/div_exp2[2] , \u4/div_exp2[3] ,
         \u4/div_exp2[4] , \u4/div_exp2[5] , \u4/div_exp2[6] ,
         \u4/div_exp2[7] , \u4/div_exp2[8] , \u4/div_exp2[9] ,
         \u4/div_exp2[10] , \u4/div_exp1[0] , \u4/div_exp1[1] ,
         \u4/div_exp1[2] , \u4/div_exp1[3] , \u4/div_exp1[4] ,
         \u4/div_exp1[5] , \u4/div_exp1[6] , \u4/div_exp1[7] ,
         \u4/div_exp1[8] , \u4/div_exp1[9] , \u4/div_exp1[10] ,
         \u4/fi_ldz_2a[0] , \u4/fi_ldz_2a[1] , \u4/fi_ldz_2a[2] ,
         \u4/fi_ldz_2a[3] , \u4/fi_ldz_2a[4] , \u4/fi_ldz_2a[5] ,
         \u4/fi_ldz_2a[6] , \u4/ldz_all[0] , \u4/ldz_all[1] , \u4/ldz_all[2] ,
         \u4/ldz_all[3] , \u4/ldz_all[4] , \u4/ldz_all[5] , \u4/ldz_all[6] ,
         \u4/N6142 , \u4/N6141 , \u4/N6140 , \u4/N6139 , \u4/N6138 ,
         \u4/N6137 , \u4/N6136 , \u4/exp_out1[0] , \u4/exp_out1[1] ,
         \u4/exp_out_pl1[0] , \u4/exp_out_pl1[1] , \u4/exp_out_pl1[2] ,
         \u4/exp_out_pl1[3] , \u4/exp_out_pl1[4] , \u4/exp_out_pl1[5] ,
         \u4/exp_out_pl1[6] , \u4/exp_out_pl1[7] , \u4/exp_out_pl1[8] ,
         \u4/exp_out_pl1[9] , \u4/exp_out_pl1[10] , \u4/fi_ldz_mi1[0] ,
         \u4/fi_ldz_mi1[1] , \u4/fi_ldz_mi1[2] , \u4/fi_ldz_mi1[3] ,
         \u4/fi_ldz_mi1[4] , \u4/fi_ldz_mi1[5] , \u4/fi_ldz_mi1[6] ,
         \u4/N6119 , \u4/N6118 , \u4/N6117 , \u4/N6116 , \u4/N6115 ,
         \u4/N6114 , \u4/N6113 , \u4/N6112 , \u4/N6111 , \u4/N6110 ,
         \u4/N6109 , \u4/N6108 , \u4/N6107 , \u4/N6106 , \u4/N6105 ,
         \u4/N6104 , \u4/N6103 , \u4/N6102 , \u4/N6101 , \u4/N6100 ,
         \u4/N6099 , \u4/N6098 , \u4/N6097 , \u4/N6096 , \u4/N6095 ,
         \u4/N6094 , \u4/N6093 , \u4/N6092 , \u4/N6091 , \u4/N6090 ,
         \u4/N6089 , \u4/N6088 , \u4/N6087 , \u4/N6086 , \u4/N6085 ,
         \u4/N6084 , \u4/N6083 , \u4/N6082 , \u4/N6081 , \u4/N6080 ,
         \u4/N6079 , \u4/N6078 , \u4/N6077 , \u4/N6076 , \u4/N6075 ,
         \u4/N6074 , \u4/N6073 , \u4/N6072 , \u4/N6071 , \u4/N6070 ,
         \u4/N6069 , \u4/N6068 , \u4/N6067 , \u4/N6066 , \u4/N6065 ,
         \u4/N6064 , \u4/N6063 , \u4/N6062 , \u4/N6061 , \u4/N6060 ,
         \u4/N6059 , \u4/N6058 , \u4/N6057 , \u4/N6056 , \u4/N6055 ,
         \u4/N6054 , \u4/N6053 , \u4/N6052 , \u4/N6051 , \u4/N6050 ,
         \u4/N6049 , \u4/N6048 , \u4/N6047 , \u4/N6046 , \u4/N6045 ,
         \u4/N6044 , \u4/N6043 , \u4/N6042 , \u4/N6041 , \u4/N6040 ,
         \u4/N6039 , \u4/N6038 , \u4/N6037 , \u4/N6036 , \u4/N6035 ,
         \u4/N6034 , \u4/N6033 , \u4/N6032 , \u4/N6031 , \u4/N6030 ,
         \u4/N6029 , \u4/N6028 , \u4/N6027 , \u4/N6026 , \u4/N6025 ,
         \u4/N6024 , \u4/N6023 , \u4/N6022 , \u4/N6021 , \u4/N6020 ,
         \u4/N6019 , \u4/N6018 , \u4/N6017 , \u4/N6016 , \u4/N6015 ,
         \u4/N6014 , \u4/N6011 , \u4/N6010 , \u4/N6009 , \u4/N6008 ,
         \u4/N6007 , \u4/N6006 , \u4/N6005 , \u4/N6004 , \u4/N6003 ,
         \u4/N6002 , \u4/N6001 , \u4/N6000 , \u4/N5999 , \u4/N5998 ,
         \u4/N5997 , \u4/N5996 , \u4/N5995 , \u4/N5994 , \u4/N5993 ,
         \u4/N5992 , \u4/N5991 , \u4/N5990 , \u4/N5989 , \u4/N5988 ,
         \u4/N5987 , \u4/N5986 , \u4/N5985 , \u4/N5984 , \u4/N5983 ,
         \u4/N5982 , \u4/N5981 , \u4/N5980 , \u4/N5979 , \u4/N5978 ,
         \u4/N5977 , \u4/N5976 , \u4/N5975 , \u4/N5974 , \u4/N5973 ,
         \u4/N5972 , \u4/N5971 , \u4/N5970 , \u4/N5969 , \u4/N5968 ,
         \u4/N5967 , \u4/N5966 , \u4/N5965 , \u4/N5964 , \u4/N5963 ,
         \u4/N5962 , \u4/N5961 , \u4/N5960 , \u4/N5959 , \u4/N5958 ,
         \u4/N5957 , \u4/N5956 , \u4/N5955 , \u4/N5954 , \u4/N5953 ,
         \u4/N5952 , \u4/N5951 , \u4/N5950 , \u4/N5949 , \u4/N5948 ,
         \u4/N5947 , \u4/N5946 , \u4/N5945 , \u4/N5944 , \u4/N5943 ,
         \u4/N5942 , \u4/N5941 , \u4/N5940 , \u4/N5939 , \u4/N5938 ,
         \u4/N5937 , \u4/N5936 , \u4/N5935 , \u4/N5934 , \u4/N5933 ,
         \u4/N5932 , \u4/N5931 , \u4/N5930 , \u4/N5929 , \u4/N5928 ,
         \u4/N5927 , \u4/N5926 , \u4/N5925 , \u4/N5924 , \u4/N5923 ,
         \u4/N5922 , \u4/N5921 , \u4/N5920 , \u4/N5919 , \u4/N5918 ,
         \u4/N5917 , \u4/N5916 , \u4/N5915 , \u4/N5914 , \u4/N5913 ,
         \u4/N5912 , \u4/N5911 , \u4/N5910 , \u4/N5909 , \u4/N5908 ,
         \u4/N5907 , \u4/N5906 , \u4/N5904 , \u4/exp_in_pl1[0] ,
         \u4/exp_in_pl1[1] , \u4/exp_in_pl1[2] , \u4/exp_in_pl1[3] ,
         \u4/exp_in_pl1[4] , \u4/exp_in_pl1[5] , \u4/exp_in_pl1[6] ,
         \u4/exp_in_pl1[7] , \u4/exp_in_pl1[8] , \u4/exp_in_pl1[9] ,
         \u4/exp_in_pl1[10] , \u4/exp_in_pl1[11] , \u4/f2i_shft[1] ,
         \u4/f2i_shft[2] , \u4/f2i_shft[3] , \u4/f2i_shft[4] ,
         \u4/f2i_shft[5] , \u4/f2i_shft[6] , \u4/f2i_shft[7] ,
         \u4/f2i_shft[8] , \u4/f2i_shft[9] , \u4/f2i_shft[10] , \u4/N5843 ,
         \u4/div_shft3[0] , \u4/div_shft3[1] , \u4/div_shft3[2] ,
         \u4/div_shft3[3] , \u4/div_shft3[4] , \u4/div_shft3[5] ,
         \u4/div_shft3[6] , \u4/div_shft3[7] , \u4/div_shft3[8] ,
         \u4/div_shft3[9] , \u4/div_shft3[10] , \u4/exp_in_mi1[1] ,
         \u4/exp_in_mi1[2] , \u4/exp_in_mi1[3] , \u4/exp_in_mi1[4] ,
         \u4/exp_in_mi1[5] , \u4/exp_in_mi1[6] , \u4/exp_in_mi1[7] ,
         \u4/exp_in_mi1[8] , \u4/exp_in_mi1[9] , \u4/exp_in_mi1[10] ,
         \u4/exp_in_mi1[11] , \u4/N5837 , \u4/N5836 , \u4/fract_out_pl1[0] ,
         \u4/fract_out_pl1[1] , \u4/fract_out_pl1[2] , \u4/fract_out_pl1[3] ,
         \u4/fract_out_pl1[4] , \u4/fract_out_pl1[5] , \u4/fract_out_pl1[6] ,
         \u4/fract_out_pl1[7] , \u4/fract_out_pl1[8] , \u4/fract_out_pl1[9] ,
         \u4/fract_out_pl1[10] , \u4/fract_out_pl1[11] ,
         \u4/fract_out_pl1[12] , \u4/fract_out_pl1[13] ,
         \u4/fract_out_pl1[14] , \u4/fract_out_pl1[15] ,
         \u4/fract_out_pl1[16] , \u4/fract_out_pl1[17] ,
         \u4/fract_out_pl1[18] , \u4/fract_out_pl1[19] ,
         \u4/fract_out_pl1[20] , \u4/fract_out_pl1[21] ,
         \u4/fract_out_pl1[22] , \u4/fract_out_pl1[23] ,
         \u4/fract_out_pl1[24] , \u4/fract_out_pl1[25] ,
         \u4/fract_out_pl1[26] , \u4/fract_out_pl1[27] ,
         \u4/fract_out_pl1[28] , \u4/fract_out_pl1[29] ,
         \u4/fract_out_pl1[30] , \u4/fract_out_pl1[31] ,
         \u4/fract_out_pl1[32] , \u4/fract_out_pl1[33] ,
         \u4/fract_out_pl1[34] , \u4/fract_out_pl1[35] ,
         \u4/fract_out_pl1[36] , \u4/fract_out_pl1[37] ,
         \u4/fract_out_pl1[38] , \u4/fract_out_pl1[39] ,
         \u4/fract_out_pl1[40] , \u4/fract_out_pl1[41] ,
         \u4/fract_out_pl1[42] , \u4/fract_out_pl1[43] ,
         \u4/fract_out_pl1[44] , \u4/fract_out_pl1[45] ,
         \u4/fract_out_pl1[46] , \u4/fract_out_pl1[47] ,
         \u4/fract_out_pl1[48] , \u4/fract_out_pl1[49] ,
         \u4/fract_out_pl1[50] , \u4/fract_out_pl1[51] ,
         \u4/fract_out_pl1[52] , \u4/exp_next_mi[0] , \u4/exp_next_mi[1] ,
         \u4/exp_next_mi[2] , \u4/exp_next_mi[3] , \u4/exp_next_mi[4] ,
         \u4/exp_next_mi[5] , \u4/exp_next_mi[6] , \u4/exp_next_mi[7] ,
         \u4/exp_next_mi[8] , \u4/exp_next_mi[9] , \u4/exp_next_mi[10] ,
         \u4/exp_next_mi[11] , \u4/fract_out[0] , \u4/fract_out[1] ,
         \u4/fract_out[2] , \u4/fract_out[3] , \u4/fract_out[4] ,
         \u4/fract_out[5] , \u4/fract_out[6] , \u4/fract_out[7] ,
         \u4/fract_out[8] , \u4/fract_out[9] , \u4/fract_out[10] ,
         \u4/fract_out[11] , \u4/fract_out[12] , \u4/fract_out[13] ,
         \u4/fract_out[14] , \u4/fract_out[15] , \u4/fract_out[16] ,
         \u4/fract_out[17] , \u4/fract_out[18] , \u4/fract_out[19] ,
         \u4/fract_out[20] , \u4/fract_out[21] , \u4/fract_out[22] ,
         \u4/fract_out[23] , \u4/fract_out[24] , \u4/fract_out[25] ,
         \u4/fract_out[26] , \u4/fract_out[27] , \u4/fract_out[28] ,
         \u4/fract_out[29] , \u4/fract_out[30] , \u4/fract_out[31] ,
         \u4/fract_out[32] , \u4/fract_out[33] , \u4/fract_out[34] ,
         \u4/fract_out[35] , \u4/fract_out[36] , \u4/fract_out[37] ,
         \u4/fract_out[38] , \u4/fract_out[39] , \u4/fract_out[40] ,
         \u4/fract_out[41] , \u4/fract_out[42] , \u4/fract_out[43] ,
         \u4/fract_out[44] , \u4/fract_out[45] , \u4/fract_out[46] ,
         \u4/fract_out[47] , \u4/fract_out[48] , \u4/fract_out[49] ,
         \u4/fract_out[50] , \u4/fract_out[51] , \u4/exp_out[0] ,
         \u4/exp_out[1] , \u4/exp_out[2] , \u4/exp_out[3] , \u4/exp_out[4] ,
         \u4/exp_out[5] , \u4/exp_out[6] , \u4/exp_out[7] , \u4/exp_out[8] ,
         \u4/exp_out[9] , \u4/exp_out[10] , \u4/fi_ldz[1] , \u4/fi_ldz[2] ,
         \u4/fi_ldz[3] , \u4/fi_ldz[4] , \u4/fi_ldz[5] , \u4/fi_ldz[6] , n203,
         n204, n205, n2388, n2389, n2390, n2391, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3621, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4194, n4195,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, \u4/ldz_dif[9] , \u4/ldz_dif[8] , \u4/ldz_dif[7] ,
         \u4/ldz_dif[6] , \u4/ldz_dif[5] , \u4/ldz_dif[4] , \u4/ldz_dif[3] ,
         \u4/ldz_dif[2] , \u4/ldz_dif[1] , \u4/ldz_dif[10] , \u4/ldz_dif[0] ,
         \u2/lt_135/A[0] , \u2/lt_135/A[5] , \u2/lt_135/A[6] ,
         \u2/lt_135/A[7] , \u2/lt_135/A[8] , \u2/lt_135/A[9] ,
         \u2/gt_145/B[11] , \u4/sub_463/carry[2] , \u4/sub_463/carry[3] ,
         \u4/sub_463/carry[4] , \u4/sub_463/carry[5] , \u4/sub_463/carry[6] ,
         \u4/sub_468/A[2] , \u4/sub_468/A[3] , \u4/sub_468/A[4] ,
         \u4/sub_468/A[5] , \u4/sub_468/A[7] , \u4/sub_468/A[9] ,
         \u4/sub_468/A[10] , \u4/sub_417/carry[2] , \u4/sub_417/carry[3] ,
         \u4/sub_417/carry[4] , \u4/sub_417/carry[5] , \u4/sub_417/carry[6] ,
         \u4/sub_417/carry[7] , \u4/sub_417/carry[8] , \u4/sub_417/carry[9] ,
         \u4/sub_417/carry[10] , \u2/sub_116/carry[2] , \u2/sub_116/carry[3] ,
         \u2/sub_116/carry[4] , \u2/sub_116/carry[5] , \u2/sub_116/carry[6] ,
         \u2/sub_116/carry[7] , \u2/sub_116/carry[8] , \u2/sub_116/carry[9] ,
         \u2/sub_116/carry[10] , \u2/sub_116/carry[11] , \u2/add_116/carry[2] ,
         \u2/add_116/carry[3] , \u2/add_116/carry[4] , \u2/add_116/carry[5] ,
         \u2/add_116/carry[6] , \u2/add_116/carry[7] , \u2/add_116/carry[8] ,
         \u2/add_116/carry[9] , \u2/add_116/carry[10] , \u2/add_116/carry[11] ,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468;
  wire   [63:52] opa_r;
  wire   [63:52] opb_r;
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  wire   [1:0] rmode_r1;
  wire   [1:0] rmode_r2;
  wire   [1:0] rmode_r3;
  wire   [2:0] fpu_op_r1;
  wire   [2:0] fpu_op_r2;
<<<<<<< HEAD
  wire   [13:0] fracta;
  wire   [13:0] fractb;
  wire   [9:0] fracta_mul;
  wire   [1:0] exp_ovf;
  wire   [2:0] underflow_fmul_d;
  wire   [14:1] fract_out_q;
  wire   [21:0] prod;
  wire   [22:0] quo;
  wire   [3:0] div_opa_ldz_r1;
  wire   [3:0] div_opa_ldz_r2;
  wire   [4:1] exp_r;
  wire   [11:4] opa_r1;
  wire   [10:9] fract_denorm;
  wire   [2:1] underflow_fmul_r;
  wire   [13:0] \u1/fractb_s ;
  wire   [13:0] \u1/fracta_s ;
  wire   [2:1] \u2/underflow_d ;
  wire   [21:0] \u5/prod1 ;
  wire   [23:0] \u6/remainder ;
  wire   [23:0] \u6/quo1 ;
  wire   [27:23] \u4/exp_f2i_1 ;
  wire   [2:0] \u4/shift_left ;
  wire   [4:0] \u4/shift_right ;
  wire   [4:3] \u4/add_407/carry ;
  wire   [4:2] \u2/add_115/carry ;
  wire   [4:2] \u2/add_113/carry ;
  wire   [4:1] \u2/add_110/carry ;
  wire   [5:1] \u2/sub_110/carry ;
  wire   [20:8] \sub_435_3/carry ;
  wire   [10:2] \sub_435_b0/carry ;
=======
  wire   [2:0] fpu_op_r3;
  wire   [55:0] fracta;
  wire   [55:0] fractb;
  wire   [10:0] exp_fasu;
  wire   [51:0] fracta_mul;
  wire   [7:2] exp_mul;
  wire   [1:0] exp_ovf;
  wire   [2:0] underflow_fmul_d;
  wire   [1:0] exp_ovf_r;
  wire   [56:0] fract_out_q;
  wire   [105:0] prod;
  wire   [4:0] div_opa_ldz_d;
  wire   [107:0] quo;
  wire   [107:0] remainder;
  wire   [4:0] div_opa_ldz_r1;
  wire   [4:0] div_opa_ldz_r2;
  wire   [6:1] exp_r;
  wire   [59:0] opa_r1;
  wire   [105:0] fract_i2f;
  wire   [105:50] fract_denorm;
  wire   [2:0] underflow_fmul_r;
  wire   [55:0] \u1/fractb_s ;
  wire   [55:0] \u1/fracta_s ;
  wire   [10:0] \u1/exp_diff2 ;
  wire   [10:0] \u1/exp_small ;
  wire   [2:0] \u2/underflow_d ;
  wire   [105:0] \u5/prod1 ;
  wire   [107:0] \u6/remainder ;
  wire   [107:0] \u6/quo1 ;
  wire   [10:0] \u4/div_exp3 ;
  wire   [117:107] \u4/exp_f2i_1 ;
  wire   [10:0] \u4/exp_fix_divb ;
  wire   [10:0] \u4/exp_fix_diva ;
  wire   [10:0] \u4/exp_out1_mi1 ;
  wire   [10:0] \u4/exp_out_mi1 ;
  wire   [6:1] \u4/fi_ldz_mi22 ;
  wire   [8:0] \u4/shift_left ;
  wire   [10:0] \u4/shift_right ;
  wire   [10:0] \u4/div_shft4 ;
  wire   [10:2] \u4/div_shft2 ;
  wire   [10:0] \u4/div_scht1a ;
  wire   [6:2] \u4/sub_481/carry ;
  wire   [10:1] \u4/sub_412/carry ;
  wire   [10:1] \u4/add_411/carry ;
  wire   [10:3] \u4/add_410/carry ;
  wire   [10:1] \u4/sub_409/carry ;
  wire   [6:2] \u4/sub_491/carry ;
  wire   [10:1] \sub_1_root_sub_0_root_u4/add_497/carry ;
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
<<<<<<< HEAD
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45;

  OR2_X2 \u4/C1739  ( .A1(\u4/N655 ), .A2(net30297), .ZN(\u4/N656 ) );
  OR2_X2 \u4/C1742  ( .A1(net85842), .A2(n2997), .ZN(\u4/N653 ) );
  OR2_X2 \u4/C1935  ( .A1(\u4/shift_right [4]), .A2(\u4/shift_right [3]), .ZN(
        \u4/N386 ) );
  AOI22_X2 U16 ( .A1(\u4/div_exp3[1] ), .A2(net15944), .B1(n3009), .B2(
        net77815), .ZN(n845) );
  OAI211_X2 U18 ( .C1(net89919), .C2(n3010), .A(n851), .B(n1669), .ZN(
        \u4/exp_out[2] ) );
  OAI221_X2 U100 ( .B1(net83296), .B2(n872), .C1(n888), .C2(net85794), .A(
        n1664), .ZN(\u4/shift_right [0]) );
  DFF_X2 \opa_r_reg[15]  ( .D(opa[15]), .CK(clk), .Q(opa_r[15]), .QN(n1569) );
  DFF_X2 \opa_r_reg[14]  ( .D(opa[14]), .CK(clk), .Q(opa_r[14]), .QN(n1594) );
  DFF_X2 \opa_r_reg[13]  ( .D(opa[13]), .CK(clk), .Q(opa_r[13]), .QN(n1560) );
  DFF_X2 \opa_r_reg[12]  ( .D(opa[12]), .CK(clk), .Q(opa_r[12]), .QN(n1573) );
  DFF_X2 \opa_r_reg[11]  ( .D(opa[11]), .CK(clk), .Q(opa_r[11]), .QN(n1725) );
  DFF_X2 \opa_r_reg[10]  ( .D(opa[10]), .CK(clk), .Q(opa_r[10]), .QN(n1723) );
  DFF_X2 \opa_r_reg[9]  ( .D(opa[9]), .CK(clk), .Q(fracta_mul[9]), .QN(n3120)
         );
  DFF_X2 \opa_r_reg[8]  ( .D(opa[8]), .CK(clk), .Q(fracta_mul[8]), .QN(n3119)
         );
  DFF_X2 \opa_r_reg[7]  ( .D(opa[7]), .CK(clk), .Q(fracta_mul[7]), .QN(n3118)
         );
  DFF_X2 \opa_r_reg[6]  ( .D(opa[6]), .CK(clk), .Q(fracta_mul[6]), .QN(n3117)
         );
  DFF_X2 \opa_r_reg[5]  ( .D(opa[5]), .CK(clk), .Q(fracta_mul[5]), .QN(n3116)
         );
  DFF_X2 \opa_r_reg[4]  ( .D(opa[4]), .CK(clk), .Q(fracta_mul[4]), .QN(n3115)
         );
  DFF_X2 \opa_r_reg[3]  ( .D(opa[3]), .CK(clk), .Q(fracta_mul[3]), .QN(n3114)
         );
  DFF_X2 \opa_r_reg[2]  ( .D(opa[2]), .CK(clk), .Q(fracta_mul[2]), .QN(n3113)
         );
  DFF_X2 \opa_r_reg[1]  ( .D(opa[1]), .CK(clk), .Q(fracta_mul[1]), .QN(n3112)
         );
  DFF_X2 \opa_r_reg[0]  ( .D(opa[0]), .CK(clk), .Q(fracta_mul[0]), .QN(n3111)
         );
  DFF_X2 \opb_r_reg[15]  ( .D(opb[15]), .CK(clk), .Q(opb_r[15]), .QN(n1686) );
  DFF_X2 \opb_r_reg[14]  ( .D(opb[14]), .CK(clk), .Q(opb_r[14]), .QN(n1734) );
  DFF_X2 \opb_r_reg[13]  ( .D(opb[13]), .CK(clk), .Q(opb_r[13]), .QN(n1728) );
  DFF_X2 \opb_r_reg[12]  ( .D(opb[12]), .CK(clk), .Q(opb_r[12]), .QN(n1727) );
  DFF_X2 \opb_r_reg[11]  ( .D(opb[11]), .CK(clk), .Q(opb_r[11]), .QN(n1730) );
  DFF_X2 \opb_r_reg[10]  ( .D(opb[10]), .CK(clk), .Q(opb_r[10]), .QN(n1726) );
  DFF_X2 \opb_r_reg[9]  ( .D(opb[9]), .CK(clk), .Q(\u6/N9 ), .QN(n3110) );
  DFF_X2 \opb_r_reg[8]  ( .D(opb[8]), .CK(clk), .Q(\u6/N8 ), .QN(n3109) );
  DFF_X2 \opb_r_reg[7]  ( .D(opb[7]), .CK(clk), .Q(\u6/N7 ), .QN(n3108) );
  DFF_X2 \opb_r_reg[6]  ( .D(opb[6]), .CK(clk), .Q(\u6/N6 ), .QN(n3107) );
  DFF_X2 \opb_r_reg[5]  ( .D(opb[5]), .CK(clk), .Q(\u6/N5 ), .QN(n3106) );
  DFF_X2 \opb_r_reg[4]  ( .D(opb[4]), .CK(clk), .Q(\u6/N4 ), .QN(n3105) );
  DFF_X2 \opb_r_reg[3]  ( .D(opb[3]), .CK(clk), .Q(\u6/N3 ), .QN(n3104) );
  DFF_X2 \opb_r_reg[2]  ( .D(opb[2]), .CK(clk), .Q(\u6/N2 ), .QN(n3103) );
  DFF_X2 \opb_r_reg[1]  ( .D(opb[1]), .CK(clk), .Q(\u6/N1 ), .QN(n3102) );
  DFF_X2 \opb_r_reg[0]  ( .D(opb[0]), .CK(clk), .Q(\u6/N0 ), .QN(n3101) );
=======
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157;

  OR2_X2 \u4/C19042  ( .A1(\u4/N6462 ), .A2(\u4/exp_out[0] ), .ZN(\u4/N6463 )
         );
  OR2_X2 \u4/C19043  ( .A1(\u4/N6461 ), .A2(\u4/exp_out[1] ), .ZN(\u4/N6462 )
         );
  OR2_X2 \u4/C19044  ( .A1(\u4/N6460 ), .A2(\u4/exp_out[2] ), .ZN(\u4/N6461 )
         );
  OR2_X2 \u4/C19045  ( .A1(\u4/N6459 ), .A2(\u4/exp_out[3] ), .ZN(\u4/N6460 )
         );
  OR2_X2 \u4/C19046  ( .A1(\u4/N6458 ), .A2(\u4/exp_out[4] ), .ZN(\u4/N6459 )
         );
  OR2_X2 \u4/C19047  ( .A1(\u4/N6457 ), .A2(\u4/exp_out[5] ), .ZN(\u4/N6458 )
         );
  OR2_X2 \u4/C19048  ( .A1(\u4/N6456 ), .A2(\u4/exp_out[6] ), .ZN(\u4/N6457 )
         );
  OR2_X2 \u4/C19049  ( .A1(\u4/N6455 ), .A2(\u4/exp_out[7] ), .ZN(\u4/N6456 )
         );
  OR2_X2 \u4/C19050  ( .A1(\u4/N6454 ), .A2(\u4/exp_out[8] ), .ZN(\u4/N6455 )
         );
  OR2_X2 \u4/C19051  ( .A1(\u4/exp_out[10] ), .A2(\u4/exp_out[9] ), .ZN(
        \u4/N6454 ) );
  OR2_X2 \u4/C19471  ( .A1(\u4/shift_right [10]), .A2(\u4/shift_right [9]), 
        .ZN(\u4/N5904 ) );
  OR2_X2 \u4/C19733  ( .A1(\u4/N6915 ), .A2(\u4/N6916 ), .ZN(\u4/N6917 ) );
  AND2_X2 \u4/C19735  ( .A1(\u4/exp_out[10] ), .A2(1'b1), .ZN(\u4/N6916 ) );
  MUX2_X2 U3 ( .A(prod[105]), .B(\fract_div[105] ), .S(fpu_op_r3[0]), .Z(n203)
         );
  MUX2_X2 U4 ( .A(fract_out_q[56]), .B(n203), .S(fpu_op_r3[1]), .Z(n204) );
  AND2_X2 U5 ( .A1(fract_i2f[105]), .A2(n4400), .ZN(n205) );
  MUX2_X2 U6 ( .A(n204), .B(n205), .S(n4661), .Z(fract_denorm[105]) );
  NAND2_X2 U8 ( .A1(n2388), .A2(n2389), .ZN(\u4/exp_out[0] ) );
  NAND2_X2 U11 ( .A1(\u4/div_exp3 [0]), .A2(n2394), .ZN(n2396) );
  AOI22_X2 U14 ( .A1(\u4/exp_f2i_1 [107]), .A2(n2400), .B1(n2401), .B2(
        \u4/exp_out1[0] ), .ZN(n2388) );
  OAI211_X2 U15 ( .C1(n5873), .C2(n4355), .A(n2402), .B(n2403), .ZN(
        \u4/exp_out[1] ) );
  AOI221_X2 U16 ( .B1(\u4/N6136 ), .B2(n2390), .C1(n2404), .C2(n6094), .A(
        n2405), .ZN(n2403) );
  NOR2_X4 U17 ( .A1(n4653), .A2(n2399), .ZN(n2404) );
  AOI22_X2 U18 ( .A1(\u4/exp_f2i_1 [108]), .A2(n2400), .B1(n2401), .B2(
        \u4/exp_out1[1] ), .ZN(n2402) );
  OAI221_X2 U19 ( .B1(n2407), .B2(n2408), .C1(n5872), .C2(n4355), .A(n2409), 
        .ZN(\u4/exp_out[2] ) );
  AOI221_X2 U20 ( .B1(\u4/exp_f2i_1 [109]), .B2(n2400), .C1(\u4/N6137 ), .C2(
        n2390), .A(n2405), .ZN(n2409) );
  OAI221_X2 U21 ( .B1(n2411), .B2(n2408), .C1(n5871), .C2(n4355), .A(n2412), 
        .ZN(\u4/exp_out[3] ) );
  AOI221_X2 U22 ( .B1(\u4/exp_f2i_1 [110]), .B2(n2400), .C1(\u4/N6138 ), .C2(
        n2390), .A(n2405), .ZN(n2412) );
  OAI221_X2 U23 ( .B1(n2414), .B2(n2408), .C1(n5870), .C2(n4355), .A(n2415), 
        .ZN(\u4/exp_out[4] ) );
  AOI221_X2 U24 ( .B1(\u4/exp_f2i_1 [111]), .B2(n2400), .C1(\u4/N6139 ), .C2(
        n2390), .A(n2405), .ZN(n2415) );
  OAI221_X2 U25 ( .B1(n2416), .B2(n2408), .C1(n5869), .C2(n4355), .A(n2417), 
        .ZN(\u4/exp_out[5] ) );
  AOI22_X2 U26 ( .A1(\u4/N6140 ), .A2(n2390), .B1(\u4/exp_f2i_1 [112]), .B2(
        n2400), .ZN(n2417) );
  OAI221_X2 U27 ( .B1(n2418), .B2(n2408), .C1(n5868), .C2(n4355), .A(n2419), 
        .ZN(\u4/exp_out[6] ) );
  AOI22_X2 U28 ( .A1(\u4/N6141 ), .A2(n2390), .B1(\u4/exp_f2i_1 [113]), .B2(
        n2400), .ZN(n2419) );
  OAI221_X2 U29 ( .B1(n2420), .B2(n2408), .C1(n5867), .C2(n4355), .A(n2421), 
        .ZN(\u4/exp_out[7] ) );
  AOI221_X2 U30 ( .B1(\u4/exp_f2i_1 [114]), .B2(n2400), .C1(\u4/N6142 ), .C2(
        n2390), .A(n2405), .ZN(n2421) );
  AND3_X2 U31 ( .A1(opas_r2), .A2(n6343), .A3(n2422), .ZN(n2405) );
  OAI221_X2 U32 ( .B1(n2424), .B2(n2408), .C1(n5866), .C2(n4355), .A(n2425), 
        .ZN(\u4/exp_out[8] ) );
  OAI221_X2 U34 ( .B1(n2428), .B2(n2408), .C1(n5865), .C2(n4355), .A(n2429), 
        .ZN(\u4/exp_out[9] ) );
  OAI221_X2 U36 ( .B1(n2431), .B2(n2408), .C1(n5864), .C2(n4355), .A(n2432), 
        .ZN(\u4/exp_out[10] ) );
  OAI211_X2 U101 ( .C1(n2442), .C2(n2443), .A(n2444), .B(n2445), .ZN(
        \u4/shift_right [9]) );
  AOI22_X2 U102 ( .A1(\u4/div_shft2 [9]), .A2(n2446), .B1(\u4/exp_in_mi1[9] ), 
        .B2(n2447), .ZN(n2445) );
  AOI22_X2 U103 ( .A1(\u4/div_shft4 [9]), .A2(n2448), .B1(\u4/div_shft3[9] ), 
        .B2(n2449), .ZN(n2444) );
  OAI211_X2 U104 ( .C1(n2442), .C2(n2450), .A(n2451), .B(n2452), .ZN(
        \u4/shift_right [8]) );
  AOI22_X2 U105 ( .A1(\u4/div_shft2 [8]), .A2(n2446), .B1(\u4/exp_in_mi1[8] ), 
        .B2(n2447), .ZN(n2452) );
  AOI22_X2 U106 ( .A1(\u4/div_shft4 [8]), .A2(n2448), .B1(\u4/div_shft3[8] ), 
        .B2(n2449), .ZN(n2451) );
  OAI211_X2 U107 ( .C1(n2442), .C2(n2453), .A(n2454), .B(n2455), .ZN(
        \u4/shift_right [7]) );
  AOI22_X2 U108 ( .A1(\u4/div_shft2 [7]), .A2(n2446), .B1(\u4/exp_in_mi1[7] ), 
        .B2(n2447), .ZN(n2455) );
  AOI22_X2 U109 ( .A1(\u4/div_shft4 [7]), .A2(n2448), .B1(\u4/div_shft3[7] ), 
        .B2(n2449), .ZN(n2454) );
  OAI211_X2 U110 ( .C1(n2442), .C2(n2456), .A(n2457), .B(n2458), .ZN(
        \u4/shift_right [6]) );
  AOI22_X2 U111 ( .A1(\u4/div_shft2 [6]), .A2(n2446), .B1(\u4/exp_in_mi1[6] ), 
        .B2(n2447), .ZN(n2458) );
  AOI22_X2 U112 ( .A1(\u4/div_shft4 [6]), .A2(n2448), .B1(\u4/div_shft3[6] ), 
        .B2(n2449), .ZN(n2457) );
  OAI211_X2 U113 ( .C1(n2442), .C2(n2459), .A(n2460), .B(n2461), .ZN(
        \u4/shift_right [5]) );
  AOI22_X2 U114 ( .A1(\u4/div_shft2 [5]), .A2(n2446), .B1(\u4/exp_in_mi1[5] ), 
        .B2(n2447), .ZN(n2461) );
  AOI22_X2 U115 ( .A1(\u4/div_shft4 [5]), .A2(n2448), .B1(\u4/div_shft3[5] ), 
        .B2(n2449), .ZN(n2460) );
  OAI211_X2 U116 ( .C1(n2442), .C2(n2462), .A(n2463), .B(n2464), .ZN(
        \u4/shift_right [4]) );
  AOI22_X2 U117 ( .A1(\u4/div_shft2 [4]), .A2(n2446), .B1(\u4/exp_in_mi1[4] ), 
        .B2(n2447), .ZN(n2464) );
  AOI22_X2 U118 ( .A1(\u4/div_shft4 [4]), .A2(n2448), .B1(\u4/div_shft3[4] ), 
        .B2(n2449), .ZN(n2463) );
  OAI211_X2 U119 ( .C1(n2442), .C2(n2465), .A(n2466), .B(n2467), .ZN(
        \u4/shift_right [3]) );
  AOI22_X2 U120 ( .A1(\u4/div_shft2 [3]), .A2(n2446), .B1(\u4/exp_in_mi1[3] ), 
        .B2(n2447), .ZN(n2467) );
  AOI22_X2 U121 ( .A1(\u4/div_shft4 [3]), .A2(n2448), .B1(\u4/div_shft3[3] ), 
        .B2(n2449), .ZN(n2466) );
  OAI211_X2 U122 ( .C1(n2442), .C2(n2468), .A(n2469), .B(n2470), .ZN(
        \u4/shift_right [2]) );
  AOI22_X2 U123 ( .A1(\u4/div_shft2 [2]), .A2(n2446), .B1(\u4/exp_in_mi1[2] ), 
        .B2(n2447), .ZN(n2470) );
  AOI22_X2 U124 ( .A1(\u4/div_shft4 [2]), .A2(n2448), .B1(\u4/div_shft3[2] ), 
        .B2(n2449), .ZN(n2469) );
  OAI211_X2 U125 ( .C1(n2442), .C2(n2471), .A(n2472), .B(n2473), .ZN(
        \u4/shift_right [1]) );
  AOI22_X2 U126 ( .A1(n4314), .A2(n2446), .B1(\u4/exp_in_mi1[1] ), .B2(n2447), 
        .ZN(n2473) );
  AOI22_X2 U127 ( .A1(\u4/div_shft4 [1]), .A2(n2448), .B1(\u4/div_shft3[1] ), 
        .B2(n2449), .ZN(n2472) );
  OAI211_X2 U128 ( .C1(\u4/N6915 ), .C2(n2442), .A(n2474), .B(n2475), .ZN(
        \u4/shift_right [10]) );
  AOI22_X2 U129 ( .A1(\u4/div_shft2 [10]), .A2(n2446), .B1(\u4/exp_in_mi1[10] ), .B2(n2447), .ZN(n2475) );
  AOI22_X2 U130 ( .A1(\u4/div_shft4 [10]), .A2(n2448), .B1(\u4/div_shft3[10] ), 
        .B2(n2449), .ZN(n2474) );
  OAI211_X2 U131 ( .C1(\u4/exp_out_mi1 [0]), .C2(n2442), .A(n2476), .B(n2477), 
        .ZN(\u4/shift_right [0]) );
  AOI22_X2 U132 ( .A1(n4600), .A2(n2446), .B1(n4349), .B2(n2447), .ZN(n2477)
         );
  AOI22_X2 U134 ( .A1(\u4/div_shft4 [0]), .A2(n2448), .B1(\u4/div_shft3[0] ), 
        .B2(n2449), .ZN(n2476) );
  NAND2_X2 U137 ( .A1(n2481), .A2(n2482), .ZN(\u4/shift_left [8]) );
  AOI22_X2 U138 ( .A1(\u4/f2i_shft[8] ), .A2(n6342), .B1(n4353), .B2(n2483), 
        .ZN(n2482) );
  AOI22_X2 U139 ( .A1(\u4/div_scht1a [8]), .A2(n2484), .B1(\u4/exp_in_pl1[8] ), 
        .B2(n2485), .ZN(n2481) );
  NAND2_X2 U140 ( .A1(n2486), .A2(n2487), .ZN(\u4/shift_left [7]) );
  AOI22_X2 U141 ( .A1(\u4/f2i_shft[7] ), .A2(n6342), .B1(n4281), .B2(n2483), 
        .ZN(n2487) );
  AOI22_X2 U142 ( .A1(\u4/div_scht1a [7]), .A2(n2484), .B1(\u4/exp_in_pl1[7] ), 
        .B2(n2485), .ZN(n2486) );
  INV_X4 U143 ( .A(n2488), .ZN(\u4/shift_left [6]) );
  AOI221_X2 U144 ( .B1(\u4/fi_ldz[6] ), .B2(n2489), .C1(n2485), .C2(
        \u4/exp_in_pl1[6] ), .A(n2490), .ZN(n2488) );
  INV_X4 U145 ( .A(n2491), .ZN(n2490) );
  INV_X4 U147 ( .A(n2492), .ZN(\u4/shift_left [5]) );
  AOI221_X2 U148 ( .B1(n2489), .B2(\u4/fi_ldz[5] ), .C1(n2485), .C2(
        \u4/exp_in_pl1[5] ), .A(n2493), .ZN(n2492) );
  INV_X4 U149 ( .A(n2494), .ZN(n2493) );
  OAI211_X2 U151 ( .C1(n2495), .C2(n6461), .A(n2496), .B(n2497), .ZN(
        \u4/shift_left [4]) );
  AOI22_X2 U153 ( .A1(\u4/div_scht1a [4]), .A2(n2484), .B1(\u4/fi_ldz[4] ), 
        .B2(n2489), .ZN(n2496) );
  OAI211_X2 U154 ( .C1(n2495), .C2(n6462), .A(n2499), .B(n2500), .ZN(
        \u4/shift_left [3]) );
  AOI22_X2 U156 ( .A1(\u4/div_scht1a [3]), .A2(n2484), .B1(\u4/fi_ldz[3] ), 
        .B2(n2489), .ZN(n2499) );
  OAI211_X2 U157 ( .C1(n2495), .C2(n6463), .A(n2501), .B(n2502), .ZN(
        \u4/shift_left [2]) );
  AOI22_X2 U159 ( .A1(\u4/div_scht1a [2]), .A2(n2484), .B1(\u4/fi_ldz[2] ), 
        .B2(n2489), .ZN(n2501) );
  NAND2_X2 U160 ( .A1(n2503), .A2(n2504), .ZN(\u4/shift_left [1]) );
  AOI221_X2 U161 ( .B1(\u4/f2i_shft[1] ), .B2(n6342), .C1(div_opa_ldz_r2[1]), 
        .C2(n2498), .A(n2505), .ZN(n2504) );
  INV_X4 U163 ( .A(n2511), .ZN(n2509) );
  OAI211_X2 U165 ( .C1(n2495), .C2(n4600), .A(n2512), .B(n2513), .ZN(
        \u4/shift_left [0]) );
  AOI22_X2 U168 ( .A1(\u4/div_scht1a [0]), .A2(n2484), .B1(\u4/fi_ldz_2a[0] ), 
        .B2(n2489), .ZN(n2512) );
  OAI211_X2 U169 ( .C1(n2508), .C2(n2511), .A(n2516), .B(n2517), .ZN(n2489) );
  INV_X4 U172 ( .A(n2485), .ZN(n2495) );
  INV_X4 U173 ( .A(n2519), .ZN(\u4/fract_out[5] ) );
  INV_X4 U174 ( .A(n2520), .ZN(\u4/fract_out[51] ) );
  INV_X4 U175 ( .A(n2521), .ZN(\u4/fract_out[50] ) );
  INV_X4 U176 ( .A(n2522), .ZN(\u4/fract_out[47] ) );
  INV_X4 U177 ( .A(n2523), .ZN(\u4/fract_out[46] ) );
  INV_X4 U178 ( .A(n2524), .ZN(\u4/fract_out[45] ) );
  INV_X4 U179 ( .A(n2525), .ZN(\u4/fract_out[40] ) );
  INV_X4 U180 ( .A(n2526), .ZN(\u4/fract_out[3] ) );
  INV_X4 U181 ( .A(n2527), .ZN(\u4/fract_out[39] ) );
  INV_X4 U182 ( .A(n2528), .ZN(\u4/fract_out[35] ) );
  INV_X4 U183 ( .A(n2529), .ZN(\u4/fract_out[34] ) );
  INV_X4 U184 ( .A(n2530), .ZN(\u4/fract_out[33] ) );
  INV_X4 U185 ( .A(n2531), .ZN(\u4/fract_out[29] ) );
  INV_X4 U186 ( .A(n2532), .ZN(\u4/fract_out[28] ) );
  INV_X4 U187 ( .A(n2533), .ZN(\u4/fract_out[27] ) );
  INV_X4 U188 ( .A(n2534), .ZN(\u4/fract_out[23] ) );
  INV_X4 U189 ( .A(n2535), .ZN(\u4/fract_out[22] ) );
  INV_X4 U190 ( .A(n2536), .ZN(\u4/fract_out[21] ) );
  INV_X4 U191 ( .A(n2537), .ZN(\u4/fract_out[17] ) );
  INV_X4 U192 ( .A(n2538), .ZN(\u4/fract_out[16] ) );
  INV_X4 U193 ( .A(n2539), .ZN(\u4/fract_out[15] ) );
  INV_X4 U194 ( .A(n2540), .ZN(\u4/fract_out[11] ) );
  INV_X4 U195 ( .A(n2541), .ZN(\u4/fract_out[10] ) );
  AND2_X2 U196 ( .A1(n2542), .A2(n6366), .ZN(\u4/fi_ldz[6] ) );
  NOR4_X2 U198 ( .A1(n2547), .A2(n2548), .A3(n2549), .A4(n2550), .ZN(n2546) );
  NOR4_X2 U199 ( .A1(n2551), .A2(n2552), .A3(n2553), .A4(n2554), .ZN(n2545) );
  NOR4_X2 U206 ( .A1(n2569), .A2(n2570), .A3(n2571), .A4(n6322), .ZN(n2568) );
  NAND4_X2 U208 ( .A1(n2574), .A2(n2575), .A3(n2576), .A4(n2577), .ZN(n2563)
         );
  NOR4_X2 U209 ( .A1(n2578), .A2(n2579), .A3(n2580), .A4(n2581), .ZN(n2577) );
  NOR4_X2 U210 ( .A1(n2582), .A2(n2583), .A3(n6333), .A4(n2584), .ZN(n2576) );
  NOR4_X2 U211 ( .A1(n2586), .A2(n2587), .A3(n2588), .A4(n2589), .ZN(n2575) );
  OAI211_X2 U215 ( .C1(n2593), .C2(n6328), .A(n2594), .B(n2595), .ZN(n2571) );
  OR3_X2 U221 ( .A1(n2604), .A2(n2605), .A3(n6332), .ZN(n2603) );
  NAND4_X2 U222 ( .A1(n2606), .A2(n2607), .A3(n2608), .A4(n2609), .ZN(n2569)
         );
  NOR4_X2 U223 ( .A1(n2610), .A2(n2611), .A3(n2612), .A4(n6330), .ZN(n2567) );
  NAND4_X2 U224 ( .A1(n2614), .A2(n2615), .A3(n2616), .A4(n2617), .ZN(n2610)
         );
  NOR4_X2 U225 ( .A1(n2618), .A2(n2619), .A3(n2620), .A4(n2621), .ZN(n2566) );
  NOR4_X2 U226 ( .A1(n2622), .A2(n2623), .A3(n2624), .A4(n2625), .ZN(n2565) );
  NOR4_X2 U228 ( .A1(n2583), .A2(n2611), .A3(n2630), .A4(n2631), .ZN(n2629) );
  AND3_X2 U231 ( .A1(fract_denorm[50]), .A2(n6403), .A3(n2637), .ZN(n2583) );
  AOI221_X2 U232 ( .B1(n2638), .B2(fract_denorm[98]), .C1(n2639), .C2(n6430), 
        .A(n2640), .ZN(n2628) );
  NAND4_X2 U241 ( .A1(n2655), .A2(n2656), .A3(n2657), .A4(n2658), .ZN(n2654)
         );
  NAND4_X2 U246 ( .A1(n2662), .A2(n6361), .A3(n6362), .A4(n4653), .ZN(n2656)
         );
  OR3_X2 U248 ( .A1(n2664), .A2(n2649), .A3(n2665), .ZN(n2653) );
  AND3_X2 U253 ( .A1(n2668), .A2(n6408), .A3(n2542), .ZN(n2586) );
  NAND4_X2 U256 ( .A1(n2672), .A2(n6323), .A3(n2673), .A4(n2674), .ZN(
        \u4/fi_ldz[1] ) );
  NOR4_X2 U257 ( .A1(n2675), .A2(n2676), .A3(n2677), .A4(n2678), .ZN(n2674) );
  OAI22_X2 U258 ( .A1(n6329), .A2(n2682), .B1(n2683), .B2(n2684), .ZN(n2675)
         );
  NAND2_X2 U259 ( .A1(n6423), .A2(n2685), .ZN(n2682) );
  OAI211_X2 U261 ( .C1(n6364), .C2(n2689), .A(n6361), .B(n6362), .ZN(n2686) );
  OR2_X2 U262 ( .A1(fract_denorm[101]), .A2(fract_denorm[102]), .ZN(n2689) );
  OR4_X2 U264 ( .A1(n2691), .A2(n2650), .A3(n6319), .A4(n2692), .ZN(n2665) );
  OR3_X2 U265 ( .A1(n2693), .A2(n2694), .A3(n2612), .ZN(n2692) );
  AND3_X2 U266 ( .A1(n2695), .A2(n6420), .A3(n2600), .ZN(n2612) );
  OR3_X2 U268 ( .A1(n2549), .A2(n2620), .A3(n2581), .ZN(n2693) );
  AND3_X2 U269 ( .A1(n2698), .A2(fract_denorm[52]), .A3(n2679), .ZN(n2581) );
  NAND4_X2 U273 ( .A1(n2602), .A2(n2702), .A3(n2703), .A4(n2704), .ZN(n2650)
         );
  AND3_X2 U275 ( .A1(n2705), .A2(fract_denorm[60]), .A3(n2562), .ZN(n2554) );
  AND3_X2 U277 ( .A1(n2706), .A2(n6406), .A3(n2542), .ZN(n2588) );
  NOR4_X2 U286 ( .A1(n6443), .A2(n2718), .A3(n2561), .A4(n6328), .ZN(n2717) );
  AOI221_X2 U289 ( .B1(n2647), .B2(fract_denorm[73]), .C1(n6336), .C2(
        fract_denorm[89]), .A(n2648), .ZN(n2713) );
  NAND4_X2 U290 ( .A1(n6321), .A2(n6320), .A3(n2719), .A4(n2720), .ZN(n2648)
         );
  AOI221_X2 U291 ( .B1(n2542), .B2(n6367), .C1(n2562), .C2(fract_denorm[65]), 
        .A(n2721), .ZN(n2720) );
  OAI221_X2 U292 ( .B1(n2593), .B2(n6328), .C1(n2722), .C2(n6332), .A(n2723), 
        .ZN(n2721) );
  AOI221_X2 U294 ( .B1(n6325), .B2(fract_denorm[81]), .C1(n6338), .C2(
        fract_denorm[97]), .A(n2701), .ZN(n2719) );
  NAND4_X2 U295 ( .A1(n2601), .A2(n2725), .A3(n2726), .A4(n2727), .ZN(n2701)
         );
  NOR4_X2 U297 ( .A1(n6334), .A2(n6388), .A3(n6387), .A4(fract_denorm[60]), 
        .ZN(n2557) );
  NAND4_X2 U298 ( .A1(n6325), .A2(n2728), .A3(fract_denorm[75]), .A4(n6381), 
        .ZN(n2617) );
  AND4_X2 U299 ( .A1(n2542), .A2(n2706), .A3(n6405), .A4(n2729), .ZN(n2589) );
  NAND4_X2 U300 ( .A1(n6338), .A2(n2707), .A3(fract_denorm[91]), .A4(n6354), 
        .ZN(n2726) );
  NAND4_X2 U301 ( .A1(n2639), .A2(n2708), .A3(n6426), .A4(n2730), .ZN(n2725)
         );
  NAND4_X2 U302 ( .A1(n2555), .A2(n2709), .A3(n6411), .A4(n2731), .ZN(n2601)
         );
  NAND4_X2 U303 ( .A1(n2606), .A2(n2732), .A3(n2733), .A4(n2734), .ZN(n2651)
         );
  AND4_X2 U305 ( .A1(n2562), .A2(n2735), .A3(fract_denorm[61]), .A4(n6389), 
        .ZN(n2553) );
  AND4_X2 U306 ( .A1(n6325), .A2(n2736), .A3(fract_denorm[77]), .A4(n6383), 
        .ZN(n2624) );
  AND4_X2 U307 ( .A1(n2542), .A2(n2668), .A3(n6407), .A4(n2737), .ZN(n2587) );
  NAND4_X2 U308 ( .A1(n6338), .A2(n2738), .A3(fract_denorm[93]), .A4(n6355), 
        .ZN(n2733) );
  NAND4_X2 U309 ( .A1(n2639), .A2(n2669), .A3(n6428), .A4(n2739), .ZN(n2732)
         );
  NAND4_X2 U310 ( .A1(n2555), .A2(n2670), .A3(n6414), .A4(n2740), .ZN(n2606)
         );
  NAND4_X2 U311 ( .A1(n2608), .A2(n2741), .A3(n2742), .A4(n2743), .ZN(n2688)
         );
  NOR4_X2 U313 ( .A1(n6334), .A2(n6392), .A3(fract_denorm[64]), .A4(
        fract_denorm[65]), .ZN(n2551) );
  NOR4_X2 U314 ( .A1(n2642), .A2(n6386), .A3(fract_denorm[80]), .A4(
        fract_denorm[81]), .ZN(n2622) );
  AND4_X2 U315 ( .A1(n2542), .A2(n6410), .A3(n2744), .A4(n2711), .ZN(n2584) );
  NAND4_X2 U316 ( .A1(n6338), .A2(fract_denorm[95]), .A3(n6356), .A4(n6358), 
        .ZN(n2742) );
  NAND4_X2 U317 ( .A1(n2639), .A2(n6432), .A3(n2681), .A4(n2722), .ZN(n2741)
         );
  NAND4_X2 U318 ( .A1(n2555), .A2(n6418), .A3(n2745), .A4(n2593), .ZN(n2608)
         );
  NAND4_X2 U321 ( .A1(n2614), .A2(n2746), .A3(n2747), .A4(n2748), .ZN(n2664)
         );
  NOR4_X2 U323 ( .A1(n6335), .A2(n6398), .A3(n6395), .A4(fract_denorm[70]), 
        .ZN(n2548) );
  AND4_X2 U324 ( .A1(n6336), .A2(n2749), .A3(fract_denorm[85]), .A4(n6376), 
        .ZN(n2619) );
  AND4_X2 U325 ( .A1(n2679), .A2(n2750), .A3(fract_denorm[53]), .A4(n6370), 
        .ZN(n2580) );
  NAND4_X2 U327 ( .A1(n6327), .A2(n2663), .A3(n6435), .A4(n2752), .ZN(n2746)
         );
  NAND4_X2 U328 ( .A1(n2600), .A2(n2660), .A3(n6421), .A4(n2753), .ZN(n2614)
         );
  NAND4_X2 U329 ( .A1(n2754), .A2(n2613), .A3(n2755), .A4(n2756), .ZN(n2691)
         );
  NOR4_X2 U330 ( .A1(n2621), .A2(n2550), .A3(n2582), .A4(n2757), .ZN(n2756) );
  NOR4_X2 U331 ( .A1(n6434), .A2(n2758), .A3(n2697), .A4(n2632), .ZN(n2757) );
  AND2_X2 U332 ( .A1(n2637), .A2(fract_denorm[51]), .ZN(n2582) );
  AND4_X2 U333 ( .A1(n2647), .A2(n2759), .A3(fract_denorm[67]), .A4(n6394), 
        .ZN(n2550) );
  AND4_X2 U334 ( .A1(n6336), .A2(n2760), .A3(fract_denorm[83]), .A4(n6374), 
        .ZN(n2621) );
  NAND4_X2 U336 ( .A1(n2600), .A2(n2695), .A3(n6419), .A4(n2762), .ZN(n2613)
         );
  NAND4_X2 U338 ( .A1(n2616), .A2(n2764), .A3(n2765), .A4(n2766), .ZN(n2690)
         );
  NOR4_X2 U340 ( .A1(n6335), .A2(n6399), .A3(fract_denorm[72]), .A4(
        fract_denorm[73]), .ZN(n2547) );
  AND4_X2 U341 ( .A1(n6336), .A2(fract_denorm[87]), .A3(n6377), .A4(n6379), 
        .ZN(n2618) );
  AND4_X2 U342 ( .A1(n2679), .A2(fract_denorm[55]), .A3(n6371), .A4(n6373), 
        .ZN(n2578) );
  OR3_X2 U343 ( .A1(n2767), .A2(n6351), .A3(n2684), .ZN(n2765) );
  NAND4_X2 U344 ( .A1(n6327), .A2(n6439), .A3(n2680), .A4(n2768), .ZN(n2764)
         );
  NAND4_X2 U345 ( .A1(n2600), .A2(n6425), .A3(n2769), .A4(n2685), .ZN(n2616)
         );
  AND3_X2 U350 ( .A1(n2698), .A2(n6400), .A3(n2679), .ZN(n2637) );
  AOI22_X2 U355 ( .A1(fract_denorm[105]), .A2(\u4/exp_in_pl1[9] ), .B1(n4654), 
        .B2(\u4/exp_next_mi[9] ), .ZN(n2428) );
  AOI22_X2 U356 ( .A1(fract_denorm[105]), .A2(\u4/exp_in_pl1[8] ), .B1(n4654), 
        .B2(\u4/exp_next_mi[8] ), .ZN(n2424) );
  AOI22_X2 U357 ( .A1(fract_denorm[105]), .A2(\u4/exp_in_pl1[7] ), .B1(n4654), 
        .B2(\u4/exp_next_mi[7] ), .ZN(n2420) );
  AOI22_X2 U358 ( .A1(fract_denorm[105]), .A2(\u4/exp_in_pl1[6] ), .B1(n4654), 
        .B2(\u4/exp_next_mi[6] ), .ZN(n2418) );
  AOI22_X2 U359 ( .A1(fract_denorm[105]), .A2(\u4/exp_in_pl1[5] ), .B1(n4654), 
        .B2(\u4/exp_next_mi[5] ), .ZN(n2416) );
  AOI22_X2 U360 ( .A1(fract_denorm[105]), .A2(\u4/exp_in_pl1[4] ), .B1(n4654), 
        .B2(\u4/exp_next_mi[4] ), .ZN(n2414) );
  AOI22_X2 U361 ( .A1(fract_denorm[105]), .A2(\u4/exp_in_pl1[3] ), .B1(n4654), 
        .B2(\u4/exp_next_mi[3] ), .ZN(n2411) );
  AOI22_X2 U362 ( .A1(fract_denorm[105]), .A2(\u4/exp_in_pl1[2] ), .B1(n4654), 
        .B2(\u4/exp_next_mi[2] ), .ZN(n2407) );
  OAI22_X2 U363 ( .A1(n4654), .A2(n6464), .B1(fract_denorm[105]), .B2(n6097), 
        .ZN(\u4/exp_out1[1] ) );
  AOI22_X2 U364 ( .A1(n4652), .A2(\u4/exp_in_pl1[10] ), .B1(n4654), .B2(
        \u4/exp_next_mi[10] ), .ZN(n2431) );
  OAI22_X2 U365 ( .A1(n4654), .A2(n4600), .B1(fract_denorm[105]), .B2(n6098), 
        .ZN(\u4/exp_out1[0] ) );
  INV_X4 U366 ( .A(\u4/exp_out[10] ), .ZN(\u4/N6915 ) );
  AOI22_X2 U368 ( .A1(n2773), .A2(n2774), .B1(n2775), .B2(n2776), .ZN(n2772)
         );
  NOR4_X2 U369 ( .A1(n2777), .A2(n6034), .A3(n6036), .A4(n6035), .ZN(n2776) );
  AND4_X2 U371 ( .A1(n2779), .A2(\u2/N27 ), .A3(\u2/N25 ), .A4(\u2/N26 ), .ZN(
        n2775) );
  AND3_X2 U372 ( .A1(\u2/N23 ), .A2(\u2/N22 ), .A3(\u2/N24 ), .ZN(n2779) );
  NOR4_X2 U373 ( .A1(n2780), .A2(n6024), .A3(\u2/N16 ), .A4(n4597), .ZN(n2774)
         );
  NOR4_X2 U375 ( .A1(n2781), .A2(n6026), .A3(n6030), .A4(n6028), .ZN(n2773) );
  OAI222_X2 U377 ( .A1(\u6/N52 ), .A2(n4268), .B1(n2782), .B2(n6274), .C1(
        n4602), .C2(n4267), .ZN(\u2/underflow_d [1]) );
  AOI22_X2 U378 ( .A1(n4603), .A2(n4267), .B1(n6303), .B2(n4268), .ZN(n2783)
         );
  AND3_X2 U379 ( .A1(n6275), .A2(n2784), .A3(\u2/N111 ), .ZN(
        \u2/underflow_d [0]) );
  AOI22_X2 U380 ( .A1(n4597), .A2(\u2/N27 ), .B1(n4598), .B2(\u2/N15 ), .ZN(
        n2795) );
  AOI22_X2 U381 ( .A1(n4597), .A2(\u2/N26 ), .B1(n4598), .B2(\u2/N14 ), .ZN(
        n2796) );
  AOI22_X2 U382 ( .A1(n4597), .A2(\u2/N25 ), .B1(n4598), .B2(\u2/N13 ), .ZN(
        n2797) );
  AOI22_X2 U383 ( .A1(n4597), .A2(\u2/N24 ), .B1(n4598), .B2(\u2/N12 ), .ZN(
        n2798) );
  AOI22_X2 U384 ( .A1(n4597), .A2(\u2/N23 ), .B1(n4598), .B2(\u2/N11 ), .ZN(
        n2799) );
  OAI22_X2 U385 ( .A1(n4599), .A2(n6033), .B1(n4597), .B2(n6024), .ZN(
        \u2/exp_tmp1[4] ) );
  OAI22_X2 U386 ( .A1(n4599), .A2(n6034), .B1(n4597), .B2(n6026), .ZN(
        \u2/exp_tmp1[3] ) );
  OAI22_X2 U387 ( .A1(n4599), .A2(n6035), .B1(n4597), .B2(n6028), .ZN(
        \u2/exp_tmp1[2] ) );
  OAI22_X2 U388 ( .A1(n4599), .A2(n6036), .B1(n4597), .B2(n6030), .ZN(
        \u2/exp_tmp1[1] ) );
  AOI22_X2 U390 ( .A1(n4597), .A2(\u2/N18 ), .B1(n4599), .B2(\u2/N6 ), .ZN(
        n2800) );
  OR3_X2 U392 ( .A1(n2803), .A2(n4599), .A3(n4363), .ZN(n2802) );
  NAND2_X2 U393 ( .A1(n4599), .A2(n4363), .ZN(n2801) );
  AOI22_X2 U394 ( .A1(\u2/N17 ), .A2(n4599), .B1(\u2/N29 ), .B2(n4597), .ZN(
        n2784) );
  OAI211_X2 U395 ( .C1(n2804), .C2(n2805), .A(n2806), .B(n2807), .ZN(\u2/N86 )
         );
  AOI22_X2 U396 ( .A1(\u2/exp_tmp3[10] ), .A2(n2808), .B1(\u2/exp_tmp4[10] ), 
        .B2(n2809), .ZN(n2807) );
  AOI22_X2 U397 ( .A1(\u2/N64 ), .A2(n2810), .B1(\u2/N75 ), .B2(n2811), .ZN(
        n2806) );
  OAI211_X2 U398 ( .C1(n2785), .C2(n2805), .A(n2812), .B(n2813), .ZN(\u2/N85 )
         );
  AOI22_X2 U399 ( .A1(\u2/exp_tmp3[9] ), .A2(n2808), .B1(n2795), .B2(n2809), 
        .ZN(n2813) );
  AOI22_X2 U400 ( .A1(\u2/N63 ), .A2(n2810), .B1(\u2/N74 ), .B2(n2811), .ZN(
        n2812) );
  AOI22_X2 U401 ( .A1(\u2/N39 ), .A2(n4599), .B1(\u2/N51 ), .B2(n4597), .ZN(
        n2785) );
  OAI211_X2 U402 ( .C1(n2786), .C2(n2805), .A(n2814), .B(n2815), .ZN(\u2/N84 )
         );
  AOI22_X2 U403 ( .A1(\u2/exp_tmp3[8] ), .A2(n2808), .B1(n2796), .B2(n2809), 
        .ZN(n2815) );
  AOI22_X2 U404 ( .A1(\u2/N62 ), .A2(n2810), .B1(\u2/N73 ), .B2(n2811), .ZN(
        n2814) );
  AOI22_X2 U405 ( .A1(\u2/N38 ), .A2(n4599), .B1(\u2/N50 ), .B2(n4597), .ZN(
        n2786) );
  OAI211_X2 U406 ( .C1(n2787), .C2(n2805), .A(n2816), .B(n2817), .ZN(\u2/N83 )
         );
  AOI22_X2 U407 ( .A1(\u2/exp_tmp3[7] ), .A2(n2808), .B1(n2797), .B2(n2809), 
        .ZN(n2817) );
  AOI22_X2 U408 ( .A1(\u2/N61 ), .A2(n2810), .B1(\u2/N72 ), .B2(n2811), .ZN(
        n2816) );
  AOI22_X2 U409 ( .A1(\u2/N37 ), .A2(n4599), .B1(\u2/N49 ), .B2(n4597), .ZN(
        n2787) );
  OAI211_X2 U410 ( .C1(n2788), .C2(n2805), .A(n2818), .B(n2819), .ZN(\u2/N82 )
         );
  AOI22_X2 U411 ( .A1(\u2/exp_tmp3[6] ), .A2(n2808), .B1(n2798), .B2(n2809), 
        .ZN(n2819) );
  AOI22_X2 U412 ( .A1(\u2/N60 ), .A2(n2810), .B1(\u2/N71 ), .B2(n2811), .ZN(
        n2818) );
  AOI22_X2 U413 ( .A1(\u2/N36 ), .A2(n4599), .B1(\u2/N48 ), .B2(n4597), .ZN(
        n2788) );
  OAI211_X2 U414 ( .C1(n2789), .C2(n2805), .A(n2820), .B(n2821), .ZN(\u2/N81 )
         );
  AOI22_X2 U415 ( .A1(\u2/exp_tmp3[5] ), .A2(n2808), .B1(n2799), .B2(n2809), 
        .ZN(n2821) );
  AOI22_X2 U416 ( .A1(\u2/N59 ), .A2(n2810), .B1(\u2/N70 ), .B2(n2811), .ZN(
        n2820) );
  AOI22_X2 U417 ( .A1(\u2/N35 ), .A2(n4599), .B1(\u2/N47 ), .B2(n4597), .ZN(
        n2789) );
  OAI211_X2 U418 ( .C1(n2790), .C2(n2805), .A(n2822), .B(n2823), .ZN(\u2/N80 )
         );
  AOI22_X2 U419 ( .A1(\u2/exp_tmp3[4] ), .A2(n2808), .B1(\u2/exp_tmp4[4] ), 
        .B2(n2809), .ZN(n2823) );
  AOI22_X2 U420 ( .A1(\u2/N58 ), .A2(n2810), .B1(\u2/N69 ), .B2(n2811), .ZN(
        n2822) );
  AOI22_X2 U421 ( .A1(\u2/N34 ), .A2(n4599), .B1(\u2/N46 ), .B2(n4597), .ZN(
        n2790) );
  OAI211_X2 U422 ( .C1(n2791), .C2(n2805), .A(n2824), .B(n2825), .ZN(\u2/N79 )
         );
  AOI22_X2 U423 ( .A1(\u2/exp_tmp3[3] ), .A2(n2808), .B1(\u2/exp_tmp4[3] ), 
        .B2(n2809), .ZN(n2825) );
  AOI22_X2 U424 ( .A1(\u2/N57 ), .A2(n2810), .B1(\u2/N68 ), .B2(n2811), .ZN(
        n2824) );
  AOI22_X2 U425 ( .A1(\u2/N33 ), .A2(n4599), .B1(\u2/N45 ), .B2(n4597), .ZN(
        n2791) );
  OAI211_X2 U426 ( .C1(n2792), .C2(n2805), .A(n2826), .B(n2827), .ZN(\u2/N78 )
         );
  AOI22_X2 U427 ( .A1(\u2/exp_tmp3[2] ), .A2(n2808), .B1(\u2/exp_tmp4[2] ), 
        .B2(n2809), .ZN(n2827) );
  AOI22_X2 U428 ( .A1(\u2/N56 ), .A2(n2810), .B1(\u2/N67 ), .B2(n2811), .ZN(
        n2826) );
  AOI22_X2 U429 ( .A1(\u2/N32 ), .A2(n4599), .B1(\u2/N44 ), .B2(n4597), .ZN(
        n2792) );
  OAI211_X2 U430 ( .C1(n2793), .C2(n2805), .A(n2828), .B(n2829), .ZN(\u2/N77 )
         );
  AOI22_X2 U431 ( .A1(\u2/exp_tmp3[1] ), .A2(n2808), .B1(\u2/exp_tmp4[1] ), 
        .B2(n2809), .ZN(n2829) );
  AOI22_X2 U432 ( .A1(\u2/N55 ), .A2(n2810), .B1(\u2/N66 ), .B2(n2811), .ZN(
        n2828) );
  AOI22_X2 U433 ( .A1(\u2/N31 ), .A2(n4599), .B1(\u2/N43 ), .B2(n4597), .ZN(
        n2793) );
  OAI211_X2 U434 ( .C1(n2794), .C2(n2805), .A(n2830), .B(n2831), .ZN(\u2/N76 )
         );
  AOI22_X2 U435 ( .A1(\u2/exp_tmp3[0] ), .A2(n2808), .B1(n2800), .B2(n2809), 
        .ZN(n2831) );
  AOI22_X2 U438 ( .A1(\u2/N54 ), .A2(n2810), .B1(\u2/lt_135/A[0] ), .B2(n2811), 
        .ZN(n2830) );
  NAND2_X2 U442 ( .A1(n2803), .A2(n2832), .ZN(\u2/exp_ovf_d[1] ) );
  AOI22_X2 U445 ( .A1(\u2/N40 ), .A2(n4599), .B1(\u2/N52 ), .B2(n4597), .ZN(
        n2804) );
  AOI22_X2 U446 ( .A1(\u2/N41 ), .A2(n4599), .B1(\u2/N53 ), .B2(n4597), .ZN(
        n2803) );
  AOI22_X2 U447 ( .A1(n2800), .A2(n4599), .B1(n2800), .B2(n4597), .ZN(n2794)
         );
  AND2_X2 U448 ( .A1(opb_r[63]), .A2(opa_r[63]), .ZN(\u2/N121 ) );
  NAND2_X2 U450 ( .A1(\u2/N113 ), .A2(n4597), .ZN(n2834) );
  NAND2_X2 U451 ( .A1(n6303), .A2(n4458), .ZN(n2833) );
  OAI22_X2 U453 ( .A1(n4636), .A2(n4533), .B1(n2835), .B2(n4643), .ZN(
        \u1/sign_d ) );
  XOR2_X2 U454 ( .A(opb_r[63]), .B(n4481), .Z(n2835) );
  OAI22_X2 U455 ( .A1(n4636), .A2(n2836), .B1(n2837), .B2(n4643), .ZN(
        \u1/fractb_s [9]) );
  OAI22_X2 U456 ( .A1(n4636), .A2(n2838), .B1(n2839), .B2(n4643), .ZN(
        \u1/fractb_s [8]) );
  OAI22_X2 U457 ( .A1(n4636), .A2(n2840), .B1(n2841), .B2(n4643), .ZN(
        \u1/fractb_s [7]) );
  OAI22_X2 U458 ( .A1(n4636), .A2(n2842), .B1(n2843), .B2(n4643), .ZN(
        \u1/fractb_s [6]) );
  OAI22_X2 U459 ( .A1(n4636), .A2(n2844), .B1(n2845), .B2(n4643), .ZN(
        \u1/fractb_s [5]) );
  OAI22_X2 U460 ( .A1(n4636), .A2(n2846), .B1(n2847), .B2(n4643), .ZN(
        \u1/fractb_s [55]) );
  OAI22_X2 U461 ( .A1(n4636), .A2(n2848), .B1(n2849), .B2(n4643), .ZN(
        \u1/fractb_s [54]) );
  OAI22_X2 U462 ( .A1(n4636), .A2(n2850), .B1(n2851), .B2(n4643), .ZN(
        \u1/fractb_s [53]) );
  OAI22_X2 U463 ( .A1(n4636), .A2(n2852), .B1(n2853), .B2(n4643), .ZN(
        \u1/fractb_s [52]) );
  OAI22_X2 U464 ( .A1(n4636), .A2(n2854), .B1(n2855), .B2(n4643), .ZN(
        \u1/fractb_s [51]) );
  OAI22_X2 U465 ( .A1(n4637), .A2(n2856), .B1(n2857), .B2(n4643), .ZN(
        \u1/fractb_s [50]) );
  OAI22_X2 U466 ( .A1(n4637), .A2(n2858), .B1(n2859), .B2(n4643), .ZN(
        \u1/fractb_s [4]) );
  OAI22_X2 U467 ( .A1(n4637), .A2(n2860), .B1(n2861), .B2(n4643), .ZN(
        \u1/fractb_s [49]) );
  OAI22_X2 U468 ( .A1(n4637), .A2(n2862), .B1(n2863), .B2(n4643), .ZN(
        \u1/fractb_s [48]) );
  OAI22_X2 U469 ( .A1(n4637), .A2(n2864), .B1(n2865), .B2(n4643), .ZN(
        \u1/fractb_s [47]) );
  OAI22_X2 U470 ( .A1(n4637), .A2(n2866), .B1(n2867), .B2(n4643), .ZN(
        \u1/fractb_s [46]) );
  OAI22_X2 U471 ( .A1(n4637), .A2(n2868), .B1(n2869), .B2(n4643), .ZN(
        \u1/fractb_s [45]) );
  OAI22_X2 U472 ( .A1(n4637), .A2(n2870), .B1(n2871), .B2(n4643), .ZN(
        \u1/fractb_s [44]) );
  OAI22_X2 U473 ( .A1(n4637), .A2(n2872), .B1(n2873), .B2(n4643), .ZN(
        \u1/fractb_s [43]) );
  OAI22_X2 U474 ( .A1(n4637), .A2(n2874), .B1(n2875), .B2(n4643), .ZN(
        \u1/fractb_s [42]) );
  OAI22_X2 U475 ( .A1(n4637), .A2(n2876), .B1(n2877), .B2(n4643), .ZN(
        \u1/fractb_s [41]) );
  OAI22_X2 U476 ( .A1(n4637), .A2(n2878), .B1(n2879), .B2(n4643), .ZN(
        \u1/fractb_s [40]) );
  OAI22_X2 U477 ( .A1(n4636), .A2(n2880), .B1(n2881), .B2(n4643), .ZN(
        \u1/fractb_s [3]) );
  OAI22_X2 U478 ( .A1(n4639), .A2(n2882), .B1(n2883), .B2(n4644), .ZN(
        \u1/fractb_s [39]) );
  OAI22_X2 U479 ( .A1(n4639), .A2(n2884), .B1(n2885), .B2(n4644), .ZN(
        \u1/fractb_s [38]) );
  OAI22_X2 U480 ( .A1(n4639), .A2(n2886), .B1(n2887), .B2(n4644), .ZN(
        \u1/fractb_s [37]) );
  OAI22_X2 U481 ( .A1(n4639), .A2(n2888), .B1(n2889), .B2(n4644), .ZN(
        \u1/fractb_s [36]) );
  OAI22_X2 U482 ( .A1(n4639), .A2(n2890), .B1(n2891), .B2(n4644), .ZN(
        \u1/fractb_s [35]) );
  OAI22_X2 U483 ( .A1(n4639), .A2(n2892), .B1(n2893), .B2(n4644), .ZN(
        \u1/fractb_s [34]) );
  OAI22_X2 U484 ( .A1(n4639), .A2(n2894), .B1(n2895), .B2(n4644), .ZN(
        \u1/fractb_s [33]) );
  OAI22_X2 U485 ( .A1(n4639), .A2(n2896), .B1(n2897), .B2(n4644), .ZN(
        \u1/fractb_s [32]) );
  OAI22_X2 U486 ( .A1(n4639), .A2(n2898), .B1(n2899), .B2(n4644), .ZN(
        \u1/fractb_s [31]) );
  OAI22_X2 U487 ( .A1(n4638), .A2(n2900), .B1(n2901), .B2(n4644), .ZN(
        \u1/fractb_s [30]) );
  OAI22_X2 U488 ( .A1(n4638), .A2(n2902), .B1(n4651), .B2(n2903), .ZN(
        \u1/fractb_s [2]) );
  OAI22_X2 U489 ( .A1(n4638), .A2(n2904), .B1(n2905), .B2(n4644), .ZN(
        \u1/fractb_s [29]) );
  OAI22_X2 U490 ( .A1(n4638), .A2(n2906), .B1(n2907), .B2(n4644), .ZN(
        \u1/fractb_s [28]) );
  OAI22_X2 U491 ( .A1(n4638), .A2(n2908), .B1(n2909), .B2(n4644), .ZN(
        \u1/fractb_s [27]) );
  OAI22_X2 U492 ( .A1(n4638), .A2(n2910), .B1(n2911), .B2(n4644), .ZN(
        \u1/fractb_s [26]) );
  OAI22_X2 U493 ( .A1(n4638), .A2(n2912), .B1(n2913), .B2(n4644), .ZN(
        \u1/fractb_s [25]) );
  OAI22_X2 U494 ( .A1(n4638), .A2(n2914), .B1(n2915), .B2(n4644), .ZN(
        \u1/fractb_s [24]) );
  OAI22_X2 U495 ( .A1(n4638), .A2(n2916), .B1(n2917), .B2(n4644), .ZN(
        \u1/fractb_s [23]) );
  OAI22_X2 U496 ( .A1(n4638), .A2(n2918), .B1(n2919), .B2(n4644), .ZN(
        \u1/fractb_s [22]) );
  OAI22_X2 U497 ( .A1(n4638), .A2(n2920), .B1(n2921), .B2(n4644), .ZN(
        \u1/fractb_s [21]) );
  OAI22_X2 U498 ( .A1(n4639), .A2(n2922), .B1(n2923), .B2(n4644), .ZN(
        \u1/fractb_s [20]) );
  OAI22_X2 U499 ( .A1(n4639), .A2(n2924), .B1(n4651), .B2(n2925), .ZN(
        \u1/fractb_s [1]) );
  OAI22_X2 U500 ( .A1(n4639), .A2(n2926), .B1(n2927), .B2(n4645), .ZN(
        \u1/fractb_s [19]) );
  OAI22_X2 U501 ( .A1(n4639), .A2(n2928), .B1(n2929), .B2(n4645), .ZN(
        \u1/fractb_s [18]) );
  OAI22_X2 U502 ( .A1(n4639), .A2(n2930), .B1(n2931), .B2(n4645), .ZN(
        \u1/fractb_s [17]) );
  OAI22_X2 U503 ( .A1(n4639), .A2(n2932), .B1(n2933), .B2(n4645), .ZN(
        \u1/fractb_s [16]) );
  OAI22_X2 U504 ( .A1(n4639), .A2(n2934), .B1(n2935), .B2(n4645), .ZN(
        \u1/fractb_s [15]) );
  OAI22_X2 U505 ( .A1(n4639), .A2(n2936), .B1(n2937), .B2(n4645), .ZN(
        \u1/fractb_s [14]) );
  OAI22_X2 U506 ( .A1(n4639), .A2(n2938), .B1(n2939), .B2(n4645), .ZN(
        \u1/fractb_s [13]) );
  OAI22_X2 U507 ( .A1(n4639), .A2(n2940), .B1(n2941), .B2(n4645), .ZN(
        \u1/fractb_s [12]) );
  OAI22_X2 U508 ( .A1(n4639), .A2(n2942), .B1(n2943), .B2(n4645), .ZN(
        \u1/fractb_s [11]) );
  OAI22_X2 U509 ( .A1(n4640), .A2(n2944), .B1(n2945), .B2(n4645), .ZN(
        \u1/fractb_s [10]) );
  OAI22_X2 U510 ( .A1(n4640), .A2(n2946), .B1(n4651), .B2(n2947), .ZN(
        \u1/fractb_s [0]) );
  OAI22_X2 U511 ( .A1(n2836), .A2(n4645), .B1(n4640), .B2(n2837), .ZN(
        \u1/fracta_s [9]) );
  AOI22_X2 U512 ( .A1(n4607), .A2(\u1/adj_op_out_sft[9] ), .B1(n4623), .B2(
        \u6/N6 ), .ZN(n2836) );
  OAI22_X2 U513 ( .A1(n2838), .A2(n4645), .B1(n4640), .B2(n2839), .ZN(
        \u1/fracta_s [8]) );
  AOI22_X2 U514 ( .A1(n4606), .A2(\u1/adj_op_out_sft[8] ), .B1(n4621), .B2(
        \u6/N5 ), .ZN(n2838) );
  OAI22_X2 U515 ( .A1(n2840), .A2(n4645), .B1(n4640), .B2(n2841), .ZN(
        \u1/fracta_s [7]) );
  AOI22_X2 U516 ( .A1(n4628), .A2(\u1/adj_op_out_sft[7] ), .B1(n4621), .B2(
        \u6/N4 ), .ZN(n2840) );
  OAI22_X2 U517 ( .A1(n2842), .A2(n4645), .B1(n4640), .B2(n2843), .ZN(
        \u1/fracta_s [6]) );
  AOI22_X2 U518 ( .A1(n4615), .A2(\u1/adj_op_out_sft[6] ), .B1(n4621), .B2(
        \u6/N3 ), .ZN(n2842) );
  OAI22_X2 U519 ( .A1(n2844), .A2(n4645), .B1(n4640), .B2(n2845), .ZN(
        \u1/fracta_s [5]) );
  AOI22_X2 U520 ( .A1(n4628), .A2(\u1/adj_op_out_sft[5] ), .B1(n4621), .B2(
        \u6/N2 ), .ZN(n2844) );
  OAI22_X2 U521 ( .A1(n2846), .A2(n4645), .B1(n4640), .B2(n2847), .ZN(
        \u1/fracta_s [55]) );
  AOI22_X2 U522 ( .A1(n4606), .A2(\u1/adj_op_out_sft[55] ), .B1(n4621), .B2(
        \u6/N52 ), .ZN(n2846) );
  OAI22_X2 U523 ( .A1(n2848), .A2(n4645), .B1(n4640), .B2(n2849), .ZN(
        \u1/fracta_s [54]) );
  AOI22_X2 U524 ( .A1(n4606), .A2(\u1/adj_op_out_sft[54] ), .B1(n4621), .B2(
        \u6/N51 ), .ZN(n2848) );
  OAI22_X2 U525 ( .A1(n2850), .A2(n4645), .B1(n4640), .B2(n2851), .ZN(
        \u1/fracta_s [53]) );
  AOI22_X2 U526 ( .A1(n4606), .A2(\u1/adj_op_out_sft[53] ), .B1(n4621), .B2(
        \u6/N50 ), .ZN(n2850) );
  OAI22_X2 U527 ( .A1(n2852), .A2(n4646), .B1(n4640), .B2(n2853), .ZN(
        \u1/fracta_s [52]) );
  AOI22_X2 U528 ( .A1(n4606), .A2(\u1/adj_op_out_sft[52] ), .B1(n4621), .B2(
        \u6/N49 ), .ZN(n2852) );
  OAI22_X2 U529 ( .A1(n2854), .A2(n4646), .B1(n4641), .B2(n2855), .ZN(
        \u1/fracta_s [51]) );
  AOI22_X2 U530 ( .A1(n4606), .A2(\u1/adj_op_out_sft[51] ), .B1(n4621), .B2(
        \u6/N48 ), .ZN(n2854) );
  OAI22_X2 U531 ( .A1(n2856), .A2(n4646), .B1(n4641), .B2(n2857), .ZN(
        \u1/fracta_s [50]) );
  AOI22_X2 U532 ( .A1(n4606), .A2(\u1/adj_op_out_sft[50] ), .B1(n4621), .B2(
        \u6/N47 ), .ZN(n2856) );
  OAI22_X2 U533 ( .A1(n2858), .A2(n4646), .B1(n4638), .B2(n2859), .ZN(
        \u1/fracta_s [4]) );
  AOI22_X2 U534 ( .A1(n4628), .A2(\u1/adj_op_out_sft[4] ), .B1(n4621), .B2(
        \u6/N1 ), .ZN(n2858) );
  OAI22_X2 U535 ( .A1(n2860), .A2(n4646), .B1(n4640), .B2(n2861), .ZN(
        \u1/fracta_s [49]) );
  AOI22_X2 U536 ( .A1(n4615), .A2(\u1/adj_op_out_sft[49] ), .B1(n4621), .B2(
        \u6/N46 ), .ZN(n2860) );
  OAI22_X2 U537 ( .A1(n2862), .A2(n4646), .B1(n4641), .B2(n2863), .ZN(
        \u1/fracta_s [48]) );
  AOI22_X2 U538 ( .A1(n4615), .A2(\u1/adj_op_out_sft[48] ), .B1(n4621), .B2(
        \u6/N45 ), .ZN(n2862) );
  OAI22_X2 U539 ( .A1(n2864), .A2(n4646), .B1(n4640), .B2(n2865), .ZN(
        \u1/fracta_s [47]) );
  AOI22_X2 U540 ( .A1(n4615), .A2(\u1/adj_op_out_sft[47] ), .B1(n4621), .B2(
        \u6/N44 ), .ZN(n2864) );
  OAI22_X2 U541 ( .A1(n2866), .A2(n4646), .B1(n4640), .B2(n2867), .ZN(
        \u1/fracta_s [46]) );
  AOI22_X2 U542 ( .A1(n4615), .A2(\u1/adj_op_out_sft[46] ), .B1(n4621), .B2(
        \u6/N43 ), .ZN(n2866) );
  OAI22_X2 U543 ( .A1(n2868), .A2(n4646), .B1(n4641), .B2(n2869), .ZN(
        \u1/fracta_s [45]) );
  AOI22_X2 U544 ( .A1(n4615), .A2(\u1/adj_op_out_sft[45] ), .B1(n4621), .B2(
        \u6/N42 ), .ZN(n2868) );
  OAI22_X2 U545 ( .A1(n2870), .A2(n4646), .B1(n4641), .B2(n2871), .ZN(
        \u1/fracta_s [44]) );
  AOI22_X2 U546 ( .A1(n4615), .A2(\u1/adj_op_out_sft[44] ), .B1(n4621), .B2(
        \u6/N41 ), .ZN(n2870) );
  OAI22_X2 U547 ( .A1(n2872), .A2(n4646), .B1(n4640), .B2(n2873), .ZN(
        \u1/fracta_s [43]) );
  AOI22_X2 U548 ( .A1(n4615), .A2(\u1/adj_op_out_sft[43] ), .B1(n4621), .B2(
        \u6/N40 ), .ZN(n2872) );
  OAI22_X2 U549 ( .A1(n2874), .A2(n4646), .B1(n4640), .B2(n2875), .ZN(
        \u1/fracta_s [42]) );
  AOI22_X2 U550 ( .A1(n4615), .A2(\u1/adj_op_out_sft[42] ), .B1(n4621), .B2(
        \u6/N39 ), .ZN(n2874) );
  OAI22_X2 U551 ( .A1(n2876), .A2(n4646), .B1(n4641), .B2(n2877), .ZN(
        \u1/fracta_s [41]) );
  AOI22_X2 U552 ( .A1(n4615), .A2(\u1/adj_op_out_sft[41] ), .B1(n4619), .B2(
        \u6/N38 ), .ZN(n2876) );
  OAI22_X2 U553 ( .A1(n2878), .A2(n4646), .B1(n4641), .B2(n2879), .ZN(
        \u1/fracta_s [40]) );
  AOI22_X2 U554 ( .A1(n4615), .A2(\u1/adj_op_out_sft[40] ), .B1(n4619), .B2(
        \u6/N37 ), .ZN(n2878) );
  OAI22_X2 U555 ( .A1(n2880), .A2(n4646), .B1(n4641), .B2(n2881), .ZN(
        \u1/fracta_s [3]) );
  AOI22_X2 U556 ( .A1(n4628), .A2(\u1/adj_op_out_sft[3] ), .B1(n4621), .B2(
        \u6/N0 ), .ZN(n2880) );
  OAI22_X2 U557 ( .A1(n2882), .A2(n4646), .B1(n4641), .B2(n2883), .ZN(
        \u1/fracta_s [39]) );
  AOI22_X2 U558 ( .A1(n4628), .A2(\u1/adj_op_out_sft[39] ), .B1(n4619), .B2(
        \u6/N36 ), .ZN(n2882) );
  OAI22_X2 U559 ( .A1(n2884), .A2(n4646), .B1(n4641), .B2(n2885), .ZN(
        \u1/fracta_s [38]) );
  AOI22_X2 U560 ( .A1(n4606), .A2(\u1/adj_op_out_sft[38] ), .B1(n4619), .B2(
        \u6/N35 ), .ZN(n2884) );
  OAI22_X2 U561 ( .A1(n2886), .A2(n4646), .B1(n4641), .B2(n2887), .ZN(
        \u1/fracta_s [37]) );
  AOI22_X2 U562 ( .A1(n4606), .A2(\u1/adj_op_out_sft[37] ), .B1(n4619), .B2(
        \u6/N34 ), .ZN(n2886) );
  OAI22_X2 U563 ( .A1(n2888), .A2(n4646), .B1(n4641), .B2(n2889), .ZN(
        \u1/fracta_s [36]) );
  AOI22_X2 U564 ( .A1(n4628), .A2(\u1/adj_op_out_sft[36] ), .B1(n4619), .B2(
        \u6/N33 ), .ZN(n2888) );
  OAI22_X2 U565 ( .A1(n2890), .A2(n4646), .B1(n4641), .B2(n2891), .ZN(
        \u1/fracta_s [35]) );
  AOI22_X2 U566 ( .A1(n4615), .A2(\u1/adj_op_out_sft[35] ), .B1(n4619), .B2(
        \u6/N32 ), .ZN(n2890) );
  OAI22_X2 U567 ( .A1(n2892), .A2(n4647), .B1(n4641), .B2(n2893), .ZN(
        \u1/fracta_s [34]) );
  AOI22_X2 U568 ( .A1(n4606), .A2(\u1/adj_op_out_sft[34] ), .B1(n4619), .B2(
        \u6/N31 ), .ZN(n2892) );
  OAI22_X2 U569 ( .A1(n2894), .A2(n4647), .B1(n4641), .B2(n2895), .ZN(
        \u1/fracta_s [33]) );
  AOI22_X2 U570 ( .A1(n4628), .A2(\u1/adj_op_out_sft[33] ), .B1(n4621), .B2(
        \u6/N30 ), .ZN(n2894) );
  OAI22_X2 U571 ( .A1(n2896), .A2(n4647), .B1(n4641), .B2(n2897), .ZN(
        \u1/fracta_s [32]) );
  AOI22_X2 U572 ( .A1(n4606), .A2(\u1/adj_op_out_sft[32] ), .B1(n4619), .B2(
        \u6/N29 ), .ZN(n2896) );
  OAI22_X2 U573 ( .A1(n2898), .A2(n4647), .B1(n4642), .B2(n2899), .ZN(
        \u1/fracta_s [31]) );
  AOI22_X2 U574 ( .A1(n4606), .A2(\u1/adj_op_out_sft[31] ), .B1(n4619), .B2(
        \u6/N28 ), .ZN(n2898) );
  OAI22_X2 U575 ( .A1(n2900), .A2(n4647), .B1(n4642), .B2(n2901), .ZN(
        \u1/fracta_s [30]) );
  AOI22_X2 U576 ( .A1(n4628), .A2(\u1/adj_op_out_sft[30] ), .B1(n4619), .B2(
        \u6/N27 ), .ZN(n2900) );
  OAI22_X2 U577 ( .A1(n4643), .A2(n2902), .B1(n4649), .B2(n2903), .ZN(
        \u1/fracta_s [2]) );
  NAND2_X2 U578 ( .A1(\u1/adj_op_out_sft[2] ), .A2(n4610), .ZN(n2902) );
  OAI22_X2 U579 ( .A1(n2904), .A2(n4647), .B1(n4642), .B2(n2905), .ZN(
        \u1/fracta_s [29]) );
  AOI22_X2 U580 ( .A1(n4615), .A2(\u1/adj_op_out_sft[29] ), .B1(n4619), .B2(
        \u6/N26 ), .ZN(n2904) );
  OAI22_X2 U581 ( .A1(n2906), .A2(n4647), .B1(n4638), .B2(n2907), .ZN(
        \u1/fracta_s [28]) );
  AOI22_X2 U582 ( .A1(n4606), .A2(\u1/adj_op_out_sft[28] ), .B1(n4619), .B2(
        \u6/N25 ), .ZN(n2906) );
  OAI22_X2 U583 ( .A1(n2908), .A2(n4645), .B1(n4638), .B2(n2909), .ZN(
        \u1/fracta_s [27]) );
  AOI22_X2 U584 ( .A1(n4606), .A2(\u1/adj_op_out_sft[27] ), .B1(n4619), .B2(
        \u6/N24 ), .ZN(n2908) );
  OAI22_X2 U585 ( .A1(n2910), .A2(n4647), .B1(n4649), .B2(n2911), .ZN(
        \u1/fracta_s [26]) );
  AOI22_X2 U586 ( .A1(n4606), .A2(\u1/adj_op_out_sft[26] ), .B1(n4619), .B2(
        \u6/N23 ), .ZN(n2910) );
  OAI22_X2 U587 ( .A1(n2912), .A2(n4647), .B1(n4649), .B2(n2913), .ZN(
        \u1/fracta_s [25]) );
  AOI22_X2 U588 ( .A1(n4606), .A2(\u1/adj_op_out_sft[25] ), .B1(n4619), .B2(
        \u6/N22 ), .ZN(n2912) );
  OAI22_X2 U589 ( .A1(n2914), .A2(n4647), .B1(n4642), .B2(n2915), .ZN(
        \u1/fracta_s [24]) );
  AOI22_X2 U590 ( .A1(n4606), .A2(\u1/adj_op_out_sft[24] ), .B1(n4619), .B2(
        \u6/N21 ), .ZN(n2914) );
  OAI22_X2 U591 ( .A1(n2916), .A2(n4647), .B1(n4638), .B2(n2917), .ZN(
        \u1/fracta_s [23]) );
  AOI22_X2 U592 ( .A1(n4606), .A2(\u1/adj_op_out_sft[23] ), .B1(n4619), .B2(
        \u6/N20 ), .ZN(n2916) );
  OAI22_X2 U593 ( .A1(n2918), .A2(n4647), .B1(n4642), .B2(n2919), .ZN(
        \u1/fracta_s [22]) );
  AOI22_X2 U594 ( .A1(n4628), .A2(\u1/adj_op_out_sft[22] ), .B1(n4622), .B2(
        \u6/N19 ), .ZN(n2918) );
  OAI22_X2 U595 ( .A1(n2920), .A2(n4647), .B1(n4642), .B2(n2921), .ZN(
        \u1/fracta_s [21]) );
  AOI22_X2 U596 ( .A1(n4606), .A2(\u1/adj_op_out_sft[21] ), .B1(n4622), .B2(
        \u6/N18 ), .ZN(n2920) );
  OAI22_X2 U597 ( .A1(n2922), .A2(n4647), .B1(n4642), .B2(n2923), .ZN(
        \u1/fracta_s [20]) );
  AOI22_X2 U598 ( .A1(n4615), .A2(\u1/adj_op_out_sft[20] ), .B1(n4622), .B2(
        \u6/N17 ), .ZN(n2922) );
  OAI22_X2 U599 ( .A1(n4643), .A2(n2924), .B1(n4642), .B2(n2925), .ZN(
        \u1/fracta_s [1]) );
  NAND2_X2 U600 ( .A1(\u1/adj_op_out_sft[1] ), .A2(n4628), .ZN(n2924) );
  OAI22_X2 U601 ( .A1(n2926), .A2(n4647), .B1(n4642), .B2(n2927), .ZN(
        \u1/fracta_s [19]) );
  AOI22_X2 U602 ( .A1(n4606), .A2(\u1/adj_op_out_sft[19] ), .B1(n4622), .B2(
        \u6/N16 ), .ZN(n2926) );
  OAI22_X2 U603 ( .A1(n2928), .A2(n4647), .B1(n4642), .B2(n2929), .ZN(
        \u1/fracta_s [18]) );
  AOI22_X2 U604 ( .A1(n4628), .A2(\u1/adj_op_out_sft[18] ), .B1(n4622), .B2(
        \u6/N15 ), .ZN(n2928) );
  OAI22_X2 U605 ( .A1(n2930), .A2(n4647), .B1(n4642), .B2(n2931), .ZN(
        \u1/fracta_s [17]) );
  AOI22_X2 U606 ( .A1(n4606), .A2(\u1/adj_op_out_sft[17] ), .B1(n4622), .B2(
        \u6/N14 ), .ZN(n2930) );
  OAI22_X2 U607 ( .A1(n2932), .A2(n4647), .B1(n4642), .B2(n2933), .ZN(
        \u1/fracta_s [16]) );
  AOI22_X2 U608 ( .A1(n4606), .A2(\u1/adj_op_out_sft[16] ), .B1(n4622), .B2(
        \u6/N13 ), .ZN(n2932) );
  OAI22_X2 U609 ( .A1(n2934), .A2(n4647), .B1(n4642), .B2(n2935), .ZN(
        \u1/fracta_s [15]) );
  AOI22_X2 U610 ( .A1(n4606), .A2(\u1/adj_op_out_sft[15] ), .B1(n4622), .B2(
        \u6/N12 ), .ZN(n2934) );
  OAI22_X2 U611 ( .A1(n2936), .A2(n4647), .B1(n4642), .B2(n2937), .ZN(
        \u1/fracta_s [14]) );
  AOI22_X2 U612 ( .A1(n4606), .A2(\u1/adj_op_out_sft[14] ), .B1(n4622), .B2(
        \u6/N11 ), .ZN(n2936) );
  OAI22_X2 U613 ( .A1(n2938), .A2(n4651), .B1(n4642), .B2(n2939), .ZN(
        \u1/fracta_s [13]) );
  AOI22_X2 U614 ( .A1(n4606), .A2(\u1/adj_op_out_sft[13] ), .B1(n4621), .B2(
        \u6/N10 ), .ZN(n2938) );
  OAI22_X2 U615 ( .A1(n2940), .A2(n4651), .B1(n4642), .B2(n2941), .ZN(
        \u1/fracta_s [12]) );
  AOI22_X2 U616 ( .A1(n4606), .A2(\u1/adj_op_out_sft[12] ), .B1(n4622), .B2(
        \u6/N9 ), .ZN(n2940) );
  OAI22_X2 U617 ( .A1(n2942), .A2(n4651), .B1(n4649), .B2(n2943), .ZN(
        \u1/fracta_s [11]) );
  AOI22_X2 U618 ( .A1(n4606), .A2(\u1/adj_op_out_sft[11] ), .B1(n4622), .B2(
        \u6/N8 ), .ZN(n2942) );
  OAI22_X2 U619 ( .A1(n2944), .A2(n4645), .B1(n4649), .B2(n2945), .ZN(
        \u1/fracta_s [10]) );
  AOI22_X2 U620 ( .A1(n4606), .A2(\u1/adj_op_out_sft[10] ), .B1(n4622), .B2(
        \u6/N7 ), .ZN(n2944) );
  OAI22_X2 U621 ( .A1(n4643), .A2(n2946), .B1(n4649), .B2(n2947), .ZN(
        \u1/fracta_s [0]) );
  NAND2_X2 U622 ( .A1(n4611), .A2(n2948), .ZN(n2946) );
  AOI22_X2 U623 ( .A1(n4622), .A2(\u1/adj_op_out_sft[9] ), .B1(fracta_mul[6]), 
        .B2(n4612), .ZN(n2837) );
  AOI22_X2 U624 ( .A1(n4622), .A2(\u1/adj_op_out_sft[8] ), .B1(n4615), .B2(
        fracta_mul[5]), .ZN(n2839) );
  AOI22_X2 U625 ( .A1(n4622), .A2(\u1/adj_op_out_sft[7] ), .B1(n4628), .B2(
        fracta_mul[4]), .ZN(n2841) );
  AOI22_X2 U626 ( .A1(n4622), .A2(\u1/adj_op_out_sft[6] ), .B1(n4628), .B2(
        fracta_mul[3]), .ZN(n2843) );
  AOI22_X2 U627 ( .A1(n4622), .A2(\u1/adj_op_out_sft[5] ), .B1(n4615), .B2(
        fracta_mul[2]), .ZN(n2845) );
  AOI22_X2 U628 ( .A1(n4621), .A2(\u1/adj_op_out_sft[55] ), .B1(n4602), .B2(
        n4612), .ZN(n2847) );
  AOI22_X2 U629 ( .A1(n4621), .A2(\u1/adj_op_out_sft[54] ), .B1(n4615), .B2(
        fracta_mul[51]), .ZN(n2849) );
  AOI22_X2 U630 ( .A1(n4621), .A2(\u1/adj_op_out_sft[53] ), .B1(n4606), .B2(
        fracta_mul[50]), .ZN(n2851) );
  AOI22_X2 U631 ( .A1(n4621), .A2(\u1/adj_op_out_sft[52] ), .B1(n4615), .B2(
        fracta_mul[49]), .ZN(n2853) );
  AOI22_X2 U632 ( .A1(n4621), .A2(\u1/adj_op_out_sft[51] ), .B1(n4615), .B2(
        fracta_mul[48]), .ZN(n2855) );
  AOI22_X2 U633 ( .A1(n4621), .A2(\u1/adj_op_out_sft[50] ), .B1(n4615), .B2(
        fracta_mul[47]), .ZN(n2857) );
  AOI22_X2 U634 ( .A1(n4621), .A2(\u1/adj_op_out_sft[4] ), .B1(n4628), .B2(
        fracta_mul[1]), .ZN(n2859) );
  AOI22_X2 U635 ( .A1(n4621), .A2(\u1/adj_op_out_sft[49] ), .B1(n4606), .B2(
        fracta_mul[46]), .ZN(n2861) );
  AOI22_X2 U636 ( .A1(n4621), .A2(\u1/adj_op_out_sft[48] ), .B1(n4615), .B2(
        fracta_mul[45]), .ZN(n2863) );
  AOI22_X2 U637 ( .A1(n4621), .A2(\u1/adj_op_out_sft[47] ), .B1(n4615), .B2(
        fracta_mul[44]), .ZN(n2865) );
  AOI22_X2 U638 ( .A1(n4621), .A2(\u1/adj_op_out_sft[46] ), .B1(n4615), .B2(
        fracta_mul[43]), .ZN(n2867) );
  AOI22_X2 U639 ( .A1(n4621), .A2(\u1/adj_op_out_sft[45] ), .B1(n4615), .B2(
        fracta_mul[42]), .ZN(n2869) );
  AOI22_X2 U640 ( .A1(n4621), .A2(\u1/adj_op_out_sft[44] ), .B1(n4615), .B2(
        fracta_mul[41]), .ZN(n2871) );
  AOI22_X2 U641 ( .A1(n4621), .A2(\u1/adj_op_out_sft[43] ), .B1(n4615), .B2(
        fracta_mul[40]), .ZN(n2873) );
  AOI22_X2 U642 ( .A1(n4621), .A2(\u1/adj_op_out_sft[42] ), .B1(n4615), .B2(
        fracta_mul[39]), .ZN(n2875) );
  AOI22_X2 U643 ( .A1(n4621), .A2(\u1/adj_op_out_sft[41] ), .B1(n4615), .B2(
        fracta_mul[38]), .ZN(n2877) );
  AOI22_X2 U644 ( .A1(n4621), .A2(\u1/adj_op_out_sft[40] ), .B1(n4615), .B2(
        fracta_mul[37]), .ZN(n2879) );
  AOI22_X2 U645 ( .A1(n4621), .A2(\u1/adj_op_out_sft[3] ), .B1(n4615), .B2(
        fracta_mul[0]), .ZN(n2881) );
  AOI22_X2 U646 ( .A1(n4619), .A2(\u1/adj_op_out_sft[39] ), .B1(n4606), .B2(
        fracta_mul[36]), .ZN(n2883) );
  AOI22_X2 U647 ( .A1(n4622), .A2(\u1/adj_op_out_sft[38] ), .B1(n4606), .B2(
        fracta_mul[35]), .ZN(n2885) );
  AOI22_X2 U648 ( .A1(n4621), .A2(\u1/adj_op_out_sft[37] ), .B1(n4606), .B2(
        fracta_mul[34]), .ZN(n2887) );
  AOI22_X2 U649 ( .A1(n4621), .A2(\u1/adj_op_out_sft[36] ), .B1(n4606), .B2(
        fracta_mul[33]), .ZN(n2889) );
  AOI22_X2 U650 ( .A1(n4621), .A2(\u1/adj_op_out_sft[35] ), .B1(n4606), .B2(
        fracta_mul[32]), .ZN(n2891) );
  AOI22_X2 U651 ( .A1(n4621), .A2(\u1/adj_op_out_sft[34] ), .B1(n4606), .B2(
        fracta_mul[31]), .ZN(n2893) );
  AOI22_X2 U652 ( .A1(n4621), .A2(\u1/adj_op_out_sft[33] ), .B1(n4606), .B2(
        fracta_mul[30]), .ZN(n2895) );
  AOI22_X2 U653 ( .A1(n4621), .A2(\u1/adj_op_out_sft[32] ), .B1(n4606), .B2(
        fracta_mul[29]), .ZN(n2897) );
  AOI22_X2 U654 ( .A1(n4621), .A2(\u1/adj_op_out_sft[31] ), .B1(n4611), .B2(
        fracta_mul[28]), .ZN(n2899) );
  AOI22_X2 U655 ( .A1(n4619), .A2(\u1/adj_op_out_sft[30] ), .B1(n4606), .B2(
        fracta_mul[27]), .ZN(n2901) );
  NAND2_X2 U656 ( .A1(\u1/adj_op_out_sft[2] ), .A2(n4626), .ZN(n2903) );
  AOI22_X2 U657 ( .A1(n4619), .A2(\u1/adj_op_out_sft[29] ), .B1(n4606), .B2(
        fracta_mul[26]), .ZN(n2905) );
  AOI22_X2 U658 ( .A1(n4619), .A2(\u1/adj_op_out_sft[28] ), .B1(n4611), .B2(
        fracta_mul[25]), .ZN(n2907) );
  AOI22_X2 U659 ( .A1(n4619), .A2(\u1/adj_op_out_sft[27] ), .B1(n4628), .B2(
        fracta_mul[24]), .ZN(n2909) );
  AOI22_X2 U660 ( .A1(n4619), .A2(\u1/adj_op_out_sft[26] ), .B1(n4611), .B2(
        fracta_mul[23]), .ZN(n2911) );
  AOI22_X2 U661 ( .A1(n4619), .A2(\u1/adj_op_out_sft[25] ), .B1(n4611), .B2(
        fracta_mul[22]), .ZN(n2913) );
  AOI22_X2 U662 ( .A1(n4619), .A2(\u1/adj_op_out_sft[24] ), .B1(n4611), .B2(
        fracta_mul[21]), .ZN(n2915) );
  AOI22_X2 U663 ( .A1(n4619), .A2(\u1/adj_op_out_sft[23] ), .B1(n4611), .B2(
        fracta_mul[20]), .ZN(n2917) );
  AOI22_X2 U664 ( .A1(n4619), .A2(\u1/adj_op_out_sft[22] ), .B1(n4611), .B2(
        fracta_mul[19]), .ZN(n2919) );
  AOI22_X2 U665 ( .A1(n4619), .A2(\u1/adj_op_out_sft[21] ), .B1(n4611), .B2(
        fracta_mul[18]), .ZN(n2921) );
  AOI22_X2 U666 ( .A1(n4619), .A2(\u1/adj_op_out_sft[20] ), .B1(n4611), .B2(
        fracta_mul[17]), .ZN(n2923) );
  NAND2_X2 U667 ( .A1(\u1/adj_op_out_sft[1] ), .A2(n4626), .ZN(n2925) );
  AOI22_X2 U668 ( .A1(n4619), .A2(\u1/adj_op_out_sft[19] ), .B1(n4615), .B2(
        fracta_mul[16]), .ZN(n2927) );
  AOI22_X2 U669 ( .A1(n4619), .A2(\u1/adj_op_out_sft[18] ), .B1(n4610), .B2(
        fracta_mul[15]), .ZN(n2929) );
  AOI22_X2 U670 ( .A1(n4619), .A2(\u1/adj_op_out_sft[17] ), .B1(n4610), .B2(
        fracta_mul[14]), .ZN(n2931) );
  AOI22_X2 U671 ( .A1(n4619), .A2(\u1/adj_op_out_sft[16] ), .B1(n4610), .B2(
        fracta_mul[13]), .ZN(n2933) );
  AOI22_X2 U672 ( .A1(n4621), .A2(\u1/adj_op_out_sft[15] ), .B1(n4610), .B2(
        fracta_mul[12]), .ZN(n2935) );
  AOI22_X2 U673 ( .A1(n4621), .A2(\u1/adj_op_out_sft[14] ), .B1(n4610), .B2(
        fracta_mul[11]), .ZN(n2937) );
  AOI22_X2 U674 ( .A1(n4621), .A2(\u1/adj_op_out_sft[13] ), .B1(n4610), .B2(
        fracta_mul[10]), .ZN(n2939) );
  AOI22_X2 U675 ( .A1(n4621), .A2(\u1/adj_op_out_sft[12] ), .B1(n4610), .B2(
        fracta_mul[9]), .ZN(n2941) );
  AOI22_X2 U676 ( .A1(n4621), .A2(\u1/adj_op_out_sft[11] ), .B1(n4610), .B2(
        fracta_mul[8]), .ZN(n2943) );
  AOI22_X2 U677 ( .A1(n4621), .A2(\u1/adj_op_out_sft[10] ), .B1(n4610), .B2(
        fracta_mul[7]), .ZN(n2945) );
  NAND2_X2 U678 ( .A1(n2948), .A2(n4626), .ZN(n2947) );
  OR3_X2 U679 ( .A1(\u1/adj_op_out_sft[0] ), .A2(n2949), .A3(n2950), .ZN(n2948) );
  AOI221_X2 U681 ( .B1(n6214), .B2(n2954), .C1(n6218), .C2(n2955), .A(n2956), 
        .ZN(n2952) );
  OAI22_X2 U682 ( .A1(n2957), .A2(n2958), .B1(n2959), .B2(n2960), .ZN(n2956)
         );
  AOI221_X2 U683 ( .B1(n6213), .B2(n2962), .C1(n6222), .C2(n2963), .A(n2964), 
        .ZN(n2951) );
  OAI22_X2 U684 ( .A1(n2965), .A2(n2966), .B1(n2967), .B2(n2968), .ZN(n2964)
         );
  OAI22_X2 U687 ( .A1(n2975), .A2(n2976), .B1(n2961), .B2(n2977), .ZN(n2974)
         );
  AOI22_X2 U688 ( .A1(n6216), .A2(n2978), .B1(n6220), .B2(n2979), .ZN(n2969)
         );
  OAI222_X2 U691 ( .A1(n2985), .A2(n2966), .B1(n2986), .B2(n2968), .C1(n2987), 
        .C2(n2980), .ZN(n2984) );
  OAI221_X2 U692 ( .B1(n2988), .B2(n2975), .C1(n2989), .C2(n2961), .A(n2990), 
        .ZN(n2983) );
  AOI22_X2 U693 ( .A1(n6216), .A2(n2991), .B1(n6220), .B2(n2992), .ZN(n2990)
         );
  OAI221_X2 U695 ( .B1(n2996), .B2(n2966), .C1(n2997), .C2(n2980), .A(n2998), 
        .ZN(n2994) );
  AOI22_X2 U696 ( .A1(n6220), .A2(n2999), .B1(n6212), .B2(n3000), .ZN(n2998)
         );
  NAND4_X2 U699 ( .A1(n6217), .A2(n6224), .A3(n6225), .A4(n3004), .ZN(n2980)
         );
  OAI221_X2 U701 ( .B1(n3005), .B2(n2961), .C1(n3006), .C2(n2960), .A(n3007), 
        .ZN(n2993) );
  AOI22_X2 U702 ( .A1(n3008), .A2(n3009), .B1(n6214), .B2(n3010), .ZN(n3007)
         );
  NAND2_X2 U703 ( .A1(n6217), .A2(n3011), .ZN(n2975) );
  NAND2_X2 U707 ( .A1(n2988), .A2(n3013), .ZN(n2954) );
  NAND2_X2 U709 ( .A1(n2977), .A2(n3014), .ZN(n3010) );
  NAND2_X2 U711 ( .A1(n2989), .A2(n3015), .ZN(n2955) );
  AND2_X2 U712 ( .A1(n3005), .A2(n3016), .ZN(n2989) );
  NAND2_X2 U715 ( .A1(n3011), .A2(n3003), .ZN(n2961) );
  NAND2_X2 U718 ( .A1(n2959), .A2(n3017), .ZN(n2978) );
  NAND2_X2 U720 ( .A1(n3006), .A2(n3018), .ZN(n2991) );
  NAND2_X2 U722 ( .A1(n2957), .A2(n3019), .ZN(n2979) );
  OR2_X2 U724 ( .A1(n2999), .A2(\u1/adj_op[37] ), .ZN(n2992) );
  OR2_X2 U725 ( .A1(n2972), .A2(\u1/adj_op[36] ), .ZN(n2999) );
  NAND2_X2 U726 ( .A1(n2967), .A2(n3020), .ZN(n2972) );
  AND2_X2 U727 ( .A1(n2986), .A2(n3021), .ZN(n2967) );
  OR2_X2 U729 ( .A1(n2973), .A2(\u1/adj_op[32] ), .ZN(n3000) );
  NAND2_X2 U730 ( .A1(n2965), .A2(n3022), .ZN(n2973) );
  AND2_X2 U731 ( .A1(n2985), .A2(n3023), .ZN(n2965) );
  AND2_X2 U732 ( .A1(n2996), .A2(n3024), .ZN(n2985) );
  OR2_X2 U734 ( .A1(n2962), .A2(\u1/adj_op[27] ), .ZN(n2971) );
  NAND2_X2 U735 ( .A1(n2987), .A2(n3025), .ZN(n2962) );
  AND2_X2 U736 ( .A1(n2997), .A2(n3026), .ZN(n2987) );
  AND4_X2 U737 ( .A1(n3027), .A2(n3028), .A3(n3029), .A4(n3030), .ZN(n2997) );
  NOR4_X2 U738 ( .A1(n3031), .A2(\u1/adj_op[3] ), .A3(n6233), .A4(n6235), .ZN(
        n3030) );
  NAND4_X2 U739 ( .A1(n3032), .A2(n3033), .A3(n3034), .A4(n3035), .ZN(n3031)
         );
  NOR4_X2 U740 ( .A1(n3036), .A2(\u1/adj_op[20] ), .A3(\u1/adj_op[22] ), .A4(
        \u1/adj_op[21] ), .ZN(n3029) );
  NOR4_X2 U742 ( .A1(n3040), .A2(\u1/adj_op[15] ), .A3(\u1/adj_op[17] ), .A4(
        \u1/adj_op[16] ), .ZN(n3028) );
  NOR4_X2 U744 ( .A1(n3044), .A2(\u1/adj_op[0] ), .A3(\u1/adj_op[11] ), .A4(
        \u1/adj_op[10] ), .ZN(n3027) );
  AOI22_X2 U746 ( .A1(n4606), .A2(opb_r[61]), .B1(n4623), .B2(opa_r[61]), .ZN(
        n3048) );
  AOI22_X2 U747 ( .A1(n4606), .A2(opb_r[60]), .B1(n4623), .B2(opa_r[60]), .ZN(
        n3049) );
  OAI22_X2 U748 ( .A1(n4625), .A2(n4340), .B1(n4614), .B2(n4442), .ZN(
        \u1/exp_small [7]) );
  OAI22_X2 U749 ( .A1(n4624), .A2(n4399), .B1(n4613), .B2(n4454), .ZN(
        \u1/exp_small [6]) );
  OAI22_X2 U750 ( .A1(n4625), .A2(n4296), .B1(n4613), .B2(n4453), .ZN(
        \u1/exp_small [5]) );
  OAI22_X2 U751 ( .A1(n4624), .A2(n4359), .B1(n4613), .B2(n4456), .ZN(
        \u1/exp_small [4]) );
  OAI22_X2 U752 ( .A1(n4625), .A2(n4321), .B1(n4614), .B2(n4358), .ZN(
        \u1/exp_small [3]) );
  OAI22_X2 U753 ( .A1(n4624), .A2(n4457), .B1(n4613), .B2(n4451), .ZN(
        \u1/exp_small [2]) );
  OAI22_X2 U754 ( .A1(n4625), .A2(n4275), .B1(n4614), .B2(n4450), .ZN(
        \u1/exp_small [1]) );
  OAI22_X2 U755 ( .A1(n4363), .A2(n4626), .B1(n4614), .B2(n4458), .ZN(
        \u1/exp_small [10]) );
  OAI22_X2 U756 ( .A1(n4625), .A2(n4270), .B1(n4614), .B2(n4449), .ZN(
        \u1/exp_small [0]) );
  NAND2_X2 U760 ( .A1(\u1/exp_diff[2] ), .A2(n6223), .ZN(n3003) );
  NAND2_X2 U761 ( .A1(\u1/exp_diff[1] ), .A2(n6223), .ZN(n2953) );
  NAND2_X2 U762 ( .A1(\u1/exp_diff[0] ), .A2(n6223), .ZN(n2995) );
  AND2_X2 U763 ( .A1(\u1/exp_diff2 [9]), .A2(n3052), .ZN(\u1/exp_diff[9] ) );
  AND2_X2 U764 ( .A1(\u1/exp_diff2 [8]), .A2(n3052), .ZN(\u1/exp_diff[8] ) );
  AND2_X2 U765 ( .A1(\u1/exp_diff2 [7]), .A2(n3052), .ZN(\u1/exp_diff[7] ) );
  AND2_X2 U766 ( .A1(\u1/exp_diff2 [6]), .A2(n3052), .ZN(\u1/exp_diff[6] ) );
  AND2_X2 U767 ( .A1(\u1/exp_diff2 [5]), .A2(n3052), .ZN(\u1/exp_diff[5] ) );
  AND2_X2 U768 ( .A1(\u1/exp_diff2 [4]), .A2(n3052), .ZN(\u1/exp_diff[4] ) );
  AND2_X2 U769 ( .A1(\u1/exp_diff2 [3]), .A2(n3052), .ZN(\u1/exp_diff[3] ) );
  AND2_X2 U770 ( .A1(\u1/exp_diff2 [2]), .A2(n3052), .ZN(\u1/exp_diff[2] ) );
  AND2_X2 U771 ( .A1(\u1/exp_diff2 [1]), .A2(n3052), .ZN(\u1/exp_diff[1] ) );
  AND2_X2 U772 ( .A1(\u1/exp_diff2 [10]), .A2(n3052), .ZN(\u1/exp_diff[10] )
         );
  AND2_X2 U773 ( .A1(\u1/exp_diff2 [0]), .A2(n3052), .ZN(\u1/exp_diff[0] ) );
  AOI22_X2 U775 ( .A1(n4606), .A2(\u6/N9 ), .B1(n4623), .B2(fracta_mul[9]), 
        .ZN(n3035) );
  AOI22_X2 U776 ( .A1(n4607), .A2(\u6/N8 ), .B1(n4623), .B2(fracta_mul[8]), 
        .ZN(n3034) );
  AOI22_X2 U777 ( .A1(n4607), .A2(\u6/N7 ), .B1(n4623), .B2(fracta_mul[7]), 
        .ZN(n3033) );
  AOI22_X2 U778 ( .A1(n4607), .A2(\u6/N6 ), .B1(n4623), .B2(fracta_mul[6]), 
        .ZN(n3032) );
  AOI22_X2 U779 ( .A1(n4607), .A2(\u6/N5 ), .B1(n4623), .B2(fracta_mul[5]), 
        .ZN(n3053) );
  OAI22_X2 U780 ( .A1(n4625), .A2(n4459), .B1(n4613), .B2(n4273), .ZN(
        \u1/adj_op[51] ) );
  AOI22_X2 U781 ( .A1(n4609), .A2(\u6/N50 ), .B1(n4623), .B2(fracta_mul[50]), 
        .ZN(n3013) );
  AOI22_X2 U782 ( .A1(n4609), .A2(\u6/N4 ), .B1(n4623), .B2(fracta_mul[4]), 
        .ZN(n3054) );
  AOI22_X2 U783 ( .A1(n4609), .A2(\u6/N49 ), .B1(n4623), .B2(fracta_mul[49]), 
        .ZN(n3055) );
  AOI22_X2 U784 ( .A1(n4609), .A2(\u6/N48 ), .B1(n4623), .B2(fracta_mul[48]), 
        .ZN(n3014) );
  AOI22_X2 U785 ( .A1(n4609), .A2(\u6/N47 ), .B1(n4624), .B2(fracta_mul[47]), 
        .ZN(n3056) );
  AOI22_X2 U786 ( .A1(n4609), .A2(\u6/N46 ), .B1(n4623), .B2(fracta_mul[46]), 
        .ZN(n3015) );
  AOI22_X2 U787 ( .A1(n4609), .A2(\u6/N45 ), .B1(n4624), .B2(fracta_mul[45]), 
        .ZN(n3016) );
  OAI22_X2 U788 ( .A1(n4625), .A2(n4468), .B1(n4613), .B2(n4277), .ZN(
        \u1/adj_op[44] ) );
  AOI22_X2 U789 ( .A1(n4609), .A2(\u6/N43 ), .B1(n4624), .B2(fracta_mul[43]), 
        .ZN(n3017) );
  OAI22_X2 U790 ( .A1(n4625), .A2(n4467), .B1(n4613), .B2(n4286), .ZN(
        \u1/adj_op[42] ) );
  AOI22_X2 U791 ( .A1(n4609), .A2(\u6/N41 ), .B1(n4623), .B2(fracta_mul[41]), 
        .ZN(n3018) );
  AOI22_X2 U792 ( .A1(n4609), .A2(\u6/N40 ), .B1(n4623), .B2(fracta_mul[40]), 
        .ZN(n3057) );
  OAI22_X2 U793 ( .A1(n4624), .A2(n4463), .B1(n4612), .B2(n4360), .ZN(
        \u1/adj_op[3] ) );
  AOI22_X2 U794 ( .A1(n4608), .A2(\u6/N39 ), .B1(n4623), .B2(fracta_mul[39]), 
        .ZN(n3019) );
  OAI22_X2 U795 ( .A1(n4625), .A2(n4465), .B1(n4612), .B2(n4284), .ZN(
        \u1/adj_op[38] ) );
  OAI22_X2 U796 ( .A1(n4625), .A2(n4471), .B1(n4613), .B2(n4272), .ZN(
        \u1/adj_op[37] ) );
  OAI22_X2 U797 ( .A1(n4625), .A2(n4470), .B1(n4613), .B2(n4276), .ZN(
        \u1/adj_op[36] ) );
  AOI22_X2 U798 ( .A1(n4608), .A2(\u6/N35 ), .B1(n4623), .B2(fracta_mul[35]), 
        .ZN(n3020) );
  AOI22_X2 U799 ( .A1(n4608), .A2(\u6/N34 ), .B1(n4624), .B2(fracta_mul[34]), 
        .ZN(n3021) );
  AOI22_X2 U800 ( .A1(n4608), .A2(\u6/N33 ), .B1(n4623), .B2(fracta_mul[33]), 
        .ZN(n3058) );
  OAI22_X2 U801 ( .A1(n4625), .A2(n4464), .B1(n4613), .B2(n4287), .ZN(
        \u1/adj_op[32] ) );
  AOI22_X2 U802 ( .A1(n4608), .A2(\u6/N31 ), .B1(n4623), .B2(fracta_mul[31]), 
        .ZN(n3022) );
  AOI22_X2 U803 ( .A1(n4608), .A2(\u6/N30 ), .B1(n4624), .B2(fracta_mul[30]), 
        .ZN(n3023) );
  AOI22_X2 U804 ( .A1(n4608), .A2(\u6/N2 ), .B1(n4623), .B2(fracta_mul[2]), 
        .ZN(n3038) );
  AOI22_X2 U805 ( .A1(n4608), .A2(\u6/N29 ), .B1(n4624), .B2(fracta_mul[29]), 
        .ZN(n3024) );
  OAI22_X2 U806 ( .A1(n4625), .A2(n4469), .B1(n4615), .B2(n4285), .ZN(
        \u1/adj_op[28] ) );
  OAI22_X2 U807 ( .A1(n4625), .A2(n4466), .B1(n4613), .B2(n4301), .ZN(
        \u1/adj_op[27] ) );
  AOI22_X2 U808 ( .A1(n4609), .A2(\u6/N26 ), .B1(n4624), .B2(fracta_mul[26]), 
        .ZN(n3025) );
  AOI22_X2 U809 ( .A1(n4608), .A2(\u6/N25 ), .B1(n4624), .B2(fracta_mul[25]), 
        .ZN(n3026) );
  AOI22_X2 U810 ( .A1(n4608), .A2(\u6/N24 ), .B1(n4624), .B2(fracta_mul[24]), 
        .ZN(n3037) );
  AOI22_X2 U811 ( .A1(n4608), .A2(\u6/N23 ), .B1(n4624), .B2(fracta_mul[23]), 
        .ZN(n3039) );
  OAI22_X2 U812 ( .A1(n4625), .A2(n4462), .B1(n4614), .B2(n4283), .ZN(
        \u1/adj_op[22] ) );
  OAI22_X2 U813 ( .A1(n4625), .A2(n4325), .B1(n4613), .B2(n4292), .ZN(
        \u1/adj_op[21] ) );
  OAI22_X2 U814 ( .A1(n4625), .A2(n4366), .B1(n4614), .B2(n4320), .ZN(
        \u1/adj_op[20] ) );
  AOI22_X2 U815 ( .A1(n4607), .A2(\u6/N1 ), .B1(n4624), .B2(fracta_mul[1]), 
        .ZN(n3042) );
  AOI22_X2 U816 ( .A1(n4607), .A2(\u6/N19 ), .B1(n4624), .B2(fracta_mul[19]), 
        .ZN(n3041) );
  AOI22_X2 U817 ( .A1(n4607), .A2(\u6/N18 ), .B1(n4624), .B2(fracta_mul[18]), 
        .ZN(n3043) );
  OAI22_X2 U818 ( .A1(n4625), .A2(n4461), .B1(n4614), .B2(n4319), .ZN(
        \u1/adj_op[17] ) );
  OAI22_X2 U819 ( .A1(n4625), .A2(n4324), .B1(n4614), .B2(n4362), .ZN(
        \u1/adj_op[16] ) );
  OAI22_X2 U820 ( .A1(n4625), .A2(n4365), .B1(n4615), .B2(n4318), .ZN(
        \u1/adj_op[15] ) );
  AOI22_X2 U821 ( .A1(n4607), .A2(\u6/N14 ), .B1(n4624), .B2(fracta_mul[14]), 
        .ZN(n3046) );
  AOI22_X2 U822 ( .A1(n4607), .A2(\u6/N13 ), .B1(n4624), .B2(fracta_mul[13]), 
        .ZN(n3045) );
  AOI22_X2 U823 ( .A1(n4607), .A2(\u6/N12 ), .B1(n4624), .B2(fracta_mul[12]), 
        .ZN(n3047) );
  OAI22_X2 U824 ( .A1(n4626), .A2(n4460), .B1(n4614), .B2(n4361), .ZN(
        \u1/adj_op[11] ) );
  OAI22_X2 U825 ( .A1(n4626), .A2(n4323), .B1(n4614), .B2(n4300), .ZN(
        \u1/adj_op[10] ) );
  OAI22_X2 U826 ( .A1(n4626), .A2(n4364), .B1(n4615), .B2(n4322), .ZN(
        \u1/adj_op[0] ) );
  OAI22_X2 U828 ( .A1(n4612), .A2(n4363), .B1(n4458), .B2(n4626), .ZN(
        \u1/exp_large[10] ) );
  AOI22_X2 U830 ( .A1(n4622), .A2(opb_r[61]), .B1(n4610), .B2(opa_r[61]), .ZN(
        n3050) );
  AOI22_X2 U832 ( .A1(n4622), .A2(opb_r[60]), .B1(n4610), .B2(opa_r[60]), .ZN(
        n3051) );
  OAI22_X2 U834 ( .A1(n4611), .A2(n4340), .B1(n4626), .B2(n4442), .ZN(
        \u1/exp_large[7] ) );
  OAI22_X2 U836 ( .A1(n4612), .A2(n4399), .B1(n4626), .B2(n4454), .ZN(
        \u1/exp_large[6] ) );
  OAI22_X2 U838 ( .A1(n4611), .A2(n4296), .B1(n4626), .B2(n4453), .ZN(
        \u1/exp_large[5] ) );
  OAI22_X2 U840 ( .A1(n4612), .A2(n4359), .B1(n4626), .B2(n4456), .ZN(
        \u1/exp_large[4] ) );
  OAI22_X2 U842 ( .A1(n4612), .A2(n4321), .B1(n4626), .B2(n4358), .ZN(
        \u1/exp_large[3] ) );
  OAI22_X2 U844 ( .A1(n4612), .A2(n4457), .B1(n4626), .B2(n4451), .ZN(
        \u1/exp_large[2] ) );
  OAI22_X2 U846 ( .A1(n4612), .A2(n4275), .B1(n4626), .B2(n4450), .ZN(
        \u1/exp_large[1] ) );
  OAI22_X2 U848 ( .A1(n4612), .A2(n4270), .B1(n4626), .B2(n4449), .ZN(
        \u1/exp_large[0] ) );
  NAND2_X2 U850 ( .A1(\u6/N52 ), .A2(n4602), .ZN(\u1/N46 ) );
  XOR2_X2 U851 ( .A(n4481), .B(\u2/sign_d ), .Z(\u1/N232 ) );
  XOR2_X2 U852 ( .A(opa_r[63]), .B(opb_r[63]), .Z(\u2/sign_d ) );
  AOI221_X2 U856 ( .B1(opb_nan), .B2(n3063), .C1(n3064), .C2(
        \u1/fracta_lt_fractb ), .A(\u1/signa_r ), .ZN(n3060) );
  NAND2_X2 U858 ( .A1(opa_nan), .A2(opb_nan), .ZN(n3063) );
  OAI22_X2 U859 ( .A1(n4490), .A2(n3065), .B1(n3066), .B2(n3067), .ZN(
        \u1/N218 ) );
  XOR2_X2 U860 ( .A(\u1/signb_r ), .B(\u1/add_r ), .Z(n3067) );
  AND2_X2 U861 ( .A1(n3065), .A2(n4490), .ZN(n3066) );
  AOI22_X2 U862 ( .A1(\u0/snan_r_a ), .A2(\u0/expa_ff ), .B1(\u0/snan_r_b ), 
        .B2(\u0/expb_ff ), .ZN(n3068) );
  AOI22_X2 U863 ( .A1(\u0/qnan_r_a ), .A2(\u0/expa_ff ), .B1(\u0/qnan_r_b ), 
        .B2(\u0/expb_ff ), .ZN(n3069) );
  NAND2_X2 U864 ( .A1(n3070), .A2(n3071), .ZN(\u0/N7 ) );
  AND2_X2 U866 ( .A1(n4459), .A2(n3072), .ZN(\u0/N5 ) );
  AND2_X2 U868 ( .A1(\u0/fractb_00 ), .A2(\u0/expb_00 ), .ZN(\u0/N17 ) );
  AND2_X2 U869 ( .A1(\u0/fracta_00 ), .A2(\u0/expa_00 ), .ZN(\u0/N16 ) );
  NAND2_X2 U870 ( .A1(\u0/infb_f_r ), .A2(\u0/expb_ff ), .ZN(n3070) );
  NAND2_X2 U871 ( .A1(\u0/infa_f_r ), .A2(\u0/expa_ff ), .ZN(n3071) );
  NAND4_X2 U874 ( .A1(opb_r[52]), .A2(opb_r[53]), .A3(n3076), .A4(n3077), .ZN(
        n3074) );
  NOR4_X2 U875 ( .A1(n3078), .A2(n4296), .A3(n4340), .A4(n4399), .ZN(n3077) );
  NAND4_X2 U878 ( .A1(opa_r[52]), .A2(opa_r[53]), .A3(n3079), .A4(n3080), .ZN(
        n3075) );
  NOR4_X2 U879 ( .A1(n3081), .A2(n4453), .A3(n4442), .A4(n4454), .ZN(n3080) );
  OAI22_X2 U882 ( .A1(n6303), .A2(n4626), .B1(n4614), .B2(n4603), .ZN(n4266)
         );
  AND2_X2 U883 ( .A1(n3073), .A2(n4273), .ZN(n4267) );
  AND4_X2 U884 ( .A1(n3082), .A2(n3083), .A3(n3084), .A4(n3085), .ZN(n3073) );
  NOR4_X2 U885 ( .A1(n3086), .A2(n3087), .A3(fracta_mul[2]), .A4(
        fracta_mul[23]), .ZN(n3085) );
  NAND4_X2 U887 ( .A1(n4277), .A2(n4367), .A3(n4478), .A4(n3088), .ZN(n3086)
         );
  NOR4_X2 U889 ( .A1(n3089), .A2(fracta_mul[20]), .A3(fracta_mul[22]), .A4(
        fracta_mul[21]), .ZN(n3084) );
  NAND2_X2 U890 ( .A1(n4322), .A2(n4373), .ZN(n3089) );
  AND2_X2 U892 ( .A1(n3091), .A2(n3092), .ZN(n3082) );
  NAND4_X2 U893 ( .A1(n4270), .A2(n4275), .A3(n3093), .A4(n3094), .ZN(\u6/N52 ) );
  NOR4_X2 U894 ( .A1(n3095), .A2(opb_r[60]), .A3(opb_r[62]), .A4(opb_r[61]), 
        .ZN(n3094) );
  NAND4_X2 U898 ( .A1(n3096), .A2(n3097), .A3(n3098), .A4(n3099), .ZN(n3072)
         );
  NOR4_X2 U899 ( .A1(n3100), .A2(n3101), .A3(n3102), .A4(n3103), .ZN(n3099) );
  NAND4_X2 U900 ( .A1(n4323), .A2(n4460), .A3(n4364), .A4(n3104), .ZN(n3103)
         );
  NAND4_X2 U902 ( .A1(n4324), .A2(n4461), .A3(n4365), .A4(n3105), .ZN(n3102)
         );
  NAND4_X2 U904 ( .A1(n4325), .A2(n4462), .A3(n4366), .A4(n3106), .ZN(n3101)
         );
  OR4_X2 U906 ( .A1(\u6/N27 ), .A2(\u6/N28 ), .A3(\u6/N26 ), .A4(n3107), .ZN(
        n3100) );
  OR4_X2 U907 ( .A1(\u6/N31 ), .A2(\u6/N30 ), .A3(\u6/N2 ), .A4(\u6/N29 ), 
        .ZN(n3107) );
  OR3_X2 U909 ( .A1(\u6/N50 ), .A2(\u6/N5 ), .A3(\u6/N4 ), .ZN(n3110) );
  OR4_X2 U910 ( .A1(\u6/N6 ), .A2(\u6/N7 ), .A3(\u6/N8 ), .A4(\u6/N9 ), .ZN(
        n3109) );
  OR4_X2 U911 ( .A1(\u6/N45 ), .A2(\u6/N46 ), .A3(\u6/N44 ), .A4(n3111), .ZN(
        n3108) );
  OR3_X2 U912 ( .A1(\u6/N47 ), .A2(\u6/N49 ), .A3(\u6/N48 ), .ZN(n3111) );
  NOR4_X2 U913 ( .A1(n3112), .A2(\u6/N38 ), .A3(\u6/N3 ), .A4(\u6/N39 ), .ZN(
        n3097) );
  OR4_X2 U914 ( .A1(\u6/N40 ), .A2(\u6/N41 ), .A3(\u6/N42 ), .A4(\u6/N43 ), 
        .ZN(n3112) );
  NOR4_X2 U915 ( .A1(n3113), .A2(\u6/N32 ), .A3(\u6/N34 ), .A4(\u6/N33 ), .ZN(
        n3096) );
  OR3_X2 U916 ( .A1(\u6/N36 ), .A2(\u6/N37 ), .A3(\u6/N35 ), .ZN(n3113) );
  AOI22_X2 U917 ( .A1(\u3/N69 ), .A2(n4659), .B1(\u3/N12 ), .B2(n4657), .ZN(
        n3114) );
  AOI22_X2 U918 ( .A1(\u3/N68 ), .A2(n4659), .B1(\u3/N11 ), .B2(n4658), .ZN(
        n3115) );
  AOI22_X2 U919 ( .A1(\u3/N67 ), .A2(n4659), .B1(\u3/N10 ), .B2(n4657), .ZN(
        n3116) );
  AOI22_X2 U920 ( .A1(\u3/N66 ), .A2(n4305), .B1(\u3/N9 ), .B2(n4658), .ZN(
        n3117) );
  AOI22_X2 U921 ( .A1(\u3/N65 ), .A2(n4659), .B1(\u3/N8 ), .B2(n4657), .ZN(
        n3118) );
  AOI22_X2 U922 ( .A1(\u3/N115 ), .A2(n4305), .B1(\u3/N58 ), .B2(n4658), .ZN(
        n3119) );
  AOI22_X2 U923 ( .A1(\u3/N114 ), .A2(n4659), .B1(\u3/N57 ), .B2(n4657), .ZN(
        n3120) );
  AOI22_X2 U924 ( .A1(\u3/N113 ), .A2(n4305), .B1(\u3/N56 ), .B2(n4658), .ZN(
        n3121) );
  AOI22_X2 U925 ( .A1(\u3/N112 ), .A2(n4659), .B1(\u3/N55 ), .B2(n4657), .ZN(
        n3122) );
  AOI22_X2 U926 ( .A1(\u3/N111 ), .A2(n4305), .B1(\u3/N54 ), .B2(n4658), .ZN(
        n3123) );
  AOI22_X2 U927 ( .A1(\u3/N110 ), .A2(n4659), .B1(\u3/N53 ), .B2(n4657), .ZN(
        n3124) );
  AOI22_X2 U928 ( .A1(\u3/N64 ), .A2(n4305), .B1(\u3/N7 ), .B2(n4657), .ZN(
        n3125) );
  AOI22_X2 U929 ( .A1(\u3/N109 ), .A2(n4659), .B1(\u3/N52 ), .B2(n4657), .ZN(
        n3126) );
  AOI22_X2 U930 ( .A1(\u3/N108 ), .A2(n4305), .B1(\u3/N51 ), .B2(n4657), .ZN(
        n3127) );
  AOI22_X2 U931 ( .A1(\u3/N107 ), .A2(n4659), .B1(\u3/N50 ), .B2(n4657), .ZN(
        n3128) );
  AOI22_X2 U932 ( .A1(\u3/N106 ), .A2(n4305), .B1(\u3/N49 ), .B2(n4657), .ZN(
        n3129) );
  AOI22_X2 U933 ( .A1(\u3/N105 ), .A2(n4659), .B1(\u3/N48 ), .B2(n4657), .ZN(
        n3130) );
  AOI22_X2 U934 ( .A1(\u3/N104 ), .A2(n4305), .B1(\u3/N47 ), .B2(n4657), .ZN(
        n3131) );
  AOI22_X2 U935 ( .A1(\u3/N103 ), .A2(n4305), .B1(\u3/N46 ), .B2(n4657), .ZN(
        n3132) );
  AOI22_X2 U936 ( .A1(\u3/N102 ), .A2(n4305), .B1(\u3/N45 ), .B2(n4657), .ZN(
        n3133) );
  AOI22_X2 U937 ( .A1(\u3/N101 ), .A2(n4305), .B1(\u3/N44 ), .B2(n4657), .ZN(
        n3134) );
  AOI22_X2 U938 ( .A1(\u3/N100 ), .A2(n4305), .B1(\u3/N43 ), .B2(n4657), .ZN(
        n3135) );
  AOI22_X2 U939 ( .A1(\u3/N63 ), .A2(n4305), .B1(\u3/N6 ), .B2(n4658), .ZN(
        n3136) );
  AOI22_X2 U940 ( .A1(\u3/N99 ), .A2(n4305), .B1(\u3/N42 ), .B2(n4658), .ZN(
        n3137) );
  AOI22_X2 U941 ( .A1(\u3/N98 ), .A2(n4305), .B1(\u3/N41 ), .B2(n4658), .ZN(
        n3138) );
  AOI22_X2 U942 ( .A1(\u3/N97 ), .A2(n4305), .B1(\u3/N40 ), .B2(n4658), .ZN(
        n3139) );
  AOI22_X2 U943 ( .A1(\u3/N96 ), .A2(n4305), .B1(\u3/N39 ), .B2(n4658), .ZN(
        n3140) );
  AOI22_X2 U944 ( .A1(\u3/N95 ), .A2(n4305), .B1(\u3/N38 ), .B2(n4658), .ZN(
        n3141) );
  AOI22_X2 U945 ( .A1(\u3/N94 ), .A2(n4305), .B1(\u3/N37 ), .B2(n4658), .ZN(
        n3142) );
  AOI22_X2 U946 ( .A1(\u3/N93 ), .A2(n4305), .B1(\u3/N36 ), .B2(n4658), .ZN(
        n3143) );
  AOI22_X2 U947 ( .A1(\u3/N92 ), .A2(n4305), .B1(\u3/N35 ), .B2(n4658), .ZN(
        n3144) );
  AOI22_X2 U948 ( .A1(\u3/N91 ), .A2(n4305), .B1(\u3/N34 ), .B2(n4658), .ZN(
        n3145) );
  AOI22_X2 U949 ( .A1(\u3/N90 ), .A2(n4305), .B1(\u3/N33 ), .B2(n4658), .ZN(
        n3146) );
  AOI22_X2 U950 ( .A1(\u3/N62 ), .A2(n4305), .B1(\u3/N5 ), .B2(n4657), .ZN(
        n3147) );
  AOI22_X2 U951 ( .A1(\u3/N89 ), .A2(n4305), .B1(\u3/N32 ), .B2(n4658), .ZN(
        n3148) );
  AOI22_X2 U952 ( .A1(\u3/N88 ), .A2(n4659), .B1(\u3/N31 ), .B2(n4657), .ZN(
        n3149) );
  AOI22_X2 U953 ( .A1(\u3/N87 ), .A2(n4659), .B1(\u3/N30 ), .B2(n4658), .ZN(
        n3150) );
  AOI22_X2 U954 ( .A1(\u3/N86 ), .A2(n4659), .B1(\u3/N29 ), .B2(n4657), .ZN(
        n3151) );
  AOI22_X2 U955 ( .A1(\u3/N85 ), .A2(n4659), .B1(\u3/N28 ), .B2(n4658), .ZN(
        n3152) );
  AOI22_X2 U956 ( .A1(\u3/N84 ), .A2(n4659), .B1(\u3/N27 ), .B2(n4657), .ZN(
        n3153) );
  AOI22_X2 U957 ( .A1(\u3/N83 ), .A2(n4659), .B1(\u3/N26 ), .B2(n4658), .ZN(
        n3154) );
  AOI22_X2 U958 ( .A1(\u3/N82 ), .A2(n4659), .B1(\u3/N25 ), .B2(n4657), .ZN(
        n3155) );
  AOI22_X2 U959 ( .A1(\u3/N81 ), .A2(n4659), .B1(\u3/N24 ), .B2(n4658), .ZN(
        n3156) );
  AOI22_X2 U960 ( .A1(\u3/N80 ), .A2(n4659), .B1(\u3/N23 ), .B2(n4658), .ZN(
        n3157) );
  AOI22_X2 U961 ( .A1(\u3/N61 ), .A2(n4659), .B1(\u3/N4 ), .B2(fasu_op), .ZN(
        n3158) );
  AOI22_X2 U962 ( .A1(\u3/N79 ), .A2(n4659), .B1(\u3/N22 ), .B2(fasu_op), .ZN(
        n3159) );
  AOI22_X2 U963 ( .A1(\u3/N78 ), .A2(n4659), .B1(\u3/N21 ), .B2(fasu_op), .ZN(
        n3160) );
  AOI22_X2 U964 ( .A1(\u3/N77 ), .A2(n4659), .B1(\u3/N20 ), .B2(fasu_op), .ZN(
        n3161) );
  AOI22_X2 U965 ( .A1(\u3/N76 ), .A2(n4659), .B1(\u3/N19 ), .B2(fasu_op), .ZN(
        n3162) );
  AOI22_X2 U966 ( .A1(\u3/N75 ), .A2(n4659), .B1(\u3/N18 ), .B2(fasu_op), .ZN(
        n3163) );
  AOI22_X2 U967 ( .A1(\u3/N74 ), .A2(n4659), .B1(\u3/N17 ), .B2(fasu_op), .ZN(
        n3164) );
  AOI22_X2 U968 ( .A1(\u3/N73 ), .A2(n4659), .B1(\u3/N16 ), .B2(fasu_op), .ZN(
        n3165) );
  AOI22_X2 U969 ( .A1(\u3/N72 ), .A2(n4659), .B1(\u3/N15 ), .B2(fasu_op), .ZN(
        n3166) );
  AOI22_X2 U970 ( .A1(\u3/N71 ), .A2(n4659), .B1(\u3/N14 ), .B2(fasu_op), .ZN(
        n3167) );
  AOI22_X2 U971 ( .A1(\u3/N70 ), .A2(n4659), .B1(\u3/N13 ), .B2(fasu_op), .ZN(
        n3168) );
  AOI22_X2 U972 ( .A1(\u3/N60 ), .A2(n4659), .B1(\u3/N3 ), .B2(n4660), .ZN(
        n3169) );
  NAND2_X2 U974 ( .A1(quo[107]), .A2(opb_dn), .ZN(n3170) );
  OAI22_X2 U975 ( .A1(n4601), .A2(n4277), .B1(n4602), .B2(n5878), .ZN(\u6/N99 ) );
  AOI22_X2 U976 ( .A1(n4602), .A2(fracta_mul[43]), .B1(n4603), .B2(N299), .ZN(
        n3181) );
  OAI22_X2 U977 ( .A1(n4601), .A2(n4286), .B1(n4602), .B2(n5879), .ZN(\u6/N97 ) );
  OAI22_X2 U978 ( .A1(n4601), .A2(n4472), .B1(n4602), .B2(n5880), .ZN(\u6/N96 ) );
  AOI22_X2 U979 ( .A1(n4602), .A2(fracta_mul[40]), .B1(n4603), .B2(N296), .ZN(
        n3182) );
  OAI22_X2 U980 ( .A1(n4601), .A2(n4478), .B1(n4602), .B2(n5881), .ZN(\u6/N94 ) );
  OAI22_X2 U981 ( .A1(n4601), .A2(n4284), .B1(n4602), .B2(n5882), .ZN(\u6/N93 ) );
  OAI22_X2 U982 ( .A1(n4601), .A2(n4272), .B1(n4602), .B2(n5883), .ZN(\u6/N92 ) );
  OAI22_X2 U983 ( .A1(n4601), .A2(n4276), .B1(n4602), .B2(n5884), .ZN(\u6/N91 ) );
  OAI22_X2 U984 ( .A1(n4601), .A2(n4474), .B1(n4602), .B2(n5885), .ZN(\u6/N90 ) );
  AOI22_X2 U985 ( .A1(n4602), .A2(fracta_mul[34]), .B1(n4603), .B2(N290), .ZN(
        n3183) );
  AOI22_X2 U986 ( .A1(n4602), .A2(fracta_mul[33]), .B1(n4603), .B2(N289), .ZN(
        n3184) );
  OAI22_X2 U987 ( .A1(n4601), .A2(n4287), .B1(n4602), .B2(n5886), .ZN(\u6/N87 ) );
  OAI22_X2 U988 ( .A1(n4601), .A2(n4370), .B1(n4602), .B2(n5887), .ZN(\u6/N86 ) );
  OAI22_X2 U989 ( .A1(n4601), .A2(n4479), .B1(n4602), .B2(n5888), .ZN(\u6/N85 ) );
  OAI22_X2 U990 ( .A1(n4601), .A2(n4475), .B1(n4602), .B2(n5889), .ZN(\u6/N84 ) );
  OAI22_X2 U991 ( .A1(n4601), .A2(n4285), .B1(n4602), .B2(n5890), .ZN(\u6/N83 ) );
  OAI22_X2 U992 ( .A1(n4601), .A2(n4301), .B1(n4602), .B2(n5891), .ZN(\u6/N82 ) );
  AOI22_X2 U993 ( .A1(n4602), .A2(fracta_mul[26]), .B1(n4603), .B2(N282), .ZN(
        n3185) );
  OAI22_X2 U994 ( .A1(n4601), .A2(n4473), .B1(n4602), .B2(n5892), .ZN(\u6/N80 ) );
  AOI22_X2 U995 ( .A1(n4602), .A2(fracta_mul[24]), .B1(n4603), .B2(N280), .ZN(
        n3186) );
  AOI22_X2 U996 ( .A1(n4602), .A2(fracta_mul[23]), .B1(n4603), .B2(N279), .ZN(
        n3187) );
  OAI22_X2 U997 ( .A1(n4603), .A2(n4283), .B1(n4602), .B2(n5893), .ZN(\u6/N77 ) );
  OAI22_X2 U998 ( .A1(n4603), .A2(n4292), .B1(n4602), .B2(n5894), .ZN(\u6/N76 ) );
  OAI22_X2 U999 ( .A1(n4603), .A2(n4320), .B1(n4602), .B2(n5895), .ZN(\u6/N75 ) );
  AOI22_X2 U1000 ( .A1(n4602), .A2(fracta_mul[19]), .B1(n4603), .B2(N275), 
        .ZN(n3188) );
  OAI22_X2 U1001 ( .A1(n4601), .A2(n4369), .B1(n4602), .B2(n5896), .ZN(
        \u6/N73 ) );
  OAI22_X2 U1002 ( .A1(n4601), .A2(n4319), .B1(n4602), .B2(n5897), .ZN(
        \u6/N72 ) );
  OAI22_X2 U1003 ( .A1(n4601), .A2(n4362), .B1(n4602), .B2(n5898), .ZN(
        \u6/N71 ) );
  OAI22_X2 U1004 ( .A1(n4601), .A2(n4318), .B1(n4602), .B2(n5899), .ZN(
        \u6/N70 ) );
  OAI22_X2 U1005 ( .A1(n4601), .A2(n4372), .B1(n4602), .B2(n5900), .ZN(
        \u6/N69 ) );
  AOI22_X2 U1006 ( .A1(n4602), .A2(fracta_mul[13]), .B1(n4603), .B2(N269), 
        .ZN(n3189) );
  OAI22_X2 U1007 ( .A1(n4601), .A2(n4374), .B1(n4602), .B2(n5901), .ZN(
        \u6/N67 ) );
  OAI22_X2 U1008 ( .A1(n4601), .A2(n4361), .B1(n4602), .B2(n5902), .ZN(
        \u6/N66 ) );
  OAI22_X2 U1009 ( .A1(n4601), .A2(n4300), .B1(n4602), .B2(n5903), .ZN(
        \u6/N65 ) );
  OAI22_X2 U1010 ( .A1(n4601), .A2(n4368), .B1(n4602), .B2(n5904), .ZN(
        \u6/N64 ) );
  OAI22_X2 U1011 ( .A1(n4601), .A2(n4326), .B1(n4602), .B2(n5905), .ZN(
        \u6/N63 ) );
  OAI22_X2 U1012 ( .A1(n4601), .A2(n4376), .B1(n4602), .B2(n5906), .ZN(
        \u6/N62 ) );
  OAI22_X2 U1013 ( .A1(n4601), .A2(n4375), .B1(n4602), .B2(n5907), .ZN(
        \u6/N61 ) );
  OAI22_X2 U1014 ( .A1(n4601), .A2(n4371), .B1(n4602), .B2(n5908), .ZN(
        \u6/N60 ) );
  AOI22_X2 U1015 ( .A1(n4602), .A2(fracta_mul[4]), .B1(n4603), .B2(N260), .ZN(
        n3190) );
  OAI22_X2 U1016 ( .A1(n4601), .A2(n4360), .B1(n4602), .B2(n5909), .ZN(
        \u6/N58 ) );
  AOI22_X2 U1017 ( .A1(n4602), .A2(fracta_mul[2]), .B1(n4603), .B2(N258), .ZN(
        n3191) );
  OAI22_X2 U1018 ( .A1(n4601), .A2(n4373), .B1(n4602), .B2(n5910), .ZN(
        \u6/N56 ) );
  OAI22_X2 U1019 ( .A1(n4601), .A2(n4322), .B1(n4602), .B2(n5911), .ZN(
        \u6/N55 ) );
  OR2_X2 U1020 ( .A1(N308), .A2(n4602), .ZN(\u6/N107 ) );
  OAI22_X2 U1021 ( .A1(n4601), .A2(n4273), .B1(n4602), .B2(n5874), .ZN(
        \u6/N106 ) );
  OAI22_X2 U1022 ( .A1(n4601), .A2(n4480), .B1(n4602), .B2(n5875), .ZN(
        \u6/N105 ) );
  AOI22_X2 U1023 ( .A1(n4602), .A2(fracta_mul[49]), .B1(n4603), .B2(N305), 
        .ZN(n3192) );
  AOI22_X2 U1024 ( .A1(n4602), .A2(fracta_mul[48]), .B1(n4603), .B2(N304), 
        .ZN(n3193) );
  AOI22_X2 U1025 ( .A1(n4602), .A2(fracta_mul[47]), .B1(n4603), .B2(N303), 
        .ZN(n3194) );
  OAI22_X2 U1026 ( .A1(n4601), .A2(n4477), .B1(n4602), .B2(n5876), .ZN(
        \u6/N101 ) );
  OAI22_X2 U1027 ( .A1(n4601), .A2(n4367), .B1(n4602), .B2(n5877), .ZN(
        \u6/N100 ) );
  NAND4_X2 U1028 ( .A1(n4449), .A2(n4450), .A3(n3195), .A4(n3196), .ZN(
        \u2/N157 ) );
  NOR4_X2 U1029 ( .A1(n3197), .A2(opa_r[60]), .A3(opa_r[62]), .A4(opa_r[61]), 
        .ZN(n3196) );
  NAND4_X2 U1032 ( .A1(n6282), .A2(n3198), .A3(n6280), .A4(n3199), .ZN(
        div_opa_ldz_d[4]) );
  NOR4_X2 U1033 ( .A1(n6292), .A2(n3200), .A3(n3201), .A4(n3202), .ZN(n3199)
         );
  NAND4_X2 U1038 ( .A1(n3210), .A2(n3211), .A3(n3212), .A4(n3213), .ZN(
        div_opa_ldz_d[3]) );
  NOR4_X2 U1039 ( .A1(n3214), .A2(n3215), .A3(n6294), .A4(n3216), .ZN(n3213)
         );
  NOR4_X2 U1040 ( .A1(fracta_mul[29]), .A2(n3217), .A3(n4285), .A4(n6279), 
        .ZN(n3216) );
  OAI22_X2 U1042 ( .A1(n4301), .A2(n3220), .B1(n3221), .B2(n3204), .ZN(n3214)
         );
  NAND2_X2 U1047 ( .A1(n3231), .A2(n3232), .ZN(div_opa_ldz_d[2]) );
  NOR4_X2 U1048 ( .A1(n3233), .A2(n3234), .A3(n6285), .A4(n3235), .ZN(n3232)
         );
  NOR4_X2 U1049 ( .A1(fracta_mul[33]), .A2(n6298), .A3(n4287), .A4(n6279), 
        .ZN(n3235) );
  AND3_X2 U1050 ( .A1(fracta_mul[48]), .A2(n4273), .A3(n3237), .ZN(n3234) );
  OAI222_X2 U1053 ( .A1(fracta_mul[26]), .A2(n3228), .B1(n3243), .B2(n3218), 
        .C1(n3244), .C2(n3204), .ZN(n3241) );
  AOI221_X2 U1054 ( .B1(n3223), .B2(n3245), .C1(fracta_mul[14]), .C2(n3246), 
        .A(n3247), .ZN(n3244) );
  OR2_X2 U1055 ( .A1(fracta_mul[18]), .A2(fracta_mul[19]), .ZN(n3248) );
  OR4_X2 U1059 ( .A1(n3249), .A2(n3250), .A3(n3251), .A4(n3252), .ZN(
        div_opa_ldz_d[1]) );
  NAND4_X2 U1060 ( .A1(n3207), .A2(n3253), .A3(n3254), .A4(n3255), .ZN(n3252)
         );
  NOR4_X2 U1061 ( .A1(n3256), .A2(n6291), .A3(n3257), .A4(n3258), .ZN(n3255)
         );
  NAND4_X2 U1063 ( .A1(n3260), .A2(fracta_mul[30]), .A3(n3261), .A4(n4370), 
        .ZN(n3207) );
  OAI211_X2 U1064 ( .C1(fracta_mul[51]), .C2(n3237), .A(n3230), .B(n3210), 
        .ZN(n3251) );
  AND4_X2 U1065 ( .A1(n3238), .A2(n6289), .A3(n3236), .A4(n3262), .ZN(n3210)
         );
  NOR4_X2 U1066 ( .A1(n3263), .A2(n3264), .A3(n3265), .A4(n6286), .ZN(n3262)
         );
  NAND2_X2 U1068 ( .A1(n3269), .A2(fracta_mul[38]), .ZN(n3238) );
  NAND2_X2 U1070 ( .A1(n3271), .A2(fracta_mul[22]), .ZN(n3239) );
  NAND4_X2 U1074 ( .A1(n6277), .A2(n3211), .A3(n3276), .A4(n3277), .ZN(
        div_opa_ldz_d[0]) );
  NOR4_X2 U1075 ( .A1(n3278), .A2(n3270), .A3(fracta_mul[51]), .A4(n3263), 
        .ZN(n3277) );
  NAND2_X2 U1078 ( .A1(n6284), .A2(n4301), .ZN(n3272) );
  NAND4_X2 U1083 ( .A1(n3253), .A2(n3259), .A3(n3280), .A4(n3281), .ZN(n3209)
         );
  AOI22_X2 U1084 ( .A1(n6284), .A2(fracta_mul[27]), .B1(n3260), .B2(
        fracta_mul[35]), .ZN(n3281) );
  OR4_X2 U1087 ( .A1(n3204), .A2(n4373), .A3(n3090), .A4(fracta_mul[2]), .ZN(
        n3253) );
  NAND2_X2 U1088 ( .A1(n3282), .A2(n4360), .ZN(n3090) );
  AOI22_X2 U1090 ( .A1(fracta_mul[43]), .A2(n3226), .B1(fracta_mul[11]), .B2(
        n6287), .ZN(n3211) );
  NAND4_X2 U1091 ( .A1(n6278), .A2(n3198), .A3(n3285), .A4(n3286), .ZN(n3242)
         );
  NAND2_X2 U1094 ( .A1(n3267), .A2(n4375), .ZN(n3205) );
  OR3_X2 U1097 ( .A1(n3264), .A2(n3256), .A3(n6283), .ZN(n3287) );
  AND3_X2 U1104 ( .A1(fracta_mul[31]), .A2(n3261), .A3(n3260), .ZN(n3291) );
  AND3_X2 U1106 ( .A1(fracta_mul[21]), .A2(n4283), .A3(n3271), .ZN(n3265) );
  NAND2_X2 U1109 ( .A1(n6288), .A2(n3222), .ZN(n3284) );
  NOR4_X2 U1112 ( .A1(fracta_mul[16]), .A2(fracta_mul[17]), .A3(fracta_mul[18]), .A4(fracta_mul[19]), .ZN(n3246) );
  NAND2_X2 U1115 ( .A1(n3260), .A2(n3091), .ZN(n3220) );
  NAND2_X2 U1121 ( .A1(n3269), .A2(n4284), .ZN(n3206) );
  NOR4_X2 U1123 ( .A1(fracta_mul[24]), .A2(fracta_mul[25]), .A3(fracta_mul[26]), .A4(fracta_mul[27]), .ZN(n3289) );
  OR2_X2 U1125 ( .A1(fracta_mul[42]), .A2(fracta_mul[43]), .ZN(n3243) );
  OR3_X2 U1127 ( .A1(fracta_mul[46]), .A2(fracta_mul[47]), .A3(n6295), .ZN(
        n3219) );
  AOI22_X2 U1130 ( .A1(\u3/N116 ), .A2(n4659), .B1(\u3/N59 ), .B2(n4660), .ZN(
        n3292) );
  NOR4_X2 U1131 ( .A1(n3293), .A2(n3294), .A3(n4489), .A4(n4384), .ZN(N923) );
  NAND4_X2 U1133 ( .A1(exp_mul[3]), .A2(exp_mul[2]), .A3(exp_mul[4]), .A4(
        n3295), .ZN(n3293) );
  AND4_X2 U1135 ( .A1(opb_00), .A2(opa_nan_r), .A3(n4486), .A4(n4382), .ZN(
        N913) );
  OAI211_X2 U1137 ( .C1(n3297), .C2(n3298), .A(n3299), .B(n3300), .ZN(N911) );
  NOR4_X2 U1139 ( .A1(n3304), .A2(n3305), .A3(n2507), .A4(n3306), .ZN(n3301)
         );
  OR2_X2 U1140 ( .A1(inf_mul2), .A2(inf_mul_r), .ZN(n3305) );
  NAND4_X2 U1141 ( .A1(n6341), .A2(n3307), .A3(n3308), .A4(n3309), .ZN(n3299)
         );
  OAI221_X2 U1143 ( .B1(n3310), .B2(n3311), .C1(n3312), .C2(n6458), .A(n3313), 
        .ZN(N906) );
  AND3_X2 U1146 ( .A1(fasu_op_r2), .A2(n3315), .A3(inf_d), .ZN(n3317) );
  NAND4_X2 U1148 ( .A1(n3321), .A2(n3322), .A3(n3323), .A4(n3324), .ZN(n3318)
         );
  NOR4_X2 U1149 ( .A1(n3325), .A2(n3326), .A3(n3327), .A4(n3328), .ZN(n3324)
         );
  NAND4_X2 U1150 ( .A1(n3329), .A2(n3330), .A3(n3331), .A4(n3332), .ZN(n3325)
         );
  NOR4_X2 U1151 ( .A1(n3333), .A2(n3334), .A3(n3335), .A4(n3336), .ZN(n3323)
         );
  NAND4_X2 U1152 ( .A1(n3337), .A2(n3338), .A3(n3339), .A4(n3340), .ZN(n3333)
         );
  AOI22_X2 U1153 ( .A1(opb_00), .A2(n4486), .B1(opa_inf), .B2(n4327), .ZN(
        n3310) );
  AOI221_X2 U1155 ( .B1(underflow_fmul_r[2]), .B2(n3345), .C1(
        underflow_fmul_r[1]), .C2(n3346), .A(n3347), .ZN(n3344) );
  OR2_X2 U1156 ( .A1(underflow_fmul_r[0]), .A2(n3348), .ZN(n3347) );
  NOR4_X2 U1157 ( .A1(n6447), .A2(n3304), .A3(n3349), .A4(n4485), .ZN(n3348)
         );
  NOR4_X2 U1158 ( .A1(n3350), .A2(n3351), .A3(n3352), .A4(n3353), .ZN(n3349)
         );
  NAND4_X2 U1159 ( .A1(n3354), .A2(n3355), .A3(n3356), .A4(n3357), .ZN(n3353)
         );
  NOR4_X2 U1160 ( .A1(n3358), .A2(prod[21]), .A3(prod[23]), .A4(prod[22]), 
        .ZN(n3357) );
  OR4_X2 U1161 ( .A1(prod[24]), .A2(prod[25]), .A3(prod[26]), .A4(prod[27]), 
        .ZN(n3358) );
  NOR4_X2 U1162 ( .A1(n3359), .A2(prod[16]), .A3(prod[18]), .A4(prod[17]), 
        .ZN(n3356) );
  OR3_X2 U1163 ( .A1(prod[1]), .A2(prod[20]), .A3(prod[19]), .ZN(n3359) );
  NOR4_X2 U1164 ( .A1(n3360), .A2(prod[105]), .A3(prod[11]), .A4(prod[10]), 
        .ZN(n3355) );
  OR4_X2 U1165 ( .A1(prod[12]), .A2(prod[13]), .A3(prod[14]), .A4(prod[15]), 
        .ZN(n3360) );
  NOR4_X2 U1166 ( .A1(n3361), .A2(prod[0]), .A3(prod[101]), .A4(prod[100]), 
        .ZN(n3354) );
  NAND4_X2 U1168 ( .A1(n3362), .A2(n3363), .A3(n3364), .A4(n3365), .ZN(n3352)
         );
  NOR4_X2 U1169 ( .A1(n3366), .A2(prod[46]), .A3(prod[48]), .A4(prod[47]), 
        .ZN(n3365) );
  OR4_X2 U1170 ( .A1(prod[49]), .A2(prod[4]), .A3(prod[50]), .A4(prod[51]), 
        .ZN(n3366) );
  NOR4_X2 U1171 ( .A1(n3367), .A2(prod[3]), .A3(prod[41]), .A4(prod[40]), .ZN(
        n3364) );
  OR4_X2 U1172 ( .A1(prod[42]), .A2(prod[43]), .A3(prod[44]), .A4(prod[45]), 
        .ZN(n3367) );
  NOR4_X2 U1173 ( .A1(n3368), .A2(prod[33]), .A3(prod[35]), .A4(prod[34]), 
        .ZN(n3363) );
  OR4_X2 U1174 ( .A1(prod[36]), .A2(prod[37]), .A3(prod[38]), .A4(prod[39]), 
        .ZN(n3368) );
  NOR4_X2 U1175 ( .A1(n3369), .A2(prod[28]), .A3(prod[2]), .A4(prod[29]), .ZN(
        n3362) );
  OR3_X2 U1176 ( .A1(prod[31]), .A2(prod[32]), .A3(prod[30]), .ZN(n3369) );
  NAND4_X2 U1177 ( .A1(n3370), .A2(n3371), .A3(n3372), .A4(n3373), .ZN(n3351)
         );
  NOR4_X2 U1178 ( .A1(n3374), .A2(prod[6]), .A3(prod[71]), .A4(prod[70]), .ZN(
        n3373) );
  NAND4_X2 U1179 ( .A1(n4313), .A2(n4407), .A3(n4298), .A4(n4343), .ZN(n3374)
         );
  NOR4_X2 U1180 ( .A1(n3375), .A2(prod[64]), .A3(prod[66]), .A4(prod[65]), 
        .ZN(n3372) );
  NOR4_X2 U1182 ( .A1(n3376), .A2(prod[58]), .A3(prod[5]), .A4(prod[59]), .ZN(
        n3371) );
  NAND4_X2 U1183 ( .A1(n4346), .A2(n4406), .A3(n4312), .A4(n4297), .ZN(n3376)
         );
  NOR4_X2 U1184 ( .A1(n3377), .A2(prod[52]), .A3(prod[54]), .A4(prod[53]), 
        .ZN(n3370) );
  NAND4_X2 U1186 ( .A1(n3378), .A2(n3379), .A3(n3380), .A4(n3381), .ZN(n3350)
         );
  NOR4_X2 U1187 ( .A1(n3382), .A2(prod[94]), .A3(prod[96]), .A4(prod[95]), 
        .ZN(n3381) );
  OR4_X2 U1188 ( .A1(prod[97]), .A2(prod[98]), .A3(prod[99]), .A4(prod[9]), 
        .ZN(n3382) );
  NOR4_X2 U1189 ( .A1(n3383), .A2(prod[88]), .A3(prod[8]), .A4(prod[89]), .ZN(
        n3380) );
  NAND4_X2 U1190 ( .A1(n4345), .A2(n4405), .A3(n4308), .A4(n4295), .ZN(n3383)
         );
  NOR4_X2 U1191 ( .A1(n3384), .A2(prod[81]), .A3(prod[83]), .A4(prod[82]), 
        .ZN(n3379) );
  NAND4_X2 U1192 ( .A1(n4344), .A2(n4404), .A3(n4307), .A4(n4294), .ZN(n3384)
         );
  NOR4_X2 U1193 ( .A1(n3385), .A2(prod[76]), .A3(prod[78]), .A4(prod[77]), 
        .ZN(n3378) );
  OR3_X2 U1194 ( .A1(prod[7]), .A2(prod[80]), .A3(prod[79]), .ZN(n3385) );
  NAND4_X2 U1196 ( .A1(n3388), .A2(n3389), .A3(n3390), .A4(n3391), .ZN(n3387)
         );
  NOR4_X2 U1197 ( .A1(n3392), .A2(n3393), .A3(n3394), .A4(n3395), .ZN(n3391)
         );
  AND3_X2 U1198 ( .A1(n3396), .A2(n3397), .A3(n3398), .ZN(n3390) );
  NAND4_X2 U1199 ( .A1(n3399), .A2(n3400), .A3(n3401), .A4(n3402), .ZN(n3319)
         );
  NOR4_X2 U1200 ( .A1(n3403), .A2(n3404), .A3(n3405), .A4(n3406), .ZN(n3402)
         );
  NAND4_X2 U1201 ( .A1(n3407), .A2(n3408), .A3(n3409), .A4(n3410), .ZN(n3403)
         );
  NOR4_X2 U1202 ( .A1(n3411), .A2(n3412), .A3(n3413), .A4(n3414), .ZN(n3401)
         );
  NOR4_X2 U1204 ( .A1(n3418), .A2(n3419), .A3(n3420), .A4(n3421), .ZN(n3400)
         );
  NAND4_X2 U1205 ( .A1(n3422), .A2(n3423), .A3(n3424), .A4(n3425), .ZN(n3418)
         );
  NOR4_X2 U1206 ( .A1(n3426), .A2(n3427), .A3(n3428), .A4(n3429), .ZN(n3399)
         );
  NAND4_X2 U1208 ( .A1(n3321), .A2(n3322), .A3(n3433), .A4(n3434), .ZN(n3386)
         );
  NOR4_X2 U1209 ( .A1(n3435), .A2(n3436), .A3(n3328), .A4(n3326), .ZN(n3434)
         );
  NAND4_X2 U1210 ( .A1(n3437), .A2(n3329), .A3(n3330), .A4(n3331), .ZN(n3435)
         );
  NOR4_X2 U1211 ( .A1(n3438), .A2(n3334), .A3(n3335), .A4(n3336), .ZN(n3433)
         );
  NOR4_X2 U1213 ( .A1(n3439), .A2(n3440), .A3(n3441), .A4(n3442), .ZN(n3322)
         );
  NAND4_X2 U1214 ( .A1(n3443), .A2(n3444), .A3(n3445), .A4(n3446), .ZN(n3439)
         );
  NOR4_X2 U1215 ( .A1(n3447), .A2(n3448), .A3(n3449), .A4(n3450), .ZN(n3321)
         );
  OAI221_X2 U1218 ( .B1(n3460), .B2(n6449), .C1(n3461), .C2(n4291), .A(n3462), 
        .ZN(N889) );
  AOI22_X2 U1221 ( .A1(n3464), .A2(n6316), .B1(n4540), .B2(n3463), .ZN(n3460)
         );
  AND2_X2 U1223 ( .A1(n3320), .A2(n3304), .ZN(n3466) );
  NAND2_X2 U1226 ( .A1(n4327), .A2(n4382), .ZN(n3306) );
  INV_X4 U1229 ( .A(n3346), .ZN(n3342) );
  NAND2_X2 U1231 ( .A1(n6316), .A2(n3472), .ZN(n3471) );
  NOR4_X2 U1232 ( .A1(exp_ovf_r[1]), .A2(n6465), .A3(\u4/exp_in_mi1[11] ), 
        .A4(n3476), .ZN(n3474) );
  OR3_X2 U1233 ( .A1(n4355), .A2(n3477), .A3(n3478), .ZN(n3470) );
  OAI211_X2 U1234 ( .C1(n3479), .C2(n3480), .A(n3481), .B(n3482), .ZN(n3469)
         );
  AOI221_X2 U1239 ( .B1(\u4/N6279 ), .B2(n3490), .C1(n3491), .C2(exp_ovf_r[1]), 
        .A(n3492), .ZN(n3483) );
  INV_X4 U1240 ( .A(n3493), .ZN(n3492) );
  AND4_X2 U1242 ( .A1(\u4/N6286 ), .A2(n3496), .A3(n3497), .A4(n3498), .ZN(
        n3494) );
  NOR4_X2 U1243 ( .A1(n3499), .A2(exp_r[3]), .A3(n4290), .A4(n4282), .ZN(n3498) );
  OR3_X2 U1244 ( .A1(n4281), .A2(n4353), .A3(exp_r[6]), .ZN(n3499) );
  INV_X4 U1246 ( .A(n2518), .ZN(n3496) );
  XOR2_X2 U1249 ( .A(n4656), .B(n5864), .Z(n3503) );
  NOR4_X2 U1250 ( .A1(n3505), .A2(n5868), .A3(n5870), .A4(n5869), .ZN(n3502)
         );
  NAND2_X2 U1252 ( .A1(\u4/div_exp3 [5]), .A2(n2394), .ZN(n3508) );
  NAND2_X2 U1255 ( .A1(\u4/div_exp3 [4]), .A2(n2394), .ZN(n3511) );
  NAND2_X2 U1258 ( .A1(\u4/div_exp3 [6]), .A2(n4542), .ZN(n3514) );
  NAND2_X2 U1262 ( .A1(\u4/div_exp3 [3]), .A2(n2394), .ZN(n3516) );
  NAND2_X2 U1265 ( .A1(\u4/div_exp3 [1]), .A2(n2394), .ZN(n3518) );
  NAND2_X2 U1268 ( .A1(\u4/div_exp3 [2]), .A2(n2394), .ZN(n3520) );
  NOR4_X2 U1270 ( .A1(n3504), .A2(n3521), .A3(n2430), .A4(n2427), .ZN(n3501)
         );
  NAND2_X2 U1272 ( .A1(\u4/div_exp3 [8]), .A2(n2394), .ZN(n3523) );
  NAND2_X2 U1275 ( .A1(\u4/div_exp3 [9]), .A2(n4542), .ZN(n3525) );
  NAND2_X2 U1277 ( .A1(n6465), .A2(n2423), .ZN(n3521) );
  NAND2_X2 U1279 ( .A1(\u4/div_exp3 [7]), .A2(n4542), .ZN(n3527) );
  NAND2_X2 U1282 ( .A1(\u4/div_exp3 [10]), .A2(n2394), .ZN(n3529) );
  OAI22_X2 U1287 ( .A1(exp_ovf_r[1]), .A2(n3530), .B1(n4452), .B2(n3531), .ZN(
        n3490) );
  AND2_X2 U1289 ( .A1(\u4/N6280 ), .A2(n3495), .ZN(n3532) );
  INV_X4 U1290 ( .A(n3533), .ZN(n3530) );
  NAND4_X2 U1291 ( .A1(n3397), .A2(n3534), .A3(n3535), .A4(n3536), .ZN(n3480)
         );
  NAND4_X2 U1292 ( .A1(n3537), .A2(n3392), .A3(n3538), .A4(n3393), .ZN(n3479)
         );
  INV_X4 U1294 ( .A(n3541), .ZN(n3461) );
  OAI221_X2 U1295 ( .B1(n2433), .B2(n3475), .C1(n3542), .C2(n2434), .A(n3543), 
        .ZN(n3541) );
  AOI221_X2 U1296 ( .B1(n3544), .B2(n3545), .C1(n4540), .C2(n3495), .A(n3477), 
        .ZN(n3543) );
  NOR4_X2 U1299 ( .A1(n4656), .A2(n6307), .A3(n4441), .A4(n4351), .ZN(n3546)
         );
  INV_X4 U1300 ( .A(n3485), .ZN(n3475) );
  AOI22_X2 U1301 ( .A1(n3549), .A2(n4540), .B1(n4355), .B2(n3550), .ZN(n3456)
         );
  OAI211_X2 U1303 ( .C1(n3551), .C2(n4356), .A(n3553), .B(n3554), .ZN(n3549)
         );
  AND3_X2 U1305 ( .A1(n4352), .A2(n3488), .A3(n3557), .ZN(n3555) );
  NAND4_X2 U1307 ( .A1(n3302), .A2(n3303), .A3(opas_r2), .A4(n6308), .ZN(n3559) );
  AOI22_X2 U1308 ( .A1(n6314), .A2(n3560), .B1(n3561), .B2(n3343), .ZN(n3558)
         );
  OAI22_X2 U1309 ( .A1(n6341), .A2(n3562), .B1(n3563), .B2(n3311), .ZN(n3561)
         );
  AOI22_X2 U1310 ( .A1(n3564), .A2(n6455), .B1(n3565), .B2(n4491), .ZN(n3563)
         );
  NAND2_X2 U1312 ( .A1(opb_inf), .A2(opa_inf), .ZN(n3309) );
  NAND2_X2 U1313 ( .A1(n4491), .A2(n3308), .ZN(n3564) );
  AOI22_X2 U1314 ( .A1(n3314), .A2(n3566), .B1(nan_sign_d), .B2(n6457), .ZN(
        n3562) );
  INV_X4 U1315 ( .A(n3567), .ZN(n3566) );
  AOI22_X2 U1316 ( .A1(sign_fasu_r), .A2(n3298), .B1(result_zero_sign_d), .B2(
        n3568), .ZN(n3567) );
  INV_X4 U1317 ( .A(n3568), .ZN(n3298) );
  NAND2_X2 U1321 ( .A1(n3303), .A2(n4540), .ZN(n3311) );
  XOR2_X2 U1322 ( .A(sign_mul_r), .B(n3569), .Z(n3560) );
  NAND2_X2 U1324 ( .A1(n3303), .A2(n6316), .ZN(n3343) );
  NAND4_X2 U1326 ( .A1(n3570), .A2(n3571), .A3(n3572), .A4(n3573), .ZN(n3304)
         );
  NOR4_X2 U1327 ( .A1(n3574), .A2(n3575), .A3(n3576), .A4(n3577), .ZN(n3573)
         );
  NAND4_X2 U1328 ( .A1(n3445), .A2(n3446), .A3(n3578), .A4(n3579), .ZN(n3577)
         );
  NAND4_X2 U1329 ( .A1(n3580), .A2(n3337), .A3(n3338), .A4(n3339), .ZN(n3576)
         );
  NAND4_X2 U1330 ( .A1(n3340), .A2(n3581), .A3(n3582), .A4(n3437), .ZN(n3575)
         );
  NAND4_X2 U1331 ( .A1(n3329), .A2(n3330), .A3(n3331), .A4(n3397), .ZN(n3574)
         );
  NOR4_X2 U1333 ( .A1(n3586), .A2(n3587), .A3(n3588), .A4(n3589), .ZN(n3572)
         );
  NAND4_X2 U1335 ( .A1(n3410), .A2(n3590), .A3(n3591), .A4(n3592), .ZN(n3588)
         );
  NAND4_X2 U1336 ( .A1(n3453), .A2(n3451), .A3(n3452), .A4(n3593), .ZN(n3587)
         );
  NAND4_X2 U1337 ( .A1(n3594), .A2(n3595), .A3(n3443), .A4(n3444), .ZN(n3586)
         );
  NOR4_X2 U1338 ( .A1(n3596), .A2(n3597), .A3(n3598), .A4(n3599), .ZN(n3571)
         );
  NAND4_X2 U1340 ( .A1(n3423), .A2(n3424), .A3(n3425), .A4(n3602), .ZN(n3598)
         );
  NAND4_X2 U1341 ( .A1(n3603), .A2(n3604), .A3(n3417), .A4(n3415), .ZN(n3597)
         );
  NAND4_X2 U1342 ( .A1(n3416), .A2(n3605), .A3(n3606), .A4(n3607), .ZN(n3596)
         );
  NAND4_X2 U1344 ( .A1(n3398), .A2(n3611), .A3(n3612), .A4(n3613), .ZN(n3610)
         );
  NAND4_X2 U1345 ( .A1(n3432), .A2(n3430), .A3(n3431), .A4(n3614), .ZN(n3609)
         );
  NAND4_X2 U1346 ( .A1(n3540), .A2(n3615), .A3(n3539), .A4(n3616), .ZN(n3608)
         );
  NOR4_X2 U1347 ( .A1(n3535), .A2(n3536), .A3(n3537), .A4(n3392), .ZN(n3616)
         );
  INV_X4 U1348 ( .A(n3617), .ZN(n3392) );
  INV_X4 U1349 ( .A(n3388), .ZN(n3537) );
  INV_X4 U1350 ( .A(n3389), .ZN(n3536) );
  INV_X4 U1351 ( .A(n3396), .ZN(n3535) );
  NAND2_X2 U1352 ( .A1(n3618), .A2(n3619), .ZN(N855) );
  OR2_X2 U1353 ( .A1(n3583), .A2(n6310), .ZN(N854) );
  OR2_X2 U1354 ( .A1(n3584), .A2(n6310), .ZN(N853) );
  NAND2_X2 U1355 ( .A1(n3539), .A2(n3619), .ZN(N852) );
  NAND2_X2 U1356 ( .A1(n3540), .A2(n3619), .ZN(N851) );
  NAND2_X2 U1357 ( .A1(n3615), .A2(n3619), .ZN(N850) );
  NAND2_X2 U1358 ( .A1(n3617), .A2(n3619), .ZN(N849) );
  NAND2_X2 U1359 ( .A1(n3388), .A2(n3619), .ZN(N848) );
  NAND2_X2 U1360 ( .A1(n3389), .A2(n3619), .ZN(N847) );
  NAND2_X2 U1361 ( .A1(n3396), .A2(n3619), .ZN(N846) );
  NAND2_X2 U1362 ( .A1(n3398), .A2(n3619), .ZN(N845) );
  INV_X4 U1364 ( .A(n3427), .ZN(n3611) );
  OAI221_X2 U1365 ( .B1(n4593), .B2(n3621), .C1(n2520), .C2(n4591), .A(n4588), 
        .ZN(n3427) );
  INV_X4 U1366 ( .A(\u4/fract_out_pl1[51] ), .ZN(n3621) );
  INV_X4 U1368 ( .A(n3429), .ZN(n3612) );
  OAI221_X2 U1369 ( .B1(n4593), .B2(n3624), .C1(n2521), .C2(n4591), .A(n4588), 
        .ZN(n3429) );
  INV_X4 U1370 ( .A(\u4/fract_out_pl1[50] ), .ZN(n3624) );
  INV_X4 U1372 ( .A(n3428), .ZN(n3613) );
  OAI221_X2 U1373 ( .B1(n4593), .B2(n3625), .C1(n3626), .C2(n4591), .A(n4588), 
        .ZN(n3428) );
  INV_X4 U1374 ( .A(\u4/fract_out_pl1[49] ), .ZN(n3625) );
  INV_X4 U1376 ( .A(n3627), .ZN(n3432) );
  OAI221_X2 U1377 ( .B1(n4593), .B2(n3628), .C1(n3629), .C2(n4591), .A(n4588), 
        .ZN(n3627) );
  INV_X4 U1378 ( .A(\u4/fract_out_pl1[48] ), .ZN(n3628) );
  INV_X4 U1380 ( .A(n3630), .ZN(n3430) );
  OAI221_X2 U1381 ( .B1(n4593), .B2(n3631), .C1(n2522), .C2(n4591), .A(n4588), 
        .ZN(n3630) );
  INV_X4 U1382 ( .A(\u4/fract_out_pl1[47] ), .ZN(n3631) );
  INV_X4 U1384 ( .A(n3632), .ZN(n3431) );
  OAI221_X2 U1385 ( .B1(n4593), .B2(n3633), .C1(n2523), .C2(n4591), .A(n4588), 
        .ZN(n3632) );
  INV_X4 U1386 ( .A(\u4/fract_out_pl1[46] ), .ZN(n3633) );
  INV_X4 U1388 ( .A(n3419), .ZN(n3614) );
  OAI221_X2 U1389 ( .B1(n4593), .B2(n3634), .C1(n2524), .C2(n4591), .A(n4588), 
        .ZN(n3419) );
  INV_X4 U1390 ( .A(\u4/fract_out_pl1[45] ), .ZN(n3634) );
  INV_X4 U1392 ( .A(n3421), .ZN(n3601) );
  OAI221_X2 U1393 ( .B1(n4593), .B2(n3635), .C1(n3636), .C2(n4591), .A(n4587), 
        .ZN(n3421) );
  INV_X4 U1394 ( .A(\u4/fract_out_pl1[44] ), .ZN(n3635) );
  INV_X4 U1396 ( .A(n3420), .ZN(n3600) );
  OAI221_X2 U1397 ( .B1(n4594), .B2(n3637), .C1(n3638), .C2(n4590), .A(n4588), 
        .ZN(n3420) );
  INV_X4 U1398 ( .A(\u4/fract_out_pl1[43] ), .ZN(n3637) );
  INV_X4 U1400 ( .A(n3639), .ZN(n3422) );
  OAI221_X2 U1401 ( .B1(n4594), .B2(n3640), .C1(n3641), .C2(n4590), .A(n4588), 
        .ZN(n3639) );
  INV_X4 U1402 ( .A(\u4/fract_out_pl1[42] ), .ZN(n3640) );
  INV_X4 U1404 ( .A(n3642), .ZN(n3423) );
  OAI221_X2 U1405 ( .B1(n4594), .B2(n3643), .C1(n3644), .C2(n4590), .A(n4588), 
        .ZN(n3642) );
  INV_X4 U1406 ( .A(\u4/fract_out_pl1[41] ), .ZN(n3643) );
  INV_X4 U1408 ( .A(n3645), .ZN(n3424) );
  OAI221_X2 U1409 ( .B1(n4594), .B2(n3646), .C1(n2525), .C2(n4590), .A(n4588), 
        .ZN(n3645) );
  INV_X4 U1410 ( .A(\u4/fract_out_pl1[40] ), .ZN(n3646) );
  INV_X4 U1412 ( .A(n3647), .ZN(n3425) );
  OAI221_X2 U1413 ( .B1(n4594), .B2(n3648), .C1(n2527), .C2(n4590), .A(n4588), 
        .ZN(n3647) );
  INV_X4 U1414 ( .A(\u4/fract_out_pl1[39] ), .ZN(n3648) );
  INV_X4 U1416 ( .A(n3412), .ZN(n3602) );
  OAI221_X2 U1417 ( .B1(n4594), .B2(n3649), .C1(n3650), .C2(n4590), .A(n4588), 
        .ZN(n3412) );
  INV_X4 U1418 ( .A(\u4/fract_out_pl1[38] ), .ZN(n3649) );
  INV_X4 U1420 ( .A(n3414), .ZN(n3603) );
  OAI221_X2 U1421 ( .B1(n4594), .B2(n3651), .C1(n3652), .C2(n4590), .A(n4588), 
        .ZN(n3414) );
  INV_X4 U1422 ( .A(\u4/fract_out_pl1[37] ), .ZN(n3651) );
  INV_X4 U1424 ( .A(n3413), .ZN(n3604) );
  OAI221_X2 U1425 ( .B1(n4594), .B2(n3653), .C1(n3654), .C2(n4590), .A(n4588), 
        .ZN(n3413) );
  INV_X4 U1426 ( .A(\u4/fract_out_pl1[36] ), .ZN(n3653) );
  INV_X4 U1428 ( .A(n3655), .ZN(n3417) );
  OAI221_X2 U1429 ( .B1(n4594), .B2(n3656), .C1(n2528), .C2(n4590), .A(n4588), 
        .ZN(n3655) );
  INV_X4 U1430 ( .A(\u4/fract_out_pl1[35] ), .ZN(n3656) );
  INV_X4 U1432 ( .A(n3657), .ZN(n3415) );
  OAI221_X2 U1433 ( .B1(n4594), .B2(n3658), .C1(n2529), .C2(n4590), .A(n4588), 
        .ZN(n3657) );
  INV_X4 U1434 ( .A(\u4/fract_out_pl1[34] ), .ZN(n3658) );
  INV_X4 U1436 ( .A(n3659), .ZN(n3416) );
  OAI221_X2 U1437 ( .B1(n4594), .B2(n3660), .C1(n2530), .C2(n4590), .A(n4588), 
        .ZN(n3659) );
  INV_X4 U1438 ( .A(\u4/fract_out_pl1[33] ), .ZN(n3660) );
  INV_X4 U1440 ( .A(n3404), .ZN(n3605) );
  OAI221_X2 U1441 ( .B1(n4593), .B2(n3661), .C1(n3662), .C2(n4589), .A(n4587), 
        .ZN(n3404) );
  INV_X4 U1442 ( .A(\u4/fract_out_pl1[32] ), .ZN(n3661) );
  INV_X4 U1444 ( .A(n3406), .ZN(n3606) );
  OAI221_X2 U1445 ( .B1(n4593), .B2(n3663), .C1(n3664), .C2(n4589), .A(n4587), 
        .ZN(n3406) );
  INV_X4 U1446 ( .A(\u4/fract_out_pl1[31] ), .ZN(n3663) );
  INV_X4 U1448 ( .A(n3405), .ZN(n3607) );
  OAI221_X2 U1449 ( .B1(n4593), .B2(n3665), .C1(n3666), .C2(n4589), .A(n4587), 
        .ZN(n3405) );
  INV_X4 U1450 ( .A(\u4/fract_out_pl1[30] ), .ZN(n3665) );
  INV_X4 U1452 ( .A(n3667), .ZN(n3407) );
  OAI221_X2 U1453 ( .B1(n4593), .B2(n3668), .C1(n2531), .C2(n4589), .A(n4587), 
        .ZN(n3667) );
  INV_X4 U1454 ( .A(\u4/fract_out_pl1[29] ), .ZN(n3668) );
  INV_X4 U1456 ( .A(n3669), .ZN(n3408) );
  OAI221_X2 U1457 ( .B1(n4593), .B2(n3670), .C1(n2532), .C2(n4589), .A(n4587), 
        .ZN(n3669) );
  INV_X4 U1458 ( .A(\u4/fract_out_pl1[28] ), .ZN(n3670) );
  INV_X4 U1460 ( .A(n3671), .ZN(n3409) );
  OAI221_X2 U1461 ( .B1(n4593), .B2(n3672), .C1(n2533), .C2(n4589), .A(n4587), 
        .ZN(n3671) );
  INV_X4 U1462 ( .A(\u4/fract_out_pl1[27] ), .ZN(n3672) );
  INV_X4 U1464 ( .A(n3673), .ZN(n3410) );
  OAI221_X2 U1465 ( .B1(n4593), .B2(n3674), .C1(n3675), .C2(n4589), .A(n4587), 
        .ZN(n3673) );
  INV_X4 U1466 ( .A(\u4/fract_out_pl1[26] ), .ZN(n3674) );
  INV_X4 U1468 ( .A(n3448), .ZN(n3590) );
  OAI221_X2 U1469 ( .B1(n4593), .B2(n3676), .C1(n3677), .C2(n4589), .A(n4587), 
        .ZN(n3448) );
  INV_X4 U1470 ( .A(\u4/fract_out_pl1[25] ), .ZN(n3676) );
  INV_X4 U1472 ( .A(n3450), .ZN(n3591) );
  OAI221_X2 U1473 ( .B1(n4593), .B2(n3678), .C1(n3679), .C2(n4589), .A(n4587), 
        .ZN(n3450) );
  INV_X4 U1474 ( .A(\u4/fract_out_pl1[24] ), .ZN(n3678) );
  INV_X4 U1476 ( .A(n3449), .ZN(n3592) );
  OAI221_X2 U1477 ( .B1(n4593), .B2(n3680), .C1(n2534), .C2(n4589), .A(n4587), 
        .ZN(n3449) );
  INV_X4 U1478 ( .A(\u4/fract_out_pl1[23] ), .ZN(n3680) );
  INV_X4 U1480 ( .A(n3681), .ZN(n3453) );
  OAI221_X2 U1481 ( .B1(n4593), .B2(n3682), .C1(n2535), .C2(n4589), .A(n4587), 
        .ZN(n3681) );
  INV_X4 U1482 ( .A(\u4/fract_out_pl1[22] ), .ZN(n3682) );
  INV_X4 U1484 ( .A(n3683), .ZN(n3451) );
  OAI221_X2 U1485 ( .B1(n4594), .B2(n3684), .C1(n2536), .C2(n4591), .A(n4586), 
        .ZN(n3683) );
  INV_X4 U1486 ( .A(\u4/fract_out_pl1[21] ), .ZN(n3684) );
  INV_X4 U1488 ( .A(n3685), .ZN(n3452) );
  OAI221_X2 U1489 ( .B1(n4592), .B2(n3686), .C1(n3687), .C2(n4591), .A(n4586), 
        .ZN(n3685) );
  INV_X4 U1490 ( .A(\u4/fract_out_pl1[20] ), .ZN(n3686) );
  INV_X4 U1492 ( .A(n3440), .ZN(n3593) );
  OAI221_X2 U1493 ( .B1(n4592), .B2(n3688), .C1(n3689), .C2(n4591), .A(n4586), 
        .ZN(n3440) );
  INV_X4 U1494 ( .A(\u4/fract_out_pl1[19] ), .ZN(n3688) );
  INV_X4 U1496 ( .A(n3442), .ZN(n3594) );
  OAI221_X2 U1497 ( .B1(n4594), .B2(n3690), .C1(n3691), .C2(n4591), .A(n4586), 
        .ZN(n3442) );
  INV_X4 U1498 ( .A(\u4/fract_out_pl1[18] ), .ZN(n3690) );
  INV_X4 U1500 ( .A(n3441), .ZN(n3595) );
  OAI221_X2 U1501 ( .B1(n4592), .B2(n3692), .C1(n2537), .C2(n4589), .A(n4586), 
        .ZN(n3441) );
  INV_X4 U1502 ( .A(\u4/fract_out_pl1[17] ), .ZN(n3692) );
  INV_X4 U1504 ( .A(n3693), .ZN(n3443) );
  OAI221_X2 U1505 ( .B1(n4592), .B2(n3694), .C1(n2538), .C2(n4589), .A(n4586), 
        .ZN(n3693) );
  INV_X4 U1506 ( .A(\u4/fract_out_pl1[16] ), .ZN(n3694) );
  INV_X4 U1508 ( .A(n3695), .ZN(n3444) );
  OAI221_X2 U1509 ( .B1(n4592), .B2(n3696), .C1(n2539), .C2(n4589), .A(n4586), 
        .ZN(n3695) );
  INV_X4 U1510 ( .A(\u4/fract_out_pl1[15] ), .ZN(n3696) );
  INV_X4 U1512 ( .A(n3697), .ZN(n3445) );
  OAI221_X2 U1513 ( .B1(n4594), .B2(n3698), .C1(n3699), .C2(n4591), .A(n4586), 
        .ZN(n3697) );
  INV_X4 U1514 ( .A(\u4/fract_out_pl1[14] ), .ZN(n3698) );
  INV_X4 U1516 ( .A(n3700), .ZN(n3446) );
  OAI221_X2 U1517 ( .B1(n4594), .B2(n3701), .C1(n3702), .C2(n4591), .A(n4586), 
        .ZN(n3700) );
  INV_X4 U1518 ( .A(\u4/fract_out_pl1[13] ), .ZN(n3701) );
  INV_X4 U1520 ( .A(n3334), .ZN(n3578) );
  OAI221_X2 U1521 ( .B1(n4594), .B2(n3703), .C1(n3704), .C2(n4591), .A(n4586), 
        .ZN(n3334) );
  INV_X4 U1522 ( .A(\u4/fract_out_pl1[12] ), .ZN(n3703) );
  INV_X4 U1524 ( .A(n3336), .ZN(n3579) );
  OAI221_X2 U1525 ( .B1(n4594), .B2(n3705), .C1(n2540), .C2(n4591), .A(n4586), 
        .ZN(n3336) );
  INV_X4 U1526 ( .A(\u4/fract_out_pl1[11] ), .ZN(n3705) );
  INV_X4 U1528 ( .A(n3335), .ZN(n3580) );
  OAI221_X2 U1529 ( .B1(n4592), .B2(n3706), .C1(n2541), .C2(n4590), .A(n4586), 
        .ZN(n3335) );
  INV_X4 U1530 ( .A(\u4/fract_out_pl1[10] ), .ZN(n3706) );
  INV_X4 U1532 ( .A(n3707), .ZN(n3337) );
  OAI221_X2 U1533 ( .B1(n4592), .B2(n3708), .C1(n3709), .C2(n4591), .A(n4586), 
        .ZN(n3707) );
  INV_X4 U1534 ( .A(\u4/fract_out_pl1[9] ), .ZN(n3708) );
  INV_X4 U1536 ( .A(n3710), .ZN(n3338) );
  OAI221_X2 U1537 ( .B1(n4592), .B2(n3711), .C1(n3712), .C2(n4589), .A(n4586), 
        .ZN(n3710) );
  INV_X4 U1538 ( .A(\u4/fract_out_pl1[8] ), .ZN(n3711) );
  INV_X4 U1540 ( .A(n3713), .ZN(n3339) );
  OAI221_X2 U1541 ( .B1(n4592), .B2(n3714), .C1(n3715), .C2(n4591), .A(n4586), 
        .ZN(n3713) );
  INV_X4 U1542 ( .A(\u4/fract_out_pl1[7] ), .ZN(n3714) );
  INV_X4 U1544 ( .A(n3436), .ZN(n3340) );
  OAI221_X2 U1545 ( .B1(n4592), .B2(n3716), .C1(n3717), .C2(n4590), .A(n4586), 
        .ZN(n3436) );
  INV_X4 U1546 ( .A(\u4/fract_out_pl1[6] ), .ZN(n3716) );
  INV_X4 U1548 ( .A(n3326), .ZN(n3581) );
  OAI221_X2 U1549 ( .B1(n4592), .B2(n3718), .C1(n2519), .C2(n4590), .A(n4586), 
        .ZN(n3326) );
  INV_X4 U1550 ( .A(\u4/fract_out_pl1[5] ), .ZN(n3718) );
  INV_X4 U1552 ( .A(n3328), .ZN(n3582) );
  OAI221_X2 U1553 ( .B1(n4592), .B2(n3719), .C1(n3720), .C2(n4590), .A(n4586), 
        .ZN(n3328) );
  INV_X4 U1554 ( .A(\u4/fract_out_pl1[4] ), .ZN(n3719) );
  INV_X4 U1556 ( .A(n3327), .ZN(n3437) );
  OAI221_X2 U1557 ( .B1(n4592), .B2(n3721), .C1(n2526), .C2(n4590), .A(n4586), 
        .ZN(n3327) );
  INV_X4 U1558 ( .A(\u4/fract_out_pl1[3] ), .ZN(n3721) );
  INV_X4 U1560 ( .A(n3722), .ZN(n3329) );
  OAI221_X2 U1561 ( .B1(n4592), .B2(n3723), .C1(n3724), .C2(n4589), .A(n4586), 
        .ZN(n3722) );
  INV_X4 U1562 ( .A(\u4/fract_out_pl1[2] ), .ZN(n3723) );
  INV_X4 U1564 ( .A(n3725), .ZN(n3330) );
  OAI221_X2 U1565 ( .B1(n4592), .B2(n3726), .C1(n3727), .C2(n4590), .A(n4586), 
        .ZN(n3725) );
  INV_X4 U1566 ( .A(\u4/fract_out_pl1[1] ), .ZN(n3726) );
  OAI22_X2 U1567 ( .A1(n6310), .A2(n3331), .B1(n3341), .B2(n3619), .ZN(N793)
         );
  OAI22_X2 U1569 ( .A1(n3308), .A2(n4355), .B1(n2507), .B2(n3468), .ZN(n3728)
         );
  AOI22_X2 U1570 ( .A1(opb_00), .A2(opa_inf), .B1(opb_inf), .B2(opa_00), .ZN(
        n3468) );
  NAND2_X2 U1571 ( .A1(opa_00), .A2(opb_00), .ZN(n3308) );
  INV_X4 U1572 ( .A(n3729), .ZN(n3331) );
  OAI221_X2 U1573 ( .B1(n4592), .B2(n3730), .C1(n3731), .C2(n4590), .A(n4586), 
        .ZN(n3729) );
  OAI221_X2 U1580 ( .B1(n4351), .B2(n3739), .C1(\u4/N6410 ), .C2(n3740), .A(
        n3741), .ZN(n3738) );
  INV_X4 U1581 ( .A(\u4/fract_out_pl1[0] ), .ZN(n3730) );
  OAI22_X2 U1583 ( .A1(\u4/N6410 ), .A2(n3743), .B1(n3744), .B2(n4351), .ZN(
        n3742) );
  INV_X4 U1584 ( .A(n3739), .ZN(n3744) );
  AND3_X2 U1585 ( .A1(n3745), .A2(n3552), .A3(n3554), .ZN(n3734) );
  AND4_X2 U1587 ( .A1(n3584), .A2(n3583), .A3(n3746), .A4(n3747), .ZN(n3332)
         );
  NOR4_X2 U1588 ( .A1(n3748), .A2(n3389), .A3(n3617), .A4(n3388), .ZN(n3747)
         );
  INV_X4 U1593 ( .A(n3615), .ZN(n3393) );
  INV_X4 U1595 ( .A(n3539), .ZN(n3395) );
  INV_X4 U1597 ( .A(n3540), .ZN(n3394) );
  INV_X4 U1600 ( .A(n3534), .ZN(n3398) );
  INV_X4 U1604 ( .A(n3585), .ZN(n3618) );
  NAND2_X2 U1608 ( .A1(n6315), .A2(n3765), .ZN(n3758) );
  NAND2_X2 U1609 ( .A1(n3761), .A2(n6315), .ZN(n3757) );
  NAND2_X2 U1610 ( .A1(n3745), .A2(n3766), .ZN(n3760) );
  OAI211_X2 U1614 ( .C1(n3769), .C2(n3556), .A(\u4/N6410 ), .B(n3297), .ZN(
        n3768) );
  AND4_X2 U1615 ( .A1(n3770), .A2(n6466), .A3(\u4/N6249 ), .A4(n3771), .ZN(
        n3769) );
  OR4_X2 U1616 ( .A1(\u4/exp_out[0] ), .A2(\u4/exp_out[8] ), .A3(
        \u4/exp_out[9] ), .A4(n3772), .ZN(n3770) );
  AND4_X2 U1618 ( .A1(sign), .A2(rmode_r3[1]), .A3(n3775), .A4(n4452), .ZN(
        n3774) );
  OAI221_X2 U1619 ( .B1(n3776), .B2(n2514), .C1(n3777), .C2(n4653), .A(n3778), 
        .ZN(n3775) );
  NAND4_X2 U1620 ( .A1(n3762), .A2(n4656), .A3(n3779), .A4(n3780), .ZN(n3778)
         );
  OR4_X2 U1621 ( .A1(n3772), .A2(n2450), .A3(n2443), .A4(\u4/exp_out_mi1 [0]), 
        .ZN(n3779) );
  INV_X4 U1623 ( .A(\u4/exp_out[9] ), .ZN(n2443) );
  NAND2_X2 U1624 ( .A1(n3781), .A2(n3782), .ZN(n3772) );
  NOR4_X2 U1625 ( .A1(\u4/exp_out[10] ), .A2(n2453), .A3(n2456), .A4(n2459), 
        .ZN(n3782) );
  NOR4_X2 U1626 ( .A1(n2462), .A2(n2465), .A3(n2468), .A4(n2471), .ZN(n3781)
         );
  OAI211_X2 U1630 ( .C1(n4355), .C2(n3481), .A(n6306), .B(n3554), .ZN(n3765)
         );
  INV_X4 U1631 ( .A(n3478), .ZN(n3554) );
  AOI22_X2 U1632 ( .A1(n4540), .A2(n3785), .B1(n3786), .B2(n3297), .ZN(n3784)
         );
  NAND4_X2 U1636 ( .A1(\u4/N6249 ), .A2(n6466), .A3(n3791), .A4(n3488), .ZN(
        n3790) );
  NAND4_X2 U1637 ( .A1(n3762), .A2(n3763), .A3(n3792), .A4(n3793), .ZN(n3791)
         );
  AND4_X2 U1638 ( .A1(n3794), .A2(n3752), .A3(n3751), .A4(n3749), .ZN(n3793)
         );
  OAI211_X2 U1639 ( .C1(n3795), .C2(n2465), .A(n3796), .B(n3797), .ZN(n3749)
         );
  AOI221_X2 U1640 ( .B1(\u4/exp_fix_divb [3]), .B2(n3798), .C1(
        \u4/exp_fix_diva [3]), .C2(n3799), .A(n3800), .ZN(n3797) );
  INV_X4 U1641 ( .A(n3801), .ZN(n3800) );
  AOI22_X2 U1642 ( .A1(\u4/exp_next_mi[3] ), .A2(n3802), .B1(exp_r[3]), .B2(
        n3803), .ZN(n3801) );
  AOI22_X2 U1643 ( .A1(\u4/exp_out_mi1 [3]), .A2(n3804), .B1(
        \u4/exp_out_pl1[3] ), .B2(n3805), .ZN(n3796) );
  OAI211_X2 U1644 ( .C1(n3795), .C2(n2462), .A(n3806), .B(n3807), .ZN(n3751)
         );
  AOI221_X2 U1645 ( .B1(\u4/exp_fix_divb [4]), .B2(n3798), .C1(
        \u4/exp_fix_diva [4]), .C2(n3799), .A(n3808), .ZN(n3807) );
  INV_X4 U1646 ( .A(n3809), .ZN(n3808) );
  AOI22_X2 U1647 ( .A1(\u4/exp_next_mi[4] ), .A2(n3802), .B1(n4282), .B2(n3803), .ZN(n3809) );
  AOI22_X2 U1648 ( .A1(\u4/exp_out_mi1 [4]), .A2(n3804), .B1(
        \u4/exp_out_pl1[4] ), .B2(n3805), .ZN(n3806) );
  OAI211_X2 U1649 ( .C1(n3795), .C2(n2468), .A(n3810), .B(n3811), .ZN(n3752)
         );
  AOI221_X2 U1650 ( .B1(\u4/exp_fix_divb [2]), .B2(n3798), .C1(
        \u4/exp_fix_diva [2]), .C2(n3799), .A(n3812), .ZN(n3811) );
  INV_X4 U1651 ( .A(n3813), .ZN(n3812) );
  AOI22_X2 U1652 ( .A1(\u4/exp_next_mi[2] ), .A2(n3802), .B1(n4315), .B2(n3803), .ZN(n3813) );
  AOI22_X2 U1653 ( .A1(\u4/exp_out_mi1 [2]), .A2(n3804), .B1(
        \u4/exp_out_pl1[2] ), .B2(n3805), .ZN(n3810) );
  INV_X4 U1654 ( .A(\u4/exp_out[2] ), .ZN(n2468) );
  AND3_X2 U1655 ( .A1(n3755), .A2(n3754), .A3(n3753), .ZN(n3794) );
  OAI211_X2 U1656 ( .C1(n3795), .C2(n2459), .A(n3814), .B(n3815), .ZN(n3753)
         );
  AOI221_X2 U1657 ( .B1(\u4/exp_fix_divb [5]), .B2(n3798), .C1(
        \u4/exp_fix_diva [5]), .C2(n3799), .A(n3816), .ZN(n3815) );
  INV_X4 U1658 ( .A(n3817), .ZN(n3816) );
  AOI22_X2 U1659 ( .A1(\u4/exp_next_mi[5] ), .A2(n3802), .B1(n4290), .B2(n3803), .ZN(n3817) );
  AOI22_X2 U1660 ( .A1(\u4/exp_out_mi1 [5]), .A2(n3804), .B1(
        \u4/exp_out_pl1[5] ), .B2(n3805), .ZN(n3814) );
  OAI211_X2 U1661 ( .C1(n3795), .C2(n2453), .A(n3818), .B(n3819), .ZN(n3754)
         );
  AOI221_X2 U1662 ( .B1(\u4/exp_fix_divb [7]), .B2(n3798), .C1(
        \u4/exp_fix_diva [7]), .C2(n3799), .A(n3820), .ZN(n3819) );
  INV_X4 U1663 ( .A(n3821), .ZN(n3820) );
  AOI22_X2 U1664 ( .A1(\u4/exp_next_mi[7] ), .A2(n3802), .B1(n4281), .B2(n3803), .ZN(n3821) );
  AOI22_X2 U1665 ( .A1(\u4/exp_out_mi1 [7]), .A2(n3804), .B1(
        \u4/exp_out_pl1[7] ), .B2(n3805), .ZN(n3818) );
  OAI211_X2 U1666 ( .C1(n3795), .C2(n2456), .A(n3822), .B(n3823), .ZN(n3755)
         );
  AOI221_X2 U1667 ( .B1(\u4/exp_fix_divb [6]), .B2(n3798), .C1(
        \u4/exp_fix_diva [6]), .C2(n3799), .A(n3824), .ZN(n3823) );
  INV_X4 U1668 ( .A(n3825), .ZN(n3824) );
  AOI22_X2 U1669 ( .A1(\u4/exp_next_mi[6] ), .A2(n3802), .B1(exp_r[6]), .B2(
        n3803), .ZN(n3825) );
  AOI22_X2 U1670 ( .A1(\u4/exp_out_mi1 [6]), .A2(n3804), .B1(
        \u4/exp_out_pl1[6] ), .B2(n3805), .ZN(n3822) );
  AND3_X2 U1671 ( .A1(n3764), .A2(n3759), .A3(n3756), .ZN(n3792) );
  AND3_X2 U1672 ( .A1(n3826), .A2(n3827), .A3(n3828), .ZN(n3756) );
  AOI22_X2 U1674 ( .A1(\u4/exp_fix_divb [0]), .A2(n3798), .B1(
        \u4/exp_fix_diva [0]), .B2(n3799), .ZN(n3827) );
  AOI22_X2 U1675 ( .A1(\u4/exp_out_mi1 [0]), .A2(n3804), .B1(n3803), .B2(n4600), .ZN(n3826) );
  OAI211_X2 U1676 ( .C1(n3795), .C2(n2471), .A(n3830), .B(n3831), .ZN(n3759)
         );
  AOI221_X2 U1677 ( .B1(\u4/exp_fix_divb [1]), .B2(n3798), .C1(
        \u4/exp_fix_diva [1]), .C2(n3799), .A(n3832), .ZN(n3831) );
  INV_X4 U1678 ( .A(n3833), .ZN(n3832) );
  AOI22_X2 U1679 ( .A1(\u4/exp_next_mi[1] ), .A2(n3802), .B1(exp_r[1]), .B2(
        n3803), .ZN(n3833) );
  AOI22_X2 U1680 ( .A1(\u4/exp_out_mi1 [1]), .A2(n3804), .B1(
        \u4/exp_out_pl1[1] ), .B2(n3805), .ZN(n3830) );
  INV_X4 U1681 ( .A(\u4/exp_out[1] ), .ZN(n2471) );
  INV_X4 U1683 ( .A(n3836), .ZN(n3835) );
  AND3_X2 U1684 ( .A1(n3837), .A2(n3838), .A3(n3839), .ZN(n3763) );
  AOI22_X2 U1686 ( .A1(\u4/exp_fix_divb [9]), .A2(n3798), .B1(
        \u4/exp_fix_diva [9]), .B2(n3799), .ZN(n3838) );
  AOI22_X2 U1687 ( .A1(\u4/exp_out_mi1 [9]), .A2(n3804), .B1(n3803), .B2(n4289), .ZN(n3837) );
  AND3_X2 U1688 ( .A1(n3840), .A2(n3841), .A3(n3842), .ZN(n3762) );
  AOI22_X2 U1690 ( .A1(\u4/exp_fix_divb [10]), .A2(n3798), .B1(
        \u4/exp_fix_diva [10]), .B2(n3799), .ZN(n3841) );
  AOI22_X2 U1691 ( .A1(\u4/exp_out_mi1 [10]), .A2(n3804), .B1(n3803), .B2(
        n4656), .ZN(n3840) );
  OAI22_X2 U1695 ( .A1(opas_r2), .A2(n6467), .B1(n6308), .B2(n3843), .ZN(n2435) );
  NAND2_X2 U1696 ( .A1(n3556), .A2(n4823), .ZN(n3481) );
  AND3_X2 U1698 ( .A1(n3844), .A2(n3845), .A3(n3846), .ZN(n3764) );
  INV_X4 U1701 ( .A(n3848), .ZN(n2440) );
  NAND2_X2 U1703 ( .A1(n3836), .A2(n3850), .ZN(n3829) );
  AOI22_X2 U1706 ( .A1(n4823), .A2(n3847), .B1(n6305), .B2(n3852), .ZN(n3836)
         );
  INV_X4 U1708 ( .A(n3551), .ZN(n3557) );
  NAND2_X2 U1709 ( .A1(n3740), .A2(\u4/fract_out_pl1[52] ), .ZN(n3847) );
  INV_X4 U1710 ( .A(n3743), .ZN(n3740) );
  AOI22_X2 U1712 ( .A1(\u4/exp_fix_divb [8]), .A2(n3798), .B1(
        \u4/exp_fix_diva [8]), .B2(n3799), .ZN(n3845) );
  AOI22_X2 U1716 ( .A1(\u4/exp_out_mi1 [8]), .A2(n3804), .B1(n3803), .B2(n4353), .ZN(n3844) );
  NAND4_X2 U1718 ( .A1(\u4/exp_out[1] ), .A2(\u4/exp_out[2] ), .A3(n3856), 
        .A4(n3857), .ZN(n3551) );
  NOR4_X2 U1719 ( .A1(n3858), .A2(n2456), .A3(n2450), .A4(n2453), .ZN(n3857)
         );
  INV_X4 U1720 ( .A(\u4/exp_out[7] ), .ZN(n2453) );
  INV_X4 U1721 ( .A(\u4/exp_out[8] ), .ZN(n2450) );
  INV_X4 U1722 ( .A(\u4/exp_out[6] ), .ZN(n2456) );
  INV_X4 U1725 ( .A(\u4/exp_out[4] ), .ZN(n2462) );
  INV_X4 U1726 ( .A(\u4/exp_out[5] ), .ZN(n2459) );
  INV_X4 U1727 ( .A(\u4/exp_out[3] ), .ZN(n2465) );
  AND4_X2 U1728 ( .A1(n3854), .A2(n6466), .A3(\u4/fract_out[0] ), .A4(n3853), 
        .ZN(n3849) );
  INV_X4 U1729 ( .A(n3731), .ZN(\u4/fract_out[0] ) );
  NAND4_X2 U1730 ( .A1(n4289), .A2(n4600), .A3(n3859), .A4(n3860), .ZN(n3787)
         );
  NOR4_X2 U1731 ( .A1(n3861), .A2(n4299), .A3(n4317), .A4(n4347), .ZN(n3860)
         );
  AND3_X2 U1733 ( .A1(exp_r[1]), .A2(n4655), .A3(n4315), .ZN(n3859) );
  NAND2_X2 U1736 ( .A1(\u4/fract_out_pl1[52] ), .A2(n3739), .ZN(n3834) );
  OAI211_X2 U1738 ( .C1(n3864), .C2(n3485), .A(n4441), .B(n6342), .ZN(n3863)
         );
  NAND2_X2 U1739 ( .A1(n3865), .A2(n3866), .ZN(n3485) );
  NAND4_X2 U1744 ( .A1(n6404), .A2(n6403), .A3(n2763), .A4(n3872), .ZN(n3869)
         );
  NOR4_X2 U1746 ( .A1(n3874), .A2(n3875), .A3(n2634), .A4(n2771), .ZN(n3867)
         );
  OR3_X2 U1747 ( .A1(n2635), .A2(n2561), .A3(n2604), .ZN(n3875) );
  NAND4_X2 U1748 ( .A1(n3876), .A2(n2636), .A3(n3877), .A4(n3878), .ZN(n3874)
         );
  AND4_X2 U1751 ( .A1(\u4/N6917 ), .A2(n6317), .A3(n3544), .A4(n2434), .ZN(
        n3881) );
  OAI211_X2 U1754 ( .C1(n4540), .C2(n3488), .A(n3473), .B(n3882), .ZN(n3885)
         );
  NAND2_X2 U1755 ( .A1(n3886), .A2(n3887), .ZN(n3473) );
  NOR4_X2 U1756 ( .A1(n3888), .A2(n3889), .A3(n3890), .A4(n3891), .ZN(n3887)
         );
  NAND4_X2 U1757 ( .A1(n2529), .A2(n2528), .A3(n2530), .A4(n3892), .ZN(n3891)
         );
  INV_X4 U1759 ( .A(n3652), .ZN(\u4/fract_out[37] ) );
  AOI22_X2 U1760 ( .A1(\u4/N5997 ), .A2(n4578), .B1(\u4/N6105 ), .B2(n4576), 
        .ZN(n3652) );
  INV_X4 U1761 ( .A(n3650), .ZN(\u4/fract_out[38] ) );
  AOI22_X2 U1762 ( .A1(\u4/N5998 ), .A2(n4582), .B1(\u4/N6106 ), .B2(n4577), 
        .ZN(n3650) );
  INV_X4 U1763 ( .A(n3654), .ZN(\u4/fract_out[36] ) );
  AOI22_X2 U1764 ( .A1(\u4/N5996 ), .A2(n4582), .B1(\u4/N6104 ), .B2(n4577), 
        .ZN(n3654) );
  AOI22_X2 U1765 ( .A1(\u4/N5993 ), .A2(n4582), .B1(\u4/N6101 ), .B2(n4577), 
        .ZN(n2530) );
  AOI22_X2 U1766 ( .A1(\u4/N5995 ), .A2(n4582), .B1(\u4/N6103 ), .B2(n4577), 
        .ZN(n2528) );
  AOI22_X2 U1767 ( .A1(\u4/N5994 ), .A2(n4582), .B1(\u4/N6102 ), .B2(n4577), 
        .ZN(n2529) );
  NAND4_X2 U1768 ( .A1(n2526), .A2(n2525), .A3(n2527), .A4(n3895), .ZN(n3890)
         );
  NOR4_X2 U1769 ( .A1(\u4/fract_out[44] ), .A2(\u4/fract_out[43] ), .A3(
        \u4/fract_out[42] ), .A4(\u4/fract_out[41] ), .ZN(n3895) );
  INV_X4 U1770 ( .A(n3644), .ZN(\u4/fract_out[41] ) );
  AOI22_X2 U1771 ( .A1(\u4/N6001 ), .A2(n4582), .B1(\u4/N6109 ), .B2(n4577), 
        .ZN(n3644) );
  INV_X4 U1772 ( .A(n3641), .ZN(\u4/fract_out[42] ) );
  AOI22_X2 U1773 ( .A1(\u4/N6002 ), .A2(n4582), .B1(\u4/N6110 ), .B2(n4577), 
        .ZN(n3641) );
  INV_X4 U1774 ( .A(n3638), .ZN(\u4/fract_out[43] ) );
  AOI22_X2 U1775 ( .A1(\u4/N6003 ), .A2(n4582), .B1(\u4/N6111 ), .B2(n4577), 
        .ZN(n3638) );
  INV_X4 U1776 ( .A(n3636), .ZN(\u4/fract_out[44] ) );
  AOI22_X2 U1777 ( .A1(\u4/N6004 ), .A2(n4582), .B1(\u4/N6112 ), .B2(n4577), 
        .ZN(n3636) );
  AOI22_X2 U1778 ( .A1(\u4/N5999 ), .A2(n4582), .B1(\u4/N6107 ), .B2(n4577), 
        .ZN(n2527) );
  AOI22_X2 U1779 ( .A1(\u4/N6000 ), .A2(n4581), .B1(\u4/N6108 ), .B2(n4577), 
        .ZN(n2525) );
  AOI22_X2 U1780 ( .A1(\u4/N5963 ), .A2(n4581), .B1(\u4/N6071 ), .B2(n4577), 
        .ZN(n2526) );
  NAND4_X2 U1781 ( .A1(n2523), .A2(n2522), .A3(n2524), .A4(n3896), .ZN(n3889)
         );
  INV_X4 U1783 ( .A(n3626), .ZN(\u4/fract_out[49] ) );
  AOI22_X2 U1784 ( .A1(\u4/N6009 ), .A2(n4581), .B1(\u4/N6117 ), .B2(n4577), 
        .ZN(n3626) );
  INV_X4 U1785 ( .A(n3720), .ZN(\u4/fract_out[4] ) );
  AOI22_X2 U1786 ( .A1(\u4/N5964 ), .A2(n4581), .B1(\u4/N6072 ), .B2(n4577), 
        .ZN(n3720) );
  INV_X4 U1787 ( .A(n3629), .ZN(\u4/fract_out[48] ) );
  AOI22_X2 U1788 ( .A1(\u4/N6008 ), .A2(n4581), .B1(\u4/N6116 ), .B2(n4577), 
        .ZN(n3629) );
  AOI22_X2 U1789 ( .A1(\u4/N6005 ), .A2(n4581), .B1(\u4/N6113 ), .B2(n4577), 
        .ZN(n2524) );
  AOI22_X2 U1790 ( .A1(\u4/N6007 ), .A2(n4581), .B1(\u4/N6115 ), .B2(n4577), 
        .ZN(n2522) );
  AOI22_X2 U1791 ( .A1(\u4/N6006 ), .A2(n4581), .B1(\u4/N6114 ), .B2(n4577), 
        .ZN(n2523) );
  NAND4_X2 U1792 ( .A1(n2520), .A2(n2519), .A3(n2521), .A4(n3897), .ZN(n3888)
         );
  NOR4_X2 U1793 ( .A1(\u4/fract_out[9] ), .A2(\u4/fract_out[8] ), .A3(
        \u4/fract_out[7] ), .A4(\u4/fract_out[6] ), .ZN(n3897) );
  INV_X4 U1794 ( .A(n3717), .ZN(\u4/fract_out[6] ) );
  AOI22_X2 U1795 ( .A1(\u4/N5966 ), .A2(n4581), .B1(\u4/N6074 ), .B2(n4577), 
        .ZN(n3717) );
  INV_X4 U1796 ( .A(n3715), .ZN(\u4/fract_out[7] ) );
  AOI22_X2 U1797 ( .A1(\u4/N5967 ), .A2(n4581), .B1(\u4/N6075 ), .B2(n4577), 
        .ZN(n3715) );
  INV_X4 U1798 ( .A(n3712), .ZN(\u4/fract_out[8] ) );
  AOI22_X2 U1799 ( .A1(\u4/N5968 ), .A2(n4581), .B1(\u4/N6076 ), .B2(n3894), 
        .ZN(n3712) );
  INV_X4 U1800 ( .A(n3709), .ZN(\u4/fract_out[9] ) );
  AOI22_X2 U1801 ( .A1(\u4/N5969 ), .A2(n4580), .B1(\u4/N6077 ), .B2(n3894), 
        .ZN(n3709) );
  AOI22_X2 U1802 ( .A1(\u4/N6010 ), .A2(n4580), .B1(\u4/N6118 ), .B2(n3894), 
        .ZN(n2521) );
  AOI22_X2 U1803 ( .A1(\u4/N5965 ), .A2(n4580), .B1(\u4/N6073 ), .B2(n3894), 
        .ZN(n2519) );
  AOI22_X2 U1804 ( .A1(\u4/N6011 ), .A2(n4580), .B1(\u4/N6119 ), .B2(n3894), 
        .ZN(n2520) );
  NOR4_X2 U1805 ( .A1(n3898), .A2(n3899), .A3(n3900), .A4(n3901), .ZN(n3886)
         );
  NAND4_X2 U1806 ( .A1(n2541), .A2(n2540), .A3(n3731), .A4(n3902), .ZN(n3901)
         );
  INV_X4 U1808 ( .A(n3702), .ZN(\u4/fract_out[13] ) );
  AOI22_X2 U1809 ( .A1(\u4/N5973 ), .A2(n4580), .B1(\u4/N6081 ), .B2(n3894), 
        .ZN(n3702) );
  INV_X4 U1810 ( .A(n3699), .ZN(\u4/fract_out[14] ) );
  AOI22_X2 U1811 ( .A1(\u4/N5974 ), .A2(n4580), .B1(\u4/N6082 ), .B2(n3894), 
        .ZN(n3699) );
  INV_X4 U1812 ( .A(n3704), .ZN(\u4/fract_out[12] ) );
  AOI22_X2 U1813 ( .A1(\u4/N5972 ), .A2(n4580), .B1(\u4/N6080 ), .B2(n3894), 
        .ZN(n3704) );
  AOI22_X2 U1814 ( .A1(\u4/N5960 ), .A2(n4580), .B1(\u4/N6068 ), .B2(n3894), 
        .ZN(n3731) );
  AOI22_X2 U1815 ( .A1(\u4/N5971 ), .A2(n4580), .B1(\u4/N6079 ), .B2(n3894), 
        .ZN(n2540) );
  AOI22_X2 U1816 ( .A1(\u4/N5970 ), .A2(n4580), .B1(\u4/N6078 ), .B2(n4576), 
        .ZN(n2541) );
  NAND4_X2 U1817 ( .A1(n2538), .A2(n2537), .A3(n2539), .A4(n3903), .ZN(n3900)
         );
  NOR4_X2 U1818 ( .A1(\u4/fract_out[20] ), .A2(\u4/fract_out[1] ), .A3(
        \u4/fract_out[19] ), .A4(\u4/fract_out[18] ), .ZN(n3903) );
  INV_X4 U1819 ( .A(n3691), .ZN(\u4/fract_out[18] ) );
  AOI22_X2 U1820 ( .A1(\u4/N5978 ), .A2(n4579), .B1(\u4/N6086 ), .B2(n4576), 
        .ZN(n3691) );
  INV_X4 U1821 ( .A(n3689), .ZN(\u4/fract_out[19] ) );
  AOI22_X2 U1822 ( .A1(\u4/N5979 ), .A2(n4579), .B1(\u4/N6087 ), .B2(n4576), 
        .ZN(n3689) );
  INV_X4 U1823 ( .A(n3727), .ZN(\u4/fract_out[1] ) );
  AOI22_X2 U1824 ( .A1(\u4/N5961 ), .A2(n4579), .B1(\u4/N6069 ), .B2(n4576), 
        .ZN(n3727) );
  INV_X4 U1825 ( .A(n3687), .ZN(\u4/fract_out[20] ) );
  AOI22_X2 U1826 ( .A1(\u4/N5980 ), .A2(n4579), .B1(\u4/N6088 ), .B2(n4576), 
        .ZN(n3687) );
  AOI22_X2 U1827 ( .A1(\u4/N5975 ), .A2(n4579), .B1(\u4/N6083 ), .B2(n4576), 
        .ZN(n2539) );
  AOI22_X2 U1828 ( .A1(\u4/N5977 ), .A2(n4579), .B1(\u4/N6085 ), .B2(n4576), 
        .ZN(n2537) );
  AOI22_X2 U1829 ( .A1(\u4/N5976 ), .A2(n4579), .B1(\u4/N6084 ), .B2(n4576), 
        .ZN(n2538) );
  NAND4_X2 U1830 ( .A1(n2535), .A2(n2534), .A3(n2536), .A4(n3904), .ZN(n3899)
         );
  INV_X4 U1832 ( .A(n3677), .ZN(\u4/fract_out[25] ) );
  AOI22_X2 U1833 ( .A1(\u4/N5985 ), .A2(n4579), .B1(\u4/N6093 ), .B2(n4576), 
        .ZN(n3677) );
  INV_X4 U1834 ( .A(n3675), .ZN(\u4/fract_out[26] ) );
  AOI22_X2 U1835 ( .A1(\u4/N5986 ), .A2(n4579), .B1(\u4/N6094 ), .B2(n4576), 
        .ZN(n3675) );
  INV_X4 U1836 ( .A(n3679), .ZN(\u4/fract_out[24] ) );
  AOI22_X2 U1837 ( .A1(\u4/N5984 ), .A2(n4579), .B1(\u4/N6092 ), .B2(n4576), 
        .ZN(n3679) );
  AOI22_X2 U1838 ( .A1(\u4/N5981 ), .A2(n4579), .B1(\u4/N6089 ), .B2(n4577), 
        .ZN(n2536) );
  AOI22_X2 U1839 ( .A1(\u4/N5983 ), .A2(n4578), .B1(\u4/N6091 ), .B2(n4576), 
        .ZN(n2534) );
  AOI22_X2 U1840 ( .A1(\u4/N5982 ), .A2(n4578), .B1(\u4/N6090 ), .B2(n4576), 
        .ZN(n2535) );
  NAND4_X2 U1841 ( .A1(n2532), .A2(n2531), .A3(n2533), .A4(n3905), .ZN(n3898)
         );
  NOR4_X2 U1842 ( .A1(\u4/fract_out[32] ), .A2(\u4/fract_out[31] ), .A3(
        \u4/fract_out[30] ), .A4(\u4/fract_out[2] ), .ZN(n3905) );
  INV_X4 U1843 ( .A(n3724), .ZN(\u4/fract_out[2] ) );
  AOI22_X2 U1844 ( .A1(\u4/N5962 ), .A2(n4578), .B1(\u4/N6070 ), .B2(n4576), 
        .ZN(n3724) );
  INV_X4 U1845 ( .A(n3666), .ZN(\u4/fract_out[30] ) );
  AOI22_X2 U1846 ( .A1(\u4/N5990 ), .A2(n4578), .B1(\u4/N6098 ), .B2(n4576), 
        .ZN(n3666) );
  INV_X4 U1847 ( .A(n3664), .ZN(\u4/fract_out[31] ) );
  AOI22_X2 U1848 ( .A1(\u4/N5991 ), .A2(n4578), .B1(\u4/N6099 ), .B2(n4577), 
        .ZN(n3664) );
  INV_X4 U1849 ( .A(n3662), .ZN(\u4/fract_out[32] ) );
  AOI22_X2 U1850 ( .A1(\u4/N5992 ), .A2(n4578), .B1(\u4/N6100 ), .B2(n4576), 
        .ZN(n3662) );
  AOI22_X2 U1851 ( .A1(\u4/N5987 ), .A2(n4578), .B1(\u4/N6095 ), .B2(n4576), 
        .ZN(n2533) );
  AOI22_X2 U1852 ( .A1(\u4/N5989 ), .A2(n4578), .B1(\u4/N6097 ), .B2(n4576), 
        .ZN(n2531) );
  AOI22_X2 U1853 ( .A1(\u4/N5988 ), .A2(n4578), .B1(\u4/N6096 ), .B2(n4576), 
        .ZN(n2532) );
  OAI22_X2 U1856 ( .A1(exp_ovf_r[0]), .A2(n6095), .B1(exp_ovf_r[1]), .B2(n3780), .ZN(n3906) );
  NAND4_X2 U1857 ( .A1(n4656), .A2(n4349), .A3(n3907), .A4(n3908), .ZN(n3780)
         );
  NOR4_X2 U1858 ( .A1(n3909), .A2(n4282), .A3(exp_r[6]), .A4(n4290), .ZN(n3908) );
  OR3_X2 U1859 ( .A1(n4353), .A2(n4289), .A3(n4281), .ZN(n3909) );
  OR2_X2 U1862 ( .A1(n3853), .A2(n3854), .ZN(n3544) );
  AND4_X2 U1864 ( .A1(\u4/N5843 ), .A2(n6369), .A3(n6352), .A4(n2761), .ZN(
        n3911) );
  AND4_X2 U1865 ( .A1(n6365), .A2(n6360), .A3(n6359), .A4(n2449), .ZN(n3910)
         );
  AOI22_X2 U1868 ( .A1(n3914), .A2(n4577), .B1(n3915), .B2(n4578), .ZN(n3866)
         );
  OR4_X2 U1869 ( .A1(n3916), .A2(n3917), .A3(n3918), .A4(n3919), .ZN(n3915) );
  NAND4_X2 U1870 ( .A1(n3920), .A2(n3921), .A3(n3922), .A4(n3923), .ZN(n3919)
         );
  NOR4_X2 U1871 ( .A1(\u4/N5918 ), .A2(\u4/N5917 ), .A3(\u4/N5916 ), .A4(
        \u4/N5915 ), .ZN(n3923) );
  NAND4_X2 U1875 ( .A1(n3924), .A2(n3925), .A3(n3926), .A4(n3927), .ZN(n3918)
         );
  NOR4_X2 U1876 ( .A1(\u4/N5931 ), .A2(\u4/N5930 ), .A3(\u4/N5929 ), .A4(
        \u4/N5928 ), .ZN(n3927) );
  NAND4_X2 U1880 ( .A1(n3928), .A2(n3929), .A3(n3930), .A4(n3931), .ZN(n3917)
         );
  NOR4_X2 U1881 ( .A1(\u4/N5944 ), .A2(\u4/N5943 ), .A3(\u4/N5942 ), .A4(
        \u4/N5941 ), .ZN(n3931) );
  NAND4_X2 U1885 ( .A1(n3932), .A2(n3933), .A3(n3934), .A4(n3935), .ZN(n3916)
         );
  NOR4_X2 U1886 ( .A1(\u4/N5958 ), .A2(\u4/N5957 ), .A3(\u4/N5956 ), .A4(
        \u4/N5955 ), .ZN(n3935) );
  NOR4_X2 U1888 ( .A1(\u4/N5951 ), .A2(\u4/N5950 ), .A3(\u4/N5949 ), .A4(
        \u4/N5948 ), .ZN(n3933) );
  OR4_X2 U1890 ( .A1(n3936), .A2(n3937), .A3(n3938), .A4(n3939), .ZN(n3914) );
  NAND4_X2 U1891 ( .A1(n3940), .A2(n3941), .A3(n3942), .A4(n3943), .ZN(n3939)
         );
  NOR4_X2 U1892 ( .A1(\u4/N6026 ), .A2(\u4/N6025 ), .A3(\u4/N6024 ), .A4(
        \u4/N6023 ), .ZN(n3943) );
  NAND4_X2 U1896 ( .A1(n3944), .A2(n3945), .A3(n3946), .A4(n3947), .ZN(n3938)
         );
  NOR4_X2 U1897 ( .A1(\u4/N6039 ), .A2(\u4/N6038 ), .A3(\u4/N6037 ), .A4(
        \u4/N6036 ), .ZN(n3947) );
  NAND4_X2 U1901 ( .A1(n3948), .A2(n3949), .A3(n3950), .A4(n3951), .ZN(n3937)
         );
  NOR4_X2 U1902 ( .A1(\u4/N6052 ), .A2(\u4/N6051 ), .A3(\u4/N6050 ), .A4(
        \u4/N6049 ), .ZN(n3951) );
  NAND4_X2 U1906 ( .A1(n3952), .A2(n3953), .A3(n3954), .A4(n3955), .ZN(n3936)
         );
  NOR4_X2 U1907 ( .A1(\u4/N6066 ), .A2(\u4/N6065 ), .A3(\u4/N6064 ), .A4(
        \u4/N6063 ), .ZN(n3955) );
  NOR4_X2 U1909 ( .A1(\u4/N6059 ), .A2(\u4/N6058 ), .A3(\u4/N6057 ), .A4(
        \u4/N6056 ), .ZN(n3953) );
  AOI22_X2 U1911 ( .A1(\u4/N5959 ), .A2(n4580), .B1(\u4/N6067 ), .B2(n3894), 
        .ZN(n3865) );
  INV_X4 U1912 ( .A(n3956), .ZN(n3894) );
  OAI211_X2 U1913 ( .C1(n3957), .C2(n2434), .A(n3958), .B(n3959), .ZN(n3956)
         );
  OAI22_X2 U1915 ( .A1(n2506), .A2(n2507), .B1(n2508), .B2(n3962), .ZN(n2485)
         );
  NAND2_X2 U1916 ( .A1(n2511), .A2(n2514), .ZN(n3962) );
  NAND2_X2 U1917 ( .A1(\u4/N6463 ), .A2(n3545), .ZN(n2511) );
  NAND2_X2 U1918 ( .A1(n6317), .A2(n3963), .ZN(n3545) );
  NAND2_X2 U1922 ( .A1(n6095), .A2(\u4/N6463 ), .ZN(n3476) );
  NAND2_X2 U1924 ( .A1(\u4/exp_in_pl1[11] ), .A2(fract_denorm[105]), .ZN(n3964) );
  OR2_X2 U1925 ( .A1(\u4/exp_in_pl1[9] ), .A2(\u4/exp_in_pl1[10] ), .ZN(n3961)
         );
  OR2_X2 U1926 ( .A1(\u4/div_scht1a [10]), .A2(\u4/div_scht1a [9]), .ZN(n3960)
         );
  AOI22_X2 U1928 ( .A1(n3489), .A2(n6448), .B1(n4356), .B2(n3533), .ZN(n2515)
         );
  NOR2_X4 U1929 ( .A1(n6447), .A2(\u4/N6463 ), .ZN(n3533) );
  INV_X4 U1932 ( .A(\u4/N6463 ), .ZN(n3489) );
  AOI22_X2 U1934 ( .A1(opas_r2), .A2(\u4/N5837 ), .B1(n3843), .B2(\u4/N5836 ), 
        .ZN(n3548) );
  NAND4_X2 U1935 ( .A1(rmode_r3[1]), .A2(rmode_r3[0]), .A3(opas_r2), .A4(n6337), .ZN(n3843) );
  AOI221_X2 U1937 ( .B1(n4575), .B2(quo[2]), .C1(n4569), .C2(prod[0]), .A(
        n3967), .ZN(n3877) );
  AND2_X2 U1938 ( .A1(fract_i2f[0]), .A2(n4662), .ZN(n3967) );
  AND3_X2 U1940 ( .A1(n3873), .A2(n2763), .A3(n2700), .ZN(n2630) );
  AND3_X2 U1941 ( .A1(n3171), .A2(n2751), .A3(n2659), .ZN(n2700) );
  NAND4_X2 U1943 ( .A1(n3968), .A2(n3969), .A3(n3970), .A4(n3971), .ZN(n2684)
         );
  NOR4_X2 U1944 ( .A1(n6444), .A2(fract_denorm[51]), .A3(fract_denorm[50]), 
        .A4(n6445), .ZN(n3971) );
  AOI221_X2 U1945 ( .B1(n4571), .B2(quo[44]), .C1(n4569), .C2(prod[42]), .A(
        n3972), .ZN(n2770) );
  AND2_X2 U1946 ( .A1(fract_i2f[42]), .A2(n4662), .ZN(n3972) );
  OAI211_X2 U1947 ( .C1(n3973), .C2(n4434), .A(n3974), .B(n3975), .ZN(
        fract_denorm[50]) );
  AOI22_X2 U1948 ( .A1(fract_out_q[1]), .A2(n4595), .B1(fract_i2f[50]), .B2(
        n4661), .ZN(n3975) );
  AOI22_X2 U1949 ( .A1(quo[0]), .A2(n4563), .B1(quo[52]), .B2(n4572), .ZN(
        n3974) );
  OAI211_X2 U1950 ( .C1(n3973), .C2(n4432), .A(n3977), .B(n3978), .ZN(
        fract_denorm[51]) );
  AOI22_X2 U1951 ( .A1(fract_out_q[2]), .A2(n4595), .B1(fract_i2f[51]), .B2(
        n4661), .ZN(n3978) );
  AOI221_X2 U1953 ( .B1(n4571), .B2(quo[11]), .C1(n4569), .C2(prod[9]), .A(
        n3979), .ZN(n2718) );
  AND2_X2 U1954 ( .A1(fract_i2f[9]), .A2(n4662), .ZN(n3979) );
  NOR4_X2 U1955 ( .A1(n6440), .A2(n6441), .A3(n6442), .A4(n6443), .ZN(n3970)
         );
  AOI221_X2 U1956 ( .B1(n4571), .B2(quo[12]), .C1(n4569), .C2(prod[10]), .A(
        n3980), .ZN(n3876) );
  AND2_X2 U1957 ( .A1(fract_i2f[10]), .A2(n4662), .ZN(n3980) );
  AOI221_X2 U1958 ( .B1(n4571), .B2(quo[20]), .C1(n4569), .C2(prod[18]), .A(
        n3981), .ZN(n2636) );
  AND2_X2 U1959 ( .A1(fract_i2f[18]), .A2(n4662), .ZN(n3981) );
  AOI221_X2 U1960 ( .B1(n4571), .B2(quo[28]), .C1(n4569), .C2(prod[26]), .A(
        n3982), .ZN(n2605) );
  AND2_X2 U1961 ( .A1(fract_i2f[26]), .A2(n4662), .ZN(n3982) );
  AOI221_X2 U1962 ( .B1(n4571), .B2(quo[36]), .C1(n4569), .C2(prod[34]), .A(
        n3983), .ZN(n2633) );
  AND2_X2 U1963 ( .A1(fract_i2f[34]), .A2(n4662), .ZN(n3983) );
  NOR4_X2 U1964 ( .A1(n2561), .A2(n2635), .A3(n2604), .A4(n2634), .ZN(n3969)
         );
  OR3_X2 U1965 ( .A1(n6433), .A2(n6434), .A3(n2697), .ZN(n2634) );
  AOI221_X2 U1968 ( .B1(n4571), .B2(quo[41]), .C1(n4569), .C2(prod[39]), .A(
        n3985), .ZN(n3984) );
  AND2_X2 U1969 ( .A1(fract_i2f[39]), .A2(n4662), .ZN(n3985) );
  AOI221_X2 U1970 ( .B1(n4571), .B2(quo[43]), .C1(n4568), .C2(prod[41]), .A(
        n3986), .ZN(n2768) );
  AND2_X2 U1971 ( .A1(fract_i2f[41]), .A2(n4662), .ZN(n3986) );
  AOI221_X2 U1972 ( .B1(n4571), .B2(quo[42]), .C1(n4568), .C2(prod[40]), .A(
        n3987), .ZN(n2680) );
  AND2_X2 U1973 ( .A1(fract_i2f[40]), .A2(n4662), .ZN(n3987) );
  AOI221_X2 U1974 ( .B1(n4571), .B2(quo[40]), .C1(n4568), .C2(prod[38]), .A(
        n3988), .ZN(n2752) );
  AND2_X2 U1975 ( .A1(fract_i2f[38]), .A2(n4662), .ZN(n3988) );
  AOI221_X2 U1976 ( .B1(n4575), .B2(quo[39]), .C1(n4568), .C2(prod[37]), .A(
        n3989), .ZN(n3174) );
  AND2_X2 U1977 ( .A1(fract_i2f[37]), .A2(n4662), .ZN(n3989) );
  AOI221_X2 U1978 ( .B1(n4575), .B2(quo[38]), .C1(n4568), .C2(prod[36]), .A(
        n3990), .ZN(n2696) );
  AND2_X2 U1979 ( .A1(fract_i2f[36]), .A2(n4662), .ZN(n3990) );
  AOI221_X2 U1980 ( .B1(n4575), .B2(quo[37]), .C1(n4568), .C2(prod[35]), .A(
        n3991), .ZN(n2758) );
  AND2_X2 U1981 ( .A1(fract_i2f[35]), .A2(n4662), .ZN(n3991) );
  AND3_X2 U1983 ( .A1(n3175), .A2(n2739), .A3(n2669), .ZN(n2708) );
  AOI221_X2 U1985 ( .B1(n4575), .B2(quo[33]), .C1(n4568), .C2(prod[31]), .A(
        n3993), .ZN(n3992) );
  AND2_X2 U1986 ( .A1(fract_i2f[31]), .A2(n4662), .ZN(n3993) );
  AOI221_X2 U1987 ( .B1(n4575), .B2(quo[35]), .C1(n4568), .C2(prod[33]), .A(
        n3994), .ZN(n2722) );
  AND2_X2 U1988 ( .A1(fract_i2f[33]), .A2(n4662), .ZN(n3994) );
  AOI221_X2 U1989 ( .B1(n4575), .B2(quo[34]), .C1(n4568), .C2(prod[32]), .A(
        n3995), .ZN(n2681) );
  AND2_X2 U1990 ( .A1(fract_i2f[32]), .A2(n4662), .ZN(n3995) );
  AOI221_X2 U1991 ( .B1(n4575), .B2(quo[32]), .C1(n4568), .C2(prod[30]), .A(
        n3996), .ZN(n2739) );
  AND2_X2 U1992 ( .A1(fract_i2f[30]), .A2(n4662), .ZN(n3996) );
  AOI221_X2 U1993 ( .B1(n4575), .B2(quo[31]), .C1(n4568), .C2(prod[29]), .A(
        n3997), .ZN(n3175) );
  AND2_X2 U1994 ( .A1(fract_i2f[29]), .A2(n4662), .ZN(n3997) );
  AOI221_X2 U1995 ( .B1(n4575), .B2(quo[30]), .C1(n4568), .C2(prod[28]), .A(
        n3998), .ZN(n2730) );
  AND2_X2 U1996 ( .A1(fract_i2f[28]), .A2(n4662), .ZN(n3998) );
  AOI221_X2 U1997 ( .B1(n4575), .B2(quo[29]), .C1(n4568), .C2(prod[27]), .A(
        n3999), .ZN(n3176) );
  AND2_X2 U1998 ( .A1(fract_i2f[27]), .A2(n4662), .ZN(n3999) );
  AND3_X2 U2000 ( .A1(n3177), .A2(n2753), .A3(n2660), .ZN(n2695) );
  AOI221_X2 U2002 ( .B1(n4575), .B2(quo[25]), .C1(n4568), .C2(prod[23]), .A(
        n4001), .ZN(n4000) );
  AND2_X2 U2003 ( .A1(fract_i2f[23]), .A2(n4662), .ZN(n4001) );
  AOI221_X2 U2004 ( .B1(n4572), .B2(quo[27]), .C1(n4568), .C2(prod[25]), .A(
        n4002), .ZN(n2685) );
  AND2_X2 U2005 ( .A1(fract_i2f[25]), .A2(n4662), .ZN(n4002) );
  AOI221_X2 U2006 ( .B1(n4572), .B2(quo[26]), .C1(n4568), .C2(prod[24]), .A(
        n4003), .ZN(n2769) );
  AND2_X2 U2007 ( .A1(fract_i2f[24]), .A2(n4662), .ZN(n4003) );
  AOI221_X2 U2008 ( .B1(n4572), .B2(quo[24]), .C1(n4568), .C2(prod[22]), .A(
        n4004), .ZN(n2753) );
  AND2_X2 U2009 ( .A1(fract_i2f[22]), .A2(n4662), .ZN(n4004) );
  AOI221_X2 U2010 ( .B1(n4572), .B2(quo[23]), .C1(n4568), .C2(prod[21]), .A(
        n4005), .ZN(n3177) );
  AND2_X2 U2011 ( .A1(fract_i2f[21]), .A2(n4662), .ZN(n4005) );
  AOI221_X2 U2012 ( .B1(n4572), .B2(quo[22]), .C1(n4568), .C2(prod[20]), .A(
        n4006), .ZN(n2762) );
  AND2_X2 U2013 ( .A1(fract_i2f[20]), .A2(n4662), .ZN(n4006) );
  AOI221_X2 U2014 ( .B1(n4572), .B2(quo[21]), .C1(n4568), .C2(prod[19]), .A(
        n4007), .ZN(n3178) );
  AND2_X2 U2015 ( .A1(fract_i2f[19]), .A2(n4662), .ZN(n4007) );
  AND3_X2 U2017 ( .A1(n3179), .A2(n2740), .A3(n2670), .ZN(n2709) );
  AOI221_X2 U2019 ( .B1(n4572), .B2(quo[17]), .C1(n4568), .C2(prod[15]), .A(
        n4009), .ZN(n4008) );
  AND2_X2 U2020 ( .A1(fract_i2f[15]), .A2(n4662), .ZN(n4009) );
  AOI221_X2 U2021 ( .B1(n4572), .B2(quo[19]), .C1(n4568), .C2(prod[17]), .A(
        n4010), .ZN(n2593) );
  AND2_X2 U2022 ( .A1(fract_i2f[17]), .A2(n4662), .ZN(n4010) );
  AOI221_X2 U2023 ( .B1(n4572), .B2(quo[18]), .C1(n4568), .C2(prod[16]), .A(
        n4011), .ZN(n2745) );
  AND2_X2 U2024 ( .A1(fract_i2f[16]), .A2(n4662), .ZN(n4011) );
  AOI221_X2 U2025 ( .B1(n4572), .B2(quo[16]), .C1(n4568), .C2(prod[14]), .A(
        n4012), .ZN(n2740) );
  AND2_X2 U2026 ( .A1(fract_i2f[14]), .A2(n4662), .ZN(n4012) );
  AOI221_X2 U2027 ( .B1(n4572), .B2(quo[15]), .C1(n4568), .C2(prod[13]), .A(
        n4013), .ZN(n3179) );
  AND2_X2 U2028 ( .A1(fract_i2f[13]), .A2(n4662), .ZN(n4013) );
  AOI221_X2 U2029 ( .B1(n4574), .B2(quo[14]), .C1(n4568), .C2(prod[12]), .A(
        n4014), .ZN(n2731) );
  AND2_X2 U2030 ( .A1(fract_i2f[12]), .A2(n4662), .ZN(n4014) );
  AOI221_X2 U2031 ( .B1(n4572), .B2(quo[13]), .C1(n4568), .C2(prod[11]), .A(
        n4015), .ZN(n3180) );
  AND2_X2 U2032 ( .A1(fract_i2f[11]), .A2(fpu_op_r3[2]), .ZN(n4015) );
  NAND4_X2 U2034 ( .A1(n2698), .A2(n2644), .A3(n4016), .A4(n4017), .ZN(n3912)
         );
  NOR4_X2 U2035 ( .A1(n4018), .A2(fract_denorm[66]), .A3(fract_denorm[82]), 
        .A4(fract_denorm[74]), .ZN(n4017) );
  OAI211_X2 U2036 ( .C1(n3973), .C2(n4298), .A(n4019), .B(n4020), .ZN(
        fract_denorm[74]) );
  AOI22_X2 U2037 ( .A1(fract_out_q[25]), .A2(n4595), .B1(fract_i2f[74]), .B2(
        n4661), .ZN(n4020) );
  AOI22_X2 U2038 ( .A1(quo[24]), .A2(n4563), .B1(quo[76]), .B2(n4575), .ZN(
        n4019) );
  OAI211_X2 U2039 ( .C1(n3973), .C2(n4416), .A(n4021), .B(n4022), .ZN(
        fract_denorm[82]) );
  AOI22_X2 U2040 ( .A1(fract_out_q[33]), .A2(n4595), .B1(fract_i2f[82]), .B2(
        n4661), .ZN(n4022) );
  AOI22_X2 U2041 ( .A1(quo[32]), .A2(n4563), .B1(quo[84]), .B2(n4575), .ZN(
        n4021) );
  OAI211_X2 U2042 ( .C1(n3973), .C2(n4423), .A(n4023), .B(n4024), .ZN(
        fract_denorm[66]) );
  AOI22_X2 U2043 ( .A1(fract_out_q[17]), .A2(n4595), .B1(fract_i2f[66]), .B2(
        n4661), .ZN(n4024) );
  AOI22_X2 U2044 ( .A1(quo[16]), .A2(n4563), .B1(quo[68]), .B2(n4574), .ZN(
        n4023) );
  NAND2_X2 U2045 ( .A1(n6400), .A2(n6401), .ZN(n4018) );
  OAI211_X2 U2046 ( .C1(n3973), .C2(n4430), .A(n4025), .B(n4026), .ZN(
        fract_denorm[58]) );
  AOI22_X2 U2047 ( .A1(fract_out_q[9]), .A2(n4595), .B1(fract_i2f[58]), .B2(
        n4661), .ZN(n4026) );
  AOI22_X2 U2048 ( .A1(quo[8]), .A2(n4563), .B1(quo[60]), .B2(n4575), .ZN(
        n4025) );
  OAI211_X2 U2049 ( .C1(n3973), .C2(n4429), .A(n4027), .B(n4028), .ZN(
        fract_denorm[52]) );
  AOI22_X2 U2050 ( .A1(fract_out_q[3]), .A2(n4595), .B1(fract_i2f[52]), .B2(
        n4661), .ZN(n4028) );
  OAI211_X2 U2056 ( .C1(n3973), .C2(n4422), .A(n4029), .B(n4030), .ZN(
        fract_denorm[71]) );
  AOI22_X2 U2057 ( .A1(fract_out_q[22]), .A2(n4595), .B1(fract_i2f[71]), .B2(
        n4661), .ZN(n4030) );
  AOI22_X2 U2058 ( .A1(quo[21]), .A2(n4563), .B1(quo[73]), .B2(n4571), .ZN(
        n4029) );
  OAI211_X2 U2059 ( .C1(n3973), .C2(n4407), .A(n4031), .B(n4032), .ZN(
        fract_denorm[73]) );
  AOI22_X2 U2060 ( .A1(fract_out_q[24]), .A2(n4595), .B1(fract_i2f[73]), .B2(
        n4661), .ZN(n4032) );
  AOI22_X2 U2061 ( .A1(quo[23]), .A2(n4563), .B1(quo[75]), .B2(n4574), .ZN(
        n4031) );
  OAI211_X2 U2062 ( .C1(n3973), .C2(n4313), .A(n4033), .B(n4034), .ZN(
        fract_denorm[72]) );
  AOI22_X2 U2063 ( .A1(fract_out_q[23]), .A2(n4595), .B1(fract_i2f[72]), .B2(
        n4661), .ZN(n4034) );
  AOI22_X2 U2064 ( .A1(quo[22]), .A2(n4563), .B1(quo[74]), .B2(n4575), .ZN(
        n4033) );
  OAI211_X2 U2065 ( .C1(n3973), .C2(n4415), .A(n4035), .B(n4036), .ZN(
        fract_denorm[70]) );
  AOI22_X2 U2066 ( .A1(fract_out_q[21]), .A2(n4595), .B1(fract_i2f[70]), .B2(
        n4661), .ZN(n4036) );
  AOI22_X2 U2067 ( .A1(quo[20]), .A2(n4563), .B1(quo[72]), .B2(n4574), .ZN(
        n4035) );
  OAI211_X2 U2068 ( .C1(n4567), .C2(n4342), .A(n4037), .B(n4038), .ZN(
        fract_denorm[69]) );
  AOI22_X2 U2069 ( .A1(fract_out_q[20]), .A2(n4595), .B1(fract_i2f[69]), .B2(
        n4661), .ZN(n4038) );
  AOI22_X2 U2070 ( .A1(quo[19]), .A2(n4563), .B1(quo[71]), .B2(n4574), .ZN(
        n4037) );
  OAI211_X2 U2071 ( .C1(n4567), .C2(n4402), .A(n4039), .B(n4040), .ZN(
        fract_denorm[68]) );
  AOI22_X2 U2072 ( .A1(fract_out_q[19]), .A2(n4595), .B1(fract_i2f[68]), .B2(
        n4661), .ZN(n4040) );
  AOI22_X2 U2073 ( .A1(quo[18]), .A2(n4563), .B1(quo[70]), .B2(n4574), .ZN(
        n4039) );
  OAI211_X2 U2074 ( .C1(n4567), .C2(n4311), .A(n4041), .B(n4042), .ZN(
        fract_denorm[67]) );
  AOI22_X2 U2075 ( .A1(fract_out_q[18]), .A2(n4595), .B1(fract_i2f[67]), .B2(
        n4661), .ZN(n4042) );
  AOI22_X2 U2076 ( .A1(quo[17]), .A2(n4563), .B1(quo[69]), .B2(n4575), .ZN(
        n4041) );
  OR3_X2 U2077 ( .A1(fract_denorm[59]), .A2(fract_denorm[60]), .A3(n6388), 
        .ZN(n2592) );
  OAI211_X2 U2080 ( .C1(n4567), .C2(n4297), .A(n4043), .B(n4044), .ZN(
        fract_denorm[63]) );
  AOI22_X2 U2081 ( .A1(fract_out_q[14]), .A2(n4595), .B1(fract_i2f[63]), .B2(
        n4661), .ZN(n4044) );
  AOI22_X2 U2082 ( .A1(quo[13]), .A2(n4563), .B1(quo[65]), .B2(n4574), .ZN(
        n4043) );
  OAI211_X2 U2083 ( .C1(n4567), .C2(n4414), .A(n4045), .B(n4046), .ZN(
        fract_denorm[65]) );
  AOI22_X2 U2084 ( .A1(fract_out_q[16]), .A2(n4595), .B1(fract_i2f[65]), .B2(
        n4662), .ZN(n4046) );
  AOI22_X2 U2085 ( .A1(quo[15]), .A2(n4563), .B1(quo[67]), .B2(n4574), .ZN(
        n4045) );
  OAI211_X2 U2086 ( .C1(n4567), .C2(n4428), .A(n4047), .B(n4048), .ZN(
        fract_denorm[64]) );
  AOI22_X2 U2087 ( .A1(fract_out_q[15]), .A2(n4595), .B1(fract_i2f[64]), .B2(
        n4662), .ZN(n4048) );
  AOI22_X2 U2088 ( .A1(quo[14]), .A2(n4563), .B1(quo[66]), .B2(n4574), .ZN(
        n4047) );
  OAI211_X2 U2089 ( .C1(n4567), .C2(n4312), .A(n4049), .B(n4050), .ZN(
        fract_denorm[62]) );
  AOI22_X2 U2090 ( .A1(fract_out_q[13]), .A2(n4595), .B1(fract_i2f[62]), .B2(
        n4662), .ZN(n4050) );
  AOI22_X2 U2091 ( .A1(quo[12]), .A2(n4563), .B1(quo[64]), .B2(n4574), .ZN(
        n4049) );
  OAI211_X2 U2092 ( .C1(n4567), .C2(n4406), .A(n4051), .B(n4052), .ZN(
        fract_denorm[61]) );
  AOI22_X2 U2093 ( .A1(fract_out_q[12]), .A2(n4595), .B1(fract_i2f[61]), .B2(
        n4662), .ZN(n4052) );
  AOI22_X2 U2094 ( .A1(quo[11]), .A2(n4563), .B1(quo[63]), .B2(n4573), .ZN(
        n4051) );
  OAI211_X2 U2095 ( .C1(n4567), .C2(n4346), .A(n4053), .B(n4054), .ZN(
        fract_denorm[60]) );
  AOI22_X2 U2096 ( .A1(fract_out_q[11]), .A2(n4595), .B1(fract_i2f[60]), .B2(
        n4662), .ZN(n4054) );
  AOI22_X2 U2097 ( .A1(quo[10]), .A2(n4563), .B1(quo[62]), .B2(n4575), .ZN(
        n4053) );
  OAI211_X2 U2098 ( .C1(n4567), .C2(n4413), .A(n4055), .B(n4056), .ZN(
        fract_denorm[59]) );
  AOI22_X2 U2099 ( .A1(fract_out_q[10]), .A2(n4595), .B1(fract_i2f[59]), .B2(
        n4662), .ZN(n4056) );
  AOI22_X2 U2100 ( .A1(quo[9]), .A2(n4563), .B1(quo[61]), .B2(n4573), .ZN(
        n4055) );
  OAI211_X2 U2104 ( .C1(n4567), .C2(n4436), .A(n4057), .B(n4058), .ZN(
        fract_denorm[79]) );
  AOI22_X2 U2105 ( .A1(fract_out_q[30]), .A2(n4595), .B1(fract_i2f[79]), .B2(
        n4662), .ZN(n4058) );
  AOI22_X2 U2106 ( .A1(quo[29]), .A2(n4563), .B1(quo[81]), .B2(n4571), .ZN(
        n4057) );
  OAI211_X2 U2107 ( .C1(n4566), .C2(n4427), .A(n4059), .B(n4060), .ZN(
        fract_denorm[81]) );
  AOI22_X2 U2108 ( .A1(fract_out_q[32]), .A2(n4595), .B1(fract_i2f[81]), .B2(
        n4662), .ZN(n4060) );
  AOI22_X2 U2109 ( .A1(quo[31]), .A2(n4563), .B1(quo[83]), .B2(n4573), .ZN(
        n4059) );
  OAI211_X2 U2110 ( .C1(n4566), .C2(n4437), .A(n4061), .B(n4062), .ZN(
        fract_denorm[80]) );
  AOI22_X2 U2111 ( .A1(fract_out_q[31]), .A2(n4595), .B1(fract_i2f[80]), .B2(
        n4662), .ZN(n4062) );
  AOI22_X2 U2112 ( .A1(quo[30]), .A2(n4563), .B1(quo[82]), .B2(n4574), .ZN(
        n4061) );
  OAI211_X2 U2113 ( .C1(n4566), .C2(n4421), .A(n4063), .B(n4064), .ZN(
        fract_denorm[78]) );
  AOI22_X2 U2114 ( .A1(fract_out_q[29]), .A2(n4595), .B1(fract_i2f[78]), .B2(
        n4662), .ZN(n4064) );
  AOI22_X2 U2115 ( .A1(quo[28]), .A2(n4563), .B1(quo[80]), .B2(n4573), .ZN(
        n4063) );
  OAI211_X2 U2116 ( .C1(n3973), .C2(n4412), .A(n4065), .B(n4066), .ZN(
        fract_denorm[77]) );
  AOI22_X2 U2117 ( .A1(fract_out_q[28]), .A2(n4595), .B1(fract_i2f[77]), .B2(
        n4662), .ZN(n4066) );
  AOI22_X2 U2118 ( .A1(quo[27]), .A2(n4563), .B1(quo[79]), .B2(n4575), .ZN(
        n4065) );
  OAI211_X2 U2119 ( .C1(n3973), .C2(n4426), .A(n4067), .B(n4068), .ZN(
        fract_denorm[76]) );
  AOI22_X2 U2120 ( .A1(fract_out_q[27]), .A2(n4595), .B1(fract_i2f[76]), .B2(
        n4662), .ZN(n4068) );
  AOI22_X2 U2121 ( .A1(quo[26]), .A2(n4563), .B1(quo[78]), .B2(n4573), .ZN(
        n4067) );
  OAI211_X2 U2122 ( .C1(n3973), .C2(n4343), .A(n4069), .B(n4070), .ZN(
        fract_denorm[75]) );
  AOI22_X2 U2123 ( .A1(fract_out_q[26]), .A2(n4595), .B1(fract_i2f[75]), .B2(
        n4662), .ZN(n4070) );
  AOI22_X2 U2124 ( .A1(quo[25]), .A2(n4563), .B1(quo[77]), .B2(n4575), .ZN(
        n4069) );
  OAI211_X2 U2128 ( .C1(n3973), .C2(n4294), .A(n4071), .B(n4072), .ZN(
        fract_denorm[87]) );
  AOI22_X2 U2129 ( .A1(fract_out_q[38]), .A2(n4595), .B1(fract_i2f[87]), .B2(
        n4662), .ZN(n4072) );
  AOI22_X2 U2130 ( .A1(quo[37]), .A2(n4563), .B1(quo[89]), .B2(n4571), .ZN(
        n4071) );
  OAI211_X2 U2131 ( .C1(n3973), .C2(n4411), .A(n4073), .B(n4074), .ZN(
        fract_denorm[89]) );
  AOI22_X2 U2132 ( .A1(fract_out_q[40]), .A2(n4595), .B1(fract_i2f[89]), .B2(
        n4662), .ZN(n4074) );
  AOI22_X2 U2133 ( .A1(quo[39]), .A2(n4563), .B1(quo[91]), .B2(n4574), .ZN(
        n4073) );
  OAI211_X2 U2134 ( .C1(n3973), .C2(n4425), .A(n4075), .B(n4076), .ZN(
        fract_denorm[88]) );
  AOI22_X2 U2135 ( .A1(fract_out_q[39]), .A2(n4595), .B1(fract_i2f[88]), .B2(
        n4662), .ZN(n4076) );
  AOI22_X2 U2136 ( .A1(quo[38]), .A2(n4563), .B1(quo[90]), .B2(n4572), .ZN(
        n4075) );
  OAI211_X2 U2137 ( .C1(n3973), .C2(n4307), .A(n4077), .B(n4078), .ZN(
        fract_denorm[86]) );
  AOI22_X2 U2138 ( .A1(fract_out_q[37]), .A2(n4595), .B1(fract_i2f[86]), .B2(
        n4662), .ZN(n4078) );
  AOI22_X2 U2139 ( .A1(quo[36]), .A2(n4563), .B1(quo[88]), .B2(n4574), .ZN(
        n4077) );
  OAI211_X2 U2140 ( .C1(n3973), .C2(n4404), .A(n4079), .B(n4080), .ZN(
        fract_denorm[85]) );
  AOI22_X2 U2141 ( .A1(fract_out_q[36]), .A2(n4595), .B1(fract_i2f[85]), .B2(
        n4662), .ZN(n4080) );
  AOI22_X2 U2142 ( .A1(quo[35]), .A2(n4563), .B1(quo[87]), .B2(n4571), .ZN(
        n4079) );
  OAI211_X2 U2143 ( .C1(n4567), .C2(n4344), .A(n4081), .B(n4082), .ZN(
        fract_denorm[84]) );
  AOI22_X2 U2144 ( .A1(fract_out_q[35]), .A2(n4595), .B1(fract_i2f[84]), .B2(
        n4662), .ZN(n4082) );
  AOI22_X2 U2145 ( .A1(quo[34]), .A2(n4564), .B1(quo[86]), .B2(n4573), .ZN(
        n4081) );
  OAI211_X2 U2146 ( .C1(n4567), .C2(n4420), .A(n4083), .B(n4084), .ZN(
        fract_denorm[83]) );
  AOI22_X2 U2147 ( .A1(fract_out_q[34]), .A2(n4595), .B1(fract_i2f[83]), .B2(
        n4662), .ZN(n4084) );
  AOI22_X2 U2148 ( .A1(quo[33]), .A2(n4564), .B1(quo[85]), .B2(n4571), .ZN(
        n4083) );
  OAI211_X2 U2151 ( .C1(n4567), .C2(n4310), .A(n4085), .B(n4086), .ZN(
        fract_denorm[55]) );
  AOI22_X2 U2152 ( .A1(fract_out_q[6]), .A2(n4595), .B1(fract_i2f[55]), .B2(
        n4662), .ZN(n4086) );
  AOI22_X2 U2153 ( .A1(quo[5]), .A2(n4564), .B1(quo[57]), .B2(n4575), .ZN(
        n4085) );
  OAI211_X2 U2154 ( .C1(n4567), .C2(n4341), .A(n4087), .B(n4088), .ZN(
        fract_denorm[57]) );
  AOI22_X2 U2155 ( .A1(fract_out_q[8]), .A2(n4595), .B1(fract_i2f[57]), .B2(
        n4662), .ZN(n4088) );
  AOI22_X2 U2156 ( .A1(quo[7]), .A2(n4564), .B1(quo[59]), .B2(n4575), .ZN(
        n4087) );
  OAI211_X2 U2157 ( .C1(n4567), .C2(n4401), .A(n4089), .B(n4090), .ZN(
        fract_denorm[56]) );
  AOI22_X2 U2158 ( .A1(fract_out_q[7]), .A2(n4595), .B1(fract_i2f[56]), .B2(
        n4662), .ZN(n4090) );
  AOI22_X2 U2159 ( .A1(quo[6]), .A2(n4564), .B1(quo[58]), .B2(n4575), .ZN(
        n4089) );
  OAI211_X2 U2160 ( .C1(n4567), .C2(n4419), .A(n4091), .B(n4092), .ZN(
        fract_denorm[54]) );
  AOI22_X2 U2161 ( .A1(fract_out_q[5]), .A2(n4595), .B1(fract_i2f[54]), .B2(
        n4662), .ZN(n4092) );
  AOI22_X2 U2162 ( .A1(quo[4]), .A2(n4564), .B1(quo[56]), .B2(n4575), .ZN(
        n4091) );
  OAI211_X2 U2163 ( .C1(n4567), .C2(n4410), .A(n4093), .B(n4094), .ZN(
        fract_denorm[53]) );
  AOI22_X2 U2164 ( .A1(fract_out_q[4]), .A2(n4595), .B1(fract_i2f[53]), .B2(
        fpu_op_r3[2]), .ZN(n4094) );
  AOI22_X2 U2165 ( .A1(quo[3]), .A2(n4564), .B1(quo[55]), .B2(n4571), .ZN(
        n4093) );
  AND3_X2 U2167 ( .A1(n3172), .A2(n2737), .A3(n2668), .ZN(n2706) );
  AOI221_X2 U2169 ( .B1(n4571), .B2(quo[49]), .C1(n4568), .C2(prod[47]), .A(
        n4096), .ZN(n4095) );
  AND2_X2 U2170 ( .A1(fract_i2f[47]), .A2(fpu_op_r3[2]), .ZN(n4096) );
  AOI221_X2 U2171 ( .B1(n4573), .B2(quo[51]), .C1(n4568), .C2(prod[49]), .A(
        n6368), .ZN(n2711) );
  AOI22_X2 U2172 ( .A1(fract_out_q[0]), .A2(n4595), .B1(fract_i2f[49]), .B2(
        fpu_op_r3[2]), .ZN(n4097) );
  AOI221_X2 U2173 ( .B1(n4573), .B2(quo[50]), .C1(n4568), .C2(prod[48]), .A(
        n4098), .ZN(n2744) );
  AND2_X2 U2174 ( .A1(fract_i2f[48]), .A2(fpu_op_r3[2]), .ZN(n4098) );
  AOI221_X2 U2175 ( .B1(n4573), .B2(quo[48]), .C1(n4568), .C2(prod[46]), .A(
        n4099), .ZN(n2737) );
  AND2_X2 U2176 ( .A1(fract_i2f[46]), .A2(fpu_op_r3[2]), .ZN(n4099) );
  AOI221_X2 U2177 ( .B1(n4571), .B2(quo[47]), .C1(n4568), .C2(prod[45]), .A(
        n4100), .ZN(n3172) );
  AND2_X2 U2178 ( .A1(fract_i2f[45]), .A2(fpu_op_r3[2]), .ZN(n4100) );
  AOI221_X2 U2179 ( .B1(n4573), .B2(quo[46]), .C1(n4568), .C2(prod[44]), .A(
        n4101), .ZN(n2729) );
  AND2_X2 U2180 ( .A1(fract_i2f[44]), .A2(fpu_op_r3[2]), .ZN(n4101) );
  AOI221_X2 U2181 ( .B1(n4573), .B2(quo[45]), .C1(n4568), .C2(prod[43]), .A(
        n4102), .ZN(n3173) );
  AND2_X2 U2182 ( .A1(fract_i2f[43]), .A2(fpu_op_r3[2]), .ZN(n4102) );
  NAND2_X2 U2184 ( .A1(n2638), .A2(n6365), .ZN(n2598) );
  OAI211_X2 U2185 ( .C1(n4566), .C2(n4435), .A(n4103), .B(n4104), .ZN(
        fract_denorm[98]) );
  AOI22_X2 U2186 ( .A1(fract_out_q[49]), .A2(n3315), .B1(fract_i2f[98]), .B2(
        n4661), .ZN(n4104) );
  AOI22_X2 U2187 ( .A1(quo[48]), .A2(n4564), .B1(quo[100]), .B2(n4571), .ZN(
        n4103) );
  AND3_X2 U2188 ( .A1(n6360), .A2(n4654), .A3(n2761), .ZN(n2638) );
  OR3_X2 U2190 ( .A1(fract_denorm[101]), .A2(fract_denorm[102]), .A3(
        fract_denorm[100]), .ZN(n2662) );
  OAI211_X2 U2191 ( .C1(n4566), .C2(n4409), .A(n4105), .B(n4106), .ZN(
        fract_denorm[100]) );
  AOI22_X2 U2192 ( .A1(fract_out_q[51]), .A2(n3315), .B1(fract_i2f[100]), .B2(
        n4661), .ZN(n4106) );
  AOI22_X2 U2193 ( .A1(quo[50]), .A2(n4309), .B1(quo[102]), .B2(n4570), .ZN(
        n4105) );
  OAI211_X2 U2194 ( .C1(n4566), .C2(n4306), .A(n4107), .B(n4108), .ZN(
        fract_denorm[102]) );
  AOI22_X2 U2195 ( .A1(fract_out_q[53]), .A2(n3315), .B1(fract_i2f[102]), .B2(
        n4661), .ZN(n4108) );
  AOI22_X2 U2196 ( .A1(quo[52]), .A2(n4309), .B1(quo[104]), .B2(n4570), .ZN(
        n4107) );
  OAI211_X2 U2197 ( .C1(n4566), .C2(n4418), .A(n4109), .B(n4110), .ZN(
        fract_denorm[101]) );
  AOI22_X2 U2198 ( .A1(fract_out_q[52]), .A2(n3315), .B1(fract_i2f[101]), .B2(
        n4662), .ZN(n4110) );
  AOI22_X2 U2199 ( .A1(quo[51]), .A2(n4309), .B1(quo[103]), .B2(n4570), .ZN(
        n4109) );
  OAI211_X2 U2200 ( .C1(n4566), .C2(n4338), .A(n4111), .B(n4112), .ZN(
        fract_denorm[104]) );
  AOI22_X2 U2201 ( .A1(fract_out_q[55]), .A2(n3315), .B1(fract_i2f[104]), .B2(
        n4661), .ZN(n4112) );
  OAI211_X2 U2203 ( .C1(n4566), .C2(n4403), .A(n4113), .B(n4114), .ZN(
        fract_denorm[103]) );
  AOI22_X2 U2204 ( .A1(fract_out_q[54]), .A2(n3315), .B1(fract_i2f[103]), .B2(
        n4661), .ZN(n4114) );
  OAI211_X2 U2206 ( .C1(n4566), .C2(n4433), .A(n4115), .B(n4116), .ZN(
        fract_denorm[99]) );
  AOI22_X2 U2207 ( .A1(fract_out_q[50]), .A2(n4595), .B1(fract_i2f[99]), .B2(
        n4662), .ZN(n4116) );
  AOI22_X2 U2208 ( .A1(quo[49]), .A2(n4564), .B1(quo[101]), .B2(n4571), .ZN(
        n4115) );
  OAI211_X2 U2209 ( .C1(n4566), .C2(n4345), .A(n4117), .B(n4118), .ZN(
        fract_denorm[90]) );
  AOI22_X2 U2210 ( .A1(fract_out_q[41]), .A2(n3315), .B1(fract_i2f[90]), .B2(
        n4661), .ZN(n4118) );
  AOI22_X2 U2211 ( .A1(quo[40]), .A2(n4564), .B1(quo[92]), .B2(n4571), .ZN(
        n4117) );
  OAI211_X2 U2215 ( .C1(n4566), .C2(n4408), .A(n4119), .B(n4120), .ZN(
        fract_denorm[95]) );
  AOI22_X2 U2216 ( .A1(fract_out_q[46]), .A2(n3315), .B1(fract_i2f[95]), .B2(
        n4661), .ZN(n4120) );
  AOI22_X2 U2217 ( .A1(quo[45]), .A2(n4564), .B1(quo[97]), .B2(n4572), .ZN(
        n4119) );
  OAI211_X2 U2218 ( .C1(n4566), .C2(n4431), .A(n4121), .B(n4122), .ZN(
        fract_denorm[97]) );
  AOI22_X2 U2219 ( .A1(fract_out_q[48]), .A2(n3315), .B1(fract_i2f[97]), .B2(
        n4661), .ZN(n4122) );
  AOI22_X2 U2220 ( .A1(quo[47]), .A2(n4564), .B1(quo[99]), .B2(n4573), .ZN(
        n4121) );
  OAI211_X2 U2221 ( .C1(n4566), .C2(n4417), .A(n4123), .B(n4124), .ZN(
        fract_denorm[96]) );
  AOI22_X2 U2222 ( .A1(fract_out_q[47]), .A2(n4595), .B1(fract_i2f[96]), .B2(
        n4661), .ZN(n4124) );
  AOI22_X2 U2223 ( .A1(quo[46]), .A2(n4564), .B1(quo[98]), .B2(n4571), .ZN(
        n4123) );
  OAI211_X2 U2224 ( .C1(n4566), .C2(n4424), .A(n4125), .B(n4126), .ZN(
        fract_denorm[94]) );
  AOI22_X2 U2225 ( .A1(fract_out_q[45]), .A2(n3315), .B1(fract_i2f[94]), .B2(
        n4661), .ZN(n4126) );
  AOI22_X2 U2226 ( .A1(quo[44]), .A2(n4564), .B1(quo[96]), .B2(n4572), .ZN(
        n4125) );
  OAI211_X2 U2227 ( .C1(n4566), .C2(n4295), .A(n4127), .B(n4128), .ZN(
        fract_denorm[93]) );
  AOI22_X2 U2228 ( .A1(fract_out_q[44]), .A2(n3315), .B1(fract_i2f[93]), .B2(
        n4661), .ZN(n4128) );
  AOI22_X2 U2229 ( .A1(quo[43]), .A2(n4564), .B1(quo[95]), .B2(n4572), .ZN(
        n4127) );
  OAI211_X2 U2230 ( .C1(n4566), .C2(n4308), .A(n4129), .B(n4130), .ZN(
        fract_denorm[92]) );
  AOI22_X2 U2231 ( .A1(fract_out_q[43]), .A2(n3315), .B1(fract_i2f[92]), .B2(
        n4662), .ZN(n4130) );
  AOI22_X2 U2232 ( .A1(quo[42]), .A2(n4564), .B1(quo[94]), .B2(n4575), .ZN(
        n4129) );
  OAI211_X2 U2233 ( .C1(n4566), .C2(n4405), .A(n4131), .B(n4132), .ZN(
        fract_denorm[91]) );
  AOI22_X2 U2234 ( .A1(fract_out_q[42]), .A2(n4595), .B1(fract_i2f[91]), .B2(
        n4661), .ZN(n4132) );
  AOI22_X2 U2236 ( .A1(quo[41]), .A2(n4564), .B1(quo[93]), .B2(n4571), .ZN(
        n4131) );
  AOI221_X2 U2238 ( .B1(n4571), .B2(quo[10]), .C1(n4568), .C2(prod[8]), .A(
        n4133), .ZN(n2683) );
  AND2_X2 U2239 ( .A1(fract_i2f[8]), .A2(fpu_op_r3[2]), .ZN(n4133) );
  AOI221_X2 U2240 ( .B1(n4573), .B2(quo[9]), .C1(n4568), .C2(prod[7]), .A(
        n4134), .ZN(n2767) );
  AND2_X2 U2241 ( .A1(fract_i2f[7]), .A2(fpu_op_r3[2]), .ZN(n4134) );
  AOI221_X2 U2242 ( .B1(n4573), .B2(quo[8]), .C1(n4568), .C2(prod[6]), .A(
        n4135), .ZN(n2751) );
  AND2_X2 U2243 ( .A1(fract_i2f[6]), .A2(fpu_op_r3[2]), .ZN(n4135) );
  AOI221_X2 U2244 ( .B1(n4573), .B2(quo[7]), .C1(n4568), .C2(prod[5]), .A(
        n4136), .ZN(n3171) );
  AND2_X2 U2245 ( .A1(fract_i2f[5]), .A2(fpu_op_r3[2]), .ZN(n4136) );
  AOI221_X2 U2246 ( .B1(n4574), .B2(quo[6]), .C1(n4568), .C2(prod[4]), .A(
        n4137), .ZN(n2763) );
  AND2_X2 U2247 ( .A1(fract_i2f[4]), .A2(n4662), .ZN(n4137) );
  AOI221_X2 U2248 ( .B1(n4573), .B2(quo[5]), .C1(n4568), .C2(prod[3]), .A(
        n4138), .ZN(n3873) );
  AND2_X2 U2249 ( .A1(fract_i2f[3]), .A2(n4662), .ZN(n4138) );
  AOI221_X2 U2250 ( .B1(n4572), .B2(quo[4]), .C1(n4569), .C2(prod[2]), .A(
        n4139), .ZN(n2724) );
  AND2_X2 U2251 ( .A1(fract_i2f[2]), .A2(n4662), .ZN(n4139) );
  AOI221_X2 U2252 ( .B1(n4571), .B2(quo[3]), .C1(n4568), .C2(prod[1]), .A(
        n4140), .ZN(n3879) );
  AND2_X2 U2253 ( .A1(fract_i2f[1]), .A2(n4662), .ZN(n4140) );
  OAI221_X2 U2256 ( .B1(n6340), .B2(n6460), .C1(n2441), .C2(n4540), .A(n4141), 
        .ZN(n3958) );
  AND2_X2 U2258 ( .A1(n2479), .A2(n3913), .ZN(n2478) );
  NAND2_X2 U2259 ( .A1(exp_ovf_r[1]), .A2(n3488), .ZN(n3913) );
  NAND4_X2 U2265 ( .A1(n4299), .A2(n4347), .A3(n4142), .A4(n4143), .ZN(n2514)
         );
  NOR4_X2 U2266 ( .A1(n4144), .A2(exp_r[1]), .A3(n4655), .A4(n4315), .ZN(n4143) );
  NAND2_X2 U2267 ( .A1(n3965), .A2(n4349), .ZN(n4144) );
  NAND2_X2 U2270 ( .A1(n4145), .A2(n4146), .ZN(n3495) );
  NOR4_X2 U2271 ( .A1(n4147), .A2(n4148), .A3(n4149), .A4(n4150), .ZN(n4146)
         );
  NAND4_X2 U2272 ( .A1(n4151), .A2(n4152), .A3(n4153), .A4(n4154), .ZN(n4150)
         );
  NOR4_X2 U2273 ( .A1(remainder[62]), .A2(remainder[61]), .A3(remainder[60]), 
        .A4(remainder[5]), .ZN(n4154) );
  NAND4_X2 U2277 ( .A1(n4155), .A2(n4156), .A3(n4157), .A4(n4158), .ZN(n4149)
         );
  NOR4_X2 U2278 ( .A1(remainder[75]), .A2(remainder[74]), .A3(remainder[73]), 
        .A4(remainder[72]), .ZN(n4158) );
  NOR4_X2 U2280 ( .A1(remainder[69]), .A2(remainder[68]), .A3(remainder[67]), 
        .A4(remainder[66]), .ZN(n4156) );
  NAND4_X2 U2282 ( .A1(n4159), .A2(n4160), .A3(n4161), .A4(n4162), .ZN(n4148)
         );
  NOR4_X2 U2283 ( .A1(remainder[87]), .A2(remainder[86]), .A3(remainder[85]), 
        .A4(remainder[84]), .ZN(n4162) );
  NAND4_X2 U2287 ( .A1(n4163), .A2(n4164), .A3(n4165), .A4(n4166), .ZN(n4147)
         );
  NOR4_X2 U2288 ( .A1(remainder[9]), .A2(remainder[99]), .A3(remainder[98]), 
        .A4(remainder[97]), .ZN(n4166) );
  NOR4_X2 U2290 ( .A1(remainder[93]), .A2(remainder[92]), .A3(remainder[91]), 
        .A4(remainder[90]), .ZN(n4164) );
  NOR4_X2 U2292 ( .A1(n4167), .A2(n4168), .A3(n4169), .A4(n4170), .ZN(n4145)
         );
  NAND4_X2 U2293 ( .A1(n4171), .A2(n4172), .A3(n4173), .A4(n4174), .ZN(n4170)
         );
  NOR4_X2 U2294 ( .A1(remainder[13]), .A2(remainder[12]), .A3(remainder[11]), 
        .A4(remainder[10]), .ZN(n4174) );
  NAND4_X2 U2298 ( .A1(n4175), .A2(n4176), .A3(n4177), .A4(n4178), .ZN(n4169)
         );
  NOR4_X2 U2299 ( .A1(remainder[26]), .A2(remainder[25]), .A3(remainder[24]), 
        .A4(remainder[23]), .ZN(n4178) );
  NOR4_X2 U2301 ( .A1(remainder[1]), .A2(remainder[19]), .A3(remainder[18]), 
        .A4(remainder[17]), .ZN(n4176) );
  NAND4_X2 U2303 ( .A1(n4179), .A2(n4180), .A3(n4181), .A4(n4182), .ZN(n4168)
         );
  NOR4_X2 U2304 ( .A1(remainder[38]), .A2(remainder[37]), .A3(remainder[36]), 
        .A4(remainder[35]), .ZN(n4182) );
  NAND4_X2 U2308 ( .A1(n4183), .A2(n4184), .A3(n4185), .A4(n4186), .ZN(n4167)
         );
  NOR4_X2 U2309 ( .A1(remainder[50]), .A2(remainder[4]), .A3(remainder[49]), 
        .A4(remainder[48]), .ZN(n4186) );
  NOR4_X2 U2311 ( .A1(remainder[44]), .A2(remainder[43]), .A3(remainder[42]), 
        .A4(remainder[41]), .ZN(n4184) );
  NAND2_X2 U2313 ( .A1(rmode_r3[0]), .A2(n4351), .ZN(n3741) );
  NAND2_X2 U2315 ( .A1(n2507), .A2(n4355), .ZN(n3297) );
  OAI211_X2 U2318 ( .C1(n4355), .C2(n4382), .A(n3303), .B(n4188), .ZN(n4187)
         );
  NAND2_X2 U2320 ( .A1(n4569), .A2(n4291), .ZN(n2507) );
  NAND2_X2 U2321 ( .A1(fpu_op_r3[1]), .A2(n4274), .ZN(n3973) );
  NAND2_X2 U2325 ( .A1(n2434), .A2(n4355), .ZN(n2439) );
  NAND2_X2 U2329 ( .A1(fpu_op_r3[1]), .A2(fpu_op_r3[0]), .ZN(n3458) );
  XOR2_X2 U2330 ( .A(n3065), .B(n4190), .Z(N789) );
  NAND2_X2 U2331 ( .A1(rmode_r2[1]), .A2(rmode_r2[0]), .ZN(n3065) );
  OAI221_X2 U2332 ( .B1(n4561), .B2(n4336), .C1(n4559), .C2(n5958), .A(n4554), 
        .ZN(N769) );
  OAI221_X2 U2333 ( .B1(n4561), .B2(n4335), .C1(n4560), .C2(n5959), .A(n4554), 
        .ZN(N768) );
  OAI221_X2 U2334 ( .B1(n4191), .B2(n4334), .C1(n4559), .C2(n5960), .A(n4554), 
        .ZN(N767) );
  OAI221_X2 U2335 ( .B1(n4191), .B2(n4332), .C1(n4560), .C2(n5961), .A(n4554), 
        .ZN(N766) );
  OAI221_X2 U2336 ( .B1(n4191), .B2(n4331), .C1(n4560), .C2(n5962), .A(n4554), 
        .ZN(N765) );
  OAI221_X2 U2337 ( .B1(n4191), .B2(n4333), .C1(n4560), .C2(n5963), .A(n4554), 
        .ZN(N764) );
  OAI221_X2 U2338 ( .B1(n4191), .B2(n4329), .C1(n4560), .C2(n5964), .A(n4554), 
        .ZN(N763) );
  OAI221_X2 U2339 ( .B1(n4191), .B2(n4483), .C1(n4560), .C2(n5965), .A(n4554), 
        .ZN(N762) );
  OAI221_X2 U2340 ( .B1(n4191), .B2(n4532), .C1(n4560), .C2(n5966), .A(n4554), 
        .ZN(N761) );
  OAI221_X2 U2341 ( .B1(n4191), .B2(n4531), .C1(n4560), .C2(n5967), .A(n4554), 
        .ZN(N760) );
  OAI221_X2 U2342 ( .B1(n4561), .B2(n4530), .C1(n4560), .C2(n5968), .A(n4554), 
        .ZN(N759) );
  OAI221_X2 U2343 ( .B1(n4561), .B2(n4529), .C1(n4560), .C2(n5969), .A(n4555), 
        .ZN(N758) );
  OAI221_X2 U2344 ( .B1(n4561), .B2(n4528), .C1(n4560), .C2(n5970), .A(n4555), 
        .ZN(N757) );
  OAI221_X2 U2345 ( .B1(n4561), .B2(n4527), .C1(n4560), .C2(n5971), .A(n4555), 
        .ZN(N756) );
  OAI221_X2 U2346 ( .B1(n4561), .B2(n4526), .C1(n4559), .C2(n5972), .A(n4555), 
        .ZN(N755) );
  OAI221_X2 U2347 ( .B1(n4561), .B2(n4525), .C1(n4559), .C2(n5973), .A(n4555), 
        .ZN(N754) );
  OAI221_X2 U2348 ( .B1(n4561), .B2(n4524), .C1(n4559), .C2(n5974), .A(n4555), 
        .ZN(N753) );
  OAI221_X2 U2349 ( .B1(n4561), .B2(n4523), .C1(n4559), .C2(n5975), .A(n4555), 
        .ZN(N752) );
  OAI221_X2 U2350 ( .B1(n4561), .B2(n4522), .C1(n4559), .C2(n5976), .A(n4555), 
        .ZN(N751) );
  OAI221_X2 U2351 ( .B1(n4561), .B2(n4521), .C1(n4559), .C2(n5977), .A(n4555), 
        .ZN(N750) );
  OAI221_X2 U2352 ( .B1(n4561), .B2(n4520), .C1(n4559), .C2(n5978), .A(n4555), 
        .ZN(N749) );
  OAI221_X2 U2353 ( .B1(n4561), .B2(n4519), .C1(n4559), .C2(n5979), .A(n4555), 
        .ZN(N748) );
  OAI221_X2 U2354 ( .B1(n4561), .B2(n4518), .C1(n4559), .C2(n5980), .A(n4556), 
        .ZN(N747) );
  OAI221_X2 U2355 ( .B1(n4561), .B2(n4517), .C1(n4559), .C2(n5981), .A(n4556), 
        .ZN(N746) );
  OAI221_X2 U2356 ( .B1(n4561), .B2(n4516), .C1(n4559), .C2(n5982), .A(n4556), 
        .ZN(N745) );
  OAI221_X2 U2357 ( .B1(n4561), .B2(n4515), .C1(n4558), .C2(n5983), .A(n4556), 
        .ZN(N744) );
  OAI221_X2 U2358 ( .B1(n4561), .B2(n4514), .C1(n4557), .C2(n5984), .A(n4556), 
        .ZN(N743) );
  OAI221_X2 U2359 ( .B1(n4561), .B2(n4513), .C1(n4558), .C2(n5985), .A(n4556), 
        .ZN(N742) );
  OAI221_X2 U2360 ( .B1(n4561), .B2(n4512), .C1(n4557), .C2(n5986), .A(n4556), 
        .ZN(N741) );
  OAI221_X2 U2361 ( .B1(n4561), .B2(n4511), .C1(n4558), .C2(n5987), .A(n4556), 
        .ZN(N740) );
  OAI221_X2 U2362 ( .B1(n4561), .B2(n4510), .C1(n4557), .C2(n5988), .A(n4556), 
        .ZN(N739) );
  OAI221_X2 U2363 ( .B1(n4561), .B2(n4509), .C1(n4558), .C2(n5989), .A(n4556), 
        .ZN(N738) );
  OAI221_X2 U2364 ( .B1(n4561), .B2(n4508), .C1(n4557), .C2(n5990), .A(n4556), 
        .ZN(N737) );
  OAI221_X2 U2365 ( .B1(n4561), .B2(n4507), .C1(n4558), .C2(n5991), .A(n4554), 
        .ZN(N736) );
  OAI221_X2 U2366 ( .B1(n4561), .B2(n4506), .C1(n4557), .C2(n5992), .A(n4555), 
        .ZN(N735) );
  OAI221_X2 U2367 ( .B1(n4561), .B2(n4505), .C1(n4558), .C2(n5993), .A(n4556), 
        .ZN(N734) );
  OAI221_X2 U2368 ( .B1(n4561), .B2(n4504), .C1(n4558), .C2(n5994), .A(n4554), 
        .ZN(N733) );
  OAI221_X2 U2369 ( .B1(n4561), .B2(n4503), .C1(n4558), .C2(n5995), .A(n4555), 
        .ZN(N732) );
  OAI221_X2 U2370 ( .B1(n4561), .B2(n4502), .C1(n4558), .C2(n5996), .A(n4556), 
        .ZN(N731) );
  OAI221_X2 U2371 ( .B1(n4561), .B2(n4501), .C1(n4558), .C2(n5997), .A(n4554), 
        .ZN(N730) );
  OAI221_X2 U2372 ( .B1(n4561), .B2(n4500), .C1(n4558), .C2(n5998), .A(n4555), 
        .ZN(N729) );
  OAI221_X2 U2373 ( .B1(n4561), .B2(n4499), .C1(n4558), .C2(n5999), .A(n4556), 
        .ZN(N728) );
  OAI221_X2 U2374 ( .B1(n4561), .B2(n4498), .C1(n4558), .C2(n6000), .A(n4554), 
        .ZN(N727) );
  OAI221_X2 U2375 ( .B1(n4561), .B2(n4497), .C1(n4558), .C2(n6001), .A(n4555), 
        .ZN(N726) );
  OAI221_X2 U2376 ( .B1(n4191), .B2(n4397), .C1(n4558), .C2(n6002), .A(n4556), 
        .ZN(N725) );
  OAI221_X2 U2377 ( .B1(n4191), .B2(n4396), .C1(n4558), .C2(n6003), .A(n4554), 
        .ZN(N724) );
  OAI221_X2 U2378 ( .B1(n4191), .B2(n4395), .C1(n4558), .C2(n6004), .A(n4555), 
        .ZN(N723) );
  OAI221_X2 U2379 ( .B1(n4191), .B2(n4394), .C1(n4557), .C2(n6005), .A(n4554), 
        .ZN(N722) );
  OAI221_X2 U2380 ( .B1(n4191), .B2(n4393), .C1(n4557), .C2(n6006), .A(n4556), 
        .ZN(N721) );
  OAI221_X2 U2381 ( .B1(n4191), .B2(n4392), .C1(n4557), .C2(n6007), .A(n4554), 
        .ZN(N720) );
  OAI221_X2 U2382 ( .B1(n4191), .B2(n4391), .C1(n4557), .C2(n6008), .A(n4555), 
        .ZN(N719) );
  OAI221_X2 U2383 ( .B1(n4191), .B2(n4390), .C1(n4557), .C2(n6009), .A(n4555), 
        .ZN(N718) );
  OAI221_X2 U2384 ( .B1(n4191), .B2(n4389), .C1(n4557), .C2(n6010), .A(n4556), 
        .ZN(N717) );
  OAI221_X2 U2386 ( .B1(n4191), .B2(n4388), .C1(n4557), .C2(n6011), .A(n4195), 
        .ZN(N716) );
  AOI22_X2 U2387 ( .A1(n4552), .A2(N340), .B1(N395), .B2(n4197), .ZN(n4195) );
  OAI221_X2 U2388 ( .B1(n4191), .B2(n4387), .C1(n4557), .C2(n6012), .A(n4198), 
        .ZN(N715) );
  AOI22_X2 U2389 ( .A1(n4552), .A2(opa_r1[51]), .B1(N394), .B2(n4197), .ZN(
        n4198) );
  OAI221_X2 U2390 ( .B1(n4191), .B2(n4386), .C1(n4557), .C2(n6013), .A(n4199), 
        .ZN(N714) );
  AOI22_X2 U2391 ( .A1(n4551), .A2(opa_r1[50]), .B1(N393), .B2(n4197), .ZN(
        n4199) );
  OAI221_X2 U2392 ( .B1(n4191), .B2(n4385), .C1(n4557), .C2(n6014), .A(n4200), 
        .ZN(N713) );
  AOI22_X2 U2393 ( .A1(n4552), .A2(opa_r1[49]), .B1(N392), .B2(n4197), .ZN(
        n4200) );
  OAI221_X2 U2394 ( .B1(n4191), .B2(n4496), .C1(n4557), .C2(n4380), .A(n4201), 
        .ZN(N712) );
  AOI22_X2 U2395 ( .A1(n4550), .A2(opa_r1[48]), .B1(N391), .B2(n4197), .ZN(
        n4201) );
  AOI22_X2 U2397 ( .A1(n4552), .A2(opa_r1[47]), .B1(N390), .B2(n4197), .ZN(
        n4202) );
  AOI22_X2 U2399 ( .A1(n4552), .A2(opa_r1[46]), .B1(N389), .B2(n4197), .ZN(
        n4203) );
  NAND2_X2 U2400 ( .A1(n4190), .A2(n6312), .ZN(n4191) );
  AOI22_X2 U2450 ( .A1(sign_fasu), .A2(n4303), .B1(sign_mul), .B2(fpu_op_r2[1]), .ZN(n4190) );
  NAND4_X2 U2451 ( .A1(n4483), .A2(n4329), .A3(n4250), .A4(n4251), .ZN(N340)
         );
  NOR4_X2 U2452 ( .A1(n4252), .A2(opa_r1[57]), .A3(opa_r1[59]), .A4(opa_r1[58]), .ZN(n4251) );
  OAI221_X2 U2455 ( .B1(n6312), .B2(n4381), .C1(n4330), .C2(n3296), .A(n4253), 
        .ZN(N337) );
  NAND2_X2 U2456 ( .A1(exp_fasu[10]), .A2(n4254), .ZN(n4253) );
  OAI221_X2 U2457 ( .B1(n6312), .B2(n4484), .C1(n4384), .C2(n3296), .A(n4255), 
        .ZN(N336) );
  NAND2_X2 U2458 ( .A1(exp_fasu[9]), .A2(n4254), .ZN(n4255) );
  OAI221_X2 U2459 ( .B1(n6312), .B2(n4328), .C1(n4489), .C2(n3296), .A(n4256), 
        .ZN(N335) );
  NAND2_X2 U2460 ( .A1(exp_fasu[8]), .A2(n4254), .ZN(n4256) );
  OAI221_X2 U2461 ( .B1(n6312), .B2(n4336), .C1(n4534), .C2(n3296), .A(n4257), 
        .ZN(N334) );
  NAND2_X2 U2462 ( .A1(exp_fasu[7]), .A2(n4254), .ZN(n4257) );
  OAI221_X2 U2463 ( .B1(n6312), .B2(n4335), .C1(n4536), .C2(n3296), .A(n4258), 
        .ZN(N333) );
  NAND2_X2 U2464 ( .A1(exp_fasu[6]), .A2(n4254), .ZN(n4258) );
  OAI221_X2 U2465 ( .B1(n6312), .B2(n4334), .C1(n4535), .C2(n3296), .A(n4259), 
        .ZN(N332) );
  NAND2_X2 U2466 ( .A1(exp_fasu[5]), .A2(n4254), .ZN(n4259) );
  OAI221_X2 U2467 ( .B1(n6312), .B2(n4332), .C1(n4537), .C2(n3296), .A(n4260), 
        .ZN(N331) );
  NAND2_X2 U2468 ( .A1(exp_fasu[4]), .A2(n4254), .ZN(n4260) );
  OAI221_X2 U2469 ( .B1(n6312), .B2(n4331), .C1(n4538), .C2(n3296), .A(n4261), 
        .ZN(N330) );
  NAND2_X2 U2470 ( .A1(exp_fasu[3]), .A2(n4254), .ZN(n4261) );
  OAI221_X2 U2473 ( .B1(n4262), .B2(n4333), .C1(n4539), .C2(n4303), .A(n4263), 
        .ZN(N329) );
  NAND2_X2 U2474 ( .A1(exp_fasu[2]), .A2(n4254), .ZN(n4263) );
  OAI221_X2 U2475 ( .B1(n4262), .B2(n4329), .C1(n4487), .C2(n4303), .A(n4264), 
        .ZN(N328) );
  NAND2_X2 U2476 ( .A1(exp_fasu[1]), .A2(n4254), .ZN(n4264) );
  OAI221_X2 U2477 ( .B1(n4262), .B2(n4483), .C1(n4383), .C2(n4303), .A(n4265), 
        .ZN(N327) );
  NAND2_X2 U2478 ( .A1(exp_fasu[0]), .A2(n4254), .ZN(n4265) );
  NAND2_X2 U2480 ( .A1(fpu_op_r2[2]), .A2(fpu_op_r2[0]), .ZN(n4262) );
  OAI33_X1 U3364 ( .A1(n6464), .A2(n2506), .A3(n2507), .B1(n2508), .B2(n2509), 
        .B3(n2510), .ZN(n2505) );
  OAI33_X1 U3366 ( .A1(n2598), .A2(n6355), .A3(n6357), .B1(n2671), .B2(n6376), 
        .B3(n6378), .ZN(n2652) );
  OAI33_X1 U3367 ( .A1(n2642), .A2(fract_denorm[81]), .A3(n6384), .B1(n6335), 
        .B2(fract_denorm[73]), .B3(n6397), .ZN(n2678) );
  OAI33_X1 U3368 ( .A1(n6334), .A2(fract_denorm[65]), .A3(n6390), .B1(n6326), 
        .B2(fract_denorm[57]), .B3(n6371), .ZN(n2677) );
  OAI33_X1 U3369 ( .A1(n2632), .A2(n6438), .A3(n2680), .B1(n6332), .B2(n6431), 
        .B3(n2681), .ZN(n2676) );
  OAI33_X1 U3370 ( .A1(n2598), .A2(fract_denorm[97]), .A3(n6356), .B1(n2671), 
        .B2(fract_denorm[89]), .B3(n6377), .ZN(n2687) );
  OAI33_X1 U3371 ( .A1(n3090), .A2(fracta_mul[2]), .A3(fracta_mul[1]), .B1(
        n3248), .B2(fracta_mul[17]), .B3(n4362), .ZN(n3247) );
  OAI33_X1 U3372 ( .A1(n6295), .A2(fracta_mul[47]), .A3(n4477), .B1(n6293), 
        .B2(fracta_mul[43]), .B3(n4286), .ZN(n3250) );
  OAI33_X1 U3373 ( .A1(n4372), .A2(fracta_mul[15]), .A3(n6300), .B1(n4300), 
        .B2(fracta_mul[11]), .B3(n6302), .ZN(n3274) );
  OAI33_X1 U3374 ( .A1(n6293), .A2(n6297), .A3(n4478), .B1(n3284), .B2(n3288), 
        .B3(n4376), .ZN(n3227) );
  OAI33_X1 U3375 ( .A1(n6449), .A2(n3342), .A3(n4274), .B1(n3343), .B2(
        inf_mul_r), .B3(n3344), .ZN(N902) );
  OAI33_X1 U3376 ( .A1(n3343), .A2(inf_d), .A3(n3454), .B1(n3455), .B2(
        fpu_op_r3[2]), .B3(n3456), .ZN(N899) );
  OAI33_X1 U3377 ( .A1(n3473), .A2(n2422), .A3(n4452), .B1(n3474), .B2(n6466), 
        .B3(n3475), .ZN(n3472) );
  OAI33_X1 U3378 ( .A1(n3783), .A2(\u4/N6410 ), .A3(n4355), .B1(n4351), .B2(
        sign), .B3(n3784), .ZN(n3478) );
  DFF_X2 \opa_r_reg[63]  ( .D(opa[63]), .CK(clk), .Q(opa_r[63]), .QN(n4533) );
  DFF_X2 \opa_r_reg[62]  ( .D(opa[62]), .CK(clk), .Q(opa_r[62]), .QN(n4458) );
  DFF_X2 \opa_r_reg[61]  ( .D(opa[61]), .CK(clk), .Q(opa_r[61]), .QN(n4448) );
  DFF_X2 \opa_r_reg[60]  ( .D(opa[60]), .CK(clk), .Q(opa_r[60]), .QN(n4357) );
  DFF_X2 \opa_r_reg[59]  ( .D(opa[59]), .CK(clk), .Q(opa_r[59]), .QN(n4442) );
  DFF_X2 \opa_r_reg[58]  ( .D(opa[58]), .CK(clk), .Q(opa_r[58]), .QN(n4454) );
  DFF_X2 \opa_r_reg[57]  ( .D(opa[57]), .CK(clk), .Q(opa_r[57]), .QN(n4453) );
  DFF_X2 \opa_r_reg[56]  ( .D(opa[56]), .CK(clk), .Q(opa_r[56]), .QN(n4456) );
  DFF_X2 \opa_r_reg[55]  ( .D(opa[55]), .CK(clk), .Q(opa_r[55]), .QN(n4358) );
  DFF_X2 \opa_r_reg[54]  ( .D(opa[54]), .CK(clk), .Q(opa_r[54]), .QN(n4451) );
  DFF_X2 \opa_r_reg[53]  ( .D(opa[53]), .CK(clk), .Q(opa_r[53]), .QN(n4450) );
  DFF_X2 \opa_r_reg[52]  ( .D(opa[52]), .CK(clk), .Q(opa_r[52]), .QN(n4449) );
  DFF_X2 \opa_r_reg[51]  ( .D(opa[51]), .CK(clk), .Q(fracta_mul[51]), .QN(
        n4273) );
  DFF_X2 \opa_r_reg[50]  ( .D(opa[50]), .CK(clk), .Q(fracta_mul[50]), .QN(
        n4480) );
  DFF_X2 \opa_r_reg[49]  ( .D(opa[49]), .CK(clk), .Q(fracta_mul[49]) );
  DFF_X2 \opa_r_reg[48]  ( .D(opa[48]), .CK(clk), .Q(fracta_mul[48]) );
  DFF_X2 \opa_r_reg[47]  ( .D(opa[47]), .CK(clk), .Q(fracta_mul[47]) );
  DFF_X2 \opa_r_reg[46]  ( .D(opa[46]), .CK(clk), .Q(fracta_mul[46]), .QN(
        n4477) );
  DFF_X2 \opa_r_reg[45]  ( .D(opa[45]), .CK(clk), .Q(fracta_mul[45]), .QN(
        n4367) );
  DFF_X2 \opa_r_reg[44]  ( .D(opa[44]), .CK(clk), .Q(fracta_mul[44]), .QN(
        n4277) );
  DFF_X2 \opa_r_reg[43]  ( .D(opa[43]), .CK(clk), .Q(fracta_mul[43]) );
  DFF_X2 \opa_r_reg[42]  ( .D(opa[42]), .CK(clk), .Q(fracta_mul[42]), .QN(
        n4286) );
  DFF_X2 \opa_r_reg[41]  ( .D(opa[41]), .CK(clk), .Q(fracta_mul[41]), .QN(
        n4472) );
  DFF_X2 \opa_r_reg[40]  ( .D(opa[40]), .CK(clk), .Q(fracta_mul[40]) );
  DFF_X2 \opa_r_reg[39]  ( .D(opa[39]), .CK(clk), .Q(fracta_mul[39]), .QN(
        n4478) );
  DFF_X2 \opa_r_reg[38]  ( .D(opa[38]), .CK(clk), .Q(fracta_mul[38]), .QN(
        n4284) );
  DFF_X2 \opa_r_reg[37]  ( .D(opa[37]), .CK(clk), .Q(fracta_mul[37]), .QN(
        n4272) );
  DFF_X2 \opa_r_reg[36]  ( .D(opa[36]), .CK(clk), .Q(fracta_mul[36]), .QN(
        n4276) );
  DFF_X2 \opa_r_reg[35]  ( .D(opa[35]), .CK(clk), .Q(fracta_mul[35]), .QN(
        n4474) );
  DFF_X2 \opa_r_reg[34]  ( .D(opa[34]), .CK(clk), .Q(fracta_mul[34]) );
  DFF_X2 \opa_r_reg[33]  ( .D(opa[33]), .CK(clk), .Q(fracta_mul[33]) );
  DFF_X2 \opa_r_reg[32]  ( .D(opa[32]), .CK(clk), .Q(fracta_mul[32]), .QN(
        n4287) );
  DFF_X2 \opa_r_reg[31]  ( .D(opa[31]), .CK(clk), .Q(fracta_mul[31]), .QN(
        n4370) );
  DFF_X2 \opa_r_reg[30]  ( .D(opa[30]), .CK(clk), .Q(fracta_mul[30]), .QN(
        n4479) );
  DFF_X2 \opa_r_reg[29]  ( .D(opa[29]), .CK(clk), .Q(fracta_mul[29]), .QN(
        n4475) );
  DFF_X2 \opa_r_reg[28]  ( .D(opa[28]), .CK(clk), .Q(fracta_mul[28]), .QN(
        n4285) );
  DFF_X2 \opa_r_reg[27]  ( .D(opa[27]), .CK(clk), .Q(fracta_mul[27]), .QN(
        n4301) );
  DFF_X2 \opa_r_reg[26]  ( .D(opa[26]), .CK(clk), .Q(fracta_mul[26]) );
  DFF_X2 \opa_r_reg[25]  ( .D(opa[25]), .CK(clk), .Q(fracta_mul[25]), .QN(
        n4473) );
  DFF_X2 \opa_r_reg[24]  ( .D(opa[24]), .CK(clk), .Q(fracta_mul[24]) );
  DFF_X2 \opa_r_reg[23]  ( .D(opa[23]), .CK(clk), .Q(fracta_mul[23]) );
  DFF_X2 \opa_r_reg[22]  ( .D(opa[22]), .CK(clk), .Q(fracta_mul[22]), .QN(
        n4283) );
  DFF_X2 \opa_r_reg[21]  ( .D(opa[21]), .CK(clk), .Q(fracta_mul[21]), .QN(
        n4292) );
  DFF_X2 \opa_r_reg[20]  ( .D(opa[20]), .CK(clk), .Q(fracta_mul[20]), .QN(
        n4320) );
  DFF_X2 \opa_r_reg[19]  ( .D(opa[19]), .CK(clk), .Q(fracta_mul[19]) );
  DFF_X2 \opa_r_reg[18]  ( .D(opa[18]), .CK(clk), .Q(fracta_mul[18]), .QN(
        n4369) );
  DFF_X2 \opa_r_reg[17]  ( .D(opa[17]), .CK(clk), .Q(fracta_mul[17]), .QN(
        n4319) );
  DFF_X2 \opa_r_reg[16]  ( .D(opa[16]), .CK(clk), .Q(fracta_mul[16]), .QN(
        n4362) );
  DFF_X2 \opa_r_reg[15]  ( .D(opa[15]), .CK(clk), .Q(fracta_mul[15]), .QN(
        n4318) );
  DFF_X2 \opa_r_reg[14]  ( .D(opa[14]), .CK(clk), .Q(fracta_mul[14]), .QN(
        n4372) );
  DFF_X2 \opa_r_reg[13]  ( .D(opa[13]), .CK(clk), .Q(fracta_mul[13]), .QN(
        n4476) );
  DFF_X2 \opa_r_reg[12]  ( .D(opa[12]), .CK(clk), .Q(fracta_mul[12]), .QN(
        n4374) );
  DFF_X2 \opa_r_reg[11]  ( .D(opa[11]), .CK(clk), .Q(fracta_mul[11]), .QN(
        n4361) );
  DFF_X2 \opa_r_reg[10]  ( .D(opa[10]), .CK(clk), .Q(fracta_mul[10]), .QN(
        n4300) );
  DFF_X2 \opa_r_reg[9]  ( .D(opa[9]), .CK(clk), .Q(fracta_mul[9]), .QN(n4368)
         );
  DFF_X2 \opa_r_reg[8]  ( .D(opa[8]), .CK(clk), .Q(fracta_mul[8]), .QN(n4326)
         );
  DFF_X2 \opa_r_reg[7]  ( .D(opa[7]), .CK(clk), .Q(fracta_mul[7]), .QN(n4376)
         );
  DFF_X2 \opa_r_reg[6]  ( .D(opa[6]), .CK(clk), .Q(fracta_mul[6]), .QN(n4375)
         );
  DFF_X2 \opa_r_reg[5]  ( .D(opa[5]), .CK(clk), .Q(fracta_mul[5]), .QN(n4371)
         );
  DFF_X2 \opa_r_reg[4]  ( .D(opa[4]), .CK(clk), .Q(fracta_mul[4]) );
  DFF_X2 \opa_r_reg[3]  ( .D(opa[3]), .CK(clk), .Q(fracta_mul[3]), .QN(n4360)
         );
  DFF_X2 \opa_r_reg[2]  ( .D(opa[2]), .CK(clk), .Q(fracta_mul[2]) );
  DFF_X2 \opa_r_reg[1]  ( .D(opa[1]), .CK(clk), .Q(fracta_mul[1]), .QN(n4373)
         );
  DFF_X2 \opa_r_reg[0]  ( .D(opa[0]), .CK(clk), .Q(fracta_mul[0]), .QN(n4322)
         );
  DFF_X2 \opb_r_reg[63]  ( .D(opb[63]), .CK(clk), .Q(opb_r[63]) );
  DFF_X2 \opb_r_reg[62]  ( .D(opb[62]), .CK(clk), .Q(opb_r[62]), .QN(n4363) );
  DFF_X2 \opb_r_reg[61]  ( .D(opb[61]), .CK(clk), .Q(opb_r[61]) );
  DFF_X2 \opb_r_reg[60]  ( .D(opb[60]), .CK(clk), .Q(opb_r[60]) );
  DFF_X2 \opb_r_reg[59]  ( .D(opb[59]), .CK(clk), .Q(opb_r[59]), .QN(n4340) );
  DFF_X2 \opb_r_reg[58]  ( .D(opb[58]), .CK(clk), .Q(opb_r[58]), .QN(n4399) );
  DFF_X2 \opb_r_reg[57]  ( .D(opb[57]), .CK(clk), .Q(opb_r[57]), .QN(n4296) );
  DFF_X2 \opb_r_reg[56]  ( .D(opb[56]), .CK(clk), .Q(opb_r[56]), .QN(n4359) );
  DFF_X2 \opb_r_reg[55]  ( .D(opb[55]), .CK(clk), .Q(opb_r[55]), .QN(n4321) );
  DFF_X2 \opb_r_reg[54]  ( .D(opb[54]), .CK(clk), .Q(opb_r[54]), .QN(n4457) );
  DFF_X2 \opb_r_reg[53]  ( .D(opb[53]), .CK(clk), .Q(opb_r[53]), .QN(n4275) );
  DFF_X2 \opb_r_reg[52]  ( .D(opb[52]), .CK(clk), .Q(opb_r[52]), .QN(n4270) );
  DFF_X2 \opb_r_reg[51]  ( .D(opb[51]), .CK(clk), .Q(\u6/N51 ), .QN(n4459) );
  DFF_X2 \opb_r_reg[50]  ( .D(opb[50]), .CK(clk), .Q(\u6/N50 ) );
  DFF_X2 \opb_r_reg[49]  ( .D(opb[49]), .CK(clk), .Q(\u6/N49 ) );
  DFF_X2 \opb_r_reg[48]  ( .D(opb[48]), .CK(clk), .Q(\u6/N48 ) );
  DFF_X2 \opb_r_reg[47]  ( .D(opb[47]), .CK(clk), .Q(\u6/N47 ) );
  DFF_X2 \opb_r_reg[46]  ( .D(opb[46]), .CK(clk), .Q(\u6/N46 ) );
  DFF_X2 \opb_r_reg[45]  ( .D(opb[45]), .CK(clk), .Q(\u6/N45 ) );
  DFF_X2 \opb_r_reg[44]  ( .D(opb[44]), .CK(clk), .Q(\u6/N44 ), .QN(n4468) );
  DFF_X2 \opb_r_reg[43]  ( .D(opb[43]), .CK(clk), .Q(\u6/N43 ) );
  DFF_X2 \opb_r_reg[42]  ( .D(opb[42]), .CK(clk), .Q(\u6/N42 ), .QN(n4467) );
  DFF_X2 \opb_r_reg[41]  ( .D(opb[41]), .CK(clk), .Q(\u6/N41 ) );
  DFF_X2 \opb_r_reg[40]  ( .D(opb[40]), .CK(clk), .Q(\u6/N40 ) );
  DFF_X2 \opb_r_reg[39]  ( .D(opb[39]), .CK(clk), .Q(\u6/N39 ) );
  DFF_X2 \opb_r_reg[38]  ( .D(opb[38]), .CK(clk), .Q(\u6/N38 ), .QN(n4465) );
  DFF_X2 \opb_r_reg[37]  ( .D(opb[37]), .CK(clk), .Q(\u6/N37 ), .QN(n4471) );
  DFF_X2 \opb_r_reg[36]  ( .D(opb[36]), .CK(clk), .Q(\u6/N36 ), .QN(n4470) );
  DFF_X2 \opb_r_reg[35]  ( .D(opb[35]), .CK(clk), .Q(\u6/N35 ) );
  DFF_X2 \opb_r_reg[34]  ( .D(opb[34]), .CK(clk), .Q(\u6/N34 ) );
  DFF_X2 \opb_r_reg[33]  ( .D(opb[33]), .CK(clk), .Q(\u6/N33 ) );
  DFF_X2 \opb_r_reg[32]  ( .D(opb[32]), .CK(clk), .Q(\u6/N32 ), .QN(n4464) );
  DFF_X2 \opb_r_reg[31]  ( .D(opb[31]), .CK(clk), .Q(\u6/N31 ) );
  DFF_X2 \opb_r_reg[30]  ( .D(opb[30]), .CK(clk), .Q(\u6/N30 ) );
  DFF_X2 \opb_r_reg[29]  ( .D(opb[29]), .CK(clk), .Q(\u6/N29 ) );
  DFF_X2 \opb_r_reg[28]  ( .D(opb[28]), .CK(clk), .Q(\u6/N28 ), .QN(n4469) );
  DFF_X2 \opb_r_reg[27]  ( .D(opb[27]), .CK(clk), .Q(\u6/N27 ), .QN(n4466) );
  DFF_X2 \opb_r_reg[26]  ( .D(opb[26]), .CK(clk), .Q(\u6/N26 ) );
  DFF_X2 \opb_r_reg[25]  ( .D(opb[25]), .CK(clk), .Q(\u6/N25 ) );
  DFF_X2 \opb_r_reg[24]  ( .D(opb[24]), .CK(clk), .Q(\u6/N24 ) );
  DFF_X2 \opb_r_reg[23]  ( .D(opb[23]), .CK(clk), .Q(\u6/N23 ) );
  DFF_X2 \opb_r_reg[22]  ( .D(opb[22]), .CK(clk), .Q(\u6/N22 ), .QN(n4462) );
  DFF_X2 \opb_r_reg[21]  ( .D(opb[21]), .CK(clk), .Q(\u6/N21 ), .QN(n4325) );
  DFF_X2 \opb_r_reg[20]  ( .D(opb[20]), .CK(clk), .Q(\u6/N20 ), .QN(n4366) );
  DFF_X2 \opb_r_reg[19]  ( .D(opb[19]), .CK(clk), .Q(\u6/N19 ) );
  DFF_X2 \opb_r_reg[18]  ( .D(opb[18]), .CK(clk), .Q(\u6/N18 ) );
  DFF_X2 \opb_r_reg[17]  ( .D(opb[17]), .CK(clk), .Q(\u6/N17 ), .QN(n4461) );
  DFF_X2 \opb_r_reg[16]  ( .D(opb[16]), .CK(clk), .Q(\u6/N16 ), .QN(n4324) );
  DFF_X2 \opb_r_reg[15]  ( .D(opb[15]), .CK(clk), .Q(\u6/N15 ), .QN(n4365) );
  DFF_X2 \opb_r_reg[14]  ( .D(opb[14]), .CK(clk), .Q(\u6/N14 ) );
  DFF_X2 \opb_r_reg[13]  ( .D(opb[13]), .CK(clk), .Q(\u6/N13 ) );
  DFF_X2 \opb_r_reg[12]  ( .D(opb[12]), .CK(clk), .Q(\u6/N12 ) );
  DFF_X2 \opb_r_reg[11]  ( .D(opb[11]), .CK(clk), .Q(\u6/N11 ), .QN(n4460) );
  DFF_X2 \opb_r_reg[10]  ( .D(opb[10]), .CK(clk), .Q(\u6/N10 ), .QN(n4323) );
  DFF_X2 \opb_r_reg[9]  ( .D(opb[9]), .CK(clk), .Q(\u6/N9 ) );
  DFF_X2 \opb_r_reg[8]  ( .D(opb[8]), .CK(clk), .Q(\u6/N8 ) );
  DFF_X2 \opb_r_reg[7]  ( .D(opb[7]), .CK(clk), .Q(\u6/N7 ) );
  DFF_X2 \opb_r_reg[6]  ( .D(opb[6]), .CK(clk), .Q(\u6/N6 ) );
  DFF_X2 \opb_r_reg[5]  ( .D(opb[5]), .CK(clk), .Q(\u6/N5 ) );
  DFF_X2 \opb_r_reg[4]  ( .D(opb[4]), .CK(clk), .Q(\u6/N4 ) );
  DFF_X2 \opb_r_reg[3]  ( .D(opb[3]), .CK(clk), .Q(\u6/N3 ), .QN(n4463) );
  DFF_X2 \opb_r_reg[2]  ( .D(opb[2]), .CK(clk), .Q(\u6/N2 ) );
  DFF_X2 \opb_r_reg[1]  ( .D(opb[1]), .CK(clk), .Q(\u6/N1 ) );
  DFF_X2 \opb_r_reg[0]  ( .D(opb[0]), .CK(clk), .Q(\u6/N0 ), .QN(n4364) );
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  DFF_X2 \rmode_r1_reg[1]  ( .D(rmode[1]), .CK(clk), .Q(rmode_r1[1]) );
  DFF_X2 \rmode_r1_reg[0]  ( .D(rmode[0]), .CK(clk), .Q(rmode_r1[0]) );
  DFF_X2 \rmode_r2_reg[1]  ( .D(rmode_r1[1]), .CK(clk), .Q(rmode_r2[1]) );
  DFF_X2 \rmode_r2_reg[0]  ( .D(rmode_r1[0]), .CK(clk), .Q(rmode_r2[0]) );
  DFF_X2 \rmode_r3_reg[1]  ( .D(rmode_r2[1]), .CK(clk), .Q(rmode_r3[1]), .QN(
<<<<<<< HEAD
        n1768) );
  DFF_X2 \rmode_r3_reg[0]  ( .D(rmode_r2[0]), .CK(clk), .Q(rmode_r3[0]), .QN(
        n1614) );
  DFF_X2 \fpu_op_r1_reg[2]  ( .D(fpu_op[2]), .CK(clk), .Q(fpu_op_r1[2]), .QN(
        n3100) );
  DFF_X2 \fpu_op_r1_reg[1]  ( .D(fpu_op[1]), .CK(clk), .Q(fpu_op_r1[1]) );
  DFF_X2 \fpu_op_r1_reg[0]  ( .D(fpu_op[0]), .CK(clk), .Q(fpu_op_r1[0]), .QN(
        n3317) );
  DFF_X2 \fpu_op_r2_reg[2]  ( .D(fpu_op_r1[2]), .CK(clk), .Q(fpu_op_r2[2]), 
        .QN(n3099) );
  DFF_X2 \fpu_op_r2_reg[1]  ( .D(fpu_op_r1[1]), .CK(clk), .Q(fpu_op_r2[1]), 
        .QN(n3098) );
  DFF_X2 \fpu_op_r2_reg[0]  ( .D(fpu_op_r1[0]), .CK(clk), .Q(fpu_op_r2[0]), 
        .QN(n3097) );
  DFF_X2 \fpu_op_r3_reg[2]  ( .D(fpu_op_r2[2]), .CK(clk), .Q(net86090), .QN(
        net11677) );
  DFF_X2 \fpu_op_r3_reg[1]  ( .D(fpu_op_r2[1]), .CK(clk), .Q(net86006), .QN(
        net11676) );
  DFF_X2 \fpu_op_r3_reg[0]  ( .D(fpu_op_r2[0]), .CK(clk), .Q(net88695), .QN(
        net11675) );
  DFF_X2 \div_opa_ldz_r1_reg[3]  ( .D(N34), .CK(clk), .Q(div_opa_ldz_r1[3]) );
  DFF_X2 \div_opa_ldz_r1_reg[2]  ( .D(N44), .CK(clk), .Q(div_opa_ldz_r1[2]) );
  DFF_X2 \div_opa_ldz_r1_reg[1]  ( .D(N56), .CK(clk), .Q(div_opa_ldz_r1[1]) );
  DFF_X2 \div_opa_ldz_r1_reg[0]  ( .D(N65), .CK(clk), .Q(div_opa_ldz_r1[0]) );
  DFF_X2 \div_opa_ldz_r2_reg[3]  ( .D(div_opa_ldz_r1[3]), .CK(clk), .Q(
        div_opa_ldz_r2[3]), .QN(n1663) );
  DFF_X2 \div_opa_ldz_r2_reg[2]  ( .D(div_opa_ldz_r1[2]), .CK(clk), .Q(
        div_opa_ldz_r2[2]), .QN(n3096) );
  DFF_X2 \div_opa_ldz_r2_reg[1]  ( .D(div_opa_ldz_r1[1]), .CK(clk), .Q(
        div_opa_ldz_r2[1]), .QN(net11671) );
  DFF_X2 \div_opa_ldz_r2_reg[0]  ( .D(div_opa_ldz_r1[0]), .CK(clk), .Q(
        div_opa_ldz_r2[0]), .QN(net11670) );
  DFF_X2 \opa_r1_reg[14]  ( .D(opa_r[14]), .CK(clk), .QN(n1635) );
  DFF_X2 \opa_r1_reg[13]  ( .D(opa_r[13]), .CK(clk), .QN(n1636) );
  DFF_X2 \opa_r1_reg[12]  ( .D(opa_r[12]), .CK(clk), .QN(n1637) );
  DFF_X2 \opa_r1_reg[11]  ( .D(opa_r[11]), .CK(clk), .Q(opa_r1[11]), .QN(n1672) );
  DFF_X2 \opa_r1_reg[10]  ( .D(opa_r[10]), .CK(clk), .Q(opa_r1[10]), .QN(n1673) );
  DFF_X2 \opa_r1_reg[9]  ( .D(fracta_mul[9]), .CK(clk), .QN(n1624) );
  DFF_X2 \opa_r1_reg[8]  ( .D(fracta_mul[8]), .CK(clk), .QN(n1625) );
  DFF_X2 \opa_r1_reg[7]  ( .D(fracta_mul[7]), .CK(clk), .QN(n1626) );
  DFF_X2 \opa_r1_reg[6]  ( .D(fracta_mul[6]), .CK(clk), .QN(n1627) );
  DFF_X2 \opa_r1_reg[5]  ( .D(fracta_mul[5]), .CK(clk), .Q(opa_r1[5]), .QN(
        n1678) );
  DFF_X2 \opa_r1_reg[4]  ( .D(fracta_mul[4]), .CK(clk), .Q(opa_r1[4]), .QN(
        n1679) );
  DFF_X2 \opa_r1_reg[3]  ( .D(fracta_mul[3]), .CK(clk), .QN(n1674) );
  DFF_X2 \opa_r1_reg[2]  ( .D(fracta_mul[2]), .CK(clk), .QN(n1675) );
  DFF_X2 \opa_r1_reg[1]  ( .D(fracta_mul[1]), .CK(clk), .QN(n1676) );
  DFF_X2 \opa_r1_reg[0]  ( .D(fracta_mul[0]), .CK(clk), .Q(N106), .QN(n1680)
         );
  DFF_X2 opas_r1_reg ( .D(opa_r[15]), .CK(clk), .Q(opas_r1) );
  DFF_X2 opas_r2_reg ( .D(opas_r1), .CK(clk), .Q(opas_r2), .QN(n1608) );
  DFF_X2 \u0/fractb_00_reg  ( .D(n3316), .CK(clk), .QN(n3095) );
  DFF_X2 \u0/fracta_00_reg  ( .D(n3314), .CK(clk), .QN(n3094) );
  DFF_X2 \u0/expb_00_reg  ( .D(n3013), .CK(clk), .Q(\u0/expb_00 ), .QN(n3093)
         );
  DFF_X2 \u0/opb_dn_reg  ( .D(\u0/expb_00 ), .CK(clk), .Q(opb_dn), .QN(
        net85974) );
  DFF_X2 \u0/opb_00_reg  ( .D(\u0/N17 ), .CK(clk), .Q(opb_00), .QN(n1570) );
  DFF_X2 \u0/expa_00_reg  ( .D(n3012), .CK(clk), .Q(\u0/expa_00 ), .QN(n3092)
         );
  DFF_X2 \u0/opa_dn_reg  ( .D(\u0/expa_00 ), .CK(clk), .Q(opa_dn), .QN(n1641)
         );
  DFF_X2 \u0/opa_00_reg  ( .D(\u0/N16 ), .CK(clk), .Q(opa_00), .QN(n1615) );
  DFF_X2 \u0/opb_nan_reg  ( .D(\u0/N11 ), .CK(clk), .Q(opb_nan), .QN(n1684) );
  DFF_X2 \u0/opa_nan_reg  ( .D(\u0/N10 ), .CK(clk), .Q(opa_nan), .QN(n1681) );
  DFF_X2 opa_nan_r_reg ( .D(N291), .CK(clk), .QN(n3091) );
  DFF_X2 \u0/snan_r_b_reg  ( .D(\u0/N5 ), .CK(clk), .QN(n3090) );
  DFF_X2 \u0/qnan_r_b_reg  ( .D(\u6/N9 ), .CK(clk), .QN(n3089) );
  DFF_X2 \u0/snan_r_a_reg  ( .D(\u0/N4 ), .CK(clk), .QN(n3088) );
  DFF_X2 \u0/qnan_r_a_reg  ( .D(fracta_mul[9]), .CK(clk), .QN(n3087) );
  DFF_X2 \u0/infb_f_r_reg  ( .D(n3316), .CK(clk), .Q(\u0/infb_f_r ) );
  DFF_X2 \u0/infa_f_r_reg  ( .D(n3314), .CK(clk), .Q(\u0/infa_f_r ) );
  DFF_X2 \u0/expb_ff_reg  ( .D(n3315), .CK(clk), .Q(\u0/expb_ff ), .QN(n1677)
         );
  DFF_X2 \u0/opb_inf_reg  ( .D(n3322), .CK(clk), .Q(opb_inf), .QN(n1595) );
  DFF_X2 \u0/expa_ff_reg  ( .D(n3312), .CK(clk), .Q(\u0/expa_ff ), .QN(n1591)
         );
  DFF_X2 \u0/snan_reg  ( .D(n3320), .CK(clk), .Q(snan_d), .QN(n3086) );
  DFF_X2 snan_reg ( .D(snan_d), .CK(clk), .Q(snan) );
  DFF_X2 \u0/qnan_reg  ( .D(n3321), .CK(clk), .QN(n3085) );
  DFF_X2 \u0/opa_inf_reg  ( .D(n3323), .CK(clk), .Q(opa_inf), .QN(n1572) );
  DFF_X2 div_by_zero_reg ( .D(N292), .CK(clk), .Q(div_by_zero) );
  DFF_X2 \u0/inf_reg  ( .D(\u0/N7 ), .CK(clk), .Q(n1576) );
  DFF_X2 \u0/ind_reg  ( .D(\u0/N6 ), .CK(clk), .Q(n1611) );
  DFF_X2 \u1/fasu_op_reg  ( .D(n3299), .CK(clk), .Q(fasu_op), .QN(n3084) );
  DFF_X2 fasu_op_r1_reg ( .D(fasu_op), .CK(clk), .Q(fasu_op_r1) );
  DFF_X2 fasu_op_r2_reg ( .D(fasu_op_r1), .CK(clk), .QN(net11627) );
  DFF_X2 qnan_reg ( .D(N283), .CK(clk), .Q(qnan) );
  DFF_X2 \u1/fracta_eq_fractb_reg  ( .D(\u1/N124 ), .CK(clk), .Q(
        \u1/fracta_eq_fractb ) );
  DFF_X2 \u1/fracta_lt_fractb_reg  ( .D(\u1/N123 ), .CK(clk), .Q(
        \u1/fracta_lt_fractb ), .QN(n1683) );
  DFF_X2 \u1/add_r_reg  ( .D(n3317), .CK(clk), .Q(\u1/add_r ) );
  DFF_X2 \u1/signb_r_reg  ( .D(opb_r[15]), .CK(clk), .QN(n1671) );
  DFF_X2 \u1/signa_r_reg  ( .D(opa_r[15]), .CK(clk), .Q(\u1/signa_r ), .QN(
        n1682) );
  DFF_X2 \u1/result_zero_sign_reg  ( .D(\u1/N122 ), .CK(clk), .Q(
        result_zero_sign_d) );
  DFF_X2 \u1/nan_sign_reg  ( .D(\u1/N133 ), .CK(clk), .Q(nan_sign_d) );
  DFF_X2 sign_fasu_r_reg ( .D(sign_fasu), .CK(clk), .Q(sign_fasu_r), .QN(n1685) );
  DFF_X2 \u1/fractb_out_reg[4]  ( .D(\u1/fractb_s [4]), .CK(clk), .Q(fractb[4]) );
  DFF_X2 \u1/fracta_out_reg[0]  ( .D(\u1/fracta_s [0]), .CK(clk), .Q(fracta[0]) );
  DFF_X2 \u1/fracta_out_reg[2]  ( .D(\u1/fracta_s [2]), .CK(clk), .Q(fracta[2]) );
  DFF_X2 \u1/fracta_out_reg[3]  ( .D(\u1/fracta_s [3]), .CK(clk), .Q(fracta[3]) );
  DFF_X2 \u1/fracta_out_reg[4]  ( .D(\u1/fracta_s [4]), .CK(clk), .Q(fracta[4]) );
  DFF_X2 \u1/fracta_out_reg[13]  ( .D(\u1/fracta_s [13]), .CK(clk), .Q(
        fracta[13]) );
  DFF_X2 \fract_out_q_reg[1]  ( .D(n3297), .CK(clk), .Q(fract_out_q[1]) );
  DFF_X2 \fract_out_q_reg[2]  ( .D(n3296), .CK(clk), .Q(fract_out_q[2]) );
  DFF_X2 \fract_out_q_reg[3]  ( .D(n3295), .CK(clk), .Q(fract_out_q[3]) );
  DFF_X2 \fract_out_q_reg[4]  ( .D(n3294), .CK(clk), .Q(fract_out_q[4]) );
  DFF_X2 \fract_out_q_reg[5]  ( .D(n3293), .CK(clk), .Q(fract_out_q[5]) );
  DFF_X2 \fract_out_q_reg[6]  ( .D(n3292), .CK(clk), .Q(fract_out_q[6]) );
  DFF_X2 \fract_out_q_reg[7]  ( .D(n3291), .CK(clk), .Q(fract_out_q[7]) );
  DFF_X2 \fract_out_q_reg[8]  ( .D(n3290), .CK(clk), .Q(fract_out_q[8]) );
  DFF_X2 \fract_out_q_reg[9]  ( .D(n3289), .CK(clk), .Q(fract_out_q[9]) );
  DFF_X2 \fract_out_q_reg[13]  ( .D(n3285), .CK(clk), .Q(fract_out_q[13]) );
  DFF_X2 \u1/exp_dn_out_reg[0]  ( .D(\u1/N35 ), .CK(clk), .QN(n3083) );
  DFF_X2 \u1/exp_dn_out_reg[1]  ( .D(\u1/N36 ), .CK(clk), .QN(n3082) );
  DFF_X2 \u1/exp_dn_out_reg[2]  ( .D(\u1/N37 ), .CK(clk), .QN(n3081) );
  DFF_X2 \u1/exp_dn_out_reg[3]  ( .D(\u1/N38 ), .CK(clk), .QN(n3080) );
  DFF_X2 \u1/exp_dn_out_reg[4]  ( .D(\u1/N39 ), .CK(clk), .QN(n3079) );
  DFF_X2 \u2/sign_exe_reg  ( .D(\u2/N73 ), .CK(clk), .Q(sign_exe) );
  DFF_X2 sign_exe_r_reg ( .D(sign_exe), .CK(clk), .Q(sign_exe_r), .QN(n1617)
         );
  DFF_X2 \u2/sign_reg  ( .D(\u2/sign_d ), .CK(clk), .Q(sign_mul) );
  DFF_X2 sign_mul_r_reg ( .D(sign_mul), .CK(clk), .Q(sign_mul_r), .QN(n1644)
         );
  DFF_X2 sign_reg ( .D(N216), .CK(clk), .Q(sign), .QN(net86016) );
  DFF_X2 \fract_i2f_reg[20]  ( .D(N195), .CK(clk), .Q(n1609) );
  DFF_X2 \fract_i2f_reg[18]  ( .D(N193), .CK(clk), .QN(n3078) );
  DFF_X2 \fract_i2f_reg[16]  ( .D(N191), .CK(clk), .QN(n3077) );
  DFF_X2 \fract_i2f_reg[14]  ( .D(N189), .CK(clk), .QN(n3076) );
  DFF_X2 \fract_i2f_reg[13]  ( .D(N188), .CK(clk), .QN(n3075) );
  DFF_X2 \fract_i2f_reg[10]  ( .D(N185), .CK(clk), .QN(net11582) );
  DFF_X2 \fract_i2f_reg[8]  ( .D(N183), .CK(clk), .QN(n3074) );
  DFF_X2 \fract_i2f_reg[7]  ( .D(N182), .CK(clk), .Q(\fract_i2f[7] ) );
  DFF_X2 \fract_i2f_reg[4]  ( .D(N179), .CK(clk), .QN(net11576) );
  DFF_X2 \fract_i2f_reg[3]  ( .D(n3281), .CK(clk), .QN(n3073) );
  DFF_X2 \fract_i2f_reg[1]  ( .D(n3283), .CK(clk), .QN(n3072) );
  DFF_X2 \u2/inf_reg  ( .D(\u2/N66 ), .CK(clk), .Q(inf_mul) );
  DFF_X2 inf_mul_r_reg ( .D(inf_mul), .CK(clk), .Q(n1631), .QN(n3071) );
  DFF_X2 \u2/underflow_reg[0]  ( .D(n1655), .CK(clk), .Q(underflow_fmul_d[0])
         );
  DFF_X2 \underflow_fmul_r_reg[0]  ( .D(underflow_fmul_d[0]), .CK(clk), .Q(
        n1612) );
=======
        n4351) );
  DFF_X2 \rmode_r3_reg[0]  ( .D(rmode_r2[0]), .CK(clk), .Q(rmode_r3[0]), .QN(
        n4441) );
  DFF_X2 \fpu_op_r1_reg[2]  ( .D(fpu_op[2]), .CK(clk), .Q(fpu_op_r1[2]), .QN(
        n4377) );
  DFF_X2 \fpu_op_r1_reg[1]  ( .D(fpu_op[1]), .CK(clk), .Q(fpu_op_r1[1]) );
  DFF_X2 \fpu_op_r1_reg[0]  ( .D(fpu_op[0]), .CK(clk), .Q(fpu_op_r1[0]), .QN(
        n4481) );
  DFF_X2 \fpu_op_r2_reg[2]  ( .D(fpu_op_r1[2]), .CK(clk), .Q(fpu_op_r2[2]) );
  DFF_X2 \fpu_op_r2_reg[1]  ( .D(fpu_op_r1[1]), .CK(clk), .Q(fpu_op_r2[1]), 
        .QN(n4303) );
  DFF_X2 \fpu_op_r2_reg[0]  ( .D(fpu_op_r1[0]), .CK(clk), .Q(fpu_op_r2[0]), 
        .QN(n4493) );
  DFF_X2 \fpu_op_r3_reg[2]  ( .D(fpu_op_r2[2]), .CK(clk), .Q(fpu_op_r3[2]), 
        .QN(n4291) );
  DFF_X2 \fpu_op_r3_reg[1]  ( .D(fpu_op_r2[1]), .CK(clk), .Q(fpu_op_r3[1]), 
        .QN(n4400) );
  DFF_X2 \fpu_op_r3_reg[0]  ( .D(fpu_op_r2[0]), .CK(clk), .Q(fpu_op_r3[0]), 
        .QN(n4274) );
  DFF_X2 \div_opa_ldz_r1_reg[4]  ( .D(div_opa_ldz_d[4]), .CK(clk), .Q(
        div_opa_ldz_r1[4]) );
  DFF_X2 \div_opa_ldz_r1_reg[3]  ( .D(div_opa_ldz_d[3]), .CK(clk), .Q(
        div_opa_ldz_r1[3]) );
  DFF_X2 \div_opa_ldz_r1_reg[2]  ( .D(div_opa_ldz_d[2]), .CK(clk), .Q(
        div_opa_ldz_r1[2]) );
  DFF_X2 \div_opa_ldz_r1_reg[1]  ( .D(div_opa_ldz_d[1]), .CK(clk), .Q(
        div_opa_ldz_r1[1]) );
  DFF_X2 \div_opa_ldz_r1_reg[0]  ( .D(div_opa_ldz_d[0]), .CK(clk), .Q(
        div_opa_ldz_r1[0]) );
  DFF_X2 \div_opa_ldz_r2_reg[4]  ( .D(div_opa_ldz_r1[4]), .CK(clk), .Q(
        div_opa_ldz_r2[4]), .QN(n4445) );
  DFF_X2 \div_opa_ldz_r2_reg[3]  ( .D(div_opa_ldz_r1[3]), .CK(clk), .Q(
        div_opa_ldz_r2[3]), .QN(n4443) );
  DFF_X2 \div_opa_ldz_r2_reg[2]  ( .D(div_opa_ldz_r1[2]), .CK(clk), .Q(
        div_opa_ldz_r2[2]), .QN(n4444) );
  DFF_X2 \div_opa_ldz_r2_reg[1]  ( .D(div_opa_ldz_r1[1]), .CK(clk), .Q(
        div_opa_ldz_r2[1]), .QN(n4446) );
  DFF_X2 \div_opa_ldz_r2_reg[0]  ( .D(div_opa_ldz_r1[0]), .CK(clk), .Q(
        div_opa_ldz_r2[0]), .QN(n4447) );
  DFF_X2 \opa_r1_reg[62]  ( .D(opa_r[62]), .CK(clk), .QN(n4381) );
  DFF_X2 \opa_r1_reg[61]  ( .D(opa_r[61]), .CK(clk), .QN(n4484) );
  DFF_X2 \opa_r1_reg[60]  ( .D(opa_r[60]), .CK(clk), .QN(n4328) );
  DFF_X2 \opa_r1_reg[59]  ( .D(opa_r[59]), .CK(clk), .Q(opa_r1[59]), .QN(n4336) );
  DFF_X2 \opa_r1_reg[58]  ( .D(opa_r[58]), .CK(clk), .Q(opa_r1[58]), .QN(n4335) );
  DFF_X2 \opa_r1_reg[57]  ( .D(opa_r[57]), .CK(clk), .Q(opa_r1[57]), .QN(n4334) );
  DFF_X2 \opa_r1_reg[56]  ( .D(opa_r[56]), .CK(clk), .Q(opa_r1[56]), .QN(n4332) );
  DFF_X2 \opa_r1_reg[55]  ( .D(opa_r[55]), .CK(clk), .Q(opa_r1[55]), .QN(n4331) );
  DFF_X2 \opa_r1_reg[54]  ( .D(opa_r[54]), .CK(clk), .Q(opa_r1[54]), .QN(n4333) );
  DFF_X2 \opa_r1_reg[53]  ( .D(opa_r[53]), .CK(clk), .Q(opa_r1[53]), .QN(n4329) );
  DFF_X2 \opa_r1_reg[52]  ( .D(opa_r[52]), .CK(clk), .Q(opa_r1[52]), .QN(n4483) );
  DFF_X2 \opa_r1_reg[51]  ( .D(fracta_mul[51]), .CK(clk), .Q(opa_r1[51]), .QN(
        n4532) );
  DFF_X2 \opa_r1_reg[50]  ( .D(fracta_mul[50]), .CK(clk), .Q(opa_r1[50]), .QN(
        n4531) );
  DFF_X2 \opa_r1_reg[49]  ( .D(fracta_mul[49]), .CK(clk), .Q(opa_r1[49]), .QN(
        n4530) );
  DFF_X2 \opa_r1_reg[48]  ( .D(fracta_mul[48]), .CK(clk), .Q(opa_r1[48]), .QN(
        n4529) );
  DFF_X2 \opa_r1_reg[47]  ( .D(fracta_mul[47]), .CK(clk), .Q(opa_r1[47]), .QN(
        n4528) );
  DFF_X2 \opa_r1_reg[46]  ( .D(fracta_mul[46]), .CK(clk), .Q(opa_r1[46]), .QN(
        n4527) );
  DFF_X2 \opa_r1_reg[45]  ( .D(fracta_mul[45]), .CK(clk), .Q(opa_r1[45]), .QN(
        n4526) );
  DFF_X2 \opa_r1_reg[44]  ( .D(fracta_mul[44]), .CK(clk), .Q(opa_r1[44]), .QN(
        n4525) );
  DFF_X2 \opa_r1_reg[43]  ( .D(fracta_mul[43]), .CK(clk), .Q(opa_r1[43]), .QN(
        n4524) );
  DFF_X2 \opa_r1_reg[42]  ( .D(fracta_mul[42]), .CK(clk), .Q(opa_r1[42]), .QN(
        n4523) );
  DFF_X2 \opa_r1_reg[41]  ( .D(fracta_mul[41]), .CK(clk), .Q(opa_r1[41]), .QN(
        n4522) );
  DFF_X2 \opa_r1_reg[40]  ( .D(fracta_mul[40]), .CK(clk), .Q(opa_r1[40]), .QN(
        n4521) );
  DFF_X2 \opa_r1_reg[39]  ( .D(fracta_mul[39]), .CK(clk), .Q(opa_r1[39]), .QN(
        n4520) );
  DFF_X2 \opa_r1_reg[38]  ( .D(fracta_mul[38]), .CK(clk), .Q(opa_r1[38]), .QN(
        n4519) );
  DFF_X2 \opa_r1_reg[37]  ( .D(fracta_mul[37]), .CK(clk), .Q(opa_r1[37]), .QN(
        n4518) );
  DFF_X2 \opa_r1_reg[36]  ( .D(fracta_mul[36]), .CK(clk), .Q(opa_r1[36]), .QN(
        n4517) );
  DFF_X2 \opa_r1_reg[35]  ( .D(fracta_mul[35]), .CK(clk), .Q(opa_r1[35]), .QN(
        n4516) );
  DFF_X2 \opa_r1_reg[34]  ( .D(fracta_mul[34]), .CK(clk), .Q(opa_r1[34]), .QN(
        n4515) );
  DFF_X2 \opa_r1_reg[33]  ( .D(fracta_mul[33]), .CK(clk), .Q(opa_r1[33]), .QN(
        n4514) );
  DFF_X2 \opa_r1_reg[32]  ( .D(fracta_mul[32]), .CK(clk), .Q(opa_r1[32]), .QN(
        n4513) );
  DFF_X2 \opa_r1_reg[31]  ( .D(fracta_mul[31]), .CK(clk), .Q(opa_r1[31]), .QN(
        n4512) );
  DFF_X2 \opa_r1_reg[30]  ( .D(fracta_mul[30]), .CK(clk), .Q(opa_r1[30]), .QN(
        n4511) );
  DFF_X2 \opa_r1_reg[29]  ( .D(fracta_mul[29]), .CK(clk), .Q(opa_r1[29]), .QN(
        n4510) );
  DFF_X2 \opa_r1_reg[28]  ( .D(fracta_mul[28]), .CK(clk), .Q(opa_r1[28]), .QN(
        n4509) );
  DFF_X2 \opa_r1_reg[27]  ( .D(fracta_mul[27]), .CK(clk), .Q(opa_r1[27]), .QN(
        n4508) );
  DFF_X2 \opa_r1_reg[26]  ( .D(fracta_mul[26]), .CK(clk), .Q(opa_r1[26]), .QN(
        n4507) );
  DFF_X2 \opa_r1_reg[25]  ( .D(fracta_mul[25]), .CK(clk), .Q(opa_r1[25]), .QN(
        n4506) );
  DFF_X2 \opa_r1_reg[24]  ( .D(fracta_mul[24]), .CK(clk), .Q(opa_r1[24]), .QN(
        n4505) );
  DFF_X2 \opa_r1_reg[23]  ( .D(fracta_mul[23]), .CK(clk), .Q(opa_r1[23]), .QN(
        n4504) );
  DFF_X2 \opa_r1_reg[22]  ( .D(fracta_mul[22]), .CK(clk), .Q(opa_r1[22]), .QN(
        n4503) );
  DFF_X2 \opa_r1_reg[21]  ( .D(fracta_mul[21]), .CK(clk), .Q(opa_r1[21]), .QN(
        n4502) );
  DFF_X2 \opa_r1_reg[20]  ( .D(fracta_mul[20]), .CK(clk), .Q(opa_r1[20]), .QN(
        n4501) );
  DFF_X2 \opa_r1_reg[19]  ( .D(fracta_mul[19]), .CK(clk), .Q(opa_r1[19]), .QN(
        n4500) );
  DFF_X2 \opa_r1_reg[18]  ( .D(fracta_mul[18]), .CK(clk), .Q(opa_r1[18]), .QN(
        n4499) );
  DFF_X2 \opa_r1_reg[17]  ( .D(fracta_mul[17]), .CK(clk), .Q(opa_r1[17]), .QN(
        n4498) );
  DFF_X2 \opa_r1_reg[16]  ( .D(fracta_mul[16]), .CK(clk), .Q(opa_r1[16]), .QN(
        n4497) );
  DFF_X2 \opa_r1_reg[15]  ( .D(fracta_mul[15]), .CK(clk), .Q(opa_r1[15]), .QN(
        n4397) );
  DFF_X2 \opa_r1_reg[14]  ( .D(fracta_mul[14]), .CK(clk), .Q(opa_r1[14]), .QN(
        n4396) );
  DFF_X2 \opa_r1_reg[13]  ( .D(fracta_mul[13]), .CK(clk), .Q(opa_r1[13]), .QN(
        n4395) );
  DFF_X2 \opa_r1_reg[12]  ( .D(fracta_mul[12]), .CK(clk), .Q(opa_r1[12]), .QN(
        n4394) );
  DFF_X2 \opa_r1_reg[11]  ( .D(fracta_mul[11]), .CK(clk), .Q(opa_r1[11]), .QN(
        n4393) );
  DFF_X2 \opa_r1_reg[10]  ( .D(fracta_mul[10]), .CK(clk), .Q(opa_r1[10]), .QN(
        n4392) );
  DFF_X2 \opa_r1_reg[9]  ( .D(fracta_mul[9]), .CK(clk), .Q(opa_r1[9]), .QN(
        n4391) );
  DFF_X2 \opa_r1_reg[8]  ( .D(fracta_mul[8]), .CK(clk), .Q(opa_r1[8]), .QN(
        n4390) );
  DFF_X2 \opa_r1_reg[7]  ( .D(fracta_mul[7]), .CK(clk), .Q(opa_r1[7]), .QN(
        n4389) );
  DFF_X2 \opa_r1_reg[6]  ( .D(fracta_mul[6]), .CK(clk), .Q(opa_r1[6]), .QN(
        n4388) );
  DFF_X2 \opa_r1_reg[5]  ( .D(fracta_mul[5]), .CK(clk), .Q(opa_r1[5]), .QN(
        n4387) );
  DFF_X2 \opa_r1_reg[4]  ( .D(fracta_mul[4]), .CK(clk), .Q(opa_r1[4]), .QN(
        n4386) );
  DFF_X2 \opa_r1_reg[3]  ( .D(fracta_mul[3]), .CK(clk), .Q(opa_r1[3]), .QN(
        n4385) );
  DFF_X2 \opa_r1_reg[2]  ( .D(fracta_mul[2]), .CK(clk), .Q(opa_r1[2]), .QN(
        n4496) );
  DFF_X2 \opa_r1_reg[1]  ( .D(fracta_mul[1]), .CK(clk), .Q(opa_r1[1]), .QN(
        n4488) );
  DFF_X2 \opa_r1_reg[0]  ( .D(fracta_mul[0]), .CK(clk), .Q(opa_r1[0]), .QN(
        n4380) );
  DFF_X2 opas_r1_reg ( .D(opa_r[63]), .CK(clk), .Q(opas_r1) );
  DFF_X2 opas_r2_reg ( .D(opas_r1), .CK(clk), .Q(opas_r2) );
  DFF_X2 \u0/fractb_00_reg  ( .D(n4268), .CK(clk), .Q(\u0/fractb_00 ) );
  DFF_X2 \u0/fracta_00_reg  ( .D(n4267), .CK(clk), .Q(\u0/fracta_00 ) );
  DFF_X2 \u0/expb_00_reg  ( .D(n6303), .CK(clk), .Q(\u0/expb_00 ) );
  DFF_X2 \u0/opb_dn_reg  ( .D(\u0/expb_00 ), .CK(clk), .Q(opb_dn), .QN(n4269)
         );
  DFF_X2 \u0/opb_00_reg  ( .D(\u0/N17 ), .CK(clk), .Q(opb_00) );
  DFF_X2 \u0/expa_00_reg  ( .D(n4601), .CK(clk), .Q(\u0/expa_00 ) );
  DFF_X2 \u0/opa_dn_reg  ( .D(\u0/expa_00 ), .CK(clk), .QN(n4271) );
  DFF_X2 \u0/opa_00_reg  ( .D(\u0/N16 ), .CK(clk), .Q(opa_00), .QN(n4486) );
  DFF_X2 \u0/opb_nan_reg  ( .D(\u0/N11 ), .CK(clk), .Q(opb_nan), .QN(n4492) );
  DFF_X2 \u0/opa_nan_reg  ( .D(\u0/N10 ), .CK(clk), .Q(opa_nan) );
  DFF_X2 opa_nan_r_reg ( .D(N912), .CK(clk), .Q(opa_nan_r) );
  DFF_X2 \u0/snan_r_b_reg  ( .D(\u0/N5 ), .CK(clk), .Q(\u0/snan_r_b ) );
  DFF_X2 \u0/qnan_r_b_reg  ( .D(\u6/N51 ), .CK(clk), .Q(\u0/qnan_r_b ) );
  DFF_X2 \u0/snan_r_a_reg  ( .D(\u0/N4 ), .CK(clk), .Q(\u0/snan_r_a ) );
  DFF_X2 \u0/qnan_r_a_reg  ( .D(fracta_mul[51]), .CK(clk), .Q(\u0/qnan_r_a )
         );
  DFF_X2 \u0/infb_f_r_reg  ( .D(n4268), .CK(clk), .Q(\u0/infb_f_r ) );
  DFF_X2 \u0/infa_f_r_reg  ( .D(n4267), .CK(clk), .Q(\u0/infa_f_r ) );
  DFF_X2 \u0/expb_ff_reg  ( .D(n6304), .CK(clk), .Q(\u0/expb_ff ) );
  DFF_X2 \u0/opb_inf_reg  ( .D(n6452), .CK(clk), .Q(opb_inf), .QN(n4327) );
  DFF_X2 \u0/expa_ff_reg  ( .D(n6276), .CK(clk), .Q(\u0/expa_ff ) );
  DFF_X2 \u0/snan_reg  ( .D(n6450), .CK(clk), .Q(snan_d) );
  DFF_X2 snan_reg ( .D(snan_d), .CK(clk), .Q(snan) );
  DFF_X2 \u0/qnan_reg  ( .D(n6451), .CK(clk), .Q(qnan_d) );
  DFF_X2 \u0/opa_inf_reg  ( .D(n6453), .CK(clk), .Q(opa_inf), .QN(n4382) );
  DFF_X2 div_by_zero_reg ( .D(N913), .CK(clk), .Q(div_by_zero) );
  DFF_X2 \u0/inf_reg  ( .D(\u0/N7 ), .CK(clk), .Q(inf_d) );
  DFF_X2 \u0/ind_reg  ( .D(\u0/N6 ), .CK(clk), .Q(ind_d) );
  DFF_X2 \u1/fasu_op_reg  ( .D(\u1/N232 ), .CK(clk), .Q(fasu_op), .QN(n4305)
         );
  DFF_X2 fasu_op_r1_reg ( .D(n4660), .CK(clk), .Q(fasu_op_r1) );
  DFF_X2 fasu_op_r2_reg ( .D(fasu_op_r1), .CK(clk), .Q(fasu_op_r2), .QN(n4494)
         );
  DFF_X2 qnan_reg ( .D(N904), .CK(clk), .Q(qnan) );
  DFF_X2 \u1/fracta_eq_fractb_reg  ( .D(\u1/N220 ), .CK(clk), .Q(
        \u1/fracta_eq_fractb ) );
  DFF_X2 \u1/fracta_lt_fractb_reg  ( .D(\u1/N219 ), .CK(clk), .Q(
        \u1/fracta_lt_fractb ) );
  DFF_X2 \u1/add_r_reg  ( .D(n4481), .CK(clk), .Q(\u1/add_r ) );
  DFF_X2 \u1/signb_r_reg  ( .D(opb_r[63]), .CK(clk), .Q(\u1/signb_r ), .QN(
        n4495) );
  DFF_X2 \u1/signa_r_reg  ( .D(opa_r[63]), .CK(clk), .Q(\u1/signa_r ), .QN(
        n4490) );
  DFF_X2 \u1/result_zero_sign_reg  ( .D(\u1/N218 ), .CK(clk), .Q(
        result_zero_sign_d) );
  DFF_X2 \u1/nan_sign_reg  ( .D(\u1/N229 ), .CK(clk), .Q(nan_sign_d) );
  DFF_X2 \u1/sign_reg  ( .D(\u1/sign_d ), .CK(clk), .Q(sign_fasu) );
  DFF_X2 sign_fasu_r_reg ( .D(sign_fasu), .CK(clk), .Q(sign_fasu_r) );
  DFF_X2 \u1/fractb_out_reg[0]  ( .D(\u1/fractb_s [0]), .CK(clk), .Q(fractb[0]) );
  DFF_X2 \u1/fractb_out_reg[1]  ( .D(\u1/fractb_s [1]), .CK(clk), .Q(fractb[1]) );
  DFF_X2 \u1/fractb_out_reg[2]  ( .D(\u1/fractb_s [2]), .CK(clk), .Q(fractb[2]) );
  DFF_X2 \u1/fractb_out_reg[3]  ( .D(\u1/fractb_s [3]), .CK(clk), .Q(fractb[3]) );
  DFF_X2 \u1/fractb_out_reg[4]  ( .D(\u1/fractb_s [4]), .CK(clk), .Q(fractb[4]) );
  DFF_X2 \u1/fractb_out_reg[5]  ( .D(\u1/fractb_s [5]), .CK(clk), .Q(fractb[5]) );
  DFF_X2 \u1/fractb_out_reg[6]  ( .D(\u1/fractb_s [6]), .CK(clk), .Q(fractb[6]) );
  DFF_X2 \u1/fractb_out_reg[7]  ( .D(\u1/fractb_s [7]), .CK(clk), .Q(fractb[7]) );
  DFF_X2 \u1/fractb_out_reg[8]  ( .D(\u1/fractb_s [8]), .CK(clk), .Q(fractb[8]) );
  DFF_X2 \u1/fractb_out_reg[9]  ( .D(\u1/fractb_s [9]), .CK(clk), .Q(fractb[9]) );
  DFF_X2 \u1/fractb_out_reg[10]  ( .D(\u1/fractb_s [10]), .CK(clk), .Q(
        fractb[10]) );
  DFF_X2 \u1/fractb_out_reg[11]  ( .D(\u1/fractb_s [11]), .CK(clk), .Q(
        fractb[11]) );
  DFF_X2 \u1/fractb_out_reg[12]  ( .D(\u1/fractb_s [12]), .CK(clk), .Q(
        fractb[12]) );
  DFF_X2 \u1/fractb_out_reg[13]  ( .D(\u1/fractb_s [13]), .CK(clk), .Q(
        fractb[13]) );
  DFF_X2 \u1/fractb_out_reg[14]  ( .D(\u1/fractb_s [14]), .CK(clk), .Q(
        fractb[14]) );
  DFF_X2 \u1/fractb_out_reg[15]  ( .D(\u1/fractb_s [15]), .CK(clk), .Q(
        fractb[15]) );
  DFF_X2 \u1/fractb_out_reg[16]  ( .D(\u1/fractb_s [16]), .CK(clk), .Q(
        fractb[16]) );
  DFF_X2 \u1/fractb_out_reg[17]  ( .D(\u1/fractb_s [17]), .CK(clk), .Q(
        fractb[17]) );
  DFF_X2 \u1/fractb_out_reg[18]  ( .D(\u1/fractb_s [18]), .CK(clk), .Q(
        fractb[18]) );
  DFF_X2 \u1/fractb_out_reg[19]  ( .D(\u1/fractb_s [19]), .CK(clk), .Q(
        fractb[19]) );
  DFF_X2 \u1/fractb_out_reg[20]  ( .D(\u1/fractb_s [20]), .CK(clk), .Q(
        fractb[20]) );
  DFF_X2 \u1/fractb_out_reg[21]  ( .D(\u1/fractb_s [21]), .CK(clk), .Q(
        fractb[21]) );
  DFF_X2 \u1/fractb_out_reg[22]  ( .D(\u1/fractb_s [22]), .CK(clk), .Q(
        fractb[22]) );
  DFF_X2 \u1/fractb_out_reg[23]  ( .D(\u1/fractb_s [23]), .CK(clk), .Q(
        fractb[23]) );
  DFF_X2 \u1/fractb_out_reg[24]  ( .D(\u1/fractb_s [24]), .CK(clk), .Q(
        fractb[24]) );
  DFF_X2 \u1/fractb_out_reg[25]  ( .D(\u1/fractb_s [25]), .CK(clk), .Q(
        fractb[25]) );
  DFF_X2 \u1/fractb_out_reg[26]  ( .D(\u1/fractb_s [26]), .CK(clk), .Q(
        fractb[26]) );
  DFF_X2 \u1/fractb_out_reg[27]  ( .D(\u1/fractb_s [27]), .CK(clk), .Q(
        fractb[27]) );
  DFF_X2 \u1/fractb_out_reg[28]  ( .D(\u1/fractb_s [28]), .CK(clk), .Q(
        fractb[28]) );
  DFF_X2 \u1/fractb_out_reg[29]  ( .D(\u1/fractb_s [29]), .CK(clk), .Q(
        fractb[29]) );
  DFF_X2 \u1/fractb_out_reg[30]  ( .D(\u1/fractb_s [30]), .CK(clk), .Q(
        fractb[30]) );
  DFF_X2 \u1/fractb_out_reg[31]  ( .D(\u1/fractb_s [31]), .CK(clk), .Q(
        fractb[31]) );
  DFF_X2 \u1/fractb_out_reg[32]  ( .D(\u1/fractb_s [32]), .CK(clk), .Q(
        fractb[32]) );
  DFF_X2 \u1/fractb_out_reg[33]  ( .D(\u1/fractb_s [33]), .CK(clk), .Q(
        fractb[33]) );
  DFF_X2 \u1/fractb_out_reg[34]  ( .D(\u1/fractb_s [34]), .CK(clk), .Q(
        fractb[34]) );
  DFF_X2 \u1/fractb_out_reg[35]  ( .D(\u1/fractb_s [35]), .CK(clk), .Q(
        fractb[35]) );
  DFF_X2 \u1/fractb_out_reg[36]  ( .D(\u1/fractb_s [36]), .CK(clk), .Q(
        fractb[36]) );
  DFF_X2 \u1/fractb_out_reg[37]  ( .D(\u1/fractb_s [37]), .CK(clk), .Q(
        fractb[37]) );
  DFF_X2 \u1/fractb_out_reg[38]  ( .D(\u1/fractb_s [38]), .CK(clk), .Q(
        fractb[38]) );
  DFF_X2 \u1/fractb_out_reg[39]  ( .D(\u1/fractb_s [39]), .CK(clk), .Q(
        fractb[39]) );
  DFF_X2 \u1/fractb_out_reg[40]  ( .D(\u1/fractb_s [40]), .CK(clk), .Q(
        fractb[40]) );
  DFF_X2 \u1/fractb_out_reg[41]  ( .D(\u1/fractb_s [41]), .CK(clk), .Q(
        fractb[41]) );
  DFF_X2 \u1/fractb_out_reg[42]  ( .D(\u1/fractb_s [42]), .CK(clk), .Q(
        fractb[42]) );
  DFF_X2 \u1/fractb_out_reg[43]  ( .D(\u1/fractb_s [43]), .CK(clk), .Q(
        fractb[43]) );
  DFF_X2 \u1/fractb_out_reg[44]  ( .D(\u1/fractb_s [44]), .CK(clk), .Q(
        fractb[44]) );
  DFF_X2 \u1/fractb_out_reg[45]  ( .D(\u1/fractb_s [45]), .CK(clk), .Q(
        fractb[45]) );
  DFF_X2 \u1/fractb_out_reg[46]  ( .D(\u1/fractb_s [46]), .CK(clk), .Q(
        fractb[46]) );
  DFF_X2 \u1/fractb_out_reg[47]  ( .D(\u1/fractb_s [47]), .CK(clk), .Q(
        fractb[47]) );
  DFF_X2 \u1/fractb_out_reg[48]  ( .D(\u1/fractb_s [48]), .CK(clk), .Q(
        fractb[48]) );
  DFF_X2 \u1/fractb_out_reg[49]  ( .D(\u1/fractb_s [49]), .CK(clk), .Q(
        fractb[49]) );
  DFF_X2 \u1/fractb_out_reg[50]  ( .D(\u1/fractb_s [50]), .CK(clk), .Q(
        fractb[50]) );
  DFF_X2 \u1/fractb_out_reg[51]  ( .D(\u1/fractb_s [51]), .CK(clk), .Q(
        fractb[51]) );
  DFF_X2 \u1/fractb_out_reg[52]  ( .D(\u1/fractb_s [52]), .CK(clk), .Q(
        fractb[52]) );
  DFF_X2 \u1/fractb_out_reg[53]  ( .D(\u1/fractb_s [53]), .CK(clk), .Q(
        fractb[53]) );
  DFF_X2 \u1/fractb_out_reg[54]  ( .D(\u1/fractb_s [54]), .CK(clk), .Q(
        fractb[54]) );
  DFF_X2 \u1/fractb_out_reg[55]  ( .D(\u1/fractb_s [55]), .CK(clk), .Q(
        fractb[55]) );
  DFF_X2 \u1/fracta_out_reg[0]  ( .D(\u1/fracta_s [0]), .CK(clk), .Q(fracta[0]) );
  DFF_X2 \u1/fracta_out_reg[1]  ( .D(\u1/fracta_s [1]), .CK(clk), .Q(fracta[1]) );
  DFF_X2 \u1/fracta_out_reg[2]  ( .D(\u1/fracta_s [2]), .CK(clk), .Q(fracta[2]) );
  DFF_X2 \u1/fracta_out_reg[3]  ( .D(\u1/fracta_s [3]), .CK(clk), .Q(fracta[3]) );
  DFF_X2 \u1/fracta_out_reg[4]  ( .D(\u1/fracta_s [4]), .CK(clk), .Q(fracta[4]) );
  DFF_X2 \u1/fracta_out_reg[5]  ( .D(\u1/fracta_s [5]), .CK(clk), .Q(fracta[5]) );
  DFF_X2 \u1/fracta_out_reg[6]  ( .D(\u1/fracta_s [6]), .CK(clk), .Q(fracta[6]) );
  DFF_X2 \u1/fracta_out_reg[7]  ( .D(\u1/fracta_s [7]), .CK(clk), .Q(fracta[7]) );
  DFF_X2 \u1/fracta_out_reg[8]  ( .D(\u1/fracta_s [8]), .CK(clk), .Q(fracta[8]) );
  DFF_X2 \u1/fracta_out_reg[9]  ( .D(\u1/fracta_s [9]), .CK(clk), .Q(fracta[9]) );
  DFF_X2 \u1/fracta_out_reg[10]  ( .D(\u1/fracta_s [10]), .CK(clk), .Q(
        fracta[10]) );
  DFF_X2 \u1/fracta_out_reg[11]  ( .D(\u1/fracta_s [11]), .CK(clk), .Q(
        fracta[11]) );
  DFF_X2 \u1/fracta_out_reg[12]  ( .D(\u1/fracta_s [12]), .CK(clk), .Q(
        fracta[12]) );
  DFF_X2 \u1/fracta_out_reg[13]  ( .D(\u1/fracta_s [13]), .CK(clk), .Q(
        fracta[13]) );
  DFF_X2 \u1/fracta_out_reg[14]  ( .D(\u1/fracta_s [14]), .CK(clk), .Q(
        fracta[14]) );
  DFF_X2 \u1/fracta_out_reg[15]  ( .D(\u1/fracta_s [15]), .CK(clk), .Q(
        fracta[15]) );
  DFF_X2 \u1/fracta_out_reg[16]  ( .D(\u1/fracta_s [16]), .CK(clk), .Q(
        fracta[16]) );
  DFF_X2 \u1/fracta_out_reg[17]  ( .D(\u1/fracta_s [17]), .CK(clk), .Q(
        fracta[17]) );
  DFF_X2 \u1/fracta_out_reg[18]  ( .D(\u1/fracta_s [18]), .CK(clk), .Q(
        fracta[18]) );
  DFF_X2 \u1/fracta_out_reg[19]  ( .D(\u1/fracta_s [19]), .CK(clk), .Q(
        fracta[19]) );
  DFF_X2 \u1/fracta_out_reg[20]  ( .D(\u1/fracta_s [20]), .CK(clk), .Q(
        fracta[20]) );
  DFF_X2 \u1/fracta_out_reg[21]  ( .D(\u1/fracta_s [21]), .CK(clk), .Q(
        fracta[21]) );
  DFF_X2 \u1/fracta_out_reg[22]  ( .D(\u1/fracta_s [22]), .CK(clk), .Q(
        fracta[22]) );
  DFF_X2 \u1/fracta_out_reg[23]  ( .D(\u1/fracta_s [23]), .CK(clk), .Q(
        fracta[23]) );
  DFF_X2 \u1/fracta_out_reg[24]  ( .D(\u1/fracta_s [24]), .CK(clk), .Q(
        fracta[24]) );
  DFF_X2 \u1/fracta_out_reg[25]  ( .D(\u1/fracta_s [25]), .CK(clk), .Q(
        fracta[25]) );
  DFF_X2 \u1/fracta_out_reg[26]  ( .D(\u1/fracta_s [26]), .CK(clk), .Q(
        fracta[26]) );
  DFF_X2 \u1/fracta_out_reg[27]  ( .D(\u1/fracta_s [27]), .CK(clk), .Q(
        fracta[27]) );
  DFF_X2 \u1/fracta_out_reg[28]  ( .D(\u1/fracta_s [28]), .CK(clk), .Q(
        fracta[28]) );
  DFF_X2 \u1/fracta_out_reg[29]  ( .D(\u1/fracta_s [29]), .CK(clk), .Q(
        fracta[29]) );
  DFF_X2 \u1/fracta_out_reg[30]  ( .D(\u1/fracta_s [30]), .CK(clk), .Q(
        fracta[30]) );
  DFF_X2 \u1/fracta_out_reg[31]  ( .D(\u1/fracta_s [31]), .CK(clk), .Q(
        fracta[31]) );
  DFF_X2 \u1/fracta_out_reg[32]  ( .D(\u1/fracta_s [32]), .CK(clk), .Q(
        fracta[32]) );
  DFF_X2 \u1/fracta_out_reg[33]  ( .D(\u1/fracta_s [33]), .CK(clk), .Q(
        fracta[33]) );
  DFF_X2 \u1/fracta_out_reg[34]  ( .D(\u1/fracta_s [34]), .CK(clk), .Q(
        fracta[34]) );
  DFF_X2 \u1/fracta_out_reg[35]  ( .D(\u1/fracta_s [35]), .CK(clk), .Q(
        fracta[35]) );
  DFF_X2 \u1/fracta_out_reg[36]  ( .D(\u1/fracta_s [36]), .CK(clk), .Q(
        fracta[36]) );
  DFF_X2 \u1/fracta_out_reg[37]  ( .D(\u1/fracta_s [37]), .CK(clk), .Q(
        fracta[37]) );
  DFF_X2 \u1/fracta_out_reg[38]  ( .D(\u1/fracta_s [38]), .CK(clk), .Q(
        fracta[38]) );
  DFF_X2 \u1/fracta_out_reg[39]  ( .D(\u1/fracta_s [39]), .CK(clk), .Q(
        fracta[39]) );
  DFF_X2 \u1/fracta_out_reg[40]  ( .D(\u1/fracta_s [40]), .CK(clk), .Q(
        fracta[40]) );
  DFF_X2 \u1/fracta_out_reg[41]  ( .D(\u1/fracta_s [41]), .CK(clk), .Q(
        fracta[41]) );
  DFF_X2 \u1/fracta_out_reg[42]  ( .D(\u1/fracta_s [42]), .CK(clk), .Q(
        fracta[42]) );
  DFF_X2 \u1/fracta_out_reg[43]  ( .D(\u1/fracta_s [43]), .CK(clk), .Q(
        fracta[43]) );
  DFF_X2 \u1/fracta_out_reg[44]  ( .D(\u1/fracta_s [44]), .CK(clk), .Q(
        fracta[44]) );
  DFF_X2 \u1/fracta_out_reg[45]  ( .D(\u1/fracta_s [45]), .CK(clk), .Q(
        fracta[45]) );
  DFF_X2 \u1/fracta_out_reg[46]  ( .D(\u1/fracta_s [46]), .CK(clk), .Q(
        fracta[46]) );
  DFF_X2 \u1/fracta_out_reg[47]  ( .D(\u1/fracta_s [47]), .CK(clk), .Q(
        fracta[47]) );
  DFF_X2 \u1/fracta_out_reg[48]  ( .D(\u1/fracta_s [48]), .CK(clk), .Q(
        fracta[48]) );
  DFF_X2 \u1/fracta_out_reg[49]  ( .D(\u1/fracta_s [49]), .CK(clk), .Q(
        fracta[49]) );
  DFF_X2 \u1/fracta_out_reg[50]  ( .D(\u1/fracta_s [50]), .CK(clk), .Q(
        fracta[50]) );
  DFF_X2 \u1/fracta_out_reg[51]  ( .D(\u1/fracta_s [51]), .CK(clk), .Q(
        fracta[51]) );
  DFF_X2 \u1/fracta_out_reg[52]  ( .D(\u1/fracta_s [52]), .CK(clk), .Q(
        fracta[52]) );
  DFF_X2 \u1/fracta_out_reg[53]  ( .D(\u1/fracta_s [53]), .CK(clk), .Q(
        fracta[53]) );
  DFF_X2 \u1/fracta_out_reg[54]  ( .D(\u1/fracta_s [54]), .CK(clk), .Q(
        fracta[54]) );
  DFF_X2 \u1/fracta_out_reg[55]  ( .D(\u1/fracta_s [55]), .CK(clk), .Q(
        fracta[55]) );
  DFF_X2 \fract_out_q_reg[0]  ( .D(n6093), .CK(clk), .Q(fract_out_q[0]) );
  DFF_X2 \fract_out_q_reg[1]  ( .D(n6092), .CK(clk), .Q(fract_out_q[1]) );
  DFF_X2 \fract_out_q_reg[2]  ( .D(n6091), .CK(clk), .Q(fract_out_q[2]) );
  DFF_X2 \fract_out_q_reg[3]  ( .D(n6090), .CK(clk), .Q(fract_out_q[3]) );
  DFF_X2 \fract_out_q_reg[4]  ( .D(n6089), .CK(clk), .Q(fract_out_q[4]) );
  DFF_X2 \fract_out_q_reg[5]  ( .D(n6088), .CK(clk), .Q(fract_out_q[5]) );
  DFF_X2 \fract_out_q_reg[6]  ( .D(n6087), .CK(clk), .Q(fract_out_q[6]) );
  DFF_X2 \fract_out_q_reg[7]  ( .D(n6086), .CK(clk), .Q(fract_out_q[7]) );
  DFF_X2 \fract_out_q_reg[8]  ( .D(n6085), .CK(clk), .Q(fract_out_q[8]) );
  DFF_X2 \fract_out_q_reg[9]  ( .D(n6084), .CK(clk), .Q(fract_out_q[9]) );
  DFF_X2 \fract_out_q_reg[10]  ( .D(n6083), .CK(clk), .Q(fract_out_q[10]) );
  DFF_X2 \fract_out_q_reg[11]  ( .D(n6082), .CK(clk), .Q(fract_out_q[11]) );
  DFF_X2 \fract_out_q_reg[12]  ( .D(n6081), .CK(clk), .Q(fract_out_q[12]) );
  DFF_X2 \fract_out_q_reg[13]  ( .D(n6080), .CK(clk), .Q(fract_out_q[13]) );
  DFF_X2 \fract_out_q_reg[14]  ( .D(n6079), .CK(clk), .Q(fract_out_q[14]) );
  DFF_X2 \fract_out_q_reg[15]  ( .D(n6078), .CK(clk), .Q(fract_out_q[15]) );
  DFF_X2 \fract_out_q_reg[16]  ( .D(n6077), .CK(clk), .Q(fract_out_q[16]) );
  DFF_X2 \fract_out_q_reg[17]  ( .D(n6076), .CK(clk), .Q(fract_out_q[17]) );
  DFF_X2 \fract_out_q_reg[18]  ( .D(n6075), .CK(clk), .Q(fract_out_q[18]) );
  DFF_X2 \fract_out_q_reg[19]  ( .D(n6074), .CK(clk), .Q(fract_out_q[19]) );
  DFF_X2 \fract_out_q_reg[20]  ( .D(n6073), .CK(clk), .Q(fract_out_q[20]) );
  DFF_X2 \fract_out_q_reg[21]  ( .D(n6072), .CK(clk), .Q(fract_out_q[21]) );
  DFF_X2 \fract_out_q_reg[22]  ( .D(n6071), .CK(clk), .Q(fract_out_q[22]) );
  DFF_X2 \fract_out_q_reg[23]  ( .D(n6070), .CK(clk), .Q(fract_out_q[23]) );
  DFF_X2 \fract_out_q_reg[24]  ( .D(n6069), .CK(clk), .Q(fract_out_q[24]) );
  DFF_X2 \fract_out_q_reg[25]  ( .D(n6068), .CK(clk), .Q(fract_out_q[25]) );
  DFF_X2 \fract_out_q_reg[26]  ( .D(n6067), .CK(clk), .Q(fract_out_q[26]) );
  DFF_X2 \fract_out_q_reg[27]  ( .D(n6066), .CK(clk), .Q(fract_out_q[27]) );
  DFF_X2 \fract_out_q_reg[28]  ( .D(n6065), .CK(clk), .Q(fract_out_q[28]) );
  DFF_X2 \fract_out_q_reg[29]  ( .D(n6064), .CK(clk), .Q(fract_out_q[29]) );
  DFF_X2 \fract_out_q_reg[30]  ( .D(n6063), .CK(clk), .Q(fract_out_q[30]) );
  DFF_X2 \fract_out_q_reg[31]  ( .D(n6062), .CK(clk), .Q(fract_out_q[31]) );
  DFF_X2 \fract_out_q_reg[32]  ( .D(n6061), .CK(clk), .Q(fract_out_q[32]) );
  DFF_X2 \fract_out_q_reg[33]  ( .D(n6060), .CK(clk), .Q(fract_out_q[33]) );
  DFF_X2 \fract_out_q_reg[34]  ( .D(n6059), .CK(clk), .Q(fract_out_q[34]) );
  DFF_X2 \fract_out_q_reg[35]  ( .D(n6058), .CK(clk), .Q(fract_out_q[35]) );
  DFF_X2 \fract_out_q_reg[36]  ( .D(n6057), .CK(clk), .Q(fract_out_q[36]) );
  DFF_X2 \fract_out_q_reg[37]  ( .D(n6056), .CK(clk), .Q(fract_out_q[37]) );
  DFF_X2 \fract_out_q_reg[38]  ( .D(n6055), .CK(clk), .Q(fract_out_q[38]) );
  DFF_X2 \fract_out_q_reg[39]  ( .D(n6054), .CK(clk), .Q(fract_out_q[39]) );
  DFF_X2 \fract_out_q_reg[40]  ( .D(n6053), .CK(clk), .Q(fract_out_q[40]) );
  DFF_X2 \fract_out_q_reg[41]  ( .D(n6052), .CK(clk), .Q(fract_out_q[41]) );
  DFF_X2 \fract_out_q_reg[42]  ( .D(n6051), .CK(clk), .Q(fract_out_q[42]) );
  DFF_X2 \fract_out_q_reg[43]  ( .D(n6050), .CK(clk), .Q(fract_out_q[43]) );
  DFF_X2 \fract_out_q_reg[44]  ( .D(n6049), .CK(clk), .Q(fract_out_q[44]) );
  DFF_X2 \fract_out_q_reg[45]  ( .D(n6048), .CK(clk), .Q(fract_out_q[45]) );
  DFF_X2 \fract_out_q_reg[46]  ( .D(n6047), .CK(clk), .Q(fract_out_q[46]) );
  DFF_X2 \fract_out_q_reg[47]  ( .D(n6046), .CK(clk), .Q(fract_out_q[47]) );
  DFF_X2 \fract_out_q_reg[48]  ( .D(n6045), .CK(clk), .Q(fract_out_q[48]) );
  DFF_X2 \fract_out_q_reg[49]  ( .D(n6044), .CK(clk), .Q(fract_out_q[49]) );
  DFF_X2 \fract_out_q_reg[50]  ( .D(n6043), .CK(clk), .Q(fract_out_q[50]) );
  DFF_X2 \fract_out_q_reg[51]  ( .D(n6042), .CK(clk), .Q(fract_out_q[51]) );
  DFF_X2 \fract_out_q_reg[52]  ( .D(n6041), .CK(clk), .Q(fract_out_q[52]) );
  DFF_X2 \fract_out_q_reg[53]  ( .D(n6040), .CK(clk), .Q(fract_out_q[53]) );
  DFF_X2 \fract_out_q_reg[54]  ( .D(n6039), .CK(clk), .Q(fract_out_q[54]) );
  DFF_X2 \fract_out_q_reg[55]  ( .D(n6038), .CK(clk), .Q(fract_out_q[55]) );
  DFF_X2 \fract_out_q_reg[56]  ( .D(n6037), .CK(clk), .Q(fract_out_q[56]) );
  DFF_X2 \u1/exp_dn_out_reg[0]  ( .D(\u1/N52 ), .CK(clk), .Q(exp_fasu[0]) );
  DFF_X2 \u1/exp_dn_out_reg[1]  ( .D(\u1/N53 ), .CK(clk), .Q(exp_fasu[1]) );
  DFF_X2 \u1/exp_dn_out_reg[2]  ( .D(\u1/N54 ), .CK(clk), .Q(exp_fasu[2]) );
  DFF_X2 \u1/exp_dn_out_reg[3]  ( .D(\u1/N55 ), .CK(clk), .Q(exp_fasu[3]) );
  DFF_X2 \u1/exp_dn_out_reg[4]  ( .D(\u1/N56 ), .CK(clk), .Q(exp_fasu[4]) );
  DFF_X2 \u1/exp_dn_out_reg[5]  ( .D(\u1/N57 ), .CK(clk), .Q(exp_fasu[5]) );
  DFF_X2 \u1/exp_dn_out_reg[6]  ( .D(\u1/N58 ), .CK(clk), .Q(exp_fasu[6]) );
  DFF_X2 \u1/exp_dn_out_reg[7]  ( .D(\u1/N59 ), .CK(clk), .Q(exp_fasu[7]) );
  DFF_X2 \u1/exp_dn_out_reg[8]  ( .D(\u1/N60 ), .CK(clk), .Q(exp_fasu[8]) );
  DFF_X2 \u1/exp_dn_out_reg[9]  ( .D(\u1/N61 ), .CK(clk), .Q(exp_fasu[9]) );
  DFF_X2 \u1/exp_dn_out_reg[10]  ( .D(\u1/N62 ), .CK(clk), .Q(exp_fasu[10]) );
  DFF_X2 \u2/sign_exe_reg  ( .D(\u2/N121 ), .CK(clk), .Q(sign_exe) );
  DFF_X2 sign_exe_r_reg ( .D(sign_exe), .CK(clk), .QN(n4482) );
  DFF_X2 \u2/sign_reg  ( .D(\u2/sign_d ), .CK(clk), .Q(sign_mul) );
  DFF_X2 sign_mul_r_reg ( .D(sign_mul), .CK(clk), .Q(sign_mul_r), .QN(n4491)
         );
  DFF_X2 sign_reg ( .D(N789), .CK(clk), .Q(sign), .QN(n4485) );
  DFF_X2 \fract_i2f_reg[105]  ( .D(N769), .CK(clk), .Q(fract_i2f[105]) );
  DFF_X2 \fract_i2f_reg[104]  ( .D(N768), .CK(clk), .Q(fract_i2f[104]) );
  DFF_X2 \fract_i2f_reg[103]  ( .D(N767), .CK(clk), .Q(fract_i2f[103]) );
  DFF_X2 \fract_i2f_reg[102]  ( .D(N766), .CK(clk), .Q(fract_i2f[102]) );
  DFF_X2 \fract_i2f_reg[101]  ( .D(N765), .CK(clk), .Q(fract_i2f[101]) );
  DFF_X2 \fract_i2f_reg[100]  ( .D(N764), .CK(clk), .Q(fract_i2f[100]) );
  DFF_X2 \fract_i2f_reg[99]  ( .D(N763), .CK(clk), .Q(fract_i2f[99]) );
  DFF_X2 \fract_i2f_reg[98]  ( .D(N762), .CK(clk), .Q(fract_i2f[98]) );
  DFF_X2 \fract_i2f_reg[97]  ( .D(N761), .CK(clk), .Q(fract_i2f[97]) );
  DFF_X2 \fract_i2f_reg[96]  ( .D(N760), .CK(clk), .Q(fract_i2f[96]) );
  DFF_X2 \fract_i2f_reg[95]  ( .D(N759), .CK(clk), .Q(fract_i2f[95]) );
  DFF_X2 \fract_i2f_reg[94]  ( .D(N758), .CK(clk), .Q(fract_i2f[94]) );
  DFF_X2 \fract_i2f_reg[93]  ( .D(N757), .CK(clk), .Q(fract_i2f[93]) );
  DFF_X2 \fract_i2f_reg[92]  ( .D(N756), .CK(clk), .Q(fract_i2f[92]) );
  DFF_X2 \fract_i2f_reg[91]  ( .D(N755), .CK(clk), .Q(fract_i2f[91]) );
  DFF_X2 \fract_i2f_reg[90]  ( .D(N754), .CK(clk), .Q(fract_i2f[90]) );
  DFF_X2 \fract_i2f_reg[89]  ( .D(N753), .CK(clk), .Q(fract_i2f[89]) );
  DFF_X2 \fract_i2f_reg[88]  ( .D(N752), .CK(clk), .Q(fract_i2f[88]) );
  DFF_X2 \fract_i2f_reg[87]  ( .D(N751), .CK(clk), .Q(fract_i2f[87]) );
  DFF_X2 \fract_i2f_reg[86]  ( .D(N750), .CK(clk), .Q(fract_i2f[86]) );
  DFF_X2 \fract_i2f_reg[85]  ( .D(N749), .CK(clk), .Q(fract_i2f[85]) );
  DFF_X2 \fract_i2f_reg[84]  ( .D(N748), .CK(clk), .Q(fract_i2f[84]) );
  DFF_X2 \fract_i2f_reg[83]  ( .D(N747), .CK(clk), .Q(fract_i2f[83]) );
  DFF_X2 \fract_i2f_reg[82]  ( .D(N746), .CK(clk), .Q(fract_i2f[82]) );
  DFF_X2 \fract_i2f_reg[81]  ( .D(N745), .CK(clk), .Q(fract_i2f[81]) );
  DFF_X2 \fract_i2f_reg[80]  ( .D(N744), .CK(clk), .Q(fract_i2f[80]) );
  DFF_X2 \fract_i2f_reg[79]  ( .D(N743), .CK(clk), .Q(fract_i2f[79]) );
  DFF_X2 \fract_i2f_reg[78]  ( .D(N742), .CK(clk), .Q(fract_i2f[78]) );
  DFF_X2 \fract_i2f_reg[77]  ( .D(N741), .CK(clk), .Q(fract_i2f[77]) );
  DFF_X2 \fract_i2f_reg[76]  ( .D(N740), .CK(clk), .Q(fract_i2f[76]) );
  DFF_X2 \fract_i2f_reg[75]  ( .D(N739), .CK(clk), .Q(fract_i2f[75]) );
  DFF_X2 \fract_i2f_reg[74]  ( .D(N738), .CK(clk), .Q(fract_i2f[74]) );
  DFF_X2 \fract_i2f_reg[73]  ( .D(N737), .CK(clk), .Q(fract_i2f[73]) );
  DFF_X2 \fract_i2f_reg[72]  ( .D(N736), .CK(clk), .Q(fract_i2f[72]) );
  DFF_X2 \fract_i2f_reg[71]  ( .D(N735), .CK(clk), .Q(fract_i2f[71]) );
  DFF_X2 \fract_i2f_reg[70]  ( .D(N734), .CK(clk), .Q(fract_i2f[70]) );
  DFF_X2 \fract_i2f_reg[69]  ( .D(N733), .CK(clk), .Q(fract_i2f[69]) );
  DFF_X2 \fract_i2f_reg[68]  ( .D(N732), .CK(clk), .Q(fract_i2f[68]) );
  DFF_X2 \fract_i2f_reg[67]  ( .D(N731), .CK(clk), .Q(fract_i2f[67]) );
  DFF_X2 \fract_i2f_reg[66]  ( .D(N730), .CK(clk), .Q(fract_i2f[66]) );
  DFF_X2 \fract_i2f_reg[65]  ( .D(N729), .CK(clk), .Q(fract_i2f[65]) );
  DFF_X2 \fract_i2f_reg[64]  ( .D(N728), .CK(clk), .Q(fract_i2f[64]) );
  DFF_X2 \fract_i2f_reg[63]  ( .D(N727), .CK(clk), .Q(fract_i2f[63]) );
  DFF_X2 \fract_i2f_reg[62]  ( .D(N726), .CK(clk), .Q(fract_i2f[62]) );
  DFF_X2 \fract_i2f_reg[61]  ( .D(N725), .CK(clk), .Q(fract_i2f[61]) );
  DFF_X2 \fract_i2f_reg[60]  ( .D(N724), .CK(clk), .Q(fract_i2f[60]) );
  DFF_X2 \fract_i2f_reg[59]  ( .D(N723), .CK(clk), .Q(fract_i2f[59]) );
  DFF_X2 \fract_i2f_reg[58]  ( .D(N722), .CK(clk), .Q(fract_i2f[58]) );
  DFF_X2 \fract_i2f_reg[57]  ( .D(N721), .CK(clk), .Q(fract_i2f[57]) );
  DFF_X2 \fract_i2f_reg[56]  ( .D(N720), .CK(clk), .Q(fract_i2f[56]) );
  DFF_X2 \fract_i2f_reg[55]  ( .D(N719), .CK(clk), .Q(fract_i2f[55]) );
  DFF_X2 \fract_i2f_reg[54]  ( .D(N718), .CK(clk), .Q(fract_i2f[54]) );
  DFF_X2 \fract_i2f_reg[53]  ( .D(N717), .CK(clk), .Q(fract_i2f[53]) );
  DFF_X2 \fract_i2f_reg[52]  ( .D(N716), .CK(clk), .Q(fract_i2f[52]) );
  DFF_X2 \fract_i2f_reg[51]  ( .D(N715), .CK(clk), .Q(fract_i2f[51]) );
  DFF_X2 \fract_i2f_reg[50]  ( .D(N714), .CK(clk), .Q(fract_i2f[50]) );
  DFF_X2 \fract_i2f_reg[49]  ( .D(N713), .CK(clk), .Q(fract_i2f[49]) );
  DFF_X2 \fract_i2f_reg[48]  ( .D(N712), .CK(clk), .Q(fract_i2f[48]) );
  DFF_X2 \fract_i2f_reg[47]  ( .D(N711), .CK(clk), .Q(fract_i2f[47]) );
  DFF_X2 \fract_i2f_reg[46]  ( .D(N710), .CK(clk), .Q(fract_i2f[46]) );
  DFF_X2 \fract_i2f_reg[45]  ( .D(n5913), .CK(clk), .Q(fract_i2f[45]) );
  DFF_X2 \fract_i2f_reg[44]  ( .D(n5914), .CK(clk), .Q(fract_i2f[44]) );
  DFF_X2 \fract_i2f_reg[43]  ( .D(n5915), .CK(clk), .Q(fract_i2f[43]) );
  DFF_X2 \fract_i2f_reg[42]  ( .D(n5916), .CK(clk), .Q(fract_i2f[42]) );
  DFF_X2 \fract_i2f_reg[41]  ( .D(n5917), .CK(clk), .Q(fract_i2f[41]) );
  DFF_X2 \fract_i2f_reg[40]  ( .D(n5918), .CK(clk), .Q(fract_i2f[40]) );
  DFF_X2 \fract_i2f_reg[39]  ( .D(n5919), .CK(clk), .Q(fract_i2f[39]) );
  DFF_X2 \fract_i2f_reg[38]  ( .D(n5920), .CK(clk), .Q(fract_i2f[38]) );
  DFF_X2 \fract_i2f_reg[37]  ( .D(n5921), .CK(clk), .Q(fract_i2f[37]) );
  DFF_X2 \fract_i2f_reg[36]  ( .D(n5922), .CK(clk), .Q(fract_i2f[36]) );
  DFF_X2 \fract_i2f_reg[35]  ( .D(n5923), .CK(clk), .Q(fract_i2f[35]) );
  DFF_X2 \fract_i2f_reg[34]  ( .D(n5924), .CK(clk), .Q(fract_i2f[34]) );
  DFF_X2 \fract_i2f_reg[33]  ( .D(n5925), .CK(clk), .Q(fract_i2f[33]) );
  DFF_X2 \fract_i2f_reg[32]  ( .D(n5926), .CK(clk), .Q(fract_i2f[32]) );
  DFF_X2 \fract_i2f_reg[31]  ( .D(n5927), .CK(clk), .Q(fract_i2f[31]) );
  DFF_X2 \fract_i2f_reg[30]  ( .D(n5928), .CK(clk), .Q(fract_i2f[30]) );
  DFF_X2 \fract_i2f_reg[29]  ( .D(n5929), .CK(clk), .Q(fract_i2f[29]) );
  DFF_X2 \fract_i2f_reg[28]  ( .D(n5930), .CK(clk), .Q(fract_i2f[28]) );
  DFF_X2 \fract_i2f_reg[27]  ( .D(n5931), .CK(clk), .Q(fract_i2f[27]) );
  DFF_X2 \fract_i2f_reg[26]  ( .D(n5932), .CK(clk), .Q(fract_i2f[26]) );
  DFF_X2 \fract_i2f_reg[25]  ( .D(n5933), .CK(clk), .Q(fract_i2f[25]) );
  DFF_X2 \fract_i2f_reg[24]  ( .D(n5934), .CK(clk), .Q(fract_i2f[24]) );
  DFF_X2 \fract_i2f_reg[23]  ( .D(n5935), .CK(clk), .Q(fract_i2f[23]) );
  DFF_X2 \fract_i2f_reg[22]  ( .D(n5936), .CK(clk), .Q(fract_i2f[22]) );
  DFF_X2 \fract_i2f_reg[21]  ( .D(n5937), .CK(clk), .Q(fract_i2f[21]) );
  DFF_X2 \fract_i2f_reg[20]  ( .D(n5938), .CK(clk), .Q(fract_i2f[20]) );
  DFF_X2 \fract_i2f_reg[19]  ( .D(n5939), .CK(clk), .Q(fract_i2f[19]) );
  DFF_X2 \fract_i2f_reg[18]  ( .D(n5940), .CK(clk), .Q(fract_i2f[18]) );
  DFF_X2 \fract_i2f_reg[17]  ( .D(n5941), .CK(clk), .Q(fract_i2f[17]) );
  DFF_X2 \fract_i2f_reg[16]  ( .D(n5942), .CK(clk), .Q(fract_i2f[16]) );
  DFF_X2 \fract_i2f_reg[15]  ( .D(n5943), .CK(clk), .Q(fract_i2f[15]) );
  DFF_X2 \fract_i2f_reg[14]  ( .D(n5944), .CK(clk), .Q(fract_i2f[14]) );
  DFF_X2 \fract_i2f_reg[13]  ( .D(n5945), .CK(clk), .Q(fract_i2f[13]) );
  DFF_X2 \fract_i2f_reg[12]  ( .D(n5946), .CK(clk), .Q(fract_i2f[12]) );
  DFF_X2 \fract_i2f_reg[11]  ( .D(n5947), .CK(clk), .Q(fract_i2f[11]) );
  DFF_X2 \fract_i2f_reg[10]  ( .D(n5948), .CK(clk), .Q(fract_i2f[10]) );
  DFF_X2 \fract_i2f_reg[9]  ( .D(n5949), .CK(clk), .Q(fract_i2f[9]) );
  DFF_X2 \fract_i2f_reg[8]  ( .D(n5950), .CK(clk), .Q(fract_i2f[8]) );
  DFF_X2 \fract_i2f_reg[7]  ( .D(n5951), .CK(clk), .Q(fract_i2f[7]) );
  DFF_X2 \fract_i2f_reg[6]  ( .D(n5952), .CK(clk), .Q(fract_i2f[6]) );
  DFF_X2 \fract_i2f_reg[5]  ( .D(n5953), .CK(clk), .Q(fract_i2f[5]) );
  DFF_X2 \fract_i2f_reg[4]  ( .D(n5954), .CK(clk), .Q(fract_i2f[4]) );
  DFF_X2 \fract_i2f_reg[3]  ( .D(n5955), .CK(clk), .Q(fract_i2f[3]) );
  DFF_X2 \fract_i2f_reg[2]  ( .D(n5956), .CK(clk), .Q(fract_i2f[2]) );
  DFF_X2 \fract_i2f_reg[1]  ( .D(n5957), .CK(clk), .Q(fract_i2f[1]) );
  DFF_X2 \fract_i2f_reg[0]  ( .D(n6311), .CK(clk), .Q(fract_i2f[0]) );
  DFF_X2 \u2/inf_reg  ( .D(\u2/N114 ), .CK(clk), .Q(inf_mul) );
  DFF_X2 inf_mul_r_reg ( .D(inf_mul), .CK(clk), .Q(inf_mul_r) );
  DFF_X2 \u2/underflow_reg[0]  ( .D(\u2/underflow_d [0]), .CK(clk), .Q(
        underflow_fmul_d[0]) );
  DFF_X2 \underflow_fmul_r_reg[0]  ( .D(underflow_fmul_d[0]), .CK(clk), .Q(
        underflow_fmul_r[0]) );
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  DFF_X2 \u2/underflow_reg[1]  ( .D(\u2/underflow_d [1]), .CK(clk), .Q(
        underflow_fmul_d[1]) );
  DFF_X2 \underflow_fmul_r_reg[1]  ( .D(underflow_fmul_d[1]), .CK(clk), .Q(
        underflow_fmul_r[1]) );
  DFF_X2 \u2/underflow_reg[2]  ( .D(\u2/underflow_d [2]), .CK(clk), .Q(
        underflow_fmul_d[2]) );
  DFF_X2 \underflow_fmul_r_reg[2]  ( .D(underflow_fmul_d[2]), .CK(clk), .Q(
        underflow_fmul_r[2]) );
  DFF_X2 \u2/exp_ovf_reg[0]  ( .D(\u2/exp_ovf_d[0] ), .CK(clk), .Q(exp_ovf[0])
         );
<<<<<<< HEAD
  DFF_X2 \exp_ovf_r_reg[0]  ( .D(exp_ovf[0]), .CK(clk), .Q(n1596), .QN(
        net11567) );
  DFF_X2 \u2/exp_ovf_reg[1]  ( .D(\u2/exp_ovf_d[1] ), .CK(clk), .Q(exp_ovf[1])
         );
  DFF_X2 \exp_ovf_r_reg[1]  ( .D(exp_ovf[1]), .CK(clk), .Q(n1571), .QN(
        net11566) );
  DFF_X2 \u2/exp_out_reg[0]  ( .D(\u2/N40 ), .CK(clk), .QN(n3070) );
  DFF_X2 \exp_r_reg[0]  ( .D(N96), .CK(clk), .Q(\u4/div_shft2[0] ), .QN(
        net11564) );
  DFF_X2 \u2/exp_out_reg[1]  ( .D(\u2/N41 ), .CK(clk), .QN(n3069) );
  DFF_X2 \exp_r_reg[1]  ( .D(N97), .CK(clk), .Q(exp_r[1]), .QN(net11562) );
  DFF_X2 \u2/exp_out_reg[2]  ( .D(\u2/N42 ), .CK(clk), .QN(n3068) );
  DFF_X2 \exp_r_reg[2]  ( .D(N98), .CK(clk), .Q(exp_r[2]), .QN(net11560) );
  DFF_X2 \u2/exp_out_reg[3]  ( .D(\u2/N43 ), .CK(clk), .QN(n3067) );
  DFF_X2 \exp_r_reg[3]  ( .D(N99), .CK(clk), .Q(exp_r[3]), .QN(net11558) );
  DFF_X2 \u2/exp_out_reg[4]  ( .D(\u2/N44 ), .CK(clk), .QN(n3066) );
  DFF_X2 inf_mul2_reg ( .D(N296), .CK(clk), .QN(n3065) );
  DFF_X2 \exp_r_reg[4]  ( .D(N100), .CK(clk), .Q(exp_r[4]), .QN(net11555) );
=======
  DFF_X2 \exp_ovf_r_reg[0]  ( .D(exp_ovf[0]), .CK(clk), .Q(exp_ovf_r[0]), .QN(
        n4356) );
  DFF_X2 \u2/exp_ovf_reg[1]  ( .D(\u2/exp_ovf_d[1] ), .CK(clk), .Q(exp_ovf[1])
         );
  DFF_X2 \exp_ovf_r_reg[1]  ( .D(exp_ovf[1]), .CK(clk), .Q(exp_ovf_r[1]), .QN(
        n4452) );
  DFF_X2 \u2/exp_out_reg[0]  ( .D(\u2/N76 ), .CK(clk), .QN(n4383) );
  DFF_X2 \exp_r_reg[0]  ( .D(N327), .CK(clk), .QN(n4349) );
  DFF_X2 \u2/exp_out_reg[1]  ( .D(\u2/N77 ), .CK(clk), .QN(n4487) );
  DFF_X2 \exp_r_reg[1]  ( .D(N328), .CK(clk), .Q(exp_r[1]), .QN(n4314) );
  DFF_X2 \u2/exp_out_reg[2]  ( .D(\u2/N78 ), .CK(clk), .Q(exp_mul[2]), .QN(
        n4539) );
  DFF_X2 \exp_r_reg[2]  ( .D(N329), .CK(clk), .Q(n4315), .QN(n4438) );
  DFF_X2 \u2/exp_out_reg[3]  ( .D(\u2/N79 ), .CK(clk), .Q(exp_mul[3]), .QN(
        n4538) );
  DFF_X2 \exp_r_reg[3]  ( .D(N330), .CK(clk), .Q(exp_r[3]), .QN(n4316) );
  DFF_X2 \u2/exp_out_reg[4]  ( .D(\u2/N80 ), .CK(clk), .Q(exp_mul[4]), .QN(
        n4537) );
  DFF_X2 \exp_r_reg[4]  ( .D(N331), .CK(clk), .Q(n4282), .QN(n4299) );
  DFF_X2 \u2/exp_out_reg[5]  ( .D(\u2/N81 ), .CK(clk), .Q(exp_mul[5]), .QN(
        n4535) );
  DFF_X2 \exp_r_reg[5]  ( .D(N332), .CK(clk), .Q(n4290), .QN(n4347) );
  DFF_X2 \u2/exp_out_reg[6]  ( .D(\u2/N82 ), .CK(clk), .Q(exp_mul[6]), .QN(
        n4536) );
  DFF_X2 \exp_r_reg[6]  ( .D(N333), .CK(clk), .Q(exp_r[6]), .QN(n4317) );
  DFF_X2 \u2/exp_out_reg[7]  ( .D(\u2/N83 ), .CK(clk), .Q(exp_mul[7]), .QN(
        n4534) );
  DFF_X2 \exp_r_reg[7]  ( .D(N334), .CK(clk), .Q(n4281), .QN(n4348) );
  DFF_X2 \u2/exp_out_reg[8]  ( .D(\u2/N84 ), .CK(clk), .QN(n4489) );
  DFF_X2 \exp_r_reg[8]  ( .D(N335), .CK(clk), .Q(n4353), .QN(n4439) );
  DFF_X2 \u2/exp_out_reg[9]  ( .D(\u2/N85 ), .CK(clk), .QN(n4384) );
  DFF_X2 \exp_r_reg[9]  ( .D(N336), .CK(clk), .Q(n4289), .QN(n4350) );
  DFF_X2 \u2/exp_out_reg[10]  ( .D(\u2/N86 ), .CK(clk), .QN(n4330) );
  DFF_X2 inf_mul2_reg ( .D(N923), .CK(clk), .Q(inf_mul2) );
  DFF_X2 \exp_r_reg[10]  ( .D(N337), .CK(clk), .Q(n4352), .QN(n4440) );
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  DFF_X2 \u5/prod1_reg[0]  ( .D(\u5/N0 ), .CK(clk), .Q(\u5/prod1 [0]) );
  DFF_X2 \u5/prod_reg[0]  ( .D(\u5/prod1 [0]), .CK(clk), .Q(prod[0]) );
  DFF_X2 \u5/prod1_reg[1]  ( .D(\u5/N1 ), .CK(clk), .Q(\u5/prod1 [1]) );
  DFF_X2 \u5/prod_reg[1]  ( .D(\u5/prod1 [1]), .CK(clk), .Q(prod[1]) );
  DFF_X2 \u5/prod1_reg[2]  ( .D(\u5/N2 ), .CK(clk), .Q(\u5/prod1 [2]) );
  DFF_X2 \u5/prod_reg[2]  ( .D(\u5/prod1 [2]), .CK(clk), .Q(prod[2]) );
  DFF_X2 \u5/prod1_reg[3]  ( .D(\u5/N3 ), .CK(clk), .Q(\u5/prod1 [3]) );
<<<<<<< HEAD
  DFF_X2 \u5/prod_reg[3]  ( .D(\u5/prod1 [3]), .CK(clk), .Q(prod[3]), .QN(
        net89543) );
  DFF_X2 \u5/prod1_reg[4]  ( .D(\u5/N4 ), .CK(clk), .Q(\u5/prod1 [4]) );
  DFF_X2 \u5/prod_reg[4]  ( .D(\u5/prod1 [4]), .CK(clk), .Q(prod[4]), .QN(
        net88972) );
=======
  DFF_X2 \u5/prod_reg[3]  ( .D(\u5/prod1 [3]), .CK(clk), .Q(prod[3]) );
  DFF_X2 \u5/prod1_reg[4]  ( .D(\u5/N4 ), .CK(clk), .Q(\u5/prod1 [4]) );
  DFF_X2 \u5/prod_reg[4]  ( .D(\u5/prod1 [4]), .CK(clk), .Q(prod[4]) );
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  DFF_X2 \u5/prod1_reg[5]  ( .D(\u5/N5 ), .CK(clk), .Q(\u5/prod1 [5]) );
  DFF_X2 \u5/prod_reg[5]  ( .D(\u5/prod1 [5]), .CK(clk), .Q(prod[5]) );
  DFF_X2 \u5/prod1_reg[6]  ( .D(\u5/N6 ), .CK(clk), .Q(\u5/prod1 [6]) );
  DFF_X2 \u5/prod_reg[6]  ( .D(\u5/prod1 [6]), .CK(clk), .Q(prod[6]) );
  DFF_X2 \u5/prod1_reg[7]  ( .D(\u5/N7 ), .CK(clk), .Q(\u5/prod1 [7]) );
<<<<<<< HEAD
  DFF_X2 \u5/prod_reg[7]  ( .D(\u5/prod1 [7]), .CK(clk), .Q(prod[7]), .QN(
        n1604) );
  DFF_X2 \u5/prod_reg[8]  ( .D(\u5/prod1 [8]), .CK(clk), .Q(prod[8]) );
  DFF_X2 \u5/prod1_reg[9]  ( .D(\u5/N9 ), .CK(clk), .Q(\u5/prod1 [9]) );
  DFF_X2 \u5/prod_reg[9]  ( .D(\u5/prod1 [9]), .CK(clk), .Q(prod[9]) );
  DFF_X2 \u5/prod_reg[10]  ( .D(\u5/prod1 [10]), .CK(clk), .Q(prod[10]) );
  DFF_X2 \u5/prod_reg[11]  ( .D(\u5/prod1 [11]), .CK(clk), .Q(prod[11]) );
  DFF_X2 \u5/prod1_reg[12]  ( .D(\u5/N12 ), .CK(clk), .Q(\u5/prod1 [12]) );
  DFF_X2 \u5/prod_reg[12]  ( .D(\u5/prod1 [12]), .CK(clk), .Q(prod[12]) );
=======
  DFF_X2 \u5/prod_reg[7]  ( .D(\u5/prod1 [7]), .CK(clk), .Q(prod[7]) );
  DFF_X2 \u5/prod1_reg[8]  ( .D(\u5/N8 ), .CK(clk), .Q(\u5/prod1 [8]) );
  DFF_X2 \u5/prod_reg[8]  ( .D(\u5/prod1 [8]), .CK(clk), .Q(prod[8]) );
  DFF_X2 \u5/prod1_reg[9]  ( .D(\u5/N9 ), .CK(clk), .Q(\u5/prod1 [9]) );
  DFF_X2 \u5/prod_reg[9]  ( .D(\u5/prod1 [9]), .CK(clk), .Q(prod[9]) );
  DFF_X2 \u5/prod1_reg[10]  ( .D(\u5/N10 ), .CK(clk), .Q(\u5/prod1 [10]) );
  DFF_X2 \u5/prod_reg[10]  ( .D(\u5/prod1 [10]), .CK(clk), .Q(prod[10]) );
  DFF_X2 \u5/prod1_reg[11]  ( .D(\u5/N11 ), .CK(clk), .Q(\u5/prod1 [11]) );
  DFF_X2 \u5/prod_reg[11]  ( .D(\u5/prod1 [11]), .CK(clk), .Q(prod[11]) );
  DFF_X2 \u5/prod1_reg[12]  ( .D(\u5/N12 ), .CK(clk), .Q(\u5/prod1 [12]) );
  DFF_X2 \u5/prod_reg[12]  ( .D(\u5/prod1 [12]), .CK(clk), .Q(prod[12]) );
  DFF_X2 \u5/prod1_reg[13]  ( .D(\u5/N13 ), .CK(clk), .Q(\u5/prod1 [13]) );
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  DFF_X2 \u5/prod_reg[13]  ( .D(\u5/prod1 [13]), .CK(clk), .Q(prod[13]) );
  DFF_X2 \u5/prod1_reg[14]  ( .D(\u5/N14 ), .CK(clk), .Q(\u5/prod1 [14]) );
  DFF_X2 \u5/prod_reg[14]  ( .D(\u5/prod1 [14]), .CK(clk), .Q(prod[14]) );
  DFF_X2 \u5/prod1_reg[15]  ( .D(\u5/N15 ), .CK(clk), .Q(\u5/prod1 [15]) );
  DFF_X2 \u5/prod_reg[15]  ( .D(\u5/prod1 [15]), .CK(clk), .Q(prod[15]) );
  DFF_X2 \u5/prod1_reg[16]  ( .D(\u5/N16 ), .CK(clk), .Q(\u5/prod1 [16]) );
  DFF_X2 \u5/prod_reg[16]  ( .D(\u5/prod1 [16]), .CK(clk), .Q(prod[16]) );
<<<<<<< HEAD
=======
  DFF_X2 \u5/prod1_reg[17]  ( .D(\u5/N17 ), .CK(clk), .Q(\u5/prod1 [17]) );
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  DFF_X2 \u5/prod_reg[17]  ( .D(\u5/prod1 [17]), .CK(clk), .Q(prod[17]) );
  DFF_X2 \u5/prod1_reg[18]  ( .D(\u5/N18 ), .CK(clk), .Q(\u5/prod1 [18]) );
  DFF_X2 \u5/prod_reg[18]  ( .D(\u5/prod1 [18]), .CK(clk), .Q(prod[18]) );
  DFF_X2 \u5/prod1_reg[19]  ( .D(\u5/N19 ), .CK(clk), .Q(\u5/prod1 [19]) );
  DFF_X2 \u5/prod_reg[19]  ( .D(\u5/prod1 [19]), .CK(clk), .Q(prod[19]) );
  DFF_X2 \u5/prod1_reg[20]  ( .D(\u5/N20 ), .CK(clk), .Q(\u5/prod1 [20]) );
  DFF_X2 \u5/prod_reg[20]  ( .D(\u5/prod1 [20]), .CK(clk), .Q(prod[20]) );
  DFF_X2 \u5/prod1_reg[21]  ( .D(\u5/N21 ), .CK(clk), .Q(\u5/prod1 [21]) );
  DFF_X2 \u5/prod_reg[21]  ( .D(\u5/prod1 [21]), .CK(clk), .Q(prod[21]) );
<<<<<<< HEAD
  DFF_X2 \u6/remainder_reg[0]  ( .D(\u6/N0 ), .CK(clk), .Q(\u6/remainder [0])
         );
  DFF_X2 \u6/rem_reg[0]  ( .D(\u6/remainder [0]), .CK(clk), .QN(n1568) );
  DFF_X2 \u6/remainder_reg[1]  ( .D(\u6/N1 ), .CK(clk), .Q(\u6/remainder [1])
         );
  DFF_X2 \u6/rem_reg[1]  ( .D(\u6/remainder [1]), .CK(clk), .QN(n3064) );
  DFF_X2 \u6/remainder_reg[2]  ( .D(\u6/N2 ), .CK(clk), .Q(\u6/remainder [2])
         );
  DFF_X2 \u6/rem_reg[2]  ( .D(\u6/remainder [2]), .CK(clk), .QN(n3063) );
  DFF_X2 \u6/remainder_reg[3]  ( .D(\u6/N3 ), .CK(clk), .Q(\u6/remainder [3])
         );
  DFF_X2 \u6/rem_reg[3]  ( .D(\u6/remainder [3]), .CK(clk), .QN(n3062) );
  DFF_X2 \u6/remainder_reg[4]  ( .D(\u6/N4 ), .CK(clk), .Q(\u6/remainder [4])
         );
  DFF_X2 \u6/rem_reg[4]  ( .D(\u6/remainder [4]), .CK(clk), .QN(n1587) );
  DFF_X2 \u6/remainder_reg[5]  ( .D(\u6/N5 ), .CK(clk), .Q(\u6/remainder [5])
         );
  DFF_X2 \u6/rem_reg[5]  ( .D(\u6/remainder [5]), .CK(clk), .QN(n1620) );
  DFF_X2 \u6/remainder_reg[6]  ( .D(\u6/N6 ), .CK(clk), .Q(\u6/remainder [6])
         );
  DFF_X2 \u6/rem_reg[6]  ( .D(\u6/remainder [6]), .CK(clk), .QN(n1584) );
  DFF_X2 \u6/remainder_reg[7]  ( .D(\u6/N7 ), .CK(clk), .Q(\u6/remainder [7])
         );
  DFF_X2 \u6/rem_reg[7]  ( .D(\u6/remainder [7]), .CK(clk), .QN(n3061) );
  DFF_X2 \u6/remainder_reg[8]  ( .D(\u6/N8 ), .CK(clk), .Q(\u6/remainder [8])
         );
  DFF_X2 \u6/rem_reg[8]  ( .D(\u6/remainder [8]), .CK(clk), .QN(n3060) );
  DFF_X2 \u6/remainder_reg[9]  ( .D(\u6/N9 ), .CK(clk), .Q(\u6/remainder [9])
         );
  DFF_X2 \u6/rem_reg[9]  ( .D(\u6/remainder [9]), .CK(clk), .QN(n3059) );
  DFF_X2 \u6/remainder_reg[10]  ( .D(n1731), .CK(clk), .Q(\u6/remainder [10])
         );
  DFF_X2 \u6/rem_reg[10]  ( .D(\u6/remainder [10]), .CK(clk), .QN(n1616) );
  DFF_X2 \u6/remainder_reg[13]  ( .D(\u6/N13 ), .CK(clk), .Q(
        \u6/remainder [13]) );
  DFF_X2 \u6/rem_reg[13]  ( .D(\u6/remainder [13]), .CK(clk), .QN(n3058) );
  DFF_X2 \u6/remainder_reg[14]  ( .D(\u6/N14 ), .CK(clk), .Q(
        \u6/remainder [14]) );
  DFF_X2 \u6/rem_reg[14]  ( .D(\u6/remainder [14]), .CK(clk), .QN(n3057) );
  DFF_X2 \u6/remainder_reg[15]  ( .D(\u6/N15 ), .CK(clk), .Q(
        \u6/remainder [15]) );
  DFF_X2 \u6/rem_reg[15]  ( .D(\u6/remainder [15]), .CK(clk), .QN(n1566) );
  DFF_X2 \u6/remainder_reg[16]  ( .D(\u6/N16 ), .CK(clk), .Q(
        \u6/remainder [16]) );
  DFF_X2 \u6/rem_reg[16]  ( .D(\u6/remainder [16]), .CK(clk), .QN(n1585) );
  DFF_X2 \u6/remainder_reg[17]  ( .D(\u6/N17 ), .CK(clk), .Q(
        \u6/remainder [17]) );
  DFF_X2 \u6/rem_reg[17]  ( .D(\u6/remainder [17]), .CK(clk), .QN(n1618) );
  DFF_X2 \u6/remainder_reg[18]  ( .D(\u6/N18 ), .CK(clk), .Q(
        \u6/remainder [18]) );
  DFF_X2 \u6/rem_reg[18]  ( .D(\u6/remainder [18]), .CK(clk), .QN(n3056) );
  DFF_X2 \u6/remainder_reg[19]  ( .D(\u6/N19 ), .CK(clk), .Q(
        \u6/remainder [19]) );
  DFF_X2 \u6/rem_reg[19]  ( .D(\u6/remainder [19]), .CK(clk), .QN(n3055) );
  DFF_X2 \u6/remainder_reg[20]  ( .D(\u6/N20 ), .CK(clk), .Q(
        \u6/remainder [20]) );
  DFF_X2 \u6/rem_reg[20]  ( .D(\u6/remainder [20]), .CK(clk), .QN(n1567) );
  DFF_X2 \u6/remainder_reg[21]  ( .D(\u6/N21 ), .CK(clk), .Q(
        \u6/remainder [21]) );
  DFF_X2 \u6/rem_reg[21]  ( .D(\u6/remainder [21]), .CK(clk), .QN(n1586) );
  DFF_X2 \u6/remainder_reg[22]  ( .D(\u6/N22 ), .CK(clk), .Q(
        \u6/remainder [22]) );
  DFF_X2 \u6/rem_reg[22]  ( .D(\u6/remainder [22]), .CK(clk), .QN(n1619) );
  DFF_X2 \u6/remainder_reg[23]  ( .D(\u6/N23 ), .CK(clk), .Q(
        \u6/remainder [23]) );
  DFF_X2 \u6/rem_reg[23]  ( .D(\u6/remainder [23]), .CK(clk), .QN(n3054) );
=======
  DFF_X2 \u5/prod1_reg[22]  ( .D(\u5/N22 ), .CK(clk), .Q(\u5/prod1 [22]) );
  DFF_X2 \u5/prod_reg[22]  ( .D(\u5/prod1 [22]), .CK(clk), .Q(prod[22]) );
  DFF_X2 \u5/prod1_reg[23]  ( .D(\u5/N23 ), .CK(clk), .Q(\u5/prod1 [23]) );
  DFF_X2 \u5/prod_reg[23]  ( .D(\u5/prod1 [23]), .CK(clk), .Q(prod[23]) );
  DFF_X2 \u5/prod1_reg[24]  ( .D(\u5/N24 ), .CK(clk), .Q(\u5/prod1 [24]) );
  DFF_X2 \u5/prod_reg[24]  ( .D(\u5/prod1 [24]), .CK(clk), .Q(prod[24]) );
  DFF_X2 \u5/prod1_reg[25]  ( .D(\u5/N25 ), .CK(clk), .Q(\u5/prod1 [25]) );
  DFF_X2 \u5/prod_reg[25]  ( .D(\u5/prod1 [25]), .CK(clk), .Q(prod[25]) );
  DFF_X2 \u5/prod1_reg[26]  ( .D(\u5/N26 ), .CK(clk), .Q(\u5/prod1 [26]) );
  DFF_X2 \u5/prod_reg[26]  ( .D(\u5/prod1 [26]), .CK(clk), .Q(prod[26]) );
  DFF_X2 \u5/prod1_reg[27]  ( .D(\u5/N27 ), .CK(clk), .Q(\u5/prod1 [27]) );
  DFF_X2 \u5/prod_reg[27]  ( .D(\u5/prod1 [27]), .CK(clk), .Q(prod[27]) );
  DFF_X2 \u5/prod1_reg[28]  ( .D(\u5/N28 ), .CK(clk), .Q(\u5/prod1 [28]) );
  DFF_X2 \u5/prod_reg[28]  ( .D(\u5/prod1 [28]), .CK(clk), .Q(prod[28]) );
  DFF_X2 \u5/prod1_reg[29]  ( .D(\u5/N29 ), .CK(clk), .Q(\u5/prod1 [29]) );
  DFF_X2 \u5/prod_reg[29]  ( .D(\u5/prod1 [29]), .CK(clk), .Q(prod[29]) );
  DFF_X2 \u5/prod1_reg[30]  ( .D(\u5/N30 ), .CK(clk), .Q(\u5/prod1 [30]) );
  DFF_X2 \u5/prod_reg[30]  ( .D(\u5/prod1 [30]), .CK(clk), .Q(prod[30]) );
  DFF_X2 \u5/prod1_reg[31]  ( .D(\u5/N31 ), .CK(clk), .Q(\u5/prod1 [31]) );
  DFF_X2 \u5/prod_reg[31]  ( .D(\u5/prod1 [31]), .CK(clk), .Q(prod[31]) );
  DFF_X2 \u5/prod1_reg[32]  ( .D(\u5/N32 ), .CK(clk), .Q(\u5/prod1 [32]) );
  DFF_X2 \u5/prod_reg[32]  ( .D(\u5/prod1 [32]), .CK(clk), .Q(prod[32]) );
  DFF_X2 \u5/prod1_reg[33]  ( .D(\u5/N33 ), .CK(clk), .Q(\u5/prod1 [33]) );
  DFF_X2 \u5/prod_reg[33]  ( .D(\u5/prod1 [33]), .CK(clk), .Q(prod[33]) );
  DFF_X2 \u5/prod1_reg[34]  ( .D(\u5/N34 ), .CK(clk), .Q(\u5/prod1 [34]) );
  DFF_X2 \u5/prod_reg[34]  ( .D(\u5/prod1 [34]), .CK(clk), .Q(prod[34]) );
  DFF_X2 \u5/prod1_reg[35]  ( .D(\u5/N35 ), .CK(clk), .Q(\u5/prod1 [35]) );
  DFF_X2 \u5/prod_reg[35]  ( .D(\u5/prod1 [35]), .CK(clk), .Q(prod[35]) );
  DFF_X2 \u5/prod1_reg[36]  ( .D(\u5/N36 ), .CK(clk), .Q(\u5/prod1 [36]) );
  DFF_X2 \u5/prod_reg[36]  ( .D(\u5/prod1 [36]), .CK(clk), .Q(prod[36]) );
  DFF_X2 \u5/prod1_reg[37]  ( .D(\u5/N37 ), .CK(clk), .Q(\u5/prod1 [37]) );
  DFF_X2 \u5/prod_reg[37]  ( .D(\u5/prod1 [37]), .CK(clk), .Q(prod[37]) );
  DFF_X2 \u5/prod1_reg[38]  ( .D(\u5/N38 ), .CK(clk), .Q(\u5/prod1 [38]) );
  DFF_X2 \u5/prod_reg[38]  ( .D(\u5/prod1 [38]), .CK(clk), .Q(prod[38]) );
  DFF_X2 \u5/prod1_reg[39]  ( .D(\u5/N39 ), .CK(clk), .Q(\u5/prod1 [39]) );
  DFF_X2 \u5/prod_reg[39]  ( .D(\u5/prod1 [39]), .CK(clk), .Q(prod[39]) );
  DFF_X2 \u5/prod1_reg[40]  ( .D(\u5/N40 ), .CK(clk), .Q(\u5/prod1 [40]) );
  DFF_X2 \u5/prod_reg[40]  ( .D(\u5/prod1 [40]), .CK(clk), .Q(prod[40]) );
  DFF_X2 \u5/prod1_reg[41]  ( .D(\u5/N41 ), .CK(clk), .Q(\u5/prod1 [41]) );
  DFF_X2 \u5/prod_reg[41]  ( .D(\u5/prod1 [41]), .CK(clk), .Q(prod[41]) );
  DFF_X2 \u5/prod1_reg[42]  ( .D(\u5/N42 ), .CK(clk), .Q(\u5/prod1 [42]) );
  DFF_X2 \u5/prod_reg[42]  ( .D(\u5/prod1 [42]), .CK(clk), .Q(prod[42]) );
  DFF_X2 \u5/prod1_reg[43]  ( .D(\u5/N43 ), .CK(clk), .Q(\u5/prod1 [43]) );
  DFF_X2 \u5/prod_reg[43]  ( .D(\u5/prod1 [43]), .CK(clk), .Q(prod[43]) );
  DFF_X2 \u5/prod1_reg[44]  ( .D(\u5/N44 ), .CK(clk), .Q(\u5/prod1 [44]) );
  DFF_X2 \u5/prod_reg[44]  ( .D(\u5/prod1 [44]), .CK(clk), .Q(prod[44]) );
  DFF_X2 \u5/prod1_reg[45]  ( .D(\u5/N45 ), .CK(clk), .Q(\u5/prod1 [45]) );
  DFF_X2 \u5/prod_reg[45]  ( .D(\u5/prod1 [45]), .CK(clk), .Q(prod[45]) );
  DFF_X2 \u5/prod1_reg[46]  ( .D(\u5/N46 ), .CK(clk), .Q(\u5/prod1 [46]) );
  DFF_X2 \u5/prod_reg[46]  ( .D(\u5/prod1 [46]), .CK(clk), .Q(prod[46]) );
  DFF_X2 \u5/prod1_reg[47]  ( .D(\u5/N47 ), .CK(clk), .Q(\u5/prod1 [47]) );
  DFF_X2 \u5/prod_reg[47]  ( .D(\u5/prod1 [47]), .CK(clk), .Q(prod[47]) );
  DFF_X2 \u5/prod1_reg[48]  ( .D(\u5/N48 ), .CK(clk), .Q(\u5/prod1 [48]) );
  DFF_X2 \u5/prod_reg[48]  ( .D(\u5/prod1 [48]), .CK(clk), .Q(prod[48]) );
  DFF_X2 \u5/prod1_reg[49]  ( .D(\u5/N49 ), .CK(clk), .Q(\u5/prod1 [49]) );
  DFF_X2 \u5/prod_reg[49]  ( .D(\u5/prod1 [49]), .CK(clk), .Q(prod[49]) );
  DFF_X2 \u5/prod1_reg[50]  ( .D(\u5/N50 ), .CK(clk), .Q(\u5/prod1 [50]) );
  DFF_X2 \u5/prod_reg[50]  ( .D(\u5/prod1 [50]), .CK(clk), .Q(prod[50]), .QN(
        n4434) );
  DFF_X2 \u5/prod1_reg[51]  ( .D(\u5/N51 ), .CK(clk), .Q(\u5/prod1 [51]) );
  DFF_X2 \u5/prod_reg[51]  ( .D(\u5/prod1 [51]), .CK(clk), .Q(prod[51]), .QN(
        n4432) );
  DFF_X2 \u5/prod1_reg[52]  ( .D(\u5/N52 ), .CK(clk), .Q(\u5/prod1 [52]) );
  DFF_X2 \u5/prod_reg[52]  ( .D(\u5/prod1 [52]), .CK(clk), .Q(prod[52]), .QN(
        n4429) );
  DFF_X2 \u5/prod1_reg[53]  ( .D(\u5/N53 ), .CK(clk), .Q(\u5/prod1 [53]) );
  DFF_X2 \u5/prod_reg[53]  ( .D(\u5/prod1 [53]), .CK(clk), .Q(prod[53]), .QN(
        n4410) );
  DFF_X2 \u5/prod1_reg[54]  ( .D(\u5/N54 ), .CK(clk), .Q(\u5/prod1 [54]) );
  DFF_X2 \u5/prod_reg[54]  ( .D(\u5/prod1 [54]), .CK(clk), .Q(prod[54]), .QN(
        n4419) );
  DFF_X2 \u5/prod1_reg[55]  ( .D(\u5/N55 ), .CK(clk), .Q(\u5/prod1 [55]) );
  DFF_X2 \u5/prod_reg[55]  ( .D(\u5/prod1 [55]), .CK(clk), .QN(n4310) );
  DFF_X2 \u5/prod1_reg[56]  ( .D(\u5/N56 ), .CK(clk), .Q(\u5/prod1 [56]) );
  DFF_X2 \u5/prod_reg[56]  ( .D(\u5/prod1 [56]), .CK(clk), .QN(n4401) );
  DFF_X2 \u5/prod1_reg[57]  ( .D(\u5/N57 ), .CK(clk), .Q(\u5/prod1 [57]) );
  DFF_X2 \u5/prod_reg[57]  ( .D(\u5/prod1 [57]), .CK(clk), .QN(n4341) );
  DFF_X2 \u5/prod1_reg[58]  ( .D(\u5/N58 ), .CK(clk), .Q(\u5/prod1 [58]) );
  DFF_X2 \u5/prod_reg[58]  ( .D(\u5/prod1 [58]), .CK(clk), .Q(prod[58]), .QN(
        n4430) );
  DFF_X2 \u5/prod1_reg[59]  ( .D(\u5/N59 ), .CK(clk), .Q(\u5/prod1 [59]) );
  DFF_X2 \u5/prod_reg[59]  ( .D(\u5/prod1 [59]), .CK(clk), .Q(prod[59]), .QN(
        n4413) );
  DFF_X2 \u5/prod1_reg[60]  ( .D(\u5/N60 ), .CK(clk), .Q(\u5/prod1 [60]) );
  DFF_X2 \u5/prod_reg[60]  ( .D(\u5/prod1 [60]), .CK(clk), .QN(n4346) );
  DFF_X2 \u5/prod1_reg[61]  ( .D(\u5/N61 ), .CK(clk), .Q(\u5/prod1 [61]) );
  DFF_X2 \u5/prod_reg[61]  ( .D(\u5/prod1 [61]), .CK(clk), .QN(n4406) );
  DFF_X2 \u5/prod1_reg[62]  ( .D(\u5/N62 ), .CK(clk), .Q(\u5/prod1 [62]) );
  DFF_X2 \u5/prod_reg[62]  ( .D(\u5/prod1 [62]), .CK(clk), .QN(n4312) );
  DFF_X2 \u5/prod1_reg[63]  ( .D(\u5/N63 ), .CK(clk), .Q(\u5/prod1 [63]) );
  DFF_X2 \u5/prod_reg[63]  ( .D(\u5/prod1 [63]), .CK(clk), .QN(n4297) );
  DFF_X2 \u5/prod1_reg[64]  ( .D(\u5/N64 ), .CK(clk), .Q(\u5/prod1 [64]) );
  DFF_X2 \u5/prod_reg[64]  ( .D(\u5/prod1 [64]), .CK(clk), .Q(prod[64]), .QN(
        n4428) );
  DFF_X2 \u5/prod1_reg[65]  ( .D(\u5/N65 ), .CK(clk), .Q(\u5/prod1 [65]) );
  DFF_X2 \u5/prod_reg[65]  ( .D(\u5/prod1 [65]), .CK(clk), .Q(prod[65]), .QN(
        n4414) );
  DFF_X2 \u5/prod1_reg[66]  ( .D(\u5/N66 ), .CK(clk), .Q(\u5/prod1 [66]) );
  DFF_X2 \u5/prod_reg[66]  ( .D(\u5/prod1 [66]), .CK(clk), .Q(prod[66]), .QN(
        n4423) );
  DFF_X2 \u5/prod1_reg[67]  ( .D(\u5/N67 ), .CK(clk), .Q(\u5/prod1 [67]) );
  DFF_X2 \u5/prod_reg[67]  ( .D(\u5/prod1 [67]), .CK(clk), .QN(n4311) );
  DFF_X2 \u5/prod1_reg[68]  ( .D(\u5/N68 ), .CK(clk), .Q(\u5/prod1 [68]) );
  DFF_X2 \u5/prod_reg[68]  ( .D(\u5/prod1 [68]), .CK(clk), .QN(n4402) );
  DFF_X2 \u5/prod1_reg[69]  ( .D(\u5/N69 ), .CK(clk), .Q(\u5/prod1 [69]) );
  DFF_X2 \u5/prod_reg[69]  ( .D(\u5/prod1 [69]), .CK(clk), .QN(n4342) );
  DFF_X2 \u5/prod1_reg[70]  ( .D(\u5/N70 ), .CK(clk), .Q(\u5/prod1 [70]) );
  DFF_X2 \u5/prod_reg[70]  ( .D(\u5/prod1 [70]), .CK(clk), .Q(prod[70]), .QN(
        n4415) );
  DFF_X2 \u5/prod1_reg[71]  ( .D(\u5/N71 ), .CK(clk), .Q(\u5/prod1 [71]) );
  DFF_X2 \u5/prod_reg[71]  ( .D(\u5/prod1 [71]), .CK(clk), .Q(prod[71]), .QN(
        n4422) );
  DFF_X2 \u5/prod1_reg[72]  ( .D(\u5/N72 ), .CK(clk), .Q(\u5/prod1 [72]) );
  DFF_X2 \u5/prod_reg[72]  ( .D(\u5/prod1 [72]), .CK(clk), .QN(n4313) );
  DFF_X2 \u5/prod1_reg[73]  ( .D(\u5/N73 ), .CK(clk), .Q(\u5/prod1 [73]) );
  DFF_X2 \u5/prod_reg[73]  ( .D(\u5/prod1 [73]), .CK(clk), .QN(n4407) );
  DFF_X2 \u5/prod1_reg[74]  ( .D(\u5/N74 ), .CK(clk), .Q(\u5/prod1 [74]) );
  DFF_X2 \u5/prod_reg[74]  ( .D(\u5/prod1 [74]), .CK(clk), .QN(n4298) );
  DFF_X2 \u5/prod1_reg[75]  ( .D(\u5/N75 ), .CK(clk), .Q(\u5/prod1 [75]) );
  DFF_X2 \u5/prod_reg[75]  ( .D(\u5/prod1 [75]), .CK(clk), .QN(n4343) );
  DFF_X2 \u5/prod1_reg[76]  ( .D(\u5/N76 ), .CK(clk), .Q(\u5/prod1 [76]) );
  DFF_X2 \u5/prod_reg[76]  ( .D(\u5/prod1 [76]), .CK(clk), .Q(prod[76]), .QN(
        n4426) );
  DFF_X2 \u5/prod1_reg[77]  ( .D(\u5/N77 ), .CK(clk), .Q(\u5/prod1 [77]) );
  DFF_X2 \u5/prod_reg[77]  ( .D(\u5/prod1 [77]), .CK(clk), .Q(prod[77]), .QN(
        n4412) );
  DFF_X2 \u5/prod1_reg[78]  ( .D(\u5/N78 ), .CK(clk), .Q(\u5/prod1 [78]) );
  DFF_X2 \u5/prod_reg[78]  ( .D(\u5/prod1 [78]), .CK(clk), .Q(prod[78]), .QN(
        n4421) );
  DFF_X2 \u5/prod1_reg[79]  ( .D(\u5/N79 ), .CK(clk), .Q(\u5/prod1 [79]) );
  DFF_X2 \u5/prod_reg[79]  ( .D(\u5/prod1 [79]), .CK(clk), .Q(prod[79]), .QN(
        n4436) );
  DFF_X2 \u5/prod1_reg[80]  ( .D(\u5/N80 ), .CK(clk), .Q(\u5/prod1 [80]) );
  DFF_X2 \u5/prod_reg[80]  ( .D(\u5/prod1 [80]), .CK(clk), .Q(prod[80]), .QN(
        n4437) );
  DFF_X2 \u5/prod1_reg[81]  ( .D(\u5/N81 ), .CK(clk), .Q(\u5/prod1 [81]) );
  DFF_X2 \u5/prod_reg[81]  ( .D(\u5/prod1 [81]), .CK(clk), .Q(prod[81]), .QN(
        n4427) );
  DFF_X2 \u5/prod1_reg[82]  ( .D(\u5/N82 ), .CK(clk), .Q(\u5/prod1 [82]) );
  DFF_X2 \u5/prod_reg[82]  ( .D(\u5/prod1 [82]), .CK(clk), .Q(prod[82]), .QN(
        n4416) );
  DFF_X2 \u5/prod1_reg[83]  ( .D(\u5/N83 ), .CK(clk), .Q(\u5/prod1 [83]) );
  DFF_X2 \u5/prod_reg[83]  ( .D(\u5/prod1 [83]), .CK(clk), .Q(prod[83]), .QN(
        n4420) );
  DFF_X2 \u5/prod1_reg[84]  ( .D(\u5/N84 ), .CK(clk), .Q(\u5/prod1 [84]) );
  DFF_X2 \u5/prod_reg[84]  ( .D(\u5/prod1 [84]), .CK(clk), .QN(n4344) );
  DFF_X2 \u5/prod1_reg[85]  ( .D(\u5/N85 ), .CK(clk), .Q(\u5/prod1 [85]) );
  DFF_X2 \u5/prod_reg[85]  ( .D(\u5/prod1 [85]), .CK(clk), .QN(n4404) );
  DFF_X2 \u5/prod1_reg[86]  ( .D(\u5/N86 ), .CK(clk), .Q(\u5/prod1 [86]) );
  DFF_X2 \u5/prod_reg[86]  ( .D(\u5/prod1 [86]), .CK(clk), .QN(n4307) );
  DFF_X2 \u5/prod1_reg[87]  ( .D(\u5/N87 ), .CK(clk), .Q(\u5/prod1 [87]) );
  DFF_X2 \u5/prod_reg[87]  ( .D(\u5/prod1 [87]), .CK(clk), .QN(n4294) );
  DFF_X2 \u5/prod1_reg[88]  ( .D(\u5/N88 ), .CK(clk), .Q(\u5/prod1 [88]) );
  DFF_X2 \u5/prod_reg[88]  ( .D(\u5/prod1 [88]), .CK(clk), .Q(prod[88]), .QN(
        n4425) );
  DFF_X2 \u5/prod1_reg[89]  ( .D(\u5/N89 ), .CK(clk), .Q(\u5/prod1 [89]) );
  DFF_X2 \u5/prod_reg[89]  ( .D(\u5/prod1 [89]), .CK(clk), .Q(prod[89]), .QN(
        n4411) );
  DFF_X2 \u5/prod1_reg[90]  ( .D(\u5/N90 ), .CK(clk), .Q(\u5/prod1 [90]) );
  DFF_X2 \u5/prod_reg[90]  ( .D(\u5/prod1 [90]), .CK(clk), .QN(n4345) );
  DFF_X2 \u5/prod1_reg[91]  ( .D(\u5/N91 ), .CK(clk), .Q(\u5/prod1 [91]) );
  DFF_X2 \u5/prod_reg[91]  ( .D(\u5/prod1 [91]), .CK(clk), .QN(n4405) );
  DFF_X2 \u5/prod1_reg[92]  ( .D(\u5/N92 ), .CK(clk), .Q(\u5/prod1 [92]) );
  DFF_X2 \u5/prod_reg[92]  ( .D(\u5/prod1 [92]), .CK(clk), .QN(n4308) );
  DFF_X2 \u5/prod1_reg[93]  ( .D(\u5/N93 ), .CK(clk), .Q(\u5/prod1 [93]) );
  DFF_X2 \u5/prod_reg[93]  ( .D(\u5/prod1 [93]), .CK(clk), .QN(n4295) );
  DFF_X2 \u5/prod1_reg[94]  ( .D(\u5/N94 ), .CK(clk), .Q(\u5/prod1 [94]) );
  DFF_X2 \u5/prod_reg[94]  ( .D(\u5/prod1 [94]), .CK(clk), .Q(prod[94]), .QN(
        n4424) );
  DFF_X2 \u5/prod1_reg[95]  ( .D(\u5/N95 ), .CK(clk), .Q(\u5/prod1 [95]) );
  DFF_X2 \u5/prod_reg[95]  ( .D(\u5/prod1 [95]), .CK(clk), .Q(prod[95]), .QN(
        n4408) );
  DFF_X2 \u5/prod1_reg[96]  ( .D(\u5/N96 ), .CK(clk), .Q(\u5/prod1 [96]) );
  DFF_X2 \u5/prod_reg[96]  ( .D(\u5/prod1 [96]), .CK(clk), .Q(prod[96]), .QN(
        n4417) );
  DFF_X2 \u5/prod1_reg[97]  ( .D(\u5/N97 ), .CK(clk), .Q(\u5/prod1 [97]) );
  DFF_X2 \u5/prod_reg[97]  ( .D(\u5/prod1 [97]), .CK(clk), .Q(prod[97]), .QN(
        n4431) );
  DFF_X2 \u5/prod1_reg[98]  ( .D(\u5/N98 ), .CK(clk), .Q(\u5/prod1 [98]) );
  DFF_X2 \u5/prod_reg[98]  ( .D(\u5/prod1 [98]), .CK(clk), .Q(prod[98]), .QN(
        n4435) );
  DFF_X2 \u5/prod1_reg[99]  ( .D(\u5/N99 ), .CK(clk), .Q(\u5/prod1 [99]) );
  DFF_X2 \u5/prod_reg[99]  ( .D(\u5/prod1 [99]), .CK(clk), .Q(prod[99]), .QN(
        n4433) );
  DFF_X2 \u5/prod1_reg[100]  ( .D(\u5/N100 ), .CK(clk), .Q(\u5/prod1 [100]) );
  DFF_X2 \u5/prod_reg[100]  ( .D(\u5/prod1 [100]), .CK(clk), .Q(prod[100]), 
        .QN(n4409) );
  DFF_X2 \u5/prod1_reg[101]  ( .D(\u5/N101 ), .CK(clk), .Q(\u5/prod1 [101]) );
  DFF_X2 \u5/prod_reg[101]  ( .D(\u5/prod1 [101]), .CK(clk), .Q(prod[101]), 
        .QN(n4418) );
  DFF_X2 \u5/prod1_reg[102]  ( .D(\u5/N102 ), .CK(clk), .Q(\u5/prod1 [102]) );
  DFF_X2 \u5/prod_reg[102]  ( .D(\u5/prod1 [102]), .CK(clk), .QN(n4306) );
  DFF_X2 \u5/prod1_reg[103]  ( .D(\u5/N103 ), .CK(clk), .Q(\u5/prod1 [103]) );
  DFF_X2 \u5/prod_reg[103]  ( .D(\u5/prod1 [103]), .CK(clk), .QN(n4403) );
  DFF_X2 \u5/prod1_reg[104]  ( .D(\u5/N104 ), .CK(clk), .Q(\u5/prod1 [104]) );
  DFF_X2 \u5/prod_reg[104]  ( .D(\u5/prod1 [104]), .CK(clk), .QN(n4338) );
  DFF_X2 \u5/prod1_reg[105]  ( .D(\u5/N105 ), .CK(clk), .Q(\u5/prod1 [105]) );
  DFF_X2 \u5/prod_reg[105]  ( .D(\u5/prod1 [105]), .CK(clk), .Q(prod[105]) );
  DFF_X2 \u6/remainder_reg[0]  ( .D(\u6/N0 ), .CK(clk), .Q(\u6/remainder [0])
         );
  DFF_X2 \u6/rem_reg[0]  ( .D(\u6/remainder [0]), .CK(clk), .Q(remainder[0])
         );
  DFF_X2 \u6/remainder_reg[1]  ( .D(\u6/N1 ), .CK(clk), .Q(\u6/remainder [1])
         );
  DFF_X2 \u6/rem_reg[1]  ( .D(\u6/remainder [1]), .CK(clk), .Q(remainder[1])
         );
  DFF_X2 \u6/remainder_reg[2]  ( .D(\u6/N2 ), .CK(clk), .Q(\u6/remainder [2])
         );
  DFF_X2 \u6/rem_reg[2]  ( .D(\u6/remainder [2]), .CK(clk), .Q(remainder[2])
         );
  DFF_X2 \u6/remainder_reg[3]  ( .D(\u6/N3 ), .CK(clk), .Q(\u6/remainder [3])
         );
  DFF_X2 \u6/rem_reg[3]  ( .D(\u6/remainder [3]), .CK(clk), .Q(remainder[3])
         );
  DFF_X2 \u6/remainder_reg[4]  ( .D(\u6/N4 ), .CK(clk), .Q(\u6/remainder [4])
         );
  DFF_X2 \u6/rem_reg[4]  ( .D(\u6/remainder [4]), .CK(clk), .Q(remainder[4])
         );
  DFF_X2 \u6/remainder_reg[5]  ( .D(\u6/N5 ), .CK(clk), .Q(\u6/remainder [5])
         );
  DFF_X2 \u6/rem_reg[5]  ( .D(\u6/remainder [5]), .CK(clk), .Q(remainder[5])
         );
  DFF_X2 \u6/remainder_reg[6]  ( .D(\u6/N6 ), .CK(clk), .Q(\u6/remainder [6])
         );
  DFF_X2 \u6/rem_reg[6]  ( .D(\u6/remainder [6]), .CK(clk), .Q(remainder[6])
         );
  DFF_X2 \u6/remainder_reg[7]  ( .D(\u6/N7 ), .CK(clk), .Q(\u6/remainder [7])
         );
  DFF_X2 \u6/rem_reg[7]  ( .D(\u6/remainder [7]), .CK(clk), .Q(remainder[7])
         );
  DFF_X2 \u6/remainder_reg[8]  ( .D(\u6/N8 ), .CK(clk), .Q(\u6/remainder [8])
         );
  DFF_X2 \u6/rem_reg[8]  ( .D(\u6/remainder [8]), .CK(clk), .Q(remainder[8])
         );
  DFF_X2 \u6/remainder_reg[9]  ( .D(\u6/N9 ), .CK(clk), .Q(\u6/remainder [9])
         );
  DFF_X2 \u6/rem_reg[9]  ( .D(\u6/remainder [9]), .CK(clk), .Q(remainder[9])
         );
  DFF_X2 \u6/remainder_reg[10]  ( .D(\u6/N10 ), .CK(clk), .Q(
        \u6/remainder [10]) );
  DFF_X2 \u6/rem_reg[10]  ( .D(\u6/remainder [10]), .CK(clk), .Q(remainder[10]) );
  DFF_X2 \u6/remainder_reg[11]  ( .D(\u6/N11 ), .CK(clk), .Q(
        \u6/remainder [11]) );
  DFF_X2 \u6/rem_reg[11]  ( .D(\u6/remainder [11]), .CK(clk), .Q(remainder[11]) );
  DFF_X2 \u6/remainder_reg[12]  ( .D(\u6/N12 ), .CK(clk), .Q(
        \u6/remainder [12]) );
  DFF_X2 \u6/rem_reg[12]  ( .D(\u6/remainder [12]), .CK(clk), .Q(remainder[12]) );
  DFF_X2 \u6/remainder_reg[13]  ( .D(\u6/N13 ), .CK(clk), .Q(
        \u6/remainder [13]) );
  DFF_X2 \u6/rem_reg[13]  ( .D(\u6/remainder [13]), .CK(clk), .Q(remainder[13]) );
  DFF_X2 \u6/remainder_reg[14]  ( .D(\u6/N14 ), .CK(clk), .Q(
        \u6/remainder [14]) );
  DFF_X2 \u6/rem_reg[14]  ( .D(\u6/remainder [14]), .CK(clk), .Q(remainder[14]) );
  DFF_X2 \u6/remainder_reg[15]  ( .D(\u6/N15 ), .CK(clk), .Q(
        \u6/remainder [15]) );
  DFF_X2 \u6/rem_reg[15]  ( .D(\u6/remainder [15]), .CK(clk), .Q(remainder[15]) );
  DFF_X2 \u6/remainder_reg[16]  ( .D(\u6/N16 ), .CK(clk), .Q(
        \u6/remainder [16]) );
  DFF_X2 \u6/rem_reg[16]  ( .D(\u6/remainder [16]), .CK(clk), .Q(remainder[16]) );
  DFF_X2 \u6/remainder_reg[17]  ( .D(\u6/N17 ), .CK(clk), .Q(
        \u6/remainder [17]) );
  DFF_X2 \u6/rem_reg[17]  ( .D(\u6/remainder [17]), .CK(clk), .Q(remainder[17]) );
  DFF_X2 \u6/remainder_reg[18]  ( .D(\u6/N18 ), .CK(clk), .Q(
        \u6/remainder [18]) );
  DFF_X2 \u6/rem_reg[18]  ( .D(\u6/remainder [18]), .CK(clk), .Q(remainder[18]) );
  DFF_X2 \u6/remainder_reg[19]  ( .D(\u6/N19 ), .CK(clk), .Q(
        \u6/remainder [19]) );
  DFF_X2 \u6/rem_reg[19]  ( .D(\u6/remainder [19]), .CK(clk), .Q(remainder[19]) );
  DFF_X2 \u6/remainder_reg[20]  ( .D(\u6/N20 ), .CK(clk), .Q(
        \u6/remainder [20]) );
  DFF_X2 \u6/rem_reg[20]  ( .D(\u6/remainder [20]), .CK(clk), .Q(remainder[20]) );
  DFF_X2 \u6/remainder_reg[21]  ( .D(\u6/N21 ), .CK(clk), .Q(
        \u6/remainder [21]) );
  DFF_X2 \u6/rem_reg[21]  ( .D(\u6/remainder [21]), .CK(clk), .Q(remainder[21]) );
  DFF_X2 \u6/remainder_reg[22]  ( .D(\u6/N22 ), .CK(clk), .Q(
        \u6/remainder [22]) );
  DFF_X2 \u6/rem_reg[22]  ( .D(\u6/remainder [22]), .CK(clk), .Q(remainder[22]) );
  DFF_X2 \u6/remainder_reg[23]  ( .D(\u6/N23 ), .CK(clk), .Q(
        \u6/remainder [23]) );
  DFF_X2 \u6/rem_reg[23]  ( .D(\u6/remainder [23]), .CK(clk), .Q(remainder[23]) );
  DFF_X2 \u6/remainder_reg[24]  ( .D(\u6/N24 ), .CK(clk), .Q(
        \u6/remainder [24]) );
  DFF_X2 \u6/rem_reg[24]  ( .D(\u6/remainder [24]), .CK(clk), .Q(remainder[24]) );
  DFF_X2 \u6/remainder_reg[25]  ( .D(\u6/N25 ), .CK(clk), .Q(
        \u6/remainder [25]) );
  DFF_X2 \u6/rem_reg[25]  ( .D(\u6/remainder [25]), .CK(clk), .Q(remainder[25]) );
  DFF_X2 \u6/remainder_reg[26]  ( .D(\u6/N26 ), .CK(clk), .Q(
        \u6/remainder [26]) );
  DFF_X2 \u6/rem_reg[26]  ( .D(\u6/remainder [26]), .CK(clk), .Q(remainder[26]) );
  DFF_X2 \u6/remainder_reg[27]  ( .D(\u6/N27 ), .CK(clk), .Q(
        \u6/remainder [27]) );
  DFF_X2 \u6/rem_reg[27]  ( .D(\u6/remainder [27]), .CK(clk), .Q(remainder[27]) );
  DFF_X2 \u6/remainder_reg[28]  ( .D(\u6/N28 ), .CK(clk), .Q(
        \u6/remainder [28]) );
  DFF_X2 \u6/rem_reg[28]  ( .D(\u6/remainder [28]), .CK(clk), .Q(remainder[28]) );
  DFF_X2 \u6/remainder_reg[29]  ( .D(\u6/N29 ), .CK(clk), .Q(
        \u6/remainder [29]) );
  DFF_X2 \u6/rem_reg[29]  ( .D(\u6/remainder [29]), .CK(clk), .Q(remainder[29]) );
  DFF_X2 \u6/remainder_reg[30]  ( .D(\u6/N30 ), .CK(clk), .Q(
        \u6/remainder [30]) );
  DFF_X2 \u6/rem_reg[30]  ( .D(\u6/remainder [30]), .CK(clk), .Q(remainder[30]) );
  DFF_X2 \u6/remainder_reg[31]  ( .D(\u6/N31 ), .CK(clk), .Q(
        \u6/remainder [31]) );
  DFF_X2 \u6/rem_reg[31]  ( .D(\u6/remainder [31]), .CK(clk), .Q(remainder[31]) );
  DFF_X2 \u6/remainder_reg[32]  ( .D(\u6/N32 ), .CK(clk), .Q(
        \u6/remainder [32]) );
  DFF_X2 \u6/rem_reg[32]  ( .D(\u6/remainder [32]), .CK(clk), .Q(remainder[32]) );
  DFF_X2 \u6/remainder_reg[33]  ( .D(\u6/N33 ), .CK(clk), .Q(
        \u6/remainder [33]) );
  DFF_X2 \u6/rem_reg[33]  ( .D(\u6/remainder [33]), .CK(clk), .Q(remainder[33]) );
  DFF_X2 \u6/remainder_reg[34]  ( .D(\u6/N34 ), .CK(clk), .Q(
        \u6/remainder [34]) );
  DFF_X2 \u6/rem_reg[34]  ( .D(\u6/remainder [34]), .CK(clk), .Q(remainder[34]) );
  DFF_X2 \u6/remainder_reg[35]  ( .D(\u6/N35 ), .CK(clk), .Q(
        \u6/remainder [35]) );
  DFF_X2 \u6/rem_reg[35]  ( .D(\u6/remainder [35]), .CK(clk), .Q(remainder[35]) );
  DFF_X2 \u6/remainder_reg[36]  ( .D(\u6/N36 ), .CK(clk), .Q(
        \u6/remainder [36]) );
  DFF_X2 \u6/rem_reg[36]  ( .D(\u6/remainder [36]), .CK(clk), .Q(remainder[36]) );
  DFF_X2 \u6/remainder_reg[37]  ( .D(\u6/N37 ), .CK(clk), .Q(
        \u6/remainder [37]) );
  DFF_X2 \u6/rem_reg[37]  ( .D(\u6/remainder [37]), .CK(clk), .Q(remainder[37]) );
  DFF_X2 \u6/remainder_reg[38]  ( .D(\u6/N38 ), .CK(clk), .Q(
        \u6/remainder [38]) );
  DFF_X2 \u6/rem_reg[38]  ( .D(\u6/remainder [38]), .CK(clk), .Q(remainder[38]) );
  DFF_X2 \u6/remainder_reg[39]  ( .D(\u6/N39 ), .CK(clk), .Q(
        \u6/remainder [39]) );
  DFF_X2 \u6/rem_reg[39]  ( .D(\u6/remainder [39]), .CK(clk), .Q(remainder[39]) );
  DFF_X2 \u6/remainder_reg[40]  ( .D(\u6/N40 ), .CK(clk), .Q(
        \u6/remainder [40]) );
  DFF_X2 \u6/rem_reg[40]  ( .D(\u6/remainder [40]), .CK(clk), .Q(remainder[40]) );
  DFF_X2 \u6/remainder_reg[41]  ( .D(\u6/N41 ), .CK(clk), .Q(
        \u6/remainder [41]) );
  DFF_X2 \u6/rem_reg[41]  ( .D(\u6/remainder [41]), .CK(clk), .Q(remainder[41]) );
  DFF_X2 \u6/remainder_reg[42]  ( .D(\u6/N42 ), .CK(clk), .Q(
        \u6/remainder [42]) );
  DFF_X2 \u6/rem_reg[42]  ( .D(\u6/remainder [42]), .CK(clk), .Q(remainder[42]) );
  DFF_X2 \u6/remainder_reg[43]  ( .D(\u6/N43 ), .CK(clk), .Q(
        \u6/remainder [43]) );
  DFF_X2 \u6/rem_reg[43]  ( .D(\u6/remainder [43]), .CK(clk), .Q(remainder[43]) );
  DFF_X2 \u6/remainder_reg[44]  ( .D(\u6/N44 ), .CK(clk), .Q(
        \u6/remainder [44]) );
  DFF_X2 \u6/rem_reg[44]  ( .D(\u6/remainder [44]), .CK(clk), .Q(remainder[44]) );
  DFF_X2 \u6/remainder_reg[45]  ( .D(\u6/N45 ), .CK(clk), .Q(
        \u6/remainder [45]) );
  DFF_X2 \u6/rem_reg[45]  ( .D(\u6/remainder [45]), .CK(clk), .Q(remainder[45]) );
  DFF_X2 \u6/remainder_reg[46]  ( .D(\u6/N46 ), .CK(clk), .Q(
        \u6/remainder [46]) );
  DFF_X2 \u6/rem_reg[46]  ( .D(\u6/remainder [46]), .CK(clk), .Q(remainder[46]) );
  DFF_X2 \u6/remainder_reg[47]  ( .D(\u6/N47 ), .CK(clk), .Q(
        \u6/remainder [47]) );
  DFF_X2 \u6/rem_reg[47]  ( .D(\u6/remainder [47]), .CK(clk), .Q(remainder[47]) );
  DFF_X2 \u6/remainder_reg[48]  ( .D(\u6/N48 ), .CK(clk), .Q(
        \u6/remainder [48]) );
  DFF_X2 \u6/rem_reg[48]  ( .D(\u6/remainder [48]), .CK(clk), .Q(remainder[48]) );
  DFF_X2 \u6/remainder_reg[49]  ( .D(\u6/N49 ), .CK(clk), .Q(
        \u6/remainder [49]) );
  DFF_X2 \u6/rem_reg[49]  ( .D(\u6/remainder [49]), .CK(clk), .Q(remainder[49]) );
  DFF_X2 \u6/remainder_reg[50]  ( .D(\u6/N50 ), .CK(clk), .Q(
        \u6/remainder [50]) );
  DFF_X2 \u6/rem_reg[50]  ( .D(\u6/remainder [50]), .CK(clk), .Q(remainder[50]) );
  DFF_X2 \u6/remainder_reg[51]  ( .D(\u6/N51 ), .CK(clk), .Q(
        \u6/remainder [51]) );
  DFF_X2 \u6/rem_reg[51]  ( .D(\u6/remainder [51]), .CK(clk), .Q(remainder[51]) );
  DFF_X2 \u6/remainder_reg[52]  ( .D(\u6/N52 ), .CK(clk), .Q(
        \u6/remainder [52]) );
  DFF_X2 \u6/rem_reg[52]  ( .D(\u6/remainder [52]), .CK(clk), .Q(remainder[52]) );
  DFF_X2 \u6/remainder_reg[55]  ( .D(\u6/N55 ), .CK(clk), .Q(
        \u6/remainder [55]) );
  DFF_X2 \u6/rem_reg[55]  ( .D(\u6/remainder [55]), .CK(clk), .Q(remainder[55]) );
  DFF_X2 \u6/remainder_reg[56]  ( .D(\u6/N56 ), .CK(clk), .Q(
        \u6/remainder [56]) );
  DFF_X2 \u6/rem_reg[56]  ( .D(\u6/remainder [56]), .CK(clk), .Q(remainder[56]) );
  DFF_X2 \u6/remainder_reg[57]  ( .D(\u6/N57 ), .CK(clk), .Q(
        \u6/remainder [57]) );
  DFF_X2 \u6/rem_reg[57]  ( .D(\u6/remainder [57]), .CK(clk), .Q(remainder[57]) );
  DFF_X2 \u6/remainder_reg[58]  ( .D(\u6/N58 ), .CK(clk), .Q(
        \u6/remainder [58]) );
  DFF_X2 \u6/rem_reg[58]  ( .D(\u6/remainder [58]), .CK(clk), .Q(remainder[58]) );
  DFF_X2 \u6/remainder_reg[59]  ( .D(\u6/N59 ), .CK(clk), .Q(
        \u6/remainder [59]) );
  DFF_X2 \u6/rem_reg[59]  ( .D(\u6/remainder [59]), .CK(clk), .Q(remainder[59]) );
  DFF_X2 \u6/remainder_reg[60]  ( .D(\u6/N60 ), .CK(clk), .Q(
        \u6/remainder [60]) );
  DFF_X2 \u6/rem_reg[60]  ( .D(\u6/remainder [60]), .CK(clk), .Q(remainder[60]) );
  DFF_X2 \u6/remainder_reg[61]  ( .D(\u6/N61 ), .CK(clk), .Q(
        \u6/remainder [61]) );
  DFF_X2 \u6/rem_reg[61]  ( .D(\u6/remainder [61]), .CK(clk), .Q(remainder[61]) );
  DFF_X2 \u6/remainder_reg[62]  ( .D(\u6/N62 ), .CK(clk), .Q(
        \u6/remainder [62]) );
  DFF_X2 \u6/rem_reg[62]  ( .D(\u6/remainder [62]), .CK(clk), .Q(remainder[62]) );
  DFF_X2 \u6/remainder_reg[63]  ( .D(\u6/N63 ), .CK(clk), .Q(
        \u6/remainder [63]) );
  DFF_X2 \u6/rem_reg[63]  ( .D(\u6/remainder [63]), .CK(clk), .Q(remainder[63]) );
  DFF_X2 \u6/remainder_reg[64]  ( .D(\u6/N64 ), .CK(clk), .Q(
        \u6/remainder [64]) );
  DFF_X2 \u6/rem_reg[64]  ( .D(\u6/remainder [64]), .CK(clk), .Q(remainder[64]) );
  DFF_X2 \u6/remainder_reg[65]  ( .D(\u6/N65 ), .CK(clk), .Q(
        \u6/remainder [65]) );
  DFF_X2 \u6/rem_reg[65]  ( .D(\u6/remainder [65]), .CK(clk), .Q(remainder[65]) );
  DFF_X2 \u6/remainder_reg[66]  ( .D(\u6/N66 ), .CK(clk), .Q(
        \u6/remainder [66]) );
  DFF_X2 \u6/rem_reg[66]  ( .D(\u6/remainder [66]), .CK(clk), .Q(remainder[66]) );
  DFF_X2 \u6/remainder_reg[67]  ( .D(\u6/N67 ), .CK(clk), .Q(
        \u6/remainder [67]) );
  DFF_X2 \u6/rem_reg[67]  ( .D(\u6/remainder [67]), .CK(clk), .Q(remainder[67]) );
  DFF_X2 \u6/remainder_reg[68]  ( .D(\u6/N68 ), .CK(clk), .Q(
        \u6/remainder [68]) );
  DFF_X2 \u6/rem_reg[68]  ( .D(\u6/remainder [68]), .CK(clk), .Q(remainder[68]) );
  DFF_X2 \u6/remainder_reg[69]  ( .D(\u6/N69 ), .CK(clk), .Q(
        \u6/remainder [69]) );
  DFF_X2 \u6/rem_reg[69]  ( .D(\u6/remainder [69]), .CK(clk), .Q(remainder[69]) );
  DFF_X2 \u6/remainder_reg[70]  ( .D(\u6/N70 ), .CK(clk), .Q(
        \u6/remainder [70]) );
  DFF_X2 \u6/rem_reg[70]  ( .D(\u6/remainder [70]), .CK(clk), .Q(remainder[70]) );
  DFF_X2 \u6/remainder_reg[71]  ( .D(\u6/N71 ), .CK(clk), .Q(
        \u6/remainder [71]) );
  DFF_X2 \u6/rem_reg[71]  ( .D(\u6/remainder [71]), .CK(clk), .Q(remainder[71]) );
  DFF_X2 \u6/remainder_reg[72]  ( .D(\u6/N72 ), .CK(clk), .Q(
        \u6/remainder [72]) );
  DFF_X2 \u6/rem_reg[72]  ( .D(\u6/remainder [72]), .CK(clk), .Q(remainder[72]) );
  DFF_X2 \u6/remainder_reg[73]  ( .D(\u6/N73 ), .CK(clk), .Q(
        \u6/remainder [73]) );
  DFF_X2 \u6/rem_reg[73]  ( .D(\u6/remainder [73]), .CK(clk), .Q(remainder[73]) );
  DFF_X2 \u6/remainder_reg[74]  ( .D(\u6/N74 ), .CK(clk), .Q(
        \u6/remainder [74]) );
  DFF_X2 \u6/rem_reg[74]  ( .D(\u6/remainder [74]), .CK(clk), .Q(remainder[74]) );
  DFF_X2 \u6/remainder_reg[75]  ( .D(\u6/N75 ), .CK(clk), .Q(
        \u6/remainder [75]) );
  DFF_X2 \u6/rem_reg[75]  ( .D(\u6/remainder [75]), .CK(clk), .Q(remainder[75]) );
  DFF_X2 \u6/remainder_reg[76]  ( .D(\u6/N76 ), .CK(clk), .Q(
        \u6/remainder [76]) );
  DFF_X2 \u6/rem_reg[76]  ( .D(\u6/remainder [76]), .CK(clk), .Q(remainder[76]) );
  DFF_X2 \u6/remainder_reg[77]  ( .D(\u6/N77 ), .CK(clk), .Q(
        \u6/remainder [77]) );
  DFF_X2 \u6/rem_reg[77]  ( .D(\u6/remainder [77]), .CK(clk), .Q(remainder[77]) );
  DFF_X2 \u6/remainder_reg[78]  ( .D(\u6/N78 ), .CK(clk), .Q(
        \u6/remainder [78]) );
  DFF_X2 \u6/rem_reg[78]  ( .D(\u6/remainder [78]), .CK(clk), .Q(remainder[78]) );
  DFF_X2 \u6/remainder_reg[79]  ( .D(\u6/N79 ), .CK(clk), .Q(
        \u6/remainder [79]) );
  DFF_X2 \u6/rem_reg[79]  ( .D(\u6/remainder [79]), .CK(clk), .Q(remainder[79]) );
  DFF_X2 \u6/remainder_reg[80]  ( .D(\u6/N80 ), .CK(clk), .Q(
        \u6/remainder [80]) );
  DFF_X2 \u6/rem_reg[80]  ( .D(\u6/remainder [80]), .CK(clk), .Q(remainder[80]) );
  DFF_X2 \u6/remainder_reg[81]  ( .D(\u6/N81 ), .CK(clk), .Q(
        \u6/remainder [81]) );
  DFF_X2 \u6/rem_reg[81]  ( .D(\u6/remainder [81]), .CK(clk), .Q(remainder[81]) );
  DFF_X2 \u6/remainder_reg[82]  ( .D(\u6/N82 ), .CK(clk), .Q(
        \u6/remainder [82]) );
  DFF_X2 \u6/rem_reg[82]  ( .D(\u6/remainder [82]), .CK(clk), .Q(remainder[82]) );
  DFF_X2 \u6/remainder_reg[83]  ( .D(\u6/N83 ), .CK(clk), .Q(
        \u6/remainder [83]) );
  DFF_X2 \u6/rem_reg[83]  ( .D(\u6/remainder [83]), .CK(clk), .Q(remainder[83]) );
  DFF_X2 \u6/remainder_reg[84]  ( .D(\u6/N84 ), .CK(clk), .Q(
        \u6/remainder [84]) );
  DFF_X2 \u6/rem_reg[84]  ( .D(\u6/remainder [84]), .CK(clk), .Q(remainder[84]) );
  DFF_X2 \u6/remainder_reg[85]  ( .D(\u6/N85 ), .CK(clk), .Q(
        \u6/remainder [85]) );
  DFF_X2 \u6/rem_reg[85]  ( .D(\u6/remainder [85]), .CK(clk), .Q(remainder[85]) );
  DFF_X2 \u6/remainder_reg[86]  ( .D(\u6/N86 ), .CK(clk), .Q(
        \u6/remainder [86]) );
  DFF_X2 \u6/rem_reg[86]  ( .D(\u6/remainder [86]), .CK(clk), .Q(remainder[86]) );
  DFF_X2 \u6/remainder_reg[87]  ( .D(\u6/N87 ), .CK(clk), .Q(
        \u6/remainder [87]) );
  DFF_X2 \u6/rem_reg[87]  ( .D(\u6/remainder [87]), .CK(clk), .Q(remainder[87]) );
  DFF_X2 \u6/remainder_reg[88]  ( .D(\u6/N88 ), .CK(clk), .Q(
        \u6/remainder [88]) );
  DFF_X2 \u6/rem_reg[88]  ( .D(\u6/remainder [88]), .CK(clk), .Q(remainder[88]) );
  DFF_X2 \u6/remainder_reg[89]  ( .D(\u6/N89 ), .CK(clk), .Q(
        \u6/remainder [89]) );
  DFF_X2 \u6/rem_reg[89]  ( .D(\u6/remainder [89]), .CK(clk), .Q(remainder[89]) );
  DFF_X2 \u6/remainder_reg[90]  ( .D(\u6/N90 ), .CK(clk), .Q(
        \u6/remainder [90]) );
  DFF_X2 \u6/rem_reg[90]  ( .D(\u6/remainder [90]), .CK(clk), .Q(remainder[90]) );
  DFF_X2 \u6/remainder_reg[91]  ( .D(\u6/N91 ), .CK(clk), .Q(
        \u6/remainder [91]) );
  DFF_X2 \u6/rem_reg[91]  ( .D(\u6/remainder [91]), .CK(clk), .Q(remainder[91]) );
  DFF_X2 \u6/remainder_reg[92]  ( .D(\u6/N92 ), .CK(clk), .Q(
        \u6/remainder [92]) );
  DFF_X2 \u6/rem_reg[92]  ( .D(\u6/remainder [92]), .CK(clk), .Q(remainder[92]) );
  DFF_X2 \u6/remainder_reg[93]  ( .D(\u6/N93 ), .CK(clk), .Q(
        \u6/remainder [93]) );
  DFF_X2 \u6/rem_reg[93]  ( .D(\u6/remainder [93]), .CK(clk), .Q(remainder[93]) );
  DFF_X2 \u6/remainder_reg[94]  ( .D(\u6/N94 ), .CK(clk), .Q(
        \u6/remainder [94]) );
  DFF_X2 \u6/rem_reg[94]  ( .D(\u6/remainder [94]), .CK(clk), .Q(remainder[94]) );
  DFF_X2 \u6/remainder_reg[95]  ( .D(\u6/N95 ), .CK(clk), .Q(
        \u6/remainder [95]) );
  DFF_X2 \u6/rem_reg[95]  ( .D(\u6/remainder [95]), .CK(clk), .Q(remainder[95]) );
  DFF_X2 \u6/remainder_reg[96]  ( .D(\u6/N96 ), .CK(clk), .Q(
        \u6/remainder [96]) );
  DFF_X2 \u6/rem_reg[96]  ( .D(\u6/remainder [96]), .CK(clk), .Q(remainder[96]) );
  DFF_X2 \u6/remainder_reg[97]  ( .D(\u6/N97 ), .CK(clk), .Q(
        \u6/remainder [97]) );
  DFF_X2 \u6/rem_reg[97]  ( .D(\u6/remainder [97]), .CK(clk), .Q(remainder[97]) );
  DFF_X2 \u6/remainder_reg[98]  ( .D(\u6/N98 ), .CK(clk), .Q(
        \u6/remainder [98]) );
  DFF_X2 \u6/rem_reg[98]  ( .D(\u6/remainder [98]), .CK(clk), .Q(remainder[98]) );
  DFF_X2 \u6/remainder_reg[99]  ( .D(\u6/N99 ), .CK(clk), .Q(
        \u6/remainder [99]) );
  DFF_X2 \u6/rem_reg[99]  ( .D(\u6/remainder [99]), .CK(clk), .Q(remainder[99]) );
  DFF_X2 \u6/remainder_reg[100]  ( .D(\u6/N100 ), .CK(clk), .Q(
        \u6/remainder [100]) );
  DFF_X2 \u6/rem_reg[100]  ( .D(\u6/remainder [100]), .CK(clk), .Q(
        remainder[100]) );
  DFF_X2 \u6/remainder_reg[101]  ( .D(\u6/N101 ), .CK(clk), .Q(
        \u6/remainder [101]) );
  DFF_X2 \u6/rem_reg[101]  ( .D(\u6/remainder [101]), .CK(clk), .Q(
        remainder[101]) );
  DFF_X2 \u6/remainder_reg[102]  ( .D(\u6/N102 ), .CK(clk), .Q(
        \u6/remainder [102]) );
  DFF_X2 \u6/rem_reg[102]  ( .D(\u6/remainder [102]), .CK(clk), .Q(
        remainder[102]) );
  DFF_X2 \u6/remainder_reg[103]  ( .D(\u6/N103 ), .CK(clk), .Q(
        \u6/remainder [103]) );
  DFF_X2 \u6/rem_reg[103]  ( .D(\u6/remainder [103]), .CK(clk), .Q(
        remainder[103]) );
  DFF_X2 \u6/remainder_reg[104]  ( .D(\u6/N104 ), .CK(clk), .Q(
        \u6/remainder [104]) );
  DFF_X2 \u6/rem_reg[104]  ( .D(\u6/remainder [104]), .CK(clk), .Q(
        remainder[104]) );
  DFF_X2 \u6/remainder_reg[105]  ( .D(\u6/N105 ), .CK(clk), .Q(
        \u6/remainder [105]) );
  DFF_X2 \u6/rem_reg[105]  ( .D(\u6/remainder [105]), .CK(clk), .Q(
        remainder[105]) );
  DFF_X2 \u6/remainder_reg[106]  ( .D(\u6/N106 ), .CK(clk), .Q(
        \u6/remainder [106]) );
  DFF_X2 \u6/rem_reg[106]  ( .D(\u6/remainder [106]), .CK(clk), .Q(
        remainder[106]) );
  DFF_X2 \u6/remainder_reg[107]  ( .D(\u6/N107 ), .CK(clk), .Q(
        \u6/remainder [107]) );
  DFF_X2 \u6/rem_reg[107]  ( .D(\u6/remainder [107]), .CK(clk), .Q(
        remainder[107]) );
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  DFF_X2 \u6/quo1_reg[0]  ( .D(\u6/N0 ), .CK(clk), .Q(\u6/quo1 [0]) );
  DFF_X2 \u6/quo_reg[0]  ( .D(\u6/quo1 [0]), .CK(clk), .Q(quo[0]) );
  DFF_X2 \u6/quo1_reg[1]  ( .D(\u6/N1 ), .CK(clk), .Q(\u6/quo1 [1]) );
  DFF_X2 \u6/quo_reg[1]  ( .D(\u6/quo1 [1]), .CK(clk), .Q(quo[1]) );
  DFF_X2 \u6/quo1_reg[2]  ( .D(\u6/N2 ), .CK(clk), .Q(\u6/quo1 [2]) );
<<<<<<< HEAD
  DFF_X2 \u6/quo_reg[2]  ( .D(\u6/quo1 [2]), .CK(clk), .Q(quo[2]), .QN(n1642)
         );
=======
  DFF_X2 \u6/quo_reg[2]  ( .D(\u6/quo1 [2]), .CK(clk), .Q(quo[2]) );
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  DFF_X2 \u6/quo1_reg[3]  ( .D(\u6/N3 ), .CK(clk), .Q(\u6/quo1 [3]) );
  DFF_X2 \u6/quo_reg[3]  ( .D(\u6/quo1 [3]), .CK(clk), .Q(quo[3]) );
  DFF_X2 \u6/quo1_reg[4]  ( .D(\u6/N4 ), .CK(clk), .Q(\u6/quo1 [4]) );
  DFF_X2 \u6/quo_reg[4]  ( .D(\u6/quo1 [4]), .CK(clk), .Q(quo[4]) );
  DFF_X2 \u6/quo1_reg[5]  ( .D(\u6/N5 ), .CK(clk), .Q(\u6/quo1 [5]) );
<<<<<<< HEAD
  DFF_X2 \u6/quo_reg[5]  ( .D(\u6/quo1 [5]), .CK(clk), .Q(quo[5]), .QN(n1650)
         );
=======
  DFF_X2 \u6/quo_reg[5]  ( .D(\u6/quo1 [5]), .CK(clk), .Q(quo[5]) );
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  DFF_X2 \u6/quo1_reg[6]  ( .D(\u6/N6 ), .CK(clk), .Q(\u6/quo1 [6]) );
  DFF_X2 \u6/quo_reg[6]  ( .D(\u6/quo1 [6]), .CK(clk), .Q(quo[6]) );
  DFF_X2 \u6/quo1_reg[7]  ( .D(\u6/N7 ), .CK(clk), .Q(\u6/quo1 [7]) );
  DFF_X2 \u6/quo_reg[7]  ( .D(\u6/quo1 [7]), .CK(clk), .Q(quo[7]) );
  DFF_X2 \u6/quo1_reg[8]  ( .D(\u6/N8 ), .CK(clk), .Q(\u6/quo1 [8]) );
  DFF_X2 \u6/quo_reg[8]  ( .D(\u6/quo1 [8]), .CK(clk), .Q(quo[8]) );
  DFF_X2 \u6/quo1_reg[9]  ( .D(\u6/N9 ), .CK(clk), .Q(\u6/quo1 [9]) );
<<<<<<< HEAD
  DFF_X2 \u6/quo_reg[9]  ( .D(\u6/quo1 [9]), .CK(clk), .Q(quo[9]), .QN(n1937)
         );
  DFF_X2 \u6/quo1_reg[10]  ( .D(n1731), .CK(clk), .Q(\u6/quo1 [10]) );
  DFF_X2 \u6/quo_reg[10]  ( .D(\u6/quo1 [10]), .CK(clk), .Q(quo[10]) );
  DFF_X2 \u6/quo1_reg[13]  ( .D(\u6/N13 ), .CK(clk), .Q(\u6/quo1 [13]) );
  DFF_X2 \u6/quo_reg[13]  ( .D(\u6/quo1 [13]), .CK(clk), .Q(quo[13]), .QN(
        net86061) );
=======
  DFF_X2 \u6/quo_reg[9]  ( .D(\u6/quo1 [9]), .CK(clk), .Q(quo[9]) );
  DFF_X2 \u6/quo1_reg[10]  ( .D(\u6/N10 ), .CK(clk), .Q(\u6/quo1 [10]) );
  DFF_X2 \u6/quo_reg[10]  ( .D(\u6/quo1 [10]), .CK(clk), .Q(quo[10]) );
  DFF_X2 \u6/quo1_reg[11]  ( .D(\u6/N11 ), .CK(clk), .Q(\u6/quo1 [11]) );
  DFF_X2 \u6/quo_reg[11]  ( .D(\u6/quo1 [11]), .CK(clk), .Q(quo[11]) );
  DFF_X2 \u6/quo1_reg[12]  ( .D(\u6/N12 ), .CK(clk), .Q(\u6/quo1 [12]) );
  DFF_X2 \u6/quo_reg[12]  ( .D(\u6/quo1 [12]), .CK(clk), .Q(quo[12]) );
  DFF_X2 \u6/quo1_reg[13]  ( .D(\u6/N13 ), .CK(clk), .Q(\u6/quo1 [13]) );
  DFF_X2 \u6/quo_reg[13]  ( .D(\u6/quo1 [13]), .CK(clk), .Q(quo[13]) );
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
  DFF_X2 \u6/quo1_reg[14]  ( .D(\u6/N14 ), .CK(clk), .Q(\u6/quo1 [14]) );
  DFF_X2 \u6/quo_reg[14]  ( .D(\u6/quo1 [14]), .CK(clk), .Q(quo[14]) );
  DFF_X2 \u6/quo1_reg[15]  ( .D(\u6/N15 ), .CK(clk), .Q(\u6/quo1 [15]) );
  DFF_X2 \u6/quo_reg[15]  ( .D(\u6/quo1 [15]), .CK(clk), .Q(quo[15]) );
  DFF_X2 \u6/quo1_reg[16]  ( .D(\u6/N16 ), .CK(clk), .Q(\u6/quo1 [16]) );
  DFF_X2 \u6/quo_reg[16]  ( .D(\u6/quo1 [16]), .CK(clk), .Q(quo[16]) );
  DFF_X2 \u6/quo1_reg[17]  ( .D(\u6/N17 ), .CK(clk), .Q(\u6/quo1 [17]) );
  DFF_X2 \u6/quo_reg[17]  ( .D(\u6/quo1 [17]), .CK(clk), .Q(quo[17]) );
  DFF_X2 \u6/quo1_reg[18]  ( .D(\u6/N18 ), .CK(clk), .Q(\u6/quo1 [18]) );
  DFF_X2 \u6/quo_reg[18]  ( .D(\u6/quo1 [18]), .CK(clk), .Q(quo[18]) );
  DFF_X2 \u6/quo1_reg[19]  ( .D(\u6/N19 ), .CK(clk), .Q(\u6/quo1 [19]) );
  DFF_X2 \u6/quo_reg[19]  ( .D(\u6/quo1 [19]), .CK(clk), .Q(quo[19]) );
  DFF_X2 \u6/quo1_reg[20]  ( .D(\u6/N20 ), .CK(clk), .Q(\u6/quo1 [20]) );
  DFF_X2 \u6/quo_reg[20]  ( .D(\u6/quo1 [20]), .CK(clk), .Q(quo[20]) );
  DFF_X2 \u6/quo1_reg[21]  ( .D(\u6/N21 ), .CK(clk), .Q(\u6/quo1 [21]) );
  DFF_X2 \u6/quo_reg[21]  ( .D(\u6/quo1 [21]), .CK(clk), .Q(quo[21]) );
  DFF_X2 \u6/quo1_reg[22]  ( .D(\u6/N22 ), .CK(clk), .Q(\u6/quo1 [22]) );
  DFF_X2 \u6/quo_reg[22]  ( .D(\u6/quo1 [22]), .CK(clk), .Q(quo[22]) );
<<<<<<< HEAD
  DFF_X2 \out_reg[13]  ( .D(N233), .CK(clk), .Q(out[13]) );
  DFF_X2 \out_reg[14]  ( .D(N234), .CK(clk), .Q(out[14]) );
  DFF_X2 \u6/quo1_reg[23]  ( .D(\u6/N23 ), .CK(clk), .Q(\u6/quo1 [23]) );
  DFF_X2 \u6/quo_reg[23]  ( .D(\u6/quo1 [23]), .CK(clk), .QN(net11485) );
  fpu_DW01_ash_1 \u4/sll_479  ( .A({net85786, net85786, net85786, net85786, 
        net85786, net85786, net85786, net85786, net85786, net86263, net77045, 
        net77161, n3003, net76254, net89624, n3002, n3004, net76672, n3005, 
        fract_denorm, net76926, net77073, net77637, net90292, net10316, n3001, 
        net76048, net90080, n3319}), .DATA_TC(1'b0), .SH({\u4/f2i_shft[4] , 
        \u4/f2i_shft[3] , \u4/f2i_shft[2] , net85710, net11564}), .SH_TC(1'b0), 
        .B({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, \u4/exp_f2i_1 , 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24}) );
  fpu_DW01_sub_7 \u3/sub_59  ( .A({1'b0, fracta}), .B({1'b0, fractb}), .CI(
        1'b0), .DIFF({\u3/N32 , \u3/N31 , \u3/N30 , \u3/N29 , \u3/N28 , 
        \u3/N27 , \u3/N26 , \u3/N25 , \u3/N24 , \u3/N23 , \u3/N22 , \u3/N21 , 
        \u3/N20 , \u3/N19 , \u3/N18 }) );
  fpu_DW01_add_5 \u3/add_59  ( .A({1'b0, fracta}), .B({1'b0, fractb}), .CI(
        1'b0), .SUM({\u3/N17 , \u3/N16 , \u3/N15 , \u3/N14 , \u3/N13 , 
        \u3/N12 , \u3/N11 , \u3/N10 , \u3/N9 , \u3/N8 , \u3/N7 , \u3/N6 , 
        \u3/N5 , \u3/N4 , \u3/N3 }) );
  fpu_DW01_ash_2 sll_385 ( .A({n3313, fracta_mul}), .DATA_TC(1'b0), .SH({N34, 
        N44, N56, N65}), .SH_TC(1'b0), .B({N77, N76, N75, N74, N73, N72, N71, 
        N70, N69, N68, N67}) );
  fpu_DW02_mult_0 \u5/mult_78  ( .A({n3313, fracta_mul[9:3], n2848, n3014, 
        n3015}), .B({\u6/N10 , \u6/N9 , \u6/N8 , \u6/N7 , \u6/N6 , \u6/N5 , 
        \u6/N4 , \u6/N3 , \u6/N2 , \u6/N1 , \u6/N0 }), .TC(1'b0), .PRODUCT({
        \u5/N21 , \u5/N20 , \u5/N19 , \u5/N18 , \u5/N17 , \u5/N16 , \u5/N15 , 
        \u5/N14 , \u5/N13 , \u5/N12 , \u5/N11 , \u5/N10 , \u5/N9 , \u5/N8 , 
        \u5/N7 , \u5/N6 , \u5/N5 , \u5/N4 , \u5/N3 , \u5/N2 , \u5/N1 , \u5/N0 }) );
  HA_X1 \u2/add_115/U1_1_1  ( .A(\u2/exp_tmp4[1] ), .B(\u2/exp_tmp4[0] ), .CO(
        \u2/add_115/carry [2]), .S(\u2/N31 ) );
  HA_X1 \u2/add_115/U1_1_2  ( .A(\u2/exp_tmp4[2] ), .B(\u2/add_115/carry [2]), 
        .CO(\u2/add_115/carry [3]), .S(\u2/N32 ) );
  HA_X1 \u2/add_115/U1_1_3  ( .A(\u2/exp_tmp4[3] ), .B(\u2/add_115/carry [3]), 
        .CO(\u2/add_115/carry [4]), .S(\u2/N33 ) );
  HA_X1 \u2/add_113/U1_1_1  ( .A(\u2/add_113/A[1] ), .B(\u2/add_113/A[0] ), 
        .CO(\u2/add_113/carry [2]), .S(\u2/exp_tmp3[1] ) );
  HA_X1 \u2/add_113/U1_1_2  ( .A(\u2/add_113/A[2] ), .B(\u2/add_113/carry [2]), 
        .CO(\u2/add_113/carry [3]), .S(\u2/exp_tmp3[2] ) );
  HA_X1 \u2/add_113/U1_1_3  ( .A(\u2/add_113/A[3] ), .B(\u2/add_113/carry [3]), 
        .CO(\u2/add_113/carry [4]), .S(\u2/exp_tmp3[3] ) );
  FA_X1 \u2/add_110/U1_1  ( .A(opa_r[11]), .B(opb_r[11]), .CI(
        \u2/add_110/carry [1]), .CO(\u2/add_110/carry [2]), .S(\u2/N13 ) );
  FA_X1 \u2/add_110/U1_2  ( .A(opa_r[12]), .B(opb_r[12]), .CI(
        \u2/add_110/carry [2]), .CO(\u2/add_110/carry [3]), .S(\u2/N14 ) );
  FA_X1 \u2/add_110/U1_3  ( .A(opa_r[13]), .B(opb_r[13]), .CI(
        \u2/add_110/carry [3]), .CO(\u2/add_110/carry [4]), .S(\u2/N15 ) );
  FA_X1 \u2/add_110/U1_4  ( .A(opa_r[14]), .B(n1733), .CI(
        \u2/add_110/carry [4]), .CO(\u2/N17 ), .S(\u2/N16 ) );
  FA_X1 \u2/sub_110/U2_1  ( .A(opa_r[11]), .B(n3016), .CI(
        \u2/sub_110/carry [1]), .CO(\u2/sub_110/carry [2]), .S(\u2/N7 ) );
  FA_X1 \u2/sub_110/U2_2  ( .A(opa_r[12]), .B(n2799), .CI(
        \u2/sub_110/carry [2]), .CO(\u2/sub_110/carry [3]), .S(\u2/N8 ) );
  FA_X1 \u2/sub_110/U2_3  ( .A(opa_r[13]), .B(n3017), .CI(
        \u2/sub_110/carry [3]), .CO(\u2/sub_110/carry [4]), .S(\u2/N9 ) );
  FA_X1 \u2/sub_110/U2_4  ( .A(opa_r[14]), .B(n1541), .CI(
        \u2/sub_110/carry [4]), .CO(\u2/sub_110/carry [5]), .S(\u2/N10 ) );
  fpu_DW01_inc_5 \u4/add_393  ( .A({1'b0, net91299, net90252, 
        \u4/fract_out[7] , net91512, n1528, net89933, net99874, n3006, n1920, 
        net60630}), .SUM({\u4/fract_out_pl1[10] , \u4/fract_out_pl1[9] , 
        \u4/fract_out_pl1[8] , \u4/fract_out_pl1[7] , \u4/fract_out_pl1[6] , 
        \u4/fract_out_pl1[5] , \u4/fract_out_pl1[4] , \u4/fract_out_pl1[3] , 
        \u4/fract_out_pl1[2] , \u4/fract_out_pl1[1] , \u4/fract_out_pl1[0] })
         );
  fpu_DW_rash_2 \u4/srl_450  ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, net85786, net86263, net91070, net90115, n3003, 
        net86004, net89624, n3002, n3004, net90007, n3005, fract_denorm[10], 
        net90211, net90037, n1883, net90290, n2998, net10316, n3001, n2999, 
        n1926, n3319}), .DATA_TC(1'b0), .SH(\u4/shift_right [2:0]), .SH_TC(
        1'b0), .B({SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, \u4/N409 , 
        \u4/N408 , \u4/N407 , \u4/N406 , \u4/N405 , \u4/N404 , \u4/N403 , 
        \u4/N402 , \u4/N401 , \u4/N400 , \u4/N399 , \u4/N398 , \u4/N397 , 
        \u4/N396 , \u4/N395 , \u4/N394 , \u4/N393 , \u4/N392 , \u4/N391 , 
        \u4/N390 , \u4/N389 , \u4/N388 }) );
  fpu_DW01_ash_4 \u4/sll_451  ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, net85786, net86263, net91070, net90115, n3003, 
        net86004, net89624, n3002, n3004, net90007, n3005, fract_denorm[10], 
        net90211, net90037, n1883, net90290, n2998, net10316, n3001, n2999, 
        n3000, n3319}), .DATA_TC(1'b0), .SH(\u4/shift_left ), .SH_TC(1'b0), 
        .B({SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, \u4/N433 , 
        \u4/N432 , \u4/N431 , \u4/N430 , \u4/N429 , \u4/N428 , \u4/N427 , 
        \u4/N426 , \u4/N425 , \u4/N424 , \u4/N423 , \u4/N422 , \u4/N421 , 
        \u4/N420 , \u4/N419 , \u4/N418 , \u4/N417 , \u4/N416 , \u4/N415 , 
        \u4/N414 , \u4/N413 , \u4/N412 }) );
  fpu_DW01_sub_23 \u4/sub_467  ( .A({1'b0, \u4/exp_in_pl1[5] , 
        \u4/exp_in_pl1[4] , \u4/exp_in_pl1[3] , \u4/exp_in_pl1[2] , net85712, 
        net15448}), .B({1'b0, 1'b0, n3008, \u4/fi_ldz_mi1[3] , 
        \u4/fi_ldz_mi1[2] , net33278, net89965}), .CI(1'b0), .DIFF({
        SYNOPSYS_UNCONNECTED__45, \u4/exp_next_mi[5] , \u4/exp_next_mi[4] , 
        \u4/exp_next_mi[3] , \u4/exp_next_mi[2] , \u4/exp_next_mi[1] , 
        \u4/exp_next_mi[0] }) );
  fpu_DW_rash_11 \u1/srl_146  ( .A({n1521, \u1/adj_op[9] , n3303, n3304, n3305, 
        n3306, n3307, n3308, n3309, n3310, n3311, 1'b0, 1'b0, 1'b0}), 
        .DATA_TC(1'b0), .SH({n3302, n3301, n3300, n1718}), .SH_TC(1'b0), .B({
=======
  DFF_X2 \u6/quo1_reg[23]  ( .D(\u6/N23 ), .CK(clk), .Q(\u6/quo1 [23]) );
  DFF_X2 \u6/quo_reg[23]  ( .D(\u6/quo1 [23]), .CK(clk), .Q(quo[23]) );
  DFF_X2 \u6/quo1_reg[24]  ( .D(\u6/N24 ), .CK(clk), .Q(\u6/quo1 [24]) );
  DFF_X2 \u6/quo_reg[24]  ( .D(\u6/quo1 [24]), .CK(clk), .Q(quo[24]) );
  DFF_X2 \u6/quo1_reg[25]  ( .D(\u6/N25 ), .CK(clk), .Q(\u6/quo1 [25]) );
  DFF_X2 \u6/quo_reg[25]  ( .D(\u6/quo1 [25]), .CK(clk), .Q(quo[25]) );
  DFF_X2 \u6/quo1_reg[26]  ( .D(\u6/N26 ), .CK(clk), .Q(\u6/quo1 [26]) );
  DFF_X2 \u6/quo_reg[26]  ( .D(\u6/quo1 [26]), .CK(clk), .Q(quo[26]) );
  DFF_X2 \u6/quo1_reg[27]  ( .D(\u6/N27 ), .CK(clk), .Q(\u6/quo1 [27]) );
  DFF_X2 \u6/quo_reg[27]  ( .D(\u6/quo1 [27]), .CK(clk), .Q(quo[27]) );
  DFF_X2 \u6/quo1_reg[28]  ( .D(\u6/N28 ), .CK(clk), .Q(\u6/quo1 [28]) );
  DFF_X2 \u6/quo_reg[28]  ( .D(\u6/quo1 [28]), .CK(clk), .Q(quo[28]) );
  DFF_X2 \u6/quo1_reg[29]  ( .D(\u6/N29 ), .CK(clk), .Q(\u6/quo1 [29]) );
  DFF_X2 \u6/quo_reg[29]  ( .D(\u6/quo1 [29]), .CK(clk), .Q(quo[29]) );
  DFF_X2 \u6/quo1_reg[30]  ( .D(\u6/N30 ), .CK(clk), .Q(\u6/quo1 [30]) );
  DFF_X2 \u6/quo_reg[30]  ( .D(\u6/quo1 [30]), .CK(clk), .Q(quo[30]) );
  DFF_X2 \u6/quo1_reg[31]  ( .D(\u6/N31 ), .CK(clk), .Q(\u6/quo1 [31]) );
  DFF_X2 \u6/quo_reg[31]  ( .D(\u6/quo1 [31]), .CK(clk), .Q(quo[31]) );
  DFF_X2 \u6/quo1_reg[32]  ( .D(\u6/N32 ), .CK(clk), .Q(\u6/quo1 [32]) );
  DFF_X2 \u6/quo_reg[32]  ( .D(\u6/quo1 [32]), .CK(clk), .Q(quo[32]) );
  DFF_X2 \u6/quo1_reg[33]  ( .D(\u6/N33 ), .CK(clk), .Q(\u6/quo1 [33]) );
  DFF_X2 \u6/quo_reg[33]  ( .D(\u6/quo1 [33]), .CK(clk), .Q(quo[33]) );
  DFF_X2 \u6/quo1_reg[34]  ( .D(\u6/N34 ), .CK(clk), .Q(\u6/quo1 [34]) );
  DFF_X2 \u6/quo_reg[34]  ( .D(\u6/quo1 [34]), .CK(clk), .Q(quo[34]) );
  DFF_X2 \u6/quo1_reg[35]  ( .D(\u6/N35 ), .CK(clk), .Q(\u6/quo1 [35]) );
  DFF_X2 \u6/quo_reg[35]  ( .D(\u6/quo1 [35]), .CK(clk), .Q(quo[35]) );
  DFF_X2 \u6/quo1_reg[36]  ( .D(\u6/N36 ), .CK(clk), .Q(\u6/quo1 [36]) );
  DFF_X2 \u6/quo_reg[36]  ( .D(\u6/quo1 [36]), .CK(clk), .Q(quo[36]) );
  DFF_X2 \u6/quo1_reg[37]  ( .D(\u6/N37 ), .CK(clk), .Q(\u6/quo1 [37]) );
  DFF_X2 \u6/quo_reg[37]  ( .D(\u6/quo1 [37]), .CK(clk), .Q(quo[37]) );
  DFF_X2 \u6/quo1_reg[38]  ( .D(\u6/N38 ), .CK(clk), .Q(\u6/quo1 [38]) );
  DFF_X2 \u6/quo_reg[38]  ( .D(\u6/quo1 [38]), .CK(clk), .Q(quo[38]) );
  DFF_X2 \u6/quo1_reg[39]  ( .D(\u6/N39 ), .CK(clk), .Q(\u6/quo1 [39]) );
  DFF_X2 \u6/quo_reg[39]  ( .D(\u6/quo1 [39]), .CK(clk), .Q(quo[39]) );
  DFF_X2 \u6/quo1_reg[40]  ( .D(\u6/N40 ), .CK(clk), .Q(\u6/quo1 [40]) );
  DFF_X2 \u6/quo_reg[40]  ( .D(\u6/quo1 [40]), .CK(clk), .Q(quo[40]) );
  DFF_X2 \u6/quo1_reg[41]  ( .D(\u6/N41 ), .CK(clk), .Q(\u6/quo1 [41]) );
  DFF_X2 \u6/quo_reg[41]  ( .D(\u6/quo1 [41]), .CK(clk), .Q(quo[41]) );
  DFF_X2 \u6/quo1_reg[42]  ( .D(\u6/N42 ), .CK(clk), .Q(\u6/quo1 [42]) );
  DFF_X2 \u6/quo_reg[42]  ( .D(\u6/quo1 [42]), .CK(clk), .Q(quo[42]) );
  DFF_X2 \u6/quo1_reg[43]  ( .D(\u6/N43 ), .CK(clk), .Q(\u6/quo1 [43]) );
  DFF_X2 \u6/quo_reg[43]  ( .D(\u6/quo1 [43]), .CK(clk), .Q(quo[43]) );
  DFF_X2 \u6/quo1_reg[44]  ( .D(\u6/N44 ), .CK(clk), .Q(\u6/quo1 [44]) );
  DFF_X2 \u6/quo_reg[44]  ( .D(\u6/quo1 [44]), .CK(clk), .Q(quo[44]) );
  DFF_X2 \u6/quo1_reg[45]  ( .D(\u6/N45 ), .CK(clk), .Q(\u6/quo1 [45]) );
  DFF_X2 \u6/quo_reg[45]  ( .D(\u6/quo1 [45]), .CK(clk), .Q(quo[45]) );
  DFF_X2 \u6/quo1_reg[46]  ( .D(\u6/N46 ), .CK(clk), .Q(\u6/quo1 [46]) );
  DFF_X2 \u6/quo_reg[46]  ( .D(\u6/quo1 [46]), .CK(clk), .Q(quo[46]) );
  DFF_X2 \u6/quo1_reg[47]  ( .D(\u6/N47 ), .CK(clk), .Q(\u6/quo1 [47]) );
  DFF_X2 \u6/quo_reg[47]  ( .D(\u6/quo1 [47]), .CK(clk), .Q(quo[47]) );
  DFF_X2 \u6/quo1_reg[48]  ( .D(\u6/N48 ), .CK(clk), .Q(\u6/quo1 [48]) );
  DFF_X2 \u6/quo_reg[48]  ( .D(\u6/quo1 [48]), .CK(clk), .Q(quo[48]) );
  DFF_X2 \u6/quo1_reg[49]  ( .D(\u6/N49 ), .CK(clk), .Q(\u6/quo1 [49]) );
  DFF_X2 \u6/quo_reg[49]  ( .D(\u6/quo1 [49]), .CK(clk), .Q(quo[49]) );
  DFF_X2 \u6/quo1_reg[50]  ( .D(\u6/N50 ), .CK(clk), .Q(\u6/quo1 [50]) );
  DFF_X2 \u6/quo_reg[50]  ( .D(\u6/quo1 [50]), .CK(clk), .Q(quo[50]) );
  DFF_X2 \u6/quo1_reg[51]  ( .D(\u6/N51 ), .CK(clk), .Q(\u6/quo1 [51]) );
  DFF_X2 \u6/quo_reg[51]  ( .D(\u6/quo1 [51]), .CK(clk), .Q(quo[51]) );
  DFF_X2 \u6/quo1_reg[52]  ( .D(\u6/N52 ), .CK(clk), .Q(\u6/quo1 [52]) );
  DFF_X2 \u6/quo_reg[52]  ( .D(\u6/quo1 [52]), .CK(clk), .Q(quo[52]) );
  DFF_X2 \u6/quo1_reg[55]  ( .D(\u6/N55 ), .CK(clk), .Q(\u6/quo1 [55]) );
  DFF_X2 \u6/quo_reg[55]  ( .D(\u6/quo1 [55]), .CK(clk), .Q(quo[55]), .QN(
        n4398) );
  DFF_X2 \u6/quo1_reg[56]  ( .D(\u6/N56 ), .CK(clk), .Q(\u6/quo1 [56]) );
  DFF_X2 \u6/quo_reg[56]  ( .D(\u6/quo1 [56]), .CK(clk), .Q(quo[56]) );
  DFF_X2 \u6/quo1_reg[57]  ( .D(\u6/N57 ), .CK(clk), .Q(\u6/quo1 [57]) );
  DFF_X2 \u6/quo_reg[57]  ( .D(\u6/quo1 [57]), .CK(clk), .Q(quo[57]) );
  DFF_X2 \u6/quo1_reg[58]  ( .D(\u6/N58 ), .CK(clk), .Q(\u6/quo1 [58]) );
  DFF_X2 \u6/quo_reg[58]  ( .D(\u6/quo1 [58]), .CK(clk), .Q(quo[58]) );
  DFF_X2 \u6/quo1_reg[59]  ( .D(\u6/N59 ), .CK(clk), .Q(\u6/quo1 [59]) );
  DFF_X2 \u6/quo_reg[59]  ( .D(\u6/quo1 [59]), .CK(clk), .Q(quo[59]) );
  DFF_X2 \u6/quo1_reg[60]  ( .D(\u6/N60 ), .CK(clk), .Q(\u6/quo1 [60]) );
  DFF_X2 \u6/quo_reg[60]  ( .D(\u6/quo1 [60]), .CK(clk), .Q(quo[60]) );
  DFF_X2 \u6/quo1_reg[61]  ( .D(\u6/N61 ), .CK(clk), .Q(\u6/quo1 [61]) );
  DFF_X2 \u6/quo_reg[61]  ( .D(\u6/quo1 [61]), .CK(clk), .Q(quo[61]) );
  DFF_X2 \u6/quo1_reg[62]  ( .D(\u6/N62 ), .CK(clk), .Q(\u6/quo1 [62]) );
  DFF_X2 \u6/quo_reg[62]  ( .D(\u6/quo1 [62]), .CK(clk), .Q(quo[62]) );
  DFF_X2 \u6/quo1_reg[63]  ( .D(\u6/N63 ), .CK(clk), .Q(\u6/quo1 [63]) );
  DFF_X2 \u6/quo_reg[63]  ( .D(\u6/quo1 [63]), .CK(clk), .Q(quo[63]) );
  DFF_X2 \u6/quo1_reg[64]  ( .D(\u6/N64 ), .CK(clk), .Q(\u6/quo1 [64]) );
  DFF_X2 \u6/quo_reg[64]  ( .D(\u6/quo1 [64]), .CK(clk), .Q(quo[64]) );
  DFF_X2 \u6/quo1_reg[65]  ( .D(\u6/N65 ), .CK(clk), .Q(\u6/quo1 [65]) );
  DFF_X2 \u6/quo_reg[65]  ( .D(\u6/quo1 [65]), .CK(clk), .Q(quo[65]) );
  DFF_X2 \u6/quo1_reg[66]  ( .D(\u6/N66 ), .CK(clk), .Q(\u6/quo1 [66]) );
  DFF_X2 \u6/quo_reg[66]  ( .D(\u6/quo1 [66]), .CK(clk), .Q(quo[66]) );
  DFF_X2 \u6/quo1_reg[67]  ( .D(\u6/N67 ), .CK(clk), .Q(\u6/quo1 [67]) );
  DFF_X2 \u6/quo_reg[67]  ( .D(\u6/quo1 [67]), .CK(clk), .Q(quo[67]) );
  DFF_X2 \u6/quo1_reg[68]  ( .D(\u6/N68 ), .CK(clk), .Q(\u6/quo1 [68]) );
  DFF_X2 \u6/quo_reg[68]  ( .D(\u6/quo1 [68]), .CK(clk), .Q(quo[68]) );
  DFF_X2 \u6/quo1_reg[69]  ( .D(\u6/N69 ), .CK(clk), .Q(\u6/quo1 [69]) );
  DFF_X2 \u6/quo_reg[69]  ( .D(\u6/quo1 [69]), .CK(clk), .Q(quo[69]) );
  DFF_X2 \u6/quo1_reg[70]  ( .D(\u6/N70 ), .CK(clk), .Q(\u6/quo1 [70]) );
  DFF_X2 \u6/quo_reg[70]  ( .D(\u6/quo1 [70]), .CK(clk), .Q(quo[70]) );
  DFF_X2 \u6/quo1_reg[71]  ( .D(\u6/N71 ), .CK(clk), .Q(\u6/quo1 [71]) );
  DFF_X2 \u6/quo_reg[71]  ( .D(\u6/quo1 [71]), .CK(clk), .Q(quo[71]) );
  DFF_X2 \u6/quo1_reg[72]  ( .D(\u6/N72 ), .CK(clk), .Q(\u6/quo1 [72]) );
  DFF_X2 \u6/quo_reg[72]  ( .D(\u6/quo1 [72]), .CK(clk), .Q(quo[72]) );
  DFF_X2 \u6/quo1_reg[73]  ( .D(\u6/N73 ), .CK(clk), .Q(\u6/quo1 [73]) );
  DFF_X2 \u6/quo_reg[73]  ( .D(\u6/quo1 [73]), .CK(clk), .Q(quo[73]) );
  DFF_X2 \u6/quo1_reg[74]  ( .D(\u6/N74 ), .CK(clk), .Q(\u6/quo1 [74]) );
  DFF_X2 \u6/quo_reg[74]  ( .D(\u6/quo1 [74]), .CK(clk), .Q(quo[74]) );
  DFF_X2 \u6/quo1_reg[75]  ( .D(\u6/N75 ), .CK(clk), .Q(\u6/quo1 [75]) );
  DFF_X2 \u6/quo_reg[75]  ( .D(\u6/quo1 [75]), .CK(clk), .Q(quo[75]) );
  DFF_X2 \u6/quo1_reg[76]  ( .D(\u6/N76 ), .CK(clk), .Q(\u6/quo1 [76]) );
  DFF_X2 \u6/quo_reg[76]  ( .D(\u6/quo1 [76]), .CK(clk), .Q(quo[76]) );
  DFF_X2 \u6/quo1_reg[77]  ( .D(\u6/N77 ), .CK(clk), .Q(\u6/quo1 [77]) );
  DFF_X2 \u6/quo_reg[77]  ( .D(\u6/quo1 [77]), .CK(clk), .Q(quo[77]) );
  DFF_X2 \u6/quo1_reg[78]  ( .D(\u6/N78 ), .CK(clk), .Q(\u6/quo1 [78]) );
  DFF_X2 \u6/quo_reg[78]  ( .D(\u6/quo1 [78]), .CK(clk), .Q(quo[78]) );
  DFF_X2 \u6/quo1_reg[79]  ( .D(\u6/N79 ), .CK(clk), .Q(\u6/quo1 [79]) );
  DFF_X2 \u6/quo_reg[79]  ( .D(\u6/quo1 [79]), .CK(clk), .Q(quo[79]) );
  DFF_X2 \u6/quo1_reg[80]  ( .D(\u6/N80 ), .CK(clk), .Q(\u6/quo1 [80]) );
  DFF_X2 \u6/quo_reg[80]  ( .D(\u6/quo1 [80]), .CK(clk), .Q(quo[80]) );
  DFF_X2 \u6/quo1_reg[81]  ( .D(\u6/N81 ), .CK(clk), .Q(\u6/quo1 [81]) );
  DFF_X2 \u6/quo_reg[81]  ( .D(\u6/quo1 [81]), .CK(clk), .Q(quo[81]) );
  DFF_X2 \u6/quo1_reg[82]  ( .D(\u6/N82 ), .CK(clk), .Q(\u6/quo1 [82]) );
  DFF_X2 \u6/quo_reg[82]  ( .D(\u6/quo1 [82]), .CK(clk), .Q(quo[82]) );
  DFF_X2 \u6/quo1_reg[83]  ( .D(\u6/N83 ), .CK(clk), .Q(\u6/quo1 [83]) );
  DFF_X2 \u6/quo_reg[83]  ( .D(\u6/quo1 [83]), .CK(clk), .Q(quo[83]) );
  DFF_X2 \u6/quo1_reg[84]  ( .D(\u6/N84 ), .CK(clk), .Q(\u6/quo1 [84]) );
  DFF_X2 \u6/quo_reg[84]  ( .D(\u6/quo1 [84]), .CK(clk), .Q(quo[84]) );
  DFF_X2 \u6/quo1_reg[85]  ( .D(\u6/N85 ), .CK(clk), .Q(\u6/quo1 [85]) );
  DFF_X2 \u6/quo_reg[85]  ( .D(\u6/quo1 [85]), .CK(clk), .Q(quo[85]) );
  DFF_X2 \u6/quo1_reg[86]  ( .D(\u6/N86 ), .CK(clk), .Q(\u6/quo1 [86]) );
  DFF_X2 \u6/quo_reg[86]  ( .D(\u6/quo1 [86]), .CK(clk), .Q(quo[86]) );
  DFF_X2 \u6/quo1_reg[87]  ( .D(\u6/N87 ), .CK(clk), .Q(\u6/quo1 [87]) );
  DFF_X2 \u6/quo_reg[87]  ( .D(\u6/quo1 [87]), .CK(clk), .Q(quo[87]) );
  DFF_X2 \u6/quo1_reg[88]  ( .D(\u6/N88 ), .CK(clk), .Q(\u6/quo1 [88]) );
  DFF_X2 \u6/quo_reg[88]  ( .D(\u6/quo1 [88]), .CK(clk), .Q(quo[88]) );
  DFF_X2 \u6/quo1_reg[89]  ( .D(\u6/N89 ), .CK(clk), .Q(\u6/quo1 [89]) );
  DFF_X2 \u6/quo_reg[89]  ( .D(\u6/quo1 [89]), .CK(clk), .Q(quo[89]) );
  DFF_X2 \u6/quo1_reg[90]  ( .D(\u6/N90 ), .CK(clk), .Q(\u6/quo1 [90]) );
  DFF_X2 \u6/quo_reg[90]  ( .D(\u6/quo1 [90]), .CK(clk), .Q(quo[90]) );
  DFF_X2 \u6/quo1_reg[91]  ( .D(\u6/N91 ), .CK(clk), .Q(\u6/quo1 [91]) );
  DFF_X2 \u6/quo_reg[91]  ( .D(\u6/quo1 [91]), .CK(clk), .Q(quo[91]) );
  DFF_X2 \u6/quo1_reg[92]  ( .D(\u6/N92 ), .CK(clk), .Q(\u6/quo1 [92]) );
  DFF_X2 \u6/quo_reg[92]  ( .D(\u6/quo1 [92]), .CK(clk), .Q(quo[92]) );
  DFF_X2 \u6/quo1_reg[93]  ( .D(\u6/N93 ), .CK(clk), .Q(\u6/quo1 [93]) );
  DFF_X2 \u6/quo_reg[93]  ( .D(\u6/quo1 [93]), .CK(clk), .Q(quo[93]) );
  DFF_X2 \u6/quo1_reg[94]  ( .D(\u6/N94 ), .CK(clk), .Q(\u6/quo1 [94]) );
  DFF_X2 \u6/quo_reg[94]  ( .D(\u6/quo1 [94]), .CK(clk), .Q(quo[94]) );
  DFF_X2 \u6/quo1_reg[95]  ( .D(\u6/N95 ), .CK(clk), .Q(\u6/quo1 [95]) );
  DFF_X2 \u6/quo_reg[95]  ( .D(\u6/quo1 [95]), .CK(clk), .Q(quo[95]) );
  DFF_X2 \u6/quo1_reg[96]  ( .D(\u6/N96 ), .CK(clk), .Q(\u6/quo1 [96]) );
  DFF_X2 \u6/quo_reg[96]  ( .D(\u6/quo1 [96]), .CK(clk), .Q(quo[96]) );
  DFF_X2 \u6/quo1_reg[97]  ( .D(\u6/N97 ), .CK(clk), .Q(\u6/quo1 [97]) );
  DFF_X2 \u6/quo_reg[97]  ( .D(\u6/quo1 [97]), .CK(clk), .Q(quo[97]) );
  DFF_X2 \u6/quo1_reg[98]  ( .D(\u6/N98 ), .CK(clk), .Q(\u6/quo1 [98]) );
  DFF_X2 \u6/quo_reg[98]  ( .D(\u6/quo1 [98]), .CK(clk), .Q(quo[98]) );
  DFF_X2 \u6/quo1_reg[99]  ( .D(\u6/N99 ), .CK(clk), .Q(\u6/quo1 [99]) );
  DFF_X2 \u6/quo_reg[99]  ( .D(\u6/quo1 [99]), .CK(clk), .Q(quo[99]) );
  DFF_X2 \u6/quo1_reg[100]  ( .D(\u6/N100 ), .CK(clk), .Q(\u6/quo1 [100]) );
  DFF_X2 \u6/quo_reg[100]  ( .D(\u6/quo1 [100]), .CK(clk), .Q(quo[100]) );
  DFF_X2 \u6/quo1_reg[101]  ( .D(\u6/N101 ), .CK(clk), .Q(\u6/quo1 [101]) );
  DFF_X2 \u6/quo_reg[101]  ( .D(\u6/quo1 [101]), .CK(clk), .Q(quo[101]) );
  DFF_X2 \u6/quo1_reg[102]  ( .D(\u6/N102 ), .CK(clk), .Q(\u6/quo1 [102]) );
  DFF_X2 \u6/quo_reg[102]  ( .D(\u6/quo1 [102]), .CK(clk), .Q(quo[102]) );
  DFF_X2 \u6/quo1_reg[103]  ( .D(\u6/N103 ), .CK(clk), .Q(\u6/quo1 [103]) );
  DFF_X2 \u6/quo_reg[103]  ( .D(\u6/quo1 [103]), .CK(clk), .Q(quo[103]) );
  DFF_X2 \u6/quo1_reg[104]  ( .D(\u6/N104 ), .CK(clk), .Q(\u6/quo1 [104]) );
  DFF_X2 \u6/quo_reg[104]  ( .D(\u6/quo1 [104]), .CK(clk), .Q(quo[104]) );
  DFF_X2 \u6/quo1_reg[105]  ( .D(\u6/N105 ), .CK(clk), .Q(\u6/quo1 [105]) );
  DFF_X2 \u6/quo_reg[105]  ( .D(\u6/quo1 [105]), .CK(clk), .Q(quo[105]) );
  DFF_X2 \u6/quo1_reg[106]  ( .D(\u6/N106 ), .CK(clk), .Q(\u6/quo1 [106]) );
  DFF_X2 \u6/quo_reg[106]  ( .D(\u6/quo1 [106]), .CK(clk), .Q(quo[106]) );
  DFF_X2 \out_reg[55]  ( .D(N848), .CK(clk), .Q(out[55]) );
  DFF_X2 \out_reg[56]  ( .D(N849), .CK(clk), .Q(out[56]) );
  DFF_X2 \out_reg[54]  ( .D(N847), .CK(clk), .Q(out[54]) );
  DFF_X2 \out_reg[57]  ( .D(N850), .CK(clk), .Q(out[57]) );
  DFF_X2 \out_reg[59]  ( .D(N852), .CK(clk), .Q(out[59]) );
  DFF_X2 \out_reg[58]  ( .D(N851), .CK(clk), .Q(out[58]) );
  DFF_X2 \out_reg[53]  ( .D(N846), .CK(clk), .Q(out[53]) );
  DFF_X2 \out_reg[52]  ( .D(N845), .CK(clk), .Q(out[52]) );
  DFF_X2 \out_reg[62]  ( .D(N855), .CK(clk), .Q(out[62]) );
  DFF_X2 \out_reg[61]  ( .D(N854), .CK(clk), .Q(out[61]) );
  DFF_X2 \out_reg[60]  ( .D(N853), .CK(clk), .Q(out[60]) );
  DFF_X2 overflow_reg ( .D(N899), .CK(clk), .Q(overflow) );
  DFF_X2 \out_reg[51]  ( .D(N844), .CK(clk), .Q(out[51]) );
  DFF_X2 \out_reg[50]  ( .D(N843), .CK(clk), .Q(out[50]) );
  DFF_X2 \out_reg[49]  ( .D(N842), .CK(clk), .Q(out[49]) );
  DFF_X2 \out_reg[48]  ( .D(N841), .CK(clk), .Q(out[48]) );
  DFF_X2 \out_reg[47]  ( .D(N840), .CK(clk), .Q(out[47]) );
  DFF_X2 \out_reg[46]  ( .D(N839), .CK(clk), .Q(out[46]) );
  DFF_X2 \out_reg[45]  ( .D(N838), .CK(clk), .Q(out[45]) );
  DFF_X2 \out_reg[44]  ( .D(N837), .CK(clk), .Q(out[44]) );
  DFF_X2 \out_reg[43]  ( .D(N836), .CK(clk), .Q(out[43]) );
  DFF_X2 \out_reg[42]  ( .D(N835), .CK(clk), .Q(out[42]) );
  DFF_X2 \out_reg[41]  ( .D(N834), .CK(clk), .Q(out[41]) );
  DFF_X2 \out_reg[40]  ( .D(N833), .CK(clk), .Q(out[40]) );
  DFF_X2 \out_reg[39]  ( .D(N832), .CK(clk), .Q(out[39]) );
  DFF_X2 \out_reg[38]  ( .D(N831), .CK(clk), .Q(out[38]) );
  DFF_X2 \out_reg[37]  ( .D(N830), .CK(clk), .Q(out[37]) );
  DFF_X2 \out_reg[36]  ( .D(N829), .CK(clk), .Q(out[36]) );
  DFF_X2 \out_reg[35]  ( .D(N828), .CK(clk), .Q(out[35]) );
  DFF_X2 \out_reg[34]  ( .D(N827), .CK(clk), .Q(out[34]) );
  DFF_X2 \out_reg[33]  ( .D(N826), .CK(clk), .Q(out[33]) );
  DFF_X2 \out_reg[32]  ( .D(N825), .CK(clk), .Q(out[32]) );
  DFF_X2 \out_reg[31]  ( .D(N824), .CK(clk), .Q(out[31]) );
  DFF_X2 \out_reg[30]  ( .D(N823), .CK(clk), .Q(out[30]) );
  DFF_X2 \out_reg[29]  ( .D(N822), .CK(clk), .Q(out[29]) );
  DFF_X2 \out_reg[28]  ( .D(N821), .CK(clk), .Q(out[28]) );
  DFF_X2 \out_reg[27]  ( .D(N820), .CK(clk), .Q(out[27]) );
  DFF_X2 \out_reg[26]  ( .D(N819), .CK(clk), .Q(out[26]) );
  DFF_X2 \out_reg[25]  ( .D(N818), .CK(clk), .Q(out[25]) );
  DFF_X2 \out_reg[24]  ( .D(N817), .CK(clk), .Q(out[24]) );
  DFF_X2 \out_reg[23]  ( .D(N816), .CK(clk), .Q(out[23]) );
  DFF_X2 \out_reg[22]  ( .D(N815), .CK(clk), .Q(out[22]) );
  DFF_X2 \out_reg[21]  ( .D(N814), .CK(clk), .Q(out[21]) );
  DFF_X2 \out_reg[20]  ( .D(N813), .CK(clk), .Q(out[20]) );
  DFF_X2 \out_reg[19]  ( .D(N812), .CK(clk), .Q(out[19]) );
  DFF_X2 \out_reg[18]  ( .D(N811), .CK(clk), .Q(out[18]) );
  DFF_X2 \out_reg[17]  ( .D(N810), .CK(clk), .Q(out[17]) );
  DFF_X2 \out_reg[16]  ( .D(N809), .CK(clk), .Q(out[16]) );
  DFF_X2 \out_reg[15]  ( .D(N808), .CK(clk), .Q(out[15]) );
  DFF_X2 \out_reg[14]  ( .D(N807), .CK(clk), .Q(out[14]) );
  DFF_X2 \out_reg[13]  ( .D(N806), .CK(clk), .Q(out[13]) );
  DFF_X2 \out_reg[12]  ( .D(N805), .CK(clk), .Q(out[12]) );
  DFF_X2 \out_reg[11]  ( .D(N804), .CK(clk), .Q(out[11]) );
  DFF_X2 \out_reg[10]  ( .D(N803), .CK(clk), .Q(out[10]) );
  DFF_X2 \out_reg[9]  ( .D(N802), .CK(clk), .Q(out[9]) );
  DFF_X2 \out_reg[8]  ( .D(N801), .CK(clk), .Q(out[8]) );
  DFF_X2 \out_reg[7]  ( .D(N800), .CK(clk), .Q(out[7]) );
  DFF_X2 \out_reg[6]  ( .D(N799), .CK(clk), .Q(out[6]) );
  DFF_X2 \out_reg[5]  ( .D(N798), .CK(clk), .Q(out[5]) );
  DFF_X2 \out_reg[4]  ( .D(N797), .CK(clk), .Q(out[4]) );
  DFF_X2 \out_reg[3]  ( .D(N796), .CK(clk), .Q(out[3]) );
  DFF_X2 \out_reg[2]  ( .D(N795), .CK(clk), .Q(out[2]) );
  DFF_X2 \out_reg[1]  ( .D(N794), .CK(clk), .Q(out[1]) );
  DFF_X2 inf_reg ( .D(N906), .CK(clk), .Q(inf) );
  DFF_X2 underflow_reg ( .D(N902), .CK(clk), .Q(underflow) );
  DFF_X2 ine_reg ( .D(N889), .CK(clk), .Q(ine) );
  DFF_X2 zero_reg ( .D(N911), .CK(clk), .Q(zero) );
  DFF_X2 \out_reg[63]  ( .D(N875), .CK(clk), .Q(out[63]) );
  DFF_X2 \out_reg[0]  ( .D(N793), .CK(clk), .Q(out[0]) );
  DFF_X2 \u6/quo1_reg[107]  ( .D(\u6/N107 ), .CK(clk), .Q(\u6/quo1 [107]) );
  DFF_X2 \u6/quo_reg[107]  ( .D(\u6/quo1 [107]), .CK(clk), .Q(quo[107]) );
  fpu_DW01_sub_0 \u4/sub_473  ( .A({n4656, n4289, n4353, n4281, exp_r[6], 
        n4290, n4282, n4655, n4315, exp_r[1], n4600}), .B({1'b0, 1'b0, 1'b0, 
        1'b0, \u4/fi_ldz_mi1[6] , \u4/fi_ldz_mi1[5] , \u4/fi_ldz_mi1[4] , 
        \u4/fi_ldz_mi1[3] , \u4/fi_ldz_mi1[2] , \u4/fi_ldz_mi1[1] , 
        \u4/fi_ldz_mi1[0] }), .CI(1'b0), .DIFF(\u4/exp_fix_divb ) );
  fpu_DW01_sub_1 \u4/sub_472  ( .A({n4656, n4289, n4353, n4281, exp_r[6], 
        n4290, n4282, n4655, n4315, exp_r[1], n4600}), .B({1'b0, 1'b0, 1'b0, 
        1'b0, \u4/fi_ldz_mi22 , \u4/fi_ldz_mi1[0] }), .CI(1'b0), .DIFF(
        \u4/exp_fix_diva ) );
  fpu_DW01_inc_0 \u4/add_464  ( .A({\u4/exp_out[10] , \u4/exp_out[9] , 
        \u4/exp_out[8] , \u4/exp_out[7] , \u4/exp_out[6] , \u4/exp_out[5] , 
        \u4/exp_out[4] , \u4/exp_out[3] , \u4/exp_out[2] , \u4/exp_out[1] , 
        \u4/exp_out[0] }), .SUM({\u4/exp_out_pl1[10] , \u4/exp_out_pl1[9] , 
        \u4/exp_out_pl1[8] , \u4/exp_out_pl1[7] , \u4/exp_out_pl1[6] , 
        \u4/exp_out_pl1[5] , \u4/exp_out_pl1[4] , \u4/exp_out_pl1[3] , 
        \u4/exp_out_pl1[2] , \u4/exp_out_pl1[1] , \u4/exp_out_pl1[0] }) );
  fpu_DW01_ash_0 \u4/sll_454  ( .A({fract_denorm, n6367, n6409, n6410, n6408, 
        n6407, n6406, n6405, n6445, n6438, n6437, n6439, n6436, n6435, n6434, 
        n6433, n6440, n6431, n6430, n6432, n6429, n6428, n6427, n6426, n6441, 
        n6424, n6423, n6425, n6422, n6421, n6420, n6419, n6442, n6417, n6416, 
        n6418, n6415, n6414, n6413, n6411, n6443, n6444, n6351, n6350, n6349, 
        n6348, n6347, n6346, n6345, n6344, n6446}), .DATA_TC(1'b0), .SH(
        \u4/shift_left ), .SH_TC(1'b0), .B({\u4/N6119 , \u4/N6118 , \u4/N6117 , 
        \u4/N6116 , \u4/N6115 , \u4/N6114 , \u4/N6113 , \u4/N6112 , \u4/N6111 , 
        \u4/N6110 , \u4/N6109 , \u4/N6108 , \u4/N6107 , \u4/N6106 , \u4/N6105 , 
        \u4/N6104 , \u4/N6103 , \u4/N6102 , \u4/N6101 , \u4/N6100 , \u4/N6099 , 
        \u4/N6098 , \u4/N6097 , \u4/N6096 , \u4/N6095 , \u4/N6094 , \u4/N6093 , 
        \u4/N6092 , \u4/N6091 , \u4/N6090 , \u4/N6089 , \u4/N6088 , \u4/N6087 , 
        \u4/N6086 , \u4/N6085 , \u4/N6084 , \u4/N6083 , \u4/N6082 , \u4/N6081 , 
        \u4/N6080 , \u4/N6079 , \u4/N6078 , \u4/N6077 , \u4/N6076 , \u4/N6075 , 
        \u4/N6074 , \u4/N6073 , \u4/N6072 , \u4/N6071 , \u4/N6070 , \u4/N6069 , 
        \u4/N6068 , \u4/N6067 , \u4/N6066 , \u4/N6065 , \u4/N6064 , \u4/N6063 , 
        \u4/N6062 , \u4/N6061 , \u4/N6060 , \u4/N6059 , \u4/N6058 , \u4/N6057 , 
        \u4/N6056 , \u4/N6055 , \u4/N6054 , \u4/N6053 , \u4/N6052 , \u4/N6051 , 
        \u4/N6050 , \u4/N6049 , \u4/N6048 , \u4/N6047 , \u4/N6046 , \u4/N6045 , 
        \u4/N6044 , \u4/N6043 , \u4/N6042 , \u4/N6041 , \u4/N6040 , \u4/N6039 , 
        \u4/N6038 , \u4/N6037 , \u4/N6036 , \u4/N6035 , \u4/N6034 , \u4/N6033 , 
        \u4/N6032 , \u4/N6031 , \u4/N6030 , \u4/N6029 , \u4/N6028 , \u4/N6027 , 
        \u4/N6026 , \u4/N6025 , \u4/N6024 , \u4/N6023 , \u4/N6022 , \u4/N6021 , 
        \u4/N6020 , \u4/N6019 , \u4/N6018 , \u4/N6017 , \u4/N6016 , \u4/N6015 , 
        \u4/N6014 }) );
  fpu_DW_rash_0 \u4/srl_453  ( .A({n4652, fract_denorm[104:50], n6367, n6409, 
        n6410, n6408, n6407, n6406, n6405, n6445, n6438, n6437, n6439, n6436, 
        n6435, n6434, n6433, n6440, n6431, n6430, n6432, n6429, n6428, n6427, 
        n6426, n6441, n6424, n6423, n6425, n6422, n6421, n6420, n6419, n6442, 
        n6417, n6416, n6418, n6415, n6414, n6413, n6411, n6443, n6444, n6351, 
        n6350, n6349, n6348, n6347, n6346, n6345, n6344, n6446}), .DATA_TC(
        1'b0), .SH(\u4/shift_right [8:0]), .SH_TC(1'b0), .B({\u4/N6011 , 
        \u4/N6010 , \u4/N6009 , \u4/N6008 , \u4/N6007 , \u4/N6006 , \u4/N6005 , 
        \u4/N6004 , \u4/N6003 , \u4/N6002 , \u4/N6001 , \u4/N6000 , \u4/N5999 , 
        \u4/N5998 , \u4/N5997 , \u4/N5996 , \u4/N5995 , \u4/N5994 , \u4/N5993 , 
        \u4/N5992 , \u4/N5991 , \u4/N5990 , \u4/N5989 , \u4/N5988 , \u4/N5987 , 
        \u4/N5986 , \u4/N5985 , \u4/N5984 , \u4/N5983 , \u4/N5982 , \u4/N5981 , 
        \u4/N5980 , \u4/N5979 , \u4/N5978 , \u4/N5977 , \u4/N5976 , \u4/N5975 , 
        \u4/N5974 , \u4/N5973 , \u4/N5972 , \u4/N5971 , \u4/N5970 , \u4/N5969 , 
        \u4/N5968 , \u4/N5967 , \u4/N5966 , \u4/N5965 , \u4/N5964 , \u4/N5963 , 
        \u4/N5962 , \u4/N5961 , \u4/N5960 , \u4/N5959 , \u4/N5958 , \u4/N5957 , 
        \u4/N5956 , \u4/N5955 , \u4/N5954 , \u4/N5953 , \u4/N5952 , \u4/N5951 , 
        \u4/N5950 , \u4/N5949 , \u4/N5948 , \u4/N5947 , \u4/N5946 , \u4/N5945 , 
        \u4/N5944 , \u4/N5943 , \u4/N5942 , \u4/N5941 , \u4/N5940 , \u4/N5939 , 
        \u4/N5938 , \u4/N5937 , \u4/N5936 , \u4/N5935 , \u4/N5934 , \u4/N5933 , 
        \u4/N5932 , \u4/N5931 , \u4/N5930 , \u4/N5929 , \u4/N5928 , \u4/N5927 , 
        \u4/N5926 , \u4/N5925 , \u4/N5924 , \u4/N5923 , \u4/N5922 , \u4/N5921 , 
        \u4/N5920 , \u4/N5919 , \u4/N5918 , \u4/N5917 , \u4/N5916 , \u4/N5915 , 
        \u4/N5914 , \u4/N5913 , \u4/N5912 , \u4/N5911 , \u4/N5910 , \u4/N5909 , 
        \u4/N5908 , \u4/N5907 , \u4/N5906 }) );
  fpu_DW01_ash_1 \u4/sll_482  ( .A({1'b0, 1'b0, 1'b0, 1'b0, fract_denorm[105], 
        fract_denorm[105], fract_denorm[105], fract_denorm[105], 
        fract_denorm[105], n4652, n4652, fract_denorm[105], fract_denorm, 
        n6367, n6409, n6410, n6408, n6407, n6406, n6405, n6445, n6438, n6437, 
        n6439, n6436, n6435, n6434, n6433, n6440, n6431, n6430, n6432, n6429, 
        n6428, n6427, n6426, n6441, n6424, n6423, n6425, n6422, n6421, n6420, 
        n6419, n6442, n6417, n6416, n6418, n6415, n6414, n6413, n6411, n6443, 
        n6444, n6351, n6350, n6349, n6348, n6347, n6346, n6345, n6344, n6446}), 
        .DATA_TC(1'b0), .SH({\u4/f2i_shft[10] , \u4/f2i_shft[9] , 
        \u4/f2i_shft[8] , \u4/f2i_shft[7] , \u4/f2i_shft[6] , \u4/f2i_shft[5] , 
        \u4/f2i_shft[4] , \u4/f2i_shft[3] , \u4/f2i_shft[2] , \u4/f2i_shft[1] , 
        n4349}), .SH_TC(1'b0), .B({\u4/exp_f2i_1 , SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, 
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, 
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, 
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, 
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, 
        SYNOPSYS_UNCONNECTED__61, SYNOPSYS_UNCONNECTED__62, 
        SYNOPSYS_UNCONNECTED__63, SYNOPSYS_UNCONNECTED__64, 
        SYNOPSYS_UNCONNECTED__65, SYNOPSYS_UNCONNECTED__66, 
        SYNOPSYS_UNCONNECTED__67, SYNOPSYS_UNCONNECTED__68, 
        SYNOPSYS_UNCONNECTED__69, SYNOPSYS_UNCONNECTED__70, 
        SYNOPSYS_UNCONNECTED__71, SYNOPSYS_UNCONNECTED__72, 
        SYNOPSYS_UNCONNECTED__73, SYNOPSYS_UNCONNECTED__74, 
        SYNOPSYS_UNCONNECTED__75, SYNOPSYS_UNCONNECTED__76, 
        SYNOPSYS_UNCONNECTED__77, SYNOPSYS_UNCONNECTED__78, 
        SYNOPSYS_UNCONNECTED__79, SYNOPSYS_UNCONNECTED__80, 
        SYNOPSYS_UNCONNECTED__81, SYNOPSYS_UNCONNECTED__82, 
        SYNOPSYS_UNCONNECTED__83, SYNOPSYS_UNCONNECTED__84, 
        SYNOPSYS_UNCONNECTED__85, SYNOPSYS_UNCONNECTED__86, 
        SYNOPSYS_UNCONNECTED__87, SYNOPSYS_UNCONNECTED__88, 
        SYNOPSYS_UNCONNECTED__89, SYNOPSYS_UNCONNECTED__90, 
        SYNOPSYS_UNCONNECTED__91, SYNOPSYS_UNCONNECTED__92, 
        SYNOPSYS_UNCONNECTED__93, SYNOPSYS_UNCONNECTED__94, 
        SYNOPSYS_UNCONNECTED__95, SYNOPSYS_UNCONNECTED__96, 
        SYNOPSYS_UNCONNECTED__97, SYNOPSYS_UNCONNECTED__98, 
        SYNOPSYS_UNCONNECTED__99, SYNOPSYS_UNCONNECTED__100, 
        SYNOPSYS_UNCONNECTED__101, SYNOPSYS_UNCONNECTED__102, 
        SYNOPSYS_UNCONNECTED__103, SYNOPSYS_UNCONNECTED__104, 
        SYNOPSYS_UNCONNECTED__105, SYNOPSYS_UNCONNECTED__106}) );
  fpu_DW01_sub_4 \u4/sub_470  ( .A({\u4/exp_in_pl1[11] , \u4/exp_in_pl1[10] , 
        \u4/exp_in_pl1[9] , \u4/exp_in_pl1[8] , \u4/exp_in_pl1[7] , 
        \u4/exp_in_pl1[6] , \u4/exp_in_pl1[5] , \u4/exp_in_pl1[4] , 
        \u4/exp_in_pl1[3] , \u4/exp_in_pl1[2] , \u4/exp_in_pl1[1] , 
        \u4/exp_in_pl1[0] }), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \u4/fi_ldz_mi1[6] , \u4/fi_ldz_mi1[5] , \u4/fi_ldz_mi1[4] , 
        \u4/fi_ldz_mi1[3] , \u4/fi_ldz_mi1[2] , \u4/fi_ldz_mi1[1] , 
        \u4/fi_ldz_mi1[0] }), .CI(1'b0), .DIFF({\u4/exp_next_mi[11] , 
        \u4/exp_next_mi[10] , \u4/exp_next_mi[9] , \u4/exp_next_mi[8] , 
        \u4/exp_next_mi[7] , \u4/exp_next_mi[6] , \u4/exp_next_mi[5] , 
        \u4/exp_next_mi[4] , \u4/exp_next_mi[3] , \u4/exp_next_mi[2] , 
        \u4/exp_next_mi[1] , \u4/exp_next_mi[0] }) );
  fpu_DW01_sub_5 \u4/sub_496  ( .A({\u4/exp_in_pl1[11] , \u4/exp_in_pl1[10] , 
        \u4/exp_in_pl1[9] , \u4/exp_in_pl1[8] , \u4/exp_in_pl1[7] , 
        \u4/exp_in_pl1[6] , \u4/exp_in_pl1[5] , \u4/exp_in_pl1[4] , 
        \u4/exp_in_pl1[3] , \u4/exp_in_pl1[2] , \u4/exp_in_pl1[1] , 
        \u4/exp_in_pl1[0] }), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \u4/ldz_all[6] , \u4/ldz_all[5] , \u4/ldz_all[4] , \u4/ldz_all[3] , 
        \u4/ldz_all[2] , \u4/ldz_all[1] , \u4/ldz_all[0] }), .CI(1'b0), .DIFF(
        {SYNOPSYS_UNCONNECTED__107, \u4/div_exp2[10] , \u4/div_exp2[9] , 
        \u4/div_exp2[8] , \u4/div_exp2[7] , \u4/div_exp2[6] , \u4/div_exp2[5] , 
        \u4/div_exp2[4] , \u4/div_exp2[3] , \u4/div_exp2[2] , \u4/div_exp2[1] , 
        \u4/div_exp2[0] }) );
  fpu_DW01_add_0 \u4/add_489  ( .A({1'b0, 1'b0, div_opa_ldz_r2}), .B({
        \u4/fi_ldz[6] , \u4/fi_ldz[5] , \u4/fi_ldz[4] , \u4/fi_ldz[3] , 
        \u4/fi_ldz[2] , \u4/fi_ldz[1] , \u4/fi_ldz_2a[0] }), .CI(1'b0), .SUM({
        \u4/ldz_all[6] , \u4/ldz_all[5] , \u4/ldz_all[4] , \u4/ldz_all[3] , 
        \u4/ldz_all[2] , \u4/ldz_all[1] , \u4/ldz_all[0] }) );
  fpu_DW01_inc_1 \u4/add_466  ( .A({1'b0, n4656, n4289, n4353, n4281, exp_r[6], 
        n4290, n4282, n4655, n4315, exp_r[1], n4600}), .SUM({
        \u4/exp_in_pl1[11] , \u4/exp_in_pl1[10] , \u4/exp_in_pl1[9] , 
        \u4/exp_in_pl1[8] , \u4/exp_in_pl1[7] , \u4/exp_in_pl1[6] , 
        \u4/exp_in_pl1[5] , \u4/exp_in_pl1[4] , \u4/exp_in_pl1[3] , 
        \u4/exp_in_pl1[2] , \u4/exp_in_pl1[1] , \u4/exp_in_pl1[0] }) );
  fpu_DW01_add_1 \u4/add_494  ( .A({\u4/exp_in_mi1[11] , \u4/exp_in_mi1[10] , 
        \u4/exp_in_mi1[9] , \u4/exp_in_mi1[8] , \u4/exp_in_mi1[7] , 
        \u4/exp_in_mi1[6] , \u4/exp_in_mi1[5] , \u4/exp_in_mi1[4] , 
        \u4/exp_in_mi1[3] , \u4/exp_in_mi1[2] , \u4/exp_in_mi1[1] , n4349}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, \u4/fi_ldz_2a[6] , \u4/fi_ldz_2a[6] , 
        \u4/fi_ldz_2a[5] , \u4/fi_ldz_2a[4] , \u4/fi_ldz_2a[3] , 
        \u4/fi_ldz_2a[2] , \u4/fi_ldz_2a[1] , \u4/fi_ldz_2a[0] }), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__108, \u4/div_exp1[10] , \u4/div_exp1[9] , 
        \u4/div_exp1[8] , \u4/div_exp1[7] , \u4/div_exp1[6] , \u4/div_exp1[5] , 
        \u4/div_exp1[4] , \u4/div_exp1[3] , \u4/div_exp1[2] , \u4/div_exp1[1] , 
        \u4/div_exp1[0] }) );
  fpu_DW01_inc_2 \u4/add_396  ( .A({1'b0, \u4/fract_out[51] , 
        \u4/fract_out[50] , \u4/fract_out[49] , \u4/fract_out[48] , 
        \u4/fract_out[47] , \u4/fract_out[46] , \u4/fract_out[45] , 
        \u4/fract_out[44] , \u4/fract_out[43] , \u4/fract_out[42] , 
        \u4/fract_out[41] , \u4/fract_out[40] , \u4/fract_out[39] , 
        \u4/fract_out[38] , \u4/fract_out[37] , \u4/fract_out[36] , 
        \u4/fract_out[35] , \u4/fract_out[34] , \u4/fract_out[33] , 
        \u4/fract_out[32] , \u4/fract_out[31] , \u4/fract_out[30] , 
        \u4/fract_out[29] , \u4/fract_out[28] , \u4/fract_out[27] , 
        \u4/fract_out[26] , \u4/fract_out[25] , \u4/fract_out[24] , 
        \u4/fract_out[23] , \u4/fract_out[22] , \u4/fract_out[21] , 
        \u4/fract_out[20] , \u4/fract_out[19] , \u4/fract_out[18] , 
        \u4/fract_out[17] , \u4/fract_out[16] , \u4/fract_out[15] , 
        \u4/fract_out[14] , \u4/fract_out[13] , \u4/fract_out[12] , 
        \u4/fract_out[11] , \u4/fract_out[10] , \u4/fract_out[9] , 
        \u4/fract_out[8] , \u4/fract_out[7] , \u4/fract_out[6] , 
        \u4/fract_out[5] , \u4/fract_out[4] , \u4/fract_out[3] , 
        \u4/fract_out[2] , \u4/fract_out[1] , \u4/fract_out[0] }), .SUM({
        \u4/fract_out_pl1[52] , \u4/fract_out_pl1[51] , \u4/fract_out_pl1[50] , 
        \u4/fract_out_pl1[49] , \u4/fract_out_pl1[48] , \u4/fract_out_pl1[47] , 
        \u4/fract_out_pl1[46] , \u4/fract_out_pl1[45] , \u4/fract_out_pl1[44] , 
        \u4/fract_out_pl1[43] , \u4/fract_out_pl1[42] , \u4/fract_out_pl1[41] , 
        \u4/fract_out_pl1[40] , \u4/fract_out_pl1[39] , \u4/fract_out_pl1[38] , 
        \u4/fract_out_pl1[37] , \u4/fract_out_pl1[36] , \u4/fract_out_pl1[35] , 
        \u4/fract_out_pl1[34] , \u4/fract_out_pl1[33] , \u4/fract_out_pl1[32] , 
        \u4/fract_out_pl1[31] , \u4/fract_out_pl1[30] , \u4/fract_out_pl1[29] , 
        \u4/fract_out_pl1[28] , \u4/fract_out_pl1[27] , \u4/fract_out_pl1[26] , 
        \u4/fract_out_pl1[25] , \u4/fract_out_pl1[24] , \u4/fract_out_pl1[23] , 
        \u4/fract_out_pl1[22] , \u4/fract_out_pl1[21] , \u4/fract_out_pl1[20] , 
        \u4/fract_out_pl1[19] , \u4/fract_out_pl1[18] , \u4/fract_out_pl1[17] , 
        \u4/fract_out_pl1[16] , \u4/fract_out_pl1[15] , \u4/fract_out_pl1[14] , 
        \u4/fract_out_pl1[13] , \u4/fract_out_pl1[12] , \u4/fract_out_pl1[11] , 
        \u4/fract_out_pl1[10] , \u4/fract_out_pl1[9] , \u4/fract_out_pl1[8] , 
        \u4/fract_out_pl1[7] , \u4/fract_out_pl1[6] , \u4/fract_out_pl1[5] , 
        \u4/fract_out_pl1[4] , \u4/fract_out_pl1[3] , \u4/fract_out_pl1[2] , 
        \u4/fract_out_pl1[1] , \u4/fract_out_pl1[0] }) );
  fpu_DW01_sub_9 \u3/sub_63  ( .A({1'b0, fracta}), .B({1'b0, fractb}), .CI(
        1'b0), .DIFF({\u3/N116 , \u3/N115 , \u3/N114 , \u3/N113 , \u3/N112 , 
        \u3/N111 , \u3/N110 , \u3/N109 , \u3/N108 , \u3/N107 , \u3/N106 , 
        \u3/N105 , \u3/N104 , \u3/N103 , \u3/N102 , \u3/N101 , \u3/N100 , 
        \u3/N99 , \u3/N98 , \u3/N97 , \u3/N96 , \u3/N95 , \u3/N94 , \u3/N93 , 
        \u3/N92 , \u3/N91 , \u3/N90 , \u3/N89 , \u3/N88 , \u3/N87 , \u3/N86 , 
        \u3/N85 , \u3/N84 , \u3/N83 , \u3/N82 , \u3/N81 , \u3/N80 , \u3/N79 , 
        \u3/N78 , \u3/N77 , \u3/N76 , \u3/N75 , \u3/N74 , \u3/N73 , \u3/N72 , 
        \u3/N71 , \u3/N70 , \u3/N69 , \u3/N68 , \u3/N67 , \u3/N66 , \u3/N65 , 
        \u3/N64 , \u3/N63 , \u3/N62 , \u3/N61 , \u3/N60 }) );
  fpu_DW01_add_4 \u3/add_63  ( .A({1'b0, fracta}), .B({1'b0, fractb}), .CI(
        1'b0), .SUM({\u3/N59 , \u3/N58 , \u3/N57 , \u3/N56 , \u3/N55 , 
        \u3/N54 , \u3/N53 , \u3/N52 , \u3/N51 , \u3/N50 , \u3/N49 , \u3/N48 , 
        \u3/N47 , \u3/N46 , \u3/N45 , \u3/N44 , \u3/N43 , \u3/N42 , \u3/N41 , 
        \u3/N40 , \u3/N39 , \u3/N38 , \u3/N37 , \u3/N36 , \u3/N35 , \u3/N34 , 
        \u3/N33 , \u3/N32 , \u3/N31 , \u3/N30 , \u3/N29 , \u3/N28 , \u3/N27 , 
        \u3/N26 , \u3/N25 , \u3/N24 , \u3/N23 , \u3/N22 , \u3/N21 , \u3/N20 , 
        \u3/N19 , \u3/N18 , \u3/N17 , \u3/N16 , \u3/N15 , \u3/N14 , \u3/N13 , 
        \u3/N12 , \u3/N11 , \u3/N10 , \u3/N9 , \u3/N8 , \u3/N7 , \u3/N6 , 
        \u3/N5 , \u3/N4 , \u3/N3 }) );
  fpu_DW01_inc_3 \u2/add_120  ( .A({\u2/exp_tmp4[10] , n2795, n2796, n2797, 
        n2798, n2799, \u2/exp_tmp4[4] , \u2/exp_tmp4[3] , \u2/exp_tmp4[2] , 
        \u2/exp_tmp4[1] , n2800}), .SUM({\u2/N64 , \u2/N63 , \u2/N62 , 
        \u2/N61 , \u2/N60 , \u2/N59 , \u2/N58 , \u2/N57 , \u2/N56 , \u2/N55 , 
        \u2/N54 }) );
  fpu_DW01_inc_4 \u2/add_118  ( .A({n6016, n6018, n6019, n6020, n6021, n6022, 
        n6023, n6025, n6027, n6029, n6031}), .SUM({\u2/exp_tmp3[10] , 
        \u2/exp_tmp3[9] , \u2/exp_tmp3[8] , \u2/exp_tmp3[7] , \u2/exp_tmp3[6] , 
        \u2/exp_tmp3[5] , \u2/exp_tmp3[4] , \u2/exp_tmp3[3] , \u2/exp_tmp3[2] , 
        \u2/exp_tmp3[1] , \u2/exp_tmp3[0] }) );
  fpu_DW01_add_6 \u2/add_115  ( .A({1'b0, opa_r[62:52]}), .B({1'b0, 
        opb_r[62:52]}), .CI(1'b0), .SUM({\u2/N29 , \u2/N28 , \u2/N27 , 
        \u2/N26 , \u2/N25 , \u2/N24 , \u2/N23 , \u2/N22 , \u2/N21 , \u2/N20 , 
        \u2/N19 , \u2/N18 }) );
  fpu_DW01_sub_12 \u2/sub_115  ( .A({1'b0, opa_r[62:52]}), .B({1'b0, 
        opb_r[62:52]}), .CI(1'b0), .DIFF({\u2/N17 , \u2/N16 , \u2/N15 , 
        \u2/N14 , \u2/N13 , \u2/N12 , \u2/N11 , \u2/N10 , \u2/N9 , \u2/N8 , 
        \u2/N7 , \u2/N6 }) );
  fpu_DW01_cmp2_13 \u1/gt_239  ( .A({n6158, n6159, n6160, n6161, n6162, n6163, 
        n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, 
        n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, 
        n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, 
        n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, 
        n6153, n6154, n6155, n6156, n6157, n6164, n6175, n6186, n6197, n6208}), 
        .B({n6105, n6106, n6107, n6108, n6109, n6110, n6112, n6113, n6114, 
        n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6123, n6124, n6125, 
        n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, 
        n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, 
        n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6100, n6101, n6102, 
        n6103, n6104, n6111, n6122, n6211, n6210, n6209}), .LEQ(1'b0), .TC(
        1'b0), .LT_LE(\u1/fractb_lt_fracta ) );
  fpu_DW_rash_1 \u1/srl_151  ( .A({n4266, \u1/adj_op[51] , n6234, n6236, n6237, 
        n6238, n6239, n6240, \u1/adj_op[44] , n6241, \u1/adj_op[42] , n6242, 
        n6243, n6244, \u1/adj_op[38] , \u1/adj_op[37] , \u1/adj_op[36] , n6245, 
        n6246, n6247, \u1/adj_op[32] , n6248, n6249, n6251, \u1/adj_op[28] , 
        \u1/adj_op[27] , n6252, n6253, n6254, n6255, \u1/adj_op[22] , 
        \u1/adj_op[21] , \u1/adj_op[20] , n6257, n6258, \u1/adj_op[17] , 
        \u1/adj_op[16] , \u1/adj_op[15] , n6259, n6260, n6261, \u1/adj_op[11] , 
        \u1/adj_op[10] , n6229, n6230, n6231, n6232, n6233, n6235, 
        \u1/adj_op[3] , n6250, n6256, \u1/adj_op[0] , 1'b0, 1'b0, 1'b0}), 
        .DATA_TC(1'b0), .SH({n6226, n6225, n6224, n6217, n6221, n6222}), 
        .SH_TC(1'b0), .B({\u1/adj_op_out_sft[55] , \u1/adj_op_out_sft[54] , 
        \u1/adj_op_out_sft[53] , \u1/adj_op_out_sft[52] , 
        \u1/adj_op_out_sft[51] , \u1/adj_op_out_sft[50] , 
        \u1/adj_op_out_sft[49] , \u1/adj_op_out_sft[48] , 
        \u1/adj_op_out_sft[47] , \u1/adj_op_out_sft[46] , 
        \u1/adj_op_out_sft[45] , \u1/adj_op_out_sft[44] , 
        \u1/adj_op_out_sft[43] , \u1/adj_op_out_sft[42] , 
        \u1/adj_op_out_sft[41] , \u1/adj_op_out_sft[40] , 
        \u1/adj_op_out_sft[39] , \u1/adj_op_out_sft[38] , 
        \u1/adj_op_out_sft[37] , \u1/adj_op_out_sft[36] , 
        \u1/adj_op_out_sft[35] , \u1/adj_op_out_sft[34] , 
        \u1/adj_op_out_sft[33] , \u1/adj_op_out_sft[32] , 
        \u1/adj_op_out_sft[31] , \u1/adj_op_out_sft[30] , 
        \u1/adj_op_out_sft[29] , \u1/adj_op_out_sft[28] , 
        \u1/adj_op_out_sft[27] , \u1/adj_op_out_sft[26] , 
        \u1/adj_op_out_sft[25] , \u1/adj_op_out_sft[24] , 
        \u1/adj_op_out_sft[23] , \u1/adj_op_out_sft[22] , 
        \u1/adj_op_out_sft[21] , \u1/adj_op_out_sft[20] , 
        \u1/adj_op_out_sft[19] , \u1/adj_op_out_sft[18] , 
        \u1/adj_op_out_sft[17] , \u1/adj_op_out_sft[16] , 
        \u1/adj_op_out_sft[15] , \u1/adj_op_out_sft[14] , 
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
        \u1/adj_op_out_sft[13] , \u1/adj_op_out_sft[12] , 
        \u1/adj_op_out_sft[11] , \u1/adj_op_out_sft[10] , 
        \u1/adj_op_out_sft[9] , \u1/adj_op_out_sft[8] , \u1/adj_op_out_sft[7] , 
        \u1/adj_op_out_sft[6] , \u1/adj_op_out_sft[5] , \u1/adj_op_out_sft[4] , 
        \u1/adj_op_out_sft[3] , \u1/adj_op_out_sft[2] , \u1/adj_op_out_sft[1] , 
        \u1/adj_op_out_sft[0] }) );
<<<<<<< HEAD
  DFF_X1 inf_reg ( .D(N285), .CK(clk), .Q(inf) );
  DFF_X1 \out_reg[4]  ( .D(N224), .CK(clk), .Q(out[4]) );
  DFF_X1 \out_reg[3]  ( .D(N223), .CK(clk), .Q(out[3]) );
  DFF_X1 \out_reg[2]  ( .D(N222), .CK(clk), .Q(out[2]) );
  DFF_X1 \out_reg[1]  ( .D(N221), .CK(clk), .Q(out[1]) );
  DFF_X1 \out_reg[5]  ( .D(N225), .CK(clk), .Q(out[5]) );
  DFF_X1 zero_reg ( .D(N290), .CK(clk), .Q(zero) );
  DFF_X1 ine_reg ( .D(n3007), .CK(clk), .Q(ine) );
  DFF_X1 underflow_reg ( .D(N281), .CK(clk), .Q(underflow) );
  DFF_X1 \out_reg[15]  ( .D(N254), .CK(clk), .Q(out[15]) );
  DFF_X2 \fract_i2f_reg[9]  ( .D(N184), .CK(clk), .QN(net90064) );
  DFF_X1 overflow_reg ( .D(N278), .CK(clk), .Q(overflow) );
  DFF_X1 \out_reg[6]  ( .D(N226), .CK(clk), .Q(out[6]) );
  DFF_X1 \out_reg[7]  ( .D(N227), .CK(clk), .Q(out[7]) );
  DFF_X1 \out_reg[8]  ( .D(N228), .CK(clk), .Q(out[8]) );
  DFF_X1 \out_reg[9]  ( .D(N229), .CK(clk), .Q(out[9]) );
  DFF_X1 \out_reg[12]  ( .D(N232), .CK(clk), .Q(out[12]) );
  DFF_X1 \u5/prod1_reg[13]  ( .D(\u5/N13 ), .CK(clk), .Q(\u5/prod1 [13]) );
  DFF_X1 \u5/prod1_reg[11]  ( .D(\u5/N11 ), .CK(clk), .Q(\u5/prod1 [11]) );
  DFF_X1 \u1/fracta_out_reg[5]  ( .D(\u1/fracta_s [5]), .CK(clk), .Q(fracta[5]) );
  DFF_X1 \u1/fractb_out_reg[13]  ( .D(\u1/fractb_s [13]), .CK(clk), .Q(
        fractb[13]) );
  DFF_X1 \u1/fractb_out_reg[10]  ( .D(\u1/fractb_s [10]), .CK(clk), .Q(
        fractb[10]) );
  DFF_X1 \u1/fractb_out_reg[6]  ( .D(\u1/fractb_s [6]), .CK(clk), .Q(fractb[6]) );
  DFF_X1 \u1/fractb_out_reg[9]  ( .D(\u1/fractb_s [9]), .CK(clk), .Q(fractb[9]) );
  DFF_X1 \u1/fractb_out_reg[11]  ( .D(\u1/fractb_s [11]), .CK(clk), .Q(
        fractb[11]) );
  DFF_X1 \u1/fracta_out_reg[1]  ( .D(\u1/fracta_s [1]), .CK(clk), .Q(fracta[1]) );
  DFF_X1 \u1/fractb_out_reg[8]  ( .D(\u1/fractb_s [8]), .CK(clk), .Q(fractb[8]) );
  DFF_X1 \u1/fracta_out_reg[6]  ( .D(\u1/fracta_s [6]), .CK(clk), .Q(fracta[6]) );
  DFF_X1 \u1/fractb_out_reg[5]  ( .D(\u1/fractb_s [5]), .CK(clk), .Q(fractb[5]) );
  DFF_X1 \u1/fractb_out_reg[2]  ( .D(\u1/fractb_s [2]), .CK(clk), .Q(fractb[2]) );
  DFF_X1 \u1/fractb_out_reg[1]  ( .D(\u1/fractb_s [1]), .CK(clk), .Q(fractb[1]) );
  DFF_X1 \u1/fractb_out_reg[7]  ( .D(\u1/fractb_s [7]), .CK(clk), .Q(fractb[7]) );
  DFF_X1 \u1/fractb_out_reg[3]  ( .D(\u1/fractb_s [3]), .CK(clk), .Q(fractb[3]) );
  DFF_X1 \u1/sign_reg  ( .D(\u1/sign_d ), .CK(clk), .Q(sign_fasu) );
  DFF_X1 \u1/fracta_out_reg[9]  ( .D(\u1/fracta_s [9]), .CK(clk), .Q(fracta[9]) );
  DFF_X1 \u1/fracta_out_reg[10]  ( .D(\u1/fracta_s [10]), .CK(clk), .Q(
        fracta[10]) );
  DFF_X1 \u1/fracta_out_reg[12]  ( .D(\u1/fracta_s [12]), .CK(clk), .Q(
        fracta[12]) );
  DFF_X1 \u1/fracta_out_reg[8]  ( .D(\u1/fracta_s [8]), .CK(clk), .Q(fracta[8]) );
  DFF_X1 \u1/fractb_out_reg[12]  ( .D(\u1/fractb_s [12]), .CK(clk), .Q(
        fractb[12]) );
  DFF_X1 \u1/fracta_out_reg[11]  ( .D(\u1/fracta_s [11]), .CK(clk), .Q(
        fracta[11]) );
  DFF_X1 \u1/fracta_out_reg[7]  ( .D(\u1/fracta_s [7]), .CK(clk), .Q(fracta[7]) );
  DFF_X1 \fract_out_q_reg[14]  ( .D(n3284), .CK(clk), .Q(fract_out_q[14]) );
  DFF_X1 \u5/prod1_reg[10]  ( .D(\u5/N10 ), .CK(clk), .Q(\u5/prod1 [10]) );
  DFF_X1 \fract_out_q_reg[11]  ( .D(n3287), .CK(clk), .Q(fract_out_q[11]) );
  DFF_X1 \fract_out_q_reg[10]  ( .D(n3288), .CK(clk), .Q(fract_out_q[10]) );
  DFF_X1 \u5/prod1_reg[8]  ( .D(\u5/N8 ), .CK(clk), .Q(\u5/prod1 [8]) );
  DFF_X1 \fract_i2f_reg[2]  ( .D(n3282), .CK(clk), .Q(n1668) );
  DFF_X1 \fract_i2f_reg[15]  ( .D(N190), .CK(clk), .Q(n1667) );
  DFF_X1 \fract_i2f_reg[0]  ( .D(n3318), .CK(clk), .Q(n1660) );
  DFF_X1 \fract_i2f_reg[11]  ( .D(N186), .CK(clk), .Q(n1659) );
  DFF_X1 \fract_i2f_reg[12]  ( .D(N187), .CK(clk), .Q(n1658) );
  DFF_X1 \fract_i2f_reg[6]  ( .D(N181), .CK(clk), .Q(n1657) );
  DFF_X1 \fract_out_q_reg[0]  ( .D(n3298), .CK(clk), .Q(n1656) );
  DFF_X1 \fract_i2f_reg[5]  ( .D(N180), .CK(clk), .Q(n1652) );
  DFF_X1 \fract_i2f_reg[21]  ( .D(N196), .CK(clk), .Q(n1643) );
  DFF_X1 \fract_i2f_reg[17]  ( .D(N192), .CK(clk), .Q(n1634) );
  DFF_X1 \fract_i2f_reg[19]  ( .D(N194), .CK(clk), .Q(n1633) );
  DFF_X1 \out_reg[0]  ( .D(N220), .CK(clk), .Q(out[0]) );
  DFF_X1 \out_reg[11]  ( .D(N231), .CK(clk), .Q(out[11]) );
  DFF_X1 \out_reg[10]  ( .D(N230), .CK(clk), .Q(out[10]) );
  DFF_X1 \u5/prod1_reg[17]  ( .D(\u5/N17 ), .CK(clk), .Q(\u5/prod1 [17]) );
  DFF_X2 \u1/fractb_out_reg[0]  ( .D(\u1/fractb_s [0]), .CK(clk), .Q(fractb[0]) );
  DFF_X1 \fract_out_q_reg[12]  ( .D(n3286), .CK(clk), .Q(fract_out_q[12]) );
  INV_X4 U1188 ( .A(net85292), .ZN(net90110) );
  INV_X4 U1189 ( .A(net85292), .ZN(net85160) );
  INV_X4 U1190 ( .A(net85263), .ZN(net85357) );
  NAND4_X2 U1191 ( .A1(net85260), .A2(n1743), .A3(net85263), .A4(1'b1), .ZN(
        net85187) );
  NAND2_X2 U1192 ( .A1(net85349), .A2(n1839), .ZN(n1838) );
  NAND2_X2 U1193 ( .A1(n3058), .A2(n3057), .ZN(n2177) );
  NAND2_X2 U1194 ( .A1(n1616), .A2(n1584), .ZN(n2173) );
  INV_X4 U1195 ( .A(net83963), .ZN(n2213) );
  INV_X4 U1196 ( .A(exp_r[4]), .ZN(n2115) );
  NAND2_X2 U1197 ( .A1(fract_out_q[13]), .A2(net83780), .ZN(net91059) );
  NAND2_X2 U1198 ( .A1(net83780), .A2(fract_out_q[13]), .ZN(net85247) );
  INV_X4 U1199 ( .A(exp_r[4]), .ZN(n2288) );
  INV_X4 U1200 ( .A(net91112), .ZN(n2200) );
  NAND2_X2 U1201 ( .A1(n2214), .A2(n2213), .ZN(net84722) );
  OAI211_X2 U1202 ( .C1(n2117), .C2(1'b0), .A(n2115), .B(n2114), .ZN(n2634) );
  NOR2_X1 U1203 ( .A1(n2099), .A2(n1527), .ZN(n1524) );
  NOR2_X2 U1204 ( .A1(n1524), .A2(n1525), .ZN(n1552) );
  AND2_X2 U1205 ( .A1(n1526), .A2(n1549), .ZN(n1525) );
  INV_X4 U1206 ( .A(n1825), .ZN(n1526) );
  OR2_X4 U1207 ( .A1(net88293), .A2(n1825), .ZN(n1527) );
  OAI21_X4 U1208 ( .B1(net84778), .B2(n2161), .A(n2160), .ZN(n1528) );
  INV_X8 U1209 ( .A(\u4/fract_out[6] ), .ZN(net84113) );
  INV_X8 U1210 ( .A(net91299), .ZN(net84118) );
  INV_X2 U1211 ( .A(n1752), .ZN(net91298) );
  NOR2_X4 U1212 ( .A1(\u4/fract_out[1] ), .A2(\u4/fract_out[4] ), .ZN(n1798)
         );
  NAND2_X4 U1213 ( .A1(n1873), .A2(net83959), .ZN(n1745) );
  NAND2_X2 U1214 ( .A1(net84069), .A2(net84070), .ZN(net84055) );
  NAND2_X2 U1215 ( .A1(net84071), .A2(net84072), .ZN(net83860) );
  INV_X2 U1216 ( .A(net83860), .ZN(net84070) );
  OAI21_X2 U1217 ( .B1(n2627), .B2(net83860), .A(net83861), .ZN(n2708) );
  INV_X2 U1218 ( .A(n2453), .ZN(n2455) );
  AOI21_X2 U1219 ( .B1(n2695), .B2(n2694), .A(n2615), .ZN(n2616) );
  OAI21_X4 U1220 ( .B1(net84575), .B2(net84574), .A(net84576), .ZN(n1529) );
  OAI21_X2 U1221 ( .B1(net84575), .B2(net84574), .A(net84576), .ZN(net91511)
         );
  OAI211_X2 U1222 ( .C1(net91015), .C2(net85018), .A(net85020), .B(net85021), 
        .ZN(n1530) );
  NOR2_X2 U1223 ( .A1(net84374), .A2(net84373), .ZN(n1536) );
  INV_X1 U1224 ( .A(n2625), .ZN(n1531) );
  INV_X2 U1225 ( .A(net84373), .ZN(n1532) );
  INV_X4 U1226 ( .A(n1532), .ZN(n1533) );
  NOR3_X2 U1227 ( .A1(n2359), .A2(n2360), .A3(n1597), .ZN(net84373) );
  INV_X2 U1228 ( .A(n1749), .ZN(n1534) );
  INV_X2 U1229 ( .A(n1534), .ZN(n1535) );
  NOR2_X4 U1230 ( .A1(net84372), .A2(n1537), .ZN(net86174) );
  INV_X4 U1231 ( .A(n1536), .ZN(n1537) );
  INV_X4 U1232 ( .A(n2926), .ZN(n2924) );
  NAND2_X4 U1233 ( .A1(opa_r[12]), .A2(n2799), .ZN(n2773) );
  INV_X4 U1234 ( .A(n2809), .ZN(n1539) );
  INV_X2 U1235 ( .A(n2817), .ZN(n2806) );
  OAI21_X2 U1236 ( .B1(n2820), .B2(n2818), .A(n2817), .ZN(n2822) );
  AOI211_X4 U1237 ( .C1(n2894), .C2(n2893), .A(n2892), .B(n2891), .ZN(n2903)
         );
  NOR2_X1 U1238 ( .A1(opa_r[14]), .A2(opb_r[14]), .ZN(n2815) );
  NOR2_X2 U1239 ( .A1(\u1/adj_op_out_sft[13] ), .A2(n2791), .ZN(n2928) );
  NOR2_X1 U1240 ( .A1(opa_r[13]), .A2(opa_r[14]), .ZN(n1984) );
  INV_X4 U1241 ( .A(n1733), .ZN(n1541) );
  NAND2_X4 U1242 ( .A1(n1734), .A2(n1730), .ZN(n1729) );
  BUF_X32 U1243 ( .A(n1728), .Z(n1543) );
  AND2_X2 U1244 ( .A1(fracta_mul[0]), .A2(n3045), .ZN(n3022) );
  OAI21_X4 U1245 ( .B1(net84211), .B2(n2339), .A(net91542), .ZN(net84169) );
  NAND2_X4 U1246 ( .A1(n2527), .A2(n2526), .ZN(net84060) );
  INV_X2 U1247 ( .A(net83736), .ZN(net83856) );
  NAND2_X4 U1248 ( .A1(net83871), .A2(n1736), .ZN(N230) );
  NAND2_X4 U1249 ( .A1(n2457), .A2(n2458), .ZN(n2520) );
  NAND2_X2 U1250 ( .A1(n2433), .A2(n2707), .ZN(N234) );
  BUF_X4 U1251 ( .A(net83765), .Z(n1546) );
  INV_X8 U1252 ( .A(net83765), .ZN(net83800) );
  INV_X8 U1253 ( .A(n2460), .ZN(n2528) );
  NAND3_X4 U1254 ( .A1(n1832), .A2(net84253), .A3(net84254), .ZN(net84096) );
  AOI21_X4 U1255 ( .B1(n2705), .B2(n2704), .A(n2703), .ZN(N278) );
  INV_X8 U1256 ( .A(n2618), .ZN(n2656) );
  AND3_X2 U1257 ( .A1(n2656), .A2(n1742), .A3(net83806), .ZN(N290) );
  BUF_X32 U1258 ( .A(n1751), .Z(n1548) );
  INV_X8 U1259 ( .A(net84138), .ZN(net84211) );
  OAI21_X1 U1260 ( .B1(n1548), .B2(net83429), .A(n2963), .ZN(n3010) );
  NAND2_X4 U1261 ( .A1(n1746), .A2(net84472), .ZN(n1597) );
  INV_X2 U1262 ( .A(n1747), .ZN(n1746) );
  OAI211_X1 U1263 ( .C1(n1554), .C2(net84312), .A(net85842), .B(net84133), 
        .ZN(n1842) );
  NAND4_X1 U1264 ( .A1(net91511), .A2(n1749), .A3(net84128), .A4(n1580), .ZN(
        n2359) );
  INV_X16 U1265 ( .A(net85853), .ZN(net86067) );
  NAND2_X4 U1266 ( .A1(net85317), .A2(net86067), .ZN(n1878) );
  INV_X8 U1267 ( .A(n2065), .ZN(n2043) );
  AOI22_X4 U1268 ( .A1(net89998), .A2(n1609), .B1(net85077), .B2(prod[20]), 
        .ZN(net90019) );
  NAND2_X4 U1269 ( .A1(n1896), .A2(net85071), .ZN(net90080) );
  NOR2_X4 U1270 ( .A1(net85752), .A2(net85730), .ZN(n2015) );
  INV_X4 U1271 ( .A(net77637), .ZN(net84910) );
  INV_X8 U1272 ( .A(net84910), .ZN(net90290) );
  INV_X8 U1273 ( .A(net85331), .ZN(net85203) );
  OR2_X4 U1274 ( .A1(net85832), .A2(net86037), .ZN(n1549) );
  AND2_X2 U1275 ( .A1(n2653), .A2(net86038), .ZN(n1550) );
  AND2_X4 U1276 ( .A1(net85107), .A2(net85108), .ZN(n1551) );
  INV_X8 U1277 ( .A(n2139), .ZN(n1940) );
  OAI21_X4 U1278 ( .B1(net84754), .B2(net84755), .A(n1905), .ZN(n1761) );
  INV_X1 U1279 ( .A(net83945), .ZN(net84672) );
  INV_X2 U1280 ( .A(net84672), .ZN(net88500) );
  INV_X16 U1281 ( .A(net91404), .ZN(net84150) );
  INV_X8 U1282 ( .A(net84995), .ZN(net85015) );
  INV_X8 U1283 ( .A(net84994), .ZN(net89753) );
  AND2_X2 U1284 ( .A1(net83959), .A2(n1593), .ZN(n1553) );
  INV_X8 U1285 ( .A(net91298), .ZN(net91299) );
  NAND2_X4 U1286 ( .A1(net84366), .A2(net84453), .ZN(n2437) );
  AND2_X4 U1287 ( .A1(net84474), .A2(net84475), .ZN(n1554) );
  AND2_X2 U1288 ( .A1(n1754), .A2(n2170), .ZN(n1555) );
  NAND2_X4 U1289 ( .A1(net84133), .A2(n2437), .ZN(n2490) );
  INV_X16 U1290 ( .A(net84135), .ZN(net84133) );
  INV_X1 U1291 ( .A(net83875), .ZN(net84085) );
  NAND2_X4 U1292 ( .A1(net84136), .A2(rmode_r3[1]), .ZN(n2496) );
  AOI21_X4 U1293 ( .B1(net86174), .B2(net84075), .A(net84206), .ZN(net84204)
         );
  NAND2_X1 U1294 ( .A1(net89856), .A2(net85041), .ZN(net10316) );
  INV_X16 U1295 ( .A(net85097), .ZN(net85089) );
  NAND2_X4 U1296 ( .A1(net84757), .A2(net84758), .ZN(net91555) );
  NAND2_X2 U1297 ( .A1(net84757), .A2(net84758), .ZN(net84301) );
  NAND3_X2 U1298 ( .A1(net85730), .A2(net85716), .A3(fract_out_q[4]), .ZN(
        n2068) );
  NOR2_X4 U1299 ( .A1(net11576), .A2(net85718), .ZN(n1556) );
  NAND3_X2 U1300 ( .A1(n2070), .A2(n2068), .A3(n2069), .ZN(net85197) );
  INV_X4 U1301 ( .A(n2070), .ZN(n2071) );
  NAND2_X2 U1302 ( .A1(net85144), .A2(n2053), .ZN(n1954) );
  OAI21_X1 U1303 ( .B1(n2055), .B2(net89677), .A(net85105), .ZN(n2057) );
  INV_X8 U1304 ( .A(n1912), .ZN(n1909) );
  AND2_X4 U1305 ( .A1(net86090), .A2(n1893), .ZN(n1891) );
  INV_X16 U1306 ( .A(net85010), .ZN(net83959) );
  BUF_X16 U1307 ( .A(net85095), .Z(net89078) );
  NOR2_X4 U1308 ( .A1(\u4/N656 ), .A2(n1571), .ZN(net85010) );
  BUF_X16 U1309 ( .A(net84609), .Z(net90122) );
  INV_X8 U1310 ( .A(n1792), .ZN(net89657) );
  NOR2_X4 U1311 ( .A1(\u4/exp_out[2] ), .A2(\u4/N653 ), .ZN(n1787) );
  INV_X2 U1312 ( .A(net86112), .ZN(net85038) );
  NAND2_X2 U1313 ( .A1(n1652), .A2(net85720), .ZN(net86096) );
  NOR2_X4 U1314 ( .A1(net76619), .A2(net85204), .ZN(n2047) );
  NAND2_X2 U1315 ( .A1(net85043), .A2(net85042), .ZN(net76619) );
  XNOR2_X1 U1316 ( .A(net84668), .B(net84610), .ZN(net84667) );
  INV_X4 U1317 ( .A(net85082), .ZN(net88618) );
  INV_X8 U1318 ( .A(net84299), .ZN(net88877) );
  NAND2_X4 U1319 ( .A1(net88895), .A2(n1777), .ZN(n1776) );
  NAND2_X2 U1320 ( .A1(n1794), .A2(net89658), .ZN(net83395) );
  NAND2_X2 U1321 ( .A1(net88646), .A2(n1792), .ZN(net89658) );
  NAND2_X2 U1322 ( .A1(n1951), .A2(n1950), .ZN(n1557) );
  INV_X8 U1323 ( .A(n2383), .ZN(n2385) );
  INV_X8 U1324 ( .A(net85720), .ZN(net88319) );
  INV_X2 U1325 ( .A(\u4/N424 ), .ZN(net84830) );
  NAND2_X4 U1326 ( .A1(\u4/N424 ), .A2(net84522), .ZN(n1869) );
  OAI21_X2 U1327 ( .B1(net84761), .B2(net85712), .A(net84610), .ZN(n1781) );
  NAND3_X1 U1328 ( .A1(net85712), .A2(n2099), .A3(net86038), .ZN(n2090) );
  NOR2_X1 U1329 ( .A1(rmode_r3[0]), .A2(net85847), .ZN(n2279) );
  AOI21_X2 U1330 ( .B1(n2221), .B2(n2261), .A(n2220), .ZN(n2224) );
  AOI21_X2 U1331 ( .B1(net83941), .B2(n1813), .A(n1814), .ZN(n1812) );
  NOR2_X2 U1332 ( .A1(net84206), .A2(net83864), .ZN(n1833) );
  NOR2_X1 U1333 ( .A1(n1720), .A2(n2948), .ZN(n2851) );
  OAI21_X1 U1334 ( .B1(net83849), .B2(n1596), .A(net83439), .ZN(n1906) );
  NAND3_X2 U1335 ( .A1(net84524), .A2(net84518), .A3(net84519), .ZN(net84458)
         );
  NAND3_X2 U1336 ( .A1(n2300), .A2(n2299), .A3(n2298), .ZN(net84524) );
  NOR2_X1 U1337 ( .A1(net85794), .A2(net83439), .ZN(n2299) );
  NOR2_X2 U1338 ( .A1(n2084), .A2(n2083), .ZN(n2085) );
  NAND2_X1 U1339 ( .A1(net89372), .A2(net85832), .ZN(net84160) );
  NOR2_X1 U1340 ( .A1(n2415), .A2(net83878), .ZN(n2325) );
  NOR2_X1 U1341 ( .A1(net11560), .A2(net84167), .ZN(n2562) );
  NAND3_X2 U1342 ( .A1(net84518), .A2(net85790), .A3(net84519), .ZN(net83946)
         );
  AOI21_X2 U1343 ( .B1(n2127), .B2(net85790), .A(n2126), .ZN(n2129) );
  NOR2_X1 U1344 ( .A1(n2306), .A2(n2991), .ZN(n2126) );
  NAND2_X2 U1345 ( .A1(n1842), .A2(net84385), .ZN(n1845) );
  INV_X4 U1346 ( .A(net86015), .ZN(net84394) );
  NAND3_X2 U1347 ( .A1(n2857), .A2(n2856), .A3(n2855), .ZN(n2864) );
  NOR2_X2 U1348 ( .A1(n2904), .A2(n2937), .ZN(n2908) );
  INV_X4 U1349 ( .A(n2190), .ZN(n2054) );
  NOR2_X1 U1350 ( .A1(net11671), .A2(net83993), .ZN(n2207) );
  NAND2_X2 U1351 ( .A1(n2498), .A2(net84128), .ZN(n2499) );
  NOR3_X1 U1352 ( .A1(n2472), .A2(n2471), .A3(n2470), .ZN(n2473) );
  NAND3_X1 U1353 ( .A1(net84343), .A2(net85790), .A3(n2317), .ZN(n2318) );
  AOI21_X1 U1354 ( .B1(n2316), .B2(net85790), .A(n2315), .ZN(n2319) );
  NAND2_X2 U1355 ( .A1(n2372), .A2(n2374), .ZN(n1932) );
  NOR2_X2 U1356 ( .A1(net83791), .A2(n1576), .ZN(net83747) );
  INV_X4 U1357 ( .A(net11567), .ZN(net85827) );
  NAND3_X2 U1358 ( .A1(n1984), .A2(n1573), .A3(n1983), .ZN(n3313) );
  INV_X4 U1359 ( .A(n1911), .ZN(n1910) );
  NOR2_X1 U1360 ( .A1(\u4/exp_in_pl1[3] ), .A2(n2551), .ZN(n2195) );
  NOR2_X2 U1361 ( .A1(n2943), .A2(n2890), .ZN(n2891) );
  NOR2_X1 U1362 ( .A1(net83995), .A2(net83974), .ZN(net83971) );
  AOI21_X1 U1363 ( .B1(n2562), .B2(net85832), .A(net83968), .ZN(n2563) );
  NAND3_X1 U1364 ( .A1(n2141), .A2(n872), .A3(n2140), .ZN(n2142) );
  NOR2_X2 U1365 ( .A1(n2263), .A2(n2243), .ZN(n2150) );
  NOR2_X2 U1366 ( .A1(n2573), .A2(n2546), .ZN(n2547) );
  NAND3_X2 U1367 ( .A1(n2181), .A2(n2180), .A3(n2179), .ZN(n2548) );
  NOR2_X2 U1368 ( .A1(n2172), .A2(n2171), .ZN(n2181) );
  NOR2_X2 U1369 ( .A1(n2174), .A2(n2173), .ZN(n2180) );
  NOR2_X2 U1370 ( .A1(n2469), .A2(n2486), .ZN(n2470) );
  AOI21_X1 U1371 ( .B1(n2305), .B2(net83927), .A(net83969), .ZN(n2312) );
  NAND3_X1 U1372 ( .A1(net83813), .A2(net84501), .A3(net84498), .ZN(net84500)
         );
  NOR2_X2 U1373 ( .A1(net86169), .A2(net84220), .ZN(n2321) );
  AOI211_X2 U1374 ( .C1(\u4/exp_next_mi[3] ), .C2(net84157), .A(net84220), .B(
        net83878), .ZN(n1877) );
  OAI21_X2 U1375 ( .B1(n2121), .B2(n2132), .A(n2120), .ZN(n2281) );
  NOR2_X1 U1376 ( .A1(prod[20]), .A2(n2650), .ZN(n2652) );
  NAND3_X1 U1377 ( .A1(net83940), .A2(net83941), .A3(net83936), .ZN(n2601) );
  NOR2_X1 U1378 ( .A1(n2573), .A2(net83950), .ZN(n2574) );
  NOR2_X2 U1379 ( .A1(n1613), .A2(n1575), .ZN(n2353) );
  OAI21_X1 U1380 ( .B1(n2876), .B2(n2863), .A(n2862), .ZN(n2865) );
  NOR2_X2 U1381 ( .A1(n2928), .A2(n2929), .ZN(n2917) );
  NOR2_X2 U1382 ( .A1(n1927), .A2(n3319), .ZN(net84912) );
  OAI21_X2 U1383 ( .B1(n2105), .B2(n2104), .A(n2103), .ZN(n2106) );
  NAND2_X1 U1384 ( .A1(net84672), .A2(net84673), .ZN(net84602) );
  OAI21_X1 U1385 ( .B1(net83427), .B2(net84600), .A(net83408), .ZN(net84598)
         );
  NOR2_X1 U1386 ( .A1(net83438), .A2(net83427), .ZN(net84599) );
  NOR2_X2 U1387 ( .A1(n1822), .A2(n1823), .ZN(n1824) );
  NOR2_X2 U1388 ( .A1(n1859), .A2(n1617), .ZN(n1858) );
  NOR3_X2 U1389 ( .A1(net84043), .A2(n1561), .A3(net84033), .ZN(n1861) );
  NAND3_X2 U1390 ( .A1(opa_inf), .A2(opb_inf), .A3(sign_exe_r), .ZN(net84047)
         );
  AOI21_X2 U1391 ( .B1(net85778), .B2(net84326), .A(n2303), .ZN(n2158) );
  NAND4_X2 U1392 ( .A1(n2523), .A2(n2527), .A3(n2526), .A4(n2524), .ZN(n2502)
         );
  NOR2_X2 U1393 ( .A1(opa_inf), .A2(opb_00), .ZN(n2376) );
  NOR2_X1 U1394 ( .A1(net84076), .A2(n2531), .ZN(net84073) );
  NOR2_X2 U1395 ( .A1(n3143), .A2(n2767), .ZN(n2730) );
  NOR2_X1 U1396 ( .A1(net83849), .A2(net83933), .ZN(n2114) );
  OAI21_X1 U1397 ( .B1(div_opa_ldz_r2[3]), .B2(net83968), .A(n2292), .ZN(n2285) );
  OAI21_X1 U1398 ( .B1(net83968), .B2(n2225), .A(exp_r[4]), .ZN(n2227) );
  AOI211_X2 U1399 ( .C1(n2258), .C2(n2257), .A(n2256), .B(net83423), .ZN(n2267) );
  AOI21_X1 U1400 ( .B1(n2255), .B2(net84639), .A(net83408), .ZN(n2256) );
  OAI21_X1 U1401 ( .B1(net11555), .B2(net83849), .A(net85828), .ZN(n2597) );
  OAI21_X2 U1402 ( .B1(n2700), .B2(net86010), .A(n2699), .ZN(n2701) );
  NOR2_X2 U1403 ( .A1(n1574), .A2(n1629), .ZN(n2700) );
  INV_X16 U1404 ( .A(net85846), .ZN(net85847) );
  NAND3_X2 U1405 ( .A1(n2538), .A2(n2537), .A3(n2536), .ZN(n2540) );
  NAND3_X2 U1406 ( .A1(n1575), .A2(net84021), .A3(n2535), .ZN(n2537) );
  NOR2_X2 U1407 ( .A1(n3143), .A2(n2833), .ZN(n2759) );
  NOR2_X2 U1408 ( .A1(net84249), .A2(net83791), .ZN(n2430) );
  NOR2_X2 U1409 ( .A1(n2889), .A2(n2896), .ZN(n1993) );
  INV_X8 U1410 ( .A(net85832), .ZN(net85778) );
  NOR3_X2 U1411 ( .A1(net84643), .A2(net84445), .A3(n1852), .ZN(net84645) );
  NAND2_X2 U1412 ( .A1(net84654), .A2(n1788), .ZN(net90079) );
  NOR2_X1 U1413 ( .A1(net83993), .A2(net83994), .ZN(n2560) );
  AOI21_X2 U1414 ( .B1(n2297), .B2(n2296), .A(n2295), .ZN(n2298) );
  INV_X4 U1415 ( .A(net86006), .ZN(net85732) );
  INV_X4 U1416 ( .A(net85071), .ZN(net85211) );
  NOR2_X2 U1417 ( .A1(n1642), .A2(opb_dn), .ZN(n1760) );
  NOR2_X2 U1418 ( .A1(net85847), .A2(n2077), .ZN(n2079) );
  OAI21_X2 U1419 ( .B1(n2260), .B2(n2195), .A(n2194), .ZN(n2202) );
  OAI21_X2 U1420 ( .B1(n2241), .B2(n2240), .A(n2239), .ZN(n2245) );
  NOR2_X2 U1421 ( .A1(n2238), .A2(n2263), .ZN(n2240) );
  NOR3_X1 U1422 ( .A1(n2019), .A2(net84290), .A3(net84305), .ZN(
        \u4/exp_in_pl1[5] ) );
  NAND3_X2 U1423 ( .A1(n1620), .A2(n1587), .A3(n1568), .ZN(n2174) );
  NAND3_X2 U1424 ( .A1(n1619), .A2(n1586), .A3(n1567), .ZN(n2171) );
  NAND3_X2 U1425 ( .A1(n1618), .A2(n1585), .A3(n1566), .ZN(n2172) );
  NAND3_X1 U1426 ( .A1(net83942), .A2(n1817), .A3(net84858), .ZN(n1813) );
  NOR2_X2 U1427 ( .A1(n2836), .A2(n2835), .ZN(n2838) );
  NOR2_X1 U1428 ( .A1(net11670), .A2(net85832), .ZN(n2208) );
  NOR2_X2 U1429 ( .A1(net85137), .A2(net77161), .ZN(net85136) );
  INV_X8 U1430 ( .A(net85196), .ZN(n1865) );
  INV_X4 U1431 ( .A(net85360), .ZN(net85159) );
  NOR2_X2 U1432 ( .A1(net83969), .A2(n2561), .ZN(n2569) );
  AOI21_X2 U1433 ( .B1(net84133), .B2(net84134), .A(net84128), .ZN(n2495) );
  NOR2_X1 U1434 ( .A1(net11560), .A2(n2461), .ZN(n2463) );
  NOR2_X1 U1435 ( .A1(n2466), .A2(n2482), .ZN(n2471) );
  OAI21_X2 U1436 ( .B1(net84884), .B2(n1571), .A(n2145), .ZN(net84853) );
  OAI21_X1 U1437 ( .B1(n2580), .B2(net84675), .A(net85794), .ZN(n2145) );
  NOR2_X1 U1438 ( .A1(net84886), .A2(n1596), .ZN(net84884) );
  AOI21_X1 U1439 ( .B1(n2314), .B2(n2313), .A(net84468), .ZN(n2315) );
  OAI21_X1 U1440 ( .B1(net83933), .B2(net83963), .A(net84465), .ZN(n2313) );
  NAND2_X2 U1441 ( .A1(n2339), .A2(net84421), .ZN(n2498) );
  NOR2_X2 U1442 ( .A1(n2409), .A2(n2408), .ZN(n2410) );
  AOI21_X2 U1443 ( .B1(n2403), .B2(n2444), .A(n2402), .ZN(n2412) );
  NOR2_X1 U1444 ( .A1(\u4/exp_in_pl1[3] ), .A2(n2401), .ZN(n2402) );
  NOR2_X1 U1445 ( .A1(net11555), .A2(n1571), .ZN(net84278) );
  NAND3_X1 U1446 ( .A1(n2304), .A2(net85832), .A3(net83963), .ZN(net83927) );
  NOR2_X1 U1447 ( .A1(opa_dn), .A2(net88427), .ZN(net84506) );
  NAND3_X2 U1448 ( .A1(n2859), .A2(n2862), .A3(n2858), .ZN(n2866) );
  NOR2_X2 U1449 ( .A1(opb_r[11]), .A2(n1725), .ZN(n2771) );
  NOR2_X2 U1450 ( .A1(n2204), .A2(n2203), .ZN(n2212) );
  NOR2_X1 U1451 ( .A1(n3096), .A2(net83994), .ZN(n2203) );
  NOR2_X1 U1452 ( .A1(n1663), .A2(net83968), .ZN(n2204) );
  NOR2_X1 U1453 ( .A1(net11558), .A2(n2209), .ZN(n2210) );
  NAND3_X2 U1454 ( .A1(n2184), .A2(n2183), .A3(n2182), .ZN(n2301) );
  NAND3_X2 U1455 ( .A1(net83934), .A2(n1853), .A3(net83936), .ZN(net83836) );
  NOR2_X2 U1456 ( .A1(n2425), .A2(n2387), .ZN(n2389) );
  NOR3_X2 U1457 ( .A1(n2458), .A2(n2343), .A3(n2342), .ZN(n2344) );
  AOI21_X2 U1458 ( .B1(n1583), .B2(n2418), .A(net85794), .ZN(net84265) );
  OAI21_X2 U1459 ( .B1(net84465), .B2(n2324), .A(n2323), .ZN(net84080) );
  NOR2_X1 U1460 ( .A1(net84468), .A2(net84343), .ZN(n2323) );
  NOR3_X2 U1461 ( .A1(net84469), .A2(net83927), .A3(n2322), .ZN(n2324) );
  AOI21_X2 U1462 ( .B1(n2362), .B2(net84368), .A(n1768), .ZN(n2371) );
  OAI21_X2 U1463 ( .B1(n1628), .B2(n2368), .A(n2367), .ZN(n2369) );
  NAND3_X1 U1464 ( .A1(net85828), .A2(net85790), .A3(n1571), .ZN(n1835) );
  OAI21_X2 U1465 ( .B1(n2100), .B2(n2076), .A(n2102), .ZN(n2108) );
  INV_X4 U1466 ( .A(net89411), .ZN(net89412) );
  INV_X4 U1467 ( .A(net89446), .ZN(net89447) );
  NOR2_X1 U1468 ( .A1(net83968), .A2(n1663), .ZN(n2113) );
  OAI21_X2 U1469 ( .B1(n2284), .B2(n2283), .A(n2282), .ZN(n2292) );
  NOR2_X1 U1470 ( .A1(div_opa_ldz_r2[2]), .A2(exp_r[2]), .ZN(n2283) );
  NOR2_X1 U1471 ( .A1(n2266), .A2(net83427), .ZN(net84617) );
  NOR2_X1 U1472 ( .A1(net84445), .A2(net83402), .ZN(n2258) );
  NOR2_X1 U1473 ( .A1(net84632), .A2(net83403), .ZN(n2257) );
  AOI211_X1 U1474 ( .C1(net84823), .C2(net11566), .A(net84571), .B(net85790), 
        .ZN(n2169) );
  NOR2_X1 U1475 ( .A1(net11555), .A2(net84279), .ZN(net84823) );
  NOR2_X1 U1476 ( .A1(n2307), .A2(net88427), .ZN(net84664) );
  NAND2_X2 U1477 ( .A1(\u1/adj_op_out_sft[1] ), .A2(n2791), .ZN(n2923) );
  NOR2_X2 U1478 ( .A1(n1561), .A2(n1581), .ZN(net84064) );
  NOR2_X2 U1479 ( .A1(net83791), .A2(n1631), .ZN(n2653) );
  NOR3_X1 U1480 ( .A1(prod[17]), .A2(prod[18]), .A3(prod[19]), .ZN(n2651) );
  OAI21_X2 U1481 ( .B1(n2591), .B2(n2590), .A(n2619), .ZN(n2592) );
  NOR2_X2 U1482 ( .A1(n2589), .A2(n2588), .ZN(n2590) );
  NOR3_X2 U1483 ( .A1(n1605), .A2(n2603), .A3(n2602), .ZN(n2607) );
  NOR2_X2 U1484 ( .A1(opa_inf), .A2(net83791), .ZN(n2535) );
  NOR2_X2 U1485 ( .A1(net83791), .A2(n2698), .ZN(n2534) );
  NOR2_X2 U1486 ( .A1(net84326), .A2(net84327), .ZN(n2384) );
  NAND3_X1 U1487 ( .A1(net84465), .A2(net84343), .A3(net85790), .ZN(n2320) );
  INV_X4 U1488 ( .A(n2770), .ZN(n2784) );
  INV_X2 U1489 ( .A(\u1/adj_op_out_sft[4] ), .ZN(n1721) );
  NOR2_X1 U1490 ( .A1(net85794), .A2(n1570), .ZN(n2428) );
  INV_X4 U1491 ( .A(net83419), .ZN(n1783) );
  OAI21_X1 U1492 ( .B1(n2973), .B2(n2972), .A(n2971), .ZN(n2974) );
  AOI21_X1 U1493 ( .B1(n2270), .B2(net84604), .A(net83403), .ZN(n2274) );
  NOR2_X1 U1494 ( .A1(n1852), .A2(net84579), .ZN(n1851) );
  NOR2_X2 U1495 ( .A1(net84913), .A2(n1608), .ZN(net84906) );
  NOR2_X2 U1496 ( .A1(result_zero_sign_d), .A2(n1803), .ZN(n1807) );
  AOI21_X2 U1497 ( .B1(n1561), .B2(n1860), .A(n1861), .ZN(n1855) );
  NOR2_X1 U1498 ( .A1(net84048), .A2(n1863), .ZN(net84028) );
  OAI21_X1 U1499 ( .B1(net85794), .B2(n2376), .A(net83779), .ZN(n2377) );
  INV_X4 U1500 ( .A(n2666), .ZN(n2670) );
  OAI21_X2 U1501 ( .B1(net83791), .B2(n2662), .A(n2661), .ZN(n2669) );
  OAI21_X2 U1502 ( .B1(n2660), .B2(n2659), .A(n1561), .ZN(n2661) );
  NOR2_X2 U1503 ( .A1(opb_inf), .A2(n1572), .ZN(n2660) );
  NOR2_X2 U1504 ( .A1(opa_00), .A2(n1570), .ZN(n2659) );
  NAND2_X2 U1505 ( .A1(n3192), .A2(n3174), .ZN(n3159) );
  NAND2_X2 U1506 ( .A1(n3188), .A2(n3165), .ZN(n3180) );
  NAND2_X2 U1507 ( .A1(n3174), .A2(n3165), .ZN(n3181) );
  NAND2_X2 U1508 ( .A1(n1653), .A2(n3182), .ZN(n3175) );
  NOR3_X2 U1509 ( .A1(n1990), .A2(n2895), .A3(n1989), .ZN(n2959) );
  NOR2_X1 U1510 ( .A1(n1725), .A2(n1723), .ZN(n1987) );
  NOR2_X1 U1511 ( .A1(n1541), .A2(n3017), .ZN(n1986) );
  NOR2_X1 U1512 ( .A1(net83402), .A2(net83403), .ZN(net83394) );
  INV_X8 U1513 ( .A(\u4/f2i_shft[1] ), .ZN(net85712) );
  OAI21_X2 U1514 ( .B1(n2986), .B2(n2976), .A(n2975), .ZN(n2977) );
  NOR2_X1 U1515 ( .A1(\u4/sub_409/net10540 ), .A2(div_opa_ldz_r2[3]), .ZN(
        n2976) );
  NOR2_X1 U1516 ( .A1(net84445), .A2(net84643), .ZN(n2268) );
  OAI211_X2 U1517 ( .C1(net83754), .C2(net83819), .A(net83820), .B(n1546), 
        .ZN(net83802) );
  NOR2_X1 U1518 ( .A1(net85847), .A2(net83791), .ZN(n2539) );
  NOR2_X2 U1519 ( .A1(n2737), .A2(n2736), .ZN(n2741) );
  NOR2_X2 U1520 ( .A1(n2744), .A2(n2743), .ZN(n2747) );
  NOR2_X2 U1521 ( .A1(n2749), .A2(n2748), .ZN(n2752) );
  NOR2_X2 U1522 ( .A1(n2756), .A2(n2755), .ZN(n2762) );
  NOR2_X2 U1523 ( .A1(n3121), .A2(n2765), .ZN(\u2/underflow_d [2]) );
  NOR2_X2 U1524 ( .A1(n2957), .A2(net86010), .ZN(N283) );
  NOR2_X2 U1525 ( .A1(n3156), .A2(fracta_mul[9]), .ZN(\u0/N4 ) );
  NOR2_X2 U1526 ( .A1(n2959), .A2(n2958), .ZN(\u0/N5 ) );
  INV_X1 U1527 ( .A(n3313), .ZN(n3012) );
  OAI21_X2 U1528 ( .B1(n1999), .B2(fracta_mul[8]), .A(n3120), .ZN(N65) );
  AOI21_X2 U1529 ( .B1(n3117), .B2(n1998), .A(fracta_mul[7]), .ZN(n1999) );
  OAI21_X2 U1530 ( .B1(n1997), .B2(n2896), .A(n3116), .ZN(n1998) );
  AOI21_X1 U1531 ( .B1(n3113), .B2(fracta_mul[1]), .A(n2889), .ZN(n1997) );
  OAI21_X2 U1532 ( .B1(n1995), .B2(n1994), .A(n3120), .ZN(n1996) );
  AOI21_X2 U1533 ( .B1(n1993), .B2(n1992), .A(n1991), .ZN(n1995) );
  NOR2_X2 U1534 ( .A1(n2961), .A2(n2960), .ZN(n888) );
  NOR2_X1 U1535 ( .A1(net83438), .A2(n2989), .ZN(n2961) );
  NOR2_X1 U1536 ( .A1(n2962), .A2(net83432), .ZN(n2963) );
  OAI21_X1 U1537 ( .B1(n872), .B2(n2996), .A(n2995), .ZN(\u4/shift_right [3])
         );
  AOI21_X1 U1538 ( .B1(n2994), .B2(net85790), .A(n2993), .ZN(n2995) );
  NOR2_X1 U1539 ( .A1(n2992), .A2(n2991), .ZN(n2993) );
  OAI21_X1 U1540 ( .B1(n872), .B2(net84393), .A(net83368), .ZN(
        \u4/shift_right [4]) );
  AOI21_X1 U1541 ( .B1(n2984), .B2(net85790), .A(n2983), .ZN(net83368) );
  NOR2_X1 U1542 ( .A1(n2982), .A2(n2991), .ZN(n2983) );
  INV_X4 U1543 ( .A(net84030), .ZN(net84027) );
  NAND2_X1 U1544 ( .A1(n2695), .A2(n2676), .ZN(n2677) );
  NAND2_X1 U1545 ( .A1(n2695), .A2(n2682), .ZN(n2684) );
  NAND2_X2 U1546 ( .A1(n1944), .A2(n2695), .ZN(n2668) );
  AND2_X2 U1547 ( .A1(n1749), .A2(net84128), .ZN(n1603) );
  INV_X8 U1548 ( .A(n1748), .ZN(n1749) );
  INV_X4 U1549 ( .A(n2520), .ZN(n2522) );
  NOR3_X2 U1550 ( .A1(n1809), .A2(n1810), .A3(n1811), .ZN(net84051) );
  OAI21_X4 U1551 ( .B1(n2529), .B2(net84083), .A(n1685), .ZN(net84050) );
  NAND2_X1 U1552 ( .A1(n2433), .A2(n1531), .ZN(N232) );
  NAND2_X4 U1553 ( .A1(n1751), .A2(net84409), .ZN(n1748) );
  INV_X4 U1554 ( .A(net84401), .ZN(n1751) );
  NAND2_X4 U1555 ( .A1(net91375), .A2(n1552), .ZN(net84950) );
  NAND2_X2 U1556 ( .A1(net84468), .A2(net84588), .ZN(net84584) );
  OAI22_X2 U1557 ( .A1(n2513), .A2(n2510), .B1(net89485), .B2(n1961), .ZN(
        n2678) );
  AOI21_X2 U1558 ( .B1(net84071), .B2(net84072), .A(net84206), .ZN(n1834) );
  NOR3_X2 U1559 ( .A1(n2595), .A2(n2594), .A3(n2593), .ZN(n2610) );
  INV_X8 U1560 ( .A(net83853), .ZN(net83906) );
  INV_X1 U1561 ( .A(net89657), .ZN(net89919) );
  OAI21_X1 U1562 ( .B1(n2702), .B2(net85794), .A(n2701), .ZN(n2703) );
  NAND3_X2 U1563 ( .A1(n2657), .A2(net83802), .A3(n2658), .ZN(N281) );
  NAND3_X2 U1564 ( .A1(n2656), .A2(net83806), .A3(n2655), .ZN(n2657) );
  AOI21_X2 U1565 ( .B1(n2647), .B2(n2646), .A(n2645), .ZN(n2658) );
  NAND2_X2 U1566 ( .A1(net83395), .A2(net83394), .ZN(net83393) );
  INV_X4 U1567 ( .A(net89054), .ZN(net89055) );
  INV_X4 U1568 ( .A(net84554), .ZN(net84575) );
  BUF_X8 U1569 ( .A(n1535), .Z(net91542) );
  NAND2_X2 U1570 ( .A1(net84329), .A2(net86171), .ZN(net84136) );
  NAND2_X2 U1571 ( .A1(net84329), .A2(rmode_r3[1]), .ZN(n2383) );
  OAI21_X2 U1572 ( .B1(sign), .B2(net84401), .A(net84403), .ZN(net84329) );
  NOR3_X4 U1573 ( .A1(n2709), .A2(n2626), .A3(n2625), .ZN(n2647) );
  NAND2_X4 U1574 ( .A1(net84026), .A2(net84025), .ZN(N254) );
  NAND2_X2 U1575 ( .A1(net84483), .A2(n1654), .ZN(net84554) );
  NAND4_X4 U1576 ( .A1(net90035), .A2(net84912), .A3(net84911), .A4(net84910), 
        .ZN(net84561) );
  INV_X4 U1577 ( .A(net85114), .ZN(net85113) );
  NAND4_X2 U1578 ( .A1(net89943), .A2(n1910), .A3(net85131), .A4(net85180), 
        .ZN(net85114) );
  AND4_X4 U1579 ( .A1(n1636), .A2(n1635), .A3(n1637), .A4(n3193), .ZN(n1558)
         );
  XNOR2_X2 U1580 ( .A(n1676), .B(n1680), .ZN(n1559) );
  INV_X1 U1581 ( .A(n2924), .ZN(n1977) );
  INV_X16 U1582 ( .A(n2926), .ZN(n1975) );
  AND2_X2 U1583 ( .A1(net83779), .A2(net85790), .ZN(n1561) );
  XNOR2_X2 U1584 ( .A(n1625), .B(\sub_435_3/carry [14]), .ZN(n1562) );
  AND2_X2 U1585 ( .A1(\u1/adj_op_out_sft[2] ), .A2(n2791), .ZN(n1563) );
  XNOR2_X2 U1586 ( .A(n1674), .B(\sub_435_b0/carry [3]), .ZN(n1564) );
  XNOR2_X2 U1587 ( .A(n1675), .B(\sub_435_b0/carry [2]), .ZN(n1565) );
  AND2_X4 U1588 ( .A1(net83747), .A2(n1570), .ZN(n1574) );
  AND2_X2 U1589 ( .A1(opb_inf), .A2(net85790), .ZN(n1575) );
  XNOR2_X2 U1590 ( .A(n1624), .B(\sub_435_3/carry [15]), .ZN(n1577) );
  XNOR2_X2 U1591 ( .A(n1637), .B(\sub_435_3/carry [18]), .ZN(n1578) );
  XOR2_X1 U1592 ( .A(div_opa_ldz_r2[3]), .B(net83968), .Z(n1579) );
  AND2_X4 U1593 ( .A1(net84475), .A2(net84150), .ZN(n1580) );
  OR2_X4 U1594 ( .A1(net83791), .A2(n1611), .ZN(n1581) );
  INV_X4 U1595 ( .A(net84079), .ZN(net84157) );
  OR2_X4 U1596 ( .A1(n1731), .A2(n3316), .ZN(n1582) );
  AND2_X2 U1597 ( .A1(n2417), .A2(n2416), .ZN(n1583) );
  AND2_X2 U1598 ( .A1(net84081), .A2(net91404), .ZN(n1588) );
  AND2_X2 U1599 ( .A1(n2187), .A2(net88500), .ZN(n1589) );
  AND2_X2 U1600 ( .A1(\u1/adj_op_out_sft[2] ), .A2(n2793), .ZN(n1590) );
  INV_X2 U1601 ( .A(net85832), .ZN(net15448) );
  INV_X4 U1602 ( .A(net85831), .ZN(net85832) );
  NAND2_X2 U1603 ( .A1(net89863), .A2(net85126), .ZN(n2276) );
  INV_X2 U1604 ( .A(n1977), .ZN(n1976) );
  INV_X8 U1605 ( .A(net91375), .ZN(net89842) );
  XNOR2_X2 U1606 ( .A(n2133), .B(n2100), .ZN(n1592) );
  INV_X4 U1607 ( .A(opb_r[12]), .ZN(n2799) );
  AND2_X2 U1608 ( .A1(n2226), .A2(net84236), .ZN(n1593) );
  INV_X2 U1609 ( .A(\u4/N404 ), .ZN(n1800) );
  XNOR2_X2 U1610 ( .A(n1672), .B(\sub_435_3/carry [17]), .ZN(n1598) );
  XNOR2_X2 U1611 ( .A(n1673), .B(\sub_435_3/carry [16]), .ZN(n1599) );
  XNOR2_X2 U1612 ( .A(n1626), .B(\sub_435_3/carry [13]), .ZN(n1600) );
  XNOR2_X2 U1613 ( .A(n1627), .B(\sub_435_3/carry [12]), .ZN(n1601) );
  XNOR2_X2 U1614 ( .A(n1678), .B(\sub_435_3/carry [11]), .ZN(n1602) );
  AND2_X4 U1615 ( .A1(n2575), .A2(net88500), .ZN(n1605) );
  AND3_X4 U1616 ( .A1(net83941), .A2(net83942), .A3(net84488), .ZN(n1606) );
  AND2_X4 U1617 ( .A1(net84265), .A2(net84266), .ZN(n1607) );
  NAND2_X1 U1618 ( .A1(n1821), .A2(net84015), .ZN(net84651) );
  INV_X4 U1619 ( .A(net84651), .ZN(net84649) );
  CLKBUF_X2 U1620 ( .A(n1761), .Z(net89537) );
  AND2_X2 U1621 ( .A1(n2545), .A2(net83946), .ZN(n1610) );
  AND2_X2 U1622 ( .A1(net86038), .A2(opb_00), .ZN(n1613) );
  INV_X4 U1623 ( .A(n2276), .ZN(n1930) );
  INV_X4 U1624 ( .A(net85140), .ZN(net88566) );
  INV_X2 U1625 ( .A(n2938), .ZN(n2904) );
  OR2_X2 U1626 ( .A1(net84984), .A2(net83933), .ZN(n1621) );
  XNOR2_X2 U1627 ( .A(n1689), .B(n3021), .ZN(n1622) );
  NAND2_X2 U1628 ( .A1(n1757), .A2(net89615), .ZN(n1623) );
  AND2_X2 U1629 ( .A1(n2482), .A2(n2486), .ZN(n1628) );
  AND2_X4 U1630 ( .A1(net83747), .A2(net90287), .ZN(n1629) );
  XOR2_X2 U1631 ( .A(\u2/exp_tmp4[3] ), .B(n3020), .Z(n1630) );
  AND2_X2 U1632 ( .A1(n2425), .A2(net85790), .ZN(n1632) );
  AND2_X2 U1633 ( .A1(net84482), .A2(net84551), .ZN(n1638) );
  OR2_X2 U1634 ( .A1(n2488), .A2(n2489), .ZN(n1639) );
  AND2_X2 U1635 ( .A1(net84673), .A2(net85794), .ZN(n1640) );
  INV_X4 U1636 ( .A(n3124), .ZN(n3136) );
  NAND3_X2 U1637 ( .A1(fpu_op_r1[0]), .A2(fpu_op_r1[1]), .A3(n3100), .ZN(n3124) );
  AND2_X2 U1638 ( .A1(\u1/adj_op_out_sft[1] ), .A2(n1976), .ZN(n1645) );
  AND2_X2 U1639 ( .A1(n2565), .A2(net11558), .ZN(n1646) );
  AND2_X2 U1640 ( .A1(net85786), .A2(net85712), .ZN(n1647) );
  AND3_X4 U1641 ( .A1(n2338), .A2(n2494), .A3(n2490), .ZN(n1648) );
  AND2_X2 U1642 ( .A1(n2928), .A2(n2929), .ZN(n1649) );
  AND2_X4 U1643 ( .A1(n1550), .A2(n1612), .ZN(n1651) );
  NAND2_X2 U1644 ( .A1(\sub_435_b0/carry [10]), .A2(n1558), .ZN(n1653) );
  NAND2_X1 U1645 ( .A1(net89073), .A2(net84568), .ZN(n1654) );
  AND3_X4 U1646 ( .A1(n3132), .A2(n3131), .A3(n2767), .ZN(n1655) );
  INV_X4 U1647 ( .A(net84984), .ZN(net85006) );
  AND4_X4 U1648 ( .A1(n1769), .A2(n1770), .A3(n1771), .A4(net84118), .ZN(n1661) );
  AND3_X4 U1649 ( .A1(n2565), .A2(net83963), .A3(n2564), .ZN(n1662) );
  OR2_X4 U1650 ( .A1(n2991), .A2(net85832), .ZN(n1664) );
  AND2_X2 U1651 ( .A1(\u4/exp_f2i_1 [26]), .A2(n1606), .ZN(n1665) );
  NAND2_X2 U1652 ( .A1(\sub_435_3/carry [20]), .A2(n1635), .ZN(n1666) );
  NAND3_X2 U1653 ( .A1(n2872), .A2(n2854), .A3(n2853), .ZN(n2869) );
  AND2_X2 U1654 ( .A1(net83393), .A2(net83392), .ZN(n1669) );
  OR2_X4 U1655 ( .A1(underflow_fmul_r[1]), .A2(n1612), .ZN(n1670) );
  NAND3_X2 U1656 ( .A1(n2169), .A2(n2168), .A3(n2322), .ZN(net84774) );
  NAND2_X2 U1657 ( .A1(n3085), .A2(n3086), .ZN(net83791) );
  XNOR2_X1 U1658 ( .A(net83968), .B(\u4/add_407/carry [3]), .ZN(n1687) );
  XNOR2_X1 U1659 ( .A(exp_r[4]), .B(\u4/add_407/carry [4]), .ZN(n1688) );
  NAND3_X1 U1660 ( .A1(n3134), .A2(n3136), .A3(n2833), .ZN(n2757) );
  MUX2_X2 U1661 ( .A(\u2/N29 ), .B(\u2/N23 ), .S(n3136), .Z(n3134) );
  NAND3_X2 U1662 ( .A1(n2733), .A2(n2734), .A3(n2735), .ZN(\u2/N44 ) );
  NOR2_X2 U1663 ( .A1(n3142), .A2(n2754), .ZN(n2755) );
  NOR2_X2 U1664 ( .A1(n3141), .A2(n2754), .ZN(n2748) );
  NOR2_X2 U1665 ( .A1(n3140), .A2(n2754), .ZN(n2743) );
  NOR2_X2 U1666 ( .A1(n3139), .A2(n2754), .ZN(n2736) );
  NOR2_X2 U1667 ( .A1(n3138), .A2(n2754), .ZN(n2731) );
  INV_X2 U1668 ( .A(n3143), .ZN(\u2/exp_ovf_d[1] ) );
  INV_X2 U1669 ( .A(\u2/lt_130/A[3] ), .ZN(\u2/exp_tmp4[3] ) );
  OR2_X2 U1670 ( .A1(\u2/lt_130/A[3] ), .A2(\u2/add_111/carry[3] ), .ZN(
        \u2/add_111/carry[4] ) );
  AND2_X2 U1671 ( .A1(\u2/sub_111/carry[3] ), .A2(\u2/lt_130/A[3] ), .ZN(
        \u2/sub_111/carry[4] ) );
  MUX2_X2 U1672 ( .A(\u2/N15 ), .B(\u2/N9 ), .S(n3136), .Z(\u2/lt_130/A[3] )
         );
  MUX2_X2 U1673 ( .A(\u2/N10 ), .B(\u2/N16 ), .S(n3124), .Z(n1689) );
  OR2_X2 U1674 ( .A1(n1689), .A2(\u2/sub_111/carry[4] ), .ZN(
        \u2/sub_111/carry[5] ) );
  AND2_X2 U1675 ( .A1(\u2/add_111/carry[4] ), .A2(\u2/exp_tmp4[4] ), .ZN(
        \u2/add_111/carry[5] ) );
  NOR2_X1 U1676 ( .A1(n2753), .A2(n1622), .ZN(n2732) );
  NOR2_X2 U1677 ( .A1(n2753), .A2(n1630), .ZN(n2737) );
  NOR2_X2 U1678 ( .A1(n2753), .A2(n2742), .ZN(n2744) );
  NOR2_X2 U1679 ( .A1(n2753), .A2(n3018), .ZN(n2749) );
  NOR2_X2 U1680 ( .A1(n2753), .A2(\u2/exp_tmp4[0] ), .ZN(n2756) );
  NAND2_X4 U1681 ( .A1(n2730), .A2(n3124), .ZN(n2753) );
  NOR2_X2 U1682 ( .A1(n2732), .A2(n2731), .ZN(n2735) );
  MUX2_X2 U1683 ( .A(\u2/N10 ), .B(\u2/N16 ), .S(n3124), .Z(\u2/exp_tmp4[4] )
         );
  NOR4_X2 U1684 ( .A1(n3138), .A2(n3136), .A3(opa_r[14]), .A4(n1733), .ZN(
        n3144) );
  NOR2_X4 U1685 ( .A1(n3134), .A2(n3144), .ZN(n3143) );
  NOR3_X1 U1686 ( .A1(n2785), .A2(n2783), .A3(n2784), .ZN(n2786) );
  INV_X8 U1687 ( .A(n2954), .ZN(n1980) );
  INV_X8 U1688 ( .A(n2875), .ZN(n1718) );
  INV_X4 U1689 ( .A(n2875), .ZN(\u1/exp_diff_sft[0] ) );
  AOI21_X2 U1690 ( .B1(n2868), .B2(n2867), .A(n2874), .ZN(n2880) );
  INV_X2 U1691 ( .A(n1718), .ZN(n1719) );
  NOR2_X1 U1692 ( .A1(n1594), .A2(n1560), .ZN(n1988) );
  NOR2_X2 U1693 ( .A1(n2763), .A2(n1594), .ZN(\u2/exp_ovf_d[0] ) );
  NAND2_X2 U1694 ( .A1(opb_r[12]), .A2(n1573), .ZN(n2770) );
  NAND2_X4 U1695 ( .A1(n2822), .A2(n2821), .ZN(n2823) );
  MUX2_X2 U1696 ( .A(n1721), .B(n3102), .S(n1976), .Z(n1720) );
  INV_X4 U1697 ( .A(n1720), .ZN(n2947) );
  OAI21_X4 U1698 ( .B1(n2836), .B2(n2829), .A(n1722), .ZN(n3301) );
  CLKBUF_X2 U1699 ( .A(n2837), .Z(n1722) );
  INV_X4 U1700 ( .A(n3300), .ZN(n2876) );
  NAND2_X1 U1701 ( .A1(n2866), .A2(n3300), .ZN(n2867) );
  AOI21_X1 U1702 ( .B1(n2870), .B2(n2857), .A(n3302), .ZN(n2878) );
  NAND2_X4 U1703 ( .A1(n2837), .A2(n2838), .ZN(n2875) );
  NAND2_X1 U1704 ( .A1(opa_r[14]), .A2(n1734), .ZN(n2789) );
  NAND2_X4 U1705 ( .A1(n1594), .A2(opb_r[14]), .ZN(n2780) );
  NOR2_X2 U1706 ( .A1(opb_r[10]), .A2(n1723), .ZN(n2772) );
  NAND3_X1 U1707 ( .A1(opa_r[12]), .A2(n1988), .A3(n1987), .ZN(n3158) );
  OAI211_X4 U1708 ( .C1(n2883), .C2(n2950), .A(n2925), .B(n2923), .ZN(n2886)
         );
  NOR2_X2 U1709 ( .A1(n2887), .A2(n2945), .ZN(n2892) );
  OAI211_X4 U1710 ( .C1(n2886), .C2(n1563), .A(n2885), .B(n2884), .ZN(n2893)
         );
  OAI211_X4 U1711 ( .C1(n2903), .C2(n2902), .A(n2901), .B(n2900), .ZN(n2909)
         );
  INV_X8 U1712 ( .A(n2791), .ZN(n2793) );
  MUX2_X1 U1713 ( .A(n2878), .B(n2877), .S(n2876), .Z(n2879) );
  NOR2_X2 U1714 ( .A1(opa_r[10]), .A2(opa_r[11]), .ZN(n1983) );
  NAND2_X4 U1715 ( .A1(n2790), .A2(n2789), .ZN(n2926) );
  INV_X1 U1716 ( .A(fracta_mul[1]), .ZN(n3049) );
  INV_X16 U1717 ( .A(n1980), .ZN(n1979) );
  NOR2_X1 U1718 ( .A1(n3016), .A2(n1726), .ZN(n1985) );
  OR2_X4 U1719 ( .A1(n1726), .A2(opa_r[10]), .ZN(\u2/sub_110/carry [1]) );
  AND2_X2 U1720 ( .A1(n1727), .A2(n1728), .ZN(n1981) );
  NOR2_X1 U1721 ( .A1(n2779), .A2(n2791), .ZN(n2787) );
  NOR2_X1 U1722 ( .A1(n2927), .A2(n2791), .ZN(n2953) );
  NAND2_X4 U1723 ( .A1(n2882), .A2(n2791), .ZN(n2925) );
  AOI21_X1 U1724 ( .B1(n1718), .B2(n2865), .A(n2864), .ZN(n2868) );
  NAND2_X1 U1725 ( .A1(n1718), .A2(n3308), .ZN(n2870) );
  INV_X4 U1726 ( .A(n1729), .ZN(n1982) );
  NAND3_X1 U1727 ( .A1(n1982), .A2(n1726), .A3(n1981), .ZN(n1731) );
  NAND3_X2 U1728 ( .A1(n1982), .A2(n1726), .A3(n1981), .ZN(\u6/N10 ) );
  NAND2_X1 U1729 ( .A1(opb_r[10]), .A2(n1723), .ZN(n2781) );
  AND2_X2 U1730 ( .A1(opa_r[10]), .A2(opb_r[10]), .ZN(\u2/add_110/carry [1])
         );
  INV_X1 U1731 ( .A(opb_r[14]), .ZN(n1732) );
  INV_X4 U1732 ( .A(n1732), .ZN(n1733) );
  INV_X1 U1733 ( .A(n1731), .ZN(n3013) );
  NOR2_X1 U1734 ( .A1(n3313), .A2(n1731), .ZN(n2836) );
  NOR2_X1 U1735 ( .A1(opa_r[14]), .A2(n1731), .ZN(n2768) );
  OAI22_X1 U1736 ( .A1(n3130), .A2(n1731), .B1(n3129), .B2(n3313), .ZN(n2765)
         );
  NAND2_X1 U1737 ( .A1(n3313), .A2(n1731), .ZN(n2833) );
  NOR2_X1 U1738 ( .A1(opb_r[13]), .A2(n1560), .ZN(n2778) );
  NAND2_X1 U1739 ( .A1(opb_r[13]), .A2(n1560), .ZN(n2769) );
  NAND3_X1 U1740 ( .A1(opb_r[12]), .A2(n1986), .A3(n1985), .ZN(n3157) );
  NOR2_X1 U1741 ( .A1(opa_r[14]), .A2(n1733), .ZN(n2766) );
  INV_X1 U1742 ( .A(opb_r[13]), .ZN(n3017) );
  AOI21_X2 U1743 ( .B1(net83863), .B2(net83862), .A(net83864), .ZN(n2627) );
  INV_X8 U1744 ( .A(n2708), .ZN(n2665) );
  INV_X4 U1745 ( .A(n2707), .ZN(n2626) );
  AND2_X2 U1746 ( .A1(n2623), .A2(n2433), .ZN(n1736) );
  AOI211_X4 U1747 ( .C1(n2337), .C2(n1925), .A(n2335), .B(n2334), .ZN(n2348)
         );
  NAND3_X2 U1748 ( .A1(net84315), .A2(net84263), .A3(net84366), .ZN(n2419) );
  OAI211_X1 U1749 ( .C1(n2422), .C2(n2421), .A(n1597), .B(net84263), .ZN(n2423) );
  NAND2_X4 U1750 ( .A1(n2358), .A2(n2357), .ZN(net84263) );
  OAI21_X2 U1751 ( .B1(n2596), .B2(n2326), .A(n2325), .ZN(n2329) );
  INV_X2 U1752 ( .A(n2596), .ZN(n2613) );
  OR3_X4 U1753 ( .A1(n2540), .A2(net84012), .A3(n2539), .ZN(n1742) );
  NAND2_X4 U1754 ( .A1(n2524), .A2(n2523), .ZN(net84059) );
  NAND3_X4 U1755 ( .A1(fract_out_q[5]), .A2(net85730), .A3(net85718), .ZN(
        n2023) );
  OAI21_X4 U1756 ( .B1(net88618), .B2(net89546), .A(net84758), .ZN(n1900) );
  NAND3_X4 U1757 ( .A1(net85227), .A2(n1744), .A3(net85678), .ZN(net85061) );
  INV_X32 U1758 ( .A(net85754), .ZN(net85752) );
  INV_X4 U1759 ( .A(net84677), .ZN(net86171) );
  INV_X8 U1760 ( .A(\u4/fract_out_pl1[10] ), .ZN(net84677) );
  NAND2_X2 U1761 ( .A1(net83863), .A2(net83862), .ZN(net83870) );
  INV_X8 U1762 ( .A(net85290), .ZN(net85240) );
  OAI21_X4 U1763 ( .B1(n2672), .B2(n2673), .A(n2671), .ZN(N285) );
  INV_X2 U1764 ( .A(n1915), .ZN(n2365) );
  NAND3_X2 U1765 ( .A1(n1915), .A2(n2425), .A3(net85794), .ZN(net84079) );
  NAND3_X2 U1766 ( .A1(n1915), .A2(n2566), .A3(n1632), .ZN(n2486) );
  NAND3_X2 U1767 ( .A1(n2555), .A2(n1915), .A3(n1632), .ZN(n2482) );
  INV_X8 U1768 ( .A(n2997), .ZN(n2996) );
  NAND2_X4 U1769 ( .A1(n2456), .A2(n2997), .ZN(net84072) );
  NAND2_X4 U1770 ( .A1(n2358), .A2(n2357), .ZN(n2997) );
  NOR2_X4 U1771 ( .A1(net84055), .A2(n1806), .ZN(n1805) );
  NAND2_X1 U1772 ( .A1(n2433), .A2(n2689), .ZN(n2690) );
  NAND2_X4 U1773 ( .A1(net89595), .A2(net84584), .ZN(net84553) );
  INV_X8 U1774 ( .A(net84553), .ZN(net84574) );
  OAI211_X4 U1775 ( .C1(n1841), .C2(n1843), .A(net84149), .B(net85842), .ZN(
        n1840) );
  INV_X32 U1776 ( .A(n1960), .ZN(n1961) );
  NAND2_X4 U1777 ( .A1(net83934), .A2(net84571), .ZN(net84648) );
  NAND2_X4 U1778 ( .A1(net84552), .A2(n1638), .ZN(n2356) );
  NOR2_X2 U1779 ( .A1(net85736), .A2(net85720), .ZN(net85297) );
  XNOR2_X2 U1780 ( .A(net84136), .B(net30297), .ZN(n2370) );
  INV_X1 U1781 ( .A(net85998), .ZN(net90217) );
  NAND3_X2 U1782 ( .A1(n1942), .A2(quo[1]), .A3(net85684), .ZN(n1743) );
  NAND3_X2 U1783 ( .A1(n1894), .A2(quo[1]), .A3(net85684), .ZN(net85261) );
  OAI21_X4 U1784 ( .B1(net85373), .B2(net85676), .A(net85374), .ZN(n1914) );
  NAND2_X4 U1785 ( .A1(net89129), .A2(quo[7]), .ZN(net85373) );
  INV_X4 U1786 ( .A(net85748), .ZN(n1744) );
  NOR2_X1 U1787 ( .A1(net84060), .A2(net83875), .ZN(n1804) );
  INV_X1 U1788 ( .A(net84471), .ZN(n1747) );
  AOI21_X4 U1789 ( .B1(n2355), .B2(net84214), .A(n2354), .ZN(n2374) );
  NAND3_X1 U1790 ( .A1(net85847), .A2(n2588), .A3(net83861), .ZN(n2354) );
  INV_X4 U1791 ( .A(net86171), .ZN(net91353) );
  NAND3_X4 U1792 ( .A1(net84343), .A2(net86171), .A3(net84334), .ZN(net84371)
         );
  NOR2_X2 U1793 ( .A1(n2350), .A2(n2349), .ZN(n2355) );
  OAI21_X4 U1794 ( .B1(net90047), .B2(n1623), .A(n1756), .ZN(net85021) );
  INV_X8 U1795 ( .A(net86165), .ZN(net90047) );
  NOR2_X1 U1796 ( .A1(n2541), .A2(n2441), .ZN(net83862) );
  NAND2_X1 U1797 ( .A1(n1849), .A2(net88721), .ZN(n1750) );
  OAI22_X4 U1798 ( .A1(net84322), .A2(n1961), .B1(n1928), .B2(n2386), .ZN(
        n2515) );
  OAI22_X4 U1799 ( .A1(net89716), .A2(n1961), .B1(n1928), .B2(n2508), .ZN(
        n2685) );
  INV_X4 U1800 ( .A(net84523), .ZN(n1766) );
  NOR3_X4 U1801 ( .A1(n2678), .A2(n2676), .A3(n2680), .ZN(n2517) );
  NAND2_X4 U1802 ( .A1(net84846), .A2(n1753), .ZN(n1752) );
  OR2_X2 U1803 ( .A1(net84778), .A2(net84845), .ZN(n1753) );
  NAND2_X2 U1804 ( .A1(\u4/N426 ), .A2(net84522), .ZN(n1754) );
  NAND2_X4 U1805 ( .A1(\u4/N426 ), .A2(net84522), .ZN(n1899) );
  NAND2_X1 U1806 ( .A1(div_opa_ldz_r2[1]), .A2(net84901), .ZN(n2103) );
  INV_X16 U1807 ( .A(net84982), .ZN(net83933) );
  NAND2_X4 U1808 ( .A1(net11555), .A2(net85033), .ZN(net84982) );
  INV_X8 U1809 ( .A(net83421), .ZN(\u4/exp_in_pl1[2] ) );
  NAND2_X2 U1810 ( .A1(net88636), .A2(net85089), .ZN(n1755) );
  INV_X8 U1811 ( .A(net86026), .ZN(net88636) );
  INV_X1 U1812 ( .A(net84895), .ZN(n1757) );
  INV_X1 U1813 ( .A(net85790), .ZN(n1758) );
  NAND2_X1 U1814 ( .A1(n1757), .A2(n1758), .ZN(n1756) );
  NAND2_X4 U1815 ( .A1(net85296), .A2(n1759), .ZN(net85161) );
  NAND2_X2 U1816 ( .A1(n2001), .A2(n1760), .ZN(n1759) );
  INV_X16 U1817 ( .A(n1880), .ZN(n1879) );
  BUF_X32 U1818 ( .A(net84909), .Z(net90035) );
  NAND4_X4 U1819 ( .A1(net85061), .A2(n2043), .A3(n2067), .A4(n2066), .ZN(
        n3004) );
  AOI21_X2 U1820 ( .B1(net90302), .B2(net89372), .A(net83407), .ZN(net84502)
         );
  INV_X2 U1821 ( .A(net89965), .ZN(net89372) );
  INV_X2 U1822 ( .A(net84755), .ZN(net89121) );
  OAI22_X4 U1823 ( .A1(n1928), .A2(n2506), .B1(net84118), .B2(n1961), .ZN(
        n2691) );
  OAI22_X4 U1824 ( .A1(net84103), .A2(n1961), .B1(n1928), .B2(n2512), .ZN(
        n2674) );
  OAI22_X4 U1825 ( .A1(n1555), .A2(n1961), .B1(n2513), .B2(n2509), .ZN(n2676)
         );
  NAND2_X2 U1826 ( .A1(net84199), .A2(net84200), .ZN(n2457) );
  AOI21_X4 U1827 ( .B1(n1580), .B2(n1529), .A(net84390), .ZN(n1762) );
  AOI211_X2 U1828 ( .C1(net85842), .C2(net84386), .A(net84387), .B(n1762), 
        .ZN(net84199) );
  INV_X1 U1829 ( .A(net84808), .ZN(n1771) );
  INV_X8 U1830 ( .A(net84014), .ZN(net85846) );
  NAND2_X4 U1831 ( .A1(net85028), .A2(n1744), .ZN(net84014) );
  BUF_X16 U1832 ( .A(net84570), .Z(net89029) );
  INV_X2 U1833 ( .A(net84059), .ZN(n1808) );
  NAND4_X1 U1834 ( .A1(n2164), .A2(n2166), .A3(n2167), .A4(n2165), .ZN(n1763)
         );
  INV_X4 U1835 ( .A(net84565), .ZN(n1764) );
  NAND4_X2 U1836 ( .A1(n2165), .A2(n2166), .A3(n2167), .A4(n2164), .ZN(
        net84523) );
  INV_X4 U1837 ( .A(n1763), .ZN(net84565) );
  INV_X4 U1838 ( .A(net84472), .ZN(net89664) );
  NAND2_X4 U1839 ( .A1(net84674), .A2(net83429), .ZN(net84472) );
  INV_X4 U1840 ( .A(net83787), .ZN(net83819) );
  NAND4_X2 U1841 ( .A1(net84569), .A2(net84648), .A3(net99831), .A4(net84649), 
        .ZN(net84644) );
  NAND2_X4 U1842 ( .A1(net84381), .A2(n1554), .ZN(net30297) );
  OAI21_X4 U1843 ( .B1(net84574), .B2(net84575), .A(net84576), .ZN(net84381)
         );
  NAND3_X2 U1844 ( .A1(net84554), .A2(net84553), .A3(net84403), .ZN(net84552)
         );
  OAI21_X4 U1845 ( .B1(net91375), .B2(net85017), .A(net84967), .ZN(net84870)
         );
  NAND2_X4 U1846 ( .A1(n2520), .A2(n2459), .ZN(n2460) );
  INV_X1 U1847 ( .A(n2521), .ZN(n2459) );
  OAI21_X4 U1848 ( .B1(n2528), .B2(n2502), .A(net83861), .ZN(net84010) );
  NAND2_X4 U1849 ( .A1(n2351), .A2(net84149), .ZN(net84214) );
  OAI21_X4 U1850 ( .B1(n1766), .B2(n1765), .A(net84649), .ZN(net84573) );
  INV_X1 U1851 ( .A(net91325), .ZN(n1765) );
  NOR2_X2 U1852 ( .A1(net89664), .A2(net84676), .ZN(net89663) );
  AOI21_X2 U1853 ( .B1(net84070), .B2(net84069), .A(sign_fasu_r), .ZN(n1810)
         );
  INV_X4 U1854 ( .A(net83868), .ZN(net84069) );
  NAND4_X1 U1855 ( .A1(net84150), .A2(net84081), .A3(n2478), .A4(net84169), 
        .ZN(n2345) );
  INV_X8 U1856 ( .A(net84220), .ZN(net84081) );
  NAND3_X1 U1857 ( .A1(net83950), .A2(n2302), .A3(\u4/fract_out_pl1[10] ), 
        .ZN(net84398) );
  INV_X8 U1858 ( .A(net84458), .ZN(net83950) );
  OAI21_X4 U1859 ( .B1(net89663), .B2(\u4/exp_out[4] ), .A(net84014), .ZN(
        net84588) );
  NAND3_X2 U1860 ( .A1(n1767), .A2(net85337), .A3(net85210), .ZN(n3001) );
  INV_X1 U1861 ( .A(net85336), .ZN(n1767) );
  NAND2_X4 U1862 ( .A1(n1951), .A2(n1950), .ZN(net84753) );
  NAND3_X4 U1863 ( .A1(n1768), .A2(n2365), .A3(rmode_r3[0]), .ZN(net84135) );
  AND2_X2 U1864 ( .A1(n1764), .A2(net84522), .ZN(n1823) );
  AOI211_X4 U1865 ( .C1(sign), .C2(net84403), .A(net84480), .B(net84675), .ZN(
        net84409) );
  INV_X1 U1866 ( .A(net84456), .ZN(n1769) );
  INV_X1 U1867 ( .A(\u4/fract_out[8] ), .ZN(n1770) );
  INV_X4 U1868 ( .A(net84676), .ZN(net84471) );
  NAND2_X4 U1869 ( .A1(n1772), .A2(net89842), .ZN(net89224) );
  INV_X1 U1870 ( .A(net84956), .ZN(n1772) );
  AOI21_X4 U1871 ( .B1(net84588), .B2(net84468), .A(n1824), .ZN(net84483) );
  INV_X8 U1872 ( .A(net84015), .ZN(net84468) );
  AOI211_X4 U1873 ( .C1(\u4/exp_f2i_1 [25]), .C2(n1606), .A(net83406), .B(
        n1773), .ZN(net83392) );
  OAI21_X4 U1874 ( .B1(n1774), .B2(n1775), .A(n1776), .ZN(n1773) );
  NOR2_X1 U1875 ( .A1(net88427), .A2(net83403), .ZN(n1777) );
  INV_X8 U1876 ( .A(opb_dn), .ZN(net88427) );
  NAND2_X2 U1877 ( .A1(net83416), .A2(net83417), .ZN(n1775) );
  INV_X4 U1878 ( .A(net83403), .ZN(net83417) );
  AOI211_X2 U1879 ( .C1(net83417), .C2(net84615), .A(n1665), .B(net84617), 
        .ZN(net84614) );
  AOI211_X4 U1880 ( .C1(net84655), .C2(net83417), .A(net84656), .B(net84657), 
        .ZN(net84654) );
  INV_X4 U1881 ( .A(net84611), .ZN(net83416) );
  NAND2_X2 U1882 ( .A1(net83416), .A2(net84667), .ZN(net84660) );
  NAND2_X2 U1883 ( .A1(net83416), .A2(net84629), .ZN(net84625) );
  NAND2_X4 U1884 ( .A1(n1785), .A2(n1786), .ZN(n1774) );
  NAND2_X4 U1885 ( .A1(n1783), .A2(n1784), .ZN(n1786) );
  INV_X8 U1886 ( .A(n1778), .ZN(n1784) );
  INV_X2 U1887 ( .A(n1784), .ZN(net90268) );
  INV_X8 U1888 ( .A(n1780), .ZN(n1778) );
  NAND2_X2 U1889 ( .A1(n1778), .A2(net83419), .ZN(n1785) );
  OAI21_X4 U1890 ( .B1(net85710), .B2(n1779), .A(n1781), .ZN(n1780) );
  NAND2_X4 U1891 ( .A1(net85313), .A2(n1782), .ZN(\u4/f2i_shft[1] ) );
  INV_X4 U1892 ( .A(net85030), .ZN(n1782) );
  INV_X4 U1893 ( .A(net84761), .ZN(n1779) );
  NOR2_X1 U1894 ( .A1(net89924), .A2(n1779), .ZN(net83987) );
  XNOR2_X2 U1895 ( .A(n1779), .B(net85710), .ZN(net84668) );
  INV_X32 U1896 ( .A(net85712), .ZN(net85710) );
  NAND2_X2 U1897 ( .A1(n1787), .A2(net91144), .ZN(\u4/N655 ) );
  INV_X4 U1898 ( .A(net90079), .ZN(net91144) );
  BUF_X32 U1899 ( .A(net90079), .Z(net91404) );
  NOR2_X4 U1900 ( .A1(n1789), .A2(n1790), .ZN(n1788) );
  NAND2_X4 U1901 ( .A1(n845), .A2(net84637), .ZN(n1790) );
  NOR2_X4 U1902 ( .A1(n1791), .A2(net83945), .ZN(n1789) );
  OR2_X4 U1903 ( .A1(net85788), .A2(net83951), .ZN(n1791) );
  INV_X16 U1904 ( .A(net76872), .ZN(net85788) );
  INV_X4 U1905 ( .A(net84658), .ZN(net84657) );
  NAND2_X4 U1906 ( .A1(\u4/exp_f2i_1 [24]), .A2(n1606), .ZN(net84658) );
  INV_X4 U1907 ( .A(net85847), .ZN(net83941) );
  AOI22_X1 U1908 ( .A1(n1574), .A2(n1744), .B1(n1550), .B2(n1670), .ZN(
        net83827) );
  INV_X1 U1909 ( .A(n1744), .ZN(net90287) );
  INV_X16 U1910 ( .A(net85752), .ZN(net85746) );
  INV_X32 U1911 ( .A(net85752), .ZN(net85744) );
  INV_X16 U1912 ( .A(net85756), .ZN(net85754) );
  INV_X4 U1913 ( .A(net11675), .ZN(net85756) );
  INV_X4 U1914 ( .A(net85323), .ZN(net85028) );
  NAND2_X1 U1915 ( .A1(net85028), .A2(net91548), .ZN(net84341) );
  NAND2_X4 U1916 ( .A1(net85028), .A2(n1643), .ZN(net85320) );
  NAND2_X4 U1917 ( .A1(net85730), .A2(net85722), .ZN(net85323) );
  INV_X16 U1918 ( .A(net85724), .ZN(net85722) );
  INV_X16 U1919 ( .A(net85726), .ZN(net85724) );
  INV_X16 U1920 ( .A(net85724), .ZN(net85720) );
  INV_X4 U1921 ( .A(net11677), .ZN(net85726) );
  INV_X16 U1922 ( .A(net85738), .ZN(net85730) );
  INV_X32 U1923 ( .A(net85740), .ZN(net85738) );
  INV_X16 U1924 ( .A(net85742), .ZN(net85740) );
  INV_X8 U1925 ( .A(net85740), .ZN(net85736) );
  INV_X4 U1926 ( .A(net11676), .ZN(net85742) );
  NAND2_X4 U1927 ( .A1(net84471), .A2(net84472), .ZN(\u4/exp_out[4] ) );
  NAND2_X4 U1928 ( .A1(net89657), .A2(net89736), .ZN(n1794) );
  NAND2_X4 U1929 ( .A1(n1793), .A2(net83398), .ZN(net89736) );
  INV_X4 U1930 ( .A(net89736), .ZN(net88646) );
  INV_X4 U1931 ( .A(net84606), .ZN(net83398) );
  AOI21_X2 U1932 ( .B1(net84663), .B2(net83398), .A(net84664), .ZN(net84662)
         );
  NOR3_X1 U1933 ( .A1(net85790), .A2(net83398), .A3(net83951), .ZN(net84591)
         );
  NAND3_X1 U1934 ( .A1(net89919), .A2(net84766), .A3(net83398), .ZN(net84642)
         );
  AOI21_X4 U1935 ( .B1(\u4/exp_next_mi[1] ), .B2(net85788), .A(n1647), .ZN(
        n1793) );
  INV_X32 U1936 ( .A(net85788), .ZN(net85786) );
  AOI22_X4 U1937 ( .A1(\u4/exp_in_pl1[2] ), .A2(net85786), .B1(
        \u4/exp_next_mi[2] ), .B2(net85788), .ZN(n1792) );
  NAND2_X1 U1938 ( .A1(\u4/exp_in_pl1[2] ), .A2(net110951), .ZN(net84298) );
  NOR2_X1 U1939 ( .A1(\u4/exp_in_pl1[2] ), .A2(net110951), .ZN(net84297) );
  NAND3_X1 U1940 ( .A1(net77815), .A2(net84606), .A3(net84633), .ZN(net84661)
         );
  NOR2_X1 U1941 ( .A1(net83402), .A2(net84606), .ZN(net84605) );
  BUF_X32 U1942 ( .A(\u4/exp_next_mi[1] ), .Z(net89692) );
  NAND2_X2 U1943 ( .A1(\u4/exp_next_mi[1] ), .A2(net85788), .ZN(net91056) );
  INV_X4 U1944 ( .A(net85313), .ZN(net85316) );
  XNOR2_X2 U1945 ( .A(net85313), .B(net11560), .ZN(net83421) );
  NOR2_X1 U1946 ( .A1(net85030), .A2(net11560), .ZN(net84916) );
  BUF_X32 U1947 ( .A(\u4/exp_next_mi[2] ), .Z(net89948) );
  MUX2_X2 U1948 ( .A(\u4/exp_next_mi[0] ), .B(net85778), .S(net76872), .Z(
        net84606) );
  NAND2_X1 U1949 ( .A1(net85712), .A2(net76872), .ZN(net91057) );
  BUF_X32 U1950 ( .A(\u4/exp_out[2] ), .Z(net86169) );
  NAND2_X2 U1951 ( .A1(net83849), .A2(net84236), .ZN(net83402) );
  INV_X8 U1952 ( .A(net83813), .ZN(net83849) );
  NAND2_X2 U1953 ( .A1(net84669), .A2(net86067), .ZN(net83403) );
  INV_X4 U1954 ( .A(net84452), .ZN(net84674) );
  OAI21_X4 U1955 ( .B1(net84678), .B2(net84677), .A(net84451), .ZN(net84676)
         );
  INV_X4 U1956 ( .A(net84679), .ZN(net84451) );
  NAND2_X2 U1957 ( .A1(net84451), .A2(net84452), .ZN(net84450) );
  OAI21_X2 U1958 ( .B1(net85794), .B2(net83995), .A(n1795), .ZN(net84679) );
  AOI21_X2 U1959 ( .B1(\u4/exp_f2i_1 [27]), .B2(n1606), .A(n1796), .ZN(n1795)
         );
  NAND2_X1 U1960 ( .A1(n1797), .A2(net84637), .ZN(n1796) );
  NAND3_X1 U1961 ( .A1(net84639), .A2(net83990), .A3(net84683), .ZN(n1797) );
  INV_X4 U1962 ( .A(net83408), .ZN(net84683) );
  NAND2_X1 U1963 ( .A1(net84683), .A2(net90302), .ZN(net84659) );
  NAND2_X4 U1964 ( .A1(net84586), .A2(net84569), .ZN(net84769) );
  OAI21_X4 U1965 ( .B1(net84769), .B2(net84573), .A(net84770), .ZN(net84678)
         );
  NAND3_X2 U1966 ( .A1(net84570), .A2(net84572), .A3(net84571), .ZN(net84586)
         );
  INV_X4 U1967 ( .A(net84829), .ZN(net84571) );
  NAND2_X2 U1968 ( .A1(net83936), .A2(n1571), .ZN(net84829) );
  NOR4_X4 U1969 ( .A1(net84808), .A2(\u4/fract_out[8] ), .A3(n1752), .A4(
        net84456), .ZN(net84572) );
  INV_X4 U1970 ( .A(net84811), .ZN(net84570) );
  NAND3_X2 U1971 ( .A1(n1798), .A2(n1799), .A3(n1801), .ZN(net84811) );
  INV_X4 U1972 ( .A(net84814), .ZN(n1801) );
  NOR2_X4 U1973 ( .A1(\u4/fract_out[5] ), .A2(n1924), .ZN(n1799) );
  NAND2_X2 U1974 ( .A1(net89819), .A2(net84842), .ZN(\u4/fract_out[7] ) );
  NAND2_X4 U1975 ( .A1(net84836), .A2(n1802), .ZN(\u4/fract_out[4] ) );
  NAND2_X2 U1976 ( .A1(net91150), .A2(\u4/N404 ), .ZN(n1802) );
  OAI21_X4 U1977 ( .B1(net84778), .B2(n1800), .A(net84836), .ZN(net89933) );
  INV_X1 U1978 ( .A(net84778), .ZN(net91150) );
  NAND2_X4 U1979 ( .A1(\u4/N428 ), .A2(net84522), .ZN(net84836) );
  INV_X16 U1980 ( .A(net84566), .ZN(net84522) );
  NAND2_X4 U1981 ( .A1(net84774), .A2(net84775), .ZN(net84569) );
  NAND3_X1 U1982 ( .A1(net89073), .A2(net84568), .A3(net84569), .ZN(net84484)
         );
  NAND2_X4 U1983 ( .A1(net84908), .A2(net91112), .ZN(net83936) );
  INV_X4 U1984 ( .A(net84561), .ZN(net84908) );
  NAND2_X4 U1985 ( .A1(net84110), .A2(net84113), .ZN(net84808) );
  NAND4_X2 U1986 ( .A1(n1750), .A2(net84050), .A3(net84051), .A4(net84052), 
        .ZN(net84025) );
  NAND4_X2 U1987 ( .A1(net84024), .A2(n1804), .A3(n1805), .A4(net83819), .ZN(
        net84052) );
  NOR2_X4 U1988 ( .A1(sign_fasu_r), .A2(net83819), .ZN(n1809) );
  NAND2_X2 U1989 ( .A1(net84024), .A2(net83819), .ZN(net83883) );
  NAND2_X2 U1990 ( .A1(n1807), .A2(n1808), .ZN(n1806) );
  INV_X4 U1991 ( .A(net83747), .ZN(n1803) );
  NOR2_X1 U1992 ( .A1(net84015), .A2(n1803), .ZN(net84012) );
  NAND2_X2 U1993 ( .A1(net84064), .A2(net84044), .ZN(n1811) );
  NAND2_X2 U1994 ( .A1(nan_sign_d), .A2(n1581), .ZN(net84043) );
  NAND2_X2 U1995 ( .A1(net11627), .A2(n1611), .ZN(net83781) );
  INV_X32 U1996 ( .A(net85794), .ZN(net85790) );
  INV_X16 U1997 ( .A(net86067), .ZN(net85794) );
  NAND2_X2 U1998 ( .A1(net84619), .A2(net86067), .ZN(net83427) );
  INV_X4 U1999 ( .A(net83791), .ZN(net83779) );
  NAND2_X4 U2000 ( .A1(\u4/N433 ), .A2(net84522), .ZN(net84846) );
  NAND3_X2 U2001 ( .A1(net84847), .A2(net84848), .A3(n1812), .ZN(net84566) );
  NOR2_X1 U2002 ( .A1(net84565), .A2(net84566), .ZN(net84555) );
  OAI21_X4 U2003 ( .B1(net84830), .B2(net84566), .A(net84810), .ZN(net60630)
         );
  NAND2_X2 U2004 ( .A1(net84564), .A2(net84566), .ZN(net84519) );
  NAND2_X2 U2005 ( .A1(n1815), .A2(net84853), .ZN(n1814) );
  NAND2_X2 U2006 ( .A1(net84854), .A2(n1816), .ZN(n1815) );
  NAND2_X2 U2007 ( .A1(net11555), .A2(net11558), .ZN(n1816) );
  INV_X2 U2008 ( .A(net84856), .ZN(net84854) );
  INV_X4 U2009 ( .A(\u4/f2i_shft[4] ), .ZN(n1817) );
  NAND2_X1 U2010 ( .A1(n1818), .A2(net83439), .ZN(net89615) );
  OAI21_X1 U2011 ( .B1(net85828), .B2(net83849), .A(net83974), .ZN(n1818) );
  INV_X32 U2012 ( .A(net85827), .ZN(net85828) );
  INV_X4 U2013 ( .A(\u4/N656 ), .ZN(net86165) );
  NAND2_X2 U2014 ( .A1(net90997), .A2(net86165), .ZN(net110929) );
  NOR2_X4 U2015 ( .A1(net86165), .A2(n1621), .ZN(net91177) );
  NAND2_X4 U2016 ( .A1(net83813), .A2(n1571), .ZN(net83439) );
  NAND2_X2 U2017 ( .A1(net83849), .A2(n1571), .ZN(net83974) );
  OAI21_X4 U2018 ( .B1(net83973), .B2(net83974), .A(net83975), .ZN(net83972)
         );
  NAND2_X2 U2019 ( .A1(n1641), .A2(net88427), .ZN(net83813) );
  OAI211_X1 U2020 ( .C1(net83811), .C2(net83812), .A(net86038), .B(net83813), 
        .ZN(net83807) );
  NAND2_X1 U2021 ( .A1(opa_dn), .A2(net85676), .ZN(net84669) );
  NAND2_X2 U2022 ( .A1(opa_dn), .A2(net84722), .ZN(net84611) );
  NOR2_X4 U2023 ( .A1(net85718), .A2(net11582), .ZN(n1819) );
  AOI21_X4 U2024 ( .B1(net85297), .B2(fract_out_q[3]), .A(n1819), .ZN(net85296) );
  INV_X32 U2025 ( .A(net85720), .ZN(net85718) );
  AND2_X2 U2026 ( .A1(net99831), .A2(net84649), .ZN(net89073) );
  NAND2_X1 U2027 ( .A1(net91325), .A2(n1763), .ZN(net99831) );
  NAND2_X4 U2028 ( .A1(net84483), .A2(net84484), .ZN(net84401) );
  INV_X4 U2029 ( .A(n1820), .ZN(n1822) );
  AOI21_X1 U2030 ( .B1(net84518), .B2(net84519), .A(net84015), .ZN(n1820) );
  NAND3_X2 U2031 ( .A1(net84571), .A2(net83849), .A3(net85794), .ZN(n1821) );
  NAND3_X4 U2032 ( .A1(net84948), .A2(net89224), .A3(net84950), .ZN(
        \u4/shift_left [0]) );
  NOR2_X4 U2033 ( .A1(net85832), .A2(net84867), .ZN(n1825) );
  INV_X1 U2034 ( .A(\u4/div_shft2[0] ), .ZN(net85831) );
  NAND4_X2 U2035 ( .A1(net11562), .A2(net85831), .A3(net11558), .A4(net11560), 
        .ZN(net84279) );
  NOR2_X4 U2036 ( .A1(net88292), .A2(n1549), .ZN(net84953) );
  INV_X8 U2037 ( .A(net88287), .ZN(net86037) );
  NAND4_X1 U2038 ( .A1(net84996), .A2(net11566), .A3(net85788), .A4(net91375), 
        .ZN(net84990) );
  BUF_X32 U2039 ( .A(\u4/exp_next_mi[5] ), .Z(net91375) );
  NOR2_X4 U2040 ( .A1(net84957), .A2(net89055), .ZN(net84948) );
  NOR2_X4 U2041 ( .A1(n1827), .A2(n1826), .ZN(net89054) );
  NOR2_X2 U2042 ( .A1(net85778), .A2(net84856), .ZN(n1826) );
  NAND2_X4 U2043 ( .A1(net84960), .A2(n1828), .ZN(n1827) );
  NAND2_X4 U2044 ( .A1(net85015), .A2(net84963), .ZN(n1828) );
  INV_X4 U2045 ( .A(net11670), .ZN(net84963) );
  NAND2_X4 U2046 ( .A1(net84202), .A2(net88374), .ZN(net84201) );
  INV_X8 U2047 ( .A(net84201), .ZN(net88721) );
  NAND2_X4 U2048 ( .A1(net83875), .A2(n1829), .ZN(net88374) );
  INV_X8 U2049 ( .A(n1830), .ZN(n1829) );
  NAND3_X4 U2050 ( .A1(n1829), .A2(net83874), .A3(net83875), .ZN(net83871) );
  NAND2_X4 U2051 ( .A1(n1832), .A2(net83861), .ZN(n1830) );
  INV_X4 U2052 ( .A(net84206), .ZN(net83861) );
  NAND2_X2 U2053 ( .A1(net84085), .A2(net83736), .ZN(net84083) );
  AOI211_X4 U2054 ( .C1(n1833), .C2(net83870), .A(n1834), .B(net84204), .ZN(
        net84202) );
  NAND3_X4 U2055 ( .A1(net84074), .A2(n1607), .A3(net84200), .ZN(n1832) );
  NAND2_X4 U2056 ( .A1(n1832), .A2(n1831), .ZN(net83853) );
  AOI21_X2 U2057 ( .B1(n1607), .B2(net84003), .A(net83878), .ZN(n1831) );
  NOR3_X4 U2058 ( .A1(net84372), .A2(n1533), .A3(net84374), .ZN(net84074) );
  NAND2_X2 U2059 ( .A1(net84414), .A2(n1835), .ZN(net84206) );
  NAND2_X2 U2060 ( .A1(n1580), .A2(n1529), .ZN(net84138) );
  INV_X4 U2061 ( .A(net84473), .ZN(net84576) );
  NAND2_X2 U2062 ( .A1(net84474), .A2(net84475), .ZN(net84453) );
  NAND2_X2 U2063 ( .A1(n1554), .A2(net84473), .ZN(net84315) );
  XNOR2_X2 U2064 ( .A(net91555), .B(net11671), .ZN(net84763) );
  AOI22_X4 U2065 ( .A1(net85080), .A2(net85079), .B1(net85081), .B2(net91555), 
        .ZN(net33278) );
  INV_X8 U2066 ( .A(net85174), .ZN(net84758) );
  NAND2_X4 U2067 ( .A1(n1836), .A2(net85108), .ZN(net85174) );
  INV_X8 U2068 ( .A(net85178), .ZN(net85108) );
  NAND2_X2 U2069 ( .A1(net85108), .A2(net84550), .ZN(net85127) );
  NAND3_X4 U2070 ( .A1(net85112), .A2(net85113), .A3(net85108), .ZN(net85111)
         );
  NAND3_X4 U2071 ( .A1(net85176), .A2(net86262), .A3(net85128), .ZN(n1836) );
  INV_X8 U2072 ( .A(net85181), .ZN(net85128) );
  NAND2_X1 U2073 ( .A1(net85128), .A2(net86262), .ZN(net85115) );
  NAND2_X2 U2074 ( .A1(net86262), .A2(net85128), .ZN(net85133) );
  NAND4_X4 U2075 ( .A1(net85128), .A2(net86262), .A3(net85179), .A4(net85180), 
        .ZN(net85084) );
  NAND2_X4 U2076 ( .A1(n1837), .A2(net85220), .ZN(net85181) );
  INV_X8 U2077 ( .A(n1838), .ZN(n1837) );
  NAND2_X4 U2078 ( .A1(net85220), .A2(n1837), .ZN(net77045) );
  NAND3_X4 U2079 ( .A1(net85076), .A2(net85676), .A3(quo[21]), .ZN(n1839) );
  INV_X16 U2080 ( .A(net85678), .ZN(net85676) );
  INV_X16 U2081 ( .A(net85975), .ZN(net85678) );
  INV_X16 U2082 ( .A(net85678), .ZN(net85674) );
  NAND3_X4 U2083 ( .A1(net85342), .A2(quo[3]), .A3(net85678), .ZN(net85051) );
  INV_X4 U2084 ( .A(net85974), .ZN(net85975) );
  INV_X8 U2085 ( .A(net85975), .ZN(net85684) );
  INV_X8 U2086 ( .A(net85351), .ZN(net85076) );
  NAND2_X4 U2087 ( .A1(fract_out_q[12]), .A2(net83780), .ZN(net85349) );
  INV_X8 U2088 ( .A(net85387), .ZN(net83780) );
  NAND2_X4 U2089 ( .A1(net85998), .A2(net85718), .ZN(net85387) );
  NAND2_X4 U2090 ( .A1(net85083), .A2(net85082), .ZN(net84757) );
  INV_X2 U2091 ( .A(net84757), .ZN(net89411) );
  INV_X8 U2092 ( .A(net85084), .ZN(net85082) );
  INV_X8 U2093 ( .A(net76645), .ZN(net85180) );
  INV_X4 U2094 ( .A(n1909), .ZN(net89624) );
  INV_X4 U2095 ( .A(net76254), .ZN(net85179) );
  INV_X1 U2096 ( .A(net85179), .ZN(net86004) );
  INV_X8 U2097 ( .A(net76352), .ZN(net86262) );
  NAND3_X2 U2098 ( .A1(net85247), .A2(net90019), .A3(net85248), .ZN(net76352)
         );
  NAND3_X2 U2099 ( .A1(net85076), .A2(net85676), .A3(quo[22]), .ZN(net85248)
         );
  INV_X4 U2100 ( .A(net85384), .ZN(net85077) );
  NAND2_X2 U2101 ( .A1(net85738), .A2(net85748), .ZN(net85384) );
  INV_X16 U2102 ( .A(net85752), .ZN(net85748) );
  OAI21_X4 U2103 ( .B1(net84974), .B2(net84975), .A(net89372), .ZN(net84956)
         );
  OAI211_X4 U2104 ( .C1(net84967), .C2(net84956), .A(net84968), .B(net84969), 
        .ZN(net84957) );
  NAND2_X4 U2105 ( .A1(\u4/exp_next_mi[5] ), .A2(net85788), .ZN(net84983) );
  INV_X2 U2106 ( .A(n1530), .ZN(net84967) );
  INV_X1 U2107 ( .A(net84975), .ZN(net85017) );
  MUX2_X2 U2108 ( .A(net84598), .B(net84599), .S(net89965), .Z(net84595) );
  NAND2_X1 U2109 ( .A1(net89965), .A2(net85778), .ZN(net84166) );
  NAND2_X4 U2110 ( .A1(net89917), .A2(net89077), .ZN(net84372) );
  INV_X4 U2111 ( .A(net89076), .ZN(net89077) );
  NAND2_X4 U2112 ( .A1(n1840), .A2(n1846), .ZN(net89076) );
  INV_X4 U2113 ( .A(n1845), .ZN(n1846) );
  OAI211_X2 U2114 ( .C1(net86169), .C2(net84408), .A(net84409), .B(net85842), 
        .ZN(net84385) );
  INV_X16 U2115 ( .A(net86160), .ZN(net85842) );
  INV_X8 U2116 ( .A(n1597), .ZN(net86160) );
  INV_X4 U2117 ( .A(net84445), .ZN(net84408) );
  NOR2_X4 U2118 ( .A1(net84408), .A2(net84642), .ZN(net84765) );
  OAI211_X2 U2119 ( .C1(net84408), .C2(net84624), .A(net84625), .B(net84626), 
        .ZN(net84615) );
  INV_X4 U2120 ( .A(n1844), .ZN(n1843) );
  OAI211_X1 U2121 ( .C1(n1841), .C2(n1843), .A(net84421), .B(net85842), .ZN(
        net89975) );
  NOR2_X1 U2122 ( .A1(n1554), .A2(net84312), .ZN(n1844) );
  INV_X4 U2123 ( .A(net84263), .ZN(n1841) );
  NOR3_X2 U2124 ( .A1(net84312), .A2(n1841), .A3(net84314), .ZN(net84276) );
  AOI211_X4 U2125 ( .C1(net84386), .C2(net85842), .A(net84387), .B(n1762), 
        .ZN(net89917) );
  NAND2_X4 U2126 ( .A1(net88721), .A2(n1849), .ZN(net84030) );
  AOI22_X4 U2127 ( .A1(net84027), .A2(net84028), .B1(net84030), .B2(net84029), 
        .ZN(net84026) );
  INV_X4 U2128 ( .A(n1848), .ZN(n1849) );
  NAND2_X4 U2129 ( .A1(net84010), .A2(n1847), .ZN(n1848) );
  NOR2_X4 U2130 ( .A1(net83787), .A2(net85847), .ZN(n1847) );
  NAND2_X4 U2131 ( .A1(net88332), .A2(net85048), .ZN(net85186) );
  NOR3_X4 U2132 ( .A1(net86027), .A2(net85186), .A3(net85285), .ZN(net88605)
         );
  OAI211_X4 U2133 ( .C1(net85186), .C2(net85187), .A(net85143), .B(net85142), 
        .ZN(net85185) );
  INV_X4 U2134 ( .A(net90110), .ZN(net85048) );
  INV_X8 U2135 ( .A(net85161), .ZN(net88332) );
  NAND4_X4 U2136 ( .A1(net88332), .A2(net85159), .A3(net85158), .A4(net85157), 
        .ZN(net85155) );
  OR2_X4 U2137 ( .A1(net85161), .A2(net90110), .ZN(fract_denorm[10]) );
  NAND2_X2 U2138 ( .A1(net84522), .A2(n1764), .ZN(net88950) );
  NAND2_X2 U2139 ( .A1(net84564), .A2(n1850), .ZN(net84518) );
  INV_X2 U2140 ( .A(\u4/N423 ), .ZN(n1850) );
  NOR2_X4 U2141 ( .A1(net84783), .A2(net84519), .ZN(net84777) );
  NAND2_X2 U2142 ( .A1(net86037), .A2(net85854), .ZN(net84015) );
  NOR2_X4 U2143 ( .A1(net84452), .A2(net84490), .ZN(net84770) );
  NAND2_X2 U2144 ( .A1(net84448), .A2(net84764), .ZN(net84452) );
  NAND2_X1 U2145 ( .A1(n1851), .A2(\u4/fract_out_pl1[10] ), .ZN(net84473) );
  INV_X4 U2146 ( .A(net84449), .ZN(n1852) );
  AND2_X2 U2147 ( .A1(net84774), .A2(net84775), .ZN(net89595) );
  INV_X4 U2148 ( .A(net84579), .ZN(net84590) );
  NAND2_X2 U2149 ( .A1(net84448), .A2(net84449), .ZN(net83432) );
  BUF_X32 U2150 ( .A(net84113), .Z(net89716) );
  NAND2_X4 U2151 ( .A1(net84839), .A2(net84840), .ZN(\u4/fract_out[6] ) );
  INV_X8 U2152 ( .A(\u4/fract_out[3] ), .ZN(net84110) );
  INV_X4 U2153 ( .A(net84110), .ZN(net99874) );
  NAND2_X4 U2154 ( .A1(n1749), .A2(net85842), .ZN(net84390) );
  INV_X1 U2155 ( .A(n1535), .ZN(net89987) );
  OAI22_X2 U2156 ( .A1(net84402), .A2(net86016), .B1(n1751), .B2(net84402), 
        .ZN(net86015) );
  INV_X4 U2157 ( .A(net84675), .ZN(n1853) );
  NOR2_X1 U2158 ( .A1(net84480), .A2(n1853), .ZN(net84551) );
  NAND2_X2 U2159 ( .A1(net85828), .A2(n1853), .ZN(net83429) );
  OAI211_X4 U2160 ( .C1(net91015), .C2(net85018), .A(net85020), .B(net85021), 
        .ZN(net84974) );
  INV_X4 U2161 ( .A(net84913), .ZN(net84895) );
  NAND2_X2 U2162 ( .A1(net84895), .A2(net83936), .ZN(net83408) );
  NAND2_X2 U2163 ( .A1(net83951), .A2(net85847), .ZN(net84913) );
  NAND2_X4 U2164 ( .A1(net91177), .A2(net85786), .ZN(net85020) );
  AOI21_X1 U2165 ( .B1(net84822), .B2(net85786), .A(n1571), .ZN(net85018) );
  NAND2_X1 U2166 ( .A1(net84081), .A2(net86174), .ZN(net84347) );
  NAND3_X2 U2167 ( .A1(net84073), .A2(net86174), .A3(net84075), .ZN(net83868)
         );
  NAND2_X2 U2168 ( .A1(n1854), .A2(net83963), .ZN(net84075) );
  INV_X4 U2169 ( .A(net11555), .ZN(net83963) );
  INV_X4 U2170 ( .A(net84168), .ZN(n1854) );
  INV_X4 U2171 ( .A(net84333), .ZN(net84414) );
  OAI21_X2 U2172 ( .B1(net84901), .B2(net84168), .A(net84169), .ZN(net84151)
         );
  NOR2_X4 U2173 ( .A1(net85778), .A2(net84168), .ZN(net84352) );
  OAI21_X4 U2174 ( .B1(net11558), .B2(net84168), .A(net84214), .ZN(net84213)
         );
  NOR2_X4 U2175 ( .A1(net84332), .A2(net84333), .ZN(net84095) );
  NOR2_X4 U2176 ( .A1(net85744), .A2(net85998), .ZN(net85342) );
  INV_X32 U2177 ( .A(net85738), .ZN(net85998) );
  NAND2_X2 U2178 ( .A1(n1855), .A2(n1856), .ZN(net84029) );
  NAND2_X2 U2179 ( .A1(net84033), .A2(n1857), .ZN(n1856) );
  XNOR2_X2 U2180 ( .A(n1858), .B(n1644), .ZN(n1857) );
  INV_X4 U2181 ( .A(net83925), .ZN(n1859) );
  INV_X4 U2182 ( .A(net84044), .ZN(net84033) );
  MUX2_X2 U2183 ( .A(n1862), .B(net84047), .S(sign_mul_r), .Z(n1860) );
  NAND2_X2 U2184 ( .A1(net84047), .A2(net84021), .ZN(n1862) );
  NAND2_X2 U2185 ( .A1(net83779), .A2(opas_r2), .ZN(n1863) );
  OAI211_X4 U2186 ( .C1(net85182), .C2(n1866), .A(net85184), .B(net85185), 
        .ZN(net85083) );
  NOR3_X4 U2187 ( .A1(net85197), .A2(net85199), .A3(n1867), .ZN(net85142) );
  INV_X8 U2188 ( .A(n1864), .ZN(n1867) );
  NOR3_X4 U2189 ( .A1(net85197), .A2(net85199), .A3(n1867), .ZN(n1868) );
  NOR3_X4 U2190 ( .A1(net85234), .A2(n1867), .A3(net88699), .ZN(net85232) );
  INV_X2 U2191 ( .A(n1867), .ZN(net88440) );
  NAND3_X4 U2192 ( .A1(net85369), .A2(quo[13]), .A3(net85674), .ZN(n1864) );
  INV_X4 U2193 ( .A(net85051), .ZN(net85199) );
  INV_X2 U2194 ( .A(net85199), .ZN(net88421) );
  INV_X8 U2195 ( .A(net85193), .ZN(net85143) );
  NAND3_X2 U2196 ( .A1(net85188), .A2(net85143), .A3(n1868), .ZN(n1866) );
  NAND2_X2 U2197 ( .A1(n1868), .A2(net85143), .ZN(net84549) );
  NAND3_X4 U2198 ( .A1(n1865), .A2(net85195), .A3(net85194), .ZN(net85193) );
  INV_X8 U2199 ( .A(n1865), .ZN(net90215) );
  NAND2_X1 U2200 ( .A1(n1865), .A2(net85059), .ZN(net76672) );
  BUF_X32 U2201 ( .A(net84110), .Z(net89485) );
  OAI21_X4 U2202 ( .B1(net84778), .B2(n1870), .A(n1871), .ZN(\u4/fract_out[3] ) );
  NAND2_X4 U2203 ( .A1(\u4/N427 ), .A2(net84522), .ZN(n1871) );
  INV_X4 U2204 ( .A(\u4/N403 ), .ZN(n1870) );
  NAND2_X4 U2205 ( .A1(net84844), .A2(net89250), .ZN(\u4/fract_out[8] ) );
  NAND2_X4 U2206 ( .A1(\u4/N432 ), .A2(net84522), .ZN(net84844) );
  INV_X4 U2207 ( .A(\u4/N409 ), .ZN(net84845) );
  NAND2_X4 U2208 ( .A1(n1869), .A2(net84810), .ZN(net84456) );
  INV_X1 U2209 ( .A(net84456), .ZN(net84322) );
  NAND2_X2 U2210 ( .A1(net84839), .A2(net84840), .ZN(net91512) );
  NAND2_X2 U2211 ( .A1(net84844), .A2(net89250), .ZN(net90252) );
  NAND2_X4 U2212 ( .A1(net84882), .A2(n1872), .ZN(net84778) );
  INV_X4 U2213 ( .A(\u4/N386 ), .ZN(n1872) );
  INV_X4 U2214 ( .A(net84853), .ZN(net84882) );
  NAND2_X4 U2215 ( .A1(n1873), .A2(net83959), .ZN(net91015) );
  OAI21_X4 U2216 ( .B1(n1745), .B2(net85027), .A(net90207), .ZN(net84975) );
  AND2_X2 U2217 ( .A1(net86038), .A2(n1593), .ZN(n1873) );
  NAND3_X2 U2218 ( .A1(net84394), .A2(n1874), .A3(n1875), .ZN(net84386) );
  AOI22_X1 U2219 ( .A1(rmode_r3[1]), .A2(net91353), .B1(net84343), .B2(
        net84398), .ZN(n1875) );
  INV_X4 U2220 ( .A(net84326), .ZN(net84343) );
  NAND2_X2 U2221 ( .A1(net84133), .A2(net84134), .ZN(n1874) );
  NOR3_X4 U2222 ( .A1(net84135), .A2(net84148), .A3(net84393), .ZN(net84387)
         );
  INV_X4 U2223 ( .A(n1597), .ZN(net84393) );
  INV_X4 U2224 ( .A(net83870), .ZN(net83869) );
  NOR2_X4 U2225 ( .A1(n1876), .A2(net84213), .ZN(net84071) );
  NAND4_X2 U2226 ( .A1(net84215), .A2(net84216), .A3(n1877), .A4(net84218), 
        .ZN(n1876) );
  INV_X4 U2227 ( .A(net84080), .ZN(net83878) );
  NAND3_X4 U2228 ( .A1(n1879), .A2(n1878), .A3(net85216), .ZN(net76872) );
  INV_X4 U2229 ( .A(net86060), .ZN(net85317) );
  MUX2_X2 U2230 ( .A(net11485), .B(net86061), .S(net85974), .Z(net86060) );
  NAND3_X4 U2231 ( .A1(n1878), .A2(net85216), .A3(n1879), .ZN(net85178) );
  NAND2_X4 U2232 ( .A1(net85320), .A2(n1881), .ZN(n1880) );
  NAND2_X4 U2233 ( .A1(fract_out_q[14]), .A2(net83780), .ZN(n1881) );
  INV_X8 U2234 ( .A(net85083), .ZN(net89546) );
  NOR2_X2 U2235 ( .A1(net85140), .A2(net85141), .ZN(net85184) );
  NOR2_X4 U2236 ( .A1(net85190), .A2(net85189), .ZN(net85188) );
  NAND3_X2 U2237 ( .A1(net85191), .A2(net86106), .A3(net85192), .ZN(net85190)
         );
  INV_X8 U2238 ( .A(net85150), .ZN(net85192) );
  INV_X4 U2239 ( .A(net99862), .ZN(net85079) );
  OAI21_X4 U2240 ( .B1(net89546), .B2(net88618), .A(net84758), .ZN(net99862)
         );
  OAI21_X2 U2241 ( .B1(net90047), .B2(net84867), .A(net85847), .ZN(n1885) );
  NOR2_X1 U2242 ( .A1(n2151), .A2(net110929), .ZN(n2152) );
  INV_X2 U2243 ( .A(n2632), .ZN(n2633) );
  NOR2_X2 U2244 ( .A1(net83933), .A2(n2632), .ZN(n2582) );
  INV_X4 U2245 ( .A(net77073), .ZN(n1882) );
  INV_X4 U2246 ( .A(n1882), .ZN(n1883) );
  INV_X2 U2247 ( .A(net85115), .ZN(net85112) );
  INV_X4 U2248 ( .A(net88877), .ZN(net110951) );
  INV_X1 U2249 ( .A(net85080), .ZN(net90026) );
  INV_X4 U2250 ( .A(net110929), .ZN(net91467) );
  NAND2_X4 U2251 ( .A1(net88636), .A2(net85089), .ZN(net85085) );
  NAND3_X4 U2252 ( .A1(net85085), .A2(net85215), .A3(net85087), .ZN(net84503)
         );
  AND3_X4 U2253 ( .A1(n1755), .A2(net88551), .A3(net85087), .ZN(net89965) );
  INV_X4 U2254 ( .A(net85089), .ZN(net91109) );
  NAND3_X2 U2255 ( .A1(net85089), .A2(net89935), .A3(net88605), .ZN(net85214)
         );
  OAI21_X4 U2256 ( .B1(n1884), .B2(fract_denorm[9]), .A(net89300), .ZN(
        net85097) );
  INV_X4 U2257 ( .A(net76926), .ZN(n1884) );
  INV_X4 U2258 ( .A(n1884), .ZN(net90037) );
  NAND2_X4 U2259 ( .A1(net85159), .A2(net85158), .ZN(fract_denorm[9]) );
  INV_X8 U2260 ( .A(fract_denorm[9]), .ZN(net90210) );
  INV_X4 U2261 ( .A(net85357), .ZN(net85158) );
  NAND2_X4 U2262 ( .A1(net85260), .A2(net85261), .ZN(net85360) );
  AND3_X4 U2263 ( .A1(net91059), .A2(net90019), .A3(net85248), .ZN(net89300)
         );
  OAI211_X4 U2264 ( .C1(net85137), .C2(net85240), .A(net89300), .B(net85177), 
        .ZN(net85239) );
  NAND2_X4 U2265 ( .A1(net89753), .A2(net84600), .ZN(net84960) );
  NAND2_X2 U2266 ( .A1(n1885), .A2(net85778), .ZN(net84969) );
  NAND2_X4 U2267 ( .A1(net88605), .A2(net89935), .ZN(net86026) );
  OAI211_X4 U2268 ( .C1(net86026), .C2(net91109), .A(net88551), .B(net85087), 
        .ZN(net85081) );
  NAND2_X4 U2269 ( .A1(net85283), .A2(net85240), .ZN(net86027) );
  NAND4_X2 U2270 ( .A1(net85168), .A2(net85171), .A3(net85169), .A4(net85170), 
        .ZN(net85290) );
  NOR3_X4 U2271 ( .A1(n1887), .A2(net90215), .A3(net85060), .ZN(net85283) );
  NAND4_X4 U2272 ( .A1(net85068), .A2(n1886), .A3(net85067), .A4(net85069), 
        .ZN(n1887) );
  NOR2_X4 U2273 ( .A1(n1888), .A2(net85310), .ZN(n1886) );
  INV_X4 U2274 ( .A(n1889), .ZN(n1888) );
  NOR2_X4 U2275 ( .A1(n1888), .A2(net85310), .ZN(net90144) );
  NAND3_X2 U2276 ( .A1(net85736), .A2(net85744), .A3(prod[14]), .ZN(n1889) );
  OAI221_X4 U2277 ( .B1(net85250), .B2(net85251), .C1(net85252), .C2(net85253), 
        .A(net85254), .ZN(net89935) );
  NOR2_X4 U2278 ( .A1(n1890), .A2(n1891), .ZN(net85260) );
  INV_X2 U2279 ( .A(net90064), .ZN(n1893) );
  INV_X4 U2280 ( .A(n1892), .ZN(n1890) );
  NAND3_X2 U2281 ( .A1(net85998), .A2(net85716), .A3(fract_out_q[2]), .ZN(
        n1892) );
  INV_X32 U2282 ( .A(net85722), .ZN(net85716) );
  XNOR2_X2 U2283 ( .A(net84503), .B(net84762), .ZN(net84609) );
  NAND2_X4 U2284 ( .A1(net84503), .A2(div_opa_ldz_r2[0]), .ZN(net84755) );
  INV_X8 U2285 ( .A(net84503), .ZN(net85080) );
  NAND3_X4 U2286 ( .A1(net84503), .A2(net89412), .A3(net89447), .ZN(net84684)
         );
  NAND2_X4 U2287 ( .A1(net85099), .A2(net85098), .ZN(net85215) );
  NAND3_X2 U2288 ( .A1(net85215), .A2(net85214), .A3(net85087), .ZN(net85213)
         );
  INV_X8 U2289 ( .A(net85239), .ZN(net85098) );
  NAND2_X4 U2290 ( .A1(net85098), .A2(net85099), .ZN(net88551) );
  INV_X8 U2291 ( .A(net85285), .ZN(net85177) );
  NAND2_X4 U2292 ( .A1(net85177), .A2(net89943), .ZN(net85176) );
  AOI21_X4 U2293 ( .B1(net77045), .B2(net86262), .A(net85178), .ZN(net85087)
         );
  INV_X2 U2294 ( .A(net91177), .ZN(net90207) );
  NAND2_X2 U2295 ( .A1(net84468), .A2(net84673), .ZN(net84984) );
  INV_X4 U2296 ( .A(net83951), .ZN(net84673) );
  NAND3_X1 U2297 ( .A1(net85786), .A2(net84915), .A3(net84673), .ZN(net84887)
         );
  INV_X4 U2298 ( .A(net84279), .ZN(net85033) );
  NAND3_X4 U2299 ( .A1(net84278), .A2(net84279), .A3(net84280), .ZN(net84277)
         );
  INV_X16 U2300 ( .A(net86037), .ZN(net86038) );
  NOR2_X4 U2301 ( .A1(net85187), .A2(net85189), .ZN(net85254) );
  NOR2_X4 U2302 ( .A1(net85744), .A2(net85728), .ZN(n1894) );
  INV_X16 U2303 ( .A(net85738), .ZN(net85728) );
  NAND2_X4 U2304 ( .A1(net85265), .A2(net85264), .ZN(net85253) );
  INV_X4 U2305 ( .A(net85251), .ZN(net85264) );
  INV_X2 U2306 ( .A(net85163), .ZN(net85265) );
  AOI21_X4 U2307 ( .B1(net85270), .B2(net90080), .A(net85272), .ZN(net85252)
         );
  INV_X8 U2308 ( .A(net85212), .ZN(n1896) );
  CLKBUF_X3 U2309 ( .A(n1896), .Z(net89266) );
  NOR2_X4 U2310 ( .A1(net85039), .A2(net86112), .ZN(net85270) );
  INV_X4 U2311 ( .A(net90292), .ZN(net85250) );
  NAND3_X2 U2312 ( .A1(net85205), .A2(net85280), .A3(net85281), .ZN(net85251)
         );
  NAND3_X4 U2313 ( .A1(n1895), .A2(net85046), .A3(net85045), .ZN(net85189) );
  INV_X8 U2314 ( .A(n1897), .ZN(n1895) );
  NAND3_X2 U2315 ( .A1(n1895), .A2(net85045), .A3(net85046), .ZN(net77073) );
  OAI21_X4 U2316 ( .B1(n1604), .B2(net90031), .A(net85257), .ZN(n1897) );
  OAI21_X4 U2317 ( .B1(n1604), .B2(net90031), .A(net85257), .ZN(net99868) );
  NAND2_X4 U2318 ( .A1(net89856), .A2(net85041), .ZN(net85163) );
  NOR3_X4 U2319 ( .A1(net85163), .A2(net90072), .A3(net85165), .ZN(net84909)
         );
  NAND2_X4 U2320 ( .A1(n1898), .A2(net85210), .ZN(net85272) );
  AOI211_X4 U2321 ( .C1(net85207), .C2(net85206), .A(net89314), .B(net85272), 
        .ZN(net85200) );
  INV_X1 U2322 ( .A(net85272), .ZN(net85162) );
  NOR2_X4 U2323 ( .A1(net85335), .A2(net85336), .ZN(n1898) );
  NAND2_X4 U2324 ( .A1(n2088), .A2(net84990), .ZN(n2093) );
  AOI22_X4 U2325 ( .A1(net85015), .A2(net84992), .B1(net89753), .B2(n1592), 
        .ZN(n2088) );
  INV_X4 U2326 ( .A(net85213), .ZN(net85116) );
  NAND2_X4 U2327 ( .A1(\fract_i2f[7] ), .A2(net85720), .ZN(net85257) );
  INV_X2 U2328 ( .A(net88695), .ZN(net91548) );
  NOR3_X2 U2329 ( .A1(\u4/N414 ), .A2(\u4/N413 ), .A3(\u4/N412 ), .ZN(n2167)
         );
  NAND2_X2 U2330 ( .A1(net91159), .A2(net84870), .ZN(n2097) );
  NAND2_X2 U2331 ( .A1(n1947), .A2(net85131), .ZN(n2055) );
  NOR2_X4 U2332 ( .A1(n1901), .A2(n1556), .ZN(net89856) );
  INV_X8 U2333 ( .A(n1903), .ZN(n1901) );
  NOR2_X4 U2334 ( .A1(n1901), .A2(n1902), .ZN(net85040) );
  NAND3_X4 U2335 ( .A1(net85736), .A2(net85744), .A3(n1904), .ZN(n1903) );
  INV_X4 U2336 ( .A(net88972), .ZN(n1904) );
  NOR2_X4 U2337 ( .A1(net11576), .A2(net85718), .ZN(n1902) );
  INV_X4 U2338 ( .A(net84643), .ZN(net84448) );
  XNOR2_X2 U2339 ( .A(net88896), .B(net84511), .ZN(net88895) );
  BUF_X32 U2340 ( .A(net88895), .Z(net89679) );
  NAND3_X2 U2341 ( .A1(net84910), .A2(net85162), .A3(net84909), .ZN(net85147)
         );
  INV_X4 U2342 ( .A(net85042), .ZN(net85165) );
  INV_X1 U2343 ( .A(net85165), .ZN(net90074) );
  NAND2_X2 U2344 ( .A1(net85393), .A2(net86096), .ZN(net90072) );
  INV_X1 U2345 ( .A(net90072), .ZN(net88585) );
  NAND3_X4 U2346 ( .A1(net85361), .A2(quo[7]), .A3(net85674), .ZN(net85042) );
  NAND2_X4 U2347 ( .A1(net85043), .A2(net85042), .ZN(net90292) );
  NAND2_X4 U2348 ( .A1(net85040), .A2(net85041), .ZN(net89314) );
  NAND2_X4 U2349 ( .A1(net85393), .A2(net86096), .ZN(net85164) );
  NAND3_X2 U2350 ( .A1(net85361), .A2(quo[8]), .A3(net85684), .ZN(net85168) );
  XNOR2_X2 U2351 ( .A(n1761), .B(net84753), .ZN(net83420) );
  INV_X4 U2352 ( .A(net83420), .ZN(net88503) );
  XNOR2_X2 U2353 ( .A(n1761), .B(n1557), .ZN(net90299) );
  NAND3_X2 U2354 ( .A1(net89412), .A2(div_opa_ldz_r2[1]), .A3(net89447), .ZN(
        n1905) );
  INV_X2 U2355 ( .A(net84758), .ZN(net89446) );
  NAND2_X4 U2356 ( .A1(net91467), .A2(net84982), .ZN(net84994) );
  NAND2_X4 U2357 ( .A1(net91467), .A2(net83933), .ZN(net84995) );
  NOR2_X1 U2358 ( .A1(net85854), .A2(n1907), .ZN(net90997) );
  INV_X4 U2359 ( .A(n1906), .ZN(n1907) );
  NAND2_X2 U2360 ( .A1(n1571), .A2(n1596), .ZN(net83844) );
  NAND4_X4 U2361 ( .A1(net85135), .A2(net85147), .A3(net85126), .A4(net85125), 
        .ZN(net85120) );
  INV_X8 U2362 ( .A(net85337), .ZN(net85335) );
  NAND3_X4 U2363 ( .A1(net85736), .A2(net85746), .A3(n1908), .ZN(net85337) );
  INV_X4 U2364 ( .A(net89543), .ZN(n1908) );
  NAND2_X4 U2365 ( .A1(net85203), .A2(net85205), .ZN(net77637) );
  NAND2_X4 U2366 ( .A1(net85032), .A2(n1551), .ZN(net90126) );
  NAND2_X2 U2367 ( .A1(n1551), .A2(net85032), .ZN(net85093) );
  NAND2_X4 U2368 ( .A1(net85032), .A2(n1551), .ZN(net84299) );
  INV_X4 U2369 ( .A(net85133), .ZN(net85107) );
  NAND3_X2 U2370 ( .A1(net85104), .A2(net85105), .A3(net85107), .ZN(net85095)
         );
  INV_X8 U2371 ( .A(net85120), .ZN(net85144) );
  INV_X8 U2372 ( .A(net85155), .ZN(net85125) );
  INV_X1 U2373 ( .A(net85125), .ZN(net89862) );
  INV_X4 U2374 ( .A(net85160), .ZN(net85157) );
  INV_X8 U2375 ( .A(net85166), .ZN(net85135) );
  OAI211_X4 U2376 ( .C1(net84549), .C2(net85124), .A(net85135), .B(net85136), 
        .ZN(net85105) );
  NAND2_X4 U2377 ( .A1(n1909), .A2(n1910), .ZN(net85166) );
  NAND4_X2 U2378 ( .A1(net85168), .A2(net85171), .A3(net85170), .A4(net85169), 
        .ZN(n1911) );
  NAND2_X4 U2379 ( .A1(net85224), .A2(n1913), .ZN(n1912) );
  INV_X8 U2380 ( .A(n1914), .ZN(n1913) );
  NAND2_X4 U2381 ( .A1(net85224), .A2(n1913), .ZN(net76645) );
  NOR2_X4 U2382 ( .A1(net83407), .A2(net83408), .ZN(net83406) );
  INV_X8 U2383 ( .A(net76048), .ZN(net85207) );
  INV_X8 U2384 ( .A(net84301), .ZN(net91159) );
  INV_X1 U2385 ( .A(net85144), .ZN(net89677) );
  AOI211_X4 U2386 ( .C1(net88950), .C2(n1610), .A(net84322), .B(n1916), .ZN(
        n1915) );
  OR2_X2 U2387 ( .A1(net83927), .A2(net84458), .ZN(n1916) );
  NAND3_X2 U2388 ( .A1(net84199), .A2(net89975), .A3(net84200), .ZN(net83863)
         );
  AOI21_X2 U2389 ( .B1(n2346), .B2(n2345), .A(n2344), .ZN(n2347) );
  OR2_X4 U2390 ( .A1(n2099), .A2(net88293), .ZN(n1917) );
  INV_X4 U2391 ( .A(n1571), .ZN(net88293) );
  NOR2_X1 U2392 ( .A1(net11560), .A2(net84856), .ZN(n2078) );
  NOR2_X2 U2393 ( .A1(net84901), .A2(net84856), .ZN(n2091) );
  NOR2_X2 U2394 ( .A1(n1662), .A2(n2567), .ZN(n2568) );
  NAND3_X2 U2395 ( .A1(net83849), .A2(n2554), .A3(n2553), .ZN(n2556) );
  NAND2_X4 U2396 ( .A1(net83861), .A2(net84220), .ZN(n2623) );
  NAND3_X2 U2397 ( .A1(n2436), .A2(n2435), .A3(n2623), .ZN(n2373) );
  OAI21_X4 U2398 ( .B1(n2501), .B2(n2500), .A(n2499), .ZN(n2523) );
  NAND3_X1 U2399 ( .A1(net85342), .A2(quo[0]), .A3(net85684), .ZN(net86106) );
  INV_X16 U2400 ( .A(net86262), .ZN(net86263) );
  NAND2_X2 U2401 ( .A1(n1900), .A2(net85116), .ZN(n1948) );
  NAND3_X2 U2402 ( .A1(quo[10]), .A2(net85752), .A3(net85738), .ZN(n1918) );
  NOR2_X4 U2403 ( .A1(net85744), .A2(net85728), .ZN(n1942) );
  NAND2_X1 U2404 ( .A1(net89266), .A2(net85071), .ZN(n3000) );
  NOR2_X2 U2405 ( .A1(net77815), .A2(net83402), .ZN(net84663) );
  NOR2_X4 U2406 ( .A1(net85730), .A2(net88695), .ZN(n2005) );
  NAND2_X4 U2407 ( .A1(n1754), .A2(n2170), .ZN(n3006) );
  NAND2_X4 U2408 ( .A1(net89819), .A2(net84842), .ZN(n1924) );
  NAND2_X4 U2409 ( .A1(\u4/N431 ), .A2(net84522), .ZN(net84842) );
  NOR3_X4 U2410 ( .A1(\u4/N416 ), .A2(\u4/N417 ), .A3(\u4/N415 ), .ZN(n2166)
         );
  NAND2_X4 U2411 ( .A1(n2162), .A2(n1952), .ZN(\u4/fract_out[1] ) );
  NAND2_X4 U2412 ( .A1(\u4/N429 ), .A2(net84522), .ZN(n2160) );
  INV_X2 U2413 ( .A(net84299), .ZN(net89681) );
  NAND2_X4 U2414 ( .A1(n3096), .A2(net90126), .ZN(n1950) );
  NAND4_X2 U2415 ( .A1(n2491), .A2(n2496), .A3(n1588), .A4(n2477), .ZN(n2480)
         );
  NOR2_X2 U2416 ( .A1(n2707), .A2(net83800), .ZN(n2664) );
  AND2_X2 U2417 ( .A1(net84522), .A2(net84774), .ZN(net91325) );
  NOR2_X4 U2418 ( .A1(div_opa_ldz_r2[1]), .A2(net91159), .ZN(net84754) );
  NAND2_X2 U2419 ( .A1(net85722), .A2(n1657), .ZN(net85281) );
  NOR2_X1 U2420 ( .A1(net88618), .A2(net89546), .ZN(n2056) );
  NOR2_X2 U2421 ( .A1(net85137), .A2(net76645), .ZN(n2045) );
  NAND2_X2 U2422 ( .A1(net89029), .A2(n1661), .ZN(net84652) );
  NAND4_X4 U2423 ( .A1(n2709), .A2(net88319), .A3(n2665), .A4(net83779), .ZN(
        n2666) );
  AOI21_X2 U2424 ( .B1(net84211), .B2(net84128), .A(net89987), .ZN(n2453) );
  NAND2_X4 U2425 ( .A1(net85116), .A2(n1900), .ZN(n2139) );
  NAND2_X4 U2426 ( .A1(\u4/N430 ), .A2(net84522), .ZN(net84839) );
  INV_X8 U2427 ( .A(net91128), .ZN(net83407) );
  CLKBUF_X3 U2428 ( .A(net84702), .Z(net91128) );
  NOR2_X4 U2429 ( .A1(net99868), .A2(n2049), .ZN(n2051) );
  NAND2_X2 U2430 ( .A1(net85720), .A2(n1658), .ZN(n2022) );
  NAND2_X1 U2431 ( .A1(net85720), .A2(n1667), .ZN(net85374) );
  AND2_X2 U2432 ( .A1(net84869), .A2(n2054), .ZN(net91112) );
  OAI21_X4 U2433 ( .B1(n2216), .B2(n2250), .A(n2215), .ZN(net84511) );
  NOR2_X4 U2434 ( .A1(net85710), .A2(net89964), .ZN(n2216) );
  AOI22_X4 U2435 ( .A1(n2018), .A2(net85684), .B1(n2017), .B2(fract_out_q[10]), 
        .ZN(n2038) );
  NAND4_X4 U2436 ( .A1(n2051), .A2(n1970), .A3(net85045), .A4(net85046), .ZN(
        n2052) );
  NAND2_X1 U2437 ( .A1(net85722), .A2(n1668), .ZN(n2029) );
  NAND2_X2 U2438 ( .A1(net85722), .A2(n1659), .ZN(n2069) );
  NAND2_X4 U2439 ( .A1(net89680), .A2(net89681), .ZN(n1935) );
  INV_X1 U2440 ( .A(net83407), .ZN(net91095) );
  AND4_X4 U2441 ( .A1(net85061), .A2(n2043), .A3(n2067), .A4(n2066), .ZN(n1971) );
  INV_X1 U2442 ( .A(net86263), .ZN(net84601) );
  INV_X4 U2443 ( .A(net90031), .ZN(net86125) );
  NAND2_X4 U2444 ( .A1(net85144), .A2(n2053), .ZN(net85104) );
  NOR2_X4 U2445 ( .A1(n2035), .A2(net89998), .ZN(net88287) );
  BUF_X8 U2446 ( .A(net83780), .Z(net91075) );
  INV_X4 U2447 ( .A(net77045), .ZN(net91069) );
  INV_X8 U2448 ( .A(net91069), .ZN(net91070) );
  NAND2_X4 U2449 ( .A1(net84749), .A2(n2190), .ZN(n2443) );
  NAND3_X4 U2450 ( .A1(n1930), .A2(net85123), .A3(net84531), .ZN(n2190) );
  NAND2_X4 U2451 ( .A1(net85091), .A2(net85095), .ZN(n1972) );
  NAND4_X2 U2452 ( .A1(net85192), .A2(net85191), .A3(n1969), .A4(n2050), .ZN(
        net76926) );
  NAND2_X4 U2453 ( .A1(net91056), .A2(net91057), .ZN(net77815) );
  BUF_X32 U2454 ( .A(\u4/fi_ldz_mi1[3] ), .Z(n1919) );
  INV_X4 U2455 ( .A(n2448), .ZN(\u4/fi_ldz_mi1[3] ) );
  NAND3_X1 U2456 ( .A1(n2040), .A2(quo[0]), .A3(net85684), .ZN(n1970) );
  XNOR2_X1 U2457 ( .A(net91112), .B(n2410), .ZN(n2411) );
  BUF_X32 U2458 ( .A(net84869), .Z(net91047) );
  NAND2_X2 U2459 ( .A1(net84953), .A2(n2099), .ZN(net84968) );
  NAND2_X4 U2460 ( .A1(n2162), .A2(n1952), .ZN(n1920) );
  NAND2_X4 U2461 ( .A1(net85778), .A2(net90026), .ZN(n2250) );
  NAND2_X2 U2462 ( .A1(net84600), .A2(net90026), .ZN(n2968) );
  INV_X2 U2463 ( .A(net85081), .ZN(net85096) );
  NAND2_X2 U2464 ( .A1(n2009), .A2(prod[15]), .ZN(n2008) );
  INV_X4 U2465 ( .A(net84310), .ZN(net90302) );
  NOR3_X4 U2466 ( .A1(n1937), .A2(net85748), .A3(net85998), .ZN(n2018) );
  NOR2_X4 U2467 ( .A1(net85748), .A2(net85730), .ZN(n2040) );
  INV_X8 U2468 ( .A(net90210), .ZN(net90211) );
  INV_X4 U2469 ( .A(n1918), .ZN(n1921) );
  NAND3_X2 U2470 ( .A1(net85369), .A2(quo[20]), .A3(net85674), .ZN(n2027) );
  NAND2_X2 U2471 ( .A1(n2047), .A2(net85203), .ZN(n2048) );
  NOR2_X1 U2472 ( .A1(net84672), .A2(net85004), .ZN(n2154) );
  OAI21_X1 U2473 ( .B1(n2154), .B2(net84867), .A(n2153), .ZN(n2157) );
  NOR3_X1 U2474 ( .A1(net83421), .A2(net84867), .A3(n2154), .ZN(n2084) );
  NOR2_X1 U2475 ( .A1(n2580), .A2(n2579), .ZN(n2581) );
  NAND3_X2 U2476 ( .A1(n2095), .A2(net85006), .A3(n2094), .ZN(n2096) );
  OAI21_X2 U2477 ( .B1(net91095), .B2(n2219), .A(n2218), .ZN(n2261) );
  NOR2_X4 U2478 ( .A1(net85744), .A2(net85998), .ZN(n1922) );
  NAND2_X4 U2479 ( .A1(net84609), .A2(net85832), .ZN(net84610) );
  NAND3_X2 U2480 ( .A1(net84662), .A2(net84661), .A3(net84660), .ZN(net84655)
         );
  NAND2_X4 U2481 ( .A1(net83969), .A2(net85853), .ZN(n872) );
  NAND2_X4 U2482 ( .A1(net84236), .A2(net85853), .ZN(n2991) );
  NAND3_X4 U2483 ( .A1(net85736), .A2(net85752), .A3(net85716), .ZN(net85853)
         );
  INV_X4 U2484 ( .A(net85192), .ZN(net90124) );
  INV_X1 U2485 ( .A(net85131), .ZN(net90115) );
  INV_X8 U2486 ( .A(net77161), .ZN(net85131) );
  INV_X8 U2487 ( .A(net11562), .ZN(net83993) );
  INV_X1 U2488 ( .A(exp_r[1]), .ZN(net84901) );
  INV_X1 U2489 ( .A(exp_r[1]), .ZN(net84167) );
  NOR2_X4 U2490 ( .A1(net85744), .A2(net85730), .ZN(n2001) );
  NOR2_X2 U2491 ( .A1(n3077), .A2(net85716), .ZN(n2003) );
  OAI21_X2 U2492 ( .B1(net88319), .B2(n2607), .A(n2606), .ZN(n2614) );
  NAND3_X2 U2493 ( .A1(net85998), .A2(net85716), .A3(fract_out_q[9]), .ZN(
        net85169) );
  NOR3_X4 U2494 ( .A1(n2052), .A2(net90124), .A3(n1921), .ZN(net85126) );
  NOR2_X4 U2495 ( .A1(net85744), .A2(net85728), .ZN(n2016) );
  NAND3_X2 U2496 ( .A1(n2098), .A2(n2097), .A3(n2096), .ZN(\u4/shift_left [1])
         );
  INV_X2 U2497 ( .A(net84684), .ZN(net89680) );
  INV_X1 U2498 ( .A(net89964), .ZN(net84310) );
  INV_X2 U2499 ( .A(net84549), .ZN(net85123) );
  NOR2_X1 U2500 ( .A1(net84548), .A2(net84549), .ZN(n2300) );
  NAND3_X1 U2501 ( .A1(net84322), .A2(net88950), .A3(n1610), .ZN(n2302) );
  NAND3_X1 U2502 ( .A1(net83946), .A2(net88950), .A3(n2574), .ZN(n2575) );
  NAND2_X4 U2503 ( .A1(net85738), .A2(net85748), .ZN(net90031) );
  NAND3_X2 U2504 ( .A1(n2034), .A2(quo[10]), .A3(net85684), .ZN(n1923) );
  INV_X2 U2505 ( .A(net89933), .ZN(net84107) );
  BUF_X4 U2506 ( .A(net76672), .Z(net90007) );
  INV_X8 U2507 ( .A(net85718), .ZN(net89998) );
  NOR2_X2 U2508 ( .A1(net85114), .A2(net85115), .ZN(net84550) );
  NAND3_X1 U2509 ( .A1(n2321), .A2(n2474), .A3(n2498), .ZN(n1925) );
  NAND3_X2 U2510 ( .A1(net89029), .A2(net84571), .A3(n1661), .ZN(net84568) );
  NAND2_X4 U2511 ( .A1(net84684), .A2(n1948), .ZN(net89964) );
  NAND3_X2 U2512 ( .A1(n2068), .A2(n2070), .A3(n2069), .ZN(net85234) );
  OAI22_X4 U2513 ( .A1(net84107), .A2(n1961), .B1(n2513), .B2(n2511), .ZN(
        n2680) );
  NOR2_X4 U2514 ( .A1(net85744), .A2(net85730), .ZN(n2024) );
  NOR2_X4 U2515 ( .A1(net85744), .A2(net85728), .ZN(net85361) );
  INV_X2 U2516 ( .A(n1924), .ZN(n2503) );
  OAI21_X2 U2517 ( .B1(n2143), .B2(net84890), .A(n2142), .ZN(n2144) );
  NOR2_X1 U2518 ( .A1(net84191), .A2(net84079), .ZN(n2472) );
  NAND2_X1 U2519 ( .A1(net89266), .A2(net85071), .ZN(n1926) );
  NAND2_X1 U2520 ( .A1(net89266), .A2(net85071), .ZN(n1927) );
  NOR3_X1 U2521 ( .A1(net84146), .A2(net84312), .A3(net86016), .ZN(n2362) );
  NAND3_X1 U2522 ( .A1(n2478), .A2(net84150), .A3(net84081), .ZN(n2479) );
  AND3_X4 U2523 ( .A1(n2036), .A2(n2038), .A3(n2037), .ZN(net89943) );
  OAI21_X4 U2524 ( .B1(n2385), .B2(n2384), .A(net84095), .ZN(n1928) );
  BUF_X32 U2525 ( .A(\u4/fi_ldz_mi1[2] ), .Z(n1929) );
  BUF_X32 U2526 ( .A(n845), .Z(net89926) );
  INV_X1 U2527 ( .A(net88503), .ZN(net89924) );
  INV_X1 U2528 ( .A(n1919), .ZN(n1931) );
  INV_X2 U2529 ( .A(net89862), .ZN(net89863) );
  NAND2_X4 U2530 ( .A1(opas_r2), .A2(net83936), .ZN(n2159) );
  NAND2_X4 U2531 ( .A1(net85194), .A2(net85195), .ZN(net85060) );
  NAND2_X4 U2532 ( .A1(net89817), .A2(\u4/N407 ), .ZN(net89819) );
  INV_X1 U2533 ( .A(net84778), .ZN(net89817) );
  INV_X1 U2534 ( .A(\u4/fract_out[1] ), .ZN(net84103) );
  NOR2_X4 U2535 ( .A1(\u4/N421 ), .A2(\u4/N422 ), .ZN(n2164) );
  INV_X4 U2536 ( .A(net84763), .ZN(net89120) );
  XNOR2_X2 U2537 ( .A(net84702), .B(n2306), .ZN(net88896) );
  NOR2_X4 U2538 ( .A1(net84151), .A2(n1639), .ZN(n2527) );
  NOR2_X1 U2539 ( .A1(n2483), .A2(n2482), .ZN(n2489) );
  OAI21_X1 U2540 ( .B1(n2487), .B2(n2486), .A(n2485), .ZN(n2488) );
  NAND3_X2 U2541 ( .A1(net84315), .A2(net84263), .A3(net84366), .ZN(n2596) );
  NAND2_X4 U2542 ( .A1(n2341), .A2(n2340), .ZN(n2521) );
  NAND2_X4 U2543 ( .A1(n2330), .A2(n2416), .ZN(n2341) );
  INV_X1 U2544 ( .A(net89753), .ZN(net89741) );
  INV_X8 U2545 ( .A(net30297), .ZN(net83296) );
  NAND2_X1 U2546 ( .A1(n2433), .A2(n2515), .ZN(n2434) );
  NOR2_X4 U2547 ( .A1(n2515), .A2(n2674), .ZN(n2516) );
  NAND2_X2 U2548 ( .A1(net84421), .A2(n2360), .ZN(n2361) );
  NAND2_X4 U2549 ( .A1(n2356), .A2(net84371), .ZN(net84149) );
  NAND2_X2 U2550 ( .A1(net84010), .A2(net88721), .ZN(n2618) );
  INV_X4 U2551 ( .A(n2706), .ZN(n2625) );
  NAND3_X2 U2552 ( .A1(net84347), .A2(n2373), .A3(n1933), .ZN(n2375) );
  INV_X4 U2553 ( .A(n1932), .ZN(n1933) );
  NAND2_X1 U2554 ( .A1(net83878), .A2(n2623), .ZN(n2372) );
  NAND2_X4 U2555 ( .A1(n2336), .A2(n2454), .ZN(n2333) );
  NOR2_X1 U2556 ( .A1(n2706), .A2(net83736), .ZN(n2663) );
  NAND2_X2 U2557 ( .A1(net84684), .A2(net90126), .ZN(n1934) );
  NAND2_X4 U2558 ( .A1(n1935), .A2(n1934), .ZN(net84702) );
  NAND2_X2 U2559 ( .A1(net84755), .A2(net84763), .ZN(n1945) );
  NOR3_X1 U2560 ( .A1(n2080), .A2(n2079), .A3(n2078), .ZN(n2086) );
  INV_X1 U2561 ( .A(net89679), .ZN(net83414) );
  INV_X1 U2562 ( .A(net90047), .ZN(net85004) );
  NOR2_X1 U2563 ( .A1(net90268), .A2(net83421), .ZN(n2188) );
  NOR2_X4 U2564 ( .A1(net85998), .A2(net85752), .ZN(n1936) );
  NAND2_X2 U2565 ( .A1(\u4/N423 ), .A2(net84522), .ZN(n2275) );
  NAND2_X4 U2566 ( .A1(n1949), .A2(net88877), .ZN(n1951) );
  OAI21_X2 U2567 ( .B1(n2468), .B2(net84297), .A(net84298), .ZN(n2444) );
  INV_X1 U2568 ( .A(n2253), .ZN(n2254) );
  INV_X2 U2569 ( .A(n2196), .ZN(n2199) );
  NAND2_X1 U2570 ( .A1(n2401), .A2(n2222), .ZN(n2223) );
  NOR2_X4 U2571 ( .A1(net85744), .A2(net85998), .ZN(net85369) );
  OAI21_X1 U2572 ( .B1(net85676), .B2(n2572), .A(n2571), .ZN(n2629) );
  NAND2_X1 U2573 ( .A1(net85676), .A2(n2309), .ZN(net84626) );
  AOI22_X1 U2574 ( .A1(net83416), .A2(n2269), .B1(net85676), .B2(n2366), .ZN(
        n2270) );
  NAND3_X1 U2575 ( .A1(net85076), .A2(net85676), .A3(quo[2]), .ZN(n2063) );
  INV_X4 U2576 ( .A(net85365), .ZN(net85224) );
  INV_X4 U2577 ( .A(net85676), .ZN(net86113) );
  AOI21_X4 U2578 ( .B1(net89078), .B2(n1940), .A(net83990), .ZN(n3008) );
  NOR2_X2 U2579 ( .A1(n3078), .A2(net85716), .ZN(n2012) );
  OAI21_X4 U2580 ( .B1(n2670), .B2(n2669), .A(n2668), .ZN(n2672) );
  NAND4_X2 U2581 ( .A1(net90144), .A2(net85067), .A3(net85068), .A4(net85069), 
        .ZN(n3002) );
  NOR2_X2 U2582 ( .A1(net85730), .A2(n1650), .ZN(net85227) );
  NAND2_X4 U2583 ( .A1(\u4/N425 ), .A2(net84522), .ZN(n2162) );
  NAND2_X1 U2584 ( .A1(n2695), .A2(n2674), .ZN(n2675) );
  NOR2_X2 U2585 ( .A1(n1768), .A2(net84329), .ZN(n2382) );
  NAND2_X1 U2586 ( .A1(net84371), .A2(net83296), .ZN(n1938) );
  NAND2_X1 U2587 ( .A1(n1648), .A2(net30297), .ZN(n1939) );
  NAND2_X2 U2588 ( .A1(n1938), .A2(n1939), .ZN(n2435) );
  AOI21_X2 U2589 ( .B1(n2675), .B2(n1546), .A(n2683), .ZN(N221) );
  NAND3_X2 U2590 ( .A1(n2425), .A2(net85842), .A3(n2365), .ZN(n2461) );
  INV_X8 U2591 ( .A(net85164), .ZN(net85043) );
  INV_X1 U2592 ( .A(net90252), .ZN(net84119) );
  NOR2_X4 U2593 ( .A1(net85998), .A2(net85752), .ZN(n2039) );
  AOI21_X1 U2594 ( .B1(net91047), .B2(net84870), .A(n2152), .ZN(net84847) );
  NOR2_X1 U2595 ( .A1(n2234), .A2(net89741), .ZN(n2080) );
  NAND2_X2 U2596 ( .A1(net91150), .A2(\u4/N408 ), .ZN(net89250) );
  NAND3_X2 U2597 ( .A1(n2087), .A2(n2086), .A3(n2085), .ZN(\u4/shift_left [2])
         );
  NAND2_X4 U2598 ( .A1(n2356), .A2(net84371), .ZN(net84421) );
  AOI21_X2 U2599 ( .B1(n2644), .B2(n2643), .A(net83827), .ZN(n2645) );
  NAND3_X2 U2600 ( .A1(n2321), .A2(n2474), .A3(n2498), .ZN(n2336) );
  NAND2_X1 U2601 ( .A1(n2667), .A2(net83787), .ZN(n1943) );
  INV_X4 U2602 ( .A(n1943), .ZN(n1944) );
  NAND2_X1 U2603 ( .A1(net91542), .A2(net84138), .ZN(n2497) );
  NAND3_X2 U2604 ( .A1(net85790), .A2(net85010), .A3(net83849), .ZN(net84856)
         );
  NAND3_X2 U2605 ( .A1(net85716), .A2(n1656), .A3(net85728), .ZN(net85045) );
  AOI21_X2 U2606 ( .B1(n2681), .B2(n1546), .A(n2683), .ZN(N224) );
  AOI21_X2 U2607 ( .B1(n2677), .B2(n1546), .A(n2683), .ZN(N222) );
  AOI21_X2 U2608 ( .B1(n2679), .B2(n1546), .A(n2683), .ZN(N223) );
  AOI21_X2 U2609 ( .B1(n2684), .B2(n1546), .A(n2683), .ZN(N225) );
  NAND4_X4 U2610 ( .A1(net85061), .A2(n2043), .A3(n2067), .A4(n2066), .ZN(
        net85141) );
  INV_X1 U2611 ( .A(net85205), .ZN(net85204) );
  NAND2_X4 U2612 ( .A1(net85037), .A2(net85038), .ZN(n2999) );
  NOR2_X4 U2613 ( .A1(net85744), .A2(net85732), .ZN(net89129) );
  NAND2_X4 U2614 ( .A1(net89120), .A2(net89121), .ZN(n1946) );
  NAND2_X4 U2615 ( .A1(n1945), .A2(n1946), .ZN(net84761) );
  INV_X4 U2616 ( .A(n2035), .ZN(n1955) );
  NAND2_X4 U2617 ( .A1(net85194), .A2(net85195), .ZN(n2041) );
  NAND2_X2 U2618 ( .A1(n2621), .A2(n2620), .ZN(n3007) );
  NOR2_X2 U2619 ( .A1(n2616), .A2(n2617), .ZN(n2621) );
  NAND2_X4 U2620 ( .A1(net84421), .A2(net83296), .ZN(n2491) );
  OAI22_X4 U2621 ( .A1(n2186), .A2(net84777), .B1(net84778), .B2(n2185), .ZN(
        net84775) );
  AND3_X4 U2622 ( .A1(n2036), .A2(n2037), .A3(n2038), .ZN(n1947) );
  INV_X8 U2623 ( .A(n1947), .ZN(n3003) );
  OAI21_X2 U2624 ( .B1(n2233), .B2(n2968), .A(n2232), .ZN(n2965) );
  OAI21_X1 U2625 ( .B1(net85832), .B2(net90122), .A(net84610), .ZN(n2269) );
  OAI21_X2 U2626 ( .B1(n2422), .B2(net84502), .A(n2421), .ZN(net84469) );
  NAND4_X2 U2627 ( .A1(net85171), .A2(net85168), .A3(net85169), .A4(net85170), 
        .ZN(net76254) );
  NAND2_X2 U2628 ( .A1(net90299), .A2(net83421), .ZN(n1958) );
  INV_X4 U2629 ( .A(n3096), .ZN(n1949) );
  NAND2_X4 U2630 ( .A1(net90074), .A2(net88585), .ZN(n2998) );
  NAND4_X4 U2631 ( .A1(n2519), .A2(n2518), .A3(n2517), .A4(n2516), .ZN(
        net83787) );
  NAND2_X4 U2632 ( .A1(n1899), .A2(n2170), .ZN(net84814) );
  OR2_X4 U2633 ( .A1(net84778), .A2(n2163), .ZN(n1952) );
  NAND3_X2 U2634 ( .A1(n2040), .A2(quo[10]), .A3(net85684), .ZN(n2025) );
  NAND2_X4 U2635 ( .A1(n2462), .A2(n2363), .ZN(net84168) );
  INV_X8 U2636 ( .A(net85051), .ZN(net88699) );
  NOR3_X1 U2637 ( .A1(prod[0]), .A2(prod[10]), .A3(prod[1]), .ZN(n2648) );
  INV_X1 U2638 ( .A(n1528), .ZN(net84115) );
  NAND2_X4 U2639 ( .A1(net88503), .A2(\u4/exp_in_pl1[2] ), .ZN(n1959) );
  NAND2_X1 U2640 ( .A1(net84983), .A2(net84822), .ZN(n2579) );
  INV_X16 U2641 ( .A(net84858), .ZN(\u4/f2i_shft[3] ) );
  NAND2_X4 U2642 ( .A1(n2029), .A2(n2030), .ZN(net85039) );
  NAND2_X4 U2643 ( .A1(n1956), .A2(net88566), .ZN(n1957) );
  NAND2_X4 U2644 ( .A1(n1957), .A2(n2045), .ZN(net85099) );
  INV_X4 U2645 ( .A(n2046), .ZN(n1956) );
  NOR2_X4 U2646 ( .A1(n2044), .A2(net85141), .ZN(n2046) );
  OAI21_X1 U2647 ( .B1(n2192), .B2(net110951), .A(n2191), .ZN(n2196) );
  NAND2_X4 U2648 ( .A1(n1959), .A2(n1958), .ZN(net83419) );
  XNOR2_X1 U2649 ( .A(net84167), .B(net90302), .ZN(n2481) );
  NAND2_X1 U2650 ( .A1(net90302), .A2(net84167), .ZN(n2393) );
  NAND2_X1 U2651 ( .A1(net84511), .A2(n2217), .ZN(n2218) );
  NOR2_X1 U2652 ( .A1(net84511), .A2(n2217), .ZN(n2219) );
  NOR2_X1 U2653 ( .A1(n1592), .A2(net89964), .ZN(n2233) );
  NAND2_X1 U2654 ( .A1(n1592), .A2(net89964), .ZN(n2232) );
  XNOR2_X1 U2655 ( .A(net89964), .B(net85710), .ZN(n2251) );
  INV_X1 U2656 ( .A(net85207), .ZN(net88545) );
  NAND2_X4 U2657 ( .A1(net83993), .A2(net83967), .ZN(net85313) );
  NOR2_X2 U2658 ( .A1(net85211), .A2(net85212), .ZN(net85206) );
  INV_X1 U2659 ( .A(net91159), .ZN(net88510) );
  INV_X1 U2660 ( .A(net89948), .ZN(net84191) );
  NOR2_X4 U2661 ( .A1(net85738), .A2(net85722), .ZN(n2017) );
  AOI21_X2 U2662 ( .B1(n2398), .B2(n2449), .A(n2397), .ZN(n2399) );
  NAND2_X4 U2663 ( .A1(n2005), .A2(prod[2]), .ZN(n2030) );
  NOR3_X1 U2664 ( .A1(prod[14]), .A2(prod[15]), .A3(prod[16]), .ZN(n2649) );
  NOR2_X1 U2665 ( .A1(n3001), .A2(net88545), .ZN(net84911) );
  NAND3_X2 U2666 ( .A1(n2006), .A2(n2007), .A3(n2008), .ZN(net85365) );
  NAND2_X1 U2667 ( .A1(n1919), .A2(net84305), .ZN(n2398) );
  NOR2_X1 U2668 ( .A1(n1919), .A2(net84305), .ZN(n2397) );
  NOR2_X1 U2669 ( .A1(net84601), .A2(net84602), .ZN(n2273) );
  NOR2_X1 U2670 ( .A1(net83414), .A2(n2307), .ZN(n2308) );
  NAND2_X4 U2671 ( .A1(n2061), .A2(n2405), .ZN(\u4/f2i_shft[4] ) );
  NAND3_X2 U2672 ( .A1(n2075), .A2(net84290), .A3(net84305), .ZN(n2226) );
  NAND2_X4 U2673 ( .A1(net11566), .A2(net83933), .ZN(net84236) );
  NOR2_X2 U2674 ( .A1(net85730), .A2(net85752), .ZN(n2009) );
  AND2_X2 U2675 ( .A1(exp_r[2]), .A2(net83993), .ZN(\u4/add_407/carry [3]) );
  AOI22_X1 U2676 ( .A1(n2393), .A2(net84166), .B1(net84310), .B2(net83993), 
        .ZN(n2465) );
  XOR2_X1 U2677 ( .A(exp_r[2]), .B(net83993), .Z(n2119) );
  NOR2_X1 U2678 ( .A1(div_opa_ldz_r2[1]), .A2(net83993), .ZN(n2121) );
  NAND2_X1 U2679 ( .A1(net83993), .A2(div_opa_ldz_r2[1]), .ZN(n2120) );
  NAND2_X1 U2680 ( .A1(net83993), .A2(net11671), .ZN(n2102) );
  XNOR2_X1 U2681 ( .A(div_opa_ldz_r2[1]), .B(net83993), .ZN(n2133) );
  NAND2_X1 U2682 ( .A1(net85030), .A2(net11560), .ZN(n2225) );
  NAND3_X4 U2683 ( .A1(n2074), .A2(net88440), .A3(net88421), .ZN(n3005) );
  OAI211_X1 U2684 ( .C1(net83987), .C2(n2551), .A(n2550), .B(net83990), .ZN(
        n2557) );
  OAI21_X1 U2685 ( .B1(n2364), .B2(n2443), .A(net83990), .ZN(n2566) );
  NAND2_X1 U2686 ( .A1(n2223), .A2(net83990), .ZN(n2242) );
  NAND3_X2 U2687 ( .A1(net85736), .A2(net85746), .A3(prod[1]), .ZN(n2032) );
  NAND3_X2 U2688 ( .A1(net85744), .A2(net85736), .A3(prod[18]), .ZN(n2011) );
  NAND3_X2 U2689 ( .A1(net85746), .A2(net85736), .A3(prod[13]), .ZN(n2042) );
  NAND3_X2 U2690 ( .A1(net85998), .A2(net85716), .A3(fract_out_q[6]), .ZN(
        n2066) );
  NOR2_X2 U2691 ( .A1(net85744), .A2(net85728), .ZN(n2033) );
  NOR2_X2 U2692 ( .A1(net91548), .A2(net85728), .ZN(n2034) );
  NOR2_X2 U2693 ( .A1(net85748), .A2(net85728), .ZN(n2014) );
  NAND3_X2 U2694 ( .A1(net85998), .A2(net85716), .A3(fract_out_q[7]), .ZN(
        net85069) );
  NAND3_X2 U2695 ( .A1(net85998), .A2(net85716), .A3(fract_out_q[11]), .ZN(
        n2026) );
  NAND2_X2 U2696 ( .A1(fract_out_q[8]), .A2(n2017), .ZN(n2007) );
  AND3_X4 U2697 ( .A1(n2426), .A2(net85794), .A3(net88500), .ZN(n2392) );
  NAND2_X1 U2698 ( .A1(net86169), .A2(net91404), .ZN(net84312) );
  OAI21_X1 U2699 ( .B1(net88500), .B2(net84887), .A(n2144), .ZN(
        \u4/shift_right [1]) );
  NAND3_X1 U2700 ( .A1(net90047), .A2(net84982), .A3(net84983), .ZN(n2094) );
  NOR2_X4 U2701 ( .A1(n2099), .A2(net88293), .ZN(net88292) );
  INV_X1 U2702 ( .A(n2068), .ZN(n2073) );
  AOI22_X1 U2703 ( .A1(n2400), .A2(net84160), .B1(net88510), .B2(net85712), 
        .ZN(n2468) );
  NAND2_X1 U2706 ( .A1(net90126), .A2(net84684), .ZN(n2222) );
  NOR2_X1 U2707 ( .A1(net110951), .A2(net84684), .ZN(n2253) );
  NOR2_X2 U2708 ( .A1(n3076), .A2(net85718), .ZN(net85310) );
  AOI21_X2 U2709 ( .B1(n2664), .B2(n2663), .A(n2669), .ZN(n2673) );
  NAND4_X4 U2710 ( .A1(n2598), .A2(net83844), .A3(net83855), .A4(net83906), 
        .ZN(n2702) );
  XNOR2_X1 U2711 ( .A(n1931), .B(net83968), .ZN(n2450) );
  NAND2_X4 U2712 ( .A1(net84869), .A2(n2054), .ZN(net83990) );
  INV_X1 U2713 ( .A(fract_denorm[10]), .ZN(net84532) );
  AOI22_X4 U2714 ( .A1(net89998), .A2(n1633), .B1(prod[19]), .B2(net86125), 
        .ZN(net85220) );
  AOI21_X1 U2715 ( .B1(net90268), .B2(net83421), .A(net89924), .ZN(n2189) );
  NOR2_X1 U2716 ( .A1(\u4/fract_out_pl1[10] ), .A2(net83429), .ZN(n2962) );
  INV_X8 U2717 ( .A(n2514), .ZN(n1960) );
  OAI21_X2 U2718 ( .B1(net83754), .B2(n2693), .A(n2692), .ZN(N229) );
  OAI21_X2 U2719 ( .B1(net83754), .B2(n2690), .A(n2692), .ZN(N228) );
  OAI21_X2 U2720 ( .B1(net83754), .B2(n2688), .A(n2692), .ZN(N227) );
  OAI21_X2 U2721 ( .B1(net83754), .B2(n2686), .A(n2692), .ZN(N226) );
  OAI21_X2 U2722 ( .B1(net83754), .B2(n2434), .A(n2692), .ZN(N220) );
  NAND2_X4 U2723 ( .A1(n2702), .A2(net85790), .ZN(n2609) );
  AOI21_X4 U2724 ( .B1(n2609), .B2(n2610), .A(n2608), .ZN(n2617) );
  NAND2_X1 U2725 ( .A1(net84421), .A2(net30297), .ZN(n2478) );
  NAND2_X1 U2726 ( .A1(net84421), .A2(net84150), .ZN(n2493) );
  NOR2_X2 U2727 ( .A1(net83853), .A2(n2628), .ZN(n2642) );
  AOI21_X2 U2728 ( .B1(n1648), .B2(n2496), .A(n2996), .ZN(n2350) );
  NAND4_X1 U2729 ( .A1(n2496), .A2(n2491), .A3(net84081), .A4(net86169), .ZN(
        n2337) );
  NAND2_X4 U2730 ( .A1(net84983), .A2(net84982), .ZN(n2081) );
  NAND3_X2 U2731 ( .A1(net85116), .A2(n2057), .A3(n2056), .ZN(n2059) );
  INV_X1 U2732 ( .A(net86169), .ZN(net84128) );
  INV_X2 U2733 ( .A(net85060), .ZN(net85059) );
  INV_X1 U2734 ( .A(n1929), .ZN(n2394) );
  NAND2_X1 U2735 ( .A1(exp_r[2]), .A2(n2394), .ZN(n2395) );
  NOR2_X1 U2736 ( .A1(exp_r[2]), .A2(n2394), .ZN(n2396) );
  INV_X8 U2737 ( .A(net85103), .ZN(net85032) );
  NAND2_X4 U2738 ( .A1(n1954), .A2(net85105), .ZN(net85103) );
  NAND2_X4 U2739 ( .A1(net85738), .A2(net85752), .ZN(net85351) );
  NAND2_X1 U2740 ( .A1(opa_00), .A2(net84015), .ZN(n2352) );
  OAI21_X2 U2741 ( .B1(n2378), .B2(n2377), .A(net84341), .ZN(n2380) );
  OAI21_X2 U2742 ( .B1(n2429), .B2(n2428), .A(opa_00), .ZN(n2431) );
  NAND2_X4 U2743 ( .A1(net85738), .A2(net85748), .ZN(n2035) );
  OAI211_X1 U2744 ( .C1(n2276), .C2(net84561), .A(net11555), .B(n1608), .ZN(
        n2277) );
  NAND3_X2 U2745 ( .A1(fract_out_q[1]), .A2(net85716), .A3(net85732), .ZN(
        n1969) );
  INV_X4 U2746 ( .A(n1969), .ZN(n2049) );
  NAND2_X4 U2747 ( .A1(n2015), .A2(prod[10]), .ZN(net85292) );
  NOR2_X4 U2748 ( .A1(n2031), .A2(net86113), .ZN(net86112) );
  NAND2_X4 U2749 ( .A1(n1921), .A2(net85676), .ZN(net85191) );
  NAND3_X2 U2750 ( .A1(n2034), .A2(quo[0]), .A3(net85684), .ZN(n2050) );
  NAND2_X4 U2751 ( .A1(n2039), .A2(prod[11]), .ZN(n2070) );
  OAI211_X4 U2752 ( .C1(n2031), .C2(net85684), .A(n2030), .B(n2029), .ZN(
        net76048) );
  NAND4_X4 U2753 ( .A1(n2028), .A2(n2027), .A3(n2026), .A4(n2025), .ZN(
        net85285) );
  NAND2_X4 U2754 ( .A1(net85280), .A2(net85281), .ZN(net85331) );
  NAND2_X4 U2755 ( .A1(n2033), .A2(quo[4]), .ZN(n2031) );
  NAND3_X1 U2756 ( .A1(net88319), .A2(n1744), .A3(net90217), .ZN(net85854) );
  NAND2_X4 U2757 ( .A1(n2015), .A2(prod[9]), .ZN(net85263) );
  NAND3_X4 U2758 ( .A1(net85076), .A2(net85674), .A3(quo[18]), .ZN(net85170)
         );
  NAND2_X4 U2759 ( .A1(n1936), .A2(prod[6]), .ZN(net85280) );
  NAND2_X4 U2760 ( .A1(n1973), .A2(net85096), .ZN(n2060) );
  INV_X4 U2761 ( .A(n1972), .ZN(n1973) );
  NAND2_X4 U2762 ( .A1(n1971), .A2(net88566), .ZN(net85124) );
  NAND2_X4 U2763 ( .A1(n2436), .A2(n2435), .ZN(net83875) );
  NAND2_X1 U2764 ( .A1(rmode_r3[1]), .A2(net84403), .ZN(net84402) );
  NAND3_X2 U2765 ( .A1(n2656), .A2(n2619), .A3(net83806), .ZN(n2620) );
  INV_X1 U2766 ( .A(net88319), .ZN(net86010) );
  NAND3_X2 U2767 ( .A1(net85744), .A2(net86006), .A3(prod[16]), .ZN(n2002) );
  XNOR2_X1 U2768 ( .A(net89681), .B(net83421), .ZN(n2467) );
  AOI22_X1 U2769 ( .A1(net85015), .A2(n1949), .B1(net89681), .B2(net84870), 
        .ZN(n2087) );
  AOI22_X4 U2770 ( .A1(net89998), .A2(n1634), .B1(n1955), .B2(prod[17]), .ZN(
        n2036) );
  NAND3_X2 U2771 ( .A1(net85736), .A2(net85746), .A3(prod[8]), .ZN(n2010) );
  NAND3_X2 U2772 ( .A1(net85746), .A2(net85736), .A3(prod[5]), .ZN(net85393)
         );
  INV_X2 U2773 ( .A(n2695), .ZN(n2696) );
  NAND2_X1 U2774 ( .A1(n2695), .A2(n2678), .ZN(n2679) );
  NAND2_X1 U2775 ( .A1(n2695), .A2(n2680), .ZN(n2681) );
  NOR2_X1 U2776 ( .A1(net86037), .A2(n1595), .ZN(n2429) );
  NOR2_X1 U2777 ( .A1(net86037), .A2(net83925), .ZN(n2587) );
  NOR2_X1 U2778 ( .A1(net86037), .A2(n2585), .ZN(n2378) );
  NOR2_X1 U2779 ( .A1(net86037), .A2(net85710), .ZN(net84996) );
  NAND4_X4 U2780 ( .A1(n2028), .A2(n2026), .A3(n2027), .A4(n1923), .ZN(
        net77161) );
  NAND3_X2 U2781 ( .A1(n2036), .A2(n2037), .A3(n2038), .ZN(net85137) );
  NAND2_X1 U2782 ( .A1(net84983), .A2(n1553), .ZN(n2082) );
  XNOR2_X1 U2783 ( .A(n1929), .B(net11560), .ZN(n2464) );
  NAND2_X1 U2784 ( .A1(n2613), .A2(net85842), .ZN(n2694) );
  NAND3_X1 U2785 ( .A1(n2597), .A2(net85842), .A3(n2613), .ZN(n2598) );
  NAND3_X1 U2786 ( .A1(n2425), .A2(net11566), .A3(net85842), .ZN(n2418) );
  XNOR2_X1 U2787 ( .A(net91159), .B(net85710), .ZN(n2484) );
  NAND2_X1 U2788 ( .A1(net91159), .A2(net85710), .ZN(n2400) );
  NOR2_X1 U2789 ( .A1(net89681), .A2(net91159), .ZN(n2364) );
  NOR2_X1 U2790 ( .A1(div_opa_ldz_r2[2]), .A2(net89537), .ZN(n2192) );
  NAND2_X1 U2791 ( .A1(div_opa_ldz_r2[2]), .A2(net89537), .ZN(n2191) );
  AOI22_X4 U2792 ( .A1(net83800), .A2(n2433), .B1(n2683), .B2(n2956), .ZN(
        n2692) );
  NAND3_X1 U2793 ( .A1(net11566), .A2(net85786), .A3(n2327), .ZN(n2543) );
  NAND2_X1 U2794 ( .A1(\u4/exp_in_pl1[5] ), .A2(net85786), .ZN(net84822) );
  NOR3_X1 U2795 ( .A1(net83849), .A2(net83959), .A3(n2566), .ZN(n2567) );
  NOR2_X1 U2796 ( .A1(net83968), .A2(net83959), .ZN(n2553) );
  NAND2_X4 U2797 ( .A1(n2081), .A2(net84468), .ZN(net83945) );
  NAND2_X4 U2798 ( .A1(n2611), .A2(n2612), .ZN(n2695) );
  NAND2_X1 U2799 ( .A1(\u4/exp_next_mi[0] ), .A2(net84157), .ZN(n2367) );
  AOI21_X1 U2800 ( .B1(net86038), .B2(n2698), .A(net85790), .ZN(n2704) );
  NAND4_X1 U2801 ( .A1(net86038), .A2(n1572), .A3(n1595), .A4(n2534), .ZN(
        n2538) );
  NAND2_X4 U2802 ( .A1(net83871), .A2(n2623), .ZN(n2709) );
  NAND2_X1 U2803 ( .A1(net83779), .A2(net86038), .ZN(net84044) );
  NAND4_X1 U2804 ( .A1(n2584), .A2(net83927), .A3(n2583), .A4(net86038), .ZN(
        n2639) );
  NAND3_X1 U2805 ( .A1(n1574), .A2(net86038), .A3(n1615), .ZN(n2605) );
  NAND2_X1 U2806 ( .A1(net86038), .A2(n2579), .ZN(n2187) );
  NAND2_X1 U2807 ( .A1(net86038), .A2(n1571), .ZN(net84675) );
  NAND2_X4 U2808 ( .A1(net88287), .A2(prod[21]), .ZN(net85216) );
  NAND2_X1 U2809 ( .A1(\u4/fract_out_pl1[10] ), .A2(rmode_r3[1]), .ZN(net84480) );
  NAND3_X1 U2810 ( .A1(n1917), .A2(n2082), .A3(net86038), .ZN(n2153) );
  NAND2_X4 U2811 ( .A1(net84096), .A2(net84095), .ZN(net83765) );
  INV_X32 U2812 ( .A(n1980), .ZN(n1978) );
  INV_X4 U2813 ( .A(opb_r[11]), .ZN(n3016) );
  INV_X4 U2814 ( .A(n3112), .ZN(n3014) );
  INV_X4 U2815 ( .A(n3111), .ZN(n3015) );
  NAND4_X2 U2816 ( .A1(n3103), .A2(n3104), .A3(n3101), .A4(n3102), .ZN(n1990)
         );
  INV_X4 U2817 ( .A(n3105), .ZN(n2895) );
  NAND4_X2 U2818 ( .A1(n3109), .A2(n3107), .A3(n3108), .A4(n3106), .ZN(n1989)
         );
  NAND2_X2 U2819 ( .A1(n2959), .A2(n3110), .ZN(n3130) );
  INV_X4 U2820 ( .A(n3114), .ZN(n2889) );
  INV_X4 U2821 ( .A(n3115), .ZN(n2896) );
  NAND2_X2 U2822 ( .A1(n3113), .A2(n3112), .ZN(n1992) );
  NAND2_X2 U2823 ( .A1(n3117), .A2(n3116), .ZN(n1991) );
  NAND2_X2 U2824 ( .A1(n3119), .A2(n3118), .ZN(n1994) );
  INV_X4 U2825 ( .A(n1996), .ZN(N56) );
  INV_X4 U2826 ( .A(N77), .ZN(n2000) );
  NAND2_X2 U2827 ( .A1(n2000), .A2(n3012), .ZN(\u6/N23 ) );
  NOR2_X4 U2828 ( .A1(exp_r[1]), .A2(\u4/div_shft2[0] ), .ZN(net85030) );
  INV_X4 U2829 ( .A(n2002), .ZN(n2004) );
  NOR2_X4 U2830 ( .A1(n2004), .A2(n2003), .ZN(net85171) );
  NAND3_X2 U2831 ( .A1(n2040), .A2(quo[17]), .A3(net85674), .ZN(n2006) );
  OAI21_X4 U2832 ( .B1(n3074), .B2(net88319), .A(n2010), .ZN(net85150) );
  INV_X4 U2833 ( .A(n2011), .ZN(n2013) );
  NOR2_X4 U2834 ( .A1(n2013), .A2(n2012), .ZN(n2028) );
  NOR2_X4 U2835 ( .A1(n3073), .A2(net85716), .ZN(net85336) );
  NAND3_X4 U2836 ( .A1(n1894), .A2(quo[5]), .A3(net85676), .ZN(net85210) );
  NAND3_X4 U2837 ( .A1(n1922), .A2(quo[8]), .A3(net85674), .ZN(net85205) );
  NAND3_X2 U2838 ( .A1(net85076), .A2(net85676), .A3(quo[19]), .ZN(n2037) );
  NAND2_X2 U2839 ( .A1(net85316), .A2(exp_r[2]), .ZN(n2019) );
  INV_X4 U2840 ( .A(exp_r[4]), .ZN(net84290) );
  INV_X4 U2841 ( .A(exp_r[3]), .ZN(net84305) );
  NAND2_X2 U2842 ( .A1(exp_r[3]), .A2(net84290), .ZN(n2404) );
  INV_X4 U2843 ( .A(n2019), .ZN(n2406) );
  MUX2_X2 U2844 ( .A(net84290), .B(n2404), .S(n2406), .Z(n2020) );
  NAND2_X2 U2845 ( .A1(exp_r[4]), .A2(net84305), .ZN(n2405) );
  NAND2_X2 U2846 ( .A1(n2020), .A2(n2405), .ZN(\u4/exp_in_pl1[4] ) );
  XNOR2_X2 U2847 ( .A(net83968), .B(n2406), .ZN(n2442) );
  INV_X4 U2848 ( .A(n2442), .ZN(\u4/exp_in_pl1[3] ) );
  NAND3_X4 U2850 ( .A1(quo[6]), .A2(net85684), .A3(net85076), .ZN(net85067) );
  NAND3_X4 U2851 ( .A1(n2024), .A2(quo[16]), .A3(net85676), .ZN(net85068) );
  NAND3_X4 U2852 ( .A1(net85736), .A2(prod[12]), .A3(net85744), .ZN(n2021) );
  NAND3_X4 U2853 ( .A1(n2023), .A2(n2022), .A3(n2021), .ZN(net85196) );
  NAND3_X4 U2854 ( .A1(net89129), .A2(quo[4]), .A3(net88427), .ZN(net85194) );
  NAND3_X4 U2855 ( .A1(n1942), .A2(quo[14]), .A3(net85676), .ZN(net85195) );
  OAI21_X4 U2856 ( .B1(n3072), .B2(net88319), .A(n2032), .ZN(net85212) );
  NAND3_X4 U2857 ( .A1(n2001), .A2(quo[3]), .A3(net85674), .ZN(net85071) );
  NAND3_X4 U2858 ( .A1(n2016), .A2(quo[6]), .A3(net85674), .ZN(net85041) );
  NAND3_X4 U2859 ( .A1(n2014), .A2(quo[9]), .A3(net85676), .ZN(net85046) );
  NOR3_X4 U2860 ( .A1(net85232), .A2(n2041), .A3(net85196), .ZN(n2044) );
  NAND3_X4 U2861 ( .A1(n2024), .A2(quo[15]), .A3(net85676), .ZN(n2067) );
  OAI21_X4 U2862 ( .B1(n3075), .B2(net88319), .A(n2042), .ZN(n2065) );
  NAND4_X2 U2863 ( .A1(net90144), .A2(net85068), .A3(net85069), .A4(net85067), 
        .ZN(net85140) );
  NOR2_X4 U2864 ( .A1(net85200), .A2(n2048), .ZN(net85182) );
  INV_X4 U2865 ( .A(n2055), .ZN(n2053) );
  INV_X4 U2866 ( .A(net85127), .ZN(net84869) );
  INV_X4 U2867 ( .A(net85124), .ZN(net84531) );
  INV_X4 U2868 ( .A(net85111), .ZN(net84749) );
  NAND2_X2 U2869 ( .A1(net84749), .A2(n2190), .ZN(n2058) );
  XNOR2_X2 U2870 ( .A(n2059), .B(n2058), .ZN(n2448) );
  OAI21_X4 U2871 ( .B1(net89546), .B2(net88618), .A(net84758), .ZN(net85091)
         );
  OAI21_X4 U2872 ( .B1(n1940), .B2(net85093), .A(n2060), .ZN(
        \u4/fi_ldz_mi1[2] ) );
  MUX2_X2 U2873 ( .A(net84290), .B(n2404), .S(net84916), .Z(n2061) );
  NAND2_X2 U2874 ( .A1(prod[0]), .A2(net86125), .ZN(n2064) );
  NAND2_X2 U2875 ( .A1(net89998), .A2(n1660), .ZN(n2062) );
  NAND3_X4 U2876 ( .A1(n2064), .A2(n2063), .A3(n2062), .ZN(n3319) );
  INV_X4 U2877 ( .A(n2069), .ZN(n2072) );
  NOR3_X4 U2878 ( .A1(n2073), .A2(n2072), .A3(n2071), .ZN(n2074) );
  INV_X4 U2879 ( .A(net85039), .ZN(net85037) );
  XNOR2_X2 U2880 ( .A(exp_r[2]), .B(net85030), .ZN(\u4/f2i_shft[2] ) );
  INV_X4 U2881 ( .A(net84822), .ZN(net85027) );
  INV_X4 U2882 ( .A(n2225), .ZN(n2075) );
  NAND3_X4 U2883 ( .A1(net83959), .A2(n2226), .A3(net84236), .ZN(n2099) );
  NAND2_X2 U2884 ( .A1(net84341), .A2(net85847), .ZN(net83951) );
  XNOR2_X2 U2885 ( .A(div_opa_ldz_r2[2]), .B(exp_r[2]), .ZN(n2122) );
  INV_X4 U2886 ( .A(div_opa_ldz_r2[0]), .ZN(net84762) );
  NOR2_X4 U2887 ( .A1(net85832), .A2(net84762), .ZN(n2100) );
  INV_X4 U2888 ( .A(n2103), .ZN(n2076) );
  XNOR2_X2 U2889 ( .A(n2122), .B(n2108), .ZN(n2234) );
  INV_X4 U2890 ( .A(\u4/f2i_shft[2] ), .ZN(n2077) );
  NAND2_X2 U2891 ( .A1(net85006), .A2(net84982), .ZN(net84867) );
  NOR2_X4 U2892 ( .A1(net83421), .A2(n2153), .ZN(n2083) );
  INV_X4 U2893 ( .A(net11671), .ZN(net84992) );
  NAND2_X2 U2894 ( .A1(net83941), .A2(net85710), .ZN(n2089) );
  NAND2_X2 U2895 ( .A1(n2090), .A2(n2089), .ZN(n2092) );
  NOR3_X4 U2896 ( .A1(n2093), .A2(n2092), .A3(n2091), .ZN(n2098) );
  NAND2_X2 U2897 ( .A1(net85710), .A2(net84982), .ZN(n2095) );
  NAND2_X2 U2898 ( .A1(net85832), .A2(net84762), .ZN(n2131) );
  INV_X4 U2899 ( .A(n2100), .ZN(n2101) );
  NAND2_X2 U2900 ( .A1(n2131), .A2(n2101), .ZN(net84600) );
  INV_X4 U2901 ( .A(net84236), .ZN(net83969) );
  INV_X4 U2902 ( .A(n2102), .ZN(n2105) );
  INV_X4 U2903 ( .A(n2131), .ZN(n2104) );
  INV_X4 U2904 ( .A(n2106), .ZN(n2972) );
  INV_X4 U2905 ( .A(n2122), .ZN(n2107) );
  XNOR2_X2 U2906 ( .A(n2972), .B(n2107), .ZN(n2125) );
  INV_X4 U2907 ( .A(n2108), .ZN(n2110) );
  NAND2_X2 U2908 ( .A1(div_opa_ldz_r2[2]), .A2(net11560), .ZN(n2971) );
  INV_X4 U2909 ( .A(n2971), .ZN(n2109) );
  NAND2_X2 U2910 ( .A1(exp_r[2]), .A2(n3096), .ZN(n2970) );
  OAI21_X4 U2911 ( .B1(n2110), .B2(n2109), .A(n2970), .ZN(n2111) );
  INV_X4 U2912 ( .A(n2111), .ZN(n2146) );
  NAND2_X2 U2913 ( .A1(net83968), .A2(n1663), .ZN(n2112) );
  OAI21_X4 U2914 ( .B1(n2146), .B2(n2113), .A(n2112), .ZN(n2148) );
  INV_X4 U2915 ( .A(n2148), .ZN(n2117) );
  INV_X4 U2916 ( .A(n2634), .ZN(n2118) );
  NAND2_X2 U2917 ( .A1(n2118), .A2(net83439), .ZN(n2989) );
  NAND2_X2 U2918 ( .A1(n2634), .A2(net83439), .ZN(net83361) );
  INV_X4 U2919 ( .A(net83361), .ZN(net84886) );
  NAND2_X2 U2920 ( .A1(net84886), .A2(n2119), .ZN(n2124) );
  INV_X4 U2921 ( .A(net83439), .ZN(net83364) );
  NAND2_X2 U2922 ( .A1(div_opa_ldz_r2[0]), .A2(net85832), .ZN(n2132) );
  XNOR2_X2 U2923 ( .A(n2122), .B(n2281), .ZN(n2289) );
  NAND2_X2 U2924 ( .A1(net83364), .A2(n2289), .ZN(n2123) );
  OAI211_X2 U2925 ( .C1(n2125), .C2(n2989), .A(n2124), .B(n2123), .ZN(n2127)
         );
  INV_X4 U2926 ( .A(net84916), .ZN(net84921) );
  NAND2_X2 U2927 ( .A1(net84921), .A2(n2225), .ZN(n2217) );
  INV_X4 U2928 ( .A(n2217), .ZN(n2306) );
  INV_X4 U2929 ( .A(n872), .ZN(net84915) );
  NAND2_X2 U2930 ( .A1(net86169), .A2(net84915), .ZN(n2128) );
  NAND2_X2 U2931 ( .A1(n2129), .A2(n2128), .ZN(\u4/shift_right [2]) );
  XNOR2_X2 U2932 ( .A(net83968), .B(net84916), .ZN(net84858) );
  INV_X4 U2933 ( .A(n2991), .ZN(n2130) );
  NAND2_X2 U2934 ( .A1(n2130), .A2(net85710), .ZN(n2140) );
  INV_X4 U2935 ( .A(net83936), .ZN(net84907) );
  NAND2_X2 U2936 ( .A1(net84906), .A2(net84907), .ZN(net84637) );
  XNOR2_X2 U2937 ( .A(n2133), .B(n2131), .ZN(n2137) );
  XNOR2_X2 U2938 ( .A(n2133), .B(n2132), .ZN(n2290) );
  INV_X4 U2939 ( .A(n2290), .ZN(n2134) );
  NAND2_X2 U2940 ( .A1(net83364), .A2(n2134), .ZN(n2136) );
  INV_X4 U2941 ( .A(net83361), .ZN(net84900) );
  NAND2_X2 U2942 ( .A1(net84900), .A2(net84901), .ZN(n2135) );
  OAI211_X2 U2943 ( .C1(n2989), .C2(n2137), .A(n2136), .B(n2135), .ZN(n2138)
         );
  NAND2_X2 U2944 ( .A1(net85790), .A2(n2138), .ZN(n2141) );
  NAND4_X2 U2945 ( .A1(n2140), .A2(net84637), .A3(n2141), .A4(net84659), .ZN(
        n2143) );
  INV_X4 U2946 ( .A(net89926), .ZN(net84890) );
  INV_X4 U2947 ( .A(n2226), .ZN(n2580) );
  XNOR2_X2 U2948 ( .A(n2146), .B(n1579), .ZN(n2147) );
  INV_X4 U2949 ( .A(n2147), .ZN(n2263) );
  XNOR2_X2 U2950 ( .A(n2288), .B(n2148), .ZN(n2149) );
  INV_X4 U2951 ( .A(n2149), .ZN(n2243) );
  MUX2_X2 U2952 ( .A(n2150), .B(n1663), .S(net83933), .Z(n2151) );
  INV_X4 U2953 ( .A(\u4/exp_in_pl1[4] ), .ZN(n2155) );
  NAND2_X2 U2954 ( .A1(n2442), .A2(n2155), .ZN(n2156) );
  NAND2_X2 U2955 ( .A1(n2157), .A2(n2156), .ZN(net84848) );
  NAND2_X2 U2956 ( .A1(rmode_r3[1]), .A2(rmode_r3[0]), .ZN(n2248) );
  NAND2_X2 U2957 ( .A1(n1614), .A2(n1768), .ZN(net84326) );
  INV_X4 U2958 ( .A(net11558), .ZN(net83968) );
  NAND2_X2 U2959 ( .A1(n2562), .A2(net83968), .ZN(n2303) );
  NOR2_X4 U2960 ( .A1(n2158), .A2(net83963), .ZN(net84048) );
  OAI21_X4 U2961 ( .B1(n2159), .B2(n2248), .A(net84048), .ZN(net83942) );
  INV_X4 U2962 ( .A(net84778), .ZN(net84520) );
  NAND2_X2 U2963 ( .A1(\u4/N406 ), .A2(net84520), .ZN(net84840) );
  INV_X4 U2964 ( .A(\u4/N405 ), .ZN(n2161) );
  OAI21_X4 U2965 ( .B1(net84778), .B2(n2161), .A(n2160), .ZN(\u4/fract_out[5] ) );
  NAND2_X2 U2966 ( .A1(\u4/N402 ), .A2(net84520), .ZN(n2170) );
  INV_X4 U2967 ( .A(\u4/N401 ), .ZN(n2163) );
  NAND2_X2 U2968 ( .A1(\u4/N400 ), .A2(net84520), .ZN(net84810) );
  NOR3_X4 U2969 ( .A1(\u4/N419 ), .A2(\u4/N420 ), .A3(\u4/N418 ), .ZN(n2165)
         );
  NAND2_X2 U2970 ( .A1(net85828), .A2(n2579), .ZN(n2168) );
  NAND2_X2 U2971 ( .A1(net85828), .A2(net11566), .ZN(n2322) );
  NAND2_X2 U2972 ( .A1(\u4/N399 ), .A2(net84520), .ZN(net84564) );
  INV_X4 U2973 ( .A(net84564), .ZN(net84784) );
  NAND3_X2 U2974 ( .A1(n3055), .A2(n3056), .A3(n3054), .ZN(n2178) );
  NAND3_X2 U2975 ( .A1(n3060), .A2(n3061), .A3(n3059), .ZN(n2176) );
  NAND3_X2 U2976 ( .A1(n3063), .A2(n3064), .A3(n3062), .ZN(n2175) );
  NOR4_X2 U2977 ( .A1(n2178), .A2(n2177), .A3(n2176), .A4(n2175), .ZN(n2179)
         );
  NAND2_X2 U2978 ( .A1(n2548), .A2(net85790), .ZN(net83913) );
  INV_X4 U2979 ( .A(net83913), .ZN(net84783) );
  NOR3_X4 U2980 ( .A1(\u4/N423 ), .A2(net84783), .A3(net84784), .ZN(n2186) );
  NOR3_X4 U2981 ( .A1(\u4/N390 ), .A2(\u4/N392 ), .A3(\u4/N388 ), .ZN(n2184)
         );
  NOR4_X2 U2982 ( .A1(\u4/N394 ), .A2(\u4/N395 ), .A3(\u4/N389 ), .A4(
        \u4/N391 ), .ZN(n2183) );
  NOR4_X2 U2983 ( .A1(\u4/N398 ), .A2(\u4/N396 ), .A3(\u4/N393 ), .A4(
        \u4/N397 ), .ZN(n2182) );
  INV_X4 U2984 ( .A(n2301), .ZN(n2185) );
  NAND2_X2 U2985 ( .A1(n1640), .A2(n1589), .ZN(net84643) );
  MUX2_X2 U2986 ( .A(\u4/exp_in_pl1[4] ), .B(\u4/exp_next_mi[4] ), .S(net85788), .Z(net84764) );
  NAND2_X2 U2987 ( .A1(rmode_r3[1]), .A2(net86016), .ZN(net84490) );
  INV_X4 U2988 ( .A(net83402), .ZN(net84633) );
  INV_X4 U2989 ( .A(\u4/exp_next_mi[3] ), .ZN(net84768) );
  MUX2_X2 U2990 ( .A(n2442), .B(net84768), .S(net85788), .Z(net84445) );
  MUX2_X2 U2991 ( .A(net85712), .B(net89692), .S(net85788), .Z(net84767) );
  INV_X4 U2992 ( .A(net84767), .ZN(net84766) );
  XOR2_X2 U2993 ( .A(net84764), .B(net84765), .Z(n2231) );
  NOR2_X4 U2994 ( .A1(n2189), .A2(n2188), .ZN(n2260) );
  XNOR2_X2 U2995 ( .A(n2443), .B(div_opa_ldz_r2[3]), .ZN(n2193) );
  XNOR2_X2 U2996 ( .A(n2193), .B(n2196), .ZN(n2551) );
  NAND2_X2 U2997 ( .A1(\u4/exp_in_pl1[3] ), .A2(n2551), .ZN(n2194) );
  INV_X4 U2998 ( .A(n2443), .ZN(n2401) );
  NOR2_X4 U2999 ( .A1(div_opa_ldz_r2[3]), .A2(n2401), .ZN(n2198) );
  NAND2_X2 U3000 ( .A1(n2401), .A2(div_opa_ldz_r2[3]), .ZN(n2197) );
  OAI21_X4 U3001 ( .B1(n2199), .B2(n2198), .A(n2197), .ZN(n2549) );
  XNOR2_X2 U3002 ( .A(n2549), .B(n2200), .ZN(n2552) );
  XNOR2_X2 U3003 ( .A(n2552), .B(\u4/exp_in_pl1[4] ), .ZN(n2201) );
  XNOR2_X2 U3004 ( .A(n2202), .B(n2201), .ZN(n2229) );
  INV_X4 U3005 ( .A(net11560), .ZN(net83994) );
  INV_X4 U3006 ( .A(net11564), .ZN(net83967) );
  NAND2_X2 U3007 ( .A1(n3096), .A2(net83994), .ZN(n2206) );
  NAND2_X2 U3008 ( .A1(net11671), .A2(net83993), .ZN(n2205) );
  OAI211_X2 U3009 ( .C1(n2208), .C2(n2207), .A(n2206), .B(n2205), .ZN(n2211)
         );
  INV_X4 U3010 ( .A(n1663), .ZN(n2209) );
  AOI21_X2 U3011 ( .B1(n2212), .B2(n2211), .A(n2210), .ZN(n2214) );
  XNOR2_X2 U3012 ( .A(n2222), .B(n2443), .ZN(n2422) );
  XNOR2_X2 U3013 ( .A(n2225), .B(net84305), .ZN(n2992) );
  NAND2_X2 U3014 ( .A1(n2422), .A2(n2992), .ZN(n2221) );
  NAND2_X2 U3015 ( .A1(net89964), .A2(net85710), .ZN(n2215) );
  NOR2_X4 U3016 ( .A1(n2422), .A2(n2992), .ZN(n2220) );
  XNOR2_X2 U3017 ( .A(n2224), .B(n2242), .ZN(n2228) );
  NAND2_X2 U3018 ( .A1(n2227), .A2(n2226), .ZN(n2981) );
  XNOR2_X2 U3019 ( .A(n2228), .B(n2981), .ZN(n2311) );
  OAI22_X2 U3020 ( .A1(n2229), .A2(net84611), .B1(n2311), .B2(net88427), .ZN(
        n2230) );
  AOI21_X2 U3021 ( .B1(net84633), .B2(n2231), .A(n2230), .ZN(n2247) );
  INV_X4 U3022 ( .A(n2965), .ZN(n2237) );
  INV_X4 U3023 ( .A(n2234), .ZN(n2964) );
  NOR2_X4 U3024 ( .A1(net83407), .A2(n2964), .ZN(n2236) );
  NAND2_X2 U3025 ( .A1(n2964), .A2(net83407), .ZN(n2235) );
  OAI21_X4 U3026 ( .B1(n2237), .B2(n2236), .A(n2235), .ZN(n2264) );
  INV_X4 U3027 ( .A(n2264), .ZN(n2241) );
  INV_X4 U3028 ( .A(n2422), .ZN(n2238) );
  NAND2_X2 U3029 ( .A1(n2263), .A2(n2238), .ZN(n2239) );
  INV_X4 U3030 ( .A(n2242), .ZN(n2421) );
  XNOR2_X2 U3031 ( .A(n2243), .B(n2421), .ZN(n2244) );
  XNOR2_X2 U3032 ( .A(n2245), .B(n2244), .ZN(n2246) );
  INV_X4 U3033 ( .A(net84669), .ZN(net84619) );
  MUX2_X2 U3034 ( .A(n2247), .B(n2246), .S(net84619), .Z(net83995) );
  INV_X4 U3035 ( .A(n2248), .ZN(n2249) );
  NAND4_X2 U3036 ( .A1(n2249), .A2(opas_r2), .A3(net83936), .A4(net84048), 
        .ZN(net84488) );
  NAND2_X2 U3037 ( .A1(n2401), .A2(n2253), .ZN(net84639) );
  XNOR2_X2 U3038 ( .A(n2251), .B(n2250), .ZN(n2307) );
  INV_X4 U3039 ( .A(net84659), .ZN(net84656) );
  INV_X4 U3040 ( .A(net84652), .ZN(net83934) );
  INV_X4 U3041 ( .A(net83429), .ZN(net84647) );
  NAND2_X2 U3042 ( .A1(net84647), .A2(net84490), .ZN(net84449) );
  INV_X4 U3043 ( .A(n2962), .ZN(n2252) );
  NAND3_X4 U3044 ( .A1(net84644), .A2(net84645), .A3(n2252), .ZN(n2358) );
  INV_X4 U3045 ( .A(net84642), .ZN(net84632) );
  NAND2_X2 U3046 ( .A1(n2254), .A2(n2443), .ZN(n2255) );
  INV_X4 U3047 ( .A(net84637), .ZN(net83423) );
  NAND2_X2 U3048 ( .A1(net84632), .A2(net84633), .ZN(net84624) );
  XNOR2_X2 U3049 ( .A(n2551), .B(n2442), .ZN(n2259) );
  XNOR2_X2 U3050 ( .A(n2260), .B(n2259), .ZN(net84629) );
  XNOR2_X2 U3051 ( .A(n2422), .B(n2992), .ZN(n2262) );
  XNOR2_X2 U3052 ( .A(n2262), .B(n2261), .ZN(n2309) );
  XNOR2_X2 U3053 ( .A(n2263), .B(n2422), .ZN(n2265) );
  XNOR2_X2 U3054 ( .A(n2265), .B(n2264), .ZN(n2266) );
  NAND2_X2 U3055 ( .A1(n2267), .A2(net84614), .ZN(n2331) );
  OAI21_X4 U3056 ( .B1(n2268), .B2(n2331), .A(net83429), .ZN(n2357) );
  NAND2_X2 U3057 ( .A1(net84160), .A2(net84166), .ZN(n2366) );
  INV_X4 U3058 ( .A(net84605), .ZN(net84604) );
  INV_X4 U3059 ( .A(net84600), .ZN(net83438) );
  NAND2_X2 U3060 ( .A1(\u4/exp_f2i_1 [23]), .A2(n1606), .ZN(n2271) );
  INV_X4 U3061 ( .A(n2271), .ZN(n2272) );
  NOR4_X2 U3062 ( .A1(n2274), .A2(n2273), .A3(net84595), .A4(n2272), .ZN(
        net84474) );
  NAND2_X2 U3063 ( .A1(net84591), .A2(n1589), .ZN(net84579) );
  NAND2_X2 U3064 ( .A1(net84590), .A2(net83429), .ZN(net84475) );
  NAND2_X2 U3065 ( .A1(n2275), .A2(net84564), .ZN(n2546) );
  INV_X4 U3066 ( .A(n2546), .ZN(n2278) );
  NAND2_X2 U3067 ( .A1(n2278), .A2(n2277), .ZN(n2280) );
  OAI21_X4 U3068 ( .B1(net84555), .B2(n2280), .A(n2279), .ZN(net84403) );
  NAND2_X2 U3069 ( .A1(sign), .A2(net84403), .ZN(net84482) );
  INV_X4 U3070 ( .A(net84550), .ZN(net84548) );
  NAND2_X2 U3071 ( .A1(net83968), .A2(div_opa_ldz_r2[3]), .ZN(n2286) );
  INV_X4 U3072 ( .A(n2281), .ZN(n2284) );
  NAND2_X2 U3073 ( .A1(exp_r[2]), .A2(div_opa_ldz_r2[2]), .ZN(n2282) );
  NAND2_X2 U3074 ( .A1(n2286), .A2(n2285), .ZN(n2287) );
  XNOR2_X2 U3075 ( .A(n2288), .B(n2287), .ZN(n2978) );
  INV_X4 U3076 ( .A(n2978), .ZN(n2297) );
  INV_X4 U3077 ( .A(n2289), .ZN(n2291) );
  NAND2_X2 U3078 ( .A1(n2291), .A2(n2290), .ZN(n2294) );
  INV_X4 U3079 ( .A(n2292), .ZN(n2293) );
  XNOR2_X2 U3080 ( .A(n1579), .B(n2293), .ZN(n2987) );
  NAND2_X2 U3081 ( .A1(n2294), .A2(n2987), .ZN(n2296) );
  NAND2_X2 U3082 ( .A1(net84531), .A2(net84532), .ZN(n2295) );
  NAND2_X2 U3083 ( .A1(net84520), .A2(n2301), .ZN(n2545) );
  NAND2_X2 U3084 ( .A1(net83950), .A2(n2302), .ZN(net84327) );
  INV_X4 U3085 ( .A(net84327), .ZN(net84334) );
  INV_X4 U3086 ( .A(n2322), .ZN(n2305) );
  INV_X4 U3087 ( .A(n2303), .ZN(n2304) );
  NAND3_X2 U3088 ( .A1(n2309), .A2(n2366), .A3(n2308), .ZN(n2310) );
  NAND3_X4 U3089 ( .A1(n2311), .A2(n2310), .A3(net84506), .ZN(n2420) );
  INV_X4 U3090 ( .A(net84469), .ZN(net84501) );
  INV_X4 U3091 ( .A(net83927), .ZN(net84498) );
  OAI21_X4 U3092 ( .B1(n2312), .B2(n2420), .A(net84500), .ZN(n2316) );
  NAND2_X2 U3093 ( .A1(net84498), .A2(net85794), .ZN(n2314) );
  INV_X4 U3094 ( .A(net83844), .ZN(net84465) );
  INV_X4 U3095 ( .A(n2420), .ZN(n2317) );
  OAI21_X4 U3096 ( .B1(n2319), .B2(net84490), .A(n2318), .ZN(net84332) );
  INV_X4 U3097 ( .A(net84332), .ZN(net83855) );
  INV_X4 U3098 ( .A(net84488), .ZN(net84487) );
  NAND2_X2 U3099 ( .A1(net84487), .A2(net83941), .ZN(n2600) );
  NAND3_X4 U3100 ( .A1(net83855), .A2(n2600), .A3(n2320), .ZN(net84220) );
  NAND2_X2 U3101 ( .A1(n1603), .A2(net84211), .ZN(n2474) );
  NOR2_X4 U3102 ( .A1(net83296), .A2(net84150), .ZN(n2339) );
  INV_X4 U3103 ( .A(net84312), .ZN(net84366) );
  NAND2_X2 U3104 ( .A1(n2437), .A2(n2420), .ZN(n2424) );
  NAND2_X2 U3105 ( .A1(rmode_r3[0]), .A2(n1768), .ZN(n2588) );
  INV_X4 U3106 ( .A(n2588), .ZN(n2425) );
  NAND2_X2 U3107 ( .A1(n2425), .A2(n1597), .ZN(n2326) );
  NOR2_X4 U3108 ( .A1(n2420), .A2(n2588), .ZN(n2415) );
  OAI21_X4 U3109 ( .B1(net85828), .B2(net83927), .A(n2420), .ZN(n2327) );
  INV_X4 U3110 ( .A(n2543), .ZN(n2328) );
  AOI211_X4 U3111 ( .C1(net83969), .C2(n2424), .A(n2329), .B(n2328), .ZN(n2458) );
  INV_X4 U3112 ( .A(n2329), .ZN(n2330) );
  NAND2_X2 U3113 ( .A1(sign), .A2(rmode_r3[1]), .ZN(n2416) );
  NAND2_X2 U3114 ( .A1(net84080), .A2(net85794), .ZN(n2340) );
  NOR2_X4 U3115 ( .A1(n2458), .A2(n2521), .ZN(n2335) );
  NAND2_X2 U3116 ( .A1(net84343), .A2(net84398), .ZN(n2494) );
  NAND2_X2 U3117 ( .A1(net84450), .A2(net85847), .ZN(net84134) );
  INV_X4 U3118 ( .A(net84134), .ZN(net84368) );
  INV_X4 U3119 ( .A(n2331), .ZN(n2332) );
  OAI21_X4 U3120 ( .B1(net84445), .B2(net83432), .A(n2332), .ZN(net84148) );
  NAND2_X2 U3121 ( .A1(net84368), .A2(net84148), .ZN(n2388) );
  NAND3_X4 U3122 ( .A1(n2490), .A2(n2494), .A3(n2338), .ZN(n2454) );
  INV_X4 U3123 ( .A(n2333), .ZN(n2334) );
  NAND2_X2 U3124 ( .A1(net84133), .A2(n2388), .ZN(n2338) );
  NAND4_X2 U3125 ( .A1(n1648), .A2(n2496), .A3(n1588), .A4(n2491), .ZN(n2346)
         );
  INV_X4 U3126 ( .A(n2340), .ZN(n2343) );
  INV_X4 U3127 ( .A(n2341), .ZN(n2342) );
  NOR2_X4 U3128 ( .A1(n2348), .A2(n2347), .ZN(n2612) );
  NAND3_X4 U3129 ( .A1(n1603), .A2(n2996), .A3(net84211), .ZN(net84218) );
  NAND2_X2 U3130 ( .A1(net84081), .A2(net84218), .ZN(n2349) );
  INV_X4 U3131 ( .A(n2437), .ZN(n2426) );
  XNOR2_X2 U3132 ( .A(n2996), .B(n2426), .ZN(n2351) );
  NAND2_X2 U3133 ( .A1(n2353), .A2(n2352), .ZN(net84333) );
  NAND2_X2 U3134 ( .A1(n2358), .A2(n2357), .ZN(n2360) );
  NOR3_X4 U3135 ( .A1(n2361), .A2(n2437), .A3(n1597), .ZN(net84374) );
  INV_X4 U3136 ( .A(n2419), .ZN(n2462) );
  INV_X4 U3137 ( .A(n2461), .ZN(n2363) );
  INV_X4 U3138 ( .A(n2566), .ZN(n2555) );
  INV_X4 U3139 ( .A(n2366), .ZN(n2368) );
  AOI211_X4 U3140 ( .C1(n2370), .C2(n2371), .A(net84352), .B(n2369), .ZN(n2436) );
  INV_X4 U3141 ( .A(n2375), .ZN(n2611) );
  NAND2_X2 U3142 ( .A1(n2611), .A2(n2612), .ZN(net84344) );
  INV_X4 U3143 ( .A(net84344), .ZN(net83754) );
  NAND2_X2 U3144 ( .A1(n3065), .A2(n3071), .ZN(n2698) );
  NAND2_X2 U3145 ( .A1(net84343), .A2(n2698), .ZN(n2585) );
  NAND2_X2 U3146 ( .A1(n1640), .A2(n1576), .ZN(n2379) );
  NAND2_X2 U3147 ( .A1(n2380), .A2(n2379), .ZN(n2683) );
  OAI21_X4 U3148 ( .B1(net84334), .B2(net84326), .A(n2588), .ZN(n2381) );
  OAI21_X4 U3149 ( .B1(n2382), .B2(n2381), .A(net84095), .ZN(n2514) );
  OAI21_X4 U3150 ( .B1(n2385), .B2(n2384), .A(net84095), .ZN(n2513) );
  INV_X4 U3151 ( .A(\u4/fract_out_pl1[0] ), .ZN(n2386) );
  INV_X4 U3152 ( .A(n2416), .ZN(n2387) );
  NOR2_X4 U3153 ( .A1(n2389), .A2(n2388), .ZN(n2391) );
  INV_X4 U3154 ( .A(n2600), .ZN(n2390) );
  AOI211_X4 U3155 ( .C1(n2392), .C2(n2391), .A(net83878), .B(n2390), .ZN(
        net84253) );
  INV_X4 U3156 ( .A(net84315), .ZN(net84314) );
  OAI21_X4 U3157 ( .B1(n2465), .B2(n2396), .A(n2395), .ZN(n2449) );
  XNOR2_X2 U3158 ( .A(exp_r[4]), .B(n2399), .ZN(n2414) );
  NAND2_X2 U3159 ( .A1(\u4/exp_in_pl1[3] ), .A2(n2401), .ZN(n2403) );
  INV_X4 U3160 ( .A(n2404), .ZN(n2409) );
  INV_X4 U3161 ( .A(n2405), .ZN(n2407) );
  MUX2_X2 U3162 ( .A(n2407), .B(net84290), .S(n2406), .Z(n2408) );
  XNOR2_X2 U3163 ( .A(n2412), .B(n2411), .ZN(n2413) );
  OAI22_X2 U3164 ( .A1(n2414), .A2(n2482), .B1(n2413), .B2(n2486), .ZN(
        net84076) );
  INV_X4 U3165 ( .A(net84076), .ZN(net84280) );
  NOR2_X4 U3166 ( .A1(net84276), .A2(net84277), .ZN(net84200) );
  INV_X4 U3167 ( .A(n2415), .ZN(n2417) );
  NAND2_X2 U3168 ( .A1(n1583), .A2(n2419), .ZN(net84266) );
  NAND2_X2 U3169 ( .A1(net84265), .A2(net84266), .ZN(net83864) );
  INV_X4 U3170 ( .A(net83864), .ZN(net83876) );
  INV_X4 U3171 ( .A(n2420), .ZN(n2438) );
  INV_X4 U3172 ( .A(n2423), .ZN(n2439) );
  OAI211_X2 U3173 ( .C1(n2438), .C2(n2439), .A(n2424), .B(net83969), .ZN(n2427) );
  OAI21_X4 U3174 ( .B1(n2438), .B2(n2426), .A(n2425), .ZN(n2542) );
  NAND3_X2 U3175 ( .A1(n2427), .A2(n2542), .A3(n2543), .ZN(n2622) );
  NAND2_X2 U3176 ( .A1(net83876), .A2(n2622), .ZN(net84254) );
  INV_X4 U3177 ( .A(n2683), .ZN(n2433) );
  NAND2_X2 U3178 ( .A1(opa_inf), .A2(n1613), .ZN(n2432) );
  INV_X4 U3179 ( .A(net83781), .ZN(net84249) );
  NAND3_X2 U3180 ( .A1(n2432), .A2(n2431), .A3(n2430), .ZN(n2956) );
  AOI21_X4 U3181 ( .B1(n2439), .B2(n2426), .A(n2438), .ZN(n2440) );
  NOR2_X4 U3182 ( .A1(n2440), .A2(net84236), .ZN(n2541) );
  NAND2_X2 U3183 ( .A1(n2543), .A2(n2542), .ZN(n2441) );
  INV_X4 U3184 ( .A(n2486), .ZN(n2447) );
  XNOR2_X2 U3185 ( .A(n2443), .B(n2442), .ZN(n2445) );
  XNOR2_X2 U3186 ( .A(n2445), .B(n2444), .ZN(n2446) );
  NAND2_X2 U3187 ( .A1(n2447), .A2(n2446), .ZN(net84215) );
  INV_X4 U3188 ( .A(n2482), .ZN(n2452) );
  XNOR2_X2 U3189 ( .A(n2450), .B(n2449), .ZN(n2451) );
  NAND2_X2 U3190 ( .A1(n2452), .A2(n2451), .ZN(net84216) );
  INV_X4 U3191 ( .A(n2454), .ZN(n2477) );
  NAND3_X2 U3192 ( .A1(n2455), .A2(n2496), .A3(n2477), .ZN(n2456) );
  NAND2_X2 U3193 ( .A1(n2463), .A2(n2462), .ZN(n2475) );
  XNOR2_X2 U3194 ( .A(n2465), .B(n2464), .ZN(n2466) );
  XNOR2_X2 U3195 ( .A(n2468), .B(n2467), .ZN(n2469) );
  NAND4_X2 U3196 ( .A1(n2475), .A2(n2474), .A3(net84081), .A4(n2473), .ZN(
        n2476) );
  INV_X4 U3197 ( .A(n2476), .ZN(n2524) );
  NAND2_X2 U3198 ( .A1(n2480), .A2(n2479), .ZN(n2526) );
  INV_X4 U3199 ( .A(net84166), .ZN(net84165) );
  XNOR2_X2 U3200 ( .A(n2481), .B(net84165), .ZN(n2483) );
  INV_X4 U3201 ( .A(net84160), .ZN(net84159) );
  XNOR2_X2 U3202 ( .A(n2484), .B(net84159), .ZN(n2487) );
  NAND2_X2 U3203 ( .A1(net89692), .A2(net84157), .ZN(n2485) );
  INV_X4 U3204 ( .A(net84148), .ZN(net84146) );
  NAND2_X2 U3205 ( .A1(net84146), .A2(net84133), .ZN(n2492) );
  NAND4_X2 U3206 ( .A1(n2493), .A2(n2492), .A3(n2491), .A4(n2490), .ZN(n2501)
         );
  NAND4_X2 U3207 ( .A1(n2497), .A2(n2496), .A3(n2495), .A4(n2494), .ZN(n2500)
         );
  INV_X4 U3208 ( .A(\u4/fract_out_pl1[7] ), .ZN(n2504) );
  OAI22_X2 U3209 ( .A1(n1928), .A2(n2504), .B1(n2503), .B2(n1961), .ZN(n2687)
         );
  INV_X4 U3210 ( .A(\u4/fract_out_pl1[8] ), .ZN(n2505) );
  OAI22_X2 U3211 ( .A1(net84119), .A2(n1961), .B1(n2513), .B2(n2505), .ZN(
        n2689) );
  INV_X4 U3212 ( .A(\u4/fract_out_pl1[9] ), .ZN(n2506) );
  NOR3_X4 U3213 ( .A1(n2687), .A2(n2689), .A3(n2691), .ZN(n2519) );
  INV_X4 U3214 ( .A(\u4/fract_out_pl1[5] ), .ZN(n2507) );
  OAI22_X2 U3215 ( .A1(net84115), .A2(n1961), .B1(n2513), .B2(n2507), .ZN(
        n2682) );
  INV_X4 U3216 ( .A(\u4/fract_out_pl1[6] ), .ZN(n2508) );
  NOR2_X4 U3217 ( .A1(n2682), .A2(n2685), .ZN(n2518) );
  INV_X4 U3218 ( .A(\u4/fract_out_pl1[2] ), .ZN(n2509) );
  INV_X4 U3219 ( .A(\u4/fract_out_pl1[3] ), .ZN(n2510) );
  INV_X4 U3220 ( .A(\u4/fract_out_pl1[4] ), .ZN(n2511) );
  INV_X4 U3221 ( .A(\u4/fract_out_pl1[1] ), .ZN(n2512) );
  NAND2_X2 U3222 ( .A1(net84095), .A2(net84096), .ZN(net84024) );
  NOR2_X4 U3223 ( .A1(n2522), .A2(n2521), .ZN(n2525) );
  OAI21_X4 U3224 ( .B1(n2525), .B2(net84059), .A(net83861), .ZN(n2706) );
  NAND3_X2 U3225 ( .A1(net83747), .A2(net84024), .A3(n2706), .ZN(n2529) );
  OAI21_X4 U3226 ( .B1(n2528), .B2(net84060), .A(net83861), .ZN(net83736) );
  INV_X4 U3227 ( .A(\u4/exp_next_mi[4] ), .ZN(n2530) );
  OAI211_X2 U3228 ( .C1(n2530), .C2(net84079), .A(net84080), .B(net84081), 
        .ZN(n2531) );
  NAND2_X2 U3229 ( .A1(opa_00), .A2(opb_00), .ZN(net84021) );
  NAND2_X2 U3230 ( .A1(opa_00), .A2(opb_inf), .ZN(n2533) );
  NAND2_X2 U3231 ( .A1(opa_inf), .A2(opb_00), .ZN(n2532) );
  NAND2_X2 U3232 ( .A1(n2533), .A2(n2532), .ZN(net83925) );
  NAND3_X2 U3233 ( .A1(n1561), .A2(n1570), .A3(n1595), .ZN(n2536) );
  INV_X4 U3234 ( .A(n2541), .ZN(n2544) );
  NAND3_X2 U3235 ( .A1(n2544), .A2(n2543), .A3(n2542), .ZN(net84003) );
  INV_X4 U3236 ( .A(n2545), .ZN(n2573) );
  NAND2_X2 U3237 ( .A1(n2547), .A2(net88950), .ZN(n2583) );
  INV_X4 U3238 ( .A(n2583), .ZN(n2572) );
  INV_X4 U3239 ( .A(n2548), .ZN(n2570) );
  INV_X4 U3240 ( .A(net83995), .ZN(net83973) );
  INV_X4 U3241 ( .A(n2549), .ZN(n2550) );
  INV_X4 U3242 ( .A(n2552), .ZN(n2554) );
  NAND2_X2 U3243 ( .A1(n2555), .A2(net83364), .ZN(n2558) );
  OAI21_X4 U3244 ( .B1(n2557), .B2(n2556), .A(n2558), .ZN(n2559) );
  INV_X4 U3245 ( .A(n2558), .ZN(n2565) );
  AOI21_X4 U3246 ( .B1(n2560), .B2(n2559), .A(n1646), .ZN(net83975) );
  MUX2_X2 U3247 ( .A(net83971), .B(net83972), .S(net11555), .Z(n2561) );
  INV_X4 U3248 ( .A(n2563), .ZN(n2564) );
  OAI21_X4 U3249 ( .B1(n2570), .B2(n2569), .A(n2568), .ZN(n2630) );
  NAND2_X2 U3250 ( .A1(net85828), .A2(n2630), .ZN(n2571) );
  NAND2_X2 U3251 ( .A1(n2629), .A2(net85790), .ZN(n2578) );
  NAND2_X2 U3252 ( .A1(n2583), .A2(net83951), .ZN(n2599) );
  INV_X4 U3253 ( .A(net83942), .ZN(net83940) );
  INV_X4 U3254 ( .A(n2601), .ZN(n2576) );
  NOR2_X4 U3255 ( .A1(n1605), .A2(n2576), .ZN(n2577) );
  NAND4_X2 U3256 ( .A1(net83906), .A2(n2578), .A3(n2599), .A4(n2577), .ZN(
        n2595) );
  NAND2_X2 U3257 ( .A1(net90047), .A2(net11566), .ZN(n2632) );
  NAND2_X2 U3258 ( .A1(n2582), .A2(n2581), .ZN(n2584) );
  NAND2_X2 U3259 ( .A1(net83836), .A2(n2639), .ZN(n2594) );
  NAND3_X2 U3260 ( .A1(n2585), .A2(n1572), .A3(n1595), .ZN(n2586) );
  NAND2_X2 U3261 ( .A1(n2587), .A2(n2586), .ZN(n2662) );
  INV_X4 U3262 ( .A(n2662), .ZN(n2591) );
  INV_X4 U3263 ( .A(n2698), .ZN(n2589) );
  INV_X4 U3264 ( .A(n2605), .ZN(n2619) );
  NAND3_X2 U3265 ( .A1(n2592), .A2(n2600), .A3(net83913), .ZN(n2593) );
  INV_X4 U3266 ( .A(n2599), .ZN(n2603) );
  NAND2_X2 U3267 ( .A1(n2601), .A2(n2600), .ZN(n2602) );
  NAND2_X2 U3268 ( .A1(net83747), .A2(net91075), .ZN(n2699) );
  NAND2_X2 U3269 ( .A1(n1574), .A2(net85790), .ZN(n2604) );
  AND3_X2 U3270 ( .A1(n2605), .A2(n2699), .A3(n2604), .ZN(n2606) );
  INV_X4 U3271 ( .A(n2614), .ZN(n2608) );
  NAND2_X2 U3272 ( .A1(n2614), .A2(net85794), .ZN(n2615) );
  INV_X4 U3273 ( .A(net83883), .ZN(net83806) );
  AOI21_X2 U3274 ( .B1(net83876), .B2(n2622), .A(net83878), .ZN(net83874) );
  NOR2_X4 U3275 ( .A1(net83869), .A2(net83864), .ZN(n2624) );
  OAI21_X4 U3276 ( .B1(n2624), .B2(net83868), .A(net83861), .ZN(n2707) );
  NAND2_X2 U3277 ( .A1(underflow_fmul_r[2]), .A2(n1550), .ZN(net83821) );
  NOR3_X4 U3278 ( .A1(net83856), .A2(n2665), .A3(net83821), .ZN(n2646) );
  NAND2_X2 U3279 ( .A1(net83855), .A2(net85790), .ZN(n2628) );
  INV_X4 U3280 ( .A(n2629), .ZN(n2638) );
  INV_X4 U3281 ( .A(n2630), .ZN(n2631) );
  MUX2_X2 U3282 ( .A(net83849), .B(n2631), .S(net85828), .Z(n2635) );
  NAND3_X2 U3283 ( .A1(n2635), .A2(n2634), .A3(n2633), .ZN(n2636) );
  NAND2_X2 U3284 ( .A1(n2636), .A2(net83844), .ZN(n2637) );
  NOR2_X4 U3285 ( .A1(n2638), .A2(n2637), .ZN(n2641) );
  INV_X4 U3286 ( .A(n2639), .ZN(n2640) );
  AOI21_X4 U3287 ( .B1(n2642), .B2(n2641), .A(n2640), .ZN(n2644) );
  INV_X4 U3288 ( .A(net83836), .ZN(net83833) );
  NOR2_X4 U3289 ( .A1(net83833), .A2(n1651), .ZN(n2643) );
  INV_X4 U3290 ( .A(net83821), .ZN(net83820) );
  NAND2_X2 U3291 ( .A1(n2649), .A2(n2648), .ZN(net83811) );
  INV_X4 U3292 ( .A(n3170), .ZN(n2650) );
  NAND4_X2 U3293 ( .A1(n3172), .A2(n3171), .A3(n2652), .A4(n2651), .ZN(
        net83812) );
  INV_X4 U3294 ( .A(n2653), .ZN(n2654) );
  NOR3_X2 U3295 ( .A1(net83807), .A2(net86016), .A3(n2654), .ZN(n2655) );
  INV_X4 U3296 ( .A(n2669), .ZN(n2667) );
  NAND4_X2 U3297 ( .A1(net83779), .A2(net91075), .A3(net83781), .A4(n1576), 
        .ZN(n2671) );
  NAND2_X2 U3298 ( .A1(n2433), .A2(n2685), .ZN(n2686) );
  NAND2_X2 U3299 ( .A1(n2433), .A2(n2687), .ZN(n2688) );
  NAND2_X2 U3300 ( .A1(n2433), .A2(n2691), .ZN(n2693) );
  INV_X4 U3301 ( .A(n2694), .ZN(n2697) );
  NOR2_X4 U3302 ( .A1(n2697), .A2(n2696), .ZN(n2705) );
  NAND2_X2 U3303 ( .A1(net83736), .A2(n2433), .ZN(N231) );
  NAND2_X2 U3304 ( .A1(n2708), .A2(n2433), .ZN(N233) );
  INV_X4 U3305 ( .A(N76), .ZN(n2710) );
  MUX2_X2 U3306 ( .A(n3120), .B(n2710), .S(n3012), .Z(n2711) );
  INV_X4 U3307 ( .A(n2711), .ZN(\u6/N22 ) );
  INV_X4 U3308 ( .A(N75), .ZN(n2712) );
  MUX2_X2 U3309 ( .A(n3119), .B(n2712), .S(n3012), .Z(n2713) );
  INV_X4 U3310 ( .A(n2713), .ZN(\u6/N21 ) );
  INV_X4 U3311 ( .A(N74), .ZN(n2714) );
  MUX2_X2 U3312 ( .A(n3118), .B(n2714), .S(n3012), .Z(n2715) );
  INV_X4 U3313 ( .A(n2715), .ZN(\u6/N20 ) );
  INV_X4 U3314 ( .A(N73), .ZN(n2716) );
  MUX2_X2 U3315 ( .A(n3117), .B(n2716), .S(n3012), .Z(n2717) );
  INV_X4 U3316 ( .A(n2717), .ZN(\u6/N19 ) );
  INV_X4 U3317 ( .A(N72), .ZN(n2718) );
  MUX2_X2 U3318 ( .A(n3116), .B(n2718), .S(n3012), .Z(n2719) );
  INV_X4 U3319 ( .A(n2719), .ZN(\u6/N18 ) );
  INV_X4 U3320 ( .A(N71), .ZN(n2720) );
  MUX2_X2 U3321 ( .A(n3115), .B(n2720), .S(n3012), .Z(n2721) );
  INV_X4 U3322 ( .A(n2721), .ZN(\u6/N17 ) );
  INV_X4 U3323 ( .A(N70), .ZN(n2722) );
  MUX2_X2 U3324 ( .A(n3114), .B(n2722), .S(n3012), .Z(n2723) );
  INV_X4 U3325 ( .A(n2723), .ZN(\u6/N16 ) );
  INV_X4 U3326 ( .A(N69), .ZN(n2724) );
  MUX2_X2 U3327 ( .A(n3113), .B(n2724), .S(n3012), .Z(n2725) );
  INV_X4 U3328 ( .A(n2725), .ZN(\u6/N15 ) );
  INV_X4 U3329 ( .A(N68), .ZN(n2726) );
  MUX2_X2 U3330 ( .A(n3112), .B(n2726), .S(n3012), .Z(n2727) );
  INV_X4 U3331 ( .A(n2727), .ZN(\u6/N14 ) );
  INV_X4 U3332 ( .A(N67), .ZN(n2728) );
  MUX2_X2 U3333 ( .A(n3111), .B(n2728), .S(n3012), .Z(n2729) );
  INV_X4 U3334 ( .A(n2729), .ZN(\u6/N13 ) );
  INV_X4 U3335 ( .A(n2833), .ZN(n2767) );
  NAND2_X2 U3336 ( .A1(n3143), .A2(n2767), .ZN(n2754) );
  NAND2_X2 U3337 ( .A1(\u2/N34 ), .A2(n2738), .ZN(n2734) );
  NOR2_X4 U3338 ( .A1(\u2/exp_ovf_d[1] ), .A2(n2767), .ZN(n2758) );
  AOI22_X2 U3339 ( .A1(n2759), .A2(n1689), .B1(\u2/exp_tmp3[4] ), .B2(n2758), 
        .ZN(n2733) );
  INV_X4 U3340 ( .A(n2757), .ZN(n2738) );
  NAND2_X2 U3341 ( .A1(\u2/N33 ), .A2(n2738), .ZN(n2740) );
  AOI22_X2 U3342 ( .A1(\u2/exp_tmp4[3] ), .A2(n2759), .B1(\u2/exp_tmp3[3] ), 
        .B2(n2758), .ZN(n2739) );
  NAND3_X4 U3343 ( .A1(n2741), .A2(n2740), .A3(n2739), .ZN(\u2/N43 ) );
  INV_X4 U3344 ( .A(\u2/N37 ), .ZN(n2742) );
  NAND2_X2 U3345 ( .A1(\u2/N32 ), .A2(n2738), .ZN(n2746) );
  AOI22_X2 U3346 ( .A1(\u2/exp_tmp4[2] ), .A2(n2759), .B1(\u2/exp_tmp3[2] ), 
        .B2(n2758), .ZN(n2745) );
  NAND3_X4 U3347 ( .A1(n2747), .A2(n2746), .A3(n2745), .ZN(\u2/N42 ) );
  NAND2_X2 U3348 ( .A1(\u2/N31 ), .A2(n2738), .ZN(n2751) );
  AOI22_X2 U3349 ( .A1(\u2/exp_tmp4[1] ), .A2(n2759), .B1(\u2/exp_tmp3[1] ), 
        .B2(n2758), .ZN(n2750) );
  NAND3_X4 U3350 ( .A1(n2752), .A2(n2751), .A3(n2750), .ZN(\u2/N41 ) );
  NAND2_X2 U3351 ( .A1(\u2/lt_130/A[0] ), .A2(n2738), .ZN(n2761) );
  AOI22_X2 U3352 ( .A1(\u2/exp_tmp4[0] ), .A2(n2759), .B1(n3142), .B2(n2758), 
        .ZN(n2760) );
  NAND3_X4 U3353 ( .A1(n2762), .A2(n2761), .A3(n2760), .ZN(\u2/N40 ) );
  MUX2_X2 U3354 ( .A(n3124), .B(n3133), .S(n1733), .Z(n2763) );
  NAND2_X2 U3355 ( .A1(n3129), .A2(n3012), .ZN(n2764) );
  OAI211_X2 U3356 ( .C1(n2766), .C2(n2765), .A(n1582), .B(n2764), .ZN(
        \u2/underflow_d [1]) );
  MUX2_X2 U3357 ( .A(n2768), .B(n3135), .S(n3124), .Z(\u2/N66 ) );
  INV_X4 U3358 ( .A(n2769), .ZN(n2779) );
  NAND2_X2 U3359 ( .A1(opb_r[11]), .A2(n1725), .ZN(n2782) );
  AOI21_X4 U3360 ( .B1(n2772), .B2(n2782), .A(n2771), .ZN(n2774) );
  OAI21_X4 U3361 ( .B1(n2784), .B2(n2774), .A(n2773), .ZN(n2777) );
  INV_X4 U3362 ( .A(n2780), .ZN(n2775) );
  NOR2_X4 U3363 ( .A1(n2775), .A2(n2779), .ZN(n2776) );
  OAI21_X4 U3364 ( .B1(n2777), .B2(n2778), .A(n2776), .ZN(n2790) );
  NAND2_X2 U3365 ( .A1(n2781), .A2(n2780), .ZN(n2785) );
  INV_X4 U3366 ( .A(n2782), .ZN(n2783) );
  NAND4_X2 U3367 ( .A1(\u1/N124 ), .A2(n3145), .A3(n2787), .A4(n2786), .ZN(
        n2792) );
  INV_X4 U3368 ( .A(n2815), .ZN(n2788) );
  AND2_X2 U3369 ( .A1(n2792), .A2(n2788), .ZN(\u1/N39 ) );
  MUX2_X2 U3370 ( .A(n1560), .B(n1543), .S(n1975), .Z(n2819) );
  AND2_X2 U3371 ( .A1(n2792), .A2(n2818), .ZN(\u1/N38 ) );
  MUX2_X2 U3372 ( .A(n1573), .B(n2799), .S(n1975), .Z(n2811) );
  INV_X4 U3373 ( .A(n2811), .ZN(n2800) );
  AND2_X2 U3374 ( .A1(n2792), .A2(n2800), .ZN(\u1/N37 ) );
  MUX2_X2 U3375 ( .A(n1725), .B(n3016), .S(n1975), .Z(n2807) );
  INV_X4 U3376 ( .A(n2807), .ZN(n2796) );
  AND2_X2 U3377 ( .A1(n2792), .A2(n2796), .ZN(\u1/N36 ) );
  NAND2_X2 U3378 ( .A1(n2790), .A2(n2789), .ZN(n2791) );
  MUX2_X2 U3379 ( .A(n1723), .B(n1726), .S(n1975), .Z(n2794) );
  INV_X4 U3380 ( .A(n2794), .ZN(n2832) );
  AND2_X2 U3381 ( .A1(n2792), .A2(n2832), .ZN(\u1/N35 ) );
  MUX2_X2 U3382 ( .A(\u3/N17 ), .B(\u3/N32 ), .S(n3084), .Z(n3284) );
  MUX2_X2 U3383 ( .A(\u3/N16 ), .B(\u3/N31 ), .S(n3084), .Z(n3285) );
  MUX2_X2 U3384 ( .A(\u3/N15 ), .B(\u3/N30 ), .S(n3084), .Z(n3286) );
  MUX2_X2 U3385 ( .A(\u3/N14 ), .B(\u3/N29 ), .S(n3084), .Z(n3287) );
  MUX2_X2 U3386 ( .A(\u3/N13 ), .B(\u3/N28 ), .S(n3084), .Z(n3288) );
  MUX2_X2 U3387 ( .A(\u3/N12 ), .B(\u3/N27 ), .S(n3084), .Z(n3289) );
  MUX2_X2 U3388 ( .A(\u3/N11 ), .B(\u3/N26 ), .S(n3084), .Z(n3290) );
  MUX2_X2 U3389 ( .A(\u3/N10 ), .B(\u3/N25 ), .S(n3084), .Z(n3291) );
  MUX2_X2 U3390 ( .A(\u3/N9 ), .B(\u3/N24 ), .S(n3084), .Z(n3292) );
  MUX2_X2 U3391 ( .A(\u3/N8 ), .B(\u3/N23 ), .S(n3084), .Z(n3293) );
  MUX2_X2 U3392 ( .A(\u3/N7 ), .B(\u3/N22 ), .S(n3084), .Z(n3294) );
  MUX2_X2 U3393 ( .A(\u3/N6 ), .B(\u3/N21 ), .S(n3084), .Z(n3295) );
  MUX2_X2 U3394 ( .A(\u3/N5 ), .B(\u3/N20 ), .S(n3084), .Z(n3296) );
  MUX2_X2 U3395 ( .A(\u3/N4 ), .B(\u3/N19 ), .S(n3084), .Z(n3297) );
  MUX2_X2 U3396 ( .A(\u3/N3 ), .B(\u3/N18 ), .S(n3084), .Z(n3298) );
  MUX2_X2 U3397 ( .A(n1731), .B(n3313), .S(n2793), .Z(n1521) );
  INV_X4 U3398 ( .A(n3110), .ZN(n2958) );
  MUX2_X2 U3399 ( .A(n2958), .B(fracta_mul[9]), .S(n2793), .Z(\u1/adj_op[9] )
         );
  INV_X4 U3400 ( .A(n3109), .ZN(n2911) );
  MUX2_X2 U3401 ( .A(n2911), .B(fracta_mul[8]), .S(n1975), .Z(n3303) );
  INV_X4 U3402 ( .A(n3108), .ZN(n2905) );
  MUX2_X2 U3403 ( .A(n2905), .B(fracta_mul[7]), .S(n1975), .Z(n3304) );
  INV_X4 U3404 ( .A(n3107), .ZN(n2844) );
  INV_X4 U3405 ( .A(n3117), .ZN(n2843) );
  MUX2_X2 U3406 ( .A(n2844), .B(n2843), .S(n1975), .Z(n3305) );
  INV_X4 U3407 ( .A(n3106), .ZN(n2841) );
  INV_X4 U3408 ( .A(n3116), .ZN(n2842) );
  MUX2_X2 U3409 ( .A(n2841), .B(n2842), .S(n1975), .Z(n3306) );
  MUX2_X2 U3410 ( .A(n2895), .B(n2896), .S(n1975), .Z(n3307) );
  INV_X4 U3411 ( .A(n3104), .ZN(n2888) );
  MUX2_X2 U3412 ( .A(n2888), .B(n2889), .S(n1975), .Z(n3308) );
  INV_X4 U3413 ( .A(n3103), .ZN(n2847) );
  INV_X4 U3414 ( .A(n3113), .ZN(n2848) );
  MUX2_X2 U3415 ( .A(n2847), .B(n2848), .S(n2924), .Z(n3309) );
  INV_X4 U3416 ( .A(n3102), .ZN(n2846) );
  MUX2_X2 U3417 ( .A(n2846), .B(n3014), .S(n2924), .Z(n3310) );
  INV_X4 U3418 ( .A(n3101), .ZN(n2852) );
  MUX2_X2 U3419 ( .A(n2852), .B(n3015), .S(n2924), .Z(n3311) );
  MUX2_X2 U3420 ( .A(n1726), .B(n1723), .S(n1975), .Z(n2831) );
  INV_X4 U3421 ( .A(n2831), .ZN(n2795) );
  OAI21_X4 U3422 ( .B1(n2795), .B2(n2833), .A(n2794), .ZN(n2809) );
  MUX2_X2 U3423 ( .A(n3016), .B(n1725), .S(n1975), .Z(n2808) );
  NOR2_X4 U3424 ( .A1(n2808), .A2(n2796), .ZN(n2798) );
  NAND2_X2 U3425 ( .A1(n2796), .A2(n2808), .ZN(n2797) );
  OAI21_X4 U3426 ( .B1(n1539), .B2(n2798), .A(n2797), .ZN(n2813) );
  INV_X4 U3427 ( .A(n2813), .ZN(n2803) );
  MUX2_X2 U3428 ( .A(n2799), .B(n1573), .S(n2924), .Z(n2812) );
  NOR2_X4 U3429 ( .A1(n2812), .A2(n2800), .ZN(n2802) );
  NAND2_X2 U3430 ( .A1(n2800), .A2(n2812), .ZN(n2801) );
  OAI21_X4 U3431 ( .B1(n2803), .B2(n2802), .A(n2801), .ZN(n2817) );
  MUX2_X2 U3432 ( .A(n1543), .B(n1560), .S(n2924), .Z(n2820) );
  INV_X4 U3433 ( .A(n2820), .ZN(n2804) );
  XNOR2_X2 U3434 ( .A(n2804), .B(n2819), .ZN(n2805) );
  XNOR2_X2 U3435 ( .A(n2806), .B(n2805), .ZN(n2828) );
  XNOR2_X2 U3436 ( .A(n2808), .B(n2807), .ZN(n2810) );
  XNOR2_X2 U3437 ( .A(n2810), .B(n2809), .ZN(n2830) );
  XNOR2_X2 U3438 ( .A(n2812), .B(n2811), .ZN(n2814) );
  XNOR2_X2 U3439 ( .A(n2813), .B(n2814), .ZN(n2829) );
  NOR3_X4 U3440 ( .A1(n2828), .A2(n2830), .A3(n2829), .ZN(n2827) );
  MUX2_X2 U3441 ( .A(opb_r[14]), .B(opa_r[14]), .S(n2924), .Z(n2816) );
  NOR2_X4 U3442 ( .A1(n2816), .A2(n2815), .ZN(n2824) );
  INV_X4 U3443 ( .A(n2819), .ZN(n2818) );
  NAND2_X2 U3444 ( .A1(n2818), .A2(n2820), .ZN(n2821) );
  XNOR2_X2 U3445 ( .A(n2823), .B(n2824), .ZN(n2826) );
  INV_X4 U3446 ( .A(n2836), .ZN(n2825) );
  OAI21_X4 U3447 ( .B1(n2827), .B2(n2826), .A(n2825), .ZN(n2837) );
  OAI21_X4 U3448 ( .B1(n2836), .B2(n2828), .A(n2837), .ZN(n3302) );
  OAI21_X4 U3449 ( .B1(n2836), .B2(n2830), .A(n2837), .ZN(n3300) );
  XNOR2_X2 U3450 ( .A(n2832), .B(n2831), .ZN(n2834) );
  XNOR2_X2 U3451 ( .A(n2834), .B(n2833), .ZN(n2835) );
  MUX2_X2 U3452 ( .A(\u1/adj_op_out_sft[13] ), .B(n1731), .S(n1976), .Z(n2929)
         );
  INV_X4 U3453 ( .A(n2929), .ZN(n2839) );
  NAND2_X2 U3454 ( .A1(n2839), .A2(n2928), .ZN(\u1/fracta_s [13]) );
  MUX2_X2 U3455 ( .A(\u1/adj_op_out_sft[12] ), .B(n2958), .S(n1976), .Z(n2931)
         );
  MUX2_X2 U3456 ( .A(fracta_mul[9]), .B(\u1/adj_op_out_sft[12] ), .S(n1976), 
        .Z(n2932) );
  INV_X4 U3457 ( .A(n2932), .ZN(n2840) );
  NAND2_X2 U3458 ( .A1(n2840), .A2(n2931), .ZN(n2919) );
  MUX2_X2 U3459 ( .A(\u1/adj_op_out_sft[8] ), .B(n2841), .S(n1976), .Z(n2939)
         );
  MUX2_X2 U3460 ( .A(n2842), .B(\u1/adj_op_out_sft[8] ), .S(n1976), .Z(n2940)
         );
  INV_X4 U3461 ( .A(n2940), .ZN(n2845) );
  MUX2_X2 U3462 ( .A(n2843), .B(\u1/adj_op_out_sft[9] ), .S(n1976), .Z(n2938)
         );
  MUX2_X2 U3463 ( .A(\u1/adj_op_out_sft[9] ), .B(n2844), .S(n1976), .Z(n2937)
         );
  AOI22_X2 U3464 ( .A1(n2939), .A2(n2845), .B1(n2904), .B2(n2937), .ZN(n2910)
         );
  MUX2_X2 U3465 ( .A(n3014), .B(\u1/adj_op_out_sft[4] ), .S(n1976), .Z(n2948)
         );
  MUX2_X2 U3466 ( .A(\u1/adj_op_out_sft[5] ), .B(n2847), .S(n1976), .Z(n2945)
         );
  INV_X4 U3467 ( .A(n2945), .ZN(n2849) );
  MUX2_X2 U3468 ( .A(fracta_mul[2]), .B(\u1/adj_op_out_sft[5] ), .S(n1976), 
        .Z(n2946) );
  NOR2_X4 U3469 ( .A1(n2849), .A2(n2946), .ZN(n2850) );
  NOR2_X4 U3470 ( .A1(n2851), .A2(n2850), .ZN(n2894) );
  MUX2_X2 U3471 ( .A(\u1/adj_op_out_sft[3] ), .B(n2852), .S(n1976), .Z(n2949)
         );
  INV_X4 U3472 ( .A(n2949), .ZN(n2883) );
  MUX2_X2 U3473 ( .A(fracta_mul[0]), .B(\u1/adj_op_out_sft[3] ), .S(n1976), 
        .Z(n2950) );
  INV_X4 U3474 ( .A(n3311), .ZN(n2872) );
  INV_X4 U3475 ( .A(n3310), .ZN(n2854) );
  INV_X4 U3476 ( .A(n3309), .ZN(n2853) );
  INV_X4 U3477 ( .A(n2869), .ZN(n2857) );
  INV_X4 U3478 ( .A(n3308), .ZN(n2856) );
  INV_X4 U3479 ( .A(n3307), .ZN(n2855) );
  INV_X4 U3480 ( .A(n2864), .ZN(n2859) );
  INV_X4 U3481 ( .A(n3306), .ZN(n2862) );
  INV_X4 U3482 ( .A(n3305), .ZN(n2858) );
  INV_X4 U3483 ( .A(n2866), .ZN(n2861) );
  INV_X4 U3484 ( .A(n3304), .ZN(n2860) );
  NAND2_X2 U3485 ( .A1(n2861), .A2(n2860), .ZN(n2871) );
  INV_X4 U3486 ( .A(n2871), .ZN(n2863) );
  INV_X4 U3487 ( .A(n3302), .ZN(n2874) );
  AOI211_X4 U3488 ( .C1(\u1/exp_diff_sft[0] ), .C2(\u1/adj_op[9] ), .A(n3303), 
        .B(n2871), .ZN(n2873) );
  OAI221_X2 U3489 ( .B1(n2854), .B2(n1719), .C1(n2874), .C2(n2873), .A(n2872), 
        .ZN(n2877) );
  MUX2_X2 U3490 ( .A(n2880), .B(n2879), .S(n3301), .Z(n2881) );
  NOR2_X4 U3491 ( .A1(\u1/adj_op_out_sft[0] ), .A2(n2881), .ZN(n2927) );
  INV_X4 U3492 ( .A(n2927), .ZN(n2882) );
  NAND2_X2 U3493 ( .A1(n1720), .A2(n2948), .ZN(n2885) );
  NAND2_X2 U3494 ( .A1(n2883), .A2(n2950), .ZN(n2884) );
  INV_X4 U3495 ( .A(n2946), .ZN(n2887) );
  MUX2_X2 U3496 ( .A(\u1/adj_op_out_sft[6] ), .B(n2888), .S(n1976), .Z(n2943)
         );
  MUX2_X2 U3497 ( .A(n2889), .B(\u1/adj_op_out_sft[6] ), .S(n1976), .Z(n2944)
         );
  INV_X4 U3498 ( .A(n2944), .ZN(n2890) );
  MUX2_X2 U3499 ( .A(\u1/adj_op_out_sft[7] ), .B(n2895), .S(n1976), .Z(n2941)
         );
  INV_X4 U3500 ( .A(n2941), .ZN(n2899) );
  MUX2_X2 U3501 ( .A(n2896), .B(\u1/adj_op_out_sft[7] ), .S(n1976), .Z(n2942)
         );
  INV_X4 U3502 ( .A(n2943), .ZN(n2897) );
  OAI22_X2 U3503 ( .A1(n2899), .A2(n2942), .B1(n2944), .B2(n2897), .ZN(n2902)
         );
  INV_X4 U3504 ( .A(n2939), .ZN(n2898) );
  NAND2_X2 U3505 ( .A1(n2940), .A2(n2898), .ZN(n2901) );
  NAND2_X2 U3506 ( .A1(n2899), .A2(n2942), .ZN(n2900) );
  MUX2_X2 U3507 ( .A(\u1/adj_op_out_sft[10] ), .B(n2905), .S(n1976), .Z(n2935)
         );
  MUX2_X2 U3508 ( .A(fracta_mul[7]), .B(\u1/adj_op_out_sft[10] ), .S(n1976), 
        .Z(n2936) );
  INV_X4 U3509 ( .A(n2936), .ZN(n2906) );
  NOR2_X4 U3510 ( .A1(n2935), .A2(n2906), .ZN(n2907) );
  AOI211_X4 U3511 ( .C1(n2909), .C2(n2910), .A(n2908), .B(n2907), .ZN(n2916)
         );
  MUX2_X2 U3512 ( .A(fracta_mul[8]), .B(\u1/adj_op_out_sft[11] ), .S(n1976), 
        .Z(n2934) );
  MUX2_X2 U3513 ( .A(\u1/adj_op_out_sft[11] ), .B(n2911), .S(n1976), .Z(n2933)
         );
  INV_X4 U3514 ( .A(n2933), .ZN(n2913) );
  INV_X4 U3515 ( .A(n2935), .ZN(n2912) );
  OAI22_X2 U3516 ( .A1(n2934), .A2(n2913), .B1(n2936), .B2(n2912), .ZN(n2915)
         );
  NAND2_X2 U3517 ( .A1(n2934), .A2(n2913), .ZN(n2914) );
  OAI21_X4 U3518 ( .B1(n2916), .B2(n2915), .A(n2914), .ZN(n2918) );
  AOI21_X4 U3519 ( .B1(n2918), .B2(n2919), .A(n2917), .ZN(n2922) );
  INV_X4 U3520 ( .A(n2931), .ZN(n2920) );
  NAND2_X2 U3521 ( .A1(n2920), .A2(n2932), .ZN(n2921) );
  AOI21_X4 U3522 ( .B1(n2922), .B2(n2921), .A(n1649), .ZN(n2954) );
  MUX2_X2 U3523 ( .A(n2931), .B(n2932), .S(n1979), .Z(\u1/fracta_s [12]) );
  MUX2_X2 U3524 ( .A(n2933), .B(n2934), .S(n1979), .Z(\u1/fracta_s [11]) );
  MUX2_X2 U3525 ( .A(n2935), .B(n2936), .S(n1979), .Z(\u1/fracta_s [10]) );
  MUX2_X2 U3526 ( .A(n2937), .B(n2938), .S(n1979), .Z(\u1/fracta_s [9]) );
  MUX2_X2 U3527 ( .A(n2939), .B(n2940), .S(n1979), .Z(\u1/fracta_s [8]) );
  MUX2_X2 U3528 ( .A(n2941), .B(n2942), .S(n1979), .Z(\u1/fracta_s [7]) );
  MUX2_X2 U3529 ( .A(n2943), .B(n2944), .S(n1978), .Z(\u1/fracta_s [6]) );
  MUX2_X2 U3530 ( .A(n2945), .B(n2946), .S(n1978), .Z(\u1/fracta_s [5]) );
  MUX2_X2 U3531 ( .A(n2947), .B(n2948), .S(n1979), .Z(\u1/fracta_s [4]) );
  MUX2_X2 U3532 ( .A(n2949), .B(n2950), .S(n1979), .Z(\u1/fracta_s [3]) );
  MUX2_X2 U3533 ( .A(n1563), .B(n1590), .S(n1979), .Z(\u1/fracta_s [2]) );
  INV_X4 U3534 ( .A(n2923), .ZN(n2951) );
  MUX2_X2 U3535 ( .A(n2951), .B(n1645), .S(n1978), .Z(\u1/fracta_s [1]) );
  INV_X4 U3536 ( .A(n2925), .ZN(n2952) );
  MUX2_X2 U3537 ( .A(n2952), .B(n2953), .S(n1978), .Z(\u1/fracta_s [0]) );
  INV_X4 U3538 ( .A(n2928), .ZN(n2930) );
  MUX2_X2 U3539 ( .A(n2930), .B(n2929), .S(n1978), .Z(\u1/fractb_s [13]) );
  MUX2_X2 U3540 ( .A(n2932), .B(n2931), .S(n1979), .Z(\u1/fractb_s [12]) );
  MUX2_X2 U3541 ( .A(n2934), .B(n2933), .S(n1978), .Z(\u1/fractb_s [11]) );
  MUX2_X2 U3542 ( .A(n2936), .B(n2935), .S(n1978), .Z(\u1/fractb_s [10]) );
  MUX2_X2 U3543 ( .A(n2938), .B(n2937), .S(n1978), .Z(\u1/fractb_s [9]) );
  MUX2_X2 U3544 ( .A(n2940), .B(n2939), .S(n1978), .Z(\u1/fractb_s [8]) );
  MUX2_X2 U3545 ( .A(n2942), .B(n2941), .S(n1978), .Z(\u1/fractb_s [7]) );
  MUX2_X2 U3546 ( .A(n2944), .B(n2943), .S(n1978), .Z(\u1/fractb_s [6]) );
  MUX2_X2 U3547 ( .A(n2946), .B(n2945), .S(n1978), .Z(\u1/fractb_s [5]) );
  MUX2_X2 U3548 ( .A(n2948), .B(n2947), .S(n1978), .Z(\u1/fractb_s [4]) );
  MUX2_X2 U3549 ( .A(n2950), .B(n2949), .S(n1978), .Z(\u1/fractb_s [3]) );
  MUX2_X2 U3550 ( .A(n1590), .B(n1563), .S(n1978), .Z(\u1/fractb_s [2]) );
  MUX2_X2 U3551 ( .A(n1645), .B(n2951), .S(n1978), .Z(\u1/fractb_s [1]) );
  MUX2_X2 U3552 ( .A(n2953), .B(n2952), .S(n1978), .Z(\u1/fractb_s [0]) );
  XNOR2_X2 U3553 ( .A(n3317), .B(opb_r[15]), .ZN(n2955) );
  MUX2_X2 U3554 ( .A(n2955), .B(opa_r[15]), .S(n1978), .Z(\u1/sign_d ) );
  INV_X4 U3555 ( .A(n2956), .ZN(n2957) );
  INV_X4 U3556 ( .A(n3158), .ZN(n3312) );
  INV_X4 U3557 ( .A(n3157), .ZN(n3315) );
  OAI22_X2 U3558 ( .A1(net85778), .A2(net83361), .B1(net83438), .B2(net83439), 
        .ZN(n2960) );
  INV_X4 U3559 ( .A(net83427), .ZN(net15944) );
  XNOR2_X2 U3560 ( .A(net83407), .B(n2964), .ZN(n2966) );
  XNOR2_X2 U3561 ( .A(n2966), .B(n2965), .ZN(n2967) );
  AOI21_X4 U3562 ( .B1(net15944), .B2(n2967), .A(net83423), .ZN(n851) );
  INV_X4 U3563 ( .A(n2968), .ZN(n2969) );
  FA_X1 U3564 ( .A(n1592), .B(n2969), .CI(net89964), .S(\u4/div_exp3[1] ) );
  INV_X4 U3565 ( .A(n3010), .ZN(n3009) );
  INV_X4 U3566 ( .A(n2970), .ZN(n2973) );
  INV_X4 U3567 ( .A(n2974), .ZN(n2986) );
  NAND2_X2 U3568 ( .A1(\u4/sub_409/net10540 ), .A2(div_opa_ldz_r2[3]), .ZN(
        n2975) );
  XNOR2_X2 U3569 ( .A(net11555), .B(n2977), .ZN(n2980) );
  NAND2_X2 U3570 ( .A1(net83364), .A2(n2978), .ZN(n2979) );
  OAI221_X2 U3571 ( .B1(n2980), .B2(n2989), .C1(net83361), .C2(n1688), .A(
        n2979), .ZN(n2984) );
  INV_X4 U3572 ( .A(n2981), .ZN(n2982) );
  XNOR2_X2 U3573 ( .A(\u4/sub_409/net10540 ), .B(div_opa_ldz_r2[3]), .ZN(n2985) );
  XNOR2_X2 U3574 ( .A(n2986), .B(n2985), .ZN(n2990) );
  NAND2_X2 U3575 ( .A1(net83364), .A2(n2987), .ZN(n2988) );
  OAI221_X2 U3576 ( .B1(n2990), .B2(n2989), .C1(net83361), .C2(n1687), .A(
        n2988), .ZN(n2994) );
  AND2_X1 U3577 ( .A1(net83968), .A2(\u4/add_407/carry [3]), .ZN(
        \u4/add_407/carry [4]) );
  XOR2_X1 U3578 ( .A(\u2/gt_140/B[5] ), .B(\u2/add_111/carry[5] ), .Z(\u2/N23 ) );
  XOR2_X1 U3579 ( .A(\u2/exp_tmp4[4] ), .B(\u2/add_111/carry[4] ), .Z(\u2/N22 ) );
  XNOR2_X1 U3580 ( .A(\u2/add_111/carry[3] ), .B(\u2/lt_130/A[3] ), .ZN(
        \u2/N21 ) );
  OR2_X1 U3581 ( .A1(\u2/lt_130/A[2] ), .A2(\u2/add_111/carry[2] ), .ZN(
        \u2/add_111/carry[3] ) );
  XNOR2_X1 U3582 ( .A(\u2/add_111/carry[2] ), .B(\u2/lt_130/A[2] ), .ZN(
        \u2/N20 ) );
  OR2_X1 U3583 ( .A1(\u2/lt_130/A[1] ), .A2(\u2/lt_130/A[0] ), .ZN(
        \u2/add_111/carry[2] ) );
  XNOR2_X1 U3584 ( .A(\u2/lt_130/A[0] ), .B(\u2/lt_130/A[1] ), .ZN(\u2/N19 )
         );
  XNOR2_X1 U3585 ( .A(\u2/gt_140/B[5] ), .B(\u2/sub_111/carry[5] ), .ZN(
        \u2/N29 ) );
  XNOR2_X1 U3586 ( .A(\u2/sub_111/carry[4] ), .B(\u2/exp_tmp4[4] ), .ZN(
        \u2/N28 ) );
  XOR2_X1 U3587 ( .A(\u2/lt_130/A[3] ), .B(\u2/sub_111/carry[3] ), .Z(\u2/N27 ) );
  AND2_X1 U3588 ( .A1(\u2/sub_111/carry[2] ), .A2(\u2/lt_130/A[2] ), .ZN(
        \u2/sub_111/carry[3] ) );
  XOR2_X1 U3589 ( .A(\u2/lt_130/A[2] ), .B(\u2/sub_111/carry[2] ), .Z(\u2/N26 ) );
  AND2_X1 U3590 ( .A1(\u2/lt_130/A[0] ), .A2(\u2/lt_130/A[1] ), .ZN(
        \u2/sub_111/carry[2] ) );
  XOR2_X1 U3591 ( .A(\u2/lt_130/A[1] ), .B(\u2/lt_130/A[0] ), .Z(\u2/N25 ) );
  XOR2_X1 U3592 ( .A(opb_r[10]), .B(opa_r[10]), .Z(\u2/N12 ) );
  XNOR2_X1 U3593 ( .A(n1726), .B(opa_r[10]), .ZN(\u2/N6 ) );
  XOR2_X1 U3594 ( .A(n1635), .B(\sub_435_3/carry [20]), .Z(N151) );
  AND2_X1 U3595 ( .A1(\sub_435_3/carry [19]), .A2(n1636), .ZN(
        \sub_435_3/carry [20]) );
  XOR2_X1 U3596 ( .A(n1636), .B(\sub_435_3/carry [19]), .Z(N150) );
  AND2_X1 U3597 ( .A1(\sub_435_3/carry [18]), .A2(n1637), .ZN(
        \sub_435_3/carry [19]) );
  AND2_X1 U3598 ( .A1(\sub_435_3/carry [17]), .A2(n1672), .ZN(
        \sub_435_3/carry [18]) );
  AND2_X1 U3599 ( .A1(\sub_435_3/carry [16]), .A2(n1673), .ZN(
        \sub_435_3/carry [17]) );
  AND2_X1 U3600 ( .A1(\sub_435_3/carry [15]), .A2(n1624), .ZN(
        \sub_435_3/carry [16]) );
  AND2_X1 U3601 ( .A1(\sub_435_3/carry [14]), .A2(n1625), .ZN(
        \sub_435_3/carry [15]) );
  AND2_X1 U3602 ( .A1(\sub_435_3/carry [13]), .A2(n1626), .ZN(
        \sub_435_3/carry [14]) );
  AND2_X1 U3603 ( .A1(\sub_435_3/carry [12]), .A2(n1627), .ZN(
        \sub_435_3/carry [13]) );
  AND2_X1 U3604 ( .A1(\sub_435_3/carry [11]), .A2(n1678), .ZN(
        \sub_435_3/carry [12]) );
  AND2_X1 U3605 ( .A1(\sub_435_3/carry [10]), .A2(n1679), .ZN(
        \sub_435_3/carry [11]) );
  XOR2_X1 U3606 ( .A(n1679), .B(\sub_435_3/carry [10]), .Z(N141) );
  AND2_X1 U3607 ( .A1(\sub_435_3/carry [9]), .A2(n1674), .ZN(
        \sub_435_3/carry [10]) );
  XOR2_X1 U3608 ( .A(n1674), .B(\sub_435_3/carry [9]), .Z(N140) );
  AND2_X1 U3609 ( .A1(\sub_435_3/carry [8]), .A2(n1675), .ZN(
        \sub_435_3/carry [9]) );
  XOR2_X1 U3610 ( .A(n1675), .B(\sub_435_3/carry [8]), .Z(N139) );
  AND2_X1 U3611 ( .A1(n1680), .A2(n1676), .ZN(\sub_435_3/carry [8]) );
  XOR2_X1 U3612 ( .A(n1676), .B(n1680), .Z(N138) );
  XOR2_X1 U3613 ( .A(n1558), .B(\sub_435_b0/carry [10]), .Z(N116) );
  AND2_X1 U3614 ( .A1(\sub_435_b0/carry [9]), .A2(n1624), .ZN(
        \sub_435_b0/carry [10]) );
  XOR2_X1 U3615 ( .A(n1624), .B(\sub_435_b0/carry [9]), .Z(N115) );
  AND2_X1 U3616 ( .A1(\sub_435_b0/carry [8]), .A2(n1625), .ZN(
        \sub_435_b0/carry [9]) );
  XOR2_X1 U3617 ( .A(n1625), .B(\sub_435_b0/carry [8]), .Z(N114) );
  AND2_X1 U3618 ( .A1(\sub_435_b0/carry [7]), .A2(n1626), .ZN(
        \sub_435_b0/carry [8]) );
  XOR2_X1 U3619 ( .A(n1626), .B(\sub_435_b0/carry [7]), .Z(N113) );
  AND2_X1 U3620 ( .A1(\sub_435_b0/carry [6]), .A2(n1627), .ZN(
        \sub_435_b0/carry [7]) );
  XOR2_X1 U3621 ( .A(n1627), .B(\sub_435_b0/carry [6]), .Z(N112) );
  AND2_X1 U3622 ( .A1(\sub_435_b0/carry [5]), .A2(n1678), .ZN(
        \sub_435_b0/carry [6]) );
  XOR2_X1 U3623 ( .A(n1678), .B(\sub_435_b0/carry [5]), .Z(N111) );
  AND2_X1 U3624 ( .A1(\sub_435_b0/carry [4]), .A2(n1679), .ZN(
        \sub_435_b0/carry [5]) );
  XOR2_X1 U3625 ( .A(n1679), .B(\sub_435_b0/carry [4]), .Z(N110) );
  AND2_X1 U3626 ( .A1(\sub_435_b0/carry [3]), .A2(n1674), .ZN(
        \sub_435_b0/carry [4]) );
  AND2_X1 U3627 ( .A1(\sub_435_b0/carry [2]), .A2(n1675), .ZN(
        \sub_435_b0/carry [3]) );
  AND2_X1 U3628 ( .A1(n1680), .A2(n1676), .ZN(\sub_435_b0/carry [2]) );
  INV_X4 U3629 ( .A(\u2/sub_110/carry [5]), .ZN(\u2/N11 ) );
  XOR2_X1 U3630 ( .A(\u2/add_113/carry [4]), .B(\u2/add_113/A[4] ), .Z(
        \u2/exp_tmp3[4] ) );
  INV_X4 U3631 ( .A(\u2/lt_130/A[0] ), .ZN(\u2/exp_tmp4[0] ) );
  INV_X4 U3632 ( .A(\u2/lt_130/A[1] ), .ZN(\u2/exp_tmp4[1] ) );
  INV_X4 U3633 ( .A(\u2/lt_130/A[2] ), .ZN(\u2/exp_tmp4[2] ) );
  XOR2_X1 U3634 ( .A(\u2/add_115/carry [4]), .B(n1689), .Z(\u2/N34 ) );
  NOR2_X1 U3635 ( .A1(\u2/exp_tmp4[1] ), .A2(\u2/exp_tmp4[0] ), .ZN(n3019) );
  AOI21_X1 U3636 ( .B1(\u2/exp_tmp4[0] ), .B2(\u2/exp_tmp4[1] ), .A(n3019), 
        .ZN(n3018) );
  NAND2_X1 U3637 ( .A1(n3019), .A2(\u2/lt_130/A[2] ), .ZN(n3020) );
  OAI21_X1 U3638 ( .B1(n3019), .B2(\u2/lt_130/A[2] ), .A(n3020), .ZN(\u2/N37 )
         );
  NOR2_X1 U3639 ( .A1(\u2/exp_tmp4[3] ), .A2(n3020), .ZN(n3021) );
  INV_X4 U3640 ( .A(net83968), .ZN(\u4/sub_409/net10540 ) );
  OAI22_X1 U3641 ( .A1(fracta_mul[1]), .A2(n3022), .B1(n3022), .B2(n3046), 
        .ZN(n3024) );
  NAND2_X1 U3642 ( .A1(fracta_mul[7]), .A2(n3108), .ZN(n3025) );
  NAND2_X1 U3643 ( .A1(fracta_mul[5]), .A2(n3106), .ZN(n3033) );
  NAND2_X1 U3644 ( .A1(fracta_mul[6]), .A2(n3107), .ZN(n3034) );
  AND2_X1 U3645 ( .A1(n3033), .A2(n3034), .ZN(n3023) );
  OR2_X1 U3646 ( .A1(n3119), .A2(\u6/N8 ), .ZN(n3026) );
  NAND4_X1 U3647 ( .A1(n3024), .A2(n3025), .A3(n3023), .A4(n3026), .ZN(n3044)
         );
  NAND2_X1 U3648 ( .A1(fracta_mul[9]), .A2(n3110), .ZN(n3040) );
  AND2_X1 U3649 ( .A1(n3026), .A2(n3025), .ZN(n3037) );
  NAND2_X1 U3650 ( .A1(fracta_mul[4]), .A2(n3105), .ZN(n3042) );
  NAND2_X1 U3651 ( .A1(fracta_mul[3]), .A2(n3104), .ZN(n3041) );
  NOR2_X1 U3652 ( .A1(n3045), .A2(fracta_mul[0]), .ZN(n3028) );
  OAI21_X1 U3653 ( .B1(fracta_mul[1]), .B2(n3048), .A(n3046), .ZN(n3027) );
  NAND2_X1 U3654 ( .A1(fracta_mul[2]), .A2(n3047), .ZN(n3039) );
  OAI211_X1 U3655 ( .C1(n3028), .C2(n3049), .A(n3027), .B(n3039), .ZN(n3029)
         );
  OAI221_X1 U3656 ( .B1(fracta_mul[2]), .B2(n3047), .C1(fracta_mul[3]), .C2(
        n3104), .A(n3029), .ZN(n3030) );
  NAND3_X1 U3657 ( .A1(n3042), .A2(n3041), .A3(n3030), .ZN(n3031) );
  OAI221_X1 U3658 ( .B1(fracta_mul[4]), .B2(n3105), .C1(fracta_mul[5]), .C2(
        n3106), .A(n3031), .ZN(n3032) );
  NAND3_X1 U3659 ( .A1(n3034), .A2(n3033), .A3(n3032), .ZN(n3035) );
  OAI221_X1 U3660 ( .B1(fracta_mul[6]), .B2(n3107), .C1(fracta_mul[7]), .C2(
        n3108), .A(n3035), .ZN(n3036) );
  AOI22_X1 U3661 ( .A1(\u6/N8 ), .A2(n3119), .B1(n3037), .B2(n3036), .ZN(n3038) );
  OAI22_X1 U3662 ( .A1(fracta_mul[9]), .A2(n3110), .B1(n3052), .B2(n3038), 
        .ZN(\u1/N123 ) );
  NAND3_X1 U3663 ( .A1(n3040), .A2(n3053), .A3(n3039), .ZN(n3043) );
  NOR4_X1 U3664 ( .A1(n3044), .A2(n3043), .A3(n3050), .A4(n3051), .ZN(
        \u1/N124 ) );
  INV_X4 U3665 ( .A(\u6/N0 ), .ZN(n3045) );
  INV_X4 U3666 ( .A(\u6/N1 ), .ZN(n3046) );
  INV_X4 U3667 ( .A(\u6/N2 ), .ZN(n3047) );
  INV_X4 U3668 ( .A(n3028), .ZN(n3048) );
  INV_X4 U3669 ( .A(n3041), .ZN(n3050) );
  INV_X4 U3670 ( .A(n3042), .ZN(n3051) );
  INV_X4 U3671 ( .A(n3040), .ZN(n3052) );
  INV_X4 U3672 ( .A(\u1/N123 ), .ZN(n3053) );
  MUX2_X1 U3673 ( .A(n3122), .B(n3123), .S(n3124), .Z(n3121) );
  NAND4_X1 U3674 ( .A1(\u2/N15 ), .A2(\u2/N14 ), .A3(n3125), .A4(\u2/N13 ), 
        .ZN(n3123) );
  NOR2_X1 U3675 ( .A1(\u2/N16 ), .A2(n3126), .ZN(n3125) );
  INV_X1 U3676 ( .A(\u2/N12 ), .ZN(n3126) );
  NAND4_X1 U3677 ( .A1(\u2/N9 ), .A2(\u2/N8 ), .A3(n3127), .A4(\u2/N7 ), .ZN(
        n3122) );
  NOR2_X1 U3678 ( .A1(\u2/N10 ), .A2(n3128), .ZN(n3127) );
  INV_X1 U3679 ( .A(\u2/N6 ), .ZN(n3128) );
  NAND2_X1 U3680 ( .A1(n3134), .A2(n3124), .ZN(n3133) );
  NOR2_X1 U3681 ( .A1(n1686), .A2(n1569), .ZN(\u2/N73 ) );
  NOR2_X1 U3682 ( .A1(n3131), .A2(n3132), .ZN(n3135) );
  INV_X1 U3683 ( .A(\u2/gt_140/B[5] ), .ZN(n3132) );
  MUX2_X1 U3684 ( .A(\u2/N17 ), .B(\u2/N11 ), .S(n3136), .Z(\u2/gt_140/B[5] )
         );
  NOR2_X1 U3685 ( .A1(n1689), .A2(n3137), .ZN(n3131) );
  AND4_X1 U3686 ( .A1(\u2/lt_130/A[3] ), .A2(\u2/lt_130/A[2] ), .A3(
        \u2/lt_130/A[0] ), .A4(\u2/lt_130/A[1] ), .ZN(n3137) );
  MUX2_X1 U3687 ( .A(\u2/N13 ), .B(\u2/N7 ), .S(n3136), .Z(\u2/lt_130/A[1] )
         );
  MUX2_X1 U3688 ( .A(\u2/N12 ), .B(\u2/N6 ), .S(n3136), .Z(\u2/lt_130/A[0] )
         );
  MUX2_X1 U3689 ( .A(\u2/N14 ), .B(\u2/N8 ), .S(n3136), .Z(\u2/lt_130/A[2] )
         );
  INV_X1 U3690 ( .A(\u2/add_113/A[3] ), .ZN(n3139) );
  INV_X1 U3691 ( .A(\u2/add_113/A[2] ), .ZN(n3140) );
  INV_X1 U3692 ( .A(\u2/add_113/A[1] ), .ZN(n3141) );
  INV_X1 U3693 ( .A(\u2/add_113/A[4] ), .ZN(n3138) );
  INV_X1 U3694 ( .A(\u2/add_113/A[0] ), .ZN(n3142) );
  OAI21_X1 U3695 ( .B1(n3146), .B2(n1671), .A(n3147), .ZN(\u1/N133 ) );
  OAI21_X1 U3696 ( .B1(n3148), .B2(n1684), .A(\u1/signa_r ), .ZN(n3147) );
  NOR3_X1 U3697 ( .A1(n1681), .A2(\u1/fracta_lt_fractb ), .A3(
        \u1/fracta_eq_fractb ), .ZN(n3148) );
  AOI21_X1 U3698 ( .B1(opb_nan), .B2(n3149), .A(\u1/signa_r ), .ZN(n3146) );
  OAI21_X1 U3699 ( .B1(\u1/fracta_eq_fractb ), .B2(n1683), .A(opa_nan), .ZN(
        n3149) );
  OAI22_X1 U3700 ( .A1(n1682), .A2(n3150), .B1(n3151), .B2(n3152), .ZN(
        \u1/N122 ) );
  XNOR2_X1 U3701 ( .A(n1671), .B(\u1/add_r ), .ZN(n3152) );
  NOR2_X1 U3702 ( .A1(n3153), .A2(\u1/signa_r ), .ZN(n3151) );
  NAND2_X1 U3703 ( .A1(n3154), .A2(n3155), .ZN(\u0/N7 ) );
  NOR2_X1 U3704 ( .A1(n3155), .A2(n3154), .ZN(\u0/N6 ) );
  NOR2_X1 U3705 ( .A1(n3093), .A2(n3095), .ZN(\u0/N17 ) );
  NOR2_X1 U3706 ( .A1(n3092), .A2(n3094), .ZN(\u0/N16 ) );
  NOR2_X1 U3707 ( .A1(n3316), .A2(n3157), .ZN(\u0/N11 ) );
  NOR2_X1 U3708 ( .A1(n3314), .A2(n3158), .ZN(\u0/N10 ) );
  OAI22_X1 U3709 ( .A1(n3159), .A2(n1674), .B1(n3160), .B2(n1564), .ZN(n3281)
         );
  OAI22_X1 U3710 ( .A1(n3159), .A2(n1675), .B1(n3160), .B2(n1565), .ZN(n3282)
         );
  OAI22_X1 U3711 ( .A1(n3159), .A2(n1676), .B1(n3160), .B2(n1559), .ZN(n3283)
         );
  MUX2_X1 U3712 ( .A(\u2/N22 ), .B(\u2/N28 ), .S(n3124), .Z(\u2/add_113/A[4] )
         );
  MUX2_X1 U3713 ( .A(\u2/N21 ), .B(\u2/N27 ), .S(n3124), .Z(\u2/add_113/A[3] )
         );
  MUX2_X1 U3714 ( .A(\u2/N26 ), .B(\u2/N20 ), .S(n3136), .Z(\u2/add_113/A[2] )
         );
  MUX2_X1 U3715 ( .A(\u2/N19 ), .B(\u2/N25 ), .S(n3124), .Z(\u2/add_113/A[1] )
         );
  MUX2_X1 U3716 ( .A(\u2/exp_tmp4[0] ), .B(\u2/exp_tmp4[0] ), .S(n3136), .Z(
        \u2/add_113/A[0] ) );
  INV_X1 U3717 ( .A(n3145), .ZN(n3299) );
  XOR2_X1 U3718 ( .A(fpu_op_r1[0]), .B(\u2/sign_d ), .Z(n3145) );
  XNOR2_X1 U3719 ( .A(n1569), .B(opb_r[15]), .ZN(\u2/sign_d ) );
  INV_X1 U3720 ( .A(n3129), .ZN(n3314) );
  NAND2_X1 U3721 ( .A1(n3120), .A2(n3156), .ZN(n3129) );
  AND4_X1 U3722 ( .A1(n3118), .A2(n3113), .A3(n3119), .A4(n3161), .ZN(n3156)
         );
  NOR3_X1 U3723 ( .A1(n3014), .A2(n3162), .A3(n3015), .ZN(n3161) );
  INV_X1 U3724 ( .A(n3130), .ZN(n3316) );
  OAI22_X1 U3725 ( .A1(n3159), .A2(n1680), .B1(n3160), .B2(n1680), .ZN(n3318)
         );
  OAI22_X1 U3726 ( .A1(n1677), .A2(n3090), .B1(n1591), .B2(n3088), .ZN(n3320)
         );
  OAI22_X1 U3727 ( .A1(n1677), .A2(n3089), .B1(n1591), .B2(n3087), .ZN(n3321)
         );
  INV_X1 U3728 ( .A(n3154), .ZN(n3322) );
  NAND2_X1 U3729 ( .A1(\u0/infb_f_r ), .A2(\u0/expb_ff ), .ZN(n3154) );
  INV_X1 U3730 ( .A(n3155), .ZN(n3323) );
  NAND2_X1 U3731 ( .A1(\u0/infa_f_r ), .A2(\u0/expa_ff ), .ZN(n3155) );
  OAI222_X1 U3732 ( .A1(n3080), .A2(n3163), .B1(n3067), .B2(n3164), .C1(n3165), 
        .C2(n1636), .ZN(N99) );
  OAI222_X1 U3733 ( .A1(n3081), .A2(n3163), .B1(n3166), .B2(n1637), .C1(n3098), 
        .C2(n3068), .ZN(N98) );
  OAI222_X1 U3734 ( .A1(n3082), .A2(n3163), .B1(n3166), .B2(n1672), .C1(n3098), 
        .C2(n3069), .ZN(N97) );
  OAI222_X1 U3735 ( .A1(n3083), .A2(n3163), .B1(n3166), .B2(n1673), .C1(n3098), 
        .C2(n3070), .ZN(N96) );
  NOR2_X1 U3736 ( .A1(n3167), .A2(n3168), .ZN(N44) );
  INV_X1 U3737 ( .A(n3162), .ZN(n3167) );
  NOR2_X1 U3738 ( .A1(n3162), .A2(n3168), .ZN(N34) );
  NAND3_X1 U3739 ( .A1(n3119), .A2(n3118), .A3(n3120), .ZN(n3168) );
  NAND4_X1 U3740 ( .A1(n3117), .A2(n3116), .A3(n3115), .A4(n3114), .ZN(n3162)
         );
  NOR4_X1 U3741 ( .A1(n3169), .A2(n3068), .A3(n3070), .A4(n3069), .ZN(N296) );
  OR2_X1 U3742 ( .A1(n3066), .A2(n3067), .ZN(n3169) );
  NOR4_X1 U3743 ( .A1(opa_inf), .A2(opa_00), .A3(n3091), .A4(n1570), .ZN(N292)
         );
  NOR3_X1 U3744 ( .A1(n3164), .A2(opa_nan), .A3(n3097), .ZN(N291) );
  NOR3_X1 U3745 ( .A1(prod[11]), .A2(prod[13]), .A3(prod[12]), .ZN(n3170) );
  NOR4_X1 U3746 ( .A1(n3173), .A2(prod[4]), .A3(prod[6]), .A4(prod[5]), .ZN(
        n3172) );
  OR3_X1 U3747 ( .A1(prod[8]), .A2(prod[9]), .A3(prod[7]), .ZN(n3173) );
  NOR3_X1 U3748 ( .A1(prod[21]), .A2(prod[3]), .A3(prod[2]), .ZN(n3171) );
  XNOR2_X1 U3749 ( .A(n3174), .B(n3153), .ZN(N216) );
  INV_X1 U3750 ( .A(n3150), .ZN(n3153) );
  NAND2_X1 U3751 ( .A1(rmode_r2[1]), .A2(rmode_r2[0]), .ZN(n3150) );
  NAND2_X1 U3752 ( .A1(n3175), .A2(n3176), .ZN(N196) );
  NAND2_X1 U3753 ( .A1(n1666), .A2(n3177), .ZN(n3176) );
  NAND2_X1 U3754 ( .A1(n3175), .A2(n3178), .ZN(N195) );
  NAND2_X1 U3755 ( .A1(N151), .A2(n3177), .ZN(n3178) );
  NAND2_X1 U3756 ( .A1(n3175), .A2(n3179), .ZN(N194) );
  NAND2_X1 U3757 ( .A1(N150), .A2(n3177), .ZN(n3179) );
  OAI221_X1 U3758 ( .B1(n3180), .B2(n1578), .C1(n3181), .C2(n1635), .A(n3175), 
        .ZN(N193) );
  OAI221_X1 U3759 ( .B1(n3180), .B2(n1598), .C1(n1636), .C2(n3181), .A(n3175), 
        .ZN(N192) );
  OAI221_X1 U3760 ( .B1(n3180), .B2(n1599), .C1(n1637), .C2(n3181), .A(n3175), 
        .ZN(N191) );
  OAI221_X1 U3761 ( .B1(n3180), .B2(n1577), .C1(n1672), .C2(n3181), .A(n3175), 
        .ZN(N190) );
  OAI221_X1 U3762 ( .B1(n3180), .B2(n1562), .C1(n1673), .C2(n3181), .A(n3175), 
        .ZN(N189) );
  OAI221_X1 U3763 ( .B1(n3180), .B2(n1600), .C1(n3181), .C2(n1624), .A(n3175), 
        .ZN(N188) );
  OAI221_X1 U3764 ( .B1(n3180), .B2(n1601), .C1(n3181), .C2(n1625), .A(n3175), 
        .ZN(N187) );
  OAI221_X1 U3765 ( .B1(n3180), .B2(n1602), .C1(n3181), .C2(n1626), .A(n3175), 
        .ZN(N186) );
  OAI221_X1 U3766 ( .B1(n1558), .B2(n3159), .C1(n3181), .C2(n1627), .A(n3183), 
        .ZN(N185) );
  AOI22_X1 U3767 ( .A1(N141), .A2(n3177), .B1(N116), .B2(n3182), .ZN(n3183) );
  OAI221_X1 U3768 ( .B1(n3159), .B2(n1624), .C1(n3181), .C2(n1678), .A(n3184), 
        .ZN(N184) );
  AOI22_X1 U3769 ( .A1(N140), .A2(n3177), .B1(N115), .B2(n3182), .ZN(n3184) );
  OAI221_X1 U3770 ( .B1(n3159), .B2(n1625), .C1(n3181), .C2(n1679), .A(n3185), 
        .ZN(N183) );
  AOI22_X1 U3771 ( .A1(N139), .A2(n3177), .B1(N114), .B2(n3182), .ZN(n3185) );
  OAI221_X1 U3772 ( .B1(n3159), .B2(n1626), .C1(n1674), .C2(n3181), .A(n3186), 
        .ZN(N182) );
  AOI22_X1 U3773 ( .A1(N138), .A2(n3177), .B1(N113), .B2(n3182), .ZN(n3186) );
  OAI221_X1 U3774 ( .B1(n3159), .B2(n1627), .C1(n1675), .C2(n3181), .A(n3187), 
        .ZN(N181) );
  AOI22_X1 U3775 ( .A1(n3177), .A2(N106), .B1(N112), .B2(n3182), .ZN(n3187) );
  INV_X1 U3776 ( .A(n3180), .ZN(n3177) );
  OAI21_X1 U3777 ( .B1(n1676), .B2(n3181), .A(n3189), .ZN(N180) );
  AOI22_X1 U3778 ( .A1(N111), .A2(n3182), .B1(opa_r1[5]), .B2(n3190), .ZN(
        n3189) );
  OAI21_X1 U3779 ( .B1(n1680), .B2(n3181), .A(n3191), .ZN(N179) );
  AOI22_X1 U3780 ( .A1(N110), .A2(n3182), .B1(opa_r1[4]), .B2(n3190), .ZN(
        n3191) );
  INV_X1 U3781 ( .A(n3159), .ZN(n3190) );
  INV_X1 U3782 ( .A(n3160), .ZN(n3182) );
  NAND2_X1 U3783 ( .A1(n3192), .A2(n3188), .ZN(n3160) );
  INV_X1 U3784 ( .A(n3188), .ZN(n3174) );
  MUX2_X1 U3785 ( .A(sign_fasu), .B(sign_mul), .S(fpu_op_r2[1]), .Z(n3188) );
  NOR2_X1 U3786 ( .A1(opa_r1[11]), .A2(opa_r1[10]), .ZN(n3193) );
  OAI222_X1 U3787 ( .A1(n3079), .A2(n3163), .B1(n3066), .B2(n3164), .C1(n3165), 
        .C2(n1635), .ZN(N100) );
  INV_X1 U3788 ( .A(n3192), .ZN(n3165) );
  NOR2_X1 U3789 ( .A1(fpu_op_r2[1]), .A2(n3166), .ZN(n3192) );
  OR2_X1 U3790 ( .A1(n3097), .A2(n3099), .ZN(n3166) );
  NAND2_X1 U3791 ( .A1(n3099), .A2(fpu_op_r2[1]), .ZN(n3164) );
  NAND2_X1 U3792 ( .A1(n3099), .A2(n3098), .ZN(n3163) );
=======
  fpu_DW01_sub_13 \sub_1_root_u1/sub_133_aco  ( .A({\u1/exp_large[10] , n6263, 
        n6264, \u1/exp_large[7] , \u1/exp_large[6] , \u1/exp_large[5] , 
        \u1/exp_large[4] , \u1/exp_large[3] , \u1/exp_large[2] , 
        \u1/exp_large[1] , \u1/exp_large[0] }), .B({\u1/exp_small [10], n6227, 
        n6228, \u1/exp_small [7:0]}), .CI(\u1/N46 ), .DIFF(\u1/exp_diff2 ) );
  fpu_DW01_sub_14 sub_436_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b1}), .B({opa_r1[57:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .CI(1'b0), .DIFF({N557, 
        N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, 
        N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, 
        N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, 
        N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, 
        N508, N507, N506, N505, N504, N503, N502, N501, 
        SYNOPSYS_UNCONNECTED__109, SYNOPSYS_UNCONNECTED__110, 
        SYNOPSYS_UNCONNECTED__111, SYNOPSYS_UNCONNECTED__112, 
        SYNOPSYS_UNCONNECTED__113, SYNOPSYS_UNCONNECTED__114, 
        SYNOPSYS_UNCONNECTED__115, SYNOPSYS_UNCONNECTED__116, 
        SYNOPSYS_UNCONNECTED__117, SYNOPSYS_UNCONNECTED__118, 
        SYNOPSYS_UNCONNECTED__119, SYNOPSYS_UNCONNECTED__120, 
        SYNOPSYS_UNCONNECTED__121, SYNOPSYS_UNCONNECTED__122, 
        SYNOPSYS_UNCONNECTED__123, SYNOPSYS_UNCONNECTED__124, 
        SYNOPSYS_UNCONNECTED__125, SYNOPSYS_UNCONNECTED__126, 
        SYNOPSYS_UNCONNECTED__127, SYNOPSYS_UNCONNECTED__128, 
        SYNOPSYS_UNCONNECTED__129, SYNOPSYS_UNCONNECTED__130, 
        SYNOPSYS_UNCONNECTED__131, SYNOPSYS_UNCONNECTED__132, 
        SYNOPSYS_UNCONNECTED__133, SYNOPSYS_UNCONNECTED__134, 
        SYNOPSYS_UNCONNECTED__135, SYNOPSYS_UNCONNECTED__136, 
        SYNOPSYS_UNCONNECTED__137, SYNOPSYS_UNCONNECTED__138, 
        SYNOPSYS_UNCONNECTED__139, SYNOPSYS_UNCONNECTED__140, 
        SYNOPSYS_UNCONNECTED__141, SYNOPSYS_UNCONNECTED__142, 
        SYNOPSYS_UNCONNECTED__143, SYNOPSYS_UNCONNECTED__144, 
        SYNOPSYS_UNCONNECTED__145, SYNOPSYS_UNCONNECTED__146, 
        SYNOPSYS_UNCONNECTED__147, SYNOPSYS_UNCONNECTED__148, 
        SYNOPSYS_UNCONNECTED__149, SYNOPSYS_UNCONNECTED__150, 
        SYNOPSYS_UNCONNECTED__151, SYNOPSYS_UNCONNECTED__152, 
        SYNOPSYS_UNCONNECTED__153, SYNOPSYS_UNCONNECTED__154, 
        SYNOPSYS_UNCONNECTED__155, SYNOPSYS_UNCONNECTED__156, 
        SYNOPSYS_UNCONNECTED__157}) );
  fpu_DW01_sub_15 sub_436_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({1'b0, N340, opa_r1[51:0]}), .CI(1'b0), .DIFF({N396, N395, N394, 
        N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, 
        N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, 
        N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, 
        N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, 
        N345, N344, N343}) );
  fpu_DW01_ash_2 sll_386 ( .A({n4602, fracta_mul}), .DATA_TC(1'b0), .SH(
        div_opa_ldz_d), .SH_TC(1'b0), .B({N308, N307, N306, N305, N304, N303, 
        N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, 
        N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, 
        N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, 
        N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256}) );
  fpu_DW01_cmp6_0 r471 ( .A(fracta_mul), .B({\u6/N51 , \u6/N50 , \u6/N49 , 
        \u6/N48 , \u6/N47 , \u6/N46 , \u6/N45 , \u6/N44 , \u6/N43 , \u6/N42 , 
        \u6/N41 , \u6/N40 , \u6/N39 , \u6/N38 , \u6/N37 , \u6/N36 , \u6/N35 , 
        \u6/N34 , \u6/N33 , \u6/N32 , \u6/N31 , \u6/N30 , \u6/N29 , \u6/N28 , 
        \u6/N27 , \u6/N26 , \u6/N25 , \u6/N24 , \u6/N23 , \u6/N22 , \u6/N21 , 
        \u6/N20 , \u6/N19 , \u6/N18 , \u6/N17 , \u6/N16 , \u6/N15 , \u6/N14 , 
        \u6/N13 , \u6/N12 , \u6/N11 , \u6/N10 , \u6/N9 , \u6/N8 , \u6/N7 , 
        \u6/N6 , \u6/N5 , \u6/N4 , \u6/N3 , \u6/N2 , \u6/N1 , \u6/N0 }), .TC(
        1'b0), .LT(\u1/N219 ), .EQ(\u1/N220 ) );
  fpu_DW01_add_9 \add_0_root_sub_0_root_u4/add_497  ( .A({\u4/ldz_dif[10] , 
        \u4/ldz_dif[9] , \u4/ldz_dif[8] , \u4/ldz_dif[7] , \u4/ldz_dif[6] , 
        \u4/ldz_dif[5] , \u4/ldz_dif[4] , \u4/ldz_dif[3] , \u4/ldz_dif[2] , 
        \u4/ldz_dif[1] , \u4/ldz_dif[0] }), .B({1'b0, 1'b0, 1'b0, 
        \u4/fi_ldz_2a[6] , \u4/fi_ldz_2a[6] , \u4/fi_ldz_2a[5] , 
        \u4/fi_ldz_2a[4] , \u4/fi_ldz_2a[3] , \u4/fi_ldz_2a[2] , 
        \u4/fi_ldz_2a[1] , \u4/fi_ldz_2a[0] }), .CI(1'b0), .SUM(\u4/div_exp3 )
         );
  fpu_DW02_mult_0 \u5/mult_82  ( .A({n4602, fracta_mul}), .B({\u6/N52 , 
        \u6/N51 , \u6/N50 , \u6/N49 , \u6/N48 , \u6/N47 , \u6/N46 , \u6/N45 , 
        \u6/N44 , \u6/N43 , \u6/N42 , \u6/N41 , \u6/N40 , \u6/N39 , \u6/N38 , 
        \u6/N37 , \u6/N36 , \u6/N35 , \u6/N34 , \u6/N33 , \u6/N32 , \u6/N31 , 
        \u6/N30 , \u6/N29 , \u6/N28 , \u6/N27 , \u6/N26 , \u6/N25 , \u6/N24 , 
        \u6/N23 , \u6/N22 , \u6/N21 , \u6/N20 , \u6/N19 , \u6/N18 , \u6/N17 , 
        \u6/N16 , \u6/N15 , \u6/N14 , \u6/N13 , \u6/N12 , \u6/N11 , \u6/N10 , 
        \u6/N9 , \u6/N8 , \u6/N7 , \u6/N6 , \u6/N5 , \u6/N4 , \u6/N3 , \u6/N2 , 
        \u6/N1 , \u6/N0 }), .TC(1'b0), .PRODUCT({\u5/N105 , \u5/N104 , 
        \u5/N103 , \u5/N102 , \u5/N101 , \u5/N100 , \u5/N99 , \u5/N98 , 
        \u5/N97 , \u5/N96 , \u5/N95 , \u5/N94 , \u5/N93 , \u5/N92 , \u5/N91 , 
        \u5/N90 , \u5/N89 , \u5/N88 , \u5/N87 , \u5/N86 , \u5/N85 , \u5/N84 , 
        \u5/N83 , \u5/N82 , \u5/N81 , \u5/N80 , \u5/N79 , \u5/N78 , \u5/N77 , 
        \u5/N76 , \u5/N75 , \u5/N74 , \u5/N73 , \u5/N72 , \u5/N71 , \u5/N70 , 
        \u5/N69 , \u5/N68 , \u5/N67 , \u5/N66 , \u5/N65 , \u5/N64 , \u5/N63 , 
        \u5/N62 , \u5/N61 , \u5/N60 , \u5/N59 , \u5/N58 , \u5/N57 , \u5/N56 , 
        \u5/N55 , \u5/N54 , \u5/N53 , \u5/N52 , \u5/N51 , \u5/N50 , \u5/N49 , 
        \u5/N48 , \u5/N47 , \u5/N46 , \u5/N45 , \u5/N44 , \u5/N43 , \u5/N42 , 
        \u5/N41 , \u5/N40 , \u5/N39 , \u5/N38 , \u5/N37 , \u5/N36 , \u5/N35 , 
        \u5/N34 , \u5/N33 , \u5/N32 , \u5/N31 , \u5/N30 , \u5/N29 , \u5/N28 , 
        \u5/N27 , \u5/N26 , \u5/N25 , \u5/N24 , \u5/N23 , \u5/N22 , \u5/N21 , 
        \u5/N20 , \u5/N19 , \u5/N18 , \u5/N17 , \u5/N16 , \u5/N15 , \u5/N14 , 
        \u5/N13 , \u5/N12 , \u5/N11 , \u5/N10 , \u5/N9 , \u5/N8 , \u5/N7 , 
        \u5/N6 , \u5/N5 , \u5/N4 , \u5/N3 , \u5/N2 , \u5/N1 , \u5/N0 }) );
  FA_X1 \u4/sub_412/U2_1  ( .A(div_opa_ldz_r2[1]), .B(n4314), .CI(
        \u4/sub_412/carry [1]), .CO(\u4/sub_412/carry [2]), .S(
        \u4/div_shft4 [1]) );
  FA_X1 \u4/sub_412/U2_2  ( .A(div_opa_ldz_r2[2]), .B(n4438), .CI(
        \u4/sub_412/carry [2]), .CO(\u4/sub_412/carry [3]), .S(
        \u4/div_shft4 [2]) );
  FA_X1 \u4/sub_412/U2_3  ( .A(div_opa_ldz_r2[3]), .B(n4316), .CI(
        \u4/sub_412/carry [3]), .CO(\u4/sub_412/carry [4]), .S(
        \u4/div_shft4 [3]) );
  FA_X1 \u4/sub_412/U2_4  ( .A(div_opa_ldz_r2[4]), .B(n4299), .CI(
        \u4/sub_412/carry [4]), .CO(\u4/sub_412/carry [5]), .S(
        \u4/div_shft4 [4]) );
  FA_X1 \u4/add_411/U1_1  ( .A(div_opa_ldz_r2[1]), .B(exp_r[1]), .CI(
        \u4/add_411/carry [1]), .CO(\u4/add_411/carry [2]), .S(
        \u4/div_shft3[1] ) );
  FA_X1 \u4/add_411/U1_2  ( .A(div_opa_ldz_r2[2]), .B(n4315), .CI(
        \u4/add_411/carry [2]), .CO(\u4/add_411/carry [3]), .S(
        \u4/div_shft3[2] ) );
  FA_X1 \u4/add_411/U1_3  ( .A(div_opa_ldz_r2[3]), .B(n4655), .CI(
        \u4/add_411/carry [3]), .CO(\u4/add_411/carry [4]), .S(
        \u4/div_shft3[3] ) );
  FA_X1 \u4/add_411/U1_4  ( .A(div_opa_ldz_r2[4]), .B(n4282), .CI(
        \u4/add_411/carry [4]), .CO(\u4/add_411/carry [5]), .S(
        \u4/div_shft3[4] ) );
  FA_X1 \u4/sub_409/U2_1  ( .A(exp_r[1]), .B(n4446), .CI(\u4/sub_409/carry [1]), .CO(\u4/sub_409/carry [2]), .S(\u4/div_scht1a [1]) );
  FA_X1 \u4/sub_409/U2_2  ( .A(n4315), .B(n4444), .CI(\u4/sub_409/carry [2]), 
        .CO(\u4/sub_409/carry [3]), .S(\u4/div_scht1a [2]) );
  FA_X1 \u4/sub_409/U2_3  ( .A(n4655), .B(n4443), .CI(\u4/sub_409/carry [3]), 
        .CO(\u4/sub_409/carry [4]), .S(\u4/div_scht1a [3]) );
  FA_X1 \u4/sub_409/U2_4  ( .A(n4282), .B(n4445), .CI(\u4/sub_409/carry [4]), 
        .CO(\u4/sub_409/carry [5]), .S(\u4/div_scht1a [4]) );
  FA_X1 \sub_1_root_sub_0_root_u4/add_497/U2_1  ( .A(exp_r[1]), .B(n4446), 
        .CI(\sub_1_root_sub_0_root_u4/add_497/carry [1]), .CO(
        \sub_1_root_sub_0_root_u4/add_497/carry [2]), .S(\u4/ldz_dif[1] ) );
  FA_X1 \sub_1_root_sub_0_root_u4/add_497/U2_2  ( .A(n4315), .B(n4444), .CI(
        \sub_1_root_sub_0_root_u4/add_497/carry [2]), .CO(
        \sub_1_root_sub_0_root_u4/add_497/carry [3]), .S(\u4/ldz_dif[2] ) );
  FA_X1 \sub_1_root_sub_0_root_u4/add_497/U2_3  ( .A(n4655), .B(n4443), .CI(
        \sub_1_root_sub_0_root_u4/add_497/carry [3]), .CO(
        \sub_1_root_sub_0_root_u4/add_497/carry [4]), .S(\u4/ldz_dif[3] ) );
  FA_X1 \sub_1_root_sub_0_root_u4/add_497/U2_4  ( .A(n4282), .B(n4445), .CI(
        \sub_1_root_sub_0_root_u4/add_497/carry [4]), .CO(
        \sub_1_root_sub_0_root_u4/add_497/carry [5]), .S(\u4/ldz_dif[4] ) );
  NAND2_X2 U3379 ( .A1(quo[2]), .A2(n4563), .ZN(n4027) );
  NAND2_X2 U3380 ( .A1(quo[106]), .A2(n4575), .ZN(n4111) );
  NAND2_X2 U3381 ( .A1(quo[1]), .A2(n4563), .ZN(n3977) );
  NAND2_X2 U3382 ( .A1(quo[105]), .A2(n4574), .ZN(n4113) );
  NOR2_X4 U3383 ( .A1(remainder[56]), .A2(remainder[55]), .ZN(n4152) );
  NOR2_X4 U3384 ( .A1(remainder[51]), .A2(remainder[52]), .ZN(n4151) );
  NOR3_X2 U3385 ( .A1(n3741), .A2(n3849), .A3(n3551), .ZN(n3803) );
  NAND3_X2 U3386 ( .A1(n3851), .A2(n3834), .A3(rmode_r3[1]), .ZN(n3850) );
  NAND3_X2 U3387 ( .A1(n3557), .A2(n2434), .A3(sign), .ZN(n3851) );
  AOI222_X1 U3388 ( .A1(n4600), .A2(n2483), .B1(n4349), .B2(n6342), .C1(
        div_opa_ldz_r2[0]), .C2(n2498), .ZN(n2513) );
  AOI222_X1 U3389 ( .A1(\u4/fi_ldz[1] ), .A2(n2489), .B1(exp_r[1]), .B2(n2483), 
        .C1(\u4/div_scht1a [1]), .C2(n2484), .ZN(n2503) );
  OAI21_X2 U3390 ( .B1(n3767), .B2(n4355), .A(n3768), .ZN(n3477) );
  AOI21_X2 U3391 ( .B1(n6305), .B2(n3773), .A(n3774), .ZN(n3767) );
  NOR3_X2 U3392 ( .A1(n2465), .A2(n2459), .A3(n2462), .ZN(n3856) );
  NAND3_X2 U3393 ( .A1(\u4/exp_out[0] ), .A2(\u4/exp_out[10] ), .A3(
        \u4/exp_out[9] ), .ZN(n3858) );
  NOR3_X2 U3394 ( .A1(fract_denorm[93]), .A2(fract_denorm[94]), .A3(n6357), 
        .ZN(n2707) );
  AOI21_X2 U3395 ( .B1(n2434), .B2(n3557), .A(n3849), .ZN(n3852) );
  NOR3_X2 U3396 ( .A1(n2514), .A2(n2515), .A3(n4355), .ZN(n2498) );
  NAND3_X2 U3397 ( .A1(n2709), .A2(n6413), .A3(n2555), .ZN(n2602) );
  NOR3_X2 U3398 ( .A1(fract_denorm[83]), .A2(fract_denorm[84]), .A3(n6375), 
        .ZN(n2644) );
  AOI21_X2 U3399 ( .B1(n2700), .B2(n6347), .A(n2701), .ZN(n2699) );
  NAND3_X2 U3400 ( .A1(n2660), .A2(n6422), .A3(n2600), .ZN(n2615) );
  NOR3_X2 U3401 ( .A1(fract_denorm[96]), .A2(fract_denorm[97]), .A3(
        fract_denorm[95]), .ZN(n2738) );
  NOR3_X2 U3402 ( .A1(n2635), .A2(n6442), .A3(n6329), .ZN(n2555) );
  AOI21_X2 U3403 ( .B1(n6466), .B2(exp_ovf_r[0]), .A(n5912), .ZN(n3777) );
  AOI21_X2 U3404 ( .B1(\u4/N6251 ), .B2(n3557), .A(n5912), .ZN(n3776) );
  AOI222_X1 U3405 ( .A1(n3829), .A2(\u4/exp_out[10] ), .B1(n3802), .B2(
        \u4/exp_next_mi[10] ), .C1(\u4/exp_out_pl1[10] ), .C2(n3805), .ZN(
        n3842) );
  AOI222_X1 U3406 ( .A1(n3829), .A2(\u4/exp_out[0] ), .B1(n3802), .B2(
        \u4/exp_next_mi[0] ), .C1(\u4/exp_out_pl1[0] ), .C2(n3805), .ZN(n3828)
         );
  AOI211_X2 U3407 ( .C1(n4452), .C2(n3476), .A(n2480), .B(\u4/exp_in_mi1[11] ), 
        .ZN(n2506) );
  NAND3_X2 U3408 ( .A1(n4452), .A2(n3489), .A3(n6447), .ZN(n2518) );
  NOR3_X2 U3409 ( .A1(n6393), .A2(fract_denorm[66]), .A3(n6335), .ZN(n2562) );
  NAND3_X2 U3410 ( .A1(n2609), .A2(n2585), .A3(n2710), .ZN(n2641) );
  NOR3_X2 U3411 ( .A1(n2634), .A2(n6440), .A3(n2632), .ZN(n2639) );
  NOR3_X2 U3412 ( .A1(n2635), .A2(n2636), .A3(n6329), .ZN(n2611) );
  NOR3_X2 U3413 ( .A1(n2648), .A2(n2649), .A3(n2650), .ZN(n2626) );
  NOR3_X2 U3414 ( .A1(fract_denorm[103]), .A2(fract_denorm[104]), .A3(n2662), 
        .ZN(n2761) );
  OAI21_X2 U3415 ( .B1(n4540), .B2(n3787), .A(n3788), .ZN(n3786) );
  OAI21_X2 U3416 ( .B1(n3789), .B2(n3783), .A(n3790), .ZN(n3785) );
  NOR3_X2 U3417 ( .A1(n2515), .A2(n6465), .A3(n4355), .ZN(n2484) );
  AOI211_X2 U3418 ( .C1(n2686), .C2(n4653), .A(n2687), .B(n2688), .ZN(n2673)
         );
  OAI21_X2 U3419 ( .B1(fract_denorm[105]), .B2(n6096), .A(n2514), .ZN(n3963)
         );
  NOR3_X2 U3420 ( .A1(n3608), .A2(n3609), .A3(n3610), .ZN(n3570) );
  NOR2_X2 U3421 ( .A1(n2434), .A2(n3304), .ZN(n3302) );
  NAND3_X2 U3422 ( .A1(n3456), .A2(n3461), .A3(n3342), .ZN(n3463) );
  AOI21_X2 U3423 ( .B1(n6305), .B2(n6459), .A(n3463), .ZN(n3465) );
  OAI21_X2 U3424 ( .B1(n3318), .B2(n3319), .A(n3320), .ZN(n3316) );
  OAI21_X2 U3425 ( .B1(n3551), .B2(n6094), .A(n3552), .ZN(n3550) );
  NOR3_X2 U3426 ( .A1(n3555), .A2(n3556), .A3(n3477), .ZN(n3553) );
  AOI222_X1 U3427 ( .A1(n2679), .A2(fract_denorm[57]), .B1(n2600), .B2(n6424), 
        .C1(n6327), .C2(n6438), .ZN(n2714) );
  NOR3_X2 U3428 ( .A1(n2690), .A2(n2691), .A3(n2664), .ZN(n2712) );
  AOI211_X2 U3429 ( .C1(n2716), .C2(n6362), .A(n4652), .B(n2717), .ZN(n2715)
         );
  NOR2_X2 U3430 ( .A1(n6362), .A2(n2399), .ZN(n2391) );
  NOR2_X2 U3431 ( .A1(n2399), .A2(n6094), .ZN(n2401) );
  INV_X4 U3432 ( .A(n4619), .ZN(n4608) );
  NOR3_X2 U3433 ( .A1(n6440), .A2(n6445), .A3(n6346), .ZN(n3872) );
  AOI21_X2 U3434 ( .B1(n3495), .B2(n4540), .A(n3544), .ZN(n3882) );
  NOR3_X2 U3435 ( .A1(exp_r[1]), .A2(n4655), .A3(n4315), .ZN(n3907) );
  INV_X4 U3436 ( .A(n4616), .ZN(n4613) );
  INV_X4 U3437 ( .A(n4627), .ZN(n4625) );
  INV_X4 U3438 ( .A(n4619), .ZN(n4609) );
  INV_X4 U3439 ( .A(n4627), .ZN(n4624) );
  INV_X4 U3440 ( .A(n4616), .ZN(n4614) );
  NAND2_X2 U3441 ( .A1(n4603), .A2(n6303), .ZN(n3052) );
  NOR2_X2 U3442 ( .A1(n2955), .A2(n6238), .ZN(n2977) );
  NAND3_X2 U3443 ( .A1(n3037), .A2(n3038), .A3(n3039), .ZN(n3036) );
  NAND3_X2 U3444 ( .A1(n3041), .A2(n3042), .A3(n3043), .ZN(n3040) );
  NAND3_X2 U3445 ( .A1(n3045), .A2(n3046), .A3(n3047), .ZN(n3044) );
  NOR2_X2 U3446 ( .A1(\u1/exp_lt_27 ), .A2(\u1/exp_diff[4] ), .ZN(n3012) );
  NOR2_X2 U3447 ( .A1(n2954), .A2(\u1/adj_op[51] ), .ZN(n2976) );
  NOR2_X2 U3448 ( .A1(\u1/exp_lt_27 ), .A2(\u1/exp_diff[3] ), .ZN(n3001) );
  NOR2_X2 U3449 ( .A1(n3004), .A2(n6225), .ZN(n3002) );
  NOR3_X2 U3450 ( .A1(n3004), .A2(n6224), .A3(n3012), .ZN(n3011) );
  NOR3_X2 U3451 ( .A1(fract_denorm[77]), .A2(fract_denorm[78]), .A3(n6385), 
        .ZN(n2728) );
  NAND3_X2 U3452 ( .A1(n6353), .A2(n6354), .A3(n2707), .ZN(n2599) );
  NOR3_X2 U3453 ( .A1(n6409), .A2(n6367), .A3(n6410), .ZN(n2668) );
  NOR3_X2 U3454 ( .A1(n6344), .A2(n6345), .A3(n6441), .ZN(n3878) );
  NOR3_X2 U3455 ( .A1(n3869), .A2(n3870), .A3(n3871), .ZN(n3868) );
  NAND3_X2 U3456 ( .A1(n2683), .A2(n2718), .A3(n2767), .ZN(n3870) );
  NAND3_X2 U3457 ( .A1(n3171), .A2(n2751), .A3(n6400), .ZN(n3871) );
  OAI21_X2 U3458 ( .B1(n3882), .B2(n3883), .A(n3884), .ZN(n3880) );
  NOR3_X2 U3459 ( .A1(n3906), .A2(n3771), .A3(n4540), .ZN(n3883) );
  NAND3_X2 U3460 ( .A1(n3885), .A2(n6337), .A3(exp_ovf_r[1]), .ZN(n3884) );
  NOR3_X2 U3461 ( .A1(n6416), .A2(n6417), .A3(n6418), .ZN(n2670) );
  NOR3_X2 U3462 ( .A1(fract_denorm[53]), .A2(fract_denorm[54]), .A3(n6372), 
        .ZN(n2698) );
  NOR3_X2 U3463 ( .A1(n6380), .A2(n2592), .A3(n6393), .ZN(n4016) );
  NOR3_X2 U3464 ( .A1(fract_denorm[75]), .A2(fract_denorm[76]), .A3(n6382), 
        .ZN(n2560) );
  NOR3_X2 U3465 ( .A1(\u4/N6040 ), .A2(\u4/N6042 ), .A3(\u4/N6041 ), .ZN(n3948) );
  NOR3_X2 U3466 ( .A1(\u4/N6043 ), .A2(\u4/N6045 ), .A3(\u4/N6044 ), .ZN(n3949) );
  NOR3_X2 U3467 ( .A1(\u4/N6046 ), .A2(\u4/N6048 ), .A3(\u4/N6047 ), .ZN(n3950) );
  NOR3_X2 U3468 ( .A1(\u4/N6053 ), .A2(\u4/N6055 ), .A3(\u4/N6054 ), .ZN(n3952) );
  NOR3_X2 U3469 ( .A1(\u4/N6060 ), .A2(\u4/N6062 ), .A3(\u4/N6061 ), .ZN(n3954) );
  NOR3_X2 U3470 ( .A1(\u4/N6027 ), .A2(\u4/N6029 ), .A3(\u4/N6028 ), .ZN(n3944) );
  NOR3_X2 U3471 ( .A1(\u4/N6030 ), .A2(\u4/N6032 ), .A3(\u4/N6031 ), .ZN(n3945) );
  NOR3_X2 U3472 ( .A1(\u4/N6033 ), .A2(\u4/N6035 ), .A3(\u4/N6034 ), .ZN(n3946) );
  NOR3_X2 U3473 ( .A1(\u4/N6014 ), .A2(\u4/N6016 ), .A3(\u4/N6015 ), .ZN(n3940) );
  NOR3_X2 U3474 ( .A1(\u4/N6017 ), .A2(\u4/N6019 ), .A3(\u4/N6018 ), .ZN(n3941) );
  NOR3_X2 U3475 ( .A1(\u4/N6020 ), .A2(\u4/N6022 ), .A3(\u4/N6021 ), .ZN(n3942) );
  NAND3_X2 U3476 ( .A1(n2410), .A2(n2406), .A3(n2413), .ZN(n3505) );
  NOR3_X2 U3477 ( .A1(\u4/fract_out[12] ), .A2(\u4/fract_out[14] ), .A3(
        \u4/fract_out[13] ), .ZN(n3902) );
  NOR3_X2 U3478 ( .A1(\u4/fract_out[36] ), .A2(\u4/fract_out[38] ), .A3(
        \u4/fract_out[37] ), .ZN(n3892) );
  NOR3_X2 U3479 ( .A1(\u4/fract_out[48] ), .A2(\u4/fract_out[4] ), .A3(
        \u4/fract_out[49] ), .ZN(n3896) );
  NOR3_X2 U3480 ( .A1(\u4/fract_out[24] ), .A2(\u4/fract_out[26] ), .A3(
        \u4/fract_out[25] ), .ZN(n3904) );
  OAI21_X2 U3481 ( .B1(\u4/fract_out[0] ), .B2(n3853), .A(n3854), .ZN(n3743)
         );
  AOI21_X2 U3482 ( .B1(sign), .B2(rmode_r3[1]), .A(n6305), .ZN(n3736) );
  NOR3_X2 U3483 ( .A1(n4789), .A2(\u4/fi_ldz_2a[6] ), .A3(\u4/fi_ldz_2a[5] ), 
        .ZN(\u4/N6251 ) );
  NOR2_X2 U3484 ( .A1(n2434), .A2(n6307), .ZN(n3737) );
  NAND3_X2 U3485 ( .A1(n6305), .A2(n4540), .A3(n3849), .ZN(n3855) );
  AOI222_X1 U3486 ( .A1(n4540), .A2(opb_inf), .B1(n3297), .B2(opa_00), .C1(
        n6316), .C2(opb_00), .ZN(n3745) );
  NOR2_X2 U3487 ( .A1(\u1/exp_lt_27 ), .A2(\u1/exp_diff[5] ), .ZN(n3004) );
  INV_X4 U3488 ( .A(n4604), .ZN(n4632) );
  INV_X4 U3489 ( .A(n4605), .ZN(n4604) );
  INV_X4 U3490 ( .A(\u1/expa_lt_expb ), .ZN(n4605) );
  AOI222_X1 U3491 ( .A1(n6213), .A2(n2971), .B1(n6212), .B2(n2972), .C1(n6219), 
        .C2(n2973), .ZN(n2970) );
  NOR2_X2 U3492 ( .A1(n2991), .A2(\u1/adj_op[42] ), .ZN(n2959) );
  NOR2_X2 U3493 ( .A1(n2992), .A2(\u1/adj_op[38] ), .ZN(n2957) );
  NAND3_X2 U3494 ( .A1(n6224), .A2(n3003), .A3(n3002), .ZN(n2958) );
  NOR2_X2 U3495 ( .A1(n2971), .A2(\u1/adj_op[28] ), .ZN(n2996) );
  NAND3_X2 U3496 ( .A1(n6217), .A2(n6224), .A3(n3002), .ZN(n2960) );
  AOI21_X2 U3497 ( .B1(n2976), .B2(n6273), .A(n3001), .ZN(n3008) );
  NOR3_X2 U3498 ( .A1(n3012), .A2(n6217), .A3(n3004), .ZN(n3009) );
  NOR2_X2 U3499 ( .A1(n2978), .A2(\u1/adj_op[44] ), .ZN(n3005) );
  NOR2_X2 U3500 ( .A1(n2979), .A2(n6243), .ZN(n3006) );
  NOR2_X2 U3501 ( .A1(n3010), .A2(n6236), .ZN(n2988) );
  NOR2_X2 U3502 ( .A1(n3000), .A2(n6247), .ZN(n2986) );
  NAND3_X2 U3503 ( .A1(n6217), .A2(n3001), .A3(n3002), .ZN(n2968) );
  NAND3_X2 U3504 ( .A1(n3003), .A2(n3001), .A3(n3002), .ZN(n2966) );
  AOI222_X1 U3505 ( .A1(n4655), .A2(n2483), .B1(\u4/f2i_shft[3] ), .B2(n6342), 
        .C1(div_opa_ldz_r2[3]), .C2(n2498), .ZN(n2500) );
  NOR2_X2 U3506 ( .A1(n6465), .A2(\u4/exp_in_pl1[1] ), .ZN(n2510) );
  AOI222_X1 U3507 ( .A1(n4315), .A2(n2483), .B1(\u4/f2i_shft[2] ), .B2(n6342), 
        .C1(div_opa_ldz_r2[2]), .C2(n2498), .ZN(n2502) );
  AOI222_X1 U3508 ( .A1(n4282), .A2(n2483), .B1(\u4/f2i_shft[4] ), .B2(n6342), 
        .C1(div_opa_ldz_r2[4]), .C2(n2498), .ZN(n2497) );
  AOI222_X1 U3509 ( .A1(\u4/div_scht1a [5]), .A2(n2484), .B1(\u4/f2i_shft[5] ), 
        .B2(n6342), .C1(n4290), .C2(n2483), .ZN(n2494) );
  NAND3_X2 U3510 ( .A1(n3173), .A2(n2729), .A3(n2706), .ZN(n2771) );
  AOI21_X2 U3511 ( .B1(n6371), .B2(n6373), .A(n6326), .ZN(n2591) );
  NOR3_X2 U3512 ( .A1(n6334), .A2(n6401), .A3(n2592), .ZN(n2590) );
  NOR3_X2 U3513 ( .A1(fract_denorm[64]), .A2(fract_denorm[65]), .A3(
        fract_denorm[63]), .ZN(n2735) );
  NOR3_X2 U3514 ( .A1(fract_denorm[61]), .A2(fract_denorm[62]), .A3(n6391), 
        .ZN(n2705) );
  NAND3_X2 U3515 ( .A1(n2560), .A2(fract_denorm[74]), .A3(n6325), .ZN(n2559)
         );
  NOR3_X2 U3516 ( .A1(fract_denorm[80]), .A2(fract_denorm[81]), .A3(
        fract_denorm[79]), .ZN(n2736) );
  OAI21_X2 U3517 ( .B1(n6424), .B2(n6423), .A(n2600), .ZN(n2594) );
  AOI21_X2 U3518 ( .B1(n6336), .B2(n2596), .A(n2597), .ZN(n2595) );
  NAND3_X2 U3519 ( .A1(n6377), .A2(n6379), .A3(n6376), .ZN(n2596) );
  NOR3_X2 U3520 ( .A1(n2598), .A2(n6359), .A3(n2599), .ZN(n2597) );
  AOI211_X2 U3521 ( .C1(fract_denorm[81]), .C2(n6325), .A(n2563), .B(n2573), 
        .ZN(n2572) );
  NAND3_X2 U3522 ( .A1(n6409), .A2(n2711), .A3(n2542), .ZN(n2585) );
  NAND3_X2 U3523 ( .A1(n6416), .A2(n2593), .A3(n2555), .ZN(n2609) );
  NOR3_X2 U3524 ( .A1(fract_denorm[67]), .A2(fract_denorm[68]), .A3(n6396), 
        .ZN(n2646) );
  NOR3_X2 U3525 ( .A1(n2632), .A2(n2696), .A3(n2697), .ZN(n2694) );
  NAND3_X2 U3526 ( .A1(n2707), .A2(fract_denorm[92]), .A3(n6338), .ZN(n2703)
         );
  NOR3_X2 U3527 ( .A1(n2588), .A2(n2625), .A3(n2554), .ZN(n2704) );
  NAND3_X2 U3528 ( .A1(n2708), .A2(n6427), .A3(n2639), .ZN(n2702) );
  NAND3_X2 U3529 ( .A1(n2670), .A2(n6415), .A3(n2555), .ZN(n2607) );
  NOR3_X2 U3530 ( .A1(n6372), .A2(n6370), .A3(n6326), .ZN(n2579) );
  NOR3_X2 U3531 ( .A1(fract_denorm[72]), .A2(fract_denorm[73]), .A3(
        fract_denorm[71]), .ZN(n2661) );
  NOR3_X2 U3532 ( .A1(n6430), .A2(n6431), .A3(n6432), .ZN(n2669) );
  OAI21_X2 U3533 ( .B1(sign), .B2(n3862), .A(n3863), .ZN(n3739) );
  AOI21_X2 U3534 ( .B1(n3880), .B2(n3297), .A(n3881), .ZN(n3862) );
  AOI211_X2 U3535 ( .C1(n3867), .C2(n3868), .A(opas_r2), .B(n4656), .ZN(n3864)
         );
  NAND3_X2 U3536 ( .A1(n3174), .A2(n2752), .A3(n2663), .ZN(n2697) );
  NOR3_X2 U3537 ( .A1(fract_denorm[69]), .A2(fract_denorm[70]), .A3(n6398), 
        .ZN(n2759) );
  NOR3_X2 U3538 ( .A1(fract_denorm[85]), .A2(fract_denorm[86]), .A3(n6378), 
        .ZN(n2760) );
  NOR3_X2 U3539 ( .A1(fract_denorm[56]), .A2(fract_denorm[57]), .A3(
        fract_denorm[55]), .ZN(n2750) );
  NOR3_X2 U3540 ( .A1(fract_denorm[88]), .A2(fract_denorm[89]), .A3(
        fract_denorm[87]), .ZN(n2749) );
  NOR3_X2 U3541 ( .A1(n6423), .A2(n6424), .A3(n6425), .ZN(n2660) );
  NAND3_X2 U3542 ( .A1(n3178), .A2(n2762), .A3(n2695), .ZN(n2635) );
  NOR3_X2 U3543 ( .A1(n2671), .A2(n2771), .A3(n3912), .ZN(n3968) );
  NAND3_X2 U3544 ( .A1(n2644), .A2(n6402), .A3(n6336), .ZN(n2642) );
  NOR3_X2 U3545 ( .A1(n2589), .A2(n6324), .A3(n2557), .ZN(n2727) );
  NAND3_X2 U3546 ( .A1(n6344), .A2(n2724), .A3(n2630), .ZN(n2723) );
  OAI21_X2 U3547 ( .B1(n3865), .B2(n4355), .A(n3866), .ZN(n3853) );
  AOI21_X2 U3548 ( .B1(n3910), .B2(n3911), .A(n3865), .ZN(n3854) );
  NOR3_X2 U3549 ( .A1(remainder[94]), .A2(remainder[96]), .A3(remainder[95]), 
        .ZN(n4165) );
  NOR3_X2 U3550 ( .A1(remainder[88]), .A2(remainder[8]), .A3(remainder[89]), 
        .ZN(n4163) );
  NOR3_X2 U3551 ( .A1(remainder[0]), .A2(remainder[101]), .A3(remainder[100]), 
        .ZN(n4171) );
  NOR3_X2 U3552 ( .A1(remainder[102]), .A2(remainder[104]), .A3(remainder[103]), .ZN(n4172) );
  NOR3_X2 U3553 ( .A1(remainder[105]), .A2(remainder[107]), .A3(remainder[106]), .ZN(n4173) );
  NOR3_X2 U3554 ( .A1(remainder[14]), .A2(remainder[16]), .A3(remainder[15]), 
        .ZN(n4175) );
  NOR3_X2 U3555 ( .A1(remainder[20]), .A2(remainder[22]), .A3(remainder[21]), 
        .ZN(n4177) );
  NOR3_X2 U3556 ( .A1(remainder[27]), .A2(remainder[29]), .A3(remainder[28]), 
        .ZN(n4179) );
  NOR3_X2 U3557 ( .A1(remainder[2]), .A2(remainder[31]), .A3(remainder[30]), 
        .ZN(n4180) );
  NOR3_X2 U3558 ( .A1(remainder[32]), .A2(remainder[34]), .A3(remainder[33]), 
        .ZN(n4181) );
  NOR3_X2 U3559 ( .A1(remainder[39]), .A2(remainder[40]), .A3(remainder[3]), 
        .ZN(n4183) );
  NOR3_X2 U3560 ( .A1(remainder[45]), .A2(remainder[47]), .A3(remainder[46]), 
        .ZN(n4185) );
  NOR3_X2 U3561 ( .A1(remainder[57]), .A2(remainder[59]), .A3(remainder[58]), 
        .ZN(n4153) );
  NOR3_X2 U3562 ( .A1(remainder[63]), .A2(remainder[65]), .A3(remainder[64]), 
        .ZN(n4155) );
  NOR3_X2 U3563 ( .A1(remainder[6]), .A2(remainder[71]), .A3(remainder[70]), 
        .ZN(n4157) );
  NOR3_X2 U3564 ( .A1(remainder[76]), .A2(remainder[78]), .A3(remainder[77]), 
        .ZN(n4159) );
  NOR3_X2 U3565 ( .A1(remainder[79]), .A2(remainder[80]), .A3(remainder[7]), 
        .ZN(n4160) );
  NOR3_X2 U3566 ( .A1(remainder[81]), .A2(remainder[83]), .A3(remainder[82]), 
        .ZN(n4161) );
  NAND3_X2 U3567 ( .A1(n2479), .A2(n4452), .A3(n3487), .ZN(n3486) );
  AOI21_X2 U3568 ( .B1(exp_ovf_r[0]), .B2(n3488), .A(n3489), .ZN(n3487) );
  OAI21_X2 U3569 ( .B1(n2480), .B2(n3494), .A(n3495), .ZN(n3493) );
  NOR3_X2 U3570 ( .A1(n6468), .A2(n4315), .A3(exp_r[1]), .ZN(n3497) );
  OAI21_X2 U3571 ( .B1(n3532), .B2(\u4/N6278 ), .A(n3488), .ZN(n3531) );
  NOR2_X2 U3572 ( .A1(n3488), .A2(n3500), .ZN(n3491) );
  AOI222_X1 U3573 ( .A1(\u4/N6284 ), .A2(\u4/N6283 ), .B1(n3501), .B2(n3502), 
        .C1(n3503), .C2(n3495), .ZN(n3500) );
  NAND3_X2 U3574 ( .A1(opb_dn), .A2(n4271), .A3(\u4/N6194 ), .ZN(n3783) );
  AOI21_X2 U3575 ( .B1(n3771), .B2(n3787), .A(n2480), .ZN(n3789) );
  NAND3_X2 U3576 ( .A1(n4353), .A2(n4656), .A3(n4281), .ZN(n3861) );
  OAI21_X2 U3577 ( .B1(n6465), .B2(n4656), .A(n3556), .ZN(n3788) );
  NAND3_X2 U3578 ( .A1(n4403), .A2(n4338), .A3(n4306), .ZN(n3361) );
  NAND3_X2 U3579 ( .A1(n3734), .A2(n3557), .A3(n3735), .ZN(n3733) );
  OAI21_X2 U3580 ( .B1(n3737), .B2(n3477), .A(n3734), .ZN(n3732) );
  NOR3_X2 U3581 ( .A1(n2439), .A2(n6094), .A3(n3736), .ZN(n3735) );
  NOR2_X2 U3582 ( .A1(exp_ovf_r[0]), .A2(exp_ovf_r[1]), .ZN(n3771) );
  OAI21_X2 U3583 ( .B1(exp_ovf_r[1]), .B2(n3551), .A(n3783), .ZN(n3773) );
  NOR3_X2 U3584 ( .A1(n3618), .A2(n3396), .A3(n3398), .ZN(n3746) );
  NAND3_X2 U3585 ( .A1(n3394), .A2(n3395), .A3(n3393), .ZN(n3748) );
  AOI21_X2 U3586 ( .B1(n3834), .B2(rmode_r3[1]), .A(n3835), .ZN(n3795) );
  OAI22_X2 U3587 ( .A1(\u4/N6410 ), .A2(n3847), .B1(n2441), .B2(n2440), .ZN(
        n3805) );
  NOR2_X2 U3588 ( .A1(n3855), .A2(\u4/N6203 ), .ZN(n3798) );
  NOR2_X2 U3589 ( .A1(n6318), .A2(n3855), .ZN(n3799) );
  NOR2_X2 U3590 ( .A1(n3765), .A2(n3477), .ZN(n3761) );
  NAND3_X2 U3591 ( .A1(exp_ovf_r[1]), .A2(n4356), .A3(n4540), .ZN(n3766) );
  INV_X4 U3592 ( .A(n4631), .ZN(n4616) );
  INV_X4 U3593 ( .A(n4632), .ZN(n4631) );
  INV_X4 U3594 ( .A(n4604), .ZN(n4633) );
  NAND3_X2 U3595 ( .A1(n2969), .A2(n6215), .A3(n2970), .ZN(n2963) );
  OAI21_X2 U3596 ( .B1(n2993), .B2(n2994), .A(n2995), .ZN(n2981) );
  OAI21_X2 U3597 ( .B1(n2983), .B2(n2984), .A(n6222), .ZN(n2982) );
  INV_X4 U3598 ( .A(n4633), .ZN(n4627) );
  NOR3_X2 U3599 ( .A1(\u6/N12 ), .A2(\u6/N14 ), .A3(\u6/N13 ), .ZN(n3104) );
  NOR3_X2 U3600 ( .A1(\u6/N18 ), .A2(\u6/N1 ), .A3(\u6/N19 ), .ZN(n3105) );
  NOR3_X2 U3601 ( .A1(\u6/N23 ), .A2(\u6/N25 ), .A3(\u6/N24 ), .ZN(n3106) );
  NOR2_X2 U3602 ( .A1(fracta_mul[34]), .A2(fracta_mul[35]), .ZN(n3283) );
  NOR3_X2 U3603 ( .A1(n3288), .A2(fracta_mul[7]), .A3(n6302), .ZN(n3267) );
  NOR3_X2 U3604 ( .A1(n6297), .A2(fracta_mul[39]), .A3(n6293), .ZN(n3269) );
  NAND3_X2 U3605 ( .A1(n2434), .A2(n2433), .A3(n6317), .ZN(n2508) );
  AOI222_X1 U3606 ( .A1(\u4/div_scht1a [6]), .A2(n2484), .B1(\u4/f2i_shft[6] ), 
        .B2(n6342), .C1(exp_r[6]), .C2(n2483), .ZN(n2491) );
  AOI21_X2 U3607 ( .B1(n2506), .B2(n6316), .A(n6343), .ZN(n2517) );
  NAND3_X2 U3608 ( .A1(n4540), .A2(n2518), .A3(n2515), .ZN(n2516) );
  INV_X4 U3609 ( .A(n2434), .ZN(n6342) );
  NOR2_X2 U3610 ( .A1(n4289), .A2(n4656), .ZN(n3965) );
  AOI211_X2 U3611 ( .C1(n2542), .C2(n6367), .A(n2590), .B(n2591), .ZN(n2574)
         );
  NOR3_X2 U3612 ( .A1(n6391), .A2(n6389), .A3(n6334), .ZN(n2552) );
  NOR3_X2 U3613 ( .A1(n6396), .A2(n6394), .A3(n6335), .ZN(n2549) );
  AOI211_X2 U3614 ( .C1(n2555), .C2(n6412), .A(n2556), .B(n2557), .ZN(n2544)
         );
  OAI21_X2 U3615 ( .B1(n2558), .B2(n6335), .A(n2559), .ZN(n2556) );
  NOR3_X2 U3616 ( .A1(fract_denorm[70]), .A2(fract_denorm[73]), .A3(
        fract_denorm[72]), .ZN(n2558) );
  NOR3_X2 U3617 ( .A1(n6382), .A2(n6381), .A3(n2642), .ZN(n2625) );
  NOR3_X2 U3618 ( .A1(n6385), .A2(n6383), .A3(n2642), .ZN(n2623) );
  NOR3_X2 U3619 ( .A1(n6375), .A2(n6374), .A3(n2671), .ZN(n2620) );
  NAND3_X2 U3620 ( .A1(n2601), .A2(n2602), .A3(n2603), .ZN(n2570) );
  OAI21_X2 U3621 ( .B1(n6384), .B2(n2642), .A(n2643), .ZN(n2573) );
  NAND3_X2 U3622 ( .A1(n2644), .A2(fract_denorm[82]), .A3(n6336), .ZN(n2643)
         );
  NOR3_X2 U3623 ( .A1(n2632), .A2(n2633), .A3(n2634), .ZN(n2631) );
  AOI21_X2 U3624 ( .B1(n6355), .B2(n6356), .A(n2598), .ZN(n2640) );
  OAI21_X2 U3625 ( .B1(n6390), .B2(n6334), .A(n2645), .ZN(n2564) );
  NAND3_X2 U3626 ( .A1(n2646), .A2(fract_denorm[66]), .A3(n2647), .ZN(n2645)
         );
  NAND3_X2 U3627 ( .A1(n2607), .A2(n2666), .A3(n2667), .ZN(n2649) );
  NOR3_X2 U3628 ( .A1(n2586), .A2(n2623), .A3(n2552), .ZN(n2667) );
  NAND3_X2 U3629 ( .A1(n2669), .A2(n6429), .A3(n2639), .ZN(n2666) );
  AOI211_X2 U3630 ( .C1(n2659), .C2(n6349), .A(n2579), .B(n6331), .ZN(n2658)
         );
  NAND3_X2 U3631 ( .A1(n2663), .A2(n6436), .A3(n6327), .ZN(n2655) );
  NAND3_X2 U3632 ( .A1(n2661), .A2(fract_denorm[70]), .A3(n2647), .ZN(n2657)
         );
  NAND3_X2 U3633 ( .A1(n6352), .A2(n6359), .A3(n6338), .ZN(n2671) );
  NOR3_X2 U3634 ( .A1(n2587), .A2(n2624), .A3(n2553), .ZN(n2734) );
  NOR3_X2 U3635 ( .A1(n2584), .A2(n2622), .A3(n2551), .ZN(n2743) );
  NOR2_X2 U3636 ( .A1(n2641), .A2(n2665), .ZN(n2672) );
  NAND3_X2 U3637 ( .A1(n3180), .A2(n2731), .A3(n2709), .ZN(n2561) );
  NOR3_X2 U3638 ( .A1(n6437), .A2(n6438), .A3(n6439), .ZN(n2663) );
  NOR3_X2 U3639 ( .A1(n6350), .A2(n6351), .A3(n2684), .ZN(n2659) );
  NAND3_X2 U3640 ( .A1(n3176), .A2(n2730), .A3(n2708), .ZN(n2604) );
  NAND3_X2 U3641 ( .A1(n6366), .A2(n2770), .A3(n2542), .ZN(n2632) );
  NOR3_X2 U3642 ( .A1(n6380), .A2(fract_denorm[74]), .A3(n2642), .ZN(n2647) );
  NAND3_X2 U3643 ( .A1(n3879), .A2(n2724), .A3(n2630), .ZN(n2710) );
  NOR2_X2 U3644 ( .A1(n3309), .A2(n4482), .ZN(n3565) );
  NOR2_X2 U3645 ( .A1(n6456), .A2(n3304), .ZN(n3568) );
  NAND3_X2 U3646 ( .A1(n3408), .A2(n3409), .A3(n3407), .ZN(n3589) );
  NAND3_X2 U3647 ( .A1(n3600), .A2(n3422), .A3(n3601), .ZN(n3599) );
  AOI211_X2 U3648 ( .C1(n4656), .C2(opas_r2), .A(n2422), .B(n3548), .ZN(n3547)
         );
  NOR2_X2 U3649 ( .A1(n3539), .A2(n3540), .ZN(n3538) );
  OAI21_X2 U3650 ( .B1(exp_ovf_r[0]), .B2(n3483), .A(n3484), .ZN(n3482) );
  NAND3_X2 U3651 ( .A1(n3485), .A2(n4269), .A3(n3486), .ZN(n3484) );
  NAND3_X2 U3652 ( .A1(n4402), .A2(n4342), .A3(n4311), .ZN(n3375) );
  NAND3_X2 U3653 ( .A1(n4401), .A2(n4341), .A3(n4310), .ZN(n3377) );
  NAND3_X2 U3654 ( .A1(n3338), .A2(n3339), .A3(n3337), .ZN(n3438) );
  NOR3_X2 U3655 ( .A1(n3583), .A2(n3584), .A3(n3585), .ZN(n3397) );
  NAND3_X2 U3656 ( .A1(n3430), .A2(n3431), .A3(n3432), .ZN(n3426) );
  NAND3_X2 U3657 ( .A1(n3415), .A2(n3416), .A3(n3417), .ZN(n3411) );
  NAND3_X2 U3658 ( .A1(n6316), .A2(n3467), .A3(n3468), .ZN(n3320) );
  OAI21_X2 U3659 ( .B1(\u4/N6410 ), .B2(n3454), .A(n6454), .ZN(n3467) );
  NAND3_X2 U3660 ( .A1(n3451), .A2(n3452), .A3(n3453), .ZN(n3447) );
  NOR2_X2 U3661 ( .A1(n4356), .A2(n4452), .ZN(n3556) );
  NAND3_X2 U3662 ( .A1(n2434), .A2(n3741), .A3(n3332), .ZN(n3552) );
  AOI222_X1 U3663 ( .A1(\u4/exp_out[8] ), .A2(n3829), .B1(n3802), .B2(
        \u4/exp_next_mi[8] ), .C1(\u4/exp_out_pl1[8] ), .C2(n3805), .ZN(n3846)
         );
  AOI222_X1 U3664 ( .A1(\u4/exp_out[9] ), .A2(n3829), .B1(n3802), .B2(
        \u4/exp_next_mi[9] ), .C1(\u4/exp_out_pl1[9] ), .C2(n3805), .ZN(n3839)
         );
  OAI21_X2 U3665 ( .B1(n3762), .B2(n3757), .A(n3758), .ZN(n3585) );
  OAI21_X2 U3666 ( .B1(n3756), .B2(n3757), .A(n3758), .ZN(n3534) );
  NOR2_X2 U3667 ( .A1(n3760), .A2(n3761), .ZN(n3750) );
  INV_X4 U3668 ( .A(n3760), .ZN(n6315) );
  NOR2_X2 U3669 ( .A1(n4262), .A2(fpu_op_r2[1]), .ZN(n4194) );
  INV_X4 U3670 ( .A(n4628), .ZN(n4623) );
  INV_X4 U3671 ( .A(n4619), .ZN(n4607) );
  INV_X4 U3672 ( .A(n4617), .ZN(n4612) );
  INV_X4 U3673 ( .A(n4629), .ZN(n4622) );
  INV_X4 U3674 ( .A(n4618), .ZN(n4610) );
  INV_X4 U3675 ( .A(n4617), .ZN(n4611) );
  AOI21_X2 U3676 ( .B1(n2981), .B2(n2982), .A(n6221), .ZN(n2949) );
  AOI21_X2 U3677 ( .B1(n2951), .B2(n2952), .A(n2953), .ZN(n2950) );
  INV_X4 U3678 ( .A(n4627), .ZN(n4626) );
  INV_X4 U3679 ( .A(\u1/fractb_lt_fracta ), .ZN(n4635) );
  NOR3_X2 U3680 ( .A1(fracta_mul[40]), .A2(fracta_mul[41]), .A3(n3243), .ZN(
        n3092) );
  NOR3_X2 U3681 ( .A1(fracta_mul[28]), .A2(fracta_mul[29]), .A3(n3217), .ZN(
        n3091) );
  NOR3_X2 U3682 ( .A1(fracta_mul[46]), .A2(fracta_mul[48]), .A3(fracta_mul[47]), .ZN(n3088) );
  NAND3_X2 U3683 ( .A1(n4272), .A2(n4284), .A3(n4276), .ZN(n3087) );
  NOR3_X2 U3684 ( .A1(n6299), .A2(n6296), .A3(n3090), .ZN(n3083) );
  NOR2_X2 U3685 ( .A1(n3219), .A2(n4367), .ZN(n3256) );
  NOR3_X2 U3686 ( .A1(n6299), .A2(fracta_mul[23]), .A3(n3220), .ZN(n3271) );
  NOR3_X2 U3687 ( .A1(n3204), .A2(n6300), .A3(n4318), .ZN(n3290) );
  NOR3_X2 U3688 ( .A1(n4476), .A2(n3225), .A3(n3204), .ZN(n3258) );
  NOR2_X2 U3689 ( .A1(fracta_mul[10]), .A2(fracta_mul[11]), .ZN(n3245) );
  NAND3_X2 U3690 ( .A1(fracta_mul[9]), .A2(n3245), .A3(n6287), .ZN(n3266) );
  NOR2_X2 U3691 ( .A1(n3206), .A2(n4272), .ZN(n3264) );
  NOR3_X2 U3692 ( .A1(n4371), .A2(n3205), .A3(n3204), .ZN(n3268) );
  NAND3_X2 U3693 ( .A1(fracta_mul[6]), .A2(n3267), .A3(n6288), .ZN(n3236) );
  NAND3_X2 U3694 ( .A1(n4326), .A2(n4368), .A3(n3245), .ZN(n3288) );
  NAND3_X2 U3695 ( .A1(n4372), .A2(n4318), .A3(n3246), .ZN(n3225) );
  NOR3_X2 U3696 ( .A1(fracta_mul[12]), .A2(fracta_mul[13]), .A3(n3225), .ZN(
        n3222) );
  NOR3_X2 U3697 ( .A1(n6302), .A2(fracta_mul[9]), .A3(n4326), .ZN(n3223) );
  NAND3_X2 U3698 ( .A1(n4479), .A2(n4370), .A3(n3261), .ZN(n3217) );
  NAND3_X2 U3699 ( .A1(fracta_mul[40]), .A2(n4472), .A3(n3226), .ZN(n3218) );
  NAND3_X2 U3700 ( .A1(fracta_mul[33]), .A2(n3283), .A3(n3260), .ZN(n3259) );
  NOR3_X2 U3701 ( .A1(fracta_mul[4]), .A2(fracta_mul[5]), .A3(n3205), .ZN(
        n3282) );
  NAND3_X2 U3702 ( .A1(fracta_mul[23]), .A2(n3289), .A3(n6284), .ZN(n3229) );
  AOI211_X2 U3703 ( .C1(fracta_mul[26]), .C2(n6281), .A(n6290), .B(n3270), 
        .ZN(n3230) );
  NAND3_X2 U3704 ( .A1(fracta_mul[24]), .A2(n4473), .A3(n6281), .ZN(n3228) );
  NOR3_X2 U3705 ( .A1(fracta_mul[32]), .A2(fracta_mul[33]), .A3(n6298), .ZN(
        n3261) );
  NOR3_X2 U3706 ( .A1(fracta_mul[36]), .A2(fracta_mul[37]), .A3(n3206), .ZN(
        n3260) );
  NOR3_X2 U3707 ( .A1(n4475), .A2(n3217), .A3(n6279), .ZN(n3257) );
  OAI21_X2 U3708 ( .B1(exp_ovf_r[0]), .B2(n2478), .A(n4452), .ZN(n4141) );
  NOR3_X2 U3709 ( .A1(exp_r[6]), .A2(n4353), .A3(n4281), .ZN(n4142) );
  AOI211_X2 U3710 ( .C1(n2562), .C2(fract_denorm[65]), .A(n2563), .B(n2564), 
        .ZN(n2543) );
  NAND2_X2 U3711 ( .A1(n4269), .A2(n4271), .ZN(n3488) );
  NOR3_X2 U3712 ( .A1(n2641), .A2(n2564), .A3(n2573), .ZN(n2627) );
  NOR2_X2 U3713 ( .A1(n3834), .A2(n4351), .ZN(n3848) );
  OAI21_X2 U3714 ( .B1(opb_dn), .B2(n4398), .A(n3170), .ZN(\fract_div[105] )
         );
  NAND3_X2 U3715 ( .A1(n3488), .A2(n2514), .A3(n4455), .ZN(n2479) );
  OAI21_X2 U3716 ( .B1(n2394), .B2(n3528), .A(n3529), .ZN(n3504) );
  AOI222_X1 U3717 ( .A1(\u4/div_exp1[10] ), .A2(opb_dn), .B1(
        \u4/exp_out1_mi1 [10]), .B2(n2397), .C1(\u4/div_exp2[10] ), .C2(n2398), 
        .ZN(n3528) );
  OAI21_X2 U3718 ( .B1(fract_denorm[102]), .B2(n6363), .A(n6361), .ZN(n2716)
         );
  NAND3_X2 U3719 ( .A1(fract_denorm[99]), .A2(n4653), .A3(n2761), .ZN(n2755)
         );
  NAND3_X2 U3720 ( .A1(n6346), .A2(n2763), .A3(n2700), .ZN(n2754) );
  NAND3_X2 U3721 ( .A1(n6348), .A2(n2751), .A3(n2659), .ZN(n2747) );
  NOR3_X2 U3722 ( .A1(n2580), .A2(n2619), .A3(n2548), .ZN(n2748) );
  NOR3_X2 U3723 ( .A1(n2578), .A2(n2618), .A3(n2547), .ZN(n2766) );
  NOR3_X2 U3724 ( .A1(n2604), .A2(n6441), .A3(n6332), .ZN(n2600) );
  NOR3_X2 U3725 ( .A1(n2592), .A2(fract_denorm[58]), .A3(n6334), .ZN(n2679) );
  NOR2_X2 U3726 ( .A1(n2710), .A2(n6446), .ZN(n2422) );
  NOR2_X2 U3727 ( .A1(n3468), .A2(n4482), .ZN(n3569) );
  NOR2_X2 U3728 ( .A1(qnan_d), .A2(snan_d), .ZN(n3303) );
  NOR3_X2 U3729 ( .A1(n3485), .A2(n3546), .A3(n3547), .ZN(n3542) );
  OAI21_X2 U3730 ( .B1(n3469), .B2(n3470), .A(n3471), .ZN(n3346) );
  NOR2_X2 U3731 ( .A1(n6458), .A2(ind_d), .ZN(n3314) );
  NOR2_X2 U3732 ( .A1(n6458), .A2(inf_d), .ZN(n3457) );
  NOR2_X2 U3733 ( .A1(inf_mul_r), .A2(inf_mul2), .ZN(n3454) );
  NOR2_X2 U3734 ( .A1(n6456), .A2(opb_00), .ZN(n3459) );
  OAI21_X2 U3735 ( .B1(n3764), .B2(n3757), .A(n3758), .ZN(n3584) );
  OAI21_X2 U3736 ( .B1(n3763), .B2(n3757), .A(n3758), .ZN(n3583) );
  AOI21_X2 U3737 ( .B1(n3759), .B2(n6315), .A(n3750), .ZN(n3396) );
  AOI21_X2 U3738 ( .B1(n3755), .B2(n6315), .A(n3750), .ZN(n3540) );
  AOI21_X2 U3739 ( .B1(n3754), .B2(n6315), .A(n3750), .ZN(n3539) );
  AOI21_X2 U3740 ( .B1(n3753), .B2(n6315), .A(n3750), .ZN(n3615) );
  AOI21_X2 U3741 ( .B1(n3752), .B2(n6315), .A(n3750), .ZN(n3389) );
  AOI21_X2 U3742 ( .B1(n3751), .B2(n6315), .A(n3750), .ZN(n3617) );
  AOI21_X2 U3743 ( .B1(n3749), .B2(n6315), .A(n3750), .ZN(n3388) );
  AOI222_X1 U3744 ( .A1(inf_d), .A2(n6339), .B1(opb_00), .B2(n4540), .C1(n4189), .C2(n6316), .ZN(n4188) );
  NOR2_X2 U3745 ( .A1(\u4/N6410 ), .A2(n3454), .ZN(n4189) );
  INV_X4 U3746 ( .A(n4194), .ZN(n6312) );
  NOR2_X2 U3747 ( .A1(fpu_op_r2[1]), .A2(fpu_op_r2[2]), .ZN(n4254) );
  NOR3_X2 U3748 ( .A1(n6275), .A2(n4598), .A3(n6015), .ZN(n2811) );
  NOR3_X2 U3749 ( .A1(n2803), .A2(n6275), .A3(n4597), .ZN(n2810) );
  NOR2_X2 U3750 ( .A1(n6015), .A2(\u1/N46 ), .ZN(n2809) );
  NOR2_X2 U3751 ( .A1(\u2/exp_ovf_d[1] ), .A2(n6275), .ZN(n2808) );
  NAND2_X2 U3752 ( .A1(n6015), .A2(n6275), .ZN(n2805) );
  NAND3_X2 U3753 ( .A1(\u2/N15 ), .A2(\u2/N14 ), .A3(\u2/N6 ), .ZN(n2781) );
  NAND3_X2 U3754 ( .A1(n4597), .A2(n6032), .A3(\u2/N18 ), .ZN(n2777) );
  NAND3_X2 U3755 ( .A1(\u2/N12 ), .A2(\u2/N11 ), .A3(\u2/N13 ), .ZN(n2780) );
  NOR2_X2 U3756 ( .A1(opb_r[62]), .A2(opa_r[62]), .ZN(n2782) );
  OAI22_X2 U3757 ( .A1(n4599), .A2(n6032), .B1(n4597), .B2(n6017), .ZN(
        \u2/exp_tmp4[10] ) );
  NOR3_X2 U3758 ( .A1(opa_r1[54]), .A2(opa_r1[56]), .A3(opa_r1[55]), .ZN(n4250) );
  NAND3_X2 U3759 ( .A1(n4484), .A2(n4381), .A3(n4328), .ZN(n4252) );
  INV_X4 U3760 ( .A(n4648), .ZN(n4647) );
  INV_X4 U3761 ( .A(n4648), .ZN(n4646) );
  NOR2_X2 U3762 ( .A1(\u1/fracta_eq_fractb ), .A2(n3063), .ZN(n3064) );
  AOI211_X2 U3763 ( .C1(n4494), .C2(ind_d), .A(n6458), .B(n3728), .ZN(n3341)
         );
  NOR3_X2 U3764 ( .A1(n4451), .A2(n4456), .A3(n4358), .ZN(n3079) );
  NAND3_X2 U3765 ( .A1(opa_r[61]), .A2(opa_r[62]), .A3(opa_r[60]), .ZN(n3081)
         );
  NOR3_X2 U3766 ( .A1(n4457), .A2(n4359), .A3(n4321), .ZN(n3076) );
  NAND3_X2 U3767 ( .A1(opb_r[61]), .A2(opb_r[62]), .A3(opb_r[60]), .ZN(n3078)
         );
  NOR3_X2 U3768 ( .A1(opa_r[54]), .A2(opa_r[56]), .A3(opa_r[55]), .ZN(n3195)
         );
  NAND3_X2 U3769 ( .A1(n4454), .A2(n4442), .A3(n4453), .ZN(n3197) );
  NOR3_X2 U3770 ( .A1(n3108), .A2(n3109), .A3(n3110), .ZN(n3098) );
  OAI21_X2 U3771 ( .B1(n3279), .B2(n3204), .A(n3266), .ZN(n3278) );
  AOI21_X2 U3772 ( .B1(fracta_mul[17]), .B2(n4369), .A(fracta_mul[19]), .ZN(
        n3279) );
  NOR3_X2 U3773 ( .A1(n4473), .A2(fracta_mul[26]), .A3(n3272), .ZN(n3270) );
  NOR3_X2 U3774 ( .A1(n4472), .A2(n3243), .A3(n6293), .ZN(n3263) );
  NAND3_X2 U3775 ( .A1(fracta_mul[34]), .A2(n4474), .A3(n3260), .ZN(n3254) );
  NAND3_X2 U3776 ( .A1(n4320), .A2(n4283), .A3(n3271), .ZN(n3204) );
  AOI211_X2 U3777 ( .C1(fracta_mul[2]), .C2(n6301), .A(n3274), .B(n3275), .ZN(
        n3273) );
  AOI21_X2 U3778 ( .B1(n4369), .B2(n4319), .A(fracta_mul[19]), .ZN(n3275) );
  NOR2_X2 U3779 ( .A1(fracta_mul[50]), .A2(fracta_mul[49]), .ZN(n3237) );
  AOI21_X2 U3780 ( .B1(n3240), .B2(fracta_mul[47]), .A(n3290), .ZN(n3285) );
  NOR3_X2 U3781 ( .A1(n3287), .A2(n3258), .A3(n3268), .ZN(n3286) );
  NOR3_X2 U3782 ( .A1(fracta_mul[48]), .A2(fracta_mul[51]), .A3(n6296), .ZN(
        n3240) );
  NAND3_X2 U3783 ( .A1(n3207), .A2(n3238), .A3(n3239), .ZN(n3233) );
  NOR3_X2 U3784 ( .A1(fracta_mul[44]), .A2(fracta_mul[45]), .A3(n3219), .ZN(
        n3226) );
  AOI211_X2 U3785 ( .C1(fracta_mul[10]), .C2(n3222), .A(n3223), .B(n3224), 
        .ZN(n3221) );
  NOR3_X2 U3786 ( .A1(n4374), .A2(fracta_mul[13]), .A3(n3225), .ZN(n3224) );
  NAND3_X2 U3787 ( .A1(fracta_mul[3]), .A2(n3282), .A3(n6288), .ZN(n3280) );
  NOR3_X2 U3788 ( .A1(n3204), .A2(fracta_mul[5]), .A3(n3205), .ZN(n3201) );
  NOR2_X2 U3789 ( .A1(n3203), .A2(n6279), .ZN(n3202) );
  NOR3_X2 U3790 ( .A1(fracta_mul[32]), .A2(fracta_mul[34]), .A3(fracta_mul[28]), .ZN(n3203) );
  NOR3_X2 U3791 ( .A1(n3206), .A2(fracta_mul[37]), .A3(n4276), .ZN(n3200) );
  NAND3_X2 U3792 ( .A1(n3228), .A2(n3229), .A3(n3230), .ZN(n3208) );
  NOR3_X2 U3793 ( .A1(n3265), .A2(n3257), .A3(n3291), .ZN(n3198) );
  INV_X4 U3794 ( .A(n3893), .ZN(n4585) );
  NOR2_X2 U3795 ( .A1(\u4/N5904 ), .A2(n3958), .ZN(n3893) );
  NOR3_X2 U3796 ( .A1(n6309), .A2(\u4/f2i_shft[9] ), .A3(\u4/f2i_shft[10] ), 
        .ZN(n3957) );
  AOI222_X1 U3797 ( .A1(n2483), .A2(n6468), .B1(n2484), .B2(n3960), .C1(n3961), 
        .C2(n2485), .ZN(n3959) );
  INV_X4 U3798 ( .A(n4584), .ZN(n4583) );
  INV_X4 U3799 ( .A(n4585), .ZN(n4584) );
  INV_X4 U3800 ( .A(n4349), .ZN(n4600) );
  NOR2_X2 U3801 ( .A1(n2514), .A2(exp_ovf_r[1]), .ZN(n2480) );
  OAI21_X2 U3802 ( .B1(n4542), .B2(n3522), .A(n3523), .ZN(n2427) );
  AOI222_X1 U3803 ( .A1(\u4/div_exp1[8] ), .A2(opb_dn), .B1(
        \u4/exp_out1_mi1 [8]), .B2(n2397), .C1(\u4/div_exp2[8] ), .C2(n2398), 
        .ZN(n3522) );
  OAI21_X2 U3804 ( .B1(n4542), .B2(n3526), .A(n3527), .ZN(n2423) );
  AOI222_X1 U3805 ( .A1(\u4/div_exp1[7] ), .A2(opb_dn), .B1(
        \u4/exp_out1_mi1 [7]), .B2(n2397), .C1(\u4/div_exp2[7] ), .C2(n2398), 
        .ZN(n3526) );
  OAI21_X2 U3806 ( .B1(n2394), .B2(n3515), .A(n3516), .ZN(n2413) );
  AOI222_X1 U3807 ( .A1(\u4/div_exp1[3] ), .A2(opb_dn), .B1(
        \u4/exp_out1_mi1 [3]), .B2(n2397), .C1(\u4/div_exp2[3] ), .C2(n2398), 
        .ZN(n3515) );
  OAI21_X2 U3808 ( .B1(n2394), .B2(n3519), .A(n3520), .ZN(n2410) );
  AOI222_X1 U3809 ( .A1(\u4/div_exp1[2] ), .A2(opb_dn), .B1(
        \u4/exp_out1_mi1 [2]), .B2(n2397), .C1(\u4/div_exp2[2] ), .C2(n2398), 
        .ZN(n3519) );
  NAND3_X2 U3810 ( .A1(fpu_op_r3[0]), .A2(n4400), .A3(n4661), .ZN(n2434) );
  OAI21_X2 U3811 ( .B1(fract_denorm[105]), .B2(n6096), .A(n3964), .ZN(n2438)
         );
  NOR2_X2 U3812 ( .A1(n4452), .A2(n2507), .ZN(n2441) );
  NAND3_X2 U3813 ( .A1(n4274), .A2(n4400), .A3(n4661), .ZN(n2433) );
  INV_X4 U3814 ( .A(n4440), .ZN(n4656) );
  NOR2_X2 U3815 ( .A1(n4355), .A2(n3913), .ZN(n2449) );
  NOR2_X2 U3816 ( .A1(n4540), .A2(n2480), .ZN(n2447) );
  NOR3_X2 U3817 ( .A1(n4355), .A2(n6448), .A3(n2479), .ZN(n2448) );
  OAI21_X2 U3818 ( .B1(n2394), .B2(n3524), .A(n3525), .ZN(n2430) );
  AOI222_X1 U3819 ( .A1(\u4/div_exp1[9] ), .A2(opb_dn), .B1(
        \u4/exp_out1_mi1 [9]), .B2(n2397), .C1(\u4/div_exp2[9] ), .C2(n2398), 
        .ZN(n3524) );
  OAI21_X2 U3820 ( .B1(n4542), .B2(n3517), .A(n3518), .ZN(n2406) );
  AOI222_X1 U3821 ( .A1(\u4/div_exp1[1] ), .A2(opb_dn), .B1(
        \u4/exp_out1_mi1 [1]), .B2(n2397), .C1(\u4/div_exp2[1] ), .C2(n2398), 
        .ZN(n3517) );
  OAI21_X2 U3822 ( .B1(n4542), .B2(n2395), .A(n2396), .ZN(n2393) );
  AOI222_X1 U3823 ( .A1(\u4/div_exp1[0] ), .A2(opb_dn), .B1(
        \u4/exp_out1_mi1 [0]), .B2(n2397), .C1(\u4/div_exp2[0] ), .C2(n2398), 
        .ZN(n2395) );
  NOR2_X2 U3824 ( .A1(n2422), .A2(n2433), .ZN(n2390) );
  OAI21_X2 U3825 ( .B1(n3302), .B2(n3558), .A(n3559), .ZN(N875) );
  OAI21_X2 U3826 ( .B1(n3301), .B2(n3302), .A(n3303), .ZN(n3300) );
  OAI21_X2 U3827 ( .B1(opb_00), .B2(n3304), .A(n4327), .ZN(n3307) );
  NAND3_X2 U3828 ( .A1(n4595), .A2(n3463), .A3(n3457), .ZN(n3462) );
  AOI21_X2 U3829 ( .B1(n3465), .B2(n3466), .A(opa_00), .ZN(n3464) );
  OAI21_X2 U3830 ( .B1(n3386), .B2(n3319), .A(n3387), .ZN(n3345) );
  NAND3_X2 U3831 ( .A1(n3314), .A2(n4595), .A3(inf_d), .ZN(n3313) );
  AOI21_X2 U3832 ( .B1(n3316), .B2(n4291), .A(n3317), .ZN(n3312) );
  NOR2_X2 U3833 ( .A1(n6310), .A2(n3330), .ZN(N794) );
  NOR2_X2 U3834 ( .A1(n6310), .A2(n3329), .ZN(N795) );
  NOR2_X2 U3835 ( .A1(n4545), .A2(n3437), .ZN(N796) );
  NOR2_X2 U3836 ( .A1(n6310), .A2(n3582), .ZN(N797) );
  NOR2_X2 U3837 ( .A1(n4545), .A2(n3581), .ZN(N798) );
  NOR2_X2 U3838 ( .A1(n4545), .A2(n3340), .ZN(N799) );
  NOR2_X2 U3839 ( .A1(n4545), .A2(n3339), .ZN(N800) );
  NOR2_X2 U3840 ( .A1(n4545), .A2(n3338), .ZN(N801) );
  NOR2_X2 U3841 ( .A1(n4545), .A2(n3337), .ZN(N802) );
  NOR2_X2 U3842 ( .A1(n4545), .A2(n3580), .ZN(N803) );
  NOR2_X2 U3843 ( .A1(n4545), .A2(n3579), .ZN(N804) );
  NOR2_X2 U3844 ( .A1(n4545), .A2(n3578), .ZN(N805) );
  NOR2_X2 U3845 ( .A1(n4545), .A2(n3446), .ZN(N806) );
  NOR2_X2 U3846 ( .A1(n4545), .A2(n3445), .ZN(N807) );
  NOR2_X2 U3847 ( .A1(n4545), .A2(n3444), .ZN(N808) );
  NOR2_X2 U3848 ( .A1(n4544), .A2(n3443), .ZN(N809) );
  NOR2_X2 U3849 ( .A1(n4544), .A2(n3595), .ZN(N810) );
  NOR2_X2 U3850 ( .A1(n4544), .A2(n3594), .ZN(N811) );
  NOR2_X2 U3851 ( .A1(n4544), .A2(n3593), .ZN(N812) );
  NOR2_X2 U3852 ( .A1(n4544), .A2(n3452), .ZN(N813) );
  NOR2_X2 U3853 ( .A1(n4544), .A2(n3451), .ZN(N814) );
  NOR2_X2 U3854 ( .A1(n4544), .A2(n3453), .ZN(N815) );
  NOR2_X2 U3855 ( .A1(n4544), .A2(n3592), .ZN(N816) );
  NOR2_X2 U3856 ( .A1(n4544), .A2(n3591), .ZN(N817) );
  NOR2_X2 U3857 ( .A1(n4544), .A2(n3590), .ZN(N818) );
  NOR2_X2 U3858 ( .A1(n4544), .A2(n3410), .ZN(N819) );
  NOR2_X2 U3859 ( .A1(n4544), .A2(n3409), .ZN(N820) );
  NOR2_X2 U3860 ( .A1(n4543), .A2(n3408), .ZN(N821) );
  NOR2_X2 U3861 ( .A1(n4545), .A2(n3407), .ZN(N822) );
  NOR2_X2 U3862 ( .A1(n4545), .A2(n3607), .ZN(N823) );
  NOR2_X2 U3863 ( .A1(n4543), .A2(n3606), .ZN(N824) );
  NOR2_X2 U3864 ( .A1(n4543), .A2(n3605), .ZN(N825) );
  NOR2_X2 U3865 ( .A1(n4545), .A2(n3416), .ZN(N826) );
  NOR2_X2 U3866 ( .A1(n4544), .A2(n3415), .ZN(N827) );
  NOR2_X2 U3867 ( .A1(n4543), .A2(n3417), .ZN(N828) );
  NOR2_X2 U3868 ( .A1(n4544), .A2(n3604), .ZN(N829) );
  NOR2_X2 U3869 ( .A1(n4544), .A2(n3603), .ZN(N830) );
  NOR2_X2 U3870 ( .A1(n4545), .A2(n3602), .ZN(N831) );
  NOR2_X2 U3871 ( .A1(n4543), .A2(n3425), .ZN(N832) );
  NOR2_X2 U3872 ( .A1(n4543), .A2(n3424), .ZN(N833) );
  NOR2_X2 U3873 ( .A1(n4544), .A2(n3423), .ZN(N834) );
  NOR2_X2 U3874 ( .A1(n4543), .A2(n3422), .ZN(N835) );
  NOR2_X2 U3875 ( .A1(n4543), .A2(n3600), .ZN(N836) );
  NOR2_X2 U3876 ( .A1(n4543), .A2(n3601), .ZN(N837) );
  NOR2_X2 U3877 ( .A1(n4543), .A2(n3614), .ZN(N838) );
  NOR2_X2 U3878 ( .A1(n4543), .A2(n3431), .ZN(N839) );
  NOR2_X2 U3879 ( .A1(n4543), .A2(n3430), .ZN(N840) );
  NOR2_X2 U3880 ( .A1(n4543), .A2(n3432), .ZN(N841) );
  NOR2_X2 U3881 ( .A1(n4543), .A2(n3613), .ZN(N842) );
  NOR2_X2 U3882 ( .A1(n4543), .A2(n3612), .ZN(N843) );
  NOR2_X2 U3883 ( .A1(n4543), .A2(n3611), .ZN(N844) );
  AOI21_X2 U3884 ( .B1(n3457), .B2(n3458), .A(n3459), .ZN(n3455) );
  NOR3_X2 U3885 ( .A1(opb_r[54]), .A2(opb_r[56]), .A3(opb_r[55]), .ZN(n3093)
         );
  NAND3_X2 U3886 ( .A1(n4399), .A2(n4340), .A3(n4296), .ZN(n3095) );
  NAND3_X2 U3887 ( .A1(exp_mul[6]), .A2(exp_mul[5]), .A3(exp_mul[7]), .ZN(
        n3294) );
  NOR3_X2 U3888 ( .A1(n4487), .A2(n4383), .A3(n4330), .ZN(n3295) );
  NAND3_X2 U3889 ( .A1(n6016), .A2(n4597), .A3(n2782), .ZN(n2832) );
  AOI21_X2 U3890 ( .B1(n2801), .B2(n2802), .A(n4458), .ZN(\u2/exp_ovf_d[0] )
         );
  NOR2_X2 U3891 ( .A1(n2772), .A2(n6274), .ZN(\u2/underflow_d [2]) );
  OAI21_X2 U3892 ( .B1(n4597), .B2(n2833), .A(n2834), .ZN(\u2/N114 ) );
  OAI21_X2 U3893 ( .B1(n4191), .B2(n4380), .A(n4203), .ZN(N710) );
  OAI21_X2 U3894 ( .B1(n4191), .B2(n4488), .A(n4202), .ZN(N711) );
  NOR2_X2 U3895 ( .A1(n3059), .A2(n6262), .ZN(\u1/N62 ) );
  NOR2_X2 U3896 ( .A1(n3059), .A2(n3050), .ZN(\u1/N61 ) );
  NOR2_X2 U3897 ( .A1(n3059), .A2(n3051), .ZN(\u1/N60 ) );
  NOR2_X2 U3898 ( .A1(n3059), .A2(n6265), .ZN(\u1/N59 ) );
  NOR2_X2 U3899 ( .A1(n3059), .A2(n6266), .ZN(\u1/N58 ) );
  NOR2_X2 U3900 ( .A1(n3059), .A2(n6267), .ZN(\u1/N57 ) );
  NOR2_X2 U3901 ( .A1(n3059), .A2(n6268), .ZN(\u1/N56 ) );
  NOR2_X2 U3902 ( .A1(n3059), .A2(n6269), .ZN(\u1/N55 ) );
  NOR2_X2 U3903 ( .A1(n3059), .A2(n6270), .ZN(\u1/N54 ) );
  NOR2_X2 U3904 ( .A1(n3059), .A2(n6271), .ZN(\u1/N53 ) );
  NOR2_X2 U3905 ( .A1(n3059), .A2(n6272), .ZN(\u1/N52 ) );
  OAI21_X2 U3906 ( .B1(n3060), .B2(n4495), .A(n3061), .ZN(\u1/N229 ) );
  OAI21_X2 U3907 ( .B1(n3062), .B2(n4492), .A(\u1/signa_r ), .ZN(n3061) );
  NOR3_X2 U3908 ( .A1(n3063), .A2(\u1/fracta_lt_fractb ), .A3(
        \u1/fracta_eq_fractb ), .ZN(n3062) );
  NOR2_X2 U3909 ( .A1(n4661), .A2(n3341), .ZN(N904) );
  NOR2_X2 U3910 ( .A1(n3071), .A2(n3070), .ZN(\u0/N6 ) );
  NOR2_X2 U3911 ( .A1(fracta_mul[51]), .A2(n3073), .ZN(\u0/N4 ) );
  NOR3_X2 U3912 ( .A1(n4493), .A2(opa_nan), .A3(n3296), .ZN(N912) );
  NOR2_X2 U3913 ( .A1(n4267), .A2(n3075), .ZN(\u0/N10 ) );
  NOR2_X2 U3914 ( .A1(n4268), .A2(n3074), .ZN(\u0/N11 ) );
  NOR2_X2 U3915 ( .A1(n3072), .A2(\u6/N51 ), .ZN(n4268) );
  AOI21_X2 U3916 ( .B1(fracta_mul[49]), .B2(n4480), .A(n3209), .ZN(n3276) );
  NOR2_X2 U3917 ( .A1(n3273), .A2(n3204), .ZN(n3249) );
  AOI211_X2 U3918 ( .C1(n3240), .C2(fracta_mul[46]), .A(n3241), .B(n3242), 
        .ZN(n3231) );
  AOI211_X2 U3919 ( .C1(n3226), .C2(fracta_mul[42]), .A(n3227), .B(n3208), 
        .ZN(n3212) );
  NOR3_X2 U3920 ( .A1(n3219), .A2(fracta_mul[45]), .A3(n4277), .ZN(n3215) );
  INV_X4 U3921 ( .A(n4583), .ZN(n4579) );
  INV_X4 U3922 ( .A(n4585), .ZN(n4580) );
  INV_X4 U3923 ( .A(n4583), .ZN(n4581) );
  INV_X4 U3924 ( .A(n4585), .ZN(n4582) );
  INV_X4 U3925 ( .A(n4583), .ZN(n4578) );
  NAND2_X2 U3926 ( .A1(n2480), .A2(n4355), .ZN(n2442) );
  OAI21_X2 U3927 ( .B1(n4542), .B2(n3513), .A(n3514), .ZN(n3512) );
  AOI222_X1 U3928 ( .A1(\u4/div_exp1[6] ), .A2(opb_dn), .B1(
        \u4/exp_out1_mi1 [6]), .B2(n2397), .C1(\u4/div_exp2[6] ), .C2(n2398), 
        .ZN(n3513) );
  OAI21_X2 U3929 ( .B1(n2394), .B2(n3507), .A(n3508), .ZN(n3506) );
  AOI222_X1 U3930 ( .A1(\u4/div_exp1[5] ), .A2(opb_dn), .B1(
        \u4/exp_out1_mi1 [5]), .B2(n2397), .C1(\u4/div_exp2[5] ), .C2(n2398), 
        .ZN(n3507) );
  OAI21_X2 U3931 ( .B1(n2394), .B2(n3510), .A(n3511), .ZN(n3509) );
  AOI222_X1 U3932 ( .A1(\u4/div_exp1[4] ), .A2(opb_dn), .B1(
        \u4/exp_out1_mi1 [4]), .B2(n2397), .C1(\u4/div_exp2[4] ), .C2(n2398), 
        .ZN(n3510) );
  INV_X4 U3933 ( .A(n2401), .ZN(n2408) );
  NOR3_X2 U3934 ( .A1(n2434), .A2(n6309), .A3(n2435), .ZN(n2400) );
  NAND3_X2 U3935 ( .A1(n2436), .A2(n2433), .A3(n2437), .ZN(n2399) );
  AOI21_X2 U3936 ( .B1(n6316), .B2(n2438), .A(n2439), .ZN(n2437) );
  NAND3_X2 U3937 ( .A1(n2440), .A2(n4356), .A3(n2441), .ZN(n2436) );
  AOI222_X1 U3938 ( .A1(\u4/fi_ldz_2a[0] ), .A2(n2390), .B1(n2391), .B2(n6094), 
        .C1(n4540), .C2(n2393), .ZN(n2389) );
  NOR3_X2 U3939 ( .A1(\u4/N5945 ), .A2(\u4/N5947 ), .A3(\u4/N5946 ), .ZN(n3932) );
  NOR3_X2 U3940 ( .A1(\u4/N5952 ), .A2(\u4/N5954 ), .A3(\u4/N5953 ), .ZN(n3934) );
  NOR3_X2 U3941 ( .A1(\u4/N5932 ), .A2(\u4/N5934 ), .A3(\u4/N5933 ), .ZN(n3928) );
  NOR3_X2 U3942 ( .A1(\u4/N5935 ), .A2(\u4/N5937 ), .A3(\u4/N5936 ), .ZN(n3929) );
  NOR3_X2 U3943 ( .A1(\u4/N5938 ), .A2(\u4/N5940 ), .A3(\u4/N5939 ), .ZN(n3930) );
  NOR3_X2 U3944 ( .A1(\u4/N5919 ), .A2(\u4/N5921 ), .A3(\u4/N5920 ), .ZN(n3924) );
  NOR3_X2 U3945 ( .A1(\u4/N5922 ), .A2(\u4/N5924 ), .A3(\u4/N5923 ), .ZN(n3925) );
  NOR3_X2 U3946 ( .A1(\u4/N5925 ), .A2(\u4/N5927 ), .A3(\u4/N5926 ), .ZN(n3926) );
  NOR3_X2 U3947 ( .A1(\u4/N5906 ), .A2(\u4/N5908 ), .A3(\u4/N5907 ), .ZN(n3920) );
  NOR3_X2 U3948 ( .A1(\u4/N5909 ), .A2(\u4/N5911 ), .A3(\u4/N5910 ), .ZN(n3921) );
  NOR3_X2 U3949 ( .A1(\u4/N5912 ), .A2(\u4/N5914 ), .A3(\u4/N5913 ), .ZN(n3922) );
  INV_X4 U3950 ( .A(n4620), .ZN(n4606) );
  INV_X4 U3951 ( .A(n4650), .ZN(n4642) );
  INV_X4 U3952 ( .A(n4630), .ZN(n4619) );
  INV_X4 U3953 ( .A(n4616), .ZN(n4615) );
  INV_X4 U3954 ( .A(n4569), .ZN(n4566) );
  INV_X4 U3955 ( .A(n4568), .ZN(n4567) );
  INV_X4 U3956 ( .A(n4632), .ZN(n4630) );
  INV_X4 U3957 ( .A(n4660), .ZN(n4659) );
  INV_X4 U3958 ( .A(n4632), .ZN(n4629) );
  AND2_X4 U3959 ( .A1(n3734), .A2(n3742), .ZN(n4278) );
  AND2_X4 U3960 ( .A1(n3734), .A2(n3738), .ZN(n4279) );
  OR2_X4 U3961 ( .A1(n4269), .A2(n3458), .ZN(n4280) );
  INV_X4 U3962 ( .A(n4634), .ZN(n4650) );
  INV_X4 U3963 ( .A(n4635), .ZN(n4634) );
  INV_X4 U3964 ( .A(n4633), .ZN(n4628) );
  INV_X4 U3965 ( .A(n4629), .ZN(n4621) );
  NAND2_X2 U3966 ( .A1(n3732), .A2(n3733), .ZN(n4288) );
  INV_X4 U3967 ( .A(n4565), .ZN(n4564) );
  INV_X4 U3968 ( .A(n4634), .ZN(n4645) );
  INV_X4 U3969 ( .A(n4634), .ZN(n4644) );
  INV_X4 U3970 ( .A(n4634), .ZN(n4643) );
  NOR2_X2 U3971 ( .A1(n4271), .A2(n4269), .ZN(n2394) );
  INV_X4 U3972 ( .A(n4541), .ZN(n4542) );
  INV_X4 U3973 ( .A(n4631), .ZN(n4618) );
  NAND2_X2 U3974 ( .A1(n4187), .A2(n2433), .ZN(n3619) );
  AND2_X4 U3975 ( .A1(n6312), .A2(n6313), .ZN(n4293) );
  INV_X4 U3976 ( .A(n4291), .ZN(n4661) );
  NOR3_X2 U3977 ( .A1(\u4/N6172 ), .A2(\u4/N6171 ), .A3(n4271), .ZN(n2398) );
  INV_X4 U3978 ( .A(n4280), .ZN(n4572) );
  INV_X4 U3979 ( .A(n3973), .ZN(n4569) );
  INV_X4 U3980 ( .A(n4650), .ZN(n4639) );
  INV_X4 U3981 ( .A(n4644), .ZN(n4637) );
  INV_X4 U3982 ( .A(n4645), .ZN(n4636) );
  AND3_X4 U3983 ( .A1(n4194), .A2(n6313), .A3(N396), .ZN(n4302) );
  OR2_X4 U3984 ( .A1(n6312), .A2(n6313), .ZN(n4304) );
  NOR2_X2 U3985 ( .A1(n3458), .A2(opb_dn), .ZN(n4309) );
  INV_X4 U3986 ( .A(n4280), .ZN(n4570) );
  INV_X4 U3987 ( .A(n3956), .ZN(n4576) );
  NOR2_X2 U3988 ( .A1(n3488), .A2(n2480), .ZN(n2397) );
  INV_X4 U3989 ( .A(n4650), .ZN(n4641) );
  INV_X4 U3990 ( .A(n4650), .ZN(n4640) );
  INV_X4 U3991 ( .A(n4650), .ZN(n4638) );
  INV_X4 U3992 ( .A(\u2/N157 ), .ZN(n4601) );
  INV_X8 U3993 ( .A(n4603), .ZN(n4602) );
  INV_X4 U3994 ( .A(\u2/N157 ), .ZN(n4603) );
  INV_X4 U3995 ( .A(n4631), .ZN(n4617) );
  INV_X4 U3996 ( .A(n4302), .ZN(n4556) );
  INV_X4 U3997 ( .A(n4302), .ZN(n4554) );
  INV_X4 U3998 ( .A(n4302), .ZN(n4555) );
  INV_X4 U3999 ( .A(n3619), .ZN(n4545) );
  INV_X4 U4000 ( .A(n3619), .ZN(n4543) );
  INV_X4 U4001 ( .A(n3619), .ZN(n4544) );
  INV_X4 U4002 ( .A(n4379), .ZN(n4598) );
  INV_X4 U4003 ( .A(n4598), .ZN(n4597) );
  INV_X4 U4004 ( .A(n4562), .ZN(n4561) );
  NOR2_X2 U4005 ( .A1(n6312), .A2(n4190), .ZN(n4197) );
  OR2_X4 U4006 ( .A1(n4720), .A2(\u4/exp_out[4] ), .ZN(n4337) );
  OR2_X4 U4007 ( .A1(n4713), .A2(\u4/sub_468/A[4] ), .ZN(n4339) );
  NOR2_X2 U4008 ( .A1(fpu_op_r3[1]), .A2(n4661), .ZN(n3315) );
  INV_X4 U4009 ( .A(n4278), .ZN(n4593) );
  INV_X4 U4010 ( .A(n4288), .ZN(n4586) );
  INV_X4 U4011 ( .A(n4280), .ZN(n4574) );
  INV_X4 U4012 ( .A(n4280), .ZN(n4573) );
  INV_X4 U4013 ( .A(n4309), .ZN(n4565) );
  INV_X4 U4014 ( .A(n4291), .ZN(n4662) );
  INV_X4 U4015 ( .A(n4653), .ZN(n4652) );
  INV_X4 U4016 ( .A(n4652), .ZN(n4654) );
  INV_X4 U4017 ( .A(fract_denorm[105]), .ZN(n4653) );
  INV_X4 U4018 ( .A(n3973), .ZN(n4568) );
  OR2_X4 U4019 ( .A1(n4692), .A2(exp_r[6]), .ZN(n4354) );
  INV_X4 U4020 ( .A(n4316), .ZN(n4655) );
  OR2_X4 U4021 ( .A1(n3458), .A2(n4661), .ZN(n4355) );
  INV_X4 U4022 ( .A(n4651), .ZN(n4648) );
  INV_X4 U4023 ( .A(n4634), .ZN(n4651) );
  NAND4_X2 U4024 ( .A1(n2712), .A2(n2713), .A3(n2714), .A4(n2715), .ZN(
        \u4/fi_ldz_2a[0] ) );
  OR2_X4 U4025 ( .A1(n4679), .A2(\u2/exp_tmp4[4] ), .ZN(n4378) );
  NAND3_X2 U4026 ( .A1(fpu_op_r1[0]), .A2(n4377), .A3(fpu_op_r1[1]), .ZN(n4379) );
  INV_X4 U4027 ( .A(n4191), .ZN(n4562) );
  INV_X4 U4028 ( .A(n4304), .ZN(n4552) );
  INV_X4 U4029 ( .A(n4293), .ZN(n4558) );
  INV_X4 U4030 ( .A(n4293), .ZN(n4557) );
  INV_X4 U4031 ( .A(n4305), .ZN(n4657) );
  INV_X4 U4032 ( .A(n4305), .ZN(n4658) );
  NOR2_X2 U4033 ( .A1(n2518), .A2(n4355), .ZN(n2483) );
  INV_X4 U4034 ( .A(n4279), .ZN(n4590) );
  INV_X4 U4035 ( .A(n4279), .ZN(n4591) );
  INV_X4 U4036 ( .A(n4279), .ZN(n4589) );
  INV_X4 U4037 ( .A(n4278), .ZN(n4592) );
  INV_X4 U4038 ( .A(n4278), .ZN(n4594) );
  INV_X4 U4039 ( .A(n4288), .ZN(n4587) );
  INV_X4 U4040 ( .A(n4288), .ZN(n4588) );
  INV_X4 U4041 ( .A(n3315), .ZN(n4596) );
  INV_X4 U4042 ( .A(n4596), .ZN(n4595) );
  NAND4_X2 U4043 ( .A1(n2626), .A2(n2627), .A3(n2628), .A4(n2629), .ZN(
        \u4/fi_ldz[3] ) );
  INV_X4 U4044 ( .A(n4280), .ZN(n4571) );
  INV_X4 U4045 ( .A(n4280), .ZN(n4575) );
  INV_X4 U4046 ( .A(n4565), .ZN(n4563) );
  NAND4_X2 U4047 ( .A1(n2565), .A2(n2566), .A3(n2567), .A4(n2568), .ZN(
        \u4/fi_ldz[4] ) );
  NAND4_X2 U4048 ( .A1(n2543), .A2(n2544), .A3(n2545), .A4(n2546), .ZN(
        \u4/fi_ldz[5] ) );
  INV_X4 U4049 ( .A(n3956), .ZN(n4577) );
  NOR2_X2 U4050 ( .A1(n4352), .A2(\u4/sub_409/carry [10]), .ZN(n4455) );
  INV_X4 U4051 ( .A(n2394), .ZN(n4541) );
  INV_X4 U4052 ( .A(n4650), .ZN(n4649) );
  INV_X4 U4053 ( .A(n4355), .ZN(n4540) );
  INV_X4 U4054 ( .A(n4630), .ZN(n4620) );
  NAND2_X2 U4055 ( .A1(n4351), .A2(n4441), .ZN(\u4/N6410 ) );
  INV_X4 U4056 ( .A(n2800), .ZN(\u2/lt_135/A[0] ) );
  INV_X4 U4057 ( .A(n4304), .ZN(n4553) );
  INV_X4 U4058 ( .A(n4304), .ZN(n4550) );
  INV_X4 U4059 ( .A(n4304), .ZN(n4551) );
  INV_X4 U4060 ( .A(n4197), .ZN(n4549) );
  INV_X4 U4061 ( .A(n4549), .ZN(n4546) );
  INV_X4 U4062 ( .A(n4549), .ZN(n4547) );
  INV_X4 U4063 ( .A(n4549), .ZN(n4548) );
  INV_X4 U4064 ( .A(n4293), .ZN(n4559) );
  INV_X4 U4065 ( .A(n4293), .ZN(n4560) );
  INV_X4 U4066 ( .A(n4305), .ZN(n4660) );
  INV_X4 U4067 ( .A(n4379), .ZN(n4599) );
  OAI22_X2 U4068 ( .A1(\u4/fi_ldz_2a[6] ), .A2(n4812), .B1(\u4/fi_ldz_2a[6] ), 
        .B2(\u4/fi_ldz_2a[5] ), .ZN(\u4/N6249 ) );
  OR2_X4 U4069 ( .A1(n4303), .A2(fpu_op_r2[2]), .ZN(n3296) );
  AND2_X4 U4070 ( .A1(n3848), .A2(n2441), .ZN(n3804) );
  AND3_X4 U4071 ( .A1(n6305), .A2(n4355), .A3(n3849), .ZN(n3802) );
  AND3_X4 U4072 ( .A1(\u1/N220 ), .A2(n6099), .A3(\u1/N49 ), .ZN(n3059) );
  AND3_X4 U4073 ( .A1(n6404), .A2(n6403), .A3(n2637), .ZN(n2542) );
  OR4_X4 U4074 ( .A1(n2651), .A2(n2652), .A3(n2653), .A4(n2654), .ZN(
        \u4/fi_ldz[2] ) );
  AND2_X4 U4075 ( .A1(n2478), .A2(n4540), .ZN(n2446) );
  XNOR2_X1 U4076 ( .A(\u4/fi_ldz[6] ), .B(\u4/sub_463/carry[6] ), .ZN(
        \u4/fi_ldz_mi22 [6]) );
  AND2_X1 U4077 ( .A1(\u4/sub_463/carry[5] ), .A2(\u4/fi_ldz[5] ), .ZN(
        \u4/sub_463/carry[6] ) );
  XOR2_X1 U4078 ( .A(\u4/fi_ldz[5] ), .B(\u4/sub_463/carry[5] ), .Z(
        \u4/fi_ldz_mi22 [5]) );
  AND2_X1 U4079 ( .A1(\u4/sub_463/carry[4] ), .A2(\u4/fi_ldz[4] ), .ZN(
        \u4/sub_463/carry[5] ) );
  XOR2_X1 U4080 ( .A(\u4/fi_ldz[4] ), .B(\u4/sub_463/carry[4] ), .Z(
        \u4/fi_ldz_mi22 [4]) );
  OR2_X1 U4081 ( .A1(\u4/fi_ldz[3] ), .A2(\u4/sub_463/carry[3] ), .ZN(
        \u4/sub_463/carry[4] ) );
  XNOR2_X1 U4082 ( .A(\u4/sub_463/carry[3] ), .B(\u4/fi_ldz[3] ), .ZN(
        \u4/fi_ldz_mi22 [3]) );
  OR2_X1 U4083 ( .A1(\u4/fi_ldz[2] ), .A2(\u4/sub_463/carry[2] ), .ZN(
        \u4/sub_463/carry[3] ) );
  XNOR2_X1 U4084 ( .A(\u4/sub_463/carry[2] ), .B(\u4/fi_ldz[2] ), .ZN(
        \u4/fi_ldz_mi22 [2]) );
  AND2_X1 U4085 ( .A1(\u4/fi_ldz_2a[0] ), .A2(\u4/fi_ldz[1] ), .ZN(
        \u4/sub_463/carry[2] ) );
  XOR2_X1 U4086 ( .A(\u4/fi_ldz[1] ), .B(\u4/fi_ldz_2a[0] ), .Z(
        \u4/fi_ldz_mi22 [1]) );
  XOR2_X1 U4087 ( .A(n4656), .B(\u4/add_410/carry [10]), .Z(\u4/div_shft2 [10]) );
  AND2_X1 U4088 ( .A1(n4289), .A2(\u4/add_410/carry [9]), .ZN(
        \u4/add_410/carry [10]) );
  XOR2_X1 U4089 ( .A(n4289), .B(\u4/add_410/carry [9]), .Z(\u4/div_shft2 [9])
         );
  XOR2_X1 U4090 ( .A(n4656), .B(\u4/add_411/carry [10]), .Z(\u4/div_shft3[10] ) );
  AND2_X1 U4091 ( .A1(n4289), .A2(\u4/add_411/carry [9]), .ZN(
        \u4/add_411/carry [10]) );
  XOR2_X1 U4092 ( .A(n4289), .B(\u4/add_411/carry [9]), .Z(\u4/div_shft3[9] )
         );
  XOR2_X1 U4093 ( .A(n4440), .B(\u4/sub_412/carry [10]), .Z(\u4/div_shft4 [10]) );
  AND2_X1 U4094 ( .A1(\u4/sub_412/carry [9]), .A2(n4350), .ZN(
        \u4/sub_412/carry [10]) );
  XOR2_X1 U4095 ( .A(n4350), .B(\u4/sub_412/carry [9]), .Z(\u4/div_shft4 [9])
         );
  XNOR2_X1 U4096 ( .A(n4656), .B(\sub_1_root_sub_0_root_u4/add_497/carry [10]), 
        .ZN(\u4/ldz_dif[10] ) );
  OR2_X1 U4097 ( .A1(n4289), .A2(\sub_1_root_sub_0_root_u4/add_497/carry [9]), 
        .ZN(\sub_1_root_sub_0_root_u4/add_497/carry [10]) );
  XNOR2_X1 U4098 ( .A(\sub_1_root_sub_0_root_u4/add_497/carry [9]), .B(n4289), 
        .ZN(\u4/ldz_dif[9] ) );
  AND2_X1 U4099 ( .A1(n4353), .A2(\u4/add_410/carry [8]), .ZN(
        \u4/add_410/carry [9]) );
  XOR2_X1 U4100 ( .A(n4353), .B(\u4/add_410/carry [8]), .Z(\u4/div_shft2 [8])
         );
  AND2_X1 U4101 ( .A1(n4353), .A2(\u4/add_411/carry [8]), .ZN(
        \u4/add_411/carry [9]) );
  XOR2_X1 U4102 ( .A(n4353), .B(\u4/add_411/carry [8]), .Z(\u4/div_shft3[8] )
         );
  AND2_X1 U4103 ( .A1(\u4/sub_412/carry [8]), .A2(n4439), .ZN(
        \u4/sub_412/carry [9]) );
  XOR2_X1 U4104 ( .A(n4439), .B(\u4/sub_412/carry [8]), .Z(\u4/div_shft4 [8])
         );
  OR2_X1 U4105 ( .A1(n4353), .A2(\sub_1_root_sub_0_root_u4/add_497/carry [8]), 
        .ZN(\sub_1_root_sub_0_root_u4/add_497/carry [9]) );
  XNOR2_X1 U4106 ( .A(\sub_1_root_sub_0_root_u4/add_497/carry [8]), .B(n4353), 
        .ZN(\u4/ldz_dif[8] ) );
  AND2_X1 U4107 ( .A1(n4281), .A2(\u4/add_410/carry [7]), .ZN(
        \u4/add_410/carry [8]) );
  XOR2_X1 U4108 ( .A(n4281), .B(\u4/add_410/carry [7]), .Z(\u4/div_shft2 [7])
         );
  AND2_X1 U4109 ( .A1(n4281), .A2(\u4/add_411/carry [7]), .ZN(
        \u4/add_411/carry [8]) );
  XOR2_X1 U4110 ( .A(n4281), .B(\u4/add_411/carry [7]), .Z(\u4/div_shft3[7] )
         );
  AND2_X1 U4111 ( .A1(\u4/sub_412/carry [7]), .A2(n4348), .ZN(
        \u4/sub_412/carry [8]) );
  XOR2_X1 U4112 ( .A(n4348), .B(\u4/sub_412/carry [7]), .Z(\u4/div_shft4 [7])
         );
  OR2_X1 U4113 ( .A1(n4281), .A2(\sub_1_root_sub_0_root_u4/add_497/carry [7]), 
        .ZN(\sub_1_root_sub_0_root_u4/add_497/carry [8]) );
  XNOR2_X1 U4114 ( .A(\sub_1_root_sub_0_root_u4/add_497/carry [7]), .B(n4281), 
        .ZN(\u4/ldz_dif[7] ) );
  AND2_X1 U4115 ( .A1(exp_r[6]), .A2(\u4/add_410/carry [6]), .ZN(
        \u4/add_410/carry [7]) );
  XOR2_X1 U4116 ( .A(exp_r[6]), .B(\u4/add_410/carry [6]), .Z(
        \u4/div_shft2 [6]) );
  AND2_X1 U4117 ( .A1(n4290), .A2(\u4/add_410/carry [5]), .ZN(
        \u4/add_410/carry [6]) );
  XOR2_X1 U4118 ( .A(n4290), .B(\u4/add_410/carry [5]), .Z(\u4/div_shft2 [5])
         );
  AND2_X1 U4119 ( .A1(n4282), .A2(\u4/add_410/carry [4]), .ZN(
        \u4/add_410/carry [5]) );
  XOR2_X1 U4120 ( .A(n4282), .B(\u4/add_410/carry [4]), .Z(\u4/div_shft2 [4])
         );
  AND2_X1 U4121 ( .A1(n4655), .A2(\u4/add_410/carry [3]), .ZN(
        \u4/add_410/carry [4]) );
  XOR2_X1 U4122 ( .A(exp_r[3]), .B(\u4/add_410/carry [3]), .Z(
        \u4/div_shft2 [3]) );
  AND2_X1 U4123 ( .A1(n4315), .A2(exp_r[1]), .ZN(\u4/add_410/carry [3]) );
  XOR2_X1 U4124 ( .A(n4315), .B(exp_r[1]), .Z(\u4/div_shft2 [2]) );
  AND2_X1 U4125 ( .A1(exp_r[6]), .A2(\u4/add_411/carry [6]), .ZN(
        \u4/add_411/carry [7]) );
  XOR2_X1 U4126 ( .A(exp_r[6]), .B(\u4/add_411/carry [6]), .Z(
        \u4/div_shft3[6] ) );
  AND2_X1 U4127 ( .A1(n4290), .A2(\u4/add_411/carry [5]), .ZN(
        \u4/add_411/carry [6]) );
  XOR2_X1 U4128 ( .A(n4290), .B(\u4/add_411/carry [5]), .Z(\u4/div_shft3[5] )
         );
  AND2_X1 U4129 ( .A1(n4600), .A2(div_opa_ldz_r2[0]), .ZN(
        \u4/add_411/carry [1]) );
  XOR2_X1 U4130 ( .A(n4600), .B(div_opa_ldz_r2[0]), .Z(\u4/div_shft3[0] ) );
  XNOR2_X1 U4131 ( .A(\u4/sub_409/carry [10]), .B(n4656), .ZN(
        \u4/div_scht1a [10]) );
  OR2_X1 U4132 ( .A1(n4289), .A2(\u4/sub_409/carry [9]), .ZN(
        \u4/sub_409/carry [10]) );
  XNOR2_X1 U4133 ( .A(\u4/sub_409/carry [9]), .B(n4289), .ZN(
        \u4/div_scht1a [9]) );
  OR2_X1 U4134 ( .A1(n4353), .A2(\u4/sub_409/carry [8]), .ZN(
        \u4/sub_409/carry [9]) );
  XNOR2_X1 U4135 ( .A(\u4/sub_409/carry [8]), .B(n4353), .ZN(
        \u4/div_scht1a [8]) );
  OR2_X1 U4136 ( .A1(n4281), .A2(\u4/sub_409/carry [7]), .ZN(
        \u4/sub_409/carry [8]) );
  XNOR2_X1 U4137 ( .A(\u4/sub_409/carry [7]), .B(n4281), .ZN(
        \u4/div_scht1a [7]) );
  OR2_X1 U4138 ( .A1(exp_r[6]), .A2(\u4/sub_409/carry [6]), .ZN(
        \u4/sub_409/carry [7]) );
  XNOR2_X1 U4139 ( .A(\u4/sub_409/carry [6]), .B(exp_r[6]), .ZN(
        \u4/div_scht1a [6]) );
  OR2_X1 U4140 ( .A1(n4290), .A2(\u4/sub_409/carry [5]), .ZN(
        \u4/sub_409/carry [6]) );
  XNOR2_X1 U4141 ( .A(\u4/sub_409/carry [5]), .B(n4290), .ZN(
        \u4/div_scht1a [5]) );
  OR2_X1 U4142 ( .A1(n4447), .A2(n4600), .ZN(\u4/sub_409/carry [1]) );
  XNOR2_X1 U4143 ( .A(n4600), .B(n4447), .ZN(\u4/div_scht1a [0]) );
  AND2_X1 U4144 ( .A1(\u4/sub_412/carry [6]), .A2(n4317), .ZN(
        \u4/sub_412/carry [7]) );
  XOR2_X1 U4145 ( .A(n4317), .B(\u4/sub_412/carry [6]), .Z(\u4/div_shft4 [6])
         );
  AND2_X1 U4146 ( .A1(\u4/sub_412/carry [5]), .A2(n4347), .ZN(
        \u4/sub_412/carry [6]) );
  XOR2_X1 U4147 ( .A(n4347), .B(\u4/sub_412/carry [5]), .Z(\u4/div_shft4 [5])
         );
  OR2_X1 U4148 ( .A1(n4349), .A2(div_opa_ldz_r2[0]), .ZN(\u4/sub_412/carry [1]) );
  XNOR2_X1 U4149 ( .A(div_opa_ldz_r2[0]), .B(n4349), .ZN(\u4/div_shft4 [0]) );
  XNOR2_X1 U4150 ( .A(n4656), .B(\u4/sub_417/carry[10] ), .ZN(
        \u4/f2i_shft[10] ) );
  OR2_X1 U4151 ( .A1(n4289), .A2(\u4/sub_417/carry[9] ), .ZN(
        \u4/sub_417/carry[10] ) );
  XNOR2_X1 U4152 ( .A(\u4/sub_417/carry[9] ), .B(n4289), .ZN(\u4/f2i_shft[9] )
         );
  OR2_X1 U4153 ( .A1(n4353), .A2(\u4/sub_417/carry[8] ), .ZN(
        \u4/sub_417/carry[9] ) );
  XNOR2_X1 U4154 ( .A(\u4/sub_417/carry[8] ), .B(n4353), .ZN(\u4/f2i_shft[8] )
         );
  OR2_X1 U4155 ( .A1(n4281), .A2(\u4/sub_417/carry[7] ), .ZN(
        \u4/sub_417/carry[8] ) );
  XNOR2_X1 U4156 ( .A(\u4/sub_417/carry[7] ), .B(n4281), .ZN(\u4/f2i_shft[7] )
         );
  AND2_X1 U4157 ( .A1(\u4/sub_417/carry[6] ), .A2(exp_r[6]), .ZN(
        \u4/sub_417/carry[7] ) );
  XOR2_X1 U4158 ( .A(exp_r[6]), .B(\u4/sub_417/carry[6] ), .Z(\u4/f2i_shft[6] ) );
  AND2_X1 U4159 ( .A1(\u4/sub_417/carry[5] ), .A2(n4290), .ZN(
        \u4/sub_417/carry[6] ) );
  XOR2_X1 U4160 ( .A(n4290), .B(\u4/sub_417/carry[5] ), .Z(\u4/f2i_shft[5] )
         );
  AND2_X1 U4161 ( .A1(\u4/sub_417/carry[4] ), .A2(n4282), .ZN(
        \u4/sub_417/carry[5] ) );
  XOR2_X1 U4162 ( .A(n4282), .B(\u4/sub_417/carry[4] ), .Z(\u4/f2i_shft[4] )
         );
  AND2_X1 U4163 ( .A1(\u4/sub_417/carry[3] ), .A2(n4655), .ZN(
        \u4/sub_417/carry[4] ) );
  XOR2_X1 U4164 ( .A(n4655), .B(\u4/sub_417/carry[3] ), .Z(\u4/f2i_shft[3] )
         );
  AND2_X1 U4165 ( .A1(\u4/sub_417/carry[2] ), .A2(n4315), .ZN(
        \u4/sub_417/carry[3] ) );
  XOR2_X1 U4166 ( .A(n4315), .B(\u4/sub_417/carry[2] ), .Z(\u4/f2i_shft[2] )
         );
  OR2_X1 U4167 ( .A1(exp_r[1]), .A2(n4600), .ZN(\u4/sub_417/carry[2] ) );
  XNOR2_X1 U4168 ( .A(n4600), .B(exp_r[1]), .ZN(\u4/f2i_shft[1] ) );
  AND2_X1 U4169 ( .A1(\u4/sub_481/carry [6]), .A2(n4663), .ZN(\u4/N6142 ) );
  XOR2_X1 U4170 ( .A(n4663), .B(\u4/sub_481/carry [6]), .Z(\u4/N6141 ) );
  AND2_X1 U4171 ( .A1(\u4/sub_481/carry [5]), .A2(n4664), .ZN(
        \u4/sub_481/carry [6]) );
  XOR2_X1 U4172 ( .A(n4664), .B(\u4/sub_481/carry [5]), .Z(\u4/N6140 ) );
  OR2_X1 U4173 ( .A1(n4665), .A2(\u4/sub_481/carry [4]), .ZN(
        \u4/sub_481/carry [5]) );
  XNOR2_X1 U4174 ( .A(\u4/sub_481/carry [4]), .B(n4665), .ZN(\u4/N6139 ) );
  OR2_X1 U4175 ( .A1(n4714), .A2(\u4/sub_481/carry [3]), .ZN(
        \u4/sub_481/carry [4]) );
  XNOR2_X1 U4176 ( .A(\u4/sub_481/carry [3]), .B(n4714), .ZN(\u4/N6138 ) );
  OR2_X1 U4177 ( .A1(n4715), .A2(\u4/sub_481/carry [2]), .ZN(
        \u4/sub_481/carry [3]) );
  XNOR2_X1 U4178 ( .A(\u4/sub_481/carry [2]), .B(n4715), .ZN(\u4/N6137 ) );
  OR2_X1 U4179 ( .A1(n4666), .A2(\u4/fi_ldz_mi1[0] ), .ZN(
        \u4/sub_481/carry [2]) );
  XNOR2_X1 U4180 ( .A(\u4/fi_ldz_mi1[0] ), .B(n4666), .ZN(\u4/N6136 ) );
  OR2_X1 U4181 ( .A1(exp_r[6]), .A2(
        \sub_1_root_sub_0_root_u4/add_497/carry [6]), .ZN(
        \sub_1_root_sub_0_root_u4/add_497/carry [7]) );
  XNOR2_X1 U4182 ( .A(\sub_1_root_sub_0_root_u4/add_497/carry [6]), .B(
        exp_r[6]), .ZN(\u4/ldz_dif[6] ) );
  OR2_X1 U4183 ( .A1(n4290), .A2(\sub_1_root_sub_0_root_u4/add_497/carry [5]), 
        .ZN(\sub_1_root_sub_0_root_u4/add_497/carry [6]) );
  XNOR2_X1 U4184 ( .A(\sub_1_root_sub_0_root_u4/add_497/carry [5]), .B(n4290), 
        .ZN(\u4/ldz_dif[5] ) );
  OR2_X1 U4185 ( .A1(n4447), .A2(n4600), .ZN(
        \sub_1_root_sub_0_root_u4/add_497/carry [1]) );
  XNOR2_X1 U4186 ( .A(n4600), .B(n4447), .ZN(\u4/ldz_dif[0] ) );
  XOR2_X1 U4187 ( .A(n4663), .B(\u4/sub_491/carry [6]), .Z(\u4/fi_ldz_2a[6] )
         );
  OR2_X1 U4188 ( .A1(n4664), .A2(\u4/sub_491/carry [5]), .ZN(
        \u4/sub_491/carry [6]) );
  XNOR2_X1 U4189 ( .A(\u4/sub_491/carry [5]), .B(n4664), .ZN(\u4/fi_ldz_2a[5] ) );
  OR2_X1 U4190 ( .A1(n4665), .A2(\u4/sub_491/carry [4]), .ZN(
        \u4/sub_491/carry [5]) );
  XNOR2_X1 U4191 ( .A(\u4/sub_491/carry [4]), .B(n4665), .ZN(\u4/fi_ldz_2a[4] ) );
  AND2_X1 U4192 ( .A1(\u4/sub_491/carry [3]), .A2(n4714), .ZN(
        \u4/sub_491/carry [4]) );
  XOR2_X1 U4193 ( .A(n4714), .B(\u4/sub_491/carry [3]), .Z(\u4/fi_ldz_2a[3] )
         );
  OR2_X1 U4194 ( .A1(n4715), .A2(\u4/sub_491/carry [2]), .ZN(
        \u4/sub_491/carry [3]) );
  XNOR2_X1 U4195 ( .A(\u4/sub_491/carry [2]), .B(n4715), .ZN(\u4/fi_ldz_2a[2] ) );
  AND2_X1 U4196 ( .A1(\u4/fi_ldz_mi1[0] ), .A2(n4666), .ZN(
        \u4/sub_491/carry [2]) );
  XOR2_X1 U4197 ( .A(n4666), .B(\u4/fi_ldz_mi1[0] ), .Z(\u4/fi_ldz_2a[1] ) );
  XNOR2_X1 U4198 ( .A(\u2/gt_145/B[11] ), .B(\u2/sub_116/carry[11] ), .ZN(
        \u2/N53 ) );
  OR2_X1 U4199 ( .A1(\u2/exp_tmp4[10] ), .A2(\u2/sub_116/carry[10] ), .ZN(
        \u2/sub_116/carry[11] ) );
  XNOR2_X1 U4200 ( .A(\u2/sub_116/carry[10] ), .B(\u2/exp_tmp4[10] ), .ZN(
        \u2/N52 ) );
  AND2_X1 U4201 ( .A1(\u2/sub_116/carry[9] ), .A2(\u2/lt_135/A[9] ), .ZN(
        \u2/sub_116/carry[10] ) );
  XOR2_X1 U4202 ( .A(\u2/lt_135/A[9] ), .B(\u2/sub_116/carry[9] ), .Z(\u2/N51 ) );
  AND2_X1 U4203 ( .A1(\u2/sub_116/carry[8] ), .A2(\u2/lt_135/A[8] ), .ZN(
        \u2/sub_116/carry[9] ) );
  XOR2_X1 U4204 ( .A(\u2/lt_135/A[8] ), .B(\u2/sub_116/carry[8] ), .Z(\u2/N50 ) );
  AND2_X1 U4205 ( .A1(\u2/sub_116/carry[7] ), .A2(\u2/lt_135/A[7] ), .ZN(
        \u2/sub_116/carry[8] ) );
  XOR2_X1 U4206 ( .A(\u2/lt_135/A[7] ), .B(\u2/sub_116/carry[7] ), .Z(\u2/N49 ) );
  AND2_X1 U4207 ( .A1(\u2/sub_116/carry[6] ), .A2(\u2/lt_135/A[6] ), .ZN(
        \u2/sub_116/carry[7] ) );
  XOR2_X1 U4208 ( .A(\u2/lt_135/A[6] ), .B(\u2/sub_116/carry[6] ), .Z(\u2/N48 ) );
  AND2_X1 U4209 ( .A1(\u2/sub_116/carry[5] ), .A2(\u2/lt_135/A[5] ), .ZN(
        \u2/sub_116/carry[6] ) );
  XOR2_X1 U4210 ( .A(\u2/lt_135/A[5] ), .B(\u2/sub_116/carry[5] ), .Z(\u2/N47 ) );
  AND2_X1 U4211 ( .A1(\u2/sub_116/carry[4] ), .A2(\u2/exp_tmp1[4] ), .ZN(
        \u2/sub_116/carry[5] ) );
  XOR2_X1 U4212 ( .A(\u2/exp_tmp1[4] ), .B(\u2/sub_116/carry[4] ), .Z(\u2/N46 ) );
  AND2_X1 U4213 ( .A1(\u2/sub_116/carry[3] ), .A2(\u2/exp_tmp1[3] ), .ZN(
        \u2/sub_116/carry[4] ) );
  XOR2_X1 U4214 ( .A(\u2/exp_tmp1[3] ), .B(\u2/sub_116/carry[3] ), .Z(\u2/N45 ) );
  AND2_X1 U4215 ( .A1(\u2/sub_116/carry[2] ), .A2(\u2/exp_tmp1[2] ), .ZN(
        \u2/sub_116/carry[3] ) );
  XOR2_X1 U4216 ( .A(\u2/exp_tmp1[2] ), .B(\u2/sub_116/carry[2] ), .Z(\u2/N44 ) );
  AND2_X1 U4217 ( .A1(\u2/lt_135/A[0] ), .A2(\u2/exp_tmp1[1] ), .ZN(
        \u2/sub_116/carry[2] ) );
  XOR2_X1 U4218 ( .A(\u2/exp_tmp1[1] ), .B(\u2/lt_135/A[0] ), .Z(\u2/N43 ) );
  XOR2_X1 U4219 ( .A(\u2/gt_145/B[11] ), .B(\u2/add_116/carry[11] ), .Z(
        \u2/N41 ) );
  AND2_X1 U4220 ( .A1(\u2/add_116/carry[10] ), .A2(\u2/exp_tmp4[10] ), .ZN(
        \u2/add_116/carry[11] ) );
  XOR2_X1 U4221 ( .A(\u2/exp_tmp4[10] ), .B(\u2/add_116/carry[10] ), .Z(
        \u2/N40 ) );
  OR2_X1 U4222 ( .A1(\u2/lt_135/A[9] ), .A2(\u2/add_116/carry[9] ), .ZN(
        \u2/add_116/carry[10] ) );
  XNOR2_X1 U4223 ( .A(\u2/add_116/carry[9] ), .B(\u2/lt_135/A[9] ), .ZN(
        \u2/N39 ) );
  OR2_X1 U4224 ( .A1(\u2/lt_135/A[8] ), .A2(\u2/add_116/carry[8] ), .ZN(
        \u2/add_116/carry[9] ) );
  XNOR2_X1 U4225 ( .A(\u2/add_116/carry[8] ), .B(\u2/lt_135/A[8] ), .ZN(
        \u2/N38 ) );
  OR2_X1 U4226 ( .A1(\u2/lt_135/A[7] ), .A2(\u2/add_116/carry[7] ), .ZN(
        \u2/add_116/carry[8] ) );
  XNOR2_X1 U4227 ( .A(\u2/add_116/carry[7] ), .B(\u2/lt_135/A[7] ), .ZN(
        \u2/N37 ) );
  OR2_X1 U4228 ( .A1(\u2/lt_135/A[6] ), .A2(\u2/add_116/carry[6] ), .ZN(
        \u2/add_116/carry[7] ) );
  XNOR2_X1 U4229 ( .A(\u2/add_116/carry[6] ), .B(\u2/lt_135/A[6] ), .ZN(
        \u2/N36 ) );
  OR2_X1 U4230 ( .A1(\u2/lt_135/A[5] ), .A2(\u2/add_116/carry[5] ), .ZN(
        \u2/add_116/carry[6] ) );
  XNOR2_X1 U4231 ( .A(\u2/add_116/carry[5] ), .B(\u2/lt_135/A[5] ), .ZN(
        \u2/N35 ) );
  OR2_X1 U4232 ( .A1(\u2/exp_tmp1[4] ), .A2(\u2/add_116/carry[4] ), .ZN(
        \u2/add_116/carry[5] ) );
  XNOR2_X1 U4233 ( .A(\u2/add_116/carry[4] ), .B(\u2/exp_tmp1[4] ), .ZN(
        \u2/N34 ) );
  OR2_X1 U4234 ( .A1(\u2/exp_tmp1[3] ), .A2(\u2/add_116/carry[3] ), .ZN(
        \u2/add_116/carry[4] ) );
  XNOR2_X1 U4235 ( .A(\u2/add_116/carry[3] ), .B(\u2/exp_tmp1[3] ), .ZN(
        \u2/N33 ) );
  OR2_X1 U4236 ( .A1(\u2/exp_tmp1[2] ), .A2(\u2/add_116/carry[2] ), .ZN(
        \u2/add_116/carry[3] ) );
  XNOR2_X1 U4237 ( .A(\u2/add_116/carry[2] ), .B(\u2/exp_tmp1[2] ), .ZN(
        \u2/N32 ) );
  OR2_X1 U4238 ( .A1(\u2/exp_tmp1[1] ), .A2(\u2/lt_135/A[0] ), .ZN(
        \u2/add_116/carry[2] ) );
  XNOR2_X1 U4239 ( .A(\u2/lt_135/A[0] ), .B(\u2/exp_tmp1[1] ), .ZN(\u2/N31 )
         );
  INV_X4 U4240 ( .A(\u4/fi_ldz[6] ), .ZN(n4663) );
  INV_X4 U4241 ( .A(\u4/fi_ldz[5] ), .ZN(n4664) );
  INV_X4 U4242 ( .A(\u4/fi_ldz[4] ), .ZN(n4665) );
  INV_X4 U4243 ( .A(\u4/fi_ldz[1] ), .ZN(n4666) );
  INV_X4 U4244 ( .A(\u2/exp_tmp1[1] ), .ZN(\u2/exp_tmp4[1] ) );
  INV_X4 U4245 ( .A(\u2/exp_tmp1[2] ), .ZN(\u2/exp_tmp4[2] ) );
  INV_X4 U4246 ( .A(\u2/exp_tmp1[3] ), .ZN(\u2/exp_tmp4[3] ) );
  INV_X4 U4247 ( .A(\u2/exp_tmp1[4] ), .ZN(\u2/exp_tmp4[4] ) );
  NOR2_X1 U4248 ( .A1(\u2/exp_tmp4[1] ), .A2(n2800), .ZN(n4668) );
  NOR2_X1 U4249 ( .A1(n4677), .A2(\u2/exp_tmp4[2] ), .ZN(n4669) );
  NOR2_X1 U4250 ( .A1(n4678), .A2(\u2/exp_tmp4[3] ), .ZN(n4670) );
  NOR2_X1 U4251 ( .A1(n4378), .A2(n2799), .ZN(n4672) );
  NAND2_X1 U4252 ( .A1(n4672), .A2(\u2/lt_135/A[6] ), .ZN(n4673) );
  NOR2_X1 U4253 ( .A1(n4673), .A2(n2797), .ZN(n4675) );
  NAND2_X1 U4254 ( .A1(n4675), .A2(\u2/lt_135/A[8] ), .ZN(n4676) );
  NOR2_X1 U4255 ( .A1(n2795), .A2(n4676), .ZN(n4667) );
  XOR2_X1 U4256 ( .A(\u2/exp_tmp4[10] ), .B(n4667), .Z(\u2/N75 ) );
  OAI21_X1 U4257 ( .B1(\u2/lt_135/A[0] ), .B2(\u2/exp_tmp1[1] ), .A(n4677), 
        .ZN(\u2/N66 ) );
  OAI21_X1 U4258 ( .B1(n4668), .B2(\u2/exp_tmp1[2] ), .A(n4678), .ZN(\u2/N67 )
         );
  OAI21_X1 U4259 ( .B1(n4669), .B2(\u2/exp_tmp1[3] ), .A(n4679), .ZN(\u2/N68 )
         );
  OAI21_X1 U4260 ( .B1(n4670), .B2(\u2/exp_tmp1[4] ), .A(n4378), .ZN(\u2/N69 )
         );
  AOI21_X1 U4261 ( .B1(n4378), .B2(n2799), .A(n4672), .ZN(n4671) );
  OAI21_X1 U4262 ( .B1(n4672), .B2(\u2/lt_135/A[6] ), .A(n4673), .ZN(\u2/N71 )
         );
  AOI21_X1 U4263 ( .B1(n4673), .B2(n2797), .A(n4675), .ZN(n4674) );
  OAI21_X1 U4264 ( .B1(n4675), .B2(\u2/lt_135/A[8] ), .A(n4676), .ZN(\u2/N73 )
         );
  XNOR2_X1 U4265 ( .A(n2795), .B(n4676), .ZN(\u2/N74 ) );
  INV_X4 U4266 ( .A(n4668), .ZN(n4677) );
  INV_X4 U4267 ( .A(n4669), .ZN(n4678) );
  INV_X4 U4268 ( .A(n4670), .ZN(n4679) );
  INV_X4 U4269 ( .A(n4671), .ZN(\u2/N70 ) );
  INV_X4 U4270 ( .A(n4674), .ZN(\u2/N72 ) );
  NOR2_X1 U4271 ( .A1(exp_r[1]), .A2(n4600), .ZN(n4681) );
  NOR2_X1 U4272 ( .A1(\u4/sub_417/carry[2] ), .A2(n4315), .ZN(n4682) );
  NOR2_X1 U4273 ( .A1(n4689), .A2(n4655), .ZN(n4683) );
  NOR2_X1 U4274 ( .A1(n4690), .A2(n4282), .ZN(n4684) );
  NOR2_X1 U4275 ( .A1(n4691), .A2(n4290), .ZN(n4685) );
  NOR2_X1 U4276 ( .A1(n4354), .A2(n4281), .ZN(n4687) );
  NAND2_X1 U4277 ( .A1(n4687), .A2(n4439), .ZN(n4688) );
  NOR3_X1 U4278 ( .A1(n4352), .A2(n4289), .A3(n4688), .ZN(\u4/exp_in_mi1[11] )
         );
  OAI21_X1 U4279 ( .B1(n4289), .B2(n4688), .A(n4352), .ZN(n4680) );
  NAND2_X1 U4280 ( .A1(n6460), .A2(n4680), .ZN(\u4/exp_in_mi1[10] ) );
  OAI21_X1 U4281 ( .B1(n4349), .B2(n4314), .A(\u4/sub_417/carry[2] ), .ZN(
        \u4/exp_in_mi1[1] ) );
  OAI21_X1 U4282 ( .B1(n4681), .B2(n4438), .A(n4689), .ZN(\u4/exp_in_mi1[2] )
         );
  OAI21_X1 U4283 ( .B1(n4682), .B2(n4316), .A(n4690), .ZN(\u4/exp_in_mi1[3] )
         );
  OAI21_X1 U4284 ( .B1(n4683), .B2(n4299), .A(n4691), .ZN(\u4/exp_in_mi1[4] )
         );
  OAI21_X1 U4285 ( .B1(n4684), .B2(n4347), .A(n4692), .ZN(\u4/exp_in_mi1[5] )
         );
  OAI21_X1 U4286 ( .B1(n4685), .B2(n4317), .A(n4354), .ZN(\u4/exp_in_mi1[6] )
         );
  AOI21_X1 U4287 ( .B1(n4354), .B2(n4281), .A(n4687), .ZN(n4686) );
  OAI21_X1 U4288 ( .B1(n4687), .B2(n4439), .A(n4688), .ZN(\u4/exp_in_mi1[8] )
         );
  XNOR2_X1 U4289 ( .A(n4289), .B(n4688), .ZN(\u4/exp_in_mi1[9] ) );
  INV_X4 U4290 ( .A(n4682), .ZN(n4689) );
  INV_X4 U4291 ( .A(n4683), .ZN(n4690) );
  INV_X4 U4292 ( .A(n4684), .ZN(n4691) );
  INV_X4 U4293 ( .A(n4685), .ZN(n4692) );
  INV_X4 U4294 ( .A(n4686), .ZN(\u4/exp_in_mi1[7] ) );
  NOR2_X1 U4295 ( .A1(\u4/fi_ldz[1] ), .A2(\u4/fi_ldz_2a[0] ), .ZN(n4694) );
  AOI21_X1 U4296 ( .B1(\u4/fi_ldz_2a[0] ), .B2(\u4/fi_ldz[1] ), .A(n4694), 
        .ZN(n4693) );
  NAND2_X1 U4297 ( .A1(n4694), .A2(n4715), .ZN(n4695) );
  OAI21_X1 U4298 ( .B1(n4694), .B2(n4715), .A(n4695), .ZN(\u4/fi_ldz_mi1[2] )
         );
  NOR2_X1 U4299 ( .A1(n4695), .A2(\u4/fi_ldz[3] ), .ZN(n4697) );
  AOI21_X1 U4300 ( .B1(n4695), .B2(\u4/fi_ldz[3] ), .A(n4697), .ZN(n4696) );
  NAND2_X1 U4301 ( .A1(n4697), .A2(n4665), .ZN(n4698) );
  OAI21_X1 U4302 ( .B1(n4697), .B2(n4665), .A(n4698), .ZN(\u4/fi_ldz_mi1[4] )
         );
  XNOR2_X1 U4303 ( .A(\u4/fi_ldz[5] ), .B(n4698), .ZN(\u4/fi_ldz_mi1[5] ) );
  NOR2_X1 U4304 ( .A1(\u4/fi_ldz[5] ), .A2(n4698), .ZN(n4699) );
  XOR2_X1 U4305 ( .A(\u4/fi_ldz[6] ), .B(n4699), .Z(\u4/fi_ldz_mi1[6] ) );
  INV_X4 U4306 ( .A(\u4/fi_ldz_2a[0] ), .ZN(\u4/fi_ldz_mi1[0] ) );
  INV_X4 U4307 ( .A(n4693), .ZN(\u4/fi_ldz_mi1[1] ) );
  INV_X4 U4308 ( .A(n4696), .ZN(\u4/fi_ldz_mi1[3] ) );
  NOR2_X1 U4309 ( .A1(\u4/exp_out1[1] ), .A2(\u4/exp_out1[0] ), .ZN(n4701) );
  NOR2_X1 U4310 ( .A1(n4710), .A2(\u4/sub_468/A[2] ), .ZN(n4702) );
  NOR2_X1 U4311 ( .A1(n4712), .A2(\u4/sub_468/A[3] ), .ZN(n4703) );
  NOR2_X1 U4312 ( .A1(n4339), .A2(\u4/sub_468/A[5] ), .ZN(n4705) );
  NAND2_X1 U4313 ( .A1(n4705), .A2(n2418), .ZN(n4706) );
  NOR2_X1 U4314 ( .A1(n4706), .A2(\u4/sub_468/A[7] ), .ZN(n4708) );
  NAND2_X1 U4315 ( .A1(n4708), .A2(n2424), .ZN(n4709) );
  NOR2_X1 U4316 ( .A1(\u4/sub_468/A[9] ), .A2(n4709), .ZN(n4700) );
  XOR2_X1 U4317 ( .A(\u4/sub_468/A[10] ), .B(n4700), .Z(\u4/exp_out1_mi1 [10])
         );
  OAI21_X1 U4318 ( .B1(\u4/exp_out1_mi1 [0]), .B2(n4711), .A(n4710), .ZN(
        \u4/exp_out1_mi1 [1]) );
  OAI21_X1 U4319 ( .B1(n4701), .B2(n2407), .A(n4712), .ZN(\u4/exp_out1_mi1 [2]) );
  OAI21_X1 U4320 ( .B1(n4702), .B2(n2411), .A(n4713), .ZN(\u4/exp_out1_mi1 [3]) );
  OAI21_X1 U4321 ( .B1(n4703), .B2(n2414), .A(n4339), .ZN(\u4/exp_out1_mi1 [4]) );
  AOI21_X1 U4322 ( .B1(n4339), .B2(\u4/sub_468/A[5] ), .A(n4705), .ZN(n4704)
         );
  OAI21_X1 U4323 ( .B1(n4705), .B2(n2418), .A(n4706), .ZN(\u4/exp_out1_mi1 [6]) );
  AOI21_X1 U4324 ( .B1(n4706), .B2(\u4/sub_468/A[7] ), .A(n4708), .ZN(n4707)
         );
  OAI21_X1 U4325 ( .B1(n4708), .B2(n2424), .A(n4709), .ZN(\u4/exp_out1_mi1 [8]) );
  XNOR2_X1 U4326 ( .A(\u4/sub_468/A[9] ), .B(n4709), .ZN(\u4/exp_out1_mi1 [9])
         );
  INV_X4 U4327 ( .A(\u4/exp_out1[0] ), .ZN(\u4/exp_out1_mi1 [0]) );
  INV_X4 U4328 ( .A(n4701), .ZN(n4710) );
  INV_X4 U4329 ( .A(\u4/exp_out1[1] ), .ZN(n4711) );
  INV_X4 U4330 ( .A(n4702), .ZN(n4712) );
  INV_X4 U4331 ( .A(n4703), .ZN(n4713) );
  INV_X4 U4332 ( .A(n4704), .ZN(\u4/exp_out1_mi1 [5]) );
  INV_X4 U4333 ( .A(n4707), .ZN(\u4/exp_out1_mi1 [7]) );
  INV_X4 U4334 ( .A(\u4/fi_ldz[3] ), .ZN(n4714) );
  INV_X4 U4335 ( .A(\u4/fi_ldz[2] ), .ZN(n4715) );
  INV_X1 U4336 ( .A(\u4/exp_out[0] ), .ZN(\u4/exp_out_mi1 [0]) );
  NOR2_X1 U4337 ( .A1(\u4/exp_out[1] ), .A2(\u4/exp_out[0] ), .ZN(n4719) );
  INV_X1 U4338 ( .A(n4719), .ZN(n4717) );
  NOR2_X1 U4339 ( .A1(n4717), .A2(\u4/exp_out[2] ), .ZN(n4721) );
  INV_X1 U4340 ( .A(n4721), .ZN(n4718) );
  NOR2_X1 U4341 ( .A1(n4718), .A2(\u4/exp_out[3] ), .ZN(n4722) );
  INV_X1 U4342 ( .A(n4722), .ZN(n4720) );
  NOR2_X1 U4343 ( .A1(n4337), .A2(\u4/exp_out[5] ), .ZN(n4724) );
  NAND2_X1 U4344 ( .A1(n4724), .A2(n2456), .ZN(n4725) );
  NOR2_X1 U4345 ( .A1(n4725), .A2(\u4/exp_out[7] ), .ZN(n4727) );
  NAND2_X1 U4346 ( .A1(n4727), .A2(n2450), .ZN(n4728) );
  NOR2_X1 U4347 ( .A1(\u4/exp_out[9] ), .A2(n4728), .ZN(n4716) );
  XOR2_X1 U4348 ( .A(\u4/exp_out[10] ), .B(n4716), .Z(\u4/exp_out_mi1 [10]) );
  OAI21_X1 U4349 ( .B1(\u4/exp_out_mi1 [0]), .B2(n2471), .A(n4717), .ZN(
        \u4/exp_out_mi1 [1]) );
  OAI21_X1 U4350 ( .B1(n4719), .B2(n2468), .A(n4718), .ZN(\u4/exp_out_mi1 [2])
         );
  OAI21_X1 U4351 ( .B1(n4721), .B2(n2465), .A(n4720), .ZN(\u4/exp_out_mi1 [3])
         );
  OAI21_X1 U4352 ( .B1(n4722), .B2(n2462), .A(n4337), .ZN(\u4/exp_out_mi1 [4])
         );
  AOI21_X1 U4353 ( .B1(n4337), .B2(\u4/exp_out[5] ), .A(n4724), .ZN(n4723) );
  INV_X1 U4354 ( .A(n4723), .ZN(\u4/exp_out_mi1 [5]) );
  OAI21_X1 U4355 ( .B1(n4724), .B2(n2456), .A(n4725), .ZN(\u4/exp_out_mi1 [6])
         );
  AOI21_X1 U4356 ( .B1(n4725), .B2(\u4/exp_out[7] ), .A(n4727), .ZN(n4726) );
  INV_X1 U4357 ( .A(n4726), .ZN(\u4/exp_out_mi1 [7]) );
  OAI21_X1 U4358 ( .B1(n4727), .B2(n2450), .A(n4728), .ZN(\u4/exp_out_mi1 [8])
         );
  XNOR2_X1 U4359 ( .A(\u4/exp_out[9] ), .B(n4728), .ZN(\u4/exp_out_mi1 [9]) );
  NAND2_X1 U4360 ( .A1(opb_r[54]), .A2(n4451), .ZN(n4745) );
  NAND2_X1 U4361 ( .A1(opb_r[59]), .A2(n4442), .ZN(n4747) );
  NAND2_X1 U4362 ( .A1(opb_r[60]), .A2(n4357), .ZN(n4748) );
  NAND2_X1 U4363 ( .A1(opb_r[57]), .A2(n4453), .ZN(n4742) );
  NAND2_X1 U4364 ( .A1(opb_r[58]), .A2(n4454), .ZN(n4740) );
  NAND2_X1 U4365 ( .A1(opb_r[55]), .A2(n4358), .ZN(n4741) );
  NAND2_X1 U4366 ( .A1(opb_r[56]), .A2(n4456), .ZN(n4744) );
  NOR2_X1 U4367 ( .A1(n4449), .A2(opb_r[52]), .ZN(n4730) );
  OAI21_X1 U4368 ( .B1(n4756), .B2(n4450), .A(opb_r[53]), .ZN(n4729) );
  OAI211_X1 U4369 ( .C1(opa_r[53]), .C2(n4730), .A(n4729), .B(n4745), .ZN(
        n4731) );
  OAI221_X1 U4370 ( .B1(opb_r[54]), .B2(n4451), .C1(opb_r[55]), .C2(n4358), 
        .A(n4731), .ZN(n4732) );
  NAND3_X1 U4371 ( .A1(n4741), .A2(n4744), .A3(n4732), .ZN(n4733) );
  OAI221_X1 U4372 ( .B1(opb_r[56]), .B2(n4456), .C1(opb_r[57]), .C2(n4453), 
        .A(n4733), .ZN(n4734) );
  NAND3_X1 U4373 ( .A1(n4742), .A2(n4740), .A3(n4734), .ZN(n4735) );
  OAI221_X1 U4374 ( .B1(opb_r[58]), .B2(n4454), .C1(opb_r[59]), .C2(n4442), 
        .A(n4735), .ZN(n4736) );
  NAND3_X1 U4375 ( .A1(n4747), .A2(n4748), .A3(n4736), .ZN(n4737) );
  OAI221_X1 U4376 ( .B1(opb_r[60]), .B2(n4357), .C1(opb_r[61]), .C2(n4448), 
        .A(n4737), .ZN(n4738) );
  NAND2_X1 U4377 ( .A1(opb_r[61]), .A2(n4448), .ZN(n4749) );
  OAI211_X1 U4378 ( .C1(opa_r[62]), .C2(n4755), .A(n4738), .B(n4749), .ZN(
        n4739) );
  AOI21_X1 U4379 ( .B1(n4755), .B2(opa_r[62]), .A(n4757), .ZN(n4754) );
  AND3_X1 U4380 ( .A1(n4742), .A2(n4741), .A3(n4740), .ZN(n4743) );
  NAND4_X1 U4381 ( .A1(n4745), .A2(n4754), .A3(n4744), .A4(n4743), .ZN(n4753)
         );
  AND2_X1 U4382 ( .A1(opb_r[52]), .A2(n4449), .ZN(n4746) );
  OAI22_X1 U4383 ( .A1(n4746), .A2(n4450), .B1(opb_r[53]), .B2(n4746), .ZN(
        n4751) );
  AND3_X1 U4384 ( .A1(n4749), .A2(n4748), .A3(n4747), .ZN(n4750) );
  OAI211_X1 U4385 ( .C1(opa_r[62]), .C2(n4755), .A(n4751), .B(n4750), .ZN(
        n4752) );
  NOR2_X1 U4386 ( .A1(n4753), .A2(n4752), .ZN(\u1/N49 ) );
  INV_X4 U4387 ( .A(opb_r[62]), .ZN(n4755) );
  INV_X4 U4388 ( .A(n4730), .ZN(n4756) );
  INV_X4 U4389 ( .A(n4739), .ZN(n4757) );
  INV_X4 U4390 ( .A(n4754), .ZN(\u1/expa_lt_expb ) );
  NOR2_X1 U4391 ( .A1(\u1/exp_diff[6] ), .A2(\u1/exp_diff[10] ), .ZN(n4761) );
  OR3_X1 U4392 ( .A1(\u1/exp_diff[2] ), .A2(\u1/exp_diff[1] ), .A3(
        \u1/exp_diff[0] ), .ZN(n4758) );
  NAND4_X1 U4393 ( .A1(\u1/exp_diff[5] ), .A2(\u1/exp_diff[4] ), .A3(
        \u1/exp_diff[3] ), .A4(n4758), .ZN(n4760) );
  NOR3_X1 U4394 ( .A1(\u1/exp_diff[7] ), .A2(\u1/exp_diff[9] ), .A3(
        \u1/exp_diff[8] ), .ZN(n4759) );
  NAND3_X1 U4395 ( .A1(n4761), .A2(n4760), .A3(n4759), .ZN(\u1/exp_lt_27 ) );
  NOR2_X1 U4396 ( .A1(\u4/div_shft3[6] ), .A2(\u4/div_shft3[10] ), .ZN(n4764)
         );
  OAI211_X1 U4397 ( .C1(\u4/div_shft3[2] ), .C2(\u4/div_shft3[3] ), .A(
        \u4/div_shft3[4] ), .B(\u4/div_shft3[5] ), .ZN(n4763) );
  NOR3_X1 U4398 ( .A1(\u4/div_shft3[7] ), .A2(\u4/div_shft3[9] ), .A3(
        \u4/div_shft3[8] ), .ZN(n4762) );
  NAND3_X1 U4399 ( .A1(n4764), .A2(n4763), .A3(n4762), .ZN(\u4/N5843 ) );
  NAND4_X1 U4400 ( .A1(\u4/div_exp2[3] ), .A2(\u4/div_exp2[2] ), .A3(
        \u4/div_exp2[1] ), .A4(\u4/div_exp2[0] ), .ZN(n4766) );
  NAND4_X1 U4401 ( .A1(\u4/div_exp2[7] ), .A2(\u4/div_exp2[6] ), .A3(
        \u4/div_exp2[5] ), .A4(\u4/div_exp2[4] ), .ZN(n4765) );
  NOR2_X1 U4402 ( .A1(n4766), .A2(n4765), .ZN(n4767) );
  OR4_X1 U4403 ( .A1(\u4/div_exp2[10] ), .A2(n4767), .A3(\u4/div_exp2[9] ), 
        .A4(\u4/div_exp2[8] ), .ZN(\u4/N6172 ) );
  NAND3_X1 U4404 ( .A1(\u4/div_exp1[1] ), .A2(\u4/div_exp1[0] ), .A3(
        \u4/div_exp1[2] ), .ZN(n4771) );
  NAND2_X1 U4405 ( .A1(\u4/div_exp1[4] ), .A2(\u4/div_exp1[3] ), .ZN(n4770) );
  NAND3_X1 U4406 ( .A1(\u4/div_exp1[6] ), .A2(\u4/div_exp1[5] ), .A3(
        \u4/div_exp1[7] ), .ZN(n4769) );
  NAND2_X1 U4407 ( .A1(\u4/div_exp1[9] ), .A2(\u4/div_exp1[8] ), .ZN(n4768) );
  NOR4_X1 U4408 ( .A1(n4771), .A2(n4770), .A3(n4769), .A4(n4768), .ZN(n4772)
         );
  NOR2_X1 U4409 ( .A1(\u4/div_exp1[10] ), .A2(n4772), .ZN(\u4/N6194 ) );
  OAI211_X1 U4410 ( .C1(\u4/ldz_all[3] ), .C2(\u4/ldz_all[2] ), .A(
        \u4/ldz_all[4] ), .B(\u4/ldz_all[5] ), .ZN(n4773) );
  NOR2_X1 U4411 ( .A1(\u4/ldz_all[6] ), .A2(n4774), .ZN(\u4/N6286 ) );
  INV_X4 U4412 ( .A(n4773), .ZN(n4774) );
  OR3_X1 U4413 ( .A1(n4282), .A2(exp_r[3]), .A3(n4315), .ZN(n4775) );
  OR3_X1 U4414 ( .A1(exp_r[1]), .A2(n4600), .A3(n4775), .ZN(n4776) );
  AOI211_X1 U4415 ( .C1(n4290), .C2(n4776), .A(exp_r[6]), .B(n4352), .ZN(n4778) );
  NOR3_X1 U4416 ( .A1(n4281), .A2(n4289), .A3(n4353), .ZN(n4777) );
  NAND2_X1 U4417 ( .A1(n4778), .A2(n4777), .ZN(\u4/N6284 ) );
  NAND4_X1 U4418 ( .A1(exp_r[3]), .A2(n4315), .A3(exp_r[1]), .A4(n4600), .ZN(
        n4780) );
  NAND3_X1 U4419 ( .A1(n4290), .A2(n4282), .A3(exp_r[6]), .ZN(n4779) );
  OAI21_X1 U4420 ( .B1(n4780), .B2(n4779), .A(n4440), .ZN(n4781) );
  NOR4_X1 U4421 ( .A1(n4781), .A2(n4281), .A3(n4289), .A4(n4353), .ZN(
        \u4/N6283 ) );
  NOR2_X1 U4422 ( .A1(exp_r[6]), .A2(n4352), .ZN(n4783) );
  OAI211_X1 U4423 ( .C1(exp_r[3]), .C2(n4315), .A(n4282), .B(n4290), .ZN(n4782) );
  NAND2_X1 U4424 ( .A1(n4783), .A2(n4782), .ZN(n4784) );
  NOR4_X1 U4425 ( .A1(n4784), .A2(n4281), .A3(n4289), .A4(n4353), .ZN(
        \u4/N6280 ) );
  NOR2_X1 U4426 ( .A1(n4290), .A2(n4352), .ZN(n4788) );
  AND3_X1 U4427 ( .A1(exp_r[1]), .A2(n4600), .A3(n4315), .ZN(n4785) );
  OAI21_X1 U4428 ( .B1(n4785), .B2(n4655), .A(n4282), .ZN(n4787) );
  NOR4_X1 U4429 ( .A1(n4289), .A2(n4353), .A3(n4281), .A4(exp_r[6]), .ZN(n4786) );
  NAND3_X1 U4430 ( .A1(n4788), .A2(n4787), .A3(n4786), .ZN(\u4/N6278 ) );
  AND2_X1 U4431 ( .A1(\u4/fi_ldz_2a[4] ), .A2(\u4/fi_ldz_2a[3] ), .ZN(n4789)
         );
  OAI211_X1 U4432 ( .C1(\u4/fi_ldz[2] ), .C2(\u4/fi_ldz[3] ), .A(
        \u4/fi_ldz[5] ), .B(\u4/fi_ldz[4] ), .ZN(n4790) );
  NAND2_X1 U4433 ( .A1(n4663), .A2(n4790), .ZN(\u4/N6203 ) );
  OR4_X1 U4434 ( .A1(n4281), .A2(exp_r[6]), .A3(n4289), .A4(n4353), .ZN(n4797)
         );
  NOR2_X1 U4435 ( .A1(n4447), .A2(n4600), .ZN(n4791) );
  AOI21_X1 U4436 ( .B1(n4791), .B2(n4314), .A(div_opa_ldz_r2[1]), .ZN(n4792)
         );
  AOI221_X1 U4437 ( .B1(n4315), .B2(n4444), .C1(exp_r[1]), .C2(
        \u4/sub_409/carry [1]), .A(n4792), .ZN(n4793) );
  AOI221_X1 U4438 ( .B1(div_opa_ldz_r2[3]), .B2(n4316), .C1(div_opa_ldz_r2[2]), 
        .C2(n4438), .A(n4793), .ZN(n4794) );
  AOI221_X1 U4439 ( .B1(n4282), .B2(n4445), .C1(n4655), .C2(n4443), .A(n4794), 
        .ZN(n4795) );
  AOI21_X1 U4440 ( .B1(div_opa_ldz_r2[4]), .B2(n4299), .A(n4795), .ZN(n4796)
         );
  NOR4_X1 U4441 ( .A1(n4797), .A2(n4796), .A3(n4290), .A4(n4352), .ZN(
        \u4/N6171 ) );
  NAND3_X1 U4442 ( .A1(\u2/exp_tmp1[1] ), .A2(\u2/lt_135/A[0] ), .A3(
        \u2/exp_tmp1[2] ), .ZN(n4801) );
  NAND2_X1 U4443 ( .A1(\u2/exp_tmp1[4] ), .A2(\u2/exp_tmp1[3] ), .ZN(n4800) );
  NAND3_X1 U4444 ( .A1(\u2/lt_135/A[6] ), .A2(\u2/lt_135/A[5] ), .A3(
        \u2/lt_135/A[7] ), .ZN(n4799) );
  NAND2_X1 U4445 ( .A1(\u2/lt_135/A[9] ), .A2(\u2/lt_135/A[8] ), .ZN(n4798) );
  NOR4_X1 U4446 ( .A1(n4801), .A2(n4800), .A3(n4799), .A4(n4798), .ZN(n4802)
         );
  OAI21_X1 U4447 ( .B1(n4802), .B2(\u2/exp_tmp4[10] ), .A(\u2/gt_145/B[11] ), 
        .ZN(n4803) );
  INV_X4 U4448 ( .A(n4803), .ZN(\u2/N113 ) );
  NAND3_X1 U4449 ( .A1(\u2/exp_tmp1[1] ), .A2(\u2/lt_135/A[0] ), .A3(
        \u2/exp_tmp1[2] ), .ZN(n4807) );
  NAND2_X1 U4450 ( .A1(\u2/exp_tmp1[4] ), .A2(\u2/exp_tmp1[3] ), .ZN(n4806) );
  NAND3_X1 U4451 ( .A1(\u2/lt_135/A[6] ), .A2(\u2/lt_135/A[5] ), .A3(
        \u2/lt_135/A[7] ), .ZN(n4805) );
  NAND2_X1 U4452 ( .A1(\u2/lt_135/A[9] ), .A2(\u2/lt_135/A[8] ), .ZN(n4804) );
  NOR4_X1 U4453 ( .A1(n4807), .A2(n4806), .A3(n4805), .A4(n4804), .ZN(n4808)
         );
  NOR2_X1 U4454 ( .A1(\u2/exp_tmp4[10] ), .A2(n4808), .ZN(\u2/N111 ) );
  OAI211_X1 U4455 ( .C1(\u4/fi_ldz[3] ), .C2(\u4/fi_ldz[2] ), .A(
        \u4/fi_ldz[4] ), .B(\u4/fi_ldz[5] ), .ZN(n4809) );
  NOR2_X1 U4456 ( .A1(\u4/fi_ldz[6] ), .A2(n4810), .ZN(\u4/N6279 ) );
  INV_X4 U4457 ( .A(n4809), .ZN(n4810) );
  OAI21_X1 U4458 ( .B1(\u4/fi_ldz_2a[1] ), .B2(\u4/fi_ldz_2a[0] ), .A(
        \u4/fi_ldz_2a[2] ), .ZN(n4811) );
  AOI21_X1 U4459 ( .B1(n4811), .B2(n4813), .A(n4814), .ZN(n4812) );
  INV_X4 U4460 ( .A(\u4/fi_ldz_2a[3] ), .ZN(n4813) );
  INV_X4 U4461 ( .A(\u4/fi_ldz_2a[4] ), .ZN(n4814) );
  NOR2_X1 U4462 ( .A1(exp_r[6]), .A2(n4290), .ZN(n4816) );
  NAND4_X1 U4463 ( .A1(exp_r[1]), .A2(n4315), .A3(n4282), .A4(n4655), .ZN(
        n4815) );
  AOI21_X1 U4464 ( .B1(n4816), .B2(n4815), .A(n4348), .ZN(n4817) );
  OR4_X1 U4465 ( .A1(n4352), .A2(n4817), .A3(n4289), .A4(n4353), .ZN(
        \u4/N5837 ) );
  OAI211_X1 U4466 ( .C1(n4600), .C2(n4823), .A(exp_r[1]), .B(n4315), .ZN(n4821) );
  NAND2_X1 U4467 ( .A1(n4282), .A2(n4655), .ZN(n4820) );
  NAND3_X1 U4468 ( .A1(exp_r[6]), .A2(n4290), .A3(n4281), .ZN(n4819) );
  NAND2_X1 U4469 ( .A1(n4289), .A2(n4353), .ZN(n4818) );
  NOR4_X1 U4470 ( .A1(n4821), .A2(n4820), .A3(n4819), .A4(n4818), .ZN(n4822)
         );
  NOR2_X1 U4471 ( .A1(n4352), .A2(n4822), .ZN(\u4/N5836 ) );
  INV_X4 U4472 ( .A(\u4/N6410 ), .ZN(n4823) );
  NAND2_X2 U4473 ( .A1(\u4/exp_f2i_1 [116]), .A2(n2400), .ZN(n2429) );
  NAND2_X2 U4474 ( .A1(\u4/exp_f2i_1 [117]), .A2(n2400), .ZN(n2432) );
  NAND2_X2 U4475 ( .A1(\u4/exp_f2i_1 [115]), .A2(n2400), .ZN(n2425) );
  AOI22_X2 U4476 ( .A1(opa_r1[0]), .A2(n4552), .B1(N343), .B2(n4546), .ZN(
        n4249) );
  AOI22_X2 U4477 ( .A1(opa_r1[1]), .A2(n4553), .B1(N344), .B2(n4197), .ZN(
        n4248) );
  AOI22_X2 U4478 ( .A1(opa_r1[2]), .A2(n4553), .B1(N345), .B2(n4197), .ZN(
        n4247) );
  AOI22_X2 U4479 ( .A1(opa_r1[3]), .A2(n4553), .B1(N346), .B2(n4546), .ZN(
        n4246) );
  AOI22_X2 U4480 ( .A1(opa_r1[4]), .A2(n4553), .B1(N347), .B2(n4546), .ZN(
        n4245) );
  AOI22_X2 U4481 ( .A1(opa_r1[5]), .A2(n4552), .B1(N348), .B2(n4546), .ZN(
        n4244) );
  AOI22_X2 U4482 ( .A1(opa_r1[6]), .A2(n4553), .B1(N349), .B2(n4546), .ZN(
        n4243) );
  AOI22_X2 U4483 ( .A1(n4552), .A2(opa_r1[7]), .B1(N350), .B2(n4546), .ZN(
        n4242) );
  AOI22_X2 U4484 ( .A1(n4552), .A2(opa_r1[8]), .B1(N351), .B2(n4546), .ZN(
        n4241) );
  AOI22_X2 U4485 ( .A1(n4552), .A2(opa_r1[9]), .B1(N352), .B2(n4546), .ZN(
        n4240) );
  AOI22_X2 U4486 ( .A1(n4552), .A2(opa_r1[10]), .B1(N353), .B2(n4546), .ZN(
        n4239) );
  AOI22_X2 U4487 ( .A1(n4552), .A2(opa_r1[11]), .B1(N354), .B2(n4546), .ZN(
        n4238) );
  AOI22_X2 U4488 ( .A1(n4552), .A2(opa_r1[12]), .B1(N355), .B2(n4546), .ZN(
        n4237) );
  AOI22_X2 U4489 ( .A1(n4552), .A2(opa_r1[13]), .B1(N356), .B2(n4546), .ZN(
        n4236) );
  AOI22_X2 U4490 ( .A1(n4551), .A2(opa_r1[14]), .B1(N357), .B2(n4546), .ZN(
        n4235) );
  AOI22_X2 U4491 ( .A1(n4551), .A2(opa_r1[15]), .B1(N358), .B2(n4547), .ZN(
        n4234) );
  AOI22_X2 U4492 ( .A1(n4551), .A2(opa_r1[16]), .B1(N359), .B2(n4547), .ZN(
        n4233) );
  AOI22_X2 U4493 ( .A1(n4551), .A2(opa_r1[17]), .B1(N360), .B2(n4547), .ZN(
        n4232) );
  AOI22_X2 U4494 ( .A1(n4551), .A2(opa_r1[18]), .B1(N361), .B2(n4547), .ZN(
        n4231) );
  AOI22_X2 U4495 ( .A1(n4551), .A2(opa_r1[19]), .B1(N362), .B2(n4547), .ZN(
        n4230) );
  AOI22_X2 U4496 ( .A1(n4551), .A2(opa_r1[20]), .B1(N363), .B2(n4547), .ZN(
        n4229) );
  AOI22_X2 U4497 ( .A1(n4551), .A2(opa_r1[21]), .B1(N364), .B2(n4547), .ZN(
        n4228) );
  AOI22_X2 U4498 ( .A1(n4551), .A2(opa_r1[22]), .B1(N365), .B2(n4547), .ZN(
        n4227) );
  AOI22_X2 U4499 ( .A1(n4551), .A2(opa_r1[23]), .B1(N366), .B2(n4547), .ZN(
        n4226) );
  AOI22_X2 U4500 ( .A1(n4550), .A2(opa_r1[24]), .B1(N367), .B2(n4547), .ZN(
        n4225) );
  AOI22_X2 U4501 ( .A1(n4550), .A2(opa_r1[25]), .B1(N368), .B2(n4547), .ZN(
        n4224) );
  AOI22_X2 U4502 ( .A1(n4550), .A2(opa_r1[26]), .B1(N369), .B2(n4548), .ZN(
        n4223) );
  AOI22_X2 U4503 ( .A1(n4550), .A2(opa_r1[27]), .B1(N370), .B2(n4548), .ZN(
        n4222) );
  AOI22_X2 U4504 ( .A1(n4550), .A2(opa_r1[28]), .B1(N371), .B2(n4548), .ZN(
        n4221) );
  AOI22_X2 U4505 ( .A1(n4550), .A2(opa_r1[29]), .B1(N372), .B2(n4548), .ZN(
        n4220) );
  AOI22_X2 U4506 ( .A1(n4550), .A2(opa_r1[30]), .B1(N373), .B2(n4548), .ZN(
        n4219) );
  AOI22_X2 U4507 ( .A1(n4550), .A2(opa_r1[31]), .B1(N374), .B2(n4548), .ZN(
        n4218) );
  AOI22_X2 U4508 ( .A1(n4550), .A2(opa_r1[32]), .B1(N375), .B2(n4548), .ZN(
        n4217) );
  AOI22_X2 U4509 ( .A1(n4550), .A2(opa_r1[33]), .B1(N376), .B2(n4548), .ZN(
        n4216) );
  AOI22_X2 U4510 ( .A1(n4550), .A2(opa_r1[34]), .B1(N377), .B2(n4548), .ZN(
        n4215) );
  AOI22_X2 U4511 ( .A1(n4552), .A2(opa_r1[35]), .B1(N378), .B2(n4548), .ZN(
        n4214) );
  AOI22_X2 U4512 ( .A1(n4552), .A2(opa_r1[36]), .B1(N379), .B2(n4548), .ZN(
        n4213) );
  AOI22_X2 U4513 ( .A1(n4552), .A2(opa_r1[37]), .B1(N380), .B2(n4548), .ZN(
        n4212) );
  AOI22_X2 U4514 ( .A1(n4552), .A2(opa_r1[38]), .B1(N381), .B2(n4547), .ZN(
        n4211) );
  AOI22_X2 U4515 ( .A1(n4552), .A2(opa_r1[39]), .B1(N382), .B2(n4546), .ZN(
        n4210) );
  AOI22_X2 U4516 ( .A1(n4552), .A2(opa_r1[40]), .B1(N383), .B2(n4548), .ZN(
        n4209) );
  AOI22_X2 U4517 ( .A1(n4552), .A2(opa_r1[41]), .B1(N384), .B2(n4547), .ZN(
        n4208) );
  AOI22_X2 U4518 ( .A1(n4552), .A2(opa_r1[42]), .B1(N385), .B2(n4546), .ZN(
        n4207) );
  AOI22_X2 U4519 ( .A1(n4552), .A2(opa_r1[43]), .B1(N386), .B2(n4548), .ZN(
        n4206) );
  AOI22_X2 U4520 ( .A1(n4552), .A2(opa_r1[44]), .B1(N387), .B2(n4547), .ZN(
        n4205) );
  AOI22_X2 U4521 ( .A1(n4551), .A2(opa_r1[45]), .B1(N388), .B2(n4546), .ZN(
        n4204) );
  INV_X4 U4522 ( .A(n3504), .ZN(n5864) );
  INV_X4 U4523 ( .A(n2430), .ZN(n5865) );
  INV_X4 U4524 ( .A(n2427), .ZN(n5866) );
  INV_X4 U4525 ( .A(n2423), .ZN(n5867) );
  INV_X4 U4526 ( .A(n3512), .ZN(n5868) );
  INV_X4 U4527 ( .A(n3506), .ZN(n5869) );
  INV_X4 U4528 ( .A(n3509), .ZN(n5870) );
  INV_X4 U4529 ( .A(n2413), .ZN(n5871) );
  INV_X4 U4530 ( .A(n2410), .ZN(n5872) );
  INV_X4 U4531 ( .A(n2406), .ZN(n5873) );
  INV_X4 U4532 ( .A(N307), .ZN(n5874) );
  INV_X4 U4533 ( .A(N306), .ZN(n5875) );
  INV_X4 U4534 ( .A(n3192), .ZN(\u6/N104 ) );
  INV_X4 U4535 ( .A(n3193), .ZN(\u6/N103 ) );
  INV_X4 U4536 ( .A(n3194), .ZN(\u6/N102 ) );
  INV_X4 U4537 ( .A(N302), .ZN(n5876) );
  INV_X4 U4538 ( .A(N301), .ZN(n5877) );
  INV_X4 U4539 ( .A(N300), .ZN(n5878) );
  INV_X4 U4540 ( .A(n3181), .ZN(\u6/N98 ) );
  INV_X4 U4541 ( .A(N298), .ZN(n5879) );
  INV_X4 U4542 ( .A(N297), .ZN(n5880) );
  INV_X4 U4543 ( .A(n3182), .ZN(\u6/N95 ) );
  INV_X4 U4544 ( .A(N295), .ZN(n5881) );
  INV_X4 U4545 ( .A(N294), .ZN(n5882) );
  INV_X4 U4546 ( .A(N293), .ZN(n5883) );
  INV_X4 U4547 ( .A(N292), .ZN(n5884) );
  INV_X4 U4548 ( .A(N291), .ZN(n5885) );
  INV_X4 U4549 ( .A(n3183), .ZN(\u6/N89 ) );
  INV_X4 U4550 ( .A(n3184), .ZN(\u6/N88 ) );
  INV_X4 U4551 ( .A(N288), .ZN(n5886) );
  INV_X4 U4552 ( .A(N287), .ZN(n5887) );
  INV_X4 U4553 ( .A(N286), .ZN(n5888) );
  INV_X4 U4554 ( .A(N285), .ZN(n5889) );
  INV_X4 U4555 ( .A(N284), .ZN(n5890) );
  INV_X4 U4556 ( .A(N283), .ZN(n5891) );
  INV_X4 U4557 ( .A(n3185), .ZN(\u6/N81 ) );
  INV_X4 U4558 ( .A(N281), .ZN(n5892) );
  INV_X4 U4559 ( .A(n3186), .ZN(\u6/N79 ) );
  INV_X4 U4560 ( .A(n3187), .ZN(\u6/N78 ) );
  INV_X4 U4561 ( .A(N278), .ZN(n5893) );
  INV_X4 U4562 ( .A(N277), .ZN(n5894) );
  INV_X4 U4563 ( .A(N276), .ZN(n5895) );
  INV_X4 U4564 ( .A(n3188), .ZN(\u6/N74 ) );
  INV_X4 U4565 ( .A(N274), .ZN(n5896) );
  INV_X4 U4566 ( .A(N273), .ZN(n5897) );
  INV_X4 U4567 ( .A(N272), .ZN(n5898) );
  INV_X4 U4568 ( .A(N271), .ZN(n5899) );
  INV_X4 U4569 ( .A(N270), .ZN(n5900) );
  INV_X4 U4570 ( .A(n3189), .ZN(\u6/N68 ) );
  INV_X4 U4571 ( .A(N268), .ZN(n5901) );
  INV_X4 U4572 ( .A(N267), .ZN(n5902) );
  INV_X4 U4573 ( .A(N266), .ZN(n5903) );
  INV_X4 U4574 ( .A(N265), .ZN(n5904) );
  INV_X4 U4575 ( .A(N264), .ZN(n5905) );
  INV_X4 U4576 ( .A(N263), .ZN(n5906) );
  INV_X4 U4577 ( .A(N262), .ZN(n5907) );
  INV_X4 U4578 ( .A(N261), .ZN(n5908) );
  INV_X4 U4579 ( .A(n3190), .ZN(\u6/N59 ) );
  INV_X4 U4580 ( .A(N259), .ZN(n5909) );
  INV_X4 U4581 ( .A(n3191), .ZN(\u6/N57 ) );
  INV_X4 U4582 ( .A(N257), .ZN(n5910) );
  INV_X4 U4583 ( .A(N256), .ZN(n5911) );
  INV_X4 U4584 ( .A(n3783), .ZN(n5912) );
  INV_X4 U4585 ( .A(n4204), .ZN(n5913) );
  INV_X4 U4586 ( .A(n4205), .ZN(n5914) );
  INV_X4 U4587 ( .A(n4206), .ZN(n5915) );
  INV_X4 U4588 ( .A(n4207), .ZN(n5916) );
  INV_X4 U4589 ( .A(n4208), .ZN(n5917) );
  INV_X4 U4590 ( .A(n4209), .ZN(n5918) );
  INV_X4 U4591 ( .A(n4210), .ZN(n5919) );
  INV_X4 U4592 ( .A(n4211), .ZN(n5920) );
  INV_X4 U4593 ( .A(n4212), .ZN(n5921) );
  INV_X4 U4594 ( .A(n4213), .ZN(n5922) );
  INV_X4 U4595 ( .A(n4214), .ZN(n5923) );
  INV_X4 U4596 ( .A(n4215), .ZN(n5924) );
  INV_X4 U4597 ( .A(n4216), .ZN(n5925) );
  INV_X4 U4598 ( .A(n4217), .ZN(n5926) );
  INV_X4 U4599 ( .A(n4218), .ZN(n5927) );
  INV_X4 U4600 ( .A(n4219), .ZN(n5928) );
  INV_X4 U4601 ( .A(n4220), .ZN(n5929) );
  INV_X4 U4602 ( .A(n4221), .ZN(n5930) );
  INV_X4 U4603 ( .A(n4222), .ZN(n5931) );
  INV_X4 U4604 ( .A(n4223), .ZN(n5932) );
  INV_X4 U4605 ( .A(n4224), .ZN(n5933) );
  INV_X4 U4606 ( .A(n4225), .ZN(n5934) );
  INV_X4 U4607 ( .A(n4226), .ZN(n5935) );
  INV_X4 U4608 ( .A(n4227), .ZN(n5936) );
  INV_X4 U4609 ( .A(n4228), .ZN(n5937) );
  INV_X4 U4610 ( .A(n4229), .ZN(n5938) );
  INV_X4 U4611 ( .A(n4230), .ZN(n5939) );
  INV_X4 U4612 ( .A(n4231), .ZN(n5940) );
  INV_X4 U4613 ( .A(n4232), .ZN(n5941) );
  INV_X4 U4614 ( .A(n4233), .ZN(n5942) );
  INV_X4 U4615 ( .A(n4234), .ZN(n5943) );
  INV_X4 U4616 ( .A(n4235), .ZN(n5944) );
  INV_X4 U4617 ( .A(n4236), .ZN(n5945) );
  INV_X4 U4618 ( .A(n4237), .ZN(n5946) );
  INV_X4 U4619 ( .A(n4238), .ZN(n5947) );
  INV_X4 U4620 ( .A(n4239), .ZN(n5948) );
  INV_X4 U4621 ( .A(n4240), .ZN(n5949) );
  INV_X4 U4622 ( .A(n4241), .ZN(n5950) );
  INV_X4 U4623 ( .A(n4242), .ZN(n5951) );
  INV_X4 U4624 ( .A(n4243), .ZN(n5952) );
  INV_X4 U4625 ( .A(n4244), .ZN(n5953) );
  INV_X4 U4626 ( .A(n4245), .ZN(n5954) );
  INV_X4 U4627 ( .A(n4246), .ZN(n5955) );
  INV_X4 U4628 ( .A(n4247), .ZN(n5956) );
  INV_X4 U4629 ( .A(n4248), .ZN(n5957) );
  INV_X4 U4630 ( .A(N557), .ZN(n5958) );
  INV_X4 U4631 ( .A(N556), .ZN(n5959) );
  INV_X4 U4632 ( .A(N555), .ZN(n5960) );
  INV_X4 U4633 ( .A(N554), .ZN(n5961) );
  INV_X4 U4634 ( .A(N553), .ZN(n5962) );
  INV_X4 U4635 ( .A(N552), .ZN(n5963) );
  INV_X4 U4636 ( .A(N551), .ZN(n5964) );
  INV_X4 U4637 ( .A(N550), .ZN(n5965) );
  INV_X4 U4638 ( .A(N549), .ZN(n5966) );
  INV_X4 U4639 ( .A(N548), .ZN(n5967) );
  INV_X4 U4640 ( .A(N547), .ZN(n5968) );
  INV_X4 U4641 ( .A(N546), .ZN(n5969) );
  INV_X4 U4642 ( .A(N545), .ZN(n5970) );
  INV_X4 U4643 ( .A(N544), .ZN(n5971) );
  INV_X4 U4644 ( .A(N543), .ZN(n5972) );
  INV_X4 U4645 ( .A(N542), .ZN(n5973) );
  INV_X4 U4646 ( .A(N541), .ZN(n5974) );
  INV_X4 U4647 ( .A(N540), .ZN(n5975) );
  INV_X4 U4648 ( .A(N539), .ZN(n5976) );
  INV_X4 U4649 ( .A(N538), .ZN(n5977) );
  INV_X4 U4650 ( .A(N537), .ZN(n5978) );
  INV_X4 U4651 ( .A(N536), .ZN(n5979) );
  INV_X4 U4652 ( .A(N535), .ZN(n5980) );
  INV_X4 U4653 ( .A(N534), .ZN(n5981) );
  INV_X4 U4654 ( .A(N533), .ZN(n5982) );
  INV_X4 U4655 ( .A(N532), .ZN(n5983) );
  INV_X4 U4656 ( .A(N531), .ZN(n5984) );
  INV_X4 U4657 ( .A(N530), .ZN(n5985) );
  INV_X4 U4658 ( .A(N529), .ZN(n5986) );
  INV_X4 U4659 ( .A(N528), .ZN(n5987) );
  INV_X4 U4660 ( .A(N527), .ZN(n5988) );
  INV_X4 U4661 ( .A(N526), .ZN(n5989) );
  INV_X4 U4662 ( .A(N525), .ZN(n5990) );
  INV_X4 U4663 ( .A(N524), .ZN(n5991) );
  INV_X4 U4664 ( .A(N523), .ZN(n5992) );
  INV_X4 U4665 ( .A(N522), .ZN(n5993) );
  INV_X4 U4666 ( .A(N521), .ZN(n5994) );
  INV_X4 U4667 ( .A(N520), .ZN(n5995) );
  INV_X4 U4668 ( .A(N519), .ZN(n5996) );
  INV_X4 U4669 ( .A(N518), .ZN(n5997) );
  INV_X4 U4670 ( .A(N517), .ZN(n5998) );
  INV_X4 U4671 ( .A(N516), .ZN(n5999) );
  INV_X4 U4672 ( .A(N515), .ZN(n6000) );
  INV_X4 U4673 ( .A(N514), .ZN(n6001) );
  INV_X4 U4674 ( .A(N513), .ZN(n6002) );
  INV_X4 U4675 ( .A(N512), .ZN(n6003) );
  INV_X4 U4676 ( .A(N511), .ZN(n6004) );
  INV_X4 U4677 ( .A(N510), .ZN(n6005) );
  INV_X4 U4678 ( .A(N509), .ZN(n6006) );
  INV_X4 U4679 ( .A(N508), .ZN(n6007) );
  INV_X4 U4680 ( .A(N507), .ZN(n6008) );
  INV_X4 U4681 ( .A(N506), .ZN(n6009) );
  INV_X4 U4682 ( .A(N505), .ZN(n6010) );
  INV_X4 U4683 ( .A(N504), .ZN(n6011) );
  INV_X4 U4684 ( .A(N503), .ZN(n6012) );
  INV_X4 U4685 ( .A(N502), .ZN(n6013) );
  INV_X4 U4686 ( .A(N501), .ZN(n6014) );
  INV_X4 U4687 ( .A(\u2/exp_ovf_d[1] ), .ZN(n6015) );
  INV_X4 U4688 ( .A(n2784), .ZN(\u2/gt_145/B[11] ) );
  INV_X4 U4689 ( .A(n2804), .ZN(n6016) );
  INV_X4 U4690 ( .A(\u2/N16 ), .ZN(n6017) );
  INV_X4 U4691 ( .A(n2785), .ZN(n6018) );
  INV_X4 U4692 ( .A(n2795), .ZN(\u2/lt_135/A[9] ) );
  INV_X4 U4693 ( .A(n2786), .ZN(n6019) );
  INV_X4 U4694 ( .A(n2796), .ZN(\u2/lt_135/A[8] ) );
  INV_X4 U4695 ( .A(n2787), .ZN(n6020) );
  INV_X4 U4696 ( .A(n2797), .ZN(\u2/lt_135/A[7] ) );
  INV_X4 U4697 ( .A(n2788), .ZN(n6021) );
  INV_X4 U4698 ( .A(n2798), .ZN(\u2/lt_135/A[6] ) );
  INV_X4 U4699 ( .A(n2789), .ZN(n6022) );
  INV_X4 U4700 ( .A(n2799), .ZN(\u2/lt_135/A[5] ) );
  INV_X4 U4701 ( .A(n2790), .ZN(n6023) );
  INV_X4 U4702 ( .A(\u2/N10 ), .ZN(n6024) );
  INV_X4 U4703 ( .A(n2791), .ZN(n6025) );
  INV_X4 U4704 ( .A(\u2/N9 ), .ZN(n6026) );
  INV_X4 U4705 ( .A(n2792), .ZN(n6027) );
  INV_X4 U4706 ( .A(\u2/N8 ), .ZN(n6028) );
  INV_X4 U4707 ( .A(n2793), .ZN(n6029) );
  INV_X4 U4708 ( .A(\u2/N7 ), .ZN(n6030) );
  INV_X4 U4709 ( .A(n2794), .ZN(n6031) );
  INV_X4 U4710 ( .A(\u2/N28 ), .ZN(n6032) );
  INV_X4 U4711 ( .A(\u2/N22 ), .ZN(n6033) );
  INV_X4 U4712 ( .A(\u2/N21 ), .ZN(n6034) );
  INV_X4 U4713 ( .A(\u2/N20 ), .ZN(n6035) );
  INV_X4 U4714 ( .A(\u2/N19 ), .ZN(n6036) );
  INV_X4 U4715 ( .A(n3292), .ZN(n6037) );
  INV_X4 U4716 ( .A(n3119), .ZN(n6038) );
  INV_X4 U4717 ( .A(n3120), .ZN(n6039) );
  INV_X4 U4718 ( .A(n3121), .ZN(n6040) );
  INV_X4 U4719 ( .A(n3122), .ZN(n6041) );
  INV_X4 U4720 ( .A(n3123), .ZN(n6042) );
  INV_X4 U4721 ( .A(n3124), .ZN(n6043) );
  INV_X4 U4722 ( .A(n3126), .ZN(n6044) );
  INV_X4 U4723 ( .A(n3127), .ZN(n6045) );
  INV_X4 U4724 ( .A(n3128), .ZN(n6046) );
  INV_X4 U4725 ( .A(n3129), .ZN(n6047) );
  INV_X4 U4726 ( .A(n3130), .ZN(n6048) );
  INV_X4 U4727 ( .A(n3131), .ZN(n6049) );
  INV_X4 U4728 ( .A(n3132), .ZN(n6050) );
  INV_X4 U4729 ( .A(n3133), .ZN(n6051) );
  INV_X4 U4730 ( .A(n3134), .ZN(n6052) );
  INV_X4 U4731 ( .A(n3135), .ZN(n6053) );
  INV_X4 U4732 ( .A(n3137), .ZN(n6054) );
  INV_X4 U4733 ( .A(n3138), .ZN(n6055) );
  INV_X4 U4734 ( .A(n3139), .ZN(n6056) );
  INV_X4 U4735 ( .A(n3140), .ZN(n6057) );
  INV_X4 U4736 ( .A(n3141), .ZN(n6058) );
  INV_X4 U4737 ( .A(n3142), .ZN(n6059) );
  INV_X4 U4738 ( .A(n3143), .ZN(n6060) );
  INV_X4 U4739 ( .A(n3144), .ZN(n6061) );
  INV_X4 U4740 ( .A(n3145), .ZN(n6062) );
  INV_X4 U4741 ( .A(n3146), .ZN(n6063) );
  INV_X4 U4742 ( .A(n3148), .ZN(n6064) );
  INV_X4 U4743 ( .A(n3149), .ZN(n6065) );
  INV_X4 U4744 ( .A(n3150), .ZN(n6066) );
  INV_X4 U4745 ( .A(n3151), .ZN(n6067) );
  INV_X4 U4746 ( .A(n3152), .ZN(n6068) );
  INV_X4 U4747 ( .A(n3153), .ZN(n6069) );
  INV_X4 U4748 ( .A(n3154), .ZN(n6070) );
  INV_X4 U4749 ( .A(n3155), .ZN(n6071) );
  INV_X4 U4750 ( .A(n3156), .ZN(n6072) );
  INV_X4 U4751 ( .A(n3157), .ZN(n6073) );
  INV_X4 U4752 ( .A(n3159), .ZN(n6074) );
  INV_X4 U4753 ( .A(n3160), .ZN(n6075) );
  INV_X4 U4754 ( .A(n3161), .ZN(n6076) );
  INV_X4 U4755 ( .A(n3162), .ZN(n6077) );
  INV_X4 U4756 ( .A(n3163), .ZN(n6078) );
  INV_X4 U4757 ( .A(n3164), .ZN(n6079) );
  INV_X4 U4758 ( .A(n3165), .ZN(n6080) );
  INV_X4 U4759 ( .A(n3166), .ZN(n6081) );
  INV_X4 U4760 ( .A(n3167), .ZN(n6082) );
  INV_X4 U4761 ( .A(n3168), .ZN(n6083) );
  INV_X4 U4762 ( .A(n3114), .ZN(n6084) );
  INV_X4 U4763 ( .A(n3115), .ZN(n6085) );
  INV_X4 U4764 ( .A(n3116), .ZN(n6086) );
  INV_X4 U4765 ( .A(n3117), .ZN(n6087) );
  INV_X4 U4766 ( .A(n3118), .ZN(n6088) );
  INV_X4 U4767 ( .A(n3125), .ZN(n6089) );
  INV_X4 U4768 ( .A(n3136), .ZN(n6090) );
  INV_X4 U4769 ( .A(n3147), .ZN(n6091) );
  INV_X4 U4770 ( .A(n3158), .ZN(n6092) );
  INV_X4 U4771 ( .A(n3169), .ZN(n6093) );
  INV_X4 U4772 ( .A(n3545), .ZN(n6094) );
  INV_X4 U4773 ( .A(n2438), .ZN(n6095) );
  INV_X4 U4774 ( .A(\u4/exp_next_mi[11] ), .ZN(n6096) );
  INV_X4 U4775 ( .A(n2431), .ZN(\u4/sub_468/A[10] ) );
  INV_X4 U4776 ( .A(n2428), .ZN(\u4/sub_468/A[9] ) );
  INV_X4 U4777 ( .A(n2420), .ZN(\u4/sub_468/A[7] ) );
  INV_X4 U4778 ( .A(n2416), .ZN(\u4/sub_468/A[5] ) );
  INV_X4 U4779 ( .A(n2414), .ZN(\u4/sub_468/A[4] ) );
  INV_X4 U4780 ( .A(n2411), .ZN(\u4/sub_468/A[3] ) );
  INV_X4 U4781 ( .A(n2407), .ZN(\u4/sub_468/A[2] ) );
  INV_X4 U4782 ( .A(\u4/exp_next_mi[1] ), .ZN(n6097) );
  INV_X4 U4783 ( .A(\u4/exp_next_mi[0] ), .ZN(n6098) );
  INV_X4 U4784 ( .A(\u1/N232 ), .ZN(n6099) );
  INV_X4 U4785 ( .A(n2836), .ZN(n6100) );
  INV_X4 U4786 ( .A(n2838), .ZN(n6101) );
  INV_X4 U4787 ( .A(n2840), .ZN(n6102) );
  INV_X4 U4788 ( .A(n2842), .ZN(n6103) );
  INV_X4 U4789 ( .A(n2844), .ZN(n6104) );
  INV_X4 U4790 ( .A(n2846), .ZN(n6105) );
  INV_X4 U4791 ( .A(n2848), .ZN(n6106) );
  INV_X4 U4792 ( .A(n2850), .ZN(n6107) );
  INV_X4 U4793 ( .A(n2852), .ZN(n6108) );
  INV_X4 U4794 ( .A(n2854), .ZN(n6109) );
  INV_X4 U4795 ( .A(n2856), .ZN(n6110) );
  INV_X4 U4796 ( .A(n2858), .ZN(n6111) );
  INV_X4 U4797 ( .A(n2860), .ZN(n6112) );
  INV_X4 U4798 ( .A(n2862), .ZN(n6113) );
  INV_X4 U4799 ( .A(n2864), .ZN(n6114) );
  INV_X4 U4800 ( .A(n2866), .ZN(n6115) );
  INV_X4 U4801 ( .A(n2868), .ZN(n6116) );
  INV_X4 U4802 ( .A(n2870), .ZN(n6117) );
  INV_X4 U4803 ( .A(n2872), .ZN(n6118) );
  INV_X4 U4804 ( .A(n2874), .ZN(n6119) );
  INV_X4 U4805 ( .A(n2876), .ZN(n6120) );
  INV_X4 U4806 ( .A(n2878), .ZN(n6121) );
  INV_X4 U4807 ( .A(n2880), .ZN(n6122) );
  INV_X4 U4808 ( .A(n2882), .ZN(n6123) );
  INV_X4 U4809 ( .A(n2884), .ZN(n6124) );
  INV_X4 U4810 ( .A(n2886), .ZN(n6125) );
  INV_X4 U4811 ( .A(n2888), .ZN(n6126) );
  INV_X4 U4812 ( .A(n2890), .ZN(n6127) );
  INV_X4 U4813 ( .A(n2892), .ZN(n6128) );
  INV_X4 U4814 ( .A(n2894), .ZN(n6129) );
  INV_X4 U4815 ( .A(n2896), .ZN(n6130) );
  INV_X4 U4816 ( .A(n2898), .ZN(n6131) );
  INV_X4 U4817 ( .A(n2900), .ZN(n6132) );
  INV_X4 U4818 ( .A(n2904), .ZN(n6133) );
  INV_X4 U4819 ( .A(n2906), .ZN(n6134) );
  INV_X4 U4820 ( .A(n2908), .ZN(n6135) );
  INV_X4 U4821 ( .A(n2910), .ZN(n6136) );
  INV_X4 U4822 ( .A(n2912), .ZN(n6137) );
  INV_X4 U4823 ( .A(n2914), .ZN(n6138) );
  INV_X4 U4824 ( .A(n2916), .ZN(n6139) );
  INV_X4 U4825 ( .A(n2918), .ZN(n6140) );
  INV_X4 U4826 ( .A(n2920), .ZN(n6141) );
  INV_X4 U4827 ( .A(n2922), .ZN(n6142) );
  INV_X4 U4828 ( .A(n2926), .ZN(n6143) );
  INV_X4 U4829 ( .A(n2928), .ZN(n6144) );
  INV_X4 U4830 ( .A(n2930), .ZN(n6145) );
  INV_X4 U4831 ( .A(n2932), .ZN(n6146) );
  INV_X4 U4832 ( .A(n2934), .ZN(n6147) );
  INV_X4 U4833 ( .A(n2936), .ZN(n6148) );
  INV_X4 U4834 ( .A(n2938), .ZN(n6149) );
  INV_X4 U4835 ( .A(n2940), .ZN(n6150) );
  INV_X4 U4836 ( .A(n2942), .ZN(n6151) );
  INV_X4 U4837 ( .A(n2944), .ZN(n6152) );
  INV_X4 U4838 ( .A(n2837), .ZN(n6153) );
  INV_X4 U4839 ( .A(n2839), .ZN(n6154) );
  INV_X4 U4840 ( .A(n2841), .ZN(n6155) );
  INV_X4 U4841 ( .A(n2843), .ZN(n6156) );
  INV_X4 U4842 ( .A(n2845), .ZN(n6157) );
  INV_X4 U4843 ( .A(n2847), .ZN(n6158) );
  INV_X4 U4844 ( .A(n2849), .ZN(n6159) );
  INV_X4 U4845 ( .A(n2851), .ZN(n6160) );
  INV_X4 U4846 ( .A(n2853), .ZN(n6161) );
  INV_X4 U4847 ( .A(n2855), .ZN(n6162) );
  INV_X4 U4848 ( .A(n2857), .ZN(n6163) );
  INV_X4 U4849 ( .A(n2859), .ZN(n6164) );
  INV_X4 U4850 ( .A(n2861), .ZN(n6165) );
  INV_X4 U4851 ( .A(n2863), .ZN(n6166) );
  INV_X4 U4852 ( .A(n2865), .ZN(n6167) );
  INV_X4 U4853 ( .A(n2867), .ZN(n6168) );
  INV_X4 U4854 ( .A(n2869), .ZN(n6169) );
  INV_X4 U4855 ( .A(n2871), .ZN(n6170) );
  INV_X4 U4856 ( .A(n2873), .ZN(n6171) );
  INV_X4 U4857 ( .A(n2875), .ZN(n6172) );
  INV_X4 U4858 ( .A(n2877), .ZN(n6173) );
  INV_X4 U4859 ( .A(n2879), .ZN(n6174) );
  INV_X4 U4860 ( .A(n2881), .ZN(n6175) );
  INV_X4 U4861 ( .A(n2883), .ZN(n6176) );
  INV_X4 U4862 ( .A(n2885), .ZN(n6177) );
  INV_X4 U4863 ( .A(n2887), .ZN(n6178) );
  INV_X4 U4864 ( .A(n2889), .ZN(n6179) );
  INV_X4 U4865 ( .A(n2891), .ZN(n6180) );
  INV_X4 U4866 ( .A(n2893), .ZN(n6181) );
  INV_X4 U4867 ( .A(n2895), .ZN(n6182) );
  INV_X4 U4868 ( .A(n2897), .ZN(n6183) );
  INV_X4 U4869 ( .A(n2899), .ZN(n6184) );
  INV_X4 U4870 ( .A(n2901), .ZN(n6185) );
  INV_X4 U4871 ( .A(n2903), .ZN(n6186) );
  INV_X4 U4872 ( .A(n2905), .ZN(n6187) );
  INV_X4 U4873 ( .A(n2907), .ZN(n6188) );
  INV_X4 U4874 ( .A(n2909), .ZN(n6189) );
  INV_X4 U4875 ( .A(n2911), .ZN(n6190) );
  INV_X4 U4876 ( .A(n2913), .ZN(n6191) );
  INV_X4 U4877 ( .A(n2915), .ZN(n6192) );
  INV_X4 U4878 ( .A(n2917), .ZN(n6193) );
  INV_X4 U4879 ( .A(n2919), .ZN(n6194) );
  INV_X4 U4880 ( .A(n2921), .ZN(n6195) );
  INV_X4 U4881 ( .A(n2923), .ZN(n6196) );
  INV_X4 U4882 ( .A(n2925), .ZN(n6197) );
  INV_X4 U4883 ( .A(n2927), .ZN(n6198) );
  INV_X4 U4884 ( .A(n2929), .ZN(n6199) );
  INV_X4 U4885 ( .A(n2931), .ZN(n6200) );
  INV_X4 U4886 ( .A(n2933), .ZN(n6201) );
  INV_X4 U4887 ( .A(n2935), .ZN(n6202) );
  INV_X4 U4888 ( .A(n2937), .ZN(n6203) );
  INV_X4 U4889 ( .A(n2939), .ZN(n6204) );
  INV_X4 U4890 ( .A(n2941), .ZN(n6205) );
  INV_X4 U4891 ( .A(n2943), .ZN(n6206) );
  INV_X4 U4892 ( .A(n2945), .ZN(n6207) );
  INV_X4 U4893 ( .A(n2947), .ZN(n6208) );
  INV_X4 U4894 ( .A(n2946), .ZN(n6209) );
  INV_X4 U4895 ( .A(n2924), .ZN(n6210) );
  INV_X4 U4896 ( .A(n2902), .ZN(n6211) );
  INV_X4 U4897 ( .A(n2968), .ZN(n6212) );
  INV_X4 U4898 ( .A(n2980), .ZN(n6213) );
  INV_X4 U4899 ( .A(n2975), .ZN(n6214) );
  INV_X4 U4900 ( .A(n2974), .ZN(n6215) );
  INV_X4 U4901 ( .A(n2960), .ZN(n6216) );
  INV_X4 U4902 ( .A(n3003), .ZN(n6217) );
  INV_X4 U4903 ( .A(n2961), .ZN(n6218) );
  INV_X4 U4904 ( .A(n2966), .ZN(n6219) );
  INV_X4 U4905 ( .A(n2958), .ZN(n6220) );
  INV_X4 U4906 ( .A(n2953), .ZN(n6221) );
  INV_X4 U4907 ( .A(n2995), .ZN(n6222) );
  INV_X4 U4908 ( .A(\u1/exp_lt_27 ), .ZN(n6223) );
  INV_X4 U4909 ( .A(n3001), .ZN(n6224) );
  INV_X4 U4910 ( .A(n3012), .ZN(n6225) );
  INV_X4 U4911 ( .A(n3004), .ZN(n6226) );
  INV_X4 U4912 ( .A(n3048), .ZN(n6227) );
  INV_X4 U4913 ( .A(n3049), .ZN(n6228) );
  INV_X4 U4914 ( .A(n3035), .ZN(n6229) );
  INV_X4 U4915 ( .A(n3034), .ZN(n6230) );
  INV_X4 U4916 ( .A(n3033), .ZN(n6231) );
  INV_X4 U4917 ( .A(n3032), .ZN(n6232) );
  INV_X4 U4918 ( .A(n3053), .ZN(n6233) );
  INV_X4 U4919 ( .A(n3013), .ZN(n6234) );
  INV_X4 U4920 ( .A(n3054), .ZN(n6235) );
  INV_X4 U4921 ( .A(n3055), .ZN(n6236) );
  INV_X4 U4922 ( .A(n3014), .ZN(n6237) );
  INV_X4 U4923 ( .A(n3056), .ZN(n6238) );
  INV_X4 U4924 ( .A(n3015), .ZN(n6239) );
  INV_X4 U4925 ( .A(n3016), .ZN(n6240) );
  INV_X4 U4926 ( .A(n3017), .ZN(n6241) );
  INV_X4 U4927 ( .A(n3018), .ZN(n6242) );
  INV_X4 U4928 ( .A(n3057), .ZN(n6243) );
  INV_X4 U4929 ( .A(n3019), .ZN(n6244) );
  INV_X4 U4930 ( .A(n3020), .ZN(n6245) );
  INV_X4 U4931 ( .A(n3021), .ZN(n6246) );
  INV_X4 U4932 ( .A(n3058), .ZN(n6247) );
  INV_X4 U4933 ( .A(n3022), .ZN(n6248) );
  INV_X4 U4934 ( .A(n3023), .ZN(n6249) );
  INV_X4 U4935 ( .A(n3038), .ZN(n6250) );
  INV_X4 U4936 ( .A(n3024), .ZN(n6251) );
  INV_X4 U4937 ( .A(n3025), .ZN(n6252) );
  INV_X4 U4938 ( .A(n3026), .ZN(n6253) );
  INV_X4 U4939 ( .A(n3037), .ZN(n6254) );
  INV_X4 U4940 ( .A(n3039), .ZN(n6255) );
  INV_X4 U4941 ( .A(n3042), .ZN(n6256) );
  INV_X4 U4942 ( .A(n3041), .ZN(n6257) );
  INV_X4 U4943 ( .A(n3043), .ZN(n6258) );
  INV_X4 U4944 ( .A(n3046), .ZN(n6259) );
  INV_X4 U4945 ( .A(n3045), .ZN(n6260) );
  INV_X4 U4946 ( .A(n3047), .ZN(n6261) );
  INV_X4 U4947 ( .A(\u1/exp_large[10] ), .ZN(n6262) );
  INV_X4 U4948 ( .A(n3050), .ZN(n6263) );
  INV_X4 U4949 ( .A(n3051), .ZN(n6264) );
  INV_X4 U4950 ( .A(\u1/exp_large[7] ), .ZN(n6265) );
  INV_X4 U4951 ( .A(\u1/exp_large[6] ), .ZN(n6266) );
  INV_X4 U4952 ( .A(\u1/exp_large[5] ), .ZN(n6267) );
  INV_X4 U4953 ( .A(\u1/exp_large[4] ), .ZN(n6268) );
  INV_X4 U4954 ( .A(\u1/exp_large[3] ), .ZN(n6269) );
  INV_X4 U4955 ( .A(\u1/exp_large[2] ), .ZN(n6270) );
  INV_X4 U4956 ( .A(\u1/exp_large[1] ), .ZN(n6271) );
  INV_X4 U4957 ( .A(\u1/exp_large[0] ), .ZN(n6272) );
  INV_X4 U4958 ( .A(n4266), .ZN(n6273) );
  INV_X4 U4959 ( .A(n2783), .ZN(n6274) );
  INV_X4 U4960 ( .A(\u1/N46 ), .ZN(n6275) );
  INV_X4 U4961 ( .A(n3075), .ZN(n6276) );
  INV_X4 U4962 ( .A(n3242), .ZN(n6277) );
  INV_X4 U4963 ( .A(n3227), .ZN(n6278) );
  INV_X4 U4964 ( .A(n3260), .ZN(n6279) );
  INV_X4 U4965 ( .A(n3208), .ZN(n6280) );
  INV_X4 U4966 ( .A(n3272), .ZN(n6281) );
  INV_X4 U4967 ( .A(n3209), .ZN(n6282) );
  INV_X4 U4968 ( .A(n3229), .ZN(n6283) );
  INV_X4 U4969 ( .A(n3220), .ZN(n6284) );
  INV_X4 U4970 ( .A(n3236), .ZN(n6285) );
  INV_X4 U4971 ( .A(n3266), .ZN(n6286) );
  INV_X4 U4972 ( .A(n3284), .ZN(n6287) );
  INV_X4 U4973 ( .A(n3204), .ZN(n6288) );
  INV_X4 U4974 ( .A(n3268), .ZN(n6289) );
  INV_X4 U4975 ( .A(n3239), .ZN(n6290) );
  INV_X4 U4976 ( .A(n3259), .ZN(n6291) );
  INV_X4 U4977 ( .A(n3207), .ZN(n6292) );
  INV_X4 U4978 ( .A(n3226), .ZN(n6293) );
  INV_X4 U4979 ( .A(n3218), .ZN(n6294) );
  INV_X4 U4980 ( .A(n3240), .ZN(n6295) );
  INV_X4 U4981 ( .A(n3237), .ZN(n6296) );
  INV_X4 U4982 ( .A(n3092), .ZN(n6297) );
  INV_X4 U4983 ( .A(n3283), .ZN(n6298) );
  INV_X4 U4984 ( .A(n3289), .ZN(n6299) );
  INV_X4 U4985 ( .A(n3246), .ZN(n6300) );
  INV_X4 U4986 ( .A(n3090), .ZN(n6301) );
  INV_X4 U4987 ( .A(n3222), .ZN(n6302) );
  INV_X4 U4988 ( .A(\u6/N52 ), .ZN(n6303) );
  INV_X4 U4989 ( .A(n3074), .ZN(n6304) );
  INV_X4 U4990 ( .A(n3741), .ZN(n6305) );
  INV_X4 U4991 ( .A(n3737), .ZN(n6306) );
  INV_X4 U4992 ( .A(n2435), .ZN(n6307) );
  INV_X4 U4993 ( .A(\u4/N5836 ), .ZN(n6308) );
  INV_X4 U4994 ( .A(n3548), .ZN(n6309) );
  INV_X4 U4995 ( .A(n3619), .ZN(n6310) );
  INV_X4 U4996 ( .A(n4249), .ZN(n6311) );
  INV_X4 U4997 ( .A(n4190), .ZN(n6313) );
  INV_X4 U4998 ( .A(n3343), .ZN(n6314) );
  INV_X4 U4999 ( .A(n2507), .ZN(n6316) );
  INV_X4 U5000 ( .A(n3297), .ZN(n6317) );
  INV_X4 U5001 ( .A(\u4/N6203 ), .ZN(n6318) );
  INV_X4 U5002 ( .A(n2699), .ZN(n6319) );
  INV_X4 U5003 ( .A(n2651), .ZN(n6320) );
  INV_X4 U5004 ( .A(n2688), .ZN(n6321) );
  INV_X4 U5005 ( .A(n2572), .ZN(n6322) );
  INV_X4 U5006 ( .A(n2690), .ZN(n6323) );
  INV_X4 U5007 ( .A(n2617), .ZN(n6324) );
  INV_X4 U5008 ( .A(n2642), .ZN(n6325) );
  INV_X4 U5009 ( .A(n2679), .ZN(n6326) );
  INV_X4 U5010 ( .A(n2632), .ZN(n6327) );
  INV_X4 U5011 ( .A(n2555), .ZN(n6328) );
  INV_X4 U5012 ( .A(n2600), .ZN(n6329) );
  INV_X4 U5013 ( .A(n2613), .ZN(n6330) );
  INV_X4 U5014 ( .A(n2615), .ZN(n6331) );
  INV_X4 U5015 ( .A(n2639), .ZN(n6332) );
  INV_X4 U5016 ( .A(n2585), .ZN(n6333) );
  INV_X4 U5017 ( .A(n2562), .ZN(n6334) );
  INV_X4 U5018 ( .A(n2647), .ZN(n6335) );
  INV_X4 U5019 ( .A(n2671), .ZN(n6336) );
  INV_X4 U5020 ( .A(n2422), .ZN(n6337) );
  INV_X4 U5021 ( .A(n2598), .ZN(n6338) );
  INV_X4 U5022 ( .A(n2439), .ZN(n6339) );
  INV_X4 U5023 ( .A(n2447), .ZN(n6340) );
  INV_X4 U5024 ( .A(n3311), .ZN(n6341) );
  INV_X4 U5025 ( .A(n2433), .ZN(n6343) );
  INV_X4 U5026 ( .A(n3879), .ZN(n6344) );
  INV_X4 U5027 ( .A(n2724), .ZN(n6345) );
  INV_X4 U5028 ( .A(n3873), .ZN(n6346) );
  INV_X4 U5029 ( .A(n2763), .ZN(n6347) );
  INV_X4 U5030 ( .A(n3171), .ZN(n6348) );
  INV_X4 U5031 ( .A(n2751), .ZN(n6349) );
  INV_X4 U5032 ( .A(n2767), .ZN(n6350) );
  INV_X4 U5033 ( .A(n2683), .ZN(n6351) );
  INV_X4 U5034 ( .A(n2599), .ZN(n6352) );
  INV_X4 U5035 ( .A(fract_denorm[91]), .ZN(n6353) );
  INV_X4 U5036 ( .A(fract_denorm[92]), .ZN(n6354) );
  INV_X4 U5037 ( .A(fract_denorm[94]), .ZN(n6355) );
  INV_X4 U5038 ( .A(fract_denorm[96]), .ZN(n6356) );
  INV_X4 U5039 ( .A(n2738), .ZN(n6357) );
  INV_X4 U5040 ( .A(fract_denorm[97]), .ZN(n6358) );
  INV_X4 U5041 ( .A(fract_denorm[90]), .ZN(n6359) );
  INV_X4 U5042 ( .A(fract_denorm[99]), .ZN(n6360) );
  INV_X4 U5043 ( .A(fract_denorm[103]), .ZN(n6361) );
  INV_X4 U5044 ( .A(fract_denorm[104]), .ZN(n6362) );
  INV_X4 U5045 ( .A(fract_denorm[101]), .ZN(n6363) );
  INV_X4 U5046 ( .A(fract_denorm[100]), .ZN(n6364) );
  INV_X4 U5047 ( .A(fract_denorm[98]), .ZN(n6365) );
  INV_X4 U5048 ( .A(n2771), .ZN(n6366) );
  INV_X4 U5049 ( .A(n2711), .ZN(n6367) );
  INV_X4 U5050 ( .A(n4097), .ZN(n6368) );
  INV_X4 U5051 ( .A(n3912), .ZN(n6369) );
  INV_X4 U5052 ( .A(fract_denorm[54]), .ZN(n6370) );
  INV_X4 U5053 ( .A(fract_denorm[56]), .ZN(n6371) );
  INV_X4 U5054 ( .A(n2750), .ZN(n6372) );
  INV_X4 U5055 ( .A(fract_denorm[57]), .ZN(n6373) );
  INV_X4 U5056 ( .A(fract_denorm[84]), .ZN(n6374) );
  INV_X4 U5057 ( .A(n2760), .ZN(n6375) );
  INV_X4 U5058 ( .A(fract_denorm[86]), .ZN(n6376) );
  INV_X4 U5059 ( .A(fract_denorm[88]), .ZN(n6377) );
  INV_X4 U5060 ( .A(n2749), .ZN(n6378) );
  INV_X4 U5061 ( .A(fract_denorm[89]), .ZN(n6379) );
  INV_X4 U5062 ( .A(n2560), .ZN(n6380) );
  INV_X4 U5063 ( .A(fract_denorm[76]), .ZN(n6381) );
  INV_X4 U5064 ( .A(n2728), .ZN(n6382) );
  INV_X4 U5065 ( .A(fract_denorm[78]), .ZN(n6383) );
  INV_X4 U5066 ( .A(fract_denorm[80]), .ZN(n6384) );
  INV_X4 U5067 ( .A(n2736), .ZN(n6385) );
  INV_X4 U5068 ( .A(fract_denorm[79]), .ZN(n6386) );
  INV_X4 U5069 ( .A(fract_denorm[59]), .ZN(n6387) );
  INV_X4 U5070 ( .A(n2705), .ZN(n6388) );
  INV_X4 U5071 ( .A(fract_denorm[62]), .ZN(n6389) );
  INV_X4 U5072 ( .A(fract_denorm[64]), .ZN(n6390) );
  INV_X4 U5073 ( .A(n2735), .ZN(n6391) );
  INV_X4 U5074 ( .A(fract_denorm[63]), .ZN(n6392) );
  INV_X4 U5075 ( .A(n2646), .ZN(n6393) );
  INV_X4 U5076 ( .A(fract_denorm[68]), .ZN(n6394) );
  INV_X4 U5077 ( .A(fract_denorm[69]), .ZN(n6395) );
  INV_X4 U5078 ( .A(n2759), .ZN(n6396) );
  INV_X4 U5079 ( .A(fract_denorm[72]), .ZN(n6397) );
  INV_X4 U5080 ( .A(n2661), .ZN(n6398) );
  INV_X4 U5081 ( .A(fract_denorm[71]), .ZN(n6399) );
  INV_X4 U5082 ( .A(fract_denorm[52]), .ZN(n6400) );
  INV_X4 U5083 ( .A(fract_denorm[58]), .ZN(n6401) );
  INV_X4 U5084 ( .A(fract_denorm[82]), .ZN(n6402) );
  INV_X4 U5085 ( .A(fract_denorm[51]), .ZN(n6403) );
  INV_X4 U5086 ( .A(fract_denorm[50]), .ZN(n6404) );
  INV_X4 U5087 ( .A(n3173), .ZN(n6405) );
  INV_X4 U5088 ( .A(n2729), .ZN(n6406) );
  INV_X4 U5089 ( .A(n3172), .ZN(n6407) );
  INV_X4 U5090 ( .A(n2737), .ZN(n6408) );
  INV_X4 U5091 ( .A(n2744), .ZN(n6409) );
  INV_X4 U5092 ( .A(n4095), .ZN(n6410) );
  INV_X4 U5093 ( .A(n3180), .ZN(n6411) );
  INV_X4 U5094 ( .A(n2561), .ZN(n6412) );
  INV_X4 U5095 ( .A(n2731), .ZN(n6413) );
  INV_X4 U5096 ( .A(n3179), .ZN(n6414) );
  INV_X4 U5097 ( .A(n2740), .ZN(n6415) );
  INV_X4 U5098 ( .A(n2745), .ZN(n6416) );
  INV_X4 U5099 ( .A(n2593), .ZN(n6417) );
  INV_X4 U5100 ( .A(n4008), .ZN(n6418) );
  INV_X4 U5101 ( .A(n3178), .ZN(n6419) );
  INV_X4 U5102 ( .A(n2762), .ZN(n6420) );
  INV_X4 U5103 ( .A(n3177), .ZN(n6421) );
  INV_X4 U5104 ( .A(n2753), .ZN(n6422) );
  INV_X4 U5105 ( .A(n2769), .ZN(n6423) );
  INV_X4 U5106 ( .A(n2685), .ZN(n6424) );
  INV_X4 U5107 ( .A(n4000), .ZN(n6425) );
  INV_X4 U5108 ( .A(n3176), .ZN(n6426) );
  INV_X4 U5109 ( .A(n2730), .ZN(n6427) );
  INV_X4 U5110 ( .A(n3175), .ZN(n6428) );
  INV_X4 U5111 ( .A(n2739), .ZN(n6429) );
  INV_X4 U5112 ( .A(n2681), .ZN(n6430) );
  INV_X4 U5113 ( .A(n2722), .ZN(n6431) );
  INV_X4 U5114 ( .A(n3992), .ZN(n6432) );
  INV_X4 U5115 ( .A(n2758), .ZN(n6433) );
  INV_X4 U5116 ( .A(n2696), .ZN(n6434) );
  INV_X4 U5117 ( .A(n3174), .ZN(n6435) );
  INV_X4 U5118 ( .A(n2752), .ZN(n6436) );
  INV_X4 U5119 ( .A(n2680), .ZN(n6437) );
  INV_X4 U5120 ( .A(n2768), .ZN(n6438) );
  INV_X4 U5121 ( .A(n3984), .ZN(n6439) );
  INV_X4 U5122 ( .A(n2633), .ZN(n6440) );
  INV_X4 U5123 ( .A(n2605), .ZN(n6441) );
  INV_X4 U5124 ( .A(n2636), .ZN(n6442) );
  INV_X4 U5125 ( .A(n3876), .ZN(n6443) );
  INV_X4 U5126 ( .A(n2718), .ZN(n6444) );
  INV_X4 U5127 ( .A(n2770), .ZN(n6445) );
  INV_X4 U5128 ( .A(n3877), .ZN(n6446) );
  INV_X4 U5129 ( .A(n3488), .ZN(n6447) );
  INV_X4 U5130 ( .A(n3913), .ZN(n6448) );
  INV_X4 U5131 ( .A(n3459), .ZN(n6449) );
  INV_X4 U5132 ( .A(n3068), .ZN(n6450) );
  INV_X4 U5133 ( .A(n3069), .ZN(n6451) );
  INV_X4 U5134 ( .A(n3070), .ZN(n6452) );
  INV_X4 U5135 ( .A(n3071), .ZN(n6453) );
  INV_X4 U5136 ( .A(n3306), .ZN(n6454) );
  INV_X4 U5137 ( .A(n3565), .ZN(n6455) );
  INV_X4 U5138 ( .A(n3457), .ZN(n6456) );
  INV_X4 U5139 ( .A(n3314), .ZN(n6457) );
  INV_X4 U5140 ( .A(n3303), .ZN(n6458) );
  INV_X4 U5141 ( .A(n3454), .ZN(n6459) );
  INV_X4 U5142 ( .A(\u4/exp_in_mi1[11] ), .ZN(n6460) );
  INV_X4 U5143 ( .A(\u4/exp_in_pl1[4] ), .ZN(n6461) );
  INV_X4 U5144 ( .A(\u4/exp_in_pl1[3] ), .ZN(n6462) );
  INV_X4 U5145 ( .A(\u4/exp_in_pl1[2] ), .ZN(n6463) );
  INV_X4 U5146 ( .A(\u4/exp_in_pl1[1] ), .ZN(n6464) );
  INV_X4 U5147 ( .A(n2514), .ZN(n6465) );
  INV_X4 U5148 ( .A(n3787), .ZN(n6466) );
  INV_X4 U5149 ( .A(\u4/N5837 ), .ZN(n6467) );
  INV_X4 U5150 ( .A(n3965), .ZN(n6468) );
>>>>>>> 19bcd6ae7dd75d2fa45f393a96c8f1177c0bf471
endmodule

