`define BIT_SIZE 63
`define EXP_SIZE 10
`define MANT_SIZE 51
`define BIAS 1023
`define EXP_SHIFT 5
