
`timescale 1ns / 100ps
module fpu ( clk, rmode, fpu_op, opa, opb, out, inf, snan, qnan, ine, overflow, 
        underflow, zero, div_by_zero );
  input [1:0] rmode;
  input [2:0] fpu_op;
  input [31:0] opa;
  input [31:0] opb;
  output [31:0] out;
  input clk;
  output inf, snan, qnan, ine, overflow, underflow, zero, div_by_zero;
  wire   inf_d, qnan_d, snan_d, opa_nan, opb_nan, opa_00, opb_00, opa_inf,
         opb_inf, opa_dn, opb_dn, sign_fasu, nan_sign_d, result_zero_sign_d,
         fasu_op, sign_fasu_r, sign_mul, sign_exe, inf_mul, inf_mul_r, N47,
         N75, N107, N141, N170, N172, N173, N174, N175, N176, N177, N178, N179,
         N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190,
         N191, N192, N193, N194, N195, N214, N215, N216, N217, N218, N219,
         N220, N221, fract_div_47_, N224, N227, N228, N229, N230, N231, N232,
         N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243,
         N244, N245, N246, N247, N248, N249, N250, N251, N298, N299, N300,
         N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311,
         N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322,
         N323, N324, N325, N391, N392, N393, N394, N395, N396, N397, N398,
         N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409,
         N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420,
         N421, opas_r1, opas_r2, sign, N441, fasu_op_r1, fasu_op_r2, inf_mul2,
         N445, N446, N447, N448, N449, N450, N451, N452, N453, N454, N455,
         N456, N457, N458, N459, N460, N461, N462, N463, N464, N465, N466,
         N467, N468, N469, N470, N471, N472, N473, N474, N475, N495, N509,
         N519, N522, N524, N526, N531, N532, opa_nan_r, N533, N540, u0_N17,
         u0_N16, u0_fractb_00, u0_fracta_00, u0_expb_00, u0_expa_00, u0_N11,
         u0_N10, u0_N7, u0_N6, u0_snan_r_b, u0_N5, u0_qnan_r_b, u0_snan_r_a,
         u0_N4, u0_qnan_r_a, u0_infb_f_r, u0_infa_f_r, u0_expb_ff, u0_expa_ff,
         u1_N140, u1_fracta_eq_fractb, u1_N131, u1_fracta_lt_fractb, u1_N130,
         u1_N129, u1_add_r, u1_signa_r, u1_sign_d, u1_fractb_lt_fracta,
         u1_adj_op_out_sft_0_, u1_adj_op_out_sft_1_, u1_adj_op_out_sft_2_,
         u1_adj_op_out_sft_3_, u1_adj_op_out_sft_4_, u1_adj_op_out_sft_5_,
         u1_adj_op_out_sft_6_, u1_adj_op_out_sft_7_, u1_adj_op_out_sft_8_,
         u1_adj_op_out_sft_9_, u1_adj_op_out_sft_10_, u1_adj_op_out_sft_11_,
         u1_adj_op_out_sft_12_, u1_adj_op_out_sft_13_, u1_adj_op_out_sft_14_,
         u1_adj_op_out_sft_15_, u1_adj_op_out_sft_16_, u1_adj_op_out_sft_17_,
         u1_adj_op_out_sft_18_, u1_adj_op_out_sft_19_, u1_adj_op_out_sft_20_,
         u1_adj_op_out_sft_21_, u1_adj_op_out_sft_22_, u1_adj_op_out_sft_23_,
         u1_adj_op_out_sft_24_, u1_adj_op_out_sft_25_, u1_adj_op_out_sft_26_,
         u1_exp_diff_sft_4_, u1_exp_lt_27, u1_adj_op_10_, u1_adj_op_17_,
         u1_adj_op_18_, u1_adj_op_19_, u1_adj_op_20_, u1_adj_op_22_, u1_N44,
         u1_N43, u1_N42, u1_N41, u1_N40, u1_N39, u1_N38, u1_N37, u1_N34,
         u1_exp_diff_0_, u1_exp_diff_1_, u1_exp_diff_2_, u1_exp_diff_3_,
         u1_exp_diff_5_, u1_exp_diff_6_, u1_exp_diff_7_, u1_expa_lt_expb,
         u2_N124, u2_N97, u2_sign_d, u2_N90, u2_N89, u2_N87, u2_exp_ovf_d_0_,
         u2_exp_ovf_d_1_, u2_N65, u2_N64, u2_N63, u2_N62, u2_N61, u2_N60,
         u2_N59, u2_N58, u2_N57, u2_N56, u2_N55, u2_N54, u2_N53, u2_N52,
         u2_N51, u2_N49, u2_N48, u2_N47, u2_N46, u2_N45, u2_N44, u2_N43,
         u2_N42, u2_exp_tmp4_0_, u2_exp_tmp4_4_, u2_exp_tmp4_7_,
         u2_exp_tmp3_0_, u2_exp_tmp3_1_, u2_exp_tmp3_2_, u2_exp_tmp3_3_,
         u2_exp_tmp3_4_, u2_exp_tmp3_5_, u2_exp_tmp3_6_, u2_exp_tmp3_7_,
         u2_N41, u2_N40, u2_N39, u2_N38, u2_N37, u2_N36, u2_N35, u2_N34,
         u2_N32, u2_N31, u2_N30, u2_N29, u2_N28, u2_N27, u2_N26, u2_N25,
         u2_exp_tmp1_0_, u2_exp_tmp1_4_, u2_N23, u2_N22, u2_N21, u2_N20,
         u2_N19, u2_N18, u2_N17, u2_N16, u2_N15, u2_N14, u2_N13, u2_N12,
         u2_N11, u2_N10, u2_N9, u2_N8, u2_N7, u2_N6, u3_N58, u3_N57, u3_N56,
         u3_N55, u3_N54, u3_N53, u3_N52, u3_N51, u3_N50, u3_N49, u3_N48,
         u3_N47, u3_N46, u3_N45, u3_N44, u3_N43, u3_N42, u3_N41, u3_N40,
         u3_N39, u3_N38, u3_N37, u3_N36, u3_N35, u3_N34, u3_N33, u3_N32,
         u3_N31, u3_N30, u3_N29, u3_N28, u3_N27, u3_N26, u3_N25, u3_N24,
         u3_N23, u3_N22, u3_N21, u3_N20, u3_N19, u3_N18, u3_N17, u3_N16,
         u3_N15, u3_N14, u3_N13, u3_N12, u3_N11, u3_N10, u3_N9, u3_N8, u3_N7,
         u3_N6, u3_N5, u3_N4, u3_N3, u5_N47, u5_N46, u5_N45, u5_N44, u5_N43,
         u5_N42, u5_N41, u5_N40, u5_N39, u5_N38, u5_N37, u5_N36, u5_N35,
         u5_N34, u5_N33, u5_N32, u5_N31, u5_N30, u5_N29, u5_N28, u5_N27,
         u5_N26, u5_N25, u5_N24, u5_N23, u5_N22, u5_N21, u5_N20, u5_N19,
         u5_N18, u5_N17, u5_N16, u5_N15, u5_N14, u5_N13, u5_N12, u5_N11,
         u5_N10, u5_N9, u5_N8, u5_N7, u5_N6, u5_N5, u5_N4, u5_N3, u5_N2, u5_N1,
         u5_N0, u6_N49, u6_N48, u6_N47, u6_N46, u6_N45, u6_N44, u6_N43, u6_N42,
         u6_N41, u6_N40, u6_N39, u6_N38, u6_N37, u6_N36, u6_N35, u6_N34,
         u6_N33, u6_N32, u6_N31, u6_N30, u6_N29, u6_N28, u6_N27, u6_N26,
         u6_N23, u6_N22, u6_N21, u6_N20, u6_N19, u6_N18, u6_N17, u6_N16,
         u6_N15, u6_N14, u6_N13, u6_N12, u6_N11, u6_N10, u6_N9, u6_N8, u6_N7,
         u6_N6, u6_N5, u6_N4, u6_N3, u6_N2, u6_N1, u6_N0, u4_N1977, u4_N1976,
         u4_N1733, u4_N1732, u4_N1731, u4_N1730, u4_N1729, u4_N1728, u4_N1727,
         u4_N1640, u4_N1606, u4_N1604, u4_N1603, u4_N1600, u4_N1599, u4_N1598,
         u4_N1573, u4_N1572, u4_N1532, u4_N1523, u4_N1504, u4_N1503,
         u4_div_exp2_0_, u4_div_exp2_1_, u4_div_exp2_2_, u4_div_exp2_3_,
         u4_div_exp2_4_, u4_div_exp2_5_, u4_div_exp2_6_, u4_div_exp2_7_,
         u4_div_exp1_0_, u4_div_exp1_1_, u4_div_exp1_2_, u4_div_exp1_3_,
         u4_div_exp1_4_, u4_div_exp1_5_, u4_div_exp1_6_, u4_div_exp1_7_,
         u4_div_exp1_8_, u4_fi_ldz_2a_0_, u4_fi_ldz_2a_1_, u4_fi_ldz_2a_3_,
         u4_fi_ldz_2a_4_, u4_fi_ldz_2a_5_, u4_ldz_all_0_, u4_ldz_all_1_,
         u4_ldz_all_2_, u4_ldz_all_3_, u4_ldz_all_4_, u4_ldz_all_5_,
         u4_ldz_all_6_, u4_N1478, u4_N1477, u4_N1476, u4_N1475, u4_N1474,
         u4_N1473, u4_N1472, u4_N1471, u4_exp_out1_1_, u4_exp_out_pl1_0_,
         u4_exp_out_pl1_1_, u4_exp_out_pl1_2_, u4_exp_out_pl1_3_,
         u4_exp_out_pl1_4_, u4_exp_out_pl1_5_, u4_exp_out_pl1_6_,
         u4_exp_out_pl1_7_, u4_fi_ldz_mi1_1_, u4_fi_ldz_mi1_2_,
         u4_fi_ldz_mi1_3_, u4_fi_ldz_mi1_4_, u4_fi_ldz_mi1_5_,
         u4_fi_ldz_mi1_6_, u4_N1455, u4_N1454, u4_N1453, u4_N1452, u4_N1451,
         u4_N1450, u4_N1449, u4_N1448, u4_N1447, u4_N1446, u4_N1445, u4_N1444,
         u4_N1443, u4_N1442, u4_N1441, u4_N1440, u4_N1439, u4_N1438, u4_N1437,
         u4_N1436, u4_N1435, u4_N1434, u4_N1433, u4_N1432, u4_N1431, u4_N1430,
         u4_N1429, u4_N1428, u4_N1427, u4_N1426, u4_N1425, u4_N1424, u4_N1423,
         u4_N1422, u4_N1421, u4_N1420, u4_N1419, u4_N1418, u4_N1417, u4_N1416,
         u4_N1415, u4_N1414, u4_N1413, u4_N1412, u4_N1411, u4_N1410, u4_N1409,
         u4_N1408, u4_N1405, u4_N1404, u4_N1403, u4_N1402, u4_N1401, u4_N1400,
         u4_N1399, u4_N1398, u4_N1397, u4_N1396, u4_N1395, u4_N1394, u4_N1393,
         u4_N1392, u4_N1391, u4_N1390, u4_N1389, u4_N1388, u4_N1387, u4_N1386,
         u4_N1385, u4_N1384, u4_N1383, u4_N1382, u4_N1381, u4_N1380, u4_N1379,
         u4_N1378, u4_N1377, u4_N1376, u4_N1375, u4_N1374, u4_N1373, u4_N1372,
         u4_N1371, u4_N1370, u4_N1369, u4_N1368, u4_N1367, u4_N1366, u4_N1365,
         u4_N1364, u4_N1363, u4_N1362, u4_N1361, u4_N1360, u4_N1359, u4_N1358,
         u4_N1356, u4_exp_in_pl1_0_, u4_exp_in_pl1_1_, u4_exp_in_pl1_2_,
         u4_exp_in_pl1_3_, u4_exp_in_pl1_4_, u4_exp_in_pl1_5_,
         u4_exp_in_pl1_6_, u4_exp_in_pl1_7_, u4_exp_in_pl1_8_, u4_f2i_shft_1_,
         u4_f2i_shft_2_, u4_f2i_shft_3_, u4_f2i_shft_4_, u4_f2i_shft_5_,
         u4_f2i_shft_6_, u4_f2i_shft_7_, u4_N1290, u4_div_shft3_0_,
         u4_div_shft3_1_, u4_div_shft3_2_, u4_div_shft3_3_, u4_div_shft3_4_,
         u4_div_shft3_5_, u4_div_shft3_6_, u4_div_shft3_7_, u4_exp_in_mi1_1_,
         u4_exp_in_mi1_2_, u4_exp_in_mi1_3_, u4_exp_in_mi1_4_,
         u4_exp_in_mi1_5_, u4_exp_in_mi1_6_, u4_exp_in_mi1_7_,
         u4_exp_in_mi1_8_, u4_N1284, u4_N1283, u4_fract_out_pl1_0_,
         u4_fract_out_pl1_1_, u4_fract_out_pl1_2_, u4_fract_out_pl1_3_,
         u4_fract_out_pl1_4_, u4_fract_out_pl1_5_, u4_fract_out_pl1_6_,
         u4_fract_out_pl1_7_, u4_fract_out_pl1_8_, u4_fract_out_pl1_9_,
         u4_fract_out_pl1_10_, u4_fract_out_pl1_11_, u4_fract_out_pl1_12_,
         u4_fract_out_pl1_13_, u4_fract_out_pl1_14_, u4_fract_out_pl1_15_,
         u4_fract_out_pl1_16_, u4_fract_out_pl1_17_, u4_fract_out_pl1_18_,
         u4_fract_out_pl1_19_, u4_fract_out_pl1_20_, u4_fract_out_pl1_21_,
         u4_fract_out_pl1_22_, u4_fract_out_pl1_23_, u4_exp_next_mi_0_,
         u4_exp_next_mi_1_, u4_exp_next_mi_2_, u4_exp_next_mi_3_,
         u4_exp_next_mi_4_, u4_exp_next_mi_5_, u4_exp_next_mi_6_,
         u4_exp_next_mi_7_, u4_exp_next_mi_8_, u4_fract_out_0_,
         u4_fract_out_1_, u4_fract_out_2_, u4_fract_out_3_, u4_fract_out_4_,
         u4_fract_out_5_, u4_fract_out_6_, u4_fract_out_7_, u4_fract_out_8_,
         u4_fract_out_9_, u4_fract_out_10_, u4_fract_out_11_, u4_fract_out_12_,
         u4_fract_out_13_, u4_fract_out_14_, u4_fract_out_15_,
         u4_fract_out_16_, u4_fract_out_17_, u4_fract_out_18_,
         u4_fract_out_19_, u4_fract_out_20_, u4_fract_out_21_,
         u4_fract_out_22_, u4_exp_out_0_, u4_exp_out_1_, u4_exp_out_2_,
         u4_exp_out_3_, u4_exp_out_4_, u4_exp_out_5_, u4_exp_out_6_,
         u4_fi_ldz_1_, u4_fi_ldz_2_, u4_fi_ldz_4_, n202, n203, n204, n1355,
         n1356, n1357, n1358, n1359, n1360, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1388, n1389, n1390, n1391, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2393, n2394, n2395, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, u4_ldz_dif_7_, u4_ldz_dif_6_,
         u4_ldz_dif_5_, u4_ldz_dif_4_, u4_ldz_dif_3_, u4_ldz_dif_2_,
         u4_ldz_dif_1_, u4_ldz_dif_0_, r489_B_0_, r524_A_5_, u2_lt_129_A_1_,
         u2_lt_129_A_2_, u2_lt_129_A_3_, u2_lt_129_A_5_, u2_lt_129_A_6_,
         u2_gt_139_B_8_, u1_gt_234_B_1_, u1_gt_234_B_2_, u1_gt_234_B_3_,
         u1_gt_234_B_4_, u1_gt_234_B_5_, u1_gt_234_B_6_, u1_gt_234_B_7_,
         u1_gt_234_B_8_, u1_gt_234_B_9_, u1_gt_234_B_10_, u1_gt_234_B_11_,
         u1_gt_234_B_12_, u1_gt_234_B_13_, u1_gt_234_B_14_, u1_gt_234_B_15_,
         u1_gt_234_B_16_, u1_gt_234_B_17_, u1_gt_234_B_18_, u1_gt_234_B_19_,
         u1_gt_234_B_20_, u1_gt_234_B_21_, u1_gt_234_B_22_, u1_gt_234_B_23_,
         u1_gt_234_B_24_, u1_gt_234_B_25_, u1_gt_234_A_0_, u1_gt_234_A_3_,
         u1_gt_234_A_4_, u1_gt_234_A_5_, u1_gt_234_A_6_, u1_gt_234_A_7_,
         u1_gt_234_A_8_, u1_gt_234_A_9_, u1_gt_234_A_10_, u1_gt_234_A_11_,
         u1_gt_234_A_12_, u1_gt_234_A_13_, u1_gt_234_A_14_, u1_gt_234_A_15_,
         u1_gt_234_A_16_, u1_gt_234_A_17_, u1_gt_234_A_18_, u1_gt_234_A_19_,
         u1_gt_234_A_20_, u1_gt_234_A_21_, u1_gt_234_A_22_, u1_gt_234_A_23_,
         u1_gt_234_A_24_, u1_gt_234_A_25_, u1_gt_234_A_26_, u1_gt_144_B_4_,
         u4_sub_465_A_0_, u4_sub_465_A_2_, u4_sub_465_A_4_, u4_sub_465_A_6_,
         u4_sub_465_A_7_, u4_sub_414_carry_2_, u4_sub_414_carry_3_,
         u4_sub_414_carry_4_, u4_sub_414_carry_5_, u4_sub_414_carry_6_,
         u4_sub_414_carry_7_, u2_sub_110_carry_2_, u2_sub_110_carry_3_,
         u2_sub_110_carry_4_, u2_sub_110_carry_5_, u2_sub_110_carry_6_,
         u2_sub_110_carry_7_, u2_sub_110_carry_8_, u2_add_110_carry_2_,
         u2_add_110_carry_3_, u2_add_110_carry_4_, u2_add_110_carry_5_,
         u2_add_110_carry_6_, u2_add_110_carry_7_, u2_add_110_carry_8_, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, u4_sub_470_n8,
         u4_sub_470_n7, u4_sub_470_n6, u4_sub_470_n5, u4_sub_470_n4,
         u4_sub_470_n3, u4_sub_470_n2, u4_sub_470_n1, u4_sub_469_n8,
         u4_sub_469_n7, u4_sub_469_n6, u4_sub_469_n5, u4_sub_469_n4,
         u4_sub_469_n3, u4_sub_469_n2, u4_sub_469_n1, u4_sll_451_n53,
         u4_sll_451_n52, u4_sll_451_n51, u4_sll_451_n50, u4_sll_451_n49,
         u4_sll_451_n48, u4_sll_451_n47, u4_sll_451_n46, u4_sll_451_n45,
         u4_sll_451_n44, u4_sll_451_n43, u4_sll_451_n42, u4_sll_451_n41,
         u4_sll_451_n40, u4_sll_451_n39, u4_sll_451_n38, u4_sll_451_n37,
         u4_sll_451_n36, u4_sll_451_n35, u4_sll_451_n34, u4_sll_451_n33,
         u4_sll_451_n32, u4_sll_451_n31, u4_sll_451_n30, u4_sll_451_n29,
         u4_sll_451_n28, u4_sll_451_n27, u4_sll_451_n26, u4_sll_451_n25,
         u4_sll_451_n24, u4_sll_451_n23, u4_sll_451_n22, u4_sll_451_n21,
         u4_sll_451_n20, u4_sll_451_n19, u4_sll_451_n18, u4_sll_451_n17,
         u4_sll_451_n16, u4_sll_451_n15, u4_sll_451_n14, u4_sll_451_n13,
         u4_sll_451_n12, u4_sll_451_n11, u4_sll_451_n10, u4_sll_451_n9,
         u4_sll_451_n8, u4_sll_451_n7, u4_sll_451_n6, u4_sll_451_n5,
         u4_sll_451_n4, u4_sll_451_n3, u4_sll_451_n2, u4_sll_451_n1,
         u4_sll_451_ML_int_5__0_, u4_sll_451_ML_int_5__1_,
         u4_sll_451_ML_int_5__2_, u4_sll_451_ML_int_5__3_,
         u4_sll_451_ML_int_5__4_, u4_sll_451_ML_int_5__5_,
         u4_sll_451_ML_int_5__6_, u4_sll_451_ML_int_5__7_,
         u4_sll_451_ML_int_5__8_, u4_sll_451_ML_int_5__9_,
         u4_sll_451_ML_int_5__10_, u4_sll_451_ML_int_5__11_,
         u4_sll_451_ML_int_5__12_, u4_sll_451_ML_int_5__13_,
         u4_sll_451_ML_int_5__14_, u4_sll_451_ML_int_5__15_,
         u4_sll_451_ML_int_5__16_, u4_sll_451_ML_int_5__17_,
         u4_sll_451_ML_int_5__18_, u4_sll_451_ML_int_5__19_,
         u4_sll_451_ML_int_5__20_, u4_sll_451_ML_int_5__21_,
         u4_sll_451_ML_int_5__22_, u4_sll_451_ML_int_5__23_,
         u4_sll_451_ML_int_5__24_, u4_sll_451_ML_int_5__25_,
         u4_sll_451_ML_int_5__26_, u4_sll_451_ML_int_5__27_,
         u4_sll_451_ML_int_5__28_, u4_sll_451_ML_int_5__29_,
         u4_sll_451_ML_int_5__30_, u4_sll_451_ML_int_5__31_,
         u4_sll_451_ML_int_5__32_, u4_sll_451_ML_int_5__33_,
         u4_sll_451_ML_int_5__34_, u4_sll_451_ML_int_5__35_,
         u4_sll_451_ML_int_5__36_, u4_sll_451_ML_int_5__37_,
         u4_sll_451_ML_int_5__38_, u4_sll_451_ML_int_5__39_,
         u4_sll_451_ML_int_5__40_, u4_sll_451_ML_int_5__41_,
         u4_sll_451_ML_int_5__42_, u4_sll_451_ML_int_5__43_,
         u4_sll_451_ML_int_5__44_, u4_sll_451_ML_int_5__45_,
         u4_sll_451_ML_int_5__46_, u4_sll_451_ML_int_5__47_,
         u4_sll_451_ML_int_4__0_, u4_sll_451_ML_int_4__1_,
         u4_sll_451_ML_int_4__2_, u4_sll_451_ML_int_4__3_,
         u4_sll_451_ML_int_4__4_, u4_sll_451_ML_int_4__5_,
         u4_sll_451_ML_int_4__6_, u4_sll_451_ML_int_4__7_,
         u4_sll_451_ML_int_4__8_, u4_sll_451_ML_int_4__9_,
         u4_sll_451_ML_int_4__10_, u4_sll_451_ML_int_4__11_,
         u4_sll_451_ML_int_4__12_, u4_sll_451_ML_int_4__13_,
         u4_sll_451_ML_int_4__14_, u4_sll_451_ML_int_4__15_,
         u4_sll_451_ML_int_4__16_, u4_sll_451_ML_int_4__17_,
         u4_sll_451_ML_int_4__18_, u4_sll_451_ML_int_4__19_,
         u4_sll_451_ML_int_4__20_, u4_sll_451_ML_int_4__21_,
         u4_sll_451_ML_int_4__22_, u4_sll_451_ML_int_4__23_,
         u4_sll_451_ML_int_4__24_, u4_sll_451_ML_int_4__25_,
         u4_sll_451_ML_int_4__26_, u4_sll_451_ML_int_4__27_,
         u4_sll_451_ML_int_4__28_, u4_sll_451_ML_int_4__29_,
         u4_sll_451_ML_int_4__30_, u4_sll_451_ML_int_4__31_,
         u4_sll_451_ML_int_4__32_, u4_sll_451_ML_int_4__33_,
         u4_sll_451_ML_int_4__34_, u4_sll_451_ML_int_4__35_,
         u4_sll_451_ML_int_4__36_, u4_sll_451_ML_int_4__37_,
         u4_sll_451_ML_int_4__38_, u4_sll_451_ML_int_4__39_,
         u4_sll_451_ML_int_4__40_, u4_sll_451_ML_int_4__41_,
         u4_sll_451_ML_int_4__42_, u4_sll_451_ML_int_4__43_,
         u4_sll_451_ML_int_4__44_, u4_sll_451_ML_int_4__45_,
         u4_sll_451_ML_int_4__46_, u4_sll_451_ML_int_4__47_,
         u4_sll_451_ML_int_3__0_, u4_sll_451_ML_int_3__1_,
         u4_sll_451_ML_int_3__2_, u4_sll_451_ML_int_3__3_,
         u4_sll_451_ML_int_3__4_, u4_sll_451_ML_int_3__5_,
         u4_sll_451_ML_int_3__6_, u4_sll_451_ML_int_3__7_,
         u4_sll_451_ML_int_3__8_, u4_sll_451_ML_int_3__9_,
         u4_sll_451_ML_int_3__10_, u4_sll_451_ML_int_3__11_,
         u4_sll_451_ML_int_3__12_, u4_sll_451_ML_int_3__13_,
         u4_sll_451_ML_int_3__14_, u4_sll_451_ML_int_3__15_,
         u4_sll_451_ML_int_3__16_, u4_sll_451_ML_int_3__17_,
         u4_sll_451_ML_int_3__18_, u4_sll_451_ML_int_3__19_,
         u4_sll_451_ML_int_3__20_, u4_sll_451_ML_int_3__21_,
         u4_sll_451_ML_int_3__22_, u4_sll_451_ML_int_3__23_,
         u4_sll_451_ML_int_3__24_, u4_sll_451_ML_int_3__25_,
         u4_sll_451_ML_int_3__26_, u4_sll_451_ML_int_3__27_,
         u4_sll_451_ML_int_3__28_, u4_sll_451_ML_int_3__29_,
         u4_sll_451_ML_int_3__30_, u4_sll_451_ML_int_3__31_,
         u4_sll_451_ML_int_3__32_, u4_sll_451_ML_int_3__33_,
         u4_sll_451_ML_int_3__34_, u4_sll_451_ML_int_3__35_,
         u4_sll_451_ML_int_3__36_, u4_sll_451_ML_int_3__37_,
         u4_sll_451_ML_int_3__38_, u4_sll_451_ML_int_3__39_,
         u4_sll_451_ML_int_3__40_, u4_sll_451_ML_int_3__41_,
         u4_sll_451_ML_int_3__42_, u4_sll_451_ML_int_3__43_,
         u4_sll_451_ML_int_3__44_, u4_sll_451_ML_int_3__45_,
         u4_sll_451_ML_int_3__46_, u4_sll_451_ML_int_3__47_,
         u4_sll_451_ML_int_2__0_, u4_sll_451_ML_int_2__1_,
         u4_sll_451_ML_int_2__2_, u4_sll_451_ML_int_2__3_,
         u4_sll_451_ML_int_2__4_, u4_sll_451_ML_int_2__5_,
         u4_sll_451_ML_int_2__6_, u4_sll_451_ML_int_2__7_,
         u4_sll_451_ML_int_2__8_, u4_sll_451_ML_int_2__9_,
         u4_sll_451_ML_int_2__10_, u4_sll_451_ML_int_2__11_,
         u4_sll_451_ML_int_2__12_, u4_sll_451_ML_int_2__13_,
         u4_sll_451_ML_int_2__14_, u4_sll_451_ML_int_2__15_,
         u4_sll_451_ML_int_2__16_, u4_sll_451_ML_int_2__17_,
         u4_sll_451_ML_int_2__18_, u4_sll_451_ML_int_2__19_,
         u4_sll_451_ML_int_2__20_, u4_sll_451_ML_int_2__21_,
         u4_sll_451_ML_int_2__22_, u4_sll_451_ML_int_2__23_,
         u4_sll_451_ML_int_2__24_, u4_sll_451_ML_int_2__25_,
         u4_sll_451_ML_int_2__26_, u4_sll_451_ML_int_2__27_,
         u4_sll_451_ML_int_2__28_, u4_sll_451_ML_int_2__29_,
         u4_sll_451_ML_int_2__30_, u4_sll_451_ML_int_2__31_,
         u4_sll_451_ML_int_2__32_, u4_sll_451_ML_int_2__33_,
         u4_sll_451_ML_int_2__34_, u4_sll_451_ML_int_2__35_,
         u4_sll_451_ML_int_2__36_, u4_sll_451_ML_int_2__37_,
         u4_sll_451_ML_int_2__38_, u4_sll_451_ML_int_2__39_,
         u4_sll_451_ML_int_2__40_, u4_sll_451_ML_int_2__41_,
         u4_sll_451_ML_int_2__42_, u4_sll_451_ML_int_2__43_,
         u4_sll_451_ML_int_2__44_, u4_sll_451_ML_int_2__45_,
         u4_sll_451_ML_int_2__46_, u4_sll_451_ML_int_2__47_,
         u4_sll_451_ML_int_1__0_, u4_sll_451_ML_int_1__1_,
         u4_sll_451_ML_int_1__2_, u4_sll_451_ML_int_1__3_,
         u4_sll_451_ML_int_1__4_, u4_sll_451_ML_int_1__5_,
         u4_sll_451_ML_int_1__6_, u4_sll_451_ML_int_1__7_,
         u4_sll_451_ML_int_1__8_, u4_sll_451_ML_int_1__9_,
         u4_sll_451_ML_int_1__10_, u4_sll_451_ML_int_1__11_,
         u4_sll_451_ML_int_1__12_, u4_sll_451_ML_int_1__13_,
         u4_sll_451_ML_int_1__14_, u4_sll_451_ML_int_1__15_,
         u4_sll_451_ML_int_1__16_, u4_sll_451_ML_int_1__17_,
         u4_sll_451_ML_int_1__18_, u4_sll_451_ML_int_1__19_,
         u4_sll_451_ML_int_1__20_, u4_sll_451_ML_int_1__21_,
         u4_sll_451_ML_int_1__22_, u4_sll_451_ML_int_1__23_,
         u4_sll_451_ML_int_1__24_, u4_sll_451_ML_int_1__25_,
         u4_sll_451_ML_int_1__26_, u4_sll_451_ML_int_1__27_,
         u4_sll_451_ML_int_1__28_, u4_sll_451_ML_int_1__29_,
         u4_sll_451_ML_int_1__30_, u4_sll_451_ML_int_1__31_,
         u4_sll_451_ML_int_1__32_, u4_sll_451_ML_int_1__33_,
         u4_sll_451_ML_int_1__34_, u4_sll_451_ML_int_1__35_,
         u4_sll_451_ML_int_1__36_, u4_sll_451_ML_int_1__37_,
         u4_sll_451_ML_int_1__38_, u4_sll_451_ML_int_1__39_,
         u4_sll_451_ML_int_1__40_, u4_sll_451_ML_int_1__41_,
         u4_sll_451_ML_int_1__42_, u4_sll_451_ML_int_1__43_,
         u4_sll_451_ML_int_1__44_, u4_sll_451_ML_int_1__45_,
         u4_sll_451_ML_int_1__46_, u4_sll_451_ML_int_1__47_, u4_srl_450_n305,
         u4_srl_450_n304, u4_srl_450_n303, u4_srl_450_n302, u4_srl_450_n301,
         u4_srl_450_n300, u4_srl_450_n299, u4_srl_450_n298, u4_srl_450_n297,
         u4_srl_450_n296, u4_srl_450_n295, u4_srl_450_n294, u4_srl_450_n293,
         u4_srl_450_n292, u4_srl_450_n291, u4_srl_450_n290, u4_srl_450_n289,
         u4_srl_450_n288, u4_srl_450_n287, u4_srl_450_n286, u4_srl_450_n285,
         u4_srl_450_n284, u4_srl_450_n283, u4_srl_450_n282, u4_srl_450_n281,
         u4_srl_450_n280, u4_srl_450_n279, u4_srl_450_n278, u4_srl_450_n277,
         u4_srl_450_n276, u4_srl_450_n275, u4_srl_450_n274, u4_srl_450_n273,
         u4_srl_450_n272, u4_srl_450_n271, u4_srl_450_n270, u4_srl_450_n269,
         u4_srl_450_n268, u4_srl_450_n267, u4_srl_450_n266, u4_srl_450_n265,
         u4_srl_450_n264, u4_srl_450_n263, u4_srl_450_n262, u4_srl_450_n261,
         u4_srl_450_n260, u4_srl_450_n259, u4_srl_450_n258, u4_srl_450_n257,
         u4_srl_450_n256, u4_srl_450_n255, u4_srl_450_n254, u4_srl_450_n253,
         u4_srl_450_n252, u4_srl_450_n251, u4_srl_450_n250, u4_srl_450_n249,
         u4_srl_450_n248, u4_srl_450_n247, u4_srl_450_n246, u4_srl_450_n245,
         u4_srl_450_n244, u4_srl_450_n243, u4_srl_450_n242, u4_srl_450_n241,
         u4_srl_450_n240, u4_srl_450_n239, u4_srl_450_n238, u4_srl_450_n237,
         u4_srl_450_n236, u4_srl_450_n235, u4_srl_450_n234, u4_srl_450_n233,
         u4_srl_450_n232, u4_srl_450_n231, u4_srl_450_n230, u4_srl_450_n229,
         u4_srl_450_n228, u4_srl_450_n227, u4_srl_450_n226, u4_srl_450_n225,
         u4_srl_450_n224, u4_srl_450_n223, u4_srl_450_n222, u4_srl_450_n221,
         u4_srl_450_n220, u4_srl_450_n219, u4_srl_450_n218, u4_srl_450_n217,
         u4_srl_450_n216, u4_srl_450_n215, u4_srl_450_n214, u4_srl_450_n213,
         u4_srl_450_n212, u4_srl_450_n211, u4_srl_450_n210, u4_srl_450_n209,
         u4_srl_450_n208, u4_srl_450_n207, u4_srl_450_n206, u4_srl_450_n205,
         u4_srl_450_n204, u4_srl_450_n203, u4_srl_450_n202, u4_srl_450_n201,
         u4_srl_450_n200, u4_srl_450_n199, u4_srl_450_n198, u4_srl_450_n197,
         u4_srl_450_n196, u4_srl_450_n195, u4_srl_450_n194, u4_srl_450_n193,
         u4_srl_450_n192, u4_srl_450_n191, u4_srl_450_n190, u4_srl_450_n189,
         u4_srl_450_n188, u4_srl_450_n187, u4_srl_450_n186, u4_srl_450_n185,
         u4_srl_450_n184, u4_srl_450_n183, u4_srl_450_n182, u4_srl_450_n181,
         u4_srl_450_n180, u4_srl_450_n179, u4_srl_450_n178, u4_srl_450_n177,
         u4_srl_450_n176, u4_srl_450_n175, u4_srl_450_n174, u4_srl_450_n173,
         u4_srl_450_n172, u4_srl_450_n171, u4_srl_450_n170, u4_srl_450_n169,
         u4_srl_450_n168, u4_srl_450_n167, u4_srl_450_n166, u4_srl_450_n165,
         u4_srl_450_n164, u4_srl_450_n163, u4_srl_450_n162, u4_srl_450_n161,
         u4_srl_450_n160, u4_srl_450_n159, u4_srl_450_n158, u4_srl_450_n157,
         u4_srl_450_n156, u4_srl_450_n155, u4_srl_450_n154, u4_srl_450_n153,
         u4_srl_450_n152, u4_srl_450_n151, u4_srl_450_n150, u4_srl_450_n149,
         u4_srl_450_n148, u4_srl_450_n147, u4_srl_450_n146, u4_srl_450_n145,
         u4_srl_450_n144, u4_srl_450_n143, u4_srl_450_n142, u4_srl_450_n141,
         u4_srl_450_n140, u4_srl_450_n139, u4_srl_450_n138, u4_srl_450_n137,
         u4_srl_450_n136, u4_srl_450_n135, u4_srl_450_n134, u4_srl_450_n133,
         u4_srl_450_n132, u4_srl_450_n131, u4_srl_450_n130, u4_srl_450_n129,
         u4_srl_450_n128, u4_srl_450_n127, u4_srl_450_n126, u4_srl_450_n125,
         u4_srl_450_n124, u4_srl_450_n123, u4_srl_450_n122, u4_srl_450_n121,
         u4_srl_450_n120, u4_srl_450_n119, u4_srl_450_n118, u4_srl_450_n117,
         u4_srl_450_n116, u4_srl_450_n115, u4_srl_450_n114, u4_srl_450_n113,
         u4_srl_450_n112, u4_srl_450_n111, u4_srl_450_n110, u4_srl_450_n109,
         u4_srl_450_n108, u4_srl_450_n107, u4_srl_450_n106, u4_srl_450_n105,
         u4_srl_450_n104, u4_srl_450_n103, u4_srl_450_n102, u4_srl_450_n101,
         u4_srl_450_n100, u4_srl_450_n99, u4_srl_450_n98, u4_srl_450_n97,
         u4_srl_450_n96, u4_srl_450_n95, u4_srl_450_n94, u4_srl_450_n93,
         u4_srl_450_n92, u4_srl_450_n91, u4_srl_450_n90, u4_srl_450_n89,
         u4_srl_450_n88, u4_srl_450_n87, u4_srl_450_n86, u4_srl_450_n85,
         u4_srl_450_n84, u4_srl_450_n83, u4_srl_450_n82, u4_srl_450_n81,
         u4_srl_450_n80, u4_srl_450_n79, u4_srl_450_n78, u4_srl_450_n77,
         u4_srl_450_n76, u4_srl_450_n75, u4_srl_450_n74, u4_srl_450_n73,
         u4_srl_450_n72, u4_srl_450_n71, u4_srl_450_n70, u4_srl_450_n69,
         u4_srl_450_n68, u4_srl_450_n67, u4_srl_450_n66, u4_srl_450_n65,
         u4_srl_450_n64, u4_srl_450_n63, u4_srl_450_n62, u4_srl_450_n61,
         u4_srl_450_n60, u4_srl_450_n59, u4_srl_450_n58, u4_srl_450_n57,
         u4_srl_450_n56, u4_srl_450_n55, u4_srl_450_n54, u4_srl_450_n53,
         u4_srl_450_n52, u4_srl_450_n51, u4_srl_450_n50, u4_srl_450_n49,
         u4_srl_450_n48, u4_srl_450_n47, u4_srl_450_n46, u4_srl_450_n45,
         u4_srl_450_n44, u4_srl_450_n43, u4_srl_450_n42, u4_srl_450_n41,
         u4_srl_450_n40, u4_srl_450_n39, u4_srl_450_n38, u4_srl_450_n37,
         u4_srl_450_n36, u4_srl_450_n35, u4_srl_450_n34, u4_srl_450_n33,
         u4_srl_450_n32, u4_srl_450_n31, u4_srl_450_n30, u4_srl_450_n29,
         u4_srl_450_n28, u4_srl_450_n27, u4_srl_450_n26, u4_srl_450_n25,
         u4_srl_450_n24, u4_srl_450_n23, u4_srl_450_n22, u4_srl_450_n21,
         u4_srl_450_n20, u4_srl_450_n19, u4_srl_450_n18, u4_srl_450_n17,
         u4_srl_450_n16, u4_srl_450_n15, u4_srl_450_n14, u4_srl_450_n13,
         u4_srl_450_n12, u4_srl_450_n11, u4_srl_450_n10, u4_srl_450_n9,
         u4_srl_450_n8, u4_srl_450_n7, u4_srl_450_n6, u4_srl_450_n5,
         u4_srl_450_n4, u4_srl_450_n3, u4_srl_450_n2, u4_srl_450_n1,
         u4_sll_479_n27, u4_sll_479_n26, u4_sll_479_n25, u4_sll_479_n24,
         u4_sll_479_n23, u4_sll_479_n22, u4_sll_479_n21, u4_sll_479_n20,
         u4_sll_479_n19, u4_sll_479_n18, u4_sll_479_n17, u4_sll_479_n16,
         u4_sll_479_n15, u4_sll_479_n14, u4_sll_479_n13, u4_sll_479_n12,
         u4_sll_479_n11, u4_sll_479_n10, u4_sll_479_n9, u4_sll_479_n8,
         u4_sll_479_n7, u4_sll_479_n6, u4_sll_479_n5, u4_sll_479_n4,
         u4_sll_479_n3, u4_sll_479_n2, u4_sll_479_n1, u4_sll_479_ML_int_6__49_,
         u4_sll_479_ML_int_6__50_, u4_sll_479_ML_int_6__51_,
         u4_sll_479_ML_int_6__52_, u4_sll_479_ML_int_6__53_,
         u4_sll_479_ML_int_6__54_, u4_sll_479_ML_int_6__55_,
         u4_sll_479_ML_int_6__56_, u4_sll_479_ML_int_5__17_,
         u4_sll_479_ML_int_5__18_, u4_sll_479_ML_int_5__19_,
         u4_sll_479_ML_int_5__20_, u4_sll_479_ML_int_5__21_,
         u4_sll_479_ML_int_5__22_, u4_sll_479_ML_int_5__23_,
         u4_sll_479_ML_int_5__24_, u4_sll_479_ML_int_5__49_,
         u4_sll_479_ML_int_5__50_, u4_sll_479_ML_int_5__51_,
         u4_sll_479_ML_int_5__52_, u4_sll_479_ML_int_5__53_,
         u4_sll_479_ML_int_5__54_, u4_sll_479_ML_int_5__55_,
         u4_sll_479_ML_int_5__56_, u4_sll_479_ML_int_4__1_,
         u4_sll_479_ML_int_4__2_, u4_sll_479_ML_int_4__3_,
         u4_sll_479_ML_int_4__4_, u4_sll_479_ML_int_4__5_,
         u4_sll_479_ML_int_4__6_, u4_sll_479_ML_int_4__7_,
         u4_sll_479_ML_int_4__8_, u4_sll_479_ML_int_4__17_,
         u4_sll_479_ML_int_4__18_, u4_sll_479_ML_int_4__19_,
         u4_sll_479_ML_int_4__20_, u4_sll_479_ML_int_4__21_,
         u4_sll_479_ML_int_4__22_, u4_sll_479_ML_int_4__23_,
         u4_sll_479_ML_int_4__24_, u4_sll_479_ML_int_4__33_,
         u4_sll_479_ML_int_4__34_, u4_sll_479_ML_int_4__35_,
         u4_sll_479_ML_int_4__36_, u4_sll_479_ML_int_4__37_,
         u4_sll_479_ML_int_4__38_, u4_sll_479_ML_int_4__39_,
         u4_sll_479_ML_int_4__40_, u4_sll_479_ML_int_4__49_,
         u4_sll_479_ML_int_4__50_, u4_sll_479_ML_int_4__51_,
         u4_sll_479_ML_int_4__52_, u4_sll_479_ML_int_4__53_,
         u4_sll_479_ML_int_4__54_, u4_sll_479_ML_int_4__55_,
         u4_sll_479_ML_int_4__56_, u4_sll_479_ML_int_3__0_,
         u4_sll_479_ML_int_3__4_, u4_sll_479_ML_int_3__5_,
         u4_sll_479_ML_int_3__6_, u4_sll_479_ML_int_3__7_,
         u4_sll_479_ML_int_3__8_, u4_sll_479_ML_int_3__9_,
         u4_sll_479_ML_int_3__10_, u4_sll_479_ML_int_3__11_,
         u4_sll_479_ML_int_3__12_, u4_sll_479_ML_int_3__13_,
         u4_sll_479_ML_int_3__14_, u4_sll_479_ML_int_3__15_,
         u4_sll_479_ML_int_3__16_, u4_sll_479_ML_int_3__17_,
         u4_sll_479_ML_int_3__18_, u4_sll_479_ML_int_3__19_,
         u4_sll_479_ML_int_3__20_, u4_sll_479_ML_int_3__21_,
         u4_sll_479_ML_int_3__22_, u4_sll_479_ML_int_3__23_,
         u4_sll_479_ML_int_3__24_, u4_sll_479_ML_int_3__25_,
         u4_sll_479_ML_int_3__26_, u4_sll_479_ML_int_3__27_,
         u4_sll_479_ML_int_3__28_, u4_sll_479_ML_int_3__29_,
         u4_sll_479_ML_int_3__30_, u4_sll_479_ML_int_3__31_,
         u4_sll_479_ML_int_3__32_, u4_sll_479_ML_int_3__33_,
         u4_sll_479_ML_int_3__34_, u4_sll_479_ML_int_3__35_,
         u4_sll_479_ML_int_3__36_, u4_sll_479_ML_int_3__37_,
         u4_sll_479_ML_int_3__38_, u4_sll_479_ML_int_3__39_,
         u4_sll_479_ML_int_3__40_, u4_sll_479_ML_int_3__41_,
         u4_sll_479_ML_int_3__42_, u4_sll_479_ML_int_3__43_,
         u4_sll_479_ML_int_3__44_, u4_sll_479_ML_int_3__45_,
         u4_sll_479_ML_int_3__46_, u4_sll_479_ML_int_3__47_,
         u4_sll_479_ML_int_3__48_, u4_sll_479_ML_int_3__49_,
         u4_sll_479_ML_int_3__50_, u4_sll_479_ML_int_3__51_,
         u4_sll_479_ML_int_3__52_, u4_sll_479_ML_int_3__53_,
         u4_sll_479_ML_int_3__54_, u4_sll_479_ML_int_3__55_,
         u4_sll_479_ML_int_3__56_, u4_sll_479_ML_int_2__1_,
         u4_sll_479_ML_int_2__2_, u4_sll_479_ML_int_2__3_,
         u4_sll_479_ML_int_2__4_, u4_sll_479_ML_int_2__5_,
         u4_sll_479_ML_int_2__6_, u4_sll_479_ML_int_2__7_,
         u4_sll_479_ML_int_2__8_, u4_sll_479_ML_int_2__9_,
         u4_sll_479_ML_int_2__10_, u4_sll_479_ML_int_2__11_,
         u4_sll_479_ML_int_2__12_, u4_sll_479_ML_int_2__13_,
         u4_sll_479_ML_int_2__14_, u4_sll_479_ML_int_2__15_,
         u4_sll_479_ML_int_2__16_, u4_sll_479_ML_int_2__17_,
         u4_sll_479_ML_int_2__18_, u4_sll_479_ML_int_2__19_,
         u4_sll_479_ML_int_2__20_, u4_sll_479_ML_int_2__21_,
         u4_sll_479_ML_int_2__22_, u4_sll_479_ML_int_2__23_,
         u4_sll_479_ML_int_2__24_, u4_sll_479_ML_int_2__25_,
         u4_sll_479_ML_int_2__26_, u4_sll_479_ML_int_2__27_,
         u4_sll_479_ML_int_2__28_, u4_sll_479_ML_int_2__29_,
         u4_sll_479_ML_int_2__30_, u4_sll_479_ML_int_2__31_,
         u4_sll_479_ML_int_2__32_, u4_sll_479_ML_int_2__33_,
         u4_sll_479_ML_int_2__34_, u4_sll_479_ML_int_2__35_,
         u4_sll_479_ML_int_2__36_, u4_sll_479_ML_int_2__37_,
         u4_sll_479_ML_int_2__38_, u4_sll_479_ML_int_2__39_,
         u4_sll_479_ML_int_2__40_, u4_sll_479_ML_int_2__41_,
         u4_sll_479_ML_int_2__42_, u4_sll_479_ML_int_2__43_,
         u4_sll_479_ML_int_2__44_, u4_sll_479_ML_int_2__45_,
         u4_sll_479_ML_int_2__46_, u4_sll_479_ML_int_2__47_,
         u4_sll_479_ML_int_2__48_, u4_sll_479_ML_int_2__49_,
         u4_sll_479_ML_int_2__50_, u4_sll_479_ML_int_2__51_,
         u4_sll_479_ML_int_2__52_, u4_sll_479_ML_int_2__53_,
         u4_sll_479_ML_int_2__54_, u4_sll_479_ML_int_2__55_,
         u4_sll_479_ML_int_2__56_, u4_sll_479_ML_int_1__0_,
         u4_sll_479_ML_int_1__1_, u4_sll_479_ML_int_1__2_,
         u4_sll_479_ML_int_1__3_, u4_sll_479_ML_int_1__4_,
         u4_sll_479_ML_int_1__5_, u4_sll_479_ML_int_1__6_,
         u4_sll_479_ML_int_1__7_, u4_sll_479_ML_int_1__8_,
         u4_sll_479_ML_int_1__9_, u4_sll_479_ML_int_1__10_,
         u4_sll_479_ML_int_1__11_, u4_sll_479_ML_int_1__12_,
         u4_sll_479_ML_int_1__13_, u4_sll_479_ML_int_1__14_,
         u4_sll_479_ML_int_1__15_, u4_sll_479_ML_int_1__16_,
         u4_sll_479_ML_int_1__17_, u4_sll_479_ML_int_1__18_,
         u4_sll_479_ML_int_1__19_, u4_sll_479_ML_int_1__20_,
         u4_sll_479_ML_int_1__21_, u4_sll_479_ML_int_1__22_,
         u4_sll_479_ML_int_1__23_, u4_sll_479_ML_int_1__24_,
         u4_sll_479_ML_int_1__25_, u4_sll_479_ML_int_1__26_,
         u4_sll_479_ML_int_1__27_, u4_sll_479_ML_int_1__28_,
         u4_sll_479_ML_int_1__29_, u4_sll_479_ML_int_1__30_,
         u4_sll_479_ML_int_1__31_, u4_sll_479_ML_int_1__32_,
         u4_sll_479_ML_int_1__33_, u4_sll_479_ML_int_1__34_,
         u4_sll_479_ML_int_1__35_, u4_sll_479_ML_int_1__36_,
         u4_sll_479_ML_int_1__37_, u4_sll_479_ML_int_1__38_,
         u4_sll_479_ML_int_1__39_, u4_sll_479_ML_int_1__40_,
         u4_sll_479_ML_int_1__41_, u4_sll_479_ML_int_1__42_,
         u4_sll_479_ML_int_1__43_, u4_sll_479_ML_int_1__44_,
         u4_sll_479_ML_int_1__45_, u4_sll_479_ML_int_1__46_,
         u4_sll_479_ML_int_1__47_, u4_sll_479_ML_int_1__48_,
         u4_sll_479_ML_int_1__49_, u4_sll_479_ML_int_1__50_,
         u4_sll_479_ML_int_1__51_, u4_sll_479_ML_int_1__52_,
         u4_sll_479_ML_int_1__53_, u4_sll_479_ML_int_1__54_,
         u4_sll_479_ML_int_1__55_, u4_sll_479_MR_int_1__55_,
         u4_sll_479_temp_int_SH_0_, u4_sll_479_temp_int_SH_1_,
         u4_sll_479_temp_int_SH_2_, u4_sll_479_temp_int_SH_3_, u4_sub_467_n10,
         u4_sub_467_n9, u4_sub_467_n8, u4_sub_467_n7, u4_sub_467_n6,
         u4_sub_467_n5, u4_sub_467_n4, u4_sub_467_n3, u4_sub_467_n2,
         u4_sub_467_n1, u4_sub_467_carry_1_, u4_sub_467_carry_2_,
         u4_sub_467_carry_3_, u4_sub_467_carry_4_, u4_sub_467_carry_5_,
         u4_sub_467_carry_6_, u4_sub_467_carry_7_, u4_sub_467_carry_8_,
         u4_sub_493_n8, u4_sub_493_n7, u4_sub_493_n6, u4_sub_493_n5,
         u4_sub_493_n4, u4_sub_493_n3, u4_sub_493_n2, u4_sub_493_n1,
         u4_add_491_n1, u4_sub_409_n14, u4_sub_409_n13, u4_sub_409_n12,
         u4_sub_409_n11, u4_sub_409_n10, u4_sub_409_n9, u4_sub_409_n8,
         u4_sub_409_n7, u4_sub_409_n6, u4_sub_409_n5, u4_sub_409_n2,
         u4_sub_409_carry_1_, u4_sub_409_carry_2_, u4_sub_409_carry_3_,
         u4_sub_409_carry_4_, u4_sub_409_carry_5_, u4_add_408_n7,
         u4_add_408_n6, u4_add_408_n5, u4_add_408_carry_2_,
         u4_add_408_carry_3_, u4_add_408_carry_4_, u4_add_408_carry_5_,
         u3_sub_60_n29, u3_sub_60_n28, u3_sub_60_n27, u3_sub_60_n26,
         u3_sub_60_n25, u3_sub_60_n24, u3_sub_60_n23, u3_sub_60_n22,
         u3_sub_60_n21, u3_sub_60_n20, u3_sub_60_n19, u3_sub_60_n18,
         u3_sub_60_n17, u3_sub_60_n16, u3_sub_60_n15, u3_sub_60_n14,
         u3_sub_60_n13, u3_sub_60_n12, u3_sub_60_n11, u3_sub_60_n10,
         u3_sub_60_n9, u3_sub_60_n8, u3_sub_60_n7, u3_sub_60_n6, u3_sub_60_n5,
         u3_sub_60_n4, u3_sub_60_n3, u3_sub_60_n1, u3_add_60_n2, u2_add_109_n2,
         u2_sub_109_n10, u2_sub_109_n9, u2_sub_109_n8, u2_sub_109_n7,
         u2_sub_109_n6, u2_sub_109_n5, u2_sub_109_n4, u2_sub_109_n3,
         u2_sub_109_n1, u1_srl_146_n141, u1_srl_146_n140, u1_srl_146_n139,
         u1_srl_146_n138, u1_srl_146_n137, u1_srl_146_n136, u1_srl_146_n135,
         u1_srl_146_n134, u1_srl_146_n133, u1_srl_146_n132, u1_srl_146_n131,
         u1_srl_146_n130, u1_srl_146_n129, u1_srl_146_n128, u1_srl_146_n127,
         u1_srl_146_n126, u1_srl_146_n125, u1_srl_146_n124, u1_srl_146_n123,
         u1_srl_146_n122, u1_srl_146_n121, u1_srl_146_n120, u1_srl_146_n119,
         u1_srl_146_n118, u1_srl_146_n117, u1_srl_146_n116, u1_srl_146_n115,
         u1_srl_146_n114, u1_srl_146_n113, u1_srl_146_n112, u1_srl_146_n111,
         u1_srl_146_n110, u1_srl_146_n109, u1_srl_146_n108, u1_srl_146_n107,
         u1_srl_146_n106, u1_srl_146_n105, u1_srl_146_n104, u1_srl_146_n103,
         u1_srl_146_n102, u1_srl_146_n101, u1_srl_146_n100, u1_srl_146_n99,
         u1_srl_146_n98, u1_srl_146_n97, u1_srl_146_n96, u1_srl_146_n95,
         u1_srl_146_n94, u1_srl_146_n93, u1_srl_146_n92, u1_srl_146_n91,
         u1_srl_146_n90, u1_srl_146_n89, u1_srl_146_n88, u1_srl_146_n87,
         u1_srl_146_n86, u1_srl_146_n85, u1_srl_146_n84, u1_srl_146_n83,
         u1_srl_146_n82, u1_srl_146_n81, u1_srl_146_n80, u1_srl_146_n79,
         u1_srl_146_n78, u1_srl_146_n77, u1_srl_146_n76, u1_srl_146_n75,
         u1_srl_146_n74, u1_srl_146_n73, u1_srl_146_n72, u1_srl_146_n71,
         u1_srl_146_n70, u1_srl_146_n69, u1_srl_146_n68, u1_srl_146_n67,
         u1_srl_146_n66, u1_srl_146_n65, u1_srl_146_n64, u1_srl_146_n63,
         u1_srl_146_n62, u1_srl_146_n61, u1_srl_146_n60, u1_srl_146_n59,
         u1_srl_146_n58, u1_srl_146_n57, u1_srl_146_n56, u1_srl_146_n55,
         u1_srl_146_n54, u1_srl_146_n53, u1_srl_146_n52, u1_srl_146_n51,
         u1_srl_146_n50, u1_srl_146_n49, u1_srl_146_n48, u1_srl_146_n47,
         u1_srl_146_n46, u1_srl_146_n45, u1_srl_146_n44, u1_srl_146_n43,
         u1_srl_146_n42, u1_srl_146_n41, u1_srl_146_n40, u1_srl_146_n39,
         u1_srl_146_n38, u1_srl_146_n37, u1_srl_146_n36, u1_srl_146_n35,
         u1_srl_146_n34, u1_srl_146_n33, u1_srl_146_n32, u1_srl_146_n31,
         u1_srl_146_n30, u1_srl_146_n29, u1_srl_146_n28, u1_srl_146_n27,
         u1_srl_146_n26, u1_srl_146_n25, u1_srl_146_n24, u1_srl_146_n23,
         u1_srl_146_n22, u1_srl_146_n21, u1_srl_146_n20, u1_srl_146_n19,
         u1_srl_146_n18, u1_srl_146_n17, u1_srl_146_n16, u1_srl_146_n15,
         u1_srl_146_n14, u1_srl_146_n13, u1_srl_146_n12, u1_srl_146_n11,
         u1_srl_146_n10, u1_srl_146_n8, u1_srl_146_n6, u1_srl_146_n5,
         u1_srl_146_n4, u1_srl_146_n3, u1_srl_146_n2, u1_srl_146_n1,
         sub_1_root_u1_sub_128_aco_n9, sub_1_root_u1_sub_128_aco_n8,
         sub_1_root_u1_sub_128_aco_n7, sub_1_root_u1_sub_128_aco_n6,
         sub_1_root_u1_sub_128_aco_n5, sub_1_root_u1_sub_128_aco_n4,
         sub_1_root_u1_sub_128_aco_n3, sub_1_root_u1_sub_128_aco_n2,
         sub_1_root_u1_sub_128_aco_n1, sub_434_3_n84, sub_434_3_n83,
         sub_434_3_n82, sub_434_3_n81, sub_434_3_n80, sub_434_3_n79,
         sub_434_3_n78, sub_434_3_n77, sub_434_3_n76, sub_434_3_n75,
         sub_434_3_n74, sub_434_3_n73, sub_434_3_n72, sub_434_3_n71,
         sub_434_3_n70, sub_434_3_n69, sub_434_3_n68, sub_434_3_n67,
         sub_434_3_n66, sub_434_3_n65, sub_434_3_n64, sub_434_3_n63,
         sub_434_3_n62, sub_434_3_n61, sub_434_3_n60, sub_434_3_n59,
         sub_434_3_n58, sub_434_3_n57, sub_434_3_n56, sub_434_3_n42,
         sub_434_3_n41, sub_434_3_n40, sub_434_3_n39, sub_434_3_n38,
         sub_434_3_n37, sub_434_3_n36, sub_434_3_n35, sub_434_3_n30,
         sub_434_3_n29, sub_434_3_n28, sub_434_3_n27, sub_434_3_n26,
         sub_434_3_n25, sub_434_3_n24, sub_434_3_n23, sub_434_3_n22,
         sub_434_3_n21, sub_434_3_n20, sub_434_3_n19, sub_434_3_n18,
         sub_434_3_n17, sub_434_3_n16, sub_434_3_n15, sub_434_3_n14,
         sub_434_3_n13, sub_434_3_n12, sub_434_b0_n70, sub_434_b0_n69,
         sub_434_b0_n68, sub_434_b0_n67, sub_434_b0_n66, sub_434_b0_n65,
         sub_434_b0_n64, sub_434_b0_n63, sub_434_b0_n62, sub_434_b0_n61,
         sub_434_b0_n60, sub_434_b0_n59, sub_434_b0_n58, sub_434_b0_n57,
         sub_434_b0_n56, sub_434_b0_n55, sub_434_b0_n54, sub_434_b0_n53,
         sub_434_b0_n52, sub_434_b0_n51, sub_434_b0_n50, sub_434_b0_n49,
         sub_434_b0_n48, sub_434_b0_n47, sub_434_b0_n25, sub_434_b0_n24,
         sub_434_b0_n23, sub_434_b0_n22, sub_434_b0_n21, sub_434_b0_n20,
         sub_434_b0_n19, sub_434_b0_n18, sub_434_b0_n17, sub_434_b0_n16,
         sub_434_b0_n15, sub_434_b0_n11, sub_434_b0_n10, sub_434_b0_n9,
         sub_434_b0_n8, sub_434_b0_n7, sub_434_b0_n6, sub_434_b0_n5,
         sub_434_b0_n4, sub_434_b0_n3, sub_434_b0_n2, sub_434_b0_n1,
         sll_384_n22, sll_384_n21, sll_384_n20, sll_384_n19, sll_384_n18,
         sll_384_n17, sll_384_n16, sll_384_n15, sll_384_n14, sll_384_n13,
         sll_384_n12, sll_384_n11, sll_384_n10, sll_384_n9, sll_384_n8,
         sll_384_n7, sll_384_n6, sll_384_n5, sll_384_n4, sll_384_n3,
         sll_384_n2, sll_384_n1, sll_384_ML_int_4__8_, sll_384_ML_int_4__9_,
         sll_384_ML_int_4__10_, sll_384_ML_int_4__11_, sll_384_ML_int_4__12_,
         sll_384_ML_int_4__13_, sll_384_ML_int_4__14_, sll_384_ML_int_4__15_,
         sll_384_ML_int_4__16_, sll_384_ML_int_4__17_, sll_384_ML_int_4__18_,
         sll_384_ML_int_4__19_, sll_384_ML_int_4__20_, sll_384_ML_int_4__21_,
         sll_384_ML_int_4__22_, sll_384_ML_int_4__23_, sll_384_ML_int_3__0_,
         sll_384_ML_int_3__1_, sll_384_ML_int_3__2_, sll_384_ML_int_3__3_,
         sll_384_ML_int_3__4_, sll_384_ML_int_3__5_, sll_384_ML_int_3__6_,
         sll_384_ML_int_3__7_, sll_384_ML_int_3__8_, sll_384_ML_int_3__9_,
         sll_384_ML_int_3__10_, sll_384_ML_int_3__11_, sll_384_ML_int_3__12_,
         sll_384_ML_int_3__13_, sll_384_ML_int_3__14_, sll_384_ML_int_3__15_,
         sll_384_ML_int_3__16_, sll_384_ML_int_3__17_, sll_384_ML_int_3__18_,
         sll_384_ML_int_3__19_, sll_384_ML_int_3__20_, sll_384_ML_int_3__21_,
         sll_384_ML_int_3__22_, sll_384_ML_int_3__23_, sll_384_ML_int_2__0_,
         sll_384_ML_int_2__1_, sll_384_ML_int_2__2_, sll_384_ML_int_2__3_,
         sll_384_ML_int_2__4_, sll_384_ML_int_2__5_, sll_384_ML_int_2__6_,
         sll_384_ML_int_2__7_, sll_384_ML_int_2__8_, sll_384_ML_int_2__9_,
         sll_384_ML_int_2__10_, sll_384_ML_int_2__11_, sll_384_ML_int_2__12_,
         sll_384_ML_int_2__13_, sll_384_ML_int_2__14_, sll_384_ML_int_2__15_,
         sll_384_ML_int_2__16_, sll_384_ML_int_2__17_, sll_384_ML_int_2__18_,
         sll_384_ML_int_2__19_, sll_384_ML_int_2__20_, sll_384_ML_int_2__21_,
         sll_384_ML_int_2__22_, sll_384_ML_int_2__23_, sll_384_ML_int_1__0_,
         sll_384_ML_int_1__1_, sll_384_ML_int_1__2_, sll_384_ML_int_1__3_,
         sll_384_ML_int_1__4_, sll_384_ML_int_1__5_, sll_384_ML_int_1__6_,
         sll_384_ML_int_1__7_, sll_384_ML_int_1__8_, sll_384_ML_int_1__9_,
         sll_384_ML_int_1__10_, sll_384_ML_int_1__11_, sll_384_ML_int_1__12_,
         sll_384_ML_int_1__13_, sll_384_ML_int_1__14_, sll_384_ML_int_1__15_,
         sll_384_ML_int_1__16_, sll_384_ML_int_1__17_, sll_384_ML_int_1__18_,
         sll_384_ML_int_1__19_, sll_384_ML_int_1__20_, sll_384_ML_int_1__21_,
         sll_384_ML_int_1__22_, sll_384_ML_int_1__23_, r473_n81, r473_n80,
         r473_n79, r473_n78, r473_n77, r473_n76, r473_n75, r473_n74, r473_n73,
         r473_n72, r473_n71, r473_n70, r473_n69, r473_n68, r473_n67, r473_n66,
         r473_n65, r473_n64, r473_n63, r473_n62, r473_n61, r473_n60, r473_n59,
         r473_n58, r473_n57, r473_n56, r473_n55, r473_n54, r473_n53, r473_n52,
         r473_n51, r473_n50, r473_n49, r473_n48, r473_n47, r473_n46, r473_n45,
         r473_n44, r473_n43, r473_n42, r473_n41, r473_n40, r473_n39, r473_n38,
         r473_n37, r473_n36, r473_n35, r473_n34, r473_n33, r473_n32, r473_n31,
         r473_n30, r473_n29, r473_n28, r473_n27, r473_n26, r473_n25, r473_n24,
         r473_n23, r473_n22, r473_n21, r473_n20, r473_n19, r473_n18, r473_n17,
         r473_n16, r473_n15, r473_n14, r473_n13, r473_n12, r473_n11, r473_n10,
         r473_n9, r473_n8, r473_n7, r473_n6, r473_n5, r473_n4, r473_n3,
         r473_n2, sub_1_root_sub_0_root_u4_add_494_n10,
         sub_1_root_sub_0_root_u4_add_494_n9,
         sub_1_root_sub_0_root_u4_add_494_n8,
         sub_1_root_sub_0_root_u4_add_494_n7,
         sub_1_root_sub_0_root_u4_add_494_n6,
         sub_1_root_sub_0_root_u4_add_494_n5,
         sub_1_root_sub_0_root_u4_add_494_n4,
         sub_1_root_sub_0_root_u4_add_494_n3,
         sub_1_root_sub_0_root_u4_add_494_n2,
         sub_1_root_sub_0_root_u4_add_494_n1,
         sub_1_root_sub_0_root_u4_add_494_carry_1_,
         sub_1_root_sub_0_root_u4_add_494_carry_2_,
         sub_1_root_sub_0_root_u4_add_494_carry_3_,
         sub_1_root_sub_0_root_u4_add_494_carry_4_,
         sub_1_root_sub_0_root_u4_add_494_carry_5_,
         sub_1_root_sub_0_root_u4_add_494_carry_6_,
         sub_1_root_sub_0_root_u4_add_494_carry_7_,
         add_0_root_sub_0_root_u4_add_494_n1, u5_mult_79_n142, u5_mult_79_n141,
         u5_mult_79_n140, u5_mult_79_n139, u5_mult_79_n138, u5_mult_79_n137,
         u5_mult_79_n136, u5_mult_79_n135, u5_mult_79_n134, u5_mult_79_n133,
         u5_mult_79_n132, u5_mult_79_n131, u5_mult_79_n130, u5_mult_79_n129,
         u5_mult_79_n128, u5_mult_79_n127, u5_mult_79_n126, u5_mult_79_n125,
         u5_mult_79_n124, u5_mult_79_n123, u5_mult_79_n122, u5_mult_79_n121,
         u5_mult_79_n120, u5_mult_79_n119, u5_mult_79_n118, u5_mult_79_n117,
         u5_mult_79_n116, u5_mult_79_n115, u5_mult_79_n114, u5_mult_79_n113,
         u5_mult_79_n112, u5_mult_79_n111, u5_mult_79_n110, u5_mult_79_n109,
         u5_mult_79_n108, u5_mult_79_n107, u5_mult_79_n106, u5_mult_79_n105,
         u5_mult_79_n104, u5_mult_79_n103, u5_mult_79_n102, u5_mult_79_n101,
         u5_mult_79_n100, u5_mult_79_n99, u5_mult_79_n98, u5_mult_79_n97,
         u5_mult_79_n96, u5_mult_79_n95, u5_mult_79_n93, u5_mult_79_n92,
         u5_mult_79_n90, u5_mult_79_n89, u5_mult_79_n88, u5_mult_79_n87,
         u5_mult_79_n86, u5_mult_79_n85, u5_mult_79_n84, u5_mult_79_n83,
         u5_mult_79_n82, u5_mult_79_n81, u5_mult_79_n80, u5_mult_79_n79,
         u5_mult_79_n78, u5_mult_79_n77, u5_mult_79_n76, u5_mult_79_n75,
         u5_mult_79_n74, u5_mult_79_n73, u5_mult_79_n72, u5_mult_79_n71,
         u5_mult_79_n70, u5_mult_79_n69, u5_mult_79_n68, u5_mult_79_n67,
         u5_mult_79_n66, u5_mult_79_n65, u5_mult_79_n64, u5_mult_79_n63,
         u5_mult_79_n62, u5_mult_79_n61, u5_mult_79_n60, u5_mult_79_n59,
         u5_mult_79_n58, u5_mult_79_n57, u5_mult_79_n56, u5_mult_79_n55,
         u5_mult_79_n54, u5_mult_79_n53, u5_mult_79_n52, u5_mult_79_n51,
         u5_mult_79_n50, u5_mult_79_n49, u5_mult_79_n48, u5_mult_79_n47,
         u5_mult_79_n46, u5_mult_79_n45, u5_mult_79_n44, u5_mult_79_n43,
         u5_mult_79_n42, u5_mult_79_n41, u5_mult_79_n40, u5_mult_79_n39,
         u5_mult_79_n38, u5_mult_79_n37, u5_mult_79_n36, u5_mult_79_n35,
         u5_mult_79_n34, u5_mult_79_n33, u5_mult_79_n32, u5_mult_79_n31,
         u5_mult_79_n30, u5_mult_79_n29, u5_mult_79_n28, u5_mult_79_n27,
         u5_mult_79_n26, u5_mult_79_n25, u5_mult_79_n24, u5_mult_79_n23,
         u5_mult_79_n22, u5_mult_79_n21, u5_mult_79_n20, u5_mult_79_n19,
         u5_mult_79_n18, u5_mult_79_n17, u5_mult_79_n16, u5_mult_79_n15,
         u5_mult_79_n14, u5_mult_79_n13, u5_mult_79_n12, u5_mult_79_n11,
         u5_mult_79_n10, u5_mult_79_n9, u5_mult_79_n8, u5_mult_79_n7,
         u5_mult_79_n6, u5_mult_79_n5, u5_mult_79_n4, u5_mult_79_n3,
         u5_mult_79_SUMB_2__1_, u5_mult_79_SUMB_2__2_, u5_mult_79_SUMB_2__3_,
         u5_mult_79_SUMB_2__4_, u5_mult_79_SUMB_2__5_, u5_mult_79_SUMB_2__6_,
         u5_mult_79_SUMB_2__7_, u5_mult_79_SUMB_2__8_, u5_mult_79_SUMB_2__9_,
         u5_mult_79_SUMB_2__10_, u5_mult_79_SUMB_2__11_,
         u5_mult_79_SUMB_2__12_, u5_mult_79_SUMB_2__13_,
         u5_mult_79_SUMB_2__14_, u5_mult_79_SUMB_2__15_,
         u5_mult_79_SUMB_2__16_, u5_mult_79_SUMB_2__17_,
         u5_mult_79_SUMB_2__18_, u5_mult_79_SUMB_2__19_,
         u5_mult_79_SUMB_2__20_, u5_mult_79_SUMB_2__21_,
         u5_mult_79_SUMB_2__22_, u5_mult_79_SUMB_3__1_, u5_mult_79_SUMB_3__2_,
         u5_mult_79_SUMB_3__3_, u5_mult_79_SUMB_3__4_, u5_mult_79_SUMB_3__5_,
         u5_mult_79_SUMB_3__6_, u5_mult_79_SUMB_3__7_, u5_mult_79_SUMB_3__8_,
         u5_mult_79_SUMB_3__9_, u5_mult_79_SUMB_3__10_, u5_mult_79_SUMB_3__11_,
         u5_mult_79_SUMB_3__12_, u5_mult_79_SUMB_3__13_,
         u5_mult_79_SUMB_3__14_, u5_mult_79_SUMB_3__15_,
         u5_mult_79_SUMB_3__16_, u5_mult_79_SUMB_3__17_,
         u5_mult_79_SUMB_3__18_, u5_mult_79_SUMB_3__19_,
         u5_mult_79_SUMB_3__20_, u5_mult_79_SUMB_3__21_,
         u5_mult_79_SUMB_3__22_, u5_mult_79_SUMB_4__1_, u5_mult_79_SUMB_4__2_,
         u5_mult_79_SUMB_4__3_, u5_mult_79_SUMB_4__4_, u5_mult_79_SUMB_4__5_,
         u5_mult_79_SUMB_4__6_, u5_mult_79_SUMB_4__7_, u5_mult_79_SUMB_4__8_,
         u5_mult_79_SUMB_4__9_, u5_mult_79_SUMB_4__10_, u5_mult_79_SUMB_4__11_,
         u5_mult_79_SUMB_4__12_, u5_mult_79_SUMB_4__13_,
         u5_mult_79_SUMB_4__14_, u5_mult_79_SUMB_4__15_,
         u5_mult_79_SUMB_4__16_, u5_mult_79_SUMB_4__17_,
         u5_mult_79_SUMB_4__18_, u5_mult_79_SUMB_4__19_,
         u5_mult_79_SUMB_4__20_, u5_mult_79_SUMB_4__21_,
         u5_mult_79_SUMB_4__22_, u5_mult_79_SUMB_5__1_, u5_mult_79_SUMB_5__2_,
         u5_mult_79_SUMB_5__3_, u5_mult_79_SUMB_5__4_, u5_mult_79_SUMB_5__5_,
         u5_mult_79_SUMB_5__6_, u5_mult_79_SUMB_5__7_, u5_mult_79_SUMB_5__8_,
         u5_mult_79_SUMB_5__9_, u5_mult_79_SUMB_5__10_, u5_mult_79_SUMB_5__11_,
         u5_mult_79_SUMB_5__12_, u5_mult_79_SUMB_5__13_,
         u5_mult_79_SUMB_5__14_, u5_mult_79_SUMB_5__15_,
         u5_mult_79_SUMB_5__16_, u5_mult_79_SUMB_5__17_,
         u5_mult_79_SUMB_5__18_, u5_mult_79_SUMB_5__19_,
         u5_mult_79_SUMB_5__20_, u5_mult_79_SUMB_5__21_,
         u5_mult_79_SUMB_5__22_, u5_mult_79_SUMB_6__1_, u5_mult_79_SUMB_6__2_,
         u5_mult_79_SUMB_6__3_, u5_mult_79_SUMB_6__4_, u5_mult_79_SUMB_6__5_,
         u5_mult_79_SUMB_6__6_, u5_mult_79_SUMB_6__7_, u5_mult_79_SUMB_6__8_,
         u5_mult_79_SUMB_6__9_, u5_mult_79_SUMB_6__10_, u5_mult_79_SUMB_6__11_,
         u5_mult_79_SUMB_6__12_, u5_mult_79_SUMB_6__13_,
         u5_mult_79_SUMB_6__14_, u5_mult_79_SUMB_6__15_,
         u5_mult_79_SUMB_6__16_, u5_mult_79_SUMB_6__17_,
         u5_mult_79_SUMB_6__18_, u5_mult_79_SUMB_6__19_,
         u5_mult_79_SUMB_6__20_, u5_mult_79_SUMB_6__21_,
         u5_mult_79_SUMB_6__22_, u5_mult_79_SUMB_7__1_, u5_mult_79_SUMB_7__2_,
         u5_mult_79_SUMB_7__3_, u5_mult_79_SUMB_7__4_, u5_mult_79_SUMB_7__5_,
         u5_mult_79_SUMB_7__6_, u5_mult_79_SUMB_7__7_, u5_mult_79_SUMB_7__8_,
         u5_mult_79_SUMB_7__9_, u5_mult_79_SUMB_7__10_, u5_mult_79_SUMB_7__11_,
         u5_mult_79_SUMB_7__12_, u5_mult_79_SUMB_7__13_,
         u5_mult_79_SUMB_7__14_, u5_mult_79_SUMB_7__15_,
         u5_mult_79_SUMB_7__16_, u5_mult_79_SUMB_7__17_,
         u5_mult_79_SUMB_7__18_, u5_mult_79_SUMB_7__19_,
         u5_mult_79_SUMB_7__20_, u5_mult_79_SUMB_7__21_,
         u5_mult_79_SUMB_7__22_, u5_mult_79_SUMB_8__1_, u5_mult_79_SUMB_8__2_,
         u5_mult_79_SUMB_8__3_, u5_mult_79_SUMB_8__4_, u5_mult_79_SUMB_8__5_,
         u5_mult_79_SUMB_8__6_, u5_mult_79_SUMB_8__7_, u5_mult_79_SUMB_8__8_,
         u5_mult_79_SUMB_8__9_, u5_mult_79_SUMB_8__10_, u5_mult_79_SUMB_8__11_,
         u5_mult_79_SUMB_8__12_, u5_mult_79_SUMB_8__13_,
         u5_mult_79_SUMB_8__14_, u5_mult_79_SUMB_8__15_,
         u5_mult_79_SUMB_8__16_, u5_mult_79_SUMB_8__17_,
         u5_mult_79_SUMB_8__18_, u5_mult_79_SUMB_8__19_,
         u5_mult_79_SUMB_8__20_, u5_mult_79_SUMB_8__21_,
         u5_mult_79_SUMB_8__22_, u5_mult_79_SUMB_9__1_, u5_mult_79_SUMB_9__2_,
         u5_mult_79_SUMB_9__3_, u5_mult_79_SUMB_9__4_, u5_mult_79_SUMB_9__5_,
         u5_mult_79_SUMB_9__6_, u5_mult_79_SUMB_9__7_, u5_mult_79_SUMB_9__8_,
         u5_mult_79_SUMB_9__9_, u5_mult_79_SUMB_9__10_, u5_mult_79_SUMB_9__11_,
         u5_mult_79_SUMB_9__12_, u5_mult_79_SUMB_9__13_,
         u5_mult_79_SUMB_9__14_, u5_mult_79_SUMB_9__15_,
         u5_mult_79_SUMB_9__16_, u5_mult_79_SUMB_9__17_,
         u5_mult_79_SUMB_9__18_, u5_mult_79_SUMB_9__19_,
         u5_mult_79_SUMB_9__20_, u5_mult_79_SUMB_9__21_,
         u5_mult_79_SUMB_9__22_, u5_mult_79_SUMB_10__1_,
         u5_mult_79_SUMB_10__2_, u5_mult_79_SUMB_10__3_,
         u5_mult_79_SUMB_10__4_, u5_mult_79_SUMB_10__5_,
         u5_mult_79_SUMB_10__6_, u5_mult_79_SUMB_10__7_,
         u5_mult_79_SUMB_10__8_, u5_mult_79_SUMB_10__9_,
         u5_mult_79_SUMB_10__10_, u5_mult_79_SUMB_10__11_,
         u5_mult_79_SUMB_10__12_, u5_mult_79_SUMB_10__13_,
         u5_mult_79_SUMB_10__14_, u5_mult_79_SUMB_10__15_,
         u5_mult_79_SUMB_10__16_, u5_mult_79_SUMB_10__17_,
         u5_mult_79_SUMB_10__18_, u5_mult_79_SUMB_10__19_,
         u5_mult_79_SUMB_10__20_, u5_mult_79_SUMB_10__21_,
         u5_mult_79_SUMB_10__22_, u5_mult_79_SUMB_11__1_,
         u5_mult_79_SUMB_11__2_, u5_mult_79_SUMB_11__3_,
         u5_mult_79_SUMB_11__4_, u5_mult_79_SUMB_11__5_,
         u5_mult_79_SUMB_11__6_, u5_mult_79_SUMB_11__7_,
         u5_mult_79_SUMB_11__8_, u5_mult_79_SUMB_11__9_,
         u5_mult_79_SUMB_11__10_, u5_mult_79_SUMB_11__11_,
         u5_mult_79_SUMB_11__12_, u5_mult_79_SUMB_11__13_,
         u5_mult_79_SUMB_11__14_, u5_mult_79_SUMB_11__15_,
         u5_mult_79_SUMB_11__16_, u5_mult_79_SUMB_11__17_,
         u5_mult_79_SUMB_11__18_, u5_mult_79_SUMB_11__19_,
         u5_mult_79_SUMB_11__20_, u5_mult_79_SUMB_11__21_,
         u5_mult_79_SUMB_11__22_, u5_mult_79_SUMB_12__1_,
         u5_mult_79_SUMB_12__2_, u5_mult_79_SUMB_12__3_,
         u5_mult_79_SUMB_12__4_, u5_mult_79_SUMB_12__5_,
         u5_mult_79_SUMB_12__6_, u5_mult_79_SUMB_12__7_,
         u5_mult_79_SUMB_12__8_, u5_mult_79_SUMB_12__9_,
         u5_mult_79_SUMB_12__10_, u5_mult_79_SUMB_12__11_,
         u5_mult_79_SUMB_12__12_, u5_mult_79_SUMB_12__13_,
         u5_mult_79_SUMB_12__14_, u5_mult_79_SUMB_12__15_,
         u5_mult_79_SUMB_12__16_, u5_mult_79_SUMB_12__17_,
         u5_mult_79_SUMB_12__18_, u5_mult_79_SUMB_12__19_,
         u5_mult_79_SUMB_12__20_, u5_mult_79_SUMB_12__21_,
         u5_mult_79_SUMB_12__22_, u5_mult_79_SUMB_13__1_,
         u5_mult_79_SUMB_13__2_, u5_mult_79_SUMB_13__3_,
         u5_mult_79_SUMB_13__4_, u5_mult_79_SUMB_13__5_,
         u5_mult_79_SUMB_13__6_, u5_mult_79_SUMB_13__7_,
         u5_mult_79_SUMB_13__8_, u5_mult_79_SUMB_13__9_,
         u5_mult_79_SUMB_13__10_, u5_mult_79_SUMB_13__11_,
         u5_mult_79_SUMB_13__12_, u5_mult_79_SUMB_13__13_,
         u5_mult_79_SUMB_13__14_, u5_mult_79_SUMB_13__15_,
         u5_mult_79_SUMB_13__16_, u5_mult_79_SUMB_13__17_,
         u5_mult_79_SUMB_13__18_, u5_mult_79_SUMB_13__19_,
         u5_mult_79_SUMB_13__20_, u5_mult_79_SUMB_13__21_,
         u5_mult_79_SUMB_13__22_, u5_mult_79_SUMB_14__1_,
         u5_mult_79_SUMB_14__2_, u5_mult_79_SUMB_14__3_,
         u5_mult_79_SUMB_14__4_, u5_mult_79_SUMB_14__5_,
         u5_mult_79_SUMB_14__6_, u5_mult_79_SUMB_14__7_,
         u5_mult_79_SUMB_14__8_, u5_mult_79_SUMB_14__9_,
         u5_mult_79_SUMB_14__10_, u5_mult_79_SUMB_14__11_,
         u5_mult_79_SUMB_14__12_, u5_mult_79_SUMB_14__13_,
         u5_mult_79_SUMB_14__14_, u5_mult_79_SUMB_14__15_,
         u5_mult_79_SUMB_14__16_, u5_mult_79_SUMB_14__17_,
         u5_mult_79_SUMB_14__18_, u5_mult_79_SUMB_14__19_,
         u5_mult_79_SUMB_14__20_, u5_mult_79_SUMB_14__21_,
         u5_mult_79_SUMB_14__22_, u5_mult_79_SUMB_15__1_,
         u5_mult_79_SUMB_15__2_, u5_mult_79_SUMB_15__3_,
         u5_mult_79_SUMB_15__4_, u5_mult_79_SUMB_15__5_,
         u5_mult_79_SUMB_15__6_, u5_mult_79_SUMB_15__7_,
         u5_mult_79_SUMB_15__8_, u5_mult_79_SUMB_15__9_,
         u5_mult_79_SUMB_15__10_, u5_mult_79_SUMB_15__11_,
         u5_mult_79_SUMB_15__12_, u5_mult_79_SUMB_15__13_,
         u5_mult_79_SUMB_15__14_, u5_mult_79_SUMB_15__15_,
         u5_mult_79_SUMB_15__16_, u5_mult_79_SUMB_15__17_,
         u5_mult_79_SUMB_15__18_, u5_mult_79_SUMB_15__19_,
         u5_mult_79_SUMB_15__20_, u5_mult_79_SUMB_15__21_,
         u5_mult_79_SUMB_15__22_, u5_mult_79_SUMB_16__1_,
         u5_mult_79_SUMB_16__2_, u5_mult_79_SUMB_16__3_,
         u5_mult_79_SUMB_16__4_, u5_mult_79_SUMB_16__5_,
         u5_mult_79_SUMB_16__6_, u5_mult_79_SUMB_16__7_,
         u5_mult_79_SUMB_16__8_, u5_mult_79_SUMB_16__9_,
         u5_mult_79_SUMB_16__10_, u5_mult_79_SUMB_16__11_,
         u5_mult_79_SUMB_16__12_, u5_mult_79_SUMB_16__13_,
         u5_mult_79_SUMB_16__14_, u5_mult_79_SUMB_16__15_,
         u5_mult_79_SUMB_16__16_, u5_mult_79_SUMB_16__17_,
         u5_mult_79_SUMB_16__18_, u5_mult_79_SUMB_16__19_,
         u5_mult_79_SUMB_16__20_, u5_mult_79_SUMB_16__21_,
         u5_mult_79_SUMB_16__22_, u5_mult_79_SUMB_17__1_,
         u5_mult_79_SUMB_17__2_, u5_mult_79_SUMB_17__3_,
         u5_mult_79_SUMB_17__4_, u5_mult_79_SUMB_17__5_,
         u5_mult_79_SUMB_17__6_, u5_mult_79_SUMB_17__7_,
         u5_mult_79_SUMB_17__8_, u5_mult_79_SUMB_17__9_,
         u5_mult_79_SUMB_17__10_, u5_mult_79_SUMB_17__11_,
         u5_mult_79_SUMB_17__12_, u5_mult_79_SUMB_17__13_,
         u5_mult_79_SUMB_17__14_, u5_mult_79_SUMB_17__15_,
         u5_mult_79_SUMB_17__16_, u5_mult_79_SUMB_17__17_,
         u5_mult_79_SUMB_17__18_, u5_mult_79_SUMB_17__19_,
         u5_mult_79_SUMB_17__20_, u5_mult_79_SUMB_17__21_,
         u5_mult_79_SUMB_17__22_, u5_mult_79_SUMB_18__1_,
         u5_mult_79_SUMB_18__2_, u5_mult_79_SUMB_18__3_,
         u5_mult_79_SUMB_18__4_, u5_mult_79_SUMB_18__5_,
         u5_mult_79_SUMB_18__6_, u5_mult_79_SUMB_18__7_,
         u5_mult_79_SUMB_18__8_, u5_mult_79_SUMB_18__9_,
         u5_mult_79_SUMB_18__10_, u5_mult_79_SUMB_18__11_,
         u5_mult_79_SUMB_18__12_, u5_mult_79_SUMB_18__13_,
         u5_mult_79_SUMB_18__14_, u5_mult_79_SUMB_18__15_,
         u5_mult_79_SUMB_18__16_, u5_mult_79_SUMB_18__17_,
         u5_mult_79_SUMB_18__18_, u5_mult_79_SUMB_18__19_,
         u5_mult_79_SUMB_18__20_, u5_mult_79_SUMB_18__21_,
         u5_mult_79_SUMB_18__22_, u5_mult_79_SUMB_19__1_,
         u5_mult_79_SUMB_19__2_, u5_mult_79_SUMB_19__3_,
         u5_mult_79_SUMB_19__4_, u5_mult_79_SUMB_19__5_,
         u5_mult_79_SUMB_19__6_, u5_mult_79_SUMB_19__7_,
         u5_mult_79_SUMB_19__8_, u5_mult_79_SUMB_19__9_,
         u5_mult_79_SUMB_19__10_, u5_mult_79_SUMB_19__11_,
         u5_mult_79_SUMB_19__12_, u5_mult_79_SUMB_19__13_,
         u5_mult_79_SUMB_19__14_, u5_mult_79_SUMB_19__15_,
         u5_mult_79_SUMB_19__16_, u5_mult_79_SUMB_19__17_,
         u5_mult_79_SUMB_19__18_, u5_mult_79_SUMB_19__19_,
         u5_mult_79_SUMB_19__20_, u5_mult_79_SUMB_19__21_,
         u5_mult_79_SUMB_19__22_, u5_mult_79_SUMB_20__1_,
         u5_mult_79_SUMB_20__2_, u5_mult_79_SUMB_20__3_,
         u5_mult_79_SUMB_20__4_, u5_mult_79_SUMB_20__5_,
         u5_mult_79_SUMB_20__6_, u5_mult_79_SUMB_20__7_,
         u5_mult_79_SUMB_20__8_, u5_mult_79_SUMB_20__9_,
         u5_mult_79_SUMB_20__10_, u5_mult_79_SUMB_20__11_,
         u5_mult_79_SUMB_20__12_, u5_mult_79_SUMB_20__13_,
         u5_mult_79_SUMB_20__14_, u5_mult_79_SUMB_20__15_,
         u5_mult_79_SUMB_20__16_, u5_mult_79_SUMB_20__17_,
         u5_mult_79_SUMB_20__18_, u5_mult_79_SUMB_20__19_,
         u5_mult_79_SUMB_20__20_, u5_mult_79_SUMB_20__21_,
         u5_mult_79_SUMB_20__22_, u5_mult_79_SUMB_21__1_,
         u5_mult_79_SUMB_21__2_, u5_mult_79_SUMB_21__3_,
         u5_mult_79_SUMB_21__4_, u5_mult_79_SUMB_21__5_,
         u5_mult_79_SUMB_21__6_, u5_mult_79_SUMB_21__7_,
         u5_mult_79_SUMB_21__8_, u5_mult_79_SUMB_21__9_,
         u5_mult_79_SUMB_21__10_, u5_mult_79_SUMB_21__11_,
         u5_mult_79_SUMB_21__12_, u5_mult_79_SUMB_21__13_,
         u5_mult_79_SUMB_21__14_, u5_mult_79_SUMB_21__15_,
         u5_mult_79_SUMB_21__16_, u5_mult_79_SUMB_21__17_,
         u5_mult_79_SUMB_21__18_, u5_mult_79_SUMB_21__19_,
         u5_mult_79_SUMB_21__20_, u5_mult_79_SUMB_21__21_,
         u5_mult_79_SUMB_21__22_, u5_mult_79_SUMB_22__1_,
         u5_mult_79_SUMB_22__2_, u5_mult_79_SUMB_22__3_,
         u5_mult_79_SUMB_22__4_, u5_mult_79_SUMB_22__5_,
         u5_mult_79_SUMB_22__6_, u5_mult_79_SUMB_22__7_,
         u5_mult_79_SUMB_22__8_, u5_mult_79_SUMB_22__9_,
         u5_mult_79_SUMB_22__10_, u5_mult_79_SUMB_22__11_,
         u5_mult_79_SUMB_22__12_, u5_mult_79_SUMB_22__13_,
         u5_mult_79_SUMB_22__14_, u5_mult_79_SUMB_22__15_,
         u5_mult_79_SUMB_22__16_, u5_mult_79_SUMB_22__17_,
         u5_mult_79_SUMB_22__18_, u5_mult_79_SUMB_22__19_,
         u5_mult_79_SUMB_22__20_, u5_mult_79_SUMB_22__21_,
         u5_mult_79_SUMB_22__22_, u5_mult_79_SUMB_23__1_,
         u5_mult_79_SUMB_23__2_, u5_mult_79_SUMB_23__3_,
         u5_mult_79_SUMB_23__4_, u5_mult_79_SUMB_23__5_,
         u5_mult_79_SUMB_23__6_, u5_mult_79_SUMB_23__7_,
         u5_mult_79_SUMB_23__8_, u5_mult_79_SUMB_23__9_,
         u5_mult_79_SUMB_23__10_, u5_mult_79_SUMB_23__11_,
         u5_mult_79_SUMB_23__12_, u5_mult_79_SUMB_23__13_,
         u5_mult_79_SUMB_23__14_, u5_mult_79_SUMB_23__15_,
         u5_mult_79_SUMB_23__16_, u5_mult_79_SUMB_23__17_,
         u5_mult_79_SUMB_23__18_, u5_mult_79_SUMB_23__19_,
         u5_mult_79_SUMB_23__20_, u5_mult_79_SUMB_23__21_,
         u5_mult_79_SUMB_23__22_, u5_mult_79_CARRYB_2__0_,
         u5_mult_79_CARRYB_2__1_, u5_mult_79_CARRYB_2__2_,
         u5_mult_79_CARRYB_2__3_, u5_mult_79_CARRYB_2__4_,
         u5_mult_79_CARRYB_2__5_, u5_mult_79_CARRYB_2__6_,
         u5_mult_79_CARRYB_2__7_, u5_mult_79_CARRYB_2__8_,
         u5_mult_79_CARRYB_2__9_, u5_mult_79_CARRYB_2__10_,
         u5_mult_79_CARRYB_2__11_, u5_mult_79_CARRYB_2__12_,
         u5_mult_79_CARRYB_2__13_, u5_mult_79_CARRYB_2__14_,
         u5_mult_79_CARRYB_2__15_, u5_mult_79_CARRYB_2__16_,
         u5_mult_79_CARRYB_2__17_, u5_mult_79_CARRYB_2__18_,
         u5_mult_79_CARRYB_2__19_, u5_mult_79_CARRYB_2__20_,
         u5_mult_79_CARRYB_2__21_, u5_mult_79_CARRYB_2__22_,
         u5_mult_79_CARRYB_3__0_, u5_mult_79_CARRYB_3__1_,
         u5_mult_79_CARRYB_3__2_, u5_mult_79_CARRYB_3__3_,
         u5_mult_79_CARRYB_3__4_, u5_mult_79_CARRYB_3__5_,
         u5_mult_79_CARRYB_3__6_, u5_mult_79_CARRYB_3__7_,
         u5_mult_79_CARRYB_3__8_, u5_mult_79_CARRYB_3__9_,
         u5_mult_79_CARRYB_3__10_, u5_mult_79_CARRYB_3__11_,
         u5_mult_79_CARRYB_3__12_, u5_mult_79_CARRYB_3__13_,
         u5_mult_79_CARRYB_3__14_, u5_mult_79_CARRYB_3__15_,
         u5_mult_79_CARRYB_3__16_, u5_mult_79_CARRYB_3__17_,
         u5_mult_79_CARRYB_3__18_, u5_mult_79_CARRYB_3__19_,
         u5_mult_79_CARRYB_3__20_, u5_mult_79_CARRYB_3__21_,
         u5_mult_79_CARRYB_3__22_, u5_mult_79_CARRYB_4__0_,
         u5_mult_79_CARRYB_4__1_, u5_mult_79_CARRYB_4__2_,
         u5_mult_79_CARRYB_4__3_, u5_mult_79_CARRYB_4__4_,
         u5_mult_79_CARRYB_4__5_, u5_mult_79_CARRYB_4__6_,
         u5_mult_79_CARRYB_4__7_, u5_mult_79_CARRYB_4__8_,
         u5_mult_79_CARRYB_4__9_, u5_mult_79_CARRYB_4__10_,
         u5_mult_79_CARRYB_4__11_, u5_mult_79_CARRYB_4__12_,
         u5_mult_79_CARRYB_4__13_, u5_mult_79_CARRYB_4__14_,
         u5_mult_79_CARRYB_4__15_, u5_mult_79_CARRYB_4__16_,
         u5_mult_79_CARRYB_4__17_, u5_mult_79_CARRYB_4__18_,
         u5_mult_79_CARRYB_4__19_, u5_mult_79_CARRYB_4__20_,
         u5_mult_79_CARRYB_4__21_, u5_mult_79_CARRYB_4__22_,
         u5_mult_79_CARRYB_5__0_, u5_mult_79_CARRYB_5__1_,
         u5_mult_79_CARRYB_5__2_, u5_mult_79_CARRYB_5__3_,
         u5_mult_79_CARRYB_5__4_, u5_mult_79_CARRYB_5__5_,
         u5_mult_79_CARRYB_5__6_, u5_mult_79_CARRYB_5__7_,
         u5_mult_79_CARRYB_5__8_, u5_mult_79_CARRYB_5__9_,
         u5_mult_79_CARRYB_5__10_, u5_mult_79_CARRYB_5__11_,
         u5_mult_79_CARRYB_5__12_, u5_mult_79_CARRYB_5__13_,
         u5_mult_79_CARRYB_5__14_, u5_mult_79_CARRYB_5__15_,
         u5_mult_79_CARRYB_5__16_, u5_mult_79_CARRYB_5__17_,
         u5_mult_79_CARRYB_5__18_, u5_mult_79_CARRYB_5__19_,
         u5_mult_79_CARRYB_5__20_, u5_mult_79_CARRYB_5__21_,
         u5_mult_79_CARRYB_5__22_, u5_mult_79_CARRYB_6__0_,
         u5_mult_79_CARRYB_6__1_, u5_mult_79_CARRYB_6__2_,
         u5_mult_79_CARRYB_6__3_, u5_mult_79_CARRYB_6__4_,
         u5_mult_79_CARRYB_6__5_, u5_mult_79_CARRYB_6__6_,
         u5_mult_79_CARRYB_6__7_, u5_mult_79_CARRYB_6__8_,
         u5_mult_79_CARRYB_6__9_, u5_mult_79_CARRYB_6__10_,
         u5_mult_79_CARRYB_6__11_, u5_mult_79_CARRYB_6__12_,
         u5_mult_79_CARRYB_6__13_, u5_mult_79_CARRYB_6__14_,
         u5_mult_79_CARRYB_6__15_, u5_mult_79_CARRYB_6__16_,
         u5_mult_79_CARRYB_6__17_, u5_mult_79_CARRYB_6__18_,
         u5_mult_79_CARRYB_6__19_, u5_mult_79_CARRYB_6__20_,
         u5_mult_79_CARRYB_6__21_, u5_mult_79_CARRYB_6__22_,
         u5_mult_79_CARRYB_7__0_, u5_mult_79_CARRYB_7__1_,
         u5_mult_79_CARRYB_7__2_, u5_mult_79_CARRYB_7__3_,
         u5_mult_79_CARRYB_7__4_, u5_mult_79_CARRYB_7__5_,
         u5_mult_79_CARRYB_7__6_, u5_mult_79_CARRYB_7__7_,
         u5_mult_79_CARRYB_7__8_, u5_mult_79_CARRYB_7__9_,
         u5_mult_79_CARRYB_7__10_, u5_mult_79_CARRYB_7__11_,
         u5_mult_79_CARRYB_7__12_, u5_mult_79_CARRYB_7__13_,
         u5_mult_79_CARRYB_7__14_, u5_mult_79_CARRYB_7__15_,
         u5_mult_79_CARRYB_7__16_, u5_mult_79_CARRYB_7__17_,
         u5_mult_79_CARRYB_7__18_, u5_mult_79_CARRYB_7__19_,
         u5_mult_79_CARRYB_7__20_, u5_mult_79_CARRYB_7__21_,
         u5_mult_79_CARRYB_7__22_, u5_mult_79_CARRYB_8__0_,
         u5_mult_79_CARRYB_8__1_, u5_mult_79_CARRYB_8__2_,
         u5_mult_79_CARRYB_8__3_, u5_mult_79_CARRYB_8__4_,
         u5_mult_79_CARRYB_8__5_, u5_mult_79_CARRYB_8__6_,
         u5_mult_79_CARRYB_8__7_, u5_mult_79_CARRYB_8__8_,
         u5_mult_79_CARRYB_8__9_, u5_mult_79_CARRYB_8__10_,
         u5_mult_79_CARRYB_8__11_, u5_mult_79_CARRYB_8__12_,
         u5_mult_79_CARRYB_8__13_, u5_mult_79_CARRYB_8__14_,
         u5_mult_79_CARRYB_8__15_, u5_mult_79_CARRYB_8__16_,
         u5_mult_79_CARRYB_8__17_, u5_mult_79_CARRYB_8__18_,
         u5_mult_79_CARRYB_8__19_, u5_mult_79_CARRYB_8__20_,
         u5_mult_79_CARRYB_8__21_, u5_mult_79_CARRYB_8__22_,
         u5_mult_79_CARRYB_9__0_, u5_mult_79_CARRYB_9__1_,
         u5_mult_79_CARRYB_9__2_, u5_mult_79_CARRYB_9__3_,
         u5_mult_79_CARRYB_9__4_, u5_mult_79_CARRYB_9__5_,
         u5_mult_79_CARRYB_9__6_, u5_mult_79_CARRYB_9__7_,
         u5_mult_79_CARRYB_9__8_, u5_mult_79_CARRYB_9__9_,
         u5_mult_79_CARRYB_9__10_, u5_mult_79_CARRYB_9__11_,
         u5_mult_79_CARRYB_9__12_, u5_mult_79_CARRYB_9__13_,
         u5_mult_79_CARRYB_9__14_, u5_mult_79_CARRYB_9__15_,
         u5_mult_79_CARRYB_9__16_, u5_mult_79_CARRYB_9__17_,
         u5_mult_79_CARRYB_9__18_, u5_mult_79_CARRYB_9__19_,
         u5_mult_79_CARRYB_9__20_, u5_mult_79_CARRYB_9__21_,
         u5_mult_79_CARRYB_9__22_, u5_mult_79_CARRYB_10__0_,
         u5_mult_79_CARRYB_10__1_, u5_mult_79_CARRYB_10__2_,
         u5_mult_79_CARRYB_10__3_, u5_mult_79_CARRYB_10__4_,
         u5_mult_79_CARRYB_10__5_, u5_mult_79_CARRYB_10__6_,
         u5_mult_79_CARRYB_10__7_, u5_mult_79_CARRYB_10__8_,
         u5_mult_79_CARRYB_10__9_, u5_mult_79_CARRYB_10__10_,
         u5_mult_79_CARRYB_10__11_, u5_mult_79_CARRYB_10__12_,
         u5_mult_79_CARRYB_10__13_, u5_mult_79_CARRYB_10__14_,
         u5_mult_79_CARRYB_10__15_, u5_mult_79_CARRYB_10__16_,
         u5_mult_79_CARRYB_10__17_, u5_mult_79_CARRYB_10__18_,
         u5_mult_79_CARRYB_10__19_, u5_mult_79_CARRYB_10__20_,
         u5_mult_79_CARRYB_10__21_, u5_mult_79_CARRYB_10__22_,
         u5_mult_79_CARRYB_11__0_, u5_mult_79_CARRYB_11__1_,
         u5_mult_79_CARRYB_11__2_, u5_mult_79_CARRYB_11__3_,
         u5_mult_79_CARRYB_11__4_, u5_mult_79_CARRYB_11__5_,
         u5_mult_79_CARRYB_11__6_, u5_mult_79_CARRYB_11__7_,
         u5_mult_79_CARRYB_11__8_, u5_mult_79_CARRYB_11__9_,
         u5_mult_79_CARRYB_11__10_, u5_mult_79_CARRYB_11__11_,
         u5_mult_79_CARRYB_11__12_, u5_mult_79_CARRYB_11__13_,
         u5_mult_79_CARRYB_11__14_, u5_mult_79_CARRYB_11__15_,
         u5_mult_79_CARRYB_11__16_, u5_mult_79_CARRYB_11__17_,
         u5_mult_79_CARRYB_11__18_, u5_mult_79_CARRYB_11__19_,
         u5_mult_79_CARRYB_11__20_, u5_mult_79_CARRYB_11__21_,
         u5_mult_79_CARRYB_11__22_, u5_mult_79_CARRYB_12__0_,
         u5_mult_79_CARRYB_12__1_, u5_mult_79_CARRYB_12__2_,
         u5_mult_79_CARRYB_12__3_, u5_mult_79_CARRYB_12__4_,
         u5_mult_79_CARRYB_12__5_, u5_mult_79_CARRYB_12__6_,
         u5_mult_79_CARRYB_12__7_, u5_mult_79_CARRYB_12__8_,
         u5_mult_79_CARRYB_12__9_, u5_mult_79_CARRYB_12__10_,
         u5_mult_79_CARRYB_12__11_, u5_mult_79_CARRYB_12__12_,
         u5_mult_79_CARRYB_12__13_, u5_mult_79_CARRYB_12__14_,
         u5_mult_79_CARRYB_12__15_, u5_mult_79_CARRYB_12__16_,
         u5_mult_79_CARRYB_12__17_, u5_mult_79_CARRYB_12__18_,
         u5_mult_79_CARRYB_12__19_, u5_mult_79_CARRYB_12__20_,
         u5_mult_79_CARRYB_12__21_, u5_mult_79_CARRYB_12__22_,
         u5_mult_79_CARRYB_13__0_, u5_mult_79_CARRYB_13__1_,
         u5_mult_79_CARRYB_13__2_, u5_mult_79_CARRYB_13__3_,
         u5_mult_79_CARRYB_13__4_, u5_mult_79_CARRYB_13__5_,
         u5_mult_79_CARRYB_13__6_, u5_mult_79_CARRYB_13__7_,
         u5_mult_79_CARRYB_13__8_, u5_mult_79_CARRYB_13__9_,
         u5_mult_79_CARRYB_13__10_, u5_mult_79_CARRYB_13__11_,
         u5_mult_79_CARRYB_13__12_, u5_mult_79_CARRYB_13__13_,
         u5_mult_79_CARRYB_13__14_, u5_mult_79_CARRYB_13__15_,
         u5_mult_79_CARRYB_13__16_, u5_mult_79_CARRYB_13__17_,
         u5_mult_79_CARRYB_13__18_, u5_mult_79_CARRYB_13__19_,
         u5_mult_79_CARRYB_13__20_, u5_mult_79_CARRYB_13__21_,
         u5_mult_79_CARRYB_13__22_, u5_mult_79_CARRYB_14__0_,
         u5_mult_79_CARRYB_14__1_, u5_mult_79_CARRYB_14__2_,
         u5_mult_79_CARRYB_14__3_, u5_mult_79_CARRYB_14__4_,
         u5_mult_79_CARRYB_14__5_, u5_mult_79_CARRYB_14__6_,
         u5_mult_79_CARRYB_14__7_, u5_mult_79_CARRYB_14__8_,
         u5_mult_79_CARRYB_14__9_, u5_mult_79_CARRYB_14__10_,
         u5_mult_79_CARRYB_14__11_, u5_mult_79_CARRYB_14__12_,
         u5_mult_79_CARRYB_14__13_, u5_mult_79_CARRYB_14__14_,
         u5_mult_79_CARRYB_14__15_, u5_mult_79_CARRYB_14__16_,
         u5_mult_79_CARRYB_14__17_, u5_mult_79_CARRYB_14__18_,
         u5_mult_79_CARRYB_14__19_, u5_mult_79_CARRYB_14__20_,
         u5_mult_79_CARRYB_14__21_, u5_mult_79_CARRYB_14__22_,
         u5_mult_79_CARRYB_15__0_, u5_mult_79_CARRYB_15__1_,
         u5_mult_79_CARRYB_15__2_, u5_mult_79_CARRYB_15__3_,
         u5_mult_79_CARRYB_15__4_, u5_mult_79_CARRYB_15__5_,
         u5_mult_79_CARRYB_15__6_, u5_mult_79_CARRYB_15__7_,
         u5_mult_79_CARRYB_15__8_, u5_mult_79_CARRYB_15__9_,
         u5_mult_79_CARRYB_15__10_, u5_mult_79_CARRYB_15__11_,
         u5_mult_79_CARRYB_15__12_, u5_mult_79_CARRYB_15__13_,
         u5_mult_79_CARRYB_15__14_, u5_mult_79_CARRYB_15__15_,
         u5_mult_79_CARRYB_15__16_, u5_mult_79_CARRYB_15__17_,
         u5_mult_79_CARRYB_15__18_, u5_mult_79_CARRYB_15__19_,
         u5_mult_79_CARRYB_15__20_, u5_mult_79_CARRYB_15__21_,
         u5_mult_79_CARRYB_15__22_, u5_mult_79_CARRYB_16__0_,
         u5_mult_79_CARRYB_16__1_, u5_mult_79_CARRYB_16__2_,
         u5_mult_79_CARRYB_16__3_, u5_mult_79_CARRYB_16__4_,
         u5_mult_79_CARRYB_16__5_, u5_mult_79_CARRYB_16__6_,
         u5_mult_79_CARRYB_16__7_, u5_mult_79_CARRYB_16__8_,
         u5_mult_79_CARRYB_16__9_, u5_mult_79_CARRYB_16__10_,
         u5_mult_79_CARRYB_16__11_, u5_mult_79_CARRYB_16__12_,
         u5_mult_79_CARRYB_16__13_, u5_mult_79_CARRYB_16__14_,
         u5_mult_79_CARRYB_16__15_, u5_mult_79_CARRYB_16__16_,
         u5_mult_79_CARRYB_16__17_, u5_mult_79_CARRYB_16__18_,
         u5_mult_79_CARRYB_16__19_, u5_mult_79_CARRYB_16__20_,
         u5_mult_79_CARRYB_16__21_, u5_mult_79_CARRYB_16__22_,
         u5_mult_79_CARRYB_17__0_, u5_mult_79_CARRYB_17__1_,
         u5_mult_79_CARRYB_17__2_, u5_mult_79_CARRYB_17__3_,
         u5_mult_79_CARRYB_17__4_, u5_mult_79_CARRYB_17__5_,
         u5_mult_79_CARRYB_17__6_, u5_mult_79_CARRYB_17__7_,
         u5_mult_79_CARRYB_17__8_, u5_mult_79_CARRYB_17__9_,
         u5_mult_79_CARRYB_17__10_, u5_mult_79_CARRYB_17__11_,
         u5_mult_79_CARRYB_17__12_, u5_mult_79_CARRYB_17__13_,
         u5_mult_79_CARRYB_17__14_, u5_mult_79_CARRYB_17__15_,
         u5_mult_79_CARRYB_17__16_, u5_mult_79_CARRYB_17__17_,
         u5_mult_79_CARRYB_17__18_, u5_mult_79_CARRYB_17__19_,
         u5_mult_79_CARRYB_17__20_, u5_mult_79_CARRYB_17__21_,
         u5_mult_79_CARRYB_17__22_, u5_mult_79_CARRYB_18__0_,
         u5_mult_79_CARRYB_18__1_, u5_mult_79_CARRYB_18__2_,
         u5_mult_79_CARRYB_18__3_, u5_mult_79_CARRYB_18__4_,
         u5_mult_79_CARRYB_18__5_, u5_mult_79_CARRYB_18__6_,
         u5_mult_79_CARRYB_18__7_, u5_mult_79_CARRYB_18__8_,
         u5_mult_79_CARRYB_18__9_, u5_mult_79_CARRYB_18__10_,
         u5_mult_79_CARRYB_18__11_, u5_mult_79_CARRYB_18__12_,
         u5_mult_79_CARRYB_18__13_, u5_mult_79_CARRYB_18__14_,
         u5_mult_79_CARRYB_18__15_, u5_mult_79_CARRYB_18__16_,
         u5_mult_79_CARRYB_18__17_, u5_mult_79_CARRYB_18__18_,
         u5_mult_79_CARRYB_18__19_, u5_mult_79_CARRYB_18__20_,
         u5_mult_79_CARRYB_18__21_, u5_mult_79_CARRYB_18__22_,
         u5_mult_79_CARRYB_19__0_, u5_mult_79_CARRYB_19__1_,
         u5_mult_79_CARRYB_19__2_, u5_mult_79_CARRYB_19__3_,
         u5_mult_79_CARRYB_19__4_, u5_mult_79_CARRYB_19__5_,
         u5_mult_79_CARRYB_19__6_, u5_mult_79_CARRYB_19__7_,
         u5_mult_79_CARRYB_19__8_, u5_mult_79_CARRYB_19__9_,
         u5_mult_79_CARRYB_19__10_, u5_mult_79_CARRYB_19__11_,
         u5_mult_79_CARRYB_19__12_, u5_mult_79_CARRYB_19__13_,
         u5_mult_79_CARRYB_19__14_, u5_mult_79_CARRYB_19__15_,
         u5_mult_79_CARRYB_19__16_, u5_mult_79_CARRYB_19__17_,
         u5_mult_79_CARRYB_19__18_, u5_mult_79_CARRYB_19__19_,
         u5_mult_79_CARRYB_19__20_, u5_mult_79_CARRYB_19__21_,
         u5_mult_79_CARRYB_19__22_, u5_mult_79_CARRYB_20__0_,
         u5_mult_79_CARRYB_20__1_, u5_mult_79_CARRYB_20__2_,
         u5_mult_79_CARRYB_20__3_, u5_mult_79_CARRYB_20__4_,
         u5_mult_79_CARRYB_20__5_, u5_mult_79_CARRYB_20__6_,
         u5_mult_79_CARRYB_20__7_, u5_mult_79_CARRYB_20__8_,
         u5_mult_79_CARRYB_20__9_, u5_mult_79_CARRYB_20__10_,
         u5_mult_79_CARRYB_20__11_, u5_mult_79_CARRYB_20__12_,
         u5_mult_79_CARRYB_20__13_, u5_mult_79_CARRYB_20__14_,
         u5_mult_79_CARRYB_20__15_, u5_mult_79_CARRYB_20__16_,
         u5_mult_79_CARRYB_20__17_, u5_mult_79_CARRYB_20__18_,
         u5_mult_79_CARRYB_20__19_, u5_mult_79_CARRYB_20__20_,
         u5_mult_79_CARRYB_20__21_, u5_mult_79_CARRYB_20__22_,
         u5_mult_79_CARRYB_21__0_, u5_mult_79_CARRYB_21__1_,
         u5_mult_79_CARRYB_21__2_, u5_mult_79_CARRYB_21__3_,
         u5_mult_79_CARRYB_21__4_, u5_mult_79_CARRYB_21__5_,
         u5_mult_79_CARRYB_21__6_, u5_mult_79_CARRYB_21__7_,
         u5_mult_79_CARRYB_21__8_, u5_mult_79_CARRYB_21__9_,
         u5_mult_79_CARRYB_21__10_, u5_mult_79_CARRYB_21__11_,
         u5_mult_79_CARRYB_21__12_, u5_mult_79_CARRYB_21__13_,
         u5_mult_79_CARRYB_21__14_, u5_mult_79_CARRYB_21__15_,
         u5_mult_79_CARRYB_21__16_, u5_mult_79_CARRYB_21__17_,
         u5_mult_79_CARRYB_21__18_, u5_mult_79_CARRYB_21__19_,
         u5_mult_79_CARRYB_21__20_, u5_mult_79_CARRYB_21__21_,
         u5_mult_79_CARRYB_21__22_, u5_mult_79_CARRYB_22__0_,
         u5_mult_79_CARRYB_22__1_, u5_mult_79_CARRYB_22__2_,
         u5_mult_79_CARRYB_22__3_, u5_mult_79_CARRYB_22__4_,
         u5_mult_79_CARRYB_22__5_, u5_mult_79_CARRYB_22__6_,
         u5_mult_79_CARRYB_22__7_, u5_mult_79_CARRYB_22__8_,
         u5_mult_79_CARRYB_22__9_, u5_mult_79_CARRYB_22__10_,
         u5_mult_79_CARRYB_22__11_, u5_mult_79_CARRYB_22__12_,
         u5_mult_79_CARRYB_22__13_, u5_mult_79_CARRYB_22__14_,
         u5_mult_79_CARRYB_22__15_, u5_mult_79_CARRYB_22__16_,
         u5_mult_79_CARRYB_22__17_, u5_mult_79_CARRYB_22__18_,
         u5_mult_79_CARRYB_22__19_, u5_mult_79_CARRYB_22__20_,
         u5_mult_79_CARRYB_22__21_, u5_mult_79_CARRYB_22__22_,
         u5_mult_79_CARRYB_23__0_, u5_mult_79_CARRYB_23__1_,
         u5_mult_79_CARRYB_23__2_, u5_mult_79_CARRYB_23__3_,
         u5_mult_79_CARRYB_23__4_, u5_mult_79_CARRYB_23__5_,
         u5_mult_79_CARRYB_23__6_, u5_mult_79_CARRYB_23__7_,
         u5_mult_79_CARRYB_23__8_, u5_mult_79_CARRYB_23__9_,
         u5_mult_79_CARRYB_23__10_, u5_mult_79_CARRYB_23__11_,
         u5_mult_79_CARRYB_23__12_, u5_mult_79_CARRYB_23__13_,
         u5_mult_79_CARRYB_23__14_, u5_mult_79_CARRYB_23__15_,
         u5_mult_79_CARRYB_23__16_, u5_mult_79_CARRYB_23__17_,
         u5_mult_79_CARRYB_23__18_, u5_mult_79_CARRYB_23__19_,
         u5_mult_79_CARRYB_23__20_, u5_mult_79_CARRYB_23__21_,
         u5_mult_79_CARRYB_23__22_, u5_mult_79_ab_0__1_, u5_mult_79_ab_0__2_,
         u5_mult_79_ab_0__3_, u5_mult_79_ab_0__4_, u5_mult_79_ab_0__5_,
         u5_mult_79_ab_0__6_, u5_mult_79_ab_0__7_, u5_mult_79_ab_0__8_,
         u5_mult_79_ab_0__9_, u5_mult_79_ab_0__10_, u5_mult_79_ab_0__11_,
         u5_mult_79_ab_0__12_, u5_mult_79_ab_0__13_, u5_mult_79_ab_0__14_,
         u5_mult_79_ab_0__15_, u5_mult_79_ab_0__16_, u5_mult_79_ab_0__17_,
         u5_mult_79_ab_0__18_, u5_mult_79_ab_0__19_, u5_mult_79_ab_0__20_,
         u5_mult_79_ab_0__21_, u5_mult_79_ab_0__22_, u5_mult_79_ab_0__23_,
         u5_mult_79_ab_1__0_, u5_mult_79_ab_1__1_, u5_mult_79_ab_1__2_,
         u5_mult_79_ab_1__3_, u5_mult_79_ab_1__4_, u5_mult_79_ab_1__5_,
         u5_mult_79_ab_1__6_, u5_mult_79_ab_1__7_, u5_mult_79_ab_1__8_,
         u5_mult_79_ab_1__9_, u5_mult_79_ab_1__10_, u5_mult_79_ab_1__11_,
         u5_mult_79_ab_1__12_, u5_mult_79_ab_1__13_, u5_mult_79_ab_1__14_,
         u5_mult_79_ab_1__15_, u5_mult_79_ab_1__16_, u5_mult_79_ab_1__17_,
         u5_mult_79_ab_1__18_, u5_mult_79_ab_1__19_, u5_mult_79_ab_1__20_,
         u5_mult_79_ab_1__21_, u5_mult_79_ab_1__22_, u5_mult_79_ab_1__23_,
         u5_mult_79_ab_2__0_, u5_mult_79_ab_2__1_, u5_mult_79_ab_2__2_,
         u5_mult_79_ab_2__3_, u5_mult_79_ab_2__4_, u5_mult_79_ab_2__5_,
         u5_mult_79_ab_2__6_, u5_mult_79_ab_2__7_, u5_mult_79_ab_2__8_,
         u5_mult_79_ab_2__9_, u5_mult_79_ab_2__10_, u5_mult_79_ab_2__11_,
         u5_mult_79_ab_2__12_, u5_mult_79_ab_2__13_, u5_mult_79_ab_2__14_,
         u5_mult_79_ab_2__15_, u5_mult_79_ab_2__16_, u5_mult_79_ab_2__17_,
         u5_mult_79_ab_2__18_, u5_mult_79_ab_2__19_, u5_mult_79_ab_2__20_,
         u5_mult_79_ab_2__21_, u5_mult_79_ab_2__22_, u5_mult_79_ab_2__23_,
         u5_mult_79_ab_3__0_, u5_mult_79_ab_3__1_, u5_mult_79_ab_3__2_,
         u5_mult_79_ab_3__3_, u5_mult_79_ab_3__4_, u5_mult_79_ab_3__5_,
         u5_mult_79_ab_3__6_, u5_mult_79_ab_3__7_, u5_mult_79_ab_3__8_,
         u5_mult_79_ab_3__9_, u5_mult_79_ab_3__10_, u5_mult_79_ab_3__11_,
         u5_mult_79_ab_3__12_, u5_mult_79_ab_3__13_, u5_mult_79_ab_3__14_,
         u5_mult_79_ab_3__15_, u5_mult_79_ab_3__16_, u5_mult_79_ab_3__17_,
         u5_mult_79_ab_3__18_, u5_mult_79_ab_3__19_, u5_mult_79_ab_3__20_,
         u5_mult_79_ab_3__21_, u5_mult_79_ab_3__22_, u5_mult_79_ab_3__23_,
         u5_mult_79_ab_4__0_, u5_mult_79_ab_4__1_, u5_mult_79_ab_4__2_,
         u5_mult_79_ab_4__3_, u5_mult_79_ab_4__4_, u5_mult_79_ab_4__5_,
         u5_mult_79_ab_4__6_, u5_mult_79_ab_4__7_, u5_mult_79_ab_4__8_,
         u5_mult_79_ab_4__9_, u5_mult_79_ab_4__10_, u5_mult_79_ab_4__11_,
         u5_mult_79_ab_4__12_, u5_mult_79_ab_4__13_, u5_mult_79_ab_4__14_,
         u5_mult_79_ab_4__15_, u5_mult_79_ab_4__16_, u5_mult_79_ab_4__17_,
         u5_mult_79_ab_4__18_, u5_mult_79_ab_4__19_, u5_mult_79_ab_4__20_,
         u5_mult_79_ab_4__21_, u5_mult_79_ab_4__22_, u5_mult_79_ab_4__23_,
         u5_mult_79_ab_5__0_, u5_mult_79_ab_5__1_, u5_mult_79_ab_5__2_,
         u5_mult_79_ab_5__3_, u5_mult_79_ab_5__4_, u5_mult_79_ab_5__5_,
         u5_mult_79_ab_5__6_, u5_mult_79_ab_5__7_, u5_mult_79_ab_5__8_,
         u5_mult_79_ab_5__9_, u5_mult_79_ab_5__10_, u5_mult_79_ab_5__11_,
         u5_mult_79_ab_5__12_, u5_mult_79_ab_5__13_, u5_mult_79_ab_5__14_,
         u5_mult_79_ab_5__15_, u5_mult_79_ab_5__16_, u5_mult_79_ab_5__17_,
         u5_mult_79_ab_5__18_, u5_mult_79_ab_5__19_, u5_mult_79_ab_5__20_,
         u5_mult_79_ab_5__21_, u5_mult_79_ab_5__22_, u5_mult_79_ab_5__23_,
         u5_mult_79_ab_6__0_, u5_mult_79_ab_6__1_, u5_mult_79_ab_6__2_,
         u5_mult_79_ab_6__3_, u5_mult_79_ab_6__4_, u5_mult_79_ab_6__5_,
         u5_mult_79_ab_6__6_, u5_mult_79_ab_6__7_, u5_mult_79_ab_6__8_,
         u5_mult_79_ab_6__9_, u5_mult_79_ab_6__10_, u5_mult_79_ab_6__11_,
         u5_mult_79_ab_6__12_, u5_mult_79_ab_6__13_, u5_mult_79_ab_6__14_,
         u5_mult_79_ab_6__15_, u5_mult_79_ab_6__16_, u5_mult_79_ab_6__17_,
         u5_mult_79_ab_6__18_, u5_mult_79_ab_6__19_, u5_mult_79_ab_6__20_,
         u5_mult_79_ab_6__21_, u5_mult_79_ab_6__22_, u5_mult_79_ab_6__23_,
         u5_mult_79_ab_7__0_, u5_mult_79_ab_7__1_, u5_mult_79_ab_7__2_,
         u5_mult_79_ab_7__3_, u5_mult_79_ab_7__4_, u5_mult_79_ab_7__5_,
         u5_mult_79_ab_7__6_, u5_mult_79_ab_7__7_, u5_mult_79_ab_7__8_,
         u5_mult_79_ab_7__9_, u5_mult_79_ab_7__10_, u5_mult_79_ab_7__11_,
         u5_mult_79_ab_7__12_, u5_mult_79_ab_7__13_, u5_mult_79_ab_7__14_,
         u5_mult_79_ab_7__15_, u5_mult_79_ab_7__16_, u5_mult_79_ab_7__17_,
         u5_mult_79_ab_7__18_, u5_mult_79_ab_7__19_, u5_mult_79_ab_7__20_,
         u5_mult_79_ab_7__21_, u5_mult_79_ab_7__22_, u5_mult_79_ab_7__23_,
         u5_mult_79_ab_8__0_, u5_mult_79_ab_8__1_, u5_mult_79_ab_8__2_,
         u5_mult_79_ab_8__3_, u5_mult_79_ab_8__4_, u5_mult_79_ab_8__5_,
         u5_mult_79_ab_8__6_, u5_mult_79_ab_8__7_, u5_mult_79_ab_8__8_,
         u5_mult_79_ab_8__9_, u5_mult_79_ab_8__10_, u5_mult_79_ab_8__11_,
         u5_mult_79_ab_8__12_, u5_mult_79_ab_8__13_, u5_mult_79_ab_8__14_,
         u5_mult_79_ab_8__15_, u5_mult_79_ab_8__16_, u5_mult_79_ab_8__17_,
         u5_mult_79_ab_8__18_, u5_mult_79_ab_8__19_, u5_mult_79_ab_8__20_,
         u5_mult_79_ab_8__21_, u5_mult_79_ab_8__22_, u5_mult_79_ab_8__23_,
         u5_mult_79_ab_9__0_, u5_mult_79_ab_9__1_, u5_mult_79_ab_9__2_,
         u5_mult_79_ab_9__3_, u5_mult_79_ab_9__4_, u5_mult_79_ab_9__5_,
         u5_mult_79_ab_9__6_, u5_mult_79_ab_9__7_, u5_mult_79_ab_9__8_,
         u5_mult_79_ab_9__9_, u5_mult_79_ab_9__10_, u5_mult_79_ab_9__11_,
         u5_mult_79_ab_9__12_, u5_mult_79_ab_9__13_, u5_mult_79_ab_9__14_,
         u5_mult_79_ab_9__15_, u5_mult_79_ab_9__16_, u5_mult_79_ab_9__17_,
         u5_mult_79_ab_9__18_, u5_mult_79_ab_9__19_, u5_mult_79_ab_9__20_,
         u5_mult_79_ab_9__21_, u5_mult_79_ab_9__22_, u5_mult_79_ab_9__23_,
         u5_mult_79_ab_10__0_, u5_mult_79_ab_10__1_, u5_mult_79_ab_10__2_,
         u5_mult_79_ab_10__3_, u5_mult_79_ab_10__4_, u5_mult_79_ab_10__5_,
         u5_mult_79_ab_10__6_, u5_mult_79_ab_10__7_, u5_mult_79_ab_10__8_,
         u5_mult_79_ab_10__9_, u5_mult_79_ab_10__10_, u5_mult_79_ab_10__11_,
         u5_mult_79_ab_10__12_, u5_mult_79_ab_10__13_, u5_mult_79_ab_10__14_,
         u5_mult_79_ab_10__15_, u5_mult_79_ab_10__16_, u5_mult_79_ab_10__17_,
         u5_mult_79_ab_10__18_, u5_mult_79_ab_10__19_, u5_mult_79_ab_10__20_,
         u5_mult_79_ab_10__21_, u5_mult_79_ab_10__22_, u5_mult_79_ab_10__23_,
         u5_mult_79_ab_11__0_, u5_mult_79_ab_11__1_, u5_mult_79_ab_11__2_,
         u5_mult_79_ab_11__3_, u5_mult_79_ab_11__4_, u5_mult_79_ab_11__5_,
         u5_mult_79_ab_11__6_, u5_mult_79_ab_11__7_, u5_mult_79_ab_11__8_,
         u5_mult_79_ab_11__9_, u5_mult_79_ab_11__10_, u5_mult_79_ab_11__11_,
         u5_mult_79_ab_11__12_, u5_mult_79_ab_11__13_, u5_mult_79_ab_11__14_,
         u5_mult_79_ab_11__15_, u5_mult_79_ab_11__16_, u5_mult_79_ab_11__17_,
         u5_mult_79_ab_11__18_, u5_mult_79_ab_11__19_, u5_mult_79_ab_11__20_,
         u5_mult_79_ab_11__21_, u5_mult_79_ab_11__22_, u5_mult_79_ab_11__23_,
         u5_mult_79_ab_12__0_, u5_mult_79_ab_12__1_, u5_mult_79_ab_12__2_,
         u5_mult_79_ab_12__3_, u5_mult_79_ab_12__4_, u5_mult_79_ab_12__5_,
         u5_mult_79_ab_12__6_, u5_mult_79_ab_12__7_, u5_mult_79_ab_12__8_,
         u5_mult_79_ab_12__9_, u5_mult_79_ab_12__10_, u5_mult_79_ab_12__11_,
         u5_mult_79_ab_12__12_, u5_mult_79_ab_12__13_, u5_mult_79_ab_12__14_,
         u5_mult_79_ab_12__15_, u5_mult_79_ab_12__16_, u5_mult_79_ab_12__17_,
         u5_mult_79_ab_12__18_, u5_mult_79_ab_12__19_, u5_mult_79_ab_12__20_,
         u5_mult_79_ab_12__21_, u5_mult_79_ab_12__22_, u5_mult_79_ab_12__23_,
         u5_mult_79_ab_13__0_, u5_mult_79_ab_13__1_, u5_mult_79_ab_13__2_,
         u5_mult_79_ab_13__3_, u5_mult_79_ab_13__4_, u5_mult_79_ab_13__5_,
         u5_mult_79_ab_13__6_, u5_mult_79_ab_13__7_, u5_mult_79_ab_13__8_,
         u5_mult_79_ab_13__9_, u5_mult_79_ab_13__10_, u5_mult_79_ab_13__11_,
         u5_mult_79_ab_13__12_, u5_mult_79_ab_13__13_, u5_mult_79_ab_13__14_,
         u5_mult_79_ab_13__15_, u5_mult_79_ab_13__16_, u5_mult_79_ab_13__17_,
         u5_mult_79_ab_13__18_, u5_mult_79_ab_13__19_, u5_mult_79_ab_13__20_,
         u5_mult_79_ab_13__21_, u5_mult_79_ab_13__22_, u5_mult_79_ab_13__23_,
         u5_mult_79_ab_14__0_, u5_mult_79_ab_14__1_, u5_mult_79_ab_14__2_,
         u5_mult_79_ab_14__3_, u5_mult_79_ab_14__4_, u5_mult_79_ab_14__5_,
         u5_mult_79_ab_14__6_, u5_mult_79_ab_14__7_, u5_mult_79_ab_14__8_,
         u5_mult_79_ab_14__9_, u5_mult_79_ab_14__10_, u5_mult_79_ab_14__11_,
         u5_mult_79_ab_14__12_, u5_mult_79_ab_14__13_, u5_mult_79_ab_14__14_,
         u5_mult_79_ab_14__15_, u5_mult_79_ab_14__16_, u5_mult_79_ab_14__17_,
         u5_mult_79_ab_14__18_, u5_mult_79_ab_14__19_, u5_mult_79_ab_14__20_,
         u5_mult_79_ab_14__21_, u5_mult_79_ab_14__22_, u5_mult_79_ab_14__23_,
         u5_mult_79_ab_15__0_, u5_mult_79_ab_15__1_, u5_mult_79_ab_15__2_,
         u5_mult_79_ab_15__3_, u5_mult_79_ab_15__4_, u5_mult_79_ab_15__5_,
         u5_mult_79_ab_15__6_, u5_mult_79_ab_15__7_, u5_mult_79_ab_15__8_,
         u5_mult_79_ab_15__9_, u5_mult_79_ab_15__10_, u5_mult_79_ab_15__11_,
         u5_mult_79_ab_15__12_, u5_mult_79_ab_15__13_, u5_mult_79_ab_15__14_,
         u5_mult_79_ab_15__15_, u5_mult_79_ab_15__16_, u5_mult_79_ab_15__17_,
         u5_mult_79_ab_15__18_, u5_mult_79_ab_15__19_, u5_mult_79_ab_15__20_,
         u5_mult_79_ab_15__21_, u5_mult_79_ab_15__22_, u5_mult_79_ab_15__23_,
         u5_mult_79_ab_16__0_, u5_mult_79_ab_16__1_, u5_mult_79_ab_16__2_,
         u5_mult_79_ab_16__3_, u5_mult_79_ab_16__4_, u5_mult_79_ab_16__5_,
         u5_mult_79_ab_16__6_, u5_mult_79_ab_16__7_, u5_mult_79_ab_16__8_,
         u5_mult_79_ab_16__9_, u5_mult_79_ab_16__10_, u5_mult_79_ab_16__11_,
         u5_mult_79_ab_16__12_, u5_mult_79_ab_16__13_, u5_mult_79_ab_16__14_,
         u5_mult_79_ab_16__15_, u5_mult_79_ab_16__16_, u5_mult_79_ab_16__17_,
         u5_mult_79_ab_16__18_, u5_mult_79_ab_16__19_, u5_mult_79_ab_16__20_,
         u5_mult_79_ab_16__21_, u5_mult_79_ab_16__22_, u5_mult_79_ab_16__23_,
         u5_mult_79_ab_17__0_, u5_mult_79_ab_17__1_, u5_mult_79_ab_17__2_,
         u5_mult_79_ab_17__3_, u5_mult_79_ab_17__4_, u5_mult_79_ab_17__5_,
         u5_mult_79_ab_17__6_, u5_mult_79_ab_17__7_, u5_mult_79_ab_17__8_,
         u5_mult_79_ab_17__9_, u5_mult_79_ab_17__10_, u5_mult_79_ab_17__11_,
         u5_mult_79_ab_17__12_, u5_mult_79_ab_17__13_, u5_mult_79_ab_17__14_,
         u5_mult_79_ab_17__15_, u5_mult_79_ab_17__16_, u5_mult_79_ab_17__17_,
         u5_mult_79_ab_17__18_, u5_mult_79_ab_17__19_, u5_mult_79_ab_17__20_,
         u5_mult_79_ab_17__21_, u5_mult_79_ab_17__22_, u5_mult_79_ab_17__23_,
         u5_mult_79_ab_18__0_, u5_mult_79_ab_18__1_, u5_mult_79_ab_18__2_,
         u5_mult_79_ab_18__3_, u5_mult_79_ab_18__4_, u5_mult_79_ab_18__5_,
         u5_mult_79_ab_18__6_, u5_mult_79_ab_18__7_, u5_mult_79_ab_18__8_,
         u5_mult_79_ab_18__9_, u5_mult_79_ab_18__10_, u5_mult_79_ab_18__11_,
         u5_mult_79_ab_18__12_, u5_mult_79_ab_18__13_, u5_mult_79_ab_18__14_,
         u5_mult_79_ab_18__15_, u5_mult_79_ab_18__16_, u5_mult_79_ab_18__17_,
         u5_mult_79_ab_18__18_, u5_mult_79_ab_18__19_, u5_mult_79_ab_18__20_,
         u5_mult_79_ab_18__21_, u5_mult_79_ab_18__22_, u5_mult_79_ab_18__23_,
         u5_mult_79_ab_19__0_, u5_mult_79_ab_19__1_, u5_mult_79_ab_19__2_,
         u5_mult_79_ab_19__3_, u5_mult_79_ab_19__4_, u5_mult_79_ab_19__5_,
         u5_mult_79_ab_19__6_, u5_mult_79_ab_19__7_, u5_mult_79_ab_19__8_,
         u5_mult_79_ab_19__9_, u5_mult_79_ab_19__10_, u5_mult_79_ab_19__11_,
         u5_mult_79_ab_19__12_, u5_mult_79_ab_19__13_, u5_mult_79_ab_19__14_,
         u5_mult_79_ab_19__15_, u5_mult_79_ab_19__16_, u5_mult_79_ab_19__17_,
         u5_mult_79_ab_19__18_, u5_mult_79_ab_19__19_, u5_mult_79_ab_19__20_,
         u5_mult_79_ab_19__21_, u5_mult_79_ab_19__22_, u5_mult_79_ab_19__23_,
         u5_mult_79_ab_20__0_, u5_mult_79_ab_20__1_, u5_mult_79_ab_20__2_,
         u5_mult_79_ab_20__3_, u5_mult_79_ab_20__4_, u5_mult_79_ab_20__5_,
         u5_mult_79_ab_20__6_, u5_mult_79_ab_20__7_, u5_mult_79_ab_20__8_,
         u5_mult_79_ab_20__9_, u5_mult_79_ab_20__10_, u5_mult_79_ab_20__11_,
         u5_mult_79_ab_20__12_, u5_mult_79_ab_20__13_, u5_mult_79_ab_20__14_,
         u5_mult_79_ab_20__15_, u5_mult_79_ab_20__16_, u5_mult_79_ab_20__17_,
         u5_mult_79_ab_20__18_, u5_mult_79_ab_20__19_, u5_mult_79_ab_20__20_,
         u5_mult_79_ab_20__21_, u5_mult_79_ab_20__22_, u5_mult_79_ab_20__23_,
         u5_mult_79_ab_21__0_, u5_mult_79_ab_21__1_, u5_mult_79_ab_21__2_,
         u5_mult_79_ab_21__3_, u5_mult_79_ab_21__4_, u5_mult_79_ab_21__5_,
         u5_mult_79_ab_21__6_, u5_mult_79_ab_21__7_, u5_mult_79_ab_21__8_,
         u5_mult_79_ab_21__9_, u5_mult_79_ab_21__10_, u5_mult_79_ab_21__11_,
         u5_mult_79_ab_21__12_, u5_mult_79_ab_21__13_, u5_mult_79_ab_21__14_,
         u5_mult_79_ab_21__15_, u5_mult_79_ab_21__16_, u5_mult_79_ab_21__17_,
         u5_mult_79_ab_21__18_, u5_mult_79_ab_21__19_, u5_mult_79_ab_21__20_,
         u5_mult_79_ab_21__21_, u5_mult_79_ab_21__22_, u5_mult_79_ab_21__23_,
         u5_mult_79_ab_22__0_, u5_mult_79_ab_22__1_, u5_mult_79_ab_22__2_,
         u5_mult_79_ab_22__3_, u5_mult_79_ab_22__4_, u5_mult_79_ab_22__5_,
         u5_mult_79_ab_22__6_, u5_mult_79_ab_22__7_, u5_mult_79_ab_22__8_,
         u5_mult_79_ab_22__9_, u5_mult_79_ab_22__10_, u5_mult_79_ab_22__11_,
         u5_mult_79_ab_22__12_, u5_mult_79_ab_22__13_, u5_mult_79_ab_22__14_,
         u5_mult_79_ab_22__15_, u5_mult_79_ab_22__16_, u5_mult_79_ab_22__17_,
         u5_mult_79_ab_22__18_, u5_mult_79_ab_22__19_, u5_mult_79_ab_22__20_,
         u5_mult_79_ab_22__21_, u5_mult_79_ab_22__22_, u5_mult_79_ab_22__23_,
         u5_mult_79_ab_23__0_, u5_mult_79_ab_23__1_, u5_mult_79_ab_23__2_,
         u5_mult_79_ab_23__3_, u5_mult_79_ab_23__4_, u5_mult_79_ab_23__5_,
         u5_mult_79_ab_23__6_, u5_mult_79_ab_23__7_, u5_mult_79_ab_23__8_,
         u5_mult_79_ab_23__9_, u5_mult_79_ab_23__10_, u5_mult_79_ab_23__11_,
         u5_mult_79_ab_23__12_, u5_mult_79_ab_23__13_, u5_mult_79_ab_23__14_,
         u5_mult_79_ab_23__15_, u5_mult_79_ab_23__16_, u5_mult_79_ab_23__17_,
         u5_mult_79_ab_23__18_, u5_mult_79_ab_23__19_, u5_mult_79_ab_23__20_,
         u5_mult_79_ab_23__21_, u5_mult_79_ab_23__22_, u5_mult_79_ab_23__23_,
         u5_mult_79_FS_1_n110, u5_mult_79_FS_1_n109, u5_mult_79_FS_1_n108,
         u5_mult_79_FS_1_n107, u5_mult_79_FS_1_n106, u5_mult_79_FS_1_n105,
         u5_mult_79_FS_1_n104, u5_mult_79_FS_1_n103, u5_mult_79_FS_1_n102,
         u5_mult_79_FS_1_n101, u5_mult_79_FS_1_n100, u5_mult_79_FS_1_n99,
         u5_mult_79_FS_1_n98, u5_mult_79_FS_1_n97, u5_mult_79_FS_1_n96,
         u5_mult_79_FS_1_n95, u5_mult_79_FS_1_n94, u5_mult_79_FS_1_n93,
         u5_mult_79_FS_1_n92, u5_mult_79_FS_1_n91, u5_mult_79_FS_1_n90,
         u5_mult_79_FS_1_n89, u5_mult_79_FS_1_n88, u5_mult_79_FS_1_n87,
         u5_mult_79_FS_1_n86, u5_mult_79_FS_1_n85, u5_mult_79_FS_1_n84,
         u5_mult_79_FS_1_n83, u5_mult_79_FS_1_n82, u5_mult_79_FS_1_n81,
         u5_mult_79_FS_1_n80, u5_mult_79_FS_1_n79, u5_mult_79_FS_1_n78,
         u5_mult_79_FS_1_n77, u5_mult_79_FS_1_n76, u5_mult_79_FS_1_n75,
         u5_mult_79_FS_1_n74, u5_mult_79_FS_1_n73, u5_mult_79_FS_1_n72,
         u5_mult_79_FS_1_n71, u5_mult_79_FS_1_n70, u5_mult_79_FS_1_n69,
         u5_mult_79_FS_1_n68, u5_mult_79_FS_1_n67, u5_mult_79_FS_1_n66,
         u5_mult_79_FS_1_n65, u5_mult_79_FS_1_n64, u5_mult_79_FS_1_n63,
         u5_mult_79_FS_1_n62, u5_mult_79_FS_1_n61, u5_mult_79_FS_1_n60,
         u5_mult_79_FS_1_n59, u5_mult_79_FS_1_n58, u5_mult_79_FS_1_n57,
         u5_mult_79_FS_1_n56, u5_mult_79_FS_1_n55, u5_mult_79_FS_1_n54,
         u5_mult_79_FS_1_n53, u5_mult_79_FS_1_n52, u5_mult_79_FS_1_n51,
         u5_mult_79_FS_1_n50, u5_mult_79_FS_1_n49, u5_mult_79_FS_1_n48,
         u5_mult_79_FS_1_n47, u5_mult_79_FS_1_n46, u5_mult_79_FS_1_n45,
         u5_mult_79_FS_1_n44, u5_mult_79_FS_1_n43, u5_mult_79_FS_1_n42,
         u5_mult_79_FS_1_n41, u5_mult_79_FS_1_n40, u5_mult_79_FS_1_n39,
         u5_mult_79_FS_1_n38, u5_mult_79_FS_1_n37, u5_mult_79_FS_1_n36,
         u5_mult_79_FS_1_n35, u5_mult_79_FS_1_n34, u5_mult_79_FS_1_n33,
         u5_mult_79_FS_1_n32, u5_mult_79_FS_1_n31, u5_mult_79_FS_1_n30,
         u5_mult_79_FS_1_n29, u5_mult_79_FS_1_n28, u5_mult_79_FS_1_n27,
         u5_mult_79_FS_1_n26, u5_mult_79_FS_1_n25, u5_mult_79_FS_1_n24,
         u5_mult_79_FS_1_n23, u5_mult_79_FS_1_n22, u5_mult_79_FS_1_n21,
         u5_mult_79_FS_1_n20, u5_mult_79_FS_1_n19, u5_mult_79_FS_1_n18,
         u5_mult_79_FS_1_n17, u5_mult_79_FS_1_n16, u5_mult_79_FS_1_n15,
         u5_mult_79_FS_1_n14, u5_mult_79_FS_1_n13, u5_mult_79_FS_1_n12,
         u5_mult_79_FS_1_n11, u5_mult_79_FS_1_n10, u5_mult_79_FS_1_n9,
         u5_mult_79_FS_1_n8, u5_mult_79_FS_1_n7, u5_mult_79_FS_1_n6,
         u5_mult_79_FS_1_n5, u5_mult_79_FS_1_n4, u5_mult_79_FS_1_n3,
         u5_mult_79_FS_1_n1;
  wire   [31:23] opa_r;
  wire   [31:23] opb_r;
  wire   [1:0] rmode_r1;
  wire   [1:0] rmode_r2;
  wire   [1:0] rmode_r3;
  wire   [2:0] fpu_op_r1;
  wire   [2:0] fpu_op_r2;
  wire   [1:0] fpu_op_r3;
  wire   [26:0] fracta;
  wire   [26:0] fractb;
  wire   [7:0] exp_fasu;
  wire   [22:0] fracta_mul;
  wire   [7:0] exp_mul;
  wire   [1:0] exp_ovf;
  wire   [2:0] underflow_fmul_d;
  wire   [1:0] exp_ovf_r;
  wire   [27:0] fract_out_q;
  wire   [47:0] prod;
  wire   [49:0] quo;
  wire   [49:0] remainder;
  wire   [4:0] div_opa_ldz_r1;
  wire   [4:0] div_opa_ldz_r2;
  wire   [30:1] opa_r1;
  wire   [47:0] fract_i2f;
  wire   [47:21] fract_denorm;
  wire   [2:0] underflow_fmul_r;
  wire   [26:0] u1_fractb_s;
  wire   [26:0] u1_fracta_s;
  wire   [7:0] u1_exp_diff2;
  wire   [7:0] u1_exp_small;
  wire   [2:0] u2_underflow_d;
  wire   [47:0] u5_prod1;
  wire   [49:0] u6_remainder;
  wire   [49:0] u6_quo1;
  wire   [7:0] u4_div_exp3;
  wire   [56:49] u4_exp_f2i_1;
  wire   [7:0] u4_exp_fix_divb;
  wire   [7:0] u4_exp_fix_diva;
  wire   [7:1] u4_exp_out1_mi1;
  wire   [7:0] u4_exp_out_mi1;
  wire   [5:2] u4_fi_ldz_mi22;
  wire   [5:0] u4_shift_left;
  wire   [7:0] u4_shift_right;
  wire   [7:0] u4_div_shft4;
  wire   [7:2] u4_div_shft2;
  wire   [7:0] u4_div_scht1a;
  wire   [5:3] u4_sub_460_carry;
  wire   [5:2] u4_sub_478_carry;
  wire   [5:1] u4_add_486_carry;
  wire   [7:3] u4_add_407_carry;
  wire   [7:1] u4_sub_406_carry;
  wire   [5:5] u4_sub_488_carry;
  wire   [7:1] u4_sub_470_carry;
  wire   [7:1] u4_sub_469_carry;
  wire   [7:2] u4_add_461_carry;
  wire   [5:4] u4_sll_479_SHMAG;
  wire   [7:1] u4_sub_493_carry;
  wire   [7:2] u4_add_463_carry;
  wire   [8:2] u4_add_491_carry;
  wire   [22:2] u4_add_393_carry;
  wire   [27:1] u3_sub_60_carry;
  wire   [26:2] u3_add_60_carry;
  wire   [7:2] u2_add_114_carry;
  wire   [7:2] u2_add_112_carry;
  wire   [7:2] u2_add_109_carry;
  wire   [8:1] u2_sub_109_carry;
  wire   [7:1] sub_1_root_u1_sub_128_aco_carry;
  wire   [7:2] add_0_root_sub_0_root_u4_add_494_carry;

  OR2_X2 u4_C5085 ( .A1(u4_N1732), .A2(u4_exp_out_0_), .ZN(u4_N1733) );
  OR2_X2 u4_C5086 ( .A1(u4_N1731), .A2(u4_exp_out_1_), .ZN(u4_N1732) );
  OR2_X2 u4_C5087 ( .A1(u4_N1730), .A2(u4_exp_out_2_), .ZN(u4_N1731) );
  OR2_X2 u4_C5088 ( .A1(u4_N1729), .A2(u4_exp_out_3_), .ZN(u4_N1730) );
  OR2_X2 u4_C5089 ( .A1(u4_N1728), .A2(u4_exp_out_4_), .ZN(u4_N1729) );
  OR2_X2 u4_C5090 ( .A1(u4_N1727), .A2(u4_exp_out_5_), .ZN(u4_N1728) );
  OR2_X2 u4_C5091 ( .A1(u4_N1976), .A2(u4_exp_out_6_), .ZN(u4_N1727) );
  OR2_X2 u4_C5360 ( .A1(u4_shift_right[7]), .A2(u4_shift_right[6]), .ZN(
        u4_N1356) );
  OR2_X2 u4_C5564 ( .A1(u4_N1640), .A2(u4_N1976), .ZN(u4_N1977) );
  MUX2_X2 U3 ( .A(prod[47]), .B(fract_div_47_), .S(fpu_op_r3[0]), .Z(n202) );
  MUX2_X2 U4 ( .A(fract_out_q[27]), .B(n202), .S(fpu_op_r3[1]), .Z(n203) );
  AND2_X2 U5 ( .A1(fract_i2f[47]), .A2(n2532), .ZN(n204) );
  MUX2_X2 U6 ( .A(n203), .B(n204), .S(n2690), .Z(fract_denorm[47]) );
  OAI221_X2 U8 ( .B1(n1355), .B2(n3440), .C1(n1356), .C2(n1357), .A(n1358), 
        .ZN(u4_exp_out_0_) );
  NAND2_X2 U11 ( .A1(u4_div_exp3[0]), .A2(n1363), .ZN(n1365) );
  OAI211_X2 U14 ( .C1(n3352), .C2(n2649), .A(n1369), .B(n1370), .ZN(
        u4_exp_out_1_) );
  AOI221_X2 U15 ( .B1(u4_N1472), .B2(n1359), .C1(n1371), .C2(n3441), .A(n1372), 
        .ZN(n1370) );
  NOR2_X4 U16 ( .A1(n2680), .A2(n1368), .ZN(n1371) );
  AOI22_X2 U17 ( .A1(u4_exp_f2i_1[50]), .A2(n3489), .B1(n1373), .B2(
        u4_exp_out1_1_), .ZN(n1369) );
  OAI221_X2 U18 ( .B1(n1374), .B2(n1357), .C1(n3351), .C2(n2649), .A(n1375), 
        .ZN(u4_exp_out_2_) );
  AOI221_X2 U19 ( .B1(u4_exp_f2i_1[51]), .B2(n3489), .C1(u4_N1473), .C2(n1359), 
        .A(n1372), .ZN(n1375) );
  OAI221_X2 U20 ( .B1(n1376), .B2(n1357), .C1(n3350), .C2(n2649), .A(n1377), 
        .ZN(u4_exp_out_3_) );
  AOI221_X2 U21 ( .B1(u4_exp_f2i_1[52]), .B2(n3489), .C1(u4_N1474), .C2(n1359), 
        .A(n1372), .ZN(n1377) );
  OAI221_X2 U22 ( .B1(n1378), .B2(n1357), .C1(n3349), .C2(n2649), .A(n1379), 
        .ZN(u4_exp_out_4_) );
  AOI221_X2 U23 ( .B1(u4_exp_f2i_1[53]), .B2(n3489), .C1(u4_N1475), .C2(n1359), 
        .A(n1372), .ZN(n1379) );
  OAI221_X2 U24 ( .B1(n1380), .B2(n1357), .C1(n3348), .C2(n2649), .A(n1381), 
        .ZN(u4_exp_out_5_) );
  AOI22_X2 U25 ( .A1(u4_N1476), .A2(n1359), .B1(u4_exp_f2i_1[54]), .B2(n3489), 
        .ZN(n1381) );
  OAI221_X2 U26 ( .B1(n1382), .B2(n1357), .C1(n3347), .C2(n2649), .A(n1383), 
        .ZN(u4_exp_out_6_) );
  AOI22_X2 U27 ( .A1(u4_N1477), .A2(n1359), .B1(u4_exp_f2i_1[55]), .B2(n3489), 
        .ZN(n1383) );
  OAI221_X2 U28 ( .B1(n1384), .B2(n1357), .C1(n3346), .C2(n2649), .A(n1385), 
        .ZN(u4_N1976) );
  AOI221_X2 U29 ( .B1(u4_exp_f2i_1[56]), .B2(n3489), .C1(u4_N1478), .C2(n1359), 
        .A(n1372), .ZN(n1385) );
  INV_X4 U33 ( .A(n1373), .ZN(n1357) );
  NOR2_X4 U34 ( .A1(n1368), .A2(n3441), .ZN(n1373) );
  AOI22_X2 U39 ( .A1(u4_exp_in_mi1_7_), .A2(n1398), .B1(n1399), .B2(u4_N1976), 
        .ZN(n1397) );
  AOI22_X2 U97 ( .A1(u4_exp_in_mi1_6_), .A2(n1398), .B1(u4_exp_out_6_), .B2(
        n1399), .ZN(n1404) );
  AOI22_X2 U100 ( .A1(u4_exp_in_mi1_5_), .A2(n1398), .B1(u4_exp_out_5_), .B2(
        n1399), .ZN(n1406) );
  AOI22_X2 U103 ( .A1(u4_exp_in_mi1_4_), .A2(n1398), .B1(u4_exp_out_4_), .B2(
        n1399), .ZN(n1408) );
  AOI22_X2 U106 ( .A1(u4_exp_in_mi1_3_), .A2(n1398), .B1(u4_exp_out_3_), .B2(
        n1399), .ZN(n1410) );
  AOI22_X2 U109 ( .A1(u4_exp_in_mi1_2_), .A2(n1398), .B1(u4_exp_out_2_), .B2(
        n1399), .ZN(n1412) );
  AOI22_X2 U112 ( .A1(u4_exp_in_mi1_1_), .A2(n1398), .B1(u4_exp_out_1_), .B2(
        n1399), .ZN(n1414) );
  AOI22_X2 U115 ( .A1(n2473), .A2(n1398), .B1(n1399), .B2(u4_exp_out_0_), .ZN(
        n1416) );
  OAI221_X2 U120 ( .B1(n1419), .B2(n3581), .C1(n1420), .C2(n1421), .A(n1422), 
        .ZN(u4_shift_left[5]) );
  INV_X4 U122 ( .A(n1425), .ZN(n1419) );
  OAI211_X2 U123 ( .C1(n1421), .C2(n2722), .A(n1426), .B(n1427), .ZN(
        u4_shift_left[4]) );
  AOI22_X2 U125 ( .A1(u4_div_scht1a[4]), .A2(n1423), .B1(u4_exp_in_pl1_4_), 
        .B2(n1425), .ZN(n1426) );
  NAND2_X2 U126 ( .A1(n1429), .A2(n1430), .ZN(u4_shift_left[3]) );
  OAI211_X2 U129 ( .C1(n1421), .C2(n2723), .A(n1432), .B(n1433), .ZN(
        u4_shift_left[2]) );
  AOI22_X2 U131 ( .A1(u4_div_scht1a[2]), .A2(n1423), .B1(u4_exp_in_pl1_2_), 
        .B2(n1425), .ZN(n1432) );
  NAND2_X2 U132 ( .A1(n1434), .A2(n1435), .ZN(u4_shift_left[1]) );
  AOI221_X2 U133 ( .B1(u4_f2i_shft_1_), .B2(n2625), .C1(div_opa_ldz_r2[1]), 
        .C2(n1428), .A(n1436), .ZN(n1435) );
  OAI211_X2 U136 ( .C1(n1421), .C2(u4_fi_ldz_2a_0_), .A(n1441), .B(n1442), 
        .ZN(u4_shift_left[0]) );
  AOI22_X2 U139 ( .A1(u4_div_scht1a[0]), .A2(n1423), .B1(u4_exp_in_pl1_0_), 
        .B2(n1425), .ZN(n1441) );
  INV_X4 U140 ( .A(n1431), .ZN(n1421) );
  OAI211_X2 U141 ( .C1(n1438), .C2(n1445), .A(n1446), .B(n1447), .ZN(n1431) );
  INV_X4 U144 ( .A(n1439), .ZN(n1445) );
  INV_X4 U145 ( .A(n1450), .ZN(u4_fract_out_9_) );
  INV_X4 U146 ( .A(n1451), .ZN(u4_fract_out_8_) );
  INV_X4 U147 ( .A(n1452), .ZN(u4_fract_out_7_) );
  INV_X4 U148 ( .A(n1453), .ZN(u4_fract_out_3_) );
  INV_X4 U149 ( .A(n1454), .ZN(u4_fract_out_2_) );
  INV_X4 U150 ( .A(n1455), .ZN(u4_fract_out_22_) );
  INV_X4 U151 ( .A(n1456), .ZN(u4_fract_out_19_) );
  INV_X4 U152 ( .A(n1457), .ZN(u4_fract_out_18_) );
  INV_X4 U153 ( .A(n1458), .ZN(u4_fract_out_17_) );
  INV_X4 U154 ( .A(n1459), .ZN(u4_fract_out_13_) );
  INV_X4 U155 ( .A(n1460), .ZN(u4_fract_out_12_) );
  INV_X4 U156 ( .A(n1461), .ZN(u4_fract_out_11_) );
  NOR4_X2 U158 ( .A1(n3514), .A2(n1465), .A3(n1466), .A4(n1467), .ZN(n1464) );
  NOR4_X2 U159 ( .A1(fract_denorm[33]), .A2(n3544), .A3(n3547), .A4(n3513), 
        .ZN(n1467) );
  OAI211_X2 U163 ( .C1(n1477), .C2(n1478), .A(n1479), .B(n1480), .ZN(n1474) );
  AOI221_X2 U164 ( .B1(n1481), .B2(fract_denorm[36]), .C1(n1482), .C2(
        fract_denorm[40]), .A(n1483), .ZN(n1472) );
  NAND4_X2 U165 ( .A1(n1484), .A2(n1485), .A3(n1486), .A4(n1487), .ZN(n1470)
         );
  NAND4_X2 U166 ( .A1(n1469), .A2(n1488), .A3(fract_denorm[24]), .A4(n3537), 
        .ZN(n1484) );
  NOR4_X2 U168 ( .A1(n1491), .A2(n3512), .A3(n1492), .A4(n1493), .ZN(n1490) );
  NAND2_X2 U169 ( .A1(n1494), .A2(n3557), .ZN(n1486) );
  NOR4_X2 U172 ( .A1(n1499), .A2(n1500), .A3(n1501), .A4(n1502), .ZN(n1489) );
  NOR4_X2 U173 ( .A1(fract_denorm[38]), .A2(fract_denorm[37]), .A3(n3550), 
        .A4(n3513), .ZN(n1502) );
  AND4_X2 U174 ( .A1(n3542), .A2(n3540), .A3(fract_denorm[28]), .A4(n1469), 
        .ZN(n1501) );
  NAND4_X2 U176 ( .A1(n1506), .A2(n3552), .A3(n3554), .A4(n2680), .ZN(n1505)
         );
  NAND2_X2 U180 ( .A1(n1513), .A2(n3527), .ZN(n1495) );
  OAI211_X2 U183 ( .C1(n3556), .C2(n1519), .A(n3552), .B(n3554), .ZN(n1517) );
  OR2_X2 U184 ( .A1(fract_denorm[43]), .A2(fract_denorm[44]), .ZN(n1519) );
  NOR4_X2 U187 ( .A1(n3503), .A2(n3541), .A3(n3538), .A4(fract_denorm[27]), 
        .ZN(n1493) );
  AND4_X2 U188 ( .A1(n1522), .A2(n3502), .A3(n1523), .A4(n1524), .ZN(n1471) );
  AND4_X2 U189 ( .A1(n1504), .A2(n1525), .A3(n1526), .A4(n3508), .ZN(n1524) );
  OAI211_X2 U190 ( .C1(n3536), .C2(n1528), .A(n1529), .B(n1530), .ZN(n1527) );
  NAND2_X2 U194 ( .A1(n1534), .A2(n3522), .ZN(n1504) );
  NOR4_X2 U196 ( .A1(n3513), .A2(n3549), .A3(n3546), .A4(fract_denorm[35]), 
        .ZN(n1492) );
  NOR4_X2 U198 ( .A1(n1540), .A2(n1475), .A3(n1531), .A4(n1512), .ZN(n1539) );
  AND2_X2 U199 ( .A1(n1508), .A2(n3530), .ZN(n1512) );
  NAND4_X2 U202 ( .A1(n1487), .A2(n1468), .A3(n1480), .A4(n2680), .ZN(n1540)
         );
  AND2_X2 U208 ( .A1(n1498), .A2(n3524), .ZN(n1536) );
  NAND4_X2 U210 ( .A1(n1547), .A2(n1525), .A3(n1548), .A4(n1549), .ZN(n1500)
         );
  NOR4_X2 U211 ( .A1(n1550), .A2(n3509), .A3(n1465), .A4(n1520), .ZN(n1549) );
  AND3_X2 U213 ( .A1(n1551), .A2(fract_denorm[27]), .A3(n1469), .ZN(n1465) );
  NAND2_X2 U214 ( .A1(n1533), .A2(n3534), .ZN(n1485) );
  AND3_X2 U220 ( .A1(n3528), .A2(n1555), .A3(n1513), .ZN(n1518) );
  NAND2_X2 U221 ( .A1(n1556), .A2(n3559), .ZN(n1529) );
  AND2_X2 U222 ( .A1(n1557), .A2(n3563), .ZN(n1483) );
  NAND2_X2 U224 ( .A1(n1559), .A2(n3561), .ZN(n1547) );
  AOI22_X2 U225 ( .A1(n1560), .A2(n1481), .B1(n1561), .B2(n3554), .ZN(n1537)
         );
  AOI22_X2 U228 ( .A1(n2679), .A2(u4_exp_in_pl1_7_), .B1(n2680), .B2(
        u4_exp_next_mi_7_), .ZN(n1384) );
  AOI22_X2 U229 ( .A1(n2679), .A2(u4_exp_in_pl1_6_), .B1(n2680), .B2(
        u4_exp_next_mi_6_), .ZN(n1382) );
  AOI22_X2 U230 ( .A1(n2679), .A2(u4_exp_in_pl1_5_), .B1(n2680), .B2(
        u4_exp_next_mi_5_), .ZN(n1380) );
  AOI22_X2 U231 ( .A1(n2679), .A2(u4_exp_in_pl1_4_), .B1(n2680), .B2(
        u4_exp_next_mi_4_), .ZN(n1378) );
  AOI22_X2 U232 ( .A1(n2679), .A2(u4_exp_in_pl1_3_), .B1(n2680), .B2(
        u4_exp_next_mi_3_), .ZN(n1376) );
  AOI22_X2 U233 ( .A1(n2679), .A2(u4_exp_in_pl1_2_), .B1(n2680), .B2(
        u4_exp_next_mi_2_), .ZN(n1374) );
  OAI22_X2 U234 ( .A1(n2680), .A2(n3582), .B1(n2679), .B2(n3444), .ZN(
        u4_exp_out1_1_) );
  AOI22_X2 U235 ( .A1(n2679), .A2(u4_exp_in_pl1_0_), .B1(n2680), .B2(
        u4_exp_next_mi_0_), .ZN(n1356) );
  NAND4_X2 U237 ( .A1(u2_N12), .A2(u2_N11), .A3(n1565), .A4(n1566), .ZN(n1563)
         );
  AND4_X2 U238 ( .A1(u2_N6), .A2(u2_N7), .A3(u2_N8), .A4(u2_N9), .ZN(n1566) );
  NAND4_X2 U240 ( .A1(u2_N17), .A2(u2_N16), .A3(n1567), .A4(n1568), .ZN(n1562)
         );
  AND4_X2 U241 ( .A1(u2_N18), .A2(u2_N19), .A3(u2_N20), .A4(u2_N21), .ZN(n1568) );
  OAI222_X2 U243 ( .A1(u6_N23), .A2(n3486), .B1(n1570), .B2(n1564), .C1(
        u2_N124), .C2(n3480), .ZN(u2_underflow_d[1]) );
  OAI22_X2 U244 ( .A1(u2_N124), .A2(n1571), .B1(u6_N23), .B2(n1572), .ZN(n1564) );
  AND3_X2 U245 ( .A1(n1573), .A2(n1574), .A3(u2_N87), .ZN(u2_underflow_d[0])
         );
  AOI22_X2 U246 ( .A1(n3494), .A2(u2_N22), .B1(n2634), .B2(u2_N13), .ZN(n1582)
         );
  AOI22_X2 U247 ( .A1(n3494), .A2(u2_N21), .B1(n2635), .B2(u2_N12), .ZN(n1583)
         );
  AOI22_X2 U248 ( .A1(n3494), .A2(u2_N20), .B1(n2634), .B2(u2_N11), .ZN(n1584)
         );
  OAI22_X2 U249 ( .A1(n2634), .A2(n3410), .B1(n3494), .B2(n3404), .ZN(
        u2_exp_tmp1_4_) );
  AOI22_X2 U250 ( .A1(n3494), .A2(u2_N18), .B1(n2634), .B2(u2_N9), .ZN(n1585)
         );
  AOI22_X2 U251 ( .A1(n3494), .A2(u2_N17), .B1(n2634), .B2(u2_N8), .ZN(n1586)
         );
  AOI22_X2 U252 ( .A1(n3494), .A2(u2_N16), .B1(n2635), .B2(u2_N7), .ZN(n1587)
         );
  OAI22_X2 U253 ( .A1(n2635), .A2(n3411), .B1(n3494), .B2(n3409), .ZN(
        u2_exp_tmp1_0_) );
  OR3_X2 U255 ( .A1(n1590), .A2(n2634), .A3(n2466), .ZN(n1589) );
  NAND2_X2 U256 ( .A1(n2634), .A2(n2466), .ZN(n1588) );
  AOI22_X2 U257 ( .A1(u2_N14), .A2(n2634), .B1(u2_N23), .B2(n3494), .ZN(n1574)
         );
  AND2_X2 U258 ( .A1(opb_r[31]), .A2(opa_r[31]), .ZN(u2_N97) );
  NAND2_X2 U260 ( .A1(u2_N89), .A2(n3494), .ZN(n1592) );
  NAND2_X2 U261 ( .A1(n3485), .A2(n2461), .ZN(n1591) );
  OAI211_X2 U262 ( .C1(n1593), .C2(n1594), .A(n1595), .B(n1596), .ZN(u2_N65)
         );
  AOI22_X2 U263 ( .A1(u2_exp_tmp3_7_), .A2(n1597), .B1(u2_exp_tmp4_7_), .B2(
        n1598), .ZN(n1596) );
  AOI22_X2 U264 ( .A1(u2_N49), .A2(n1599), .B1(u2_N57), .B2(n1600), .ZN(n1595)
         );
  OAI211_X2 U265 ( .C1(n1575), .C2(n1594), .A(n1601), .B(n1602), .ZN(u2_N64)
         );
  AOI22_X2 U266 ( .A1(u2_exp_tmp3_6_), .A2(n1597), .B1(n1583), .B2(n1598), 
        .ZN(n1602) );
  AOI22_X2 U267 ( .A1(u2_N48), .A2(n1599), .B1(u2_N56), .B2(n1600), .ZN(n1601)
         );
  AOI22_X2 U268 ( .A1(u2_N30), .A2(n2635), .B1(u2_N39), .B2(n3494), .ZN(n1575)
         );
  OAI211_X2 U269 ( .C1(n1576), .C2(n1594), .A(n1603), .B(n1604), .ZN(u2_N63)
         );
  AOI22_X2 U270 ( .A1(u2_exp_tmp3_5_), .A2(n1597), .B1(n1584), .B2(n1598), 
        .ZN(n1604) );
  AOI22_X2 U271 ( .A1(u2_N47), .A2(n1599), .B1(u2_N55), .B2(n1600), .ZN(n1603)
         );
  AOI22_X2 U272 ( .A1(u2_N29), .A2(n2634), .B1(u2_N38), .B2(n3494), .ZN(n1576)
         );
  OAI211_X2 U273 ( .C1(n1577), .C2(n1594), .A(n1605), .B(n1606), .ZN(u2_N62)
         );
  AOI22_X2 U274 ( .A1(u2_exp_tmp3_4_), .A2(n1597), .B1(u2_exp_tmp4_4_), .B2(
        n1598), .ZN(n1606) );
  AOI22_X2 U275 ( .A1(u2_N46), .A2(n1599), .B1(u2_N54), .B2(n1600), .ZN(n1605)
         );
  AOI22_X2 U276 ( .A1(u2_N28), .A2(n2634), .B1(u2_N37), .B2(n3494), .ZN(n1577)
         );
  OAI211_X2 U277 ( .C1(n1578), .C2(n1594), .A(n1607), .B(n1608), .ZN(u2_N61)
         );
  AOI22_X2 U278 ( .A1(u2_exp_tmp3_3_), .A2(n1597), .B1(n1585), .B2(n1598), 
        .ZN(n1608) );
  AOI22_X2 U279 ( .A1(u2_N45), .A2(n1599), .B1(u2_N53), .B2(n1600), .ZN(n1607)
         );
  AOI22_X2 U280 ( .A1(u2_N27), .A2(n2635), .B1(u2_N36), .B2(n3494), .ZN(n1578)
         );
  OAI211_X2 U281 ( .C1(n1579), .C2(n1594), .A(n1609), .B(n1610), .ZN(u2_N60)
         );
  AOI22_X2 U282 ( .A1(u2_exp_tmp3_2_), .A2(n1597), .B1(n1586), .B2(n1598), 
        .ZN(n1610) );
  AOI22_X2 U283 ( .A1(u2_N44), .A2(n1599), .B1(u2_N52), .B2(n1600), .ZN(n1609)
         );
  AOI22_X2 U284 ( .A1(u2_N26), .A2(n2635), .B1(u2_N35), .B2(n3494), .ZN(n1579)
         );
  OAI211_X2 U285 ( .C1(n1580), .C2(n1594), .A(n1611), .B(n1612), .ZN(u2_N59)
         );
  AOI22_X2 U286 ( .A1(u2_exp_tmp3_1_), .A2(n1597), .B1(n1587), .B2(n1598), 
        .ZN(n1612) );
  AOI22_X2 U287 ( .A1(u2_N43), .A2(n1599), .B1(u2_N51), .B2(n1600), .ZN(n1611)
         );
  AOI22_X2 U288 ( .A1(u2_N25), .A2(n2634), .B1(u2_N34), .B2(n3494), .ZN(n1580)
         );
  OAI211_X2 U289 ( .C1(n1581), .C2(n1594), .A(n1613), .B(n1614), .ZN(u2_N58)
         );
  AOI22_X2 U290 ( .A1(u2_exp_tmp3_0_), .A2(n1597), .B1(u2_exp_tmp4_0_), .B2(
        n1598), .ZN(n1614) );
  AOI22_X2 U293 ( .A1(u2_N42), .A2(n1599), .B1(u2_exp_tmp1_0_), .B2(n1600), 
        .ZN(n1613) );
  NAND2_X2 U296 ( .A1(n3399), .A2(n1573), .ZN(n1594) );
  NAND2_X2 U297 ( .A1(n1590), .A2(n1615), .ZN(u2_exp_ovf_d_1_) );
  AOI22_X2 U300 ( .A1(u2_N31), .A2(n2634), .B1(u2_N40), .B2(n3494), .ZN(n1593)
         );
  AOI22_X2 U301 ( .A1(u2_N32), .A2(n2634), .B1(u2_N41), .B2(n3494), .ZN(n1590)
         );
  AOI22_X2 U302 ( .A1(u2_exp_tmp4_0_), .A2(n2634), .B1(u2_exp_tmp4_0_), .B2(
        n3494), .ZN(n1581) );
  OAI22_X2 U304 ( .A1(n2670), .A2(n2601), .B1(n1616), .B2(n2676), .ZN(
        u1_sign_d) );
  XNOR2_X2 U305 ( .A(opb_r[31]), .B(fpu_op_r1[0]), .ZN(n1616) );
  OAI22_X2 U306 ( .A1(n2670), .A2(n1617), .B1(n1618), .B2(n2675), .ZN(
        u1_fractb_s[9]) );
  OAI22_X2 U307 ( .A1(n2670), .A2(n1619), .B1(n1620), .B2(n2675), .ZN(
        u1_fractb_s[8]) );
  OAI22_X2 U308 ( .A1(n2670), .A2(n1621), .B1(n1622), .B2(n2675), .ZN(
        u1_fractb_s[7]) );
  OAI22_X2 U309 ( .A1(n2670), .A2(n1623), .B1(n1624), .B2(n2675), .ZN(
        u1_fractb_s[6]) );
  OAI22_X2 U310 ( .A1(n2670), .A2(n1625), .B1(n1626), .B2(n2676), .ZN(
        u1_fractb_s[5]) );
  OAI22_X2 U311 ( .A1(n2670), .A2(n1627), .B1(n1628), .B2(n2676), .ZN(
        u1_fractb_s[4]) );
  OAI22_X2 U312 ( .A1(n2670), .A2(n1629), .B1(n1630), .B2(n2676), .ZN(
        u1_fractb_s[3]) );
  OAI22_X2 U313 ( .A1(n2670), .A2(n1631), .B1(n2674), .B2(n1632), .ZN(
        u1_fractb_s[2]) );
  OAI22_X2 U314 ( .A1(n2670), .A2(n1633), .B1(n1634), .B2(n2676), .ZN(
        u1_fractb_s[26]) );
  OAI22_X2 U315 ( .A1(n2670), .A2(n1635), .B1(n1636), .B2(n2676), .ZN(
        u1_fractb_s[25]) );
  OAI22_X2 U316 ( .A1(n2670), .A2(n1637), .B1(n1638), .B2(n2676), .ZN(
        u1_fractb_s[24]) );
  OAI22_X2 U317 ( .A1(n2670), .A2(n1639), .B1(n1640), .B2(n2676), .ZN(
        u1_fractb_s[23]) );
  OAI22_X2 U318 ( .A1(n2670), .A2(n1641), .B1(n1642), .B2(n2676), .ZN(
        u1_fractb_s[22]) );
  OAI22_X2 U319 ( .A1(n2670), .A2(n1643), .B1(n1644), .B2(n2676), .ZN(
        u1_fractb_s[21]) );
  OAI22_X2 U320 ( .A1(n2670), .A2(n1645), .B1(n1646), .B2(n2676), .ZN(
        u1_fractb_s[20]) );
  OAI22_X2 U321 ( .A1(n2670), .A2(n1647), .B1(n2674), .B2(n1648), .ZN(
        u1_fractb_s[1]) );
  OAI22_X2 U322 ( .A1(n2670), .A2(n1649), .B1(n1650), .B2(n2676), .ZN(
        u1_fractb_s[19]) );
  OAI22_X2 U323 ( .A1(n2670), .A2(n1651), .B1(n1652), .B2(n2676), .ZN(
        u1_fractb_s[18]) );
  OAI22_X2 U324 ( .A1(n2670), .A2(n1653), .B1(n1654), .B2(n2676), .ZN(
        u1_fractb_s[17]) );
  OAI22_X2 U325 ( .A1(n2670), .A2(n1655), .B1(n1656), .B2(n2676), .ZN(
        u1_fractb_s[16]) );
  OAI22_X2 U326 ( .A1(n2670), .A2(n1657), .B1(n1658), .B2(n2676), .ZN(
        u1_fractb_s[15]) );
  OAI22_X2 U327 ( .A1(n2671), .A2(n1659), .B1(n1660), .B2(n2676), .ZN(
        u1_fractb_s[14]) );
  OAI22_X2 U328 ( .A1(n2671), .A2(n1661), .B1(n1662), .B2(n2676), .ZN(
        u1_fractb_s[13]) );
  OAI22_X2 U329 ( .A1(n2671), .A2(n1663), .B1(n1664), .B2(n2676), .ZN(
        u1_fractb_s[12]) );
  OAI22_X2 U330 ( .A1(n2671), .A2(n1665), .B1(n1666), .B2(n2676), .ZN(
        u1_fractb_s[11]) );
  OAI22_X2 U331 ( .A1(n2671), .A2(n1667), .B1(n1668), .B2(n2676), .ZN(
        u1_fractb_s[10]) );
  OAI22_X2 U332 ( .A1(n2671), .A2(n1669), .B1(n2674), .B2(n1670), .ZN(
        u1_fractb_s[0]) );
  OAI22_X2 U333 ( .A1(n1617), .A2(n2678), .B1(n2671), .B2(n1618), .ZN(
        u1_fracta_s[9]) );
  AOI22_X2 U334 ( .A1(n2661), .A2(u1_adj_op_out_sft_9_), .B1(n2656), .B2(u6_N6), .ZN(n1617) );
  OAI22_X2 U335 ( .A1(n1619), .A2(n2676), .B1(n2671), .B2(n1620), .ZN(
        u1_fracta_s[8]) );
  AOI22_X2 U336 ( .A1(n2660), .A2(u1_adj_op_out_sft_8_), .B1(n2655), .B2(u6_N5), .ZN(n1619) );
  OAI22_X2 U337 ( .A1(n1621), .A2(n2678), .B1(n2671), .B2(n1622), .ZN(
        u1_fracta_s[7]) );
  AOI22_X2 U338 ( .A1(n2660), .A2(u1_adj_op_out_sft_7_), .B1(n2655), .B2(u6_N4), .ZN(n1621) );
  OAI22_X2 U339 ( .A1(n1623), .A2(n2678), .B1(n2671), .B2(n1624), .ZN(
        u1_fracta_s[6]) );
  AOI22_X2 U340 ( .A1(n2660), .A2(u1_adj_op_out_sft_6_), .B1(n2656), .B2(u6_N3), .ZN(n1623) );
  OAI22_X2 U341 ( .A1(n1625), .A2(n2678), .B1(n2671), .B2(n1626), .ZN(
        u1_fracta_s[5]) );
  AOI22_X2 U342 ( .A1(n2660), .A2(u1_adj_op_out_sft_5_), .B1(n2655), .B2(u6_N2), .ZN(n1625) );
  OAI22_X2 U343 ( .A1(n1627), .A2(n2676), .B1(n2672), .B2(n1628), .ZN(
        u1_fracta_s[4]) );
  AOI22_X2 U344 ( .A1(n2660), .A2(u1_adj_op_out_sft_4_), .B1(n2655), .B2(u6_N1), .ZN(n1627) );
  OAI22_X2 U345 ( .A1(n1629), .A2(n2676), .B1(n2672), .B2(n1630), .ZN(
        u1_fracta_s[3]) );
  AOI22_X2 U346 ( .A1(n2660), .A2(u1_adj_op_out_sft_3_), .B1(n2655), .B2(u6_N0), .ZN(n1629) );
  OAI22_X2 U347 ( .A1(n2675), .A2(n1631), .B1(n2672), .B2(n1632), .ZN(
        u1_fracta_s[2]) );
  NAND2_X2 U348 ( .A1(u1_adj_op_out_sft_2_), .A2(n2664), .ZN(n1631) );
  OAI22_X2 U349 ( .A1(n1633), .A2(n2678), .B1(n2672), .B2(n1634), .ZN(
        u1_fracta_s[26]) );
  AOI22_X2 U350 ( .A1(n2660), .A2(u1_adj_op_out_sft_26_), .B1(n2656), .B2(
        u6_N23), .ZN(n1633) );
  OAI22_X2 U351 ( .A1(n1635), .A2(n2676), .B1(n2672), .B2(n1636), .ZN(
        u1_fracta_s[25]) );
  AOI22_X2 U352 ( .A1(n2661), .A2(u1_adj_op_out_sft_25_), .B1(n2655), .B2(
        u6_N22), .ZN(n1635) );
  OAI22_X2 U353 ( .A1(n1637), .A2(n2676), .B1(n2672), .B2(n1638), .ZN(
        u1_fracta_s[24]) );
  AOI22_X2 U354 ( .A1(n2661), .A2(u1_adj_op_out_sft_24_), .B1(n2655), .B2(
        u6_N21), .ZN(n1637) );
  OAI22_X2 U355 ( .A1(n1639), .A2(n2676), .B1(n2672), .B2(n1640), .ZN(
        u1_fracta_s[23]) );
  AOI22_X2 U356 ( .A1(n2661), .A2(u1_adj_op_out_sft_23_), .B1(n2655), .B2(
        u6_N20), .ZN(n1639) );
  OAI22_X2 U357 ( .A1(n1641), .A2(n2676), .B1(n2672), .B2(n1642), .ZN(
        u1_fracta_s[22]) );
  AOI22_X2 U358 ( .A1(n2661), .A2(u1_adj_op_out_sft_22_), .B1(n2656), .B2(
        u6_N19), .ZN(n1641) );
  OAI22_X2 U359 ( .A1(n1643), .A2(n2678), .B1(n2672), .B2(n1644), .ZN(
        u1_fracta_s[21]) );
  AOI22_X2 U360 ( .A1(n2661), .A2(u1_adj_op_out_sft_21_), .B1(n2655), .B2(
        u6_N18), .ZN(n1643) );
  OAI22_X2 U361 ( .A1(n1645), .A2(n2676), .B1(n2672), .B2(n1646), .ZN(
        u1_fracta_s[20]) );
  AOI22_X2 U362 ( .A1(n2661), .A2(u1_adj_op_out_sft_20_), .B1(n2655), .B2(
        u6_N17), .ZN(n1645) );
  OAI22_X2 U363 ( .A1(n2675), .A2(n1647), .B1(n2672), .B2(n1648), .ZN(
        u1_fracta_s[1]) );
  NAND2_X2 U364 ( .A1(u1_adj_op_out_sft_1_), .A2(n2664), .ZN(n1647) );
  OAI22_X2 U365 ( .A1(n1649), .A2(n2674), .B1(n2673), .B2(n1650), .ZN(
        u1_fracta_s[19]) );
  AOI22_X2 U366 ( .A1(n2661), .A2(u1_adj_op_out_sft_19_), .B1(n2655), .B2(
        u6_N16), .ZN(n1649) );
  OAI22_X2 U367 ( .A1(n1651), .A2(n2676), .B1(n2673), .B2(n1652), .ZN(
        u1_fracta_s[18]) );
  AOI22_X2 U368 ( .A1(n2661), .A2(u1_adj_op_out_sft_18_), .B1(n2656), .B2(
        u6_N15), .ZN(n1651) );
  OAI22_X2 U369 ( .A1(n1653), .A2(n2676), .B1(n2673), .B2(n1654), .ZN(
        u1_fracta_s[17]) );
  AOI22_X2 U370 ( .A1(n2661), .A2(u1_adj_op_out_sft_17_), .B1(n2655), .B2(
        u6_N14), .ZN(n1653) );
  OAI22_X2 U371 ( .A1(n1655), .A2(n2674), .B1(n2673), .B2(n1656), .ZN(
        u1_fracta_s[16]) );
  AOI22_X2 U372 ( .A1(n2661), .A2(u1_adj_op_out_sft_16_), .B1(n2656), .B2(
        u6_N13), .ZN(n1655) );
  OAI22_X2 U373 ( .A1(n1657), .A2(n2676), .B1(n2673), .B2(n1658), .ZN(
        u1_fracta_s[15]) );
  AOI22_X2 U374 ( .A1(n2661), .A2(u1_adj_op_out_sft_15_), .B1(n2656), .B2(
        u6_N12), .ZN(n1657) );
  OAI22_X2 U375 ( .A1(n1659), .A2(n2674), .B1(n2673), .B2(n1660), .ZN(
        u1_fracta_s[14]) );
  AOI22_X2 U376 ( .A1(n2661), .A2(u1_adj_op_out_sft_14_), .B1(n2656), .B2(
        u6_N11), .ZN(n1659) );
  OAI22_X2 U377 ( .A1(n1661), .A2(n2676), .B1(n2673), .B2(n1662), .ZN(
        u1_fracta_s[13]) );
  AOI22_X2 U378 ( .A1(n2661), .A2(u1_adj_op_out_sft_13_), .B1(n2656), .B2(
        u6_N10), .ZN(n1661) );
  OAI22_X2 U379 ( .A1(n1663), .A2(n2674), .B1(n2673), .B2(n1664), .ZN(
        u1_fracta_s[12]) );
  AOI22_X2 U380 ( .A1(n2661), .A2(u1_adj_op_out_sft_12_), .B1(n2656), .B2(
        u6_N9), .ZN(n1663) );
  OAI22_X2 U381 ( .A1(n1665), .A2(n2674), .B1(n2673), .B2(n1666), .ZN(
        u1_fracta_s[11]) );
  AOI22_X2 U382 ( .A1(n2661), .A2(u1_adj_op_out_sft_11_), .B1(n2656), .B2(
        u6_N8), .ZN(n1665) );
  OAI22_X2 U383 ( .A1(n1667), .A2(n2676), .B1(n2673), .B2(n1668), .ZN(
        u1_fracta_s[10]) );
  AOI22_X2 U384 ( .A1(n2661), .A2(u1_adj_op_out_sft_10_), .B1(n2656), .B2(
        u6_N7), .ZN(n1667) );
  OAI22_X2 U385 ( .A1(n2675), .A2(n1669), .B1(n2673), .B2(n1670), .ZN(
        u1_fracta_s[0]) );
  NAND2_X2 U386 ( .A1(n2664), .A2(n1671), .ZN(n1669) );
  AOI22_X2 U387 ( .A1(n2655), .A2(u1_adj_op_out_sft_9_), .B1(fracta_mul[6]), 
        .B2(n2663), .ZN(n1618) );
  AOI22_X2 U388 ( .A1(n2655), .A2(u1_adj_op_out_sft_8_), .B1(n2661), .B2(
        fracta_mul[5]), .ZN(n1620) );
  AOI22_X2 U389 ( .A1(n2655), .A2(u1_adj_op_out_sft_7_), .B1(n2662), .B2(
        fracta_mul[4]), .ZN(n1622) );
  AOI22_X2 U390 ( .A1(n2654), .A2(u1_adj_op_out_sft_6_), .B1(n2662), .B2(
        fracta_mul[3]), .ZN(n1624) );
  AOI22_X2 U391 ( .A1(n2655), .A2(u1_adj_op_out_sft_5_), .B1(n2662), .B2(
        fracta_mul[2]), .ZN(n1626) );
  AOI22_X2 U392 ( .A1(n2655), .A2(u1_adj_op_out_sft_4_), .B1(n2662), .B2(
        fracta_mul[1]), .ZN(n1628) );
  AOI22_X2 U393 ( .A1(n2655), .A2(u1_adj_op_out_sft_3_), .B1(n2662), .B2(
        fracta_mul[0]), .ZN(n1630) );
  NAND2_X2 U394 ( .A1(u1_adj_op_out_sft_2_), .A2(n2656), .ZN(n1632) );
  AOI22_X2 U395 ( .A1(n2654), .A2(u1_adj_op_out_sft_26_), .B1(n2651), .B2(
        n2663), .ZN(n1634) );
  AOI22_X2 U396 ( .A1(n2655), .A2(u1_adj_op_out_sft_25_), .B1(n2662), .B2(
        fracta_mul[22]), .ZN(n1636) );
  AOI22_X2 U397 ( .A1(n2655), .A2(u1_adj_op_out_sft_24_), .B1(n2662), .B2(
        fracta_mul[21]), .ZN(n1638) );
  AOI22_X2 U398 ( .A1(n2655), .A2(u1_adj_op_out_sft_23_), .B1(n2662), .B2(
        fracta_mul[20]), .ZN(n1640) );
  AOI22_X2 U399 ( .A1(n2655), .A2(u1_adj_op_out_sft_22_), .B1(n2662), .B2(
        fracta_mul[19]), .ZN(n1642) );
  AOI22_X2 U400 ( .A1(n2654), .A2(u1_adj_op_out_sft_21_), .B1(n2662), .B2(
        fracta_mul[18]), .ZN(n1644) );
  AOI22_X2 U401 ( .A1(n2655), .A2(u1_adj_op_out_sft_20_), .B1(n2662), .B2(
        fracta_mul[17]), .ZN(n1646) );
  NAND2_X2 U402 ( .A1(u1_adj_op_out_sft_1_), .A2(n2655), .ZN(n1648) );
  AOI22_X2 U403 ( .A1(n2655), .A2(u1_adj_op_out_sft_19_), .B1(n2662), .B2(
        fracta_mul[16]), .ZN(n1650) );
  AOI22_X2 U404 ( .A1(n2655), .A2(u1_adj_op_out_sft_18_), .B1(n2662), .B2(
        fracta_mul[15]), .ZN(n1652) );
  AOI22_X2 U405 ( .A1(n2655), .A2(u1_adj_op_out_sft_17_), .B1(n2661), .B2(
        fracta_mul[14]), .ZN(n1654) );
  AOI22_X2 U406 ( .A1(n2655), .A2(u1_adj_op_out_sft_16_), .B1(n2662), .B2(
        fracta_mul[13]), .ZN(n1656) );
  AOI22_X2 U407 ( .A1(n2655), .A2(u1_adj_op_out_sft_15_), .B1(n2661), .B2(
        fracta_mul[12]), .ZN(n1658) );
  AOI22_X2 U408 ( .A1(n2655), .A2(u1_adj_op_out_sft_14_), .B1(n2662), .B2(
        fracta_mul[11]), .ZN(n1660) );
  AOI22_X2 U409 ( .A1(n2655), .A2(u1_adj_op_out_sft_13_), .B1(n2661), .B2(
        fracta_mul[10]), .ZN(n1662) );
  AOI22_X2 U410 ( .A1(n2655), .A2(u1_adj_op_out_sft_12_), .B1(n2662), .B2(
        fracta_mul[9]), .ZN(n1664) );
  AOI22_X2 U411 ( .A1(n2655), .A2(u1_adj_op_out_sft_11_), .B1(n2661), .B2(
        fracta_mul[8]), .ZN(n1666) );
  AOI22_X2 U412 ( .A1(n2655), .A2(u1_adj_op_out_sft_10_), .B1(n2661), .B2(
        fracta_mul[7]), .ZN(n1668) );
  NAND2_X2 U413 ( .A1(n1671), .A2(n2656), .ZN(n1670) );
  AOI221_X2 U415 ( .B1(n1673), .B2(n3450), .C1(n1674), .C2(n1675), .A(n1676), 
        .ZN(n1672) );
  OAI22_X2 U418 ( .A1(n1682), .A2(n1683), .B1(n1684), .B2(n3447), .ZN(n1674)
         );
  AOI221_X2 U420 ( .B1(n1686), .B2(n3452), .C1(n3462), .C2(n3450), .A(n3469), 
        .ZN(n1682) );
  OAI211_X2 U421 ( .C1(n1687), .C2(n1688), .A(n1689), .B(n1690), .ZN(n1686) );
  NAND2_X2 U426 ( .A1(n1694), .A2(n1695), .ZN(n1680) );
  AND2_X2 U427 ( .A1(n1684), .A2(n1696), .ZN(n1694) );
  AND2_X2 U428 ( .A1(n1691), .A2(n1697), .ZN(n1684) );
  AND2_X2 U430 ( .A1(n1677), .A2(n1698), .ZN(n1691) );
  OAI22_X2 U432 ( .A1(n2466), .A2(n2658), .B1(n2663), .B2(n2461), .ZN(
        u1_exp_small[7]) );
  OAI22_X2 U433 ( .A1(n2657), .A2(n2577), .B1(n2663), .B2(n2476), .ZN(
        u1_exp_small[6]) );
  OAI22_X2 U434 ( .A1(n2658), .A2(n2494), .B1(n2663), .B2(n2574), .ZN(
        u1_exp_small[5]) );
  OAI22_X2 U435 ( .A1(n2657), .A2(n2477), .B1(n2663), .B2(n2573), .ZN(
        u1_exp_small[4]) );
  OAI22_X2 U436 ( .A1(n2658), .A2(n2495), .B1(n2663), .B2(n2572), .ZN(
        u1_exp_small[3]) );
  OAI22_X2 U437 ( .A1(n2658), .A2(n2478), .B1(n2663), .B2(n2575), .ZN(
        u1_exp_small[2]) );
  OAI22_X2 U438 ( .A1(n2657), .A2(n2576), .B1(n2663), .B2(n2570), .ZN(
        u1_exp_small[1]) );
  OAI22_X2 U439 ( .A1(n2657), .A2(n2467), .B1(n2663), .B2(n2571), .ZN(
        u1_exp_small[0]) );
  NAND2_X2 U440 ( .A1(n3449), .A2(n1707), .ZN(u1_exp_diff_sft_4_) );
  NAND2_X2 U442 ( .A1(u1_exp_diff_2_), .A2(n3449), .ZN(n1683) );
  AND2_X2 U445 ( .A1(u1_exp_diff2[7]), .A2(n1708), .ZN(u1_exp_diff_7_) );
  AND2_X2 U446 ( .A1(u1_exp_diff2[6]), .A2(n1708), .ZN(u1_exp_diff_6_) );
  AND2_X2 U447 ( .A1(u1_exp_diff2[5]), .A2(n1708), .ZN(u1_exp_diff_5_) );
  NAND2_X2 U448 ( .A1(u1_exp_diff2[4]), .A2(n1708), .ZN(n1707) );
  AND2_X2 U449 ( .A1(u1_exp_diff2[3]), .A2(n1708), .ZN(u1_exp_diff_3_) );
  AND2_X2 U450 ( .A1(u1_exp_diff2[2]), .A2(n1708), .ZN(u1_exp_diff_2_) );
  AND2_X2 U451 ( .A1(u1_exp_diff2[1]), .A2(n1708), .ZN(u1_exp_diff_1_) );
  AND2_X2 U452 ( .A1(u1_exp_diff2[0]), .A2(n1708), .ZN(u1_exp_diff_0_) );
  NAND2_X2 U453 ( .A1(n2653), .A2(n3485), .ZN(n1708) );
  AOI22_X2 U454 ( .A1(n2661), .A2(u6_N9), .B1(n2656), .B2(fracta_mul[9]), .ZN(
        n1688) );
  AOI22_X2 U455 ( .A1(n2661), .A2(u6_N8), .B1(n2655), .B2(fracta_mul[8]), .ZN(
        n1689) );
  AOI22_X2 U456 ( .A1(n2661), .A2(u6_N7), .B1(n2656), .B2(fracta_mul[7]), .ZN(
        n1709) );
  AOI22_X2 U457 ( .A1(n2661), .A2(u6_N6), .B1(n2655), .B2(fracta_mul[6]), .ZN(
        n1695) );
  AOI22_X2 U458 ( .A1(n2661), .A2(u6_N5), .B1(n2655), .B2(fracta_mul[5]), .ZN(
        n1696) );
  AOI22_X2 U459 ( .A1(n2661), .A2(u6_N4), .B1(n2657), .B2(fracta_mul[4]), .ZN(
        n1697) );
  AOI22_X2 U460 ( .A1(n2661), .A2(u6_N3), .B1(n2656), .B2(fracta_mul[3]), .ZN(
        n1698) );
  AOI22_X2 U461 ( .A1(n2661), .A2(u6_N2), .B1(n2657), .B2(fracta_mul[2]), .ZN(
        n1710) );
  OAI22_X2 U462 ( .A1(n2658), .A2(n2582), .B1(n2663), .B2(n2462), .ZN(
        u1_adj_op_22_) );
  AOI22_X2 U463 ( .A1(n2661), .A2(u6_N21), .B1(n2656), .B2(fracta_mul[21]), 
        .ZN(n1711) );
  OAI22_X2 U464 ( .A1(n2658), .A2(n2586), .B1(n2663), .B2(n2498), .ZN(
        u1_adj_op_20_) );
  AOI22_X2 U465 ( .A1(n2661), .A2(u6_N1), .B1(n2657), .B2(fracta_mul[1]), .ZN(
        n1712) );
  OAI22_X2 U466 ( .A1(n2658), .A2(n2499), .B1(n2663), .B2(n2580), .ZN(
        u1_adj_op_19_) );
  OAI22_X2 U467 ( .A1(n2658), .A2(n2583), .B1(n2664), .B2(n2496), .ZN(
        u1_adj_op_18_) );
  OAI22_X2 U468 ( .A1(n2658), .A2(n2479), .B1(n2663), .B2(n2581), .ZN(
        u1_adj_op_17_) );
  AOI22_X2 U469 ( .A1(n2661), .A2(u6_N16), .B1(n2655), .B2(fracta_mul[16]), 
        .ZN(n1713) );
  AOI22_X2 U470 ( .A1(n2661), .A2(u6_N15), .B1(n2657), .B2(fracta_mul[15]), 
        .ZN(n1714) );
  AOI22_X2 U471 ( .A1(n2661), .A2(u6_N14), .B1(n2655), .B2(fracta_mul[14]), 
        .ZN(n1715) );
  AOI22_X2 U472 ( .A1(n2661), .A2(u6_N13), .B1(n2656), .B2(fracta_mul[13]), 
        .ZN(n1716) );
  AOI22_X2 U473 ( .A1(n2661), .A2(u6_N12), .B1(n2657), .B2(fracta_mul[12]), 
        .ZN(n1717) );
  AOI22_X2 U474 ( .A1(n2661), .A2(u6_N11), .B1(n2657), .B2(fracta_mul[11]), 
        .ZN(n1718) );
  OAI22_X2 U475 ( .A1(n2658), .A2(n2585), .B1(n2663), .B2(n2497), .ZN(
        u1_adj_op_10_) );
  AOI22_X2 U476 ( .A1(n2661), .A2(u6_N0), .B1(n2657), .B2(fracta_mul[0]), .ZN(
        n1719) );
  AOI22_X2 U478 ( .A1(n2654), .A2(opb_r[30]), .B1(opa_r[30]), .B2(n2663), .ZN(
        n1699) );
  AOI22_X2 U480 ( .A1(n2654), .A2(opb_r[29]), .B1(n2662), .B2(opa_r[29]), .ZN(
        n1700) );
  AOI22_X2 U482 ( .A1(n2654), .A2(opb_r[28]), .B1(n2662), .B2(opa_r[28]), .ZN(
        n1701) );
  AOI22_X2 U484 ( .A1(n2654), .A2(opb_r[27]), .B1(n2662), .B2(opa_r[27]), .ZN(
        n1702) );
  AOI22_X2 U486 ( .A1(n2654), .A2(opb_r[26]), .B1(n2662), .B2(opa_r[26]), .ZN(
        n1703) );
  AOI22_X2 U488 ( .A1(n2654), .A2(opb_r[25]), .B1(n2663), .B2(opa_r[25]), .ZN(
        n1704) );
  AOI22_X2 U490 ( .A1(n2654), .A2(opb_r[24]), .B1(n2663), .B2(opa_r[24]), .ZN(
        n1705) );
  AOI22_X2 U492 ( .A1(n2654), .A2(opb_r[23]), .B1(n2663), .B2(opa_r[23]), .ZN(
        n1706) );
  AND3_X2 U493 ( .A1(u1_N131), .A2(n1721), .A3(u1_N34), .ZN(n1720) );
  XOR2_X2 U495 ( .A(fpu_op_r1[0]), .B(u2_sign_d), .Z(n1721) );
  XNOR2_X2 U496 ( .A(n2601), .B(opb_r[31]), .ZN(u2_sign_d) );
  AOI221_X2 U500 ( .B1(opb_nan), .B2(n1725), .C1(n1726), .C2(
        u1_fracta_lt_fractb), .A(u1_signa_r), .ZN(n1722) );
  NAND2_X2 U502 ( .A1(opa_nan), .A2(opb_nan), .ZN(n1725) );
  OAI22_X2 U503 ( .A1(n2604), .A2(n1727), .B1(n1728), .B2(n1729), .ZN(u1_N129)
         );
  XNOR2_X2 U504 ( .A(n2600), .B(u1_add_r), .ZN(n1729) );
  AND2_X2 U505 ( .A1(n1727), .A2(n2604), .ZN(n1728) );
  AOI22_X2 U506 ( .A1(u0_snan_r_a), .A2(u0_expa_ff), .B1(u0_snan_r_b), .B2(
        u0_expb_ff), .ZN(n1730) );
  AOI22_X2 U507 ( .A1(u0_qnan_r_a), .A2(u0_expa_ff), .B1(u0_qnan_r_b), .B2(
        u0_expb_ff), .ZN(n1731) );
  NAND2_X2 U508 ( .A1(n1732), .A2(n1733), .ZN(u0_N7) );
  AND2_X2 U512 ( .A1(u0_fractb_00), .A2(u0_expb_00), .ZN(u0_N17) );
  AND2_X2 U513 ( .A1(u0_fracta_00), .A2(u0_expa_00), .ZN(u0_N16) );
  NAND2_X2 U514 ( .A1(u0_infb_f_r), .A2(u0_expb_ff), .ZN(n1732) );
  NAND2_X2 U515 ( .A1(u0_infa_f_r), .A2(u0_expa_ff), .ZN(n1733) );
  NAND2_X2 U518 ( .A1(n1738), .A2(n1739), .ZN(n1736) );
  NOR4_X2 U519 ( .A1(n2466), .A2(n2577), .A3(n2494), .A4(n2477), .ZN(n1739) );
  NOR4_X2 U520 ( .A1(n2495), .A2(n2478), .A3(n2576), .A4(n2467), .ZN(n1738) );
  NAND2_X2 U521 ( .A1(n1740), .A2(n1741), .ZN(n1737) );
  NOR4_X2 U522 ( .A1(n2461), .A2(n2476), .A3(n2574), .A4(n2573), .ZN(n1741) );
  NOR4_X2 U523 ( .A1(n2572), .A2(n2575), .A3(n2570), .A4(n2571), .ZN(n1740) );
  OAI22_X2 U524 ( .A1(n3485), .A2(n2658), .B1(n2663), .B2(n2652), .ZN(n2459)
         );
  NAND2_X2 U525 ( .A1(n1735), .A2(n2462), .ZN(n1571) );
  AND4_X2 U526 ( .A1(n1742), .A2(n1743), .A3(n1744), .A4(n1745), .ZN(n1735) );
  NOR4_X2 U527 ( .A1(fracta_mul[8]), .A2(fracta_mul[6]), .A3(fracta_mul[5]), 
        .A4(fracta_mul[4]), .ZN(n1745) );
  NOR4_X2 U528 ( .A1(fracta_mul[3]), .A2(fracta_mul[2]), .A3(fracta_mul[20]), 
        .A4(fracta_mul[1]), .ZN(n1744) );
  NOR4_X2 U529 ( .A1(fracta_mul[18]), .A2(fracta_mul[16]), .A3(fracta_mul[14]), 
        .A4(fracta_mul[12]), .ZN(n1743) );
  NAND2_X2 U531 ( .A1(n1747), .A2(n1748), .ZN(u6_N23) );
  NOR4_X2 U532 ( .A1(opb_r[30]), .A2(opb_r[29]), .A3(opb_r[28]), .A4(opb_r[27]), .ZN(n1748) );
  NOR4_X2 U533 ( .A1(opb_r[26]), .A2(opb_r[25]), .A3(opb_r[24]), .A4(opb_r[23]), .ZN(n1747) );
  NAND2_X2 U534 ( .A1(n1734), .A2(n2582), .ZN(n1572) );
  AND4_X2 U535 ( .A1(n1749), .A2(n1750), .A3(n1751), .A4(n1752), .ZN(n1734) );
  NOR4_X2 U536 ( .A1(n1753), .A2(u6_N4), .A3(u6_N6), .A4(u6_N5), .ZN(n1752) );
  OR3_X2 U537 ( .A1(u6_N8), .A2(u6_N9), .A3(u6_N7), .ZN(n1753) );
  NOR4_X2 U538 ( .A1(n1754), .A2(u6_N21), .A3(u6_N3), .A4(u6_N2), .ZN(n1751)
         );
  OR2_X2 U539 ( .A1(u6_N1), .A2(u6_N20), .ZN(n1754) );
  NOR4_X2 U540 ( .A1(n1755), .A2(u6_N14), .A3(u6_N16), .A4(u6_N15), .ZN(n1750)
         );
  NOR4_X2 U542 ( .A1(n1756), .A2(u6_N11), .A3(u6_N13), .A4(u6_N12), .ZN(n1749)
         );
  OR2_X2 U543 ( .A1(u6_N0), .A2(u6_N10), .ZN(n1756) );
  AOI22_X2 U544 ( .A1(u3_N40), .A2(n2470), .B1(u3_N12), .B2(fasu_op), .ZN(
        n1757) );
  AOI22_X2 U545 ( .A1(u3_N39), .A2(n2470), .B1(u3_N11), .B2(fasu_op), .ZN(
        n1758) );
  AOI22_X2 U546 ( .A1(u3_N38), .A2(n2470), .B1(u3_N10), .B2(fasu_op), .ZN(
        n1759) );
  AOI22_X2 U547 ( .A1(u3_N37), .A2(n2470), .B1(u3_N9), .B2(fasu_op), .ZN(n1760) );
  AOI22_X2 U548 ( .A1(u3_N36), .A2(n2470), .B1(u3_N8), .B2(fasu_op), .ZN(n1761) );
  AOI22_X2 U549 ( .A1(u3_N35), .A2(n2470), .B1(u3_N7), .B2(fasu_op), .ZN(n1762) );
  AOI22_X2 U550 ( .A1(u3_N34), .A2(n2470), .B1(u3_N6), .B2(fasu_op), .ZN(n1763) );
  AOI22_X2 U551 ( .A1(u3_N33), .A2(n2470), .B1(u3_N5), .B2(fasu_op), .ZN(n1764) );
  AOI22_X2 U552 ( .A1(u3_N57), .A2(n2689), .B1(u3_N29), .B2(fasu_op), .ZN(
        n1765) );
  AOI22_X2 U553 ( .A1(u3_N56), .A2(n2689), .B1(u3_N28), .B2(n2688), .ZN(n1766)
         );
  AOI22_X2 U554 ( .A1(u3_N55), .A2(n2689), .B1(u3_N27), .B2(n2688), .ZN(n1767)
         );
  AOI22_X2 U555 ( .A1(u3_N54), .A2(n2689), .B1(u3_N26), .B2(n2688), .ZN(n1768)
         );
  AOI22_X2 U556 ( .A1(u3_N53), .A2(n2689), .B1(u3_N25), .B2(n2688), .ZN(n1769)
         );
  AOI22_X2 U557 ( .A1(u3_N52), .A2(n2689), .B1(u3_N24), .B2(n2688), .ZN(n1770)
         );
  AOI22_X2 U558 ( .A1(u3_N51), .A2(n2689), .B1(u3_N23), .B2(n2688), .ZN(n1771)
         );
  AOI22_X2 U559 ( .A1(u3_N32), .A2(n2689), .B1(u3_N4), .B2(n2688), .ZN(n1772)
         );
  AOI22_X2 U560 ( .A1(u3_N50), .A2(n2689), .B1(u3_N22), .B2(n2688), .ZN(n1773)
         );
  AOI22_X2 U561 ( .A1(u3_N49), .A2(n2689), .B1(u3_N21), .B2(n2688), .ZN(n1774)
         );
  AOI22_X2 U562 ( .A1(u3_N48), .A2(n2689), .B1(u3_N20), .B2(n2688), .ZN(n1775)
         );
  AOI22_X2 U563 ( .A1(u3_N47), .A2(n2689), .B1(u3_N19), .B2(n2688), .ZN(n1776)
         );
  AOI22_X2 U564 ( .A1(u3_N46), .A2(n2689), .B1(u3_N18), .B2(n2688), .ZN(n1777)
         );
  AOI22_X2 U565 ( .A1(u3_N45), .A2(n2689), .B1(u3_N17), .B2(n2688), .ZN(n1778)
         );
  AOI22_X2 U566 ( .A1(u3_N44), .A2(n2689), .B1(u3_N16), .B2(fasu_op), .ZN(
        n1779) );
  AOI22_X2 U567 ( .A1(u3_N43), .A2(n2689), .B1(u3_N15), .B2(fasu_op), .ZN(
        n1780) );
  AOI22_X2 U568 ( .A1(u3_N42), .A2(n2689), .B1(u3_N14), .B2(fasu_op), .ZN(
        n1781) );
  AOI22_X2 U569 ( .A1(u3_N41), .A2(n2689), .B1(u3_N13), .B2(fasu_op), .ZN(
        n1782) );
  AOI22_X2 U570 ( .A1(u3_N31), .A2(n2689), .B1(u3_N3), .B2(fasu_op), .ZN(n1783) );
  NAND2_X2 U572 ( .A1(quo[49]), .A2(opb_dn), .ZN(n1784) );
  OR2_X2 U573 ( .A1(N195), .A2(u2_N124), .ZN(u6_N49) );
  AOI22_X2 U574 ( .A1(u2_N124), .A2(fracta_mul[22]), .B1(n2653), .B2(N194), 
        .ZN(n1792) );
  AOI22_X2 U575 ( .A1(u2_N124), .A2(fracta_mul[21]), .B1(n2653), .B2(N193), 
        .ZN(n1793) );
  AOI22_X2 U576 ( .A1(u2_N124), .A2(fracta_mul[20]), .B1(n2653), .B2(N192), 
        .ZN(n1794) );
  AOI22_X2 U577 ( .A1(u2_N124), .A2(fracta_mul[19]), .B1(n2653), .B2(N191), 
        .ZN(n1795) );
  AOI22_X2 U578 ( .A1(u2_N124), .A2(fracta_mul[18]), .B1(n2653), .B2(N190), 
        .ZN(n1796) );
  AOI22_X2 U579 ( .A1(u2_N124), .A2(fracta_mul[17]), .B1(n2653), .B2(N189), 
        .ZN(n1797) );
  AOI22_X2 U580 ( .A1(u2_N124), .A2(fracta_mul[16]), .B1(n2653), .B2(N188), 
        .ZN(n1798) );
  AOI22_X2 U581 ( .A1(u2_N124), .A2(fracta_mul[15]), .B1(n2653), .B2(N187), 
        .ZN(n1799) );
  AOI22_X2 U582 ( .A1(u2_N124), .A2(fracta_mul[14]), .B1(n2653), .B2(N186), 
        .ZN(n1800) );
  AOI22_X2 U583 ( .A1(u2_N124), .A2(fracta_mul[13]), .B1(n2653), .B2(N185), 
        .ZN(n1801) );
  AOI22_X2 U584 ( .A1(u2_N124), .A2(fracta_mul[12]), .B1(n2653), .B2(N184), 
        .ZN(n1802) );
  AOI22_X2 U585 ( .A1(u2_N124), .A2(fracta_mul[11]), .B1(n2653), .B2(N183), 
        .ZN(n1803) );
  AOI22_X2 U586 ( .A1(u2_N124), .A2(fracta_mul[10]), .B1(n2652), .B2(N182), 
        .ZN(n1804) );
  AOI22_X2 U587 ( .A1(u2_N124), .A2(fracta_mul[9]), .B1(n2652), .B2(N181), 
        .ZN(n1805) );
  AOI22_X2 U588 ( .A1(u2_N124), .A2(fracta_mul[8]), .B1(n2652), .B2(N180), 
        .ZN(n1806) );
  AOI22_X2 U589 ( .A1(u2_N124), .A2(fracta_mul[7]), .B1(n2652), .B2(N179), 
        .ZN(n1807) );
  AOI22_X2 U590 ( .A1(u2_N124), .A2(fracta_mul[6]), .B1(n2652), .B2(N178), 
        .ZN(n1808) );
  AOI22_X2 U591 ( .A1(u2_N124), .A2(fracta_mul[5]), .B1(n2652), .B2(N177), 
        .ZN(n1809) );
  AOI22_X2 U592 ( .A1(u2_N124), .A2(fracta_mul[4]), .B1(n2652), .B2(N176), 
        .ZN(n1810) );
  AOI22_X2 U593 ( .A1(u2_N124), .A2(fracta_mul[3]), .B1(n2652), .B2(N175), 
        .ZN(n1811) );
  AOI22_X2 U594 ( .A1(u2_N124), .A2(fracta_mul[2]), .B1(n2652), .B2(N174), 
        .ZN(n1812) );
  AOI22_X2 U595 ( .A1(u2_N124), .A2(fracta_mul[1]), .B1(n2652), .B2(N173), 
        .ZN(n1813) );
  AOI22_X2 U596 ( .A1(u2_N124), .A2(fracta_mul[0]), .B1(n2652), .B2(N172), 
        .ZN(n1814) );
  NAND2_X2 U597 ( .A1(n1815), .A2(n1816), .ZN(u2_N124) );
  NOR4_X2 U598 ( .A1(opa_r[30]), .A2(opa_r[29]), .A3(opa_r[28]), .A4(opa_r[27]), .ZN(n1816) );
  NOR4_X2 U599 ( .A1(opa_r[26]), .A2(opa_r[25]), .A3(opa_r[24]), .A4(opa_r[23]), .ZN(n1815) );
  AOI22_X2 U600 ( .A1(u3_N58), .A2(n2689), .B1(u3_N30), .B2(fasu_op), .ZN(
        n1817) );
  NOR4_X2 U601 ( .A1(fracta_mul[16]), .A2(n1818), .A3(n1819), .A4(n1820), .ZN(
        N75) );
  NAND4_X2 U603 ( .A1(exp_mul[7]), .A2(exp_mul[6]), .A3(exp_mul[5]), .A4(
        exp_mul[4]), .ZN(n1822) );
  NAND4_X2 U604 ( .A1(exp_mul[3]), .A2(exp_mul[2]), .A3(exp_mul[1]), .A4(
        exp_mul[0]), .ZN(n1821) );
  AND4_X2 U605 ( .A1(opb_00), .A2(opa_nan_r), .A3(n2596), .A4(n2503), .ZN(N533) );
  OAI211_X2 U607 ( .C1(n3518), .C2(n1824), .A(n1825), .B(n1826), .ZN(N531) );
  NOR4_X2 U609 ( .A1(n1830), .A2(n1831), .A3(n2474), .A4(n3573), .ZN(n1827) );
  OR2_X2 U610 ( .A1(inf_mul2), .A2(inf_mul_r), .ZN(n1831) );
  NAND4_X2 U611 ( .A1(n1833), .A2(n1834), .A3(n1835), .A4(n1836), .ZN(n1825)
         );
  NAND4_X2 U618 ( .A1(n1845), .A2(n1846), .A3(n1847), .A4(n1848), .ZN(n1841)
         );
  NOR4_X2 U619 ( .A1(n1849), .A2(n1850), .A3(n1851), .A4(n1852), .ZN(n1848) );
  OR3_X2 U620 ( .A1(n1853), .A2(n1854), .A3(n1855), .ZN(n1849) );
  NOR4_X2 U621 ( .A1(n1856), .A2(n1857), .A3(n1858), .A4(n1859), .ZN(n1847) );
  NOR4_X2 U623 ( .A1(n1863), .A2(n1864), .A3(n1865), .A4(n1866), .ZN(n1846) );
  NOR4_X2 U625 ( .A1(n1870), .A2(n1871), .A3(n1872), .A4(n1873), .ZN(n1845) );
  AOI221_X2 U628 ( .B1(underflow_fmul_r[2]), .B2(n1881), .C1(
        underflow_fmul_r[1]), .C2(n1882), .A(n1883), .ZN(n1880) );
  OR2_X2 U629 ( .A1(underflow_fmul_r[0]), .A2(n1884), .ZN(n1883) );
  NAND4_X2 U632 ( .A1(n1889), .A2(n1890), .A3(n1891), .A4(n1892), .ZN(n1888)
         );
  NOR4_X2 U633 ( .A1(n1893), .A2(prod[26]), .A3(prod[28]), .A4(prod[27]), .ZN(
        n1892) );
  OR3_X2 U634 ( .A1(prod[2]), .A2(prod[30]), .A3(prod[29]), .ZN(n1893) );
  NOR4_X2 U635 ( .A1(n1894), .A2(prod[20]), .A3(prod[22]), .A4(prod[21]), .ZN(
        n1891) );
  NOR4_X2 U637 ( .A1(n1895), .A2(prod[15]), .A3(prod[17]), .A4(prod[16]), .ZN(
        n1890) );
  OR3_X2 U638 ( .A1(prod[19]), .A2(prod[1]), .A3(prod[18]), .ZN(n1895) );
  NOR4_X2 U639 ( .A1(n1896), .A2(prod[0]), .A3(prod[11]), .A4(prod[10]), .ZN(
        n1889) );
  OR3_X2 U640 ( .A1(prod[13]), .A2(prod[14]), .A3(prod[12]), .ZN(n1896) );
  NAND4_X2 U641 ( .A1(n1897), .A2(n1898), .A3(n1899), .A4(n1900), .ZN(n1887)
         );
  NOR4_X2 U642 ( .A1(n1901), .A2(prod[4]), .A3(prod[6]), .A4(prod[5]), .ZN(
        n1900) );
  OR3_X2 U643 ( .A1(prod[8]), .A2(prod[9]), .A3(prod[7]), .ZN(n1901) );
  NOR4_X2 U644 ( .A1(n1902), .A2(prod[45]), .A3(prod[47]), .A4(prod[46]), .ZN(
        n1899) );
  NOR4_X2 U646 ( .A1(n1903), .A2(prod[37]), .A3(prod[39]), .A4(prod[38]), .ZN(
        n1898) );
  OR3_X2 U647 ( .A1(prod[40]), .A2(prod[41]), .A3(prod[3]), .ZN(n1903) );
  NOR4_X2 U648 ( .A1(n1904), .A2(prod[31]), .A3(prod[33]), .A4(prod[32]), .ZN(
        n1897) );
  NAND4_X2 U651 ( .A1(n1908), .A2(n1909), .A3(n1910), .A4(n1911), .ZN(n1907)
         );
  NOR4_X2 U652 ( .A1(n1912), .A2(n1913), .A3(n1852), .A4(n1850), .ZN(n1911) );
  NOR4_X2 U654 ( .A1(n1917), .A2(n1918), .A3(n1859), .A4(n1857), .ZN(n1910) );
  NOR4_X2 U656 ( .A1(n1920), .A2(n1921), .A3(n1866), .A4(n1864), .ZN(n1909) );
  NAND4_X2 U660 ( .A1(n1925), .A2(n1926), .A3(n1927), .A4(n1928), .ZN(n1906)
         );
  NAND4_X2 U661 ( .A1(n1929), .A2(n1930), .A3(n1931), .A4(n1932), .ZN(n1905)
         );
  NAND2_X2 U662 ( .A1(n1829), .A2(n2624), .ZN(n1879) );
  OAI221_X2 U664 ( .B1(n1939), .B2(n3567), .C1(n1940), .C2(n2491), .A(n1941), 
        .ZN(N509) );
  AOI22_X2 U667 ( .A1(n1944), .A2(n2624), .B1(n2490), .B2(n1943), .ZN(n1939)
         );
  AND2_X2 U669 ( .A1(n1842), .A2(n1830), .ZN(n1946) );
  INV_X4 U675 ( .A(n1882), .ZN(n1878) );
  NAND2_X2 U676 ( .A1(n1950), .A2(n1951), .ZN(n1882) );
  NAND4_X2 U677 ( .A1(n1952), .A2(n1854), .A3(n1953), .A4(n1954), .ZN(n1951)
         );
  NAND4_X2 U685 ( .A1(u4_N1606), .A2(n1969), .A3(n1970), .A4(n2486), .ZN(n1968) );
  OR4_X2 U686 ( .A1(n2682), .A2(n2683), .A3(n2684), .A4(n2685), .ZN(n1967) );
  XNOR2_X2 U689 ( .A(n2687), .B(n1975), .ZN(n1974) );
  NOR4_X2 U690 ( .A1(n3352), .A2(n3351), .A3(n3350), .A4(n3349), .ZN(n1973) );
  NAND2_X2 U692 ( .A1(u4_div_exp3[4]), .A2(n1363), .ZN(n1978) );
  NAND2_X2 U695 ( .A1(u4_div_exp3[3]), .A2(n1363), .ZN(n1981) );
  NAND2_X2 U698 ( .A1(u4_div_exp3[2]), .A2(n1363), .ZN(n1984) );
  NAND2_X2 U701 ( .A1(u4_div_exp3[1]), .A2(n1363), .ZN(n1987) );
  NOR4_X2 U703 ( .A1(n3348), .A2(n3347), .A3(n3346), .A4(n1444), .ZN(n1972) );
  NAND2_X2 U705 ( .A1(u4_div_exp3[7]), .A2(n1363), .ZN(n1989) );
  NAND2_X2 U708 ( .A1(u4_div_exp3[6]), .A2(n1363), .ZN(n1992) );
  NAND2_X2 U711 ( .A1(u4_div_exp3[5]), .A2(n1363), .ZN(n1995) );
  OAI22_X2 U716 ( .A1(exp_ovf_r[1]), .A2(n1996), .B1(n2492), .B2(n1997), .ZN(
        n1963) );
  AND2_X2 U718 ( .A1(u4_N1600), .A2(n1966), .ZN(n1998) );
  NAND2_X2 U719 ( .A1(n2624), .A2(n1999), .ZN(n1950) );
  NOR4_X2 U720 ( .A1(u4_exp_in_mi1_8_), .A2(exp_ovf_r[1]), .A3(n3583), .A4(
        n2003), .ZN(n2001) );
  INV_X4 U721 ( .A(n2004), .ZN(n1940) );
  OAI221_X2 U722 ( .B1(n3498), .B2(n2002), .C1(n2005), .C2(n2465), .A(n2006), 
        .ZN(n2004) );
  AOI221_X2 U723 ( .B1(n2007), .B2(n2008), .C1(n2490), .C2(n1966), .A(n1956), 
        .ZN(n2006) );
  NOR4_X2 U726 ( .A1(n2687), .A2(n1389), .A3(n2584), .A4(n2500), .ZN(n2009) );
  INV_X4 U727 ( .A(n2011), .ZN(n1935) );
  OAI22_X2 U728 ( .A1(n2012), .A2(n2649), .B1(n2490), .B2(n2013), .ZN(n2011)
         );
  NOR4_X2 U730 ( .A1(n2016), .A2(n1956), .A3(n2017), .A4(n2018), .ZN(n2012) );
  INV_X4 U731 ( .A(n2019), .ZN(n2016) );
  NAND4_X2 U734 ( .A1(n1828), .A2(n1829), .A3(opas_r2), .A4(n3487), .ZN(n2021)
         );
  AOI22_X2 U735 ( .A1(n2022), .A2(n2023), .B1(n2024), .B2(n3519), .ZN(n2020)
         );
  OAI22_X2 U736 ( .A1(n1833), .A2(n2025), .B1(n2026), .B2(n3516), .ZN(n2024)
         );
  AOI22_X2 U737 ( .A1(n2027), .A2(n3572), .B1(n2028), .B2(n2599), .ZN(n2026)
         );
  NAND2_X2 U739 ( .A1(opb_inf), .A2(opa_inf), .ZN(n1836) );
  NAND2_X2 U740 ( .A1(n2599), .A2(n1835), .ZN(n2027) );
  AOI22_X2 U741 ( .A1(n3576), .A2(n2029), .B1(nan_sign_d), .B2(n2030), .ZN(
        n2025) );
  INV_X4 U742 ( .A(n2031), .ZN(n2029) );
  AOI22_X2 U743 ( .A1(sign_fasu_r), .A2(n1824), .B1(result_zero_sign_d), .B2(
        n2032), .ZN(n2031) );
  INV_X4 U744 ( .A(n2032), .ZN(n1824) );
  NAND2_X2 U747 ( .A1(n1829), .A2(n2602), .ZN(n2030) );
  XNOR2_X2 U749 ( .A(n2599), .B(n2033), .ZN(n2023) );
  NAND4_X2 U753 ( .A1(n2034), .A2(n2035), .A3(n2036), .A4(n2037), .ZN(n1830)
         );
  NOR4_X2 U754 ( .A1(n2038), .A2(n2039), .A3(n2040), .A4(n2041), .ZN(n2037) );
  NAND4_X2 U755 ( .A1(n1922), .A2(n1869), .A3(n1867), .A4(n1868), .ZN(n2041)
         );
  NAND4_X2 U756 ( .A1(n2042), .A2(n2043), .A3(n1919), .A4(n1862), .ZN(n2040)
         );
  NAND4_X2 U757 ( .A1(n1860), .A2(n1861), .A3(n2044), .A4(n2045), .ZN(n2039)
         );
  NAND4_X2 U758 ( .A1(n1916), .A2(n1914), .A3(n1915), .A4(n1932), .ZN(n2038)
         );
  AND4_X2 U759 ( .A1(n2046), .A2(n1925), .A3(n1927), .A4(n1926), .ZN(n2036) );
  AND4_X2 U760 ( .A1(n1928), .A2(n1929), .A3(n1930), .A4(n1931), .ZN(n2046) );
  NOR4_X2 U761 ( .A1(n1866), .A2(n1864), .A3(n1921), .A4(n2047), .ZN(n2035) );
  NOR4_X2 U762 ( .A1(n2048), .A2(n1872), .A3(n1873), .A4(n1871), .ZN(n2034) );
  NAND2_X2 U763 ( .A1(n1925), .A2(n2049), .ZN(N475) );
  NAND2_X2 U764 ( .A1(n1926), .A2(n2049), .ZN(N474) );
  NAND2_X2 U765 ( .A1(n1927), .A2(n2049), .ZN(N473) );
  NAND2_X2 U766 ( .A1(n1928), .A2(n2049), .ZN(N472) );
  NAND2_X2 U767 ( .A1(n1929), .A2(n2049), .ZN(N471) );
  NAND2_X2 U768 ( .A1(n1930), .A2(n2049), .ZN(N470) );
  NOR4_X2 U769 ( .A1(fracta_mul[16]), .A2(n1819), .A3(n1820), .A4(n3482), .ZN(
        N47) );
  OR3_X2 U771 ( .A1(fracta_mul[13]), .A2(fracta_mul[15]), .A3(fracta_mul[14]), 
        .ZN(n2051) );
  OR2_X2 U772 ( .A1(n2052), .A2(fracta_mul[19]), .ZN(n1820) );
  NAND2_X2 U773 ( .A1(n1931), .A2(n2049), .ZN(N469) );
  NAND2_X2 U774 ( .A1(n1932), .A2(n2049), .ZN(N468) );
  OAI22_X2 U775 ( .A1(n1877), .A2(n2049), .B1(n3490), .B2(n2053), .ZN(N467) );
  INV_X4 U776 ( .A(n1871), .ZN(n2053) );
  OAI211_X2 U777 ( .C1(n1455), .C2(n2628), .A(n2055), .B(n2632), .ZN(n1871) );
  NAND2_X2 U778 ( .A1(u4_fract_out_pl1_22_), .A2(n2057), .ZN(n2055) );
  AND2_X2 U779 ( .A1(n2049), .A2(n1873), .ZN(N466) );
  OAI211_X2 U780 ( .C1(n2058), .C2(n2627), .A(n2059), .B(n2631), .ZN(n1873) );
  NAND2_X2 U781 ( .A1(u4_fract_out_pl1_21_), .A2(n2057), .ZN(n2059) );
  INV_X4 U783 ( .A(n1872), .ZN(n1924) );
  OAI211_X2 U784 ( .C1(n2060), .C2(n2627), .A(n2061), .B(n2056), .ZN(n1872) );
  NAND2_X2 U785 ( .A1(u4_fract_out_pl1_20_), .A2(n2057), .ZN(n2061) );
  INV_X4 U787 ( .A(n2048), .ZN(n1876) );
  OAI211_X2 U788 ( .C1(n1456), .C2(n2628), .A(n2062), .B(n2632), .ZN(n2048) );
  NAND2_X2 U789 ( .A1(u4_fract_out_pl1_19_), .A2(n2630), .ZN(n2062) );
  INV_X4 U791 ( .A(n2047), .ZN(n1874) );
  OAI211_X2 U792 ( .C1(n1457), .C2(n2628), .A(n2063), .B(n2631), .ZN(n2047) );
  NAND2_X2 U793 ( .A1(u4_fract_out_pl1_18_), .A2(n2630), .ZN(n2063) );
  INV_X4 U795 ( .A(n1921), .ZN(n1875) );
  OAI211_X2 U796 ( .C1(n1458), .C2(n2627), .A(n2064), .B(n2056), .ZN(n1921) );
  NAND2_X2 U797 ( .A1(u4_fract_out_pl1_17_), .A2(n2057), .ZN(n2064) );
  AND2_X2 U798 ( .A1(n2049), .A2(n1864), .ZN(N461) );
  OAI211_X2 U799 ( .C1(n2065), .C2(n2627), .A(n2066), .B(n2632), .ZN(n1864) );
  NAND2_X2 U800 ( .A1(u4_fract_out_pl1_16_), .A2(n2057), .ZN(n2066) );
  AND2_X2 U801 ( .A1(n2049), .A2(n1866), .ZN(N460) );
  OAI211_X2 U802 ( .C1(n2067), .C2(n2628), .A(n2068), .B(n2631), .ZN(n1866) );
  NAND2_X2 U803 ( .A1(u4_fract_out_pl1_15_), .A2(n2057), .ZN(n2068) );
  INV_X4 U805 ( .A(n1865), .ZN(n1922) );
  OAI211_X2 U806 ( .C1(n2069), .C2(n2628), .A(n2070), .B(n2056), .ZN(n1865) );
  NAND2_X2 U807 ( .A1(u4_fract_out_pl1_14_), .A2(n2057), .ZN(n2070) );
  INV_X4 U809 ( .A(n2071), .ZN(n1869) );
  OAI211_X2 U810 ( .C1(n1459), .C2(n2628), .A(n2072), .B(n2632), .ZN(n2071) );
  NAND2_X2 U811 ( .A1(u4_fract_out_pl1_13_), .A2(n2630), .ZN(n2072) );
  INV_X4 U813 ( .A(n2073), .ZN(n1867) );
  OAI211_X2 U814 ( .C1(n1460), .C2(n2627), .A(n2074), .B(n2631), .ZN(n2073) );
  NAND2_X2 U815 ( .A1(u4_fract_out_pl1_12_), .A2(n2057), .ZN(n2074) );
  INV_X4 U817 ( .A(n1918), .ZN(n1868) );
  OAI211_X2 U818 ( .C1(n1461), .C2(n2627), .A(n2075), .B(n2056), .ZN(n1918) );
  NAND2_X2 U819 ( .A1(u4_fract_out_pl1_11_), .A2(n2630), .ZN(n2075) );
  INV_X4 U821 ( .A(n1857), .ZN(n2042) );
  OAI211_X2 U822 ( .C1(n2076), .C2(n2627), .A(n2077), .B(n2632), .ZN(n1857) );
  NAND2_X2 U823 ( .A1(u4_fract_out_pl1_10_), .A2(n2630), .ZN(n2077) );
  INV_X4 U825 ( .A(n1859), .ZN(n2043) );
  OAI211_X2 U826 ( .C1(n1450), .C2(n2627), .A(n2078), .B(n2631), .ZN(n1859) );
  NAND2_X2 U827 ( .A1(u4_fract_out_pl1_9_), .A2(n2630), .ZN(n2078) );
  INV_X4 U829 ( .A(n1858), .ZN(n1919) );
  OAI211_X2 U830 ( .C1(n1451), .C2(n2628), .A(n2079), .B(n2056), .ZN(n1858) );
  NAND2_X2 U831 ( .A1(u4_fract_out_pl1_8_), .A2(n2630), .ZN(n2079) );
  INV_X4 U833 ( .A(n2080), .ZN(n1862) );
  OAI211_X2 U834 ( .C1(n1452), .C2(n2628), .A(n2081), .B(n2632), .ZN(n2080) );
  NAND2_X2 U835 ( .A1(u4_fract_out_pl1_7_), .A2(n2630), .ZN(n2081) );
  INV_X4 U837 ( .A(n2082), .ZN(n1860) );
  OAI211_X2 U838 ( .C1(n2083), .C2(n2627), .A(n2084), .B(n2631), .ZN(n2082) );
  NAND2_X2 U839 ( .A1(u4_fract_out_pl1_6_), .A2(n2057), .ZN(n2084) );
  INV_X4 U841 ( .A(n1913), .ZN(n1861) );
  OAI211_X2 U842 ( .C1(n2085), .C2(n2627), .A(n2086), .B(n2056), .ZN(n1913) );
  NAND2_X2 U843 ( .A1(u4_fract_out_pl1_5_), .A2(n2057), .ZN(n2086) );
  INV_X4 U845 ( .A(n1850), .ZN(n2044) );
  OAI211_X2 U846 ( .C1(n2087), .C2(n2628), .A(n2088), .B(n2632), .ZN(n1850) );
  NAND2_X2 U847 ( .A1(u4_fract_out_pl1_4_), .A2(n2630), .ZN(n2088) );
  INV_X4 U849 ( .A(n1852), .ZN(n2045) );
  OAI211_X2 U850 ( .C1(n1453), .C2(n2628), .A(n2089), .B(n2631), .ZN(n1852) );
  NAND2_X2 U851 ( .A1(u4_fract_out_pl1_3_), .A2(n2630), .ZN(n2089) );
  INV_X4 U853 ( .A(n1851), .ZN(n1916) );
  OAI211_X2 U854 ( .C1(n1454), .C2(n2628), .A(n2090), .B(n2056), .ZN(n1851) );
  NAND2_X2 U855 ( .A1(u4_fract_out_pl1_2_), .A2(n2630), .ZN(n2090) );
  INV_X4 U857 ( .A(n1855), .ZN(n1914) );
  OAI211_X2 U858 ( .C1(n2091), .C2(n2628), .A(n2092), .B(n2632), .ZN(n1855) );
  NAND2_X2 U859 ( .A1(u4_fract_out_pl1_1_), .A2(n2057), .ZN(n2092) );
  OAI22_X2 U860 ( .A1(n1877), .A2(n2049), .B1(n3490), .B2(n1915), .ZN(N445) );
  INV_X4 U861 ( .A(n1853), .ZN(n1915) );
  OAI211_X2 U862 ( .C1(n2093), .C2(n2627), .A(n2094), .B(n2631), .ZN(n1853) );
  NAND2_X2 U868 ( .A1(u4_fract_out_pl1_0_), .A2(n2057), .ZN(n2094) );
  AOI22_X2 U870 ( .A1(n2104), .A2(n2105), .B1(n2106), .B2(rmode_r3[1]), .ZN(
        n2103) );
  INV_X4 U871 ( .A(n2097), .ZN(n2102) );
  OAI221_X2 U873 ( .B1(n2500), .B2(n2106), .C1(r489_B_0_), .C2(n2105), .A(
        n3493), .ZN(n2107) );
  NAND2_X2 U876 ( .A1(n2108), .A2(n2109), .ZN(n1854) );
  NOR4_X2 U877 ( .A1(n1925), .A2(n1926), .A3(n1927), .A4(n1928), .ZN(n2109) );
  NOR4_X2 U882 ( .A1(n1929), .A2(n1930), .A3(n1931), .A4(n1932), .ZN(n2108) );
  NAND2_X2 U883 ( .A1(n2111), .A2(n2116), .ZN(n1932) );
  AND2_X2 U888 ( .A1(n2111), .A2(n2118), .ZN(n2112) );
  NAND2_X2 U889 ( .A1(n2119), .A2(n2123), .ZN(n2118) );
  INV_X4 U890 ( .A(n1956), .ZN(n2123) );
  OAI211_X2 U892 ( .C1(n2126), .C2(n2017), .A(r489_B_0_), .B(n3518), .ZN(n2125) );
  NOR4_X2 U893 ( .A1(n2127), .A2(n2128), .A3(n3353), .A4(n3579), .ZN(n2126) );
  NOR4_X2 U896 ( .A1(exp_ovf_r[1]), .A2(n2133), .A3(n2500), .A4(n2587), .ZN(
        n2132) );
  OAI22_X2 U900 ( .A1(n2138), .A2(n2680), .B1(n2139), .B2(n1444), .ZN(n2134)
         );
  AOI22_X2 U906 ( .A1(n2490), .A2(n2143), .B1(n2144), .B2(n3518), .ZN(n2142)
         );
  OAI211_X2 U910 ( .C1(n2148), .C2(n2149), .A(n3565), .B(n2150), .ZN(n2147) );
  NAND4_X2 U912 ( .A1(n2117), .A2(n2120), .A3(n2121), .A4(n2122), .ZN(n2149)
         );
  NAND2_X2 U913 ( .A1(n2151), .A2(n2152), .ZN(n2121) );
  AOI221_X2 U914 ( .B1(u4_exp_fix_divb[2]), .B2(n2153), .C1(u4_exp_fix_diva[2]), .C2(n2154), .A(n2155), .ZN(n2152) );
  INV_X4 U915 ( .A(n2156), .ZN(n2155) );
  AOI22_X2 U916 ( .A1(u4_exp_next_mi_2_), .A2(n2157), .B1(n2682), .B2(n2158), 
        .ZN(n2156) );
  NAND2_X2 U918 ( .A1(n2162), .A2(n2163), .ZN(n2120) );
  AOI221_X2 U919 ( .B1(u4_exp_fix_divb[1]), .B2(n2153), .C1(u4_exp_fix_diva[1]), .C2(n2154), .A(n2164), .ZN(n2163) );
  INV_X4 U920 ( .A(n2165), .ZN(n2164) );
  AOI22_X2 U921 ( .A1(u4_exp_next_mi_1_), .A2(n2157), .B1(n2681), .B2(n2158), 
        .ZN(n2165) );
  AND2_X2 U923 ( .A1(n2166), .A2(n2167), .ZN(n2117) );
  AOI221_X2 U924 ( .B1(u4_exp_fix_divb[0]), .B2(n2153), .C1(u4_exp_fix_diva[0]), .C2(n2154), .A(n2168), .ZN(n2167) );
  AOI22_X2 U927 ( .A1(rmode_r3[1]), .A2(n2173), .B1(u4_exp_out_mi1[0]), .B2(
        n2160), .ZN(n2170) );
  NAND4_X2 U932 ( .A1(n2110), .A2(n2113), .A3(n2114), .A4(n2115), .ZN(n2148)
         );
  NAND2_X2 U933 ( .A1(n2177), .A2(n2178), .ZN(n2115) );
  AOI221_X2 U934 ( .B1(u4_exp_fix_divb[7]), .B2(n2153), .C1(u4_exp_fix_diva[7]), .C2(n2154), .A(n2179), .ZN(n2178) );
  INV_X4 U935 ( .A(n2180), .ZN(n2179) );
  AOI22_X2 U936 ( .A1(u4_exp_next_mi_7_), .A2(n2157), .B1(n2687), .B2(n2158), 
        .ZN(n2180) );
  NAND2_X2 U938 ( .A1(n2181), .A2(n2182), .ZN(n2114) );
  AOI221_X2 U939 ( .B1(u4_exp_fix_divb[6]), .B2(n2153), .C1(u4_exp_fix_diva[6]), .C2(n2154), .A(n2183), .ZN(n2182) );
  INV_X4 U940 ( .A(n2184), .ZN(n2183) );
  AOI22_X2 U941 ( .A1(u4_exp_next_mi_6_), .A2(n2157), .B1(n2686), .B2(n2158), 
        .ZN(n2184) );
  NAND2_X2 U943 ( .A1(n2185), .A2(n2186), .ZN(n2113) );
  AOI221_X2 U944 ( .B1(u4_exp_fix_divb[5]), .B2(n2153), .C1(u4_exp_fix_diva[5]), .C2(n2154), .A(n2187), .ZN(n2186) );
  INV_X4 U945 ( .A(n2188), .ZN(n2187) );
  AOI22_X2 U946 ( .A1(u4_exp_next_mi_5_), .A2(n2157), .B1(n2685), .B2(n2158), 
        .ZN(n2188) );
  NAND2_X2 U948 ( .A1(n2189), .A2(n2190), .ZN(n2110) );
  AOI221_X2 U949 ( .B1(u4_exp_fix_divb[4]), .B2(n2153), .C1(u4_exp_fix_diva[4]), .C2(n2154), .A(n2191), .ZN(n2190) );
  INV_X4 U950 ( .A(n2192), .ZN(n2191) );
  AOI22_X2 U951 ( .A1(u4_exp_next_mi_4_), .A2(n2157), .B1(n2684), .B2(n2158), 
        .ZN(n2192) );
  AOI22_X2 U956 ( .A1(n2567), .A2(u4_N1284), .B1(u4_N1283), .B2(n3492), .ZN(
        n1389) );
  NAND2_X2 U957 ( .A1(n2017), .A2(n2104), .ZN(n1952) );
  NAND2_X2 U961 ( .A1(n2196), .A2(n2197), .ZN(n2122) );
  AOI221_X2 U962 ( .B1(u4_exp_fix_divb[3]), .B2(n2153), .C1(u4_exp_fix_diva[3]), .C2(n2154), .A(n2198), .ZN(n2197) );
  INV_X4 U963 ( .A(n2199), .ZN(n2198) );
  AOI22_X2 U964 ( .A1(u4_exp_next_mi_3_), .A2(n2157), .B1(n2683), .B2(n2158), 
        .ZN(n2199) );
  OAI22_X2 U971 ( .A1(r489_B_0_), .A2(n2203), .B1(n1395), .B2(n1394), .ZN(
        n2161) );
  NAND2_X2 U973 ( .A1(n2174), .A2(rmode_r3[1]), .ZN(n1394) );
  INV_X4 U975 ( .A(n2176), .ZN(n2204) );
  OAI211_X2 U977 ( .C1(n2625), .C2(n2141), .A(n2201), .B(n1949), .ZN(n2205) );
  INV_X4 U978 ( .A(n2200), .ZN(n2201) );
  NOR4_X2 U979 ( .A1(n2206), .A2(n2128), .A3(n2093), .A4(n2207), .ZN(n2200) );
  NAND2_X2 U980 ( .A1(n2208), .A2(n2209), .ZN(n2128) );
  AND4_X2 U981 ( .A1(n2687), .A2(n2685), .A3(n2684), .A4(n2683), .ZN(n2209) );
  AND4_X2 U982 ( .A1(n2682), .A2(n2681), .A3(n2650), .A4(n2686), .ZN(n2208) );
  INV_X4 U983 ( .A(n2014), .ZN(n2141) );
  NAND4_X2 U985 ( .A1(u4_exp_out_2_), .A2(u4_exp_out_3_), .A3(u4_exp_out_1_), 
        .A4(n2210), .ZN(n2130) );
  AND3_X2 U986 ( .A1(u4_exp_out_4_), .A2(u4_exp_out_6_), .A3(u4_exp_out_5_), 
        .ZN(n2210) );
  INV_X4 U988 ( .A(u4_N1976), .ZN(u4_N1640) );
  INV_X4 U989 ( .A(n2203), .ZN(n2172) );
  NAND2_X2 U990 ( .A1(n2105), .A2(u4_fract_out_pl1_23_), .ZN(n2203) );
  AND2_X2 U992 ( .A1(u4_fract_out_pl1_23_), .A2(n2106), .ZN(n2174) );
  OAI211_X2 U994 ( .C1(n2213), .C2(n1959), .A(n2584), .B(n2625), .ZN(n2212) );
  INV_X4 U995 ( .A(n2002), .ZN(n1959) );
  NOR4_X2 U998 ( .A1(n2217), .A2(n2218), .A3(n2219), .A4(n2220), .ZN(n2216) );
  NAND4_X2 U999 ( .A1(n1555), .A2(n1790), .A3(n1791), .A4(n2221), .ZN(n2220)
         );
  NAND4_X2 U1001 ( .A1(n1789), .A2(n1788), .A3(n1546), .A4(n2223), .ZN(n2219)
         );
  NAND4_X2 U1003 ( .A1(n3535), .A2(n3536), .A3(n1787), .A4(n2226), .ZN(n2218)
         );
  NAND4_X2 U1005 ( .A1(n1497), .A2(n1785), .A3(n1786), .A4(n2228), .ZN(n2217)
         );
  AND4_X2 U1008 ( .A1(u4_N1977), .A2(n2232), .A3(n2007), .A4(n2465), .ZN(n2231) );
  OAI211_X2 U1010 ( .C1(n2236), .C2(n2237), .A(n1386), .B(exp_ovf_r[1]), .ZN(
        n2235) );
  NAND4_X2 U1012 ( .A1(n2238), .A2(n2239), .A3(n2240), .A4(n2241), .ZN(n2000)
         );
  NOR4_X2 U1013 ( .A1(n2242), .A2(u4_fract_out_4_), .A3(u4_fract_out_6_), .A4(
        u4_fract_out_5_), .ZN(n2241) );
  INV_X4 U1014 ( .A(n2085), .ZN(u4_fract_out_5_) );
  AOI22_X2 U1015 ( .A1(u4_N1388), .A2(n2243), .B1(u4_N1438), .B2(n2244), .ZN(
        n2085) );
  INV_X4 U1016 ( .A(n2083), .ZN(u4_fract_out_6_) );
  AOI22_X2 U1017 ( .A1(u4_N1389), .A2(n2243), .B1(u4_N1439), .B2(n2244), .ZN(
        n2083) );
  INV_X4 U1018 ( .A(n2087), .ZN(u4_fract_out_4_) );
  AOI22_X2 U1019 ( .A1(u4_N1387), .A2(n2243), .B1(u4_N1437), .B2(n2646), .ZN(
        n2087) );
  AOI22_X2 U1021 ( .A1(u4_N1390), .A2(n2243), .B1(u4_N1440), .B2(n2244), .ZN(
        n1452) );
  AOI22_X2 U1022 ( .A1(u4_N1392), .A2(n2243), .B1(u4_N1442), .B2(n2244), .ZN(
        n1450) );
  AOI22_X2 U1023 ( .A1(u4_N1391), .A2(n2243), .B1(u4_N1441), .B2(n2244), .ZN(
        n1451) );
  NOR4_X2 U1024 ( .A1(n2245), .A2(u4_fract_out_1_), .A3(u4_fract_out_21_), 
        .A4(u4_fract_out_20_), .ZN(n2240) );
  INV_X4 U1025 ( .A(n2060), .ZN(u4_fract_out_20_) );
  AOI22_X2 U1026 ( .A1(u4_N1403), .A2(n2243), .B1(u4_N1453), .B2(n2244), .ZN(
        n2060) );
  INV_X4 U1027 ( .A(n2058), .ZN(u4_fract_out_21_) );
  AOI22_X2 U1028 ( .A1(u4_N1404), .A2(n2243), .B1(u4_N1454), .B2(n2244), .ZN(
        n2058) );
  INV_X4 U1029 ( .A(n2091), .ZN(u4_fract_out_1_) );
  AOI22_X2 U1030 ( .A1(u4_N1384), .A2(n2243), .B1(u4_N1434), .B2(n2646), .ZN(
        n2091) );
  AOI22_X2 U1032 ( .A1(u4_N1405), .A2(n2243), .B1(u4_N1455), .B2(n2244), .ZN(
        n1455) );
  AOI22_X2 U1033 ( .A1(u4_N1386), .A2(n2243), .B1(u4_N1436), .B2(n2646), .ZN(
        n1453) );
  AOI22_X2 U1034 ( .A1(u4_N1385), .A2(n2243), .B1(u4_N1435), .B2(n2646), .ZN(
        n1454) );
  NOR4_X2 U1035 ( .A1(n2246), .A2(u4_fract_out_14_), .A3(u4_fract_out_16_), 
        .A4(u4_fract_out_15_), .ZN(n2239) );
  INV_X4 U1036 ( .A(n2067), .ZN(u4_fract_out_15_) );
  AOI22_X2 U1037 ( .A1(u4_N1398), .A2(n2243), .B1(u4_N1448), .B2(n2646), .ZN(
        n2067) );
  INV_X4 U1038 ( .A(n2065), .ZN(u4_fract_out_16_) );
  AOI22_X2 U1039 ( .A1(u4_N1399), .A2(n2243), .B1(u4_N1449), .B2(n2646), .ZN(
        n2065) );
  INV_X4 U1040 ( .A(n2069), .ZN(u4_fract_out_14_) );
  AOI22_X2 U1041 ( .A1(u4_N1397), .A2(n2243), .B1(u4_N1447), .B2(n2646), .ZN(
        n2069) );
  AOI22_X2 U1043 ( .A1(u4_N1400), .A2(n2243), .B1(u4_N1450), .B2(n2646), .ZN(
        n1458) );
  AOI22_X2 U1044 ( .A1(u4_N1402), .A2(n2243), .B1(u4_N1452), .B2(n2646), .ZN(
        n1456) );
  AOI22_X2 U1045 ( .A1(u4_N1401), .A2(n2243), .B1(u4_N1451), .B2(n2646), .ZN(
        n1457) );
  INV_X4 U1047 ( .A(n2093), .ZN(u4_fract_out_0_) );
  INV_X4 U1048 ( .A(n2076), .ZN(u4_fract_out_10_) );
  AOI22_X2 U1049 ( .A1(u4_N1393), .A2(n2243), .B1(u4_N1443), .B2(n2646), .ZN(
        n2076) );
  AOI22_X2 U1051 ( .A1(u4_N1394), .A2(n2243), .B1(u4_N1444), .B2(n2646), .ZN(
        n1461) );
  AOI22_X2 U1052 ( .A1(u4_N1396), .A2(n2243), .B1(u4_N1446), .B2(n2646), .ZN(
        n1459) );
  AOI22_X2 U1053 ( .A1(u4_N1395), .A2(n2243), .B1(u4_N1445), .B2(n2646), .ZN(
        n1460) );
  INV_X4 U1054 ( .A(n2233), .ZN(n2236) );
  OAI22_X2 U1057 ( .A1(exp_ovf_r[0]), .A2(n3442), .B1(exp_ovf_r[1]), .B2(n2137), .ZN(n2248) );
  NAND4_X2 U1058 ( .A1(n2687), .A2(n2473), .A3(n2249), .A4(n2250), .ZN(n2137)
         );
  NOR4_X2 U1059 ( .A1(n2686), .A2(n2685), .A3(n2684), .A4(n2683), .ZN(n2250)
         );
  NAND2_X2 U1062 ( .A1(n2207), .A2(n2206), .ZN(n2007) );
  NAND2_X2 U1063 ( .A1(n2251), .A2(n2214), .ZN(n2206) );
  NAND4_X2 U1064 ( .A1(u4_N1290), .A2(n1543), .A3(n2252), .A4(n2253), .ZN(
        n2251) );
  NOR4_X2 U1065 ( .A1(n2254), .A2(fract_denorm[39]), .A3(fract_denorm[41]), 
        .A4(fract_denorm[40]), .ZN(n2253) );
  OR3_X2 U1066 ( .A1(fract_denorm[23]), .A2(fract_denorm[31]), .A3(n2493), 
        .ZN(n2254) );
  NAND4_X2 U1071 ( .A1(n2260), .A2(n2261), .A3(n2262), .A4(n2263), .ZN(n2259)
         );
  NAND4_X2 U1076 ( .A1(n2264), .A2(n2265), .A3(n2266), .A4(n2267), .ZN(n2258)
         );
  NAND4_X2 U1082 ( .A1(n2270), .A2(n2271), .A3(n2272), .A4(n2273), .ZN(n2269)
         );
  NAND4_X2 U1087 ( .A1(n2274), .A2(n2275), .A3(n2276), .A4(n2277), .ZN(n2268)
         );
  INV_X4 U1092 ( .A(n2278), .ZN(n2214) );
  AOI22_X2 U1093 ( .A1(u4_N1382), .A2(n2243), .B1(u4_N1432), .B2(n2646), .ZN(
        n2278) );
  OR4_X2 U1094 ( .A1(n2279), .A2(n2280), .A3(n2281), .A4(n2282), .ZN(n1966) );
  NAND4_X2 U1095 ( .A1(n2283), .A2(n2284), .A3(n2285), .A4(n2286), .ZN(n2282)
         );
  NAND4_X2 U1100 ( .A1(n2287), .A2(n2288), .A3(n2289), .A4(n2290), .ZN(n2281)
         );
  NOR4_X2 U1101 ( .A1(remainder[9]), .A2(remainder[8]), .A3(remainder[7]), 
        .A4(remainder[6]), .ZN(n2290) );
  NAND4_X2 U1105 ( .A1(n2291), .A2(n2292), .A3(n2293), .A4(n2294), .ZN(n2280)
         );
  NAND4_X2 U1110 ( .A1(n2295), .A2(n2296), .A3(n2297), .A4(n2298), .ZN(n2279)
         );
  NOR4_X2 U1111 ( .A1(remainder[31]), .A2(remainder[30]), .A3(remainder[2]), 
        .A4(remainder[29]), .ZN(n2298) );
  AOI22_X2 U1117 ( .A1(u4_N1383), .A2(n2243), .B1(u4_N1433), .B2(n2244), .ZN(
        n2093) );
  INV_X4 U1118 ( .A(n2256), .ZN(n2244) );
  OAI211_X2 U1119 ( .C1(n1970), .C2(n2299), .A(n2300), .B(n2301), .ZN(n2256)
         );
  OR3_X2 U1122 ( .A1(n1439), .A2(n3583), .A3(n1438), .ZN(n2305) );
  NAND2_X2 U1125 ( .A1(n2232), .A2(n2306), .ZN(n2008) );
  NAND2_X2 U1130 ( .A1(n3442), .A2(u4_N1733), .ZN(n2003) );
  NAND2_X2 U1132 ( .A1(u4_exp_in_pl1_8_), .A2(n2679), .ZN(n2307) );
  OR2_X2 U1133 ( .A1(u4_exp_in_pl1_7_), .A2(u4_exp_in_pl1_6_), .ZN(n2304) );
  OR2_X2 U1134 ( .A1(u4_div_scht1a[6]), .A2(u4_div_scht1a[7]), .ZN(n2303) );
  INV_X4 U1136 ( .A(n2308), .ZN(n1443) );
  OAI22_X2 U1137 ( .A1(u4_N1733), .A2(n2493), .B1(exp_ovf_r[0]), .B2(n1996), 
        .ZN(n2308) );
  NAND2_X2 U1138 ( .A1(n3565), .A2(n1962), .ZN(n1996) );
  INV_X4 U1139 ( .A(u4_N1733), .ZN(n1962) );
  OR3_X2 U1140 ( .A1(u4_f2i_shft_7_), .A2(u4_f2i_shft_6_), .A3(n3488), .ZN(
        n2302) );
  AOI22_X2 U1141 ( .A1(opas_r2), .A2(u4_N1284), .B1(n2193), .B2(u4_N1283), 
        .ZN(n1388) );
  NAND4_X2 U1142 ( .A1(rmode_r3[1]), .A2(rmode_r3[0]), .A3(opas_r2), .A4(n1386), .ZN(n2193) );
  NAND2_X2 U1143 ( .A1(n1466), .A2(n1791), .ZN(n1386) );
  AOI221_X2 U1144 ( .B1(n2644), .B2(quo[2]), .C1(n2621), .C2(prod[0]), .A(
        n2311), .ZN(n1791) );
  AND2_X2 U1145 ( .A1(fract_i2f[0]), .A2(n2690), .ZN(n2311) );
  AND3_X2 U1146 ( .A1(n2224), .A2(n1558), .A3(n1534), .ZN(n1466) );
  AND2_X2 U1147 ( .A1(n1557), .A2(n2227), .ZN(n1534) );
  AOI221_X2 U1148 ( .B1(n2643), .B2(quo[5]), .C1(n2622), .C2(prod[3]), .A(
        n2312), .ZN(n2227) );
  AND2_X2 U1149 ( .A1(fract_i2f[3]), .A2(n2690), .ZN(n2312) );
  AND3_X2 U1150 ( .A1(n1786), .A2(n1497), .A3(n1498), .ZN(n1557) );
  AND2_X2 U1151 ( .A1(n1535), .A2(n1785), .ZN(n1498) );
  AOI221_X2 U1152 ( .B1(n2643), .B2(quo[8]), .C1(n2621), .C2(prod[6]), .A(
        n2313), .ZN(n1785) );
  AND2_X2 U1153 ( .A1(fract_i2f[6]), .A2(n2690), .ZN(n2313) );
  AND2_X2 U1156 ( .A1(n1559), .A2(n1790), .ZN(n1513) );
  AOI221_X2 U1157 ( .B1(n2643), .B2(quo[13]), .C1(n2621), .C2(prod[11]), .A(
        n2314), .ZN(n1790) );
  AND2_X2 U1158 ( .A1(fract_i2f[11]), .A2(n2690), .ZN(n2314) );
  AND3_X2 U1159 ( .A1(n2222), .A2(n1507), .A3(n1508), .ZN(n1559) );
  AOI221_X2 U1161 ( .B1(n2643), .B2(quo[16]), .C1(n2623), .C2(prod[14]), .A(
        n2315), .ZN(n1514) );
  AND2_X2 U1162 ( .A1(fract_i2f[14]), .A2(n2690), .ZN(n2315) );
  NAND2_X2 U1164 ( .A1(n1556), .A2(n1788), .ZN(n1420) );
  AOI221_X2 U1165 ( .B1(n2643), .B2(quo[19]), .C1(n2621), .C2(prod[17]), .A(
        n2316), .ZN(n1788) );
  AND2_X2 U1166 ( .A1(fract_i2f[17]), .A2(n2690), .ZN(n2316) );
  AND3_X2 U1167 ( .A1(n2225), .A2(n1532), .A3(n1533), .ZN(n1556) );
  AND2_X2 U1168 ( .A1(n1494), .A2(n1787), .ZN(n1533) );
  AOI221_X2 U1169 ( .B1(n2643), .B2(quo[22]), .C1(n2623), .C2(prod[20]), .A(
        n3558), .ZN(n1787) );
  AOI22_X2 U1170 ( .A1(fract_out_q[0]), .A2(n1942), .B1(fract_i2f[20]), .B2(
        n2690), .ZN(n2317) );
  OR3_X2 U1177 ( .A1(fract_denorm[43]), .A2(fract_denorm[44]), .A3(
        fract_denorm[42]), .ZN(n1506) );
  OAI211_X2 U1178 ( .C1(n2533), .C2(n2464), .A(n2318), .B(n2319), .ZN(
        fract_denorm[42]) );
  AOI22_X2 U1179 ( .A1(fract_out_q[22]), .A2(n1942), .B1(fract_i2f[42]), .B2(
        n2690), .ZN(n2319) );
  AOI22_X2 U1180 ( .A1(quo[21]), .A2(n2320), .B1(quo[44]), .B2(n2309), .ZN(
        n2318) );
  OAI211_X2 U1181 ( .C1(n2533), .C2(n2484), .A(n2321), .B(n2322), .ZN(
        fract_denorm[44]) );
  AOI22_X2 U1182 ( .A1(fract_out_q[24]), .A2(n1942), .B1(fract_i2f[44]), .B2(
        n2690), .ZN(n2322) );
  AOI22_X2 U1183 ( .A1(quo[23]), .A2(n2320), .B1(quo[46]), .B2(n2309), .ZN(
        n2321) );
  OAI211_X2 U1184 ( .C1(n2533), .C2(n2534), .A(n2323), .B(n2324), .ZN(
        fract_denorm[43]) );
  AOI22_X2 U1185 ( .A1(fract_out_q[23]), .A2(n1942), .B1(fract_i2f[43]), .B2(
        n2690), .ZN(n2324) );
  AOI22_X2 U1186 ( .A1(quo[22]), .A2(n2320), .B1(quo[45]), .B2(n2309), .ZN(
        n2323) );
  OAI211_X2 U1187 ( .C1(n2638), .C2(n2539), .A(n2325), .B(n2326), .ZN(
        fract_denorm[46]) );
  AOI22_X2 U1188 ( .A1(fract_out_q[26]), .A2(n1942), .B1(fract_i2f[46]), .B2(
        n2690), .ZN(n2326) );
  OAI211_X2 U1190 ( .C1(n2638), .C2(n2541), .A(n2327), .B(n2328), .ZN(
        fract_denorm[45]) );
  AOI22_X2 U1191 ( .A1(fract_out_q[25]), .A2(n1942), .B1(fract_i2f[45]), .B2(
        n2690), .ZN(n2328) );
  OAI211_X2 U1193 ( .C1(n2638), .C2(n2542), .A(n2329), .B(n2330), .ZN(
        fract_denorm[41]) );
  AOI22_X2 U1194 ( .A1(fract_out_q[21]), .A2(n1942), .B1(fract_i2f[41]), .B2(
        n2690), .ZN(n2330) );
  AOI22_X2 U1195 ( .A1(quo[20]), .A2(n2320), .B1(quo[43]), .B2(n2644), .ZN(
        n2329) );
  OAI211_X2 U1196 ( .C1(n2638), .C2(n2555), .A(n2331), .B(n2332), .ZN(
        fract_denorm[40]) );
  AOI22_X2 U1197 ( .A1(fract_out_q[20]), .A2(n1942), .B1(fract_i2f[40]), .B2(
        n2690), .ZN(n2332) );
  AOI22_X2 U1198 ( .A1(quo[19]), .A2(n2320), .B1(quo[42]), .B2(n2644), .ZN(
        n2331) );
  OAI211_X2 U1199 ( .C1(n2638), .C2(n2552), .A(n2333), .B(n2334), .ZN(
        fract_denorm[39]) );
  AOI22_X2 U1200 ( .A1(fract_out_q[19]), .A2(n1942), .B1(fract_i2f[39]), .B2(
        n2690), .ZN(n2334) );
  AOI22_X2 U1201 ( .A1(quo[18]), .A2(n2320), .B1(quo[41]), .B2(n2644), .ZN(
        n2333) );
  OAI211_X2 U1202 ( .C1(n2638), .C2(n2554), .A(n2335), .B(n2336), .ZN(
        fract_denorm[31]) );
  AOI22_X2 U1203 ( .A1(fract_out_q[11]), .A2(n1942), .B1(fract_i2f[31]), .B2(
        n2690), .ZN(n2336) );
  AOI22_X2 U1204 ( .A1(quo[10]), .A2(n2320), .B1(quo[33]), .B2(n2643), .ZN(
        n2335) );
  OAI211_X2 U1208 ( .C1(n2638), .C2(n2483), .A(n2337), .B(n2338), .ZN(
        fract_denorm[36]) );
  AOI22_X2 U1209 ( .A1(fract_out_q[16]), .A2(n1942), .B1(fract_i2f[36]), .B2(
        n2690), .ZN(n2338) );
  AOI22_X2 U1210 ( .A1(quo[15]), .A2(n2320), .B1(quo[38]), .B2(n2644), .ZN(
        n2337) );
  OAI211_X2 U1211 ( .C1(n2638), .C2(n2538), .A(n2339), .B(n2340), .ZN(
        fract_denorm[38]) );
  AOI22_X2 U1212 ( .A1(fract_out_q[18]), .A2(n1942), .B1(fract_i2f[38]), .B2(
        n2690), .ZN(n2340) );
  AOI22_X2 U1213 ( .A1(quo[17]), .A2(n2320), .B1(quo[40]), .B2(n2643), .ZN(
        n2339) );
  OAI211_X2 U1214 ( .C1(n2638), .C2(n2540), .A(n2341), .B(n2342), .ZN(
        fract_denorm[37]) );
  AOI22_X2 U1215 ( .A1(fract_out_q[17]), .A2(n1942), .B1(fract_i2f[37]), .B2(
        n2690), .ZN(n2342) );
  AOI22_X2 U1216 ( .A1(quo[16]), .A2(n2320), .B1(quo[39]), .B2(n2644), .ZN(
        n2341) );
  OAI211_X2 U1217 ( .C1(n2638), .C2(n2544), .A(n2343), .B(n2344), .ZN(
        fract_denorm[35]) );
  AOI22_X2 U1218 ( .A1(fract_out_q[15]), .A2(n1942), .B1(fract_i2f[35]), .B2(
        n2690), .ZN(n2344) );
  AOI22_X2 U1219 ( .A1(quo[14]), .A2(n2320), .B1(quo[37]), .B2(n2644), .ZN(
        n2343) );
  OAI211_X2 U1220 ( .C1(n2638), .C2(n2471), .A(n2345), .B(n2346), .ZN(
        fract_denorm[34]) );
  AOI22_X2 U1221 ( .A1(fract_out_q[14]), .A2(n1942), .B1(fract_i2f[34]), .B2(
        n2690), .ZN(n2346) );
  AOI22_X2 U1222 ( .A1(quo[13]), .A2(n2320), .B1(quo[36]), .B2(n2644), .ZN(
        n2345) );
  OAI211_X2 U1223 ( .C1(n2638), .C2(n2551), .A(n2347), .B(n2348), .ZN(
        fract_denorm[33]) );
  AOI22_X2 U1224 ( .A1(fract_out_q[13]), .A2(n1942), .B1(fract_i2f[33]), .B2(
        n2690), .ZN(n2348) );
  AOI22_X2 U1225 ( .A1(quo[12]), .A2(n2320), .B1(quo[35]), .B2(n2644), .ZN(
        n2347) );
  OAI211_X2 U1226 ( .C1(n2638), .C2(n2548), .A(n2349), .B(n2350), .ZN(
        fract_denorm[32]) );
  AOI22_X2 U1227 ( .A1(fract_out_q[12]), .A2(n1942), .B1(fract_i2f[32]), .B2(
        n2690), .ZN(n2350) );
  AOI22_X2 U1228 ( .A1(quo[11]), .A2(n2320), .B1(quo[34]), .B2(n2644), .ZN(
        n2349) );
  OAI211_X2 U1229 ( .C1(n2638), .C2(n2472), .A(n2351), .B(n2352), .ZN(
        fract_denorm[23]) );
  AOI22_X2 U1230 ( .A1(fract_out_q[3]), .A2(n1942), .B1(fract_i2f[23]), .B2(
        n2690), .ZN(n2352) );
  OAI211_X2 U1235 ( .C1(n2638), .C2(n2550), .A(n2353), .B(n2354), .ZN(
        fract_denorm[28]) );
  AOI22_X2 U1236 ( .A1(fract_out_q[8]), .A2(n1942), .B1(fract_i2f[28]), .B2(
        n2690), .ZN(n2354) );
  AOI22_X2 U1237 ( .A1(quo[7]), .A2(n2320), .B1(quo[30]), .B2(n2644), .ZN(
        n2353) );
  OAI211_X2 U1238 ( .C1(n2638), .C2(n2557), .A(n2355), .B(n2356), .ZN(
        fract_denorm[30]) );
  AOI22_X2 U1239 ( .A1(fract_out_q[10]), .A2(n1942), .B1(fract_i2f[30]), .B2(
        n2690), .ZN(n2356) );
  AOI22_X2 U1240 ( .A1(quo[9]), .A2(n2320), .B1(quo[32]), .B2(n2644), .ZN(
        n2355) );
  OAI211_X2 U1241 ( .C1(n2638), .C2(n2556), .A(n2357), .B(n2358), .ZN(
        fract_denorm[29]) );
  AOI22_X2 U1242 ( .A1(fract_out_q[9]), .A2(n1942), .B1(fract_i2f[29]), .B2(
        n2690), .ZN(n2358) );
  AOI22_X2 U1243 ( .A1(quo[8]), .A2(n2320), .B1(quo[31]), .B2(n2644), .ZN(
        n2357) );
  OAI211_X2 U1244 ( .C1(n2638), .C2(n2547), .A(n2359), .B(n2360), .ZN(
        fract_denorm[27]) );
  AOI22_X2 U1245 ( .A1(fract_out_q[7]), .A2(n1942), .B1(fract_i2f[27]), .B2(
        n2690), .ZN(n2360) );
  AOI22_X2 U1246 ( .A1(quo[6]), .A2(n2320), .B1(quo[29]), .B2(n2644), .ZN(
        n2359) );
  OAI211_X2 U1247 ( .C1(n2638), .C2(n2553), .A(n2361), .B(n2362), .ZN(
        fract_denorm[26]) );
  AOI22_X2 U1248 ( .A1(fract_out_q[6]), .A2(n1942), .B1(fract_i2f[26]), .B2(
        n2690), .ZN(n2362) );
  AOI22_X2 U1249 ( .A1(quo[5]), .A2(n2320), .B1(quo[28]), .B2(n2644), .ZN(
        n2361) );
  OAI211_X2 U1250 ( .C1(n2638), .C2(n2485), .A(n2363), .B(n2364), .ZN(
        fract_denorm[25]) );
  AOI22_X2 U1251 ( .A1(fract_out_q[5]), .A2(n1942), .B1(fract_i2f[25]), .B2(
        n2690), .ZN(n2364) );
  AOI22_X2 U1252 ( .A1(quo[4]), .A2(n2320), .B1(quo[27]), .B2(n2644), .ZN(
        n2363) );
  OAI211_X2 U1253 ( .C1(n2638), .C2(n2545), .A(n2365), .B(n2366), .ZN(
        fract_denorm[24]) );
  AOI22_X2 U1254 ( .A1(fract_out_q[4]), .A2(n1942), .B1(fract_i2f[24]), .B2(
        n2690), .ZN(n2366) );
  AOI22_X2 U1255 ( .A1(quo[3]), .A2(n2320), .B1(quo[26]), .B2(n2644), .ZN(
        n2365) );
  OAI211_X2 U1256 ( .C1(n2638), .C2(n2549), .A(n2367), .B(n2368), .ZN(
        fract_denorm[22]) );
  AOI22_X2 U1257 ( .A1(fract_out_q[2]), .A2(n1942), .B1(fract_i2f[22]), .B2(
        n2690), .ZN(n2368) );
  OAI211_X2 U1259 ( .C1(n2638), .C2(n2546), .A(n2369), .B(n2370), .ZN(
        fract_denorm[21]) );
  AOI22_X2 U1260 ( .A1(fract_out_q[1]), .A2(n1942), .B1(fract_i2f[21]), .B2(
        n2690), .ZN(n2370) );
  AOI22_X2 U1262 ( .A1(quo[0]), .A2(n2320), .B1(quo[23]), .B2(n2644), .ZN(
        n2369) );
  AOI221_X2 U1264 ( .B1(n2643), .B2(quo[21]), .C1(n2621), .C2(prod[19]), .A(
        n2371), .ZN(n1532) );
  AND2_X2 U1265 ( .A1(fract_i2f[19]), .A2(n2690), .ZN(n2371) );
  AOI221_X2 U1266 ( .B1(n2643), .B2(quo[20]), .C1(n2622), .C2(prod[18]), .A(
        n2372), .ZN(n2225) );
  AND2_X2 U1267 ( .A1(fract_i2f[18]), .A2(n2690), .ZN(n2372) );
  AOI221_X2 U1268 ( .B1(n2643), .B2(quo[18]), .C1(n2622), .C2(prod[16]), .A(
        n2373), .ZN(n1789) );
  AND2_X2 U1269 ( .A1(fract_i2f[16]), .A2(n2690), .ZN(n2373) );
  AOI221_X2 U1270 ( .B1(n2644), .B2(quo[17]), .C1(n2621), .C2(prod[15]), .A(
        n2374), .ZN(n1546) );
  AND2_X2 U1271 ( .A1(fract_i2f[15]), .A2(n2690), .ZN(n2374) );
  AOI221_X2 U1272 ( .B1(n2644), .B2(quo[15]), .C1(n2623), .C2(prod[13]), .A(
        n2375), .ZN(n1507) );
  AND2_X2 U1273 ( .A1(fract_i2f[13]), .A2(n2690), .ZN(n2375) );
  AOI221_X2 U1274 ( .B1(n2644), .B2(quo[14]), .C1(n2621), .C2(prod[12]), .A(
        n2376), .ZN(n2222) );
  AND2_X2 U1275 ( .A1(fract_i2f[12]), .A2(n2690), .ZN(n2376) );
  AOI221_X2 U1276 ( .B1(n2644), .B2(quo[11]), .C1(n2621), .C2(prod[9]), .A(
        n2377), .ZN(n2229) );
  AND2_X2 U1277 ( .A1(fract_i2f[9]), .A2(n2690), .ZN(n2377) );
  AOI221_X2 U1278 ( .B1(n2644), .B2(quo[12]), .C1(n2623), .C2(prod[10]), .A(
        n2378), .ZN(n1555) );
  AND2_X2 U1279 ( .A1(fract_i2f[10]), .A2(n2690), .ZN(n2378) );
  AOI221_X2 U1280 ( .B1(n2644), .B2(quo[10]), .C1(n2622), .C2(prod[8]), .A(
        n2379), .ZN(n1477) );
  AND2_X2 U1281 ( .A1(fract_i2f[8]), .A2(n2690), .ZN(n2379) );
  AOI221_X2 U1282 ( .B1(n2644), .B2(quo[9]), .C1(n2621), .C2(prod[7]), .A(
        n2380), .ZN(n1541) );
  AND2_X2 U1283 ( .A1(fract_i2f[7]), .A2(n2690), .ZN(n2380) );
  AOI221_X2 U1284 ( .B1(n2644), .B2(quo[7]), .C1(n2622), .C2(prod[5]), .A(
        n2381), .ZN(n1497) );
  AND2_X2 U1285 ( .A1(fract_i2f[5]), .A2(n2690), .ZN(n2381) );
  AOI221_X2 U1286 ( .B1(n2644), .B2(quo[6]), .C1(n2621), .C2(prod[4]), .A(
        n2382), .ZN(n1786) );
  AND2_X2 U1287 ( .A1(fract_i2f[4]), .A2(n2690), .ZN(n2382) );
  AOI221_X2 U1288 ( .B1(n2644), .B2(quo[4]), .C1(n2621), .C2(prod[2]), .A(
        n2383), .ZN(n1558) );
  AND2_X2 U1289 ( .A1(fract_i2f[2]), .A2(n2690), .ZN(n2383) );
  AOI221_X2 U1290 ( .B1(n2643), .B2(quo[3]), .C1(n2623), .C2(prod[1]), .A(
        n2384), .ZN(n2224) );
  AND2_X2 U1291 ( .A1(fract_i2f[1]), .A2(n2690), .ZN(n2384) );
  INV_X4 U1293 ( .A(n1424), .ZN(n2299) );
  INV_X4 U1295 ( .A(n1969), .ZN(n1449) );
  NAND4_X2 U1303 ( .A1(n2473), .A2(n2486), .A3(n1970), .A4(n2387), .ZN(n1444)
         );
  NOR4_X2 U1304 ( .A1(n2685), .A2(n2684), .A3(n2683), .A4(n2682), .ZN(n2387)
         );
  OAI211_X2 U1311 ( .C1(n2649), .C2(n2503), .A(n1829), .B(n2389), .ZN(n2388)
         );
  AND2_X2 U1316 ( .A1(opb_00), .A2(n2490), .ZN(n1838) );
  AOI22_X2 U1322 ( .A1(opb_00), .A2(opa_inf), .B1(opb_inf), .B2(opa_00), .ZN(
        n1948) );
  NAND2_X2 U1326 ( .A1(opa_00), .A2(opb_00), .ZN(n1835) );
  NAND2_X2 U1328 ( .A1(fpu_op_r3[1]), .A2(fpu_op_r3[0]), .ZN(n1937) );
  XNOR2_X2 U1329 ( .A(n1727), .B(n3497), .ZN(N441) );
  NAND2_X2 U1330 ( .A1(rmode_r2[1]), .A2(rmode_r2[0]), .ZN(n1727) );
  OAI221_X2 U1331 ( .B1(n2469), .B2(n2512), .C1(n2636), .C2(n3371), .A(n2393), 
        .ZN(N421) );
  OAI221_X2 U1332 ( .B1(n2469), .B2(n2513), .C1(n2637), .C2(n3372), .A(n2620), 
        .ZN(N420) );
  OAI221_X2 U1333 ( .B1(n2469), .B2(n2508), .C1(n2636), .C2(n3373), .A(n2393), 
        .ZN(N419) );
  OAI221_X2 U1334 ( .B1(n2469), .B2(n2506), .C1(n2637), .C2(n3374), .A(n2620), 
        .ZN(N418) );
  OAI221_X2 U1335 ( .B1(n2469), .B2(n2509), .C1(n2636), .C2(n3375), .A(n2393), 
        .ZN(N417) );
  OAI221_X2 U1336 ( .B1(n2469), .B2(n2510), .C1(n2637), .C2(n3376), .A(n2620), 
        .ZN(N416) );
  OAI221_X2 U1337 ( .B1(n2469), .B2(n2507), .C1(n2636), .C2(n3377), .A(n2393), 
        .ZN(N415) );
  OAI221_X2 U1338 ( .B1(n2469), .B2(n2505), .C1(n2637), .C2(n3378), .A(n2620), 
        .ZN(N414) );
  OAI221_X2 U1339 ( .B1(n2469), .B2(n2529), .C1(n2637), .C2(n3379), .A(n2393), 
        .ZN(N413) );
  OAI221_X2 U1340 ( .B1(n2469), .B2(n2528), .C1(n2637), .C2(n3380), .A(n2620), 
        .ZN(N412) );
  OAI221_X2 U1341 ( .B1(n2469), .B2(n2527), .C1(n2637), .C2(n3381), .A(n2393), 
        .ZN(N411) );
  OAI221_X2 U1342 ( .B1(n2469), .B2(n2611), .C1(n2636), .C2(n3382), .A(n2620), 
        .ZN(N410) );
  OAI221_X2 U1343 ( .B1(n2469), .B2(n2610), .C1(n2636), .C2(n3383), .A(n2393), 
        .ZN(N409) );
  OAI221_X2 U1344 ( .B1(n2469), .B2(n2609), .C1(n2636), .C2(n3384), .A(n2620), 
        .ZN(N408) );
  OAI221_X2 U1345 ( .B1(n2469), .B2(n2608), .C1(n2636), .C2(n3385), .A(n2393), 
        .ZN(N407) );
  OAI221_X2 U1346 ( .B1(n2469), .B2(n2526), .C1(n2636), .C2(n3386), .A(n2620), 
        .ZN(N406) );
  OAI221_X2 U1347 ( .B1(n2469), .B2(n2525), .C1(n2636), .C2(n3387), .A(n2393), 
        .ZN(N405) );
  OAI221_X2 U1348 ( .B1(n2469), .B2(n2524), .C1(n2636), .C2(n3388), .A(n2620), 
        .ZN(N404) );
  OAI221_X2 U1349 ( .B1(n2469), .B2(n2523), .C1(n2636), .C2(n3389), .A(n2393), 
        .ZN(N403) );
  OAI221_X2 U1350 ( .B1(n2469), .B2(n2522), .C1(n2636), .C2(n3390), .A(n2620), 
        .ZN(N402) );
  OAI221_X2 U1351 ( .B1(n2469), .B2(n2521), .C1(n2636), .C2(n3391), .A(n2393), 
        .ZN(N401) );
  OAI221_X2 U1352 ( .B1(n2469), .B2(n2520), .C1(n2636), .C2(n3392), .A(n2620), 
        .ZN(N400) );
  OAI221_X2 U1353 ( .B1(n2469), .B2(n2519), .C1(n2637), .C2(n3393), .A(n2393), 
        .ZN(N399) );
  OAI221_X2 U1354 ( .B1(n2469), .B2(n2518), .C1(n2637), .C2(n3394), .A(n2620), 
        .ZN(N398) );
  OAI221_X2 U1356 ( .B1(n2469), .B2(n2517), .C1(n2637), .C2(n3395), .A(n2395), 
        .ZN(N397) );
  AOI22_X2 U1357 ( .A1(n2641), .A2(N224), .B1(N250), .B2(n2397), .ZN(n2395) );
  OAI221_X2 U1358 ( .B1(n2469), .B2(n2516), .C1(n2637), .C2(n3396), .A(n2398), 
        .ZN(N396) );
  AOI22_X2 U1359 ( .A1(n2642), .A2(opa_r1[22]), .B1(N249), .B2(n2397), .ZN(
        n2398) );
  OAI221_X2 U1360 ( .B1(n2469), .B2(n2515), .C1(n2637), .C2(n3397), .A(n2399), 
        .ZN(N395) );
  AOI22_X2 U1361 ( .A1(n2642), .A2(opa_r1[21]), .B1(N248), .B2(n2397), .ZN(
        n2399) );
  OAI221_X2 U1362 ( .B1(n2469), .B2(n2514), .C1(n2637), .C2(n3398), .A(n2400), 
        .ZN(N394) );
  AOI22_X2 U1363 ( .A1(n2642), .A2(opa_r1[20]), .B1(N247), .B2(n2397), .ZN(
        n2400) );
  OAI221_X2 U1364 ( .B1(n2469), .B2(n2607), .C1(n2637), .C2(n2504), .A(n2401), 
        .ZN(N393) );
  AOI22_X2 U1365 ( .A1(n2642), .A2(opa_r1[19]), .B1(N246), .B2(n2397), .ZN(
        n2401) );
  AOI22_X2 U1367 ( .A1(n2642), .A2(opa_r1[18]), .B1(N245), .B2(n2397), .ZN(
        n2402) );
  AOI22_X2 U1369 ( .A1(n2642), .A2(opa_r1[17]), .B1(N244), .B2(n2397), .ZN(
        n2403) );
  AOI22_X2 U1391 ( .A1(sign_fasu), .A2(n2481), .B1(sign_mul), .B2(fpu_op_r2[1]), .ZN(n2405) );
  NAND2_X2 U1392 ( .A1(n2423), .A2(n2424), .ZN(N224) );
  NOR4_X2 U1393 ( .A1(opa_r1[30]), .A2(opa_r1[29]), .A3(opa_r1[28]), .A4(
        opa_r1[27]), .ZN(n2424) );
  NOR4_X2 U1394 ( .A1(opa_r1[26]), .A2(opa_r1[25]), .A3(opa_r1[24]), .A4(
        opa_r1[23]), .ZN(n2423) );
  OAI221_X2 U1395 ( .B1(n3496), .B2(n2512), .C1(n2617), .C2(n1823), .A(n2425), 
        .ZN(N221) );
  NAND2_X2 U1396 ( .A1(exp_fasu[7]), .A2(n2426), .ZN(n2425) );
  OAI221_X2 U1397 ( .B1(n3496), .B2(n2513), .C1(n2619), .C2(n1823), .A(n2427), 
        .ZN(N220) );
  NAND2_X2 U1398 ( .A1(exp_fasu[6]), .A2(n2426), .ZN(n2427) );
  OAI221_X2 U1399 ( .B1(n3496), .B2(n2508), .C1(n2615), .C2(n1823), .A(n2428), 
        .ZN(N219) );
  NAND2_X2 U1400 ( .A1(exp_fasu[5]), .A2(n2426), .ZN(n2428) );
  OAI221_X2 U1401 ( .B1(n3496), .B2(n2506), .C1(n2613), .C2(n1823), .A(n2429), 
        .ZN(N218) );
  NAND2_X2 U1402 ( .A1(exp_fasu[4]), .A2(n2426), .ZN(n2429) );
  OAI221_X2 U1403 ( .B1(n3496), .B2(n2509), .C1(n2616), .C2(n1823), .A(n2430), 
        .ZN(N217) );
  NAND2_X2 U1404 ( .A1(exp_fasu[3]), .A2(n2426), .ZN(n2430) );
  OR2_X2 U1405 ( .A1(n2481), .A2(fpu_op_r2[2]), .ZN(n1823) );
  OAI221_X2 U1407 ( .B1(n2431), .B2(n2510), .C1(n2618), .C2(n2481), .A(n2432), 
        .ZN(N216) );
  NAND2_X2 U1408 ( .A1(exp_fasu[2]), .A2(n2426), .ZN(n2432) );
  OAI221_X2 U1409 ( .B1(n2431), .B2(n2507), .C1(n2614), .C2(n2481), .A(n2433), 
        .ZN(N215) );
  NAND2_X2 U1410 ( .A1(exp_fasu[1]), .A2(n2426), .ZN(n2433) );
  OAI221_X2 U1411 ( .B1(n2431), .B2(n2505), .C1(n2612), .C2(n2481), .A(n2434), 
        .ZN(N214) );
  NAND2_X2 U1412 ( .A1(exp_fasu[0]), .A2(n2426), .ZN(n2434) );
  NAND2_X2 U1414 ( .A1(fpu_op_r2[2]), .A2(fpu_op_r2[0]), .ZN(n2431) );
  AOI22_X2 U1416 ( .A1(n2437), .A2(n2438), .B1(n2439), .B2(n2589), .ZN(n2436)
         );
  NOR4_X2 U1425 ( .A1(fracta_mul[15]), .A2(fracta_mul[17]), .A3(fracta_mul[19]), .A4(fracta_mul[21]), .ZN(n2437) );
  OAI22_X2 U1428 ( .A1(fracta_mul[22]), .A2(n2446), .B1(n2447), .B2(n2448), 
        .ZN(N141) );
  OAI211_X2 U1429 ( .C1(n2449), .C2(n2450), .A(n2501), .B(n2594), .ZN(n2448)
         );
  OR3_X2 U1431 ( .A1(fracta_mul[6]), .A2(fracta_mul[7]), .A3(fracta_mul[11]), 
        .ZN(n2452) );
  OR2_X2 U1432 ( .A1(fracta_mul[12]), .A2(fracta_mul[13]), .ZN(n2449) );
  AND3_X2 U1434 ( .A1(n2454), .A2(n2589), .A3(n2498), .ZN(n2446) );
  OAI211_X2 U1435 ( .C1(fracta_mul[17]), .C2(fracta_mul[16]), .A(n2580), .B(
        n2496), .ZN(n2454) );
  NOR4_X2 U1438 ( .A1(fracta_mul[19]), .A2(fracta_mul[16]), .A3(n2456), .A4(
        n1819), .ZN(n2455) );
  NAND2_X2 U1439 ( .A1(n2581), .A2(n2496), .ZN(n1819) );
  NOR4_X2 U1440 ( .A1(n2457), .A2(fracta_mul[13]), .A3(fracta_mul[15]), .A4(
        fracta_mul[14]), .ZN(n2456) );
  NOR4_X2 U1444 ( .A1(fracta_mul[7]), .A2(fracta_mul[6]), .A3(fracta_mul[5]), 
        .A4(fracta_mul[4]), .ZN(n2458) );
  OAI33_X1 U1926 ( .A1(n3582), .A2(n1437), .A3(n2474), .B1(n1438), .B2(n1439), 
        .B3(n1440), .ZN(n1436) );
  OAI33_X1 U1928 ( .A1(n3567), .A2(n1878), .A3(n2475), .B1(n1879), .B2(
        inf_mul_r), .B3(n1880), .ZN(N522) );
  OAI33_X1 U1929 ( .A1(n3519), .A2(inf_d), .A3(n1933), .B1(n1934), .B2(n2690), 
        .B3(n1935), .ZN(N519) );
  OAI33_X1 U1930 ( .A1(n2000), .A2(n3504), .A3(n2492), .B1(n2001), .B2(n3584), 
        .B3(n2002), .ZN(n1999) );
  OAI33_X1 U1931 ( .A1(n2140), .A2(r489_B_0_), .A3(n2649), .B1(n2500), .B2(
        sign), .B3(n2142), .ZN(n1955) );
  OAI33_X1 U1932 ( .A1(n2451), .A2(fracta_mul[11]), .A3(fracta_mul[10]), .B1(
        n2452), .B2(fracta_mul[10]), .B3(n2453), .ZN(n2450) );
  DFF_X2 opa_r_reg_31_ ( .D(opa[31]), .CK(clk), .Q(opa_r[31]), .QN(n2601) );
  DFF_X2 opa_r_reg_30_ ( .D(opa[30]), .CK(clk), .Q(opa_r[30]), .QN(n2461) );
  DFF_X2 opa_r_reg_29_ ( .D(opa[29]), .CK(clk), .Q(opa_r[29]), .QN(n2476) );
  DFF_X2 opa_r_reg_28_ ( .D(opa[28]), .CK(clk), .Q(opa_r[28]), .QN(n2574) );
  DFF_X2 opa_r_reg_27_ ( .D(opa[27]), .CK(clk), .Q(opa_r[27]), .QN(n2573) );
  DFF_X2 opa_r_reg_26_ ( .D(opa[26]), .CK(clk), .Q(opa_r[26]), .QN(n2572) );
  DFF_X2 opa_r_reg_25_ ( .D(opa[25]), .CK(clk), .Q(opa_r[25]), .QN(n2575) );
  DFF_X2 opa_r_reg_24_ ( .D(opa[24]), .CK(clk), .Q(opa_r[24]), .QN(n2570) );
  DFF_X2 opa_r_reg_23_ ( .D(opa[23]), .CK(clk), .Q(opa_r[23]), .QN(n2571) );
  DFF_X2 opa_r_reg_22_ ( .D(opa[22]), .CK(clk), .Q(fracta_mul[22]), .QN(n2462)
         );
  DFF_X2 opa_r_reg_21_ ( .D(opa[21]), .CK(clk), .Q(fracta_mul[21]), .QN(n2589)
         );
  DFF_X2 opa_r_reg_20_ ( .D(opa[20]), .CK(clk), .Q(fracta_mul[20]), .QN(n2498)
         );
  DFF_X2 opa_r_reg_19_ ( .D(opa[19]), .CK(clk), .Q(fracta_mul[19]), .QN(n2580)
         );
  DFF_X2 opa_r_reg_18_ ( .D(opa[18]), .CK(clk), .Q(fracta_mul[18]), .QN(n2496)
         );
  DFF_X2 opa_r_reg_17_ ( .D(opa[17]), .CK(clk), .Q(fracta_mul[17]), .QN(n2581)
         );
  DFF_X2 opa_r_reg_16_ ( .D(opa[16]), .CK(clk), .Q(fracta_mul[16]) );
  DFF_X2 opa_r_reg_15_ ( .D(opa[15]), .CK(clk), .Q(fracta_mul[15]), .QN(n2594)
         );
  DFF_X2 opa_r_reg_14_ ( .D(opa[14]), .CK(clk), .Q(fracta_mul[14]), .QN(n2501)
         );
  DFF_X2 opa_r_reg_13_ ( .D(opa[13]), .CK(clk), .Q(fracta_mul[13]) );
  DFF_X2 opa_r_reg_12_ ( .D(opa[12]), .CK(clk), .Q(fracta_mul[12]), .QN(n2590)
         );
  DFF_X2 opa_r_reg_11_ ( .D(opa[11]), .CK(clk), .Q(fracta_mul[11]), .QN(n2588)
         );
  DFF_X2 opa_r_reg_10_ ( .D(opa[10]), .CK(clk), .Q(fracta_mul[10]), .QN(n2497)
         );
  DFF_X2 opa_r_reg_9_ ( .D(opa[9]), .CK(clk), .Q(fracta_mul[9]) );
  DFF_X2 opa_r_reg_8_ ( .D(opa[8]), .CK(clk), .Q(fracta_mul[8]), .QN(n2593) );
  DFF_X2 opa_r_reg_7_ ( .D(opa[7]), .CK(clk), .Q(fracta_mul[7]) );
  DFF_X2 opa_r_reg_6_ ( .D(opa[6]), .CK(clk), .Q(fracta_mul[6]) );
  DFF_X2 opa_r_reg_5_ ( .D(opa[5]), .CK(clk), .Q(fracta_mul[5]) );
  DFF_X2 opa_r_reg_4_ ( .D(opa[4]), .CK(clk), .Q(fracta_mul[4]), .QN(n2591) );
  DFF_X2 opa_r_reg_3_ ( .D(opa[3]), .CK(clk), .Q(fracta_mul[3]), .QN(n2592) );
  DFF_X2 opa_r_reg_2_ ( .D(opa[2]), .CK(clk), .Q(fracta_mul[2]), .QN(n2502) );
  DFF_X2 opa_r_reg_1_ ( .D(opa[1]), .CK(clk), .Q(fracta_mul[1]) );
  DFF_X2 opa_r_reg_0_ ( .D(opa[0]), .CK(clk), .Q(fracta_mul[0]) );
  DFF_X2 opb_r_reg_31_ ( .D(opb[31]), .CK(clk), .Q(opb_r[31]) );
  DFF_X2 opb_r_reg_30_ ( .D(opb[30]), .CK(clk), .Q(opb_r[30]), .QN(n2466) );
  DFF_X2 opb_r_reg_29_ ( .D(opb[29]), .CK(clk), .Q(opb_r[29]), .QN(n2577) );
  DFF_X2 opb_r_reg_28_ ( .D(opb[28]), .CK(clk), .Q(opb_r[28]), .QN(n2494) );
  DFF_X2 opb_r_reg_27_ ( .D(opb[27]), .CK(clk), .Q(opb_r[27]), .QN(n2477) );
  DFF_X2 opb_r_reg_26_ ( .D(opb[26]), .CK(clk), .Q(opb_r[26]), .QN(n2495) );
  DFF_X2 opb_r_reg_25_ ( .D(opb[25]), .CK(clk), .Q(opb_r[25]), .QN(n2478) );
  DFF_X2 opb_r_reg_24_ ( .D(opb[24]), .CK(clk), .Q(opb_r[24]), .QN(n2576) );
  DFF_X2 opb_r_reg_23_ ( .D(opb[23]), .CK(clk), .Q(opb_r[23]), .QN(n2467) );
  DFF_X2 opb_r_reg_22_ ( .D(opb[22]), .CK(clk), .Q(u6_N22), .QN(n2582) );
  DFF_X2 opb_r_reg_21_ ( .D(opb[21]), .CK(clk), .Q(u6_N21) );
  DFF_X2 opb_r_reg_20_ ( .D(opb[20]), .CK(clk), .Q(u6_N20), .QN(n2586) );
  DFF_X2 opb_r_reg_19_ ( .D(opb[19]), .CK(clk), .Q(u6_N19), .QN(n2499) );
  DFF_X2 opb_r_reg_18_ ( .D(opb[18]), .CK(clk), .Q(u6_N18), .QN(n2583) );
  DFF_X2 opb_r_reg_17_ ( .D(opb[17]), .CK(clk), .Q(u6_N17), .QN(n2479) );
  DFF_X2 opb_r_reg_16_ ( .D(opb[16]), .CK(clk), .Q(u6_N16) );
  DFF_X2 opb_r_reg_15_ ( .D(opb[15]), .CK(clk), .Q(u6_N15) );
  DFF_X2 opb_r_reg_14_ ( .D(opb[14]), .CK(clk), .Q(u6_N14) );
  DFF_X2 opb_r_reg_13_ ( .D(opb[13]), .CK(clk), .Q(u6_N13) );
  DFF_X2 opb_r_reg_12_ ( .D(opb[12]), .CK(clk), .Q(u6_N12) );
  DFF_X2 opb_r_reg_11_ ( .D(opb[11]), .CK(clk), .Q(u6_N11) );
  DFF_X2 opb_r_reg_10_ ( .D(opb[10]), .CK(clk), .Q(u6_N10), .QN(n2585) );
  DFF_X2 opb_r_reg_9_ ( .D(opb[9]), .CK(clk), .Q(u6_N9) );
  DFF_X2 opb_r_reg_8_ ( .D(opb[8]), .CK(clk), .Q(u6_N8) );
  DFF_X2 opb_r_reg_7_ ( .D(opb[7]), .CK(clk), .Q(u6_N7) );
  DFF_X2 opb_r_reg_6_ ( .D(opb[6]), .CK(clk), .Q(u6_N6) );
  DFF_X2 opb_r_reg_5_ ( .D(opb[5]), .CK(clk), .Q(u6_N5) );
  DFF_X2 opb_r_reg_4_ ( .D(opb[4]), .CK(clk), .Q(u6_N4) );
  DFF_X2 opb_r_reg_3_ ( .D(opb[3]), .CK(clk), .Q(u6_N3) );
  DFF_X2 opb_r_reg_2_ ( .D(opb[2]), .CK(clk), .Q(u6_N2) );
  DFF_X2 opb_r_reg_1_ ( .D(opb[1]), .CK(clk), .Q(u6_N1) );
  DFF_X2 opb_r_reg_0_ ( .D(opb[0]), .CK(clk), .Q(u6_N0) );
  DFF_X2 rmode_r1_reg_1_ ( .D(rmode[1]), .CK(clk), .Q(rmode_r1[1]) );
  DFF_X2 rmode_r1_reg_0_ ( .D(rmode[0]), .CK(clk), .Q(rmode_r1[0]) );
  DFF_X2 rmode_r2_reg_1_ ( .D(rmode_r1[1]), .CK(clk), .Q(rmode_r2[1]) );
  DFF_X2 rmode_r2_reg_0_ ( .D(rmode_r1[0]), .CK(clk), .Q(rmode_r2[0]) );
  DFF_X2 rmode_r3_reg_1_ ( .D(rmode_r2[1]), .CK(clk), .Q(rmode_r3[1]), .QN(
        n2500) );
  DFF_X2 rmode_r3_reg_0_ ( .D(rmode_r2[0]), .CK(clk), .Q(rmode_r3[0]), .QN(
        n2584) );
  DFF_X2 fpu_op_r1_reg_2_ ( .D(fpu_op[2]), .CK(clk), .Q(fpu_op_r1[2]) );
  DFF_X2 fpu_op_r1_reg_1_ ( .D(fpu_op[1]), .CK(clk), .Q(fpu_op_r1[1]), .QN(
        n2595) );
  DFF_X2 fpu_op_r1_reg_0_ ( .D(fpu_op[0]), .CK(clk), .Q(fpu_op_r1[0]), .QN(
        n2468) );
  DFF_X2 fpu_op_r2_reg_2_ ( .D(fpu_op_r1[2]), .CK(clk), .Q(fpu_op_r2[2]) );
  DFF_X2 fpu_op_r2_reg_1_ ( .D(fpu_op_r1[1]), .CK(clk), .Q(fpu_op_r2[1]), .QN(
        n2481) );
  DFF_X2 fpu_op_r2_reg_0_ ( .D(fpu_op_r1[0]), .CK(clk), .Q(fpu_op_r2[0]), .QN(
        n2606) );
  DFF_X2 fpu_op_r3_reg_2_ ( .D(fpu_op_r2[2]), .CK(clk), .Q(n2460), .QN(n2491)
         );
  DFF_X2 fpu_op_r3_reg_1_ ( .D(fpu_op_r2[1]), .CK(clk), .Q(fpu_op_r3[1]), .QN(
        n2532) );
  DFF_X2 fpu_op_r3_reg_0_ ( .D(fpu_op_r2[0]), .CK(clk), .Q(fpu_op_r3[0]), .QN(
        n2475) );
  DFF_X2 div_opa_ldz_r1_reg_4_ ( .D(N47), .CK(clk), .Q(div_opa_ldz_r1[4]) );
  DFF_X2 div_opa_ldz_r1_reg_3_ ( .D(N75), .CK(clk), .Q(div_opa_ldz_r1[3]) );
  DFF_X2 div_opa_ldz_r1_reg_2_ ( .D(N107), .CK(clk), .Q(div_opa_ldz_r1[2]) );
  DFF_X2 div_opa_ldz_r1_reg_1_ ( .D(N141), .CK(clk), .Q(div_opa_ldz_r1[1]) );
  DFF_X2 div_opa_ldz_r1_reg_0_ ( .D(N170), .CK(clk), .Q(div_opa_ldz_r1[0]) );
  DFF_X2 div_opa_ldz_r2_reg_4_ ( .D(div_opa_ldz_r1[4]), .CK(clk), .Q(
        div_opa_ldz_r2[4]), .QN(n2569) );
  DFF_X2 div_opa_ldz_r2_reg_3_ ( .D(div_opa_ldz_r1[3]), .CK(clk), .Q(
        div_opa_ldz_r2[3]), .QN(n2565) );
  DFF_X2 div_opa_ldz_r2_reg_2_ ( .D(div_opa_ldz_r1[2]), .CK(clk), .Q(
        div_opa_ldz_r2[2]), .QN(n2566) );
  DFF_X2 div_opa_ldz_r2_reg_1_ ( .D(div_opa_ldz_r1[1]), .CK(clk), .Q(
        div_opa_ldz_r2[1]), .QN(n2564) );
  DFF_X2 div_opa_ldz_r2_reg_0_ ( .D(div_opa_ldz_r1[0]), .CK(clk), .Q(
        div_opa_ldz_r2[0]), .QN(n2563) );
  DFF_X2 opa_r1_reg_30_ ( .D(opa_r[30]), .CK(clk), .Q(opa_r1[30]), .QN(n2512)
         );
  DFF_X2 opa_r1_reg_29_ ( .D(opa_r[29]), .CK(clk), .Q(opa_r1[29]), .QN(n2513)
         );
  DFF_X2 opa_r1_reg_28_ ( .D(opa_r[28]), .CK(clk), .Q(opa_r1[28]), .QN(n2508)
         );
  DFF_X2 opa_r1_reg_27_ ( .D(opa_r[27]), .CK(clk), .Q(opa_r1[27]), .QN(n2506)
         );
  DFF_X2 opa_r1_reg_26_ ( .D(opa_r[26]), .CK(clk), .Q(opa_r1[26]), .QN(n2509)
         );
  DFF_X2 opa_r1_reg_25_ ( .D(opa_r[25]), .CK(clk), .Q(opa_r1[25]), .QN(n2510)
         );
  DFF_X2 opa_r1_reg_24_ ( .D(opa_r[24]), .CK(clk), .Q(opa_r1[24]), .QN(n2507)
         );
  DFF_X2 opa_r1_reg_23_ ( .D(opa_r[23]), .CK(clk), .Q(opa_r1[23]), .QN(n2505)
         );
  DFF_X2 opa_r1_reg_22_ ( .D(fracta_mul[22]), .CK(clk), .Q(opa_r1[22]), .QN(
        n2529) );
  DFF_X2 opa_r1_reg_21_ ( .D(fracta_mul[21]), .CK(clk), .Q(opa_r1[21]), .QN(
        n2528) );
  DFF_X2 opa_r1_reg_20_ ( .D(fracta_mul[20]), .CK(clk), .Q(opa_r1[20]), .QN(
        n2527) );
  DFF_X2 opa_r1_reg_19_ ( .D(fracta_mul[19]), .CK(clk), .Q(opa_r1[19]), .QN(
        n2611) );
  DFF_X2 opa_r1_reg_18_ ( .D(fracta_mul[18]), .CK(clk), .Q(opa_r1[18]), .QN(
        n2610) );
  DFF_X2 opa_r1_reg_17_ ( .D(fracta_mul[17]), .CK(clk), .Q(opa_r1[17]), .QN(
        n2609) );
  DFF_X2 opa_r1_reg_16_ ( .D(fracta_mul[16]), .CK(clk), .Q(opa_r1[16]), .QN(
        n2608) );
  DFF_X2 opa_r1_reg_15_ ( .D(fracta_mul[15]), .CK(clk), .Q(opa_r1[15]), .QN(
        n2526) );
  DFF_X2 opa_r1_reg_14_ ( .D(fracta_mul[14]), .CK(clk), .Q(opa_r1[14]), .QN(
        n2525) );
  DFF_X2 opa_r1_reg_13_ ( .D(fracta_mul[13]), .CK(clk), .Q(opa_r1[13]), .QN(
        n2524) );
  DFF_X2 opa_r1_reg_12_ ( .D(fracta_mul[12]), .CK(clk), .Q(opa_r1[12]), .QN(
        n2523) );
  DFF_X2 opa_r1_reg_11_ ( .D(fracta_mul[11]), .CK(clk), .Q(opa_r1[11]), .QN(
        n2522) );
  DFF_X2 opa_r1_reg_10_ ( .D(fracta_mul[10]), .CK(clk), .Q(opa_r1[10]), .QN(
        n2521) );
  DFF_X2 opa_r1_reg_9_ ( .D(fracta_mul[9]), .CK(clk), .Q(opa_r1[9]), .QN(n2520) );
  DFF_X2 opa_r1_reg_8_ ( .D(fracta_mul[8]), .CK(clk), .Q(opa_r1[8]), .QN(n2519) );
  DFF_X2 opa_r1_reg_7_ ( .D(fracta_mul[7]), .CK(clk), .Q(opa_r1[7]), .QN(n2518) );
  DFF_X2 opa_r1_reg_6_ ( .D(fracta_mul[6]), .CK(clk), .Q(opa_r1[6]), .QN(n2517) );
  DFF_X2 opa_r1_reg_5_ ( .D(fracta_mul[5]), .CK(clk), .Q(opa_r1[5]), .QN(n2516) );
  DFF_X2 opa_r1_reg_4_ ( .D(fracta_mul[4]), .CK(clk), .Q(opa_r1[4]), .QN(n2515) );
  DFF_X2 opa_r1_reg_3_ ( .D(fracta_mul[3]), .CK(clk), .Q(opa_r1[3]), .QN(n2514) );
  DFF_X2 opa_r1_reg_2_ ( .D(fracta_mul[2]), .CK(clk), .Q(opa_r1[2]), .QN(n2607) );
  DFF_X2 opa_r1_reg_1_ ( .D(fracta_mul[1]), .CK(clk), .Q(opa_r1[1]), .QN(n2603) );
  DFF_X2 opa_r1_reg_0_ ( .D(fracta_mul[0]), .CK(clk), .Q(N227), .QN(n2504) );
  DFF_X2 opas_r1_reg ( .D(opa_r[31]), .CK(clk), .Q(opas_r1) );
  DFF_X2 opas_r2_reg ( .D(opas_r1), .CK(clk), .Q(opas_r2), .QN(n2567) );
  DFF_X2 u0_fractb_00_reg ( .D(n3486), .CK(clk), .Q(u0_fractb_00) );
  DFF_X2 u0_fracta_00_reg ( .D(n3480), .CK(clk), .Q(u0_fracta_00) );
  DFF_X2 u0_expb_00_reg ( .D(n3485), .CK(clk), .Q(u0_expb_00) );
  DFF_X2 u0_opb_dn_reg ( .D(u0_expb_00), .CK(clk), .Q(opb_dn), .QN(n2463) );
  DFF_X2 u0_opb_00_reg ( .D(u0_N17), .CK(clk), .Q(opb_00) );
  DFF_X2 u0_expa_00_reg ( .D(n2652), .CK(clk), .Q(u0_expa_00) );
  DFF_X2 u0_opa_dn_reg ( .D(u0_expa_00), .CK(clk), .Q(opa_dn), .QN(n2562) );
  DFF_X2 u0_opa_00_reg ( .D(u0_N16), .CK(clk), .Q(opa_00), .QN(n2596) );
  DFF_X2 u0_opb_nan_reg ( .D(u0_N11), .CK(clk), .Q(opb_nan), .QN(n2605) );
  DFF_X2 u0_opa_nan_reg ( .D(u0_N10), .CK(clk), .Q(opa_nan) );
  DFF_X2 opa_nan_r_reg ( .D(N532), .CK(clk), .Q(opa_nan_r) );
  DFF_X2 u0_snan_r_b_reg ( .D(u0_N5), .CK(clk), .Q(u0_snan_r_b) );
  DFF_X2 u0_qnan_r_b_reg ( .D(u6_N22), .CK(clk), .Q(u0_qnan_r_b) );
  DFF_X2 u0_snan_r_a_reg ( .D(u0_N4), .CK(clk), .Q(u0_snan_r_a) );
  DFF_X2 u0_qnan_r_a_reg ( .D(fracta_mul[22]), .CK(clk), .Q(u0_qnan_r_a) );
  DFF_X2 u0_infb_f_r_reg ( .D(n3486), .CK(clk), .Q(u0_infb_f_r) );
  DFF_X2 u0_infa_f_r_reg ( .D(n3480), .CK(clk), .Q(u0_infa_f_r) );
  DFF_X2 u0_expb_ff_reg ( .D(n3484), .CK(clk), .Q(u0_expb_ff) );
  DFF_X2 u0_opb_inf_reg ( .D(n3570), .CK(clk), .Q(opb_inf), .QN(n2598) );
  DFF_X2 u0_expa_ff_reg ( .D(n3478), .CK(clk), .Q(u0_expa_ff) );
  DFF_X2 u0_snan_reg ( .D(n3568), .CK(clk), .Q(snan_d) );
  DFF_X2 snan_reg ( .D(snan_d), .CK(clk), .Q(snan) );
  DFF_X2 u0_qnan_reg ( .D(n3569), .CK(clk), .Q(qnan_d) );
  DFF_X2 u0_opa_inf_reg ( .D(n3571), .CK(clk), .Q(opa_inf), .QN(n2503) );
  DFF_X2 div_by_zero_reg ( .D(N533), .CK(clk), .Q(div_by_zero) );
  DFF_X2 u0_inf_reg ( .D(u0_N7), .CK(clk), .Q(inf_d) );
  DFF_X2 u0_ind_reg ( .D(u0_N6), .CK(clk), .QN(n2602) );
  DFF_X2 u1_fasu_op_reg ( .D(n3445), .CK(clk), .Q(fasu_op), .QN(n2470) );
  DFF_X2 fasu_op_r1_reg ( .D(fasu_op), .CK(clk), .Q(fasu_op_r1) );
  DFF_X2 fasu_op_r2_reg ( .D(fasu_op_r1), .CK(clk), .Q(fasu_op_r2) );
  DFF_X2 qnan_reg ( .D(N524), .CK(clk), .Q(qnan) );
  DFF_X2 u1_fracta_eq_fractb_reg ( .D(u1_N131), .CK(clk), .Q(
        u1_fracta_eq_fractb) );
  DFF_X2 u1_fracta_lt_fractb_reg ( .D(u1_N130), .CK(clk), .Q(
        u1_fracta_lt_fractb) );
  DFF_X2 u1_add_r_reg ( .D(n2468), .CK(clk), .Q(u1_add_r) );
  DFF_X2 u1_signb_r_reg ( .D(opb_r[31]), .CK(clk), .QN(n2600) );
  DFF_X2 u1_signa_r_reg ( .D(opa_r[31]), .CK(clk), .Q(u1_signa_r), .QN(n2604)
         );
  DFF_X2 u1_result_zero_sign_reg ( .D(u1_N129), .CK(clk), .Q(
        result_zero_sign_d) );
  DFF_X2 u1_nan_sign_reg ( .D(u1_N140), .CK(clk), .Q(nan_sign_d) );
  DFF_X2 u1_sign_reg ( .D(u1_sign_d), .CK(clk), .Q(sign_fasu) );
  DFF_X2 sign_fasu_r_reg ( .D(sign_fasu), .CK(clk), .Q(sign_fasu_r) );
  DFF_X2 u1_fractb_out_reg_0_ ( .D(u1_fractb_s[0]), .CK(clk), .Q(fractb[0]) );
  DFF_X2 u1_fractb_out_reg_1_ ( .D(u1_fractb_s[1]), .CK(clk), .Q(fractb[1]) );
  DFF_X2 u1_fractb_out_reg_2_ ( .D(u1_fractb_s[2]), .CK(clk), .Q(fractb[2]) );
  DFF_X2 u1_fractb_out_reg_3_ ( .D(u1_fractb_s[3]), .CK(clk), .Q(fractb[3]) );
  DFF_X2 u1_fractb_out_reg_4_ ( .D(u1_fractb_s[4]), .CK(clk), .Q(fractb[4]) );
  DFF_X2 u1_fractb_out_reg_5_ ( .D(u1_fractb_s[5]), .CK(clk), .Q(fractb[5]) );
  DFF_X2 u1_fractb_out_reg_6_ ( .D(u1_fractb_s[6]), .CK(clk), .Q(fractb[6]) );
  DFF_X2 u1_fractb_out_reg_7_ ( .D(u1_fractb_s[7]), .CK(clk), .Q(fractb[7]) );
  DFF_X2 u1_fractb_out_reg_8_ ( .D(u1_fractb_s[8]), .CK(clk), .Q(fractb[8]) );
  DFF_X2 u1_fractb_out_reg_9_ ( .D(u1_fractb_s[9]), .CK(clk), .Q(fractb[9]) );
  DFF_X2 u1_fractb_out_reg_10_ ( .D(u1_fractb_s[10]), .CK(clk), .Q(fractb[10])
         );
  DFF_X2 u1_fractb_out_reg_11_ ( .D(u1_fractb_s[11]), .CK(clk), .Q(fractb[11])
         );
  DFF_X2 u1_fractb_out_reg_12_ ( .D(u1_fractb_s[12]), .CK(clk), .Q(fractb[12])
         );
  DFF_X2 u1_fractb_out_reg_13_ ( .D(u1_fractb_s[13]), .CK(clk), .Q(fractb[13])
         );
  DFF_X2 u1_fractb_out_reg_14_ ( .D(u1_fractb_s[14]), .CK(clk), .Q(fractb[14])
         );
  DFF_X2 u1_fractb_out_reg_15_ ( .D(u1_fractb_s[15]), .CK(clk), .Q(fractb[15])
         );
  DFF_X2 u1_fractb_out_reg_16_ ( .D(u1_fractb_s[16]), .CK(clk), .Q(fractb[16])
         );
  DFF_X2 u1_fractb_out_reg_17_ ( .D(u1_fractb_s[17]), .CK(clk), .Q(fractb[17])
         );
  DFF_X2 u1_fractb_out_reg_18_ ( .D(u1_fractb_s[18]), .CK(clk), .Q(fractb[18])
         );
  DFF_X2 u1_fractb_out_reg_19_ ( .D(u1_fractb_s[19]), .CK(clk), .Q(fractb[19])
         );
  DFF_X2 u1_fractb_out_reg_20_ ( .D(u1_fractb_s[20]), .CK(clk), .Q(fractb[20])
         );
  DFF_X2 u1_fractb_out_reg_21_ ( .D(u1_fractb_s[21]), .CK(clk), .Q(fractb[21])
         );
  DFF_X2 u1_fractb_out_reg_22_ ( .D(u1_fractb_s[22]), .CK(clk), .Q(fractb[22])
         );
  DFF_X2 u1_fractb_out_reg_23_ ( .D(u1_fractb_s[23]), .CK(clk), .Q(fractb[23])
         );
  DFF_X2 u1_fractb_out_reg_24_ ( .D(u1_fractb_s[24]), .CK(clk), .Q(fractb[24])
         );
  DFF_X2 u1_fractb_out_reg_25_ ( .D(u1_fractb_s[25]), .CK(clk), .Q(fractb[25])
         );
  DFF_X2 u1_fractb_out_reg_26_ ( .D(u1_fractb_s[26]), .CK(clk), .Q(fractb[26])
         );
  DFF_X2 u1_fracta_out_reg_0_ ( .D(u1_fracta_s[0]), .CK(clk), .Q(fracta[0]) );
  DFF_X2 u1_fracta_out_reg_1_ ( .D(u1_fracta_s[1]), .CK(clk), .Q(fracta[1]) );
  DFF_X2 u1_fracta_out_reg_2_ ( .D(u1_fracta_s[2]), .CK(clk), .Q(fracta[2]) );
  DFF_X2 u1_fracta_out_reg_3_ ( .D(u1_fracta_s[3]), .CK(clk), .Q(fracta[3]) );
  DFF_X2 u1_fracta_out_reg_4_ ( .D(u1_fracta_s[4]), .CK(clk), .Q(fracta[4]) );
  DFF_X2 u1_fracta_out_reg_5_ ( .D(u1_fracta_s[5]), .CK(clk), .Q(fracta[5]) );
  DFF_X2 u1_fracta_out_reg_6_ ( .D(u1_fracta_s[6]), .CK(clk), .Q(fracta[6]) );
  DFF_X2 u1_fracta_out_reg_7_ ( .D(u1_fracta_s[7]), .CK(clk), .Q(fracta[7]) );
  DFF_X2 u1_fracta_out_reg_8_ ( .D(u1_fracta_s[8]), .CK(clk), .Q(fracta[8]) );
  DFF_X2 u1_fracta_out_reg_9_ ( .D(u1_fracta_s[9]), .CK(clk), .Q(fracta[9]) );
  DFF_X2 u1_fracta_out_reg_10_ ( .D(u1_fracta_s[10]), .CK(clk), .Q(fracta[10])
         );
  DFF_X2 u1_fracta_out_reg_11_ ( .D(u1_fracta_s[11]), .CK(clk), .Q(fracta[11])
         );
  DFF_X2 u1_fracta_out_reg_12_ ( .D(u1_fracta_s[12]), .CK(clk), .Q(fracta[12])
         );
  DFF_X2 u1_fracta_out_reg_13_ ( .D(u1_fracta_s[13]), .CK(clk), .Q(fracta[13])
         );
  DFF_X2 u1_fracta_out_reg_14_ ( .D(u1_fracta_s[14]), .CK(clk), .Q(fracta[14])
         );
  DFF_X2 u1_fracta_out_reg_15_ ( .D(u1_fracta_s[15]), .CK(clk), .Q(fracta[15])
         );
  DFF_X2 u1_fracta_out_reg_16_ ( .D(u1_fracta_s[16]), .CK(clk), .Q(fracta[16])
         );
  DFF_X2 u1_fracta_out_reg_17_ ( .D(u1_fracta_s[17]), .CK(clk), .Q(fracta[17])
         );
  DFF_X2 u1_fracta_out_reg_18_ ( .D(u1_fracta_s[18]), .CK(clk), .Q(fracta[18])
         );
  DFF_X2 u1_fracta_out_reg_19_ ( .D(u1_fracta_s[19]), .CK(clk), .Q(fracta[19])
         );
  DFF_X2 u1_fracta_out_reg_20_ ( .D(u1_fracta_s[20]), .CK(clk), .Q(fracta[20])
         );
  DFF_X2 u1_fracta_out_reg_21_ ( .D(u1_fracta_s[21]), .CK(clk), .Q(fracta[21])
         );
  DFF_X2 u1_fracta_out_reg_22_ ( .D(u1_fracta_s[22]), .CK(clk), .Q(fracta[22])
         );
  DFF_X2 u1_fracta_out_reg_23_ ( .D(u1_fracta_s[23]), .CK(clk), .Q(fracta[23])
         );
  DFF_X2 u1_fracta_out_reg_24_ ( .D(u1_fracta_s[24]), .CK(clk), .Q(fracta[24])
         );
  DFF_X2 u1_fracta_out_reg_25_ ( .D(u1_fracta_s[25]), .CK(clk), .Q(fracta[25])
         );
  DFF_X2 u1_fracta_out_reg_26_ ( .D(u1_fracta_s[26]), .CK(clk), .Q(fracta[26])
         );
  DFF_X2 fract_out_q_reg_0_ ( .D(n3439), .CK(clk), .Q(fract_out_q[0]) );
  DFF_X2 fract_out_q_reg_1_ ( .D(n3438), .CK(clk), .Q(fract_out_q[1]) );
  DFF_X2 fract_out_q_reg_2_ ( .D(n3437), .CK(clk), .Q(fract_out_q[2]) );
  DFF_X2 fract_out_q_reg_3_ ( .D(n3436), .CK(clk), .Q(fract_out_q[3]) );
  DFF_X2 fract_out_q_reg_4_ ( .D(n3435), .CK(clk), .Q(fract_out_q[4]) );
  DFF_X2 fract_out_q_reg_5_ ( .D(n3434), .CK(clk), .Q(fract_out_q[5]) );
  DFF_X2 fract_out_q_reg_6_ ( .D(n3433), .CK(clk), .Q(fract_out_q[6]) );
  DFF_X2 fract_out_q_reg_7_ ( .D(n3432), .CK(clk), .Q(fract_out_q[7]) );
  DFF_X2 fract_out_q_reg_8_ ( .D(n3431), .CK(clk), .Q(fract_out_q[8]) );
  DFF_X2 fract_out_q_reg_9_ ( .D(n3430), .CK(clk), .Q(fract_out_q[9]) );
  DFF_X2 fract_out_q_reg_10_ ( .D(n3429), .CK(clk), .Q(fract_out_q[10]) );
  DFF_X2 fract_out_q_reg_11_ ( .D(n3428), .CK(clk), .Q(fract_out_q[11]) );
  DFF_X2 fract_out_q_reg_12_ ( .D(n3427), .CK(clk), .Q(fract_out_q[12]) );
  DFF_X2 fract_out_q_reg_13_ ( .D(n3426), .CK(clk), .Q(fract_out_q[13]) );
  DFF_X2 fract_out_q_reg_14_ ( .D(n3425), .CK(clk), .Q(fract_out_q[14]) );
  DFF_X2 fract_out_q_reg_15_ ( .D(n3424), .CK(clk), .Q(fract_out_q[15]) );
  DFF_X2 fract_out_q_reg_16_ ( .D(n3423), .CK(clk), .Q(fract_out_q[16]) );
  DFF_X2 fract_out_q_reg_17_ ( .D(n3422), .CK(clk), .Q(fract_out_q[17]) );
  DFF_X2 fract_out_q_reg_18_ ( .D(n3421), .CK(clk), .Q(fract_out_q[18]) );
  DFF_X2 fract_out_q_reg_19_ ( .D(n3420), .CK(clk), .Q(fract_out_q[19]) );
  DFF_X2 fract_out_q_reg_20_ ( .D(n3419), .CK(clk), .Q(fract_out_q[20]) );
  DFF_X2 fract_out_q_reg_21_ ( .D(n3418), .CK(clk), .Q(fract_out_q[21]) );
  DFF_X2 fract_out_q_reg_22_ ( .D(n3417), .CK(clk), .Q(fract_out_q[22]) );
  DFF_X2 fract_out_q_reg_23_ ( .D(n3416), .CK(clk), .Q(fract_out_q[23]) );
  DFF_X2 fract_out_q_reg_24_ ( .D(n3415), .CK(clk), .Q(fract_out_q[24]) );
  DFF_X2 fract_out_q_reg_25_ ( .D(n3414), .CK(clk), .Q(fract_out_q[25]) );
  DFF_X2 fract_out_q_reg_26_ ( .D(n3413), .CK(clk), .Q(fract_out_q[26]) );
  DFF_X2 fract_out_q_reg_27_ ( .D(n3412), .CK(clk), .Q(fract_out_q[27]) );
  DFF_X2 u1_exp_dn_out_reg_0_ ( .D(u1_N37), .CK(clk), .Q(exp_fasu[0]) );
  DFF_X2 u1_exp_dn_out_reg_1_ ( .D(u1_N38), .CK(clk), .Q(exp_fasu[1]) );
  DFF_X2 u1_exp_dn_out_reg_2_ ( .D(u1_N39), .CK(clk), .Q(exp_fasu[2]) );
  DFF_X2 u1_exp_dn_out_reg_3_ ( .D(u1_N40), .CK(clk), .Q(exp_fasu[3]) );
  DFF_X2 u1_exp_dn_out_reg_4_ ( .D(u1_N41), .CK(clk), .Q(exp_fasu[4]) );
  DFF_X2 u1_exp_dn_out_reg_5_ ( .D(u1_N42), .CK(clk), .Q(exp_fasu[5]) );
  DFF_X2 u1_exp_dn_out_reg_6_ ( .D(u1_N43), .CK(clk), .Q(exp_fasu[6]) );
  DFF_X2 u1_exp_dn_out_reg_7_ ( .D(u1_N44), .CK(clk), .Q(exp_fasu[7]) );
  DFF_X2 u2_sign_exe_reg ( .D(u2_N97), .CK(clk), .Q(sign_exe) );
  DFF_X2 sign_exe_r_reg ( .D(sign_exe), .CK(clk), .QN(n2597) );
  DFF_X2 u2_sign_reg ( .D(u2_sign_d), .CK(clk), .Q(sign_mul) );
  DFF_X2 sign_mul_r_reg ( .D(sign_mul), .CK(clk), .QN(n2599) );
  DFF_X2 sign_reg ( .D(N441), .CK(clk), .Q(sign), .QN(n2587) );
  DFF_X2 fract_i2f_reg_47_ ( .D(N421), .CK(clk), .Q(fract_i2f[47]) );
  DFF_X2 fract_i2f_reg_46_ ( .D(N420), .CK(clk), .Q(fract_i2f[46]) );
  DFF_X2 fract_i2f_reg_45_ ( .D(N419), .CK(clk), .Q(fract_i2f[45]) );
  DFF_X2 fract_i2f_reg_44_ ( .D(N418), .CK(clk), .Q(fract_i2f[44]) );
  DFF_X2 fract_i2f_reg_43_ ( .D(N417), .CK(clk), .Q(fract_i2f[43]) );
  DFF_X2 fract_i2f_reg_42_ ( .D(N416), .CK(clk), .Q(fract_i2f[42]) );
  DFF_X2 fract_i2f_reg_41_ ( .D(N415), .CK(clk), .Q(fract_i2f[41]) );
  DFF_X2 fract_i2f_reg_40_ ( .D(N414), .CK(clk), .Q(fract_i2f[40]) );
  DFF_X2 fract_i2f_reg_39_ ( .D(N413), .CK(clk), .Q(fract_i2f[39]) );
  DFF_X2 fract_i2f_reg_38_ ( .D(N412), .CK(clk), .Q(fract_i2f[38]) );
  DFF_X2 fract_i2f_reg_37_ ( .D(N411), .CK(clk), .Q(fract_i2f[37]) );
  DFF_X2 fract_i2f_reg_36_ ( .D(N410), .CK(clk), .Q(fract_i2f[36]) );
  DFF_X2 fract_i2f_reg_35_ ( .D(N409), .CK(clk), .Q(fract_i2f[35]) );
  DFF_X2 fract_i2f_reg_34_ ( .D(N408), .CK(clk), .Q(fract_i2f[34]) );
  DFF_X2 fract_i2f_reg_33_ ( .D(N407), .CK(clk), .Q(fract_i2f[33]) );
  DFF_X2 fract_i2f_reg_32_ ( .D(N406), .CK(clk), .Q(fract_i2f[32]) );
  DFF_X2 fract_i2f_reg_31_ ( .D(N405), .CK(clk), .Q(fract_i2f[31]) );
  DFF_X2 fract_i2f_reg_30_ ( .D(N404), .CK(clk), .Q(fract_i2f[30]) );
  DFF_X2 fract_i2f_reg_29_ ( .D(N403), .CK(clk), .Q(fract_i2f[29]) );
  DFF_X2 fract_i2f_reg_28_ ( .D(N402), .CK(clk), .Q(fract_i2f[28]) );
  DFF_X2 fract_i2f_reg_27_ ( .D(N401), .CK(clk), .Q(fract_i2f[27]) );
  DFF_X2 fract_i2f_reg_26_ ( .D(N400), .CK(clk), .Q(fract_i2f[26]) );
  DFF_X2 fract_i2f_reg_25_ ( .D(N399), .CK(clk), .Q(fract_i2f[25]) );
  DFF_X2 fract_i2f_reg_24_ ( .D(N398), .CK(clk), .Q(fract_i2f[24]) );
  DFF_X2 fract_i2f_reg_23_ ( .D(N397), .CK(clk), .Q(fract_i2f[23]) );
  DFF_X2 fract_i2f_reg_22_ ( .D(N396), .CK(clk), .Q(fract_i2f[22]) );
  DFF_X2 fract_i2f_reg_21_ ( .D(N395), .CK(clk), .Q(fract_i2f[21]) );
  DFF_X2 fract_i2f_reg_20_ ( .D(N394), .CK(clk), .Q(fract_i2f[20]) );
  DFF_X2 fract_i2f_reg_19_ ( .D(N393), .CK(clk), .Q(fract_i2f[19]) );
  DFF_X2 fract_i2f_reg_18_ ( .D(N392), .CK(clk), .Q(fract_i2f[18]) );
  DFF_X2 fract_i2f_reg_17_ ( .D(N391), .CK(clk), .Q(fract_i2f[17]) );
  DFF_X2 fract_i2f_reg_16_ ( .D(n3355), .CK(clk), .Q(fract_i2f[16]) );
  DFF_X2 fract_i2f_reg_15_ ( .D(n3356), .CK(clk), .Q(fract_i2f[15]) );
  DFF_X2 fract_i2f_reg_14_ ( .D(n3357), .CK(clk), .Q(fract_i2f[14]) );
  DFF_X2 fract_i2f_reg_13_ ( .D(n3358), .CK(clk), .Q(fract_i2f[13]) );
  DFF_X2 fract_i2f_reg_12_ ( .D(n3359), .CK(clk), .Q(fract_i2f[12]) );
  DFF_X2 fract_i2f_reg_11_ ( .D(n3360), .CK(clk), .Q(fract_i2f[11]) );
  DFF_X2 fract_i2f_reg_10_ ( .D(n3361), .CK(clk), .Q(fract_i2f[10]) );
  DFF_X2 fract_i2f_reg_9_ ( .D(n3362), .CK(clk), .Q(fract_i2f[9]) );
  DFF_X2 fract_i2f_reg_8_ ( .D(n3363), .CK(clk), .Q(fract_i2f[8]) );
  DFF_X2 fract_i2f_reg_7_ ( .D(n3364), .CK(clk), .Q(fract_i2f[7]) );
  DFF_X2 fract_i2f_reg_6_ ( .D(n3365), .CK(clk), .Q(fract_i2f[6]) );
  DFF_X2 fract_i2f_reg_5_ ( .D(n3366), .CK(clk), .Q(fract_i2f[5]) );
  DFF_X2 fract_i2f_reg_4_ ( .D(n3367), .CK(clk), .Q(fract_i2f[4]) );
  DFF_X2 fract_i2f_reg_3_ ( .D(n3368), .CK(clk), .Q(fract_i2f[3]) );
  DFF_X2 fract_i2f_reg_2_ ( .D(n3369), .CK(clk), .Q(fract_i2f[2]) );
  DFF_X2 fract_i2f_reg_1_ ( .D(n3370), .CK(clk), .Q(fract_i2f[1]) );
  DFF_X2 fract_i2f_reg_0_ ( .D(n3495), .CK(clk), .Q(fract_i2f[0]) );
  DFF_X2 u2_inf_reg ( .D(u2_N90), .CK(clk), .Q(inf_mul) );
  DFF_X2 inf_mul_r_reg ( .D(inf_mul), .CK(clk), .Q(inf_mul_r) );
  DFF_X2 u2_underflow_reg_0_ ( .D(u2_underflow_d[0]), .CK(clk), .Q(
        underflow_fmul_d[0]) );
  DFF_X2 underflow_fmul_r_reg_0_ ( .D(underflow_fmul_d[0]), .CK(clk), .Q(
        underflow_fmul_r[0]) );
  DFF_X2 u2_underflow_reg_1_ ( .D(u2_underflow_d[1]), .CK(clk), .Q(
        underflow_fmul_d[1]) );
  DFF_X2 underflow_fmul_r_reg_1_ ( .D(underflow_fmul_d[1]), .CK(clk), .Q(
        underflow_fmul_r[1]) );
  DFF_X2 u2_underflow_reg_2_ ( .D(u2_underflow_d[2]), .CK(clk), .Q(
        underflow_fmul_d[2]) );
  DFF_X2 underflow_fmul_r_reg_2_ ( .D(underflow_fmul_d[2]), .CK(clk), .Q(
        underflow_fmul_r[2]) );
  DFF_X2 u2_exp_ovf_reg_0_ ( .D(u2_exp_ovf_d_0_), .CK(clk), .Q(exp_ovf[0]) );
  DFF_X2 exp_ovf_r_reg_0_ ( .D(exp_ovf[0]), .CK(clk), .Q(exp_ovf_r[0]), .QN(
        n2579) );
  DFF_X2 u2_exp_ovf_reg_1_ ( .D(u2_exp_ovf_d_1_), .CK(clk), .Q(exp_ovf[1]) );
  DFF_X2 exp_ovf_r_reg_1_ ( .D(exp_ovf[1]), .CK(clk), .Q(exp_ovf_r[1]), .QN(
        n2492) );
  DFF_X2 u2_exp_out_reg_0_ ( .D(u2_N58), .CK(clk), .Q(exp_mul[0]), .QN(n2612)
         );
  DFF_X2 exp_r_reg_0_ ( .D(N214), .CK(clk), .QN(n2473) );
  DFF_X2 u2_exp_out_reg_1_ ( .D(u2_N59), .CK(clk), .Q(exp_mul[1]), .QN(n2614)
         );
  DFF_X2 exp_r_reg_1_ ( .D(N215), .CK(clk), .QN(n2486) );
  DFF_X2 u2_exp_out_reg_2_ ( .D(u2_N60), .CK(clk), .Q(exp_mul[2]), .QN(n2618)
         );
  DFF_X2 exp_r_reg_2_ ( .D(N216), .CK(clk), .QN(n2559) );
  DFF_X2 u2_exp_out_reg_3_ ( .D(u2_N61), .CK(clk), .Q(exp_mul[3]), .QN(n2616)
         );
  DFF_X2 exp_r_reg_3_ ( .D(N217), .CK(clk), .QN(n2488) );
  DFF_X2 u2_exp_out_reg_4_ ( .D(u2_N62), .CK(clk), .Q(exp_mul[4]), .QN(n2613)
         );
  DFF_X2 exp_r_reg_4_ ( .D(N218), .CK(clk), .QN(n2489) );
  DFF_X2 u2_exp_out_reg_5_ ( .D(u2_N63), .CK(clk), .Q(exp_mul[5]), .QN(n2615)
         );
  DFF_X2 exp_r_reg_5_ ( .D(N219), .CK(clk), .QN(n2487) );
  DFF_X2 u2_exp_out_reg_6_ ( .D(u2_N64), .CK(clk), .Q(exp_mul[6]), .QN(n2619)
         );
  DFF_X2 exp_r_reg_6_ ( .D(N220), .CK(clk), .QN(n2560) );
  DFF_X2 u2_exp_out_reg_7_ ( .D(u2_N65), .CK(clk), .Q(exp_mul[7]), .QN(n2617)
         );
  DFF_X2 exp_r_reg_7_ ( .D(N221), .CK(clk), .QN(n2558) );
  DFF_X2 inf_mul2_reg ( .D(N540), .CK(clk), .Q(inf_mul2) );
  DFF_X2 u5_prod1_reg_0_ ( .D(u5_N0), .CK(clk), .Q(u5_prod1[0]) );
  DFF_X2 u5_prod_reg_0_ ( .D(u5_prod1[0]), .CK(clk), .Q(prod[0]) );
  DFF_X2 u5_prod1_reg_1_ ( .D(u5_N1), .CK(clk), .Q(u5_prod1[1]) );
  DFF_X2 u5_prod_reg_1_ ( .D(u5_prod1[1]), .CK(clk), .Q(prod[1]) );
  DFF_X2 u5_prod1_reg_2_ ( .D(u5_N2), .CK(clk), .Q(u5_prod1[2]) );
  DFF_X2 u5_prod_reg_2_ ( .D(u5_prod1[2]), .CK(clk), .Q(prod[2]) );
  DFF_X2 u5_prod1_reg_3_ ( .D(u5_N3), .CK(clk), .Q(u5_prod1[3]) );
  DFF_X2 u5_prod_reg_3_ ( .D(u5_prod1[3]), .CK(clk), .Q(prod[3]) );
  DFF_X2 u5_prod1_reg_4_ ( .D(u5_N4), .CK(clk), .Q(u5_prod1[4]) );
  DFF_X2 u5_prod_reg_4_ ( .D(u5_prod1[4]), .CK(clk), .Q(prod[4]) );
  DFF_X2 u5_prod1_reg_5_ ( .D(u5_N5), .CK(clk), .Q(u5_prod1[5]) );
  DFF_X2 u5_prod_reg_5_ ( .D(u5_prod1[5]), .CK(clk), .Q(prod[5]) );
  DFF_X2 u5_prod1_reg_6_ ( .D(u5_N6), .CK(clk), .Q(u5_prod1[6]) );
  DFF_X2 u5_prod_reg_6_ ( .D(u5_prod1[6]), .CK(clk), .Q(prod[6]) );
  DFF_X2 u5_prod1_reg_7_ ( .D(u5_N7), .CK(clk), .Q(u5_prod1[7]) );
  DFF_X2 u5_prod_reg_7_ ( .D(u5_prod1[7]), .CK(clk), .Q(prod[7]) );
  DFF_X2 u5_prod1_reg_8_ ( .D(u5_N8), .CK(clk), .Q(u5_prod1[8]) );
  DFF_X2 u5_prod_reg_8_ ( .D(u5_prod1[8]), .CK(clk), .Q(prod[8]) );
  DFF_X2 u5_prod1_reg_9_ ( .D(u5_N9), .CK(clk), .Q(u5_prod1[9]) );
  DFF_X2 u5_prod_reg_9_ ( .D(u5_prod1[9]), .CK(clk), .Q(prod[9]) );
  DFF_X2 u5_prod1_reg_10_ ( .D(u5_N10), .CK(clk), .Q(u5_prod1[10]) );
  DFF_X2 u5_prod_reg_10_ ( .D(u5_prod1[10]), .CK(clk), .Q(prod[10]) );
  DFF_X2 u5_prod1_reg_11_ ( .D(u5_N11), .CK(clk), .Q(u5_prod1[11]) );
  DFF_X2 u5_prod_reg_11_ ( .D(u5_prod1[11]), .CK(clk), .Q(prod[11]) );
  DFF_X2 u5_prod1_reg_12_ ( .D(u5_N12), .CK(clk), .Q(u5_prod1[12]) );
  DFF_X2 u5_prod_reg_12_ ( .D(u5_prod1[12]), .CK(clk), .Q(prod[12]) );
  DFF_X2 u5_prod1_reg_13_ ( .D(u5_N13), .CK(clk), .Q(u5_prod1[13]) );
  DFF_X2 u5_prod_reg_13_ ( .D(u5_prod1[13]), .CK(clk), .Q(prod[13]) );
  DFF_X2 u5_prod1_reg_14_ ( .D(u5_N14), .CK(clk), .Q(u5_prod1[14]) );
  DFF_X2 u5_prod_reg_14_ ( .D(u5_prod1[14]), .CK(clk), .Q(prod[14]) );
  DFF_X2 u5_prod1_reg_15_ ( .D(u5_N15), .CK(clk), .Q(u5_prod1[15]) );
  DFF_X2 u5_prod_reg_15_ ( .D(u5_prod1[15]), .CK(clk), .Q(prod[15]) );
  DFF_X2 u5_prod1_reg_16_ ( .D(u5_N16), .CK(clk), .Q(u5_prod1[16]) );
  DFF_X2 u5_prod_reg_16_ ( .D(u5_prod1[16]), .CK(clk), .Q(prod[16]) );
  DFF_X2 u5_prod1_reg_17_ ( .D(u5_N17), .CK(clk), .Q(u5_prod1[17]) );
  DFF_X2 u5_prod_reg_17_ ( .D(u5_prod1[17]), .CK(clk), .Q(prod[17]) );
  DFF_X2 u5_prod1_reg_18_ ( .D(u5_N18), .CK(clk), .Q(u5_prod1[18]) );
  DFF_X2 u5_prod_reg_18_ ( .D(u5_prod1[18]), .CK(clk), .Q(prod[18]) );
  DFF_X2 u5_prod1_reg_19_ ( .D(u5_N19), .CK(clk), .Q(u5_prod1[19]) );
  DFF_X2 u5_prod_reg_19_ ( .D(u5_prod1[19]), .CK(clk), .Q(prod[19]) );
  DFF_X2 u5_prod1_reg_20_ ( .D(u5_N20), .CK(clk), .Q(u5_prod1[20]) );
  DFF_X2 u5_prod_reg_20_ ( .D(u5_prod1[20]), .CK(clk), .Q(prod[20]) );
  DFF_X2 u5_prod1_reg_21_ ( .D(u5_N21), .CK(clk), .Q(u5_prod1[21]) );
  DFF_X2 u5_prod_reg_21_ ( .D(u5_prod1[21]), .CK(clk), .Q(prod[21]), .QN(n2546) );
  DFF_X2 u5_prod1_reg_22_ ( .D(u5_N22), .CK(clk), .Q(u5_prod1[22]) );
  DFF_X2 u5_prod_reg_22_ ( .D(u5_prod1[22]), .CK(clk), .Q(prod[22]), .QN(n2549) );
  DFF_X2 u5_prod1_reg_23_ ( .D(u5_N23), .CK(clk), .Q(u5_prod1[23]) );
  DFF_X2 u5_prod_reg_23_ ( .D(u5_prod1[23]), .CK(clk), .QN(n2472) );
  DFF_X2 u5_prod1_reg_24_ ( .D(u5_N24), .CK(clk), .Q(u5_prod1[24]) );
  DFF_X2 u5_prod_reg_24_ ( .D(u5_prod1[24]), .CK(clk), .QN(n2545) );
  DFF_X2 u5_prod1_reg_25_ ( .D(u5_N25), .CK(clk), .Q(u5_prod1[25]) );
  DFF_X2 u5_prod_reg_25_ ( .D(u5_prod1[25]), .CK(clk), .QN(n2485) );
  DFF_X2 u5_prod1_reg_26_ ( .D(u5_N26), .CK(clk), .Q(u5_prod1[26]) );
  DFF_X2 u5_prod_reg_26_ ( .D(u5_prod1[26]), .CK(clk), .Q(prod[26]), .QN(n2553) );
  DFF_X2 u5_prod1_reg_27_ ( .D(u5_N27), .CK(clk), .Q(u5_prod1[27]) );
  DFF_X2 u5_prod_reg_27_ ( .D(u5_prod1[27]), .CK(clk), .Q(prod[27]), .QN(n2547) );
  DFF_X2 u5_prod1_reg_28_ ( .D(u5_N28), .CK(clk), .Q(u5_prod1[28]) );
  DFF_X2 u5_prod_reg_28_ ( .D(u5_prod1[28]), .CK(clk), .Q(prod[28]), .QN(n2550) );
  DFF_X2 u5_prod1_reg_29_ ( .D(u5_N29), .CK(clk), .Q(u5_prod1[29]) );
  DFF_X2 u5_prod_reg_29_ ( .D(u5_prod1[29]), .CK(clk), .Q(prod[29]), .QN(n2556) );
  DFF_X2 u5_prod1_reg_30_ ( .D(u5_N30), .CK(clk), .Q(u5_prod1[30]) );
  DFF_X2 u5_prod_reg_30_ ( .D(u5_prod1[30]), .CK(clk), .Q(prod[30]), .QN(n2557) );
  DFF_X2 u5_prod1_reg_31_ ( .D(u5_N31), .CK(clk), .Q(u5_prod1[31]) );
  DFF_X2 u5_prod_reg_31_ ( .D(u5_prod1[31]), .CK(clk), .Q(prod[31]), .QN(n2554) );
  DFF_X2 u5_prod1_reg_32_ ( .D(u5_N32), .CK(clk), .Q(u5_prod1[32]) );
  DFF_X2 u5_prod_reg_32_ ( .D(u5_prod1[32]), .CK(clk), .Q(prod[32]), .QN(n2548) );
  DFF_X2 u5_prod1_reg_33_ ( .D(u5_N33), .CK(clk), .Q(u5_prod1[33]) );
  DFF_X2 u5_prod_reg_33_ ( .D(u5_prod1[33]), .CK(clk), .Q(prod[33]), .QN(n2551) );
  DFF_X2 u5_prod1_reg_34_ ( .D(u5_N34), .CK(clk), .Q(u5_prod1[34]) );
  DFF_X2 u5_prod_reg_34_ ( .D(u5_prod1[34]), .CK(clk), .QN(n2471) );
  DFF_X2 u5_prod1_reg_35_ ( .D(u5_N35), .CK(clk), .Q(u5_prod1[35]) );
  DFF_X2 u5_prod_reg_35_ ( .D(u5_prod1[35]), .CK(clk), .QN(n2544) );
  DFF_X2 u5_prod1_reg_36_ ( .D(u5_N36), .CK(clk), .Q(u5_prod1[36]) );
  DFF_X2 u5_prod_reg_36_ ( .D(u5_prod1[36]), .CK(clk), .QN(n2483) );
  DFF_X2 u5_prod1_reg_37_ ( .D(u5_N37), .CK(clk), .Q(u5_prod1[37]) );
  DFF_X2 u5_prod_reg_37_ ( .D(u5_prod1[37]), .CK(clk), .Q(prod[37]), .QN(n2540) );
  DFF_X2 u5_prod1_reg_38_ ( .D(u5_N38), .CK(clk), .Q(u5_prod1[38]) );
  DFF_X2 u5_prod_reg_38_ ( .D(u5_prod1[38]), .CK(clk), .Q(prod[38]), .QN(n2538) );
  DFF_X2 u5_prod1_reg_39_ ( .D(u5_N39), .CK(clk), .Q(u5_prod1[39]) );
  DFF_X2 u5_prod_reg_39_ ( .D(u5_prod1[39]), .CK(clk), .Q(prod[39]), .QN(n2552) );
  DFF_X2 u5_prod1_reg_40_ ( .D(u5_N40), .CK(clk), .Q(u5_prod1[40]) );
  DFF_X2 u5_prod_reg_40_ ( .D(u5_prod1[40]), .CK(clk), .Q(prod[40]), .QN(n2555) );
  DFF_X2 u5_prod1_reg_41_ ( .D(u5_N41), .CK(clk), .Q(u5_prod1[41]) );
  DFF_X2 u5_prod_reg_41_ ( .D(u5_prod1[41]), .CK(clk), .Q(prod[41]), .QN(n2542) );
  DFF_X2 u5_prod1_reg_42_ ( .D(u5_N42), .CK(clk), .Q(u5_prod1[42]) );
  DFF_X2 u5_prod_reg_42_ ( .D(u5_prod1[42]), .CK(clk), .QN(n2464) );
  DFF_X2 u5_prod1_reg_43_ ( .D(u5_N43), .CK(clk), .Q(u5_prod1[43]) );
  DFF_X2 u5_prod_reg_43_ ( .D(u5_prod1[43]), .CK(clk), .QN(n2534) );
  DFF_X2 u5_prod1_reg_44_ ( .D(u5_N44), .CK(clk), .Q(u5_prod1[44]) );
  DFF_X2 u5_prod_reg_44_ ( .D(u5_prod1[44]), .CK(clk), .QN(n2484) );
  DFF_X2 u5_prod1_reg_45_ ( .D(u5_N45), .CK(clk), .Q(u5_prod1[45]) );
  DFF_X2 u5_prod_reg_45_ ( .D(u5_prod1[45]), .CK(clk), .Q(prod[45]), .QN(n2541) );
  DFF_X2 u5_prod1_reg_46_ ( .D(u5_N46), .CK(clk), .Q(u5_prod1[46]) );
  DFF_X2 u5_prod_reg_46_ ( .D(u5_prod1[46]), .CK(clk), .Q(prod[46]), .QN(n2539) );
  DFF_X2 u5_prod1_reg_47_ ( .D(u5_N47), .CK(clk), .Q(u5_prod1[47]) );
  DFF_X2 u5_prod_reg_47_ ( .D(u5_prod1[47]), .CK(clk), .Q(prod[47]) );
  DFF_X2 u6_remainder_reg_0_ ( .D(u6_N0), .CK(clk), .Q(u6_remainder[0]) );
  DFF_X2 u6_rem_reg_0_ ( .D(u6_remainder[0]), .CK(clk), .Q(remainder[0]) );
  DFF_X2 u6_remainder_reg_1_ ( .D(u6_N1), .CK(clk), .Q(u6_remainder[1]) );
  DFF_X2 u6_rem_reg_1_ ( .D(u6_remainder[1]), .CK(clk), .Q(remainder[1]) );
  DFF_X2 u6_remainder_reg_2_ ( .D(u6_N2), .CK(clk), .Q(u6_remainder[2]) );
  DFF_X2 u6_rem_reg_2_ ( .D(u6_remainder[2]), .CK(clk), .Q(remainder[2]) );
  DFF_X2 u6_remainder_reg_3_ ( .D(u6_N3), .CK(clk), .Q(u6_remainder[3]) );
  DFF_X2 u6_rem_reg_3_ ( .D(u6_remainder[3]), .CK(clk), .Q(remainder[3]) );
  DFF_X2 u6_remainder_reg_4_ ( .D(u6_N4), .CK(clk), .Q(u6_remainder[4]) );
  DFF_X2 u6_rem_reg_4_ ( .D(u6_remainder[4]), .CK(clk), .Q(remainder[4]) );
  DFF_X2 u6_remainder_reg_5_ ( .D(u6_N5), .CK(clk), .Q(u6_remainder[5]) );
  DFF_X2 u6_rem_reg_5_ ( .D(u6_remainder[5]), .CK(clk), .Q(remainder[5]) );
  DFF_X2 u6_remainder_reg_6_ ( .D(u6_N6), .CK(clk), .Q(u6_remainder[6]) );
  DFF_X2 u6_rem_reg_6_ ( .D(u6_remainder[6]), .CK(clk), .Q(remainder[6]) );
  DFF_X2 u6_remainder_reg_7_ ( .D(u6_N7), .CK(clk), .Q(u6_remainder[7]) );
  DFF_X2 u6_rem_reg_7_ ( .D(u6_remainder[7]), .CK(clk), .Q(remainder[7]) );
  DFF_X2 u6_remainder_reg_8_ ( .D(u6_N8), .CK(clk), .Q(u6_remainder[8]) );
  DFF_X2 u6_rem_reg_8_ ( .D(u6_remainder[8]), .CK(clk), .Q(remainder[8]) );
  DFF_X2 u6_remainder_reg_9_ ( .D(u6_N9), .CK(clk), .Q(u6_remainder[9]) );
  DFF_X2 u6_rem_reg_9_ ( .D(u6_remainder[9]), .CK(clk), .Q(remainder[9]) );
  DFF_X2 u6_remainder_reg_10_ ( .D(u6_N10), .CK(clk), .Q(u6_remainder[10]) );
  DFF_X2 u6_rem_reg_10_ ( .D(u6_remainder[10]), .CK(clk), .Q(remainder[10]) );
  DFF_X2 u6_remainder_reg_11_ ( .D(u6_N11), .CK(clk), .Q(u6_remainder[11]) );
  DFF_X2 u6_rem_reg_11_ ( .D(u6_remainder[11]), .CK(clk), .Q(remainder[11]) );
  DFF_X2 u6_remainder_reg_12_ ( .D(u6_N12), .CK(clk), .Q(u6_remainder[12]) );
  DFF_X2 u6_rem_reg_12_ ( .D(u6_remainder[12]), .CK(clk), .Q(remainder[12]) );
  DFF_X2 u6_remainder_reg_13_ ( .D(u6_N13), .CK(clk), .Q(u6_remainder[13]) );
  DFF_X2 u6_rem_reg_13_ ( .D(u6_remainder[13]), .CK(clk), .Q(remainder[13]) );
  DFF_X2 u6_remainder_reg_14_ ( .D(u6_N14), .CK(clk), .Q(u6_remainder[14]) );
  DFF_X2 u6_rem_reg_14_ ( .D(u6_remainder[14]), .CK(clk), .Q(remainder[14]) );
  DFF_X2 u6_remainder_reg_15_ ( .D(u6_N15), .CK(clk), .Q(u6_remainder[15]) );
  DFF_X2 u6_rem_reg_15_ ( .D(u6_remainder[15]), .CK(clk), .Q(remainder[15]) );
  DFF_X2 u6_remainder_reg_16_ ( .D(u6_N16), .CK(clk), .Q(u6_remainder[16]) );
  DFF_X2 u6_rem_reg_16_ ( .D(u6_remainder[16]), .CK(clk), .Q(remainder[16]) );
  DFF_X2 u6_remainder_reg_17_ ( .D(u6_N17), .CK(clk), .Q(u6_remainder[17]) );
  DFF_X2 u6_rem_reg_17_ ( .D(u6_remainder[17]), .CK(clk), .Q(remainder[17]) );
  DFF_X2 u6_remainder_reg_18_ ( .D(u6_N18), .CK(clk), .Q(u6_remainder[18]) );
  DFF_X2 u6_rem_reg_18_ ( .D(u6_remainder[18]), .CK(clk), .Q(remainder[18]) );
  DFF_X2 u6_remainder_reg_19_ ( .D(u6_N19), .CK(clk), .Q(u6_remainder[19]) );
  DFF_X2 u6_rem_reg_19_ ( .D(u6_remainder[19]), .CK(clk), .Q(remainder[19]) );
  DFF_X2 u6_remainder_reg_20_ ( .D(u6_N20), .CK(clk), .Q(u6_remainder[20]) );
  DFF_X2 u6_rem_reg_20_ ( .D(u6_remainder[20]), .CK(clk), .Q(remainder[20]) );
  DFF_X2 u6_remainder_reg_21_ ( .D(u6_N21), .CK(clk), .Q(u6_remainder[21]) );
  DFF_X2 u6_rem_reg_21_ ( .D(u6_remainder[21]), .CK(clk), .Q(remainder[21]) );
  DFF_X2 u6_remainder_reg_22_ ( .D(u6_N22), .CK(clk), .Q(u6_remainder[22]) );
  DFF_X2 u6_rem_reg_22_ ( .D(u6_remainder[22]), .CK(clk), .Q(remainder[22]) );
  DFF_X2 u6_remainder_reg_23_ ( .D(u6_N23), .CK(clk), .Q(u6_remainder[23]) );
  DFF_X2 u6_rem_reg_23_ ( .D(u6_remainder[23]), .CK(clk), .Q(remainder[23]) );
  DFF_X2 u6_remainder_reg_26_ ( .D(u6_N26), .CK(clk), .Q(u6_remainder[26]) );
  DFF_X2 u6_rem_reg_26_ ( .D(u6_remainder[26]), .CK(clk), .Q(remainder[26]) );
  DFF_X2 u6_remainder_reg_27_ ( .D(u6_N27), .CK(clk), .Q(u6_remainder[27]) );
  DFF_X2 u6_rem_reg_27_ ( .D(u6_remainder[27]), .CK(clk), .Q(remainder[27]) );
  DFF_X2 u6_remainder_reg_28_ ( .D(u6_N28), .CK(clk), .Q(u6_remainder[28]) );
  DFF_X2 u6_rem_reg_28_ ( .D(u6_remainder[28]), .CK(clk), .Q(remainder[28]) );
  DFF_X2 u6_remainder_reg_29_ ( .D(u6_N29), .CK(clk), .Q(u6_remainder[29]) );
  DFF_X2 u6_rem_reg_29_ ( .D(u6_remainder[29]), .CK(clk), .Q(remainder[29]) );
  DFF_X2 u6_remainder_reg_30_ ( .D(u6_N30), .CK(clk), .Q(u6_remainder[30]) );
  DFF_X2 u6_rem_reg_30_ ( .D(u6_remainder[30]), .CK(clk), .Q(remainder[30]) );
  DFF_X2 u6_remainder_reg_31_ ( .D(u6_N31), .CK(clk), .Q(u6_remainder[31]) );
  DFF_X2 u6_rem_reg_31_ ( .D(u6_remainder[31]), .CK(clk), .Q(remainder[31]) );
  DFF_X2 u6_remainder_reg_32_ ( .D(u6_N32), .CK(clk), .Q(u6_remainder[32]) );
  DFF_X2 u6_rem_reg_32_ ( .D(u6_remainder[32]), .CK(clk), .Q(remainder[32]) );
  DFF_X2 u6_remainder_reg_33_ ( .D(u6_N33), .CK(clk), .Q(u6_remainder[33]) );
  DFF_X2 u6_rem_reg_33_ ( .D(u6_remainder[33]), .CK(clk), .Q(remainder[33]) );
  DFF_X2 u6_remainder_reg_34_ ( .D(u6_N34), .CK(clk), .Q(u6_remainder[34]) );
  DFF_X2 u6_rem_reg_34_ ( .D(u6_remainder[34]), .CK(clk), .Q(remainder[34]) );
  DFF_X2 u6_remainder_reg_35_ ( .D(u6_N35), .CK(clk), .Q(u6_remainder[35]) );
  DFF_X2 u6_rem_reg_35_ ( .D(u6_remainder[35]), .CK(clk), .Q(remainder[35]) );
  DFF_X2 u6_remainder_reg_36_ ( .D(u6_N36), .CK(clk), .Q(u6_remainder[36]) );
  DFF_X2 u6_rem_reg_36_ ( .D(u6_remainder[36]), .CK(clk), .Q(remainder[36]) );
  DFF_X2 u6_remainder_reg_37_ ( .D(u6_N37), .CK(clk), .Q(u6_remainder[37]) );
  DFF_X2 u6_rem_reg_37_ ( .D(u6_remainder[37]), .CK(clk), .Q(remainder[37]) );
  DFF_X2 u6_remainder_reg_38_ ( .D(u6_N38), .CK(clk), .Q(u6_remainder[38]) );
  DFF_X2 u6_rem_reg_38_ ( .D(u6_remainder[38]), .CK(clk), .Q(remainder[38]) );
  DFF_X2 u6_remainder_reg_39_ ( .D(u6_N39), .CK(clk), .Q(u6_remainder[39]) );
  DFF_X2 u6_rem_reg_39_ ( .D(u6_remainder[39]), .CK(clk), .Q(remainder[39]) );
  DFF_X2 u6_remainder_reg_40_ ( .D(u6_N40), .CK(clk), .Q(u6_remainder[40]) );
  DFF_X2 u6_rem_reg_40_ ( .D(u6_remainder[40]), .CK(clk), .Q(remainder[40]) );
  DFF_X2 u6_remainder_reg_41_ ( .D(u6_N41), .CK(clk), .Q(u6_remainder[41]) );
  DFF_X2 u6_rem_reg_41_ ( .D(u6_remainder[41]), .CK(clk), .Q(remainder[41]) );
  DFF_X2 u6_remainder_reg_42_ ( .D(u6_N42), .CK(clk), .Q(u6_remainder[42]) );
  DFF_X2 u6_rem_reg_42_ ( .D(u6_remainder[42]), .CK(clk), .Q(remainder[42]) );
  DFF_X2 u6_remainder_reg_43_ ( .D(u6_N43), .CK(clk), .Q(u6_remainder[43]) );
  DFF_X2 u6_rem_reg_43_ ( .D(u6_remainder[43]), .CK(clk), .Q(remainder[43]) );
  DFF_X2 u6_remainder_reg_44_ ( .D(u6_N44), .CK(clk), .Q(u6_remainder[44]) );
  DFF_X2 u6_rem_reg_44_ ( .D(u6_remainder[44]), .CK(clk), .Q(remainder[44]) );
  DFF_X2 u6_remainder_reg_45_ ( .D(u6_N45), .CK(clk), .Q(u6_remainder[45]) );
  DFF_X2 u6_rem_reg_45_ ( .D(u6_remainder[45]), .CK(clk), .Q(remainder[45]) );
  DFF_X2 u6_remainder_reg_46_ ( .D(u6_N46), .CK(clk), .Q(u6_remainder[46]) );
  DFF_X2 u6_rem_reg_46_ ( .D(u6_remainder[46]), .CK(clk), .Q(remainder[46]) );
  DFF_X2 u6_remainder_reg_47_ ( .D(u6_N47), .CK(clk), .Q(u6_remainder[47]) );
  DFF_X2 u6_rem_reg_47_ ( .D(u6_remainder[47]), .CK(clk), .Q(remainder[47]) );
  DFF_X2 u6_remainder_reg_48_ ( .D(u6_N48), .CK(clk), .Q(u6_remainder[48]) );
  DFF_X2 u6_rem_reg_48_ ( .D(u6_remainder[48]), .CK(clk), .Q(remainder[48]) );
  DFF_X2 u6_remainder_reg_49_ ( .D(u6_N49), .CK(clk), .Q(u6_remainder[49]) );
  DFF_X2 u6_rem_reg_49_ ( .D(u6_remainder[49]), .CK(clk), .Q(remainder[49]) );
  DFF_X2 u6_quo1_reg_0_ ( .D(u6_N0), .CK(clk), .Q(u6_quo1[0]) );
  DFF_X2 u6_quo_reg_0_ ( .D(u6_quo1[0]), .CK(clk), .Q(quo[0]) );
  DFF_X2 u6_quo1_reg_1_ ( .D(u6_N1), .CK(clk), .Q(u6_quo1[1]) );
  DFF_X2 u6_quo_reg_1_ ( .D(u6_quo1[1]), .CK(clk), .Q(quo[1]) );
  DFF_X2 u6_quo1_reg_2_ ( .D(u6_N2), .CK(clk), .Q(u6_quo1[2]) );
  DFF_X2 u6_quo_reg_2_ ( .D(u6_quo1[2]), .CK(clk), .Q(quo[2]) );
  DFF_X2 u6_quo1_reg_3_ ( .D(u6_N3), .CK(clk), .Q(u6_quo1[3]) );
  DFF_X2 u6_quo_reg_3_ ( .D(u6_quo1[3]), .CK(clk), .Q(quo[3]) );
  DFF_X2 u6_quo1_reg_4_ ( .D(u6_N4), .CK(clk), .Q(u6_quo1[4]) );
  DFF_X2 u6_quo_reg_4_ ( .D(u6_quo1[4]), .CK(clk), .Q(quo[4]) );
  DFF_X2 u6_quo1_reg_5_ ( .D(u6_N5), .CK(clk), .Q(u6_quo1[5]) );
  DFF_X2 u6_quo_reg_5_ ( .D(u6_quo1[5]), .CK(clk), .Q(quo[5]) );
  DFF_X2 u6_quo1_reg_6_ ( .D(u6_N6), .CK(clk), .Q(u6_quo1[6]) );
  DFF_X2 u6_quo_reg_6_ ( .D(u6_quo1[6]), .CK(clk), .Q(quo[6]) );
  DFF_X2 u6_quo1_reg_7_ ( .D(u6_N7), .CK(clk), .Q(u6_quo1[7]) );
  DFF_X2 u6_quo_reg_7_ ( .D(u6_quo1[7]), .CK(clk), .Q(quo[7]) );
  DFF_X2 u6_quo1_reg_8_ ( .D(u6_N8), .CK(clk), .Q(u6_quo1[8]) );
  DFF_X2 u6_quo_reg_8_ ( .D(u6_quo1[8]), .CK(clk), .Q(quo[8]) );
  DFF_X2 u6_quo1_reg_9_ ( .D(u6_N9), .CK(clk), .Q(u6_quo1[9]) );
  DFF_X2 u6_quo_reg_9_ ( .D(u6_quo1[9]), .CK(clk), .Q(quo[9]) );
  DFF_X2 u6_quo1_reg_10_ ( .D(u6_N10), .CK(clk), .Q(u6_quo1[10]) );
  DFF_X2 u6_quo_reg_10_ ( .D(u6_quo1[10]), .CK(clk), .Q(quo[10]) );
  DFF_X2 u6_quo1_reg_11_ ( .D(u6_N11), .CK(clk), .Q(u6_quo1[11]) );
  DFF_X2 u6_quo_reg_11_ ( .D(u6_quo1[11]), .CK(clk), .Q(quo[11]) );
  DFF_X2 u6_quo1_reg_12_ ( .D(u6_N12), .CK(clk), .Q(u6_quo1[12]) );
  DFF_X2 u6_quo_reg_12_ ( .D(u6_quo1[12]), .CK(clk), .Q(quo[12]) );
  DFF_X2 u6_quo1_reg_13_ ( .D(u6_N13), .CK(clk), .Q(u6_quo1[13]) );
  DFF_X2 u6_quo_reg_13_ ( .D(u6_quo1[13]), .CK(clk), .Q(quo[13]) );
  DFF_X2 u6_quo1_reg_14_ ( .D(u6_N14), .CK(clk), .Q(u6_quo1[14]) );
  DFF_X2 u6_quo_reg_14_ ( .D(u6_quo1[14]), .CK(clk), .Q(quo[14]) );
  DFF_X2 u6_quo1_reg_15_ ( .D(u6_N15), .CK(clk), .Q(u6_quo1[15]) );
  DFF_X2 u6_quo_reg_15_ ( .D(u6_quo1[15]), .CK(clk), .Q(quo[15]) );
  DFF_X2 u6_quo1_reg_16_ ( .D(u6_N16), .CK(clk), .Q(u6_quo1[16]) );
  DFF_X2 u6_quo_reg_16_ ( .D(u6_quo1[16]), .CK(clk), .Q(quo[16]) );
  DFF_X2 u6_quo1_reg_17_ ( .D(u6_N17), .CK(clk), .Q(u6_quo1[17]) );
  DFF_X2 u6_quo_reg_17_ ( .D(u6_quo1[17]), .CK(clk), .Q(quo[17]) );
  DFF_X2 u6_quo1_reg_18_ ( .D(u6_N18), .CK(clk), .Q(u6_quo1[18]) );
  DFF_X2 u6_quo_reg_18_ ( .D(u6_quo1[18]), .CK(clk), .Q(quo[18]) );
  DFF_X2 u6_quo1_reg_19_ ( .D(u6_N19), .CK(clk), .Q(u6_quo1[19]) );
  DFF_X2 u6_quo_reg_19_ ( .D(u6_quo1[19]), .CK(clk), .Q(quo[19]) );
  DFF_X2 u6_quo1_reg_20_ ( .D(u6_N20), .CK(clk), .Q(u6_quo1[20]) );
  DFF_X2 u6_quo_reg_20_ ( .D(u6_quo1[20]), .CK(clk), .Q(quo[20]) );
  DFF_X2 u6_quo1_reg_21_ ( .D(u6_N21), .CK(clk), .Q(u6_quo1[21]) );
  DFF_X2 u6_quo_reg_21_ ( .D(u6_quo1[21]), .CK(clk), .Q(quo[21]) );
  DFF_X2 u6_quo1_reg_22_ ( .D(u6_N22), .CK(clk), .Q(u6_quo1[22]) );
  DFF_X2 u6_quo_reg_22_ ( .D(u6_quo1[22]), .CK(clk), .Q(quo[22]) );
  DFF_X2 u6_quo1_reg_23_ ( .D(u6_N23), .CK(clk), .Q(u6_quo1[23]) );
  DFF_X2 u6_quo_reg_23_ ( .D(u6_quo1[23]), .CK(clk), .Q(quo[23]) );
  DFF_X2 u6_quo1_reg_26_ ( .D(u6_N26), .CK(clk), .Q(u6_quo1[26]) );
  DFF_X2 u6_quo_reg_26_ ( .D(u6_quo1[26]), .CK(clk), .Q(quo[26]), .QN(n2537)
         );
  DFF_X2 u6_quo1_reg_27_ ( .D(u6_N27), .CK(clk), .Q(u6_quo1[27]) );
  DFF_X2 u6_quo_reg_27_ ( .D(u6_quo1[27]), .CK(clk), .Q(quo[27]) );
  DFF_X2 u6_quo1_reg_28_ ( .D(u6_N28), .CK(clk), .Q(u6_quo1[28]) );
  DFF_X2 u6_quo_reg_28_ ( .D(u6_quo1[28]), .CK(clk), .Q(quo[28]) );
  DFF_X2 u6_quo1_reg_29_ ( .D(u6_N29), .CK(clk), .Q(u6_quo1[29]) );
  DFF_X2 u6_quo_reg_29_ ( .D(u6_quo1[29]), .CK(clk), .Q(quo[29]) );
  DFF_X2 u6_quo1_reg_30_ ( .D(u6_N30), .CK(clk), .Q(u6_quo1[30]) );
  DFF_X2 u6_quo_reg_30_ ( .D(u6_quo1[30]), .CK(clk), .Q(quo[30]) );
  DFF_X2 u6_quo1_reg_31_ ( .D(u6_N31), .CK(clk), .Q(u6_quo1[31]) );
  DFF_X2 u6_quo_reg_31_ ( .D(u6_quo1[31]), .CK(clk), .Q(quo[31]) );
  DFF_X2 u6_quo1_reg_32_ ( .D(u6_N32), .CK(clk), .Q(u6_quo1[32]) );
  DFF_X2 u6_quo_reg_32_ ( .D(u6_quo1[32]), .CK(clk), .Q(quo[32]) );
  DFF_X2 u6_quo1_reg_33_ ( .D(u6_N33), .CK(clk), .Q(u6_quo1[33]) );
  DFF_X2 u6_quo_reg_33_ ( .D(u6_quo1[33]), .CK(clk), .Q(quo[33]) );
  DFF_X2 u6_quo1_reg_34_ ( .D(u6_N34), .CK(clk), .Q(u6_quo1[34]) );
  DFF_X2 u6_quo_reg_34_ ( .D(u6_quo1[34]), .CK(clk), .Q(quo[34]) );
  DFF_X2 u6_quo1_reg_35_ ( .D(u6_N35), .CK(clk), .Q(u6_quo1[35]) );
  DFF_X2 u6_quo_reg_35_ ( .D(u6_quo1[35]), .CK(clk), .Q(quo[35]) );
  DFF_X2 u6_quo1_reg_36_ ( .D(u6_N36), .CK(clk), .Q(u6_quo1[36]) );
  DFF_X2 u6_quo_reg_36_ ( .D(u6_quo1[36]), .CK(clk), .Q(quo[36]) );
  DFF_X2 u6_quo1_reg_37_ ( .D(u6_N37), .CK(clk), .Q(u6_quo1[37]) );
  DFF_X2 u6_quo_reg_37_ ( .D(u6_quo1[37]), .CK(clk), .Q(quo[37]) );
  DFF_X2 u6_quo1_reg_38_ ( .D(u6_N38), .CK(clk), .Q(u6_quo1[38]) );
  DFF_X2 u6_quo_reg_38_ ( .D(u6_quo1[38]), .CK(clk), .Q(quo[38]) );
  DFF_X2 u6_quo1_reg_39_ ( .D(u6_N39), .CK(clk), .Q(u6_quo1[39]) );
  DFF_X2 u6_quo_reg_39_ ( .D(u6_quo1[39]), .CK(clk), .Q(quo[39]) );
  DFF_X2 u6_quo1_reg_40_ ( .D(u6_N40), .CK(clk), .Q(u6_quo1[40]) );
  DFF_X2 u6_quo_reg_40_ ( .D(u6_quo1[40]), .CK(clk), .Q(quo[40]) );
  DFF_X2 u6_quo1_reg_41_ ( .D(u6_N41), .CK(clk), .Q(u6_quo1[41]) );
  DFF_X2 u6_quo_reg_41_ ( .D(u6_quo1[41]), .CK(clk), .Q(quo[41]) );
  DFF_X2 u6_quo1_reg_42_ ( .D(u6_N42), .CK(clk), .Q(u6_quo1[42]) );
  DFF_X2 u6_quo_reg_42_ ( .D(u6_quo1[42]), .CK(clk), .Q(quo[42]) );
  DFF_X2 u6_quo1_reg_43_ ( .D(u6_N43), .CK(clk), .Q(u6_quo1[43]) );
  DFF_X2 u6_quo_reg_43_ ( .D(u6_quo1[43]), .CK(clk), .Q(quo[43]) );
  DFF_X2 u6_quo1_reg_44_ ( .D(u6_N44), .CK(clk), .Q(u6_quo1[44]) );
  DFF_X2 u6_quo_reg_44_ ( .D(u6_quo1[44]), .CK(clk), .Q(quo[44]) );
  DFF_X2 u6_quo1_reg_45_ ( .D(u6_N45), .CK(clk), .Q(u6_quo1[45]) );
  DFF_X2 u6_quo_reg_45_ ( .D(u6_quo1[45]), .CK(clk), .Q(quo[45]) );
  DFF_X2 u6_quo1_reg_46_ ( .D(u6_N46), .CK(clk), .Q(u6_quo1[46]) );
  DFF_X2 u6_quo_reg_46_ ( .D(u6_quo1[46]), .CK(clk), .Q(quo[46]) );
  DFF_X2 u6_quo1_reg_47_ ( .D(u6_N47), .CK(clk), .Q(u6_quo1[47]) );
  DFF_X2 u6_quo_reg_47_ ( .D(u6_quo1[47]), .CK(clk), .Q(quo[47]) );
  DFF_X2 u6_quo1_reg_48_ ( .D(u6_N48), .CK(clk), .Q(u6_quo1[48]) );
  DFF_X2 u6_quo_reg_48_ ( .D(u6_quo1[48]), .CK(clk), .Q(quo[48]) );
  DFF_X2 out_reg_23_ ( .D(N468), .CK(clk), .Q(out[23]) );
  DFF_X2 out_reg_27_ ( .D(N472), .CK(clk), .Q(out[27]) );
  DFF_X2 out_reg_28_ ( .D(N473), .CK(clk), .Q(out[28]) );
  DFF_X2 out_reg_29_ ( .D(N474), .CK(clk), .Q(out[29]) );
  DFF_X2 out_reg_30_ ( .D(N475), .CK(clk), .Q(out[30]) );
  DFF_X2 out_reg_24_ ( .D(N469), .CK(clk), .Q(out[24]) );
  DFF_X2 out_reg_25_ ( .D(N470), .CK(clk), .Q(out[25]) );
  DFF_X2 out_reg_26_ ( .D(N471), .CK(clk), .Q(out[26]) );
  DFF_X2 overflow_reg ( .D(N519), .CK(clk), .Q(overflow) );
  DFF_X2 out_reg_22_ ( .D(N467), .CK(clk), .Q(out[22]) );
  DFF_X2 out_reg_21_ ( .D(N466), .CK(clk), .Q(out[21]) );
  DFF_X2 out_reg_20_ ( .D(N465), .CK(clk), .Q(out[20]) );
  DFF_X2 out_reg_19_ ( .D(N464), .CK(clk), .Q(out[19]) );
  DFF_X2 out_reg_18_ ( .D(N463), .CK(clk), .Q(out[18]) );
  DFF_X2 out_reg_17_ ( .D(N462), .CK(clk), .Q(out[17]) );
  DFF_X2 out_reg_16_ ( .D(N461), .CK(clk), .Q(out[16]) );
  DFF_X2 out_reg_15_ ( .D(N460), .CK(clk), .Q(out[15]) );
  DFF_X2 out_reg_14_ ( .D(N459), .CK(clk), .Q(out[14]) );
  DFF_X2 out_reg_13_ ( .D(N458), .CK(clk), .Q(out[13]) );
  DFF_X2 out_reg_12_ ( .D(N457), .CK(clk), .Q(out[12]) );
  DFF_X2 out_reg_11_ ( .D(N456), .CK(clk), .Q(out[11]) );
  DFF_X2 out_reg_10_ ( .D(N455), .CK(clk), .Q(out[10]) );
  DFF_X2 out_reg_9_ ( .D(N454), .CK(clk), .Q(out[9]) );
  DFF_X2 out_reg_8_ ( .D(N453), .CK(clk), .Q(out[8]) );
  DFF_X2 out_reg_7_ ( .D(N452), .CK(clk), .Q(out[7]) );
  DFF_X2 out_reg_6_ ( .D(N451), .CK(clk), .Q(out[6]) );
  DFF_X2 out_reg_5_ ( .D(N450), .CK(clk), .Q(out[5]) );
  DFF_X2 out_reg_4_ ( .D(N449), .CK(clk), .Q(out[4]) );
  DFF_X2 out_reg_3_ ( .D(N448), .CK(clk), .Q(out[3]) );
  DFF_X2 out_reg_2_ ( .D(N447), .CK(clk), .Q(out[2]) );
  DFF_X2 out_reg_1_ ( .D(N446), .CK(clk), .Q(out[1]) );
  DFF_X2 inf_reg ( .D(N526), .CK(clk), .Q(inf) );
  DFF_X2 underflow_reg ( .D(N522), .CK(clk), .Q(underflow) );
  DFF_X2 ine_reg ( .D(N509), .CK(clk), .Q(ine) );
  DFF_X2 zero_reg ( .D(N531), .CK(clk), .Q(zero) );
  DFF_X2 out_reg_31_ ( .D(N495), .CK(clk), .Q(out[31]) );
  DFF_X2 out_reg_0_ ( .D(N445), .CK(clk), .Q(out[0]) );
  DFF_X2 u6_quo1_reg_49_ ( .D(u6_N49), .CK(clk), .Q(u6_quo1[49]) );
  DFF_X2 u6_quo_reg_49_ ( .D(u6_quo1[49]), .CK(clk), .Q(quo[49]) );
  FA_X1 u4_add_486_U1_1 ( .A(div_opa_ldz_r2[1]), .B(u4_fi_ldz_1_), .CI(
        u4_add_486_carry[1]), .CO(u4_add_486_carry[2]), .S(u4_ldz_all_1_) );
  FA_X1 u4_add_486_U1_2 ( .A(div_opa_ldz_r2[2]), .B(u4_fi_ldz_2_), .CI(
        u4_add_486_carry[2]), .CO(u4_add_486_carry[3]), .S(u4_ldz_all_2_) );
  FA_X1 u4_add_486_U1_3 ( .A(div_opa_ldz_r2[3]), .B(u4_fi_ldz_2a_3_), .CI(
        u4_add_486_carry[3]), .CO(u4_add_486_carry[4]), .S(u4_ldz_all_3_) );
  FA_X1 u4_add_486_U1_4 ( .A(div_opa_ldz_r2[4]), .B(u4_fi_ldz_4_), .CI(
        u4_add_486_carry[4]), .CO(u4_add_486_carry[5]), .S(u4_ldz_all_4_) );
  FA_X1 u4_sub_406_U2_1 ( .A(n2681), .B(n2564), .CI(u4_sub_406_carry[1]), .CO(
        u4_sub_406_carry[2]), .S(u4_div_scht1a[1]) );
  FA_X1 u4_sub_406_U2_2 ( .A(n2682), .B(n2566), .CI(u4_sub_406_carry[2]), .CO(
        u4_sub_406_carry[3]), .S(u4_div_scht1a[2]) );
  FA_X1 u4_sub_406_U2_3 ( .A(n2683), .B(n2565), .CI(u4_sub_406_carry[3]), .CO(
        u4_sub_406_carry[4]), .S(u4_div_scht1a[3]) );
  FA_X1 u4_sub_406_U2_4 ( .A(n2684), .B(n2569), .CI(u4_sub_406_carry[4]), .CO(
        u4_sub_406_carry[5]), .S(u4_div_scht1a[4]) );
  NAND2_X2 U1933 ( .A1(quo[48]), .A2(n2643), .ZN(n2325) );
  NAND2_X2 U1934 ( .A1(quo[2]), .A2(n2320), .ZN(n2351) );
  NAND2_X2 U1935 ( .A1(quo[47]), .A2(n2643), .ZN(n2327) );
  NAND2_X2 U1936 ( .A1(quo[1]), .A2(n2320), .ZN(n2367) );
  INV_X4 U1937 ( .A(remainder[23]), .ZN(n2296) );
  NOR3_X2 U1938 ( .A1(u4_N1429), .A2(u4_N1431), .A3(u4_N1430), .ZN(n2277) );
  NOR3_X2 U1939 ( .A1(u4_N1417), .A2(u4_N1419), .A3(u4_N1418), .ZN(n2273) );
  INV_X4 U1940 ( .A(n2659), .ZN(n2658) );
  NOR3_X2 U1941 ( .A1(n3529), .A2(n3560), .A3(n3530), .ZN(n2221) );
  NOR3_X2 U1942 ( .A1(n3533), .A2(n3521), .A3(n3534), .ZN(n2223) );
  NOR3_X2 U1943 ( .A1(n3525), .A2(n3528), .A3(n3526), .ZN(n2228) );
  NOR3_X2 U1944 ( .A1(fract_denorm[23]), .A2(n3563), .A3(n3522), .ZN(n2226) );
  AOI21_X2 U1945 ( .B1(n1966), .B2(n2490), .A(n2007), .ZN(n2233) );
  NOR2_X2 U1946 ( .A1(n2682), .A2(n2681), .ZN(n2249) );
  OAI21_X2 U1947 ( .B1(n2647), .B2(n3565), .A(n2000), .ZN(n2237) );
  NOR3_X2 U1948 ( .A1(fract_denorm[37]), .A2(fract_denorm[38]), .A3(
        fract_denorm[36]), .ZN(n1554) );
  NOR3_X2 U1949 ( .A1(fract_denorm[34]), .A2(fract_denorm[35]), .A3(n3549), 
        .ZN(n1552) );
  NOR3_X2 U1950 ( .A1(n3545), .A2(n2648), .A3(n3553), .ZN(n2252) );
  NOR3_X2 U1951 ( .A1(u4_N1420), .A2(u4_N1422), .A3(u4_N1421), .ZN(n2274) );
  NOR3_X2 U1952 ( .A1(u4_N1423), .A2(u4_N1425), .A3(u4_N1424), .ZN(n2275) );
  NOR3_X2 U1953 ( .A1(u4_N1426), .A2(u4_N1428), .A3(u4_N1427), .ZN(n2276) );
  NOR3_X2 U1954 ( .A1(u4_N1408), .A2(u4_N1410), .A3(u4_N1409), .ZN(n2270) );
  NOR3_X2 U1955 ( .A1(u4_N1411), .A2(u4_N1413), .A3(u4_N1412), .ZN(n2271) );
  NOR3_X2 U1956 ( .A1(u4_N1414), .A2(u4_N1416), .A3(u4_N1415), .ZN(n2272) );
  NOR3_X2 U1957 ( .A1(n2755), .A2(n2543), .A3(u4_fi_ldz_2a_5_), .ZN(u4_N1572)
         );
  NOR2_X2 U1958 ( .A1(exp_ovf_r[0]), .A2(exp_ovf_r[1]), .ZN(n2129) );
  AOI21_X2 U1959 ( .B1(u4_N1572), .B2(n2014), .A(n3354), .ZN(n2139) );
  AOI21_X2 U1960 ( .B1(n3584), .B2(exp_ovf_r[0]), .A(n3354), .ZN(n2138) );
  NOR3_X2 U1961 ( .A1(n2136), .A2(n2558), .A3(n2115), .ZN(n2135) );
  OAI21_X2 U1962 ( .B1(u4_exp_out_mi1[0]), .B2(n2130), .A(n2137), .ZN(n2136)
         );
  OAI21_X2 U1963 ( .B1(u4_exp_out_mi1[0]), .B2(n2174), .A(n2175), .ZN(n2173)
         );
  NAND3_X2 U1964 ( .A1(n2174), .A2(n3520), .A3(u4_exp_out_pl1_0_), .ZN(n2175)
         );
  NAND3_X2 U1965 ( .A1(n1949), .A2(n2647), .A3(n2200), .ZN(n2202) );
  NOR2_X2 U1966 ( .A1(n2128), .A2(n3353), .ZN(n2150) );
  AOI21_X2 U1967 ( .B1(n2129), .B2(n2128), .A(n1417), .ZN(n2146) );
  OAI21_X2 U1968 ( .B1(n3583), .B2(n2687), .A(n2017), .ZN(n2145) );
  NAND3_X2 U1969 ( .A1(opb_dn), .A2(n2562), .A3(u4_N1523), .ZN(n2140) );
  INV_X4 U1970 ( .A(n2659), .ZN(n2657) );
  INV_X4 U1971 ( .A(n2669), .ZN(n2668) );
  INV_X4 U1972 ( .A(u1_expa_lt_expb), .ZN(n2669) );
  NOR2_X2 U1973 ( .A1(u1_exp_lt_27), .A2(u1_exp_diff_3_), .ZN(n1685) );
  NOR2_X2 U1974 ( .A1(u1_exp_lt_27), .A2(u1_exp_diff_0_), .ZN(n1687) );
  NOR2_X2 U1975 ( .A1(n1680), .A2(n3455), .ZN(n1690) );
  NOR2_X2 U1976 ( .A1(n1685), .A2(n3448), .ZN(n1681) );
  NOR3_X2 U1977 ( .A1(n3462), .A2(n3460), .A3(n3469), .ZN(n1677) );
  AOI222_X1 U1978 ( .A1(n2650), .A2(n1424), .B1(n2473), .B2(n2625), .C1(
        div_opa_ldz_r2[0]), .C2(n1428), .ZN(n1442) );
  NOR2_X2 U1979 ( .A1(n3583), .A2(u4_exp_in_pl1_1_), .ZN(n1440) );
  AOI222_X1 U1980 ( .A1(u4_fi_ldz_2a_3_), .A2(n1431), .B1(u4_div_scht1a[3]), 
        .B2(n1423), .C1(u4_exp_in_pl1_3_), .C2(n1425), .ZN(n1429) );
  NOR3_X2 U1981 ( .A1(exp_ovf_r[1]), .A2(u4_N1733), .A3(n3565), .ZN(n1969) );
  AOI222_X1 U1982 ( .A1(n2682), .A2(n1424), .B1(u4_f2i_shft_2_), .B2(n2625), 
        .C1(div_opa_ldz_r2[2]), .C2(n1428), .ZN(n1433) );
  NOR3_X2 U1983 ( .A1(n2649), .A2(n1443), .A3(n1444), .ZN(n1428) );
  AOI21_X2 U1984 ( .B1(n1437), .B2(n2624), .A(n1448), .ZN(n1447) );
  NAND3_X2 U1985 ( .A1(n2647), .A2(n1449), .A3(n1443), .ZN(n1446) );
  OAI21_X2 U1986 ( .B1(n2233), .B2(n2234), .A(n2235), .ZN(n2230) );
  NOR3_X2 U1987 ( .A1(n2248), .A2(n2129), .A3(n2647), .ZN(n2234) );
  NOR3_X2 U1988 ( .A1(fract_denorm[29]), .A2(fract_denorm[30]), .A3(
        fract_denorm[28]), .ZN(n1551) );
  NAND3_X2 U1989 ( .A1(n1554), .A2(fract_denorm[35]), .A3(n1481), .ZN(n1479)
         );
  NOR3_X2 U1990 ( .A1(fract_denorm[26]), .A2(fract_denorm[27]), .A3(n3541), 
        .ZN(n1488) );
  NOR3_X2 U1991 ( .A1(fract_denorm[21]), .A2(fract_denorm[22]), .A3(n1528), 
        .ZN(n1494) );
  NAND3_X2 U1992 ( .A1(n3523), .A2(n1497), .A3(n1498), .ZN(n1476) );
  NAND3_X2 U1993 ( .A1(n3533), .A2(n1532), .A3(n1533), .ZN(n1496) );
  NOR3_X2 U1994 ( .A1(fract_denorm[45]), .A2(fract_denorm[46]), .A3(n1506), 
        .ZN(n1553) );
  NAND3_X2 U1995 ( .A1(n1552), .A2(fract_denorm[33]), .A3(n1481), .ZN(n1522)
         );
  OAI21_X2 U1996 ( .B1(fract_denorm[37]), .B2(fract_denorm[38]), .A(n1481), 
        .ZN(n1526) );
  NOR3_X2 U1997 ( .A1(n3525), .A2(n3526), .A3(n1478), .ZN(n1535) );
  NOR3_X2 U1998 ( .A1(fract_denorm[24]), .A2(fract_denorm[25]), .A3(n3539), 
        .ZN(n1543) );
  NOR3_X2 U1999 ( .A1(fract_denorm[32]), .A2(fract_denorm[33]), .A3(n3547), 
        .ZN(n1542) );
  NOR3_X2 U2000 ( .A1(n3539), .A2(n3537), .A3(n3503), .ZN(n1520) );
  NAND3_X2 U2001 ( .A1(n1479), .A2(n1516), .A3(n1522), .ZN(n1550) );
  NAND3_X2 U2002 ( .A1(n3521), .A2(n1558), .A3(n1534), .ZN(n1525) );
  AOI21_X2 U2003 ( .B1(n2214), .B2(n2490), .A(n2215), .ZN(n2207) );
  NOR3_X2 U2004 ( .A1(remainder[40]), .A2(remainder[42]), .A3(remainder[41]), 
        .ZN(n2286) );
  NOR3_X2 U2005 ( .A1(remainder[38]), .A2(remainder[3]), .A3(remainder[39]), 
        .ZN(n2285) );
  NOR3_X2 U2006 ( .A1(remainder[35]), .A2(remainder[37]), .A3(remainder[36]), 
        .ZN(n2284) );
  NOR3_X2 U2007 ( .A1(remainder[32]), .A2(remainder[34]), .A3(remainder[33]), 
        .ZN(n2283) );
  NOR3_X2 U2008 ( .A1(remainder[26]), .A2(remainder[28]), .A3(remainder[27]), 
        .ZN(n2297) );
  NOR3_X2 U2009 ( .A1(remainder[20]), .A2(remainder[22]), .A3(remainder[21]), 
        .ZN(n2295) );
  NOR3_X2 U2010 ( .A1(remainder[18]), .A2(remainder[1]), .A3(remainder[19]), 
        .ZN(n2294) );
  NOR3_X2 U2011 ( .A1(remainder[15]), .A2(remainder[17]), .A3(remainder[16]), 
        .ZN(n2293) );
  NOR3_X2 U2012 ( .A1(remainder[12]), .A2(remainder[14]), .A3(remainder[13]), 
        .ZN(n2292) );
  NOR3_X2 U2013 ( .A1(remainder[0]), .A2(remainder[11]), .A3(remainder[10]), 
        .ZN(n2291) );
  NOR3_X2 U2014 ( .A1(remainder[43]), .A2(remainder[45]), .A3(remainder[44]), 
        .ZN(n2287) );
  NOR3_X2 U2015 ( .A1(remainder[46]), .A2(remainder[48]), .A3(remainder[47]), 
        .ZN(n2288) );
  NOR3_X2 U2016 ( .A1(remainder[49]), .A2(remainder[5]), .A3(remainder[4]), 
        .ZN(n2289) );
  NAND3_X2 U2017 ( .A1(n1457), .A2(n1456), .A3(n1458), .ZN(n2246) );
  NAND3_X2 U2018 ( .A1(n1451), .A2(n1450), .A3(n1452), .ZN(n2242) );
  NAND3_X2 U2019 ( .A1(n1460), .A2(n1459), .A3(n1461), .ZN(n2247) );
  OAI21_X2 U2020 ( .B1(n2255), .B2(n2256), .A(n2257), .ZN(n2215) );
  OAI21_X2 U2021 ( .B1(n2258), .B2(n2259), .A(n2243), .ZN(n2257) );
  NOR2_X2 U2022 ( .A1(n2268), .A2(n2269), .ZN(n2255) );
  NAND3_X2 U2023 ( .A1(n1418), .A2(n2492), .A3(n1961), .ZN(n1960) );
  AOI21_X2 U2024 ( .B1(exp_ovf_r[0]), .B2(n3565), .A(n1962), .ZN(n1961) );
  OAI21_X2 U2025 ( .B1(n1967), .B2(n1968), .A(n3580), .ZN(n1965) );
  OAI21_X2 U2026 ( .B1(n1998), .B2(u4_N1598), .A(n3565), .ZN(n1997) );
  NOR2_X2 U2027 ( .A1(n3565), .A2(n1971), .ZN(n1964) );
  AOI222_X1 U2028 ( .A1(u4_N1604), .A2(u4_N1603), .B1(n1972), .B2(n1973), .C1(
        n1974), .C2(n1966), .ZN(n1971) );
  NAND3_X2 U2029 ( .A1(n2545), .A2(n2485), .A3(n2472), .ZN(n1894) );
  AOI21_X2 U2030 ( .B1(n2093), .B2(n2207), .A(n2206), .ZN(n2105) );
  NOR3_X2 U2031 ( .A1(n3517), .A2(n2015), .A3(n1955), .ZN(n2097) );
  OAI21_X2 U2032 ( .B1(n2101), .B2(n1956), .A(n2097), .ZN(n2095) );
  NAND3_X2 U2033 ( .A1(n2097), .A2(n2014), .A3(n2098), .ZN(n2096) );
  NOR3_X2 U2034 ( .A1(n3499), .A2(n3441), .A3(n2099), .ZN(n2098) );
  AOI21_X2 U2035 ( .B1(sign), .B2(rmode_r3[1]), .A(n1949), .ZN(n2099) );
  NOR3_X2 U2036 ( .A1(n2130), .A2(u4_exp_out_0_), .A3(u4_N1640), .ZN(n2127) );
  AOI211_X2 U2037 ( .C1(u4_N1573), .C2(n2018), .A(n2134), .B(n2135), .ZN(n2133) );
  OAI21_X2 U2038 ( .B1(exp_ovf_r[1]), .B2(n2141), .A(n2140), .ZN(n2131) );
  OAI21_X2 U2039 ( .B1(n2174), .B2(n2500), .A(n2204), .ZN(n2159) );
  NOR2_X2 U2040 ( .A1(n1394), .A2(n3520), .ZN(n2160) );
  NOR3_X2 U2041 ( .A1(n3493), .A2(n2200), .A3(n2141), .ZN(n2158) );
  OAI21_X2 U2042 ( .B1(r489_B_0_), .B2(n2172), .A(n2205), .ZN(n2176) );
  NOR3_X2 U2043 ( .A1(n3493), .A2(n2647), .A3(n2201), .ZN(n2157) );
  OAI21_X2 U2044 ( .B1(n2169), .B2(n2170), .A(n2171), .ZN(n2168) );
  NAND3_X2 U2045 ( .A1(n2172), .A2(n2104), .A3(u4_exp_out_pl1_0_), .ZN(n2171)
         );
  NOR3_X2 U2046 ( .A1(n2587), .A2(n2625), .A3(n2141), .ZN(n2169) );
  NOR2_X2 U2047 ( .A1(n2202), .A2(u4_N1532), .ZN(n2153) );
  NOR2_X2 U2048 ( .A1(n3500), .A2(n2202), .ZN(n2154) );
  OAI21_X2 U2049 ( .B1(n2647), .B2(n2128), .A(n2145), .ZN(n2144) );
  OAI21_X2 U2050 ( .B1(n2146), .B2(n2140), .A(n2147), .ZN(n2143) );
  NOR2_X2 U2051 ( .A1(n2465), .A2(n1389), .ZN(n2101) );
  AOI222_X1 U2052 ( .A1(n2647), .A2(opb_inf), .B1(n3518), .B2(opa_00), .C1(
        n2624), .C2(opb_00), .ZN(n2194) );
  NOR2_X2 U2053 ( .A1(rmode_r3[1]), .A2(rmode_r3[0]), .ZN(n2104) );
  INV_X4 U2054 ( .A(n2668), .ZN(n2665) );
  NAND3_X2 U2055 ( .A1(n3451), .A2(n1685), .A3(n3448), .ZN(n1678) );
  NAND3_X2 U2056 ( .A1(n3452), .A2(n1683), .A3(n1693), .ZN(n1692) );
  OAI21_X2 U2057 ( .B1(n1675), .B2(n1690), .A(n1694), .ZN(n1693) );
  NOR2_X2 U2058 ( .A1(u1_exp_lt_27), .A2(u1_exp_diff_1_), .ZN(n1675) );
  OAI21_X2 U2059 ( .B1(n1677), .B2(n1678), .A(n1679), .ZN(n1676) );
  NAND3_X2 U2060 ( .A1(n1680), .A2(n3451), .A3(n1681), .ZN(n1679) );
  OAI21_X2 U2061 ( .B1(n1415), .B2(n2649), .A(n1416), .ZN(u4_shift_right[0])
         );
  AOI222_X1 U2062 ( .A1(u4_div_shft3_0_), .A2(n2626), .B1(n2650), .B2(n1401), 
        .C1(u4_div_shft4[0]), .C2(n1402), .ZN(n1415) );
  OAI21_X2 U2063 ( .B1(n1413), .B2(n2649), .A(n1414), .ZN(u4_shift_right[1])
         );
  AOI222_X1 U2064 ( .A1(u4_div_shft3_1_), .A2(n2626), .B1(n2486), .B2(n1401), 
        .C1(u4_div_shft4[1]), .C2(n1402), .ZN(n1413) );
  AOI222_X1 U2065 ( .A1(u4_fi_ldz_1_), .A2(n1431), .B1(n2681), .B2(n1424), 
        .C1(u4_div_scht1a[1]), .C2(n1423), .ZN(n1434) );
  AOI222_X1 U2066 ( .A1(n2683), .A2(n1424), .B1(u4_f2i_shft_3_), .B2(n2625), 
        .C1(div_opa_ldz_r2[3]), .C2(n1428), .ZN(n1430) );
  NOR2_X2 U2067 ( .A1(n1962), .A2(n3441), .ZN(n1439) );
  AOI211_X2 U2068 ( .C1(n2492), .C2(n2003), .A(n1417), .B(u4_exp_in_mi1_8_), 
        .ZN(n1437) );
  NAND3_X2 U2069 ( .A1(n2465), .A2(n3498), .A3(n2232), .ZN(n1438) );
  AOI222_X1 U2070 ( .A1(n2684), .A2(n1424), .B1(u4_f2i_shft_4_), .B2(n2625), 
        .C1(div_opa_ldz_r2[4]), .C2(n1428), .ZN(n1427) );
  OAI21_X2 U2071 ( .B1(n1411), .B2(n2649), .A(n1412), .ZN(u4_shift_right[2])
         );
  AOI222_X1 U2072 ( .A1(u4_div_shft3_2_), .A2(n2626), .B1(u4_div_shft2[2]), 
        .B2(n1401), .C1(u4_div_shft4[2]), .C2(n1402), .ZN(n1411) );
  OAI21_X2 U2073 ( .B1(sign), .B2(n2211), .A(n2212), .ZN(n2106) );
  AOI21_X2 U2074 ( .B1(n2230), .B2(n3518), .A(n2231), .ZN(n2211) );
  NOR3_X2 U2075 ( .A1(n2216), .A2(opas_r2), .A3(n2687), .ZN(n2213) );
  NOR3_X2 U2076 ( .A1(n3545), .A2(fract_denorm[31]), .A3(n3513), .ZN(n1469) );
  NOR2_X2 U2077 ( .A1(n1531), .A2(n3511), .ZN(n1530) );
  NAND3_X2 U2078 ( .A1(n1503), .A2(n1504), .A3(n1505), .ZN(n1499) );
  NAND3_X2 U2079 ( .A1(n3529), .A2(n1507), .A3(n1508), .ZN(n1503) );
  NAND3_X2 U2080 ( .A1(n1495), .A2(n1496), .A3(n1476), .ZN(n1491) );
  NAND3_X2 U2081 ( .A1(n1546), .A2(n1789), .A3(r524_A_5_), .ZN(n1515) );
  NAND3_X2 U2082 ( .A1(fract_denorm[41]), .A2(n2680), .A3(n1553), .ZN(n1516)
         );
  NOR3_X2 U2083 ( .A1(n1520), .A2(n1493), .A3(n1521), .ZN(n1462) );
  AOI21_X2 U2084 ( .B1(n3542), .B2(n3540), .A(n3503), .ZN(n1521) );
  AOI21_X2 U2085 ( .B1(n1535), .B2(n3562), .A(n1536), .ZN(n1523) );
  NAND3_X2 U2086 ( .A1(n1555), .A2(n2229), .A3(n1513), .ZN(n1478) );
  NOR2_X2 U2087 ( .A1(n1515), .A2(n3560), .ZN(n1508) );
  NAND3_X2 U2088 ( .A1(n1543), .A2(n3543), .A3(n1469), .ZN(n1528) );
  NAND3_X2 U2089 ( .A1(fract_denorm[39]), .A2(n3551), .A3(n1482), .ZN(n1480)
         );
  NAND3_X2 U2090 ( .A1(n1543), .A2(fract_denorm[23]), .A3(n1469), .ZN(n1487)
         );
  NAND3_X2 U2091 ( .A1(n1542), .A2(fract_denorm[31]), .A3(n1481), .ZN(n1468)
         );
  NOR3_X2 U2092 ( .A1(fract_denorm[41]), .A2(n2679), .A3(n3553), .ZN(n1482) );
  NOR3_X2 U2093 ( .A1(n1483), .A2(n3507), .A3(n1518), .ZN(n1548) );
  INV_X4 U2094 ( .A(n2473), .ZN(n2650) );
  INV_X4 U2095 ( .A(n1886), .ZN(n3565) );
  INV_X4 U2096 ( .A(n2486), .ZN(n2681) );
  INV_X4 U2097 ( .A(n2489), .ZN(n2684) );
  INV_X4 U2098 ( .A(n2559), .ZN(n2682) );
  INV_X4 U2099 ( .A(n2488), .ZN(n2683) );
  NOR2_X2 U2100 ( .A1(n1836), .A2(n2597), .ZN(n2028) );
  NOR2_X2 U2101 ( .A1(n3574), .A2(n1830), .ZN(n2032) );
  AOI211_X2 U2102 ( .C1(n2687), .C2(opas_r2), .A(n3504), .B(n1388), .ZN(n2010)
         );
  NOR2_X2 U2103 ( .A1(n2584), .A2(rmode_r3[1]), .ZN(n1949) );
  NOR3_X2 U2104 ( .A1(n2247), .A2(u4_fract_out_10_), .A3(u4_fract_out_0_), 
        .ZN(n2238) );
  NOR2_X2 U2105 ( .A1(n2214), .A2(n2215), .ZN(n2002) );
  NOR3_X2 U2106 ( .A1(n1955), .A2(n1956), .A3(n2648), .ZN(n1954) );
  OAI21_X2 U2107 ( .B1(exp_ovf_r[0]), .B2(n1957), .A(n1958), .ZN(n1953) );
  AOI222_X1 U2108 ( .A1(u4_N1599), .A2(n1963), .B1(n1964), .B2(exp_ovf_r[1]), 
        .C1(n1965), .C2(n1966), .ZN(n1957) );
  NAND3_X2 U2109 ( .A1(n1959), .A2(n2463), .A3(n1960), .ZN(n1958) );
  NAND3_X2 U2110 ( .A1(n1914), .A2(n1915), .A3(n1916), .ZN(n1912) );
  NAND3_X2 U2111 ( .A1(n1869), .A2(n1867), .A3(n1922), .ZN(n1920) );
  NAND3_X2 U2112 ( .A1(n1876), .A2(n1874), .A3(n1924), .ZN(n1923) );
  NAND3_X2 U2113 ( .A1(n1862), .A2(n1860), .A3(n1919), .ZN(n1917) );
  NAND3_X2 U2114 ( .A1(n2534), .A2(n2484), .A3(n2464), .ZN(n1902) );
  NAND3_X2 U2115 ( .A1(n2544), .A2(n2483), .A3(n2471), .ZN(n1904) );
  NOR2_X2 U2116 ( .A1(opb_dn), .A2(opa_dn), .ZN(n1886) );
  NAND3_X2 U2117 ( .A1(n1867), .A2(n1868), .A3(n1869), .ZN(n1863) );
  NAND3_X2 U2118 ( .A1(n1874), .A2(n1875), .A3(n1876), .ZN(n1870) );
  NAND3_X2 U2119 ( .A1(n1860), .A2(n1861), .A3(n1862), .ZN(n1856) );
  NOR2_X2 U2120 ( .A1(opb_inf), .A2(opa_inf), .ZN(n1832) );
  NOR3_X2 U2121 ( .A1(n2625), .A2(n1949), .A3(n1854), .ZN(n2015) );
  NOR3_X2 U2122 ( .A1(u4_N1640), .A2(u4_exp_out_mi1[0]), .A3(n2130), .ZN(n2014) );
  NOR3_X2 U2123 ( .A1(n2558), .A2(n1886), .A3(n2141), .ZN(n2018) );
  AOI21_X2 U2124 ( .B1(exp_ovf_r[0]), .B2(n2014), .A(n1955), .ZN(n2019) );
  NOR2_X2 U2125 ( .A1(n2579), .A2(n2492), .ZN(n2017) );
  OAI21_X2 U2126 ( .B1(n2124), .B2(n2649), .A(n2125), .ZN(n1956) );
  AOI21_X2 U2127 ( .B1(n1949), .B2(n2131), .A(n2132), .ZN(n2124) );
  AOI222_X1 U2128 ( .A1(u4_exp_out_3_), .A2(n2159), .B1(u4_exp_out_mi1[3]), 
        .B2(n2160), .C1(u4_exp_out_pl1_3_), .C2(n2161), .ZN(n2196) );
  AOI222_X1 U2129 ( .A1(u4_exp_out_2_), .A2(n2159), .B1(u4_exp_out_mi1[2]), 
        .B2(n2160), .C1(u4_exp_out_pl1_2_), .C2(n2161), .ZN(n2151) );
  AOI222_X1 U2130 ( .A1(u4_exp_out_1_), .A2(n2159), .B1(u4_exp_out_mi1[1]), 
        .B2(n2160), .C1(u4_exp_out_pl1_1_), .C2(n2161), .ZN(n2162) );
  AOI222_X1 U2131 ( .A1(n2159), .A2(u4_N1976), .B1(u4_exp_out_mi1[7]), .B2(
        n2160), .C1(u4_exp_out_pl1_7_), .C2(n2161), .ZN(n2177) );
  AOI222_X1 U2132 ( .A1(u4_exp_out_6_), .A2(n2159), .B1(u4_exp_out_mi1[6]), 
        .B2(n2160), .C1(u4_exp_out_pl1_6_), .C2(n2161), .ZN(n2181) );
  AOI222_X1 U2133 ( .A1(u4_exp_out_5_), .A2(n2159), .B1(u4_exp_out_mi1[5]), 
        .B2(n2160), .C1(u4_exp_out_pl1_5_), .C2(n2161), .ZN(n2185) );
  AOI222_X1 U2134 ( .A1(u4_exp_out_4_), .A2(n2159), .B1(u4_exp_out_mi1[4]), 
        .B2(n2160), .C1(u4_exp_out_pl1_4_), .C2(n2161), .ZN(n2189) );
  AOI222_X1 U2135 ( .A1(n2157), .A2(u4_exp_next_mi_0_), .B1(n2158), .B2(n2650), 
        .C1(n2176), .C2(u4_exp_out_0_), .ZN(n2166) );
  AOI211_X2 U2136 ( .C1(n2647), .C2(n3491), .A(n2101), .B(n1955), .ZN(n2119)
         );
  NAND3_X2 U2137 ( .A1(exp_ovf_r[1]), .A2(n2579), .A3(n2647), .ZN(n2195) );
  NOR2_X2 U2138 ( .A1(n2431), .A2(fpu_op_r2[1]), .ZN(n2394) );
  INV_X4 U2139 ( .A(n2665), .ZN(n2663) );
  INV_X4 U2140 ( .A(n2660), .ZN(n2654) );
  INV_X4 U2141 ( .A(n2665), .ZN(n2662) );
  OAI21_X2 U2142 ( .B1(u1_exp_diff_sft_4_), .B2(n1672), .A(n3446), .ZN(n1671)
         );
  OAI21_X2 U2143 ( .B1(n1691), .B2(n1678), .A(n1692), .ZN(n1673) );
  NOR2_X2 U2144 ( .A1(fasu_op_r2), .A2(n2602), .ZN(n1844) );
  NOR3_X2 U2145 ( .A1(n1746), .A2(fracta_mul[10]), .A3(fracta_mul[0]), .ZN(
        n1742) );
  NAND3_X2 U2146 ( .A1(n2583), .A2(n2499), .A3(n2479), .ZN(n1755) );
  NAND3_X2 U2147 ( .A1(n2437), .A2(n2588), .A3(n2444), .ZN(n1746) );
  NOR3_X2 U2148 ( .A1(fracta_mul[13]), .A2(fracta_mul[9]), .A3(fracta_mul[7]), 
        .ZN(n2444) );
  NOR2_X2 U2149 ( .A1(fracta_mul[9]), .A2(fracta_mul[8]), .ZN(n2451) );
  OAI21_X2 U2150 ( .B1(n1409), .B2(n2649), .A(n1410), .ZN(u4_shift_right[3])
         );
  AOI222_X1 U2151 ( .A1(u4_div_shft3_3_), .A2(n2626), .B1(u4_div_shft2[3]), 
        .B2(n1401), .C1(u4_div_shft4[3]), .C2(n1402), .ZN(n1409) );
  OAI21_X2 U2152 ( .B1(n1407), .B2(n2649), .A(n1408), .ZN(u4_shift_right[4])
         );
  AOI222_X1 U2153 ( .A1(u4_div_shft3_4_), .A2(n2626), .B1(u4_div_shft2[4]), 
        .B2(n1401), .C1(u4_div_shft4[4]), .C2(n1402), .ZN(n1407) );
  NOR2_X2 U2154 ( .A1(n2687), .A2(n2686), .ZN(n1970) );
  NOR2_X2 U2155 ( .A1(n1449), .A2(n2649), .ZN(n1424) );
  NOR3_X2 U2156 ( .A1(n1443), .A2(n3583), .A3(n2648), .ZN(n1423) );
  OAI21_X2 U2157 ( .B1(n1437), .B2(n2474), .A(n2305), .ZN(n1425) );
  AOI222_X1 U2158 ( .A1(u4_div_scht1a[5]), .A2(n1423), .B1(u4_f2i_shft_5_), 
        .B2(n2625), .C1(n2685), .C2(n1424), .ZN(n1422) );
  NOR2_X2 U2159 ( .A1(n2624), .A2(n2647), .ZN(n2232) );
  NOR2_X2 U2160 ( .A1(n2625), .A2(n2647), .ZN(n2100) );
  NOR3_X2 U2161 ( .A1(fpu_op_r3[0]), .A2(fpu_op_r3[1]), .A3(n2491), .ZN(n1448)
         );
  INV_X4 U2162 ( .A(n2487), .ZN(n2685) );
  NAND3_X2 U2163 ( .A1(n3565), .A2(n1444), .A3(n2568), .ZN(n1418) );
  OAI21_X2 U2164 ( .B1(n1363), .B2(n1988), .A(n1989), .ZN(n1975) );
  AOI222_X1 U2165 ( .A1(u4_div_exp1_7_), .A2(opb_dn), .B1(u4_exp_out1_mi1[7]), 
        .B2(n1366), .C1(u4_div_exp2_7_), .C2(n1367), .ZN(n1988) );
  AOI21_X2 U2166 ( .B1(n1469), .B2(fract_denorm[28]), .A(n1470), .ZN(n1463) );
  NOR3_X2 U2167 ( .A1(n1474), .A2(n1475), .A3(n3505), .ZN(n1473) );
  NOR3_X2 U2168 ( .A1(n1511), .A2(n1512), .A3(n3506), .ZN(n1510) );
  AOI21_X2 U2169 ( .B1(n1517), .B2(n2680), .A(n1518), .ZN(n1509) );
  OAI21_X2 U2170 ( .B1(n1514), .B2(n1515), .A(n1516), .ZN(n1511) );
  INV_X4 U2171 ( .A(n2680), .ZN(n2679) );
  NOR3_X2 U2172 ( .A1(n1420), .A2(n3532), .A3(n1546), .ZN(n1545) );
  NOR3_X2 U2173 ( .A1(n3503), .A2(fract_denorm[30]), .A3(n3540), .ZN(n1544) );
  NOR3_X2 U2174 ( .A1(n1541), .A2(n3526), .A3(n1478), .ZN(n1475) );
  NOR3_X2 U2175 ( .A1(n3535), .A2(fract_denorm[22]), .A3(n1528), .ZN(n1531) );
  NOR3_X2 U2176 ( .A1(fract_denorm[39]), .A2(fract_denorm[40]), .A3(n3515), 
        .ZN(n1481) );
  OAI21_X2 U2177 ( .B1(fract_denorm[44]), .B2(n3555), .A(n3552), .ZN(n1561) );
  NOR2_X2 U2178 ( .A1(fract_denorm[38]), .A2(n3548), .ZN(n1560) );
  NOR3_X2 U2179 ( .A1(u4_N1504), .A2(u4_N1503), .A3(n2562), .ZN(n1367) );
  NOR2_X2 U2180 ( .A1(n3565), .A2(n1417), .ZN(n1366) );
  NOR2_X2 U2181 ( .A1(n3575), .A2(n2474), .ZN(n2022) );
  NOR2_X2 U2182 ( .A1(n1948), .A2(n2597), .ZN(n2033) );
  NOR2_X2 U2183 ( .A1(n3575), .A2(n2649), .ZN(n1833) );
  NOR2_X2 U2184 ( .A1(n2465), .A2(n1830), .ZN(n1828) );
  NOR3_X2 U2185 ( .A1(n1959), .A2(n2009), .A3(n2010), .ZN(n2005) );
  NAND3_X2 U2186 ( .A1(n1935), .A2(n1940), .A3(n1878), .ZN(n1943) );
  AOI21_X2 U2187 ( .B1(n1949), .B2(n3578), .A(n1943), .ZN(n1945) );
  NOR3_X2 U2188 ( .A1(n1923), .A2(n1873), .A3(n1871), .ZN(n1908) );
  NOR2_X2 U2189 ( .A1(qnan_d), .A2(snan_d), .ZN(n1829) );
  NOR3_X2 U2190 ( .A1(n1885), .A2(n1886), .A3(n1830), .ZN(n1884) );
  OAI21_X2 U2191 ( .B1(n1887), .B2(n1888), .A(sign), .ZN(n1885) );
  NAND3_X2 U2192 ( .A1(n2624), .A2(n1947), .A3(n1948), .ZN(n1842) );
  OAI21_X2 U2193 ( .B1(r489_B_0_), .B2(n1933), .A(n1832), .ZN(n1947) );
  NAND3_X2 U2194 ( .A1(n3577), .A2(n2532), .A3(inf_d), .ZN(n1843) );
  INV_X4 U2195 ( .A(n2049), .ZN(n3490) );
  NOR2_X2 U2196 ( .A1(n3575), .A2(inf_d), .ZN(n1936) );
  AOI21_X2 U2197 ( .B1(n2014), .B2(n2008), .A(n2015), .ZN(n2013) );
  NOR2_X2 U2198 ( .A1(inf_mul_r), .A2(inf_mul2), .ZN(n1933) );
  NOR2_X2 U2199 ( .A1(n3574), .A2(opb_00), .ZN(n1938) );
  AOI21_X2 U2200 ( .B1(n2122), .B2(n2111), .A(n2112), .ZN(n1929) );
  AOI21_X2 U2201 ( .B1(n2121), .B2(n2111), .A(n2112), .ZN(n1930) );
  AOI21_X2 U2202 ( .B1(n2120), .B2(n2111), .A(n2112), .ZN(n1931) );
  AOI21_X2 U2203 ( .B1(n2115), .B2(n2111), .A(n2112), .ZN(n1925) );
  AOI21_X2 U2204 ( .B1(n2114), .B2(n2111), .A(n2112), .ZN(n1926) );
  AOI21_X2 U2205 ( .B1(n2113), .B2(n2111), .A(n2112), .ZN(n1927) );
  AOI21_X2 U2206 ( .B1(n2110), .B2(n2111), .A(n2112), .ZN(n1928) );
  OAI21_X2 U2207 ( .B1(n2117), .B2(n2118), .A(n2119), .ZN(n2116) );
  NAND2_X2 U2208 ( .A1(n2388), .A2(n3498), .ZN(n2049) );
  AOI211_X2 U2209 ( .C1(inf_d), .C2(n2100), .A(n1838), .B(n2390), .ZN(n2389)
         );
  NOR3_X2 U2210 ( .A1(n2474), .A2(r489_B_0_), .A3(n1933), .ZN(n2390) );
  NOR2_X2 U2211 ( .A1(fpu_op_r2[1]), .A2(fpu_op_r2[2]), .ZN(n2426) );
  NOR3_X2 U2212 ( .A1(n1573), .A2(n2634), .A3(n3399), .ZN(n1600) );
  NOR3_X2 U2213 ( .A1(n1590), .A2(n1573), .A3(n3494), .ZN(n1599) );
  NOR2_X2 U2214 ( .A1(n3399), .A2(n3479), .ZN(n1598) );
  NOR2_X2 U2215 ( .A1(u2_exp_ovf_d_1_), .A2(n1573), .ZN(n1597) );
  NOR3_X2 U2216 ( .A1(n3411), .A2(u2_N22), .A3(n2634), .ZN(n1567) );
  NOR3_X2 U2217 ( .A1(n3404), .A2(u2_N13), .A3(n3494), .ZN(n1565) );
  NOR2_X2 U2218 ( .A1(opb_r[30]), .A2(opa_r[30]), .ZN(n1570) );
  NOR2_X2 U2219 ( .A1(n3485), .A2(n2653), .ZN(n1573) );
  INV_X4 U2220 ( .A(n1569), .ZN(n3494) );
  NAND3_X2 U2221 ( .A1(n2394), .A2(n3497), .A3(N251), .ZN(n2620) );
  NAND3_X2 U2222 ( .A1(n2394), .A2(n3497), .A3(N251), .ZN(n2393) );
  INV_X4 U2223 ( .A(fasu_op), .ZN(n2689) );
  INV_X4 U2224 ( .A(n2674), .ZN(n2672) );
  INV_X4 U2225 ( .A(n2674), .ZN(n2673) );
  INV_X4 U2226 ( .A(n2674), .ZN(n2671) );
  NOR2_X2 U2227 ( .A1(u1_fracta_eq_fractb), .A2(n1725), .ZN(n1726) );
  AOI211_X2 U2228 ( .C1(n2647), .C2(n3566), .A(n1844), .B(n2391), .ZN(n1877)
         );
  OAI21_X2 U2229 ( .B1(n2474), .B2(n1948), .A(n1829), .ZN(n2391) );
  AOI21_X2 U2230 ( .B1(fracta_mul[16]), .B2(n2581), .A(fracta_mul[18]), .ZN(
        n2440) );
  AOI21_X2 U2231 ( .B1(n2591), .B2(n3483), .A(fracta_mul[5]), .ZN(n2443) );
  AOI21_X2 U2232 ( .B1(n2502), .B2(fracta_mul[1]), .A(fracta_mul[3]), .ZN(
        n2445) );
  OAI21_X2 U2233 ( .B1(fracta_mul[13]), .B2(n2441), .A(n2501), .ZN(n2438) );
  AOI21_X2 U2234 ( .B1(n2442), .B2(n2588), .A(fracta_mul[12]), .ZN(n2441) );
  OAI21_X2 U2235 ( .B1(fracta_mul[9]), .B2(n2593), .A(n2497), .ZN(n2442) );
  AOI211_X2 U2236 ( .C1(n2502), .C2(n2592), .A(fracta_mul[5]), .B(
        fracta_mul[4]), .ZN(n2453) );
  NAND3_X2 U2237 ( .A1(n2497), .A2(n2588), .A3(n2451), .ZN(n2050) );
  NAND3_X2 U2238 ( .A1(n2589), .A2(n2462), .A3(n2498), .ZN(n2052) );
  NOR3_X2 U2239 ( .A1(n2050), .A2(fracta_mul[12]), .A3(n2051), .ZN(n1818) );
  OAI21_X2 U2240 ( .B1(n1405), .B2(n2649), .A(n1406), .ZN(u4_shift_right[5])
         );
  AOI222_X1 U2241 ( .A1(u4_div_shft3_5_), .A2(n2626), .B1(u4_div_shft2[5]), 
        .B2(n1401), .C1(u4_div_shft4[5]), .C2(n1402), .ZN(n1405) );
  AOI222_X1 U2242 ( .A1(n2625), .A2(n2302), .B1(n1423), .B2(n2303), .C1(n2304), 
        .C2(n1425), .ZN(n2301) );
  OAI21_X2 U2243 ( .B1(n2647), .B2(n2385), .A(n2386), .ZN(n2300) );
  NOR2_X2 U2244 ( .A1(u4_exp_in_mi1_8_), .A2(n3520), .ZN(n2385) );
  OAI21_X2 U2245 ( .B1(exp_ovf_r[0]), .B2(n1401), .A(n2492), .ZN(n2386) );
  NOR2_X2 U2246 ( .A1(n1444), .A2(exp_ovf_r[1]), .ZN(n1417) );
  OAI21_X2 U2247 ( .B1(n2679), .B2(n3443), .A(n1444), .ZN(n2306) );
  OAI21_X2 U2248 ( .B1(n2679), .B2(n3443), .A(n2307), .ZN(n1393) );
  NOR2_X2 U2249 ( .A1(n2492), .A2(n2474), .ZN(n1395) );
  OAI21_X2 U2250 ( .B1(opb_dn), .B2(n2537), .A(n1784), .ZN(fract_div_47_) );
  INV_X4 U2251 ( .A(n2560), .ZN(n2686) );
  INV_X4 U2252 ( .A(n2558), .ZN(n2687) );
  NOR2_X2 U2253 ( .A1(n1418), .A2(n2626), .ZN(n1402) );
  OAI21_X2 U2254 ( .B1(n1363), .B2(n1991), .A(n1992), .ZN(n1990) );
  AOI222_X1 U2255 ( .A1(u4_div_exp1_6_), .A2(opb_dn), .B1(u4_exp_out1_mi1[6]), 
        .B2(n1366), .C1(u4_div_exp2_6_), .C2(n1367), .ZN(n1991) );
  OAI21_X2 U2256 ( .B1(n1363), .B2(n1994), .A(n1995), .ZN(n1993) );
  AOI222_X1 U2257 ( .A1(u4_div_exp1_5_), .A2(opb_dn), .B1(u4_exp_out1_mi1[5]), 
        .B2(n1366), .C1(u4_div_exp2_5_), .C2(n1367), .ZN(n1994) );
  OAI21_X2 U2258 ( .B1(n1363), .B2(n1977), .A(n1978), .ZN(n1976) );
  AOI222_X1 U2259 ( .A1(u4_div_exp1_4_), .A2(opb_dn), .B1(u4_exp_out1_mi1[4]), 
        .B2(n1366), .C1(u4_div_exp2_4_), .C2(n1367), .ZN(n1977) );
  OAI21_X2 U2260 ( .B1(n1363), .B2(n1980), .A(n1981), .ZN(n1979) );
  AOI222_X1 U2261 ( .A1(u4_div_exp1_3_), .A2(opb_dn), .B1(u4_exp_out1_mi1[3]), 
        .B2(n1366), .C1(u4_div_exp2_3_), .C2(n1367), .ZN(n1980) );
  OAI21_X2 U2262 ( .B1(n1363), .B2(n1983), .A(n1984), .ZN(n1982) );
  AOI222_X1 U2263 ( .A1(u4_div_exp1_2_), .A2(opb_dn), .B1(u4_exp_out1_mi1[2]), 
        .B2(n1366), .C1(u4_div_exp2_2_), .C2(n1367), .ZN(n1983) );
  OAI21_X2 U2264 ( .B1(n1363), .B2(n1986), .A(n1987), .ZN(n1985) );
  AOI222_X1 U2265 ( .A1(u4_div_exp1_1_), .A2(opb_dn), .B1(u4_exp_out1_mi1[1]), 
        .B2(n1366), .C1(u4_div_exp2_1_), .C2(n1367), .ZN(n1986) );
  NOR3_X2 U2266 ( .A1(n2567), .A2(n3498), .A3(n1386), .ZN(n1372) );
  NAND3_X2 U2267 ( .A1(n2625), .A2(n1388), .A3(n1389), .ZN(n1355) );
  NOR2_X2 U2268 ( .A1(n3554), .A2(n1368), .ZN(n1360) );
  NOR3_X2 U2269 ( .A1(n1544), .A2(n1536), .A3(n1545), .ZN(n1538) );
  NOR2_X2 U2270 ( .A1(n3504), .A2(n3498), .ZN(n1359) );
  INV_X4 U2271 ( .A(n2648), .ZN(n2647) );
  OAI21_X2 U2272 ( .B1(n1363), .B2(n1364), .A(n1365), .ZN(n1362) );
  AOI222_X1 U2273 ( .A1(u4_div_exp1_0_), .A2(opb_dn), .B1(n1356), .B2(n1366), 
        .C1(u4_div_exp2_0_), .C2(n1367), .ZN(n1364) );
  OAI21_X2 U2274 ( .B1(n1828), .B2(n2020), .A(n2021), .ZN(N495) );
  OAI21_X2 U2275 ( .B1(n1827), .B2(n1828), .A(n1829), .ZN(n1826) );
  OAI21_X2 U2276 ( .B1(opb_00), .B2(n1830), .A(n2598), .ZN(n1834) );
  NAND3_X2 U2277 ( .A1(n1942), .A2(n1943), .A3(n1936), .ZN(n1941) );
  AOI21_X2 U2278 ( .B1(n1945), .B2(n1946), .A(opa_00), .ZN(n1944) );
  OAI21_X2 U2279 ( .B1(n1905), .B2(n1906), .A(n1907), .ZN(n1881) );
  NOR3_X2 U2280 ( .A1(n3575), .A2(n2690), .A3(n1837), .ZN(N526) );
  AOI211_X2 U2281 ( .C1(n1838), .C2(n2596), .A(n1839), .B(n1840), .ZN(n1837)
         );
  NOR3_X2 U2282 ( .A1(n2503), .A2(opb_inf), .A3(n2648), .ZN(n1840) );
  NAND3_X2 U2283 ( .A1(n1841), .A2(n1842), .A3(n1843), .ZN(n1839) );
  NOR2_X2 U2284 ( .A1(n3490), .A2(n1914), .ZN(N446) );
  NOR2_X2 U2285 ( .A1(n3490), .A2(n1916), .ZN(N447) );
  NOR2_X2 U2286 ( .A1(n3490), .A2(n2045), .ZN(N448) );
  NOR2_X2 U2287 ( .A1(n3490), .A2(n2044), .ZN(N449) );
  NOR2_X2 U2288 ( .A1(n3490), .A2(n1861), .ZN(N450) );
  NOR2_X2 U2289 ( .A1(n3490), .A2(n1860), .ZN(N451) );
  NOR2_X2 U2290 ( .A1(n3490), .A2(n1862), .ZN(N452) );
  NOR2_X2 U2291 ( .A1(n3490), .A2(n1919), .ZN(N453) );
  NOR2_X2 U2292 ( .A1(n3490), .A2(n2043), .ZN(N454) );
  NOR2_X2 U2293 ( .A1(n3490), .A2(n2042), .ZN(N455) );
  NOR2_X2 U2294 ( .A1(n3490), .A2(n1868), .ZN(N456) );
  NOR2_X2 U2295 ( .A1(n3490), .A2(n1867), .ZN(N457) );
  NOR2_X2 U2296 ( .A1(n3490), .A2(n1869), .ZN(N458) );
  NOR2_X2 U2297 ( .A1(n3490), .A2(n1922), .ZN(N459) );
  NOR2_X2 U2298 ( .A1(n3490), .A2(n1875), .ZN(N462) );
  NOR2_X2 U2299 ( .A1(n3490), .A2(n1874), .ZN(N463) );
  NOR2_X2 U2300 ( .A1(n3490), .A2(n1876), .ZN(N464) );
  NOR2_X2 U2301 ( .A1(n3490), .A2(n1924), .ZN(N465) );
  AOI21_X2 U2302 ( .B1(n1936), .B2(n1937), .A(n1938), .ZN(n1934) );
  NOR2_X2 U2303 ( .A1(n1821), .A2(n1822), .ZN(N540) );
  NAND3_X2 U2304 ( .A1(n3400), .A2(n3494), .A3(n1570), .ZN(n1615) );
  AOI21_X2 U2305 ( .B1(n1588), .B2(n1589), .A(n2461), .ZN(u2_exp_ovf_d_0_) );
  AOI21_X2 U2306 ( .B1(n1562), .B2(n1563), .A(n1564), .ZN(u2_underflow_d[2])
         );
  OAI21_X2 U2307 ( .B1(n3494), .B2(n1591), .A(n1592), .ZN(u2_N90) );
  OAI21_X2 U2308 ( .B1(n2469), .B2(n2504), .A(n2403), .ZN(N391) );
  OAI21_X2 U2309 ( .B1(n2469), .B2(n2603), .A(n2402), .ZN(N392) );
  NOR2_X2 U2310 ( .A1(n1720), .A2(n1699), .ZN(u1_N44) );
  NOR2_X2 U2311 ( .A1(n1720), .A2(n1700), .ZN(u1_N43) );
  NOR2_X2 U2312 ( .A1(n1720), .A2(n1701), .ZN(u1_N42) );
  NOR2_X2 U2313 ( .A1(n1720), .A2(n1702), .ZN(u1_N41) );
  NOR2_X2 U2314 ( .A1(n1720), .A2(n1703), .ZN(u1_N40) );
  NOR2_X2 U2315 ( .A1(n1720), .A2(n1704), .ZN(u1_N39) );
  NOR2_X2 U2316 ( .A1(n1720), .A2(n1705), .ZN(u1_N38) );
  NOR2_X2 U2317 ( .A1(n1720), .A2(n1706), .ZN(u1_N37) );
  OAI21_X2 U2318 ( .B1(n1722), .B2(n2600), .A(n1723), .ZN(u1_N140) );
  OAI21_X2 U2319 ( .B1(n1724), .B2(n2605), .A(u1_signa_r), .ZN(n1723) );
  NOR3_X2 U2320 ( .A1(n1725), .A2(u1_fracta_lt_fractb), .A3(
        u1_fracta_eq_fractb), .ZN(n1724) );
  NOR2_X2 U2321 ( .A1(n2690), .A2(n1877), .ZN(N524) );
  NOR2_X2 U2322 ( .A1(n1733), .A2(n1732), .ZN(u0_N6) );
  NOR2_X2 U2323 ( .A1(fracta_mul[22]), .A2(n1735), .ZN(u0_N4) );
  NOR2_X2 U2324 ( .A1(u6_N22), .A2(n1734), .ZN(u0_N5) );
  NOR3_X2 U2325 ( .A1(n2606), .A2(opa_nan), .A3(n1823), .ZN(N532) );
  NOR2_X2 U2326 ( .A1(n3480), .A2(n1737), .ZN(u0_N10) );
  NOR2_X2 U2327 ( .A1(n3486), .A2(n1736), .ZN(u0_N11) );
  NAND3_X2 U2328 ( .A1(n2435), .A2(n2462), .A3(n2436), .ZN(N170) );
  OAI21_X2 U2329 ( .B1(n2443), .B2(fracta_mul[6]), .A(n3481), .ZN(n2435) );
  OAI21_X2 U2330 ( .B1(fracta_mul[19]), .B2(n2440), .A(n2498), .ZN(n2439) );
  NAND3_X2 U2331 ( .A1(n2580), .A2(n2462), .A3(n2496), .ZN(n2447) );
  NOR2_X2 U2332 ( .A1(n2455), .A2(n2052), .ZN(N107) );
  OAI21_X2 U2333 ( .B1(n2458), .B2(n2050), .A(n2590), .ZN(n2457) );
  NOR2_X2 U2334 ( .A1(n3580), .A2(n2647), .ZN(n1399) );
  NOR2_X2 U2335 ( .A1(n2490), .A2(n1417), .ZN(n1398) );
  NAND3_X2 U2336 ( .A1(n1390), .A2(n3498), .A3(n1391), .ZN(n1368) );
  AOI21_X2 U2337 ( .B1(n2624), .B2(n1393), .A(n3499), .ZN(n1391) );
  NAND3_X2 U2338 ( .A1(n1394), .A2(n2579), .A3(n1395), .ZN(n1390) );
  OAI21_X2 U2339 ( .B1(n1403), .B2(n2649), .A(n1404), .ZN(u4_shift_right[6])
         );
  AOI222_X1 U2340 ( .A1(u4_div_shft3_6_), .A2(n2626), .B1(u4_div_shft2[6]), 
        .B2(n1401), .C1(u4_div_shft4[6]), .C2(n1402), .ZN(n1403) );
  OAI21_X2 U2341 ( .B1(n1396), .B2(n2649), .A(n1397), .ZN(u4_shift_right[7])
         );
  AOI222_X1 U2342 ( .A1(u4_div_shft3_7_), .A2(n2626), .B1(u4_div_shft2[7]), 
        .B2(n1401), .C1(u4_div_shft4[7]), .C2(n1402), .ZN(n1396) );
  AOI222_X1 U2343 ( .A1(u4_N1471), .A2(n1359), .B1(n1360), .B2(n3441), .C1(
        n2647), .C2(n1362), .ZN(n1358) );
  NOR3_X2 U2344 ( .A1(u4_N1370), .A2(u4_N1372), .A3(u4_N1371), .ZN(n2264) );
  NOR3_X2 U2345 ( .A1(u4_N1373), .A2(u4_N1375), .A3(u4_N1374), .ZN(n2265) );
  NOR3_X2 U2346 ( .A1(u4_N1376), .A2(u4_N1378), .A3(u4_N1377), .ZN(n2266) );
  NOR3_X2 U2347 ( .A1(u4_N1379), .A2(u4_N1381), .A3(u4_N1380), .ZN(n2267) );
  NOR3_X2 U2348 ( .A1(u4_N1358), .A2(u4_N1360), .A3(u4_N1359), .ZN(n2260) );
  NOR3_X2 U2349 ( .A1(u4_N1361), .A2(u4_N1363), .A3(u4_N1362), .ZN(n2261) );
  NOR3_X2 U2350 ( .A1(u4_N1364), .A2(u4_N1366), .A3(u4_N1365), .ZN(n2262) );
  NOR3_X2 U2351 ( .A1(u4_N1367), .A2(u4_N1369), .A3(u4_N1368), .ZN(n2263) );
  NAND3_X2 U2352 ( .A1(n1454), .A2(n1453), .A3(n1455), .ZN(n2245) );
  INV_X4 U2353 ( .A(n2533), .ZN(n2622) );
  INV_X4 U2354 ( .A(n2677), .ZN(n2676) );
  INV_X4 U2355 ( .A(n2668), .ZN(n2666) );
  INV_X4 U2356 ( .A(n2666), .ZN(n2661) );
  NOR3_X2 U2357 ( .A1(n2468), .A2(fpu_op_r1[2]), .A3(n2595), .ZN(n1569) );
  INV_X4 U2358 ( .A(n2533), .ZN(n2623) );
  OR3_X4 U2359 ( .A1(n2475), .A2(fpu_op_r3[1]), .A3(n2491), .ZN(n2465) );
  INV_X4 U2360 ( .A(u1_fractb_lt_fracta), .ZN(n2678) );
  INV_X4 U2361 ( .A(n2667), .ZN(n2659) );
  NAND2_X4 U2362 ( .A1(n2405), .A2(n3496), .ZN(n2469) );
  INV_X4 U2363 ( .A(n2309), .ZN(n2645) );
  INV_X4 U2364 ( .A(n2645), .ZN(n2643) );
  INV_X4 U2365 ( .A(n2623), .ZN(n2638) );
  OR2_X4 U2366 ( .A1(n2638), .A2(n2690), .ZN(n2474) );
  INV_X4 U2367 ( .A(n2490), .ZN(n2649) );
  INV_X4 U2368 ( .A(u1_fractb_lt_fracta), .ZN(n2675) );
  INV_X4 U2369 ( .A(n2675), .ZN(n2670) );
  INV_X4 U2370 ( .A(n2652), .ZN(n2651) );
  INV_X4 U2371 ( .A(n2651), .ZN(n2653) );
  INV_X4 U2372 ( .A(u2_N124), .ZN(n2652) );
  INV_X4 U2373 ( .A(n2664), .ZN(n2656) );
  OR2_X4 U2374 ( .A1(n1587), .A2(u2_exp_tmp4_0_), .ZN(n2480) );
  INV_X4 U2375 ( .A(n2633), .ZN(n2635) );
  AND2_X4 U2376 ( .A1(n2097), .A2(n2107), .ZN(n2482) );
  NOR2_X2 U2377 ( .A1(n1937), .A2(opb_dn), .ZN(n2320) );
  NOR2_X2 U2378 ( .A1(n2463), .A2(n1937), .ZN(n2309) );
  INV_X4 U2379 ( .A(n2533), .ZN(n2621) );
  NAND4_X2 U2380 ( .A1(n1537), .A2(n3501), .A3(n1538), .A4(n1539), .ZN(
        u4_N1471) );
  INV_X4 U2381 ( .A(fract_denorm[47]), .ZN(n2680) );
  NOR2_X2 U2382 ( .A1(n1937), .A2(n2690), .ZN(n2490) );
  OR2_X4 U2383 ( .A1(n2492), .A2(n1886), .ZN(n2493) );
  INV_X4 U2384 ( .A(n2666), .ZN(n2660) );
  INV_X4 U2385 ( .A(n2664), .ZN(n2655) );
  INV_X4 U2386 ( .A(n1569), .ZN(n2633) );
  INV_X4 U2387 ( .A(n2633), .ZN(n2634) );
  INV_X4 U2388 ( .A(n2470), .ZN(n2688) );
  OR2_X4 U2389 ( .A1(n3496), .A2(n3497), .ZN(n2511) );
  NOR2_X2 U2390 ( .A1(n2394), .A2(n2405), .ZN(n2530) );
  NOR2_X2 U2391 ( .A1(n3496), .A2(n2405), .ZN(n2397) );
  OR2_X4 U2392 ( .A1(u4_exp_out_1_), .A2(u4_exp_out_0_), .ZN(n2531) );
  OR2_X4 U2393 ( .A1(n2532), .A2(fpu_op_r3[0]), .ZN(n2533) );
  INV_X4 U2394 ( .A(n2482), .ZN(n2628) );
  INV_X4 U2395 ( .A(n2482), .ZN(n2627) );
  OR2_X4 U2396 ( .A1(u4_exp_out1_1_), .A2(u4_sub_465_A_0_), .ZN(n2535) );
  OR2_X4 U2397 ( .A1(n2713), .A2(u4_fi_ldz_2_), .ZN(n2536) );
  INV_X4 U2398 ( .A(n2057), .ZN(n2629) );
  NOR2_X2 U2399 ( .A1(n2102), .A2(n2103), .ZN(n2057) );
  INV_X4 U2400 ( .A(n2629), .ZN(n2630) );
  NOR2_X2 U2401 ( .A1(fpu_op_r3[1]), .A2(n2460), .ZN(n1942) );
  NAND2_X2 U2402 ( .A1(u4_sub_488_carry[5]), .A2(n1420), .ZN(n2543) );
  NAND4_X2 U2403 ( .A1(n1471), .A2(n3510), .A3(n1472), .A4(n1473), .ZN(
        u4_fi_ldz_2a_3_) );
  INV_X4 U2404 ( .A(n2645), .ZN(n2644) );
  NOR2_X2 U2405 ( .A1(u4_N1356), .A2(n2300), .ZN(n2243) );
  INV_X4 U2406 ( .A(n2491), .ZN(n2690) );
  INV_X4 U2407 ( .A(n2256), .ZN(n2646) );
  NAND2_X2 U2408 ( .A1(n1489), .A2(n1490), .ZN(u4_fi_ldz_2_) );
  OR2_X4 U2409 ( .A1(n2707), .A2(n2684), .ZN(n2561) );
  NAND4_X2 U2410 ( .A1(n1462), .A2(n3508), .A3(n1463), .A4(n1464), .ZN(
        u4_fi_ldz_4_) );
  NOR2_X2 U2411 ( .A1(n2687), .A2(u4_sub_406_carry[7]), .ZN(n2568) );
  NOR2_X2 U2412 ( .A1(n2562), .A2(n2463), .ZN(n1363) );
  INV_X4 U2413 ( .A(n2474), .ZN(n2624) );
  INV_X4 U2414 ( .A(n2465), .ZN(n2625) );
  INV_X4 U2415 ( .A(n2493), .ZN(n2626) );
  INV_X4 U2416 ( .A(n2490), .ZN(n2648) );
  INV_X4 U2417 ( .A(n2678), .ZN(n2677) );
  INV_X4 U2418 ( .A(u1_fractb_lt_fracta), .ZN(n2674) );
  NAND4_X2 U2419 ( .A1(n1471), .A2(n1462), .A3(n1509), .A4(n1510), .ZN(
        u4_fi_ldz_1_) );
  NOR2_X2 U2420 ( .A1(r524_A_5_), .A2(u4_sub_460_carry[5]), .ZN(n2578) );
  INV_X4 U2421 ( .A(n2668), .ZN(n2667) );
  INV_X4 U2422 ( .A(n2665), .ZN(n2664) );
  INV_X4 U2423 ( .A(n1420), .ZN(r524_A_5_) );
  INV_X4 U2424 ( .A(n2530), .ZN(n2637) );
  INV_X4 U2425 ( .A(n2530), .ZN(n2636) );
  INV_X4 U2426 ( .A(n2397), .ZN(n2640) );
  INV_X4 U2427 ( .A(n2640), .ZN(n2639) );
  INV_X4 U2428 ( .A(n2511), .ZN(n2642) );
  INV_X4 U2429 ( .A(n2511), .ZN(n2641) );
  AND2_X4 U2430 ( .A1(n1418), .A2(n2493), .ZN(n1401) );
  AND2_X4 U2431 ( .A1(n2194), .A2(n2195), .ZN(n2111) );
  AND2_X4 U2432 ( .A1(n2095), .A2(n2096), .ZN(n2631) );
  AND2_X4 U2433 ( .A1(n2095), .A2(n2096), .ZN(n2632) );
  AND2_X4 U2434 ( .A1(n2095), .A2(n2096), .ZN(n2056) );
  XNOR2_X1 U2435 ( .A(u4_sub_460_carry[5]), .B(r524_A_5_), .ZN(
        u4_fi_ldz_mi22[5]) );
  AND2_X1 U2436 ( .A1(u4_sub_460_carry[4]), .A2(u4_fi_ldz_4_), .ZN(
        u4_sub_460_carry[5]) );
  XOR2_X1 U2437 ( .A(u4_fi_ldz_4_), .B(u4_sub_460_carry[4]), .Z(
        u4_fi_ldz_mi22[4]) );
  OR2_X1 U2438 ( .A1(u4_fi_ldz_2a_3_), .A2(u4_sub_460_carry[3]), .ZN(
        u4_sub_460_carry[4]) );
  XNOR2_X1 U2439 ( .A(u4_sub_460_carry[3]), .B(u4_fi_ldz_2a_3_), .ZN(
        u4_fi_ldz_mi22[3]) );
  AND2_X1 U2440 ( .A1(u4_fi_ldz_1_), .A2(u4_fi_ldz_2_), .ZN(
        u4_sub_460_carry[3]) );
  XOR2_X1 U2441 ( .A(u4_fi_ldz_2_), .B(u4_fi_ldz_1_), .Z(u4_fi_ldz_mi22[2]) );
  XOR2_X1 U2442 ( .A(n2687), .B(u4_add_407_carry[7]), .Z(u4_div_shft2[7]) );
  AND2_X1 U2443 ( .A1(n2686), .A2(u4_add_407_carry[6]), .ZN(
        u4_add_407_carry[7]) );
  XOR2_X1 U2444 ( .A(n2686), .B(u4_add_407_carry[6]), .Z(u4_div_shft2[6]) );
  AND2_X1 U2445 ( .A1(u4_sub_478_carry[5]), .A2(n1420), .ZN(u4_N1478) );
  XOR2_X1 U2446 ( .A(n1420), .B(u4_sub_478_carry[5]), .Z(u4_N1476) );
  XOR2_X1 U2447 ( .A(n1420), .B(u4_sub_488_carry[5]), .Z(u4_fi_ldz_2a_5_) );
  AND2_X1 U2448 ( .A1(n2685), .A2(u4_add_407_carry[5]), .ZN(
        u4_add_407_carry[6]) );
  XOR2_X1 U2449 ( .A(n2685), .B(u4_add_407_carry[5]), .Z(u4_div_shft2[5]) );
  OR2_X1 U2450 ( .A1(n2722), .A2(u4_sub_478_carry[4]), .ZN(u4_sub_478_carry[5]) );
  XNOR2_X1 U2451 ( .A(u4_sub_478_carry[4]), .B(n2722), .ZN(u4_N1475) );
  OR2_X1 U2452 ( .A1(n2722), .A2(n2691), .ZN(u4_sub_488_carry[5]) );
  XNOR2_X1 U2453 ( .A(n2691), .B(n2722), .ZN(u4_fi_ldz_2a_4_) );
  AND2_X1 U2454 ( .A1(n2684), .A2(u4_add_407_carry[4]), .ZN(
        u4_add_407_carry[5]) );
  XOR2_X1 U2455 ( .A(n2684), .B(u4_add_407_carry[4]), .Z(u4_div_shft2[4]) );
  OR2_X1 U2456 ( .A1(n2691), .A2(u4_sub_478_carry[3]), .ZN(u4_sub_478_carry[4]) );
  XNOR2_X1 U2457 ( .A(u4_sub_478_carry[3]), .B(n2691), .ZN(u4_N1474) );
  AND2_X1 U2458 ( .A1(n2683), .A2(u4_add_407_carry[3]), .ZN(
        u4_add_407_carry[4]) );
  XOR2_X1 U2459 ( .A(n2683), .B(u4_add_407_carry[3]), .Z(u4_div_shft2[3]) );
  OR2_X1 U2460 ( .A1(n2723), .A2(u4_sub_478_carry[2]), .ZN(u4_sub_478_carry[3]) );
  XNOR2_X1 U2461 ( .A(u4_sub_478_carry[2]), .B(n2723), .ZN(u4_N1473) );
  OR2_X1 U2462 ( .A1(u4_fi_ldz_2a_1_), .A2(u4_fi_ldz_2a_0_), .ZN(
        u4_sub_478_carry[2]) );
  XNOR2_X1 U2463 ( .A(u4_fi_ldz_2a_0_), .B(u4_fi_ldz_2a_1_), .ZN(u4_N1472) );
  AND2_X1 U2464 ( .A1(n2682), .A2(n2681), .ZN(u4_add_407_carry[3]) );
  XOR2_X1 U2465 ( .A(n2682), .B(n2681), .Z(u4_div_shft2[2]) );
  XNOR2_X1 U2466 ( .A(n2687), .B(u4_sub_414_carry_7_), .ZN(u4_f2i_shft_7_) );
  AND2_X1 U2467 ( .A1(u4_sub_414_carry_6_), .A2(n2686), .ZN(
        u4_sub_414_carry_7_) );
  XOR2_X1 U2468 ( .A(n2686), .B(u4_sub_414_carry_6_), .Z(u4_f2i_shft_6_) );
  AND2_X1 U2469 ( .A1(u4_sub_414_carry_5_), .A2(n2685), .ZN(
        u4_sub_414_carry_6_) );
  XOR2_X1 U2470 ( .A(n2685), .B(u4_sub_414_carry_5_), .Z(u4_f2i_shft_5_) );
  AND2_X1 U2471 ( .A1(u4_sub_414_carry_4_), .A2(n2684), .ZN(
        u4_sub_414_carry_5_) );
  XOR2_X1 U2472 ( .A(n2684), .B(u4_sub_414_carry_4_), .Z(u4_f2i_shft_4_) );
  AND2_X1 U2473 ( .A1(u4_sub_414_carry_3_), .A2(n2683), .ZN(
        u4_sub_414_carry_4_) );
  XOR2_X1 U2474 ( .A(n2683), .B(u4_sub_414_carry_3_), .Z(u4_f2i_shft_3_) );
  AND2_X1 U2475 ( .A1(u4_sub_414_carry_2_), .A2(n2682), .ZN(
        u4_sub_414_carry_3_) );
  XOR2_X1 U2476 ( .A(n2682), .B(u4_sub_414_carry_2_), .Z(u4_f2i_shft_2_) );
  OR2_X1 U2477 ( .A1(n2681), .A2(n2650), .ZN(u4_sub_414_carry_2_) );
  XNOR2_X1 U2478 ( .A(n2650), .B(n2681), .ZN(u4_f2i_shft_1_) );
  AND2_X1 U2479 ( .A1(u4_add_486_carry[5]), .A2(r524_A_5_), .ZN(u4_ldz_all_6_)
         );
  XOR2_X1 U2480 ( .A(r524_A_5_), .B(u4_add_486_carry[5]), .Z(u4_ldz_all_5_) );
  AND2_X1 U2481 ( .A1(u4_N1471), .A2(div_opa_ldz_r2[0]), .ZN(
        u4_add_486_carry[1]) );
  XOR2_X1 U2482 ( .A(u4_N1471), .B(div_opa_ldz_r2[0]), .Z(u4_ldz_all_0_) );
  XNOR2_X1 U2483 ( .A(u4_sub_406_carry[7]), .B(n2687), .ZN(u4_div_scht1a[7])
         );
  OR2_X1 U2484 ( .A1(n2686), .A2(u4_sub_406_carry[6]), .ZN(u4_sub_406_carry[7]) );
  XNOR2_X1 U2485 ( .A(u4_sub_406_carry[6]), .B(n2686), .ZN(u4_div_scht1a[6])
         );
  OR2_X1 U2486 ( .A1(n2685), .A2(u4_sub_406_carry[5]), .ZN(u4_sub_406_carry[6]) );
  XNOR2_X1 U2487 ( .A(u4_sub_406_carry[5]), .B(n2685), .ZN(u4_div_scht1a[5])
         );
  OR2_X1 U2488 ( .A1(n2563), .A2(n2650), .ZN(u4_sub_406_carry[1]) );
  XNOR2_X1 U2489 ( .A(n2650), .B(n2563), .ZN(u4_div_scht1a[0]) );
  XNOR2_X1 U2490 ( .A(u2_gt_139_B_8_), .B(u2_sub_110_carry_8_), .ZN(u2_N41) );
  OR2_X1 U2491 ( .A1(u2_exp_tmp4_7_), .A2(u2_sub_110_carry_7_), .ZN(
        u2_sub_110_carry_8_) );
  XNOR2_X1 U2492 ( .A(u2_sub_110_carry_7_), .B(u2_exp_tmp4_7_), .ZN(u2_N40) );
  AND2_X1 U2493 ( .A1(u2_sub_110_carry_6_), .A2(u2_lt_129_A_6_), .ZN(
        u2_sub_110_carry_7_) );
  XOR2_X1 U2494 ( .A(u2_lt_129_A_6_), .B(u2_sub_110_carry_6_), .Z(u2_N39) );
  AND2_X1 U2495 ( .A1(u2_sub_110_carry_5_), .A2(u2_lt_129_A_5_), .ZN(
        u2_sub_110_carry_6_) );
  XOR2_X1 U2496 ( .A(u2_lt_129_A_5_), .B(u2_sub_110_carry_5_), .Z(u2_N38) );
  AND2_X1 U2497 ( .A1(u2_sub_110_carry_4_), .A2(u2_exp_tmp1_4_), .ZN(
        u2_sub_110_carry_5_) );
  XOR2_X1 U2498 ( .A(u2_exp_tmp1_4_), .B(u2_sub_110_carry_4_), .Z(u2_N37) );
  AND2_X1 U2499 ( .A1(u2_sub_110_carry_3_), .A2(u2_lt_129_A_3_), .ZN(
        u2_sub_110_carry_4_) );
  XOR2_X1 U2500 ( .A(u2_lt_129_A_3_), .B(u2_sub_110_carry_3_), .Z(u2_N36) );
  AND2_X1 U2501 ( .A1(u2_sub_110_carry_2_), .A2(u2_lt_129_A_2_), .ZN(
        u2_sub_110_carry_3_) );
  XOR2_X1 U2502 ( .A(u2_lt_129_A_2_), .B(u2_sub_110_carry_2_), .Z(u2_N35) );
  AND2_X1 U2503 ( .A1(u2_exp_tmp1_0_), .A2(u2_lt_129_A_1_), .ZN(
        u2_sub_110_carry_2_) );
  XOR2_X1 U2504 ( .A(u2_lt_129_A_1_), .B(u2_exp_tmp1_0_), .Z(u2_N34) );
  XOR2_X1 U2505 ( .A(u2_gt_139_B_8_), .B(u2_add_110_carry_8_), .Z(u2_N32) );
  AND2_X1 U2506 ( .A1(u2_add_110_carry_7_), .A2(u2_exp_tmp4_7_), .ZN(
        u2_add_110_carry_8_) );
  XOR2_X1 U2507 ( .A(u2_exp_tmp4_7_), .B(u2_add_110_carry_7_), .Z(u2_N31) );
  OR2_X1 U2508 ( .A1(u2_lt_129_A_6_), .A2(u2_add_110_carry_6_), .ZN(
        u2_add_110_carry_7_) );
  XNOR2_X1 U2509 ( .A(u2_add_110_carry_6_), .B(u2_lt_129_A_6_), .ZN(u2_N30) );
  OR2_X1 U2510 ( .A1(u2_lt_129_A_5_), .A2(u2_add_110_carry_5_), .ZN(
        u2_add_110_carry_6_) );
  XNOR2_X1 U2511 ( .A(u2_add_110_carry_5_), .B(u2_lt_129_A_5_), .ZN(u2_N29) );
  OR2_X1 U2512 ( .A1(u2_exp_tmp1_4_), .A2(u2_add_110_carry_4_), .ZN(
        u2_add_110_carry_5_) );
  XNOR2_X1 U2513 ( .A(u2_add_110_carry_4_), .B(u2_exp_tmp1_4_), .ZN(u2_N28) );
  OR2_X1 U2514 ( .A1(u2_lt_129_A_3_), .A2(u2_add_110_carry_3_), .ZN(
        u2_add_110_carry_4_) );
  XNOR2_X1 U2515 ( .A(u2_add_110_carry_3_), .B(u2_lt_129_A_3_), .ZN(u2_N27) );
  OR2_X1 U2516 ( .A1(u2_lt_129_A_2_), .A2(u2_add_110_carry_2_), .ZN(
        u2_add_110_carry_3_) );
  XNOR2_X1 U2517 ( .A(u2_add_110_carry_2_), .B(u2_lt_129_A_2_), .ZN(u2_N26) );
  OR2_X1 U2518 ( .A1(u2_lt_129_A_1_), .A2(u2_exp_tmp1_0_), .ZN(
        u2_add_110_carry_2_) );
  XNOR2_X1 U2519 ( .A(u2_exp_tmp1_0_), .B(u2_lt_129_A_1_), .ZN(u2_N25) );
  INV_X4 U2520 ( .A(u4_fi_ldz_2a_3_), .ZN(n2691) );
  INV_X4 U2521 ( .A(u4_N1471), .ZN(u4_fi_ldz_2a_0_) );
  INV_X4 U2522 ( .A(u4_fi_ldz_1_), .ZN(u4_fi_ldz_2a_1_) );
  INV_X4 U2523 ( .A(u2_exp_tmp1_0_), .ZN(u2_exp_tmp4_0_) );
  INV_X4 U2524 ( .A(u2_exp_tmp1_4_), .ZN(u2_exp_tmp4_4_) );
  OAI21_X1 U2525 ( .B1(u2_exp_tmp1_0_), .B2(u2_lt_129_A_1_), .A(n2480), .ZN(
        u2_N51) );
  NOR2_X1 U2526 ( .A1(n2480), .A2(n1586), .ZN(n2693) );
  AOI21_X1 U2527 ( .B1(n2480), .B2(n1586), .A(n2693), .ZN(n2692) );
  NAND2_X1 U2528 ( .A1(n2693), .A2(u2_lt_129_A_3_), .ZN(n2694) );
  OAI21_X1 U2529 ( .B1(n2693), .B2(u2_lt_129_A_3_), .A(n2694), .ZN(u2_N53) );
  NOR2_X1 U2530 ( .A1(n2694), .A2(u2_exp_tmp4_4_), .ZN(n2696) );
  AOI21_X1 U2531 ( .B1(n2694), .B2(u2_exp_tmp4_4_), .A(n2696), .ZN(n2695) );
  NAND2_X1 U2532 ( .A1(n2696), .A2(u2_lt_129_A_5_), .ZN(n2697) );
  OAI21_X1 U2533 ( .B1(n2696), .B2(u2_lt_129_A_5_), .A(n2697), .ZN(u2_N55) );
  XNOR2_X1 U2534 ( .A(n1583), .B(n2697), .ZN(u2_N56) );
  NOR2_X1 U2535 ( .A1(n1583), .A2(n2697), .ZN(n2698) );
  XOR2_X1 U2536 ( .A(u2_exp_tmp4_7_), .B(n2698), .Z(u2_N57) );
  INV_X4 U2537 ( .A(n2692), .ZN(u2_N52) );
  INV_X4 U2538 ( .A(n2695), .ZN(u2_N54) );
  NOR2_X1 U2539 ( .A1(n2681), .A2(n2650), .ZN(n2699) );
  OAI21_X1 U2540 ( .B1(n2473), .B2(n2486), .A(u4_sub_414_carry_2_), .ZN(
        u4_exp_in_mi1_1_) );
  NOR2_X1 U2541 ( .A1(u4_sub_414_carry_2_), .A2(n2682), .ZN(n2700) );
  OAI21_X1 U2542 ( .B1(n2699), .B2(n2559), .A(n2706), .ZN(u4_exp_in_mi1_2_) );
  NOR2_X1 U2543 ( .A1(n2706), .A2(n2683), .ZN(n2701) );
  OAI21_X1 U2544 ( .B1(n2700), .B2(n2488), .A(n2707), .ZN(u4_exp_in_mi1_3_) );
  OAI21_X1 U2545 ( .B1(n2701), .B2(n2489), .A(n2561), .ZN(u4_exp_in_mi1_4_) );
  NOR2_X1 U2546 ( .A1(n2561), .A2(n2685), .ZN(n2703) );
  AOI21_X1 U2547 ( .B1(n2561), .B2(n2685), .A(n2703), .ZN(n2702) );
  NAND2_X1 U2548 ( .A1(n2703), .A2(n2560), .ZN(n2704) );
  OAI21_X1 U2549 ( .B1(n2703), .B2(n2560), .A(n2704), .ZN(u4_exp_in_mi1_6_) );
  NOR2_X1 U2550 ( .A1(n2704), .A2(n2687), .ZN(u4_exp_in_mi1_8_) );
  AOI21_X1 U2551 ( .B1(n2704), .B2(n2687), .A(u4_exp_in_mi1_8_), .ZN(n2705) );
  INV_X4 U2552 ( .A(n2700), .ZN(n2706) );
  INV_X4 U2553 ( .A(n2701), .ZN(n2707) );
  INV_X4 U2554 ( .A(n2705), .ZN(u4_exp_in_mi1_7_) );
  INV_X4 U2555 ( .A(n2702), .ZN(u4_exp_in_mi1_5_) );
  NOR2_X1 U2556 ( .A1(u4_fi_ldz_1_), .A2(u4_N1471), .ZN(n2708) );
  OAI21_X1 U2557 ( .B1(u4_fi_ldz_2a_0_), .B2(u4_fi_ldz_2a_1_), .A(n2713), .ZN(
        u4_fi_ldz_mi1_1_) );
  OAI21_X1 U2558 ( .B1(n2708), .B2(n2723), .A(n2536), .ZN(u4_fi_ldz_mi1_2_) );
  NOR2_X1 U2559 ( .A1(n2536), .A2(u4_fi_ldz_2a_3_), .ZN(n2710) );
  AOI21_X1 U2560 ( .B1(n2536), .B2(u4_fi_ldz_2a_3_), .A(n2710), .ZN(n2709) );
  NAND2_X1 U2561 ( .A1(n2710), .A2(n2722), .ZN(n2711) );
  OAI21_X1 U2562 ( .B1(n2710), .B2(n2722), .A(n2711), .ZN(u4_fi_ldz_mi1_4_) );
  NOR2_X1 U2563 ( .A1(n2711), .A2(r524_A_5_), .ZN(u4_fi_ldz_mi1_6_) );
  AOI21_X1 U2564 ( .B1(n2711), .B2(r524_A_5_), .A(u4_fi_ldz_mi1_6_), .ZN(n2712) );
  INV_X4 U2565 ( .A(n2708), .ZN(n2713) );
  INV_X4 U2566 ( .A(n2712), .ZN(u4_fi_ldz_mi1_5_) );
  INV_X4 U2567 ( .A(n2709), .ZN(u4_fi_ldz_mi1_3_) );
  OAI21_X1 U2568 ( .B1(n1356), .B2(n2721), .A(n2535), .ZN(u4_exp_out1_mi1[1])
         );
  NOR2_X1 U2569 ( .A1(n2535), .A2(u4_sub_465_A_2_), .ZN(n2715) );
  AOI21_X1 U2570 ( .B1(n2535), .B2(u4_sub_465_A_2_), .A(n2715), .ZN(n2714) );
  NAND2_X1 U2571 ( .A1(n2715), .A2(n1376), .ZN(n2716) );
  OAI21_X1 U2572 ( .B1(n2715), .B2(n1376), .A(n2716), .ZN(u4_exp_out1_mi1[3])
         );
  NOR2_X1 U2573 ( .A1(n2716), .A2(u4_sub_465_A_4_), .ZN(n2718) );
  AOI21_X1 U2574 ( .B1(n2716), .B2(u4_sub_465_A_4_), .A(n2718), .ZN(n2717) );
  NAND2_X1 U2575 ( .A1(n2718), .A2(n1380), .ZN(n2719) );
  OAI21_X1 U2576 ( .B1(n2718), .B2(n1380), .A(n2719), .ZN(u4_exp_out1_mi1[5])
         );
  XNOR2_X1 U2577 ( .A(u4_sub_465_A_6_), .B(n2719), .ZN(u4_exp_out1_mi1[6]) );
  NOR2_X1 U2578 ( .A1(u4_sub_465_A_6_), .A2(n2719), .ZN(n2720) );
  XOR2_X1 U2579 ( .A(u4_sub_465_A_7_), .B(n2720), .Z(u4_exp_out1_mi1[7]) );
  INV_X4 U2580 ( .A(u4_exp_out1_1_), .ZN(n2721) );
  INV_X4 U2581 ( .A(n2714), .ZN(u4_exp_out1_mi1[2]) );
  INV_X4 U2582 ( .A(n2717), .ZN(u4_exp_out1_mi1[4]) );
  INV_X4 U2583 ( .A(u4_fi_ldz_4_), .ZN(n2722) );
  INV_X4 U2584 ( .A(u4_fi_ldz_2_), .ZN(n2723) );
  INV_X4 U2585 ( .A(u4_N1478), .ZN(u4_N1477) );
  INV_X1 U2586 ( .A(u4_exp_out_0_), .ZN(u4_exp_out_mi1[0]) );
  INV_X1 U2587 ( .A(u4_exp_out_1_), .ZN(n2724) );
  OAI21_X1 U2588 ( .B1(u4_exp_out_mi1[0]), .B2(n2724), .A(n2531), .ZN(
        u4_exp_out_mi1[1]) );
  NOR2_X1 U2589 ( .A1(n2531), .A2(u4_exp_out_2_), .ZN(n2727) );
  AOI21_X1 U2590 ( .B1(n2531), .B2(u4_exp_out_2_), .A(n2727), .ZN(n2725) );
  INV_X1 U2591 ( .A(n2725), .ZN(u4_exp_out_mi1[2]) );
  INV_X1 U2592 ( .A(u4_exp_out_3_), .ZN(n2726) );
  NAND2_X1 U2593 ( .A1(n2727), .A2(n2726), .ZN(n2728) );
  OAI21_X1 U2594 ( .B1(n2727), .B2(n2726), .A(n2728), .ZN(u4_exp_out_mi1[3])
         );
  NOR2_X1 U2595 ( .A1(n2728), .A2(u4_exp_out_4_), .ZN(n2731) );
  AOI21_X1 U2596 ( .B1(n2728), .B2(u4_exp_out_4_), .A(n2731), .ZN(n2729) );
  INV_X1 U2597 ( .A(n2729), .ZN(u4_exp_out_mi1[4]) );
  INV_X1 U2598 ( .A(u4_exp_out_5_), .ZN(n2730) );
  NAND2_X1 U2599 ( .A1(n2731), .A2(n2730), .ZN(n2732) );
  OAI21_X1 U2600 ( .B1(n2731), .B2(n2730), .A(n2732), .ZN(u4_exp_out_mi1[5])
         );
  XNOR2_X1 U2601 ( .A(u4_exp_out_6_), .B(n2732), .ZN(u4_exp_out_mi1[6]) );
  NOR2_X1 U2602 ( .A1(u4_exp_out_6_), .A2(n2732), .ZN(n2733) );
  XOR2_X1 U2603 ( .A(u4_N1976), .B(n2733), .Z(u4_exp_out_mi1[7]) );
  NAND2_X1 U2604 ( .A1(opb_r[26]), .A2(n2572), .ZN(n2744) );
  NAND2_X1 U2605 ( .A1(opb_r[25]), .A2(n2575), .ZN(n2743) );
  NAND2_X1 U2606 ( .A1(opb_r[30]), .A2(n2753), .ZN(n2742) );
  NAND2_X1 U2607 ( .A1(opb_r[28]), .A2(n2574), .ZN(n2747) );
  OR2_X1 U2608 ( .A1(n2577), .A2(opa_r[29]), .ZN(n2748) );
  AND2_X1 U2609 ( .A1(n2747), .A2(n2748), .ZN(n2740) );
  NAND2_X1 U2610 ( .A1(opb_r[27]), .A2(n2573), .ZN(n2746) );
  NOR2_X1 U2611 ( .A1(n2571), .A2(opb_r[23]), .ZN(n2735) );
  OAI21_X1 U2612 ( .B1(n2752), .B2(n2570), .A(opb_r[24]), .ZN(n2734) );
  OAI211_X1 U2613 ( .C1(opa_r[24]), .C2(n2735), .A(n2734), .B(n2743), .ZN(
        n2736) );
  OAI221_X1 U2614 ( .B1(opb_r[25]), .B2(n2575), .C1(opb_r[26]), .C2(n2572), 
        .A(n2736), .ZN(n2737) );
  NAND3_X1 U2615 ( .A1(n2746), .A2(n2744), .A3(n2737), .ZN(n2738) );
  OAI221_X1 U2616 ( .B1(opb_r[27]), .B2(n2573), .C1(opb_r[28]), .C2(n2574), 
        .A(n2738), .ZN(n2739) );
  AOI22_X1 U2617 ( .A1(opa_r[29]), .A2(n2577), .B1(n2740), .B2(n2739), .ZN(
        n2741) );
  OAI22_X1 U2618 ( .A1(opb_r[30]), .A2(n2753), .B1(n2754), .B2(n2741), .ZN(
        u1_expa_lt_expb) );
  NAND4_X1 U2619 ( .A1(n2744), .A2(n2743), .A3(n2742), .A4(n2655), .ZN(n2751)
         );
  AND2_X1 U2620 ( .A1(opb_r[23]), .A2(n2571), .ZN(n2745) );
  OAI22_X1 U2621 ( .A1(n2745), .A2(n2570), .B1(opb_r[24]), .B2(n2745), .ZN(
        n2749) );
  NAND4_X1 U2622 ( .A1(n2749), .A2(n2748), .A3(n2747), .A4(n2746), .ZN(n2750)
         );
  NOR2_X1 U2623 ( .A1(n2751), .A2(n2750), .ZN(u1_N34) );
  INV_X4 U2624 ( .A(n2735), .ZN(n2752) );
  INV_X4 U2625 ( .A(opa_r[30]), .ZN(n2753) );
  INV_X4 U2626 ( .A(n2742), .ZN(n2754) );
  AND2_X1 U2627 ( .A1(u4_fi_ldz_2a_4_), .A2(u4_fi_ldz_2a_3_), .ZN(n2755) );
  AND3_X1 U2628 ( .A1(u1_exp_diff_3_), .A2(u1_exp_diff_2_), .A3(u1_gt_144_B_4_), .ZN(n2756) );
  OR4_X1 U2629 ( .A1(u1_exp_diff_5_), .A2(n2756), .A3(u1_exp_diff_7_), .A4(
        u1_exp_diff_6_), .ZN(u1_exp_lt_27) );
  NOR2_X1 U2630 ( .A1(n1669), .A2(u1_gt_234_A_0_), .ZN(n2758) );
  AND2_X1 U2631 ( .A1(n1648), .A2(n2758), .ZN(n2757) );
  OAI222_X1 U2632 ( .A1(n2758), .A2(n1648), .B1(u1_gt_234_B_1_), .B2(n2757), 
        .C1(u1_gt_234_B_2_), .C2(n1632), .ZN(n2759) );
  AOI221_X1 U2633 ( .B1(n1632), .B2(u1_gt_234_B_2_), .C1(n1630), .C2(
        u1_gt_234_B_3_), .A(n2784), .ZN(n2760) );
  AOI221_X1 U2634 ( .B1(n1629), .B2(u1_gt_234_A_3_), .C1(n1627), .C2(
        u1_gt_234_A_4_), .A(n2760), .ZN(n2761) );
  AOI221_X1 U2635 ( .B1(n1628), .B2(u1_gt_234_B_4_), .C1(n1626), .C2(
        u1_gt_234_B_5_), .A(n2761), .ZN(n2762) );
  AOI221_X1 U2636 ( .B1(n1625), .B2(u1_gt_234_A_5_), .C1(n1623), .C2(
        u1_gt_234_A_6_), .A(n2762), .ZN(n2763) );
  AOI221_X1 U2637 ( .B1(n1624), .B2(u1_gt_234_B_6_), .C1(n1622), .C2(
        u1_gt_234_B_7_), .A(n2763), .ZN(n2764) );
  AOI221_X1 U2638 ( .B1(n1621), .B2(u1_gt_234_A_7_), .C1(n1619), .C2(
        u1_gt_234_A_8_), .A(n2764), .ZN(n2765) );
  AOI221_X1 U2639 ( .B1(n1620), .B2(u1_gt_234_B_8_), .C1(n1618), .C2(
        u1_gt_234_B_9_), .A(n2765), .ZN(n2766) );
  AOI221_X1 U2640 ( .B1(n1667), .B2(u1_gt_234_A_10_), .C1(n1617), .C2(
        u1_gt_234_A_9_), .A(n2766), .ZN(n2767) );
  AOI221_X1 U2641 ( .B1(n1668), .B2(u1_gt_234_B_10_), .C1(n1666), .C2(
        u1_gt_234_B_11_), .A(n2767), .ZN(n2768) );
  AOI221_X1 U2642 ( .B1(n1665), .B2(u1_gt_234_A_11_), .C1(n1663), .C2(
        u1_gt_234_A_12_), .A(n2768), .ZN(n2769) );
  AOI221_X1 U2643 ( .B1(n1664), .B2(u1_gt_234_B_12_), .C1(n1662), .C2(
        u1_gt_234_B_13_), .A(n2769), .ZN(n2770) );
  AOI221_X1 U2644 ( .B1(n1661), .B2(u1_gt_234_A_13_), .C1(n1659), .C2(
        u1_gt_234_A_14_), .A(n2770), .ZN(n2771) );
  AOI221_X1 U2645 ( .B1(n1660), .B2(u1_gt_234_B_14_), .C1(n1658), .C2(
        u1_gt_234_B_15_), .A(n2771), .ZN(n2772) );
  AOI221_X1 U2646 ( .B1(n1657), .B2(u1_gt_234_A_15_), .C1(n1655), .C2(
        u1_gt_234_A_16_), .A(n2772), .ZN(n2773) );
  AOI221_X1 U2647 ( .B1(n1656), .B2(u1_gt_234_B_16_), .C1(n1654), .C2(
        u1_gt_234_B_17_), .A(n2773), .ZN(n2774) );
  AOI221_X1 U2648 ( .B1(n1653), .B2(u1_gt_234_A_17_), .C1(n1651), .C2(
        u1_gt_234_A_18_), .A(n2774), .ZN(n2775) );
  AOI221_X1 U2649 ( .B1(n1652), .B2(u1_gt_234_B_18_), .C1(n1650), .C2(
        u1_gt_234_B_19_), .A(n2775), .ZN(n2776) );
  AOI221_X1 U2650 ( .B1(n1649), .B2(u1_gt_234_A_19_), .C1(n1645), .C2(
        u1_gt_234_A_20_), .A(n2776), .ZN(n2777) );
  AOI221_X1 U2651 ( .B1(n1646), .B2(u1_gt_234_B_20_), .C1(n1644), .C2(
        u1_gt_234_B_21_), .A(n2777), .ZN(n2778) );
  AOI221_X1 U2652 ( .B1(n1643), .B2(u1_gt_234_A_21_), .C1(n1641), .C2(
        u1_gt_234_A_22_), .A(n2778), .ZN(n2779) );
  AOI221_X1 U2653 ( .B1(n1642), .B2(u1_gt_234_B_22_), .C1(n1640), .C2(
        u1_gt_234_B_23_), .A(n2779), .ZN(n2780) );
  AOI221_X1 U2654 ( .B1(n1639), .B2(u1_gt_234_A_23_), .C1(n1637), .C2(
        u1_gt_234_A_24_), .A(n2780), .ZN(n2781) );
  AOI221_X1 U2655 ( .B1(n1638), .B2(u1_gt_234_B_24_), .C1(n1636), .C2(
        u1_gt_234_B_25_), .A(n2781), .ZN(n2782) );
  AOI221_X1 U2656 ( .B1(n1635), .B2(u1_gt_234_A_25_), .C1(n1633), .C2(
        u1_gt_234_A_26_), .A(n2782), .ZN(n2783) );
  OAI21_X1 U2657 ( .B1(u1_gt_234_A_26_), .B2(n1633), .A(n2785), .ZN(
        u1_fractb_lt_fracta) );
  INV_X4 U2658 ( .A(n2759), .ZN(n2784) );
  INV_X4 U2659 ( .A(n2783), .ZN(n2785) );
  AND3_X1 U2660 ( .A1(u4_div_shft3_1_), .A2(u4_div_shft3_0_), .A3(
        u4_div_shft3_2_), .ZN(n2786) );
  OAI21_X1 U2661 ( .B1(n2786), .B2(u4_div_shft3_3_), .A(u4_div_shft3_4_), .ZN(
        n2787) );
  OR4_X1 U2662 ( .A1(u4_div_shft3_5_), .A2(n2788), .A3(u4_div_shft3_7_), .A4(
        u4_div_shft3_6_), .ZN(u4_N1290) );
  INV_X4 U2663 ( .A(n2787), .ZN(n2788) );
  NAND4_X1 U2664 ( .A1(u4_div_exp2_4_), .A2(u4_div_exp2_3_), .A3(
        u4_div_exp2_7_), .A4(u4_div_exp2_6_), .ZN(n2790) );
  NAND4_X1 U2665 ( .A1(u4_div_exp2_1_), .A2(u4_div_exp2_0_), .A3(
        u4_div_exp2_5_), .A4(u4_div_exp2_2_), .ZN(n2789) );
  NOR2_X1 U2666 ( .A1(n2790), .A2(n2789), .ZN(u4_N1504) );
  AND3_X1 U2667 ( .A1(u4_ldz_all_2_), .A2(u4_ldz_all_1_), .A3(u4_ldz_all_0_), 
        .ZN(n2791) );
  OR2_X1 U2668 ( .A1(u4_ldz_all_3_), .A2(n2791), .ZN(n2792) );
  AOI211_X1 U2669 ( .C1(u4_ldz_all_4_), .C2(n2792), .A(u4_ldz_all_6_), .B(
        u4_ldz_all_5_), .ZN(u4_N1606) );
  OR3_X1 U2670 ( .A1(n2684), .A2(n2683), .A3(n2682), .ZN(n2793) );
  OR3_X1 U2671 ( .A1(n2681), .A2(n2650), .A3(n2793), .ZN(n2794) );
  AOI211_X1 U2672 ( .C1(n2685), .C2(n2794), .A(n2687), .B(n2686), .ZN(n2795)
         );
  INV_X4 U2673 ( .A(n2795), .ZN(u4_N1604) );
  AND3_X1 U2674 ( .A1(n2650), .A2(n2684), .A3(n2681), .ZN(n2797) );
  AND4_X1 U2675 ( .A1(n2683), .A2(n2682), .A3(n2686), .A4(n2685), .ZN(n2796)
         );
  AOI21_X1 U2676 ( .B1(n2797), .B2(n2796), .A(n2687), .ZN(u4_N1603) );
  AND3_X1 U2677 ( .A1(n2681), .A2(n2650), .A3(n2682), .ZN(n2798) );
  OAI21_X1 U2678 ( .B1(n2683), .B2(n2798), .A(n2684), .ZN(n2799) );
  NOR4_X1 U2679 ( .A1(n2687), .A2(n2686), .A3(n2685), .A4(n2800), .ZN(u4_N1600) );
  INV_X4 U2680 ( .A(n2799), .ZN(n2800) );
  AND3_X1 U2681 ( .A1(n2681), .A2(n2650), .A3(n2682), .ZN(n2801) );
  OAI21_X1 U2682 ( .B1(n2801), .B2(n2683), .A(n2684), .ZN(n2802) );
  OR4_X1 U2683 ( .A1(n2685), .A2(n2803), .A3(n2687), .A4(n2686), .ZN(u4_N1598)
         );
  INV_X4 U2684 ( .A(n2802), .ZN(n2803) );
  NAND4_X1 U2685 ( .A1(u4_div_exp1_1_), .A2(u4_div_exp1_0_), .A3(
        u4_div_exp1_5_), .A4(u4_div_exp1_2_), .ZN(n2805) );
  NAND4_X1 U2686 ( .A1(u4_div_exp1_4_), .A2(u4_div_exp1_3_), .A3(
        u4_div_exp1_7_), .A4(u4_div_exp1_6_), .ZN(n2804) );
  OAI21_X1 U2687 ( .B1(n2805), .B2(n2804), .A(n2806), .ZN(u4_N1573) );
  INV_X4 U2688 ( .A(u4_div_exp1_8_), .ZN(n2806) );
  AND3_X1 U2689 ( .A1(u4_fi_ldz_2_), .A2(u4_fi_ldz_1_), .A3(u4_N1471), .ZN(
        n2807) );
  OAI21_X1 U2690 ( .B1(n2807), .B2(u4_fi_ldz_2a_3_), .A(u4_fi_ldz_4_), .ZN(
        n2808) );
  NAND2_X1 U2691 ( .A1(n1420), .A2(n2808), .ZN(u4_N1532) );
  AND3_X1 U2692 ( .A1(u4_div_exp1_0_), .A2(u4_div_exp1_4_), .A3(u4_div_exp1_1_), .ZN(n2810) );
  AND4_X1 U2693 ( .A1(u4_div_exp1_3_), .A2(u4_div_exp1_2_), .A3(u4_div_exp1_6_), .A4(u4_div_exp1_5_), .ZN(n2809) );
  AOI21_X1 U2694 ( .B1(n2810), .B2(n2809), .A(u4_div_exp1_7_), .ZN(u4_N1523)
         );
  NOR2_X1 U2695 ( .A1(n2563), .A2(n2650), .ZN(n2811) );
  AOI21_X1 U2696 ( .B1(n2811), .B2(n2486), .A(div_opa_ldz_r2[1]), .ZN(n2812)
         );
  AOI221_X1 U2697 ( .B1(n2682), .B2(n2566), .C1(n2681), .C2(
        u4_sub_406_carry[1]), .A(n2812), .ZN(n2813) );
  AOI221_X1 U2698 ( .B1(div_opa_ldz_r2[3]), .B2(n2488), .C1(div_opa_ldz_r2[2]), 
        .C2(n2559), .A(n2813), .ZN(n2814) );
  AOI221_X1 U2699 ( .B1(n2684), .B2(n2569), .C1(n2683), .C2(n2565), .A(n2814), 
        .ZN(n2815) );
  AOI21_X1 U2700 ( .B1(div_opa_ldz_r2[4]), .B2(n2489), .A(n2815), .ZN(n2816)
         );
  NOR4_X1 U2701 ( .A1(n2687), .A2(n2686), .A3(n2685), .A4(n2816), .ZN(u4_N1503) );
  AND4_X1 U2702 ( .A1(u2_lt_129_A_3_), .A2(u2_lt_129_A_2_), .A3(u2_lt_129_A_6_), .A4(u2_lt_129_A_5_), .ZN(n2817) );
  AND4_X1 U2703 ( .A1(u2_exp_tmp1_0_), .A2(u2_exp_tmp1_4_), .A3(u2_lt_129_A_1_), .A4(n2817), .ZN(n2818) );
  OAI21_X1 U2704 ( .B1(n2818), .B2(u2_exp_tmp4_7_), .A(u2_gt_139_B_8_), .ZN(
        n2819) );
  INV_X4 U2705 ( .A(n2819), .ZN(u2_N89) );
  AND3_X1 U2706 ( .A1(u2_exp_tmp1_0_), .A2(u2_exp_tmp1_4_), .A3(u2_lt_129_A_1_), .ZN(n2821) );
  AND4_X1 U2707 ( .A1(u2_lt_129_A_3_), .A2(u2_lt_129_A_2_), .A3(u2_lt_129_A_6_), .A4(u2_lt_129_A_5_), .ZN(n2820) );
  AOI21_X1 U2708 ( .B1(n2821), .B2(n2820), .A(u2_exp_tmp4_7_), .ZN(u2_N87) );
  AND3_X1 U2709 ( .A1(u4_fi_ldz_2_), .A2(u4_fi_ldz_1_), .A3(u4_N1471), .ZN(
        n2822) );
  OR2_X1 U2710 ( .A1(u4_fi_ldz_2a_3_), .A2(n2822), .ZN(n2823) );
  AOI21_X1 U2711 ( .B1(u4_fi_ldz_4_), .B2(n2823), .A(r524_A_5_), .ZN(u4_N1599)
         );
  NOR2_X1 U2712 ( .A1(n2686), .A2(n2685), .ZN(n2825) );
  NAND4_X1 U2713 ( .A1(n2684), .A2(n2683), .A3(n2681), .A4(n2682), .ZN(n2824)
         );
  AOI21_X1 U2714 ( .B1(n2825), .B2(n2824), .A(n2558), .ZN(u4_N1284) );
  AND3_X1 U2715 ( .A1(n2684), .A2(n2686), .A3(n2681), .ZN(n2828) );
  NAND2_X1 U2716 ( .A1(r489_B_0_), .A2(n2473), .ZN(n2826) );
  AND4_X1 U2717 ( .A1(n2685), .A2(n2683), .A3(n2682), .A4(n2826), .ZN(n2827)
         );
  AOI21_X1 U2718 ( .B1(n2828), .B2(n2827), .A(n2687), .ZN(u4_N1283) );
  AOI22_X2 U2719 ( .A1(N227), .A2(n2641), .B1(N227), .B2(n2397), .ZN(n2422) );
  AOI22_X2 U2720 ( .A1(opa_r1[1]), .A2(n2642), .B1(N228), .B2(n2397), .ZN(
        n2421) );
  AOI22_X2 U2721 ( .A1(opa_r1[2]), .A2(n2642), .B1(N229), .B2(n2397), .ZN(
        n2420) );
  AOI22_X2 U2722 ( .A1(opa_r1[3]), .A2(n2642), .B1(N230), .B2(n2397), .ZN(
        n2419) );
  AOI22_X2 U2723 ( .A1(opa_r1[4]), .A2(n2642), .B1(N231), .B2(n2639), .ZN(
        n2418) );
  AOI22_X2 U2724 ( .A1(opa_r1[5]), .A2(n2642), .B1(N232), .B2(n2639), .ZN(
        n2417) );
  AOI22_X2 U2725 ( .A1(opa_r1[6]), .A2(n2642), .B1(N233), .B2(n2639), .ZN(
        n2416) );
  AOI22_X2 U2726 ( .A1(n2641), .A2(opa_r1[7]), .B1(N234), .B2(n2639), .ZN(
        n2415) );
  AOI22_X2 U2727 ( .A1(n2641), .A2(opa_r1[8]), .B1(N235), .B2(n2639), .ZN(
        n2414) );
  AOI22_X2 U2728 ( .A1(n2641), .A2(opa_r1[9]), .B1(N236), .B2(n2639), .ZN(
        n2413) );
  AOI22_X2 U2729 ( .A1(n2641), .A2(opa_r1[10]), .B1(N237), .B2(n2639), .ZN(
        n2412) );
  AOI22_X2 U2730 ( .A1(n2641), .A2(opa_r1[11]), .B1(N238), .B2(n2639), .ZN(
        n2411) );
  AOI22_X2 U2731 ( .A1(n2641), .A2(opa_r1[12]), .B1(N239), .B2(n2639), .ZN(
        n2410) );
  AOI22_X2 U2732 ( .A1(n2641), .A2(opa_r1[13]), .B1(N240), .B2(n2639), .ZN(
        n2409) );
  AOI22_X2 U2733 ( .A1(n2641), .A2(opa_r1[14]), .B1(N241), .B2(n2639), .ZN(
        n2408) );
  AOI22_X2 U2734 ( .A1(n2641), .A2(opa_r1[15]), .B1(N242), .B2(n2639), .ZN(
        n2407) );
  AOI22_X2 U2735 ( .A1(n2641), .A2(opa_r1[16]), .B1(N243), .B2(n2639), .ZN(
        n2406) );
  INV_X4 U2736 ( .A(n1975), .ZN(n3346) );
  INV_X4 U2737 ( .A(n1990), .ZN(n3347) );
  INV_X4 U2738 ( .A(n1993), .ZN(n3348) );
  INV_X4 U2739 ( .A(n1976), .ZN(n3349) );
  INV_X4 U2740 ( .A(n1979), .ZN(n3350) );
  INV_X4 U2741 ( .A(n1982), .ZN(n3351) );
  INV_X4 U2742 ( .A(n1985), .ZN(n3352) );
  INV_X4 U2743 ( .A(n1792), .ZN(u6_N48) );
  INV_X4 U2744 ( .A(n1793), .ZN(u6_N47) );
  INV_X4 U2745 ( .A(n1794), .ZN(u6_N46) );
  INV_X4 U2746 ( .A(n1795), .ZN(u6_N45) );
  INV_X4 U2747 ( .A(n1796), .ZN(u6_N44) );
  INV_X4 U2748 ( .A(n1797), .ZN(u6_N43) );
  INV_X4 U2749 ( .A(n1798), .ZN(u6_N42) );
  INV_X4 U2750 ( .A(n1799), .ZN(u6_N41) );
  INV_X4 U2751 ( .A(n1800), .ZN(u6_N40) );
  INV_X4 U2752 ( .A(n1801), .ZN(u6_N39) );
  INV_X4 U2753 ( .A(n1802), .ZN(u6_N38) );
  INV_X4 U2754 ( .A(n1803), .ZN(u6_N37) );
  INV_X4 U2755 ( .A(n1804), .ZN(u6_N36) );
  INV_X4 U2756 ( .A(n1805), .ZN(u6_N35) );
  INV_X4 U2757 ( .A(n1806), .ZN(u6_N34) );
  INV_X4 U2758 ( .A(n1807), .ZN(u6_N33) );
  INV_X4 U2759 ( .A(n1808), .ZN(u6_N32) );
  INV_X4 U2760 ( .A(n1809), .ZN(u6_N31) );
  INV_X4 U2761 ( .A(n1810), .ZN(u6_N30) );
  INV_X4 U2762 ( .A(n1811), .ZN(u6_N29) );
  INV_X4 U2763 ( .A(n1812), .ZN(u6_N28) );
  INV_X4 U2764 ( .A(n1813), .ZN(u6_N27) );
  INV_X4 U2765 ( .A(n1814), .ZN(u6_N26) );
  INV_X4 U2766 ( .A(u4_N1572), .ZN(n3353) );
  INV_X4 U2767 ( .A(n2140), .ZN(n3354) );
  INV_X4 U2768 ( .A(n2406), .ZN(n3355) );
  INV_X4 U2769 ( .A(n2407), .ZN(n3356) );
  INV_X4 U2770 ( .A(n2408), .ZN(n3357) );
  INV_X4 U2771 ( .A(n2409), .ZN(n3358) );
  INV_X4 U2772 ( .A(n2410), .ZN(n3359) );
  INV_X4 U2773 ( .A(n2411), .ZN(n3360) );
  INV_X4 U2774 ( .A(n2412), .ZN(n3361) );
  INV_X4 U2775 ( .A(n2413), .ZN(n3362) );
  INV_X4 U2776 ( .A(n2414), .ZN(n3363) );
  INV_X4 U2777 ( .A(n2415), .ZN(n3364) );
  INV_X4 U2778 ( .A(n2416), .ZN(n3365) );
  INV_X4 U2779 ( .A(n2417), .ZN(n3366) );
  INV_X4 U2780 ( .A(n2418), .ZN(n3367) );
  INV_X4 U2781 ( .A(n2419), .ZN(n3368) );
  INV_X4 U2782 ( .A(n2420), .ZN(n3369) );
  INV_X4 U2783 ( .A(n2421), .ZN(n3370) );
  INV_X4 U2784 ( .A(N325), .ZN(n3371) );
  INV_X4 U2785 ( .A(N324), .ZN(n3372) );
  INV_X4 U2786 ( .A(N323), .ZN(n3373) );
  INV_X4 U2787 ( .A(N322), .ZN(n3374) );
  INV_X4 U2788 ( .A(N321), .ZN(n3375) );
  INV_X4 U2789 ( .A(N320), .ZN(n3376) );
  INV_X4 U2790 ( .A(N319), .ZN(n3377) );
  INV_X4 U2791 ( .A(N318), .ZN(n3378) );
  INV_X4 U2792 ( .A(N317), .ZN(n3379) );
  INV_X4 U2793 ( .A(N316), .ZN(n3380) );
  INV_X4 U2794 ( .A(N315), .ZN(n3381) );
  INV_X4 U2795 ( .A(N314), .ZN(n3382) );
  INV_X4 U2796 ( .A(N313), .ZN(n3383) );
  INV_X4 U2797 ( .A(N312), .ZN(n3384) );
  INV_X4 U2798 ( .A(N311), .ZN(n3385) );
  INV_X4 U2799 ( .A(N310), .ZN(n3386) );
  INV_X4 U2800 ( .A(N309), .ZN(n3387) );
  INV_X4 U2801 ( .A(N308), .ZN(n3388) );
  INV_X4 U2802 ( .A(N307), .ZN(n3389) );
  INV_X4 U2803 ( .A(N306), .ZN(n3390) );
  INV_X4 U2804 ( .A(N305), .ZN(n3391) );
  INV_X4 U2805 ( .A(N304), .ZN(n3392) );
  INV_X4 U2806 ( .A(N303), .ZN(n3393) );
  INV_X4 U2807 ( .A(N302), .ZN(n3394) );
  INV_X4 U2808 ( .A(N301), .ZN(n3395) );
  INV_X4 U2809 ( .A(N300), .ZN(n3396) );
  INV_X4 U2810 ( .A(N299), .ZN(n3397) );
  INV_X4 U2811 ( .A(N298), .ZN(n3398) );
  INV_X4 U2812 ( .A(u2_exp_ovf_d_1_), .ZN(n3399) );
  INV_X4 U2813 ( .A(n1574), .ZN(u2_gt_139_B_8_) );
  INV_X4 U2814 ( .A(n1593), .ZN(n3400) );
  INV_X4 U2815 ( .A(n1582), .ZN(u2_exp_tmp4_7_) );
  INV_X4 U2816 ( .A(n1575), .ZN(n3401) );
  INV_X4 U2817 ( .A(n1583), .ZN(u2_lt_129_A_6_) );
  INV_X4 U2818 ( .A(n1576), .ZN(n3402) );
  INV_X4 U2819 ( .A(n1584), .ZN(u2_lt_129_A_5_) );
  INV_X4 U2820 ( .A(n1577), .ZN(n3403) );
  INV_X4 U2821 ( .A(u2_N10), .ZN(n3404) );
  INV_X4 U2822 ( .A(n1578), .ZN(n3405) );
  INV_X4 U2823 ( .A(n1585), .ZN(u2_lt_129_A_3_) );
  INV_X4 U2824 ( .A(n1579), .ZN(n3406) );
  INV_X4 U2825 ( .A(n1586), .ZN(u2_lt_129_A_2_) );
  INV_X4 U2826 ( .A(n1580), .ZN(n3407) );
  INV_X4 U2827 ( .A(n1587), .ZN(u2_lt_129_A_1_) );
  INV_X4 U2828 ( .A(n1581), .ZN(n3408) );
  INV_X4 U2829 ( .A(u2_N6), .ZN(n3409) );
  INV_X4 U2830 ( .A(u2_N19), .ZN(n3410) );
  INV_X4 U2831 ( .A(u2_N15), .ZN(n3411) );
  INV_X4 U2832 ( .A(n1817), .ZN(n3412) );
  INV_X4 U2833 ( .A(n1765), .ZN(n3413) );
  INV_X4 U2834 ( .A(n1766), .ZN(n3414) );
  INV_X4 U2835 ( .A(n1767), .ZN(n3415) );
  INV_X4 U2836 ( .A(n1768), .ZN(n3416) );
  INV_X4 U2837 ( .A(n1769), .ZN(n3417) );
  INV_X4 U2838 ( .A(n1770), .ZN(n3418) );
  INV_X4 U2839 ( .A(n1771), .ZN(n3419) );
  INV_X4 U2840 ( .A(n1773), .ZN(n3420) );
  INV_X4 U2841 ( .A(n1774), .ZN(n3421) );
  INV_X4 U2842 ( .A(n1775), .ZN(n3422) );
  INV_X4 U2843 ( .A(n1776), .ZN(n3423) );
  INV_X4 U2844 ( .A(n1777), .ZN(n3424) );
  INV_X4 U2845 ( .A(n1778), .ZN(n3425) );
  INV_X4 U2846 ( .A(n1779), .ZN(n3426) );
  INV_X4 U2847 ( .A(n1780), .ZN(n3427) );
  INV_X4 U2848 ( .A(n1781), .ZN(n3428) );
  INV_X4 U2849 ( .A(n1782), .ZN(n3429) );
  INV_X4 U2850 ( .A(n1757), .ZN(n3430) );
  INV_X4 U2851 ( .A(n1758), .ZN(n3431) );
  INV_X4 U2852 ( .A(n1759), .ZN(n3432) );
  INV_X4 U2853 ( .A(n1760), .ZN(n3433) );
  INV_X4 U2854 ( .A(n1761), .ZN(n3434) );
  INV_X4 U2855 ( .A(n1762), .ZN(n3435) );
  INV_X4 U2856 ( .A(n1763), .ZN(n3436) );
  INV_X4 U2857 ( .A(n1764), .ZN(n3437) );
  INV_X4 U2858 ( .A(n1772), .ZN(n3438) );
  INV_X4 U2859 ( .A(n1783), .ZN(n3439) );
  INV_X4 U2860 ( .A(u4_exp_f2i_1[49]), .ZN(n3440) );
  INV_X4 U2861 ( .A(n2008), .ZN(n3441) );
  INV_X4 U2862 ( .A(n1393), .ZN(n3442) );
  INV_X4 U2863 ( .A(u4_exp_next_mi_8_), .ZN(n3443) );
  INV_X4 U2864 ( .A(n1384), .ZN(u4_sub_465_A_7_) );
  INV_X4 U2865 ( .A(n1382), .ZN(u4_sub_465_A_6_) );
  INV_X4 U2866 ( .A(n1378), .ZN(u4_sub_465_A_4_) );
  INV_X4 U2867 ( .A(n1374), .ZN(u4_sub_465_A_2_) );
  INV_X4 U2868 ( .A(u4_exp_next_mi_1_), .ZN(n3444) );
  INV_X4 U2869 ( .A(n1356), .ZN(u4_sub_465_A_0_) );
  INV_X4 U2870 ( .A(n1721), .ZN(n3445) );
  INV_X4 U2871 ( .A(n1617), .ZN(u1_gt_234_B_9_) );
  INV_X4 U2872 ( .A(n1619), .ZN(u1_gt_234_B_8_) );
  INV_X4 U2873 ( .A(n1621), .ZN(u1_gt_234_B_7_) );
  INV_X4 U2874 ( .A(n1623), .ZN(u1_gt_234_B_6_) );
  INV_X4 U2875 ( .A(n1625), .ZN(u1_gt_234_B_5_) );
  INV_X4 U2876 ( .A(n1627), .ZN(u1_gt_234_B_4_) );
  INV_X4 U2877 ( .A(n1629), .ZN(u1_gt_234_B_3_) );
  INV_X4 U2878 ( .A(n1635), .ZN(u1_gt_234_B_25_) );
  INV_X4 U2879 ( .A(n1637), .ZN(u1_gt_234_B_24_) );
  INV_X4 U2880 ( .A(n1639), .ZN(u1_gt_234_B_23_) );
  INV_X4 U2881 ( .A(n1641), .ZN(u1_gt_234_B_22_) );
  INV_X4 U2882 ( .A(n1643), .ZN(u1_gt_234_B_21_) );
  INV_X4 U2883 ( .A(n1645), .ZN(u1_gt_234_B_20_) );
  INV_X4 U2884 ( .A(n1649), .ZN(u1_gt_234_B_19_) );
  INV_X4 U2885 ( .A(n1651), .ZN(u1_gt_234_B_18_) );
  INV_X4 U2886 ( .A(n1653), .ZN(u1_gt_234_B_17_) );
  INV_X4 U2887 ( .A(n1655), .ZN(u1_gt_234_B_16_) );
  INV_X4 U2888 ( .A(n1657), .ZN(u1_gt_234_B_15_) );
  INV_X4 U2889 ( .A(n1659), .ZN(u1_gt_234_B_14_) );
  INV_X4 U2890 ( .A(n1661), .ZN(u1_gt_234_B_13_) );
  INV_X4 U2891 ( .A(n1663), .ZN(u1_gt_234_B_12_) );
  INV_X4 U2892 ( .A(n1665), .ZN(u1_gt_234_B_11_) );
  INV_X4 U2893 ( .A(n1667), .ZN(u1_gt_234_B_10_) );
  INV_X4 U2894 ( .A(n1618), .ZN(u1_gt_234_A_9_) );
  INV_X4 U2895 ( .A(n1620), .ZN(u1_gt_234_A_8_) );
  INV_X4 U2896 ( .A(n1622), .ZN(u1_gt_234_A_7_) );
  INV_X4 U2897 ( .A(n1624), .ZN(u1_gt_234_A_6_) );
  INV_X4 U2898 ( .A(n1626), .ZN(u1_gt_234_A_5_) );
  INV_X4 U2899 ( .A(n1628), .ZN(u1_gt_234_A_4_) );
  INV_X4 U2900 ( .A(n1630), .ZN(u1_gt_234_A_3_) );
  INV_X4 U2901 ( .A(n1634), .ZN(u1_gt_234_A_26_) );
  INV_X4 U2902 ( .A(n1636), .ZN(u1_gt_234_A_25_) );
  INV_X4 U2903 ( .A(n1638), .ZN(u1_gt_234_A_24_) );
  INV_X4 U2904 ( .A(n1640), .ZN(u1_gt_234_A_23_) );
  INV_X4 U2905 ( .A(n1642), .ZN(u1_gt_234_A_22_) );
  INV_X4 U2906 ( .A(n1644), .ZN(u1_gt_234_A_21_) );
  INV_X4 U2907 ( .A(n1646), .ZN(u1_gt_234_A_20_) );
  INV_X4 U2908 ( .A(n1650), .ZN(u1_gt_234_A_19_) );
  INV_X4 U2909 ( .A(n1652), .ZN(u1_gt_234_A_18_) );
  INV_X4 U2910 ( .A(n1654), .ZN(u1_gt_234_A_17_) );
  INV_X4 U2911 ( .A(n1656), .ZN(u1_gt_234_A_16_) );
  INV_X4 U2912 ( .A(n1658), .ZN(u1_gt_234_A_15_) );
  INV_X4 U2913 ( .A(n1660), .ZN(u1_gt_234_A_14_) );
  INV_X4 U2914 ( .A(n1662), .ZN(u1_gt_234_A_13_) );
  INV_X4 U2915 ( .A(n1664), .ZN(u1_gt_234_A_12_) );
  INV_X4 U2916 ( .A(n1666), .ZN(u1_gt_234_A_11_) );
  INV_X4 U2917 ( .A(n1668), .ZN(u1_gt_234_A_10_) );
  INV_X4 U2918 ( .A(n1670), .ZN(u1_gt_234_A_0_) );
  INV_X4 U2919 ( .A(u1_adj_op_out_sft_0_), .ZN(n3446) );
  INV_X4 U2920 ( .A(n1647), .ZN(u1_gt_234_B_1_) );
  INV_X4 U2921 ( .A(n1631), .ZN(u1_gt_234_B_2_) );
  INV_X4 U2922 ( .A(n1681), .ZN(n3447) );
  INV_X4 U2923 ( .A(n1683), .ZN(n3448) );
  INV_X4 U2924 ( .A(u1_exp_lt_27), .ZN(n3449) );
  INV_X4 U2925 ( .A(n1687), .ZN(n3450) );
  INV_X4 U2926 ( .A(n1675), .ZN(n3451) );
  INV_X4 U2927 ( .A(n1685), .ZN(n3452) );
  INV_X4 U2928 ( .A(n1707), .ZN(u1_gt_144_B_4_) );
  INV_X4 U2929 ( .A(n1688), .ZN(n3453) );
  INV_X4 U2930 ( .A(n1689), .ZN(n3454) );
  INV_X4 U2931 ( .A(n1709), .ZN(n3455) );
  INV_X4 U2932 ( .A(n1695), .ZN(n3456) );
  INV_X4 U2933 ( .A(n1696), .ZN(n3457) );
  INV_X4 U2934 ( .A(n1697), .ZN(n3458) );
  INV_X4 U2935 ( .A(n1698), .ZN(n3459) );
  INV_X4 U2936 ( .A(n1710), .ZN(n3460) );
  INV_X4 U2937 ( .A(n1711), .ZN(n3461) );
  INV_X4 U2938 ( .A(n1712), .ZN(n3462) );
  INV_X4 U2939 ( .A(n1713), .ZN(n3463) );
  INV_X4 U2940 ( .A(n1714), .ZN(n3464) );
  INV_X4 U2941 ( .A(n1715), .ZN(n3465) );
  INV_X4 U2942 ( .A(n1716), .ZN(n3466) );
  INV_X4 U2943 ( .A(n1717), .ZN(n3467) );
  INV_X4 U2944 ( .A(n1718), .ZN(n3468) );
  INV_X4 U2945 ( .A(n1719), .ZN(n3469) );
  INV_X4 U2946 ( .A(n1699), .ZN(n3470) );
  INV_X4 U2947 ( .A(n1700), .ZN(n3471) );
  INV_X4 U2948 ( .A(n1701), .ZN(n3472) );
  INV_X4 U2949 ( .A(n1702), .ZN(n3473) );
  INV_X4 U2950 ( .A(n1703), .ZN(n3474) );
  INV_X4 U2951 ( .A(n1704), .ZN(n3475) );
  INV_X4 U2952 ( .A(n1705), .ZN(n3476) );
  INV_X4 U2953 ( .A(n1706), .ZN(n3477) );
  INV_X4 U2954 ( .A(n1737), .ZN(n3478) );
  INV_X4 U2955 ( .A(n1573), .ZN(n3479) );
  INV_X4 U2956 ( .A(n1571), .ZN(n3480) );
  INV_X4 U2957 ( .A(n1746), .ZN(n3481) );
  INV_X4 U2958 ( .A(n1818), .ZN(n3482) );
  INV_X4 U2959 ( .A(n2445), .ZN(n3483) );
  INV_X4 U2960 ( .A(n1736), .ZN(n3484) );
  INV_X4 U2961 ( .A(u6_N23), .ZN(n3485) );
  INV_X4 U2962 ( .A(n1572), .ZN(n3486) );
  INV_X4 U2963 ( .A(u4_N1283), .ZN(n3487) );
  INV_X4 U2964 ( .A(n1388), .ZN(n3488) );
  INV_X4 U2965 ( .A(n1355), .ZN(n3489) );
  INV_X4 U2966 ( .A(n2104), .ZN(r489_B_0_) );
  INV_X4 U2967 ( .A(n1952), .ZN(n3491) );
  INV_X4 U2968 ( .A(n2193), .ZN(n3492) );
  INV_X4 U2969 ( .A(n1949), .ZN(n3493) );
  INV_X4 U2970 ( .A(n2422), .ZN(n3495) );
  INV_X4 U2971 ( .A(n2394), .ZN(n3496) );
  INV_X4 U2972 ( .A(n2405), .ZN(n3497) );
  INV_X4 U2973 ( .A(n1448), .ZN(n3498) );
  INV_X4 U2974 ( .A(n2100), .ZN(n3499) );
  INV_X4 U2975 ( .A(u4_N1532), .ZN(n3500) );
  INV_X4 U2976 ( .A(n1500), .ZN(n3501) );
  INV_X4 U2977 ( .A(n1492), .ZN(n3502) );
  INV_X4 U2978 ( .A(n1469), .ZN(n3503) );
  INV_X4 U2979 ( .A(n1386), .ZN(n3504) );
  INV_X4 U2980 ( .A(n1476), .ZN(n3505) );
  INV_X4 U2981 ( .A(n1495), .ZN(n3506) );
  INV_X4 U2982 ( .A(n1529), .ZN(n3507) );
  INV_X4 U2983 ( .A(n1527), .ZN(n3508) );
  INV_X4 U2984 ( .A(n1485), .ZN(n3509) );
  INV_X4 U2985 ( .A(n1470), .ZN(n3510) );
  INV_X4 U2986 ( .A(n1496), .ZN(n3511) );
  INV_X4 U2987 ( .A(n1486), .ZN(n3512) );
  INV_X4 U2988 ( .A(n1481), .ZN(n3513) );
  INV_X4 U2989 ( .A(n1468), .ZN(n3514) );
  INV_X4 U2990 ( .A(n1482), .ZN(n3515) );
  INV_X4 U2991 ( .A(n1833), .ZN(n3516) );
  INV_X4 U2992 ( .A(n2194), .ZN(n3517) );
  INV_X4 U2993 ( .A(n2232), .ZN(n3518) );
  INV_X4 U2994 ( .A(n2022), .ZN(n3519) );
  INV_X4 U2995 ( .A(n1395), .ZN(n3520) );
  INV_X4 U2996 ( .A(n2224), .ZN(n3521) );
  INV_X4 U2997 ( .A(n1558), .ZN(n3522) );
  INV_X4 U2998 ( .A(n1786), .ZN(n3523) );
  INV_X4 U2999 ( .A(n1497), .ZN(n3524) );
  INV_X4 U3000 ( .A(n1541), .ZN(n3525) );
  INV_X4 U3001 ( .A(n1477), .ZN(n3526) );
  INV_X4 U3002 ( .A(n1555), .ZN(n3527) );
  INV_X4 U3003 ( .A(n2229), .ZN(n3528) );
  INV_X4 U3004 ( .A(n2222), .ZN(n3529) );
  INV_X4 U3005 ( .A(n1507), .ZN(n3530) );
  INV_X4 U3006 ( .A(n1546), .ZN(n3531) );
  INV_X4 U3007 ( .A(n1789), .ZN(n3532) );
  INV_X4 U3008 ( .A(n2225), .ZN(n3533) );
  INV_X4 U3009 ( .A(n1532), .ZN(n3534) );
  INV_X4 U3010 ( .A(fract_denorm[21]), .ZN(n3535) );
  INV_X4 U3011 ( .A(fract_denorm[22]), .ZN(n3536) );
  INV_X4 U3012 ( .A(fract_denorm[25]), .ZN(n3537) );
  INV_X4 U3013 ( .A(fract_denorm[26]), .ZN(n3538) );
  INV_X4 U3014 ( .A(n1488), .ZN(n3539) );
  INV_X4 U3015 ( .A(fract_denorm[29]), .ZN(n3540) );
  INV_X4 U3016 ( .A(n1551), .ZN(n3541) );
  INV_X4 U3017 ( .A(fract_denorm[30]), .ZN(n3542) );
  INV_X4 U3018 ( .A(fract_denorm[23]), .ZN(n3543) );
  INV_X4 U3019 ( .A(fract_denorm[32]), .ZN(n3544) );
  INV_X4 U3020 ( .A(n1542), .ZN(n3545) );
  INV_X4 U3021 ( .A(fract_denorm[34]), .ZN(n3546) );
  INV_X4 U3022 ( .A(n1552), .ZN(n3547) );
  INV_X4 U3023 ( .A(fract_denorm[37]), .ZN(n3548) );
  INV_X4 U3024 ( .A(n1554), .ZN(n3549) );
  INV_X4 U3025 ( .A(fract_denorm[36]), .ZN(n3550) );
  INV_X4 U3026 ( .A(fract_denorm[40]), .ZN(n3551) );
  INV_X4 U3027 ( .A(fract_denorm[45]), .ZN(n3552) );
  INV_X4 U3028 ( .A(n1553), .ZN(n3553) );
  INV_X4 U3029 ( .A(fract_denorm[46]), .ZN(n3554) );
  INV_X4 U3030 ( .A(fract_denorm[43]), .ZN(n3555) );
  INV_X4 U3031 ( .A(fract_denorm[42]), .ZN(n3556) );
  INV_X4 U3032 ( .A(n1787), .ZN(n3557) );
  INV_X4 U3033 ( .A(n2317), .ZN(n3558) );
  INV_X4 U3034 ( .A(n1788), .ZN(n3559) );
  INV_X4 U3035 ( .A(n1514), .ZN(n3560) );
  INV_X4 U3036 ( .A(n1790), .ZN(n3561) );
  INV_X4 U3037 ( .A(n1785), .ZN(n3562) );
  INV_X4 U3038 ( .A(n2227), .ZN(n3563) );
  INV_X4 U3039 ( .A(n1791), .ZN(n3564) );
  INV_X4 U3040 ( .A(n1835), .ZN(n3566) );
  INV_X4 U3041 ( .A(n1938), .ZN(n3567) );
  INV_X4 U3042 ( .A(n1730), .ZN(n3568) );
  INV_X4 U3043 ( .A(n1731), .ZN(n3569) );
  INV_X4 U3044 ( .A(n1732), .ZN(n3570) );
  INV_X4 U3045 ( .A(n1733), .ZN(n3571) );
  INV_X4 U3046 ( .A(n2028), .ZN(n3572) );
  INV_X4 U3047 ( .A(n1832), .ZN(n3573) );
  INV_X4 U3048 ( .A(n1936), .ZN(n3574) );
  INV_X4 U3049 ( .A(n1829), .ZN(n3575) );
  INV_X4 U3050 ( .A(n2030), .ZN(n3576) );
  INV_X4 U3051 ( .A(n1844), .ZN(n3577) );
  INV_X4 U3052 ( .A(n1933), .ZN(n3578) );
  INV_X4 U3053 ( .A(n2129), .ZN(n3579) );
  INV_X4 U3054 ( .A(n1417), .ZN(n3580) );
  INV_X4 U3055 ( .A(u4_exp_in_pl1_5_), .ZN(n3581) );
  INV_X4 U3056 ( .A(u4_exp_in_pl1_1_), .ZN(n3582) );
  INV_X4 U3057 ( .A(n1444), .ZN(n3583) );
  INV_X4 U3058 ( .A(n2128), .ZN(n3584) );
  INV_X4 u4_sub_470_U11 ( .A(u4_fi_ldz_2a_0_), .ZN(u4_sub_470_n8) );
  INV_X4 u4_sub_470_U10 ( .A(u4_fi_ldz_mi1_1_), .ZN(u4_sub_470_n7) );
  INV_X4 u4_sub_470_U9 ( .A(u4_fi_ldz_mi1_5_), .ZN(u4_sub_470_n6) );
  INV_X4 u4_sub_470_U8 ( .A(u4_fi_ldz_mi1_6_), .ZN(u4_sub_470_n5) );
  INV_X4 u4_sub_470_U7 ( .A(u4_fi_ldz_mi1_4_), .ZN(u4_sub_470_n4) );
  INV_X4 u4_sub_470_U6 ( .A(u4_fi_ldz_mi1_3_), .ZN(u4_sub_470_n3) );
  INV_X4 u4_sub_470_U5 ( .A(u4_fi_ldz_mi1_2_), .ZN(u4_sub_470_n2) );
  INV_X4 u4_sub_470_U4 ( .A(n2650), .ZN(u4_sub_470_n1) );
  XNOR2_X2 u4_sub_470_U3 ( .A(u4_sub_470_n8), .B(n2650), .ZN(
        u4_exp_fix_divb[0]) );
  NAND2_X2 u4_sub_470_U2 ( .A1(u4_fi_ldz_2a_0_), .A2(u4_sub_470_n1), .ZN(
        u4_sub_470_carry[1]) );
  XNOR2_X2 u4_sub_470_U1 ( .A(n2687), .B(u4_sub_470_carry[7]), .ZN(
        u4_exp_fix_divb[7]) );
  FA_X1 u4_sub_470_U2_1 ( .A(n2681), .B(u4_sub_470_n7), .CI(
        u4_sub_470_carry[1]), .CO(u4_sub_470_carry[2]), .S(u4_exp_fix_divb[1])
         );
  FA_X1 u4_sub_470_U2_2 ( .A(n2682), .B(u4_sub_470_n2), .CI(
        u4_sub_470_carry[2]), .CO(u4_sub_470_carry[3]), .S(u4_exp_fix_divb[2])
         );
  FA_X1 u4_sub_470_U2_3 ( .A(n2683), .B(u4_sub_470_n3), .CI(
        u4_sub_470_carry[3]), .CO(u4_sub_470_carry[4]), .S(u4_exp_fix_divb[3])
         );
  FA_X1 u4_sub_470_U2_4 ( .A(n2684), .B(u4_sub_470_n4), .CI(
        u4_sub_470_carry[4]), .CO(u4_sub_470_carry[5]), .S(u4_exp_fix_divb[4])
         );
  FA_X1 u4_sub_470_U2_5 ( .A(n2685), .B(u4_sub_470_n6), .CI(
        u4_sub_470_carry[5]), .CO(u4_sub_470_carry[6]), .S(u4_exp_fix_divb[5])
         );
  FA_X1 u4_sub_470_U2_6 ( .A(n2686), .B(u4_sub_470_n5), .CI(
        u4_sub_470_carry[6]), .CO(u4_sub_470_carry[7]), .S(u4_exp_fix_divb[6])
         );
  INV_X4 u4_sub_469_U11 ( .A(u4_N1471), .ZN(u4_sub_469_n8) );
  INV_X4 u4_sub_469_U10 ( .A(u4_fi_ldz_2a_1_), .ZN(u4_sub_469_n7) );
  INV_X4 u4_sub_469_U9 ( .A(u4_fi_ldz_mi22[2]), .ZN(u4_sub_469_n6) );
  INV_X4 u4_sub_469_U8 ( .A(u4_fi_ldz_mi22[3]), .ZN(u4_sub_469_n5) );
  INV_X4 u4_sub_469_U7 ( .A(u4_fi_ldz_mi22[4]), .ZN(u4_sub_469_n4) );
  INV_X4 u4_sub_469_U6 ( .A(u4_fi_ldz_mi22[5]), .ZN(u4_sub_469_n3) );
  INV_X4 u4_sub_469_U5 ( .A(n2578), .ZN(u4_sub_469_n2) );
  INV_X4 u4_sub_469_U4 ( .A(n2650), .ZN(u4_sub_469_n1) );
  XNOR2_X2 u4_sub_469_U3 ( .A(u4_sub_469_n8), .B(n2650), .ZN(
        u4_exp_fix_diva[0]) );
  NAND2_X2 u4_sub_469_U2 ( .A1(u4_N1471), .A2(u4_sub_469_n1), .ZN(
        u4_sub_469_carry[1]) );
  XNOR2_X2 u4_sub_469_U1 ( .A(n2687), .B(u4_sub_469_carry[7]), .ZN(
        u4_exp_fix_diva[7]) );
  FA_X1 u4_sub_469_U2_1 ( .A(n2681), .B(u4_sub_469_n7), .CI(
        u4_sub_469_carry[1]), .CO(u4_sub_469_carry[2]), .S(u4_exp_fix_diva[1])
         );
  FA_X1 u4_sub_469_U2_2 ( .A(n2682), .B(u4_sub_469_n6), .CI(
        u4_sub_469_carry[2]), .CO(u4_sub_469_carry[3]), .S(u4_exp_fix_diva[2])
         );
  FA_X1 u4_sub_469_U2_3 ( .A(n2683), .B(u4_sub_469_n5), .CI(
        u4_sub_469_carry[3]), .CO(u4_sub_469_carry[4]), .S(u4_exp_fix_diva[3])
         );
  FA_X1 u4_sub_469_U2_4 ( .A(n2684), .B(u4_sub_469_n4), .CI(
        u4_sub_469_carry[4]), .CO(u4_sub_469_carry[5]), .S(u4_exp_fix_diva[4])
         );
  FA_X1 u4_sub_469_U2_5 ( .A(n2685), .B(u4_sub_469_n3), .CI(
        u4_sub_469_carry[5]), .CO(u4_sub_469_carry[6]), .S(u4_exp_fix_diva[5])
         );
  FA_X1 u4_sub_469_U2_6 ( .A(n2686), .B(u4_sub_469_n2), .CI(
        u4_sub_469_carry[6]), .CO(u4_sub_469_carry[7]), .S(u4_exp_fix_diva[6])
         );
  INV_X1 u4_add_461_U2 ( .A(u4_exp_out_0_), .ZN(u4_exp_out_pl1_0_) );
  XOR2_X1 u4_add_461_U1 ( .A(u4_add_461_carry[7]), .B(u4_N1976), .Z(
        u4_exp_out_pl1_7_) );
  HA_X1 u4_add_461_U1_1_1 ( .A(u4_exp_out_1_), .B(u4_exp_out_0_), .CO(
        u4_add_461_carry[2]), .S(u4_exp_out_pl1_1_) );
  HA_X1 u4_add_461_U1_1_2 ( .A(u4_exp_out_2_), .B(u4_add_461_carry[2]), .CO(
        u4_add_461_carry[3]), .S(u4_exp_out_pl1_2_) );
  HA_X1 u4_add_461_U1_1_3 ( .A(u4_exp_out_3_), .B(u4_add_461_carry[3]), .CO(
        u4_add_461_carry[4]), .S(u4_exp_out_pl1_3_) );
  HA_X1 u4_add_461_U1_1_4 ( .A(u4_exp_out_4_), .B(u4_add_461_carry[4]), .CO(
        u4_add_461_carry[5]), .S(u4_exp_out_pl1_4_) );
  HA_X1 u4_add_461_U1_1_5 ( .A(u4_exp_out_5_), .B(u4_add_461_carry[5]), .CO(
        u4_add_461_carry[6]), .S(u4_exp_out_pl1_5_) );
  HA_X1 u4_add_461_U1_1_6 ( .A(u4_exp_out_6_), .B(u4_add_461_carry[6]), .CO(
        u4_add_461_carry[7]), .S(u4_exp_out_pl1_6_) );
  AND2_X1 u4_sll_451_U118 ( .A1(n3564), .A2(u4_sll_451_n33), .ZN(
        u4_sll_451_ML_int_1__0_) );
  AND2_X1 u4_sll_451_U117 ( .A1(u4_sll_451_ML_int_1__0_), .A2(u4_sll_451_n31), 
        .ZN(u4_sll_451_ML_int_2__0_) );
  AND2_X1 u4_sll_451_U116 ( .A1(u4_sll_451_ML_int_1__1_), .A2(u4_sll_451_n31), 
        .ZN(u4_sll_451_ML_int_2__1_) );
  AND2_X1 u4_sll_451_U115 ( .A1(u4_sll_451_ML_int_2__0_), .A2(u4_sll_451_n23), 
        .ZN(u4_sll_451_ML_int_3__0_) );
  AND2_X1 u4_sll_451_U114 ( .A1(u4_sll_451_ML_int_2__1_), .A2(u4_sll_451_n22), 
        .ZN(u4_sll_451_ML_int_3__1_) );
  AND2_X1 u4_sll_451_U113 ( .A1(u4_sll_451_ML_int_2__2_), .A2(u4_sll_451_n23), 
        .ZN(u4_sll_451_ML_int_3__2_) );
  AND2_X1 u4_sll_451_U112 ( .A1(u4_sll_451_ML_int_2__3_), .A2(u4_sll_451_n23), 
        .ZN(u4_sll_451_ML_int_3__3_) );
  AND2_X1 u4_sll_451_U111 ( .A1(u4_sll_451_ML_int_3__0_), .A2(u4_sll_451_n19), 
        .ZN(u4_sll_451_ML_int_4__0_) );
  AND2_X1 u4_sll_451_U110 ( .A1(u4_sll_451_ML_int_3__1_), .A2(u4_sll_451_n19), 
        .ZN(u4_sll_451_ML_int_4__1_) );
  AND2_X1 u4_sll_451_U109 ( .A1(u4_sll_451_ML_int_3__2_), .A2(u4_sll_451_n19), 
        .ZN(u4_sll_451_ML_int_4__2_) );
  AND2_X1 u4_sll_451_U108 ( .A1(u4_sll_451_ML_int_3__3_), .A2(u4_sll_451_n14), 
        .ZN(u4_sll_451_ML_int_4__3_) );
  AND2_X1 u4_sll_451_U107 ( .A1(u4_sll_451_ML_int_3__4_), .A2(u4_sll_451_n14), 
        .ZN(u4_sll_451_ML_int_4__4_) );
  AND2_X1 u4_sll_451_U106 ( .A1(u4_sll_451_ML_int_3__5_), .A2(u4_sll_451_n14), 
        .ZN(u4_sll_451_ML_int_4__5_) );
  AND2_X1 u4_sll_451_U105 ( .A1(u4_sll_451_ML_int_3__6_), .A2(u4_sll_451_n14), 
        .ZN(u4_sll_451_ML_int_4__6_) );
  AND2_X1 u4_sll_451_U104 ( .A1(u4_sll_451_ML_int_3__7_), .A2(u4_sll_451_n14), 
        .ZN(u4_sll_451_ML_int_4__7_) );
  NAND2_X1 u4_sll_451_U103 ( .A1(u4_sll_451_ML_int_4__0_), .A2(u4_sll_451_n6), 
        .ZN(u4_sll_451_n53) );
  INV_X1 u4_sll_451_U102 ( .A(u4_sll_451_n53), .ZN(u4_sll_451_ML_int_5__0_) );
  NAND2_X1 u4_sll_451_U101 ( .A1(u4_sll_451_ML_int_4__10_), .A2(u4_sll_451_n6), 
        .ZN(u4_sll_451_n52) );
  INV_X1 u4_sll_451_U100 ( .A(u4_sll_451_n52), .ZN(u4_sll_451_ML_int_5__10_)
         );
  NAND2_X1 u4_sll_451_U99 ( .A1(u4_sll_451_ML_int_4__11_), .A2(u4_sll_451_n7), 
        .ZN(u4_sll_451_n51) );
  INV_X1 u4_sll_451_U98 ( .A(u4_sll_451_n51), .ZN(u4_sll_451_ML_int_5__11_) );
  NAND2_X1 u4_sll_451_U97 ( .A1(u4_sll_451_ML_int_4__12_), .A2(u4_sll_451_n7), 
        .ZN(u4_sll_451_n50) );
  INV_X1 u4_sll_451_U96 ( .A(u4_sll_451_n50), .ZN(u4_sll_451_ML_int_5__12_) );
  NAND2_X1 u4_sll_451_U95 ( .A1(u4_sll_451_ML_int_4__13_), .A2(u4_sll_451_n7), 
        .ZN(u4_sll_451_n49) );
  INV_X1 u4_sll_451_U94 ( .A(u4_sll_451_n49), .ZN(u4_sll_451_ML_int_5__13_) );
  NAND2_X1 u4_sll_451_U93 ( .A1(u4_sll_451_ML_int_4__14_), .A2(u4_sll_451_n7), 
        .ZN(u4_sll_451_n48) );
  INV_X1 u4_sll_451_U92 ( .A(u4_sll_451_n48), .ZN(u4_sll_451_ML_int_5__14_) );
  NAND2_X1 u4_sll_451_U91 ( .A1(u4_sll_451_ML_int_4__15_), .A2(u4_sll_451_n7), 
        .ZN(u4_sll_451_n47) );
  INV_X1 u4_sll_451_U90 ( .A(u4_sll_451_n47), .ZN(u4_sll_451_ML_int_5__15_) );
  NAND2_X1 u4_sll_451_U89 ( .A1(u4_sll_451_ML_int_4__1_), .A2(u4_sll_451_n7), 
        .ZN(u4_sll_451_n46) );
  INV_X1 u4_sll_451_U88 ( .A(u4_sll_451_n46), .ZN(u4_sll_451_ML_int_5__1_) );
  NAND2_X1 u4_sll_451_U87 ( .A1(u4_sll_451_ML_int_4__2_), .A2(u4_sll_451_n7), 
        .ZN(u4_sll_451_n45) );
  INV_X1 u4_sll_451_U86 ( .A(u4_sll_451_n45), .ZN(u4_sll_451_ML_int_5__2_) );
  NAND2_X1 u4_sll_451_U85 ( .A1(u4_sll_451_ML_int_4__3_), .A2(u4_sll_451_n7), 
        .ZN(u4_sll_451_n44) );
  INV_X1 u4_sll_451_U84 ( .A(u4_sll_451_n44), .ZN(u4_sll_451_ML_int_5__3_) );
  NAND2_X1 u4_sll_451_U83 ( .A1(u4_sll_451_ML_int_4__4_), .A2(u4_sll_451_n7), 
        .ZN(u4_sll_451_n43) );
  INV_X1 u4_sll_451_U82 ( .A(u4_sll_451_n43), .ZN(u4_sll_451_ML_int_5__4_) );
  NAND2_X1 u4_sll_451_U81 ( .A1(u4_sll_451_ML_int_4__5_), .A2(u4_sll_451_n7), 
        .ZN(u4_sll_451_n42) );
  INV_X1 u4_sll_451_U80 ( .A(u4_sll_451_n42), .ZN(u4_sll_451_ML_int_5__5_) );
  NAND2_X1 u4_sll_451_U79 ( .A1(u4_sll_451_ML_int_4__6_), .A2(u4_sll_451_n7), 
        .ZN(u4_sll_451_n41) );
  INV_X1 u4_sll_451_U78 ( .A(u4_sll_451_n41), .ZN(u4_sll_451_ML_int_5__6_) );
  NAND2_X1 u4_sll_451_U77 ( .A1(u4_sll_451_ML_int_4__7_), .A2(u4_sll_451_n7), 
        .ZN(u4_sll_451_n40) );
  INV_X1 u4_sll_451_U76 ( .A(u4_sll_451_n40), .ZN(u4_sll_451_ML_int_5__7_) );
  NAND2_X1 u4_sll_451_U75 ( .A1(u4_sll_451_ML_int_4__8_), .A2(u4_sll_451_n7), 
        .ZN(u4_sll_451_n39) );
  INV_X1 u4_sll_451_U74 ( .A(u4_sll_451_n39), .ZN(u4_sll_451_ML_int_5__8_) );
  NAND2_X1 u4_sll_451_U73 ( .A1(u4_sll_451_ML_int_4__9_), .A2(u4_sll_451_n7), 
        .ZN(u4_sll_451_n38) );
  INV_X1 u4_sll_451_U72 ( .A(u4_sll_451_n38), .ZN(u4_sll_451_ML_int_5__9_) );
  NOR2_X1 u4_sll_451_U71 ( .A1(u4_sll_451_n2), .A2(u4_sll_451_n53), .ZN(
        u4_N1408) );
  NOR2_X1 u4_sll_451_U70 ( .A1(u4_sll_451_n2), .A2(u4_sll_451_n52), .ZN(
        u4_N1418) );
  NOR2_X1 u4_sll_451_U69 ( .A1(u4_sll_451_n2), .A2(u4_sll_451_n51), .ZN(
        u4_N1419) );
  NOR2_X1 u4_sll_451_U68 ( .A1(u4_sll_451_n2), .A2(u4_sll_451_n50), .ZN(
        u4_N1420) );
  NOR2_X1 u4_sll_451_U67 ( .A1(u4_sll_451_n2), .A2(u4_sll_451_n49), .ZN(
        u4_N1421) );
  NOR2_X1 u4_sll_451_U66 ( .A1(u4_sll_451_n2), .A2(u4_sll_451_n48), .ZN(
        u4_N1422) );
  NOR2_X1 u4_sll_451_U65 ( .A1(u4_sll_451_n2), .A2(u4_sll_451_n47), .ZN(
        u4_N1423) );
  AND2_X1 u4_sll_451_U64 ( .A1(u4_sll_451_ML_int_5__16_), .A2(u4_sll_451_n3), 
        .ZN(u4_N1424) );
  AND2_X1 u4_sll_451_U63 ( .A1(u4_sll_451_ML_int_5__17_), .A2(u4_sll_451_n1), 
        .ZN(u4_N1425) );
  AND2_X1 u4_sll_451_U62 ( .A1(u4_sll_451_ML_int_5__18_), .A2(u4_sll_451_n1), 
        .ZN(u4_N1426) );
  AND2_X1 u4_sll_451_U61 ( .A1(u4_sll_451_ML_int_5__19_), .A2(u4_sll_451_n3), 
        .ZN(u4_N1427) );
  NOR2_X1 u4_sll_451_U60 ( .A1(u4_sll_451_n2), .A2(u4_sll_451_n46), .ZN(
        u4_N1409) );
  AND2_X1 u4_sll_451_U59 ( .A1(u4_sll_451_ML_int_5__20_), .A2(u4_sll_451_n1), 
        .ZN(u4_N1428) );
  AND2_X1 u4_sll_451_U58 ( .A1(u4_sll_451_ML_int_5__21_), .A2(u4_sll_451_n1), 
        .ZN(u4_N1429) );
  AND2_X1 u4_sll_451_U57 ( .A1(u4_sll_451_ML_int_5__22_), .A2(u4_sll_451_n3), 
        .ZN(u4_N1430) );
  AND2_X1 u4_sll_451_U56 ( .A1(u4_sll_451_ML_int_5__23_), .A2(u4_sll_451_n3), 
        .ZN(u4_N1431) );
  AND2_X1 u4_sll_451_U55 ( .A1(u4_sll_451_ML_int_5__24_), .A2(u4_sll_451_n1), 
        .ZN(u4_N1432) );
  AND2_X1 u4_sll_451_U54 ( .A1(u4_sll_451_ML_int_5__25_), .A2(u4_sll_451_n1), 
        .ZN(u4_N1433) );
  AND2_X1 u4_sll_451_U53 ( .A1(u4_sll_451_ML_int_5__26_), .A2(u4_sll_451_n3), 
        .ZN(u4_N1434) );
  AND2_X1 u4_sll_451_U52 ( .A1(u4_sll_451_ML_int_5__27_), .A2(u4_sll_451_n3), 
        .ZN(u4_N1435) );
  AND2_X1 u4_sll_451_U51 ( .A1(u4_sll_451_ML_int_5__28_), .A2(u4_sll_451_n3), 
        .ZN(u4_N1436) );
  AND2_X1 u4_sll_451_U50 ( .A1(u4_sll_451_ML_int_5__29_), .A2(u4_sll_451_n3), 
        .ZN(u4_N1437) );
  NOR2_X1 u4_sll_451_U49 ( .A1(u4_sll_451_n2), .A2(u4_sll_451_n45), .ZN(
        u4_N1410) );
  AND2_X1 u4_sll_451_U48 ( .A1(u4_sll_451_ML_int_5__30_), .A2(u4_sll_451_n3), 
        .ZN(u4_N1438) );
  AND2_X1 u4_sll_451_U47 ( .A1(u4_sll_451_ML_int_5__31_), .A2(u4_sll_451_n3), 
        .ZN(u4_N1439) );
  NOR2_X1 u4_sll_451_U46 ( .A1(u4_sll_451_n2), .A2(u4_sll_451_n44), .ZN(
        u4_N1411) );
  NOR2_X1 u4_sll_451_U45 ( .A1(u4_sll_451_n2), .A2(u4_sll_451_n43), .ZN(
        u4_N1412) );
  NOR2_X1 u4_sll_451_U44 ( .A1(u4_sll_451_n2), .A2(u4_sll_451_n42), .ZN(
        u4_N1413) );
  NOR2_X1 u4_sll_451_U43 ( .A1(u4_sll_451_n2), .A2(u4_sll_451_n41), .ZN(
        u4_N1414) );
  NOR2_X1 u4_sll_451_U42 ( .A1(u4_sll_451_n2), .A2(u4_sll_451_n40), .ZN(
        u4_N1415) );
  NOR2_X1 u4_sll_451_U41 ( .A1(u4_sll_451_n2), .A2(u4_sll_451_n39), .ZN(
        u4_N1416) );
  NOR2_X1 u4_sll_451_U40 ( .A1(u4_sll_451_n2), .A2(u4_sll_451_n38), .ZN(
        u4_N1417) );
  INV_X4 u4_sll_451_U39 ( .A(u4_sll_451_n3), .ZN(u4_sll_451_n2) );
  INV_X4 u4_sll_451_U38 ( .A(u4_shift_left[5]), .ZN(u4_sll_451_n3) );
  INV_X4 u4_sll_451_U37 ( .A(u4_sll_451_n12), .ZN(u4_sll_451_n19) );
  INV_X4 u4_sll_451_U36 ( .A(u4_sll_451_n31), .ZN(u4_sll_451_n30) );
  INV_X4 u4_sll_451_U35 ( .A(u4_shift_left[1]), .ZN(u4_sll_451_n31) );
  INV_X4 u4_sll_451_U34 ( .A(u4_sll_451_n37), .ZN(u4_sll_451_n36) );
  INV_X4 u4_sll_451_U33 ( .A(u4_sll_451_n32), .ZN(u4_sll_451_n37) );
  INV_X4 u4_sll_451_U32 ( .A(u4_sll_451_n24), .ZN(u4_sll_451_n23) );
  INV_X4 u4_sll_451_U31 ( .A(u4_sll_451_n21), .ZN(u4_sll_451_n25) );
  INV_X4 u4_sll_451_U30 ( .A(u4_sll_451_n18), .ZN(u4_sll_451_n15) );
  INV_X4 u4_sll_451_U29 ( .A(u4_shift_left[5]), .ZN(u4_sll_451_n1) );
  INV_X4 u4_sll_451_U28 ( .A(u4_sll_451_n11), .ZN(u4_sll_451_n10) );
  INV_X4 u4_sll_451_U27 ( .A(u4_sll_451_n8), .ZN(u4_sll_451_n6) );
  INV_X4 u4_sll_451_U26 ( .A(u4_sll_451_n5), .ZN(u4_sll_451_n4) );
  INV_X4 u4_sll_451_U25 ( .A(u4_sll_451_n28), .ZN(u4_sll_451_n27) );
  INV_X4 u4_sll_451_U24 ( .A(u4_sll_451_n20), .ZN(u4_sll_451_n28) );
  INV_X4 u4_sll_451_U23 ( .A(u4_sll_451_n31), .ZN(u4_sll_451_n29) );
  INV_X4 u4_sll_451_U22 ( .A(u4_sll_451_n11), .ZN(u4_sll_451_n8) );
  INV_X4 u4_sll_451_U21 ( .A(u4_sll_451_n17), .ZN(u4_sll_451_n14) );
  INV_X4 u4_sll_451_U20 ( .A(u4_sll_451_n21), .ZN(u4_sll_451_n24) );
  INV_X4 u4_sll_451_U19 ( .A(u4_sll_451_n33), .ZN(u4_sll_451_n34) );
  INV_X4 u4_sll_451_U18 ( .A(u4_sll_451_n18), .ZN(u4_sll_451_n17) );
  INV_X4 u4_sll_451_U17 ( .A(u4_sll_451_n10), .ZN(u4_sll_451_n7) );
  INV_X4 u4_sll_451_U16 ( .A(u4_shift_left[2]), .ZN(u4_sll_451_n21) );
  INV_X4 u4_sll_451_U15 ( .A(u4_sll_451_n21), .ZN(u4_sll_451_n20) );
  INV_X4 u4_sll_451_U14 ( .A(u4_shift_left[0]), .ZN(u4_sll_451_n33) );
  INV_X4 u4_sll_451_U13 ( .A(u4_sll_451_n33), .ZN(u4_sll_451_n32) );
  INV_X4 u4_sll_451_U12 ( .A(u4_sll_451_n11), .ZN(u4_sll_451_n9) );
  INV_X4 u4_sll_451_U11 ( .A(u4_shift_left[4]), .ZN(u4_sll_451_n5) );
  INV_X4 u4_sll_451_U10 ( .A(u4_sll_451_n4), .ZN(u4_sll_451_n11) );
  INV_X4 u4_sll_451_U9 ( .A(u4_sll_451_n18), .ZN(u4_sll_451_n16) );
  INV_X4 u4_sll_451_U8 ( .A(u4_sll_451_n12), .ZN(u4_sll_451_n18) );
  INV_X4 u4_sll_451_U7 ( .A(u4_sll_451_n28), .ZN(u4_sll_451_n26) );
  INV_X4 u4_sll_451_U6 ( .A(u4_sll_451_n25), .ZN(u4_sll_451_n22) );
  INV_X4 u4_sll_451_U5 ( .A(u4_shift_left[3]), .ZN(u4_sll_451_n13) );
  INV_X4 u4_sll_451_U4 ( .A(u4_sll_451_n13), .ZN(u4_sll_451_n12) );
  INV_X4 u4_sll_451_U3 ( .A(u4_sll_451_n37), .ZN(u4_sll_451_n35) );
  MUX2_X2 u4_sll_451_M1_0_1 ( .A(n3521), .B(n3564), .S(u4_sll_451_n34), .Z(
        u4_sll_451_ML_int_1__1_) );
  MUX2_X2 u4_sll_451_M1_0_2 ( .A(n3522), .B(n3521), .S(u4_sll_451_n34), .Z(
        u4_sll_451_ML_int_1__2_) );
  MUX2_X2 u4_sll_451_M1_0_3 ( .A(n3563), .B(n3522), .S(u4_sll_451_n34), .Z(
        u4_sll_451_ML_int_1__3_) );
  MUX2_X2 u4_sll_451_M1_0_4 ( .A(n3523), .B(n3563), .S(u4_sll_451_n34), .Z(
        u4_sll_451_ML_int_1__4_) );
  MUX2_X2 u4_sll_451_M1_0_5 ( .A(n3524), .B(n3523), .S(u4_sll_451_n34), .Z(
        u4_sll_451_ML_int_1__5_) );
  MUX2_X2 u4_sll_451_M1_0_6 ( .A(n3562), .B(n3524), .S(u4_sll_451_n34), .Z(
        u4_sll_451_ML_int_1__6_) );
  MUX2_X2 u4_sll_451_M1_0_7 ( .A(n3525), .B(n3562), .S(u4_sll_451_n35), .Z(
        u4_sll_451_ML_int_1__7_) );
  MUX2_X2 u4_sll_451_M1_0_8 ( .A(n3526), .B(n3525), .S(u4_sll_451_n35), .Z(
        u4_sll_451_ML_int_1__8_) );
  MUX2_X2 u4_sll_451_M1_0_9 ( .A(n3528), .B(n3526), .S(u4_sll_451_n35), .Z(
        u4_sll_451_ML_int_1__9_) );
  MUX2_X2 u4_sll_451_M1_0_10 ( .A(n3527), .B(n3528), .S(u4_sll_451_n35), .Z(
        u4_sll_451_ML_int_1__10_) );
  MUX2_X2 u4_sll_451_M1_0_11 ( .A(n3561), .B(n3527), .S(u4_sll_451_n35), .Z(
        u4_sll_451_ML_int_1__11_) );
  MUX2_X2 u4_sll_451_M1_0_12 ( .A(n3529), .B(n3561), .S(u4_sll_451_n35), .Z(
        u4_sll_451_ML_int_1__12_) );
  MUX2_X2 u4_sll_451_M1_0_13 ( .A(n3530), .B(n3529), .S(u4_sll_451_n35), .Z(
        u4_sll_451_ML_int_1__13_) );
  MUX2_X2 u4_sll_451_M1_0_14 ( .A(n3560), .B(n3530), .S(u4_sll_451_n35), .Z(
        u4_sll_451_ML_int_1__14_) );
  MUX2_X2 u4_sll_451_M1_0_15 ( .A(n3531), .B(n3560), .S(u4_sll_451_n35), .Z(
        u4_sll_451_ML_int_1__15_) );
  MUX2_X2 u4_sll_451_M1_0_16 ( .A(n3532), .B(n3531), .S(u4_sll_451_n35), .Z(
        u4_sll_451_ML_int_1__16_) );
  MUX2_X2 u4_sll_451_M1_0_17 ( .A(n3559), .B(n3532), .S(u4_sll_451_n35), .Z(
        u4_sll_451_ML_int_1__17_) );
  MUX2_X2 u4_sll_451_M1_0_18 ( .A(n3533), .B(n3559), .S(u4_sll_451_n35), .Z(
        u4_sll_451_ML_int_1__18_) );
  MUX2_X2 u4_sll_451_M1_0_19 ( .A(n3534), .B(n3533), .S(u4_sll_451_n35), .Z(
        u4_sll_451_ML_int_1__19_) );
  MUX2_X2 u4_sll_451_M1_0_20 ( .A(n3557), .B(n3534), .S(u4_sll_451_n35), .Z(
        u4_sll_451_ML_int_1__20_) );
  MUX2_X2 u4_sll_451_M1_0_21 ( .A(fract_denorm[21]), .B(n3557), .S(
        u4_sll_451_n35), .Z(u4_sll_451_ML_int_1__21_) );
  MUX2_X2 u4_sll_451_M1_0_22 ( .A(fract_denorm[22]), .B(fract_denorm[21]), .S(
        u4_sll_451_n35), .Z(u4_sll_451_ML_int_1__22_) );
  MUX2_X2 u4_sll_451_M1_0_23 ( .A(fract_denorm[23]), .B(fract_denorm[22]), .S(
        u4_sll_451_n35), .Z(u4_sll_451_ML_int_1__23_) );
  MUX2_X2 u4_sll_451_M1_0_24 ( .A(fract_denorm[24]), .B(fract_denorm[23]), .S(
        u4_sll_451_n35), .Z(u4_sll_451_ML_int_1__24_) );
  MUX2_X2 u4_sll_451_M1_0_25 ( .A(fract_denorm[25]), .B(fract_denorm[24]), .S(
        u4_sll_451_n36), .Z(u4_sll_451_ML_int_1__25_) );
  MUX2_X2 u4_sll_451_M1_0_26 ( .A(fract_denorm[26]), .B(fract_denorm[25]), .S(
        u4_sll_451_n36), .Z(u4_sll_451_ML_int_1__26_) );
  MUX2_X2 u4_sll_451_M1_0_27 ( .A(fract_denorm[27]), .B(fract_denorm[26]), .S(
        u4_sll_451_n36), .Z(u4_sll_451_ML_int_1__27_) );
  MUX2_X2 u4_sll_451_M1_0_28 ( .A(fract_denorm[28]), .B(fract_denorm[27]), .S(
        u4_sll_451_n36), .Z(u4_sll_451_ML_int_1__28_) );
  MUX2_X2 u4_sll_451_M1_0_29 ( .A(fract_denorm[29]), .B(fract_denorm[28]), .S(
        u4_sll_451_n36), .Z(u4_sll_451_ML_int_1__29_) );
  MUX2_X2 u4_sll_451_M1_0_30 ( .A(fract_denorm[30]), .B(fract_denorm[29]), .S(
        u4_sll_451_n36), .Z(u4_sll_451_ML_int_1__30_) );
  MUX2_X2 u4_sll_451_M1_0_31 ( .A(fract_denorm[31]), .B(fract_denorm[30]), .S(
        u4_sll_451_n36), .Z(u4_sll_451_ML_int_1__31_) );
  MUX2_X2 u4_sll_451_M1_0_32 ( .A(fract_denorm[32]), .B(fract_denorm[31]), .S(
        u4_sll_451_n36), .Z(u4_sll_451_ML_int_1__32_) );
  MUX2_X2 u4_sll_451_M1_0_33 ( .A(fract_denorm[33]), .B(fract_denorm[32]), .S(
        u4_sll_451_n36), .Z(u4_sll_451_ML_int_1__33_) );
  MUX2_X2 u4_sll_451_M1_0_34 ( .A(fract_denorm[34]), .B(fract_denorm[33]), .S(
        u4_sll_451_n36), .Z(u4_sll_451_ML_int_1__34_) );
  MUX2_X2 u4_sll_451_M1_0_35 ( .A(fract_denorm[35]), .B(fract_denorm[34]), .S(
        u4_sll_451_n36), .Z(u4_sll_451_ML_int_1__35_) );
  MUX2_X2 u4_sll_451_M1_0_36 ( .A(fract_denorm[36]), .B(fract_denorm[35]), .S(
        u4_sll_451_n36), .Z(u4_sll_451_ML_int_1__36_) );
  MUX2_X2 u4_sll_451_M1_0_37 ( .A(fract_denorm[37]), .B(fract_denorm[36]), .S(
        u4_sll_451_n36), .Z(u4_sll_451_ML_int_1__37_) );
  MUX2_X2 u4_sll_451_M1_0_38 ( .A(fract_denorm[38]), .B(fract_denorm[37]), .S(
        u4_sll_451_n36), .Z(u4_sll_451_ML_int_1__38_) );
  MUX2_X2 u4_sll_451_M1_0_39 ( .A(fract_denorm[39]), .B(fract_denorm[38]), .S(
        u4_sll_451_n36), .Z(u4_sll_451_ML_int_1__39_) );
  MUX2_X2 u4_sll_451_M1_0_40 ( .A(fract_denorm[40]), .B(fract_denorm[39]), .S(
        u4_sll_451_n36), .Z(u4_sll_451_ML_int_1__40_) );
  MUX2_X2 u4_sll_451_M1_0_41 ( .A(fract_denorm[41]), .B(fract_denorm[40]), .S(
        u4_sll_451_n36), .Z(u4_sll_451_ML_int_1__41_) );
  MUX2_X2 u4_sll_451_M1_0_42 ( .A(fract_denorm[42]), .B(fract_denorm[41]), .S(
        u4_sll_451_n36), .Z(u4_sll_451_ML_int_1__42_) );
  MUX2_X2 u4_sll_451_M1_0_43 ( .A(fract_denorm[43]), .B(fract_denorm[42]), .S(
        u4_sll_451_n36), .Z(u4_sll_451_ML_int_1__43_) );
  MUX2_X2 u4_sll_451_M1_0_44 ( .A(fract_denorm[44]), .B(fract_denorm[43]), .S(
        u4_sll_451_n36), .Z(u4_sll_451_ML_int_1__44_) );
  MUX2_X2 u4_sll_451_M1_0_45 ( .A(fract_denorm[45]), .B(fract_denorm[44]), .S(
        u4_sll_451_n36), .Z(u4_sll_451_ML_int_1__45_) );
  MUX2_X2 u4_sll_451_M1_0_46 ( .A(fract_denorm[46]), .B(fract_denorm[45]), .S(
        u4_sll_451_n36), .Z(u4_sll_451_ML_int_1__46_) );
  MUX2_X2 u4_sll_451_M1_0_47 ( .A(n2679), .B(fract_denorm[46]), .S(
        u4_sll_451_n36), .Z(u4_sll_451_ML_int_1__47_) );
  MUX2_X2 u4_sll_451_M1_1_2 ( .A(u4_sll_451_ML_int_1__2_), .B(
        u4_sll_451_ML_int_1__0_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__2_) );
  MUX2_X2 u4_sll_451_M1_1_3 ( .A(u4_sll_451_ML_int_1__3_), .B(
        u4_sll_451_ML_int_1__1_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__3_) );
  MUX2_X2 u4_sll_451_M1_1_4 ( .A(u4_sll_451_ML_int_1__4_), .B(
        u4_sll_451_ML_int_1__2_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__4_) );
  MUX2_X2 u4_sll_451_M1_1_5 ( .A(u4_sll_451_ML_int_1__5_), .B(
        u4_sll_451_ML_int_1__3_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__5_) );
  MUX2_X2 u4_sll_451_M1_1_6 ( .A(u4_sll_451_ML_int_1__6_), .B(
        u4_sll_451_ML_int_1__4_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__6_) );
  MUX2_X2 u4_sll_451_M1_1_7 ( .A(u4_sll_451_ML_int_1__7_), .B(
        u4_sll_451_ML_int_1__5_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__7_) );
  MUX2_X2 u4_sll_451_M1_1_8 ( .A(u4_sll_451_ML_int_1__8_), .B(
        u4_sll_451_ML_int_1__6_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__8_) );
  MUX2_X2 u4_sll_451_M1_1_9 ( .A(u4_sll_451_ML_int_1__9_), .B(
        u4_sll_451_ML_int_1__7_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__9_) );
  MUX2_X2 u4_sll_451_M1_1_10 ( .A(u4_sll_451_ML_int_1__10_), .B(
        u4_sll_451_ML_int_1__8_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__10_) );
  MUX2_X2 u4_sll_451_M1_1_11 ( .A(u4_sll_451_ML_int_1__11_), .B(
        u4_sll_451_ML_int_1__9_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__11_) );
  MUX2_X2 u4_sll_451_M1_1_12 ( .A(u4_sll_451_ML_int_1__12_), .B(
        u4_sll_451_ML_int_1__10_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__12_) );
  MUX2_X2 u4_sll_451_M1_1_13 ( .A(u4_sll_451_ML_int_1__13_), .B(
        u4_sll_451_ML_int_1__11_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__13_) );
  MUX2_X2 u4_sll_451_M1_1_14 ( .A(u4_sll_451_ML_int_1__14_), .B(
        u4_sll_451_ML_int_1__12_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__14_) );
  MUX2_X2 u4_sll_451_M1_1_15 ( .A(u4_sll_451_ML_int_1__15_), .B(
        u4_sll_451_ML_int_1__13_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__15_) );
  MUX2_X2 u4_sll_451_M1_1_16 ( .A(u4_sll_451_ML_int_1__16_), .B(
        u4_sll_451_ML_int_1__14_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__16_) );
  MUX2_X2 u4_sll_451_M1_1_17 ( .A(u4_sll_451_ML_int_1__17_), .B(
        u4_sll_451_ML_int_1__15_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__17_) );
  MUX2_X2 u4_sll_451_M1_1_18 ( .A(u4_sll_451_ML_int_1__18_), .B(
        u4_sll_451_ML_int_1__16_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__18_) );
  MUX2_X2 u4_sll_451_M1_1_19 ( .A(u4_sll_451_ML_int_1__19_), .B(
        u4_sll_451_ML_int_1__17_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__19_) );
  MUX2_X2 u4_sll_451_M1_1_20 ( .A(u4_sll_451_ML_int_1__20_), .B(
        u4_sll_451_ML_int_1__18_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__20_) );
  MUX2_X2 u4_sll_451_M1_1_21 ( .A(u4_sll_451_ML_int_1__21_), .B(
        u4_sll_451_ML_int_1__19_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__21_) );
  MUX2_X2 u4_sll_451_M1_1_22 ( .A(u4_sll_451_ML_int_1__22_), .B(
        u4_sll_451_ML_int_1__20_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__22_) );
  MUX2_X2 u4_sll_451_M1_1_23 ( .A(u4_sll_451_ML_int_1__23_), .B(
        u4_sll_451_ML_int_1__21_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__23_) );
  MUX2_X2 u4_sll_451_M1_1_24 ( .A(u4_sll_451_ML_int_1__24_), .B(
        u4_sll_451_ML_int_1__22_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__24_) );
  MUX2_X2 u4_sll_451_M1_1_25 ( .A(u4_sll_451_ML_int_1__25_), .B(
        u4_sll_451_ML_int_1__23_), .S(u4_sll_451_n29), .Z(
        u4_sll_451_ML_int_2__25_) );
  MUX2_X2 u4_sll_451_M1_1_26 ( .A(u4_sll_451_ML_int_1__26_), .B(
        u4_sll_451_ML_int_1__24_), .S(u4_sll_451_n30), .Z(
        u4_sll_451_ML_int_2__26_) );
  MUX2_X2 u4_sll_451_M1_1_27 ( .A(u4_sll_451_ML_int_1__27_), .B(
        u4_sll_451_ML_int_1__25_), .S(u4_sll_451_n30), .Z(
        u4_sll_451_ML_int_2__27_) );
  MUX2_X2 u4_sll_451_M1_1_28 ( .A(u4_sll_451_ML_int_1__28_), .B(
        u4_sll_451_ML_int_1__26_), .S(u4_sll_451_n30), .Z(
        u4_sll_451_ML_int_2__28_) );
  MUX2_X2 u4_sll_451_M1_1_29 ( .A(u4_sll_451_ML_int_1__29_), .B(
        u4_sll_451_ML_int_1__27_), .S(u4_sll_451_n30), .Z(
        u4_sll_451_ML_int_2__29_) );
  MUX2_X2 u4_sll_451_M1_1_30 ( .A(u4_sll_451_ML_int_1__30_), .B(
        u4_sll_451_ML_int_1__28_), .S(u4_sll_451_n30), .Z(
        u4_sll_451_ML_int_2__30_) );
  MUX2_X2 u4_sll_451_M1_1_31 ( .A(u4_sll_451_ML_int_1__31_), .B(
        u4_sll_451_ML_int_1__29_), .S(u4_sll_451_n30), .Z(
        u4_sll_451_ML_int_2__31_) );
  MUX2_X2 u4_sll_451_M1_1_32 ( .A(u4_sll_451_ML_int_1__32_), .B(
        u4_sll_451_ML_int_1__30_), .S(u4_sll_451_n30), .Z(
        u4_sll_451_ML_int_2__32_) );
  MUX2_X2 u4_sll_451_M1_1_33 ( .A(u4_sll_451_ML_int_1__33_), .B(
        u4_sll_451_ML_int_1__31_), .S(u4_sll_451_n30), .Z(
        u4_sll_451_ML_int_2__33_) );
  MUX2_X2 u4_sll_451_M1_1_34 ( .A(u4_sll_451_ML_int_1__34_), .B(
        u4_sll_451_ML_int_1__32_), .S(u4_sll_451_n30), .Z(
        u4_sll_451_ML_int_2__34_) );
  MUX2_X2 u4_sll_451_M1_1_35 ( .A(u4_sll_451_ML_int_1__35_), .B(
        u4_sll_451_ML_int_1__33_), .S(u4_sll_451_n30), .Z(
        u4_sll_451_ML_int_2__35_) );
  MUX2_X2 u4_sll_451_M1_1_36 ( .A(u4_sll_451_ML_int_1__36_), .B(
        u4_sll_451_ML_int_1__34_), .S(u4_sll_451_n30), .Z(
        u4_sll_451_ML_int_2__36_) );
  MUX2_X2 u4_sll_451_M1_1_37 ( .A(u4_sll_451_ML_int_1__37_), .B(
        u4_sll_451_ML_int_1__35_), .S(u4_sll_451_n30), .Z(
        u4_sll_451_ML_int_2__37_) );
  MUX2_X2 u4_sll_451_M1_1_38 ( .A(u4_sll_451_ML_int_1__38_), .B(
        u4_sll_451_ML_int_1__36_), .S(u4_sll_451_n30), .Z(
        u4_sll_451_ML_int_2__38_) );
  MUX2_X2 u4_sll_451_M1_1_39 ( .A(u4_sll_451_ML_int_1__39_), .B(
        u4_sll_451_ML_int_1__37_), .S(u4_sll_451_n30), .Z(
        u4_sll_451_ML_int_2__39_) );
  MUX2_X2 u4_sll_451_M1_1_40 ( .A(u4_sll_451_ML_int_1__40_), .B(
        u4_sll_451_ML_int_1__38_), .S(u4_sll_451_n30), .Z(
        u4_sll_451_ML_int_2__40_) );
  MUX2_X2 u4_sll_451_M1_1_41 ( .A(u4_sll_451_ML_int_1__41_), .B(
        u4_sll_451_ML_int_1__39_), .S(u4_sll_451_n30), .Z(
        u4_sll_451_ML_int_2__41_) );
  MUX2_X2 u4_sll_451_M1_1_42 ( .A(u4_sll_451_ML_int_1__42_), .B(
        u4_sll_451_ML_int_1__40_), .S(u4_sll_451_n30), .Z(
        u4_sll_451_ML_int_2__42_) );
  MUX2_X2 u4_sll_451_M1_1_43 ( .A(u4_sll_451_ML_int_1__43_), .B(
        u4_sll_451_ML_int_1__41_), .S(u4_sll_451_n30), .Z(
        u4_sll_451_ML_int_2__43_) );
  MUX2_X2 u4_sll_451_M1_1_44 ( .A(u4_sll_451_ML_int_1__44_), .B(
        u4_sll_451_ML_int_1__42_), .S(u4_sll_451_n30), .Z(
        u4_sll_451_ML_int_2__44_) );
  MUX2_X2 u4_sll_451_M1_1_45 ( .A(u4_sll_451_ML_int_1__45_), .B(
        u4_sll_451_ML_int_1__43_), .S(u4_sll_451_n30), .Z(
        u4_sll_451_ML_int_2__45_) );
  MUX2_X2 u4_sll_451_M1_1_46 ( .A(u4_sll_451_ML_int_1__46_), .B(
        u4_sll_451_ML_int_1__44_), .S(u4_sll_451_n30), .Z(
        u4_sll_451_ML_int_2__46_) );
  MUX2_X2 u4_sll_451_M1_1_47 ( .A(u4_sll_451_ML_int_1__47_), .B(
        u4_sll_451_ML_int_1__45_), .S(u4_sll_451_n30), .Z(
        u4_sll_451_ML_int_2__47_) );
  MUX2_X2 u4_sll_451_M1_2_4 ( .A(u4_sll_451_ML_int_2__4_), .B(
        u4_sll_451_ML_int_2__0_), .S(u4_sll_451_n25), .Z(
        u4_sll_451_ML_int_3__4_) );
  MUX2_X2 u4_sll_451_M1_2_5 ( .A(u4_sll_451_ML_int_2__5_), .B(
        u4_sll_451_ML_int_2__1_), .S(u4_sll_451_n25), .Z(
        u4_sll_451_ML_int_3__5_) );
  MUX2_X2 u4_sll_451_M1_2_6 ( .A(u4_sll_451_ML_int_2__6_), .B(
        u4_sll_451_ML_int_2__2_), .S(u4_sll_451_n25), .Z(
        u4_sll_451_ML_int_3__6_) );
  MUX2_X2 u4_sll_451_M1_2_7 ( .A(u4_sll_451_ML_int_2__7_), .B(
        u4_sll_451_ML_int_2__3_), .S(u4_sll_451_n25), .Z(
        u4_sll_451_ML_int_3__7_) );
  MUX2_X2 u4_sll_451_M1_2_8 ( .A(u4_sll_451_ML_int_2__8_), .B(
        u4_sll_451_ML_int_2__4_), .S(u4_sll_451_n25), .Z(
        u4_sll_451_ML_int_3__8_) );
  MUX2_X2 u4_sll_451_M1_2_9 ( .A(u4_sll_451_ML_int_2__9_), .B(
        u4_sll_451_ML_int_2__5_), .S(u4_sll_451_n25), .Z(
        u4_sll_451_ML_int_3__9_) );
  MUX2_X2 u4_sll_451_M1_2_10 ( .A(u4_sll_451_ML_int_2__10_), .B(
        u4_sll_451_ML_int_2__6_), .S(u4_sll_451_n26), .Z(
        u4_sll_451_ML_int_3__10_) );
  MUX2_X2 u4_sll_451_M1_2_11 ( .A(u4_sll_451_ML_int_2__11_), .B(
        u4_sll_451_ML_int_2__7_), .S(u4_sll_451_n26), .Z(
        u4_sll_451_ML_int_3__11_) );
  MUX2_X2 u4_sll_451_M1_2_12 ( .A(u4_sll_451_ML_int_2__12_), .B(
        u4_sll_451_ML_int_2__8_), .S(u4_sll_451_n26), .Z(
        u4_sll_451_ML_int_3__12_) );
  MUX2_X2 u4_sll_451_M1_2_13 ( .A(u4_sll_451_ML_int_2__13_), .B(
        u4_sll_451_ML_int_2__9_), .S(u4_sll_451_n26), .Z(
        u4_sll_451_ML_int_3__13_) );
  MUX2_X2 u4_sll_451_M1_2_14 ( .A(u4_sll_451_ML_int_2__14_), .B(
        u4_sll_451_ML_int_2__10_), .S(u4_sll_451_n26), .Z(
        u4_sll_451_ML_int_3__14_) );
  MUX2_X2 u4_sll_451_M1_2_15 ( .A(u4_sll_451_ML_int_2__15_), .B(
        u4_sll_451_ML_int_2__11_), .S(u4_sll_451_n26), .Z(
        u4_sll_451_ML_int_3__15_) );
  MUX2_X2 u4_sll_451_M1_2_16 ( .A(u4_sll_451_ML_int_2__16_), .B(
        u4_sll_451_ML_int_2__12_), .S(u4_sll_451_n26), .Z(
        u4_sll_451_ML_int_3__16_) );
  MUX2_X2 u4_sll_451_M1_2_17 ( .A(u4_sll_451_ML_int_2__17_), .B(
        u4_sll_451_ML_int_2__13_), .S(u4_sll_451_n26), .Z(
        u4_sll_451_ML_int_3__17_) );
  MUX2_X2 u4_sll_451_M1_2_18 ( .A(u4_sll_451_ML_int_2__18_), .B(
        u4_sll_451_ML_int_2__14_), .S(u4_sll_451_n26), .Z(
        u4_sll_451_ML_int_3__18_) );
  MUX2_X2 u4_sll_451_M1_2_19 ( .A(u4_sll_451_ML_int_2__19_), .B(
        u4_sll_451_ML_int_2__15_), .S(u4_sll_451_n26), .Z(
        u4_sll_451_ML_int_3__19_) );
  MUX2_X2 u4_sll_451_M1_2_20 ( .A(u4_sll_451_ML_int_2__20_), .B(
        u4_sll_451_ML_int_2__16_), .S(u4_sll_451_n26), .Z(
        u4_sll_451_ML_int_3__20_) );
  MUX2_X2 u4_sll_451_M1_2_21 ( .A(u4_sll_451_ML_int_2__21_), .B(
        u4_sll_451_ML_int_2__17_), .S(u4_sll_451_n26), .Z(
        u4_sll_451_ML_int_3__21_) );
  MUX2_X2 u4_sll_451_M1_2_22 ( .A(u4_sll_451_ML_int_2__22_), .B(
        u4_sll_451_ML_int_2__18_), .S(u4_sll_451_n26), .Z(
        u4_sll_451_ML_int_3__22_) );
  MUX2_X2 u4_sll_451_M1_2_23 ( .A(u4_sll_451_ML_int_2__23_), .B(
        u4_sll_451_ML_int_2__19_), .S(u4_sll_451_n26), .Z(
        u4_sll_451_ML_int_3__23_) );
  MUX2_X2 u4_sll_451_M1_2_24 ( .A(u4_sll_451_ML_int_2__24_), .B(
        u4_sll_451_ML_int_2__20_), .S(u4_sll_451_n26), .Z(
        u4_sll_451_ML_int_3__24_) );
  MUX2_X2 u4_sll_451_M1_2_25 ( .A(u4_sll_451_ML_int_2__25_), .B(
        u4_sll_451_ML_int_2__21_), .S(u4_sll_451_n26), .Z(
        u4_sll_451_ML_int_3__25_) );
  MUX2_X2 u4_sll_451_M1_2_26 ( .A(u4_sll_451_ML_int_2__26_), .B(
        u4_sll_451_ML_int_2__22_), .S(u4_sll_451_n26), .Z(
        u4_sll_451_ML_int_3__26_) );
  MUX2_X2 u4_sll_451_M1_2_27 ( .A(u4_sll_451_ML_int_2__27_), .B(
        u4_sll_451_ML_int_2__23_), .S(u4_sll_451_n26), .Z(
        u4_sll_451_ML_int_3__27_) );
  MUX2_X2 u4_sll_451_M1_2_28 ( .A(u4_sll_451_ML_int_2__28_), .B(
        u4_sll_451_ML_int_2__24_), .S(u4_sll_451_n27), .Z(
        u4_sll_451_ML_int_3__28_) );
  MUX2_X2 u4_sll_451_M1_2_29 ( .A(u4_sll_451_ML_int_2__29_), .B(
        u4_sll_451_ML_int_2__25_), .S(u4_sll_451_n27), .Z(
        u4_sll_451_ML_int_3__29_) );
  MUX2_X2 u4_sll_451_M1_2_30 ( .A(u4_sll_451_ML_int_2__30_), .B(
        u4_sll_451_ML_int_2__26_), .S(u4_sll_451_n27), .Z(
        u4_sll_451_ML_int_3__30_) );
  MUX2_X2 u4_sll_451_M1_2_31 ( .A(u4_sll_451_ML_int_2__31_), .B(
        u4_sll_451_ML_int_2__27_), .S(u4_sll_451_n27), .Z(
        u4_sll_451_ML_int_3__31_) );
  MUX2_X2 u4_sll_451_M1_2_32 ( .A(u4_sll_451_ML_int_2__32_), .B(
        u4_sll_451_ML_int_2__28_), .S(u4_sll_451_n27), .Z(
        u4_sll_451_ML_int_3__32_) );
  MUX2_X2 u4_sll_451_M1_2_33 ( .A(u4_sll_451_ML_int_2__33_), .B(
        u4_sll_451_ML_int_2__29_), .S(u4_sll_451_n27), .Z(
        u4_sll_451_ML_int_3__33_) );
  MUX2_X2 u4_sll_451_M1_2_34 ( .A(u4_sll_451_ML_int_2__34_), .B(
        u4_sll_451_ML_int_2__30_), .S(u4_sll_451_n27), .Z(
        u4_sll_451_ML_int_3__34_) );
  MUX2_X2 u4_sll_451_M1_2_35 ( .A(u4_sll_451_ML_int_2__35_), .B(
        u4_sll_451_ML_int_2__31_), .S(u4_sll_451_n27), .Z(
        u4_sll_451_ML_int_3__35_) );
  MUX2_X2 u4_sll_451_M1_2_36 ( .A(u4_sll_451_ML_int_2__36_), .B(
        u4_sll_451_ML_int_2__32_), .S(u4_sll_451_n27), .Z(
        u4_sll_451_ML_int_3__36_) );
  MUX2_X2 u4_sll_451_M1_2_37 ( .A(u4_sll_451_ML_int_2__37_), .B(
        u4_sll_451_ML_int_2__33_), .S(u4_sll_451_n27), .Z(
        u4_sll_451_ML_int_3__37_) );
  MUX2_X2 u4_sll_451_M1_2_38 ( .A(u4_sll_451_ML_int_2__38_), .B(
        u4_sll_451_ML_int_2__34_), .S(u4_sll_451_n27), .Z(
        u4_sll_451_ML_int_3__38_) );
  MUX2_X2 u4_sll_451_M1_2_39 ( .A(u4_sll_451_ML_int_2__39_), .B(
        u4_sll_451_ML_int_2__35_), .S(u4_sll_451_n27), .Z(
        u4_sll_451_ML_int_3__39_) );
  MUX2_X2 u4_sll_451_M1_2_40 ( .A(u4_sll_451_ML_int_2__40_), .B(
        u4_sll_451_ML_int_2__36_), .S(u4_sll_451_n27), .Z(
        u4_sll_451_ML_int_3__40_) );
  MUX2_X2 u4_sll_451_M1_2_41 ( .A(u4_sll_451_ML_int_2__41_), .B(
        u4_sll_451_ML_int_2__37_), .S(u4_sll_451_n27), .Z(
        u4_sll_451_ML_int_3__41_) );
  MUX2_X2 u4_sll_451_M1_2_42 ( .A(u4_sll_451_ML_int_2__42_), .B(
        u4_sll_451_ML_int_2__38_), .S(u4_sll_451_n27), .Z(
        u4_sll_451_ML_int_3__42_) );
  MUX2_X2 u4_sll_451_M1_2_43 ( .A(u4_sll_451_ML_int_2__43_), .B(
        u4_sll_451_ML_int_2__39_), .S(u4_sll_451_n27), .Z(
        u4_sll_451_ML_int_3__43_) );
  MUX2_X2 u4_sll_451_M1_2_44 ( .A(u4_sll_451_ML_int_2__44_), .B(
        u4_sll_451_ML_int_2__40_), .S(u4_sll_451_n27), .Z(
        u4_sll_451_ML_int_3__44_) );
  MUX2_X2 u4_sll_451_M1_2_45 ( .A(u4_sll_451_ML_int_2__45_), .B(
        u4_sll_451_ML_int_2__41_), .S(u4_sll_451_n27), .Z(
        u4_sll_451_ML_int_3__45_) );
  MUX2_X2 u4_sll_451_M1_2_46 ( .A(u4_sll_451_ML_int_2__46_), .B(
        u4_sll_451_ML_int_2__42_), .S(u4_sll_451_n27), .Z(
        u4_sll_451_ML_int_3__46_) );
  MUX2_X2 u4_sll_451_M1_2_47 ( .A(u4_sll_451_ML_int_2__47_), .B(
        u4_sll_451_ML_int_2__43_), .S(u4_sll_451_n27), .Z(
        u4_sll_451_ML_int_3__47_) );
  MUX2_X2 u4_sll_451_M1_3_8 ( .A(u4_sll_451_ML_int_3__8_), .B(
        u4_sll_451_ML_int_3__0_), .S(u4_sll_451_n15), .Z(
        u4_sll_451_ML_int_4__8_) );
  MUX2_X2 u4_sll_451_M1_3_9 ( .A(u4_sll_451_ML_int_3__9_), .B(
        u4_sll_451_ML_int_3__1_), .S(u4_sll_451_n15), .Z(
        u4_sll_451_ML_int_4__9_) );
  MUX2_X2 u4_sll_451_M1_3_10 ( .A(u4_sll_451_ML_int_3__10_), .B(
        u4_sll_451_ML_int_3__2_), .S(u4_sll_451_n15), .Z(
        u4_sll_451_ML_int_4__10_) );
  MUX2_X2 u4_sll_451_M1_3_11 ( .A(u4_sll_451_ML_int_3__11_), .B(
        u4_sll_451_ML_int_3__3_), .S(u4_sll_451_n15), .Z(
        u4_sll_451_ML_int_4__11_) );
  MUX2_X2 u4_sll_451_M1_3_12 ( .A(u4_sll_451_ML_int_3__12_), .B(
        u4_sll_451_ML_int_3__4_), .S(u4_sll_451_n15), .Z(
        u4_sll_451_ML_int_4__12_) );
  MUX2_X2 u4_sll_451_M1_3_13 ( .A(u4_sll_451_ML_int_3__13_), .B(
        u4_sll_451_ML_int_3__5_), .S(u4_sll_451_n15), .Z(
        u4_sll_451_ML_int_4__13_) );
  MUX2_X2 u4_sll_451_M1_3_14 ( .A(u4_sll_451_ML_int_3__14_), .B(
        u4_sll_451_ML_int_3__6_), .S(u4_sll_451_n16), .Z(
        u4_sll_451_ML_int_4__14_) );
  MUX2_X2 u4_sll_451_M1_3_15 ( .A(u4_sll_451_ML_int_3__15_), .B(
        u4_sll_451_ML_int_3__7_), .S(u4_sll_451_n16), .Z(
        u4_sll_451_ML_int_4__15_) );
  MUX2_X2 u4_sll_451_M1_3_16 ( .A(u4_sll_451_ML_int_3__16_), .B(
        u4_sll_451_ML_int_3__8_), .S(u4_sll_451_n16), .Z(
        u4_sll_451_ML_int_4__16_) );
  MUX2_X2 u4_sll_451_M1_3_17 ( .A(u4_sll_451_ML_int_3__17_), .B(
        u4_sll_451_ML_int_3__9_), .S(u4_sll_451_n16), .Z(
        u4_sll_451_ML_int_4__17_) );
  MUX2_X2 u4_sll_451_M1_3_18 ( .A(u4_sll_451_ML_int_3__18_), .B(
        u4_sll_451_ML_int_3__10_), .S(u4_sll_451_n16), .Z(
        u4_sll_451_ML_int_4__18_) );
  MUX2_X2 u4_sll_451_M1_3_19 ( .A(u4_sll_451_ML_int_3__19_), .B(
        u4_sll_451_ML_int_3__11_), .S(u4_sll_451_n16), .Z(
        u4_sll_451_ML_int_4__19_) );
  MUX2_X2 u4_sll_451_M1_3_20 ( .A(u4_sll_451_ML_int_3__20_), .B(
        u4_sll_451_ML_int_3__12_), .S(u4_sll_451_n16), .Z(
        u4_sll_451_ML_int_4__20_) );
  MUX2_X2 u4_sll_451_M1_3_21 ( .A(u4_sll_451_ML_int_3__21_), .B(
        u4_sll_451_ML_int_3__13_), .S(u4_sll_451_n16), .Z(
        u4_sll_451_ML_int_4__21_) );
  MUX2_X2 u4_sll_451_M1_3_22 ( .A(u4_sll_451_ML_int_3__22_), .B(
        u4_sll_451_ML_int_3__14_), .S(u4_sll_451_n16), .Z(
        u4_sll_451_ML_int_4__22_) );
  MUX2_X2 u4_sll_451_M1_3_23 ( .A(u4_sll_451_ML_int_3__23_), .B(
        u4_sll_451_ML_int_3__15_), .S(u4_sll_451_n16), .Z(
        u4_sll_451_ML_int_4__23_) );
  MUX2_X2 u4_sll_451_M1_3_24 ( .A(u4_sll_451_ML_int_3__24_), .B(
        u4_sll_451_ML_int_3__16_), .S(u4_sll_451_n16), .Z(
        u4_sll_451_ML_int_4__24_) );
  MUX2_X2 u4_sll_451_M1_3_25 ( .A(u4_sll_451_ML_int_3__25_), .B(
        u4_sll_451_ML_int_3__17_), .S(u4_sll_451_n16), .Z(
        u4_sll_451_ML_int_4__25_) );
  MUX2_X2 u4_sll_451_M1_3_26 ( .A(u4_sll_451_ML_int_3__26_), .B(
        u4_sll_451_ML_int_3__18_), .S(u4_sll_451_n16), .Z(
        u4_sll_451_ML_int_4__26_) );
  MUX2_X2 u4_sll_451_M1_3_27 ( .A(u4_sll_451_ML_int_3__27_), .B(
        u4_sll_451_ML_int_3__19_), .S(u4_sll_451_n16), .Z(
        u4_sll_451_ML_int_4__27_) );
  MUX2_X2 u4_sll_451_M1_3_28 ( .A(u4_sll_451_ML_int_3__28_), .B(
        u4_sll_451_ML_int_3__20_), .S(u4_sll_451_n16), .Z(
        u4_sll_451_ML_int_4__28_) );
  MUX2_X2 u4_sll_451_M1_3_29 ( .A(u4_sll_451_ML_int_3__29_), .B(
        u4_sll_451_ML_int_3__21_), .S(u4_sll_451_n16), .Z(
        u4_sll_451_ML_int_4__29_) );
  MUX2_X2 u4_sll_451_M1_3_30 ( .A(u4_sll_451_ML_int_3__30_), .B(
        u4_sll_451_ML_int_3__22_), .S(u4_sll_451_n16), .Z(
        u4_sll_451_ML_int_4__30_) );
  MUX2_X2 u4_sll_451_M1_3_31 ( .A(u4_sll_451_ML_int_3__31_), .B(
        u4_sll_451_ML_int_3__23_), .S(u4_sll_451_n16), .Z(
        u4_sll_451_ML_int_4__31_) );
  MUX2_X2 u4_sll_451_M1_3_32 ( .A(u4_sll_451_ML_int_3__32_), .B(
        u4_sll_451_ML_int_3__24_), .S(u4_sll_451_n17), .Z(
        u4_sll_451_ML_int_4__32_) );
  MUX2_X2 u4_sll_451_M1_3_33 ( .A(u4_sll_451_ML_int_3__33_), .B(
        u4_sll_451_ML_int_3__25_), .S(u4_sll_451_n17), .Z(
        u4_sll_451_ML_int_4__33_) );
  MUX2_X2 u4_sll_451_M1_3_34 ( .A(u4_sll_451_ML_int_3__34_), .B(
        u4_sll_451_ML_int_3__26_), .S(u4_sll_451_n17), .Z(
        u4_sll_451_ML_int_4__34_) );
  MUX2_X2 u4_sll_451_M1_3_35 ( .A(u4_sll_451_ML_int_3__35_), .B(
        u4_sll_451_ML_int_3__27_), .S(u4_sll_451_n17), .Z(
        u4_sll_451_ML_int_4__35_) );
  MUX2_X2 u4_sll_451_M1_3_36 ( .A(u4_sll_451_ML_int_3__36_), .B(
        u4_sll_451_ML_int_3__28_), .S(u4_sll_451_n17), .Z(
        u4_sll_451_ML_int_4__36_) );
  MUX2_X2 u4_sll_451_M1_3_37 ( .A(u4_sll_451_ML_int_3__37_), .B(
        u4_sll_451_ML_int_3__29_), .S(u4_sll_451_n17), .Z(
        u4_sll_451_ML_int_4__37_) );
  MUX2_X2 u4_sll_451_M1_3_38 ( .A(u4_sll_451_ML_int_3__38_), .B(
        u4_sll_451_ML_int_3__30_), .S(u4_sll_451_n17), .Z(
        u4_sll_451_ML_int_4__38_) );
  MUX2_X2 u4_sll_451_M1_3_39 ( .A(u4_sll_451_ML_int_3__39_), .B(
        u4_sll_451_ML_int_3__31_), .S(u4_sll_451_n17), .Z(
        u4_sll_451_ML_int_4__39_) );
  MUX2_X2 u4_sll_451_M1_3_40 ( .A(u4_sll_451_ML_int_3__40_), .B(
        u4_sll_451_ML_int_3__32_), .S(u4_sll_451_n17), .Z(
        u4_sll_451_ML_int_4__40_) );
  MUX2_X2 u4_sll_451_M1_3_41 ( .A(u4_sll_451_ML_int_3__41_), .B(
        u4_sll_451_ML_int_3__33_), .S(u4_sll_451_n17), .Z(
        u4_sll_451_ML_int_4__41_) );
  MUX2_X2 u4_sll_451_M1_3_42 ( .A(u4_sll_451_ML_int_3__42_), .B(
        u4_sll_451_ML_int_3__34_), .S(u4_sll_451_n17), .Z(
        u4_sll_451_ML_int_4__42_) );
  MUX2_X2 u4_sll_451_M1_3_43 ( .A(u4_sll_451_ML_int_3__43_), .B(
        u4_sll_451_ML_int_3__35_), .S(u4_sll_451_n17), .Z(
        u4_sll_451_ML_int_4__43_) );
  MUX2_X2 u4_sll_451_M1_3_44 ( .A(u4_sll_451_ML_int_3__44_), .B(
        u4_sll_451_ML_int_3__36_), .S(u4_sll_451_n17), .Z(
        u4_sll_451_ML_int_4__44_) );
  MUX2_X2 u4_sll_451_M1_3_45 ( .A(u4_sll_451_ML_int_3__45_), .B(
        u4_sll_451_ML_int_3__37_), .S(u4_sll_451_n17), .Z(
        u4_sll_451_ML_int_4__45_) );
  MUX2_X2 u4_sll_451_M1_3_46 ( .A(u4_sll_451_ML_int_3__46_), .B(
        u4_sll_451_ML_int_3__38_), .S(u4_sll_451_n17), .Z(
        u4_sll_451_ML_int_4__46_) );
  MUX2_X2 u4_sll_451_M1_3_47 ( .A(u4_sll_451_ML_int_3__47_), .B(
        u4_sll_451_ML_int_3__39_), .S(u4_sll_451_n17), .Z(
        u4_sll_451_ML_int_4__47_) );
  MUX2_X2 u4_sll_451_M1_4_16 ( .A(u4_sll_451_ML_int_4__16_), .B(
        u4_sll_451_ML_int_4__0_), .S(u4_sll_451_n8), .Z(
        u4_sll_451_ML_int_5__16_) );
  MUX2_X2 u4_sll_451_M1_4_17 ( .A(u4_sll_451_ML_int_4__17_), .B(
        u4_sll_451_ML_int_4__1_), .S(u4_sll_451_n8), .Z(
        u4_sll_451_ML_int_5__17_) );
  MUX2_X2 u4_sll_451_M1_4_18 ( .A(u4_sll_451_ML_int_4__18_), .B(
        u4_sll_451_ML_int_4__2_), .S(u4_sll_451_n8), .Z(
        u4_sll_451_ML_int_5__18_) );
  MUX2_X2 u4_sll_451_M1_4_19 ( .A(u4_sll_451_ML_int_4__19_), .B(
        u4_sll_451_ML_int_4__3_), .S(u4_sll_451_n8), .Z(
        u4_sll_451_ML_int_5__19_) );
  MUX2_X2 u4_sll_451_M1_4_20 ( .A(u4_sll_451_ML_int_4__20_), .B(
        u4_sll_451_ML_int_4__4_), .S(u4_sll_451_n8), .Z(
        u4_sll_451_ML_int_5__20_) );
  MUX2_X2 u4_sll_451_M1_4_21 ( .A(u4_sll_451_ML_int_4__21_), .B(
        u4_sll_451_ML_int_4__5_), .S(u4_sll_451_n8), .Z(
        u4_sll_451_ML_int_5__21_) );
  MUX2_X2 u4_sll_451_M1_4_22 ( .A(u4_sll_451_ML_int_4__22_), .B(
        u4_sll_451_ML_int_4__6_), .S(u4_sll_451_n9), .Z(
        u4_sll_451_ML_int_5__22_) );
  MUX2_X2 u4_sll_451_M1_4_23 ( .A(u4_sll_451_ML_int_4__23_), .B(
        u4_sll_451_ML_int_4__7_), .S(u4_sll_451_n9), .Z(
        u4_sll_451_ML_int_5__23_) );
  MUX2_X2 u4_sll_451_M1_4_24 ( .A(u4_sll_451_ML_int_4__24_), .B(
        u4_sll_451_ML_int_4__8_), .S(u4_sll_451_n9), .Z(
        u4_sll_451_ML_int_5__24_) );
  MUX2_X2 u4_sll_451_M1_4_25 ( .A(u4_sll_451_ML_int_4__25_), .B(
        u4_sll_451_ML_int_4__9_), .S(u4_sll_451_n9), .Z(
        u4_sll_451_ML_int_5__25_) );
  MUX2_X2 u4_sll_451_M1_4_26 ( .A(u4_sll_451_ML_int_4__26_), .B(
        u4_sll_451_ML_int_4__10_), .S(u4_sll_451_n9), .Z(
        u4_sll_451_ML_int_5__26_) );
  MUX2_X2 u4_sll_451_M1_4_27 ( .A(u4_sll_451_ML_int_4__27_), .B(
        u4_sll_451_ML_int_4__11_), .S(u4_sll_451_n9), .Z(
        u4_sll_451_ML_int_5__27_) );
  MUX2_X2 u4_sll_451_M1_4_28 ( .A(u4_sll_451_ML_int_4__28_), .B(
        u4_sll_451_ML_int_4__12_), .S(u4_sll_451_n9), .Z(
        u4_sll_451_ML_int_5__28_) );
  MUX2_X2 u4_sll_451_M1_4_29 ( .A(u4_sll_451_ML_int_4__29_), .B(
        u4_sll_451_ML_int_4__13_), .S(u4_sll_451_n9), .Z(
        u4_sll_451_ML_int_5__29_) );
  MUX2_X2 u4_sll_451_M1_4_30 ( .A(u4_sll_451_ML_int_4__30_), .B(
        u4_sll_451_ML_int_4__14_), .S(u4_sll_451_n9), .Z(
        u4_sll_451_ML_int_5__30_) );
  MUX2_X2 u4_sll_451_M1_4_31 ( .A(u4_sll_451_ML_int_4__31_), .B(
        u4_sll_451_ML_int_4__15_), .S(u4_sll_451_n9), .Z(
        u4_sll_451_ML_int_5__31_) );
  MUX2_X2 u4_sll_451_M1_4_32 ( .A(u4_sll_451_ML_int_4__32_), .B(
        u4_sll_451_ML_int_4__16_), .S(u4_sll_451_n9), .Z(
        u4_sll_451_ML_int_5__32_) );
  MUX2_X2 u4_sll_451_M1_4_33 ( .A(u4_sll_451_ML_int_4__33_), .B(
        u4_sll_451_ML_int_4__17_), .S(u4_sll_451_n9), .Z(
        u4_sll_451_ML_int_5__33_) );
  MUX2_X2 u4_sll_451_M1_4_34 ( .A(u4_sll_451_ML_int_4__34_), .B(
        u4_sll_451_ML_int_4__18_), .S(u4_sll_451_n9), .Z(
        u4_sll_451_ML_int_5__34_) );
  MUX2_X2 u4_sll_451_M1_4_35 ( .A(u4_sll_451_ML_int_4__35_), .B(
        u4_sll_451_ML_int_4__19_), .S(u4_sll_451_n9), .Z(
        u4_sll_451_ML_int_5__35_) );
  MUX2_X2 u4_sll_451_M1_4_36 ( .A(u4_sll_451_ML_int_4__36_), .B(
        u4_sll_451_ML_int_4__20_), .S(u4_sll_451_n9), .Z(
        u4_sll_451_ML_int_5__36_) );
  MUX2_X2 u4_sll_451_M1_4_37 ( .A(u4_sll_451_ML_int_4__37_), .B(
        u4_sll_451_ML_int_4__21_), .S(u4_sll_451_n9), .Z(
        u4_sll_451_ML_int_5__37_) );
  MUX2_X2 u4_sll_451_M1_4_38 ( .A(u4_sll_451_ML_int_4__38_), .B(
        u4_sll_451_ML_int_4__22_), .S(u4_sll_451_n9), .Z(
        u4_sll_451_ML_int_5__38_) );
  MUX2_X2 u4_sll_451_M1_4_39 ( .A(u4_sll_451_ML_int_4__39_), .B(
        u4_sll_451_ML_int_4__23_), .S(u4_sll_451_n9), .Z(
        u4_sll_451_ML_int_5__39_) );
  MUX2_X2 u4_sll_451_M1_4_40 ( .A(u4_sll_451_ML_int_4__40_), .B(
        u4_sll_451_ML_int_4__24_), .S(u4_sll_451_n10), .Z(
        u4_sll_451_ML_int_5__40_) );
  MUX2_X2 u4_sll_451_M1_4_41 ( .A(u4_sll_451_ML_int_4__41_), .B(
        u4_sll_451_ML_int_4__25_), .S(u4_sll_451_n10), .Z(
        u4_sll_451_ML_int_5__41_) );
  MUX2_X2 u4_sll_451_M1_4_42 ( .A(u4_sll_451_ML_int_4__42_), .B(
        u4_sll_451_ML_int_4__26_), .S(u4_sll_451_n10), .Z(
        u4_sll_451_ML_int_5__42_) );
  MUX2_X2 u4_sll_451_M1_4_43 ( .A(u4_sll_451_ML_int_4__43_), .B(
        u4_sll_451_ML_int_4__27_), .S(u4_sll_451_n10), .Z(
        u4_sll_451_ML_int_5__43_) );
  MUX2_X2 u4_sll_451_M1_4_44 ( .A(u4_sll_451_ML_int_4__44_), .B(
        u4_sll_451_ML_int_4__28_), .S(u4_sll_451_n10), .Z(
        u4_sll_451_ML_int_5__44_) );
  MUX2_X2 u4_sll_451_M1_4_45 ( .A(u4_sll_451_ML_int_4__45_), .B(
        u4_sll_451_ML_int_4__29_), .S(u4_sll_451_n10), .Z(
        u4_sll_451_ML_int_5__45_) );
  MUX2_X2 u4_sll_451_M1_4_46 ( .A(u4_sll_451_ML_int_4__46_), .B(
        u4_sll_451_ML_int_4__30_), .S(u4_sll_451_n10), .Z(
        u4_sll_451_ML_int_5__46_) );
  MUX2_X2 u4_sll_451_M1_4_47 ( .A(u4_sll_451_ML_int_4__47_), .B(
        u4_sll_451_ML_int_4__31_), .S(u4_sll_451_n10), .Z(
        u4_sll_451_ML_int_5__47_) );
  MUX2_X2 u4_sll_451_M1_5_32 ( .A(u4_sll_451_ML_int_5__32_), .B(
        u4_sll_451_ML_int_5__0_), .S(u4_sll_451_n2), .Z(u4_N1440) );
  MUX2_X2 u4_sll_451_M1_5_33 ( .A(u4_sll_451_ML_int_5__33_), .B(
        u4_sll_451_ML_int_5__1_), .S(u4_sll_451_n2), .Z(u4_N1441) );
  MUX2_X2 u4_sll_451_M1_5_34 ( .A(u4_sll_451_ML_int_5__34_), .B(
        u4_sll_451_ML_int_5__2_), .S(u4_sll_451_n2), .Z(u4_N1442) );
  MUX2_X2 u4_sll_451_M1_5_35 ( .A(u4_sll_451_ML_int_5__35_), .B(
        u4_sll_451_ML_int_5__3_), .S(u4_sll_451_n2), .Z(u4_N1443) );
  MUX2_X2 u4_sll_451_M1_5_36 ( .A(u4_sll_451_ML_int_5__36_), .B(
        u4_sll_451_ML_int_5__4_), .S(u4_sll_451_n2), .Z(u4_N1444) );
  MUX2_X2 u4_sll_451_M1_5_37 ( .A(u4_sll_451_ML_int_5__37_), .B(
        u4_sll_451_ML_int_5__5_), .S(u4_sll_451_n2), .Z(u4_N1445) );
  MUX2_X2 u4_sll_451_M1_5_38 ( .A(u4_sll_451_ML_int_5__38_), .B(
        u4_sll_451_ML_int_5__6_), .S(u4_sll_451_n2), .Z(u4_N1446) );
  MUX2_X2 u4_sll_451_M1_5_39 ( .A(u4_sll_451_ML_int_5__39_), .B(
        u4_sll_451_ML_int_5__7_), .S(u4_sll_451_n2), .Z(u4_N1447) );
  MUX2_X2 u4_sll_451_M1_5_40 ( .A(u4_sll_451_ML_int_5__40_), .B(
        u4_sll_451_ML_int_5__8_), .S(u4_sll_451_n2), .Z(u4_N1448) );
  MUX2_X2 u4_sll_451_M1_5_41 ( .A(u4_sll_451_ML_int_5__41_), .B(
        u4_sll_451_ML_int_5__9_), .S(u4_sll_451_n2), .Z(u4_N1449) );
  MUX2_X2 u4_sll_451_M1_5_42 ( .A(u4_sll_451_ML_int_5__42_), .B(
        u4_sll_451_ML_int_5__10_), .S(u4_sll_451_n2), .Z(u4_N1450) );
  MUX2_X2 u4_sll_451_M1_5_43 ( .A(u4_sll_451_ML_int_5__43_), .B(
        u4_sll_451_ML_int_5__11_), .S(u4_sll_451_n2), .Z(u4_N1451) );
  MUX2_X2 u4_sll_451_M1_5_44 ( .A(u4_sll_451_ML_int_5__44_), .B(
        u4_sll_451_ML_int_5__12_), .S(u4_sll_451_n2), .Z(u4_N1452) );
  MUX2_X2 u4_sll_451_M1_5_45 ( .A(u4_sll_451_ML_int_5__45_), .B(
        u4_sll_451_ML_int_5__13_), .S(u4_sll_451_n2), .Z(u4_N1453) );
  MUX2_X2 u4_sll_451_M1_5_46 ( .A(u4_sll_451_ML_int_5__46_), .B(
        u4_sll_451_ML_int_5__14_), .S(u4_sll_451_n2), .Z(u4_N1454) );
  MUX2_X2 u4_sll_451_M1_5_47 ( .A(u4_sll_451_ML_int_5__47_), .B(
        u4_sll_451_ML_int_5__15_), .S(u4_sll_451_n2), .Z(u4_N1455) );
  INV_X1 u4_srl_450_U355 ( .A(u4_shift_right[2]), .ZN(u4_srl_450_n302) );
  INV_X1 u4_srl_450_U354 ( .A(u4_shift_right[3]), .ZN(u4_srl_450_n255) );
  NAND2_X1 u4_srl_450_U353 ( .A1(u4_srl_450_n302), .A2(u4_srl_450_n255), .ZN(
        u4_srl_450_n275) );
  NOR2_X1 u4_srl_450_U352 ( .A1(u4_srl_450_n275), .A2(u4_shift_right[4]), .ZN(
        u4_srl_450_n130) );
  NAND2_X1 u4_srl_450_U351 ( .A1(u4_shift_right[1]), .A2(u4_shift_right[0]), 
        .ZN(u4_srl_450_n139) );
  INV_X1 u4_srl_450_U350 ( .A(u4_shift_right[0]), .ZN(u4_srl_450_n305) );
  NAND2_X1 u4_srl_450_U349 ( .A1(u4_shift_right[1]), .A2(u4_srl_450_n305), 
        .ZN(u4_srl_450_n140) );
  NOR2_X1 u4_srl_450_U348 ( .A1(u4_srl_450_n305), .A2(u4_shift_right[1]), .ZN(
        u4_srl_450_n142) );
  NOR2_X1 u4_srl_450_U347 ( .A1(u4_shift_right[0]), .A2(u4_shift_right[1]), 
        .ZN(u4_srl_450_n143) );
  AOI22_X1 u4_srl_450_U346 ( .A1(n3521), .A2(u4_srl_450_n12), .B1(n3564), .B2(
        u4_srl_450_n143), .ZN(u4_srl_450_n304) );
  OAI221_X1 u4_srl_450_U345 ( .B1(u4_srl_450_n4), .B2(u4_srl_450_n64), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n20), .A(u4_srl_450_n304), .ZN(
        u4_srl_450_n290) );
  AOI22_X1 u4_srl_450_U344 ( .A1(n3528), .A2(u4_srl_450_n12), .B1(n3526), .B2(
        u4_srl_450_n16), .ZN(u4_srl_450_n303) );
  OAI221_X1 u4_srl_450_U343 ( .B1(u4_srl_450_n4), .B2(u4_srl_450_n62), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n25), .A(u4_srl_450_n303), .ZN(
        u4_srl_450_n87) );
  AOI22_X1 u4_srl_450_U342 ( .A1(n3530), .A2(u4_srl_450_n12), .B1(n3529), .B2(
        u4_srl_450_n16), .ZN(u4_srl_450_n301) );
  OAI221_X1 u4_srl_450_U341 ( .B1(u4_srl_450_n4), .B2(u4_srl_450_n29), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n61), .A(u4_srl_450_n301), .ZN(
        u4_srl_450_n83) );
  AOI22_X1 u4_srl_450_U340 ( .A1(n3524), .A2(u4_srl_450_n12), .B1(n3523), .B2(
        u4_srl_450_n16), .ZN(u4_srl_450_n300) );
  OAI221_X1 u4_srl_450_U339 ( .B1(u4_srl_450_n4), .B2(u4_srl_450_n23), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n63), .A(u4_srl_450_n300), .ZN(
        u4_srl_450_n117) );
  NAND2_X1 u4_srl_450_U338 ( .A1(u4_shift_right[2]), .A2(u4_srl_450_n255), 
        .ZN(u4_srl_450_n272) );
  INV_X1 u4_srl_450_U337 ( .A(u4_srl_450_n272), .ZN(u4_srl_450_n138) );
  AOI222_X1 u4_srl_450_U336 ( .A1(u4_srl_450_n87), .A2(u4_srl_450_n136), .B1(
        u4_srl_450_n83), .B2(u4_srl_450_n137), .C1(u4_srl_450_n117), .C2(
        u4_srl_450_n3), .ZN(u4_srl_450_n293) );
  AOI22_X1 u4_srl_450_U335 ( .A1(fract_denorm[29]), .A2(u4_srl_450_n12), .B1(
        fract_denorm[28]), .B2(u4_srl_450_n16), .ZN(u4_srl_450_n299) );
  OAI221_X1 u4_srl_450_U334 ( .B1(u4_srl_450_n4), .B2(u4_srl_450_n50), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n40), .A(u4_srl_450_n299), .ZN(
        u4_srl_450_n174) );
  AOI22_X1 u4_srl_450_U333 ( .A1(fract_denorm[25]), .A2(u4_srl_450_n12), .B1(
        u4_srl_450_n14), .B2(fract_denorm[24]), .ZN(u4_srl_450_n298) );
  OAI221_X1 u4_srl_450_U332 ( .B1(u4_srl_450_n4), .B2(u4_srl_450_n38), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n37), .A(u4_srl_450_n298), .ZN(
        u4_srl_450_n175) );
  AOI22_X1 u4_srl_450_U331 ( .A1(fract_denorm[21]), .A2(u4_srl_450_n12), .B1(
        n3557), .B2(u4_srl_450_n16), .ZN(u4_srl_450_n297) );
  OAI221_X1 u4_srl_450_U330 ( .B1(u4_srl_450_n4), .B2(u4_srl_450_n42), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n34), .A(u4_srl_450_n297), .ZN(
        u4_srl_450_n84) );
  AOI22_X1 u4_srl_450_U329 ( .A1(n3559), .A2(u4_srl_450_n12), .B1(n3532), .B2(
        u4_srl_450_n16), .ZN(u4_srl_450_n296) );
  OAI221_X1 u4_srl_450_U328 ( .B1(u4_srl_450_n4), .B2(u4_srl_450_n32), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n31), .A(u4_srl_450_n296), .ZN(
        u4_srl_450_n85) );
  AOI22_X1 u4_srl_450_U327 ( .A1(u4_srl_450_n3), .A2(u4_srl_450_n84), .B1(
        u4_srl_450_n17), .B2(u4_srl_450_n85), .ZN(u4_srl_450_n295) );
  INV_X1 u4_srl_450_U326 ( .A(u4_srl_450_n295), .ZN(u4_srl_450_n294) );
  AOI221_X1 u4_srl_450_U325 ( .B1(u4_srl_450_n174), .B2(u4_srl_450_n137), .C1(
        u4_srl_450_n175), .C2(u4_srl_450_n136), .A(u4_srl_450_n294), .ZN(
        u4_srl_450_n226) );
  MUX2_X1 u4_srl_450_U324 ( .A(u4_srl_450_n293), .B(u4_srl_450_n226), .S(
        u4_shift_right[4]), .Z(u4_srl_450_n292) );
  INV_X1 u4_srl_450_U323 ( .A(u4_srl_450_n292), .ZN(u4_srl_450_n291) );
  AOI21_X1 u4_srl_450_U322 ( .B1(u4_srl_450_n130), .B2(u4_srl_450_n290), .A(
        u4_srl_450_n291), .ZN(u4_srl_450_n284) );
  AOI22_X1 u4_srl_450_U321 ( .A1(fract_denorm[37]), .A2(u4_srl_450_n12), .B1(
        fract_denorm[36]), .B2(u4_srl_450_n16), .ZN(u4_srl_450_n289) );
  OAI221_X1 u4_srl_450_U320 ( .B1(u4_srl_450_n4), .B2(u4_srl_450_n51), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n48), .A(u4_srl_450_n289), .ZN(
        u4_srl_450_n202) );
  AOI22_X1 u4_srl_450_U319 ( .A1(fract_denorm[33]), .A2(u4_srl_450_n12), .B1(
        fract_denorm[32]), .B2(u4_srl_450_n16), .ZN(u4_srl_450_n288) );
  OAI221_X1 u4_srl_450_U318 ( .B1(u4_srl_450_n4), .B2(u4_srl_450_n46), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n45), .A(u4_srl_450_n288), .ZN(
        u4_srl_450_n179) );
  AOI22_X1 u4_srl_450_U317 ( .A1(fract_denorm[45]), .A2(u4_srl_450_n12), .B1(
        fract_denorm[44]), .B2(u4_srl_450_n16), .ZN(u4_srl_450_n287) );
  OAI221_X1 u4_srl_450_U316 ( .B1(u4_srl_450_n4), .B2(u4_srl_450_n19), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n55), .A(u4_srl_450_n287), .ZN(
        u4_srl_450_n173) );
  INV_X1 u4_srl_450_U315 ( .A(u4_srl_450_n173), .ZN(u4_srl_450_n123) );
  AOI22_X1 u4_srl_450_U314 ( .A1(fract_denorm[41]), .A2(u4_srl_450_n12), .B1(
        fract_denorm[40]), .B2(u4_srl_450_n16), .ZN(u4_srl_450_n286) );
  OAI221_X1 u4_srl_450_U313 ( .B1(u4_srl_450_n6), .B2(u4_srl_450_n56), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n58), .A(u4_srl_450_n286), .ZN(
        u4_srl_450_n172) );
  INV_X1 u4_srl_450_U312 ( .A(u4_srl_450_n172), .ZN(u4_srl_450_n250) );
  OAI22_X1 u4_srl_450_U311 ( .A1(u4_srl_450_n168), .A2(u4_srl_450_n123), .B1(
        u4_srl_450_n170), .B2(u4_srl_450_n250), .ZN(u4_srl_450_n285) );
  AOI221_X1 u4_srl_450_U310 ( .B1(u4_srl_450_n202), .B2(u4_srl_450_n3), .C1(
        u4_srl_450_n179), .C2(u4_srl_450_n17), .A(u4_srl_450_n285), .ZN(
        u4_srl_450_n147) );
  INV_X1 u4_srl_450_U309 ( .A(u4_shift_right[4]), .ZN(u4_srl_450_n276) );
  NAND2_X1 u4_srl_450_U308 ( .A1(u4_shift_right[5]), .A2(u4_srl_450_n276), 
        .ZN(u4_srl_450_n129) );
  OAI22_X1 u4_srl_450_U307 ( .A1(u4_shift_right[5]), .A2(u4_srl_450_n284), 
        .B1(u4_srl_450_n147), .B2(u4_srl_450_n129), .ZN(u4_N1358) );
  AOI22_X1 u4_srl_450_U306 ( .A1(fract_denorm[31]), .A2(u4_srl_450_n12), .B1(
        fract_denorm[30]), .B2(u4_srl_450_n16), .ZN(u4_srl_450_n283) );
  OAI221_X1 u4_srl_450_U305 ( .B1(u4_srl_450_n6), .B2(u4_srl_450_n44), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n43), .A(u4_srl_450_n283), .ZN(
        u4_srl_450_n197) );
  AOI22_X1 u4_srl_450_U304 ( .A1(fract_denorm[27]), .A2(u4_srl_450_n12), .B1(
        fract_denorm[26]), .B2(u4_srl_450_n143), .ZN(u4_srl_450_n282) );
  OAI221_X1 u4_srl_450_U303 ( .B1(u4_srl_450_n4), .B2(u4_srl_450_n39), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n41), .A(u4_srl_450_n282), .ZN(
        u4_srl_450_n192) );
  AOI22_X1 u4_srl_450_U302 ( .A1(fract_denorm[39]), .A2(u4_srl_450_n12), .B1(
        fract_denorm[38]), .B2(u4_srl_450_n16), .ZN(u4_srl_450_n281) );
  OAI221_X1 u4_srl_450_U301 ( .B1(u4_srl_450_n4), .B2(u4_srl_450_n53), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n52), .A(u4_srl_450_n281), .ZN(
        u4_srl_450_n191) );
  INV_X1 u4_srl_450_U300 ( .A(u4_srl_450_n191), .ZN(u4_srl_450_n235) );
  AOI22_X1 u4_srl_450_U299 ( .A1(fract_denorm[35]), .A2(u4_srl_450_n12), .B1(
        fract_denorm[34]), .B2(u4_srl_450_n16), .ZN(u4_srl_450_n280) );
  OAI221_X1 u4_srl_450_U298 ( .B1(u4_srl_450_n6), .B2(u4_srl_450_n47), .C1(
        u4_srl_450_n10), .C2(u4_srl_450_n49), .A(u4_srl_450_n280), .ZN(
        u4_srl_450_n217) );
  INV_X1 u4_srl_450_U297 ( .A(u4_srl_450_n217), .ZN(u4_srl_450_n195) );
  OAI22_X1 u4_srl_450_U296 ( .A1(u4_srl_450_n168), .A2(u4_srl_450_n235), .B1(
        u4_srl_450_n170), .B2(u4_srl_450_n195), .ZN(u4_srl_450_n279) );
  AOI221_X1 u4_srl_450_U295 ( .B1(u4_srl_450_n197), .B2(u4_srl_450_n138), .C1(
        u4_srl_450_n192), .C2(u4_srl_450_n18), .A(u4_srl_450_n279), .ZN(
        u4_srl_450_n162) );
  INV_X1 u4_srl_450_U294 ( .A(u4_shift_right[5]), .ZN(u4_srl_450_n277) );
  NAND2_X1 u4_srl_450_U293 ( .A1(u4_shift_right[4]), .A2(u4_srl_450_n277), 
        .ZN(u4_srl_450_n66) );
  INV_X1 u4_srl_450_U292 ( .A(u4_srl_450_n129), .ZN(u4_srl_450_n75) );
  AOI22_X1 u4_srl_450_U291 ( .A1(fract_denorm[43]), .A2(u4_srl_450_n12), .B1(
        fract_denorm[42]), .B2(u4_srl_450_n16), .ZN(u4_srl_450_n278) );
  OAI221_X1 u4_srl_450_U290 ( .B1(u4_srl_450_n6), .B2(u4_srl_450_n54), .C1(
        u4_srl_450_n140), .C2(u4_srl_450_n57), .A(u4_srl_450_n278), .ZN(
        u4_srl_450_n189) );
  AOI22_X1 u4_srl_450_U289 ( .A1(u4_srl_450_n16), .A2(fract_denorm[46]), .B1(
        u4_srl_450_n12), .B2(n2679), .ZN(u4_srl_450_n121) );
  INV_X1 u4_srl_450_U288 ( .A(u4_srl_450_n121), .ZN(u4_srl_450_n190) );
  AOI22_X1 u4_srl_450_U287 ( .A1(u4_srl_450_n189), .A2(u4_srl_450_n17), .B1(
        u4_srl_450_n190), .B2(u4_srl_450_n3), .ZN(u4_srl_450_n126) );
  INV_X1 u4_srl_450_U286 ( .A(u4_srl_450_n126), .ZN(u4_srl_450_n273) );
  AOI22_X1 u4_srl_450_U285 ( .A1(n3561), .A2(u4_srl_450_n12), .B1(n3527), .B2(
        u4_srl_450_n143), .ZN(u4_srl_450_n274) );
  OAI221_X1 u4_srl_450_U284 ( .B1(u4_srl_450_n6), .B2(u4_srl_450_n28), .C1(
        u4_srl_450_n140), .C2(u4_srl_450_n27), .A(u4_srl_450_n274), .ZN(
        u4_srl_450_n101) );
  AOI22_X1 u4_srl_450_U283 ( .A1(u4_srl_450_n75), .A2(u4_srl_450_n273), .B1(
        u4_srl_450_n77), .B2(u4_srl_450_n101), .ZN(u4_srl_450_n267) );
  AOI22_X1 u4_srl_450_U282 ( .A1(n3531), .A2(u4_srl_450_n12), .B1(n3560), .B2(
        u4_srl_450_n14), .ZN(u4_srl_450_n271) );
  OAI221_X1 u4_srl_450_U281 ( .B1(u4_srl_450_n6), .B2(u4_srl_450_n60), .C1(
        u4_srl_450_n140), .C2(u4_srl_450_n30), .A(u4_srl_450_n271), .ZN(
        u4_srl_450_n103) );
  AOI22_X1 u4_srl_450_U280 ( .A1(u4_srl_450_n12), .A2(fract_denorm[23]), .B1(
        u4_srl_450_n143), .B2(fract_denorm[22]), .ZN(u4_srl_450_n270) );
  OAI221_X1 u4_srl_450_U279 ( .B1(u4_srl_450_n4), .B2(u4_srl_450_n36), .C1(
        u4_srl_450_n35), .C2(u4_srl_450_n8), .A(u4_srl_450_n270), .ZN(
        u4_srl_450_n193) );
  AOI22_X1 u4_srl_450_U278 ( .A1(n3534), .A2(u4_srl_450_n12), .B1(n3533), .B2(
        u4_srl_450_n143), .ZN(u4_srl_450_n269) );
  OAI221_X1 u4_srl_450_U277 ( .B1(u4_srl_450_n6), .B2(u4_srl_450_n33), .C1(
        u4_srl_450_n140), .C2(u4_srl_450_n59), .A(u4_srl_450_n269), .ZN(
        u4_srl_450_n102) );
  AOI222_X1 u4_srl_450_U276 ( .A1(u4_srl_450_n69), .A2(u4_srl_450_n103), .B1(
        u4_srl_450_n71), .B2(u4_srl_450_n193), .C1(u4_srl_450_n73), .C2(
        u4_srl_450_n102), .ZN(u4_srl_450_n268) );
  OAI211_X1 u4_srl_450_U275 ( .C1(u4_srl_450_n162), .C2(u4_srl_450_n2), .A(
        u4_srl_450_n267), .B(u4_srl_450_n268), .ZN(u4_N1368) );
  AOI22_X1 u4_srl_450_U274 ( .A1(fract_denorm[32]), .A2(u4_srl_450_n12), .B1(
        fract_denorm[31]), .B2(u4_srl_450_n16), .ZN(u4_srl_450_n266) );
  OAI221_X1 u4_srl_450_U273 ( .B1(u4_srl_450_n6), .B2(u4_srl_450_n45), .C1(
        u4_srl_450_n140), .C2(u4_srl_450_n44), .A(u4_srl_450_n266), .ZN(
        u4_srl_450_n188) );
  AOI22_X1 u4_srl_450_U272 ( .A1(fract_denorm[28]), .A2(u4_srl_450_n12), .B1(
        fract_denorm[27]), .B2(u4_srl_450_n143), .ZN(u4_srl_450_n265) );
  OAI221_X1 u4_srl_450_U271 ( .B1(u4_srl_450_n5), .B2(u4_srl_450_n40), .C1(
        u4_srl_450_n140), .C2(u4_srl_450_n39), .A(u4_srl_450_n265), .ZN(
        u4_srl_450_n183) );
  AOI22_X1 u4_srl_450_U270 ( .A1(fract_denorm[40]), .A2(u4_srl_450_n12), .B1(
        fract_denorm[39]), .B2(u4_srl_450_n16), .ZN(u4_srl_450_n264) );
  OAI221_X1 u4_srl_450_U269 ( .B1(u4_srl_450_n5), .B2(u4_srl_450_n58), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n53), .A(u4_srl_450_n264), .ZN(
        u4_srl_450_n182) );
  AOI22_X1 u4_srl_450_U268 ( .A1(fract_denorm[36]), .A2(u4_srl_450_n142), .B1(
        fract_denorm[35]), .B2(u4_srl_450_n143), .ZN(u4_srl_450_n263) );
  OAI221_X1 u4_srl_450_U267 ( .B1(u4_srl_450_n5), .B2(u4_srl_450_n48), .C1(
        u4_srl_450_n140), .C2(u4_srl_450_n47), .A(u4_srl_450_n263), .ZN(
        u4_srl_450_n187) );
  AOI22_X1 u4_srl_450_U266 ( .A1(u4_srl_450_n137), .A2(u4_srl_450_n182), .B1(
        u4_srl_450_n136), .B2(u4_srl_450_n187), .ZN(u4_srl_450_n262) );
  INV_X1 u4_srl_450_U265 ( .A(u4_srl_450_n262), .ZN(u4_srl_450_n261) );
  AOI221_X1 u4_srl_450_U264 ( .B1(u4_srl_450_n188), .B2(u4_srl_450_n3), .C1(
        u4_srl_450_n183), .C2(u4_srl_450_n17), .A(u4_srl_450_n261), .ZN(
        u4_srl_450_n161) );
  INV_X1 u4_srl_450_U263 ( .A(u4_srl_450_n161), .ZN(u4_srl_450_n258) );
  AOI22_X1 u4_srl_450_U262 ( .A1(n3532), .A2(u4_srl_450_n12), .B1(n3531), .B2(
        u4_srl_450_n14), .ZN(u4_srl_450_n260) );
  OAI221_X1 u4_srl_450_U261 ( .B1(u4_srl_450_n5), .B2(u4_srl_450_n31), .C1(
        u4_srl_450_n140), .C2(u4_srl_450_n60), .A(u4_srl_450_n260), .ZN(
        u4_srl_450_n94) );
  AOI22_X1 u4_srl_450_U260 ( .A1(n3529), .A2(u4_srl_450_n142), .B1(n3561), 
        .B2(u4_srl_450_n14), .ZN(u4_srl_450_n259) );
  OAI221_X1 u4_srl_450_U259 ( .B1(u4_srl_450_n5), .B2(u4_srl_450_n61), .C1(
        u4_srl_450_n140), .C2(u4_srl_450_n28), .A(u4_srl_450_n259), .ZN(
        u4_srl_450_n92) );
  AOI222_X1 u4_srl_450_U258 ( .A1(u4_srl_450_n1), .A2(u4_srl_450_n258), .B1(
        u4_srl_450_n69), .B2(u4_srl_450_n94), .C1(u4_srl_450_n77), .C2(
        u4_srl_450_n92), .ZN(u4_srl_450_n251) );
  AOI22_X1 u4_srl_450_U257 ( .A1(n3557), .A2(u4_srl_450_n142), .B1(n3534), 
        .B2(u4_srl_450_n14), .ZN(u4_srl_450_n257) );
  OAI221_X1 u4_srl_450_U256 ( .B1(u4_srl_450_n5), .B2(u4_srl_450_n34), .C1(
        u4_srl_450_n140), .C2(u4_srl_450_n33), .A(u4_srl_450_n257), .ZN(
        u4_srl_450_n93) );
  AOI22_X1 u4_srl_450_U255 ( .A1(fract_denorm[44]), .A2(u4_srl_450_n142), .B1(
        fract_denorm[43]), .B2(u4_srl_450_n14), .ZN(u4_srl_450_n256) );
  OAI221_X1 u4_srl_450_U254 ( .B1(u4_srl_450_n5), .B2(u4_srl_450_n55), .C1(
        u4_srl_450_n140), .C2(u4_srl_450_n54), .A(u4_srl_450_n256), .ZN(
        u4_srl_450_n180) );
  NAND2_X1 u4_srl_450_U253 ( .A1(n2679), .A2(u4_srl_450_n16), .ZN(
        u4_srl_450_n120) );
  INV_X1 u4_srl_450_U252 ( .A(u4_srl_450_n120), .ZN(u4_srl_450_n181) );
  MUX2_X1 u4_srl_450_U251 ( .A(u4_srl_450_n180), .B(u4_srl_450_n181), .S(
        u4_shift_right[2]), .Z(u4_srl_450_n214) );
  NAND2_X1 u4_srl_450_U250 ( .A1(u4_srl_450_n214), .A2(u4_srl_450_n255), .ZN(
        u4_srl_450_n125) );
  INV_X1 u4_srl_450_U249 ( .A(u4_srl_450_n125), .ZN(u4_srl_450_n253) );
  AOI22_X1 u4_srl_450_U248 ( .A1(u4_srl_450_n12), .A2(fract_denorm[24]), .B1(
        u4_srl_450_n143), .B2(fract_denorm[23]), .ZN(u4_srl_450_n254) );
  OAI221_X1 u4_srl_450_U247 ( .B1(u4_srl_450_n5), .B2(u4_srl_450_n37), .C1(
        u4_srl_450_n140), .C2(u4_srl_450_n36), .A(u4_srl_450_n254), .ZN(
        u4_srl_450_n184) );
  AOI222_X1 u4_srl_450_U246 ( .A1(u4_srl_450_n73), .A2(u4_srl_450_n93), .B1(
        u4_srl_450_n253), .B2(u4_srl_450_n75), .C1(u4_srl_450_n71), .C2(
        u4_srl_450_n184), .ZN(u4_srl_450_n252) );
  NAND2_X1 u4_srl_450_U245 ( .A1(u4_srl_450_n251), .A2(u4_srl_450_n252), .ZN(
        u4_N1369) );
  INV_X1 u4_srl_450_U244 ( .A(u4_srl_450_n202), .ZN(u4_srl_450_n177) );
  OAI22_X1 u4_srl_450_U243 ( .A1(u4_srl_450_n168), .A2(u4_srl_450_n250), .B1(
        u4_srl_450_n170), .B2(u4_srl_450_n177), .ZN(u4_srl_450_n249) );
  AOI221_X1 u4_srl_450_U242 ( .B1(u4_srl_450_n179), .B2(u4_srl_450_n3), .C1(
        u4_srl_450_n174), .C2(u4_srl_450_n17), .A(u4_srl_450_n249), .ZN(
        u4_srl_450_n160) );
  AOI22_X1 u4_srl_450_U241 ( .A1(u4_srl_450_n69), .A2(u4_srl_450_n85), .B1(
        u4_srl_450_n77), .B2(u4_srl_450_n83), .ZN(u4_srl_450_n247) );
  AND2_X1 u4_srl_450_U240 ( .A1(u4_srl_450_n130), .A2(u4_shift_right[5]), .ZN(
        u4_srl_450_n229) );
  AOI222_X1 u4_srl_450_U239 ( .A1(u4_srl_450_n73), .A2(u4_srl_450_n84), .B1(
        u4_srl_450_n229), .B2(u4_srl_450_n173), .C1(u4_srl_450_n71), .C2(
        u4_srl_450_n175), .ZN(u4_srl_450_n248) );
  OAI211_X1 u4_srl_450_U238 ( .C1(u4_srl_450_n160), .C2(u4_srl_450_n2), .A(
        u4_srl_450_n247), .B(u4_srl_450_n248), .ZN(u4_N1370) );
  AOI22_X1 u4_srl_450_U237 ( .A1(fract_denorm[34]), .A2(u4_srl_450_n142), .B1(
        fract_denorm[33]), .B2(u4_srl_450_n14), .ZN(u4_srl_450_n246) );
  OAI221_X1 u4_srl_450_U236 ( .B1(u4_srl_450_n5), .B2(u4_srl_450_n49), .C1(
        u4_srl_450_n10), .C2(u4_srl_450_n46), .A(u4_srl_450_n246), .ZN(
        u4_srl_450_n201) );
  AOI22_X1 u4_srl_450_U235 ( .A1(fract_denorm[30]), .A2(u4_srl_450_n12), .B1(
        fract_denorm[29]), .B2(u4_srl_450_n14), .ZN(u4_srl_450_n245) );
  OAI221_X1 u4_srl_450_U234 ( .B1(u4_srl_450_n5), .B2(u4_srl_450_n43), .C1(
        u4_srl_450_n140), .C2(u4_srl_450_n50), .A(u4_srl_450_n245), .ZN(
        u4_srl_450_n165) );
  AOI22_X1 u4_srl_450_U233 ( .A1(fract_denorm[42]), .A2(u4_srl_450_n12), .B1(
        fract_denorm[41]), .B2(u4_srl_450_n14), .ZN(u4_srl_450_n244) );
  OAI221_X1 u4_srl_450_U232 ( .B1(u4_srl_450_n5), .B2(u4_srl_450_n57), .C1(
        u4_srl_450_n140), .C2(u4_srl_450_n56), .A(u4_srl_450_n244), .ZN(
        u4_srl_450_n163) );
  INV_X1 u4_srl_450_U231 ( .A(u4_srl_450_n163), .ZN(u4_srl_450_n223) );
  AOI22_X1 u4_srl_450_U230 ( .A1(fract_denorm[38]), .A2(u4_srl_450_n12), .B1(
        fract_denorm[37]), .B2(u4_srl_450_n14), .ZN(u4_srl_450_n243) );
  OAI221_X1 u4_srl_450_U229 ( .B1(u4_srl_450_n6), .B2(u4_srl_450_n52), .C1(
        u4_srl_450_n10), .C2(u4_srl_450_n51), .A(u4_srl_450_n243), .ZN(
        u4_srl_450_n198) );
  INV_X1 u4_srl_450_U228 ( .A(u4_srl_450_n198), .ZN(u4_srl_450_n169) );
  OAI22_X1 u4_srl_450_U227 ( .A1(u4_srl_450_n168), .A2(u4_srl_450_n223), .B1(
        u4_srl_450_n170), .B2(u4_srl_450_n169), .ZN(u4_srl_450_n242) );
  AOI221_X1 u4_srl_450_U226 ( .B1(u4_srl_450_n201), .B2(u4_srl_450_n3), .C1(
        u4_srl_450_n165), .C2(u4_srl_450_n18), .A(u4_srl_450_n242), .ZN(
        u4_srl_450_n159) );
  AOI22_X1 u4_srl_450_U225 ( .A1(n3533), .A2(u4_srl_450_n142), .B1(n3559), 
        .B2(u4_srl_450_n14), .ZN(u4_srl_450_n241) );
  OAI221_X1 u4_srl_450_U224 ( .B1(u4_srl_450_n6), .B2(u4_srl_450_n59), .C1(
        u4_srl_450_n140), .C2(u4_srl_450_n32), .A(u4_srl_450_n241), .ZN(
        u4_srl_450_n74) );
  AOI22_X1 u4_srl_450_U223 ( .A1(n3560), .A2(u4_srl_450_n142), .B1(n3530), 
        .B2(u4_srl_450_n14), .ZN(u4_srl_450_n240) );
  OAI221_X1 u4_srl_450_U222 ( .B1(u4_srl_450_n6), .B2(u4_srl_450_n30), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n29), .A(u4_srl_450_n240), .ZN(
        u4_srl_450_n70) );
  AOI22_X1 u4_srl_450_U221 ( .A1(u4_srl_450_n69), .A2(u4_srl_450_n74), .B1(
        u4_srl_450_n77), .B2(u4_srl_450_n70), .ZN(u4_srl_450_n236) );
  AOI22_X1 u4_srl_450_U220 ( .A1(fract_denorm[22]), .A2(u4_srl_450_n142), .B1(
        fract_denorm[21]), .B2(u4_srl_450_n14), .ZN(u4_srl_450_n239) );
  OAI221_X1 u4_srl_450_U219 ( .B1(u4_srl_450_n6), .B2(u4_srl_450_n35), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n42), .A(u4_srl_450_n239), .ZN(
        u4_srl_450_n72) );
  AOI222_X1 u4_srl_450_U218 ( .A1(u4_srl_450_n12), .A2(fract_denorm[46]), .B1(
        u4_srl_450_n9), .B2(n2679), .C1(u4_srl_450_n14), .C2(fract_denorm[45]), 
        .ZN(u4_srl_450_n122) );
  INV_X1 u4_srl_450_U217 ( .A(u4_srl_450_n122), .ZN(u4_srl_450_n164) );
  AOI22_X1 u4_srl_450_U216 ( .A1(fract_denorm[26]), .A2(u4_srl_450_n12), .B1(
        fract_denorm[25]), .B2(u4_srl_450_n14), .ZN(u4_srl_450_n238) );
  OAI221_X1 u4_srl_450_U215 ( .B1(u4_srl_450_n6), .B2(u4_srl_450_n41), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n38), .A(u4_srl_450_n238), .ZN(
        u4_srl_450_n166) );
  AOI222_X1 u4_srl_450_U214 ( .A1(u4_srl_450_n73), .A2(u4_srl_450_n72), .B1(
        u4_srl_450_n229), .B2(u4_srl_450_n164), .C1(u4_srl_450_n71), .C2(
        u4_srl_450_n166), .ZN(u4_srl_450_n237) );
  OAI211_X1 u4_srl_450_U213 ( .C1(u4_srl_450_n159), .C2(u4_srl_450_n2), .A(
        u4_srl_450_n236), .B(u4_srl_450_n237), .ZN(u4_N1371) );
  INV_X1 u4_srl_450_U212 ( .A(u4_srl_450_n189), .ZN(u4_srl_450_n219) );
  OAI22_X1 u4_srl_450_U211 ( .A1(u4_srl_450_n168), .A2(u4_srl_450_n219), .B1(
        u4_srl_450_n170), .B2(u4_srl_450_n235), .ZN(u4_srl_450_n234) );
  AOI221_X1 u4_srl_450_U210 ( .B1(u4_srl_450_n217), .B2(u4_srl_450_n3), .C1(
        u4_srl_450_n197), .C2(u4_srl_450_n17), .A(u4_srl_450_n234), .ZN(
        u4_srl_450_n150) );
  AOI22_X1 u4_srl_450_U209 ( .A1(u4_srl_450_n69), .A2(u4_srl_450_n102), .B1(
        u4_srl_450_n77), .B2(u4_srl_450_n103), .ZN(u4_srl_450_n232) );
  AOI222_X1 u4_srl_450_U208 ( .A1(u4_srl_450_n73), .A2(u4_srl_450_n193), .B1(
        u4_srl_450_n229), .B2(u4_srl_450_n190), .C1(u4_srl_450_n71), .C2(
        u4_srl_450_n192), .ZN(u4_srl_450_n233) );
  OAI211_X1 u4_srl_450_U207 ( .C1(u4_srl_450_n150), .C2(u4_srl_450_n2), .A(
        u4_srl_450_n232), .B(u4_srl_450_n233), .ZN(u4_N1372) );
  AOI22_X1 u4_srl_450_U206 ( .A1(u4_srl_450_n137), .A2(u4_srl_450_n180), .B1(
        u4_srl_450_n136), .B2(u4_srl_450_n182), .ZN(u4_srl_450_n231) );
  INV_X1 u4_srl_450_U205 ( .A(u4_srl_450_n231), .ZN(u4_srl_450_n230) );
  AOI221_X1 u4_srl_450_U204 ( .B1(u4_srl_450_n187), .B2(u4_srl_450_n3), .C1(
        u4_srl_450_n188), .C2(u4_srl_450_n18), .A(u4_srl_450_n230), .ZN(
        u4_srl_450_n148) );
  AOI22_X1 u4_srl_450_U203 ( .A1(u4_srl_450_n69), .A2(u4_srl_450_n93), .B1(
        u4_srl_450_n77), .B2(u4_srl_450_n94), .ZN(u4_srl_450_n227) );
  AOI222_X1 u4_srl_450_U202 ( .A1(u4_srl_450_n73), .A2(u4_srl_450_n184), .B1(
        u4_srl_450_n229), .B2(u4_srl_450_n181), .C1(u4_srl_450_n71), .C2(
        u4_srl_450_n183), .ZN(u4_srl_450_n228) );
  OAI211_X1 u4_srl_450_U201 ( .C1(u4_srl_450_n148), .C2(u4_srl_450_n2), .A(
        u4_srl_450_n227), .B(u4_srl_450_n228), .ZN(u4_N1373) );
  OAI22_X1 u4_srl_450_U200 ( .A1(u4_srl_450_n226), .A2(u4_srl_450_n124), .B1(
        u4_srl_450_n147), .B2(u4_srl_450_n2), .ZN(u4_N1374) );
  AOI22_X1 u4_srl_450_U199 ( .A1(u4_srl_450_n137), .A2(u4_srl_450_n165), .B1(
        u4_srl_450_n136), .B2(u4_srl_450_n166), .ZN(u4_srl_450_n225) );
  INV_X1 u4_srl_450_U198 ( .A(u4_srl_450_n225), .ZN(u4_srl_450_n224) );
  AOI221_X1 u4_srl_450_U197 ( .B1(u4_srl_450_n72), .B2(u4_srl_450_n3), .C1(
        u4_srl_450_n74), .C2(u4_srl_450_n18), .A(u4_srl_450_n224), .ZN(
        u4_srl_450_n210) );
  OAI22_X1 u4_srl_450_U196 ( .A1(u4_srl_450_n168), .A2(u4_srl_450_n122), .B1(
        u4_srl_450_n170), .B2(u4_srl_450_n223), .ZN(u4_srl_450_n222) );
  AOI221_X1 u4_srl_450_U195 ( .B1(u4_srl_450_n198), .B2(u4_srl_450_n3), .C1(
        u4_srl_450_n201), .C2(u4_srl_450_n18), .A(u4_srl_450_n222), .ZN(
        u4_srl_450_n146) );
  OAI22_X1 u4_srl_450_U194 ( .A1(u4_srl_450_n210), .A2(u4_srl_450_n124), .B1(
        u4_srl_450_n146), .B2(u4_srl_450_n2), .ZN(u4_N1375) );
  AOI22_X1 u4_srl_450_U193 ( .A1(u4_srl_450_n137), .A2(u4_srl_450_n197), .B1(
        u4_srl_450_n136), .B2(u4_srl_450_n192), .ZN(u4_srl_450_n221) );
  INV_X1 u4_srl_450_U192 ( .A(u4_srl_450_n221), .ZN(u4_srl_450_n220) );
  AOI221_X1 u4_srl_450_U191 ( .B1(u4_srl_450_n193), .B2(u4_srl_450_n3), .C1(
        u4_srl_450_n102), .C2(u4_srl_450_n18), .A(u4_srl_450_n220), .ZN(
        u4_srl_450_n156) );
  OAI22_X1 u4_srl_450_U190 ( .A1(u4_srl_450_n168), .A2(u4_srl_450_n121), .B1(
        u4_srl_450_n170), .B2(u4_srl_450_n219), .ZN(u4_srl_450_n218) );
  AOI221_X1 u4_srl_450_U189 ( .B1(u4_srl_450_n191), .B2(u4_srl_450_n3), .C1(
        u4_srl_450_n217), .C2(u4_srl_450_n17), .A(u4_srl_450_n218), .ZN(
        u4_srl_450_n145) );
  OAI22_X1 u4_srl_450_U188 ( .A1(u4_srl_450_n156), .A2(u4_srl_450_n124), .B1(
        u4_srl_450_n145), .B2(u4_srl_450_n2), .ZN(u4_N1376) );
  AOI22_X1 u4_srl_450_U187 ( .A1(u4_srl_450_n137), .A2(u4_srl_450_n188), .B1(
        u4_srl_450_n136), .B2(u4_srl_450_n183), .ZN(u4_srl_450_n216) );
  INV_X1 u4_srl_450_U186 ( .A(u4_srl_450_n216), .ZN(u4_srl_450_n215) );
  AOI221_X1 u4_srl_450_U185 ( .B1(u4_srl_450_n184), .B2(u4_srl_450_n3), .C1(
        u4_srl_450_n93), .C2(u4_srl_450_n18), .A(u4_srl_450_n215), .ZN(
        u4_srl_450_n135) );
  AOI222_X1 u4_srl_450_U184 ( .A1(u4_srl_450_n187), .A2(u4_srl_450_n17), .B1(
        u4_srl_450_n182), .B2(u4_srl_450_n3), .C1(u4_srl_450_n214), .C2(
        u4_shift_right[3]), .ZN(u4_srl_450_n128) );
  OAI22_X1 u4_srl_450_U183 ( .A1(u4_srl_450_n135), .A2(u4_srl_450_n124), .B1(
        u4_srl_450_n128), .B2(u4_srl_450_n2), .ZN(u4_N1377) );
  AOI22_X1 u4_srl_450_U182 ( .A1(n3522), .A2(u4_srl_450_n12), .B1(n3521), .B2(
        u4_srl_450_n143), .ZN(u4_srl_450_n213) );
  OAI221_X1 u4_srl_450_U181 ( .B1(u4_srl_450_n6), .B2(u4_srl_450_n21), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n64), .A(u4_srl_450_n213), .ZN(
        u4_srl_450_n206) );
  AOI22_X1 u4_srl_450_U180 ( .A1(n3527), .A2(u4_srl_450_n12), .B1(n3528), .B2(
        u4_srl_450_n143), .ZN(u4_srl_450_n212) );
  OAI221_X1 u4_srl_450_U179 ( .B1(u4_srl_450_n6), .B2(u4_srl_450_n27), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n62), .A(u4_srl_450_n212), .ZN(
        u4_srl_450_n78) );
  AOI22_X1 u4_srl_450_U178 ( .A1(n3562), .A2(u4_srl_450_n12), .B1(n3524), .B2(
        u4_srl_450_n143), .ZN(u4_srl_450_n211) );
  OAI221_X1 u4_srl_450_U177 ( .B1(u4_srl_450_n6), .B2(u4_srl_450_n24), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n23), .A(u4_srl_450_n211), .ZN(
        u4_srl_450_n111) );
  AOI222_X1 u4_srl_450_U176 ( .A1(u4_srl_450_n78), .A2(u4_srl_450_n136), .B1(
        u4_srl_450_n70), .B2(u4_srl_450_n137), .C1(u4_srl_450_n111), .C2(
        u4_srl_450_n3), .ZN(u4_srl_450_n209) );
  MUX2_X1 u4_srl_450_U175 ( .A(u4_srl_450_n209), .B(u4_srl_450_n210), .S(
        u4_shift_right[4]), .Z(u4_srl_450_n208) );
  INV_X1 u4_srl_450_U174 ( .A(u4_srl_450_n208), .ZN(u4_srl_450_n207) );
  AOI21_X1 u4_srl_450_U173 ( .B1(u4_srl_450_n130), .B2(u4_srl_450_n206), .A(
        u4_srl_450_n207), .ZN(u4_srl_450_n205) );
  OAI22_X1 u4_srl_450_U172 ( .A1(u4_shift_right[5]), .A2(u4_srl_450_n205), 
        .B1(u4_srl_450_n146), .B2(u4_srl_450_n129), .ZN(u4_N1359) );
  AOI22_X1 u4_srl_450_U171 ( .A1(u4_srl_450_n137), .A2(u4_srl_450_n179), .B1(
        u4_srl_450_n136), .B2(u4_srl_450_n174), .ZN(u4_srl_450_n204) );
  INV_X1 u4_srl_450_U170 ( .A(u4_srl_450_n204), .ZN(u4_srl_450_n203) );
  AOI221_X1 u4_srl_450_U169 ( .B1(u4_srl_450_n175), .B2(u4_srl_450_n3), .C1(
        u4_srl_450_n84), .C2(u4_srl_450_n18), .A(u4_srl_450_n203), .ZN(
        u4_srl_450_n113) );
  AOI222_X1 u4_srl_450_U168 ( .A1(u4_srl_450_n172), .A2(u4_srl_450_n3), .B1(
        u4_srl_450_n173), .B2(u4_srl_450_n136), .C1(u4_srl_450_n202), .C2(
        u4_srl_450_n17), .ZN(u4_srl_450_n118) );
  OAI22_X1 u4_srl_450_U167 ( .A1(u4_srl_450_n113), .A2(u4_srl_450_n124), .B1(
        u4_srl_450_n118), .B2(u4_srl_450_n2), .ZN(u4_N1378) );
  INV_X1 u4_srl_450_U166 ( .A(u4_srl_450_n201), .ZN(u4_srl_450_n171) );
  INV_X1 u4_srl_450_U165 ( .A(u4_srl_450_n165), .ZN(u4_srl_450_n200) );
  OAI22_X1 u4_srl_450_U164 ( .A1(u4_srl_450_n168), .A2(u4_srl_450_n171), .B1(
        u4_srl_450_n170), .B2(u4_srl_450_n200), .ZN(u4_srl_450_n199) );
  AOI221_X1 u4_srl_450_U163 ( .B1(u4_srl_450_n166), .B2(u4_srl_450_n3), .C1(
        u4_srl_450_n72), .C2(u4_srl_450_n18), .A(u4_srl_450_n199), .ZN(
        u4_srl_450_n107) );
  AOI222_X1 u4_srl_450_U162 ( .A1(u4_srl_450_n163), .A2(u4_srl_450_n3), .B1(
        u4_srl_450_n164), .B2(u4_srl_450_n136), .C1(u4_srl_450_n198), .C2(
        u4_srl_450_n17), .ZN(u4_srl_450_n112) );
  OAI22_X1 u4_srl_450_U161 ( .A1(u4_srl_450_n107), .A2(u4_srl_450_n124), .B1(
        u4_srl_450_n112), .B2(u4_srl_450_n2), .ZN(u4_N1379) );
  INV_X1 u4_srl_450_U160 ( .A(u4_srl_450_n197), .ZN(u4_srl_450_n196) );
  OAI22_X1 u4_srl_450_U159 ( .A1(u4_srl_450_n168), .A2(u4_srl_450_n195), .B1(
        u4_srl_450_n170), .B2(u4_srl_450_n196), .ZN(u4_srl_450_n194) );
  AOI221_X1 u4_srl_450_U158 ( .B1(u4_srl_450_n192), .B2(u4_srl_450_n3), .C1(
        u4_srl_450_n193), .C2(u4_srl_450_n18), .A(u4_srl_450_n194), .ZN(
        u4_srl_450_n98) );
  AOI222_X1 u4_srl_450_U157 ( .A1(u4_srl_450_n189), .A2(u4_srl_450_n3), .B1(
        u4_srl_450_n190), .B2(u4_srl_450_n136), .C1(u4_srl_450_n191), .C2(
        u4_srl_450_n17), .ZN(u4_srl_450_n106) );
  OAI22_X1 u4_srl_450_U156 ( .A1(u4_srl_450_n98), .A2(u4_srl_450_n124), .B1(
        u4_srl_450_n106), .B2(u4_srl_450_n2), .ZN(u4_N1380) );
  AOI22_X1 u4_srl_450_U155 ( .A1(u4_srl_450_n137), .A2(u4_srl_450_n187), .B1(
        u4_srl_450_n136), .B2(u4_srl_450_n188), .ZN(u4_srl_450_n186) );
  INV_X1 u4_srl_450_U154 ( .A(u4_srl_450_n186), .ZN(u4_srl_450_n185) );
  AOI221_X1 u4_srl_450_U153 ( .B1(u4_srl_450_n183), .B2(u4_srl_450_n3), .C1(
        u4_srl_450_n184), .C2(u4_srl_450_n18), .A(u4_srl_450_n185), .ZN(
        u4_srl_450_n89) );
  AOI222_X1 u4_srl_450_U152 ( .A1(u4_srl_450_n180), .A2(u4_srl_450_n3), .B1(
        u4_srl_450_n136), .B2(u4_srl_450_n181), .C1(u4_srl_450_n182), .C2(
        u4_srl_450_n17), .ZN(u4_srl_450_n97) );
  OAI22_X1 u4_srl_450_U151 ( .A1(u4_srl_450_n89), .A2(u4_srl_450_n124), .B1(
        u4_srl_450_n97), .B2(u4_srl_450_n2), .ZN(u4_N1381) );
  INV_X1 u4_srl_450_U150 ( .A(u4_srl_450_n179), .ZN(u4_srl_450_n178) );
  OAI22_X1 u4_srl_450_U149 ( .A1(u4_srl_450_n168), .A2(u4_srl_450_n177), .B1(
        u4_srl_450_n170), .B2(u4_srl_450_n178), .ZN(u4_srl_450_n176) );
  AOI221_X1 u4_srl_450_U148 ( .B1(u4_srl_450_n174), .B2(u4_srl_450_n3), .C1(
        u4_srl_450_n175), .C2(u4_srl_450_n17), .A(u4_srl_450_n176), .ZN(
        u4_srl_450_n80) );
  AOI22_X1 u4_srl_450_U147 ( .A1(u4_srl_450_n172), .A2(u4_srl_450_n17), .B1(
        u4_srl_450_n173), .B2(u4_srl_450_n138), .ZN(u4_srl_450_n88) );
  OAI22_X1 u4_srl_450_U146 ( .A1(u4_srl_450_n80), .A2(u4_srl_450_n124), .B1(
        u4_srl_450_n88), .B2(u4_srl_450_n2), .ZN(u4_N1382) );
  OAI22_X1 u4_srl_450_U145 ( .A1(u4_srl_450_n168), .A2(u4_srl_450_n169), .B1(
        u4_srl_450_n170), .B2(u4_srl_450_n171), .ZN(u4_srl_450_n167) );
  AOI221_X1 u4_srl_450_U144 ( .B1(u4_srl_450_n165), .B2(u4_srl_450_n138), .C1(
        u4_srl_450_n166), .C2(u4_srl_450_n17), .A(u4_srl_450_n167), .ZN(
        u4_srl_450_n65) );
  AOI22_X1 u4_srl_450_U143 ( .A1(u4_srl_450_n163), .A2(u4_srl_450_n18), .B1(
        u4_srl_450_n164), .B2(u4_srl_450_n138), .ZN(u4_srl_450_n79) );
  OAI22_X1 u4_srl_450_U142 ( .A1(u4_srl_450_n65), .A2(u4_srl_450_n124), .B1(
        u4_srl_450_n79), .B2(u4_srl_450_n66), .ZN(u4_N1383) );
  OAI22_X1 u4_srl_450_U141 ( .A1(u4_srl_450_n162), .A2(u4_srl_450_n124), .B1(
        u4_srl_450_n126), .B2(u4_srl_450_n66), .ZN(u4_N1384) );
  OAI22_X1 u4_srl_450_U140 ( .A1(u4_srl_450_n161), .A2(u4_srl_450_n124), .B1(
        u4_srl_450_n2), .B2(u4_srl_450_n125), .ZN(u4_N1385) );
  NAND2_X1 u4_srl_450_U139 ( .A1(u4_srl_450_n1), .A2(u4_srl_450_n17), .ZN(
        u4_srl_450_n149) );
  OAI22_X1 u4_srl_450_U138 ( .A1(u4_srl_450_n160), .A2(u4_srl_450_n124), .B1(
        u4_srl_450_n123), .B2(u4_srl_450_n149), .ZN(u4_N1386) );
  OAI22_X1 u4_srl_450_U137 ( .A1(u4_srl_450_n159), .A2(u4_srl_450_n124), .B1(
        u4_srl_450_n122), .B2(u4_srl_450_n149), .ZN(u4_N1387) );
  AOI22_X1 u4_srl_450_U136 ( .A1(n3563), .A2(u4_srl_450_n12), .B1(n3522), .B2(
        u4_srl_450_n143), .ZN(u4_srl_450_n158) );
  OAI221_X1 u4_srl_450_U135 ( .B1(u4_srl_450_n6), .B2(u4_srl_450_n22), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n21), .A(u4_srl_450_n158), .ZN(
        u4_srl_450_n152) );
  AOI22_X1 u4_srl_450_U134 ( .A1(n3525), .A2(u4_srl_450_n12), .B1(n3562), .B2(
        u4_srl_450_n143), .ZN(u4_srl_450_n157) );
  OAI221_X1 u4_srl_450_U133 ( .B1(u4_srl_450_n6), .B2(u4_srl_450_n26), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n24), .A(u4_srl_450_n157), .ZN(
        u4_srl_450_n105) );
  AOI222_X1 u4_srl_450_U132 ( .A1(u4_srl_450_n101), .A2(u4_srl_450_n136), .B1(
        u4_srl_450_n103), .B2(u4_srl_450_n137), .C1(u4_srl_450_n105), .C2(
        u4_srl_450_n3), .ZN(u4_srl_450_n155) );
  MUX2_X1 u4_srl_450_U131 ( .A(u4_srl_450_n155), .B(u4_srl_450_n156), .S(
        u4_shift_right[4]), .Z(u4_srl_450_n154) );
  INV_X1 u4_srl_450_U130 ( .A(u4_srl_450_n154), .ZN(u4_srl_450_n153) );
  AOI21_X1 u4_srl_450_U129 ( .B1(u4_srl_450_n130), .B2(u4_srl_450_n152), .A(
        u4_srl_450_n153), .ZN(u4_srl_450_n151) );
  OAI22_X1 u4_srl_450_U128 ( .A1(u4_shift_right[5]), .A2(u4_srl_450_n151), 
        .B1(u4_srl_450_n145), .B2(u4_srl_450_n129), .ZN(u4_N1360) );
  OAI22_X1 u4_srl_450_U127 ( .A1(u4_srl_450_n150), .A2(u4_srl_450_n124), .B1(
        u4_srl_450_n121), .B2(u4_srl_450_n149), .ZN(u4_N1388) );
  OAI22_X1 u4_srl_450_U126 ( .A1(u4_srl_450_n148), .A2(u4_srl_450_n124), .B1(
        u4_srl_450_n120), .B2(u4_srl_450_n149), .ZN(u4_N1389) );
  NOR2_X1 u4_srl_450_U125 ( .A1(u4_srl_450_n147), .A2(u4_srl_450_n124), .ZN(
        u4_N1390) );
  NOR2_X1 u4_srl_450_U124 ( .A1(u4_srl_450_n146), .A2(u4_srl_450_n124), .ZN(
        u4_N1391) );
  NOR2_X1 u4_srl_450_U123 ( .A1(u4_srl_450_n145), .A2(u4_srl_450_n124), .ZN(
        u4_N1392) );
  NOR2_X1 u4_srl_450_U122 ( .A1(u4_srl_450_n128), .A2(u4_srl_450_n124), .ZN(
        u4_N1393) );
  NOR2_X1 u4_srl_450_U121 ( .A1(u4_srl_450_n118), .A2(u4_srl_450_n124), .ZN(
        u4_N1394) );
  NOR2_X1 u4_srl_450_U120 ( .A1(u4_srl_450_n112), .A2(u4_srl_450_n124), .ZN(
        u4_N1395) );
  NOR2_X1 u4_srl_450_U119 ( .A1(u4_srl_450_n106), .A2(u4_srl_450_n124), .ZN(
        u4_N1396) );
  NOR2_X1 u4_srl_450_U118 ( .A1(u4_srl_450_n97), .A2(u4_srl_450_n124), .ZN(
        u4_N1397) );
  AOI22_X1 u4_srl_450_U117 ( .A1(n3523), .A2(u4_srl_450_n12), .B1(n3563), .B2(
        u4_srl_450_n143), .ZN(u4_srl_450_n144) );
  OAI221_X1 u4_srl_450_U116 ( .B1(u4_srl_450_n6), .B2(u4_srl_450_n63), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n22), .A(u4_srl_450_n144), .ZN(
        u4_srl_450_n131) );
  AOI22_X1 u4_srl_450_U115 ( .A1(n3526), .A2(u4_srl_450_n12), .B1(n3525), .B2(
        u4_srl_450_n16), .ZN(u4_srl_450_n141) );
  OAI221_X1 u4_srl_450_U114 ( .B1(u4_srl_450_n4), .B2(u4_srl_450_n25), .C1(
        u4_srl_450_n10), .C2(u4_srl_450_n26), .A(u4_srl_450_n141), .ZN(
        u4_srl_450_n96) );
  AOI222_X1 u4_srl_450_U113 ( .A1(u4_srl_450_n92), .A2(u4_srl_450_n136), .B1(
        u4_srl_450_n94), .B2(u4_srl_450_n137), .C1(u4_srl_450_n96), .C2(
        u4_srl_450_n3), .ZN(u4_srl_450_n134) );
  MUX2_X1 u4_srl_450_U112 ( .A(u4_srl_450_n134), .B(u4_srl_450_n135), .S(
        u4_shift_right[4]), .Z(u4_srl_450_n133) );
  INV_X1 u4_srl_450_U111 ( .A(u4_srl_450_n133), .ZN(u4_srl_450_n132) );
  AOI21_X1 u4_srl_450_U110 ( .B1(u4_srl_450_n130), .B2(u4_srl_450_n131), .A(
        u4_srl_450_n132), .ZN(u4_srl_450_n127) );
  OAI22_X1 u4_srl_450_U109 ( .A1(u4_shift_right[5]), .A2(u4_srl_450_n127), 
        .B1(u4_srl_450_n128), .B2(u4_srl_450_n129), .ZN(u4_N1361) );
  NOR2_X1 u4_srl_450_U108 ( .A1(u4_srl_450_n88), .A2(u4_srl_450_n124), .ZN(
        u4_N1398) );
  NOR2_X1 u4_srl_450_U107 ( .A1(u4_srl_450_n79), .A2(u4_srl_450_n124), .ZN(
        u4_N1399) );
  NOR2_X1 u4_srl_450_U106 ( .A1(u4_srl_450_n126), .A2(u4_srl_450_n124), .ZN(
        u4_N1400) );
  NOR2_X1 u4_srl_450_U105 ( .A1(u4_srl_450_n124), .A2(u4_srl_450_n125), .ZN(
        u4_N1401) );
  INV_X1 u4_srl_450_U104 ( .A(u4_srl_450_n77), .ZN(u4_srl_450_n119) );
  NOR2_X1 u4_srl_450_U103 ( .A1(u4_srl_450_n123), .A2(u4_srl_450_n119), .ZN(
        u4_N1402) );
  NOR2_X1 u4_srl_450_U102 ( .A1(u4_srl_450_n122), .A2(u4_srl_450_n119), .ZN(
        u4_N1403) );
  NOR2_X1 u4_srl_450_U101 ( .A1(u4_srl_450_n121), .A2(u4_srl_450_n119), .ZN(
        u4_N1404) );
  NOR2_X1 u4_srl_450_U100 ( .A1(u4_srl_450_n119), .A2(u4_srl_450_n120), .ZN(
        u4_N1405) );
  INV_X1 u4_srl_450_U99 ( .A(u4_srl_450_n118), .ZN(u4_srl_450_n116) );
  AOI22_X1 u4_srl_450_U98 ( .A1(u4_srl_450_n75), .A2(u4_srl_450_n116), .B1(
        u4_srl_450_n77), .B2(u4_srl_450_n117), .ZN(u4_srl_450_n114) );
  AOI222_X1 u4_srl_450_U97 ( .A1(u4_srl_450_n69), .A2(u4_srl_450_n87), .B1(
        u4_srl_450_n71), .B2(u4_srl_450_n85), .C1(u4_srl_450_n73), .C2(
        u4_srl_450_n83), .ZN(u4_srl_450_n115) );
  OAI211_X1 u4_srl_450_U96 ( .C1(u4_srl_450_n113), .C2(u4_srl_450_n2), .A(
        u4_srl_450_n114), .B(u4_srl_450_n115), .ZN(u4_N1362) );
  INV_X1 u4_srl_450_U95 ( .A(u4_srl_450_n112), .ZN(u4_srl_450_n110) );
  AOI22_X1 u4_srl_450_U94 ( .A1(u4_srl_450_n75), .A2(u4_srl_450_n110), .B1(
        u4_srl_450_n77), .B2(u4_srl_450_n111), .ZN(u4_srl_450_n108) );
  AOI222_X1 u4_srl_450_U93 ( .A1(u4_srl_450_n69), .A2(u4_srl_450_n78), .B1(
        u4_srl_450_n71), .B2(u4_srl_450_n74), .C1(u4_srl_450_n73), .C2(
        u4_srl_450_n70), .ZN(u4_srl_450_n109) );
  OAI211_X1 u4_srl_450_U92 ( .C1(u4_srl_450_n107), .C2(u4_srl_450_n2), .A(
        u4_srl_450_n108), .B(u4_srl_450_n109), .ZN(u4_N1363) );
  INV_X1 u4_srl_450_U91 ( .A(u4_srl_450_n106), .ZN(u4_srl_450_n104) );
  AOI22_X1 u4_srl_450_U90 ( .A1(u4_srl_450_n75), .A2(u4_srl_450_n104), .B1(
        u4_srl_450_n77), .B2(u4_srl_450_n105), .ZN(u4_srl_450_n99) );
  AOI222_X1 u4_srl_450_U89 ( .A1(u4_srl_450_n69), .A2(u4_srl_450_n101), .B1(
        u4_srl_450_n71), .B2(u4_srl_450_n102), .C1(u4_srl_450_n73), .C2(
        u4_srl_450_n103), .ZN(u4_srl_450_n100) );
  OAI211_X1 u4_srl_450_U88 ( .C1(u4_srl_450_n98), .C2(u4_srl_450_n2), .A(
        u4_srl_450_n99), .B(u4_srl_450_n100), .ZN(u4_N1364) );
  INV_X1 u4_srl_450_U87 ( .A(u4_srl_450_n97), .ZN(u4_srl_450_n95) );
  AOI22_X1 u4_srl_450_U86 ( .A1(u4_srl_450_n75), .A2(u4_srl_450_n95), .B1(
        u4_srl_450_n77), .B2(u4_srl_450_n96), .ZN(u4_srl_450_n90) );
  AOI222_X1 u4_srl_450_U85 ( .A1(u4_srl_450_n69), .A2(u4_srl_450_n92), .B1(
        u4_srl_450_n71), .B2(u4_srl_450_n93), .C1(u4_srl_450_n73), .C2(
        u4_srl_450_n94), .ZN(u4_srl_450_n91) );
  OAI211_X1 u4_srl_450_U84 ( .C1(u4_srl_450_n89), .C2(u4_srl_450_n2), .A(
        u4_srl_450_n90), .B(u4_srl_450_n91), .ZN(u4_N1365) );
  INV_X1 u4_srl_450_U83 ( .A(u4_srl_450_n88), .ZN(u4_srl_450_n86) );
  AOI22_X1 u4_srl_450_U82 ( .A1(u4_srl_450_n75), .A2(u4_srl_450_n86), .B1(
        u4_srl_450_n77), .B2(u4_srl_450_n87), .ZN(u4_srl_450_n81) );
  AOI222_X1 u4_srl_450_U81 ( .A1(u4_srl_450_n69), .A2(u4_srl_450_n83), .B1(
        u4_srl_450_n71), .B2(u4_srl_450_n84), .C1(u4_srl_450_n73), .C2(
        u4_srl_450_n85), .ZN(u4_srl_450_n82) );
  OAI211_X1 u4_srl_450_U80 ( .C1(u4_srl_450_n80), .C2(u4_srl_450_n2), .A(
        u4_srl_450_n81), .B(u4_srl_450_n82), .ZN(u4_N1366) );
  INV_X1 u4_srl_450_U79 ( .A(u4_srl_450_n79), .ZN(u4_srl_450_n76) );
  AOI22_X1 u4_srl_450_U78 ( .A1(u4_srl_450_n75), .A2(u4_srl_450_n76), .B1(
        u4_srl_450_n77), .B2(u4_srl_450_n78), .ZN(u4_srl_450_n67) );
  AOI222_X1 u4_srl_450_U77 ( .A1(u4_srl_450_n69), .A2(u4_srl_450_n70), .B1(
        u4_srl_450_n71), .B2(u4_srl_450_n72), .C1(u4_srl_450_n73), .C2(
        u4_srl_450_n74), .ZN(u4_srl_450_n68) );
  OAI211_X1 u4_srl_450_U76 ( .C1(u4_srl_450_n65), .C2(u4_srl_450_n2), .A(
        u4_srl_450_n67), .B(u4_srl_450_n68), .ZN(u4_N1367) );
  INV_X4 u4_srl_450_U75 ( .A(n3563), .ZN(u4_srl_450_n64) );
  INV_X4 u4_srl_450_U74 ( .A(n3562), .ZN(u4_srl_450_n63) );
  INV_X4 u4_srl_450_U73 ( .A(n3561), .ZN(u4_srl_450_n62) );
  INV_X4 u4_srl_450_U72 ( .A(n3560), .ZN(u4_srl_450_n61) );
  INV_X4 u4_srl_450_U71 ( .A(n3559), .ZN(u4_srl_450_n60) );
  INV_X4 u4_srl_450_U70 ( .A(n3557), .ZN(u4_srl_450_n59) );
  INV_X4 u4_srl_450_U69 ( .A(fract_denorm[42]), .ZN(u4_srl_450_n58) );
  INV_X4 u4_srl_450_U68 ( .A(fract_denorm[44]), .ZN(u4_srl_450_n57) );
  INV_X4 u4_srl_450_U67 ( .A(fract_denorm[43]), .ZN(u4_srl_450_n56) );
  INV_X4 u4_srl_450_U66 ( .A(fract_denorm[46]), .ZN(u4_srl_450_n55) );
  INV_X4 u4_srl_450_U65 ( .A(fract_denorm[45]), .ZN(u4_srl_450_n54) );
  INV_X4 u4_srl_450_U64 ( .A(fract_denorm[41]), .ZN(u4_srl_450_n53) );
  INV_X4 u4_srl_450_U63 ( .A(fract_denorm[40]), .ZN(u4_srl_450_n52) );
  INV_X4 u4_srl_450_U62 ( .A(fract_denorm[39]), .ZN(u4_srl_450_n51) );
  INV_X4 u4_srl_450_U61 ( .A(fract_denorm[31]), .ZN(u4_srl_450_n50) );
  INV_X4 u4_srl_450_U60 ( .A(fract_denorm[36]), .ZN(u4_srl_450_n49) );
  INV_X4 u4_srl_450_U59 ( .A(fract_denorm[38]), .ZN(u4_srl_450_n48) );
  INV_X4 u4_srl_450_U58 ( .A(fract_denorm[37]), .ZN(u4_srl_450_n47) );
  INV_X4 u4_srl_450_U57 ( .A(fract_denorm[35]), .ZN(u4_srl_450_n46) );
  INV_X4 u4_srl_450_U56 ( .A(fract_denorm[34]), .ZN(u4_srl_450_n45) );
  INV_X4 u4_srl_450_U55 ( .A(fract_denorm[33]), .ZN(u4_srl_450_n44) );
  INV_X4 u4_srl_450_U54 ( .A(fract_denorm[32]), .ZN(u4_srl_450_n43) );
  INV_X4 u4_srl_450_U53 ( .A(fract_denorm[23]), .ZN(u4_srl_450_n42) );
  INV_X4 u4_srl_450_U52 ( .A(fract_denorm[28]), .ZN(u4_srl_450_n41) );
  INV_X4 u4_srl_450_U51 ( .A(fract_denorm[30]), .ZN(u4_srl_450_n40) );
  INV_X4 u4_srl_450_U50 ( .A(fract_denorm[29]), .ZN(u4_srl_450_n39) );
  INV_X4 u4_srl_450_U49 ( .A(fract_denorm[27]), .ZN(u4_srl_450_n38) );
  INV_X4 u4_srl_450_U48 ( .A(fract_denorm[26]), .ZN(u4_srl_450_n37) );
  INV_X4 u4_srl_450_U47 ( .A(fract_denorm[25]), .ZN(u4_srl_450_n36) );
  INV_X4 u4_srl_450_U46 ( .A(fract_denorm[24]), .ZN(u4_srl_450_n35) );
  INV_X4 u4_srl_450_U45 ( .A(fract_denorm[22]), .ZN(u4_srl_450_n34) );
  INV_X4 u4_srl_450_U44 ( .A(fract_denorm[21]), .ZN(u4_srl_450_n33) );
  INV_X4 u4_srl_450_U43 ( .A(n3534), .ZN(u4_srl_450_n32) );
  INV_X4 u4_srl_450_U42 ( .A(n3533), .ZN(u4_srl_450_n31) );
  INV_X4 u4_srl_450_U41 ( .A(n3532), .ZN(u4_srl_450_n30) );
  INV_X4 u4_srl_450_U40 ( .A(n3531), .ZN(u4_srl_450_n29) );
  INV_X4 u4_srl_450_U39 ( .A(n3530), .ZN(u4_srl_450_n28) );
  INV_X4 u4_srl_450_U38 ( .A(n3529), .ZN(u4_srl_450_n27) );
  INV_X4 u4_srl_450_U37 ( .A(n3528), .ZN(u4_srl_450_n26) );
  INV_X4 u4_srl_450_U36 ( .A(n3527), .ZN(u4_srl_450_n25) );
  INV_X4 u4_srl_450_U35 ( .A(n3526), .ZN(u4_srl_450_n24) );
  INV_X4 u4_srl_450_U34 ( .A(n3525), .ZN(u4_srl_450_n23) );
  INV_X4 u4_srl_450_U33 ( .A(n3524), .ZN(u4_srl_450_n22) );
  INV_X4 u4_srl_450_U32 ( .A(n3523), .ZN(u4_srl_450_n21) );
  INV_X4 u4_srl_450_U31 ( .A(n3522), .ZN(u4_srl_450_n20) );
  INV_X4 u4_srl_450_U30 ( .A(n2679), .ZN(u4_srl_450_n19) );
  INV_X4 u4_srl_450_U29 ( .A(u4_srl_450_n7), .ZN(u4_srl_450_n4) );
  INV_X4 u4_srl_450_U28 ( .A(u4_srl_450_n139), .ZN(u4_srl_450_n7) );
  INV_X4 u4_srl_450_U27 ( .A(u4_srl_450_n1), .ZN(u4_srl_450_n2) );
  INV_X4 u4_srl_450_U26 ( .A(u4_srl_450_n142), .ZN(u4_srl_450_n13) );
  INV_X4 u4_srl_450_U25 ( .A(u4_srl_450_n15), .ZN(u4_srl_450_n16) );
  INV_X4 u4_srl_450_U24 ( .A(u4_srl_450_n275), .ZN(u4_srl_450_n17) );
  INV_X4 u4_srl_450_U23 ( .A(u4_srl_450_n275), .ZN(u4_srl_450_n18) );
  INV_X4 u4_srl_450_U22 ( .A(u4_srl_450_n272), .ZN(u4_srl_450_n3) );
  INV_X4 u4_srl_450_U21 ( .A(u4_srl_450_n13), .ZN(u4_srl_450_n12) );
  INV_X4 u4_srl_450_U20 ( .A(u4_srl_450_n9), .ZN(u4_srl_450_n8) );
  INV_X4 u4_srl_450_U19 ( .A(u4_srl_450_n10), .ZN(u4_srl_450_n9) );
  INV_X4 u4_srl_450_U18 ( .A(u4_srl_450_n11), .ZN(u4_srl_450_n10) );
  INV_X4 u4_srl_450_U17 ( .A(u4_srl_450_n66), .ZN(u4_srl_450_n1) );
  INV_X4 u4_srl_450_U16 ( .A(u4_srl_450_n15), .ZN(u4_srl_450_n14) );
  INV_X4 u4_srl_450_U15 ( .A(u4_srl_450_n143), .ZN(u4_srl_450_n15) );
  NAND2_X2 u4_srl_450_U14 ( .A1(u4_srl_450_n276), .A2(u4_srl_450_n277), .ZN(
        u4_srl_450_n124) );
  INV_X4 u4_srl_450_U13 ( .A(u4_srl_450_n140), .ZN(u4_srl_450_n11) );
  INV_X4 u4_srl_450_U12 ( .A(u4_srl_450_n7), .ZN(u4_srl_450_n6) );
  NOR2_X2 u4_srl_450_U11 ( .A1(u4_srl_450_n275), .A2(u4_srl_450_n124), .ZN(
        u4_srl_450_n77) );
  NOR2_X2 u4_srl_450_U10 ( .A1(u4_srl_450_n272), .A2(u4_srl_450_n124), .ZN(
        u4_srl_450_n69) );
  NOR2_X2 u4_srl_450_U9 ( .A1(u4_srl_450_n124), .A2(u4_srl_450_n168), .ZN(
        u4_srl_450_n71) );
  NOR2_X2 u4_srl_450_U8 ( .A1(u4_srl_450_n170), .A2(u4_srl_450_n124), .ZN(
        u4_srl_450_n73) );
  NAND2_X2 u4_srl_450_U7 ( .A1(u4_shift_right[3]), .A2(u4_shift_right[2]), 
        .ZN(u4_srl_450_n168) );
  NAND2_X2 u4_srl_450_U6 ( .A1(u4_shift_right[3]), .A2(u4_srl_450_n302), .ZN(
        u4_srl_450_n170) );
  INV_X4 u4_srl_450_U5 ( .A(u4_srl_450_n168), .ZN(u4_srl_450_n137) );
  INV_X4 u4_srl_450_U4 ( .A(u4_srl_450_n170), .ZN(u4_srl_450_n136) );
  INV_X4 u4_srl_450_U3 ( .A(u4_srl_450_n7), .ZN(u4_srl_450_n5) );
  NAND2_X1 u4_sll_479_U54 ( .A1(u4_f2i_shft_6_), .A2(u4_sll_479_n19), .ZN(
        u4_sll_479_n21) );
  OR2_X1 u4_sll_479_U53 ( .A1(u4_sll_479_n19), .A2(u4_f2i_shft_6_), .ZN(
        u4_sll_479_n20) );
  NAND2_X1 u4_sll_479_U52 ( .A1(n2473), .A2(u4_sll_479_n20), .ZN(
        u4_sll_479_n27) );
  NAND2_X1 u4_sll_479_U51 ( .A1(u4_sll_479_n21), .A2(u4_sll_479_n27), .ZN(
        u4_sll_479_temp_int_SH_0_) );
  AND2_X1 u4_sll_479_U50 ( .A1(n3564), .A2(u4_sll_479_n4), .ZN(
        u4_sll_479_ML_int_1__0_) );
  AND2_X1 u4_sll_479_U49 ( .A1(n2679), .A2(u4_sll_479_n2), .ZN(
        u4_sll_479_MR_int_1__55_) );
  NAND2_X1 u4_sll_479_U48 ( .A1(u4_f2i_shft_1_), .A2(u4_sll_479_n20), .ZN(
        u4_sll_479_n26) );
  NAND2_X1 u4_sll_479_U47 ( .A1(u4_sll_479_n21), .A2(u4_sll_479_n26), .ZN(
        u4_sll_479_temp_int_SH_1_) );
  NAND2_X1 u4_sll_479_U46 ( .A1(u4_sll_479_ML_int_1__0_), .A2(u4_sll_479_n8), 
        .ZN(u4_sll_479_n24) );
  AND2_X1 u4_sll_479_U45 ( .A1(u4_sll_479_ML_int_1__1_), .A2(u4_sll_479_n8), 
        .ZN(u4_sll_479_ML_int_2__1_) );
  NAND2_X1 u4_sll_479_U44 ( .A1(u4_f2i_shft_2_), .A2(u4_sll_479_n20), .ZN(
        u4_sll_479_n25) );
  NAND2_X1 u4_sll_479_U43 ( .A1(u4_sll_479_n21), .A2(u4_sll_479_n25), .ZN(
        u4_sll_479_temp_int_SH_2_) );
  NOR2_X1 u4_sll_479_U42 ( .A1(u4_sll_479_n10), .A2(u4_sll_479_n24), .ZN(
        u4_sll_479_ML_int_3__0_) );
  NAND2_X1 u4_sll_479_U41 ( .A1(u4_f2i_shft_3_), .A2(u4_sll_479_n20), .ZN(
        u4_sll_479_n23) );
  NAND2_X1 u4_sll_479_U40 ( .A1(u4_sll_479_n21), .A2(u4_sll_479_n23), .ZN(
        u4_sll_479_temp_int_SH_3_) );
  NOR2_X1 u4_sll_479_U39 ( .A1(u4_sll_479_n11), .A2(u4_sll_479_temp_int_SH_3_), 
        .ZN(u4_sll_479_n22) );
  AND2_X1 u4_sll_479_U38 ( .A1(u4_sll_479_n22), .A2(u4_sll_479_ML_int_2__1_), 
        .ZN(u4_sll_479_ML_int_4__1_) );
  AND2_X1 u4_sll_479_U37 ( .A1(u4_sll_479_ML_int_2__2_), .A2(u4_sll_479_n22), 
        .ZN(u4_sll_479_ML_int_4__2_) );
  AND2_X1 u4_sll_479_U36 ( .A1(u4_sll_479_ML_int_2__3_), .A2(u4_sll_479_n22), 
        .ZN(u4_sll_479_ML_int_4__3_) );
  AND2_X1 u4_sll_479_U35 ( .A1(u4_sll_479_ML_int_3__4_), .A2(u4_sll_479_n14), 
        .ZN(u4_sll_479_ML_int_4__4_) );
  AND2_X1 u4_sll_479_U34 ( .A1(u4_sll_479_ML_int_3__5_), .A2(u4_sll_479_n14), 
        .ZN(u4_sll_479_ML_int_4__5_) );
  AND2_X1 u4_sll_479_U33 ( .A1(u4_sll_479_ML_int_3__6_), .A2(u4_sll_479_n14), 
        .ZN(u4_sll_479_ML_int_4__6_) );
  AND2_X1 u4_sll_479_U32 ( .A1(u4_sll_479_ML_int_3__7_), .A2(u4_sll_479_n14), 
        .ZN(u4_sll_479_ML_int_4__7_) );
  AND2_X1 u4_sll_479_U31 ( .A1(u4_sll_479_ML_int_6__49_), .A2(u4_sll_479_n19), 
        .ZN(u4_exp_f2i_1[49]) );
  AND2_X1 u4_sll_479_U30 ( .A1(u4_sll_479_ML_int_6__50_), .A2(u4_sll_479_n19), 
        .ZN(u4_exp_f2i_1[50]) );
  AND2_X1 u4_sll_479_U29 ( .A1(u4_sll_479_ML_int_6__51_), .A2(u4_sll_479_n19), 
        .ZN(u4_exp_f2i_1[51]) );
  AND2_X1 u4_sll_479_U28 ( .A1(u4_sll_479_ML_int_6__52_), .A2(u4_sll_479_n19), 
        .ZN(u4_exp_f2i_1[52]) );
  AND2_X1 u4_sll_479_U27 ( .A1(u4_sll_479_ML_int_6__53_), .A2(u4_sll_479_n19), 
        .ZN(u4_exp_f2i_1[53]) );
  AND2_X1 u4_sll_479_U26 ( .A1(u4_sll_479_ML_int_6__54_), .A2(u4_sll_479_n19), 
        .ZN(u4_exp_f2i_1[54]) );
  AND2_X1 u4_sll_479_U25 ( .A1(u4_sll_479_ML_int_6__55_), .A2(u4_sll_479_n19), 
        .ZN(u4_exp_f2i_1[55]) );
  AND2_X1 u4_sll_479_U24 ( .A1(u4_sll_479_ML_int_6__56_), .A2(u4_sll_479_n19), 
        .ZN(u4_exp_f2i_1[56]) );
  OAI21_X1 u4_sll_479_U23 ( .B1(u4_f2i_shft_4_), .B2(u4_sll_479_n18), .A(
        u4_sll_479_n20), .ZN(u4_sll_479_SHMAG[4]) );
  OAI21_X1 u4_sll_479_U22 ( .B1(u4_f2i_shft_5_), .B2(u4_sll_479_n18), .A(
        u4_sll_479_n20), .ZN(u4_sll_479_SHMAG[5]) );
  INV_X4 u4_sll_479_U21 ( .A(u4_f2i_shft_7_), .ZN(u4_sll_479_n19) );
  INV_X4 u4_sll_479_U20 ( .A(u4_sll_479_n21), .ZN(u4_sll_479_n18) );
  INV_X4 u4_sll_479_U19 ( .A(u4_sll_479_SHMAG[5]), .ZN(u4_sll_479_n17) );
  INV_X4 u4_sll_479_U18 ( .A(u4_sll_479_SHMAG[4]), .ZN(u4_sll_479_n16) );
  INV_X4 u4_sll_479_U17 ( .A(u4_sll_479_n24), .ZN(u4_sll_479_n15) );
  INV_X4 u4_sll_479_U16 ( .A(u4_sll_479_n14), .ZN(u4_sll_479_n13) );
  INV_X4 u4_sll_479_U15 ( .A(u4_sll_479_n9), .ZN(u4_sll_479_n11) );
  INV_X4 u4_sll_479_U14 ( .A(u4_sll_479_n9), .ZN(u4_sll_479_n10) );
  INV_X4 u4_sll_479_U13 ( .A(u4_sll_479_n9), .ZN(u4_sll_479_n12) );
  INV_X4 u4_sll_479_U12 ( .A(u4_sll_479_n7), .ZN(u4_sll_479_n6) );
  INV_X4 u4_sll_479_U11 ( .A(u4_sll_479_n4), .ZN(u4_sll_479_n1) );
  INV_X4 u4_sll_479_U10 ( .A(u4_sll_479_temp_int_SH_2_), .ZN(u4_sll_479_n9) );
  INV_X4 u4_sll_479_U9 ( .A(u4_sll_479_n7), .ZN(u4_sll_479_n5) );
  INV_X4 u4_sll_479_U8 ( .A(u4_sll_479_temp_int_SH_3_), .ZN(u4_sll_479_n14) );
  INV_X4 u4_sll_479_U7 ( .A(u4_sll_479_n4), .ZN(u4_sll_479_n2) );
  INV_X4 u4_sll_479_U6 ( .A(u4_sll_479_n4), .ZN(u4_sll_479_n3) );
  INV_X4 u4_sll_479_U5 ( .A(u4_sll_479_temp_int_SH_0_), .ZN(u4_sll_479_n4) );
  INV_X4 u4_sll_479_U4 ( .A(u4_sll_479_temp_int_SH_1_), .ZN(u4_sll_479_n8) );
  INV_X4 u4_sll_479_U3 ( .A(u4_sll_479_temp_int_SH_1_), .ZN(u4_sll_479_n7) );
  MUX2_X2 u4_sll_479_M1_0_1 ( .A(n3521), .B(n3564), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_1__1_) );
  MUX2_X2 u4_sll_479_M1_0_2 ( .A(n3522), .B(n3521), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_1__2_) );
  MUX2_X2 u4_sll_479_M1_0_3 ( .A(n3563), .B(n3522), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_1__3_) );
  MUX2_X2 u4_sll_479_M1_0_4 ( .A(n3523), .B(n3563), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_1__4_) );
  MUX2_X2 u4_sll_479_M1_0_5 ( .A(n3524), .B(n3523), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_1__5_) );
  MUX2_X2 u4_sll_479_M1_0_6 ( .A(n3562), .B(n3524), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_1__6_) );
  MUX2_X2 u4_sll_479_M1_0_7 ( .A(n3525), .B(n3562), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_1__7_) );
  MUX2_X2 u4_sll_479_M1_0_8 ( .A(n3526), .B(n3525), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_1__8_) );
  MUX2_X2 u4_sll_479_M1_0_9 ( .A(n3528), .B(n3526), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_1__9_) );
  MUX2_X2 u4_sll_479_M1_0_10 ( .A(n3527), .B(n3528), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_1__10_) );
  MUX2_X2 u4_sll_479_M1_0_11 ( .A(n3561), .B(n3527), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_1__11_) );
  MUX2_X2 u4_sll_479_M1_0_12 ( .A(n3529), .B(n3561), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_1__12_) );
  MUX2_X2 u4_sll_479_M1_0_13 ( .A(n3530), .B(n3529), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_1__13_) );
  MUX2_X2 u4_sll_479_M1_0_14 ( .A(n3560), .B(n3530), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_1__14_) );
  MUX2_X2 u4_sll_479_M1_0_15 ( .A(n3531), .B(n3560), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_1__15_) );
  MUX2_X2 u4_sll_479_M1_0_16 ( .A(n3532), .B(n3531), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_1__16_) );
  MUX2_X2 u4_sll_479_M1_0_17 ( .A(n3559), .B(n3532), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_1__17_) );
  MUX2_X2 u4_sll_479_M1_0_18 ( .A(n3533), .B(n3559), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_1__18_) );
  MUX2_X2 u4_sll_479_M1_0_19 ( .A(n3534), .B(n3533), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_1__19_) );
  MUX2_X2 u4_sll_479_M1_0_20 ( .A(n3557), .B(n3534), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_1__20_) );
  MUX2_X2 u4_sll_479_M1_0_21 ( .A(fract_denorm[21]), .B(n3557), .S(
        u4_sll_479_n1), .Z(u4_sll_479_ML_int_1__21_) );
  MUX2_X2 u4_sll_479_M1_0_22 ( .A(fract_denorm[22]), .B(fract_denorm[21]), .S(
        u4_sll_479_n1), .Z(u4_sll_479_ML_int_1__22_) );
  MUX2_X2 u4_sll_479_M1_0_23 ( .A(fract_denorm[23]), .B(fract_denorm[22]), .S(
        u4_sll_479_n3), .Z(u4_sll_479_ML_int_1__23_) );
  MUX2_X2 u4_sll_479_M1_0_24 ( .A(fract_denorm[24]), .B(fract_denorm[23]), .S(
        u4_sll_479_temp_int_SH_0_), .Z(u4_sll_479_ML_int_1__24_) );
  MUX2_X2 u4_sll_479_M1_0_25 ( .A(fract_denorm[25]), .B(fract_denorm[24]), .S(
        u4_sll_479_n3), .Z(u4_sll_479_ML_int_1__25_) );
  MUX2_X2 u4_sll_479_M1_0_26 ( .A(fract_denorm[26]), .B(fract_denorm[25]), .S(
        u4_sll_479_n1), .Z(u4_sll_479_ML_int_1__26_) );
  MUX2_X2 u4_sll_479_M1_0_27 ( .A(fract_denorm[27]), .B(fract_denorm[26]), .S(
        u4_sll_479_temp_int_SH_0_), .Z(u4_sll_479_ML_int_1__27_) );
  MUX2_X2 u4_sll_479_M1_0_28 ( .A(fract_denorm[28]), .B(fract_denorm[27]), .S(
        u4_sll_479_n3), .Z(u4_sll_479_ML_int_1__28_) );
  MUX2_X2 u4_sll_479_M1_0_29 ( .A(fract_denorm[29]), .B(fract_denorm[28]), .S(
        u4_sll_479_temp_int_SH_0_), .Z(u4_sll_479_ML_int_1__29_) );
  MUX2_X2 u4_sll_479_M1_0_30 ( .A(fract_denorm[30]), .B(fract_denorm[29]), .S(
        u4_sll_479_n3), .Z(u4_sll_479_ML_int_1__30_) );
  MUX2_X2 u4_sll_479_M1_0_31 ( .A(fract_denorm[31]), .B(fract_denorm[30]), .S(
        u4_sll_479_temp_int_SH_0_), .Z(u4_sll_479_ML_int_1__31_) );
  MUX2_X2 u4_sll_479_M1_0_32 ( .A(fract_denorm[32]), .B(fract_denorm[31]), .S(
        u4_sll_479_temp_int_SH_0_), .Z(u4_sll_479_ML_int_1__32_) );
  MUX2_X2 u4_sll_479_M1_0_33 ( .A(fract_denorm[33]), .B(fract_denorm[32]), .S(
        u4_sll_479_temp_int_SH_0_), .Z(u4_sll_479_ML_int_1__33_) );
  MUX2_X2 u4_sll_479_M1_0_34 ( .A(fract_denorm[34]), .B(fract_denorm[33]), .S(
        u4_sll_479_n1), .Z(u4_sll_479_ML_int_1__34_) );
  MUX2_X2 u4_sll_479_M1_0_35 ( .A(fract_denorm[35]), .B(fract_denorm[34]), .S(
        u4_sll_479_n1), .Z(u4_sll_479_ML_int_1__35_) );
  MUX2_X2 u4_sll_479_M1_0_36 ( .A(fract_denorm[36]), .B(fract_denorm[35]), .S(
        u4_sll_479_n2), .Z(u4_sll_479_ML_int_1__36_) );
  MUX2_X2 u4_sll_479_M1_0_37 ( .A(fract_denorm[37]), .B(fract_denorm[36]), .S(
        u4_sll_479_n2), .Z(u4_sll_479_ML_int_1__37_) );
  MUX2_X2 u4_sll_479_M1_0_38 ( .A(fract_denorm[38]), .B(fract_denorm[37]), .S(
        u4_sll_479_n1), .Z(u4_sll_479_ML_int_1__38_) );
  MUX2_X2 u4_sll_479_M1_0_39 ( .A(fract_denorm[39]), .B(fract_denorm[38]), .S(
        u4_sll_479_n1), .Z(u4_sll_479_ML_int_1__39_) );
  MUX2_X2 u4_sll_479_M1_0_40 ( .A(fract_denorm[40]), .B(fract_denorm[39]), .S(
        u4_sll_479_n1), .Z(u4_sll_479_ML_int_1__40_) );
  MUX2_X2 u4_sll_479_M1_0_41 ( .A(fract_denorm[41]), .B(fract_denorm[40]), .S(
        u4_sll_479_temp_int_SH_0_), .Z(u4_sll_479_ML_int_1__41_) );
  MUX2_X2 u4_sll_479_M1_0_42 ( .A(fract_denorm[42]), .B(fract_denorm[41]), .S(
        u4_sll_479_n3), .Z(u4_sll_479_ML_int_1__42_) );
  MUX2_X2 u4_sll_479_M1_0_43 ( .A(fract_denorm[43]), .B(fract_denorm[42]), .S(
        u4_sll_479_temp_int_SH_0_), .Z(u4_sll_479_ML_int_1__43_) );
  MUX2_X2 u4_sll_479_M1_0_44 ( .A(fract_denorm[44]), .B(fract_denorm[43]), .S(
        u4_sll_479_n1), .Z(u4_sll_479_ML_int_1__44_) );
  MUX2_X2 u4_sll_479_M1_0_45 ( .A(fract_denorm[45]), .B(fract_denorm[44]), .S(
        u4_sll_479_temp_int_SH_0_), .Z(u4_sll_479_ML_int_1__45_) );
  MUX2_X2 u4_sll_479_M1_0_46 ( .A(fract_denorm[46]), .B(fract_denorm[45]), .S(
        u4_sll_479_temp_int_SH_0_), .Z(u4_sll_479_ML_int_1__46_) );
  MUX2_X2 u4_sll_479_M1_0_47 ( .A(n2679), .B(fract_denorm[46]), .S(
        u4_sll_479_n3), .Z(u4_sll_479_ML_int_1__47_) );
  MUX2_X2 u4_sll_479_M1_0_48 ( .A(n2679), .B(n2679), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_1__48_) );
  MUX2_X2 u4_sll_479_M1_0_49 ( .A(n2679), .B(n2679), .S(
        u4_sll_479_temp_int_SH_0_), .Z(u4_sll_479_ML_int_1__49_) );
  MUX2_X2 u4_sll_479_M1_0_50 ( .A(n2679), .B(n2679), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_1__50_) );
  MUX2_X2 u4_sll_479_M1_0_51 ( .A(n2679), .B(n2679), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_1__51_) );
  MUX2_X2 u4_sll_479_M1_0_52 ( .A(n2679), .B(n2679), .S(
        u4_sll_479_temp_int_SH_0_), .Z(u4_sll_479_ML_int_1__52_) );
  MUX2_X2 u4_sll_479_M1_0_53 ( .A(n2679), .B(n2679), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_1__53_) );
  MUX2_X2 u4_sll_479_M1_0_54 ( .A(n2679), .B(n2679), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_1__54_) );
  MUX2_X2 u4_sll_479_M1_0_55 ( .A(n2679), .B(n2679), .S(u4_sll_479_n3), .Z(
        u4_sll_479_ML_int_1__55_) );
  MUX2_X2 u4_sll_479_M1_1_2 ( .A(u4_sll_479_ML_int_1__2_), .B(
        u4_sll_479_ML_int_1__0_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__2_) );
  MUX2_X2 u4_sll_479_M1_1_3 ( .A(u4_sll_479_ML_int_1__3_), .B(
        u4_sll_479_ML_int_1__1_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__3_) );
  MUX2_X2 u4_sll_479_M1_1_4 ( .A(u4_sll_479_ML_int_1__4_), .B(
        u4_sll_479_ML_int_1__2_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__4_) );
  MUX2_X2 u4_sll_479_M1_1_5 ( .A(u4_sll_479_ML_int_1__5_), .B(
        u4_sll_479_ML_int_1__3_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__5_) );
  MUX2_X2 u4_sll_479_M1_1_6 ( .A(u4_sll_479_ML_int_1__6_), .B(
        u4_sll_479_ML_int_1__4_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__6_) );
  MUX2_X2 u4_sll_479_M1_1_7 ( .A(u4_sll_479_ML_int_1__7_), .B(
        u4_sll_479_ML_int_1__5_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__7_) );
  MUX2_X2 u4_sll_479_M1_1_8 ( .A(u4_sll_479_ML_int_1__8_), .B(
        u4_sll_479_ML_int_1__6_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__8_) );
  MUX2_X2 u4_sll_479_M1_1_9 ( .A(u4_sll_479_ML_int_1__9_), .B(
        u4_sll_479_ML_int_1__7_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__9_) );
  MUX2_X2 u4_sll_479_M1_1_10 ( .A(u4_sll_479_ML_int_1__10_), .B(
        u4_sll_479_ML_int_1__8_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__10_) );
  MUX2_X2 u4_sll_479_M1_1_11 ( .A(u4_sll_479_ML_int_1__11_), .B(
        u4_sll_479_ML_int_1__9_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__11_) );
  MUX2_X2 u4_sll_479_M1_1_12 ( .A(u4_sll_479_ML_int_1__12_), .B(
        u4_sll_479_ML_int_1__10_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__12_) );
  MUX2_X2 u4_sll_479_M1_1_13 ( .A(u4_sll_479_ML_int_1__13_), .B(
        u4_sll_479_ML_int_1__11_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__13_) );
  MUX2_X2 u4_sll_479_M1_1_14 ( .A(u4_sll_479_ML_int_1__14_), .B(
        u4_sll_479_ML_int_1__12_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__14_) );
  MUX2_X2 u4_sll_479_M1_1_15 ( .A(u4_sll_479_ML_int_1__15_), .B(
        u4_sll_479_ML_int_1__13_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__15_) );
  MUX2_X2 u4_sll_479_M1_1_16 ( .A(u4_sll_479_ML_int_1__16_), .B(
        u4_sll_479_ML_int_1__14_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__16_) );
  MUX2_X2 u4_sll_479_M1_1_17 ( .A(u4_sll_479_ML_int_1__17_), .B(
        u4_sll_479_ML_int_1__15_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__17_) );
  MUX2_X2 u4_sll_479_M1_1_18 ( .A(u4_sll_479_ML_int_1__18_), .B(
        u4_sll_479_ML_int_1__16_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__18_) );
  MUX2_X2 u4_sll_479_M1_1_19 ( .A(u4_sll_479_ML_int_1__19_), .B(
        u4_sll_479_ML_int_1__17_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__19_) );
  MUX2_X2 u4_sll_479_M1_1_20 ( .A(u4_sll_479_ML_int_1__20_), .B(
        u4_sll_479_ML_int_1__18_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__20_) );
  MUX2_X2 u4_sll_479_M1_1_21 ( .A(u4_sll_479_ML_int_1__21_), .B(
        u4_sll_479_ML_int_1__19_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__21_) );
  MUX2_X2 u4_sll_479_M1_1_22 ( .A(u4_sll_479_ML_int_1__22_), .B(
        u4_sll_479_ML_int_1__20_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__22_) );
  MUX2_X2 u4_sll_479_M1_1_23 ( .A(u4_sll_479_ML_int_1__23_), .B(
        u4_sll_479_ML_int_1__21_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__23_) );
  MUX2_X2 u4_sll_479_M1_1_24 ( .A(u4_sll_479_ML_int_1__24_), .B(
        u4_sll_479_ML_int_1__22_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__24_) );
  MUX2_X2 u4_sll_479_M1_1_25 ( .A(u4_sll_479_ML_int_1__25_), .B(
        u4_sll_479_ML_int_1__23_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__25_) );
  MUX2_X2 u4_sll_479_M1_1_26 ( .A(u4_sll_479_ML_int_1__26_), .B(
        u4_sll_479_ML_int_1__24_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__26_) );
  MUX2_X2 u4_sll_479_M1_1_27 ( .A(u4_sll_479_ML_int_1__27_), .B(
        u4_sll_479_ML_int_1__25_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__27_) );
  MUX2_X2 u4_sll_479_M1_1_28 ( .A(u4_sll_479_ML_int_1__28_), .B(
        u4_sll_479_ML_int_1__26_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__28_) );
  MUX2_X2 u4_sll_479_M1_1_29 ( .A(u4_sll_479_ML_int_1__29_), .B(
        u4_sll_479_ML_int_1__27_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__29_) );
  MUX2_X2 u4_sll_479_M1_1_30 ( .A(u4_sll_479_ML_int_1__30_), .B(
        u4_sll_479_ML_int_1__28_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__30_) );
  MUX2_X2 u4_sll_479_M1_1_31 ( .A(u4_sll_479_ML_int_1__31_), .B(
        u4_sll_479_ML_int_1__29_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__31_) );
  MUX2_X2 u4_sll_479_M1_1_32 ( .A(u4_sll_479_ML_int_1__32_), .B(
        u4_sll_479_ML_int_1__30_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__32_) );
  MUX2_X2 u4_sll_479_M1_1_33 ( .A(u4_sll_479_ML_int_1__33_), .B(
        u4_sll_479_ML_int_1__31_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__33_) );
  MUX2_X2 u4_sll_479_M1_1_34 ( .A(u4_sll_479_ML_int_1__34_), .B(
        u4_sll_479_ML_int_1__32_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__34_) );
  MUX2_X2 u4_sll_479_M1_1_35 ( .A(u4_sll_479_ML_int_1__35_), .B(
        u4_sll_479_ML_int_1__33_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__35_) );
  MUX2_X2 u4_sll_479_M1_1_36 ( .A(u4_sll_479_ML_int_1__36_), .B(
        u4_sll_479_ML_int_1__34_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__36_) );
  MUX2_X2 u4_sll_479_M1_1_37 ( .A(u4_sll_479_ML_int_1__37_), .B(
        u4_sll_479_ML_int_1__35_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__37_) );
  MUX2_X2 u4_sll_479_M1_1_38 ( .A(u4_sll_479_ML_int_1__38_), .B(
        u4_sll_479_ML_int_1__36_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__38_) );
  MUX2_X2 u4_sll_479_M1_1_39 ( .A(u4_sll_479_ML_int_1__39_), .B(
        u4_sll_479_ML_int_1__37_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__39_) );
  MUX2_X2 u4_sll_479_M1_1_40 ( .A(u4_sll_479_ML_int_1__40_), .B(
        u4_sll_479_ML_int_1__38_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__40_) );
  MUX2_X2 u4_sll_479_M1_1_41 ( .A(u4_sll_479_ML_int_1__41_), .B(
        u4_sll_479_ML_int_1__39_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__41_) );
  MUX2_X2 u4_sll_479_M1_1_42 ( .A(u4_sll_479_ML_int_1__42_), .B(
        u4_sll_479_ML_int_1__40_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__42_) );
  MUX2_X2 u4_sll_479_M1_1_43 ( .A(u4_sll_479_ML_int_1__43_), .B(
        u4_sll_479_ML_int_1__41_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__43_) );
  MUX2_X2 u4_sll_479_M1_1_44 ( .A(u4_sll_479_ML_int_1__44_), .B(
        u4_sll_479_ML_int_1__42_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__44_) );
  MUX2_X2 u4_sll_479_M1_1_45 ( .A(u4_sll_479_ML_int_1__45_), .B(
        u4_sll_479_ML_int_1__43_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__45_) );
  MUX2_X2 u4_sll_479_M1_1_46 ( .A(u4_sll_479_ML_int_1__46_), .B(
        u4_sll_479_ML_int_1__44_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__46_) );
  MUX2_X2 u4_sll_479_M1_1_47 ( .A(u4_sll_479_ML_int_1__47_), .B(
        u4_sll_479_ML_int_1__45_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__47_) );
  MUX2_X2 u4_sll_479_M1_1_48 ( .A(u4_sll_479_ML_int_1__48_), .B(
        u4_sll_479_ML_int_1__46_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__48_) );
  MUX2_X2 u4_sll_479_M1_1_49 ( .A(u4_sll_479_ML_int_1__49_), .B(
        u4_sll_479_ML_int_1__47_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__49_) );
  MUX2_X2 u4_sll_479_M1_1_50 ( .A(u4_sll_479_ML_int_1__50_), .B(
        u4_sll_479_ML_int_1__48_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__50_) );
  MUX2_X2 u4_sll_479_M1_1_51 ( .A(u4_sll_479_ML_int_1__51_), .B(
        u4_sll_479_ML_int_1__49_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__51_) );
  MUX2_X2 u4_sll_479_M1_1_52 ( .A(u4_sll_479_ML_int_1__52_), .B(
        u4_sll_479_ML_int_1__50_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__52_) );
  MUX2_X2 u4_sll_479_M1_1_53 ( .A(u4_sll_479_ML_int_1__53_), .B(
        u4_sll_479_ML_int_1__51_), .S(u4_sll_479_n6), .Z(
        u4_sll_479_ML_int_2__53_) );
  MUX2_X2 u4_sll_479_M1_1_54 ( .A(u4_sll_479_ML_int_1__54_), .B(
        u4_sll_479_ML_int_1__52_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__54_) );
  MUX2_X2 u4_sll_479_M1_1_55 ( .A(u4_sll_479_ML_int_1__55_), .B(
        u4_sll_479_ML_int_1__53_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__55_) );
  MUX2_X2 u4_sll_479_M1_1_56 ( .A(u4_sll_479_MR_int_1__55_), .B(
        u4_sll_479_ML_int_1__54_), .S(u4_sll_479_n5), .Z(
        u4_sll_479_ML_int_2__56_) );
  MUX2_X2 u4_sll_479_M1_2_4 ( .A(u4_sll_479_ML_int_2__4_), .B(u4_sll_479_n15), 
        .S(u4_sll_479_n11), .Z(u4_sll_479_ML_int_3__4_) );
  MUX2_X2 u4_sll_479_M1_2_5 ( .A(u4_sll_479_ML_int_2__5_), .B(
        u4_sll_479_ML_int_2__1_), .S(u4_sll_479_n10), .Z(
        u4_sll_479_ML_int_3__5_) );
  MUX2_X2 u4_sll_479_M1_2_6 ( .A(u4_sll_479_ML_int_2__6_), .B(
        u4_sll_479_ML_int_2__2_), .S(u4_sll_479_n11), .Z(
        u4_sll_479_ML_int_3__6_) );
  MUX2_X2 u4_sll_479_M1_2_7 ( .A(u4_sll_479_ML_int_2__7_), .B(
        u4_sll_479_ML_int_2__3_), .S(u4_sll_479_n10), .Z(
        u4_sll_479_ML_int_3__7_) );
  MUX2_X2 u4_sll_479_M1_2_8 ( .A(u4_sll_479_ML_int_2__8_), .B(
        u4_sll_479_ML_int_2__4_), .S(u4_sll_479_n12), .Z(
        u4_sll_479_ML_int_3__8_) );
  MUX2_X2 u4_sll_479_M1_2_9 ( .A(u4_sll_479_ML_int_2__9_), .B(
        u4_sll_479_ML_int_2__5_), .S(u4_sll_479_n11), .Z(
        u4_sll_479_ML_int_3__9_) );
  MUX2_X2 u4_sll_479_M1_2_10 ( .A(u4_sll_479_ML_int_2__10_), .B(
        u4_sll_479_ML_int_2__6_), .S(u4_sll_479_n10), .Z(
        u4_sll_479_ML_int_3__10_) );
  MUX2_X2 u4_sll_479_M1_2_11 ( .A(u4_sll_479_ML_int_2__11_), .B(
        u4_sll_479_ML_int_2__7_), .S(u4_sll_479_n10), .Z(
        u4_sll_479_ML_int_3__11_) );
  MUX2_X2 u4_sll_479_M1_2_12 ( .A(u4_sll_479_ML_int_2__12_), .B(
        u4_sll_479_ML_int_2__8_), .S(u4_sll_479_n11), .Z(
        u4_sll_479_ML_int_3__12_) );
  MUX2_X2 u4_sll_479_M1_2_13 ( .A(u4_sll_479_ML_int_2__13_), .B(
        u4_sll_479_ML_int_2__9_), .S(u4_sll_479_n12), .Z(
        u4_sll_479_ML_int_3__13_) );
  MUX2_X2 u4_sll_479_M1_2_14 ( .A(u4_sll_479_ML_int_2__14_), .B(
        u4_sll_479_ML_int_2__10_), .S(u4_sll_479_n12), .Z(
        u4_sll_479_ML_int_3__14_) );
  MUX2_X2 u4_sll_479_M1_2_15 ( .A(u4_sll_479_ML_int_2__15_), .B(
        u4_sll_479_ML_int_2__11_), .S(u4_sll_479_n12), .Z(
        u4_sll_479_ML_int_3__15_) );
  MUX2_X2 u4_sll_479_M1_2_16 ( .A(u4_sll_479_ML_int_2__16_), .B(
        u4_sll_479_ML_int_2__12_), .S(u4_sll_479_n12), .Z(
        u4_sll_479_ML_int_3__16_) );
  MUX2_X2 u4_sll_479_M1_2_17 ( .A(u4_sll_479_ML_int_2__17_), .B(
        u4_sll_479_ML_int_2__13_), .S(u4_sll_479_n12), .Z(
        u4_sll_479_ML_int_3__17_) );
  MUX2_X2 u4_sll_479_M1_2_18 ( .A(u4_sll_479_ML_int_2__18_), .B(
        u4_sll_479_ML_int_2__14_), .S(u4_sll_479_n12), .Z(
        u4_sll_479_ML_int_3__18_) );
  MUX2_X2 u4_sll_479_M1_2_19 ( .A(u4_sll_479_ML_int_2__19_), .B(
        u4_sll_479_ML_int_2__15_), .S(u4_sll_479_n12), .Z(
        u4_sll_479_ML_int_3__19_) );
  MUX2_X2 u4_sll_479_M1_2_20 ( .A(u4_sll_479_ML_int_2__20_), .B(
        u4_sll_479_ML_int_2__16_), .S(u4_sll_479_n12), .Z(
        u4_sll_479_ML_int_3__20_) );
  MUX2_X2 u4_sll_479_M1_2_21 ( .A(u4_sll_479_ML_int_2__21_), .B(
        u4_sll_479_ML_int_2__17_), .S(u4_sll_479_n12), .Z(
        u4_sll_479_ML_int_3__21_) );
  MUX2_X2 u4_sll_479_M1_2_22 ( .A(u4_sll_479_ML_int_2__22_), .B(
        u4_sll_479_ML_int_2__18_), .S(u4_sll_479_n12), .Z(
        u4_sll_479_ML_int_3__22_) );
  MUX2_X2 u4_sll_479_M1_2_23 ( .A(u4_sll_479_ML_int_2__23_), .B(
        u4_sll_479_ML_int_2__19_), .S(u4_sll_479_n12), .Z(
        u4_sll_479_ML_int_3__23_) );
  MUX2_X2 u4_sll_479_M1_2_24 ( .A(u4_sll_479_ML_int_2__24_), .B(
        u4_sll_479_ML_int_2__20_), .S(u4_sll_479_n12), .Z(
        u4_sll_479_ML_int_3__24_) );
  MUX2_X2 u4_sll_479_M1_2_25 ( .A(u4_sll_479_ML_int_2__25_), .B(
        u4_sll_479_ML_int_2__21_), .S(u4_sll_479_n11), .Z(
        u4_sll_479_ML_int_3__25_) );
  MUX2_X2 u4_sll_479_M1_2_26 ( .A(u4_sll_479_ML_int_2__26_), .B(
        u4_sll_479_ML_int_2__22_), .S(u4_sll_479_n12), .Z(
        u4_sll_479_ML_int_3__26_) );
  MUX2_X2 u4_sll_479_M1_2_27 ( .A(u4_sll_479_ML_int_2__27_), .B(
        u4_sll_479_ML_int_2__23_), .S(u4_sll_479_n11), .Z(
        u4_sll_479_ML_int_3__27_) );
  MUX2_X2 u4_sll_479_M1_2_28 ( .A(u4_sll_479_ML_int_2__28_), .B(
        u4_sll_479_ML_int_2__24_), .S(u4_sll_479_n10), .Z(
        u4_sll_479_ML_int_3__28_) );
  MUX2_X2 u4_sll_479_M1_2_29 ( .A(u4_sll_479_ML_int_2__29_), .B(
        u4_sll_479_ML_int_2__25_), .S(u4_sll_479_n12), .Z(
        u4_sll_479_ML_int_3__29_) );
  MUX2_X2 u4_sll_479_M1_2_30 ( .A(u4_sll_479_ML_int_2__30_), .B(
        u4_sll_479_ML_int_2__26_), .S(u4_sll_479_n11), .Z(
        u4_sll_479_ML_int_3__30_) );
  MUX2_X2 u4_sll_479_M1_2_31 ( .A(u4_sll_479_ML_int_2__31_), .B(
        u4_sll_479_ML_int_2__27_), .S(u4_sll_479_n10), .Z(
        u4_sll_479_ML_int_3__31_) );
  MUX2_X2 u4_sll_479_M1_2_32 ( .A(u4_sll_479_ML_int_2__32_), .B(
        u4_sll_479_ML_int_2__28_), .S(u4_sll_479_n12), .Z(
        u4_sll_479_ML_int_3__32_) );
  MUX2_X2 u4_sll_479_M1_2_33 ( .A(u4_sll_479_ML_int_2__33_), .B(
        u4_sll_479_ML_int_2__29_), .S(u4_sll_479_n12), .Z(
        u4_sll_479_ML_int_3__33_) );
  MUX2_X2 u4_sll_479_M1_2_34 ( .A(u4_sll_479_ML_int_2__34_), .B(
        u4_sll_479_ML_int_2__30_), .S(u4_sll_479_n10), .Z(
        u4_sll_479_ML_int_3__34_) );
  MUX2_X2 u4_sll_479_M1_2_35 ( .A(u4_sll_479_ML_int_2__35_), .B(
        u4_sll_479_ML_int_2__31_), .S(u4_sll_479_n11), .Z(
        u4_sll_479_ML_int_3__35_) );
  MUX2_X2 u4_sll_479_M1_2_36 ( .A(u4_sll_479_ML_int_2__36_), .B(
        u4_sll_479_ML_int_2__32_), .S(u4_sll_479_n11), .Z(
        u4_sll_479_ML_int_3__36_) );
  MUX2_X2 u4_sll_479_M1_2_37 ( .A(u4_sll_479_ML_int_2__37_), .B(
        u4_sll_479_ML_int_2__33_), .S(u4_sll_479_n11), .Z(
        u4_sll_479_ML_int_3__37_) );
  MUX2_X2 u4_sll_479_M1_2_38 ( .A(u4_sll_479_ML_int_2__38_), .B(
        u4_sll_479_ML_int_2__34_), .S(u4_sll_479_n11), .Z(
        u4_sll_479_ML_int_3__38_) );
  MUX2_X2 u4_sll_479_M1_2_39 ( .A(u4_sll_479_ML_int_2__39_), .B(
        u4_sll_479_ML_int_2__35_), .S(u4_sll_479_n11), .Z(
        u4_sll_479_ML_int_3__39_) );
  MUX2_X2 u4_sll_479_M1_2_40 ( .A(u4_sll_479_ML_int_2__40_), .B(
        u4_sll_479_ML_int_2__36_), .S(u4_sll_479_n11), .Z(
        u4_sll_479_ML_int_3__40_) );
  MUX2_X2 u4_sll_479_M1_2_41 ( .A(u4_sll_479_ML_int_2__41_), .B(
        u4_sll_479_ML_int_2__37_), .S(u4_sll_479_n11), .Z(
        u4_sll_479_ML_int_3__41_) );
  MUX2_X2 u4_sll_479_M1_2_42 ( .A(u4_sll_479_ML_int_2__42_), .B(
        u4_sll_479_ML_int_2__38_), .S(u4_sll_479_n11), .Z(
        u4_sll_479_ML_int_3__42_) );
  MUX2_X2 u4_sll_479_M1_2_43 ( .A(u4_sll_479_ML_int_2__43_), .B(
        u4_sll_479_ML_int_2__39_), .S(u4_sll_479_n11), .Z(
        u4_sll_479_ML_int_3__43_) );
  MUX2_X2 u4_sll_479_M1_2_44 ( .A(u4_sll_479_ML_int_2__44_), .B(
        u4_sll_479_ML_int_2__40_), .S(u4_sll_479_n11), .Z(
        u4_sll_479_ML_int_3__44_) );
  MUX2_X2 u4_sll_479_M1_2_45 ( .A(u4_sll_479_ML_int_2__45_), .B(
        u4_sll_479_ML_int_2__41_), .S(u4_sll_479_n11), .Z(
        u4_sll_479_ML_int_3__45_) );
  MUX2_X2 u4_sll_479_M1_2_46 ( .A(u4_sll_479_ML_int_2__46_), .B(
        u4_sll_479_ML_int_2__42_), .S(u4_sll_479_n10), .Z(
        u4_sll_479_ML_int_3__46_) );
  MUX2_X2 u4_sll_479_M1_2_47 ( .A(u4_sll_479_ML_int_2__47_), .B(
        u4_sll_479_ML_int_2__43_), .S(u4_sll_479_n10), .Z(
        u4_sll_479_ML_int_3__47_) );
  MUX2_X2 u4_sll_479_M1_2_48 ( .A(u4_sll_479_ML_int_2__48_), .B(
        u4_sll_479_ML_int_2__44_), .S(u4_sll_479_n10), .Z(
        u4_sll_479_ML_int_3__48_) );
  MUX2_X2 u4_sll_479_M1_2_49 ( .A(u4_sll_479_ML_int_2__49_), .B(
        u4_sll_479_ML_int_2__45_), .S(u4_sll_479_n10), .Z(
        u4_sll_479_ML_int_3__49_) );
  MUX2_X2 u4_sll_479_M1_2_50 ( .A(u4_sll_479_ML_int_2__50_), .B(
        u4_sll_479_ML_int_2__46_), .S(u4_sll_479_n10), .Z(
        u4_sll_479_ML_int_3__50_) );
  MUX2_X2 u4_sll_479_M1_2_51 ( .A(u4_sll_479_ML_int_2__51_), .B(
        u4_sll_479_ML_int_2__47_), .S(u4_sll_479_n10), .Z(
        u4_sll_479_ML_int_3__51_) );
  MUX2_X2 u4_sll_479_M1_2_52 ( .A(u4_sll_479_ML_int_2__52_), .B(
        u4_sll_479_ML_int_2__48_), .S(u4_sll_479_n10), .Z(
        u4_sll_479_ML_int_3__52_) );
  MUX2_X2 u4_sll_479_M1_2_53 ( .A(u4_sll_479_ML_int_2__53_), .B(
        u4_sll_479_ML_int_2__49_), .S(u4_sll_479_n10), .Z(
        u4_sll_479_ML_int_3__53_) );
  MUX2_X2 u4_sll_479_M1_2_54 ( .A(u4_sll_479_ML_int_2__54_), .B(
        u4_sll_479_ML_int_2__50_), .S(u4_sll_479_n10), .Z(
        u4_sll_479_ML_int_3__54_) );
  MUX2_X2 u4_sll_479_M1_2_55 ( .A(u4_sll_479_ML_int_2__55_), .B(
        u4_sll_479_ML_int_2__51_), .S(u4_sll_479_n10), .Z(
        u4_sll_479_ML_int_3__55_) );
  MUX2_X2 u4_sll_479_M1_2_56 ( .A(u4_sll_479_ML_int_2__56_), .B(
        u4_sll_479_ML_int_2__52_), .S(u4_sll_479_n10), .Z(
        u4_sll_479_ML_int_3__56_) );
  MUX2_X2 u4_sll_479_M1_3_8 ( .A(u4_sll_479_ML_int_3__8_), .B(
        u4_sll_479_ML_int_3__0_), .S(u4_sll_479_n13), .Z(
        u4_sll_479_ML_int_4__8_) );
  MUX2_X2 u4_sll_479_M1_3_17 ( .A(u4_sll_479_ML_int_3__17_), .B(
        u4_sll_479_ML_int_3__9_), .S(u4_sll_479_n13), .Z(
        u4_sll_479_ML_int_4__17_) );
  MUX2_X2 u4_sll_479_M1_3_18 ( .A(u4_sll_479_ML_int_3__18_), .B(
        u4_sll_479_ML_int_3__10_), .S(u4_sll_479_temp_int_SH_3_), .Z(
        u4_sll_479_ML_int_4__18_) );
  MUX2_X2 u4_sll_479_M1_3_19 ( .A(u4_sll_479_ML_int_3__19_), .B(
        u4_sll_479_ML_int_3__11_), .S(u4_sll_479_temp_int_SH_3_), .Z(
        u4_sll_479_ML_int_4__19_) );
  MUX2_X2 u4_sll_479_M1_3_20 ( .A(u4_sll_479_ML_int_3__20_), .B(
        u4_sll_479_ML_int_3__12_), .S(u4_sll_479_n13), .Z(
        u4_sll_479_ML_int_4__20_) );
  MUX2_X2 u4_sll_479_M1_3_21 ( .A(u4_sll_479_ML_int_3__21_), .B(
        u4_sll_479_ML_int_3__13_), .S(u4_sll_479_temp_int_SH_3_), .Z(
        u4_sll_479_ML_int_4__21_) );
  MUX2_X2 u4_sll_479_M1_3_22 ( .A(u4_sll_479_ML_int_3__22_), .B(
        u4_sll_479_ML_int_3__14_), .S(u4_sll_479_temp_int_SH_3_), .Z(
        u4_sll_479_ML_int_4__22_) );
  MUX2_X2 u4_sll_479_M1_3_23 ( .A(u4_sll_479_ML_int_3__23_), .B(
        u4_sll_479_ML_int_3__15_), .S(u4_sll_479_n13), .Z(
        u4_sll_479_ML_int_4__23_) );
  MUX2_X2 u4_sll_479_M1_3_24 ( .A(u4_sll_479_ML_int_3__24_), .B(
        u4_sll_479_ML_int_3__16_), .S(u4_sll_479_n13), .Z(
        u4_sll_479_ML_int_4__24_) );
  MUX2_X2 u4_sll_479_M1_3_33 ( .A(u4_sll_479_ML_int_3__33_), .B(
        u4_sll_479_ML_int_3__25_), .S(u4_sll_479_temp_int_SH_3_), .Z(
        u4_sll_479_ML_int_4__33_) );
  MUX2_X2 u4_sll_479_M1_3_34 ( .A(u4_sll_479_ML_int_3__34_), .B(
        u4_sll_479_ML_int_3__26_), .S(u4_sll_479_temp_int_SH_3_), .Z(
        u4_sll_479_ML_int_4__34_) );
  MUX2_X2 u4_sll_479_M1_3_35 ( .A(u4_sll_479_ML_int_3__35_), .B(
        u4_sll_479_ML_int_3__27_), .S(u4_sll_479_n13), .Z(
        u4_sll_479_ML_int_4__35_) );
  MUX2_X2 u4_sll_479_M1_3_36 ( .A(u4_sll_479_ML_int_3__36_), .B(
        u4_sll_479_ML_int_3__28_), .S(u4_sll_479_temp_int_SH_3_), .Z(
        u4_sll_479_ML_int_4__36_) );
  MUX2_X2 u4_sll_479_M1_3_37 ( .A(u4_sll_479_ML_int_3__37_), .B(
        u4_sll_479_ML_int_3__29_), .S(u4_sll_479_temp_int_SH_3_), .Z(
        u4_sll_479_ML_int_4__37_) );
  MUX2_X2 u4_sll_479_M1_3_38 ( .A(u4_sll_479_ML_int_3__38_), .B(
        u4_sll_479_ML_int_3__30_), .S(u4_sll_479_temp_int_SH_3_), .Z(
        u4_sll_479_ML_int_4__38_) );
  MUX2_X2 u4_sll_479_M1_3_39 ( .A(u4_sll_479_ML_int_3__39_), .B(
        u4_sll_479_ML_int_3__31_), .S(u4_sll_479_n13), .Z(
        u4_sll_479_ML_int_4__39_) );
  MUX2_X2 u4_sll_479_M1_3_40 ( .A(u4_sll_479_ML_int_3__40_), .B(
        u4_sll_479_ML_int_3__32_), .S(u4_sll_479_n13), .Z(
        u4_sll_479_ML_int_4__40_) );
  MUX2_X2 u4_sll_479_M1_3_49 ( .A(u4_sll_479_ML_int_3__49_), .B(
        u4_sll_479_ML_int_3__41_), .S(u4_sll_479_n13), .Z(
        u4_sll_479_ML_int_4__49_) );
  MUX2_X2 u4_sll_479_M1_3_50 ( .A(u4_sll_479_ML_int_3__50_), .B(
        u4_sll_479_ML_int_3__42_), .S(u4_sll_479_n13), .Z(
        u4_sll_479_ML_int_4__50_) );
  MUX2_X2 u4_sll_479_M1_3_51 ( .A(u4_sll_479_ML_int_3__51_), .B(
        u4_sll_479_ML_int_3__43_), .S(u4_sll_479_n13), .Z(
        u4_sll_479_ML_int_4__51_) );
  MUX2_X2 u4_sll_479_M1_3_52 ( .A(u4_sll_479_ML_int_3__52_), .B(
        u4_sll_479_ML_int_3__44_), .S(u4_sll_479_temp_int_SH_3_), .Z(
        u4_sll_479_ML_int_4__52_) );
  MUX2_X2 u4_sll_479_M1_3_53 ( .A(u4_sll_479_ML_int_3__53_), .B(
        u4_sll_479_ML_int_3__45_), .S(u4_sll_479_n13), .Z(
        u4_sll_479_ML_int_4__53_) );
  MUX2_X2 u4_sll_479_M1_3_54 ( .A(u4_sll_479_ML_int_3__54_), .B(
        u4_sll_479_ML_int_3__46_), .S(u4_sll_479_temp_int_SH_3_), .Z(
        u4_sll_479_ML_int_4__54_) );
  MUX2_X2 u4_sll_479_M1_3_55 ( .A(u4_sll_479_ML_int_3__55_), .B(
        u4_sll_479_ML_int_3__47_), .S(u4_sll_479_temp_int_SH_3_), .Z(
        u4_sll_479_ML_int_4__55_) );
  MUX2_X2 u4_sll_479_M1_3_56 ( .A(u4_sll_479_ML_int_3__56_), .B(
        u4_sll_479_ML_int_3__48_), .S(u4_sll_479_n13), .Z(
        u4_sll_479_ML_int_4__56_) );
  MUX2_X2 u4_sll_479_M1_4_17 ( .A(u4_sll_479_ML_int_4__17_), .B(
        u4_sll_479_ML_int_4__1_), .S(u4_sll_479_n16), .Z(
        u4_sll_479_ML_int_5__17_) );
  MUX2_X2 u4_sll_479_M1_4_18 ( .A(u4_sll_479_ML_int_4__18_), .B(
        u4_sll_479_ML_int_4__2_), .S(u4_sll_479_n16), .Z(
        u4_sll_479_ML_int_5__18_) );
  MUX2_X2 u4_sll_479_M1_4_19 ( .A(u4_sll_479_ML_int_4__19_), .B(
        u4_sll_479_ML_int_4__3_), .S(u4_sll_479_n16), .Z(
        u4_sll_479_ML_int_5__19_) );
  MUX2_X2 u4_sll_479_M1_4_20 ( .A(u4_sll_479_ML_int_4__20_), .B(
        u4_sll_479_ML_int_4__4_), .S(u4_sll_479_n16), .Z(
        u4_sll_479_ML_int_5__20_) );
  MUX2_X2 u4_sll_479_M1_4_21 ( .A(u4_sll_479_ML_int_4__21_), .B(
        u4_sll_479_ML_int_4__5_), .S(u4_sll_479_n16), .Z(
        u4_sll_479_ML_int_5__21_) );
  MUX2_X2 u4_sll_479_M1_4_22 ( .A(u4_sll_479_ML_int_4__22_), .B(
        u4_sll_479_ML_int_4__6_), .S(u4_sll_479_n16), .Z(
        u4_sll_479_ML_int_5__22_) );
  MUX2_X2 u4_sll_479_M1_4_23 ( .A(u4_sll_479_ML_int_4__23_), .B(
        u4_sll_479_ML_int_4__7_), .S(u4_sll_479_n16), .Z(
        u4_sll_479_ML_int_5__23_) );
  MUX2_X2 u4_sll_479_M1_4_24 ( .A(u4_sll_479_ML_int_4__24_), .B(
        u4_sll_479_ML_int_4__8_), .S(u4_sll_479_n16), .Z(
        u4_sll_479_ML_int_5__24_) );
  MUX2_X2 u4_sll_479_M1_4_49 ( .A(u4_sll_479_ML_int_4__49_), .B(
        u4_sll_479_ML_int_4__33_), .S(u4_sll_479_n16), .Z(
        u4_sll_479_ML_int_5__49_) );
  MUX2_X2 u4_sll_479_M1_4_50 ( .A(u4_sll_479_ML_int_4__50_), .B(
        u4_sll_479_ML_int_4__34_), .S(u4_sll_479_n16), .Z(
        u4_sll_479_ML_int_5__50_) );
  MUX2_X2 u4_sll_479_M1_4_51 ( .A(u4_sll_479_ML_int_4__51_), .B(
        u4_sll_479_ML_int_4__35_), .S(u4_sll_479_n16), .Z(
        u4_sll_479_ML_int_5__51_) );
  MUX2_X2 u4_sll_479_M1_4_52 ( .A(u4_sll_479_ML_int_4__52_), .B(
        u4_sll_479_ML_int_4__36_), .S(u4_sll_479_n16), .Z(
        u4_sll_479_ML_int_5__52_) );
  MUX2_X2 u4_sll_479_M1_4_53 ( .A(u4_sll_479_ML_int_4__53_), .B(
        u4_sll_479_ML_int_4__37_), .S(u4_sll_479_n16), .Z(
        u4_sll_479_ML_int_5__53_) );
  MUX2_X2 u4_sll_479_M1_4_54 ( .A(u4_sll_479_ML_int_4__54_), .B(
        u4_sll_479_ML_int_4__38_), .S(u4_sll_479_n16), .Z(
        u4_sll_479_ML_int_5__54_) );
  MUX2_X2 u4_sll_479_M1_4_55 ( .A(u4_sll_479_ML_int_4__55_), .B(
        u4_sll_479_ML_int_4__39_), .S(u4_sll_479_n16), .Z(
        u4_sll_479_ML_int_5__55_) );
  MUX2_X2 u4_sll_479_M1_4_56 ( .A(u4_sll_479_ML_int_4__56_), .B(
        u4_sll_479_ML_int_4__40_), .S(u4_sll_479_n16), .Z(
        u4_sll_479_ML_int_5__56_) );
  MUX2_X2 u4_sll_479_M1_5_49 ( .A(u4_sll_479_ML_int_5__49_), .B(
        u4_sll_479_ML_int_5__17_), .S(u4_sll_479_n17), .Z(
        u4_sll_479_ML_int_6__49_) );
  MUX2_X2 u4_sll_479_M1_5_50 ( .A(u4_sll_479_ML_int_5__50_), .B(
        u4_sll_479_ML_int_5__18_), .S(u4_sll_479_n17), .Z(
        u4_sll_479_ML_int_6__50_) );
  MUX2_X2 u4_sll_479_M1_5_51 ( .A(u4_sll_479_ML_int_5__51_), .B(
        u4_sll_479_ML_int_5__19_), .S(u4_sll_479_n17), .Z(
        u4_sll_479_ML_int_6__51_) );
  MUX2_X2 u4_sll_479_M1_5_52 ( .A(u4_sll_479_ML_int_5__52_), .B(
        u4_sll_479_ML_int_5__20_), .S(u4_sll_479_n17), .Z(
        u4_sll_479_ML_int_6__52_) );
  MUX2_X2 u4_sll_479_M1_5_53 ( .A(u4_sll_479_ML_int_5__53_), .B(
        u4_sll_479_ML_int_5__21_), .S(u4_sll_479_n17), .Z(
        u4_sll_479_ML_int_6__53_) );
  MUX2_X2 u4_sll_479_M1_5_54 ( .A(u4_sll_479_ML_int_5__54_), .B(
        u4_sll_479_ML_int_5__22_), .S(u4_sll_479_n17), .Z(
        u4_sll_479_ML_int_6__54_) );
  MUX2_X2 u4_sll_479_M1_5_55 ( .A(u4_sll_479_ML_int_5__55_), .B(
        u4_sll_479_ML_int_5__23_), .S(u4_sll_479_n17), .Z(
        u4_sll_479_ML_int_6__55_) );
  MUX2_X2 u4_sll_479_M1_5_56 ( .A(u4_sll_479_ML_int_5__56_), .B(
        u4_sll_479_ML_int_5__24_), .S(u4_sll_479_n17), .Z(
        u4_sll_479_ML_int_6__56_) );
  INV_X4 u4_sub_467_U15 ( .A(u4_fi_ldz_2a_0_), .ZN(u4_sub_467_n10) );
  INV_X4 u4_sub_467_U14 ( .A(u4_fi_ldz_mi1_1_), .ZN(u4_sub_467_n9) );
  INV_X4 u4_sub_467_U13 ( .A(u4_fi_ldz_mi1_5_), .ZN(u4_sub_467_n8) );
  INV_X4 u4_sub_467_U12 ( .A(u4_fi_ldz_mi1_6_), .ZN(u4_sub_467_n7) );
  INV_X4 u4_sub_467_U11 ( .A(u4_fi_ldz_mi1_4_), .ZN(u4_sub_467_n6) );
  INV_X4 u4_sub_467_U10 ( .A(u4_fi_ldz_mi1_3_), .ZN(u4_sub_467_n5) );
  INV_X4 u4_sub_467_U9 ( .A(u4_fi_ldz_mi1_2_), .ZN(u4_sub_467_n4) );
  INV_X4 u4_sub_467_U8 ( .A(u4_exp_in_pl1_0_), .ZN(u4_sub_467_n3) );
  XNOR2_X2 u4_sub_467_U7 ( .A(u4_sub_467_n10), .B(u4_exp_in_pl1_0_), .ZN(
        u4_exp_next_mi_0_) );
  NAND2_X2 u4_sub_467_U6 ( .A1(u4_fi_ldz_2a_0_), .A2(u4_sub_467_n3), .ZN(
        u4_sub_467_carry_1_) );
  XNOR2_X2 u4_sub_467_U5 ( .A(u4_exp_in_pl1_8_), .B(u4_sub_467_carry_8_), .ZN(
        u4_exp_next_mi_8_) );
  INV_X4 u4_sub_467_U4 ( .A(u4_sub_467_carry_7_), .ZN(u4_sub_467_n2) );
  INV_X4 u4_sub_467_U3 ( .A(u4_exp_in_pl1_7_), .ZN(u4_sub_467_n1) );
  XNOR2_X2 u4_sub_467_U2 ( .A(u4_exp_in_pl1_7_), .B(u4_sub_467_carry_7_), .ZN(
        u4_exp_next_mi_7_) );
  NAND2_X2 u4_sub_467_U1 ( .A1(u4_sub_467_n1), .A2(u4_sub_467_n2), .ZN(
        u4_sub_467_carry_8_) );
  FA_X1 u4_sub_467_U2_1 ( .A(u4_exp_in_pl1_1_), .B(u4_sub_467_n9), .CI(
        u4_sub_467_carry_1_), .CO(u4_sub_467_carry_2_), .S(u4_exp_next_mi_1_)
         );
  FA_X1 u4_sub_467_U2_2 ( .A(u4_exp_in_pl1_2_), .B(u4_sub_467_n4), .CI(
        u4_sub_467_carry_2_), .CO(u4_sub_467_carry_3_), .S(u4_exp_next_mi_2_)
         );
  FA_X1 u4_sub_467_U2_3 ( .A(u4_exp_in_pl1_3_), .B(u4_sub_467_n5), .CI(
        u4_sub_467_carry_3_), .CO(u4_sub_467_carry_4_), .S(u4_exp_next_mi_3_)
         );
  FA_X1 u4_sub_467_U2_4 ( .A(u4_exp_in_pl1_4_), .B(u4_sub_467_n6), .CI(
        u4_sub_467_carry_4_), .CO(u4_sub_467_carry_5_), .S(u4_exp_next_mi_4_)
         );
  FA_X1 u4_sub_467_U2_5 ( .A(u4_exp_in_pl1_5_), .B(u4_sub_467_n8), .CI(
        u4_sub_467_carry_5_), .CO(u4_sub_467_carry_6_), .S(u4_exp_next_mi_5_)
         );
  FA_X1 u4_sub_467_U2_6 ( .A(u4_exp_in_pl1_6_), .B(u4_sub_467_n7), .CI(
        u4_sub_467_carry_6_), .CO(u4_sub_467_carry_7_), .S(u4_exp_next_mi_6_)
         );
  INV_X4 u4_sub_493_U11 ( .A(u4_ldz_all_0_), .ZN(u4_sub_493_n8) );
  INV_X4 u4_sub_493_U10 ( .A(u4_ldz_all_1_), .ZN(u4_sub_493_n7) );
  INV_X4 u4_sub_493_U9 ( .A(u4_ldz_all_2_), .ZN(u4_sub_493_n6) );
  INV_X4 u4_sub_493_U8 ( .A(u4_ldz_all_3_), .ZN(u4_sub_493_n5) );
  INV_X4 u4_sub_493_U7 ( .A(u4_ldz_all_4_), .ZN(u4_sub_493_n4) );
  INV_X4 u4_sub_493_U6 ( .A(u4_ldz_all_5_), .ZN(u4_sub_493_n3) );
  INV_X4 u4_sub_493_U5 ( .A(u4_ldz_all_6_), .ZN(u4_sub_493_n2) );
  INV_X4 u4_sub_493_U4 ( .A(u4_exp_in_pl1_0_), .ZN(u4_sub_493_n1) );
  XNOR2_X2 u4_sub_493_U3 ( .A(u4_sub_493_n8), .B(u4_exp_in_pl1_0_), .ZN(
        u4_div_exp2_0_) );
  NAND2_X2 u4_sub_493_U2 ( .A1(u4_ldz_all_0_), .A2(u4_sub_493_n1), .ZN(
        u4_sub_493_carry[1]) );
  XNOR2_X2 u4_sub_493_U1 ( .A(u4_exp_in_pl1_7_), .B(u4_sub_493_carry[7]), .ZN(
        u4_div_exp2_7_) );
  FA_X1 u4_sub_493_U2_1 ( .A(u4_exp_in_pl1_1_), .B(u4_sub_493_n7), .CI(
        u4_sub_493_carry[1]), .CO(u4_sub_493_carry[2]), .S(u4_div_exp2_1_) );
  FA_X1 u4_sub_493_U2_2 ( .A(u4_exp_in_pl1_2_), .B(u4_sub_493_n6), .CI(
        u4_sub_493_carry[2]), .CO(u4_sub_493_carry[3]), .S(u4_div_exp2_2_) );
  FA_X1 u4_sub_493_U2_3 ( .A(u4_exp_in_pl1_3_), .B(u4_sub_493_n5), .CI(
        u4_sub_493_carry[3]), .CO(u4_sub_493_carry[4]), .S(u4_div_exp2_3_) );
  FA_X1 u4_sub_493_U2_4 ( .A(u4_exp_in_pl1_4_), .B(u4_sub_493_n4), .CI(
        u4_sub_493_carry[4]), .CO(u4_sub_493_carry[5]), .S(u4_div_exp2_4_) );
  FA_X1 u4_sub_493_U2_5 ( .A(u4_exp_in_pl1_5_), .B(u4_sub_493_n3), .CI(
        u4_sub_493_carry[5]), .CO(u4_sub_493_carry[6]), .S(u4_div_exp2_5_) );
  FA_X1 u4_sub_493_U2_6 ( .A(u4_exp_in_pl1_6_), .B(u4_sub_493_n2), .CI(
        u4_sub_493_carry[6]), .CO(u4_sub_493_carry[7]), .S(u4_div_exp2_6_) );
  INV_X4 u4_add_463_U1 ( .A(n2650), .ZN(u4_exp_in_pl1_0_) );
  HA_X1 u4_add_463_U1_1_1 ( .A(n2681), .B(n2650), .CO(u4_add_463_carry[2]), 
        .S(u4_exp_in_pl1_1_) );
  HA_X1 u4_add_463_U1_1_2 ( .A(n2682), .B(u4_add_463_carry[2]), .CO(
        u4_add_463_carry[3]), .S(u4_exp_in_pl1_2_) );
  HA_X1 u4_add_463_U1_1_3 ( .A(n2683), .B(u4_add_463_carry[3]), .CO(
        u4_add_463_carry[4]), .S(u4_exp_in_pl1_3_) );
  HA_X1 u4_add_463_U1_1_4 ( .A(n2684), .B(u4_add_463_carry[4]), .CO(
        u4_add_463_carry[5]), .S(u4_exp_in_pl1_4_) );
  HA_X1 u4_add_463_U1_1_5 ( .A(n2685), .B(u4_add_463_carry[5]), .CO(
        u4_add_463_carry[6]), .S(u4_exp_in_pl1_5_) );
  HA_X1 u4_add_463_U1_1_6 ( .A(n2686), .B(u4_add_463_carry[6]), .CO(
        u4_add_463_carry[7]), .S(u4_exp_in_pl1_6_) );
  HA_X1 u4_add_463_U1_1_7 ( .A(n2687), .B(u4_add_463_carry[7]), .CO(
        u4_exp_in_pl1_8_), .S(u4_exp_in_pl1_7_) );
  XOR2_X2 u4_add_491_U3 ( .A(u4_exp_in_mi1_8_), .B(u4_add_491_carry[8]), .Z(
        u4_div_exp1_8_) );
  XOR2_X2 u4_add_491_U2 ( .A(u4_fi_ldz_2a_0_), .B(n2473), .Z(u4_div_exp1_0_)
         );
  AND2_X4 u4_add_491_U1 ( .A1(u4_fi_ldz_2a_0_), .A2(n2473), .ZN(u4_add_491_n1)
         );
  FA_X1 u4_add_491_U1_1 ( .A(u4_exp_in_mi1_1_), .B(u4_fi_ldz_2a_1_), .CI(
        u4_add_491_n1), .CO(u4_add_491_carry[2]), .S(u4_div_exp1_1_) );
  FA_X1 u4_add_491_U1_2 ( .A(u4_exp_in_mi1_2_), .B(n2723), .CI(
        u4_add_491_carry[2]), .CO(u4_add_491_carry[3]), .S(u4_div_exp1_2_) );
  FA_X1 u4_add_491_U1_3 ( .A(u4_exp_in_mi1_3_), .B(u4_fi_ldz_2a_3_), .CI(
        u4_add_491_carry[3]), .CO(u4_add_491_carry[4]), .S(u4_div_exp1_3_) );
  FA_X1 u4_add_491_U1_4 ( .A(u4_exp_in_mi1_4_), .B(u4_fi_ldz_2a_4_), .CI(
        u4_add_491_carry[4]), .CO(u4_add_491_carry[5]), .S(u4_div_exp1_4_) );
  FA_X1 u4_add_491_U1_5 ( .A(u4_exp_in_mi1_5_), .B(u4_fi_ldz_2a_5_), .CI(
        u4_add_491_carry[5]), .CO(u4_add_491_carry[6]), .S(u4_div_exp1_5_) );
  FA_X1 u4_add_491_U1_6 ( .A(u4_exp_in_mi1_6_), .B(n2543), .CI(
        u4_add_491_carry[6]), .CO(u4_add_491_carry[7]), .S(u4_div_exp1_6_) );
  FA_X1 u4_add_491_U1_7 ( .A(u4_exp_in_mi1_7_), .B(n2543), .CI(
        u4_add_491_carry[7]), .CO(u4_add_491_carry[8]), .S(u4_div_exp1_7_) );
  INV_X4 u4_sub_409_U16 ( .A(div_opa_ldz_r2[0]), .ZN(u4_sub_409_n6) );
  XNOR2_X2 u4_sub_409_U15 ( .A(u4_sub_409_n7), .B(div_opa_ldz_r2[0]), .ZN(
        u4_div_shft4[0]) );
  NAND2_X2 u4_sub_409_U14 ( .A1(n2650), .A2(u4_sub_409_n6), .ZN(
        u4_sub_409_carry_1_) );
  INV_X4 u4_sub_409_U13 ( .A(n2650), .ZN(u4_sub_409_n7) );
  AND2_X4 u4_sub_409_U12 ( .A1(u4_sub_409_n13), .A2(u4_sub_409_n2), .ZN(
        u4_sub_409_n5) );
  XOR2_X2 u4_sub_409_U11 ( .A(u4_sub_409_n13), .B(u4_sub_409_n2), .Z(
        u4_div_shft4[6]) );
  XOR2_X2 u4_sub_409_U10 ( .A(u4_sub_409_n12), .B(u4_sub_409_carry_5_), .Z(
        u4_div_shft4[5]) );
  AND2_X4 u4_sub_409_U9 ( .A1(u4_sub_409_n12), .A2(u4_sub_409_carry_5_), .ZN(
        u4_sub_409_n2) );
  XOR2_X2 u4_sub_409_U8 ( .A(u4_sub_409_n14), .B(u4_sub_409_n5), .Z(
        u4_div_shft4[7]) );
  INV_X4 u4_sub_409_U7 ( .A(n2687), .ZN(u4_sub_409_n14) );
  INV_X4 u4_sub_409_U6 ( .A(n2686), .ZN(u4_sub_409_n13) );
  INV_X4 u4_sub_409_U5 ( .A(n2685), .ZN(u4_sub_409_n12) );
  INV_X4 u4_sub_409_U4 ( .A(n2684), .ZN(u4_sub_409_n11) );
  INV_X4 u4_sub_409_U3 ( .A(n2683), .ZN(u4_sub_409_n10) );
  INV_X4 u4_sub_409_U2 ( .A(n2682), .ZN(u4_sub_409_n9) );
  INV_X4 u4_sub_409_U1 ( .A(n2681), .ZN(u4_sub_409_n8) );
  FA_X1 u4_sub_409_U2_1 ( .A(div_opa_ldz_r2[1]), .B(u4_sub_409_n8), .CI(
        u4_sub_409_carry_1_), .CO(u4_sub_409_carry_2_), .S(u4_div_shft4[1]) );
  FA_X1 u4_sub_409_U2_2 ( .A(div_opa_ldz_r2[2]), .B(u4_sub_409_n9), .CI(
        u4_sub_409_carry_2_), .CO(u4_sub_409_carry_3_), .S(u4_div_shft4[2]) );
  FA_X1 u4_sub_409_U2_3 ( .A(div_opa_ldz_r2[3]), .B(u4_sub_409_n10), .CI(
        u4_sub_409_carry_3_), .CO(u4_sub_409_carry_4_), .S(u4_div_shft4[3]) );
  FA_X1 u4_sub_409_U2_4 ( .A(div_opa_ldz_r2[4]), .B(u4_sub_409_n11), .CI(
        u4_sub_409_carry_4_), .CO(u4_sub_409_carry_5_), .S(u4_div_shft4[4]) );
  AND2_X4 u4_add_408_U7 ( .A1(n2686), .A2(u4_add_408_n5), .ZN(u4_add_408_n7)
         );
  AND2_X4 u4_add_408_U6 ( .A1(n2650), .A2(div_opa_ldz_r2[0]), .ZN(
        u4_add_408_n6) );
  AND2_X4 u4_add_408_U5 ( .A1(n2685), .A2(u4_add_408_carry_5_), .ZN(
        u4_add_408_n5) );
  XOR2_X2 u4_add_408_U4 ( .A(n2650), .B(div_opa_ldz_r2[0]), .Z(u4_div_shft3_0_) );
  XOR2_X2 u4_add_408_U3 ( .A(n2686), .B(u4_add_408_n5), .Z(u4_div_shft3_6_) );
  XOR2_X2 u4_add_408_U2 ( .A(n2687), .B(u4_add_408_n7), .Z(u4_div_shft3_7_) );
  XOR2_X2 u4_add_408_U1 ( .A(n2685), .B(u4_add_408_carry_5_), .Z(
        u4_div_shft3_5_) );
  FA_X1 u4_add_408_U1_1 ( .A(div_opa_ldz_r2[1]), .B(n2681), .CI(u4_add_408_n6), 
        .CO(u4_add_408_carry_2_), .S(u4_div_shft3_1_) );
  FA_X1 u4_add_408_U1_2 ( .A(div_opa_ldz_r2[2]), .B(n2682), .CI(
        u4_add_408_carry_2_), .CO(u4_add_408_carry_3_), .S(u4_div_shft3_2_) );
  FA_X1 u4_add_408_U1_3 ( .A(div_opa_ldz_r2[3]), .B(n2683), .CI(
        u4_add_408_carry_3_), .CO(u4_add_408_carry_4_), .S(u4_div_shft3_3_) );
  FA_X1 u4_add_408_U1_4 ( .A(div_opa_ldz_r2[4]), .B(n2684), .CI(
        u4_add_408_carry_4_), .CO(u4_add_408_carry_5_), .S(u4_div_shft3_4_) );
  INV_X1 u4_add_393_U1 ( .A(u4_fract_out_0_), .ZN(u4_fract_out_pl1_0_) );
  HA_X1 u4_add_393_U1_1_1 ( .A(u4_fract_out_1_), .B(u4_fract_out_0_), .CO(
        u4_add_393_carry[2]), .S(u4_fract_out_pl1_1_) );
  HA_X1 u4_add_393_U1_1_2 ( .A(u4_fract_out_2_), .B(u4_add_393_carry[2]), .CO(
        u4_add_393_carry[3]), .S(u4_fract_out_pl1_2_) );
  HA_X1 u4_add_393_U1_1_3 ( .A(u4_fract_out_3_), .B(u4_add_393_carry[3]), .CO(
        u4_add_393_carry[4]), .S(u4_fract_out_pl1_3_) );
  HA_X1 u4_add_393_U1_1_4 ( .A(u4_fract_out_4_), .B(u4_add_393_carry[4]), .CO(
        u4_add_393_carry[5]), .S(u4_fract_out_pl1_4_) );
  HA_X1 u4_add_393_U1_1_5 ( .A(u4_fract_out_5_), .B(u4_add_393_carry[5]), .CO(
        u4_add_393_carry[6]), .S(u4_fract_out_pl1_5_) );
  HA_X1 u4_add_393_U1_1_6 ( .A(u4_fract_out_6_), .B(u4_add_393_carry[6]), .CO(
        u4_add_393_carry[7]), .S(u4_fract_out_pl1_6_) );
  HA_X1 u4_add_393_U1_1_7 ( .A(u4_fract_out_7_), .B(u4_add_393_carry[7]), .CO(
        u4_add_393_carry[8]), .S(u4_fract_out_pl1_7_) );
  HA_X1 u4_add_393_U1_1_8 ( .A(u4_fract_out_8_), .B(u4_add_393_carry[8]), .CO(
        u4_add_393_carry[9]), .S(u4_fract_out_pl1_8_) );
  HA_X1 u4_add_393_U1_1_9 ( .A(u4_fract_out_9_), .B(u4_add_393_carry[9]), .CO(
        u4_add_393_carry[10]), .S(u4_fract_out_pl1_9_) );
  HA_X1 u4_add_393_U1_1_10 ( .A(u4_fract_out_10_), .B(u4_add_393_carry[10]), 
        .CO(u4_add_393_carry[11]), .S(u4_fract_out_pl1_10_) );
  HA_X1 u4_add_393_U1_1_11 ( .A(u4_fract_out_11_), .B(u4_add_393_carry[11]), 
        .CO(u4_add_393_carry[12]), .S(u4_fract_out_pl1_11_) );
  HA_X1 u4_add_393_U1_1_12 ( .A(u4_fract_out_12_), .B(u4_add_393_carry[12]), 
        .CO(u4_add_393_carry[13]), .S(u4_fract_out_pl1_12_) );
  HA_X1 u4_add_393_U1_1_13 ( .A(u4_fract_out_13_), .B(u4_add_393_carry[13]), 
        .CO(u4_add_393_carry[14]), .S(u4_fract_out_pl1_13_) );
  HA_X1 u4_add_393_U1_1_14 ( .A(u4_fract_out_14_), .B(u4_add_393_carry[14]), 
        .CO(u4_add_393_carry[15]), .S(u4_fract_out_pl1_14_) );
  HA_X1 u4_add_393_U1_1_15 ( .A(u4_fract_out_15_), .B(u4_add_393_carry[15]), 
        .CO(u4_add_393_carry[16]), .S(u4_fract_out_pl1_15_) );
  HA_X1 u4_add_393_U1_1_16 ( .A(u4_fract_out_16_), .B(u4_add_393_carry[16]), 
        .CO(u4_add_393_carry[17]), .S(u4_fract_out_pl1_16_) );
  HA_X1 u4_add_393_U1_1_17 ( .A(u4_fract_out_17_), .B(u4_add_393_carry[17]), 
        .CO(u4_add_393_carry[18]), .S(u4_fract_out_pl1_17_) );
  HA_X1 u4_add_393_U1_1_18 ( .A(u4_fract_out_18_), .B(u4_add_393_carry[18]), 
        .CO(u4_add_393_carry[19]), .S(u4_fract_out_pl1_18_) );
  HA_X1 u4_add_393_U1_1_19 ( .A(u4_fract_out_19_), .B(u4_add_393_carry[19]), 
        .CO(u4_add_393_carry[20]), .S(u4_fract_out_pl1_19_) );
  HA_X1 u4_add_393_U1_1_20 ( .A(u4_fract_out_20_), .B(u4_add_393_carry[20]), 
        .CO(u4_add_393_carry[21]), .S(u4_fract_out_pl1_20_) );
  HA_X1 u4_add_393_U1_1_21 ( .A(u4_fract_out_21_), .B(u4_add_393_carry[21]), 
        .CO(u4_add_393_carry[22]), .S(u4_fract_out_pl1_21_) );
  HA_X1 u4_add_393_U1_1_22 ( .A(u4_fract_out_22_), .B(u4_add_393_carry[22]), 
        .CO(u4_fract_out_pl1_23_), .S(u4_fract_out_pl1_22_) );
  INV_X4 u3_sub_60_U31 ( .A(fractb[26]), .ZN(u3_sub_60_n29) );
  INV_X4 u3_sub_60_U30 ( .A(fractb[25]), .ZN(u3_sub_60_n28) );
  INV_X4 u3_sub_60_U29 ( .A(fractb[24]), .ZN(u3_sub_60_n27) );
  INV_X4 u3_sub_60_U28 ( .A(fractb[23]), .ZN(u3_sub_60_n26) );
  INV_X4 u3_sub_60_U27 ( .A(fractb[22]), .ZN(u3_sub_60_n25) );
  INV_X4 u3_sub_60_U26 ( .A(fractb[21]), .ZN(u3_sub_60_n24) );
  INV_X4 u3_sub_60_U25 ( .A(fractb[20]), .ZN(u3_sub_60_n23) );
  INV_X4 u3_sub_60_U24 ( .A(fractb[19]), .ZN(u3_sub_60_n22) );
  INV_X4 u3_sub_60_U23 ( .A(fractb[18]), .ZN(u3_sub_60_n21) );
  INV_X4 u3_sub_60_U22 ( .A(fractb[17]), .ZN(u3_sub_60_n20) );
  INV_X4 u3_sub_60_U21 ( .A(fractb[16]), .ZN(u3_sub_60_n19) );
  INV_X4 u3_sub_60_U20 ( .A(fractb[15]), .ZN(u3_sub_60_n18) );
  INV_X4 u3_sub_60_U19 ( .A(fractb[14]), .ZN(u3_sub_60_n17) );
  INV_X4 u3_sub_60_U18 ( .A(fractb[13]), .ZN(u3_sub_60_n16) );
  INV_X4 u3_sub_60_U17 ( .A(fractb[12]), .ZN(u3_sub_60_n15) );
  INV_X4 u3_sub_60_U16 ( .A(fractb[11]), .ZN(u3_sub_60_n14) );
  INV_X4 u3_sub_60_U15 ( .A(fractb[10]), .ZN(u3_sub_60_n13) );
  INV_X4 u3_sub_60_U14 ( .A(fractb[9]), .ZN(u3_sub_60_n12) );
  INV_X4 u3_sub_60_U13 ( .A(fractb[8]), .ZN(u3_sub_60_n11) );
  INV_X4 u3_sub_60_U12 ( .A(fractb[7]), .ZN(u3_sub_60_n10) );
  INV_X4 u3_sub_60_U11 ( .A(fractb[6]), .ZN(u3_sub_60_n9) );
  INV_X4 u3_sub_60_U10 ( .A(fractb[5]), .ZN(u3_sub_60_n8) );
  INV_X4 u3_sub_60_U9 ( .A(fractb[4]), .ZN(u3_sub_60_n7) );
  INV_X4 u3_sub_60_U8 ( .A(fractb[3]), .ZN(u3_sub_60_n6) );
  INV_X4 u3_sub_60_U7 ( .A(fractb[2]), .ZN(u3_sub_60_n5) );
  INV_X4 u3_sub_60_U6 ( .A(fractb[1]), .ZN(u3_sub_60_n4) );
  INV_X4 u3_sub_60_U5 ( .A(fractb[0]), .ZN(u3_sub_60_n3) );
  INV_X4 u3_sub_60_U4 ( .A(u3_sub_60_carry[27]), .ZN(u3_N58) );
  INV_X4 u3_sub_60_U3 ( .A(fracta[0]), .ZN(u3_sub_60_n1) );
  XNOR2_X2 u3_sub_60_U2 ( .A(u3_sub_60_n3), .B(fracta[0]), .ZN(u3_N31) );
  NAND2_X2 u3_sub_60_U1 ( .A1(fractb[0]), .A2(u3_sub_60_n1), .ZN(
        u3_sub_60_carry[1]) );
  FA_X1 u3_sub_60_U2_1 ( .A(fracta[1]), .B(u3_sub_60_n4), .CI(
        u3_sub_60_carry[1]), .CO(u3_sub_60_carry[2]), .S(u3_N32) );
  FA_X1 u3_sub_60_U2_2 ( .A(fracta[2]), .B(u3_sub_60_n5), .CI(
        u3_sub_60_carry[2]), .CO(u3_sub_60_carry[3]), .S(u3_N33) );
  FA_X1 u3_sub_60_U2_3 ( .A(fracta[3]), .B(u3_sub_60_n6), .CI(
        u3_sub_60_carry[3]), .CO(u3_sub_60_carry[4]), .S(u3_N34) );
  FA_X1 u3_sub_60_U2_4 ( .A(fracta[4]), .B(u3_sub_60_n7), .CI(
        u3_sub_60_carry[4]), .CO(u3_sub_60_carry[5]), .S(u3_N35) );
  FA_X1 u3_sub_60_U2_5 ( .A(fracta[5]), .B(u3_sub_60_n8), .CI(
        u3_sub_60_carry[5]), .CO(u3_sub_60_carry[6]), .S(u3_N36) );
  FA_X1 u3_sub_60_U2_6 ( .A(fracta[6]), .B(u3_sub_60_n9), .CI(
        u3_sub_60_carry[6]), .CO(u3_sub_60_carry[7]), .S(u3_N37) );
  FA_X1 u3_sub_60_U2_7 ( .A(fracta[7]), .B(u3_sub_60_n10), .CI(
        u3_sub_60_carry[7]), .CO(u3_sub_60_carry[8]), .S(u3_N38) );
  FA_X1 u3_sub_60_U2_8 ( .A(fracta[8]), .B(u3_sub_60_n11), .CI(
        u3_sub_60_carry[8]), .CO(u3_sub_60_carry[9]), .S(u3_N39) );
  FA_X1 u3_sub_60_U2_9 ( .A(fracta[9]), .B(u3_sub_60_n12), .CI(
        u3_sub_60_carry[9]), .CO(u3_sub_60_carry[10]), .S(u3_N40) );
  FA_X1 u3_sub_60_U2_10 ( .A(fracta[10]), .B(u3_sub_60_n13), .CI(
        u3_sub_60_carry[10]), .CO(u3_sub_60_carry[11]), .S(u3_N41) );
  FA_X1 u3_sub_60_U2_11 ( .A(fracta[11]), .B(u3_sub_60_n14), .CI(
        u3_sub_60_carry[11]), .CO(u3_sub_60_carry[12]), .S(u3_N42) );
  FA_X1 u3_sub_60_U2_12 ( .A(fracta[12]), .B(u3_sub_60_n15), .CI(
        u3_sub_60_carry[12]), .CO(u3_sub_60_carry[13]), .S(u3_N43) );
  FA_X1 u3_sub_60_U2_13 ( .A(fracta[13]), .B(u3_sub_60_n16), .CI(
        u3_sub_60_carry[13]), .CO(u3_sub_60_carry[14]), .S(u3_N44) );
  FA_X1 u3_sub_60_U2_14 ( .A(fracta[14]), .B(u3_sub_60_n17), .CI(
        u3_sub_60_carry[14]), .CO(u3_sub_60_carry[15]), .S(u3_N45) );
  FA_X1 u3_sub_60_U2_15 ( .A(fracta[15]), .B(u3_sub_60_n18), .CI(
        u3_sub_60_carry[15]), .CO(u3_sub_60_carry[16]), .S(u3_N46) );
  FA_X1 u3_sub_60_U2_16 ( .A(fracta[16]), .B(u3_sub_60_n19), .CI(
        u3_sub_60_carry[16]), .CO(u3_sub_60_carry[17]), .S(u3_N47) );
  FA_X1 u3_sub_60_U2_17 ( .A(fracta[17]), .B(u3_sub_60_n20), .CI(
        u3_sub_60_carry[17]), .CO(u3_sub_60_carry[18]), .S(u3_N48) );
  FA_X1 u3_sub_60_U2_18 ( .A(fracta[18]), .B(u3_sub_60_n21), .CI(
        u3_sub_60_carry[18]), .CO(u3_sub_60_carry[19]), .S(u3_N49) );
  FA_X1 u3_sub_60_U2_19 ( .A(fracta[19]), .B(u3_sub_60_n22), .CI(
        u3_sub_60_carry[19]), .CO(u3_sub_60_carry[20]), .S(u3_N50) );
  FA_X1 u3_sub_60_U2_20 ( .A(fracta[20]), .B(u3_sub_60_n23), .CI(
        u3_sub_60_carry[20]), .CO(u3_sub_60_carry[21]), .S(u3_N51) );
  FA_X1 u3_sub_60_U2_21 ( .A(fracta[21]), .B(u3_sub_60_n24), .CI(
        u3_sub_60_carry[21]), .CO(u3_sub_60_carry[22]), .S(u3_N52) );
  FA_X1 u3_sub_60_U2_22 ( .A(fracta[22]), .B(u3_sub_60_n25), .CI(
        u3_sub_60_carry[22]), .CO(u3_sub_60_carry[23]), .S(u3_N53) );
  FA_X1 u3_sub_60_U2_23 ( .A(fracta[23]), .B(u3_sub_60_n26), .CI(
        u3_sub_60_carry[23]), .CO(u3_sub_60_carry[24]), .S(u3_N54) );
  FA_X1 u3_sub_60_U2_24 ( .A(fracta[24]), .B(u3_sub_60_n27), .CI(
        u3_sub_60_carry[24]), .CO(u3_sub_60_carry[25]), .S(u3_N55) );
  FA_X1 u3_sub_60_U2_25 ( .A(fracta[25]), .B(u3_sub_60_n28), .CI(
        u3_sub_60_carry[25]), .CO(u3_sub_60_carry[26]), .S(u3_N56) );
  FA_X1 u3_sub_60_U2_26 ( .A(fracta[26]), .B(u3_sub_60_n29), .CI(
        u3_sub_60_carry[26]), .CO(u3_sub_60_carry[27]), .S(u3_N57) );
  AND2_X4 u3_add_60_U2 ( .A1(fractb[0]), .A2(fracta[0]), .ZN(u3_add_60_n2) );
  XOR2_X2 u3_add_60_U1 ( .A(fractb[0]), .B(fracta[0]), .Z(u3_N3) );
  FA_X1 u3_add_60_U1_1 ( .A(fracta[1]), .B(fractb[1]), .CI(u3_add_60_n2), .CO(
        u3_add_60_carry[2]), .S(u3_N4) );
  FA_X1 u3_add_60_U1_2 ( .A(fracta[2]), .B(fractb[2]), .CI(u3_add_60_carry[2]), 
        .CO(u3_add_60_carry[3]), .S(u3_N5) );
  FA_X1 u3_add_60_U1_3 ( .A(fracta[3]), .B(fractb[3]), .CI(u3_add_60_carry[3]), 
        .CO(u3_add_60_carry[4]), .S(u3_N6) );
  FA_X1 u3_add_60_U1_4 ( .A(fracta[4]), .B(fractb[4]), .CI(u3_add_60_carry[4]), 
        .CO(u3_add_60_carry[5]), .S(u3_N7) );
  FA_X1 u3_add_60_U1_5 ( .A(fracta[5]), .B(fractb[5]), .CI(u3_add_60_carry[5]), 
        .CO(u3_add_60_carry[6]), .S(u3_N8) );
  FA_X1 u3_add_60_U1_6 ( .A(fracta[6]), .B(fractb[6]), .CI(u3_add_60_carry[6]), 
        .CO(u3_add_60_carry[7]), .S(u3_N9) );
  FA_X1 u3_add_60_U1_7 ( .A(fracta[7]), .B(fractb[7]), .CI(u3_add_60_carry[7]), 
        .CO(u3_add_60_carry[8]), .S(u3_N10) );
  FA_X1 u3_add_60_U1_8 ( .A(fracta[8]), .B(fractb[8]), .CI(u3_add_60_carry[8]), 
        .CO(u3_add_60_carry[9]), .S(u3_N11) );
  FA_X1 u3_add_60_U1_9 ( .A(fracta[9]), .B(fractb[9]), .CI(u3_add_60_carry[9]), 
        .CO(u3_add_60_carry[10]), .S(u3_N12) );
  FA_X1 u3_add_60_U1_10 ( .A(fracta[10]), .B(fractb[10]), .CI(
        u3_add_60_carry[10]), .CO(u3_add_60_carry[11]), .S(u3_N13) );
  FA_X1 u3_add_60_U1_11 ( .A(fracta[11]), .B(fractb[11]), .CI(
        u3_add_60_carry[11]), .CO(u3_add_60_carry[12]), .S(u3_N14) );
  FA_X1 u3_add_60_U1_12 ( .A(fracta[12]), .B(fractb[12]), .CI(
        u3_add_60_carry[12]), .CO(u3_add_60_carry[13]), .S(u3_N15) );
  FA_X1 u3_add_60_U1_13 ( .A(fracta[13]), .B(fractb[13]), .CI(
        u3_add_60_carry[13]), .CO(u3_add_60_carry[14]), .S(u3_N16) );
  FA_X1 u3_add_60_U1_14 ( .A(fracta[14]), .B(fractb[14]), .CI(
        u3_add_60_carry[14]), .CO(u3_add_60_carry[15]), .S(u3_N17) );
  FA_X1 u3_add_60_U1_15 ( .A(fracta[15]), .B(fractb[15]), .CI(
        u3_add_60_carry[15]), .CO(u3_add_60_carry[16]), .S(u3_N18) );
  FA_X1 u3_add_60_U1_16 ( .A(fracta[16]), .B(fractb[16]), .CI(
        u3_add_60_carry[16]), .CO(u3_add_60_carry[17]), .S(u3_N19) );
  FA_X1 u3_add_60_U1_17 ( .A(fracta[17]), .B(fractb[17]), .CI(
        u3_add_60_carry[17]), .CO(u3_add_60_carry[18]), .S(u3_N20) );
  FA_X1 u3_add_60_U1_18 ( .A(fracta[18]), .B(fractb[18]), .CI(
        u3_add_60_carry[18]), .CO(u3_add_60_carry[19]), .S(u3_N21) );
  FA_X1 u3_add_60_U1_19 ( .A(fracta[19]), .B(fractb[19]), .CI(
        u3_add_60_carry[19]), .CO(u3_add_60_carry[20]), .S(u3_N22) );
  FA_X1 u3_add_60_U1_20 ( .A(fracta[20]), .B(fractb[20]), .CI(
        u3_add_60_carry[20]), .CO(u3_add_60_carry[21]), .S(u3_N23) );
  FA_X1 u3_add_60_U1_21 ( .A(fracta[21]), .B(fractb[21]), .CI(
        u3_add_60_carry[21]), .CO(u3_add_60_carry[22]), .S(u3_N24) );
  FA_X1 u3_add_60_U1_22 ( .A(fracta[22]), .B(fractb[22]), .CI(
        u3_add_60_carry[22]), .CO(u3_add_60_carry[23]), .S(u3_N25) );
  FA_X1 u3_add_60_U1_23 ( .A(fracta[23]), .B(fractb[23]), .CI(
        u3_add_60_carry[23]), .CO(u3_add_60_carry[24]), .S(u3_N26) );
  FA_X1 u3_add_60_U1_24 ( .A(fracta[24]), .B(fractb[24]), .CI(
        u3_add_60_carry[24]), .CO(u3_add_60_carry[25]), .S(u3_N27) );
  FA_X1 u3_add_60_U1_25 ( .A(fracta[25]), .B(fractb[25]), .CI(
        u3_add_60_carry[25]), .CO(u3_add_60_carry[26]), .S(u3_N28) );
  FA_X1 u3_add_60_U1_26 ( .A(fracta[26]), .B(fractb[26]), .CI(
        u3_add_60_carry[26]), .CO(u3_N30), .S(u3_N29) );
  XOR2_X1 u2_add_114_U2 ( .A(u2_add_114_carry[7]), .B(u2_exp_tmp4_7_), .Z(
        u2_N49) );
  INV_X4 u2_add_114_U1 ( .A(u2_exp_tmp4_0_), .ZN(u2_N42) );
  HA_X1 u2_add_114_U1_1_1 ( .A(n1587), .B(u2_exp_tmp4_0_), .CO(
        u2_add_114_carry[2]), .S(u2_N43) );
  HA_X1 u2_add_114_U1_1_2 ( .A(n1586), .B(u2_add_114_carry[2]), .CO(
        u2_add_114_carry[3]), .S(u2_N44) );
  HA_X1 u2_add_114_U1_1_3 ( .A(n1585), .B(u2_add_114_carry[3]), .CO(
        u2_add_114_carry[4]), .S(u2_N45) );
  HA_X1 u2_add_114_U1_1_4 ( .A(u2_exp_tmp4_4_), .B(u2_add_114_carry[4]), .CO(
        u2_add_114_carry[5]), .S(u2_N46) );
  HA_X1 u2_add_114_U1_1_5 ( .A(n1584), .B(u2_add_114_carry[5]), .CO(
        u2_add_114_carry[6]), .S(u2_N47) );
  HA_X1 u2_add_114_U1_1_6 ( .A(n1583), .B(u2_add_114_carry[6]), .CO(
        u2_add_114_carry[7]), .S(u2_N48) );
  XOR2_X1 u2_add_112_U2 ( .A(u2_add_112_carry[7]), .B(n3400), .Z(
        u2_exp_tmp3_7_) );
  INV_X4 u2_add_112_U1 ( .A(n3408), .ZN(u2_exp_tmp3_0_) );
  HA_X1 u2_add_112_U1_1_1 ( .A(n3407), .B(n3408), .CO(u2_add_112_carry[2]), 
        .S(u2_exp_tmp3_1_) );
  HA_X1 u2_add_112_U1_1_2 ( .A(n3406), .B(u2_add_112_carry[2]), .CO(
        u2_add_112_carry[3]), .S(u2_exp_tmp3_2_) );
  HA_X1 u2_add_112_U1_1_3 ( .A(n3405), .B(u2_add_112_carry[3]), .CO(
        u2_add_112_carry[4]), .S(u2_exp_tmp3_3_) );
  HA_X1 u2_add_112_U1_1_4 ( .A(n3403), .B(u2_add_112_carry[4]), .CO(
        u2_add_112_carry[5]), .S(u2_exp_tmp3_4_) );
  HA_X1 u2_add_112_U1_1_5 ( .A(n3402), .B(u2_add_112_carry[5]), .CO(
        u2_add_112_carry[6]), .S(u2_exp_tmp3_5_) );
  HA_X1 u2_add_112_U1_1_6 ( .A(n3401), .B(u2_add_112_carry[6]), .CO(
        u2_add_112_carry[7]), .S(u2_exp_tmp3_6_) );
  AND2_X4 u2_add_109_U2 ( .A1(opb_r[23]), .A2(opa_r[23]), .ZN(u2_add_109_n2)
         );
  XOR2_X2 u2_add_109_U1 ( .A(opb_r[23]), .B(opa_r[23]), .Z(u2_N15) );
  FA_X1 u2_add_109_U1_1 ( .A(opa_r[24]), .B(opb_r[24]), .CI(u2_add_109_n2), 
        .CO(u2_add_109_carry[2]), .S(u2_N16) );
  FA_X1 u2_add_109_U1_2 ( .A(opa_r[25]), .B(opb_r[25]), .CI(
        u2_add_109_carry[2]), .CO(u2_add_109_carry[3]), .S(u2_N17) );
  FA_X1 u2_add_109_U1_3 ( .A(opa_r[26]), .B(opb_r[26]), .CI(
        u2_add_109_carry[3]), .CO(u2_add_109_carry[4]), .S(u2_N18) );
  FA_X1 u2_add_109_U1_4 ( .A(opa_r[27]), .B(opb_r[27]), .CI(
        u2_add_109_carry[4]), .CO(u2_add_109_carry[5]), .S(u2_N19) );
  FA_X1 u2_add_109_U1_5 ( .A(opa_r[28]), .B(opb_r[28]), .CI(
        u2_add_109_carry[5]), .CO(u2_add_109_carry[6]), .S(u2_N20) );
  FA_X1 u2_add_109_U1_6 ( .A(opa_r[29]), .B(opb_r[29]), .CI(
        u2_add_109_carry[6]), .CO(u2_add_109_carry[7]), .S(u2_N21) );
  FA_X1 u2_add_109_U1_7 ( .A(opa_r[30]), .B(opb_r[30]), .CI(
        u2_add_109_carry[7]), .CO(u2_N23), .S(u2_N22) );
  INV_X4 u2_sub_109_U12 ( .A(opb_r[23]), .ZN(u2_sub_109_n10) );
  INV_X4 u2_sub_109_U11 ( .A(opb_r[24]), .ZN(u2_sub_109_n9) );
  INV_X4 u2_sub_109_U10 ( .A(opb_r[25]), .ZN(u2_sub_109_n8) );
  INV_X4 u2_sub_109_U9 ( .A(opb_r[26]), .ZN(u2_sub_109_n7) );
  INV_X4 u2_sub_109_U8 ( .A(opb_r[27]), .ZN(u2_sub_109_n6) );
  INV_X4 u2_sub_109_U7 ( .A(opb_r[28]), .ZN(u2_sub_109_n5) );
  INV_X4 u2_sub_109_U6 ( .A(opb_r[29]), .ZN(u2_sub_109_n4) );
  INV_X4 u2_sub_109_U5 ( .A(opb_r[30]), .ZN(u2_sub_109_n3) );
  INV_X4 u2_sub_109_U4 ( .A(u2_sub_109_carry[8]), .ZN(u2_N14) );
  INV_X4 u2_sub_109_U3 ( .A(opa_r[23]), .ZN(u2_sub_109_n1) );
  XNOR2_X2 u2_sub_109_U2 ( .A(u2_sub_109_n10), .B(opa_r[23]), .ZN(u2_N6) );
  NAND2_X2 u2_sub_109_U1 ( .A1(opb_r[23]), .A2(u2_sub_109_n1), .ZN(
        u2_sub_109_carry[1]) );
  FA_X1 u2_sub_109_U2_1 ( .A(opa_r[24]), .B(u2_sub_109_n9), .CI(
        u2_sub_109_carry[1]), .CO(u2_sub_109_carry[2]), .S(u2_N7) );
  FA_X1 u2_sub_109_U2_2 ( .A(opa_r[25]), .B(u2_sub_109_n8), .CI(
        u2_sub_109_carry[2]), .CO(u2_sub_109_carry[3]), .S(u2_N8) );
  FA_X1 u2_sub_109_U2_3 ( .A(opa_r[26]), .B(u2_sub_109_n7), .CI(
        u2_sub_109_carry[3]), .CO(u2_sub_109_carry[4]), .S(u2_N9) );
  FA_X1 u2_sub_109_U2_4 ( .A(opa_r[27]), .B(u2_sub_109_n6), .CI(
        u2_sub_109_carry[4]), .CO(u2_sub_109_carry[5]), .S(u2_N10) );
  FA_X1 u2_sub_109_U2_5 ( .A(opa_r[28]), .B(u2_sub_109_n5), .CI(
        u2_sub_109_carry[5]), .CO(u2_sub_109_carry[6]), .S(u2_N11) );
  FA_X1 u2_sub_109_U2_6 ( .A(opa_r[29]), .B(u2_sub_109_n4), .CI(
        u2_sub_109_carry[6]), .CO(u2_sub_109_carry[7]), .S(u2_N12) );
  FA_X1 u2_sub_109_U2_7 ( .A(opa_r[30]), .B(u2_sub_109_n3), .CI(
        u2_sub_109_carry[7]), .CO(u2_sub_109_carry[8]), .S(u2_N13) );
  NAND2_X1 u1_srl_146_U168 ( .A1(n3451), .A2(u1_srl_146_n31), .ZN(
        u1_srl_146_n91) );
  AOI22_X1 u1_srl_146_U167 ( .A1(n3458), .A2(u1_srl_146_n4), .B1(n3462), .B2(
        u1_srl_146_n1), .ZN(u1_srl_146_n141) );
  OAI221_X1 u1_srl_146_U166 ( .B1(u1_srl_146_n90), .B2(u1_srl_146_n40), .C1(
        u1_srl_146_n5), .C2(u1_srl_146_n39), .A(u1_srl_146_n141), .ZN(
        u1_srl_146_n140) );
  NOR2_X1 u1_srl_146_U165 ( .A1(u1_srl_146_n14), .A2(n3452), .ZN(
        u1_srl_146_n105) );
  AOI22_X1 u1_srl_146_U164 ( .A1(u1_srl_146_n93), .A2(u1_adj_op_20_), .B1(
        u1_adj_op_17_), .B2(u1_srl_146_n2), .ZN(u1_srl_146_n139) );
  OAI221_X1 u1_srl_146_U163 ( .B1(u1_srl_146_n90), .B2(u1_srl_146_n46), .C1(
        u1_srl_146_n45), .C2(u1_srl_146_n5), .A(u1_srl_146_n139), .ZN(
        u1_srl_146_n70) );
  OAI222_X1 u1_srl_146_U162 ( .A1(u1_srl_146_n56), .A2(u1_srl_146_n5), .B1(
        u1_srl_146_n90), .B2(u1_srl_146_n41), .C1(u1_srl_146_n16), .C2(
        u1_srl_146_n42), .ZN(u1_srl_146_n69) );
  AND2_X1 u1_srl_146_U161 ( .A1(n3452), .A2(u1_srl_146_n14), .ZN(
        u1_srl_146_n113) );
  AOI22_X1 u1_srl_146_U160 ( .A1(n3463), .A2(u1_srl_146_n4), .B1(n3466), .B2(
        u1_srl_146_n94), .ZN(u1_srl_146_n138) );
  OAI221_X1 u1_srl_146_U159 ( .B1(u1_srl_146_n90), .B2(u1_srl_146_n50), .C1(
        u1_srl_146_n5), .C2(u1_srl_146_n49), .A(u1_srl_146_n138), .ZN(
        u1_srl_146_n68) );
  NOR2_X1 u1_srl_146_U158 ( .A1(n3448), .A2(n3452), .ZN(u1_srl_146_n104) );
  AOI222_X1 u1_srl_146_U157 ( .A1(u1_srl_146_n70), .A2(u1_srl_146_n105), .B1(
        u1_srl_146_n69), .B2(u1_srl_146_n113), .C1(u1_srl_146_n68), .C2(
        u1_srl_146_n104), .ZN(u1_srl_146_n114) );
  NAND2_X1 u1_srl_146_U156 ( .A1(n3452), .A2(u1_srl_146_n12), .ZN(
        u1_srl_146_n116) );
  AOI22_X1 u1_srl_146_U155 ( .A1(n3454), .A2(u1_srl_146_n93), .B1(n3457), .B2(
        u1_srl_146_n1), .ZN(u1_srl_146_n137) );
  OAI221_X1 u1_srl_146_U154 ( .B1(u1_srl_146_n90), .B2(u1_srl_146_n36), .C1(
        u1_srl_146_n5), .C2(u1_srl_146_n35), .A(u1_srl_146_n137), .ZN(
        u1_srl_146_n71) );
  AOI22_X1 u1_srl_146_U153 ( .A1(n3467), .A2(u1_srl_146_n3), .B1(n3453), .B2(
        u1_srl_146_n2), .ZN(u1_srl_146_n136) );
  OAI221_X1 u1_srl_146_U152 ( .B1(u1_srl_146_n90), .B2(u1_srl_146_n54), .C1(
        u1_srl_146_n91), .C2(u1_srl_146_n53), .A(u1_srl_146_n136), .ZN(
        u1_srl_146_n86) );
  NOR3_X1 u1_srl_146_U151 ( .A1(u1_srl_146_n55), .A2(u1_srl_146_n30), .A3(
        u1_srl_146_n58), .ZN(u1_srl_146_n135) );
  AOI221_X1 u1_srl_146_U150 ( .B1(u1_srl_146_n60), .B2(u1_srl_146_n71), .C1(
        u1_srl_146_n64), .C2(u1_srl_146_n86), .A(u1_srl_146_n135), .ZN(
        u1_srl_146_n134) );
  OAI221_X1 u1_srl_146_U149 ( .B1(u1_srl_146_n15), .B2(u1_srl_146_n57), .C1(
        u1_srl_146_n114), .C2(u1_srl_146_n12), .A(u1_srl_146_n134), .ZN(
        u1_adj_op_out_sft_0_) );
  AOI22_X1 u1_srl_146_U148 ( .A1(n3465), .A2(u1_srl_146_n4), .B1(n3468), .B2(
        u1_srl_146_n94), .ZN(u1_srl_146_n133) );
  OAI221_X1 u1_srl_146_U147 ( .B1(u1_srl_146_n90), .B2(u1_srl_146_n52), .C1(
        u1_srl_146_n91), .C2(u1_srl_146_n51), .A(u1_srl_146_n133), .ZN(
        u1_srl_146_n78) );
  AOI22_X1 u1_srl_146_U146 ( .A1(u1_adj_op_10_), .A2(u1_srl_146_n93), .B1(
        n3455), .B2(u1_srl_146_n1), .ZN(u1_srl_146_n132) );
  OAI221_X1 u1_srl_146_U145 ( .B1(u1_srl_146_n90), .B2(u1_srl_146_n34), .C1(
        u1_srl_146_n91), .C2(u1_srl_146_n33), .A(u1_srl_146_n132), .ZN(
        u1_srl_146_n99) );
  AOI22_X1 u1_srl_146_U144 ( .A1(u1_adj_op_18_), .A2(u1_srl_146_n3), .B1(n3464), .B2(u1_srl_146_n2), .ZN(u1_srl_146_n131) );
  OAI221_X1 u1_srl_146_U143 ( .B1(u1_srl_146_n90), .B2(u1_srl_146_n48), .C1(
        u1_srl_146_n91), .C2(u1_srl_146_n47), .A(u1_srl_146_n131), .ZN(
        u1_srl_146_n80) );
  NOR2_X1 u1_srl_146_U142 ( .A1(u1_srl_146_n16), .A2(u1_srl_146_n56), .ZN(
        u1_srl_146_n103) );
  AND2_X1 u1_srl_146_U141 ( .A1(u1_exp_diff_sft_4_), .A2(u1_srl_146_n104), 
        .ZN(u1_srl_146_n62) );
  AOI22_X1 u1_srl_146_U140 ( .A1(u1_srl_146_n3), .A2(u1_adj_op_22_), .B1(
        u1_adj_op_19_), .B2(u1_srl_146_n94), .ZN(u1_srl_146_n130) );
  OAI221_X1 u1_srl_146_U139 ( .B1(u1_srl_146_n90), .B2(u1_srl_146_n43), .C1(
        u1_srl_146_n91), .C2(u1_srl_146_n42), .A(u1_srl_146_n130), .ZN(
        u1_srl_146_n112) );
  AOI222_X1 u1_srl_146_U138 ( .A1(u1_srl_146_n60), .A2(u1_srl_146_n80), .B1(
        u1_srl_146_n103), .B2(u1_srl_146_n62), .C1(u1_srl_146_n64), .C2(
        u1_srl_146_n112), .ZN(u1_srl_146_n129) );
  OAI221_X1 u1_srl_146_U137 ( .B1(u1_srl_146_n20), .B2(u1_srl_146_n57), .C1(
        u1_srl_146_n21), .C2(u1_srl_146_n58), .A(u1_srl_146_n129), .ZN(
        u1_adj_op_out_sft_10_) );
  AOI22_X1 u1_srl_146_U136 ( .A1(u1_srl_146_n4), .A2(n2459), .B1(u1_adj_op_20_), .B2(u1_srl_146_n1), .ZN(u1_srl_146_n128) );
  OAI221_X1 u1_srl_146_U135 ( .B1(u1_srl_146_n90), .B2(u1_srl_146_n42), .C1(
        u1_srl_146_n41), .C2(u1_srl_146_n5), .A(u1_srl_146_n128), .ZN(
        u1_srl_146_n74) );
  AOI22_X1 u1_srl_146_U134 ( .A1(u1_srl_146_n93), .A2(u1_adj_op_19_), .B1(
        n3463), .B2(u1_srl_146_n2), .ZN(u1_srl_146_n127) );
  OAI221_X1 u1_srl_146_U133 ( .B1(u1_srl_146_n90), .B2(u1_srl_146_n47), .C1(
        u1_srl_146_n91), .C2(u1_srl_146_n46), .A(u1_srl_146_n127), .ZN(
        u1_srl_146_n75) );
  AOI22_X1 u1_srl_146_U132 ( .A1(n3464), .A2(u1_srl_146_n4), .B1(n3467), .B2(
        u1_srl_146_n94), .ZN(u1_srl_146_n126) );
  OAI221_X1 u1_srl_146_U131 ( .B1(u1_srl_146_n90), .B2(u1_srl_146_n51), .C1(
        u1_srl_146_n91), .C2(u1_srl_146_n50), .A(u1_srl_146_n126), .ZN(
        u1_srl_146_n73) );
  AOI22_X1 u1_srl_146_U130 ( .A1(n3468), .A2(u1_srl_146_n93), .B1(n3454), .B2(
        u1_srl_146_n1), .ZN(u1_srl_146_n125) );
  OAI221_X1 u1_srl_146_U129 ( .B1(u1_srl_146_n90), .B2(u1_srl_146_n33), .C1(
        u1_srl_146_n91), .C2(u1_srl_146_n54), .A(u1_srl_146_n125), .ZN(
        u1_srl_146_n76) );
  AOI22_X1 u1_srl_146_U128 ( .A1(u1_srl_146_n10), .A2(u1_srl_146_n73), .B1(
        u1_srl_146_n11), .B2(u1_srl_146_n76), .ZN(u1_srl_146_n124) );
  AOI221_X1 u1_srl_146_U127 ( .B1(u1_srl_146_n74), .B2(u1_srl_146_n64), .C1(
        u1_srl_146_n75), .C2(u1_srl_146_n60), .A(u1_srl_146_n8), .ZN(
        u1_srl_146_n123) );
  AOI22_X1 u1_srl_146_U126 ( .A1(u1_srl_146_n64), .A2(u1_srl_146_n69), .B1(
        u1_srl_146_n60), .B2(u1_srl_146_n70), .ZN(u1_srl_146_n122) );
  OAI221_X1 u1_srl_146_U125 ( .B1(u1_srl_146_n17), .B2(u1_srl_146_n57), .C1(
        u1_srl_146_n19), .C2(u1_srl_146_n58), .A(u1_srl_146_n122), .ZN(
        u1_adj_op_out_sft_12_) );
  AOI22_X1 u1_srl_146_U124 ( .A1(u1_adj_op_17_), .A2(u1_srl_146_n3), .B1(n3465), .B2(u1_srl_146_n2), .ZN(u1_srl_146_n121) );
  OAI221_X1 u1_srl_146_U123 ( .B1(u1_srl_146_n90), .B2(u1_srl_146_n49), .C1(
        u1_srl_146_n5), .C2(u1_srl_146_n48), .A(u1_srl_146_n121), .ZN(
        u1_srl_146_n61) );
  AOI22_X1 u1_srl_146_U122 ( .A1(n3466), .A2(u1_srl_146_n4), .B1(u1_adj_op_10_), .B2(u1_srl_146_n94), .ZN(u1_srl_146_n120) );
  OAI221_X1 u1_srl_146_U121 ( .B1(u1_srl_146_n90), .B2(u1_srl_146_n53), .C1(
        u1_srl_146_n5), .C2(u1_srl_146_n52), .A(u1_srl_146_n120), .ZN(
        u1_srl_146_n83) );
  OAI22_X1 u1_srl_146_U120 ( .A1(u1_srl_146_n16), .A2(u1_srl_146_n41), .B1(
        u1_srl_146_n90), .B2(u1_srl_146_n56), .ZN(u1_srl_146_n63) );
  AOI22_X1 u1_srl_146_U119 ( .A1(n3461), .A2(u1_srl_146_n93), .B1(
        u1_adj_op_18_), .B2(u1_srl_146_n1), .ZN(u1_srl_146_n119) );
  OAI221_X1 u1_srl_146_U118 ( .B1(u1_srl_146_n90), .B2(u1_srl_146_n45), .C1(
        u1_srl_146_n5), .C2(u1_srl_146_n43), .A(u1_srl_146_n119), .ZN(
        u1_srl_146_n65) );
  AOI22_X1 u1_srl_146_U117 ( .A1(u1_srl_146_n64), .A2(u1_srl_146_n63), .B1(
        u1_srl_146_n60), .B2(u1_srl_146_n65), .ZN(u1_srl_146_n118) );
  OAI221_X1 u1_srl_146_U116 ( .B1(u1_srl_146_n24), .B2(u1_srl_146_n57), .C1(
        u1_srl_146_n25), .C2(u1_srl_146_n58), .A(u1_srl_146_n118), .ZN(
        u1_adj_op_out_sft_13_) );
  MUX2_X1 u1_srl_146_U115 ( .A(u1_srl_146_n103), .B(u1_srl_146_n112), .S(
        u1_srl_146_n14), .Z(u1_srl_146_n117) );
  OAI222_X1 u1_srl_146_U114 ( .A1(u1_srl_146_n22), .A2(u1_srl_146_n57), .B1(
        u1_srl_146_n13), .B2(u1_srl_146_n116), .C1(u1_srl_146_n20), .C2(
        u1_srl_146_n58), .ZN(u1_adj_op_out_sft_14_) );
  AOI222_X1 u1_srl_146_U113 ( .A1(u1_srl_146_n75), .A2(u1_srl_146_n10), .B1(
        u1_srl_146_n74), .B2(u1_srl_146_n60), .C1(u1_srl_146_n73), .C2(
        u1_srl_146_n11), .ZN(u1_srl_146_n115) );
  NOR2_X1 u1_srl_146_U112 ( .A1(u1_exp_diff_sft_4_), .A2(u1_srl_146_n114), 
        .ZN(u1_adj_op_out_sft_16_) );
  AOI222_X1 u1_srl_146_U111 ( .A1(u1_srl_146_n65), .A2(u1_srl_146_n105), .B1(
        u1_srl_146_n63), .B2(u1_srl_146_n113), .C1(u1_srl_146_n61), .C2(
        u1_srl_146_n104), .ZN(u1_srl_146_n106) );
  NOR2_X1 u1_srl_146_U110 ( .A1(u1_exp_diff_sft_4_), .A2(u1_srl_146_n106), 
        .ZN(u1_adj_op_out_sft_17_) );
  AOI222_X1 u1_srl_146_U109 ( .A1(u1_srl_146_n112), .A2(u1_srl_146_n105), .B1(
        u1_srl_146_n103), .B2(u1_srl_146_n113), .C1(u1_srl_146_n80), .C2(
        u1_srl_146_n104), .ZN(u1_srl_146_n97) );
  NOR2_X1 u1_srl_146_U108 ( .A1(u1_exp_diff_sft_4_), .A2(u1_srl_146_n97), .ZN(
        u1_adj_op_out_sft_18_) );
  AOI22_X1 u1_srl_146_U107 ( .A1(u1_srl_146_n75), .A2(u1_srl_146_n104), .B1(
        u1_srl_146_n74), .B2(u1_srl_146_n105), .ZN(u1_srl_146_n87) );
  NOR2_X1 u1_srl_146_U106 ( .A1(u1_exp_diff_sft_4_), .A2(u1_srl_146_n87), .ZN(
        u1_adj_op_out_sft_19_) );
  AOI22_X1 u1_srl_146_U105 ( .A1(n3457), .A2(u1_srl_146_n3), .B1(n3460), .B2(
        u1_srl_146_n2), .ZN(u1_srl_146_n111) );
  OAI221_X1 u1_srl_146_U104 ( .B1(u1_srl_146_n90), .B2(u1_srl_146_n39), .C1(
        u1_srl_146_n5), .C2(u1_srl_146_n38), .A(u1_srl_146_n111), .ZN(
        u1_srl_146_n110) );
  AOI22_X1 u1_srl_146_U103 ( .A1(n3453), .A2(u1_srl_146_n4), .B1(n3456), .B2(
        u1_srl_146_n94), .ZN(u1_srl_146_n109) );
  OAI221_X1 u1_srl_146_U102 ( .B1(u1_srl_146_n90), .B2(u1_srl_146_n35), .C1(
        u1_srl_146_n5), .C2(u1_srl_146_n34), .A(u1_srl_146_n109), .ZN(
        u1_srl_146_n66) );
  OAI22_X1 u1_srl_146_U101 ( .A1(u1_srl_146_n30), .A2(u1_srl_146_n44), .B1(
        u1_srl_146_n5), .B2(u1_srl_146_n55), .ZN(u1_srl_146_n108) );
  AOI222_X1 u1_srl_146_U100 ( .A1(u1_srl_146_n60), .A2(u1_srl_146_n66), .B1(
        u1_srl_146_n11), .B2(u1_srl_146_n108), .C1(u1_srl_146_n64), .C2(
        u1_srl_146_n83), .ZN(u1_srl_146_n107) );
  OAI221_X1 u1_srl_146_U99 ( .B1(u1_srl_146_n26), .B2(u1_srl_146_n57), .C1(
        u1_srl_146_n106), .C2(u1_srl_146_n12), .A(u1_srl_146_n107), .ZN(
        u1_adj_op_out_sft_1_) );
  AOI22_X1 u1_srl_146_U98 ( .A1(u1_srl_146_n70), .A2(u1_srl_146_n104), .B1(
        u1_srl_146_n69), .B2(u1_srl_146_n105), .ZN(u1_srl_146_n84) );
  NOR2_X1 u1_srl_146_U97 ( .A1(u1_exp_diff_sft_4_), .A2(u1_srl_146_n84), .ZN(
        u1_adj_op_out_sft_20_) );
  AOI22_X1 u1_srl_146_U96 ( .A1(u1_srl_146_n65), .A2(u1_srl_146_n104), .B1(
        u1_srl_146_n63), .B2(u1_srl_146_n105), .ZN(u1_srl_146_n81) );
  NOR2_X1 u1_srl_146_U95 ( .A1(u1_exp_diff_sft_4_), .A2(u1_srl_146_n81), .ZN(
        u1_adj_op_out_sft_21_) );
  NOR3_X1 u1_srl_146_U94 ( .A1(u1_srl_146_n13), .A2(u1_exp_diff_sft_4_), .A3(
        n3452), .ZN(u1_adj_op_out_sft_22_) );
  AND2_X1 u1_srl_146_U93 ( .A1(u1_srl_146_n74), .A2(u1_srl_146_n11), .ZN(
        u1_adj_op_out_sft_23_) );
  AND2_X1 u1_srl_146_U92 ( .A1(u1_srl_146_n69), .A2(u1_srl_146_n11), .ZN(
        u1_adj_op_out_sft_24_) );
  AND2_X1 u1_srl_146_U91 ( .A1(u1_srl_146_n63), .A2(u1_srl_146_n11), .ZN(
        u1_adj_op_out_sft_25_) );
  AND2_X1 u1_srl_146_U90 ( .A1(u1_srl_146_n11), .A2(u1_srl_146_n103), .ZN(
        u1_adj_op_out_sft_26_) );
  AOI22_X1 u1_srl_146_U89 ( .A1(n3456), .A2(u1_srl_146_n93), .B1(n3459), .B2(
        u1_srl_146_n1), .ZN(u1_srl_146_n102) );
  OAI221_X1 u1_srl_146_U88 ( .B1(u1_srl_146_n90), .B2(u1_srl_146_n38), .C1(
        u1_srl_146_n5), .C2(u1_srl_146_n37), .A(u1_srl_146_n102), .ZN(
        u1_srl_146_n101) );
  OAI222_X1 u1_srl_146_U87 ( .A1(u1_srl_146_n5), .A2(u1_srl_146_n44), .B1(
        u1_srl_146_n90), .B2(u1_srl_146_n55), .C1(u1_srl_146_n30), .C2(
        u1_srl_146_n40), .ZN(u1_srl_146_n100) );
  AOI222_X1 u1_srl_146_U86 ( .A1(u1_srl_146_n60), .A2(u1_srl_146_n99), .B1(
        u1_srl_146_n11), .B2(u1_srl_146_n100), .C1(u1_srl_146_n64), .C2(
        u1_srl_146_n78), .ZN(u1_srl_146_n98) );
  OAI221_X1 u1_srl_146_U85 ( .B1(u1_srl_146_n28), .B2(u1_srl_146_n57), .C1(
        u1_srl_146_n97), .C2(u1_srl_146_n12), .A(u1_srl_146_n98), .ZN(
        u1_adj_op_out_sft_2_) );
  AOI22_X1 u1_srl_146_U84 ( .A1(n3455), .A2(u1_srl_146_n3), .B1(n3458), .B2(
        u1_srl_146_n2), .ZN(u1_srl_146_n96) );
  OAI221_X1 u1_srl_146_U83 ( .B1(u1_srl_146_n90), .B2(u1_srl_146_n37), .C1(
        u1_srl_146_n5), .C2(u1_srl_146_n36), .A(u1_srl_146_n96), .ZN(
        u1_srl_146_n95) );
  AOI22_X1 u1_srl_146_U82 ( .A1(n3459), .A2(u1_srl_146_n4), .B1(n3469), .B2(
        u1_srl_146_n94), .ZN(u1_srl_146_n92) );
  OAI221_X1 u1_srl_146_U81 ( .B1(u1_srl_146_n90), .B2(u1_srl_146_n44), .C1(
        u1_srl_146_n91), .C2(u1_srl_146_n40), .A(u1_srl_146_n92), .ZN(
        u1_srl_146_n89) );
  AOI222_X1 u1_srl_146_U80 ( .A1(u1_srl_146_n60), .A2(u1_srl_146_n76), .B1(
        u1_srl_146_n11), .B2(u1_srl_146_n89), .C1(u1_srl_146_n64), .C2(
        u1_srl_146_n73), .ZN(u1_srl_146_n88) );
  OAI221_X1 u1_srl_146_U79 ( .B1(u1_srl_146_n29), .B2(u1_srl_146_n57), .C1(
        u1_srl_146_n87), .C2(u1_srl_146_n12), .A(u1_srl_146_n88), .ZN(
        u1_adj_op_out_sft_3_) );
  AOI222_X1 u1_srl_146_U78 ( .A1(u1_srl_146_n10), .A2(u1_srl_146_n71), .B1(
        u1_srl_146_n64), .B2(u1_srl_146_n68), .C1(u1_srl_146_n60), .C2(
        u1_srl_146_n86), .ZN(u1_srl_146_n85) );
  OAI221_X1 u1_srl_146_U77 ( .B1(u1_srl_146_n15), .B2(u1_srl_146_n58), .C1(
        u1_srl_146_n84), .C2(u1_srl_146_n12), .A(u1_srl_146_n85), .ZN(
        u1_adj_op_out_sft_4_) );
  AOI222_X1 u1_srl_146_U76 ( .A1(u1_srl_146_n10), .A2(u1_srl_146_n66), .B1(
        u1_srl_146_n64), .B2(u1_srl_146_n61), .C1(u1_srl_146_n60), .C2(
        u1_srl_146_n83), .ZN(u1_srl_146_n82) );
  OAI221_X1 u1_srl_146_U75 ( .B1(u1_srl_146_n26), .B2(u1_srl_146_n58), .C1(
        u1_srl_146_n81), .C2(u1_srl_146_n12), .A(u1_srl_146_n82), .ZN(
        u1_adj_op_out_sft_5_) );
  NOR2_X1 u1_srl_146_U74 ( .A1(n3452), .A2(u1_srl_146_n13), .ZN(u1_srl_146_n79) );
  AOI222_X1 u1_srl_146_U73 ( .A1(u1_srl_146_n60), .A2(u1_srl_146_n78), .B1(
        u1_srl_146_n79), .B2(u1_exp_diff_sft_4_), .C1(u1_srl_146_n64), .C2(
        u1_srl_146_n80), .ZN(u1_srl_146_n77) );
  OAI221_X1 u1_srl_146_U72 ( .B1(u1_srl_146_n21), .B2(u1_srl_146_n57), .C1(
        u1_srl_146_n28), .C2(u1_srl_146_n58), .A(u1_srl_146_n77), .ZN(
        u1_adj_op_out_sft_6_) );
  AOI222_X1 u1_srl_146_U71 ( .A1(u1_srl_146_n60), .A2(u1_srl_146_n73), .B1(
        u1_srl_146_n62), .B2(u1_srl_146_n74), .C1(u1_srl_146_n64), .C2(
        u1_srl_146_n75), .ZN(u1_srl_146_n72) );
  OAI221_X1 u1_srl_146_U70 ( .B1(u1_srl_146_n23), .B2(u1_srl_146_n57), .C1(
        u1_srl_146_n29), .C2(u1_srl_146_n58), .A(u1_srl_146_n72), .ZN(
        u1_adj_op_out_sft_7_) );
  AOI222_X1 u1_srl_146_U69 ( .A1(u1_srl_146_n60), .A2(u1_srl_146_n68), .B1(
        u1_srl_146_n62), .B2(u1_srl_146_n69), .C1(u1_srl_146_n64), .C2(
        u1_srl_146_n70), .ZN(u1_srl_146_n67) );
  OAI221_X1 u1_srl_146_U68 ( .B1(u1_srl_146_n19), .B2(u1_srl_146_n57), .C1(
        u1_srl_146_n18), .C2(u1_srl_146_n58), .A(u1_srl_146_n67), .ZN(
        u1_adj_op_out_sft_8_) );
  AOI222_X1 u1_srl_146_U67 ( .A1(u1_srl_146_n60), .A2(u1_srl_146_n61), .B1(
        u1_srl_146_n62), .B2(u1_srl_146_n63), .C1(u1_srl_146_n64), .C2(
        u1_srl_146_n65), .ZN(u1_srl_146_n59) );
  OAI221_X1 u1_srl_146_U66 ( .B1(u1_srl_146_n25), .B2(u1_srl_146_n57), .C1(
        u1_srl_146_n27), .C2(u1_srl_146_n58), .A(u1_srl_146_n59), .ZN(
        u1_adj_op_out_sft_9_) );
  INV_X4 u1_srl_146_U65 ( .A(n2459), .ZN(u1_srl_146_n56) );
  INV_X4 u1_srl_146_U64 ( .A(n3469), .ZN(u1_srl_146_n55) );
  INV_X4 u1_srl_146_U63 ( .A(u1_adj_op_10_), .ZN(u1_srl_146_n54) );
  INV_X4 u1_srl_146_U62 ( .A(n3468), .ZN(u1_srl_146_n53) );
  INV_X4 u1_srl_146_U61 ( .A(n3467), .ZN(u1_srl_146_n52) );
  INV_X4 u1_srl_146_U60 ( .A(n3466), .ZN(u1_srl_146_n51) );
  INV_X4 u1_srl_146_U59 ( .A(n3465), .ZN(u1_srl_146_n50) );
  INV_X4 u1_srl_146_U58 ( .A(n3464), .ZN(u1_srl_146_n49) );
  INV_X4 u1_srl_146_U57 ( .A(n3463), .ZN(u1_srl_146_n48) );
  INV_X4 u1_srl_146_U56 ( .A(u1_adj_op_17_), .ZN(u1_srl_146_n47) );
  INV_X4 u1_srl_146_U55 ( .A(u1_adj_op_18_), .ZN(u1_srl_146_n46) );
  INV_X4 u1_srl_146_U54 ( .A(u1_adj_op_19_), .ZN(u1_srl_146_n45) );
  INV_X4 u1_srl_146_U53 ( .A(n3462), .ZN(u1_srl_146_n44) );
  INV_X4 u1_srl_146_U52 ( .A(u1_adj_op_20_), .ZN(u1_srl_146_n43) );
  INV_X4 u1_srl_146_U51 ( .A(n3461), .ZN(u1_srl_146_n42) );
  INV_X4 u1_srl_146_U50 ( .A(u1_adj_op_22_), .ZN(u1_srl_146_n41) );
  INV_X4 u1_srl_146_U49 ( .A(n3460), .ZN(u1_srl_146_n40) );
  INV_X4 u1_srl_146_U48 ( .A(n3459), .ZN(u1_srl_146_n39) );
  INV_X4 u1_srl_146_U47 ( .A(n3458), .ZN(u1_srl_146_n38) );
  INV_X4 u1_srl_146_U46 ( .A(n3457), .ZN(u1_srl_146_n37) );
  INV_X4 u1_srl_146_U45 ( .A(n3456), .ZN(u1_srl_146_n36) );
  INV_X4 u1_srl_146_U44 ( .A(n3455), .ZN(u1_srl_146_n35) );
  INV_X4 u1_srl_146_U43 ( .A(n3454), .ZN(u1_srl_146_n34) );
  INV_X4 u1_srl_146_U42 ( .A(n3453), .ZN(u1_srl_146_n33) );
  INV_X4 u1_srl_146_U41 ( .A(n3451), .ZN(u1_srl_146_n32) );
  INV_X4 u1_srl_146_U40 ( .A(n3450), .ZN(u1_srl_146_n31) );
  INV_X4 u1_srl_146_U39 ( .A(u1_srl_146_n3), .ZN(u1_srl_146_n30) );
  INV_X4 u1_srl_146_U38 ( .A(u1_srl_146_n95), .ZN(u1_srl_146_n29) );
  INV_X4 u1_srl_146_U37 ( .A(u1_srl_146_n101), .ZN(u1_srl_146_n28) );
  INV_X4 u1_srl_146_U36 ( .A(u1_srl_146_n66), .ZN(u1_srl_146_n27) );
  INV_X4 u1_srl_146_U35 ( .A(u1_srl_146_n110), .ZN(u1_srl_146_n26) );
  INV_X4 u1_srl_146_U34 ( .A(u1_srl_146_n83), .ZN(u1_srl_146_n25) );
  INV_X4 u1_srl_146_U33 ( .A(u1_srl_146_n61), .ZN(u1_srl_146_n24) );
  INV_X4 u1_srl_146_U32 ( .A(u1_srl_146_n76), .ZN(u1_srl_146_n23) );
  INV_X4 u1_srl_146_U31 ( .A(u1_srl_146_n80), .ZN(u1_srl_146_n22) );
  INV_X4 u1_srl_146_U30 ( .A(u1_srl_146_n99), .ZN(u1_srl_146_n21) );
  INV_X4 u1_srl_146_U29 ( .A(u1_srl_146_n78), .ZN(u1_srl_146_n20) );
  INV_X4 u1_srl_146_U28 ( .A(u1_srl_146_n86), .ZN(u1_srl_146_n19) );
  INV_X4 u1_srl_146_U27 ( .A(u1_srl_146_n71), .ZN(u1_srl_146_n18) );
  INV_X4 u1_srl_146_U26 ( .A(u1_srl_146_n68), .ZN(u1_srl_146_n17) );
  INV_X4 u1_srl_146_U25 ( .A(u1_srl_146_n1), .ZN(u1_srl_146_n16) );
  INV_X4 u1_srl_146_U24 ( .A(u1_srl_146_n140), .ZN(u1_srl_146_n15) );
  INV_X4 u1_srl_146_U23 ( .A(n3448), .ZN(u1_srl_146_n14) );
  INV_X4 u1_srl_146_U22 ( .A(u1_srl_146_n117), .ZN(u1_srl_146_n13) );
  INV_X4 u1_srl_146_U21 ( .A(u1_srl_146_n57), .ZN(u1_srl_146_n10) );
  INV_X4 u1_srl_146_U20 ( .A(u1_srl_146_n115), .ZN(u1_adj_op_out_sft_15_) );
  INV_X4 u1_srl_146_U19 ( .A(u1_srl_146_n124), .ZN(u1_srl_146_n8) );
  INV_X4 u1_srl_146_U18 ( .A(u1_srl_146_n123), .ZN(u1_adj_op_out_sft_11_) );
  INV_X4 u1_srl_146_U17 ( .A(u1_srl_146_n6), .ZN(u1_srl_146_n5) );
  INV_X4 u1_srl_146_U16 ( .A(u1_srl_146_n91), .ZN(u1_srl_146_n6) );
  NAND2_X2 u1_srl_146_U15 ( .A1(n3450), .A2(u1_srl_146_n32), .ZN(
        u1_srl_146_n90) );
  INV_X4 u1_srl_146_U14 ( .A(u1_srl_146_n58), .ZN(u1_srl_146_n11) );
  NAND2_X2 u1_srl_146_U13 ( .A1(u1_srl_146_n105), .A2(u1_srl_146_n12), .ZN(
        u1_srl_146_n57) );
  INV_X4 u1_srl_146_U12 ( .A(u1_exp_diff_sft_4_), .ZN(u1_srl_146_n12) );
  NOR2_X2 u1_srl_146_U11 ( .A1(u1_srl_146_n14), .A2(u1_srl_146_n116), .ZN(
        u1_srl_146_n64) );
  NOR2_X2 u1_srl_146_U10 ( .A1(u1_srl_146_n116), .A2(n3448), .ZN(
        u1_srl_146_n60) );
  NOR2_X2 u1_srl_146_U9 ( .A1(u1_srl_146_n32), .A2(u1_srl_146_n31), .ZN(
        u1_srl_146_n4) );
  NOR2_X2 u1_srl_146_U8 ( .A1(n3450), .A2(n3451), .ZN(u1_srl_146_n94) );
  NAND2_X2 u1_srl_146_U7 ( .A1(u1_srl_146_n104), .A2(u1_srl_146_n12), .ZN(
        u1_srl_146_n58) );
  NOR2_X2 u1_srl_146_U6 ( .A1(n3450), .A2(n3451), .ZN(u1_srl_146_n2) );
  NOR2_X2 u1_srl_146_U5 ( .A1(u1_srl_146_n32), .A2(u1_srl_146_n31), .ZN(
        u1_srl_146_n3) );
  NOR2_X2 u1_srl_146_U4 ( .A1(n3450), .A2(n3451), .ZN(u1_srl_146_n1) );
  NOR2_X2 u1_srl_146_U3 ( .A1(u1_srl_146_n32), .A2(u1_srl_146_n31), .ZN(
        u1_srl_146_n93) );
  INV_X4 sub_1_root_u1_sub_128_aco_U9 ( .A(n3479), .ZN(
        sub_1_root_u1_sub_128_aco_n9) );
  INV_X4 sub_1_root_u1_sub_128_aco_U8 ( .A(u1_exp_small[0]), .ZN(
        sub_1_root_u1_sub_128_aco_n8) );
  INV_X4 sub_1_root_u1_sub_128_aco_U7 ( .A(u1_exp_small[1]), .ZN(
        sub_1_root_u1_sub_128_aco_n7) );
  INV_X4 sub_1_root_u1_sub_128_aco_U6 ( .A(u1_exp_small[2]), .ZN(
        sub_1_root_u1_sub_128_aco_n6) );
  INV_X4 sub_1_root_u1_sub_128_aco_U5 ( .A(u1_exp_small[3]), .ZN(
        sub_1_root_u1_sub_128_aco_n5) );
  INV_X4 sub_1_root_u1_sub_128_aco_U4 ( .A(u1_exp_small[4]), .ZN(
        sub_1_root_u1_sub_128_aco_n4) );
  INV_X4 sub_1_root_u1_sub_128_aco_U3 ( .A(u1_exp_small[5]), .ZN(
        sub_1_root_u1_sub_128_aco_n3) );
  INV_X4 sub_1_root_u1_sub_128_aco_U2 ( .A(u1_exp_small[6]), .ZN(
        sub_1_root_u1_sub_128_aco_n2) );
  INV_X4 sub_1_root_u1_sub_128_aco_U1 ( .A(u1_exp_small[7]), .ZN(
        sub_1_root_u1_sub_128_aco_n1) );
  FA_X1 sub_1_root_u1_sub_128_aco_U2_0 ( .A(n3477), .B(
        sub_1_root_u1_sub_128_aco_n8), .CI(sub_1_root_u1_sub_128_aco_n9), .CO(
        sub_1_root_u1_sub_128_aco_carry[1]), .S(u1_exp_diff2[0]) );
  FA_X1 sub_1_root_u1_sub_128_aco_U2_1 ( .A(n3476), .B(
        sub_1_root_u1_sub_128_aco_n7), .CI(sub_1_root_u1_sub_128_aco_carry[1]), 
        .CO(sub_1_root_u1_sub_128_aco_carry[2]), .S(u1_exp_diff2[1]) );
  FA_X1 sub_1_root_u1_sub_128_aco_U2_2 ( .A(n3475), .B(
        sub_1_root_u1_sub_128_aco_n6), .CI(sub_1_root_u1_sub_128_aco_carry[2]), 
        .CO(sub_1_root_u1_sub_128_aco_carry[3]), .S(u1_exp_diff2[2]) );
  FA_X1 sub_1_root_u1_sub_128_aco_U2_3 ( .A(n3474), .B(
        sub_1_root_u1_sub_128_aco_n5), .CI(sub_1_root_u1_sub_128_aco_carry[3]), 
        .CO(sub_1_root_u1_sub_128_aco_carry[4]), .S(u1_exp_diff2[3]) );
  FA_X1 sub_1_root_u1_sub_128_aco_U2_4 ( .A(n3473), .B(
        sub_1_root_u1_sub_128_aco_n4), .CI(sub_1_root_u1_sub_128_aco_carry[4]), 
        .CO(sub_1_root_u1_sub_128_aco_carry[5]), .S(u1_exp_diff2[4]) );
  FA_X1 sub_1_root_u1_sub_128_aco_U2_5 ( .A(n3472), .B(
        sub_1_root_u1_sub_128_aco_n3), .CI(sub_1_root_u1_sub_128_aco_carry[5]), 
        .CO(sub_1_root_u1_sub_128_aco_carry[6]), .S(u1_exp_diff2[5]) );
  FA_X1 sub_1_root_u1_sub_128_aco_U2_6 ( .A(n3471), .B(
        sub_1_root_u1_sub_128_aco_n2), .CI(sub_1_root_u1_sub_128_aco_carry[6]), 
        .CO(sub_1_root_u1_sub_128_aco_carry[7]), .S(u1_exp_diff2[6]) );
  FA_X1 sub_1_root_u1_sub_128_aco_U2_7 ( .A(n3470), .B(
        sub_1_root_u1_sub_128_aco_n1), .CI(sub_1_root_u1_sub_128_aco_carry[7]), 
        .S(u1_exp_diff2[7]) );
  INV_X4 sub_434_3_U84 ( .A(N227), .ZN(sub_434_3_n84) );
  INV_X4 sub_434_3_U83 ( .A(opa_r1[1]), .ZN(sub_434_3_n83) );
  INV_X4 sub_434_3_U82 ( .A(opa_r1[2]), .ZN(sub_434_3_n82) );
  INV_X4 sub_434_3_U81 ( .A(opa_r1[3]), .ZN(sub_434_3_n81) );
  INV_X4 sub_434_3_U80 ( .A(opa_r1[4]), .ZN(sub_434_3_n80) );
  INV_X4 sub_434_3_U79 ( .A(opa_r1[5]), .ZN(sub_434_3_n79) );
  INV_X4 sub_434_3_U78 ( .A(opa_r1[6]), .ZN(sub_434_3_n78) );
  INV_X4 sub_434_3_U77 ( .A(opa_r1[7]), .ZN(sub_434_3_n77) );
  INV_X4 sub_434_3_U76 ( .A(opa_r1[8]), .ZN(sub_434_3_n76) );
  INV_X4 sub_434_3_U75 ( .A(opa_r1[9]), .ZN(sub_434_3_n75) );
  INV_X4 sub_434_3_U74 ( .A(opa_r1[10]), .ZN(sub_434_3_n74) );
  INV_X4 sub_434_3_U73 ( .A(opa_r1[11]), .ZN(sub_434_3_n73) );
  INV_X4 sub_434_3_U72 ( .A(opa_r1[12]), .ZN(sub_434_3_n72) );
  INV_X4 sub_434_3_U71 ( .A(opa_r1[13]), .ZN(sub_434_3_n71) );
  INV_X4 sub_434_3_U70 ( .A(opa_r1[14]), .ZN(sub_434_3_n70) );
  INV_X4 sub_434_3_U69 ( .A(opa_r1[15]), .ZN(sub_434_3_n69) );
  INV_X4 sub_434_3_U68 ( .A(opa_r1[16]), .ZN(sub_434_3_n68) );
  INV_X4 sub_434_3_U67 ( .A(opa_r1[17]), .ZN(sub_434_3_n67) );
  INV_X4 sub_434_3_U66 ( .A(opa_r1[18]), .ZN(sub_434_3_n66) );
  INV_X4 sub_434_3_U65 ( .A(opa_r1[19]), .ZN(sub_434_3_n65) );
  INV_X4 sub_434_3_U64 ( .A(opa_r1[20]), .ZN(sub_434_3_n64) );
  INV_X4 sub_434_3_U63 ( .A(opa_r1[21]), .ZN(sub_434_3_n63) );
  INV_X4 sub_434_3_U62 ( .A(opa_r1[22]), .ZN(sub_434_3_n62) );
  INV_X4 sub_434_3_U61 ( .A(opa_r1[23]), .ZN(sub_434_3_n61) );
  INV_X4 sub_434_3_U60 ( .A(opa_r1[24]), .ZN(sub_434_3_n60) );
  INV_X4 sub_434_3_U59 ( .A(opa_r1[25]), .ZN(sub_434_3_n59) );
  INV_X4 sub_434_3_U58 ( .A(opa_r1[26]), .ZN(sub_434_3_n58) );
  INV_X4 sub_434_3_U57 ( .A(opa_r1[27]), .ZN(sub_434_3_n57) );
  INV_X4 sub_434_3_U56 ( .A(opa_r1[28]), .ZN(sub_434_3_n56) );
  XOR2_X2 sub_434_3_U55 ( .A(sub_434_3_n71), .B(sub_434_3_n25), .Z(N310) );
  XOR2_X2 sub_434_3_U54 ( .A(sub_434_3_n72), .B(sub_434_3_n19), .Z(N309) );
  XOR2_X2 sub_434_3_U53 ( .A(sub_434_3_n73), .B(sub_434_3_n17), .Z(N308) );
  XOR2_X2 sub_434_3_U52 ( .A(sub_434_3_n74), .B(sub_434_3_n20), .Z(N307) );
  XOR2_X2 sub_434_3_U51 ( .A(sub_434_3_n75), .B(sub_434_3_n18), .Z(N306) );
  XOR2_X2 sub_434_3_U50 ( .A(sub_434_3_n81), .B(sub_434_3_n14), .Z(N300) );
  XOR2_X2 sub_434_3_U49 ( .A(sub_434_3_n82), .B(sub_434_3_n24), .Z(N299) );
  XOR2_X2 sub_434_3_U48 ( .A(sub_434_3_n76), .B(sub_434_3_n21), .Z(N305) );
  XOR2_X2 sub_434_3_U47 ( .A(sub_434_3_n77), .B(sub_434_3_n12), .Z(N304) );
  XOR2_X2 sub_434_3_U46 ( .A(sub_434_3_n78), .B(sub_434_3_n22), .Z(N303) );
  XOR2_X2 sub_434_3_U45 ( .A(sub_434_3_n79), .B(sub_434_3_n13), .Z(N302) );
  XOR2_X2 sub_434_3_U44 ( .A(sub_434_3_n80), .B(sub_434_3_n23), .Z(N301) );
  XOR2_X2 sub_434_3_U43 ( .A(sub_434_3_n83), .B(sub_434_3_n84), .Z(N298) );
  AND2_X4 sub_434_3_U42 ( .A1(sub_434_3_n57), .A2(sub_434_3_n28), .ZN(
        sub_434_3_n42) );
  AND2_X4 sub_434_3_U41 ( .A1(sub_434_3_n61), .A2(sub_434_3_n26), .ZN(
        sub_434_3_n41) );
  AND2_X4 sub_434_3_U40 ( .A1(sub_434_3_n59), .A2(sub_434_3_n29), .ZN(
        sub_434_3_n40) );
  AND2_X4 sub_434_3_U39 ( .A1(sub_434_3_n71), .A2(sub_434_3_n25), .ZN(
        sub_434_3_n39) );
  AND2_X4 sub_434_3_U38 ( .A1(sub_434_3_n69), .A2(sub_434_3_n16), .ZN(
        sub_434_3_n38) );
  AND2_X4 sub_434_3_U37 ( .A1(sub_434_3_n67), .A2(sub_434_3_n15), .ZN(
        sub_434_3_n37) );
  AND2_X4 sub_434_3_U36 ( .A1(sub_434_3_n65), .A2(sub_434_3_n30), .ZN(
        sub_434_3_n36) );
  AND2_X4 sub_434_3_U35 ( .A1(sub_434_3_n63), .A2(sub_434_3_n27), .ZN(
        sub_434_3_n35) );
  XOR2_X2 sub_434_3_U34 ( .A(sub_434_3_n69), .B(sub_434_3_n16), .Z(N312) );
  XOR2_X2 sub_434_3_U33 ( .A(sub_434_3_n70), .B(sub_434_3_n39), .Z(N311) );
  XOR2_X2 sub_434_3_U32 ( .A(sub_434_3_n67), .B(sub_434_3_n15), .Z(N314) );
  XOR2_X2 sub_434_3_U31 ( .A(sub_434_3_n68), .B(sub_434_3_n38), .Z(N313) );
  AND2_X4 sub_434_3_U30 ( .A1(sub_434_3_n66), .A2(sub_434_3_n37), .ZN(
        sub_434_3_n30) );
  AND2_X4 sub_434_3_U29 ( .A1(sub_434_3_n60), .A2(sub_434_3_n41), .ZN(
        sub_434_3_n29) );
  AND2_X4 sub_434_3_U28 ( .A1(sub_434_3_n58), .A2(sub_434_3_n40), .ZN(
        sub_434_3_n28) );
  AND2_X4 sub_434_3_U27 ( .A1(sub_434_3_n64), .A2(sub_434_3_n36), .ZN(
        sub_434_3_n27) );
  AND2_X4 sub_434_3_U26 ( .A1(sub_434_3_n62), .A2(sub_434_3_n35), .ZN(
        sub_434_3_n26) );
  AND2_X4 sub_434_3_U25 ( .A1(sub_434_3_n72), .A2(sub_434_3_n19), .ZN(
        sub_434_3_n25) );
  AND2_X4 sub_434_3_U24 ( .A1(sub_434_3_n83), .A2(sub_434_3_n84), .ZN(
        sub_434_3_n24) );
  AND2_X4 sub_434_3_U23 ( .A1(sub_434_3_n81), .A2(sub_434_3_n14), .ZN(
        sub_434_3_n23) );
  AND2_X4 sub_434_3_U22 ( .A1(sub_434_3_n79), .A2(sub_434_3_n13), .ZN(
        sub_434_3_n22) );
  AND2_X4 sub_434_3_U21 ( .A1(sub_434_3_n77), .A2(sub_434_3_n12), .ZN(
        sub_434_3_n21) );
  AND2_X4 sub_434_3_U20 ( .A1(sub_434_3_n75), .A2(sub_434_3_n18), .ZN(
        sub_434_3_n20) );
  AND2_X4 sub_434_3_U19 ( .A1(sub_434_3_n73), .A2(sub_434_3_n17), .ZN(
        sub_434_3_n19) );
  AND2_X4 sub_434_3_U18 ( .A1(sub_434_3_n76), .A2(sub_434_3_n21), .ZN(
        sub_434_3_n18) );
  AND2_X4 sub_434_3_U17 ( .A1(sub_434_3_n74), .A2(sub_434_3_n20), .ZN(
        sub_434_3_n17) );
  AND2_X4 sub_434_3_U16 ( .A1(sub_434_3_n70), .A2(sub_434_3_n39), .ZN(
        sub_434_3_n16) );
  AND2_X4 sub_434_3_U15 ( .A1(sub_434_3_n68), .A2(sub_434_3_n38), .ZN(
        sub_434_3_n15) );
  AND2_X4 sub_434_3_U14 ( .A1(sub_434_3_n82), .A2(sub_434_3_n24), .ZN(
        sub_434_3_n14) );
  AND2_X4 sub_434_3_U13 ( .A1(sub_434_3_n80), .A2(sub_434_3_n23), .ZN(
        sub_434_3_n13) );
  AND2_X4 sub_434_3_U12 ( .A1(sub_434_3_n78), .A2(sub_434_3_n22), .ZN(
        sub_434_3_n12) );
  XOR2_X2 sub_434_3_U11 ( .A(sub_434_3_n58), .B(sub_434_3_n40), .Z(N323) );
  XOR2_X2 sub_434_3_U10 ( .A(sub_434_3_n59), .B(sub_434_3_n29), .Z(N322) );
  XOR2_X2 sub_434_3_U9 ( .A(sub_434_3_n61), .B(sub_434_3_n26), .Z(N320) );
  XOR2_X2 sub_434_3_U8 ( .A(sub_434_3_n64), .B(sub_434_3_n36), .Z(N317) );
  XOR2_X2 sub_434_3_U7 ( .A(sub_434_3_n65), .B(sub_434_3_n30), .Z(N316) );
  XOR2_X2 sub_434_3_U6 ( .A(sub_434_3_n60), .B(sub_434_3_n41), .Z(N321) );
  XOR2_X2 sub_434_3_U5 ( .A(sub_434_3_n62), .B(sub_434_3_n35), .Z(N319) );
  XOR2_X2 sub_434_3_U4 ( .A(sub_434_3_n63), .B(sub_434_3_n27), .Z(N318) );
  XOR2_X2 sub_434_3_U3 ( .A(sub_434_3_n66), .B(sub_434_3_n37), .Z(N315) );
  XOR2_X2 sub_434_3_U2 ( .A(sub_434_3_n56), .B(sub_434_3_n42), .Z(N325) );
  XOR2_X2 sub_434_3_U1 ( .A(sub_434_3_n57), .B(sub_434_3_n28), .Z(N324) );
  INV_X4 sub_434_b0_U70 ( .A(N227), .ZN(sub_434_b0_n70) );
  INV_X4 sub_434_b0_U69 ( .A(opa_r1[1]), .ZN(sub_434_b0_n69) );
  INV_X4 sub_434_b0_U68 ( .A(opa_r1[2]), .ZN(sub_434_b0_n68) );
  INV_X4 sub_434_b0_U67 ( .A(opa_r1[3]), .ZN(sub_434_b0_n67) );
  INV_X4 sub_434_b0_U66 ( .A(opa_r1[4]), .ZN(sub_434_b0_n66) );
  INV_X4 sub_434_b0_U65 ( .A(opa_r1[5]), .ZN(sub_434_b0_n65) );
  INV_X4 sub_434_b0_U64 ( .A(opa_r1[6]), .ZN(sub_434_b0_n64) );
  INV_X4 sub_434_b0_U63 ( .A(opa_r1[7]), .ZN(sub_434_b0_n63) );
  INV_X4 sub_434_b0_U62 ( .A(opa_r1[8]), .ZN(sub_434_b0_n62) );
  INV_X4 sub_434_b0_U61 ( .A(opa_r1[9]), .ZN(sub_434_b0_n61) );
  INV_X4 sub_434_b0_U60 ( .A(opa_r1[10]), .ZN(sub_434_b0_n60) );
  INV_X4 sub_434_b0_U59 ( .A(opa_r1[11]), .ZN(sub_434_b0_n59) );
  INV_X4 sub_434_b0_U58 ( .A(opa_r1[12]), .ZN(sub_434_b0_n58) );
  INV_X4 sub_434_b0_U57 ( .A(opa_r1[13]), .ZN(sub_434_b0_n57) );
  INV_X4 sub_434_b0_U56 ( .A(opa_r1[14]), .ZN(sub_434_b0_n56) );
  INV_X4 sub_434_b0_U55 ( .A(opa_r1[15]), .ZN(sub_434_b0_n55) );
  INV_X4 sub_434_b0_U54 ( .A(opa_r1[16]), .ZN(sub_434_b0_n54) );
  INV_X4 sub_434_b0_U53 ( .A(opa_r1[17]), .ZN(sub_434_b0_n53) );
  INV_X4 sub_434_b0_U52 ( .A(opa_r1[18]), .ZN(sub_434_b0_n52) );
  INV_X4 sub_434_b0_U51 ( .A(opa_r1[19]), .ZN(sub_434_b0_n51) );
  INV_X4 sub_434_b0_U50 ( .A(opa_r1[20]), .ZN(sub_434_b0_n50) );
  INV_X4 sub_434_b0_U49 ( .A(opa_r1[21]), .ZN(sub_434_b0_n49) );
  INV_X4 sub_434_b0_U48 ( .A(opa_r1[22]), .ZN(sub_434_b0_n48) );
  INV_X4 sub_434_b0_U47 ( .A(N224), .ZN(sub_434_b0_n47) );
  NAND2_X2 sub_434_b0_U46 ( .A1(sub_434_b0_n47), .A2(sub_434_b0_n1), .ZN(N251)
         );
  XOR2_X2 sub_434_b0_U45 ( .A(sub_434_b0_n57), .B(sub_434_b0_n4), .Z(N240) );
  XOR2_X2 sub_434_b0_U44 ( .A(sub_434_b0_n58), .B(sub_434_b0_n20), .Z(N239) );
  XOR2_X2 sub_434_b0_U43 ( .A(sub_434_b0_n59), .B(sub_434_b0_n5), .Z(N238) );
  XOR2_X2 sub_434_b0_U42 ( .A(sub_434_b0_n60), .B(sub_434_b0_n21), .Z(N237) );
  XOR2_X2 sub_434_b0_U41 ( .A(sub_434_b0_n61), .B(sub_434_b0_n6), .Z(N236) );
  XOR2_X2 sub_434_b0_U40 ( .A(sub_434_b0_n62), .B(sub_434_b0_n22), .Z(N235) );
  XOR2_X2 sub_434_b0_U39 ( .A(sub_434_b0_n63), .B(sub_434_b0_n7), .Z(N234) );
  XOR2_X2 sub_434_b0_U38 ( .A(sub_434_b0_n65), .B(sub_434_b0_n2), .Z(N232) );
  XOR2_X2 sub_434_b0_U37 ( .A(sub_434_b0_n66), .B(sub_434_b0_n24), .Z(N231) );
  XOR2_X2 sub_434_b0_U36 ( .A(sub_434_b0_n67), .B(sub_434_b0_n8), .Z(N230) );
  XOR2_X2 sub_434_b0_U35 ( .A(sub_434_b0_n68), .B(sub_434_b0_n25), .Z(N229) );
  XOR2_X2 sub_434_b0_U34 ( .A(sub_434_b0_n69), .B(sub_434_b0_n70), .Z(N228) );
  XOR2_X2 sub_434_b0_U33 ( .A(sub_434_b0_n48), .B(sub_434_b0_n15), .Z(N249) );
  XOR2_X2 sub_434_b0_U32 ( .A(sub_434_b0_n49), .B(sub_434_b0_n3), .Z(N248) );
  XOR2_X2 sub_434_b0_U31 ( .A(sub_434_b0_n50), .B(sub_434_b0_n16), .Z(N247) );
  XOR2_X2 sub_434_b0_U30 ( .A(sub_434_b0_n51), .B(sub_434_b0_n9), .Z(N246) );
  XOR2_X2 sub_434_b0_U29 ( .A(sub_434_b0_n52), .B(sub_434_b0_n17), .Z(N245) );
  XOR2_X2 sub_434_b0_U28 ( .A(sub_434_b0_n53), .B(sub_434_b0_n10), .Z(N244) );
  XOR2_X2 sub_434_b0_U27 ( .A(sub_434_b0_n56), .B(sub_434_b0_n19), .Z(N241) );
  XOR2_X2 sub_434_b0_U26 ( .A(sub_434_b0_n47), .B(sub_434_b0_n1), .Z(N250) );
  AND2_X4 sub_434_b0_U25 ( .A1(sub_434_b0_n69), .A2(sub_434_b0_n70), .ZN(
        sub_434_b0_n25) );
  AND2_X4 sub_434_b0_U24 ( .A1(sub_434_b0_n67), .A2(sub_434_b0_n8), .ZN(
        sub_434_b0_n24) );
  AND2_X4 sub_434_b0_U23 ( .A1(sub_434_b0_n65), .A2(sub_434_b0_n2), .ZN(
        sub_434_b0_n23) );
  AND2_X4 sub_434_b0_U22 ( .A1(sub_434_b0_n63), .A2(sub_434_b0_n7), .ZN(
        sub_434_b0_n22) );
  AND2_X4 sub_434_b0_U21 ( .A1(sub_434_b0_n61), .A2(sub_434_b0_n6), .ZN(
        sub_434_b0_n21) );
  AND2_X4 sub_434_b0_U20 ( .A1(sub_434_b0_n59), .A2(sub_434_b0_n5), .ZN(
        sub_434_b0_n20) );
  AND2_X4 sub_434_b0_U19 ( .A1(sub_434_b0_n57), .A2(sub_434_b0_n4), .ZN(
        sub_434_b0_n19) );
  AND2_X4 sub_434_b0_U18 ( .A1(sub_434_b0_n55), .A2(sub_434_b0_n11), .ZN(
        sub_434_b0_n18) );
  AND2_X4 sub_434_b0_U17 ( .A1(sub_434_b0_n53), .A2(sub_434_b0_n10), .ZN(
        sub_434_b0_n17) );
  AND2_X4 sub_434_b0_U16 ( .A1(sub_434_b0_n51), .A2(sub_434_b0_n9), .ZN(
        sub_434_b0_n16) );
  AND2_X4 sub_434_b0_U15 ( .A1(sub_434_b0_n49), .A2(sub_434_b0_n3), .ZN(
        sub_434_b0_n15) );
  XOR2_X2 sub_434_b0_U14 ( .A(sub_434_b0_n64), .B(sub_434_b0_n23), .Z(N233) );
  XOR2_X2 sub_434_b0_U13 ( .A(sub_434_b0_n54), .B(sub_434_b0_n18), .Z(N243) );
  XOR2_X2 sub_434_b0_U12 ( .A(sub_434_b0_n55), .B(sub_434_b0_n11), .Z(N242) );
  AND2_X4 sub_434_b0_U11 ( .A1(sub_434_b0_n56), .A2(sub_434_b0_n19), .ZN(
        sub_434_b0_n11) );
  AND2_X4 sub_434_b0_U10 ( .A1(sub_434_b0_n54), .A2(sub_434_b0_n18), .ZN(
        sub_434_b0_n10) );
  AND2_X4 sub_434_b0_U9 ( .A1(sub_434_b0_n52), .A2(sub_434_b0_n17), .ZN(
        sub_434_b0_n9) );
  AND2_X4 sub_434_b0_U8 ( .A1(sub_434_b0_n68), .A2(sub_434_b0_n25), .ZN(
        sub_434_b0_n8) );
  AND2_X4 sub_434_b0_U7 ( .A1(sub_434_b0_n64), .A2(sub_434_b0_n23), .ZN(
        sub_434_b0_n7) );
  AND2_X4 sub_434_b0_U6 ( .A1(sub_434_b0_n62), .A2(sub_434_b0_n22), .ZN(
        sub_434_b0_n6) );
  AND2_X4 sub_434_b0_U5 ( .A1(sub_434_b0_n60), .A2(sub_434_b0_n21), .ZN(
        sub_434_b0_n5) );
  AND2_X4 sub_434_b0_U4 ( .A1(sub_434_b0_n58), .A2(sub_434_b0_n20), .ZN(
        sub_434_b0_n4) );
  AND2_X4 sub_434_b0_U3 ( .A1(sub_434_b0_n50), .A2(sub_434_b0_n16), .ZN(
        sub_434_b0_n3) );
  AND2_X4 sub_434_b0_U2 ( .A1(sub_434_b0_n66), .A2(sub_434_b0_n24), .ZN(
        sub_434_b0_n2) );
  AND2_X4 sub_434_b0_U1 ( .A1(sub_434_b0_n48), .A2(sub_434_b0_n15), .ZN(
        sub_434_b0_n1) );
  AND2_X1 sll_384_U47 ( .A1(fracta_mul[0]), .A2(sll_384_n2), .ZN(
        sll_384_ML_int_1__0_) );
  AND2_X1 sll_384_U46 ( .A1(sll_384_ML_int_1__0_), .A2(sll_384_n4), .ZN(
        sll_384_ML_int_2__0_) );
  AND2_X1 sll_384_U45 ( .A1(sll_384_ML_int_1__1_), .A2(sll_384_n4), .ZN(
        sll_384_ML_int_2__1_) );
  AND2_X1 sll_384_U44 ( .A1(sll_384_ML_int_2__0_), .A2(sll_384_n1), .ZN(
        sll_384_ML_int_3__0_) );
  AND2_X1 sll_384_U43 ( .A1(sll_384_ML_int_2__1_), .A2(sll_384_n1), .ZN(
        sll_384_ML_int_3__1_) );
  AND2_X1 sll_384_U42 ( .A1(sll_384_ML_int_2__2_), .A2(sll_384_n1), .ZN(
        sll_384_ML_int_3__2_) );
  AND2_X1 sll_384_U41 ( .A1(sll_384_ML_int_2__3_), .A2(sll_384_n1), .ZN(
        sll_384_ML_int_3__3_) );
  NAND2_X1 sll_384_U40 ( .A1(sll_384_ML_int_3__0_), .A2(sll_384_n14), .ZN(
        sll_384_n22) );
  NAND2_X1 sll_384_U39 ( .A1(sll_384_ML_int_3__1_), .A2(sll_384_n14), .ZN(
        sll_384_n21) );
  NAND2_X1 sll_384_U38 ( .A1(sll_384_ML_int_3__2_), .A2(sll_384_n14), .ZN(
        sll_384_n20) );
  NAND2_X1 sll_384_U37 ( .A1(sll_384_ML_int_3__3_), .A2(sll_384_n14), .ZN(
        sll_384_n19) );
  NAND2_X1 sll_384_U36 ( .A1(sll_384_ML_int_3__4_), .A2(sll_384_n14), .ZN(
        sll_384_n18) );
  NAND2_X1 sll_384_U35 ( .A1(sll_384_ML_int_3__5_), .A2(sll_384_n14), .ZN(
        sll_384_n17) );
  NAND2_X1 sll_384_U34 ( .A1(sll_384_ML_int_3__6_), .A2(sll_384_n14), .ZN(
        sll_384_n16) );
  NAND2_X1 sll_384_U33 ( .A1(sll_384_ML_int_3__7_), .A2(sll_384_n14), .ZN(
        sll_384_n15) );
  NOR2_X1 sll_384_U32 ( .A1(N47), .A2(sll_384_n22), .ZN(N172) );
  AND2_X1 sll_384_U31 ( .A1(sll_384_ML_int_4__10_), .A2(sll_384_n13), .ZN(N182) );
  AND2_X1 sll_384_U30 ( .A1(sll_384_ML_int_4__11_), .A2(sll_384_n13), .ZN(N183) );
  AND2_X1 sll_384_U29 ( .A1(sll_384_ML_int_4__12_), .A2(sll_384_n13), .ZN(N184) );
  AND2_X1 sll_384_U28 ( .A1(sll_384_ML_int_4__13_), .A2(sll_384_n13), .ZN(N185) );
  AND2_X1 sll_384_U27 ( .A1(sll_384_ML_int_4__14_), .A2(sll_384_n13), .ZN(N186) );
  AND2_X1 sll_384_U26 ( .A1(sll_384_ML_int_4__15_), .A2(sll_384_n13), .ZN(N187) );
  NOR2_X1 sll_384_U25 ( .A1(N47), .A2(sll_384_n21), .ZN(N173) );
  NOR2_X1 sll_384_U24 ( .A1(N47), .A2(sll_384_n20), .ZN(N174) );
  NOR2_X1 sll_384_U23 ( .A1(N47), .A2(sll_384_n19), .ZN(N175) );
  NOR2_X1 sll_384_U22 ( .A1(N47), .A2(sll_384_n18), .ZN(N176) );
  NOR2_X1 sll_384_U21 ( .A1(N47), .A2(sll_384_n17), .ZN(N177) );
  NOR2_X1 sll_384_U20 ( .A1(N47), .A2(sll_384_n16), .ZN(N178) );
  NOR2_X1 sll_384_U19 ( .A1(N47), .A2(sll_384_n15), .ZN(N179) );
  AND2_X1 sll_384_U18 ( .A1(sll_384_ML_int_4__8_), .A2(sll_384_n13), .ZN(N180)
         );
  AND2_X1 sll_384_U17 ( .A1(sll_384_ML_int_4__9_), .A2(sll_384_n13), .ZN(N181)
         );
  INV_X4 sll_384_U16 ( .A(N75), .ZN(sll_384_n14) );
  INV_X4 sll_384_U15 ( .A(N47), .ZN(sll_384_n13) );
  INV_X4 sll_384_U14 ( .A(sll_384_n15), .ZN(sll_384_n12) );
  INV_X4 sll_384_U13 ( .A(sll_384_n19), .ZN(sll_384_n11) );
  INV_X4 sll_384_U12 ( .A(sll_384_n17), .ZN(sll_384_n10) );
  INV_X4 sll_384_U11 ( .A(sll_384_n21), .ZN(sll_384_n9) );
  INV_X4 sll_384_U10 ( .A(sll_384_n16), .ZN(sll_384_n8) );
  INV_X4 sll_384_U9 ( .A(sll_384_n20), .ZN(sll_384_n7) );
  INV_X4 sll_384_U8 ( .A(sll_384_n18), .ZN(sll_384_n6) );
  INV_X4 sll_384_U7 ( .A(sll_384_n22), .ZN(sll_384_n5) );
  INV_X4 sll_384_U6 ( .A(N107), .ZN(sll_384_n1) );
  INV_X4 sll_384_U5 ( .A(N141), .ZN(sll_384_n4) );
  INV_X4 sll_384_U4 ( .A(sll_384_n2), .ZN(sll_384_n3) );
  INV_X4 sll_384_U3 ( .A(N170), .ZN(sll_384_n2) );
  MUX2_X2 sll_384_M1_0_1 ( .A(fracta_mul[1]), .B(fracta_mul[0]), .S(sll_384_n3), .Z(sll_384_ML_int_1__1_) );
  MUX2_X2 sll_384_M1_0_2 ( .A(fracta_mul[2]), .B(fracta_mul[1]), .S(sll_384_n3), .Z(sll_384_ML_int_1__2_) );
  MUX2_X2 sll_384_M1_0_3 ( .A(fracta_mul[3]), .B(fracta_mul[2]), .S(sll_384_n3), .Z(sll_384_ML_int_1__3_) );
  MUX2_X2 sll_384_M1_0_4 ( .A(fracta_mul[4]), .B(fracta_mul[3]), .S(sll_384_n3), .Z(sll_384_ML_int_1__4_) );
  MUX2_X2 sll_384_M1_0_5 ( .A(fracta_mul[5]), .B(fracta_mul[4]), .S(sll_384_n3), .Z(sll_384_ML_int_1__5_) );
  MUX2_X2 sll_384_M1_0_6 ( .A(fracta_mul[6]), .B(fracta_mul[5]), .S(sll_384_n3), .Z(sll_384_ML_int_1__6_) );
  MUX2_X2 sll_384_M1_0_7 ( .A(fracta_mul[7]), .B(fracta_mul[6]), .S(sll_384_n3), .Z(sll_384_ML_int_1__7_) );
  MUX2_X2 sll_384_M1_0_8 ( .A(fracta_mul[8]), .B(fracta_mul[7]), .S(sll_384_n3), .Z(sll_384_ML_int_1__8_) );
  MUX2_X2 sll_384_M1_0_9 ( .A(fracta_mul[9]), .B(fracta_mul[8]), .S(sll_384_n3), .Z(sll_384_ML_int_1__9_) );
  MUX2_X2 sll_384_M1_0_10 ( .A(fracta_mul[10]), .B(fracta_mul[9]), .S(
        sll_384_n3), .Z(sll_384_ML_int_1__10_) );
  MUX2_X2 sll_384_M1_0_11 ( .A(fracta_mul[11]), .B(fracta_mul[10]), .S(
        sll_384_n3), .Z(sll_384_ML_int_1__11_) );
  MUX2_X2 sll_384_M1_0_12 ( .A(fracta_mul[12]), .B(fracta_mul[11]), .S(
        sll_384_n3), .Z(sll_384_ML_int_1__12_) );
  MUX2_X2 sll_384_M1_0_13 ( .A(fracta_mul[13]), .B(fracta_mul[12]), .S(
        sll_384_n3), .Z(sll_384_ML_int_1__13_) );
  MUX2_X2 sll_384_M1_0_14 ( .A(fracta_mul[14]), .B(fracta_mul[13]), .S(N170), 
        .Z(sll_384_ML_int_1__14_) );
  MUX2_X2 sll_384_M1_0_15 ( .A(fracta_mul[15]), .B(fracta_mul[14]), .S(N170), 
        .Z(sll_384_ML_int_1__15_) );
  MUX2_X2 sll_384_M1_0_16 ( .A(fracta_mul[16]), .B(fracta_mul[15]), .S(
        sll_384_n3), .Z(sll_384_ML_int_1__16_) );
  MUX2_X2 sll_384_M1_0_17 ( .A(fracta_mul[17]), .B(fracta_mul[16]), .S(N170), 
        .Z(sll_384_ML_int_1__17_) );
  MUX2_X2 sll_384_M1_0_18 ( .A(fracta_mul[18]), .B(fracta_mul[17]), .S(N170), 
        .Z(sll_384_ML_int_1__18_) );
  MUX2_X2 sll_384_M1_0_19 ( .A(fracta_mul[19]), .B(fracta_mul[18]), .S(N170), 
        .Z(sll_384_ML_int_1__19_) );
  MUX2_X2 sll_384_M1_0_20 ( .A(fracta_mul[20]), .B(fracta_mul[19]), .S(N170), 
        .Z(sll_384_ML_int_1__20_) );
  MUX2_X2 sll_384_M1_0_21 ( .A(fracta_mul[21]), .B(fracta_mul[20]), .S(N170), 
        .Z(sll_384_ML_int_1__21_) );
  MUX2_X2 sll_384_M1_0_22 ( .A(fracta_mul[22]), .B(fracta_mul[21]), .S(N170), 
        .Z(sll_384_ML_int_1__22_) );
  MUX2_X2 sll_384_M1_0_23 ( .A(u2_N124), .B(fracta_mul[22]), .S(N170), .Z(
        sll_384_ML_int_1__23_) );
  MUX2_X2 sll_384_M1_1_2 ( .A(sll_384_ML_int_1__2_), .B(sll_384_ML_int_1__0_), 
        .S(N141), .Z(sll_384_ML_int_2__2_) );
  MUX2_X2 sll_384_M1_1_3 ( .A(sll_384_ML_int_1__3_), .B(sll_384_ML_int_1__1_), 
        .S(N141), .Z(sll_384_ML_int_2__3_) );
  MUX2_X2 sll_384_M1_1_4 ( .A(sll_384_ML_int_1__4_), .B(sll_384_ML_int_1__2_), 
        .S(N141), .Z(sll_384_ML_int_2__4_) );
  MUX2_X2 sll_384_M1_1_5 ( .A(sll_384_ML_int_1__5_), .B(sll_384_ML_int_1__3_), 
        .S(N141), .Z(sll_384_ML_int_2__5_) );
  MUX2_X2 sll_384_M1_1_6 ( .A(sll_384_ML_int_1__6_), .B(sll_384_ML_int_1__4_), 
        .S(N141), .Z(sll_384_ML_int_2__6_) );
  MUX2_X2 sll_384_M1_1_7 ( .A(sll_384_ML_int_1__7_), .B(sll_384_ML_int_1__5_), 
        .S(N141), .Z(sll_384_ML_int_2__7_) );
  MUX2_X2 sll_384_M1_1_8 ( .A(sll_384_ML_int_1__8_), .B(sll_384_ML_int_1__6_), 
        .S(N141), .Z(sll_384_ML_int_2__8_) );
  MUX2_X2 sll_384_M1_1_9 ( .A(sll_384_ML_int_1__9_), .B(sll_384_ML_int_1__7_), 
        .S(N141), .Z(sll_384_ML_int_2__9_) );
  MUX2_X2 sll_384_M1_1_10 ( .A(sll_384_ML_int_1__10_), .B(sll_384_ML_int_1__8_), .S(N141), .Z(sll_384_ML_int_2__10_) );
  MUX2_X2 sll_384_M1_1_11 ( .A(sll_384_ML_int_1__11_), .B(sll_384_ML_int_1__9_), .S(N141), .Z(sll_384_ML_int_2__11_) );
  MUX2_X2 sll_384_M1_1_12 ( .A(sll_384_ML_int_1__12_), .B(
        sll_384_ML_int_1__10_), .S(N141), .Z(sll_384_ML_int_2__12_) );
  MUX2_X2 sll_384_M1_1_13 ( .A(sll_384_ML_int_1__13_), .B(
        sll_384_ML_int_1__11_), .S(N141), .Z(sll_384_ML_int_2__13_) );
  MUX2_X2 sll_384_M1_1_14 ( .A(sll_384_ML_int_1__14_), .B(
        sll_384_ML_int_1__12_), .S(N141), .Z(sll_384_ML_int_2__14_) );
  MUX2_X2 sll_384_M1_1_15 ( .A(sll_384_ML_int_1__15_), .B(
        sll_384_ML_int_1__13_), .S(N141), .Z(sll_384_ML_int_2__15_) );
  MUX2_X2 sll_384_M1_1_16 ( .A(sll_384_ML_int_1__16_), .B(
        sll_384_ML_int_1__14_), .S(N141), .Z(sll_384_ML_int_2__16_) );
  MUX2_X2 sll_384_M1_1_17 ( .A(sll_384_ML_int_1__17_), .B(
        sll_384_ML_int_1__15_), .S(N141), .Z(sll_384_ML_int_2__17_) );
  MUX2_X2 sll_384_M1_1_18 ( .A(sll_384_ML_int_1__18_), .B(
        sll_384_ML_int_1__16_), .S(N141), .Z(sll_384_ML_int_2__18_) );
  MUX2_X2 sll_384_M1_1_19 ( .A(sll_384_ML_int_1__19_), .B(
        sll_384_ML_int_1__17_), .S(N141), .Z(sll_384_ML_int_2__19_) );
  MUX2_X2 sll_384_M1_1_20 ( .A(sll_384_ML_int_1__20_), .B(
        sll_384_ML_int_1__18_), .S(N141), .Z(sll_384_ML_int_2__20_) );
  MUX2_X2 sll_384_M1_1_21 ( .A(sll_384_ML_int_1__21_), .B(
        sll_384_ML_int_1__19_), .S(N141), .Z(sll_384_ML_int_2__21_) );
  MUX2_X2 sll_384_M1_1_22 ( .A(sll_384_ML_int_1__22_), .B(
        sll_384_ML_int_1__20_), .S(N141), .Z(sll_384_ML_int_2__22_) );
  MUX2_X2 sll_384_M1_1_23 ( .A(sll_384_ML_int_1__23_), .B(
        sll_384_ML_int_1__21_), .S(N141), .Z(sll_384_ML_int_2__23_) );
  MUX2_X2 sll_384_M1_2_4 ( .A(sll_384_ML_int_2__4_), .B(sll_384_ML_int_2__0_), 
        .S(N107), .Z(sll_384_ML_int_3__4_) );
  MUX2_X2 sll_384_M1_2_5 ( .A(sll_384_ML_int_2__5_), .B(sll_384_ML_int_2__1_), 
        .S(N107), .Z(sll_384_ML_int_3__5_) );
  MUX2_X2 sll_384_M1_2_6 ( .A(sll_384_ML_int_2__6_), .B(sll_384_ML_int_2__2_), 
        .S(N107), .Z(sll_384_ML_int_3__6_) );
  MUX2_X2 sll_384_M1_2_7 ( .A(sll_384_ML_int_2__7_), .B(sll_384_ML_int_2__3_), 
        .S(N107), .Z(sll_384_ML_int_3__7_) );
  MUX2_X2 sll_384_M1_2_8 ( .A(sll_384_ML_int_2__8_), .B(sll_384_ML_int_2__4_), 
        .S(N107), .Z(sll_384_ML_int_3__8_) );
  MUX2_X2 sll_384_M1_2_9 ( .A(sll_384_ML_int_2__9_), .B(sll_384_ML_int_2__5_), 
        .S(N107), .Z(sll_384_ML_int_3__9_) );
  MUX2_X2 sll_384_M1_2_10 ( .A(sll_384_ML_int_2__10_), .B(sll_384_ML_int_2__6_), .S(N107), .Z(sll_384_ML_int_3__10_) );
  MUX2_X2 sll_384_M1_2_11 ( .A(sll_384_ML_int_2__11_), .B(sll_384_ML_int_2__7_), .S(N107), .Z(sll_384_ML_int_3__11_) );
  MUX2_X2 sll_384_M1_2_12 ( .A(sll_384_ML_int_2__12_), .B(sll_384_ML_int_2__8_), .S(N107), .Z(sll_384_ML_int_3__12_) );
  MUX2_X2 sll_384_M1_2_13 ( .A(sll_384_ML_int_2__13_), .B(sll_384_ML_int_2__9_), .S(N107), .Z(sll_384_ML_int_3__13_) );
  MUX2_X2 sll_384_M1_2_14 ( .A(sll_384_ML_int_2__14_), .B(
        sll_384_ML_int_2__10_), .S(N107), .Z(sll_384_ML_int_3__14_) );
  MUX2_X2 sll_384_M1_2_15 ( .A(sll_384_ML_int_2__15_), .B(
        sll_384_ML_int_2__11_), .S(N107), .Z(sll_384_ML_int_3__15_) );
  MUX2_X2 sll_384_M1_2_16 ( .A(sll_384_ML_int_2__16_), .B(
        sll_384_ML_int_2__12_), .S(N107), .Z(sll_384_ML_int_3__16_) );
  MUX2_X2 sll_384_M1_2_17 ( .A(sll_384_ML_int_2__17_), .B(
        sll_384_ML_int_2__13_), .S(N107), .Z(sll_384_ML_int_3__17_) );
  MUX2_X2 sll_384_M1_2_18 ( .A(sll_384_ML_int_2__18_), .B(
        sll_384_ML_int_2__14_), .S(N107), .Z(sll_384_ML_int_3__18_) );
  MUX2_X2 sll_384_M1_2_19 ( .A(sll_384_ML_int_2__19_), .B(
        sll_384_ML_int_2__15_), .S(N107), .Z(sll_384_ML_int_3__19_) );
  MUX2_X2 sll_384_M1_2_20 ( .A(sll_384_ML_int_2__20_), .B(
        sll_384_ML_int_2__16_), .S(N107), .Z(sll_384_ML_int_3__20_) );
  MUX2_X2 sll_384_M1_2_21 ( .A(sll_384_ML_int_2__21_), .B(
        sll_384_ML_int_2__17_), .S(N107), .Z(sll_384_ML_int_3__21_) );
  MUX2_X2 sll_384_M1_2_22 ( .A(sll_384_ML_int_2__22_), .B(
        sll_384_ML_int_2__18_), .S(N107), .Z(sll_384_ML_int_3__22_) );
  MUX2_X2 sll_384_M1_2_23 ( .A(sll_384_ML_int_2__23_), .B(
        sll_384_ML_int_2__19_), .S(N107), .Z(sll_384_ML_int_3__23_) );
  MUX2_X2 sll_384_M1_3_8 ( .A(sll_384_ML_int_3__8_), .B(sll_384_ML_int_3__0_), 
        .S(N75), .Z(sll_384_ML_int_4__8_) );
  MUX2_X2 sll_384_M1_3_9 ( .A(sll_384_ML_int_3__9_), .B(sll_384_ML_int_3__1_), 
        .S(N75), .Z(sll_384_ML_int_4__9_) );
  MUX2_X2 sll_384_M1_3_10 ( .A(sll_384_ML_int_3__10_), .B(sll_384_ML_int_3__2_), .S(N75), .Z(sll_384_ML_int_4__10_) );
  MUX2_X2 sll_384_M1_3_11 ( .A(sll_384_ML_int_3__11_), .B(sll_384_ML_int_3__3_), .S(N75), .Z(sll_384_ML_int_4__11_) );
  MUX2_X2 sll_384_M1_3_12 ( .A(sll_384_ML_int_3__12_), .B(sll_384_ML_int_3__4_), .S(N75), .Z(sll_384_ML_int_4__12_) );
  MUX2_X2 sll_384_M1_3_13 ( .A(sll_384_ML_int_3__13_), .B(sll_384_ML_int_3__5_), .S(N75), .Z(sll_384_ML_int_4__13_) );
  MUX2_X2 sll_384_M1_3_14 ( .A(sll_384_ML_int_3__14_), .B(sll_384_ML_int_3__6_), .S(N75), .Z(sll_384_ML_int_4__14_) );
  MUX2_X2 sll_384_M1_3_15 ( .A(sll_384_ML_int_3__15_), .B(sll_384_ML_int_3__7_), .S(N75), .Z(sll_384_ML_int_4__15_) );
  MUX2_X2 sll_384_M1_3_16 ( .A(sll_384_ML_int_3__16_), .B(sll_384_ML_int_3__8_), .S(N75), .Z(sll_384_ML_int_4__16_) );
  MUX2_X2 sll_384_M1_3_17 ( .A(sll_384_ML_int_3__17_), .B(sll_384_ML_int_3__9_), .S(N75), .Z(sll_384_ML_int_4__17_) );
  MUX2_X2 sll_384_M1_3_18 ( .A(sll_384_ML_int_3__18_), .B(
        sll_384_ML_int_3__10_), .S(N75), .Z(sll_384_ML_int_4__18_) );
  MUX2_X2 sll_384_M1_3_19 ( .A(sll_384_ML_int_3__19_), .B(
        sll_384_ML_int_3__11_), .S(N75), .Z(sll_384_ML_int_4__19_) );
  MUX2_X2 sll_384_M1_3_20 ( .A(sll_384_ML_int_3__20_), .B(
        sll_384_ML_int_3__12_), .S(N75), .Z(sll_384_ML_int_4__20_) );
  MUX2_X2 sll_384_M1_3_21 ( .A(sll_384_ML_int_3__21_), .B(
        sll_384_ML_int_3__13_), .S(N75), .Z(sll_384_ML_int_4__21_) );
  MUX2_X2 sll_384_M1_3_22 ( .A(sll_384_ML_int_3__22_), .B(
        sll_384_ML_int_3__14_), .S(N75), .Z(sll_384_ML_int_4__22_) );
  MUX2_X2 sll_384_M1_3_23 ( .A(sll_384_ML_int_3__23_), .B(
        sll_384_ML_int_3__15_), .S(N75), .Z(sll_384_ML_int_4__23_) );
  MUX2_X2 sll_384_M1_4_16 ( .A(sll_384_ML_int_4__16_), .B(sll_384_n5), .S(N47), 
        .Z(N188) );
  MUX2_X2 sll_384_M1_4_17 ( .A(sll_384_ML_int_4__17_), .B(sll_384_n9), .S(N47), 
        .Z(N189) );
  MUX2_X2 sll_384_M1_4_18 ( .A(sll_384_ML_int_4__18_), .B(sll_384_n7), .S(N47), 
        .Z(N190) );
  MUX2_X2 sll_384_M1_4_19 ( .A(sll_384_ML_int_4__19_), .B(sll_384_n11), .S(N47), .Z(N191) );
  MUX2_X2 sll_384_M1_4_20 ( .A(sll_384_ML_int_4__20_), .B(sll_384_n6), .S(N47), 
        .Z(N192) );
  MUX2_X2 sll_384_M1_4_21 ( .A(sll_384_ML_int_4__21_), .B(sll_384_n10), .S(N47), .Z(N193) );
  MUX2_X2 sll_384_M1_4_22 ( .A(sll_384_ML_int_4__22_), .B(sll_384_n8), .S(N47), 
        .Z(N194) );
  MUX2_X2 sll_384_M1_4_23 ( .A(sll_384_ML_int_4__23_), .B(sll_384_n12), .S(N47), .Z(N195) );
  NAND2_X1 r473_U82 ( .A1(fracta_mul[2]), .A2(r473_n25), .ZN(r473_n53) );
  NAND2_X1 r473_U81 ( .A1(fracta_mul[20]), .A2(r473_n7), .ZN(r473_n37) );
  NAND2_X1 r473_U80 ( .A1(fracta_mul[19]), .A2(r473_n8), .ZN(r473_n36) );
  NAND2_X1 r473_U79 ( .A1(fracta_mul[18]), .A2(r473_n9), .ZN(r473_n41) );
  NAND2_X1 r473_U78 ( .A1(fracta_mul[17]), .A2(r473_n10), .ZN(r473_n39) );
  NAND2_X1 r473_U77 ( .A1(fracta_mul[16]), .A2(r473_n11), .ZN(r473_n40) );
  NAND2_X1 r473_U76 ( .A1(fracta_mul[15]), .A2(r473_n12), .ZN(r473_n43) );
  NAND2_X1 r473_U75 ( .A1(fracta_mul[14]), .A2(r473_n13), .ZN(r473_n45) );
  NAND2_X1 r473_U74 ( .A1(fracta_mul[13]), .A2(r473_n14), .ZN(r473_n44) );
  NAND2_X1 r473_U73 ( .A1(fracta_mul[12]), .A2(r473_n15), .ZN(r473_n48) );
  NAND2_X1 r473_U72 ( .A1(fracta_mul[11]), .A2(r473_n16), .ZN(r473_n46) );
  NAND2_X1 r473_U71 ( .A1(fracta_mul[10]), .A2(r473_n17), .ZN(r473_n47) );
  NAND2_X1 r473_U70 ( .A1(fracta_mul[9]), .A2(r473_n18), .ZN(r473_n50) );
  NAND2_X1 r473_U69 ( .A1(fracta_mul[8]), .A2(r473_n19), .ZN(r473_n52) );
  NAND2_X1 r473_U68 ( .A1(fracta_mul[7]), .A2(r473_n20), .ZN(r473_n51) );
  NAND2_X1 r473_U67 ( .A1(fracta_mul[6]), .A2(r473_n21), .ZN(r473_n56) );
  NAND2_X1 r473_U66 ( .A1(fracta_mul[5]), .A2(r473_n22), .ZN(r473_n58) );
  NAND2_X1 r473_U65 ( .A1(fracta_mul[4]), .A2(r473_n23), .ZN(r473_n57) );
  NAND2_X1 r473_U64 ( .A1(fracta_mul[3]), .A2(r473_n24), .ZN(r473_n54) );
  NOR2_X1 r473_U63 ( .A1(r473_n27), .A2(fracta_mul[0]), .ZN(r473_n80) );
  AOI21_X1 r473_U62 ( .B1(r473_n5), .B2(r473_n80), .A(u6_N1), .ZN(r473_n81) );
  OAI211_X1 r473_U61 ( .C1(r473_n80), .C2(r473_n5), .A(r473_n4), .B(r473_n53), 
        .ZN(r473_n79) );
  OAI221_X1 r473_U60 ( .B1(fracta_mul[2]), .B2(r473_n25), .C1(fracta_mul[3]), 
        .C2(r473_n24), .A(r473_n79), .ZN(r473_n78) );
  NAND3_X1 r473_U59 ( .A1(r473_n57), .A2(r473_n54), .A3(r473_n78), .ZN(
        r473_n77) );
  OAI221_X1 r473_U58 ( .B1(fracta_mul[4]), .B2(r473_n23), .C1(fracta_mul[5]), 
        .C2(r473_n22), .A(r473_n77), .ZN(r473_n76) );
  NAND3_X1 r473_U57 ( .A1(r473_n56), .A2(r473_n58), .A3(r473_n76), .ZN(
        r473_n75) );
  OAI221_X1 r473_U56 ( .B1(fracta_mul[6]), .B2(r473_n21), .C1(fracta_mul[7]), 
        .C2(r473_n20), .A(r473_n75), .ZN(r473_n74) );
  NAND3_X1 r473_U55 ( .A1(r473_n52), .A2(r473_n51), .A3(r473_n74), .ZN(
        r473_n73) );
  OAI221_X1 r473_U54 ( .B1(fracta_mul[8]), .B2(r473_n19), .C1(fracta_mul[9]), 
        .C2(r473_n18), .A(r473_n73), .ZN(r473_n72) );
  NAND3_X1 r473_U53 ( .A1(r473_n47), .A2(r473_n50), .A3(r473_n72), .ZN(
        r473_n71) );
  OAI221_X1 r473_U52 ( .B1(fracta_mul[10]), .B2(r473_n17), .C1(fracta_mul[11]), 
        .C2(r473_n16), .A(r473_n71), .ZN(r473_n70) );
  NAND3_X1 r473_U51 ( .A1(r473_n48), .A2(r473_n46), .A3(r473_n70), .ZN(
        r473_n69) );
  OAI221_X1 r473_U50 ( .B1(fracta_mul[12]), .B2(r473_n15), .C1(fracta_mul[13]), 
        .C2(r473_n14), .A(r473_n69), .ZN(r473_n68) );
  NAND3_X1 r473_U49 ( .A1(r473_n45), .A2(r473_n44), .A3(r473_n68), .ZN(
        r473_n67) );
  OAI221_X1 r473_U48 ( .B1(fracta_mul[14]), .B2(r473_n13), .C1(fracta_mul[15]), 
        .C2(r473_n12), .A(r473_n67), .ZN(r473_n66) );
  NAND3_X1 r473_U47 ( .A1(r473_n40), .A2(r473_n43), .A3(r473_n66), .ZN(
        r473_n65) );
  OAI221_X1 r473_U46 ( .B1(fracta_mul[16]), .B2(r473_n11), .C1(fracta_mul[17]), 
        .C2(r473_n10), .A(r473_n65), .ZN(r473_n64) );
  NAND3_X1 r473_U45 ( .A1(r473_n41), .A2(r473_n39), .A3(r473_n64), .ZN(
        r473_n63) );
  OAI221_X1 r473_U44 ( .B1(fracta_mul[18]), .B2(r473_n9), .C1(fracta_mul[19]), 
        .C2(r473_n8), .A(r473_n63), .ZN(r473_n62) );
  NAND3_X1 r473_U43 ( .A1(r473_n37), .A2(r473_n36), .A3(r473_n62), .ZN(
        r473_n61) );
  OAI221_X1 r473_U42 ( .B1(fracta_mul[20]), .B2(r473_n7), .C1(fracta_mul[21]), 
        .C2(r473_n6), .A(r473_n61), .ZN(r473_n60) );
  NAND2_X1 r473_U41 ( .A1(fracta_mul[21]), .A2(r473_n6), .ZN(r473_n35) );
  OAI211_X1 r473_U40 ( .C1(u6_N22), .C2(r473_n3), .A(r473_n60), .B(r473_n35), 
        .ZN(r473_n59) );
  AOI21_X1 r473_U39 ( .B1(r473_n3), .B2(u6_N22), .A(r473_n2), .ZN(r473_n28) );
  AND3_X1 r473_U38 ( .A1(r473_n56), .A2(r473_n57), .A3(r473_n58), .ZN(r473_n55) );
  NAND4_X1 r473_U37 ( .A1(r473_n53), .A2(r473_n28), .A3(r473_n54), .A4(
        r473_n55), .ZN(r473_n29) );
  AND3_X1 r473_U36 ( .A1(r473_n50), .A2(r473_n51), .A3(r473_n52), .ZN(r473_n49) );
  NAND4_X1 r473_U35 ( .A1(r473_n46), .A2(r473_n47), .A3(r473_n48), .A4(
        r473_n49), .ZN(r473_n30) );
  AND3_X1 r473_U34 ( .A1(r473_n43), .A2(r473_n44), .A3(r473_n45), .ZN(r473_n42) );
  NAND4_X1 r473_U33 ( .A1(r473_n39), .A2(r473_n40), .A3(r473_n41), .A4(
        r473_n42), .ZN(r473_n31) );
  AND2_X1 r473_U32 ( .A1(fracta_mul[0]), .A2(r473_n27), .ZN(r473_n38) );
  OAI22_X1 r473_U31 ( .A1(fracta_mul[1]), .A2(r473_n38), .B1(r473_n38), .B2(
        r473_n26), .ZN(r473_n33) );
  AND3_X1 r473_U30 ( .A1(r473_n35), .A2(r473_n36), .A3(r473_n37), .ZN(r473_n34) );
  OAI211_X1 r473_U29 ( .C1(u6_N22), .C2(r473_n3), .A(r473_n33), .B(r473_n34), 
        .ZN(r473_n32) );
  NOR4_X1 r473_U28 ( .A1(r473_n29), .A2(r473_n30), .A3(r473_n31), .A4(r473_n32), .ZN(u1_N131) );
  INV_X4 r473_U27 ( .A(u6_N0), .ZN(r473_n27) );
  INV_X4 r473_U26 ( .A(u6_N1), .ZN(r473_n26) );
  INV_X4 r473_U25 ( .A(u6_N2), .ZN(r473_n25) );
  INV_X4 r473_U24 ( .A(u6_N3), .ZN(r473_n24) );
  INV_X4 r473_U23 ( .A(u6_N4), .ZN(r473_n23) );
  INV_X4 r473_U22 ( .A(u6_N5), .ZN(r473_n22) );
  INV_X4 r473_U21 ( .A(u6_N6), .ZN(r473_n21) );
  INV_X4 r473_U20 ( .A(u6_N7), .ZN(r473_n20) );
  INV_X4 r473_U19 ( .A(u6_N8), .ZN(r473_n19) );
  INV_X4 r473_U18 ( .A(u6_N9), .ZN(r473_n18) );
  INV_X4 r473_U17 ( .A(u6_N10), .ZN(r473_n17) );
  INV_X4 r473_U16 ( .A(u6_N11), .ZN(r473_n16) );
  INV_X4 r473_U15 ( .A(u6_N12), .ZN(r473_n15) );
  INV_X4 r473_U14 ( .A(u6_N13), .ZN(r473_n14) );
  INV_X4 r473_U13 ( .A(u6_N14), .ZN(r473_n13) );
  INV_X4 r473_U12 ( .A(u6_N15), .ZN(r473_n12) );
  INV_X4 r473_U11 ( .A(u6_N16), .ZN(r473_n11) );
  INV_X4 r473_U10 ( .A(u6_N17), .ZN(r473_n10) );
  INV_X4 r473_U9 ( .A(u6_N18), .ZN(r473_n9) );
  INV_X4 r473_U8 ( .A(u6_N19), .ZN(r473_n8) );
  INV_X4 r473_U7 ( .A(u6_N20), .ZN(r473_n7) );
  INV_X4 r473_U6 ( .A(u6_N21), .ZN(r473_n6) );
  INV_X4 r473_U5 ( .A(fracta_mul[1]), .ZN(r473_n5) );
  INV_X4 r473_U4 ( .A(r473_n81), .ZN(r473_n4) );
  INV_X4 r473_U3 ( .A(fracta_mul[22]), .ZN(r473_n3) );
  INV_X4 r473_U2 ( .A(r473_n59), .ZN(r473_n2) );
  INV_X4 r473_U1 ( .A(r473_n28), .ZN(u1_N130) );
  INV_X4 sub_1_root_sub_0_root_u4_add_494_U17 ( .A(div_opa_ldz_r2[0]), .ZN(
        sub_1_root_sub_0_root_u4_add_494_n10) );
  INV_X4 sub_1_root_sub_0_root_u4_add_494_U16 ( .A(div_opa_ldz_r2[1]), .ZN(
        sub_1_root_sub_0_root_u4_add_494_n9) );
  INV_X4 sub_1_root_sub_0_root_u4_add_494_U15 ( .A(div_opa_ldz_r2[2]), .ZN(
        sub_1_root_sub_0_root_u4_add_494_n8) );
  INV_X4 sub_1_root_sub_0_root_u4_add_494_U14 ( .A(div_opa_ldz_r2[3]), .ZN(
        sub_1_root_sub_0_root_u4_add_494_n7) );
  INV_X4 sub_1_root_sub_0_root_u4_add_494_U13 ( .A(div_opa_ldz_r2[4]), .ZN(
        sub_1_root_sub_0_root_u4_add_494_n6) );
  INV_X4 sub_1_root_sub_0_root_u4_add_494_U12 ( .A(n2650), .ZN(
        sub_1_root_sub_0_root_u4_add_494_n5) );
  XNOR2_X2 sub_1_root_sub_0_root_u4_add_494_U11 ( .A(
        sub_1_root_sub_0_root_u4_add_494_n10), .B(n2650), .ZN(u4_ldz_dif_0_)
         );
  NAND2_X2 sub_1_root_sub_0_root_u4_add_494_U10 ( .A1(div_opa_ldz_r2[0]), .A2(
        sub_1_root_sub_0_root_u4_add_494_n5), .ZN(
        sub_1_root_sub_0_root_u4_add_494_carry_1_) );
  XNOR2_X2 sub_1_root_sub_0_root_u4_add_494_U9 ( .A(n2687), .B(
        sub_1_root_sub_0_root_u4_add_494_carry_7_), .ZN(u4_ldz_dif_7_) );
  INV_X4 sub_1_root_sub_0_root_u4_add_494_U8 ( .A(
        sub_1_root_sub_0_root_u4_add_494_carry_6_), .ZN(
        sub_1_root_sub_0_root_u4_add_494_n4) );
  INV_X4 sub_1_root_sub_0_root_u4_add_494_U7 ( .A(n2686), .ZN(
        sub_1_root_sub_0_root_u4_add_494_n3) );
  XNOR2_X2 sub_1_root_sub_0_root_u4_add_494_U6 ( .A(n2686), .B(
        sub_1_root_sub_0_root_u4_add_494_carry_6_), .ZN(u4_ldz_dif_6_) );
  NAND2_X2 sub_1_root_sub_0_root_u4_add_494_U5 ( .A1(
        sub_1_root_sub_0_root_u4_add_494_n3), .A2(
        sub_1_root_sub_0_root_u4_add_494_n4), .ZN(
        sub_1_root_sub_0_root_u4_add_494_carry_7_) );
  INV_X4 sub_1_root_sub_0_root_u4_add_494_U4 ( .A(
        sub_1_root_sub_0_root_u4_add_494_carry_5_), .ZN(
        sub_1_root_sub_0_root_u4_add_494_n2) );
  INV_X4 sub_1_root_sub_0_root_u4_add_494_U3 ( .A(n2685), .ZN(
        sub_1_root_sub_0_root_u4_add_494_n1) );
  XNOR2_X2 sub_1_root_sub_0_root_u4_add_494_U2 ( .A(n2685), .B(
        sub_1_root_sub_0_root_u4_add_494_carry_5_), .ZN(u4_ldz_dif_5_) );
  NAND2_X2 sub_1_root_sub_0_root_u4_add_494_U1 ( .A1(
        sub_1_root_sub_0_root_u4_add_494_n1), .A2(
        sub_1_root_sub_0_root_u4_add_494_n2), .ZN(
        sub_1_root_sub_0_root_u4_add_494_carry_6_) );
  FA_X1 sub_1_root_sub_0_root_u4_add_494_U2_1 ( .A(n2681), .B(
        sub_1_root_sub_0_root_u4_add_494_n9), .CI(
        sub_1_root_sub_0_root_u4_add_494_carry_1_), .CO(
        sub_1_root_sub_0_root_u4_add_494_carry_2_), .S(u4_ldz_dif_1_) );
  FA_X1 sub_1_root_sub_0_root_u4_add_494_U2_2 ( .A(n2682), .B(
        sub_1_root_sub_0_root_u4_add_494_n8), .CI(
        sub_1_root_sub_0_root_u4_add_494_carry_2_), .CO(
        sub_1_root_sub_0_root_u4_add_494_carry_3_), .S(u4_ldz_dif_2_) );
  FA_X1 sub_1_root_sub_0_root_u4_add_494_U2_3 ( .A(n2683), .B(
        sub_1_root_sub_0_root_u4_add_494_n7), .CI(
        sub_1_root_sub_0_root_u4_add_494_carry_3_), .CO(
        sub_1_root_sub_0_root_u4_add_494_carry_4_), .S(u4_ldz_dif_3_) );
  FA_X1 sub_1_root_sub_0_root_u4_add_494_U2_4 ( .A(n2684), .B(
        sub_1_root_sub_0_root_u4_add_494_n6), .CI(
        sub_1_root_sub_0_root_u4_add_494_carry_4_), .CO(
        sub_1_root_sub_0_root_u4_add_494_carry_5_), .S(u4_ldz_dif_4_) );
  XOR2_X2 add_0_root_sub_0_root_u4_add_494_U2 ( .A(u4_fi_ldz_2a_0_), .B(
        u4_ldz_dif_0_), .Z(u4_div_exp3[0]) );
  AND2_X4 add_0_root_sub_0_root_u4_add_494_U1 ( .A1(u4_fi_ldz_2a_0_), .A2(
        u4_ldz_dif_0_), .ZN(add_0_root_sub_0_root_u4_add_494_n1) );
  FA_X1 add_0_root_sub_0_root_u4_add_494_U1_1 ( .A(u4_ldz_dif_1_), .B(
        u4_fi_ldz_2a_1_), .CI(add_0_root_sub_0_root_u4_add_494_n1), .CO(
        add_0_root_sub_0_root_u4_add_494_carry[2]), .S(u4_div_exp3[1]) );
  FA_X1 add_0_root_sub_0_root_u4_add_494_U1_2 ( .A(u4_ldz_dif_2_), .B(n2723), 
        .CI(add_0_root_sub_0_root_u4_add_494_carry[2]), .CO(
        add_0_root_sub_0_root_u4_add_494_carry[3]), .S(u4_div_exp3[2]) );
  FA_X1 add_0_root_sub_0_root_u4_add_494_U1_3 ( .A(u4_ldz_dif_3_), .B(
        u4_fi_ldz_2a_3_), .CI(add_0_root_sub_0_root_u4_add_494_carry[3]), .CO(
        add_0_root_sub_0_root_u4_add_494_carry[4]), .S(u4_div_exp3[3]) );
  FA_X1 add_0_root_sub_0_root_u4_add_494_U1_4 ( .A(u4_ldz_dif_4_), .B(
        u4_fi_ldz_2a_4_), .CI(add_0_root_sub_0_root_u4_add_494_carry[4]), .CO(
        add_0_root_sub_0_root_u4_add_494_carry[5]), .S(u4_div_exp3[4]) );
  FA_X1 add_0_root_sub_0_root_u4_add_494_U1_5 ( .A(u4_ldz_dif_5_), .B(
        u4_fi_ldz_2a_5_), .CI(add_0_root_sub_0_root_u4_add_494_carry[5]), .CO(
        add_0_root_sub_0_root_u4_add_494_carry[6]), .S(u4_div_exp3[5]) );
  FA_X1 add_0_root_sub_0_root_u4_add_494_U1_6 ( .A(u4_ldz_dif_6_), .B(n2543), 
        .CI(add_0_root_sub_0_root_u4_add_494_carry[6]), .CO(
        add_0_root_sub_0_root_u4_add_494_carry[7]), .S(u4_div_exp3[6]) );
  FA_X1 add_0_root_sub_0_root_u4_add_494_U1_7 ( .A(u4_ldz_dif_7_), .B(n2543), 
        .CI(add_0_root_sub_0_root_u4_add_494_carry[7]), .S(u4_div_exp3[7]) );
  NOR2_X1 u5_mult_79_U718 ( .A1(u5_mult_79_n142), .A2(u5_mult_79_n118), .ZN(
        u5_N0) );
  NOR2_X1 u5_mult_79_U717 ( .A1(u5_mult_79_n132), .A2(u5_mult_79_n118), .ZN(
        u5_mult_79_ab_0__10_) );
  NOR2_X1 u5_mult_79_U716 ( .A1(u5_mult_79_n131), .A2(u5_mult_79_n118), .ZN(
        u5_mult_79_ab_0__11_) );
  NOR2_X1 u5_mult_79_U715 ( .A1(u5_mult_79_n130), .A2(u5_mult_79_n118), .ZN(
        u5_mult_79_ab_0__12_) );
  NOR2_X1 u5_mult_79_U714 ( .A1(u5_mult_79_n129), .A2(u5_mult_79_n118), .ZN(
        u5_mult_79_ab_0__13_) );
  NOR2_X1 u5_mult_79_U713 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_n118), .ZN(
        u5_mult_79_ab_0__14_) );
  NOR2_X1 u5_mult_79_U712 ( .A1(u5_mult_79_n127), .A2(u5_mult_79_n118), .ZN(
        u5_mult_79_ab_0__15_) );
  NOR2_X1 u5_mult_79_U711 ( .A1(u5_mult_79_n126), .A2(u5_mult_79_n118), .ZN(
        u5_mult_79_ab_0__16_) );
  NOR2_X1 u5_mult_79_U710 ( .A1(u5_mult_79_n125), .A2(u5_mult_79_n118), .ZN(
        u5_mult_79_ab_0__17_) );
  NOR2_X1 u5_mult_79_U709 ( .A1(u5_mult_79_n124), .A2(u5_mult_79_n118), .ZN(
        u5_mult_79_ab_0__18_) );
  NOR2_X1 u5_mult_79_U708 ( .A1(u5_mult_79_n123), .A2(u5_mult_79_n118), .ZN(
        u5_mult_79_ab_0__19_) );
  NOR2_X1 u5_mult_79_U707 ( .A1(u5_mult_79_n141), .A2(u5_mult_79_n118), .ZN(
        u5_mult_79_ab_0__1_) );
  NOR2_X1 u5_mult_79_U706 ( .A1(u5_mult_79_n122), .A2(u5_mult_79_n118), .ZN(
        u5_mult_79_ab_0__20_) );
  NOR2_X1 u5_mult_79_U705 ( .A1(u5_mult_79_n121), .A2(u5_mult_79_n118), .ZN(
        u5_mult_79_ab_0__21_) );
  NOR2_X1 u5_mult_79_U704 ( .A1(u5_mult_79_n120), .A2(u5_mult_79_n118), .ZN(
        u5_mult_79_ab_0__22_) );
  NOR2_X1 u5_mult_79_U703 ( .A1(u5_mult_79_n119), .A2(u5_mult_79_n118), .ZN(
        u5_mult_79_ab_0__23_) );
  NOR2_X1 u5_mult_79_U702 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n118), .ZN(
        u5_mult_79_ab_0__2_) );
  NOR2_X1 u5_mult_79_U701 ( .A1(u5_mult_79_n139), .A2(u5_mult_79_n118), .ZN(
        u5_mult_79_ab_0__3_) );
  NOR2_X1 u5_mult_79_U700 ( .A1(u5_mult_79_n138), .A2(u5_mult_79_n118), .ZN(
        u5_mult_79_ab_0__4_) );
  NOR2_X1 u5_mult_79_U699 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n118), .ZN(
        u5_mult_79_ab_0__5_) );
  NOR2_X1 u5_mult_79_U698 ( .A1(u5_mult_79_n136), .A2(u5_mult_79_n118), .ZN(
        u5_mult_79_ab_0__6_) );
  NOR2_X1 u5_mult_79_U697 ( .A1(u5_mult_79_n135), .A2(u5_mult_79_n118), .ZN(
        u5_mult_79_ab_0__7_) );
  NOR2_X1 u5_mult_79_U696 ( .A1(u5_mult_79_n134), .A2(u5_mult_79_n118), .ZN(
        u5_mult_79_ab_0__8_) );
  NOR2_X1 u5_mult_79_U695 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_n118), .ZN(
        u5_mult_79_ab_0__9_) );
  NOR2_X1 u5_mult_79_U694 ( .A1(u5_mult_79_n142), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__0_) );
  NOR2_X1 u5_mult_79_U693 ( .A1(u5_mult_79_n132), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__10_) );
  NOR2_X1 u5_mult_79_U692 ( .A1(u5_mult_79_n131), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__11_) );
  NOR2_X1 u5_mult_79_U691 ( .A1(u5_mult_79_n130), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__12_) );
  NOR2_X1 u5_mult_79_U690 ( .A1(u5_mult_79_n129), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__13_) );
  NOR2_X1 u5_mult_79_U689 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__14_) );
  NOR2_X1 u5_mult_79_U688 ( .A1(u5_mult_79_n127), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__15_) );
  NOR2_X1 u5_mult_79_U687 ( .A1(u5_mult_79_n126), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__16_) );
  NOR2_X1 u5_mult_79_U686 ( .A1(u5_mult_79_n125), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__17_) );
  NOR2_X1 u5_mult_79_U685 ( .A1(u5_mult_79_n124), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__18_) );
  NOR2_X1 u5_mult_79_U684 ( .A1(u5_mult_79_n123), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__19_) );
  NOR2_X1 u5_mult_79_U683 ( .A1(u5_mult_79_n141), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__1_) );
  NOR2_X1 u5_mult_79_U682 ( .A1(u5_mult_79_n122), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__20_) );
  NOR2_X1 u5_mult_79_U681 ( .A1(u5_mult_79_n121), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__21_) );
  NOR2_X1 u5_mult_79_U680 ( .A1(u5_mult_79_n120), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__22_) );
  NOR2_X1 u5_mult_79_U679 ( .A1(u5_mult_79_n119), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__23_) );
  NOR2_X1 u5_mult_79_U678 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__2_) );
  NOR2_X1 u5_mult_79_U677 ( .A1(u5_mult_79_n139), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__3_) );
  NOR2_X1 u5_mult_79_U676 ( .A1(u5_mult_79_n138), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__4_) );
  NOR2_X1 u5_mult_79_U675 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__5_) );
  NOR2_X1 u5_mult_79_U674 ( .A1(u5_mult_79_n136), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__6_) );
  NOR2_X1 u5_mult_79_U673 ( .A1(u5_mult_79_n135), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__7_) );
  NOR2_X1 u5_mult_79_U672 ( .A1(u5_mult_79_n134), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__8_) );
  NOR2_X1 u5_mult_79_U671 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_n108), .ZN(
        u5_mult_79_ab_10__9_) );
  NOR2_X1 u5_mult_79_U670 ( .A1(u5_mult_79_n142), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__0_) );
  NOR2_X1 u5_mult_79_U669 ( .A1(u5_mult_79_n132), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__10_) );
  NOR2_X1 u5_mult_79_U668 ( .A1(u5_mult_79_n131), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__11_) );
  NOR2_X1 u5_mult_79_U667 ( .A1(u5_mult_79_n130), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__12_) );
  NOR2_X1 u5_mult_79_U666 ( .A1(u5_mult_79_n129), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__13_) );
  NOR2_X1 u5_mult_79_U665 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__14_) );
  NOR2_X1 u5_mult_79_U664 ( .A1(u5_mult_79_n127), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__15_) );
  NOR2_X1 u5_mult_79_U663 ( .A1(u5_mult_79_n126), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__16_) );
  NOR2_X1 u5_mult_79_U662 ( .A1(u5_mult_79_n125), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__17_) );
  NOR2_X1 u5_mult_79_U661 ( .A1(u5_mult_79_n124), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__18_) );
  NOR2_X1 u5_mult_79_U660 ( .A1(u5_mult_79_n123), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__19_) );
  NOR2_X1 u5_mult_79_U659 ( .A1(u5_mult_79_n141), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__1_) );
  NOR2_X1 u5_mult_79_U658 ( .A1(u5_mult_79_n122), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__20_) );
  NOR2_X1 u5_mult_79_U657 ( .A1(u5_mult_79_n121), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__21_) );
  NOR2_X1 u5_mult_79_U656 ( .A1(u5_mult_79_n120), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__22_) );
  NOR2_X1 u5_mult_79_U655 ( .A1(u5_mult_79_n119), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__23_) );
  NOR2_X1 u5_mult_79_U654 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__2_) );
  NOR2_X1 u5_mult_79_U653 ( .A1(u5_mult_79_n139), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__3_) );
  NOR2_X1 u5_mult_79_U652 ( .A1(u5_mult_79_n138), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__4_) );
  NOR2_X1 u5_mult_79_U651 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__5_) );
  NOR2_X1 u5_mult_79_U650 ( .A1(u5_mult_79_n136), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__6_) );
  NOR2_X1 u5_mult_79_U649 ( .A1(u5_mult_79_n135), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__7_) );
  NOR2_X1 u5_mult_79_U648 ( .A1(u5_mult_79_n134), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__8_) );
  NOR2_X1 u5_mult_79_U647 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_n107), .ZN(
        u5_mult_79_ab_11__9_) );
  NOR2_X1 u5_mult_79_U646 ( .A1(u5_mult_79_n142), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__0_) );
  NOR2_X1 u5_mult_79_U645 ( .A1(u5_mult_79_n132), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__10_) );
  NOR2_X1 u5_mult_79_U644 ( .A1(u5_mult_79_n131), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__11_) );
  NOR2_X1 u5_mult_79_U643 ( .A1(u5_mult_79_n130), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__12_) );
  NOR2_X1 u5_mult_79_U642 ( .A1(u5_mult_79_n129), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__13_) );
  NOR2_X1 u5_mult_79_U641 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__14_) );
  NOR2_X1 u5_mult_79_U640 ( .A1(u5_mult_79_n127), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__15_) );
  NOR2_X1 u5_mult_79_U639 ( .A1(u5_mult_79_n126), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__16_) );
  NOR2_X1 u5_mult_79_U638 ( .A1(u5_mult_79_n125), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__17_) );
  NOR2_X1 u5_mult_79_U637 ( .A1(u5_mult_79_n124), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__18_) );
  NOR2_X1 u5_mult_79_U636 ( .A1(u5_mult_79_n123), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__19_) );
  NOR2_X1 u5_mult_79_U635 ( .A1(u5_mult_79_n141), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__1_) );
  NOR2_X1 u5_mult_79_U634 ( .A1(u5_mult_79_n122), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__20_) );
  NOR2_X1 u5_mult_79_U633 ( .A1(u5_mult_79_n121), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__21_) );
  NOR2_X1 u5_mult_79_U632 ( .A1(u5_mult_79_n120), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__22_) );
  NOR2_X1 u5_mult_79_U631 ( .A1(u5_mult_79_n119), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__23_) );
  NOR2_X1 u5_mult_79_U630 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__2_) );
  NOR2_X1 u5_mult_79_U629 ( .A1(u5_mult_79_n139), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__3_) );
  NOR2_X1 u5_mult_79_U628 ( .A1(u5_mult_79_n138), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__4_) );
  NOR2_X1 u5_mult_79_U627 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__5_) );
  NOR2_X1 u5_mult_79_U626 ( .A1(u5_mult_79_n136), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__6_) );
  NOR2_X1 u5_mult_79_U625 ( .A1(u5_mult_79_n135), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__7_) );
  NOR2_X1 u5_mult_79_U624 ( .A1(u5_mult_79_n134), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__8_) );
  NOR2_X1 u5_mult_79_U623 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_n106), .ZN(
        u5_mult_79_ab_12__9_) );
  NOR2_X1 u5_mult_79_U622 ( .A1(u5_mult_79_n142), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__0_) );
  NOR2_X1 u5_mult_79_U621 ( .A1(u5_mult_79_n132), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__10_) );
  NOR2_X1 u5_mult_79_U620 ( .A1(u5_mult_79_n131), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__11_) );
  NOR2_X1 u5_mult_79_U619 ( .A1(u5_mult_79_n130), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__12_) );
  NOR2_X1 u5_mult_79_U618 ( .A1(u5_mult_79_n129), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__13_) );
  NOR2_X1 u5_mult_79_U617 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__14_) );
  NOR2_X1 u5_mult_79_U616 ( .A1(u5_mult_79_n127), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__15_) );
  NOR2_X1 u5_mult_79_U615 ( .A1(u5_mult_79_n126), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__16_) );
  NOR2_X1 u5_mult_79_U614 ( .A1(u5_mult_79_n125), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__17_) );
  NOR2_X1 u5_mult_79_U613 ( .A1(u5_mult_79_n124), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__18_) );
  NOR2_X1 u5_mult_79_U612 ( .A1(u5_mult_79_n123), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__19_) );
  NOR2_X1 u5_mult_79_U611 ( .A1(u5_mult_79_n141), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__1_) );
  NOR2_X1 u5_mult_79_U610 ( .A1(u5_mult_79_n122), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__20_) );
  NOR2_X1 u5_mult_79_U609 ( .A1(u5_mult_79_n121), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__21_) );
  NOR2_X1 u5_mult_79_U608 ( .A1(u5_mult_79_n120), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__22_) );
  NOR2_X1 u5_mult_79_U607 ( .A1(u5_mult_79_n119), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__23_) );
  NOR2_X1 u5_mult_79_U606 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__2_) );
  NOR2_X1 u5_mult_79_U605 ( .A1(u5_mult_79_n139), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__3_) );
  NOR2_X1 u5_mult_79_U604 ( .A1(u5_mult_79_n138), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__4_) );
  NOR2_X1 u5_mult_79_U603 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__5_) );
  NOR2_X1 u5_mult_79_U602 ( .A1(u5_mult_79_n136), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__6_) );
  NOR2_X1 u5_mult_79_U601 ( .A1(u5_mult_79_n135), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__7_) );
  NOR2_X1 u5_mult_79_U600 ( .A1(u5_mult_79_n134), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__8_) );
  NOR2_X1 u5_mult_79_U599 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_n105), .ZN(
        u5_mult_79_ab_13__9_) );
  NOR2_X1 u5_mult_79_U598 ( .A1(u5_mult_79_n142), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__0_) );
  NOR2_X1 u5_mult_79_U597 ( .A1(u5_mult_79_n132), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__10_) );
  NOR2_X1 u5_mult_79_U596 ( .A1(u5_mult_79_n131), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__11_) );
  NOR2_X1 u5_mult_79_U595 ( .A1(u5_mult_79_n130), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__12_) );
  NOR2_X1 u5_mult_79_U594 ( .A1(u5_mult_79_n129), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__13_) );
  NOR2_X1 u5_mult_79_U593 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__14_) );
  NOR2_X1 u5_mult_79_U592 ( .A1(u5_mult_79_n127), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__15_) );
  NOR2_X1 u5_mult_79_U591 ( .A1(u5_mult_79_n126), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__16_) );
  NOR2_X1 u5_mult_79_U590 ( .A1(u5_mult_79_n125), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__17_) );
  NOR2_X1 u5_mult_79_U589 ( .A1(u5_mult_79_n124), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__18_) );
  NOR2_X1 u5_mult_79_U588 ( .A1(u5_mult_79_n123), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__19_) );
  NOR2_X1 u5_mult_79_U587 ( .A1(u5_mult_79_n141), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__1_) );
  NOR2_X1 u5_mult_79_U586 ( .A1(u5_mult_79_n122), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__20_) );
  NOR2_X1 u5_mult_79_U585 ( .A1(u5_mult_79_n121), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__21_) );
  NOR2_X1 u5_mult_79_U584 ( .A1(u5_mult_79_n120), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__22_) );
  NOR2_X1 u5_mult_79_U583 ( .A1(u5_mult_79_n119), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__23_) );
  NOR2_X1 u5_mult_79_U582 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__2_) );
  NOR2_X1 u5_mult_79_U581 ( .A1(u5_mult_79_n139), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__3_) );
  NOR2_X1 u5_mult_79_U580 ( .A1(u5_mult_79_n138), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__4_) );
  NOR2_X1 u5_mult_79_U579 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__5_) );
  NOR2_X1 u5_mult_79_U578 ( .A1(u5_mult_79_n136), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__6_) );
  NOR2_X1 u5_mult_79_U577 ( .A1(u5_mult_79_n135), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__7_) );
  NOR2_X1 u5_mult_79_U576 ( .A1(u5_mult_79_n134), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__8_) );
  NOR2_X1 u5_mult_79_U575 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_n104), .ZN(
        u5_mult_79_ab_14__9_) );
  NOR2_X1 u5_mult_79_U574 ( .A1(u5_mult_79_n142), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__0_) );
  NOR2_X1 u5_mult_79_U573 ( .A1(u5_mult_79_n132), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__10_) );
  NOR2_X1 u5_mult_79_U572 ( .A1(u5_mult_79_n131), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__11_) );
  NOR2_X1 u5_mult_79_U571 ( .A1(u5_mult_79_n130), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__12_) );
  NOR2_X1 u5_mult_79_U570 ( .A1(u5_mult_79_n129), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__13_) );
  NOR2_X1 u5_mult_79_U569 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__14_) );
  NOR2_X1 u5_mult_79_U568 ( .A1(u5_mult_79_n127), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__15_) );
  NOR2_X1 u5_mult_79_U567 ( .A1(u5_mult_79_n126), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__16_) );
  NOR2_X1 u5_mult_79_U566 ( .A1(u5_mult_79_n125), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__17_) );
  NOR2_X1 u5_mult_79_U565 ( .A1(u5_mult_79_n124), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__18_) );
  NOR2_X1 u5_mult_79_U564 ( .A1(u5_mult_79_n123), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__19_) );
  NOR2_X1 u5_mult_79_U563 ( .A1(u5_mult_79_n141), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__1_) );
  NOR2_X1 u5_mult_79_U562 ( .A1(u5_mult_79_n122), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__20_) );
  NOR2_X1 u5_mult_79_U561 ( .A1(u5_mult_79_n121), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__21_) );
  NOR2_X1 u5_mult_79_U560 ( .A1(u5_mult_79_n120), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__22_) );
  NOR2_X1 u5_mult_79_U559 ( .A1(u5_mult_79_n119), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__23_) );
  NOR2_X1 u5_mult_79_U558 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__2_) );
  NOR2_X1 u5_mult_79_U557 ( .A1(u5_mult_79_n139), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__3_) );
  NOR2_X1 u5_mult_79_U556 ( .A1(u5_mult_79_n138), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__4_) );
  NOR2_X1 u5_mult_79_U555 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__5_) );
  NOR2_X1 u5_mult_79_U554 ( .A1(u5_mult_79_n136), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__6_) );
  NOR2_X1 u5_mult_79_U553 ( .A1(u5_mult_79_n135), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__7_) );
  NOR2_X1 u5_mult_79_U552 ( .A1(u5_mult_79_n134), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__8_) );
  NOR2_X1 u5_mult_79_U551 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_n103), .ZN(
        u5_mult_79_ab_15__9_) );
  NOR2_X1 u5_mult_79_U550 ( .A1(u5_mult_79_n142), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__0_) );
  NOR2_X1 u5_mult_79_U549 ( .A1(u5_mult_79_n132), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__10_) );
  NOR2_X1 u5_mult_79_U548 ( .A1(u5_mult_79_n131), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__11_) );
  NOR2_X1 u5_mult_79_U547 ( .A1(u5_mult_79_n130), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__12_) );
  NOR2_X1 u5_mult_79_U546 ( .A1(u5_mult_79_n129), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__13_) );
  NOR2_X1 u5_mult_79_U545 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__14_) );
  NOR2_X1 u5_mult_79_U544 ( .A1(u5_mult_79_n127), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__15_) );
  NOR2_X1 u5_mult_79_U543 ( .A1(u5_mult_79_n126), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__16_) );
  NOR2_X1 u5_mult_79_U542 ( .A1(u5_mult_79_n125), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__17_) );
  NOR2_X1 u5_mult_79_U541 ( .A1(u5_mult_79_n124), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__18_) );
  NOR2_X1 u5_mult_79_U540 ( .A1(u5_mult_79_n123), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__19_) );
  NOR2_X1 u5_mult_79_U539 ( .A1(u5_mult_79_n141), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__1_) );
  NOR2_X1 u5_mult_79_U538 ( .A1(u5_mult_79_n122), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__20_) );
  NOR2_X1 u5_mult_79_U537 ( .A1(u5_mult_79_n121), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__21_) );
  NOR2_X1 u5_mult_79_U536 ( .A1(u5_mult_79_n120), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__22_) );
  NOR2_X1 u5_mult_79_U535 ( .A1(u5_mult_79_n119), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__23_) );
  NOR2_X1 u5_mult_79_U534 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__2_) );
  NOR2_X1 u5_mult_79_U533 ( .A1(u5_mult_79_n139), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__3_) );
  NOR2_X1 u5_mult_79_U532 ( .A1(u5_mult_79_n138), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__4_) );
  NOR2_X1 u5_mult_79_U531 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__5_) );
  NOR2_X1 u5_mult_79_U530 ( .A1(u5_mult_79_n136), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__6_) );
  NOR2_X1 u5_mult_79_U529 ( .A1(u5_mult_79_n135), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__7_) );
  NOR2_X1 u5_mult_79_U528 ( .A1(u5_mult_79_n134), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__8_) );
  NOR2_X1 u5_mult_79_U527 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_n102), .ZN(
        u5_mult_79_ab_16__9_) );
  NOR2_X1 u5_mult_79_U526 ( .A1(u5_mult_79_n142), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__0_) );
  NOR2_X1 u5_mult_79_U525 ( .A1(u5_mult_79_n132), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__10_) );
  NOR2_X1 u5_mult_79_U524 ( .A1(u5_mult_79_n131), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__11_) );
  NOR2_X1 u5_mult_79_U523 ( .A1(u5_mult_79_n130), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__12_) );
  NOR2_X1 u5_mult_79_U522 ( .A1(u5_mult_79_n129), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__13_) );
  NOR2_X1 u5_mult_79_U521 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__14_) );
  NOR2_X1 u5_mult_79_U520 ( .A1(u5_mult_79_n127), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__15_) );
  NOR2_X1 u5_mult_79_U519 ( .A1(u5_mult_79_n126), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__16_) );
  NOR2_X1 u5_mult_79_U518 ( .A1(u5_mult_79_n125), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__17_) );
  NOR2_X1 u5_mult_79_U517 ( .A1(u5_mult_79_n124), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__18_) );
  NOR2_X1 u5_mult_79_U516 ( .A1(u5_mult_79_n123), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__19_) );
  NOR2_X1 u5_mult_79_U515 ( .A1(u5_mult_79_n141), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__1_) );
  NOR2_X1 u5_mult_79_U514 ( .A1(u5_mult_79_n122), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__20_) );
  NOR2_X1 u5_mult_79_U513 ( .A1(u5_mult_79_n121), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__21_) );
  NOR2_X1 u5_mult_79_U512 ( .A1(u5_mult_79_n120), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__22_) );
  NOR2_X1 u5_mult_79_U511 ( .A1(u5_mult_79_n119), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__23_) );
  NOR2_X1 u5_mult_79_U510 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__2_) );
  NOR2_X1 u5_mult_79_U509 ( .A1(u5_mult_79_n139), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__3_) );
  NOR2_X1 u5_mult_79_U508 ( .A1(u5_mult_79_n138), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__4_) );
  NOR2_X1 u5_mult_79_U507 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__5_) );
  NOR2_X1 u5_mult_79_U506 ( .A1(u5_mult_79_n136), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__6_) );
  NOR2_X1 u5_mult_79_U505 ( .A1(u5_mult_79_n135), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__7_) );
  NOR2_X1 u5_mult_79_U504 ( .A1(u5_mult_79_n134), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__8_) );
  NOR2_X1 u5_mult_79_U503 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_n101), .ZN(
        u5_mult_79_ab_17__9_) );
  NOR2_X1 u5_mult_79_U502 ( .A1(u5_mult_79_n142), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__0_) );
  NOR2_X1 u5_mult_79_U501 ( .A1(u5_mult_79_n132), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__10_) );
  NOR2_X1 u5_mult_79_U500 ( .A1(u5_mult_79_n131), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__11_) );
  NOR2_X1 u5_mult_79_U499 ( .A1(u5_mult_79_n130), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__12_) );
  NOR2_X1 u5_mult_79_U498 ( .A1(u5_mult_79_n129), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__13_) );
  NOR2_X1 u5_mult_79_U497 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__14_) );
  NOR2_X1 u5_mult_79_U496 ( .A1(u5_mult_79_n127), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__15_) );
  NOR2_X1 u5_mult_79_U495 ( .A1(u5_mult_79_n126), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__16_) );
  NOR2_X1 u5_mult_79_U494 ( .A1(u5_mult_79_n125), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__17_) );
  NOR2_X1 u5_mult_79_U493 ( .A1(u5_mult_79_n124), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__18_) );
  NOR2_X1 u5_mult_79_U492 ( .A1(u5_mult_79_n123), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__19_) );
  NOR2_X1 u5_mult_79_U491 ( .A1(u5_mult_79_n141), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__1_) );
  NOR2_X1 u5_mult_79_U490 ( .A1(u5_mult_79_n122), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__20_) );
  NOR2_X1 u5_mult_79_U489 ( .A1(u5_mult_79_n121), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__21_) );
  NOR2_X1 u5_mult_79_U488 ( .A1(u5_mult_79_n120), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__22_) );
  NOR2_X1 u5_mult_79_U487 ( .A1(u5_mult_79_n119), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__23_) );
  NOR2_X1 u5_mult_79_U486 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__2_) );
  NOR2_X1 u5_mult_79_U485 ( .A1(u5_mult_79_n139), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__3_) );
  NOR2_X1 u5_mult_79_U484 ( .A1(u5_mult_79_n138), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__4_) );
  NOR2_X1 u5_mult_79_U483 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__5_) );
  NOR2_X1 u5_mult_79_U482 ( .A1(u5_mult_79_n136), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__6_) );
  NOR2_X1 u5_mult_79_U481 ( .A1(u5_mult_79_n135), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__7_) );
  NOR2_X1 u5_mult_79_U480 ( .A1(u5_mult_79_n134), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__8_) );
  NOR2_X1 u5_mult_79_U479 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_n100), .ZN(
        u5_mult_79_ab_18__9_) );
  NOR2_X1 u5_mult_79_U478 ( .A1(u5_mult_79_n142), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__0_) );
  NOR2_X1 u5_mult_79_U477 ( .A1(u5_mult_79_n132), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__10_) );
  NOR2_X1 u5_mult_79_U476 ( .A1(u5_mult_79_n131), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__11_) );
  NOR2_X1 u5_mult_79_U475 ( .A1(u5_mult_79_n130), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__12_) );
  NOR2_X1 u5_mult_79_U474 ( .A1(u5_mult_79_n129), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__13_) );
  NOR2_X1 u5_mult_79_U473 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__14_) );
  NOR2_X1 u5_mult_79_U472 ( .A1(u5_mult_79_n127), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__15_) );
  NOR2_X1 u5_mult_79_U471 ( .A1(u5_mult_79_n126), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__16_) );
  NOR2_X1 u5_mult_79_U470 ( .A1(u5_mult_79_n125), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__17_) );
  NOR2_X1 u5_mult_79_U469 ( .A1(u5_mult_79_n124), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__18_) );
  NOR2_X1 u5_mult_79_U468 ( .A1(u5_mult_79_n123), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__19_) );
  NOR2_X1 u5_mult_79_U467 ( .A1(u5_mult_79_n141), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__1_) );
  NOR2_X1 u5_mult_79_U466 ( .A1(u5_mult_79_n122), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__20_) );
  NOR2_X1 u5_mult_79_U465 ( .A1(u5_mult_79_n121), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__21_) );
  NOR2_X1 u5_mult_79_U464 ( .A1(u5_mult_79_n120), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__22_) );
  NOR2_X1 u5_mult_79_U463 ( .A1(u5_mult_79_n119), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__23_) );
  NOR2_X1 u5_mult_79_U462 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__2_) );
  NOR2_X1 u5_mult_79_U461 ( .A1(u5_mult_79_n139), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__3_) );
  NOR2_X1 u5_mult_79_U460 ( .A1(u5_mult_79_n138), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__4_) );
  NOR2_X1 u5_mult_79_U459 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__5_) );
  NOR2_X1 u5_mult_79_U458 ( .A1(u5_mult_79_n136), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__6_) );
  NOR2_X1 u5_mult_79_U457 ( .A1(u5_mult_79_n135), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__7_) );
  NOR2_X1 u5_mult_79_U456 ( .A1(u5_mult_79_n134), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__8_) );
  NOR2_X1 u5_mult_79_U455 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_n99), .ZN(
        u5_mult_79_ab_19__9_) );
  NOR2_X1 u5_mult_79_U454 ( .A1(u5_mult_79_n142), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__0_) );
  NOR2_X1 u5_mult_79_U453 ( .A1(u5_mult_79_n132), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__10_) );
  NOR2_X1 u5_mult_79_U452 ( .A1(u5_mult_79_n131), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__11_) );
  NOR2_X1 u5_mult_79_U451 ( .A1(u5_mult_79_n130), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__12_) );
  NOR2_X1 u5_mult_79_U450 ( .A1(u5_mult_79_n129), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__13_) );
  NOR2_X1 u5_mult_79_U449 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__14_) );
  NOR2_X1 u5_mult_79_U448 ( .A1(u5_mult_79_n127), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__15_) );
  NOR2_X1 u5_mult_79_U447 ( .A1(u5_mult_79_n126), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__16_) );
  NOR2_X1 u5_mult_79_U446 ( .A1(u5_mult_79_n125), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__17_) );
  NOR2_X1 u5_mult_79_U445 ( .A1(u5_mult_79_n124), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__18_) );
  NOR2_X1 u5_mult_79_U444 ( .A1(u5_mult_79_n123), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__19_) );
  NOR2_X1 u5_mult_79_U443 ( .A1(u5_mult_79_n141), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__1_) );
  NOR2_X1 u5_mult_79_U442 ( .A1(u5_mult_79_n122), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__20_) );
  NOR2_X1 u5_mult_79_U441 ( .A1(u5_mult_79_n121), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__21_) );
  NOR2_X1 u5_mult_79_U440 ( .A1(u5_mult_79_n120), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__22_) );
  NOR2_X1 u5_mult_79_U439 ( .A1(u5_mult_79_n119), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__23_) );
  NOR2_X1 u5_mult_79_U438 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__2_) );
  NOR2_X1 u5_mult_79_U437 ( .A1(u5_mult_79_n139), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__3_) );
  NOR2_X1 u5_mult_79_U436 ( .A1(u5_mult_79_n138), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__4_) );
  NOR2_X1 u5_mult_79_U435 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__5_) );
  NOR2_X1 u5_mult_79_U434 ( .A1(u5_mult_79_n136), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__6_) );
  NOR2_X1 u5_mult_79_U433 ( .A1(u5_mult_79_n135), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__7_) );
  NOR2_X1 u5_mult_79_U432 ( .A1(u5_mult_79_n134), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__8_) );
  NOR2_X1 u5_mult_79_U431 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_n117), .ZN(
        u5_mult_79_ab_1__9_) );
  NOR2_X1 u5_mult_79_U430 ( .A1(u5_mult_79_n142), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__0_) );
  NOR2_X1 u5_mult_79_U429 ( .A1(u5_mult_79_n132), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__10_) );
  NOR2_X1 u5_mult_79_U428 ( .A1(u5_mult_79_n131), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__11_) );
  NOR2_X1 u5_mult_79_U427 ( .A1(u5_mult_79_n130), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__12_) );
  NOR2_X1 u5_mult_79_U426 ( .A1(u5_mult_79_n129), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__13_) );
  NOR2_X1 u5_mult_79_U425 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__14_) );
  NOR2_X1 u5_mult_79_U424 ( .A1(u5_mult_79_n127), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__15_) );
  NOR2_X1 u5_mult_79_U423 ( .A1(u5_mult_79_n126), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__16_) );
  NOR2_X1 u5_mult_79_U422 ( .A1(u5_mult_79_n125), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__17_) );
  NOR2_X1 u5_mult_79_U421 ( .A1(u5_mult_79_n124), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__18_) );
  NOR2_X1 u5_mult_79_U420 ( .A1(u5_mult_79_n123), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__19_) );
  NOR2_X1 u5_mult_79_U419 ( .A1(u5_mult_79_n141), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__1_) );
  NOR2_X1 u5_mult_79_U418 ( .A1(u5_mult_79_n122), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__20_) );
  NOR2_X1 u5_mult_79_U417 ( .A1(u5_mult_79_n121), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__21_) );
  NOR2_X1 u5_mult_79_U416 ( .A1(u5_mult_79_n120), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__22_) );
  NOR2_X1 u5_mult_79_U415 ( .A1(u5_mult_79_n119), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__23_) );
  NOR2_X1 u5_mult_79_U414 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__2_) );
  NOR2_X1 u5_mult_79_U413 ( .A1(u5_mult_79_n139), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__3_) );
  NOR2_X1 u5_mult_79_U412 ( .A1(u5_mult_79_n138), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__4_) );
  NOR2_X1 u5_mult_79_U411 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__5_) );
  NOR2_X1 u5_mult_79_U410 ( .A1(u5_mult_79_n136), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__6_) );
  NOR2_X1 u5_mult_79_U409 ( .A1(u5_mult_79_n135), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__7_) );
  NOR2_X1 u5_mult_79_U408 ( .A1(u5_mult_79_n134), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__8_) );
  NOR2_X1 u5_mult_79_U407 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_n98), .ZN(
        u5_mult_79_ab_20__9_) );
  NOR2_X1 u5_mult_79_U406 ( .A1(u5_mult_79_n142), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__0_) );
  NOR2_X1 u5_mult_79_U405 ( .A1(u5_mult_79_n132), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__10_) );
  NOR2_X1 u5_mult_79_U404 ( .A1(u5_mult_79_n131), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__11_) );
  NOR2_X1 u5_mult_79_U403 ( .A1(u5_mult_79_n130), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__12_) );
  NOR2_X1 u5_mult_79_U402 ( .A1(u5_mult_79_n129), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__13_) );
  NOR2_X1 u5_mult_79_U401 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__14_) );
  NOR2_X1 u5_mult_79_U400 ( .A1(u5_mult_79_n127), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__15_) );
  NOR2_X1 u5_mult_79_U399 ( .A1(u5_mult_79_n126), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__16_) );
  NOR2_X1 u5_mult_79_U398 ( .A1(u5_mult_79_n125), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__17_) );
  NOR2_X1 u5_mult_79_U397 ( .A1(u5_mult_79_n124), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__18_) );
  NOR2_X1 u5_mult_79_U396 ( .A1(u5_mult_79_n123), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__19_) );
  NOR2_X1 u5_mult_79_U395 ( .A1(u5_mult_79_n141), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__1_) );
  NOR2_X1 u5_mult_79_U394 ( .A1(u5_mult_79_n122), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__20_) );
  NOR2_X1 u5_mult_79_U393 ( .A1(u5_mult_79_n121), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__21_) );
  NOR2_X1 u5_mult_79_U392 ( .A1(u5_mult_79_n120), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__22_) );
  NOR2_X1 u5_mult_79_U391 ( .A1(u5_mult_79_n119), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__23_) );
  NOR2_X1 u5_mult_79_U390 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__2_) );
  NOR2_X1 u5_mult_79_U389 ( .A1(u5_mult_79_n139), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__3_) );
  NOR2_X1 u5_mult_79_U388 ( .A1(u5_mult_79_n138), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__4_) );
  NOR2_X1 u5_mult_79_U387 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__5_) );
  NOR2_X1 u5_mult_79_U386 ( .A1(u5_mult_79_n136), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__6_) );
  NOR2_X1 u5_mult_79_U385 ( .A1(u5_mult_79_n135), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__7_) );
  NOR2_X1 u5_mult_79_U384 ( .A1(u5_mult_79_n134), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__8_) );
  NOR2_X1 u5_mult_79_U383 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_n97), .ZN(
        u5_mult_79_ab_21__9_) );
  NOR2_X1 u5_mult_79_U382 ( .A1(u5_mult_79_n142), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__0_) );
  NOR2_X1 u5_mult_79_U381 ( .A1(u5_mult_79_n132), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__10_) );
  NOR2_X1 u5_mult_79_U380 ( .A1(u5_mult_79_n131), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__11_) );
  NOR2_X1 u5_mult_79_U379 ( .A1(u5_mult_79_n130), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__12_) );
  NOR2_X1 u5_mult_79_U378 ( .A1(u5_mult_79_n129), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__13_) );
  NOR2_X1 u5_mult_79_U377 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__14_) );
  NOR2_X1 u5_mult_79_U376 ( .A1(u5_mult_79_n127), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__15_) );
  NOR2_X1 u5_mult_79_U375 ( .A1(u5_mult_79_n126), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__16_) );
  NOR2_X1 u5_mult_79_U374 ( .A1(u5_mult_79_n125), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__17_) );
  NOR2_X1 u5_mult_79_U373 ( .A1(u5_mult_79_n124), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__18_) );
  NOR2_X1 u5_mult_79_U372 ( .A1(u5_mult_79_n123), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__19_) );
  NOR2_X1 u5_mult_79_U371 ( .A1(u5_mult_79_n141), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__1_) );
  NOR2_X1 u5_mult_79_U370 ( .A1(u5_mult_79_n122), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__20_) );
  NOR2_X1 u5_mult_79_U369 ( .A1(u5_mult_79_n121), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__21_) );
  NOR2_X1 u5_mult_79_U368 ( .A1(u5_mult_79_n120), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__22_) );
  NOR2_X1 u5_mult_79_U367 ( .A1(u5_mult_79_n119), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__23_) );
  NOR2_X1 u5_mult_79_U366 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__2_) );
  NOR2_X1 u5_mult_79_U365 ( .A1(u5_mult_79_n139), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__3_) );
  NOR2_X1 u5_mult_79_U364 ( .A1(u5_mult_79_n138), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__4_) );
  NOR2_X1 u5_mult_79_U363 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__5_) );
  NOR2_X1 u5_mult_79_U362 ( .A1(u5_mult_79_n136), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__6_) );
  NOR2_X1 u5_mult_79_U361 ( .A1(u5_mult_79_n135), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__7_) );
  NOR2_X1 u5_mult_79_U360 ( .A1(u5_mult_79_n134), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__8_) );
  NOR2_X1 u5_mult_79_U359 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_n96), .ZN(
        u5_mult_79_ab_22__9_) );
  NOR2_X1 u5_mult_79_U358 ( .A1(u5_mult_79_n142), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__0_) );
  NOR2_X1 u5_mult_79_U357 ( .A1(u5_mult_79_n132), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__10_) );
  NOR2_X1 u5_mult_79_U356 ( .A1(u5_mult_79_n131), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__11_) );
  NOR2_X1 u5_mult_79_U355 ( .A1(u5_mult_79_n130), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__12_) );
  NOR2_X1 u5_mult_79_U354 ( .A1(u5_mult_79_n129), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__13_) );
  NOR2_X1 u5_mult_79_U353 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__14_) );
  NOR2_X1 u5_mult_79_U352 ( .A1(u5_mult_79_n127), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__15_) );
  NOR2_X1 u5_mult_79_U351 ( .A1(u5_mult_79_n126), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__16_) );
  NOR2_X1 u5_mult_79_U350 ( .A1(u5_mult_79_n125), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__17_) );
  NOR2_X1 u5_mult_79_U349 ( .A1(u5_mult_79_n124), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__18_) );
  NOR2_X1 u5_mult_79_U348 ( .A1(u5_mult_79_n123), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__19_) );
  NOR2_X1 u5_mult_79_U347 ( .A1(u5_mult_79_n141), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__1_) );
  NOR2_X1 u5_mult_79_U346 ( .A1(u5_mult_79_n122), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__20_) );
  NOR2_X1 u5_mult_79_U345 ( .A1(u5_mult_79_n121), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__21_) );
  NOR2_X1 u5_mult_79_U344 ( .A1(u5_mult_79_n120), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__22_) );
  NOR2_X1 u5_mult_79_U343 ( .A1(u5_mult_79_n119), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__23_) );
  NOR2_X1 u5_mult_79_U342 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__2_) );
  NOR2_X1 u5_mult_79_U341 ( .A1(u5_mult_79_n139), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__3_) );
  NOR2_X1 u5_mult_79_U340 ( .A1(u5_mult_79_n138), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__4_) );
  NOR2_X1 u5_mult_79_U339 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__5_) );
  NOR2_X1 u5_mult_79_U338 ( .A1(u5_mult_79_n136), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__6_) );
  NOR2_X1 u5_mult_79_U337 ( .A1(u5_mult_79_n135), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__7_) );
  NOR2_X1 u5_mult_79_U336 ( .A1(u5_mult_79_n134), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__8_) );
  NOR2_X1 u5_mult_79_U335 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_n95), .ZN(
        u5_mult_79_ab_23__9_) );
  NOR2_X1 u5_mult_79_U334 ( .A1(u5_mult_79_n142), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__0_) );
  NOR2_X1 u5_mult_79_U333 ( .A1(u5_mult_79_n132), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__10_) );
  NOR2_X1 u5_mult_79_U332 ( .A1(u5_mult_79_n131), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__11_) );
  NOR2_X1 u5_mult_79_U331 ( .A1(u5_mult_79_n130), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__12_) );
  NOR2_X1 u5_mult_79_U330 ( .A1(u5_mult_79_n129), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__13_) );
  NOR2_X1 u5_mult_79_U329 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__14_) );
  NOR2_X1 u5_mult_79_U328 ( .A1(u5_mult_79_n127), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__15_) );
  NOR2_X1 u5_mult_79_U327 ( .A1(u5_mult_79_n126), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__16_) );
  NOR2_X1 u5_mult_79_U326 ( .A1(u5_mult_79_n125), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__17_) );
  NOR2_X1 u5_mult_79_U325 ( .A1(u5_mult_79_n124), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__18_) );
  NOR2_X1 u5_mult_79_U324 ( .A1(u5_mult_79_n123), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__19_) );
  NOR2_X1 u5_mult_79_U323 ( .A1(u5_mult_79_n141), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__1_) );
  NOR2_X1 u5_mult_79_U322 ( .A1(u5_mult_79_n122), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__20_) );
  NOR2_X1 u5_mult_79_U321 ( .A1(u5_mult_79_n121), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__21_) );
  NOR2_X1 u5_mult_79_U320 ( .A1(u5_mult_79_n120), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__22_) );
  NOR2_X1 u5_mult_79_U319 ( .A1(u5_mult_79_n119), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__23_) );
  NOR2_X1 u5_mult_79_U318 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__2_) );
  NOR2_X1 u5_mult_79_U317 ( .A1(u5_mult_79_n139), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__3_) );
  NOR2_X1 u5_mult_79_U316 ( .A1(u5_mult_79_n138), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__4_) );
  NOR2_X1 u5_mult_79_U315 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__5_) );
  NOR2_X1 u5_mult_79_U314 ( .A1(u5_mult_79_n136), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__6_) );
  NOR2_X1 u5_mult_79_U313 ( .A1(u5_mult_79_n135), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__7_) );
  NOR2_X1 u5_mult_79_U312 ( .A1(u5_mult_79_n134), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__8_) );
  NOR2_X1 u5_mult_79_U311 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_ab_2__9_) );
  NOR2_X1 u5_mult_79_U310 ( .A1(u5_mult_79_n142), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__0_) );
  NOR2_X1 u5_mult_79_U309 ( .A1(u5_mult_79_n132), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__10_) );
  NOR2_X1 u5_mult_79_U308 ( .A1(u5_mult_79_n131), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__11_) );
  NOR2_X1 u5_mult_79_U307 ( .A1(u5_mult_79_n130), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__12_) );
  NOR2_X1 u5_mult_79_U306 ( .A1(u5_mult_79_n129), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__13_) );
  NOR2_X1 u5_mult_79_U305 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__14_) );
  NOR2_X1 u5_mult_79_U304 ( .A1(u5_mult_79_n127), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__15_) );
  NOR2_X1 u5_mult_79_U303 ( .A1(u5_mult_79_n126), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__16_) );
  NOR2_X1 u5_mult_79_U302 ( .A1(u5_mult_79_n125), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__17_) );
  NOR2_X1 u5_mult_79_U301 ( .A1(u5_mult_79_n124), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__18_) );
  NOR2_X1 u5_mult_79_U300 ( .A1(u5_mult_79_n123), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__19_) );
  NOR2_X1 u5_mult_79_U299 ( .A1(u5_mult_79_n141), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__1_) );
  NOR2_X1 u5_mult_79_U298 ( .A1(u5_mult_79_n122), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__20_) );
  NOR2_X1 u5_mult_79_U297 ( .A1(u5_mult_79_n121), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__21_) );
  NOR2_X1 u5_mult_79_U296 ( .A1(u5_mult_79_n120), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__22_) );
  NOR2_X1 u5_mult_79_U295 ( .A1(u5_mult_79_n119), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__23_) );
  NOR2_X1 u5_mult_79_U294 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__2_) );
  NOR2_X1 u5_mult_79_U293 ( .A1(u5_mult_79_n139), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__3_) );
  NOR2_X1 u5_mult_79_U292 ( .A1(u5_mult_79_n138), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__4_) );
  NOR2_X1 u5_mult_79_U291 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__5_) );
  NOR2_X1 u5_mult_79_U290 ( .A1(u5_mult_79_n136), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__6_) );
  NOR2_X1 u5_mult_79_U289 ( .A1(u5_mult_79_n135), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__7_) );
  NOR2_X1 u5_mult_79_U288 ( .A1(u5_mult_79_n134), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__8_) );
  NOR2_X1 u5_mult_79_U287 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_n115), .ZN(
        u5_mult_79_ab_3__9_) );
  NOR2_X1 u5_mult_79_U286 ( .A1(u5_mult_79_n142), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__0_) );
  NOR2_X1 u5_mult_79_U285 ( .A1(u5_mult_79_n132), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__10_) );
  NOR2_X1 u5_mult_79_U284 ( .A1(u5_mult_79_n131), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__11_) );
  NOR2_X1 u5_mult_79_U283 ( .A1(u5_mult_79_n130), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__12_) );
  NOR2_X1 u5_mult_79_U282 ( .A1(u5_mult_79_n129), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__13_) );
  NOR2_X1 u5_mult_79_U281 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__14_) );
  NOR2_X1 u5_mult_79_U280 ( .A1(u5_mult_79_n127), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__15_) );
  NOR2_X1 u5_mult_79_U279 ( .A1(u5_mult_79_n126), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__16_) );
  NOR2_X1 u5_mult_79_U278 ( .A1(u5_mult_79_n125), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__17_) );
  NOR2_X1 u5_mult_79_U277 ( .A1(u5_mult_79_n124), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__18_) );
  NOR2_X1 u5_mult_79_U276 ( .A1(u5_mult_79_n123), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__19_) );
  NOR2_X1 u5_mult_79_U275 ( .A1(u5_mult_79_n141), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__1_) );
  NOR2_X1 u5_mult_79_U274 ( .A1(u5_mult_79_n122), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__20_) );
  NOR2_X1 u5_mult_79_U273 ( .A1(u5_mult_79_n121), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__21_) );
  NOR2_X1 u5_mult_79_U272 ( .A1(u5_mult_79_n120), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__22_) );
  NOR2_X1 u5_mult_79_U271 ( .A1(u5_mult_79_n119), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__23_) );
  NOR2_X1 u5_mult_79_U270 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__2_) );
  NOR2_X1 u5_mult_79_U269 ( .A1(u5_mult_79_n139), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__3_) );
  NOR2_X1 u5_mult_79_U268 ( .A1(u5_mult_79_n138), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__4_) );
  NOR2_X1 u5_mult_79_U267 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__5_) );
  NOR2_X1 u5_mult_79_U266 ( .A1(u5_mult_79_n136), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__6_) );
  NOR2_X1 u5_mult_79_U265 ( .A1(u5_mult_79_n135), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__7_) );
  NOR2_X1 u5_mult_79_U264 ( .A1(u5_mult_79_n134), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__8_) );
  NOR2_X1 u5_mult_79_U263 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_n114), .ZN(
        u5_mult_79_ab_4__9_) );
  NOR2_X1 u5_mult_79_U262 ( .A1(u5_mult_79_n142), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__0_) );
  NOR2_X1 u5_mult_79_U261 ( .A1(u5_mult_79_n132), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__10_) );
  NOR2_X1 u5_mult_79_U260 ( .A1(u5_mult_79_n131), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__11_) );
  NOR2_X1 u5_mult_79_U259 ( .A1(u5_mult_79_n130), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__12_) );
  NOR2_X1 u5_mult_79_U258 ( .A1(u5_mult_79_n129), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__13_) );
  NOR2_X1 u5_mult_79_U257 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__14_) );
  NOR2_X1 u5_mult_79_U256 ( .A1(u5_mult_79_n127), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__15_) );
  NOR2_X1 u5_mult_79_U255 ( .A1(u5_mult_79_n126), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__16_) );
  NOR2_X1 u5_mult_79_U254 ( .A1(u5_mult_79_n125), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__17_) );
  NOR2_X1 u5_mult_79_U253 ( .A1(u5_mult_79_n124), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__18_) );
  NOR2_X1 u5_mult_79_U252 ( .A1(u5_mult_79_n123), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__19_) );
  NOR2_X1 u5_mult_79_U251 ( .A1(u5_mult_79_n141), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__1_) );
  NOR2_X1 u5_mult_79_U250 ( .A1(u5_mult_79_n122), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__20_) );
  NOR2_X1 u5_mult_79_U249 ( .A1(u5_mult_79_n121), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__21_) );
  NOR2_X1 u5_mult_79_U248 ( .A1(u5_mult_79_n120), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__22_) );
  NOR2_X1 u5_mult_79_U247 ( .A1(u5_mult_79_n119), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__23_) );
  NOR2_X1 u5_mult_79_U246 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__2_) );
  NOR2_X1 u5_mult_79_U245 ( .A1(u5_mult_79_n139), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__3_) );
  NOR2_X1 u5_mult_79_U244 ( .A1(u5_mult_79_n138), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__4_) );
  NOR2_X1 u5_mult_79_U243 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__5_) );
  NOR2_X1 u5_mult_79_U242 ( .A1(u5_mult_79_n136), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__6_) );
  NOR2_X1 u5_mult_79_U241 ( .A1(u5_mult_79_n135), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__7_) );
  NOR2_X1 u5_mult_79_U240 ( .A1(u5_mult_79_n134), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__8_) );
  NOR2_X1 u5_mult_79_U239 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_n113), .ZN(
        u5_mult_79_ab_5__9_) );
  NOR2_X1 u5_mult_79_U238 ( .A1(u5_mult_79_n142), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__0_) );
  NOR2_X1 u5_mult_79_U237 ( .A1(u5_mult_79_n132), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__10_) );
  NOR2_X1 u5_mult_79_U236 ( .A1(u5_mult_79_n131), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__11_) );
  NOR2_X1 u5_mult_79_U235 ( .A1(u5_mult_79_n130), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__12_) );
  NOR2_X1 u5_mult_79_U234 ( .A1(u5_mult_79_n129), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__13_) );
  NOR2_X1 u5_mult_79_U233 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__14_) );
  NOR2_X1 u5_mult_79_U232 ( .A1(u5_mult_79_n127), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__15_) );
  NOR2_X1 u5_mult_79_U231 ( .A1(u5_mult_79_n126), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__16_) );
  NOR2_X1 u5_mult_79_U230 ( .A1(u5_mult_79_n125), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__17_) );
  NOR2_X1 u5_mult_79_U229 ( .A1(u5_mult_79_n124), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__18_) );
  NOR2_X1 u5_mult_79_U228 ( .A1(u5_mult_79_n123), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__19_) );
  NOR2_X1 u5_mult_79_U227 ( .A1(u5_mult_79_n141), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__1_) );
  NOR2_X1 u5_mult_79_U226 ( .A1(u5_mult_79_n122), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__20_) );
  NOR2_X1 u5_mult_79_U225 ( .A1(u5_mult_79_n121), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__21_) );
  NOR2_X1 u5_mult_79_U224 ( .A1(u5_mult_79_n120), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__22_) );
  NOR2_X1 u5_mult_79_U223 ( .A1(u5_mult_79_n119), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__23_) );
  NOR2_X1 u5_mult_79_U222 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__2_) );
  NOR2_X1 u5_mult_79_U221 ( .A1(u5_mult_79_n139), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__3_) );
  NOR2_X1 u5_mult_79_U220 ( .A1(u5_mult_79_n138), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__4_) );
  NOR2_X1 u5_mult_79_U219 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__5_) );
  NOR2_X1 u5_mult_79_U218 ( .A1(u5_mult_79_n136), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__6_) );
  NOR2_X1 u5_mult_79_U217 ( .A1(u5_mult_79_n135), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__7_) );
  NOR2_X1 u5_mult_79_U216 ( .A1(u5_mult_79_n134), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__8_) );
  NOR2_X1 u5_mult_79_U215 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_n112), .ZN(
        u5_mult_79_ab_6__9_) );
  NOR2_X1 u5_mult_79_U214 ( .A1(u5_mult_79_n142), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__0_) );
  NOR2_X1 u5_mult_79_U213 ( .A1(u5_mult_79_n132), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__10_) );
  NOR2_X1 u5_mult_79_U212 ( .A1(u5_mult_79_n131), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__11_) );
  NOR2_X1 u5_mult_79_U211 ( .A1(u5_mult_79_n130), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__12_) );
  NOR2_X1 u5_mult_79_U210 ( .A1(u5_mult_79_n129), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__13_) );
  NOR2_X1 u5_mult_79_U209 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__14_) );
  NOR2_X1 u5_mult_79_U208 ( .A1(u5_mult_79_n127), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__15_) );
  NOR2_X1 u5_mult_79_U207 ( .A1(u5_mult_79_n126), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__16_) );
  NOR2_X1 u5_mult_79_U206 ( .A1(u5_mult_79_n125), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__17_) );
  NOR2_X1 u5_mult_79_U205 ( .A1(u5_mult_79_n124), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__18_) );
  NOR2_X1 u5_mult_79_U204 ( .A1(u5_mult_79_n123), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__19_) );
  NOR2_X1 u5_mult_79_U203 ( .A1(u5_mult_79_n141), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__1_) );
  NOR2_X1 u5_mult_79_U202 ( .A1(u5_mult_79_n122), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__20_) );
  NOR2_X1 u5_mult_79_U201 ( .A1(u5_mult_79_n121), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__21_) );
  NOR2_X1 u5_mult_79_U200 ( .A1(u5_mult_79_n120), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__22_) );
  NOR2_X1 u5_mult_79_U199 ( .A1(u5_mult_79_n119), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__23_) );
  NOR2_X1 u5_mult_79_U198 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__2_) );
  NOR2_X1 u5_mult_79_U197 ( .A1(u5_mult_79_n139), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__3_) );
  NOR2_X1 u5_mult_79_U196 ( .A1(u5_mult_79_n138), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__4_) );
  NOR2_X1 u5_mult_79_U195 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__5_) );
  NOR2_X1 u5_mult_79_U194 ( .A1(u5_mult_79_n136), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__6_) );
  NOR2_X1 u5_mult_79_U193 ( .A1(u5_mult_79_n135), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__7_) );
  NOR2_X1 u5_mult_79_U192 ( .A1(u5_mult_79_n134), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__8_) );
  NOR2_X1 u5_mult_79_U191 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_n111), .ZN(
        u5_mult_79_ab_7__9_) );
  NOR2_X1 u5_mult_79_U190 ( .A1(u5_mult_79_n142), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__0_) );
  NOR2_X1 u5_mult_79_U189 ( .A1(u5_mult_79_n132), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__10_) );
  NOR2_X1 u5_mult_79_U188 ( .A1(u5_mult_79_n131), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__11_) );
  NOR2_X1 u5_mult_79_U187 ( .A1(u5_mult_79_n130), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__12_) );
  NOR2_X1 u5_mult_79_U186 ( .A1(u5_mult_79_n129), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__13_) );
  NOR2_X1 u5_mult_79_U185 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__14_) );
  NOR2_X1 u5_mult_79_U184 ( .A1(u5_mult_79_n127), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__15_) );
  NOR2_X1 u5_mult_79_U183 ( .A1(u5_mult_79_n126), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__16_) );
  NOR2_X1 u5_mult_79_U182 ( .A1(u5_mult_79_n125), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__17_) );
  NOR2_X1 u5_mult_79_U181 ( .A1(u5_mult_79_n124), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__18_) );
  NOR2_X1 u5_mult_79_U180 ( .A1(u5_mult_79_n123), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__19_) );
  NOR2_X1 u5_mult_79_U179 ( .A1(u5_mult_79_n141), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__1_) );
  NOR2_X1 u5_mult_79_U178 ( .A1(u5_mult_79_n122), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__20_) );
  NOR2_X1 u5_mult_79_U177 ( .A1(u5_mult_79_n121), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__21_) );
  NOR2_X1 u5_mult_79_U176 ( .A1(u5_mult_79_n120), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__22_) );
  NOR2_X1 u5_mult_79_U175 ( .A1(u5_mult_79_n119), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__23_) );
  NOR2_X1 u5_mult_79_U174 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__2_) );
  NOR2_X1 u5_mult_79_U173 ( .A1(u5_mult_79_n139), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__3_) );
  NOR2_X1 u5_mult_79_U172 ( .A1(u5_mult_79_n138), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__4_) );
  NOR2_X1 u5_mult_79_U171 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__5_) );
  NOR2_X1 u5_mult_79_U170 ( .A1(u5_mult_79_n136), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__6_) );
  NOR2_X1 u5_mult_79_U169 ( .A1(u5_mult_79_n135), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__7_) );
  NOR2_X1 u5_mult_79_U168 ( .A1(u5_mult_79_n134), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__8_) );
  NOR2_X1 u5_mult_79_U167 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_n110), .ZN(
        u5_mult_79_ab_8__9_) );
  NOR2_X1 u5_mult_79_U166 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n142), .ZN(
        u5_mult_79_ab_9__0_) );
  NOR2_X1 u5_mult_79_U165 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n132), .ZN(
        u5_mult_79_ab_9__10_) );
  NOR2_X1 u5_mult_79_U164 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n131), .ZN(
        u5_mult_79_ab_9__11_) );
  NOR2_X1 u5_mult_79_U163 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n130), .ZN(
        u5_mult_79_ab_9__12_) );
  NOR2_X1 u5_mult_79_U162 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n129), .ZN(
        u5_mult_79_ab_9__13_) );
  NOR2_X1 u5_mult_79_U161 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n128), .ZN(
        u5_mult_79_ab_9__14_) );
  NOR2_X1 u5_mult_79_U160 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n127), .ZN(
        u5_mult_79_ab_9__15_) );
  NOR2_X1 u5_mult_79_U159 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n126), .ZN(
        u5_mult_79_ab_9__16_) );
  NOR2_X1 u5_mult_79_U158 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n125), .ZN(
        u5_mult_79_ab_9__17_) );
  NOR2_X1 u5_mult_79_U157 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n124), .ZN(
        u5_mult_79_ab_9__18_) );
  NOR2_X1 u5_mult_79_U156 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n123), .ZN(
        u5_mult_79_ab_9__19_) );
  NOR2_X1 u5_mult_79_U155 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n141), .ZN(
        u5_mult_79_ab_9__1_) );
  NOR2_X1 u5_mult_79_U154 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n122), .ZN(
        u5_mult_79_ab_9__20_) );
  NOR2_X1 u5_mult_79_U153 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n121), .ZN(
        u5_mult_79_ab_9__21_) );
  NOR2_X1 u5_mult_79_U152 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n120), .ZN(
        u5_mult_79_ab_9__22_) );
  NOR2_X1 u5_mult_79_U151 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n119), .ZN(
        u5_mult_79_ab_9__23_) );
  NOR2_X1 u5_mult_79_U150 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n140), .ZN(
        u5_mult_79_ab_9__2_) );
  NOR2_X1 u5_mult_79_U149 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n139), .ZN(
        u5_mult_79_ab_9__3_) );
  NOR2_X1 u5_mult_79_U148 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n138), .ZN(
        u5_mult_79_ab_9__4_) );
  NOR2_X1 u5_mult_79_U147 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n137), .ZN(
        u5_mult_79_ab_9__5_) );
  NOR2_X1 u5_mult_79_U146 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n136), .ZN(
        u5_mult_79_ab_9__6_) );
  NOR2_X1 u5_mult_79_U145 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n135), .ZN(
        u5_mult_79_ab_9__7_) );
  NOR2_X1 u5_mult_79_U144 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n134), .ZN(
        u5_mult_79_ab_9__8_) );
  NOR2_X1 u5_mult_79_U143 ( .A1(u5_mult_79_n109), .A2(u5_mult_79_n133), .ZN(
        u5_mult_79_ab_9__9_) );
  XOR2_X2 u5_mult_79_U141 ( .A(u5_mult_79_ab_1__0_), .B(u5_mult_79_ab_0__1_), 
        .Z(u5_N1) );
  INV_X4 u5_mult_79_U140 ( .A(n2651), .ZN(u5_mult_79_n95) );
  AND2_X4 u5_mult_79_U139 ( .A1(u5_mult_79_SUMB_23__22_), .A2(
        u5_mult_79_CARRYB_23__21_), .ZN(u5_mult_79_n93) );
  AND2_X4 u5_mult_79_U138 ( .A1(u5_mult_79_ab_23__23_), .A2(
        u5_mult_79_CARRYB_23__22_), .ZN(u5_mult_79_n92) );
  XOR2_X2 u5_mult_79_U137 ( .A(u5_mult_79_CARRYB_23__0_), .B(
        u5_mult_79_SUMB_23__1_), .Z(u5_N24) );
  AND2_X4 u5_mult_79_U136 ( .A1(u5_mult_79_SUMB_23__11_), .A2(
        u5_mult_79_CARRYB_23__10_), .ZN(u5_mult_79_n90) );
  AND2_X4 u5_mult_79_U135 ( .A1(u5_mult_79_SUMB_23__13_), .A2(
        u5_mult_79_CARRYB_23__12_), .ZN(u5_mult_79_n89) );
  AND2_X4 u5_mult_79_U134 ( .A1(u5_mult_79_SUMB_23__15_), .A2(
        u5_mult_79_CARRYB_23__14_), .ZN(u5_mult_79_n88) );
  AND2_X4 u5_mult_79_U133 ( .A1(u5_mult_79_SUMB_23__17_), .A2(
        u5_mult_79_CARRYB_23__16_), .ZN(u5_mult_79_n87) );
  AND2_X4 u5_mult_79_U132 ( .A1(u5_mult_79_SUMB_23__19_), .A2(
        u5_mult_79_CARRYB_23__18_), .ZN(u5_mult_79_n86) );
  AND2_X4 u5_mult_79_U131 ( .A1(u5_mult_79_SUMB_23__21_), .A2(
        u5_mult_79_CARRYB_23__20_), .ZN(u5_mult_79_n85) );
  AND2_X4 u5_mult_79_U130 ( .A1(u5_mult_79_SUMB_23__12_), .A2(
        u5_mult_79_CARRYB_23__11_), .ZN(u5_mult_79_n84) );
  AND2_X4 u5_mult_79_U129 ( .A1(u5_mult_79_SUMB_23__14_), .A2(
        u5_mult_79_CARRYB_23__13_), .ZN(u5_mult_79_n83) );
  AND2_X4 u5_mult_79_U128 ( .A1(u5_mult_79_SUMB_23__16_), .A2(
        u5_mult_79_CARRYB_23__15_), .ZN(u5_mult_79_n82) );
  AND2_X4 u5_mult_79_U127 ( .A1(u5_mult_79_SUMB_23__18_), .A2(
        u5_mult_79_CARRYB_23__17_), .ZN(u5_mult_79_n81) );
  AND2_X4 u5_mult_79_U126 ( .A1(u5_mult_79_SUMB_23__20_), .A2(
        u5_mult_79_CARRYB_23__19_), .ZN(u5_mult_79_n80) );
  AND2_X4 u5_mult_79_U125 ( .A1(u5_mult_79_SUMB_23__1_), .A2(
        u5_mult_79_CARRYB_23__0_), .ZN(u5_mult_79_n79) );
  AND2_X4 u5_mult_79_U124 ( .A1(u5_mult_79_SUMB_23__3_), .A2(
        u5_mult_79_CARRYB_23__2_), .ZN(u5_mult_79_n78) );
  AND2_X4 u5_mult_79_U123 ( .A1(u5_mult_79_SUMB_23__5_), .A2(
        u5_mult_79_CARRYB_23__4_), .ZN(u5_mult_79_n77) );
  AND2_X4 u5_mult_79_U122 ( .A1(u5_mult_79_SUMB_23__7_), .A2(
        u5_mult_79_CARRYB_23__6_), .ZN(u5_mult_79_n76) );
  AND2_X4 u5_mult_79_U121 ( .A1(u5_mult_79_SUMB_23__9_), .A2(
        u5_mult_79_CARRYB_23__8_), .ZN(u5_mult_79_n75) );
  AND2_X4 u5_mult_79_U120 ( .A1(u5_mult_79_SUMB_23__2_), .A2(
        u5_mult_79_CARRYB_23__1_), .ZN(u5_mult_79_n74) );
  AND2_X4 u5_mult_79_U119 ( .A1(u5_mult_79_SUMB_23__4_), .A2(
        u5_mult_79_CARRYB_23__3_), .ZN(u5_mult_79_n73) );
  AND2_X4 u5_mult_79_U118 ( .A1(u5_mult_79_SUMB_23__6_), .A2(
        u5_mult_79_CARRYB_23__5_), .ZN(u5_mult_79_n72) );
  AND2_X4 u5_mult_79_U117 ( .A1(u5_mult_79_SUMB_23__8_), .A2(
        u5_mult_79_CARRYB_23__7_), .ZN(u5_mult_79_n71) );
  AND2_X4 u5_mult_79_U116 ( .A1(u5_mult_79_SUMB_23__10_), .A2(
        u5_mult_79_CARRYB_23__9_), .ZN(u5_mult_79_n70) );
  XOR2_X2 u5_mult_79_U115 ( .A(u5_mult_79_ab_1__1_), .B(u5_mult_79_ab_0__2_), 
        .Z(u5_mult_79_n69) );
  XOR2_X2 u5_mult_79_U114 ( .A(u5_mult_79_ab_1__2_), .B(u5_mult_79_ab_0__3_), 
        .Z(u5_mult_79_n68) );
  XOR2_X2 u5_mult_79_U113 ( .A(u5_mult_79_ab_1__3_), .B(u5_mult_79_ab_0__4_), 
        .Z(u5_mult_79_n67) );
  XOR2_X2 u5_mult_79_U112 ( .A(u5_mult_79_ab_1__4_), .B(u5_mult_79_ab_0__5_), 
        .Z(u5_mult_79_n66) );
  XOR2_X2 u5_mult_79_U111 ( .A(u5_mult_79_ab_1__5_), .B(u5_mult_79_ab_0__6_), 
        .Z(u5_mult_79_n65) );
  XOR2_X2 u5_mult_79_U110 ( .A(u5_mult_79_ab_1__6_), .B(u5_mult_79_ab_0__7_), 
        .Z(u5_mult_79_n64) );
  XOR2_X2 u5_mult_79_U109 ( .A(u5_mult_79_ab_1__7_), .B(u5_mult_79_ab_0__8_), 
        .Z(u5_mult_79_n63) );
  XOR2_X2 u5_mult_79_U108 ( .A(u5_mult_79_ab_1__8_), .B(u5_mult_79_ab_0__9_), 
        .Z(u5_mult_79_n62) );
  XOR2_X2 u5_mult_79_U107 ( .A(u5_mult_79_ab_1__9_), .B(u5_mult_79_ab_0__10_), 
        .Z(u5_mult_79_n61) );
  XOR2_X2 u5_mult_79_U106 ( .A(u5_mult_79_ab_1__10_), .B(u5_mult_79_ab_0__11_), 
        .Z(u5_mult_79_n60) );
  XOR2_X2 u5_mult_79_U105 ( .A(u5_mult_79_ab_1__11_), .B(u5_mult_79_ab_0__12_), 
        .Z(u5_mult_79_n59) );
  XOR2_X2 u5_mult_79_U104 ( .A(u5_mult_79_ab_1__12_), .B(u5_mult_79_ab_0__13_), 
        .Z(u5_mult_79_n58) );
  XOR2_X2 u5_mult_79_U103 ( .A(u5_mult_79_ab_1__13_), .B(u5_mult_79_ab_0__14_), 
        .Z(u5_mult_79_n57) );
  XOR2_X2 u5_mult_79_U102 ( .A(u5_mult_79_ab_1__14_), .B(u5_mult_79_ab_0__15_), 
        .Z(u5_mult_79_n56) );
  XOR2_X2 u5_mult_79_U101 ( .A(u5_mult_79_ab_1__15_), .B(u5_mult_79_ab_0__16_), 
        .Z(u5_mult_79_n55) );
  XOR2_X2 u5_mult_79_U100 ( .A(u5_mult_79_ab_1__16_), .B(u5_mult_79_ab_0__17_), 
        .Z(u5_mult_79_n54) );
  XOR2_X2 u5_mult_79_U99 ( .A(u5_mult_79_ab_1__17_), .B(u5_mult_79_ab_0__18_), 
        .Z(u5_mult_79_n53) );
  XOR2_X2 u5_mult_79_U98 ( .A(u5_mult_79_ab_1__18_), .B(u5_mult_79_ab_0__19_), 
        .Z(u5_mult_79_n52) );
  XOR2_X2 u5_mult_79_U97 ( .A(u5_mult_79_ab_1__19_), .B(u5_mult_79_ab_0__20_), 
        .Z(u5_mult_79_n51) );
  XOR2_X2 u5_mult_79_U96 ( .A(u5_mult_79_ab_1__20_), .B(u5_mult_79_ab_0__21_), 
        .Z(u5_mult_79_n50) );
  XOR2_X2 u5_mult_79_U95 ( .A(u5_mult_79_ab_1__21_), .B(u5_mult_79_ab_0__22_), 
        .Z(u5_mult_79_n49) );
  XOR2_X2 u5_mult_79_U94 ( .A(u5_mult_79_ab_1__22_), .B(u5_mult_79_ab_0__23_), 
        .Z(u5_mult_79_n48) );
  AND2_X4 u5_mult_79_U93 ( .A1(u5_mult_79_ab_0__23_), .A2(u5_mult_79_ab_1__22_), .ZN(u5_mult_79_n47) );
  XOR2_X2 u5_mult_79_U92 ( .A(u5_mult_79_CARRYB_23__22_), .B(
        u5_mult_79_ab_23__23_), .Z(u5_mult_79_n46) );
  XOR2_X2 u5_mult_79_U91 ( .A(u5_mult_79_CARRYB_23__13_), .B(
        u5_mult_79_SUMB_23__14_), .Z(u5_mult_79_n45) );
  XOR2_X2 u5_mult_79_U90 ( .A(u5_mult_79_CARRYB_23__15_), .B(
        u5_mult_79_SUMB_23__16_), .Z(u5_mult_79_n44) );
  XOR2_X2 u5_mult_79_U89 ( .A(u5_mult_79_CARRYB_23__17_), .B(
        u5_mult_79_SUMB_23__18_), .Z(u5_mult_79_n43) );
  XOR2_X2 u5_mult_79_U88 ( .A(u5_mult_79_CARRYB_23__19_), .B(
        u5_mult_79_SUMB_23__20_), .Z(u5_mult_79_n42) );
  XOR2_X2 u5_mult_79_U87 ( .A(u5_mult_79_CARRYB_23__21_), .B(
        u5_mult_79_SUMB_23__22_), .Z(u5_mult_79_n41) );
  XOR2_X2 u5_mult_79_U86 ( .A(u5_mult_79_CARRYB_23__12_), .B(
        u5_mult_79_SUMB_23__13_), .Z(u5_mult_79_n40) );
  XOR2_X2 u5_mult_79_U85 ( .A(u5_mult_79_CARRYB_23__14_), .B(
        u5_mult_79_SUMB_23__15_), .Z(u5_mult_79_n39) );
  XOR2_X2 u5_mult_79_U84 ( .A(u5_mult_79_CARRYB_23__16_), .B(
        u5_mult_79_SUMB_23__17_), .Z(u5_mult_79_n38) );
  XOR2_X2 u5_mult_79_U83 ( .A(u5_mult_79_CARRYB_23__18_), .B(
        u5_mult_79_SUMB_23__19_), .Z(u5_mult_79_n37) );
  XOR2_X2 u5_mult_79_U82 ( .A(u5_mult_79_CARRYB_23__20_), .B(
        u5_mult_79_SUMB_23__21_), .Z(u5_mult_79_n36) );
  XOR2_X2 u5_mult_79_U81 ( .A(u5_mult_79_CARRYB_23__3_), .B(
        u5_mult_79_SUMB_23__4_), .Z(u5_mult_79_n35) );
  XOR2_X2 u5_mult_79_U80 ( .A(u5_mult_79_CARRYB_23__5_), .B(
        u5_mult_79_SUMB_23__6_), .Z(u5_mult_79_n34) );
  XOR2_X2 u5_mult_79_U79 ( .A(u5_mult_79_CARRYB_23__7_), .B(
        u5_mult_79_SUMB_23__8_), .Z(u5_mult_79_n33) );
  XOR2_X2 u5_mult_79_U78 ( .A(u5_mult_79_CARRYB_23__9_), .B(
        u5_mult_79_SUMB_23__10_), .Z(u5_mult_79_n32) );
  XOR2_X2 u5_mult_79_U77 ( .A(u5_mult_79_CARRYB_23__11_), .B(
        u5_mult_79_SUMB_23__12_), .Z(u5_mult_79_n31) );
  XOR2_X2 u5_mult_79_U76 ( .A(u5_mult_79_CARRYB_23__1_), .B(
        u5_mult_79_SUMB_23__2_), .Z(u5_mult_79_n30) );
  XOR2_X2 u5_mult_79_U75 ( .A(u5_mult_79_CARRYB_23__2_), .B(
        u5_mult_79_SUMB_23__3_), .Z(u5_mult_79_n29) );
  XOR2_X2 u5_mult_79_U74 ( .A(u5_mult_79_CARRYB_23__4_), .B(
        u5_mult_79_SUMB_23__5_), .Z(u5_mult_79_n28) );
  XOR2_X2 u5_mult_79_U73 ( .A(u5_mult_79_CARRYB_23__6_), .B(
        u5_mult_79_SUMB_23__7_), .Z(u5_mult_79_n27) );
  XOR2_X2 u5_mult_79_U72 ( .A(u5_mult_79_CARRYB_23__8_), .B(
        u5_mult_79_SUMB_23__9_), .Z(u5_mult_79_n26) );
  XOR2_X2 u5_mult_79_U71 ( .A(u5_mult_79_CARRYB_23__10_), .B(
        u5_mult_79_SUMB_23__11_), .Z(u5_mult_79_n25) );
  AND2_X4 u5_mult_79_U70 ( .A1(u5_mult_79_ab_0__1_), .A2(u5_mult_79_ab_1__0_), 
        .ZN(u5_mult_79_n24) );
  AND2_X4 u5_mult_79_U69 ( .A1(u5_mult_79_ab_0__2_), .A2(u5_mult_79_ab_1__1_), 
        .ZN(u5_mult_79_n23) );
  AND2_X4 u5_mult_79_U68 ( .A1(u5_mult_79_ab_0__3_), .A2(u5_mult_79_ab_1__2_), 
        .ZN(u5_mult_79_n22) );
  AND2_X4 u5_mult_79_U67 ( .A1(u5_mult_79_ab_0__4_), .A2(u5_mult_79_ab_1__3_), 
        .ZN(u5_mult_79_n21) );
  AND2_X4 u5_mult_79_U66 ( .A1(u5_mult_79_ab_0__5_), .A2(u5_mult_79_ab_1__4_), 
        .ZN(u5_mult_79_n20) );
  AND2_X4 u5_mult_79_U65 ( .A1(u5_mult_79_ab_0__6_), .A2(u5_mult_79_ab_1__5_), 
        .ZN(u5_mult_79_n19) );
  AND2_X4 u5_mult_79_U64 ( .A1(u5_mult_79_ab_0__7_), .A2(u5_mult_79_ab_1__6_), 
        .ZN(u5_mult_79_n18) );
  AND2_X4 u5_mult_79_U63 ( .A1(u5_mult_79_ab_0__8_), .A2(u5_mult_79_ab_1__7_), 
        .ZN(u5_mult_79_n17) );
  AND2_X4 u5_mult_79_U62 ( .A1(u5_mult_79_ab_0__9_), .A2(u5_mult_79_ab_1__8_), 
        .ZN(u5_mult_79_n16) );
  AND2_X4 u5_mult_79_U61 ( .A1(u5_mult_79_ab_0__10_), .A2(u5_mult_79_ab_1__9_), 
        .ZN(u5_mult_79_n15) );
  AND2_X4 u5_mult_79_U60 ( .A1(u5_mult_79_ab_0__11_), .A2(u5_mult_79_ab_1__10_), .ZN(u5_mult_79_n14) );
  AND2_X4 u5_mult_79_U59 ( .A1(u5_mult_79_ab_0__12_), .A2(u5_mult_79_ab_1__11_), .ZN(u5_mult_79_n13) );
  AND2_X4 u5_mult_79_U58 ( .A1(u5_mult_79_ab_0__13_), .A2(u5_mult_79_ab_1__12_), .ZN(u5_mult_79_n12) );
  AND2_X4 u5_mult_79_U57 ( .A1(u5_mult_79_ab_0__14_), .A2(u5_mult_79_ab_1__13_), .ZN(u5_mult_79_n11) );
  AND2_X4 u5_mult_79_U56 ( .A1(u5_mult_79_ab_0__15_), .A2(u5_mult_79_ab_1__14_), .ZN(u5_mult_79_n10) );
  AND2_X4 u5_mult_79_U55 ( .A1(u5_mult_79_ab_0__16_), .A2(u5_mult_79_ab_1__15_), .ZN(u5_mult_79_n9) );
  AND2_X4 u5_mult_79_U54 ( .A1(u5_mult_79_ab_0__17_), .A2(u5_mult_79_ab_1__16_), .ZN(u5_mult_79_n8) );
  AND2_X4 u5_mult_79_U53 ( .A1(u5_mult_79_ab_0__18_), .A2(u5_mult_79_ab_1__17_), .ZN(u5_mult_79_n7) );
  AND2_X4 u5_mult_79_U52 ( .A1(u5_mult_79_ab_0__19_), .A2(u5_mult_79_ab_1__18_), .ZN(u5_mult_79_n6) );
  AND2_X4 u5_mult_79_U51 ( .A1(u5_mult_79_ab_0__20_), .A2(u5_mult_79_ab_1__19_), .ZN(u5_mult_79_n5) );
  AND2_X4 u5_mult_79_U50 ( .A1(u5_mult_79_ab_0__21_), .A2(u5_mult_79_ab_1__20_), .ZN(u5_mult_79_n4) );
  AND2_X4 u5_mult_79_U49 ( .A1(u5_mult_79_ab_0__22_), .A2(u5_mult_79_ab_1__21_), .ZN(u5_mult_79_n3) );
  INV_X4 u5_mult_79_U48 ( .A(u6_N0), .ZN(u5_mult_79_n142) );
  INV_X4 u5_mult_79_U47 ( .A(fracta_mul[0]), .ZN(u5_mult_79_n118) );
  INV_X4 u5_mult_79_U46 ( .A(fracta_mul[2]), .ZN(u5_mult_79_n116) );
  INV_X4 u5_mult_79_U45 ( .A(fracta_mul[3]), .ZN(u5_mult_79_n115) );
  INV_X4 u5_mult_79_U44 ( .A(fracta_mul[4]), .ZN(u5_mult_79_n114) );
  INV_X4 u5_mult_79_U43 ( .A(fracta_mul[5]), .ZN(u5_mult_79_n113) );
  INV_X4 u5_mult_79_U42 ( .A(fracta_mul[6]), .ZN(u5_mult_79_n112) );
  INV_X4 u5_mult_79_U41 ( .A(fracta_mul[7]), .ZN(u5_mult_79_n111) );
  INV_X4 u5_mult_79_U40 ( .A(fracta_mul[8]), .ZN(u5_mult_79_n110) );
  INV_X4 u5_mult_79_U39 ( .A(fracta_mul[9]), .ZN(u5_mult_79_n109) );
  INV_X4 u5_mult_79_U38 ( .A(fracta_mul[10]), .ZN(u5_mult_79_n108) );
  INV_X4 u5_mult_79_U37 ( .A(fracta_mul[11]), .ZN(u5_mult_79_n107) );
  INV_X4 u5_mult_79_U36 ( .A(fracta_mul[12]), .ZN(u5_mult_79_n106) );
  INV_X4 u5_mult_79_U35 ( .A(fracta_mul[13]), .ZN(u5_mult_79_n105) );
  INV_X4 u5_mult_79_U34 ( .A(fracta_mul[14]), .ZN(u5_mult_79_n104) );
  INV_X4 u5_mult_79_U33 ( .A(fracta_mul[15]), .ZN(u5_mult_79_n103) );
  INV_X4 u5_mult_79_U32 ( .A(fracta_mul[16]), .ZN(u5_mult_79_n102) );
  INV_X4 u5_mult_79_U31 ( .A(fracta_mul[17]), .ZN(u5_mult_79_n101) );
  INV_X4 u5_mult_79_U30 ( .A(fracta_mul[18]), .ZN(u5_mult_79_n100) );
  INV_X4 u5_mult_79_U29 ( .A(fracta_mul[19]), .ZN(u5_mult_79_n99) );
  INV_X4 u5_mult_79_U28 ( .A(fracta_mul[20]), .ZN(u5_mult_79_n98) );
  INV_X4 u5_mult_79_U27 ( .A(fracta_mul[21]), .ZN(u5_mult_79_n97) );
  INV_X4 u5_mult_79_U26 ( .A(fracta_mul[22]), .ZN(u5_mult_79_n96) );
  INV_X4 u5_mult_79_U25 ( .A(u6_N1), .ZN(u5_mult_79_n141) );
  INV_X4 u5_mult_79_U24 ( .A(fracta_mul[1]), .ZN(u5_mult_79_n117) );
  INV_X4 u5_mult_79_U23 ( .A(u6_N2), .ZN(u5_mult_79_n140) );
  INV_X4 u5_mult_79_U22 ( .A(u6_N23), .ZN(u5_mult_79_n119) );
  INV_X4 u5_mult_79_U21 ( .A(u6_N22), .ZN(u5_mult_79_n120) );
  INV_X4 u5_mult_79_U20 ( .A(u6_N3), .ZN(u5_mult_79_n139) );
  INV_X4 u5_mult_79_U19 ( .A(u6_N4), .ZN(u5_mult_79_n138) );
  INV_X4 u5_mult_79_U18 ( .A(u6_N5), .ZN(u5_mult_79_n137) );
  INV_X4 u5_mult_79_U17 ( .A(u6_N6), .ZN(u5_mult_79_n136) );
  INV_X4 u5_mult_79_U16 ( .A(u6_N7), .ZN(u5_mult_79_n135) );
  INV_X4 u5_mult_79_U15 ( .A(u6_N8), .ZN(u5_mult_79_n134) );
  INV_X4 u5_mult_79_U14 ( .A(u6_N9), .ZN(u5_mult_79_n133) );
  INV_X4 u5_mult_79_U13 ( .A(u6_N10), .ZN(u5_mult_79_n132) );
  INV_X4 u5_mult_79_U12 ( .A(u6_N11), .ZN(u5_mult_79_n131) );
  INV_X4 u5_mult_79_U11 ( .A(u6_N12), .ZN(u5_mult_79_n130) );
  INV_X4 u5_mult_79_U10 ( .A(u6_N13), .ZN(u5_mult_79_n129) );
  INV_X4 u5_mult_79_U9 ( .A(u6_N14), .ZN(u5_mult_79_n128) );
  INV_X4 u5_mult_79_U8 ( .A(u6_N15), .ZN(u5_mult_79_n127) );
  INV_X4 u5_mult_79_U7 ( .A(u6_N16), .ZN(u5_mult_79_n126) );
  INV_X4 u5_mult_79_U6 ( .A(u6_N17), .ZN(u5_mult_79_n125) );
  INV_X4 u5_mult_79_U5 ( .A(u6_N18), .ZN(u5_mult_79_n124) );
  INV_X4 u5_mult_79_U4 ( .A(u6_N19), .ZN(u5_mult_79_n123) );
  INV_X4 u5_mult_79_U3 ( .A(u6_N20), .ZN(u5_mult_79_n122) );
  INV_X4 u5_mult_79_U2 ( .A(u6_N21), .ZN(u5_mult_79_n121) );
  FA_X1 u5_mult_79_S3_2_22 ( .A(u5_mult_79_ab_2__22_), .B(u5_mult_79_n47), 
        .CI(u5_mult_79_ab_1__23_), .CO(u5_mult_79_CARRYB_2__22_), .S(
        u5_mult_79_SUMB_2__22_) );
  FA_X1 u5_mult_79_S2_2_21 ( .A(u5_mult_79_ab_2__21_), .B(u5_mult_79_n3), .CI(
        u5_mult_79_n48), .CO(u5_mult_79_CARRYB_2__21_), .S(
        u5_mult_79_SUMB_2__21_) );
  FA_X1 u5_mult_79_S2_2_20 ( .A(u5_mult_79_ab_2__20_), .B(u5_mult_79_n4), .CI(
        u5_mult_79_n49), .CO(u5_mult_79_CARRYB_2__20_), .S(
        u5_mult_79_SUMB_2__20_) );
  FA_X1 u5_mult_79_S2_2_19 ( .A(u5_mult_79_ab_2__19_), .B(u5_mult_79_n5), .CI(
        u5_mult_79_n50), .CO(u5_mult_79_CARRYB_2__19_), .S(
        u5_mult_79_SUMB_2__19_) );
  FA_X1 u5_mult_79_S2_2_18 ( .A(u5_mult_79_ab_2__18_), .B(u5_mult_79_n6), .CI(
        u5_mult_79_n51), .CO(u5_mult_79_CARRYB_2__18_), .S(
        u5_mult_79_SUMB_2__18_) );
  FA_X1 u5_mult_79_S2_2_17 ( .A(u5_mult_79_ab_2__17_), .B(u5_mult_79_n7), .CI(
        u5_mult_79_n52), .CO(u5_mult_79_CARRYB_2__17_), .S(
        u5_mult_79_SUMB_2__17_) );
  FA_X1 u5_mult_79_S2_2_16 ( .A(u5_mult_79_ab_2__16_), .B(u5_mult_79_n8), .CI(
        u5_mult_79_n53), .CO(u5_mult_79_CARRYB_2__16_), .S(
        u5_mult_79_SUMB_2__16_) );
  FA_X1 u5_mult_79_S2_2_15 ( .A(u5_mult_79_ab_2__15_), .B(u5_mult_79_n9), .CI(
        u5_mult_79_n54), .CO(u5_mult_79_CARRYB_2__15_), .S(
        u5_mult_79_SUMB_2__15_) );
  FA_X1 u5_mult_79_S2_2_14 ( .A(u5_mult_79_ab_2__14_), .B(u5_mult_79_n10), 
        .CI(u5_mult_79_n55), .CO(u5_mult_79_CARRYB_2__14_), .S(
        u5_mult_79_SUMB_2__14_) );
  FA_X1 u5_mult_79_S2_2_13 ( .A(u5_mult_79_ab_2__13_), .B(u5_mult_79_n11), 
        .CI(u5_mult_79_n56), .CO(u5_mult_79_CARRYB_2__13_), .S(
        u5_mult_79_SUMB_2__13_) );
  FA_X1 u5_mult_79_S2_2_12 ( .A(u5_mult_79_ab_2__12_), .B(u5_mult_79_n12), 
        .CI(u5_mult_79_n57), .CO(u5_mult_79_CARRYB_2__12_), .S(
        u5_mult_79_SUMB_2__12_) );
  FA_X1 u5_mult_79_S2_2_11 ( .A(u5_mult_79_ab_2__11_), .B(u5_mult_79_n13), 
        .CI(u5_mult_79_n58), .CO(u5_mult_79_CARRYB_2__11_), .S(
        u5_mult_79_SUMB_2__11_) );
  FA_X1 u5_mult_79_S2_2_10 ( .A(u5_mult_79_ab_2__10_), .B(u5_mult_79_n14), 
        .CI(u5_mult_79_n59), .CO(u5_mult_79_CARRYB_2__10_), .S(
        u5_mult_79_SUMB_2__10_) );
  FA_X1 u5_mult_79_S2_2_9 ( .A(u5_mult_79_ab_2__9_), .B(u5_mult_79_n15), .CI(
        u5_mult_79_n60), .CO(u5_mult_79_CARRYB_2__9_), .S(
        u5_mult_79_SUMB_2__9_) );
  FA_X1 u5_mult_79_S2_2_8 ( .A(u5_mult_79_ab_2__8_), .B(u5_mult_79_n16), .CI(
        u5_mult_79_n61), .CO(u5_mult_79_CARRYB_2__8_), .S(
        u5_mult_79_SUMB_2__8_) );
  FA_X1 u5_mult_79_S2_2_7 ( .A(u5_mult_79_ab_2__7_), .B(u5_mult_79_n17), .CI(
        u5_mult_79_n62), .CO(u5_mult_79_CARRYB_2__7_), .S(
        u5_mult_79_SUMB_2__7_) );
  FA_X1 u5_mult_79_S2_2_6 ( .A(u5_mult_79_ab_2__6_), .B(u5_mult_79_n18), .CI(
        u5_mult_79_n63), .CO(u5_mult_79_CARRYB_2__6_), .S(
        u5_mult_79_SUMB_2__6_) );
  FA_X1 u5_mult_79_S2_2_5 ( .A(u5_mult_79_ab_2__5_), .B(u5_mult_79_n19), .CI(
        u5_mult_79_n64), .CO(u5_mult_79_CARRYB_2__5_), .S(
        u5_mult_79_SUMB_2__5_) );
  FA_X1 u5_mult_79_S2_2_4 ( .A(u5_mult_79_ab_2__4_), .B(u5_mult_79_n20), .CI(
        u5_mult_79_n65), .CO(u5_mult_79_CARRYB_2__4_), .S(
        u5_mult_79_SUMB_2__4_) );
  FA_X1 u5_mult_79_S2_2_3 ( .A(u5_mult_79_ab_2__3_), .B(u5_mult_79_n21), .CI(
        u5_mult_79_n66), .CO(u5_mult_79_CARRYB_2__3_), .S(
        u5_mult_79_SUMB_2__3_) );
  FA_X1 u5_mult_79_S2_2_2 ( .A(u5_mult_79_ab_2__2_), .B(u5_mult_79_n22), .CI(
        u5_mult_79_n67), .CO(u5_mult_79_CARRYB_2__2_), .S(
        u5_mult_79_SUMB_2__2_) );
  FA_X1 u5_mult_79_S2_2_1 ( .A(u5_mult_79_ab_2__1_), .B(u5_mult_79_n23), .CI(
        u5_mult_79_n68), .CO(u5_mult_79_CARRYB_2__1_), .S(
        u5_mult_79_SUMB_2__1_) );
  FA_X1 u5_mult_79_S1_2_0 ( .A(u5_mult_79_ab_2__0_), .B(u5_mult_79_n24), .CI(
        u5_mult_79_n69), .CO(u5_mult_79_CARRYB_2__0_), .S(u5_N2) );
  FA_X1 u5_mult_79_S3_3_22 ( .A(u5_mult_79_ab_3__22_), .B(
        u5_mult_79_CARRYB_2__22_), .CI(u5_mult_79_ab_2__23_), .CO(
        u5_mult_79_CARRYB_3__22_), .S(u5_mult_79_SUMB_3__22_) );
  FA_X1 u5_mult_79_S2_3_21 ( .A(u5_mult_79_ab_3__21_), .B(
        u5_mult_79_CARRYB_2__21_), .CI(u5_mult_79_SUMB_2__22_), .CO(
        u5_mult_79_CARRYB_3__21_), .S(u5_mult_79_SUMB_3__21_) );
  FA_X1 u5_mult_79_S2_3_20 ( .A(u5_mult_79_ab_3__20_), .B(
        u5_mult_79_CARRYB_2__20_), .CI(u5_mult_79_SUMB_2__21_), .CO(
        u5_mult_79_CARRYB_3__20_), .S(u5_mult_79_SUMB_3__20_) );
  FA_X1 u5_mult_79_S2_3_19 ( .A(u5_mult_79_ab_3__19_), .B(
        u5_mult_79_CARRYB_2__19_), .CI(u5_mult_79_SUMB_2__20_), .CO(
        u5_mult_79_CARRYB_3__19_), .S(u5_mult_79_SUMB_3__19_) );
  FA_X1 u5_mult_79_S2_3_18 ( .A(u5_mult_79_ab_3__18_), .B(
        u5_mult_79_CARRYB_2__18_), .CI(u5_mult_79_SUMB_2__19_), .CO(
        u5_mult_79_CARRYB_3__18_), .S(u5_mult_79_SUMB_3__18_) );
  FA_X1 u5_mult_79_S2_3_17 ( .A(u5_mult_79_ab_3__17_), .B(
        u5_mult_79_CARRYB_2__17_), .CI(u5_mult_79_SUMB_2__18_), .CO(
        u5_mult_79_CARRYB_3__17_), .S(u5_mult_79_SUMB_3__17_) );
  FA_X1 u5_mult_79_S2_3_16 ( .A(u5_mult_79_ab_3__16_), .B(
        u5_mult_79_CARRYB_2__16_), .CI(u5_mult_79_SUMB_2__17_), .CO(
        u5_mult_79_CARRYB_3__16_), .S(u5_mult_79_SUMB_3__16_) );
  FA_X1 u5_mult_79_S2_3_15 ( .A(u5_mult_79_ab_3__15_), .B(
        u5_mult_79_CARRYB_2__15_), .CI(u5_mult_79_SUMB_2__16_), .CO(
        u5_mult_79_CARRYB_3__15_), .S(u5_mult_79_SUMB_3__15_) );
  FA_X1 u5_mult_79_S2_3_14 ( .A(u5_mult_79_ab_3__14_), .B(
        u5_mult_79_CARRYB_2__14_), .CI(u5_mult_79_SUMB_2__15_), .CO(
        u5_mult_79_CARRYB_3__14_), .S(u5_mult_79_SUMB_3__14_) );
  FA_X1 u5_mult_79_S2_3_13 ( .A(u5_mult_79_ab_3__13_), .B(
        u5_mult_79_CARRYB_2__13_), .CI(u5_mult_79_SUMB_2__14_), .CO(
        u5_mult_79_CARRYB_3__13_), .S(u5_mult_79_SUMB_3__13_) );
  FA_X1 u5_mult_79_S2_3_12 ( .A(u5_mult_79_ab_3__12_), .B(
        u5_mult_79_CARRYB_2__12_), .CI(u5_mult_79_SUMB_2__13_), .CO(
        u5_mult_79_CARRYB_3__12_), .S(u5_mult_79_SUMB_3__12_) );
  FA_X1 u5_mult_79_S2_3_11 ( .A(u5_mult_79_ab_3__11_), .B(
        u5_mult_79_CARRYB_2__11_), .CI(u5_mult_79_SUMB_2__12_), .CO(
        u5_mult_79_CARRYB_3__11_), .S(u5_mult_79_SUMB_3__11_) );
  FA_X1 u5_mult_79_S2_3_10 ( .A(u5_mult_79_ab_3__10_), .B(
        u5_mult_79_CARRYB_2__10_), .CI(u5_mult_79_SUMB_2__11_), .CO(
        u5_mult_79_CARRYB_3__10_), .S(u5_mult_79_SUMB_3__10_) );
  FA_X1 u5_mult_79_S2_3_9 ( .A(u5_mult_79_ab_3__9_), .B(
        u5_mult_79_CARRYB_2__9_), .CI(u5_mult_79_SUMB_2__10_), .CO(
        u5_mult_79_CARRYB_3__9_), .S(u5_mult_79_SUMB_3__9_) );
  FA_X1 u5_mult_79_S2_3_8 ( .A(u5_mult_79_ab_3__8_), .B(
        u5_mult_79_CARRYB_2__8_), .CI(u5_mult_79_SUMB_2__9_), .CO(
        u5_mult_79_CARRYB_3__8_), .S(u5_mult_79_SUMB_3__8_) );
  FA_X1 u5_mult_79_S2_3_7 ( .A(u5_mult_79_ab_3__7_), .B(
        u5_mult_79_CARRYB_2__7_), .CI(u5_mult_79_SUMB_2__8_), .CO(
        u5_mult_79_CARRYB_3__7_), .S(u5_mult_79_SUMB_3__7_) );
  FA_X1 u5_mult_79_S2_3_6 ( .A(u5_mult_79_ab_3__6_), .B(
        u5_mult_79_CARRYB_2__6_), .CI(u5_mult_79_SUMB_2__7_), .CO(
        u5_mult_79_CARRYB_3__6_), .S(u5_mult_79_SUMB_3__6_) );
  FA_X1 u5_mult_79_S2_3_5 ( .A(u5_mult_79_ab_3__5_), .B(
        u5_mult_79_CARRYB_2__5_), .CI(u5_mult_79_SUMB_2__6_), .CO(
        u5_mult_79_CARRYB_3__5_), .S(u5_mult_79_SUMB_3__5_) );
  FA_X1 u5_mult_79_S2_3_4 ( .A(u5_mult_79_ab_3__4_), .B(
        u5_mult_79_CARRYB_2__4_), .CI(u5_mult_79_SUMB_2__5_), .CO(
        u5_mult_79_CARRYB_3__4_), .S(u5_mult_79_SUMB_3__4_) );
  FA_X1 u5_mult_79_S2_3_3 ( .A(u5_mult_79_ab_3__3_), .B(
        u5_mult_79_CARRYB_2__3_), .CI(u5_mult_79_SUMB_2__4_), .CO(
        u5_mult_79_CARRYB_3__3_), .S(u5_mult_79_SUMB_3__3_) );
  FA_X1 u5_mult_79_S2_3_2 ( .A(u5_mult_79_ab_3__2_), .B(
        u5_mult_79_CARRYB_2__2_), .CI(u5_mult_79_SUMB_2__3_), .CO(
        u5_mult_79_CARRYB_3__2_), .S(u5_mult_79_SUMB_3__2_) );
  FA_X1 u5_mult_79_S2_3_1 ( .A(u5_mult_79_ab_3__1_), .B(
        u5_mult_79_CARRYB_2__1_), .CI(u5_mult_79_SUMB_2__2_), .CO(
        u5_mult_79_CARRYB_3__1_), .S(u5_mult_79_SUMB_3__1_) );
  FA_X1 u5_mult_79_S1_3_0 ( .A(u5_mult_79_ab_3__0_), .B(
        u5_mult_79_CARRYB_2__0_), .CI(u5_mult_79_SUMB_2__1_), .CO(
        u5_mult_79_CARRYB_3__0_), .S(u5_N3) );
  FA_X1 u5_mult_79_S3_4_22 ( .A(u5_mult_79_ab_4__22_), .B(
        u5_mult_79_CARRYB_3__22_), .CI(u5_mult_79_ab_3__23_), .CO(
        u5_mult_79_CARRYB_4__22_), .S(u5_mult_79_SUMB_4__22_) );
  FA_X1 u5_mult_79_S2_4_21 ( .A(u5_mult_79_ab_4__21_), .B(
        u5_mult_79_CARRYB_3__21_), .CI(u5_mult_79_SUMB_3__22_), .CO(
        u5_mult_79_CARRYB_4__21_), .S(u5_mult_79_SUMB_4__21_) );
  FA_X1 u5_mult_79_S2_4_20 ( .A(u5_mult_79_ab_4__20_), .B(
        u5_mult_79_CARRYB_3__20_), .CI(u5_mult_79_SUMB_3__21_), .CO(
        u5_mult_79_CARRYB_4__20_), .S(u5_mult_79_SUMB_4__20_) );
  FA_X1 u5_mult_79_S2_4_19 ( .A(u5_mult_79_ab_4__19_), .B(
        u5_mult_79_CARRYB_3__19_), .CI(u5_mult_79_SUMB_3__20_), .CO(
        u5_mult_79_CARRYB_4__19_), .S(u5_mult_79_SUMB_4__19_) );
  FA_X1 u5_mult_79_S2_4_18 ( .A(u5_mult_79_ab_4__18_), .B(
        u5_mult_79_CARRYB_3__18_), .CI(u5_mult_79_SUMB_3__19_), .CO(
        u5_mult_79_CARRYB_4__18_), .S(u5_mult_79_SUMB_4__18_) );
  FA_X1 u5_mult_79_S2_4_17 ( .A(u5_mult_79_ab_4__17_), .B(
        u5_mult_79_CARRYB_3__17_), .CI(u5_mult_79_SUMB_3__18_), .CO(
        u5_mult_79_CARRYB_4__17_), .S(u5_mult_79_SUMB_4__17_) );
  FA_X1 u5_mult_79_S2_4_16 ( .A(u5_mult_79_ab_4__16_), .B(
        u5_mult_79_CARRYB_3__16_), .CI(u5_mult_79_SUMB_3__17_), .CO(
        u5_mult_79_CARRYB_4__16_), .S(u5_mult_79_SUMB_4__16_) );
  FA_X1 u5_mult_79_S2_4_15 ( .A(u5_mult_79_ab_4__15_), .B(
        u5_mult_79_CARRYB_3__15_), .CI(u5_mult_79_SUMB_3__16_), .CO(
        u5_mult_79_CARRYB_4__15_), .S(u5_mult_79_SUMB_4__15_) );
  FA_X1 u5_mult_79_S2_4_14 ( .A(u5_mult_79_ab_4__14_), .B(
        u5_mult_79_CARRYB_3__14_), .CI(u5_mult_79_SUMB_3__15_), .CO(
        u5_mult_79_CARRYB_4__14_), .S(u5_mult_79_SUMB_4__14_) );
  FA_X1 u5_mult_79_S2_4_13 ( .A(u5_mult_79_ab_4__13_), .B(
        u5_mult_79_CARRYB_3__13_), .CI(u5_mult_79_SUMB_3__14_), .CO(
        u5_mult_79_CARRYB_4__13_), .S(u5_mult_79_SUMB_4__13_) );
  FA_X1 u5_mult_79_S2_4_12 ( .A(u5_mult_79_ab_4__12_), .B(
        u5_mult_79_CARRYB_3__12_), .CI(u5_mult_79_SUMB_3__13_), .CO(
        u5_mult_79_CARRYB_4__12_), .S(u5_mult_79_SUMB_4__12_) );
  FA_X1 u5_mult_79_S2_4_11 ( .A(u5_mult_79_ab_4__11_), .B(
        u5_mult_79_CARRYB_3__11_), .CI(u5_mult_79_SUMB_3__12_), .CO(
        u5_mult_79_CARRYB_4__11_), .S(u5_mult_79_SUMB_4__11_) );
  FA_X1 u5_mult_79_S2_4_10 ( .A(u5_mult_79_ab_4__10_), .B(
        u5_mult_79_CARRYB_3__10_), .CI(u5_mult_79_SUMB_3__11_), .CO(
        u5_mult_79_CARRYB_4__10_), .S(u5_mult_79_SUMB_4__10_) );
  FA_X1 u5_mult_79_S2_4_9 ( .A(u5_mult_79_ab_4__9_), .B(
        u5_mult_79_CARRYB_3__9_), .CI(u5_mult_79_SUMB_3__10_), .CO(
        u5_mult_79_CARRYB_4__9_), .S(u5_mult_79_SUMB_4__9_) );
  FA_X1 u5_mult_79_S2_4_8 ( .A(u5_mult_79_ab_4__8_), .B(
        u5_mult_79_CARRYB_3__8_), .CI(u5_mult_79_SUMB_3__9_), .CO(
        u5_mult_79_CARRYB_4__8_), .S(u5_mult_79_SUMB_4__8_) );
  FA_X1 u5_mult_79_S2_4_7 ( .A(u5_mult_79_ab_4__7_), .B(
        u5_mult_79_CARRYB_3__7_), .CI(u5_mult_79_SUMB_3__8_), .CO(
        u5_mult_79_CARRYB_4__7_), .S(u5_mult_79_SUMB_4__7_) );
  FA_X1 u5_mult_79_S2_4_6 ( .A(u5_mult_79_ab_4__6_), .B(
        u5_mult_79_CARRYB_3__6_), .CI(u5_mult_79_SUMB_3__7_), .CO(
        u5_mult_79_CARRYB_4__6_), .S(u5_mult_79_SUMB_4__6_) );
  FA_X1 u5_mult_79_S2_4_5 ( .A(u5_mult_79_ab_4__5_), .B(
        u5_mult_79_CARRYB_3__5_), .CI(u5_mult_79_SUMB_3__6_), .CO(
        u5_mult_79_CARRYB_4__5_), .S(u5_mult_79_SUMB_4__5_) );
  FA_X1 u5_mult_79_S2_4_4 ( .A(u5_mult_79_ab_4__4_), .B(
        u5_mult_79_CARRYB_3__4_), .CI(u5_mult_79_SUMB_3__5_), .CO(
        u5_mult_79_CARRYB_4__4_), .S(u5_mult_79_SUMB_4__4_) );
  FA_X1 u5_mult_79_S2_4_3 ( .A(u5_mult_79_ab_4__3_), .B(
        u5_mult_79_CARRYB_3__3_), .CI(u5_mult_79_SUMB_3__4_), .CO(
        u5_mult_79_CARRYB_4__3_), .S(u5_mult_79_SUMB_4__3_) );
  FA_X1 u5_mult_79_S2_4_2 ( .A(u5_mult_79_ab_4__2_), .B(
        u5_mult_79_CARRYB_3__2_), .CI(u5_mult_79_SUMB_3__3_), .CO(
        u5_mult_79_CARRYB_4__2_), .S(u5_mult_79_SUMB_4__2_) );
  FA_X1 u5_mult_79_S2_4_1 ( .A(u5_mult_79_ab_4__1_), .B(
        u5_mult_79_CARRYB_3__1_), .CI(u5_mult_79_SUMB_3__2_), .CO(
        u5_mult_79_CARRYB_4__1_), .S(u5_mult_79_SUMB_4__1_) );
  FA_X1 u5_mult_79_S1_4_0 ( .A(u5_mult_79_ab_4__0_), .B(
        u5_mult_79_CARRYB_3__0_), .CI(u5_mult_79_SUMB_3__1_), .CO(
        u5_mult_79_CARRYB_4__0_), .S(u5_N4) );
  FA_X1 u5_mult_79_S3_5_22 ( .A(u5_mult_79_ab_5__22_), .B(
        u5_mult_79_CARRYB_4__22_), .CI(u5_mult_79_ab_4__23_), .CO(
        u5_mult_79_CARRYB_5__22_), .S(u5_mult_79_SUMB_5__22_) );
  FA_X1 u5_mult_79_S2_5_21 ( .A(u5_mult_79_ab_5__21_), .B(
        u5_mult_79_CARRYB_4__21_), .CI(u5_mult_79_SUMB_4__22_), .CO(
        u5_mult_79_CARRYB_5__21_), .S(u5_mult_79_SUMB_5__21_) );
  FA_X1 u5_mult_79_S2_5_20 ( .A(u5_mult_79_ab_5__20_), .B(
        u5_mult_79_CARRYB_4__20_), .CI(u5_mult_79_SUMB_4__21_), .CO(
        u5_mult_79_CARRYB_5__20_), .S(u5_mult_79_SUMB_5__20_) );
  FA_X1 u5_mult_79_S2_5_19 ( .A(u5_mult_79_ab_5__19_), .B(
        u5_mult_79_CARRYB_4__19_), .CI(u5_mult_79_SUMB_4__20_), .CO(
        u5_mult_79_CARRYB_5__19_), .S(u5_mult_79_SUMB_5__19_) );
  FA_X1 u5_mult_79_S2_5_18 ( .A(u5_mult_79_ab_5__18_), .B(
        u5_mult_79_CARRYB_4__18_), .CI(u5_mult_79_SUMB_4__19_), .CO(
        u5_mult_79_CARRYB_5__18_), .S(u5_mult_79_SUMB_5__18_) );
  FA_X1 u5_mult_79_S2_5_17 ( .A(u5_mult_79_ab_5__17_), .B(
        u5_mult_79_CARRYB_4__17_), .CI(u5_mult_79_SUMB_4__18_), .CO(
        u5_mult_79_CARRYB_5__17_), .S(u5_mult_79_SUMB_5__17_) );
  FA_X1 u5_mult_79_S2_5_16 ( .A(u5_mult_79_ab_5__16_), .B(
        u5_mult_79_CARRYB_4__16_), .CI(u5_mult_79_SUMB_4__17_), .CO(
        u5_mult_79_CARRYB_5__16_), .S(u5_mult_79_SUMB_5__16_) );
  FA_X1 u5_mult_79_S2_5_15 ( .A(u5_mult_79_ab_5__15_), .B(
        u5_mult_79_CARRYB_4__15_), .CI(u5_mult_79_SUMB_4__16_), .CO(
        u5_mult_79_CARRYB_5__15_), .S(u5_mult_79_SUMB_5__15_) );
  FA_X1 u5_mult_79_S2_5_14 ( .A(u5_mult_79_ab_5__14_), .B(
        u5_mult_79_CARRYB_4__14_), .CI(u5_mult_79_SUMB_4__15_), .CO(
        u5_mult_79_CARRYB_5__14_), .S(u5_mult_79_SUMB_5__14_) );
  FA_X1 u5_mult_79_S2_5_13 ( .A(u5_mult_79_ab_5__13_), .B(
        u5_mult_79_CARRYB_4__13_), .CI(u5_mult_79_SUMB_4__14_), .CO(
        u5_mult_79_CARRYB_5__13_), .S(u5_mult_79_SUMB_5__13_) );
  FA_X1 u5_mult_79_S2_5_12 ( .A(u5_mult_79_ab_5__12_), .B(
        u5_mult_79_CARRYB_4__12_), .CI(u5_mult_79_SUMB_4__13_), .CO(
        u5_mult_79_CARRYB_5__12_), .S(u5_mult_79_SUMB_5__12_) );
  FA_X1 u5_mult_79_S2_5_11 ( .A(u5_mult_79_ab_5__11_), .B(
        u5_mult_79_CARRYB_4__11_), .CI(u5_mult_79_SUMB_4__12_), .CO(
        u5_mult_79_CARRYB_5__11_), .S(u5_mult_79_SUMB_5__11_) );
  FA_X1 u5_mult_79_S2_5_10 ( .A(u5_mult_79_ab_5__10_), .B(
        u5_mult_79_CARRYB_4__10_), .CI(u5_mult_79_SUMB_4__11_), .CO(
        u5_mult_79_CARRYB_5__10_), .S(u5_mult_79_SUMB_5__10_) );
  FA_X1 u5_mult_79_S2_5_9 ( .A(u5_mult_79_ab_5__9_), .B(
        u5_mult_79_CARRYB_4__9_), .CI(u5_mult_79_SUMB_4__10_), .CO(
        u5_mult_79_CARRYB_5__9_), .S(u5_mult_79_SUMB_5__9_) );
  FA_X1 u5_mult_79_S2_5_8 ( .A(u5_mult_79_ab_5__8_), .B(
        u5_mult_79_CARRYB_4__8_), .CI(u5_mult_79_SUMB_4__9_), .CO(
        u5_mult_79_CARRYB_5__8_), .S(u5_mult_79_SUMB_5__8_) );
  FA_X1 u5_mult_79_S2_5_7 ( .A(u5_mult_79_ab_5__7_), .B(
        u5_mult_79_CARRYB_4__7_), .CI(u5_mult_79_SUMB_4__8_), .CO(
        u5_mult_79_CARRYB_5__7_), .S(u5_mult_79_SUMB_5__7_) );
  FA_X1 u5_mult_79_S2_5_6 ( .A(u5_mult_79_ab_5__6_), .B(
        u5_mult_79_CARRYB_4__6_), .CI(u5_mult_79_SUMB_4__7_), .CO(
        u5_mult_79_CARRYB_5__6_), .S(u5_mult_79_SUMB_5__6_) );
  FA_X1 u5_mult_79_S2_5_5 ( .A(u5_mult_79_ab_5__5_), .B(
        u5_mult_79_CARRYB_4__5_), .CI(u5_mult_79_SUMB_4__6_), .CO(
        u5_mult_79_CARRYB_5__5_), .S(u5_mult_79_SUMB_5__5_) );
  FA_X1 u5_mult_79_S2_5_4 ( .A(u5_mult_79_ab_5__4_), .B(
        u5_mult_79_CARRYB_4__4_), .CI(u5_mult_79_SUMB_4__5_), .CO(
        u5_mult_79_CARRYB_5__4_), .S(u5_mult_79_SUMB_5__4_) );
  FA_X1 u5_mult_79_S2_5_3 ( .A(u5_mult_79_ab_5__3_), .B(
        u5_mult_79_CARRYB_4__3_), .CI(u5_mult_79_SUMB_4__4_), .CO(
        u5_mult_79_CARRYB_5__3_), .S(u5_mult_79_SUMB_5__3_) );
  FA_X1 u5_mult_79_S2_5_2 ( .A(u5_mult_79_ab_5__2_), .B(
        u5_mult_79_CARRYB_4__2_), .CI(u5_mult_79_SUMB_4__3_), .CO(
        u5_mult_79_CARRYB_5__2_), .S(u5_mult_79_SUMB_5__2_) );
  FA_X1 u5_mult_79_S2_5_1 ( .A(u5_mult_79_ab_5__1_), .B(
        u5_mult_79_CARRYB_4__1_), .CI(u5_mult_79_SUMB_4__2_), .CO(
        u5_mult_79_CARRYB_5__1_), .S(u5_mult_79_SUMB_5__1_) );
  FA_X1 u5_mult_79_S1_5_0 ( .A(u5_mult_79_ab_5__0_), .B(
        u5_mult_79_CARRYB_4__0_), .CI(u5_mult_79_SUMB_4__1_), .CO(
        u5_mult_79_CARRYB_5__0_), .S(u5_N5) );
  FA_X1 u5_mult_79_S3_6_22 ( .A(u5_mult_79_ab_6__22_), .B(
        u5_mult_79_CARRYB_5__22_), .CI(u5_mult_79_ab_5__23_), .CO(
        u5_mult_79_CARRYB_6__22_), .S(u5_mult_79_SUMB_6__22_) );
  FA_X1 u5_mult_79_S2_6_21 ( .A(u5_mult_79_ab_6__21_), .B(
        u5_mult_79_CARRYB_5__21_), .CI(u5_mult_79_SUMB_5__22_), .CO(
        u5_mult_79_CARRYB_6__21_), .S(u5_mult_79_SUMB_6__21_) );
  FA_X1 u5_mult_79_S2_6_20 ( .A(u5_mult_79_ab_6__20_), .B(
        u5_mult_79_CARRYB_5__20_), .CI(u5_mult_79_SUMB_5__21_), .CO(
        u5_mult_79_CARRYB_6__20_), .S(u5_mult_79_SUMB_6__20_) );
  FA_X1 u5_mult_79_S2_6_19 ( .A(u5_mult_79_ab_6__19_), .B(
        u5_mult_79_CARRYB_5__19_), .CI(u5_mult_79_SUMB_5__20_), .CO(
        u5_mult_79_CARRYB_6__19_), .S(u5_mult_79_SUMB_6__19_) );
  FA_X1 u5_mult_79_S2_6_18 ( .A(u5_mult_79_ab_6__18_), .B(
        u5_mult_79_CARRYB_5__18_), .CI(u5_mult_79_SUMB_5__19_), .CO(
        u5_mult_79_CARRYB_6__18_), .S(u5_mult_79_SUMB_6__18_) );
  FA_X1 u5_mult_79_S2_6_17 ( .A(u5_mult_79_ab_6__17_), .B(
        u5_mult_79_CARRYB_5__17_), .CI(u5_mult_79_SUMB_5__18_), .CO(
        u5_mult_79_CARRYB_6__17_), .S(u5_mult_79_SUMB_6__17_) );
  FA_X1 u5_mult_79_S2_6_16 ( .A(u5_mult_79_ab_6__16_), .B(
        u5_mult_79_CARRYB_5__16_), .CI(u5_mult_79_SUMB_5__17_), .CO(
        u5_mult_79_CARRYB_6__16_), .S(u5_mult_79_SUMB_6__16_) );
  FA_X1 u5_mult_79_S2_6_15 ( .A(u5_mult_79_ab_6__15_), .B(
        u5_mult_79_CARRYB_5__15_), .CI(u5_mult_79_SUMB_5__16_), .CO(
        u5_mult_79_CARRYB_6__15_), .S(u5_mult_79_SUMB_6__15_) );
  FA_X1 u5_mult_79_S2_6_14 ( .A(u5_mult_79_ab_6__14_), .B(
        u5_mult_79_CARRYB_5__14_), .CI(u5_mult_79_SUMB_5__15_), .CO(
        u5_mult_79_CARRYB_6__14_), .S(u5_mult_79_SUMB_6__14_) );
  FA_X1 u5_mult_79_S2_6_13 ( .A(u5_mult_79_ab_6__13_), .B(
        u5_mult_79_CARRYB_5__13_), .CI(u5_mult_79_SUMB_5__14_), .CO(
        u5_mult_79_CARRYB_6__13_), .S(u5_mult_79_SUMB_6__13_) );
  FA_X1 u5_mult_79_S2_6_12 ( .A(u5_mult_79_ab_6__12_), .B(
        u5_mult_79_CARRYB_5__12_), .CI(u5_mult_79_SUMB_5__13_), .CO(
        u5_mult_79_CARRYB_6__12_), .S(u5_mult_79_SUMB_6__12_) );
  FA_X1 u5_mult_79_S2_6_11 ( .A(u5_mult_79_ab_6__11_), .B(
        u5_mult_79_CARRYB_5__11_), .CI(u5_mult_79_SUMB_5__12_), .CO(
        u5_mult_79_CARRYB_6__11_), .S(u5_mult_79_SUMB_6__11_) );
  FA_X1 u5_mult_79_S2_6_10 ( .A(u5_mult_79_ab_6__10_), .B(
        u5_mult_79_CARRYB_5__10_), .CI(u5_mult_79_SUMB_5__11_), .CO(
        u5_mult_79_CARRYB_6__10_), .S(u5_mult_79_SUMB_6__10_) );
  FA_X1 u5_mult_79_S2_6_9 ( .A(u5_mult_79_ab_6__9_), .B(
        u5_mult_79_CARRYB_5__9_), .CI(u5_mult_79_SUMB_5__10_), .CO(
        u5_mult_79_CARRYB_6__9_), .S(u5_mult_79_SUMB_6__9_) );
  FA_X1 u5_mult_79_S2_6_8 ( .A(u5_mult_79_ab_6__8_), .B(
        u5_mult_79_CARRYB_5__8_), .CI(u5_mult_79_SUMB_5__9_), .CO(
        u5_mult_79_CARRYB_6__8_), .S(u5_mult_79_SUMB_6__8_) );
  FA_X1 u5_mult_79_S2_6_7 ( .A(u5_mult_79_ab_6__7_), .B(
        u5_mult_79_CARRYB_5__7_), .CI(u5_mult_79_SUMB_5__8_), .CO(
        u5_mult_79_CARRYB_6__7_), .S(u5_mult_79_SUMB_6__7_) );
  FA_X1 u5_mult_79_S2_6_6 ( .A(u5_mult_79_ab_6__6_), .B(
        u5_mult_79_CARRYB_5__6_), .CI(u5_mult_79_SUMB_5__7_), .CO(
        u5_mult_79_CARRYB_6__6_), .S(u5_mult_79_SUMB_6__6_) );
  FA_X1 u5_mult_79_S2_6_5 ( .A(u5_mult_79_ab_6__5_), .B(
        u5_mult_79_CARRYB_5__5_), .CI(u5_mult_79_SUMB_5__6_), .CO(
        u5_mult_79_CARRYB_6__5_), .S(u5_mult_79_SUMB_6__5_) );
  FA_X1 u5_mult_79_S2_6_4 ( .A(u5_mult_79_ab_6__4_), .B(
        u5_mult_79_CARRYB_5__4_), .CI(u5_mult_79_SUMB_5__5_), .CO(
        u5_mult_79_CARRYB_6__4_), .S(u5_mult_79_SUMB_6__4_) );
  FA_X1 u5_mult_79_S2_6_3 ( .A(u5_mult_79_ab_6__3_), .B(
        u5_mult_79_CARRYB_5__3_), .CI(u5_mult_79_SUMB_5__4_), .CO(
        u5_mult_79_CARRYB_6__3_), .S(u5_mult_79_SUMB_6__3_) );
  FA_X1 u5_mult_79_S2_6_2 ( .A(u5_mult_79_ab_6__2_), .B(
        u5_mult_79_CARRYB_5__2_), .CI(u5_mult_79_SUMB_5__3_), .CO(
        u5_mult_79_CARRYB_6__2_), .S(u5_mult_79_SUMB_6__2_) );
  FA_X1 u5_mult_79_S2_6_1 ( .A(u5_mult_79_ab_6__1_), .B(
        u5_mult_79_CARRYB_5__1_), .CI(u5_mult_79_SUMB_5__2_), .CO(
        u5_mult_79_CARRYB_6__1_), .S(u5_mult_79_SUMB_6__1_) );
  FA_X1 u5_mult_79_S1_6_0 ( .A(u5_mult_79_ab_6__0_), .B(
        u5_mult_79_CARRYB_5__0_), .CI(u5_mult_79_SUMB_5__1_), .CO(
        u5_mult_79_CARRYB_6__0_), .S(u5_N6) );
  FA_X1 u5_mult_79_S3_7_22 ( .A(u5_mult_79_ab_7__22_), .B(
        u5_mult_79_CARRYB_6__22_), .CI(u5_mult_79_ab_6__23_), .CO(
        u5_mult_79_CARRYB_7__22_), .S(u5_mult_79_SUMB_7__22_) );
  FA_X1 u5_mult_79_S2_7_21 ( .A(u5_mult_79_ab_7__21_), .B(
        u5_mult_79_CARRYB_6__21_), .CI(u5_mult_79_SUMB_6__22_), .CO(
        u5_mult_79_CARRYB_7__21_), .S(u5_mult_79_SUMB_7__21_) );
  FA_X1 u5_mult_79_S2_7_20 ( .A(u5_mult_79_ab_7__20_), .B(
        u5_mult_79_CARRYB_6__20_), .CI(u5_mult_79_SUMB_6__21_), .CO(
        u5_mult_79_CARRYB_7__20_), .S(u5_mult_79_SUMB_7__20_) );
  FA_X1 u5_mult_79_S2_7_19 ( .A(u5_mult_79_ab_7__19_), .B(
        u5_mult_79_CARRYB_6__19_), .CI(u5_mult_79_SUMB_6__20_), .CO(
        u5_mult_79_CARRYB_7__19_), .S(u5_mult_79_SUMB_7__19_) );
  FA_X1 u5_mult_79_S2_7_18 ( .A(u5_mult_79_ab_7__18_), .B(
        u5_mult_79_CARRYB_6__18_), .CI(u5_mult_79_SUMB_6__19_), .CO(
        u5_mult_79_CARRYB_7__18_), .S(u5_mult_79_SUMB_7__18_) );
  FA_X1 u5_mult_79_S2_7_17 ( .A(u5_mult_79_ab_7__17_), .B(
        u5_mult_79_CARRYB_6__17_), .CI(u5_mult_79_SUMB_6__18_), .CO(
        u5_mult_79_CARRYB_7__17_), .S(u5_mult_79_SUMB_7__17_) );
  FA_X1 u5_mult_79_S2_7_16 ( .A(u5_mult_79_ab_7__16_), .B(
        u5_mult_79_CARRYB_6__16_), .CI(u5_mult_79_SUMB_6__17_), .CO(
        u5_mult_79_CARRYB_7__16_), .S(u5_mult_79_SUMB_7__16_) );
  FA_X1 u5_mult_79_S2_7_15 ( .A(u5_mult_79_ab_7__15_), .B(
        u5_mult_79_CARRYB_6__15_), .CI(u5_mult_79_SUMB_6__16_), .CO(
        u5_mult_79_CARRYB_7__15_), .S(u5_mult_79_SUMB_7__15_) );
  FA_X1 u5_mult_79_S2_7_14 ( .A(u5_mult_79_ab_7__14_), .B(
        u5_mult_79_CARRYB_6__14_), .CI(u5_mult_79_SUMB_6__15_), .CO(
        u5_mult_79_CARRYB_7__14_), .S(u5_mult_79_SUMB_7__14_) );
  FA_X1 u5_mult_79_S2_7_13 ( .A(u5_mult_79_ab_7__13_), .B(
        u5_mult_79_CARRYB_6__13_), .CI(u5_mult_79_SUMB_6__14_), .CO(
        u5_mult_79_CARRYB_7__13_), .S(u5_mult_79_SUMB_7__13_) );
  FA_X1 u5_mult_79_S2_7_12 ( .A(u5_mult_79_ab_7__12_), .B(
        u5_mult_79_CARRYB_6__12_), .CI(u5_mult_79_SUMB_6__13_), .CO(
        u5_mult_79_CARRYB_7__12_), .S(u5_mult_79_SUMB_7__12_) );
  FA_X1 u5_mult_79_S2_7_11 ( .A(u5_mult_79_ab_7__11_), .B(
        u5_mult_79_CARRYB_6__11_), .CI(u5_mult_79_SUMB_6__12_), .CO(
        u5_mult_79_CARRYB_7__11_), .S(u5_mult_79_SUMB_7__11_) );
  FA_X1 u5_mult_79_S2_7_10 ( .A(u5_mult_79_ab_7__10_), .B(
        u5_mult_79_CARRYB_6__10_), .CI(u5_mult_79_SUMB_6__11_), .CO(
        u5_mult_79_CARRYB_7__10_), .S(u5_mult_79_SUMB_7__10_) );
  FA_X1 u5_mult_79_S2_7_9 ( .A(u5_mult_79_ab_7__9_), .B(
        u5_mult_79_CARRYB_6__9_), .CI(u5_mult_79_SUMB_6__10_), .CO(
        u5_mult_79_CARRYB_7__9_), .S(u5_mult_79_SUMB_7__9_) );
  FA_X1 u5_mult_79_S2_7_8 ( .A(u5_mult_79_ab_7__8_), .B(
        u5_mult_79_CARRYB_6__8_), .CI(u5_mult_79_SUMB_6__9_), .CO(
        u5_mult_79_CARRYB_7__8_), .S(u5_mult_79_SUMB_7__8_) );
  FA_X1 u5_mult_79_S2_7_7 ( .A(u5_mult_79_ab_7__7_), .B(
        u5_mult_79_CARRYB_6__7_), .CI(u5_mult_79_SUMB_6__8_), .CO(
        u5_mult_79_CARRYB_7__7_), .S(u5_mult_79_SUMB_7__7_) );
  FA_X1 u5_mult_79_S2_7_6 ( .A(u5_mult_79_ab_7__6_), .B(
        u5_mult_79_CARRYB_6__6_), .CI(u5_mult_79_SUMB_6__7_), .CO(
        u5_mult_79_CARRYB_7__6_), .S(u5_mult_79_SUMB_7__6_) );
  FA_X1 u5_mult_79_S2_7_5 ( .A(u5_mult_79_ab_7__5_), .B(
        u5_mult_79_CARRYB_6__5_), .CI(u5_mult_79_SUMB_6__6_), .CO(
        u5_mult_79_CARRYB_7__5_), .S(u5_mult_79_SUMB_7__5_) );
  FA_X1 u5_mult_79_S2_7_4 ( .A(u5_mult_79_ab_7__4_), .B(
        u5_mult_79_CARRYB_6__4_), .CI(u5_mult_79_SUMB_6__5_), .CO(
        u5_mult_79_CARRYB_7__4_), .S(u5_mult_79_SUMB_7__4_) );
  FA_X1 u5_mult_79_S2_7_3 ( .A(u5_mult_79_ab_7__3_), .B(
        u5_mult_79_CARRYB_6__3_), .CI(u5_mult_79_SUMB_6__4_), .CO(
        u5_mult_79_CARRYB_7__3_), .S(u5_mult_79_SUMB_7__3_) );
  FA_X1 u5_mult_79_S2_7_2 ( .A(u5_mult_79_ab_7__2_), .B(
        u5_mult_79_CARRYB_6__2_), .CI(u5_mult_79_SUMB_6__3_), .CO(
        u5_mult_79_CARRYB_7__2_), .S(u5_mult_79_SUMB_7__2_) );
  FA_X1 u5_mult_79_S2_7_1 ( .A(u5_mult_79_ab_7__1_), .B(
        u5_mult_79_CARRYB_6__1_), .CI(u5_mult_79_SUMB_6__2_), .CO(
        u5_mult_79_CARRYB_7__1_), .S(u5_mult_79_SUMB_7__1_) );
  FA_X1 u5_mult_79_S1_7_0 ( .A(u5_mult_79_ab_7__0_), .B(
        u5_mult_79_CARRYB_6__0_), .CI(u5_mult_79_SUMB_6__1_), .CO(
        u5_mult_79_CARRYB_7__0_), .S(u5_N7) );
  FA_X1 u5_mult_79_S3_8_22 ( .A(u5_mult_79_ab_8__22_), .B(
        u5_mult_79_CARRYB_7__22_), .CI(u5_mult_79_ab_7__23_), .CO(
        u5_mult_79_CARRYB_8__22_), .S(u5_mult_79_SUMB_8__22_) );
  FA_X1 u5_mult_79_S2_8_21 ( .A(u5_mult_79_ab_8__21_), .B(
        u5_mult_79_CARRYB_7__21_), .CI(u5_mult_79_SUMB_7__22_), .CO(
        u5_mult_79_CARRYB_8__21_), .S(u5_mult_79_SUMB_8__21_) );
  FA_X1 u5_mult_79_S2_8_20 ( .A(u5_mult_79_ab_8__20_), .B(
        u5_mult_79_CARRYB_7__20_), .CI(u5_mult_79_SUMB_7__21_), .CO(
        u5_mult_79_CARRYB_8__20_), .S(u5_mult_79_SUMB_8__20_) );
  FA_X1 u5_mult_79_S2_8_19 ( .A(u5_mult_79_ab_8__19_), .B(
        u5_mult_79_CARRYB_7__19_), .CI(u5_mult_79_SUMB_7__20_), .CO(
        u5_mult_79_CARRYB_8__19_), .S(u5_mult_79_SUMB_8__19_) );
  FA_X1 u5_mult_79_S2_8_18 ( .A(u5_mult_79_ab_8__18_), .B(
        u5_mult_79_CARRYB_7__18_), .CI(u5_mult_79_SUMB_7__19_), .CO(
        u5_mult_79_CARRYB_8__18_), .S(u5_mult_79_SUMB_8__18_) );
  FA_X1 u5_mult_79_S2_8_17 ( .A(u5_mult_79_ab_8__17_), .B(
        u5_mult_79_CARRYB_7__17_), .CI(u5_mult_79_SUMB_7__18_), .CO(
        u5_mult_79_CARRYB_8__17_), .S(u5_mult_79_SUMB_8__17_) );
  FA_X1 u5_mult_79_S2_8_16 ( .A(u5_mult_79_ab_8__16_), .B(
        u5_mult_79_CARRYB_7__16_), .CI(u5_mult_79_SUMB_7__17_), .CO(
        u5_mult_79_CARRYB_8__16_), .S(u5_mult_79_SUMB_8__16_) );
  FA_X1 u5_mult_79_S2_8_15 ( .A(u5_mult_79_ab_8__15_), .B(
        u5_mult_79_CARRYB_7__15_), .CI(u5_mult_79_SUMB_7__16_), .CO(
        u5_mult_79_CARRYB_8__15_), .S(u5_mult_79_SUMB_8__15_) );
  FA_X1 u5_mult_79_S2_8_14 ( .A(u5_mult_79_ab_8__14_), .B(
        u5_mult_79_CARRYB_7__14_), .CI(u5_mult_79_SUMB_7__15_), .CO(
        u5_mult_79_CARRYB_8__14_), .S(u5_mult_79_SUMB_8__14_) );
  FA_X1 u5_mult_79_S2_8_13 ( .A(u5_mult_79_ab_8__13_), .B(
        u5_mult_79_CARRYB_7__13_), .CI(u5_mult_79_SUMB_7__14_), .CO(
        u5_mult_79_CARRYB_8__13_), .S(u5_mult_79_SUMB_8__13_) );
  FA_X1 u5_mult_79_S2_8_12 ( .A(u5_mult_79_ab_8__12_), .B(
        u5_mult_79_CARRYB_7__12_), .CI(u5_mult_79_SUMB_7__13_), .CO(
        u5_mult_79_CARRYB_8__12_), .S(u5_mult_79_SUMB_8__12_) );
  FA_X1 u5_mult_79_S2_8_11 ( .A(u5_mult_79_ab_8__11_), .B(
        u5_mult_79_CARRYB_7__11_), .CI(u5_mult_79_SUMB_7__12_), .CO(
        u5_mult_79_CARRYB_8__11_), .S(u5_mult_79_SUMB_8__11_) );
  FA_X1 u5_mult_79_S2_8_10 ( .A(u5_mult_79_ab_8__10_), .B(
        u5_mult_79_CARRYB_7__10_), .CI(u5_mult_79_SUMB_7__11_), .CO(
        u5_mult_79_CARRYB_8__10_), .S(u5_mult_79_SUMB_8__10_) );
  FA_X1 u5_mult_79_S2_8_9 ( .A(u5_mult_79_ab_8__9_), .B(
        u5_mult_79_CARRYB_7__9_), .CI(u5_mult_79_SUMB_7__10_), .CO(
        u5_mult_79_CARRYB_8__9_), .S(u5_mult_79_SUMB_8__9_) );
  FA_X1 u5_mult_79_S2_8_8 ( .A(u5_mult_79_ab_8__8_), .B(
        u5_mult_79_CARRYB_7__8_), .CI(u5_mult_79_SUMB_7__9_), .CO(
        u5_mult_79_CARRYB_8__8_), .S(u5_mult_79_SUMB_8__8_) );
  FA_X1 u5_mult_79_S2_8_7 ( .A(u5_mult_79_ab_8__7_), .B(
        u5_mult_79_CARRYB_7__7_), .CI(u5_mult_79_SUMB_7__8_), .CO(
        u5_mult_79_CARRYB_8__7_), .S(u5_mult_79_SUMB_8__7_) );
  FA_X1 u5_mult_79_S2_8_6 ( .A(u5_mult_79_ab_8__6_), .B(
        u5_mult_79_CARRYB_7__6_), .CI(u5_mult_79_SUMB_7__7_), .CO(
        u5_mult_79_CARRYB_8__6_), .S(u5_mult_79_SUMB_8__6_) );
  FA_X1 u5_mult_79_S2_8_5 ( .A(u5_mult_79_ab_8__5_), .B(
        u5_mult_79_CARRYB_7__5_), .CI(u5_mult_79_SUMB_7__6_), .CO(
        u5_mult_79_CARRYB_8__5_), .S(u5_mult_79_SUMB_8__5_) );
  FA_X1 u5_mult_79_S2_8_4 ( .A(u5_mult_79_ab_8__4_), .B(
        u5_mult_79_CARRYB_7__4_), .CI(u5_mult_79_SUMB_7__5_), .CO(
        u5_mult_79_CARRYB_8__4_), .S(u5_mult_79_SUMB_8__4_) );
  FA_X1 u5_mult_79_S2_8_3 ( .A(u5_mult_79_ab_8__3_), .B(
        u5_mult_79_CARRYB_7__3_), .CI(u5_mult_79_SUMB_7__4_), .CO(
        u5_mult_79_CARRYB_8__3_), .S(u5_mult_79_SUMB_8__3_) );
  FA_X1 u5_mult_79_S2_8_2 ( .A(u5_mult_79_ab_8__2_), .B(
        u5_mult_79_CARRYB_7__2_), .CI(u5_mult_79_SUMB_7__3_), .CO(
        u5_mult_79_CARRYB_8__2_), .S(u5_mult_79_SUMB_8__2_) );
  FA_X1 u5_mult_79_S2_8_1 ( .A(u5_mult_79_ab_8__1_), .B(
        u5_mult_79_CARRYB_7__1_), .CI(u5_mult_79_SUMB_7__2_), .CO(
        u5_mult_79_CARRYB_8__1_), .S(u5_mult_79_SUMB_8__1_) );
  FA_X1 u5_mult_79_S1_8_0 ( .A(u5_mult_79_ab_8__0_), .B(
        u5_mult_79_CARRYB_7__0_), .CI(u5_mult_79_SUMB_7__1_), .CO(
        u5_mult_79_CARRYB_8__0_), .S(u5_N8) );
  FA_X1 u5_mult_79_S3_9_22 ( .A(u5_mult_79_ab_9__22_), .B(
        u5_mult_79_CARRYB_8__22_), .CI(u5_mult_79_ab_8__23_), .CO(
        u5_mult_79_CARRYB_9__22_), .S(u5_mult_79_SUMB_9__22_) );
  FA_X1 u5_mult_79_S2_9_21 ( .A(u5_mult_79_ab_9__21_), .B(
        u5_mult_79_CARRYB_8__21_), .CI(u5_mult_79_SUMB_8__22_), .CO(
        u5_mult_79_CARRYB_9__21_), .S(u5_mult_79_SUMB_9__21_) );
  FA_X1 u5_mult_79_S2_9_20 ( .A(u5_mult_79_ab_9__20_), .B(
        u5_mult_79_CARRYB_8__20_), .CI(u5_mult_79_SUMB_8__21_), .CO(
        u5_mult_79_CARRYB_9__20_), .S(u5_mult_79_SUMB_9__20_) );
  FA_X1 u5_mult_79_S2_9_19 ( .A(u5_mult_79_ab_9__19_), .B(
        u5_mult_79_CARRYB_8__19_), .CI(u5_mult_79_SUMB_8__20_), .CO(
        u5_mult_79_CARRYB_9__19_), .S(u5_mult_79_SUMB_9__19_) );
  FA_X1 u5_mult_79_S2_9_18 ( .A(u5_mult_79_ab_9__18_), .B(
        u5_mult_79_CARRYB_8__18_), .CI(u5_mult_79_SUMB_8__19_), .CO(
        u5_mult_79_CARRYB_9__18_), .S(u5_mult_79_SUMB_9__18_) );
  FA_X1 u5_mult_79_S2_9_17 ( .A(u5_mult_79_ab_9__17_), .B(
        u5_mult_79_CARRYB_8__17_), .CI(u5_mult_79_SUMB_8__18_), .CO(
        u5_mult_79_CARRYB_9__17_), .S(u5_mult_79_SUMB_9__17_) );
  FA_X1 u5_mult_79_S2_9_16 ( .A(u5_mult_79_ab_9__16_), .B(
        u5_mult_79_CARRYB_8__16_), .CI(u5_mult_79_SUMB_8__17_), .CO(
        u5_mult_79_CARRYB_9__16_), .S(u5_mult_79_SUMB_9__16_) );
  FA_X1 u5_mult_79_S2_9_15 ( .A(u5_mult_79_ab_9__15_), .B(
        u5_mult_79_CARRYB_8__15_), .CI(u5_mult_79_SUMB_8__16_), .CO(
        u5_mult_79_CARRYB_9__15_), .S(u5_mult_79_SUMB_9__15_) );
  FA_X1 u5_mult_79_S2_9_14 ( .A(u5_mult_79_ab_9__14_), .B(
        u5_mult_79_CARRYB_8__14_), .CI(u5_mult_79_SUMB_8__15_), .CO(
        u5_mult_79_CARRYB_9__14_), .S(u5_mult_79_SUMB_9__14_) );
  FA_X1 u5_mult_79_S2_9_13 ( .A(u5_mult_79_ab_9__13_), .B(
        u5_mult_79_CARRYB_8__13_), .CI(u5_mult_79_SUMB_8__14_), .CO(
        u5_mult_79_CARRYB_9__13_), .S(u5_mult_79_SUMB_9__13_) );
  FA_X1 u5_mult_79_S2_9_12 ( .A(u5_mult_79_ab_9__12_), .B(
        u5_mult_79_CARRYB_8__12_), .CI(u5_mult_79_SUMB_8__13_), .CO(
        u5_mult_79_CARRYB_9__12_), .S(u5_mult_79_SUMB_9__12_) );
  FA_X1 u5_mult_79_S2_9_11 ( .A(u5_mult_79_ab_9__11_), .B(
        u5_mult_79_CARRYB_8__11_), .CI(u5_mult_79_SUMB_8__12_), .CO(
        u5_mult_79_CARRYB_9__11_), .S(u5_mult_79_SUMB_9__11_) );
  FA_X1 u5_mult_79_S2_9_10 ( .A(u5_mult_79_ab_9__10_), .B(
        u5_mult_79_CARRYB_8__10_), .CI(u5_mult_79_SUMB_8__11_), .CO(
        u5_mult_79_CARRYB_9__10_), .S(u5_mult_79_SUMB_9__10_) );
  FA_X1 u5_mult_79_S2_9_9 ( .A(u5_mult_79_ab_9__9_), .B(
        u5_mult_79_CARRYB_8__9_), .CI(u5_mult_79_SUMB_8__10_), .CO(
        u5_mult_79_CARRYB_9__9_), .S(u5_mult_79_SUMB_9__9_) );
  FA_X1 u5_mult_79_S2_9_8 ( .A(u5_mult_79_ab_9__8_), .B(
        u5_mult_79_CARRYB_8__8_), .CI(u5_mult_79_SUMB_8__9_), .CO(
        u5_mult_79_CARRYB_9__8_), .S(u5_mult_79_SUMB_9__8_) );
  FA_X1 u5_mult_79_S2_9_7 ( .A(u5_mult_79_ab_9__7_), .B(
        u5_mult_79_CARRYB_8__7_), .CI(u5_mult_79_SUMB_8__8_), .CO(
        u5_mult_79_CARRYB_9__7_), .S(u5_mult_79_SUMB_9__7_) );
  FA_X1 u5_mult_79_S2_9_6 ( .A(u5_mult_79_ab_9__6_), .B(
        u5_mult_79_CARRYB_8__6_), .CI(u5_mult_79_SUMB_8__7_), .CO(
        u5_mult_79_CARRYB_9__6_), .S(u5_mult_79_SUMB_9__6_) );
  FA_X1 u5_mult_79_S2_9_5 ( .A(u5_mult_79_ab_9__5_), .B(
        u5_mult_79_CARRYB_8__5_), .CI(u5_mult_79_SUMB_8__6_), .CO(
        u5_mult_79_CARRYB_9__5_), .S(u5_mult_79_SUMB_9__5_) );
  FA_X1 u5_mult_79_S2_9_4 ( .A(u5_mult_79_ab_9__4_), .B(
        u5_mult_79_CARRYB_8__4_), .CI(u5_mult_79_SUMB_8__5_), .CO(
        u5_mult_79_CARRYB_9__4_), .S(u5_mult_79_SUMB_9__4_) );
  FA_X1 u5_mult_79_S2_9_3 ( .A(u5_mult_79_ab_9__3_), .B(
        u5_mult_79_CARRYB_8__3_), .CI(u5_mult_79_SUMB_8__4_), .CO(
        u5_mult_79_CARRYB_9__3_), .S(u5_mult_79_SUMB_9__3_) );
  FA_X1 u5_mult_79_S2_9_2 ( .A(u5_mult_79_ab_9__2_), .B(
        u5_mult_79_CARRYB_8__2_), .CI(u5_mult_79_SUMB_8__3_), .CO(
        u5_mult_79_CARRYB_9__2_), .S(u5_mult_79_SUMB_9__2_) );
  FA_X1 u5_mult_79_S2_9_1 ( .A(u5_mult_79_ab_9__1_), .B(
        u5_mult_79_CARRYB_8__1_), .CI(u5_mult_79_SUMB_8__2_), .CO(
        u5_mult_79_CARRYB_9__1_), .S(u5_mult_79_SUMB_9__1_) );
  FA_X1 u5_mult_79_S1_9_0 ( .A(u5_mult_79_ab_9__0_), .B(
        u5_mult_79_CARRYB_8__0_), .CI(u5_mult_79_SUMB_8__1_), .CO(
        u5_mult_79_CARRYB_9__0_), .S(u5_N9) );
  FA_X1 u5_mult_79_S3_10_22 ( .A(u5_mult_79_ab_10__22_), .B(
        u5_mult_79_CARRYB_9__22_), .CI(u5_mult_79_ab_9__23_), .CO(
        u5_mult_79_CARRYB_10__22_), .S(u5_mult_79_SUMB_10__22_) );
  FA_X1 u5_mult_79_S2_10_21 ( .A(u5_mult_79_ab_10__21_), .B(
        u5_mult_79_CARRYB_9__21_), .CI(u5_mult_79_SUMB_9__22_), .CO(
        u5_mult_79_CARRYB_10__21_), .S(u5_mult_79_SUMB_10__21_) );
  FA_X1 u5_mult_79_S2_10_20 ( .A(u5_mult_79_ab_10__20_), .B(
        u5_mult_79_CARRYB_9__20_), .CI(u5_mult_79_SUMB_9__21_), .CO(
        u5_mult_79_CARRYB_10__20_), .S(u5_mult_79_SUMB_10__20_) );
  FA_X1 u5_mult_79_S2_10_19 ( .A(u5_mult_79_ab_10__19_), .B(
        u5_mult_79_CARRYB_9__19_), .CI(u5_mult_79_SUMB_9__20_), .CO(
        u5_mult_79_CARRYB_10__19_), .S(u5_mult_79_SUMB_10__19_) );
  FA_X1 u5_mult_79_S2_10_18 ( .A(u5_mult_79_ab_10__18_), .B(
        u5_mult_79_CARRYB_9__18_), .CI(u5_mult_79_SUMB_9__19_), .CO(
        u5_mult_79_CARRYB_10__18_), .S(u5_mult_79_SUMB_10__18_) );
  FA_X1 u5_mult_79_S2_10_17 ( .A(u5_mult_79_ab_10__17_), .B(
        u5_mult_79_CARRYB_9__17_), .CI(u5_mult_79_SUMB_9__18_), .CO(
        u5_mult_79_CARRYB_10__17_), .S(u5_mult_79_SUMB_10__17_) );
  FA_X1 u5_mult_79_S2_10_16 ( .A(u5_mult_79_ab_10__16_), .B(
        u5_mult_79_CARRYB_9__16_), .CI(u5_mult_79_SUMB_9__17_), .CO(
        u5_mult_79_CARRYB_10__16_), .S(u5_mult_79_SUMB_10__16_) );
  FA_X1 u5_mult_79_S2_10_15 ( .A(u5_mult_79_ab_10__15_), .B(
        u5_mult_79_CARRYB_9__15_), .CI(u5_mult_79_SUMB_9__16_), .CO(
        u5_mult_79_CARRYB_10__15_), .S(u5_mult_79_SUMB_10__15_) );
  FA_X1 u5_mult_79_S2_10_14 ( .A(u5_mult_79_ab_10__14_), .B(
        u5_mult_79_CARRYB_9__14_), .CI(u5_mult_79_SUMB_9__15_), .CO(
        u5_mult_79_CARRYB_10__14_), .S(u5_mult_79_SUMB_10__14_) );
  FA_X1 u5_mult_79_S2_10_13 ( .A(u5_mult_79_ab_10__13_), .B(
        u5_mult_79_CARRYB_9__13_), .CI(u5_mult_79_SUMB_9__14_), .CO(
        u5_mult_79_CARRYB_10__13_), .S(u5_mult_79_SUMB_10__13_) );
  FA_X1 u5_mult_79_S2_10_12 ( .A(u5_mult_79_ab_10__12_), .B(
        u5_mult_79_CARRYB_9__12_), .CI(u5_mult_79_SUMB_9__13_), .CO(
        u5_mult_79_CARRYB_10__12_), .S(u5_mult_79_SUMB_10__12_) );
  FA_X1 u5_mult_79_S2_10_11 ( .A(u5_mult_79_ab_10__11_), .B(
        u5_mult_79_CARRYB_9__11_), .CI(u5_mult_79_SUMB_9__12_), .CO(
        u5_mult_79_CARRYB_10__11_), .S(u5_mult_79_SUMB_10__11_) );
  FA_X1 u5_mult_79_S2_10_10 ( .A(u5_mult_79_ab_10__10_), .B(
        u5_mult_79_CARRYB_9__10_), .CI(u5_mult_79_SUMB_9__11_), .CO(
        u5_mult_79_CARRYB_10__10_), .S(u5_mult_79_SUMB_10__10_) );
  FA_X1 u5_mult_79_S2_10_9 ( .A(u5_mult_79_ab_10__9_), .B(
        u5_mult_79_CARRYB_9__9_), .CI(u5_mult_79_SUMB_9__10_), .CO(
        u5_mult_79_CARRYB_10__9_), .S(u5_mult_79_SUMB_10__9_) );
  FA_X1 u5_mult_79_S2_10_8 ( .A(u5_mult_79_ab_10__8_), .B(
        u5_mult_79_CARRYB_9__8_), .CI(u5_mult_79_SUMB_9__9_), .CO(
        u5_mult_79_CARRYB_10__8_), .S(u5_mult_79_SUMB_10__8_) );
  FA_X1 u5_mult_79_S2_10_7 ( .A(u5_mult_79_ab_10__7_), .B(
        u5_mult_79_CARRYB_9__7_), .CI(u5_mult_79_SUMB_9__8_), .CO(
        u5_mult_79_CARRYB_10__7_), .S(u5_mult_79_SUMB_10__7_) );
  FA_X1 u5_mult_79_S2_10_6 ( .A(u5_mult_79_ab_10__6_), .B(
        u5_mult_79_CARRYB_9__6_), .CI(u5_mult_79_SUMB_9__7_), .CO(
        u5_mult_79_CARRYB_10__6_), .S(u5_mult_79_SUMB_10__6_) );
  FA_X1 u5_mult_79_S2_10_5 ( .A(u5_mult_79_ab_10__5_), .B(
        u5_mult_79_CARRYB_9__5_), .CI(u5_mult_79_SUMB_9__6_), .CO(
        u5_mult_79_CARRYB_10__5_), .S(u5_mult_79_SUMB_10__5_) );
  FA_X1 u5_mult_79_S2_10_4 ( .A(u5_mult_79_ab_10__4_), .B(
        u5_mult_79_CARRYB_9__4_), .CI(u5_mult_79_SUMB_9__5_), .CO(
        u5_mult_79_CARRYB_10__4_), .S(u5_mult_79_SUMB_10__4_) );
  FA_X1 u5_mult_79_S2_10_3 ( .A(u5_mult_79_ab_10__3_), .B(
        u5_mult_79_CARRYB_9__3_), .CI(u5_mult_79_SUMB_9__4_), .CO(
        u5_mult_79_CARRYB_10__3_), .S(u5_mult_79_SUMB_10__3_) );
  FA_X1 u5_mult_79_S2_10_2 ( .A(u5_mult_79_ab_10__2_), .B(
        u5_mult_79_CARRYB_9__2_), .CI(u5_mult_79_SUMB_9__3_), .CO(
        u5_mult_79_CARRYB_10__2_), .S(u5_mult_79_SUMB_10__2_) );
  FA_X1 u5_mult_79_S2_10_1 ( .A(u5_mult_79_ab_10__1_), .B(
        u5_mult_79_CARRYB_9__1_), .CI(u5_mult_79_SUMB_9__2_), .CO(
        u5_mult_79_CARRYB_10__1_), .S(u5_mult_79_SUMB_10__1_) );
  FA_X1 u5_mult_79_S1_10_0 ( .A(u5_mult_79_ab_10__0_), .B(
        u5_mult_79_CARRYB_9__0_), .CI(u5_mult_79_SUMB_9__1_), .CO(
        u5_mult_79_CARRYB_10__0_), .S(u5_N10) );
  FA_X1 u5_mult_79_S3_11_22 ( .A(u5_mult_79_ab_11__22_), .B(
        u5_mult_79_CARRYB_10__22_), .CI(u5_mult_79_ab_10__23_), .CO(
        u5_mult_79_CARRYB_11__22_), .S(u5_mult_79_SUMB_11__22_) );
  FA_X1 u5_mult_79_S2_11_21 ( .A(u5_mult_79_ab_11__21_), .B(
        u5_mult_79_CARRYB_10__21_), .CI(u5_mult_79_SUMB_10__22_), .CO(
        u5_mult_79_CARRYB_11__21_), .S(u5_mult_79_SUMB_11__21_) );
  FA_X1 u5_mult_79_S2_11_20 ( .A(u5_mult_79_ab_11__20_), .B(
        u5_mult_79_CARRYB_10__20_), .CI(u5_mult_79_SUMB_10__21_), .CO(
        u5_mult_79_CARRYB_11__20_), .S(u5_mult_79_SUMB_11__20_) );
  FA_X1 u5_mult_79_S2_11_19 ( .A(u5_mult_79_ab_11__19_), .B(
        u5_mult_79_CARRYB_10__19_), .CI(u5_mult_79_SUMB_10__20_), .CO(
        u5_mult_79_CARRYB_11__19_), .S(u5_mult_79_SUMB_11__19_) );
  FA_X1 u5_mult_79_S2_11_18 ( .A(u5_mult_79_ab_11__18_), .B(
        u5_mult_79_CARRYB_10__18_), .CI(u5_mult_79_SUMB_10__19_), .CO(
        u5_mult_79_CARRYB_11__18_), .S(u5_mult_79_SUMB_11__18_) );
  FA_X1 u5_mult_79_S2_11_17 ( .A(u5_mult_79_ab_11__17_), .B(
        u5_mult_79_CARRYB_10__17_), .CI(u5_mult_79_SUMB_10__18_), .CO(
        u5_mult_79_CARRYB_11__17_), .S(u5_mult_79_SUMB_11__17_) );
  FA_X1 u5_mult_79_S2_11_16 ( .A(u5_mult_79_ab_11__16_), .B(
        u5_mult_79_CARRYB_10__16_), .CI(u5_mult_79_SUMB_10__17_), .CO(
        u5_mult_79_CARRYB_11__16_), .S(u5_mult_79_SUMB_11__16_) );
  FA_X1 u5_mult_79_S2_11_15 ( .A(u5_mult_79_ab_11__15_), .B(
        u5_mult_79_CARRYB_10__15_), .CI(u5_mult_79_SUMB_10__16_), .CO(
        u5_mult_79_CARRYB_11__15_), .S(u5_mult_79_SUMB_11__15_) );
  FA_X1 u5_mult_79_S2_11_14 ( .A(u5_mult_79_ab_11__14_), .B(
        u5_mult_79_CARRYB_10__14_), .CI(u5_mult_79_SUMB_10__15_), .CO(
        u5_mult_79_CARRYB_11__14_), .S(u5_mult_79_SUMB_11__14_) );
  FA_X1 u5_mult_79_S2_11_13 ( .A(u5_mult_79_ab_11__13_), .B(
        u5_mult_79_CARRYB_10__13_), .CI(u5_mult_79_SUMB_10__14_), .CO(
        u5_mult_79_CARRYB_11__13_), .S(u5_mult_79_SUMB_11__13_) );
  FA_X1 u5_mult_79_S2_11_12 ( .A(u5_mult_79_ab_11__12_), .B(
        u5_mult_79_CARRYB_10__12_), .CI(u5_mult_79_SUMB_10__13_), .CO(
        u5_mult_79_CARRYB_11__12_), .S(u5_mult_79_SUMB_11__12_) );
  FA_X1 u5_mult_79_S2_11_11 ( .A(u5_mult_79_ab_11__11_), .B(
        u5_mult_79_CARRYB_10__11_), .CI(u5_mult_79_SUMB_10__12_), .CO(
        u5_mult_79_CARRYB_11__11_), .S(u5_mult_79_SUMB_11__11_) );
  FA_X1 u5_mult_79_S2_11_10 ( .A(u5_mult_79_ab_11__10_), .B(
        u5_mult_79_CARRYB_10__10_), .CI(u5_mult_79_SUMB_10__11_), .CO(
        u5_mult_79_CARRYB_11__10_), .S(u5_mult_79_SUMB_11__10_) );
  FA_X1 u5_mult_79_S2_11_9 ( .A(u5_mult_79_ab_11__9_), .B(
        u5_mult_79_CARRYB_10__9_), .CI(u5_mult_79_SUMB_10__10_), .CO(
        u5_mult_79_CARRYB_11__9_), .S(u5_mult_79_SUMB_11__9_) );
  FA_X1 u5_mult_79_S2_11_8 ( .A(u5_mult_79_ab_11__8_), .B(
        u5_mult_79_CARRYB_10__8_), .CI(u5_mult_79_SUMB_10__9_), .CO(
        u5_mult_79_CARRYB_11__8_), .S(u5_mult_79_SUMB_11__8_) );
  FA_X1 u5_mult_79_S2_11_7 ( .A(u5_mult_79_ab_11__7_), .B(
        u5_mult_79_CARRYB_10__7_), .CI(u5_mult_79_SUMB_10__8_), .CO(
        u5_mult_79_CARRYB_11__7_), .S(u5_mult_79_SUMB_11__7_) );
  FA_X1 u5_mult_79_S2_11_6 ( .A(u5_mult_79_ab_11__6_), .B(
        u5_mult_79_CARRYB_10__6_), .CI(u5_mult_79_SUMB_10__7_), .CO(
        u5_mult_79_CARRYB_11__6_), .S(u5_mult_79_SUMB_11__6_) );
  FA_X1 u5_mult_79_S2_11_5 ( .A(u5_mult_79_ab_11__5_), .B(
        u5_mult_79_CARRYB_10__5_), .CI(u5_mult_79_SUMB_10__6_), .CO(
        u5_mult_79_CARRYB_11__5_), .S(u5_mult_79_SUMB_11__5_) );
  FA_X1 u5_mult_79_S2_11_4 ( .A(u5_mult_79_ab_11__4_), .B(
        u5_mult_79_CARRYB_10__4_), .CI(u5_mult_79_SUMB_10__5_), .CO(
        u5_mult_79_CARRYB_11__4_), .S(u5_mult_79_SUMB_11__4_) );
  FA_X1 u5_mult_79_S2_11_3 ( .A(u5_mult_79_ab_11__3_), .B(
        u5_mult_79_CARRYB_10__3_), .CI(u5_mult_79_SUMB_10__4_), .CO(
        u5_mult_79_CARRYB_11__3_), .S(u5_mult_79_SUMB_11__3_) );
  FA_X1 u5_mult_79_S2_11_2 ( .A(u5_mult_79_ab_11__2_), .B(
        u5_mult_79_CARRYB_10__2_), .CI(u5_mult_79_SUMB_10__3_), .CO(
        u5_mult_79_CARRYB_11__2_), .S(u5_mult_79_SUMB_11__2_) );
  FA_X1 u5_mult_79_S2_11_1 ( .A(u5_mult_79_ab_11__1_), .B(
        u5_mult_79_CARRYB_10__1_), .CI(u5_mult_79_SUMB_10__2_), .CO(
        u5_mult_79_CARRYB_11__1_), .S(u5_mult_79_SUMB_11__1_) );
  FA_X1 u5_mult_79_S1_11_0 ( .A(u5_mult_79_ab_11__0_), .B(
        u5_mult_79_CARRYB_10__0_), .CI(u5_mult_79_SUMB_10__1_), .CO(
        u5_mult_79_CARRYB_11__0_), .S(u5_N11) );
  FA_X1 u5_mult_79_S3_12_22 ( .A(u5_mult_79_ab_12__22_), .B(
        u5_mult_79_CARRYB_11__22_), .CI(u5_mult_79_ab_11__23_), .CO(
        u5_mult_79_CARRYB_12__22_), .S(u5_mult_79_SUMB_12__22_) );
  FA_X1 u5_mult_79_S2_12_21 ( .A(u5_mult_79_ab_12__21_), .B(
        u5_mult_79_CARRYB_11__21_), .CI(u5_mult_79_SUMB_11__22_), .CO(
        u5_mult_79_CARRYB_12__21_), .S(u5_mult_79_SUMB_12__21_) );
  FA_X1 u5_mult_79_S2_12_20 ( .A(u5_mult_79_ab_12__20_), .B(
        u5_mult_79_CARRYB_11__20_), .CI(u5_mult_79_SUMB_11__21_), .CO(
        u5_mult_79_CARRYB_12__20_), .S(u5_mult_79_SUMB_12__20_) );
  FA_X1 u5_mult_79_S2_12_19 ( .A(u5_mult_79_ab_12__19_), .B(
        u5_mult_79_CARRYB_11__19_), .CI(u5_mult_79_SUMB_11__20_), .CO(
        u5_mult_79_CARRYB_12__19_), .S(u5_mult_79_SUMB_12__19_) );
  FA_X1 u5_mult_79_S2_12_18 ( .A(u5_mult_79_ab_12__18_), .B(
        u5_mult_79_CARRYB_11__18_), .CI(u5_mult_79_SUMB_11__19_), .CO(
        u5_mult_79_CARRYB_12__18_), .S(u5_mult_79_SUMB_12__18_) );
  FA_X1 u5_mult_79_S2_12_17 ( .A(u5_mult_79_ab_12__17_), .B(
        u5_mult_79_CARRYB_11__17_), .CI(u5_mult_79_SUMB_11__18_), .CO(
        u5_mult_79_CARRYB_12__17_), .S(u5_mult_79_SUMB_12__17_) );
  FA_X1 u5_mult_79_S2_12_16 ( .A(u5_mult_79_ab_12__16_), .B(
        u5_mult_79_CARRYB_11__16_), .CI(u5_mult_79_SUMB_11__17_), .CO(
        u5_mult_79_CARRYB_12__16_), .S(u5_mult_79_SUMB_12__16_) );
  FA_X1 u5_mult_79_S2_12_15 ( .A(u5_mult_79_ab_12__15_), .B(
        u5_mult_79_CARRYB_11__15_), .CI(u5_mult_79_SUMB_11__16_), .CO(
        u5_mult_79_CARRYB_12__15_), .S(u5_mult_79_SUMB_12__15_) );
  FA_X1 u5_mult_79_S2_12_14 ( .A(u5_mult_79_ab_12__14_), .B(
        u5_mult_79_CARRYB_11__14_), .CI(u5_mult_79_SUMB_11__15_), .CO(
        u5_mult_79_CARRYB_12__14_), .S(u5_mult_79_SUMB_12__14_) );
  FA_X1 u5_mult_79_S2_12_13 ( .A(u5_mult_79_ab_12__13_), .B(
        u5_mult_79_CARRYB_11__13_), .CI(u5_mult_79_SUMB_11__14_), .CO(
        u5_mult_79_CARRYB_12__13_), .S(u5_mult_79_SUMB_12__13_) );
  FA_X1 u5_mult_79_S2_12_12 ( .A(u5_mult_79_ab_12__12_), .B(
        u5_mult_79_CARRYB_11__12_), .CI(u5_mult_79_SUMB_11__13_), .CO(
        u5_mult_79_CARRYB_12__12_), .S(u5_mult_79_SUMB_12__12_) );
  FA_X1 u5_mult_79_S2_12_11 ( .A(u5_mult_79_ab_12__11_), .B(
        u5_mult_79_CARRYB_11__11_), .CI(u5_mult_79_SUMB_11__12_), .CO(
        u5_mult_79_CARRYB_12__11_), .S(u5_mult_79_SUMB_12__11_) );
  FA_X1 u5_mult_79_S2_12_10 ( .A(u5_mult_79_ab_12__10_), .B(
        u5_mult_79_CARRYB_11__10_), .CI(u5_mult_79_SUMB_11__11_), .CO(
        u5_mult_79_CARRYB_12__10_), .S(u5_mult_79_SUMB_12__10_) );
  FA_X1 u5_mult_79_S2_12_9 ( .A(u5_mult_79_ab_12__9_), .B(
        u5_mult_79_CARRYB_11__9_), .CI(u5_mult_79_SUMB_11__10_), .CO(
        u5_mult_79_CARRYB_12__9_), .S(u5_mult_79_SUMB_12__9_) );
  FA_X1 u5_mult_79_S2_12_8 ( .A(u5_mult_79_ab_12__8_), .B(
        u5_mult_79_CARRYB_11__8_), .CI(u5_mult_79_SUMB_11__9_), .CO(
        u5_mult_79_CARRYB_12__8_), .S(u5_mult_79_SUMB_12__8_) );
  FA_X1 u5_mult_79_S2_12_7 ( .A(u5_mult_79_ab_12__7_), .B(
        u5_mult_79_CARRYB_11__7_), .CI(u5_mult_79_SUMB_11__8_), .CO(
        u5_mult_79_CARRYB_12__7_), .S(u5_mult_79_SUMB_12__7_) );
  FA_X1 u5_mult_79_S2_12_6 ( .A(u5_mult_79_ab_12__6_), .B(
        u5_mult_79_CARRYB_11__6_), .CI(u5_mult_79_SUMB_11__7_), .CO(
        u5_mult_79_CARRYB_12__6_), .S(u5_mult_79_SUMB_12__6_) );
  FA_X1 u5_mult_79_S2_12_5 ( .A(u5_mult_79_ab_12__5_), .B(
        u5_mult_79_CARRYB_11__5_), .CI(u5_mult_79_SUMB_11__6_), .CO(
        u5_mult_79_CARRYB_12__5_), .S(u5_mult_79_SUMB_12__5_) );
  FA_X1 u5_mult_79_S2_12_4 ( .A(u5_mult_79_ab_12__4_), .B(
        u5_mult_79_CARRYB_11__4_), .CI(u5_mult_79_SUMB_11__5_), .CO(
        u5_mult_79_CARRYB_12__4_), .S(u5_mult_79_SUMB_12__4_) );
  FA_X1 u5_mult_79_S2_12_3 ( .A(u5_mult_79_ab_12__3_), .B(
        u5_mult_79_CARRYB_11__3_), .CI(u5_mult_79_SUMB_11__4_), .CO(
        u5_mult_79_CARRYB_12__3_), .S(u5_mult_79_SUMB_12__3_) );
  FA_X1 u5_mult_79_S2_12_2 ( .A(u5_mult_79_ab_12__2_), .B(
        u5_mult_79_CARRYB_11__2_), .CI(u5_mult_79_SUMB_11__3_), .CO(
        u5_mult_79_CARRYB_12__2_), .S(u5_mult_79_SUMB_12__2_) );
  FA_X1 u5_mult_79_S2_12_1 ( .A(u5_mult_79_ab_12__1_), .B(
        u5_mult_79_CARRYB_11__1_), .CI(u5_mult_79_SUMB_11__2_), .CO(
        u5_mult_79_CARRYB_12__1_), .S(u5_mult_79_SUMB_12__1_) );
  FA_X1 u5_mult_79_S1_12_0 ( .A(u5_mult_79_ab_12__0_), .B(
        u5_mult_79_CARRYB_11__0_), .CI(u5_mult_79_SUMB_11__1_), .CO(
        u5_mult_79_CARRYB_12__0_), .S(u5_N12) );
  FA_X1 u5_mult_79_S3_13_22 ( .A(u5_mult_79_ab_13__22_), .B(
        u5_mult_79_CARRYB_12__22_), .CI(u5_mult_79_ab_12__23_), .CO(
        u5_mult_79_CARRYB_13__22_), .S(u5_mult_79_SUMB_13__22_) );
  FA_X1 u5_mult_79_S2_13_21 ( .A(u5_mult_79_ab_13__21_), .B(
        u5_mult_79_CARRYB_12__21_), .CI(u5_mult_79_SUMB_12__22_), .CO(
        u5_mult_79_CARRYB_13__21_), .S(u5_mult_79_SUMB_13__21_) );
  FA_X1 u5_mult_79_S2_13_20 ( .A(u5_mult_79_ab_13__20_), .B(
        u5_mult_79_CARRYB_12__20_), .CI(u5_mult_79_SUMB_12__21_), .CO(
        u5_mult_79_CARRYB_13__20_), .S(u5_mult_79_SUMB_13__20_) );
  FA_X1 u5_mult_79_S2_13_19 ( .A(u5_mult_79_ab_13__19_), .B(
        u5_mult_79_CARRYB_12__19_), .CI(u5_mult_79_SUMB_12__20_), .CO(
        u5_mult_79_CARRYB_13__19_), .S(u5_mult_79_SUMB_13__19_) );
  FA_X1 u5_mult_79_S2_13_18 ( .A(u5_mult_79_ab_13__18_), .B(
        u5_mult_79_CARRYB_12__18_), .CI(u5_mult_79_SUMB_12__19_), .CO(
        u5_mult_79_CARRYB_13__18_), .S(u5_mult_79_SUMB_13__18_) );
  FA_X1 u5_mult_79_S2_13_17 ( .A(u5_mult_79_ab_13__17_), .B(
        u5_mult_79_CARRYB_12__17_), .CI(u5_mult_79_SUMB_12__18_), .CO(
        u5_mult_79_CARRYB_13__17_), .S(u5_mult_79_SUMB_13__17_) );
  FA_X1 u5_mult_79_S2_13_16 ( .A(u5_mult_79_ab_13__16_), .B(
        u5_mult_79_CARRYB_12__16_), .CI(u5_mult_79_SUMB_12__17_), .CO(
        u5_mult_79_CARRYB_13__16_), .S(u5_mult_79_SUMB_13__16_) );
  FA_X1 u5_mult_79_S2_13_15 ( .A(u5_mult_79_ab_13__15_), .B(
        u5_mult_79_CARRYB_12__15_), .CI(u5_mult_79_SUMB_12__16_), .CO(
        u5_mult_79_CARRYB_13__15_), .S(u5_mult_79_SUMB_13__15_) );
  FA_X1 u5_mult_79_S2_13_14 ( .A(u5_mult_79_ab_13__14_), .B(
        u5_mult_79_CARRYB_12__14_), .CI(u5_mult_79_SUMB_12__15_), .CO(
        u5_mult_79_CARRYB_13__14_), .S(u5_mult_79_SUMB_13__14_) );
  FA_X1 u5_mult_79_S2_13_13 ( .A(u5_mult_79_ab_13__13_), .B(
        u5_mult_79_CARRYB_12__13_), .CI(u5_mult_79_SUMB_12__14_), .CO(
        u5_mult_79_CARRYB_13__13_), .S(u5_mult_79_SUMB_13__13_) );
  FA_X1 u5_mult_79_S2_13_12 ( .A(u5_mult_79_ab_13__12_), .B(
        u5_mult_79_CARRYB_12__12_), .CI(u5_mult_79_SUMB_12__13_), .CO(
        u5_mult_79_CARRYB_13__12_), .S(u5_mult_79_SUMB_13__12_) );
  FA_X1 u5_mult_79_S2_13_11 ( .A(u5_mult_79_ab_13__11_), .B(
        u5_mult_79_CARRYB_12__11_), .CI(u5_mult_79_SUMB_12__12_), .CO(
        u5_mult_79_CARRYB_13__11_), .S(u5_mult_79_SUMB_13__11_) );
  FA_X1 u5_mult_79_S2_13_10 ( .A(u5_mult_79_ab_13__10_), .B(
        u5_mult_79_CARRYB_12__10_), .CI(u5_mult_79_SUMB_12__11_), .CO(
        u5_mult_79_CARRYB_13__10_), .S(u5_mult_79_SUMB_13__10_) );
  FA_X1 u5_mult_79_S2_13_9 ( .A(u5_mult_79_ab_13__9_), .B(
        u5_mult_79_CARRYB_12__9_), .CI(u5_mult_79_SUMB_12__10_), .CO(
        u5_mult_79_CARRYB_13__9_), .S(u5_mult_79_SUMB_13__9_) );
  FA_X1 u5_mult_79_S2_13_8 ( .A(u5_mult_79_ab_13__8_), .B(
        u5_mult_79_CARRYB_12__8_), .CI(u5_mult_79_SUMB_12__9_), .CO(
        u5_mult_79_CARRYB_13__8_), .S(u5_mult_79_SUMB_13__8_) );
  FA_X1 u5_mult_79_S2_13_7 ( .A(u5_mult_79_ab_13__7_), .B(
        u5_mult_79_CARRYB_12__7_), .CI(u5_mult_79_SUMB_12__8_), .CO(
        u5_mult_79_CARRYB_13__7_), .S(u5_mult_79_SUMB_13__7_) );
  FA_X1 u5_mult_79_S2_13_6 ( .A(u5_mult_79_ab_13__6_), .B(
        u5_mult_79_CARRYB_12__6_), .CI(u5_mult_79_SUMB_12__7_), .CO(
        u5_mult_79_CARRYB_13__6_), .S(u5_mult_79_SUMB_13__6_) );
  FA_X1 u5_mult_79_S2_13_5 ( .A(u5_mult_79_ab_13__5_), .B(
        u5_mult_79_CARRYB_12__5_), .CI(u5_mult_79_SUMB_12__6_), .CO(
        u5_mult_79_CARRYB_13__5_), .S(u5_mult_79_SUMB_13__5_) );
  FA_X1 u5_mult_79_S2_13_4 ( .A(u5_mult_79_ab_13__4_), .B(
        u5_mult_79_CARRYB_12__4_), .CI(u5_mult_79_SUMB_12__5_), .CO(
        u5_mult_79_CARRYB_13__4_), .S(u5_mult_79_SUMB_13__4_) );
  FA_X1 u5_mult_79_S2_13_3 ( .A(u5_mult_79_ab_13__3_), .B(
        u5_mult_79_CARRYB_12__3_), .CI(u5_mult_79_SUMB_12__4_), .CO(
        u5_mult_79_CARRYB_13__3_), .S(u5_mult_79_SUMB_13__3_) );
  FA_X1 u5_mult_79_S2_13_2 ( .A(u5_mult_79_ab_13__2_), .B(
        u5_mult_79_CARRYB_12__2_), .CI(u5_mult_79_SUMB_12__3_), .CO(
        u5_mult_79_CARRYB_13__2_), .S(u5_mult_79_SUMB_13__2_) );
  FA_X1 u5_mult_79_S2_13_1 ( .A(u5_mult_79_ab_13__1_), .B(
        u5_mult_79_CARRYB_12__1_), .CI(u5_mult_79_SUMB_12__2_), .CO(
        u5_mult_79_CARRYB_13__1_), .S(u5_mult_79_SUMB_13__1_) );
  FA_X1 u5_mult_79_S1_13_0 ( .A(u5_mult_79_ab_13__0_), .B(
        u5_mult_79_CARRYB_12__0_), .CI(u5_mult_79_SUMB_12__1_), .CO(
        u5_mult_79_CARRYB_13__0_), .S(u5_N13) );
  FA_X1 u5_mult_79_S3_14_22 ( .A(u5_mult_79_ab_14__22_), .B(
        u5_mult_79_CARRYB_13__22_), .CI(u5_mult_79_ab_13__23_), .CO(
        u5_mult_79_CARRYB_14__22_), .S(u5_mult_79_SUMB_14__22_) );
  FA_X1 u5_mult_79_S2_14_21 ( .A(u5_mult_79_ab_14__21_), .B(
        u5_mult_79_CARRYB_13__21_), .CI(u5_mult_79_SUMB_13__22_), .CO(
        u5_mult_79_CARRYB_14__21_), .S(u5_mult_79_SUMB_14__21_) );
  FA_X1 u5_mult_79_S2_14_20 ( .A(u5_mult_79_ab_14__20_), .B(
        u5_mult_79_CARRYB_13__20_), .CI(u5_mult_79_SUMB_13__21_), .CO(
        u5_mult_79_CARRYB_14__20_), .S(u5_mult_79_SUMB_14__20_) );
  FA_X1 u5_mult_79_S2_14_19 ( .A(u5_mult_79_ab_14__19_), .B(
        u5_mult_79_CARRYB_13__19_), .CI(u5_mult_79_SUMB_13__20_), .CO(
        u5_mult_79_CARRYB_14__19_), .S(u5_mult_79_SUMB_14__19_) );
  FA_X1 u5_mult_79_S2_14_18 ( .A(u5_mult_79_ab_14__18_), .B(
        u5_mult_79_CARRYB_13__18_), .CI(u5_mult_79_SUMB_13__19_), .CO(
        u5_mult_79_CARRYB_14__18_), .S(u5_mult_79_SUMB_14__18_) );
  FA_X1 u5_mult_79_S2_14_17 ( .A(u5_mult_79_ab_14__17_), .B(
        u5_mult_79_CARRYB_13__17_), .CI(u5_mult_79_SUMB_13__18_), .CO(
        u5_mult_79_CARRYB_14__17_), .S(u5_mult_79_SUMB_14__17_) );
  FA_X1 u5_mult_79_S2_14_16 ( .A(u5_mult_79_ab_14__16_), .B(
        u5_mult_79_CARRYB_13__16_), .CI(u5_mult_79_SUMB_13__17_), .CO(
        u5_mult_79_CARRYB_14__16_), .S(u5_mult_79_SUMB_14__16_) );
  FA_X1 u5_mult_79_S2_14_15 ( .A(u5_mult_79_ab_14__15_), .B(
        u5_mult_79_CARRYB_13__15_), .CI(u5_mult_79_SUMB_13__16_), .CO(
        u5_mult_79_CARRYB_14__15_), .S(u5_mult_79_SUMB_14__15_) );
  FA_X1 u5_mult_79_S2_14_14 ( .A(u5_mult_79_ab_14__14_), .B(
        u5_mult_79_CARRYB_13__14_), .CI(u5_mult_79_SUMB_13__15_), .CO(
        u5_mult_79_CARRYB_14__14_), .S(u5_mult_79_SUMB_14__14_) );
  FA_X1 u5_mult_79_S2_14_13 ( .A(u5_mult_79_ab_14__13_), .B(
        u5_mult_79_CARRYB_13__13_), .CI(u5_mult_79_SUMB_13__14_), .CO(
        u5_mult_79_CARRYB_14__13_), .S(u5_mult_79_SUMB_14__13_) );
  FA_X1 u5_mult_79_S2_14_12 ( .A(u5_mult_79_ab_14__12_), .B(
        u5_mult_79_CARRYB_13__12_), .CI(u5_mult_79_SUMB_13__13_), .CO(
        u5_mult_79_CARRYB_14__12_), .S(u5_mult_79_SUMB_14__12_) );
  FA_X1 u5_mult_79_S2_14_11 ( .A(u5_mult_79_ab_14__11_), .B(
        u5_mult_79_CARRYB_13__11_), .CI(u5_mult_79_SUMB_13__12_), .CO(
        u5_mult_79_CARRYB_14__11_), .S(u5_mult_79_SUMB_14__11_) );
  FA_X1 u5_mult_79_S2_14_10 ( .A(u5_mult_79_ab_14__10_), .B(
        u5_mult_79_CARRYB_13__10_), .CI(u5_mult_79_SUMB_13__11_), .CO(
        u5_mult_79_CARRYB_14__10_), .S(u5_mult_79_SUMB_14__10_) );
  FA_X1 u5_mult_79_S2_14_9 ( .A(u5_mult_79_ab_14__9_), .B(
        u5_mult_79_CARRYB_13__9_), .CI(u5_mult_79_SUMB_13__10_), .CO(
        u5_mult_79_CARRYB_14__9_), .S(u5_mult_79_SUMB_14__9_) );
  FA_X1 u5_mult_79_S2_14_8 ( .A(u5_mult_79_ab_14__8_), .B(
        u5_mult_79_CARRYB_13__8_), .CI(u5_mult_79_SUMB_13__9_), .CO(
        u5_mult_79_CARRYB_14__8_), .S(u5_mult_79_SUMB_14__8_) );
  FA_X1 u5_mult_79_S2_14_7 ( .A(u5_mult_79_ab_14__7_), .B(
        u5_mult_79_CARRYB_13__7_), .CI(u5_mult_79_SUMB_13__8_), .CO(
        u5_mult_79_CARRYB_14__7_), .S(u5_mult_79_SUMB_14__7_) );
  FA_X1 u5_mult_79_S2_14_6 ( .A(u5_mult_79_ab_14__6_), .B(
        u5_mult_79_CARRYB_13__6_), .CI(u5_mult_79_SUMB_13__7_), .CO(
        u5_mult_79_CARRYB_14__6_), .S(u5_mult_79_SUMB_14__6_) );
  FA_X1 u5_mult_79_S2_14_5 ( .A(u5_mult_79_ab_14__5_), .B(
        u5_mult_79_CARRYB_13__5_), .CI(u5_mult_79_SUMB_13__6_), .CO(
        u5_mult_79_CARRYB_14__5_), .S(u5_mult_79_SUMB_14__5_) );
  FA_X1 u5_mult_79_S2_14_4 ( .A(u5_mult_79_ab_14__4_), .B(
        u5_mult_79_CARRYB_13__4_), .CI(u5_mult_79_SUMB_13__5_), .CO(
        u5_mult_79_CARRYB_14__4_), .S(u5_mult_79_SUMB_14__4_) );
  FA_X1 u5_mult_79_S2_14_3 ( .A(u5_mult_79_ab_14__3_), .B(
        u5_mult_79_CARRYB_13__3_), .CI(u5_mult_79_SUMB_13__4_), .CO(
        u5_mult_79_CARRYB_14__3_), .S(u5_mult_79_SUMB_14__3_) );
  FA_X1 u5_mult_79_S2_14_2 ( .A(u5_mult_79_ab_14__2_), .B(
        u5_mult_79_CARRYB_13__2_), .CI(u5_mult_79_SUMB_13__3_), .CO(
        u5_mult_79_CARRYB_14__2_), .S(u5_mult_79_SUMB_14__2_) );
  FA_X1 u5_mult_79_S2_14_1 ( .A(u5_mult_79_ab_14__1_), .B(
        u5_mult_79_CARRYB_13__1_), .CI(u5_mult_79_SUMB_13__2_), .CO(
        u5_mult_79_CARRYB_14__1_), .S(u5_mult_79_SUMB_14__1_) );
  FA_X1 u5_mult_79_S1_14_0 ( .A(u5_mult_79_ab_14__0_), .B(
        u5_mult_79_CARRYB_13__0_), .CI(u5_mult_79_SUMB_13__1_), .CO(
        u5_mult_79_CARRYB_14__0_), .S(u5_N14) );
  FA_X1 u5_mult_79_S3_15_22 ( .A(u5_mult_79_ab_15__22_), .B(
        u5_mult_79_CARRYB_14__22_), .CI(u5_mult_79_ab_14__23_), .CO(
        u5_mult_79_CARRYB_15__22_), .S(u5_mult_79_SUMB_15__22_) );
  FA_X1 u5_mult_79_S2_15_21 ( .A(u5_mult_79_ab_15__21_), .B(
        u5_mult_79_CARRYB_14__21_), .CI(u5_mult_79_SUMB_14__22_), .CO(
        u5_mult_79_CARRYB_15__21_), .S(u5_mult_79_SUMB_15__21_) );
  FA_X1 u5_mult_79_S2_15_20 ( .A(u5_mult_79_ab_15__20_), .B(
        u5_mult_79_CARRYB_14__20_), .CI(u5_mult_79_SUMB_14__21_), .CO(
        u5_mult_79_CARRYB_15__20_), .S(u5_mult_79_SUMB_15__20_) );
  FA_X1 u5_mult_79_S2_15_19 ( .A(u5_mult_79_ab_15__19_), .B(
        u5_mult_79_CARRYB_14__19_), .CI(u5_mult_79_SUMB_14__20_), .CO(
        u5_mult_79_CARRYB_15__19_), .S(u5_mult_79_SUMB_15__19_) );
  FA_X1 u5_mult_79_S2_15_18 ( .A(u5_mult_79_ab_15__18_), .B(
        u5_mult_79_CARRYB_14__18_), .CI(u5_mult_79_SUMB_14__19_), .CO(
        u5_mult_79_CARRYB_15__18_), .S(u5_mult_79_SUMB_15__18_) );
  FA_X1 u5_mult_79_S2_15_17 ( .A(u5_mult_79_ab_15__17_), .B(
        u5_mult_79_CARRYB_14__17_), .CI(u5_mult_79_SUMB_14__18_), .CO(
        u5_mult_79_CARRYB_15__17_), .S(u5_mult_79_SUMB_15__17_) );
  FA_X1 u5_mult_79_S2_15_16 ( .A(u5_mult_79_ab_15__16_), .B(
        u5_mult_79_CARRYB_14__16_), .CI(u5_mult_79_SUMB_14__17_), .CO(
        u5_mult_79_CARRYB_15__16_), .S(u5_mult_79_SUMB_15__16_) );
  FA_X1 u5_mult_79_S2_15_15 ( .A(u5_mult_79_ab_15__15_), .B(
        u5_mult_79_CARRYB_14__15_), .CI(u5_mult_79_SUMB_14__16_), .CO(
        u5_mult_79_CARRYB_15__15_), .S(u5_mult_79_SUMB_15__15_) );
  FA_X1 u5_mult_79_S2_15_14 ( .A(u5_mult_79_ab_15__14_), .B(
        u5_mult_79_CARRYB_14__14_), .CI(u5_mult_79_SUMB_14__15_), .CO(
        u5_mult_79_CARRYB_15__14_), .S(u5_mult_79_SUMB_15__14_) );
  FA_X1 u5_mult_79_S2_15_13 ( .A(u5_mult_79_ab_15__13_), .B(
        u5_mult_79_CARRYB_14__13_), .CI(u5_mult_79_SUMB_14__14_), .CO(
        u5_mult_79_CARRYB_15__13_), .S(u5_mult_79_SUMB_15__13_) );
  FA_X1 u5_mult_79_S2_15_12 ( .A(u5_mult_79_ab_15__12_), .B(
        u5_mult_79_CARRYB_14__12_), .CI(u5_mult_79_SUMB_14__13_), .CO(
        u5_mult_79_CARRYB_15__12_), .S(u5_mult_79_SUMB_15__12_) );
  FA_X1 u5_mult_79_S2_15_11 ( .A(u5_mult_79_ab_15__11_), .B(
        u5_mult_79_CARRYB_14__11_), .CI(u5_mult_79_SUMB_14__12_), .CO(
        u5_mult_79_CARRYB_15__11_), .S(u5_mult_79_SUMB_15__11_) );
  FA_X1 u5_mult_79_S2_15_10 ( .A(u5_mult_79_ab_15__10_), .B(
        u5_mult_79_CARRYB_14__10_), .CI(u5_mult_79_SUMB_14__11_), .CO(
        u5_mult_79_CARRYB_15__10_), .S(u5_mult_79_SUMB_15__10_) );
  FA_X1 u5_mult_79_S2_15_9 ( .A(u5_mult_79_ab_15__9_), .B(
        u5_mult_79_CARRYB_14__9_), .CI(u5_mult_79_SUMB_14__10_), .CO(
        u5_mult_79_CARRYB_15__9_), .S(u5_mult_79_SUMB_15__9_) );
  FA_X1 u5_mult_79_S2_15_8 ( .A(u5_mult_79_ab_15__8_), .B(
        u5_mult_79_CARRYB_14__8_), .CI(u5_mult_79_SUMB_14__9_), .CO(
        u5_mult_79_CARRYB_15__8_), .S(u5_mult_79_SUMB_15__8_) );
  FA_X1 u5_mult_79_S2_15_7 ( .A(u5_mult_79_ab_15__7_), .B(
        u5_mult_79_CARRYB_14__7_), .CI(u5_mult_79_SUMB_14__8_), .CO(
        u5_mult_79_CARRYB_15__7_), .S(u5_mult_79_SUMB_15__7_) );
  FA_X1 u5_mult_79_S2_15_6 ( .A(u5_mult_79_ab_15__6_), .B(
        u5_mult_79_CARRYB_14__6_), .CI(u5_mult_79_SUMB_14__7_), .CO(
        u5_mult_79_CARRYB_15__6_), .S(u5_mult_79_SUMB_15__6_) );
  FA_X1 u5_mult_79_S2_15_5 ( .A(u5_mult_79_ab_15__5_), .B(
        u5_mult_79_CARRYB_14__5_), .CI(u5_mult_79_SUMB_14__6_), .CO(
        u5_mult_79_CARRYB_15__5_), .S(u5_mult_79_SUMB_15__5_) );
  FA_X1 u5_mult_79_S2_15_4 ( .A(u5_mult_79_ab_15__4_), .B(
        u5_mult_79_CARRYB_14__4_), .CI(u5_mult_79_SUMB_14__5_), .CO(
        u5_mult_79_CARRYB_15__4_), .S(u5_mult_79_SUMB_15__4_) );
  FA_X1 u5_mult_79_S2_15_3 ( .A(u5_mult_79_ab_15__3_), .B(
        u5_mult_79_CARRYB_14__3_), .CI(u5_mult_79_SUMB_14__4_), .CO(
        u5_mult_79_CARRYB_15__3_), .S(u5_mult_79_SUMB_15__3_) );
  FA_X1 u5_mult_79_S2_15_2 ( .A(u5_mult_79_ab_15__2_), .B(
        u5_mult_79_CARRYB_14__2_), .CI(u5_mult_79_SUMB_14__3_), .CO(
        u5_mult_79_CARRYB_15__2_), .S(u5_mult_79_SUMB_15__2_) );
  FA_X1 u5_mult_79_S2_15_1 ( .A(u5_mult_79_ab_15__1_), .B(
        u5_mult_79_CARRYB_14__1_), .CI(u5_mult_79_SUMB_14__2_), .CO(
        u5_mult_79_CARRYB_15__1_), .S(u5_mult_79_SUMB_15__1_) );
  FA_X1 u5_mult_79_S1_15_0 ( .A(u5_mult_79_ab_15__0_), .B(
        u5_mult_79_CARRYB_14__0_), .CI(u5_mult_79_SUMB_14__1_), .CO(
        u5_mult_79_CARRYB_15__0_), .S(u5_N15) );
  FA_X1 u5_mult_79_S3_16_22 ( .A(u5_mult_79_ab_16__22_), .B(
        u5_mult_79_CARRYB_15__22_), .CI(u5_mult_79_ab_15__23_), .CO(
        u5_mult_79_CARRYB_16__22_), .S(u5_mult_79_SUMB_16__22_) );
  FA_X1 u5_mult_79_S2_16_21 ( .A(u5_mult_79_ab_16__21_), .B(
        u5_mult_79_CARRYB_15__21_), .CI(u5_mult_79_SUMB_15__22_), .CO(
        u5_mult_79_CARRYB_16__21_), .S(u5_mult_79_SUMB_16__21_) );
  FA_X1 u5_mult_79_S2_16_20 ( .A(u5_mult_79_ab_16__20_), .B(
        u5_mult_79_CARRYB_15__20_), .CI(u5_mult_79_SUMB_15__21_), .CO(
        u5_mult_79_CARRYB_16__20_), .S(u5_mult_79_SUMB_16__20_) );
  FA_X1 u5_mult_79_S2_16_19 ( .A(u5_mult_79_ab_16__19_), .B(
        u5_mult_79_CARRYB_15__19_), .CI(u5_mult_79_SUMB_15__20_), .CO(
        u5_mult_79_CARRYB_16__19_), .S(u5_mult_79_SUMB_16__19_) );
  FA_X1 u5_mult_79_S2_16_18 ( .A(u5_mult_79_ab_16__18_), .B(
        u5_mult_79_CARRYB_15__18_), .CI(u5_mult_79_SUMB_15__19_), .CO(
        u5_mult_79_CARRYB_16__18_), .S(u5_mult_79_SUMB_16__18_) );
  FA_X1 u5_mult_79_S2_16_17 ( .A(u5_mult_79_ab_16__17_), .B(
        u5_mult_79_CARRYB_15__17_), .CI(u5_mult_79_SUMB_15__18_), .CO(
        u5_mult_79_CARRYB_16__17_), .S(u5_mult_79_SUMB_16__17_) );
  FA_X1 u5_mult_79_S2_16_16 ( .A(u5_mult_79_ab_16__16_), .B(
        u5_mult_79_CARRYB_15__16_), .CI(u5_mult_79_SUMB_15__17_), .CO(
        u5_mult_79_CARRYB_16__16_), .S(u5_mult_79_SUMB_16__16_) );
  FA_X1 u5_mult_79_S2_16_15 ( .A(u5_mult_79_ab_16__15_), .B(
        u5_mult_79_CARRYB_15__15_), .CI(u5_mult_79_SUMB_15__16_), .CO(
        u5_mult_79_CARRYB_16__15_), .S(u5_mult_79_SUMB_16__15_) );
  FA_X1 u5_mult_79_S2_16_14 ( .A(u5_mult_79_ab_16__14_), .B(
        u5_mult_79_CARRYB_15__14_), .CI(u5_mult_79_SUMB_15__15_), .CO(
        u5_mult_79_CARRYB_16__14_), .S(u5_mult_79_SUMB_16__14_) );
  FA_X1 u5_mult_79_S2_16_13 ( .A(u5_mult_79_ab_16__13_), .B(
        u5_mult_79_CARRYB_15__13_), .CI(u5_mult_79_SUMB_15__14_), .CO(
        u5_mult_79_CARRYB_16__13_), .S(u5_mult_79_SUMB_16__13_) );
  FA_X1 u5_mult_79_S2_16_12 ( .A(u5_mult_79_ab_16__12_), .B(
        u5_mult_79_CARRYB_15__12_), .CI(u5_mult_79_SUMB_15__13_), .CO(
        u5_mult_79_CARRYB_16__12_), .S(u5_mult_79_SUMB_16__12_) );
  FA_X1 u5_mult_79_S2_16_11 ( .A(u5_mult_79_ab_16__11_), .B(
        u5_mult_79_CARRYB_15__11_), .CI(u5_mult_79_SUMB_15__12_), .CO(
        u5_mult_79_CARRYB_16__11_), .S(u5_mult_79_SUMB_16__11_) );
  FA_X1 u5_mult_79_S2_16_10 ( .A(u5_mult_79_ab_16__10_), .B(
        u5_mult_79_CARRYB_15__10_), .CI(u5_mult_79_SUMB_15__11_), .CO(
        u5_mult_79_CARRYB_16__10_), .S(u5_mult_79_SUMB_16__10_) );
  FA_X1 u5_mult_79_S2_16_9 ( .A(u5_mult_79_ab_16__9_), .B(
        u5_mult_79_CARRYB_15__9_), .CI(u5_mult_79_SUMB_15__10_), .CO(
        u5_mult_79_CARRYB_16__9_), .S(u5_mult_79_SUMB_16__9_) );
  FA_X1 u5_mult_79_S2_16_8 ( .A(u5_mult_79_ab_16__8_), .B(
        u5_mult_79_CARRYB_15__8_), .CI(u5_mult_79_SUMB_15__9_), .CO(
        u5_mult_79_CARRYB_16__8_), .S(u5_mult_79_SUMB_16__8_) );
  FA_X1 u5_mult_79_S2_16_7 ( .A(u5_mult_79_ab_16__7_), .B(
        u5_mult_79_CARRYB_15__7_), .CI(u5_mult_79_SUMB_15__8_), .CO(
        u5_mult_79_CARRYB_16__7_), .S(u5_mult_79_SUMB_16__7_) );
  FA_X1 u5_mult_79_S2_16_6 ( .A(u5_mult_79_ab_16__6_), .B(
        u5_mult_79_CARRYB_15__6_), .CI(u5_mult_79_SUMB_15__7_), .CO(
        u5_mult_79_CARRYB_16__6_), .S(u5_mult_79_SUMB_16__6_) );
  FA_X1 u5_mult_79_S2_16_5 ( .A(u5_mult_79_ab_16__5_), .B(
        u5_mult_79_CARRYB_15__5_), .CI(u5_mult_79_SUMB_15__6_), .CO(
        u5_mult_79_CARRYB_16__5_), .S(u5_mult_79_SUMB_16__5_) );
  FA_X1 u5_mult_79_S2_16_4 ( .A(u5_mult_79_ab_16__4_), .B(
        u5_mult_79_CARRYB_15__4_), .CI(u5_mult_79_SUMB_15__5_), .CO(
        u5_mult_79_CARRYB_16__4_), .S(u5_mult_79_SUMB_16__4_) );
  FA_X1 u5_mult_79_S2_16_3 ( .A(u5_mult_79_ab_16__3_), .B(
        u5_mult_79_CARRYB_15__3_), .CI(u5_mult_79_SUMB_15__4_), .CO(
        u5_mult_79_CARRYB_16__3_), .S(u5_mult_79_SUMB_16__3_) );
  FA_X1 u5_mult_79_S2_16_2 ( .A(u5_mult_79_ab_16__2_), .B(
        u5_mult_79_CARRYB_15__2_), .CI(u5_mult_79_SUMB_15__3_), .CO(
        u5_mult_79_CARRYB_16__2_), .S(u5_mult_79_SUMB_16__2_) );
  FA_X1 u5_mult_79_S2_16_1 ( .A(u5_mult_79_ab_16__1_), .B(
        u5_mult_79_CARRYB_15__1_), .CI(u5_mult_79_SUMB_15__2_), .CO(
        u5_mult_79_CARRYB_16__1_), .S(u5_mult_79_SUMB_16__1_) );
  FA_X1 u5_mult_79_S1_16_0 ( .A(u5_mult_79_ab_16__0_), .B(
        u5_mult_79_CARRYB_15__0_), .CI(u5_mult_79_SUMB_15__1_), .CO(
        u5_mult_79_CARRYB_16__0_), .S(u5_N16) );
  FA_X1 u5_mult_79_S3_17_22 ( .A(u5_mult_79_ab_17__22_), .B(
        u5_mult_79_CARRYB_16__22_), .CI(u5_mult_79_ab_16__23_), .CO(
        u5_mult_79_CARRYB_17__22_), .S(u5_mult_79_SUMB_17__22_) );
  FA_X1 u5_mult_79_S2_17_21 ( .A(u5_mult_79_ab_17__21_), .B(
        u5_mult_79_CARRYB_16__21_), .CI(u5_mult_79_SUMB_16__22_), .CO(
        u5_mult_79_CARRYB_17__21_), .S(u5_mult_79_SUMB_17__21_) );
  FA_X1 u5_mult_79_S2_17_20 ( .A(u5_mult_79_ab_17__20_), .B(
        u5_mult_79_CARRYB_16__20_), .CI(u5_mult_79_SUMB_16__21_), .CO(
        u5_mult_79_CARRYB_17__20_), .S(u5_mult_79_SUMB_17__20_) );
  FA_X1 u5_mult_79_S2_17_19 ( .A(u5_mult_79_ab_17__19_), .B(
        u5_mult_79_CARRYB_16__19_), .CI(u5_mult_79_SUMB_16__20_), .CO(
        u5_mult_79_CARRYB_17__19_), .S(u5_mult_79_SUMB_17__19_) );
  FA_X1 u5_mult_79_S2_17_18 ( .A(u5_mult_79_ab_17__18_), .B(
        u5_mult_79_CARRYB_16__18_), .CI(u5_mult_79_SUMB_16__19_), .CO(
        u5_mult_79_CARRYB_17__18_), .S(u5_mult_79_SUMB_17__18_) );
  FA_X1 u5_mult_79_S2_17_17 ( .A(u5_mult_79_ab_17__17_), .B(
        u5_mult_79_CARRYB_16__17_), .CI(u5_mult_79_SUMB_16__18_), .CO(
        u5_mult_79_CARRYB_17__17_), .S(u5_mult_79_SUMB_17__17_) );
  FA_X1 u5_mult_79_S2_17_16 ( .A(u5_mult_79_ab_17__16_), .B(
        u5_mult_79_CARRYB_16__16_), .CI(u5_mult_79_SUMB_16__17_), .CO(
        u5_mult_79_CARRYB_17__16_), .S(u5_mult_79_SUMB_17__16_) );
  FA_X1 u5_mult_79_S2_17_15 ( .A(u5_mult_79_ab_17__15_), .B(
        u5_mult_79_CARRYB_16__15_), .CI(u5_mult_79_SUMB_16__16_), .CO(
        u5_mult_79_CARRYB_17__15_), .S(u5_mult_79_SUMB_17__15_) );
  FA_X1 u5_mult_79_S2_17_14 ( .A(u5_mult_79_ab_17__14_), .B(
        u5_mult_79_CARRYB_16__14_), .CI(u5_mult_79_SUMB_16__15_), .CO(
        u5_mult_79_CARRYB_17__14_), .S(u5_mult_79_SUMB_17__14_) );
  FA_X1 u5_mult_79_S2_17_13 ( .A(u5_mult_79_ab_17__13_), .B(
        u5_mult_79_CARRYB_16__13_), .CI(u5_mult_79_SUMB_16__14_), .CO(
        u5_mult_79_CARRYB_17__13_), .S(u5_mult_79_SUMB_17__13_) );
  FA_X1 u5_mult_79_S2_17_12 ( .A(u5_mult_79_ab_17__12_), .B(
        u5_mult_79_CARRYB_16__12_), .CI(u5_mult_79_SUMB_16__13_), .CO(
        u5_mult_79_CARRYB_17__12_), .S(u5_mult_79_SUMB_17__12_) );
  FA_X1 u5_mult_79_S2_17_11 ( .A(u5_mult_79_ab_17__11_), .B(
        u5_mult_79_CARRYB_16__11_), .CI(u5_mult_79_SUMB_16__12_), .CO(
        u5_mult_79_CARRYB_17__11_), .S(u5_mult_79_SUMB_17__11_) );
  FA_X1 u5_mult_79_S2_17_10 ( .A(u5_mult_79_ab_17__10_), .B(
        u5_mult_79_CARRYB_16__10_), .CI(u5_mult_79_SUMB_16__11_), .CO(
        u5_mult_79_CARRYB_17__10_), .S(u5_mult_79_SUMB_17__10_) );
  FA_X1 u5_mult_79_S2_17_9 ( .A(u5_mult_79_ab_17__9_), .B(
        u5_mult_79_CARRYB_16__9_), .CI(u5_mult_79_SUMB_16__10_), .CO(
        u5_mult_79_CARRYB_17__9_), .S(u5_mult_79_SUMB_17__9_) );
  FA_X1 u5_mult_79_S2_17_8 ( .A(u5_mult_79_ab_17__8_), .B(
        u5_mult_79_CARRYB_16__8_), .CI(u5_mult_79_SUMB_16__9_), .CO(
        u5_mult_79_CARRYB_17__8_), .S(u5_mult_79_SUMB_17__8_) );
  FA_X1 u5_mult_79_S2_17_7 ( .A(u5_mult_79_ab_17__7_), .B(
        u5_mult_79_CARRYB_16__7_), .CI(u5_mult_79_SUMB_16__8_), .CO(
        u5_mult_79_CARRYB_17__7_), .S(u5_mult_79_SUMB_17__7_) );
  FA_X1 u5_mult_79_S2_17_6 ( .A(u5_mult_79_ab_17__6_), .B(
        u5_mult_79_CARRYB_16__6_), .CI(u5_mult_79_SUMB_16__7_), .CO(
        u5_mult_79_CARRYB_17__6_), .S(u5_mult_79_SUMB_17__6_) );
  FA_X1 u5_mult_79_S2_17_5 ( .A(u5_mult_79_ab_17__5_), .B(
        u5_mult_79_CARRYB_16__5_), .CI(u5_mult_79_SUMB_16__6_), .CO(
        u5_mult_79_CARRYB_17__5_), .S(u5_mult_79_SUMB_17__5_) );
  FA_X1 u5_mult_79_S2_17_4 ( .A(u5_mult_79_ab_17__4_), .B(
        u5_mult_79_CARRYB_16__4_), .CI(u5_mult_79_SUMB_16__5_), .CO(
        u5_mult_79_CARRYB_17__4_), .S(u5_mult_79_SUMB_17__4_) );
  FA_X1 u5_mult_79_S2_17_3 ( .A(u5_mult_79_ab_17__3_), .B(
        u5_mult_79_CARRYB_16__3_), .CI(u5_mult_79_SUMB_16__4_), .CO(
        u5_mult_79_CARRYB_17__3_), .S(u5_mult_79_SUMB_17__3_) );
  FA_X1 u5_mult_79_S2_17_2 ( .A(u5_mult_79_ab_17__2_), .B(
        u5_mult_79_CARRYB_16__2_), .CI(u5_mult_79_SUMB_16__3_), .CO(
        u5_mult_79_CARRYB_17__2_), .S(u5_mult_79_SUMB_17__2_) );
  FA_X1 u5_mult_79_S2_17_1 ( .A(u5_mult_79_ab_17__1_), .B(
        u5_mult_79_CARRYB_16__1_), .CI(u5_mult_79_SUMB_16__2_), .CO(
        u5_mult_79_CARRYB_17__1_), .S(u5_mult_79_SUMB_17__1_) );
  FA_X1 u5_mult_79_S1_17_0 ( .A(u5_mult_79_ab_17__0_), .B(
        u5_mult_79_CARRYB_16__0_), .CI(u5_mult_79_SUMB_16__1_), .CO(
        u5_mult_79_CARRYB_17__0_), .S(u5_N17) );
  FA_X1 u5_mult_79_S3_18_22 ( .A(u5_mult_79_ab_18__22_), .B(
        u5_mult_79_CARRYB_17__22_), .CI(u5_mult_79_ab_17__23_), .CO(
        u5_mult_79_CARRYB_18__22_), .S(u5_mult_79_SUMB_18__22_) );
  FA_X1 u5_mult_79_S2_18_21 ( .A(u5_mult_79_ab_18__21_), .B(
        u5_mult_79_CARRYB_17__21_), .CI(u5_mult_79_SUMB_17__22_), .CO(
        u5_mult_79_CARRYB_18__21_), .S(u5_mult_79_SUMB_18__21_) );
  FA_X1 u5_mult_79_S2_18_20 ( .A(u5_mult_79_ab_18__20_), .B(
        u5_mult_79_CARRYB_17__20_), .CI(u5_mult_79_SUMB_17__21_), .CO(
        u5_mult_79_CARRYB_18__20_), .S(u5_mult_79_SUMB_18__20_) );
  FA_X1 u5_mult_79_S2_18_19 ( .A(u5_mult_79_ab_18__19_), .B(
        u5_mult_79_CARRYB_17__19_), .CI(u5_mult_79_SUMB_17__20_), .CO(
        u5_mult_79_CARRYB_18__19_), .S(u5_mult_79_SUMB_18__19_) );
  FA_X1 u5_mult_79_S2_18_18 ( .A(u5_mult_79_ab_18__18_), .B(
        u5_mult_79_CARRYB_17__18_), .CI(u5_mult_79_SUMB_17__19_), .CO(
        u5_mult_79_CARRYB_18__18_), .S(u5_mult_79_SUMB_18__18_) );
  FA_X1 u5_mult_79_S2_18_17 ( .A(u5_mult_79_ab_18__17_), .B(
        u5_mult_79_CARRYB_17__17_), .CI(u5_mult_79_SUMB_17__18_), .CO(
        u5_mult_79_CARRYB_18__17_), .S(u5_mult_79_SUMB_18__17_) );
  FA_X1 u5_mult_79_S2_18_16 ( .A(u5_mult_79_ab_18__16_), .B(
        u5_mult_79_CARRYB_17__16_), .CI(u5_mult_79_SUMB_17__17_), .CO(
        u5_mult_79_CARRYB_18__16_), .S(u5_mult_79_SUMB_18__16_) );
  FA_X1 u5_mult_79_S2_18_15 ( .A(u5_mult_79_ab_18__15_), .B(
        u5_mult_79_CARRYB_17__15_), .CI(u5_mult_79_SUMB_17__16_), .CO(
        u5_mult_79_CARRYB_18__15_), .S(u5_mult_79_SUMB_18__15_) );
  FA_X1 u5_mult_79_S2_18_14 ( .A(u5_mult_79_ab_18__14_), .B(
        u5_mult_79_CARRYB_17__14_), .CI(u5_mult_79_SUMB_17__15_), .CO(
        u5_mult_79_CARRYB_18__14_), .S(u5_mult_79_SUMB_18__14_) );
  FA_X1 u5_mult_79_S2_18_13 ( .A(u5_mult_79_ab_18__13_), .B(
        u5_mult_79_CARRYB_17__13_), .CI(u5_mult_79_SUMB_17__14_), .CO(
        u5_mult_79_CARRYB_18__13_), .S(u5_mult_79_SUMB_18__13_) );
  FA_X1 u5_mult_79_S2_18_12 ( .A(u5_mult_79_ab_18__12_), .B(
        u5_mult_79_CARRYB_17__12_), .CI(u5_mult_79_SUMB_17__13_), .CO(
        u5_mult_79_CARRYB_18__12_), .S(u5_mult_79_SUMB_18__12_) );
  FA_X1 u5_mult_79_S2_18_11 ( .A(u5_mult_79_ab_18__11_), .B(
        u5_mult_79_CARRYB_17__11_), .CI(u5_mult_79_SUMB_17__12_), .CO(
        u5_mult_79_CARRYB_18__11_), .S(u5_mult_79_SUMB_18__11_) );
  FA_X1 u5_mult_79_S2_18_10 ( .A(u5_mult_79_ab_18__10_), .B(
        u5_mult_79_CARRYB_17__10_), .CI(u5_mult_79_SUMB_17__11_), .CO(
        u5_mult_79_CARRYB_18__10_), .S(u5_mult_79_SUMB_18__10_) );
  FA_X1 u5_mult_79_S2_18_9 ( .A(u5_mult_79_ab_18__9_), .B(
        u5_mult_79_CARRYB_17__9_), .CI(u5_mult_79_SUMB_17__10_), .CO(
        u5_mult_79_CARRYB_18__9_), .S(u5_mult_79_SUMB_18__9_) );
  FA_X1 u5_mult_79_S2_18_8 ( .A(u5_mult_79_ab_18__8_), .B(
        u5_mult_79_CARRYB_17__8_), .CI(u5_mult_79_SUMB_17__9_), .CO(
        u5_mult_79_CARRYB_18__8_), .S(u5_mult_79_SUMB_18__8_) );
  FA_X1 u5_mult_79_S2_18_7 ( .A(u5_mult_79_ab_18__7_), .B(
        u5_mult_79_CARRYB_17__7_), .CI(u5_mult_79_SUMB_17__8_), .CO(
        u5_mult_79_CARRYB_18__7_), .S(u5_mult_79_SUMB_18__7_) );
  FA_X1 u5_mult_79_S2_18_6 ( .A(u5_mult_79_ab_18__6_), .B(
        u5_mult_79_CARRYB_17__6_), .CI(u5_mult_79_SUMB_17__7_), .CO(
        u5_mult_79_CARRYB_18__6_), .S(u5_mult_79_SUMB_18__6_) );
  FA_X1 u5_mult_79_S2_18_5 ( .A(u5_mult_79_ab_18__5_), .B(
        u5_mult_79_CARRYB_17__5_), .CI(u5_mult_79_SUMB_17__6_), .CO(
        u5_mult_79_CARRYB_18__5_), .S(u5_mult_79_SUMB_18__5_) );
  FA_X1 u5_mult_79_S2_18_4 ( .A(u5_mult_79_ab_18__4_), .B(
        u5_mult_79_CARRYB_17__4_), .CI(u5_mult_79_SUMB_17__5_), .CO(
        u5_mult_79_CARRYB_18__4_), .S(u5_mult_79_SUMB_18__4_) );
  FA_X1 u5_mult_79_S2_18_3 ( .A(u5_mult_79_ab_18__3_), .B(
        u5_mult_79_CARRYB_17__3_), .CI(u5_mult_79_SUMB_17__4_), .CO(
        u5_mult_79_CARRYB_18__3_), .S(u5_mult_79_SUMB_18__3_) );
  FA_X1 u5_mult_79_S2_18_2 ( .A(u5_mult_79_ab_18__2_), .B(
        u5_mult_79_CARRYB_17__2_), .CI(u5_mult_79_SUMB_17__3_), .CO(
        u5_mult_79_CARRYB_18__2_), .S(u5_mult_79_SUMB_18__2_) );
  FA_X1 u5_mult_79_S2_18_1 ( .A(u5_mult_79_ab_18__1_), .B(
        u5_mult_79_CARRYB_17__1_), .CI(u5_mult_79_SUMB_17__2_), .CO(
        u5_mult_79_CARRYB_18__1_), .S(u5_mult_79_SUMB_18__1_) );
  FA_X1 u5_mult_79_S1_18_0 ( .A(u5_mult_79_ab_18__0_), .B(
        u5_mult_79_CARRYB_17__0_), .CI(u5_mult_79_SUMB_17__1_), .CO(
        u5_mult_79_CARRYB_18__0_), .S(u5_N18) );
  FA_X1 u5_mult_79_S3_19_22 ( .A(u5_mult_79_ab_19__22_), .B(
        u5_mult_79_CARRYB_18__22_), .CI(u5_mult_79_ab_18__23_), .CO(
        u5_mult_79_CARRYB_19__22_), .S(u5_mult_79_SUMB_19__22_) );
  FA_X1 u5_mult_79_S2_19_21 ( .A(u5_mult_79_ab_19__21_), .B(
        u5_mult_79_CARRYB_18__21_), .CI(u5_mult_79_SUMB_18__22_), .CO(
        u5_mult_79_CARRYB_19__21_), .S(u5_mult_79_SUMB_19__21_) );
  FA_X1 u5_mult_79_S2_19_20 ( .A(u5_mult_79_ab_19__20_), .B(
        u5_mult_79_CARRYB_18__20_), .CI(u5_mult_79_SUMB_18__21_), .CO(
        u5_mult_79_CARRYB_19__20_), .S(u5_mult_79_SUMB_19__20_) );
  FA_X1 u5_mult_79_S2_19_19 ( .A(u5_mult_79_ab_19__19_), .B(
        u5_mult_79_CARRYB_18__19_), .CI(u5_mult_79_SUMB_18__20_), .CO(
        u5_mult_79_CARRYB_19__19_), .S(u5_mult_79_SUMB_19__19_) );
  FA_X1 u5_mult_79_S2_19_18 ( .A(u5_mult_79_ab_19__18_), .B(
        u5_mult_79_CARRYB_18__18_), .CI(u5_mult_79_SUMB_18__19_), .CO(
        u5_mult_79_CARRYB_19__18_), .S(u5_mult_79_SUMB_19__18_) );
  FA_X1 u5_mult_79_S2_19_17 ( .A(u5_mult_79_ab_19__17_), .B(
        u5_mult_79_CARRYB_18__17_), .CI(u5_mult_79_SUMB_18__18_), .CO(
        u5_mult_79_CARRYB_19__17_), .S(u5_mult_79_SUMB_19__17_) );
  FA_X1 u5_mult_79_S2_19_16 ( .A(u5_mult_79_ab_19__16_), .B(
        u5_mult_79_CARRYB_18__16_), .CI(u5_mult_79_SUMB_18__17_), .CO(
        u5_mult_79_CARRYB_19__16_), .S(u5_mult_79_SUMB_19__16_) );
  FA_X1 u5_mult_79_S2_19_15 ( .A(u5_mult_79_ab_19__15_), .B(
        u5_mult_79_CARRYB_18__15_), .CI(u5_mult_79_SUMB_18__16_), .CO(
        u5_mult_79_CARRYB_19__15_), .S(u5_mult_79_SUMB_19__15_) );
  FA_X1 u5_mult_79_S2_19_14 ( .A(u5_mult_79_ab_19__14_), .B(
        u5_mult_79_CARRYB_18__14_), .CI(u5_mult_79_SUMB_18__15_), .CO(
        u5_mult_79_CARRYB_19__14_), .S(u5_mult_79_SUMB_19__14_) );
  FA_X1 u5_mult_79_S2_19_13 ( .A(u5_mult_79_ab_19__13_), .B(
        u5_mult_79_CARRYB_18__13_), .CI(u5_mult_79_SUMB_18__14_), .CO(
        u5_mult_79_CARRYB_19__13_), .S(u5_mult_79_SUMB_19__13_) );
  FA_X1 u5_mult_79_S2_19_12 ( .A(u5_mult_79_ab_19__12_), .B(
        u5_mult_79_CARRYB_18__12_), .CI(u5_mult_79_SUMB_18__13_), .CO(
        u5_mult_79_CARRYB_19__12_), .S(u5_mult_79_SUMB_19__12_) );
  FA_X1 u5_mult_79_S2_19_11 ( .A(u5_mult_79_ab_19__11_), .B(
        u5_mult_79_CARRYB_18__11_), .CI(u5_mult_79_SUMB_18__12_), .CO(
        u5_mult_79_CARRYB_19__11_), .S(u5_mult_79_SUMB_19__11_) );
  FA_X1 u5_mult_79_S2_19_10 ( .A(u5_mult_79_ab_19__10_), .B(
        u5_mult_79_CARRYB_18__10_), .CI(u5_mult_79_SUMB_18__11_), .CO(
        u5_mult_79_CARRYB_19__10_), .S(u5_mult_79_SUMB_19__10_) );
  FA_X1 u5_mult_79_S2_19_9 ( .A(u5_mult_79_ab_19__9_), .B(
        u5_mult_79_CARRYB_18__9_), .CI(u5_mult_79_SUMB_18__10_), .CO(
        u5_mult_79_CARRYB_19__9_), .S(u5_mult_79_SUMB_19__9_) );
  FA_X1 u5_mult_79_S2_19_8 ( .A(u5_mult_79_ab_19__8_), .B(
        u5_mult_79_CARRYB_18__8_), .CI(u5_mult_79_SUMB_18__9_), .CO(
        u5_mult_79_CARRYB_19__8_), .S(u5_mult_79_SUMB_19__8_) );
  FA_X1 u5_mult_79_S2_19_7 ( .A(u5_mult_79_ab_19__7_), .B(
        u5_mult_79_CARRYB_18__7_), .CI(u5_mult_79_SUMB_18__8_), .CO(
        u5_mult_79_CARRYB_19__7_), .S(u5_mult_79_SUMB_19__7_) );
  FA_X1 u5_mult_79_S2_19_6 ( .A(u5_mult_79_ab_19__6_), .B(
        u5_mult_79_CARRYB_18__6_), .CI(u5_mult_79_SUMB_18__7_), .CO(
        u5_mult_79_CARRYB_19__6_), .S(u5_mult_79_SUMB_19__6_) );
  FA_X1 u5_mult_79_S2_19_5 ( .A(u5_mult_79_ab_19__5_), .B(
        u5_mult_79_CARRYB_18__5_), .CI(u5_mult_79_SUMB_18__6_), .CO(
        u5_mult_79_CARRYB_19__5_), .S(u5_mult_79_SUMB_19__5_) );
  FA_X1 u5_mult_79_S2_19_4 ( .A(u5_mult_79_ab_19__4_), .B(
        u5_mult_79_CARRYB_18__4_), .CI(u5_mult_79_SUMB_18__5_), .CO(
        u5_mult_79_CARRYB_19__4_), .S(u5_mult_79_SUMB_19__4_) );
  FA_X1 u5_mult_79_S2_19_3 ( .A(u5_mult_79_ab_19__3_), .B(
        u5_mult_79_CARRYB_18__3_), .CI(u5_mult_79_SUMB_18__4_), .CO(
        u5_mult_79_CARRYB_19__3_), .S(u5_mult_79_SUMB_19__3_) );
  FA_X1 u5_mult_79_S2_19_2 ( .A(u5_mult_79_ab_19__2_), .B(
        u5_mult_79_CARRYB_18__2_), .CI(u5_mult_79_SUMB_18__3_), .CO(
        u5_mult_79_CARRYB_19__2_), .S(u5_mult_79_SUMB_19__2_) );
  FA_X1 u5_mult_79_S2_19_1 ( .A(u5_mult_79_ab_19__1_), .B(
        u5_mult_79_CARRYB_18__1_), .CI(u5_mult_79_SUMB_18__2_), .CO(
        u5_mult_79_CARRYB_19__1_), .S(u5_mult_79_SUMB_19__1_) );
  FA_X1 u5_mult_79_S1_19_0 ( .A(u5_mult_79_ab_19__0_), .B(
        u5_mult_79_CARRYB_18__0_), .CI(u5_mult_79_SUMB_18__1_), .CO(
        u5_mult_79_CARRYB_19__0_), .S(u5_N19) );
  FA_X1 u5_mult_79_S3_20_22 ( .A(u5_mult_79_ab_20__22_), .B(
        u5_mult_79_CARRYB_19__22_), .CI(u5_mult_79_ab_19__23_), .CO(
        u5_mult_79_CARRYB_20__22_), .S(u5_mult_79_SUMB_20__22_) );
  FA_X1 u5_mult_79_S2_20_21 ( .A(u5_mult_79_ab_20__21_), .B(
        u5_mult_79_CARRYB_19__21_), .CI(u5_mult_79_SUMB_19__22_), .CO(
        u5_mult_79_CARRYB_20__21_), .S(u5_mult_79_SUMB_20__21_) );
  FA_X1 u5_mult_79_S2_20_20 ( .A(u5_mult_79_ab_20__20_), .B(
        u5_mult_79_CARRYB_19__20_), .CI(u5_mult_79_SUMB_19__21_), .CO(
        u5_mult_79_CARRYB_20__20_), .S(u5_mult_79_SUMB_20__20_) );
  FA_X1 u5_mult_79_S2_20_19 ( .A(u5_mult_79_ab_20__19_), .B(
        u5_mult_79_CARRYB_19__19_), .CI(u5_mult_79_SUMB_19__20_), .CO(
        u5_mult_79_CARRYB_20__19_), .S(u5_mult_79_SUMB_20__19_) );
  FA_X1 u5_mult_79_S2_20_18 ( .A(u5_mult_79_ab_20__18_), .B(
        u5_mult_79_CARRYB_19__18_), .CI(u5_mult_79_SUMB_19__19_), .CO(
        u5_mult_79_CARRYB_20__18_), .S(u5_mult_79_SUMB_20__18_) );
  FA_X1 u5_mult_79_S2_20_17 ( .A(u5_mult_79_ab_20__17_), .B(
        u5_mult_79_CARRYB_19__17_), .CI(u5_mult_79_SUMB_19__18_), .CO(
        u5_mult_79_CARRYB_20__17_), .S(u5_mult_79_SUMB_20__17_) );
  FA_X1 u5_mult_79_S2_20_16 ( .A(u5_mult_79_ab_20__16_), .B(
        u5_mult_79_CARRYB_19__16_), .CI(u5_mult_79_SUMB_19__17_), .CO(
        u5_mult_79_CARRYB_20__16_), .S(u5_mult_79_SUMB_20__16_) );
  FA_X1 u5_mult_79_S2_20_15 ( .A(u5_mult_79_ab_20__15_), .B(
        u5_mult_79_CARRYB_19__15_), .CI(u5_mult_79_SUMB_19__16_), .CO(
        u5_mult_79_CARRYB_20__15_), .S(u5_mult_79_SUMB_20__15_) );
  FA_X1 u5_mult_79_S2_20_14 ( .A(u5_mult_79_ab_20__14_), .B(
        u5_mult_79_CARRYB_19__14_), .CI(u5_mult_79_SUMB_19__15_), .CO(
        u5_mult_79_CARRYB_20__14_), .S(u5_mult_79_SUMB_20__14_) );
  FA_X1 u5_mult_79_S2_20_13 ( .A(u5_mult_79_ab_20__13_), .B(
        u5_mult_79_CARRYB_19__13_), .CI(u5_mult_79_SUMB_19__14_), .CO(
        u5_mult_79_CARRYB_20__13_), .S(u5_mult_79_SUMB_20__13_) );
  FA_X1 u5_mult_79_S2_20_12 ( .A(u5_mult_79_ab_20__12_), .B(
        u5_mult_79_CARRYB_19__12_), .CI(u5_mult_79_SUMB_19__13_), .CO(
        u5_mult_79_CARRYB_20__12_), .S(u5_mult_79_SUMB_20__12_) );
  FA_X1 u5_mult_79_S2_20_11 ( .A(u5_mult_79_ab_20__11_), .B(
        u5_mult_79_CARRYB_19__11_), .CI(u5_mult_79_SUMB_19__12_), .CO(
        u5_mult_79_CARRYB_20__11_), .S(u5_mult_79_SUMB_20__11_) );
  FA_X1 u5_mult_79_S2_20_10 ( .A(u5_mult_79_ab_20__10_), .B(
        u5_mult_79_CARRYB_19__10_), .CI(u5_mult_79_SUMB_19__11_), .CO(
        u5_mult_79_CARRYB_20__10_), .S(u5_mult_79_SUMB_20__10_) );
  FA_X1 u5_mult_79_S2_20_9 ( .A(u5_mult_79_ab_20__9_), .B(
        u5_mult_79_CARRYB_19__9_), .CI(u5_mult_79_SUMB_19__10_), .CO(
        u5_mult_79_CARRYB_20__9_), .S(u5_mult_79_SUMB_20__9_) );
  FA_X1 u5_mult_79_S2_20_8 ( .A(u5_mult_79_ab_20__8_), .B(
        u5_mult_79_CARRYB_19__8_), .CI(u5_mult_79_SUMB_19__9_), .CO(
        u5_mult_79_CARRYB_20__8_), .S(u5_mult_79_SUMB_20__8_) );
  FA_X1 u5_mult_79_S2_20_7 ( .A(u5_mult_79_ab_20__7_), .B(
        u5_mult_79_CARRYB_19__7_), .CI(u5_mult_79_SUMB_19__8_), .CO(
        u5_mult_79_CARRYB_20__7_), .S(u5_mult_79_SUMB_20__7_) );
  FA_X1 u5_mult_79_S2_20_6 ( .A(u5_mult_79_ab_20__6_), .B(
        u5_mult_79_CARRYB_19__6_), .CI(u5_mult_79_SUMB_19__7_), .CO(
        u5_mult_79_CARRYB_20__6_), .S(u5_mult_79_SUMB_20__6_) );
  FA_X1 u5_mult_79_S2_20_5 ( .A(u5_mult_79_ab_20__5_), .B(
        u5_mult_79_CARRYB_19__5_), .CI(u5_mult_79_SUMB_19__6_), .CO(
        u5_mult_79_CARRYB_20__5_), .S(u5_mult_79_SUMB_20__5_) );
  FA_X1 u5_mult_79_S2_20_4 ( .A(u5_mult_79_ab_20__4_), .B(
        u5_mult_79_CARRYB_19__4_), .CI(u5_mult_79_SUMB_19__5_), .CO(
        u5_mult_79_CARRYB_20__4_), .S(u5_mult_79_SUMB_20__4_) );
  FA_X1 u5_mult_79_S2_20_3 ( .A(u5_mult_79_ab_20__3_), .B(
        u5_mult_79_CARRYB_19__3_), .CI(u5_mult_79_SUMB_19__4_), .CO(
        u5_mult_79_CARRYB_20__3_), .S(u5_mult_79_SUMB_20__3_) );
  FA_X1 u5_mult_79_S2_20_2 ( .A(u5_mult_79_ab_20__2_), .B(
        u5_mult_79_CARRYB_19__2_), .CI(u5_mult_79_SUMB_19__3_), .CO(
        u5_mult_79_CARRYB_20__2_), .S(u5_mult_79_SUMB_20__2_) );
  FA_X1 u5_mult_79_S2_20_1 ( .A(u5_mult_79_ab_20__1_), .B(
        u5_mult_79_CARRYB_19__1_), .CI(u5_mult_79_SUMB_19__2_), .CO(
        u5_mult_79_CARRYB_20__1_), .S(u5_mult_79_SUMB_20__1_) );
  FA_X1 u5_mult_79_S1_20_0 ( .A(u5_mult_79_ab_20__0_), .B(
        u5_mult_79_CARRYB_19__0_), .CI(u5_mult_79_SUMB_19__1_), .CO(
        u5_mult_79_CARRYB_20__0_), .S(u5_N20) );
  FA_X1 u5_mult_79_S3_21_22 ( .A(u5_mult_79_ab_21__22_), .B(
        u5_mult_79_CARRYB_20__22_), .CI(u5_mult_79_ab_20__23_), .CO(
        u5_mult_79_CARRYB_21__22_), .S(u5_mult_79_SUMB_21__22_) );
  FA_X1 u5_mult_79_S2_21_21 ( .A(u5_mult_79_ab_21__21_), .B(
        u5_mult_79_CARRYB_20__21_), .CI(u5_mult_79_SUMB_20__22_), .CO(
        u5_mult_79_CARRYB_21__21_), .S(u5_mult_79_SUMB_21__21_) );
  FA_X1 u5_mult_79_S2_21_20 ( .A(u5_mult_79_ab_21__20_), .B(
        u5_mult_79_CARRYB_20__20_), .CI(u5_mult_79_SUMB_20__21_), .CO(
        u5_mult_79_CARRYB_21__20_), .S(u5_mult_79_SUMB_21__20_) );
  FA_X1 u5_mult_79_S2_21_19 ( .A(u5_mult_79_ab_21__19_), .B(
        u5_mult_79_CARRYB_20__19_), .CI(u5_mult_79_SUMB_20__20_), .CO(
        u5_mult_79_CARRYB_21__19_), .S(u5_mult_79_SUMB_21__19_) );
  FA_X1 u5_mult_79_S2_21_18 ( .A(u5_mult_79_ab_21__18_), .B(
        u5_mult_79_CARRYB_20__18_), .CI(u5_mult_79_SUMB_20__19_), .CO(
        u5_mult_79_CARRYB_21__18_), .S(u5_mult_79_SUMB_21__18_) );
  FA_X1 u5_mult_79_S2_21_17 ( .A(u5_mult_79_ab_21__17_), .B(
        u5_mult_79_CARRYB_20__17_), .CI(u5_mult_79_SUMB_20__18_), .CO(
        u5_mult_79_CARRYB_21__17_), .S(u5_mult_79_SUMB_21__17_) );
  FA_X1 u5_mult_79_S2_21_16 ( .A(u5_mult_79_ab_21__16_), .B(
        u5_mult_79_CARRYB_20__16_), .CI(u5_mult_79_SUMB_20__17_), .CO(
        u5_mult_79_CARRYB_21__16_), .S(u5_mult_79_SUMB_21__16_) );
  FA_X1 u5_mult_79_S2_21_15 ( .A(u5_mult_79_ab_21__15_), .B(
        u5_mult_79_CARRYB_20__15_), .CI(u5_mult_79_SUMB_20__16_), .CO(
        u5_mult_79_CARRYB_21__15_), .S(u5_mult_79_SUMB_21__15_) );
  FA_X1 u5_mult_79_S2_21_14 ( .A(u5_mult_79_ab_21__14_), .B(
        u5_mult_79_CARRYB_20__14_), .CI(u5_mult_79_SUMB_20__15_), .CO(
        u5_mult_79_CARRYB_21__14_), .S(u5_mult_79_SUMB_21__14_) );
  FA_X1 u5_mult_79_S2_21_13 ( .A(u5_mult_79_ab_21__13_), .B(
        u5_mult_79_CARRYB_20__13_), .CI(u5_mult_79_SUMB_20__14_), .CO(
        u5_mult_79_CARRYB_21__13_), .S(u5_mult_79_SUMB_21__13_) );
  FA_X1 u5_mult_79_S2_21_12 ( .A(u5_mult_79_ab_21__12_), .B(
        u5_mult_79_CARRYB_20__12_), .CI(u5_mult_79_SUMB_20__13_), .CO(
        u5_mult_79_CARRYB_21__12_), .S(u5_mult_79_SUMB_21__12_) );
  FA_X1 u5_mult_79_S2_21_11 ( .A(u5_mult_79_ab_21__11_), .B(
        u5_mult_79_CARRYB_20__11_), .CI(u5_mult_79_SUMB_20__12_), .CO(
        u5_mult_79_CARRYB_21__11_), .S(u5_mult_79_SUMB_21__11_) );
  FA_X1 u5_mult_79_S2_21_10 ( .A(u5_mult_79_ab_21__10_), .B(
        u5_mult_79_CARRYB_20__10_), .CI(u5_mult_79_SUMB_20__11_), .CO(
        u5_mult_79_CARRYB_21__10_), .S(u5_mult_79_SUMB_21__10_) );
  FA_X1 u5_mult_79_S2_21_9 ( .A(u5_mult_79_ab_21__9_), .B(
        u5_mult_79_CARRYB_20__9_), .CI(u5_mult_79_SUMB_20__10_), .CO(
        u5_mult_79_CARRYB_21__9_), .S(u5_mult_79_SUMB_21__9_) );
  FA_X1 u5_mult_79_S2_21_8 ( .A(u5_mult_79_ab_21__8_), .B(
        u5_mult_79_CARRYB_20__8_), .CI(u5_mult_79_SUMB_20__9_), .CO(
        u5_mult_79_CARRYB_21__8_), .S(u5_mult_79_SUMB_21__8_) );
  FA_X1 u5_mult_79_S2_21_7 ( .A(u5_mult_79_ab_21__7_), .B(
        u5_mult_79_CARRYB_20__7_), .CI(u5_mult_79_SUMB_20__8_), .CO(
        u5_mult_79_CARRYB_21__7_), .S(u5_mult_79_SUMB_21__7_) );
  FA_X1 u5_mult_79_S2_21_6 ( .A(u5_mult_79_ab_21__6_), .B(
        u5_mult_79_CARRYB_20__6_), .CI(u5_mult_79_SUMB_20__7_), .CO(
        u5_mult_79_CARRYB_21__6_), .S(u5_mult_79_SUMB_21__6_) );
  FA_X1 u5_mult_79_S2_21_5 ( .A(u5_mult_79_ab_21__5_), .B(
        u5_mult_79_CARRYB_20__5_), .CI(u5_mult_79_SUMB_20__6_), .CO(
        u5_mult_79_CARRYB_21__5_), .S(u5_mult_79_SUMB_21__5_) );
  FA_X1 u5_mult_79_S2_21_4 ( .A(u5_mult_79_ab_21__4_), .B(
        u5_mult_79_CARRYB_20__4_), .CI(u5_mult_79_SUMB_20__5_), .CO(
        u5_mult_79_CARRYB_21__4_), .S(u5_mult_79_SUMB_21__4_) );
  FA_X1 u5_mult_79_S2_21_3 ( .A(u5_mult_79_ab_21__3_), .B(
        u5_mult_79_CARRYB_20__3_), .CI(u5_mult_79_SUMB_20__4_), .CO(
        u5_mult_79_CARRYB_21__3_), .S(u5_mult_79_SUMB_21__3_) );
  FA_X1 u5_mult_79_S2_21_2 ( .A(u5_mult_79_ab_21__2_), .B(
        u5_mult_79_CARRYB_20__2_), .CI(u5_mult_79_SUMB_20__3_), .CO(
        u5_mult_79_CARRYB_21__2_), .S(u5_mult_79_SUMB_21__2_) );
  FA_X1 u5_mult_79_S2_21_1 ( .A(u5_mult_79_ab_21__1_), .B(
        u5_mult_79_CARRYB_20__1_), .CI(u5_mult_79_SUMB_20__2_), .CO(
        u5_mult_79_CARRYB_21__1_), .S(u5_mult_79_SUMB_21__1_) );
  FA_X1 u5_mult_79_S1_21_0 ( .A(u5_mult_79_ab_21__0_), .B(
        u5_mult_79_CARRYB_20__0_), .CI(u5_mult_79_SUMB_20__1_), .CO(
        u5_mult_79_CARRYB_21__0_), .S(u5_N21) );
  FA_X1 u5_mult_79_S3_22_22 ( .A(u5_mult_79_ab_22__22_), .B(
        u5_mult_79_CARRYB_21__22_), .CI(u5_mult_79_ab_21__23_), .CO(
        u5_mult_79_CARRYB_22__22_), .S(u5_mult_79_SUMB_22__22_) );
  FA_X1 u5_mult_79_S2_22_21 ( .A(u5_mult_79_ab_22__21_), .B(
        u5_mult_79_CARRYB_21__21_), .CI(u5_mult_79_SUMB_21__22_), .CO(
        u5_mult_79_CARRYB_22__21_), .S(u5_mult_79_SUMB_22__21_) );
  FA_X1 u5_mult_79_S2_22_20 ( .A(u5_mult_79_ab_22__20_), .B(
        u5_mult_79_CARRYB_21__20_), .CI(u5_mult_79_SUMB_21__21_), .CO(
        u5_mult_79_CARRYB_22__20_), .S(u5_mult_79_SUMB_22__20_) );
  FA_X1 u5_mult_79_S2_22_19 ( .A(u5_mult_79_ab_22__19_), .B(
        u5_mult_79_CARRYB_21__19_), .CI(u5_mult_79_SUMB_21__20_), .CO(
        u5_mult_79_CARRYB_22__19_), .S(u5_mult_79_SUMB_22__19_) );
  FA_X1 u5_mult_79_S2_22_18 ( .A(u5_mult_79_ab_22__18_), .B(
        u5_mult_79_CARRYB_21__18_), .CI(u5_mult_79_SUMB_21__19_), .CO(
        u5_mult_79_CARRYB_22__18_), .S(u5_mult_79_SUMB_22__18_) );
  FA_X1 u5_mult_79_S2_22_17 ( .A(u5_mult_79_ab_22__17_), .B(
        u5_mult_79_CARRYB_21__17_), .CI(u5_mult_79_SUMB_21__18_), .CO(
        u5_mult_79_CARRYB_22__17_), .S(u5_mult_79_SUMB_22__17_) );
  FA_X1 u5_mult_79_S2_22_16 ( .A(u5_mult_79_ab_22__16_), .B(
        u5_mult_79_CARRYB_21__16_), .CI(u5_mult_79_SUMB_21__17_), .CO(
        u5_mult_79_CARRYB_22__16_), .S(u5_mult_79_SUMB_22__16_) );
  FA_X1 u5_mult_79_S2_22_15 ( .A(u5_mult_79_ab_22__15_), .B(
        u5_mult_79_CARRYB_21__15_), .CI(u5_mult_79_SUMB_21__16_), .CO(
        u5_mult_79_CARRYB_22__15_), .S(u5_mult_79_SUMB_22__15_) );
  FA_X1 u5_mult_79_S2_22_14 ( .A(u5_mult_79_ab_22__14_), .B(
        u5_mult_79_CARRYB_21__14_), .CI(u5_mult_79_SUMB_21__15_), .CO(
        u5_mult_79_CARRYB_22__14_), .S(u5_mult_79_SUMB_22__14_) );
  FA_X1 u5_mult_79_S2_22_13 ( .A(u5_mult_79_ab_22__13_), .B(
        u5_mult_79_CARRYB_21__13_), .CI(u5_mult_79_SUMB_21__14_), .CO(
        u5_mult_79_CARRYB_22__13_), .S(u5_mult_79_SUMB_22__13_) );
  FA_X1 u5_mult_79_S2_22_12 ( .A(u5_mult_79_ab_22__12_), .B(
        u5_mult_79_CARRYB_21__12_), .CI(u5_mult_79_SUMB_21__13_), .CO(
        u5_mult_79_CARRYB_22__12_), .S(u5_mult_79_SUMB_22__12_) );
  FA_X1 u5_mult_79_S2_22_11 ( .A(u5_mult_79_ab_22__11_), .B(
        u5_mult_79_CARRYB_21__11_), .CI(u5_mult_79_SUMB_21__12_), .CO(
        u5_mult_79_CARRYB_22__11_), .S(u5_mult_79_SUMB_22__11_) );
  FA_X1 u5_mult_79_S2_22_10 ( .A(u5_mult_79_ab_22__10_), .B(
        u5_mult_79_CARRYB_21__10_), .CI(u5_mult_79_SUMB_21__11_), .CO(
        u5_mult_79_CARRYB_22__10_), .S(u5_mult_79_SUMB_22__10_) );
  FA_X1 u5_mult_79_S2_22_9 ( .A(u5_mult_79_ab_22__9_), .B(
        u5_mult_79_CARRYB_21__9_), .CI(u5_mult_79_SUMB_21__10_), .CO(
        u5_mult_79_CARRYB_22__9_), .S(u5_mult_79_SUMB_22__9_) );
  FA_X1 u5_mult_79_S2_22_8 ( .A(u5_mult_79_ab_22__8_), .B(
        u5_mult_79_CARRYB_21__8_), .CI(u5_mult_79_SUMB_21__9_), .CO(
        u5_mult_79_CARRYB_22__8_), .S(u5_mult_79_SUMB_22__8_) );
  FA_X1 u5_mult_79_S2_22_7 ( .A(u5_mult_79_ab_22__7_), .B(
        u5_mult_79_CARRYB_21__7_), .CI(u5_mult_79_SUMB_21__8_), .CO(
        u5_mult_79_CARRYB_22__7_), .S(u5_mult_79_SUMB_22__7_) );
  FA_X1 u5_mult_79_S2_22_6 ( .A(u5_mult_79_ab_22__6_), .B(
        u5_mult_79_CARRYB_21__6_), .CI(u5_mult_79_SUMB_21__7_), .CO(
        u5_mult_79_CARRYB_22__6_), .S(u5_mult_79_SUMB_22__6_) );
  FA_X1 u5_mult_79_S2_22_5 ( .A(u5_mult_79_ab_22__5_), .B(
        u5_mult_79_CARRYB_21__5_), .CI(u5_mult_79_SUMB_21__6_), .CO(
        u5_mult_79_CARRYB_22__5_), .S(u5_mult_79_SUMB_22__5_) );
  FA_X1 u5_mult_79_S2_22_4 ( .A(u5_mult_79_ab_22__4_), .B(
        u5_mult_79_CARRYB_21__4_), .CI(u5_mult_79_SUMB_21__5_), .CO(
        u5_mult_79_CARRYB_22__4_), .S(u5_mult_79_SUMB_22__4_) );
  FA_X1 u5_mult_79_S2_22_3 ( .A(u5_mult_79_ab_22__3_), .B(
        u5_mult_79_CARRYB_21__3_), .CI(u5_mult_79_SUMB_21__4_), .CO(
        u5_mult_79_CARRYB_22__3_), .S(u5_mult_79_SUMB_22__3_) );
  FA_X1 u5_mult_79_S2_22_2 ( .A(u5_mult_79_ab_22__2_), .B(
        u5_mult_79_CARRYB_21__2_), .CI(u5_mult_79_SUMB_21__3_), .CO(
        u5_mult_79_CARRYB_22__2_), .S(u5_mult_79_SUMB_22__2_) );
  FA_X1 u5_mult_79_S2_22_1 ( .A(u5_mult_79_ab_22__1_), .B(
        u5_mult_79_CARRYB_21__1_), .CI(u5_mult_79_SUMB_21__2_), .CO(
        u5_mult_79_CARRYB_22__1_), .S(u5_mult_79_SUMB_22__1_) );
  FA_X1 u5_mult_79_S1_22_0 ( .A(u5_mult_79_ab_22__0_), .B(
        u5_mult_79_CARRYB_21__0_), .CI(u5_mult_79_SUMB_21__1_), .CO(
        u5_mult_79_CARRYB_22__0_), .S(u5_N22) );
  FA_X1 u5_mult_79_S5_22 ( .A(u5_mult_79_ab_23__22_), .B(
        u5_mult_79_CARRYB_22__22_), .CI(u5_mult_79_ab_22__23_), .CO(
        u5_mult_79_CARRYB_23__22_), .S(u5_mult_79_SUMB_23__22_) );
  FA_X1 u5_mult_79_S4_21 ( .A(u5_mult_79_ab_23__21_), .B(
        u5_mult_79_CARRYB_22__21_), .CI(u5_mult_79_SUMB_22__22_), .CO(
        u5_mult_79_CARRYB_23__21_), .S(u5_mult_79_SUMB_23__21_) );
  FA_X1 u5_mult_79_S4_20 ( .A(u5_mult_79_ab_23__20_), .B(
        u5_mult_79_CARRYB_22__20_), .CI(u5_mult_79_SUMB_22__21_), .CO(
        u5_mult_79_CARRYB_23__20_), .S(u5_mult_79_SUMB_23__20_) );
  FA_X1 u5_mult_79_S4_19 ( .A(u5_mult_79_ab_23__19_), .B(
        u5_mult_79_CARRYB_22__19_), .CI(u5_mult_79_SUMB_22__20_), .CO(
        u5_mult_79_CARRYB_23__19_), .S(u5_mult_79_SUMB_23__19_) );
  FA_X1 u5_mult_79_S4_18 ( .A(u5_mult_79_ab_23__18_), .B(
        u5_mult_79_CARRYB_22__18_), .CI(u5_mult_79_SUMB_22__19_), .CO(
        u5_mult_79_CARRYB_23__18_), .S(u5_mult_79_SUMB_23__18_) );
  FA_X1 u5_mult_79_S4_17 ( .A(u5_mult_79_ab_23__17_), .B(
        u5_mult_79_CARRYB_22__17_), .CI(u5_mult_79_SUMB_22__18_), .CO(
        u5_mult_79_CARRYB_23__17_), .S(u5_mult_79_SUMB_23__17_) );
  FA_X1 u5_mult_79_S4_16 ( .A(u5_mult_79_ab_23__16_), .B(
        u5_mult_79_CARRYB_22__16_), .CI(u5_mult_79_SUMB_22__17_), .CO(
        u5_mult_79_CARRYB_23__16_), .S(u5_mult_79_SUMB_23__16_) );
  FA_X1 u5_mult_79_S4_15 ( .A(u5_mult_79_ab_23__15_), .B(
        u5_mult_79_CARRYB_22__15_), .CI(u5_mult_79_SUMB_22__16_), .CO(
        u5_mult_79_CARRYB_23__15_), .S(u5_mult_79_SUMB_23__15_) );
  FA_X1 u5_mult_79_S4_14 ( .A(u5_mult_79_ab_23__14_), .B(
        u5_mult_79_CARRYB_22__14_), .CI(u5_mult_79_SUMB_22__15_), .CO(
        u5_mult_79_CARRYB_23__14_), .S(u5_mult_79_SUMB_23__14_) );
  FA_X1 u5_mult_79_S4_13 ( .A(u5_mult_79_ab_23__13_), .B(
        u5_mult_79_CARRYB_22__13_), .CI(u5_mult_79_SUMB_22__14_), .CO(
        u5_mult_79_CARRYB_23__13_), .S(u5_mult_79_SUMB_23__13_) );
  FA_X1 u5_mult_79_S4_12 ( .A(u5_mult_79_ab_23__12_), .B(
        u5_mult_79_CARRYB_22__12_), .CI(u5_mult_79_SUMB_22__13_), .CO(
        u5_mult_79_CARRYB_23__12_), .S(u5_mult_79_SUMB_23__12_) );
  FA_X1 u5_mult_79_S4_11 ( .A(u5_mult_79_ab_23__11_), .B(
        u5_mult_79_CARRYB_22__11_), .CI(u5_mult_79_SUMB_22__12_), .CO(
        u5_mult_79_CARRYB_23__11_), .S(u5_mult_79_SUMB_23__11_) );
  FA_X1 u5_mult_79_S4_10 ( .A(u5_mult_79_ab_23__10_), .B(
        u5_mult_79_CARRYB_22__10_), .CI(u5_mult_79_SUMB_22__11_), .CO(
        u5_mult_79_CARRYB_23__10_), .S(u5_mult_79_SUMB_23__10_) );
  FA_X1 u5_mult_79_S4_9 ( .A(u5_mult_79_ab_23__9_), .B(
        u5_mult_79_CARRYB_22__9_), .CI(u5_mult_79_SUMB_22__10_), .CO(
        u5_mult_79_CARRYB_23__9_), .S(u5_mult_79_SUMB_23__9_) );
  FA_X1 u5_mult_79_S4_8 ( .A(u5_mult_79_ab_23__8_), .B(
        u5_mult_79_CARRYB_22__8_), .CI(u5_mult_79_SUMB_22__9_), .CO(
        u5_mult_79_CARRYB_23__8_), .S(u5_mult_79_SUMB_23__8_) );
  FA_X1 u5_mult_79_S4_7 ( .A(u5_mult_79_ab_23__7_), .B(
        u5_mult_79_CARRYB_22__7_), .CI(u5_mult_79_SUMB_22__8_), .CO(
        u5_mult_79_CARRYB_23__7_), .S(u5_mult_79_SUMB_23__7_) );
  FA_X1 u5_mult_79_S4_6 ( .A(u5_mult_79_ab_23__6_), .B(
        u5_mult_79_CARRYB_22__6_), .CI(u5_mult_79_SUMB_22__7_), .CO(
        u5_mult_79_CARRYB_23__6_), .S(u5_mult_79_SUMB_23__6_) );
  FA_X1 u5_mult_79_S4_5 ( .A(u5_mult_79_ab_23__5_), .B(
        u5_mult_79_CARRYB_22__5_), .CI(u5_mult_79_SUMB_22__6_), .CO(
        u5_mult_79_CARRYB_23__5_), .S(u5_mult_79_SUMB_23__5_) );
  FA_X1 u5_mult_79_S4_4 ( .A(u5_mult_79_ab_23__4_), .B(
        u5_mult_79_CARRYB_22__4_), .CI(u5_mult_79_SUMB_22__5_), .CO(
        u5_mult_79_CARRYB_23__4_), .S(u5_mult_79_SUMB_23__4_) );
  FA_X1 u5_mult_79_S4_3 ( .A(u5_mult_79_ab_23__3_), .B(
        u5_mult_79_CARRYB_22__3_), .CI(u5_mult_79_SUMB_22__4_), .CO(
        u5_mult_79_CARRYB_23__3_), .S(u5_mult_79_SUMB_23__3_) );
  FA_X1 u5_mult_79_S4_2 ( .A(u5_mult_79_ab_23__2_), .B(
        u5_mult_79_CARRYB_22__2_), .CI(u5_mult_79_SUMB_22__3_), .CO(
        u5_mult_79_CARRYB_23__2_), .S(u5_mult_79_SUMB_23__2_) );
  FA_X1 u5_mult_79_S4_1 ( .A(u5_mult_79_ab_23__1_), .B(
        u5_mult_79_CARRYB_22__1_), .CI(u5_mult_79_SUMB_22__2_), .CO(
        u5_mult_79_CARRYB_23__1_), .S(u5_mult_79_SUMB_23__1_) );
  FA_X1 u5_mult_79_S4_0 ( .A(u5_mult_79_ab_23__0_), .B(
        u5_mult_79_CARRYB_22__0_), .CI(u5_mult_79_SUMB_22__1_), .CO(
        u5_mult_79_CARRYB_23__0_), .S(u5_N23) );
  NAND2_X1 u5_mult_79_FS_1_U133 ( .A1(u5_mult_79_n79), .A2(u5_mult_79_n30), 
        .ZN(u5_mult_79_FS_1_n110) );
  AND2_X1 u5_mult_79_FS_1_U132 ( .A1(u5_mult_79_n74), .A2(u5_mult_79_n29), 
        .ZN(u5_mult_79_FS_1_n107) );
  NOR2_X1 u5_mult_79_FS_1_U131 ( .A1(u5_mult_79_n74), .A2(u5_mult_79_n29), 
        .ZN(u5_mult_79_FS_1_n108) );
  NOR2_X1 u5_mult_79_FS_1_U130 ( .A1(u5_mult_79_FS_1_n107), .A2(
        u5_mult_79_FS_1_n108), .ZN(u5_mult_79_FS_1_n109) );
  XOR2_X1 u5_mult_79_FS_1_U129 ( .A(u5_mult_79_FS_1_n25), .B(
        u5_mult_79_FS_1_n109), .Z(u5_N26) );
  NOR2_X1 u5_mult_79_FS_1_U128 ( .A1(u5_mult_79_n78), .A2(u5_mult_79_n35), 
        .ZN(u5_mult_79_FS_1_n103) );
  NAND2_X1 u5_mult_79_FS_1_U127 ( .A1(u5_mult_79_n78), .A2(u5_mult_79_n35), 
        .ZN(u5_mult_79_FS_1_n105) );
  NAND2_X1 u5_mult_79_FS_1_U126 ( .A1(u5_mult_79_FS_1_n23), .A2(
        u5_mult_79_FS_1_n105), .ZN(u5_mult_79_FS_1_n106) );
  AOI21_X1 u5_mult_79_FS_1_U125 ( .B1(u5_mult_79_FS_1_n24), .B2(
        u5_mult_79_FS_1_n25), .A(u5_mult_79_FS_1_n107), .ZN(
        u5_mult_79_FS_1_n104) );
  XOR2_X1 u5_mult_79_FS_1_U124 ( .A(u5_mult_79_FS_1_n106), .B(
        u5_mult_79_FS_1_n104), .Z(u5_N27) );
  OAI21_X1 u5_mult_79_FS_1_U123 ( .B1(u5_mult_79_FS_1_n103), .B2(
        u5_mult_79_FS_1_n104), .A(u5_mult_79_FS_1_n105), .ZN(
        u5_mult_79_FS_1_n99) );
  AND2_X1 u5_mult_79_FS_1_U122 ( .A1(u5_mult_79_n73), .A2(u5_mult_79_n28), 
        .ZN(u5_mult_79_FS_1_n100) );
  NOR2_X1 u5_mult_79_FS_1_U121 ( .A1(u5_mult_79_n73), .A2(u5_mult_79_n28), 
        .ZN(u5_mult_79_FS_1_n101) );
  NOR2_X1 u5_mult_79_FS_1_U120 ( .A1(u5_mult_79_FS_1_n100), .A2(
        u5_mult_79_FS_1_n101), .ZN(u5_mult_79_FS_1_n102) );
  XOR2_X1 u5_mult_79_FS_1_U119 ( .A(u5_mult_79_FS_1_n99), .B(
        u5_mult_79_FS_1_n102), .Z(u5_N28) );
  NOR2_X1 u5_mult_79_FS_1_U118 ( .A1(u5_mult_79_n77), .A2(u5_mult_79_n34), 
        .ZN(u5_mult_79_FS_1_n95) );
  NAND2_X1 u5_mult_79_FS_1_U117 ( .A1(u5_mult_79_n77), .A2(u5_mult_79_n34), 
        .ZN(u5_mult_79_FS_1_n97) );
  NAND2_X1 u5_mult_79_FS_1_U116 ( .A1(u5_mult_79_FS_1_n21), .A2(
        u5_mult_79_FS_1_n97), .ZN(u5_mult_79_FS_1_n98) );
  AOI21_X1 u5_mult_79_FS_1_U115 ( .B1(u5_mult_79_FS_1_n99), .B2(
        u5_mult_79_FS_1_n22), .A(u5_mult_79_FS_1_n100), .ZN(
        u5_mult_79_FS_1_n96) );
  XOR2_X1 u5_mult_79_FS_1_U114 ( .A(u5_mult_79_FS_1_n98), .B(
        u5_mult_79_FS_1_n96), .Z(u5_N29) );
  OAI21_X1 u5_mult_79_FS_1_U113 ( .B1(u5_mult_79_FS_1_n95), .B2(
        u5_mult_79_FS_1_n96), .A(u5_mult_79_FS_1_n97), .ZN(u5_mult_79_FS_1_n91) );
  AND2_X1 u5_mult_79_FS_1_U112 ( .A1(u5_mult_79_n72), .A2(u5_mult_79_n27), 
        .ZN(u5_mult_79_FS_1_n92) );
  NOR2_X1 u5_mult_79_FS_1_U111 ( .A1(u5_mult_79_n72), .A2(u5_mult_79_n27), 
        .ZN(u5_mult_79_FS_1_n93) );
  NOR2_X1 u5_mult_79_FS_1_U110 ( .A1(u5_mult_79_FS_1_n92), .A2(
        u5_mult_79_FS_1_n93), .ZN(u5_mult_79_FS_1_n94) );
  XOR2_X1 u5_mult_79_FS_1_U109 ( .A(u5_mult_79_FS_1_n91), .B(
        u5_mult_79_FS_1_n94), .Z(u5_N30) );
  NOR2_X1 u5_mult_79_FS_1_U108 ( .A1(u5_mult_79_n76), .A2(u5_mult_79_n33), 
        .ZN(u5_mult_79_FS_1_n87) );
  NAND2_X1 u5_mult_79_FS_1_U107 ( .A1(u5_mult_79_n76), .A2(u5_mult_79_n33), 
        .ZN(u5_mult_79_FS_1_n89) );
  NAND2_X1 u5_mult_79_FS_1_U106 ( .A1(u5_mult_79_FS_1_n19), .A2(
        u5_mult_79_FS_1_n89), .ZN(u5_mult_79_FS_1_n90) );
  AOI21_X1 u5_mult_79_FS_1_U105 ( .B1(u5_mult_79_FS_1_n20), .B2(
        u5_mult_79_FS_1_n91), .A(u5_mult_79_FS_1_n92), .ZN(u5_mult_79_FS_1_n88) );
  XOR2_X1 u5_mult_79_FS_1_U104 ( .A(u5_mult_79_FS_1_n90), .B(
        u5_mult_79_FS_1_n88), .Z(u5_N31) );
  OAI21_X1 u5_mult_79_FS_1_U103 ( .B1(u5_mult_79_FS_1_n87), .B2(
        u5_mult_79_FS_1_n88), .A(u5_mult_79_FS_1_n89), .ZN(u5_mult_79_FS_1_n83) );
  AND2_X1 u5_mult_79_FS_1_U102 ( .A1(u5_mult_79_n71), .A2(u5_mult_79_n26), 
        .ZN(u5_mult_79_FS_1_n84) );
  NOR2_X1 u5_mult_79_FS_1_U101 ( .A1(u5_mult_79_n71), .A2(u5_mult_79_n26), 
        .ZN(u5_mult_79_FS_1_n85) );
  NOR2_X1 u5_mult_79_FS_1_U100 ( .A1(u5_mult_79_FS_1_n84), .A2(
        u5_mult_79_FS_1_n85), .ZN(u5_mult_79_FS_1_n86) );
  XOR2_X1 u5_mult_79_FS_1_U99 ( .A(u5_mult_79_FS_1_n83), .B(
        u5_mult_79_FS_1_n86), .Z(u5_N32) );
  NOR2_X1 u5_mult_79_FS_1_U98 ( .A1(u5_mult_79_n75), .A2(u5_mult_79_n32), .ZN(
        u5_mult_79_FS_1_n79) );
  NAND2_X1 u5_mult_79_FS_1_U97 ( .A1(u5_mult_79_n75), .A2(u5_mult_79_n32), 
        .ZN(u5_mult_79_FS_1_n81) );
  NAND2_X1 u5_mult_79_FS_1_U96 ( .A1(u5_mult_79_FS_1_n17), .A2(
        u5_mult_79_FS_1_n81), .ZN(u5_mult_79_FS_1_n82) );
  AOI21_X1 u5_mult_79_FS_1_U95 ( .B1(u5_mult_79_FS_1_n18), .B2(
        u5_mult_79_FS_1_n83), .A(u5_mult_79_FS_1_n84), .ZN(u5_mult_79_FS_1_n80) );
  XOR2_X1 u5_mult_79_FS_1_U94 ( .A(u5_mult_79_FS_1_n82), .B(
        u5_mult_79_FS_1_n80), .Z(u5_N33) );
  OAI21_X1 u5_mult_79_FS_1_U93 ( .B1(u5_mult_79_FS_1_n79), .B2(
        u5_mult_79_FS_1_n80), .A(u5_mult_79_FS_1_n81), .ZN(u5_mult_79_FS_1_n75) );
  AND2_X1 u5_mult_79_FS_1_U92 ( .A1(u5_mult_79_n70), .A2(u5_mult_79_n25), .ZN(
        u5_mult_79_FS_1_n76) );
  NOR2_X1 u5_mult_79_FS_1_U91 ( .A1(u5_mult_79_n70), .A2(u5_mult_79_n25), .ZN(
        u5_mult_79_FS_1_n77) );
  NOR2_X1 u5_mult_79_FS_1_U90 ( .A1(u5_mult_79_FS_1_n76), .A2(
        u5_mult_79_FS_1_n77), .ZN(u5_mult_79_FS_1_n78) );
  XOR2_X1 u5_mult_79_FS_1_U89 ( .A(u5_mult_79_FS_1_n75), .B(
        u5_mult_79_FS_1_n78), .Z(u5_N34) );
  NOR2_X1 u5_mult_79_FS_1_U88 ( .A1(u5_mult_79_n90), .A2(u5_mult_79_n31), .ZN(
        u5_mult_79_FS_1_n71) );
  NAND2_X1 u5_mult_79_FS_1_U87 ( .A1(u5_mult_79_n90), .A2(u5_mult_79_n31), 
        .ZN(u5_mult_79_FS_1_n73) );
  NAND2_X1 u5_mult_79_FS_1_U86 ( .A1(u5_mult_79_FS_1_n15), .A2(
        u5_mult_79_FS_1_n73), .ZN(u5_mult_79_FS_1_n74) );
  AOI21_X1 u5_mult_79_FS_1_U85 ( .B1(u5_mult_79_FS_1_n16), .B2(
        u5_mult_79_FS_1_n75), .A(u5_mult_79_FS_1_n76), .ZN(u5_mult_79_FS_1_n72) );
  XOR2_X1 u5_mult_79_FS_1_U84 ( .A(u5_mult_79_FS_1_n74), .B(
        u5_mult_79_FS_1_n72), .Z(u5_N35) );
  OAI21_X1 u5_mult_79_FS_1_U83 ( .B1(u5_mult_79_FS_1_n71), .B2(
        u5_mult_79_FS_1_n72), .A(u5_mult_79_FS_1_n73), .ZN(u5_mult_79_FS_1_n67) );
  AND2_X1 u5_mult_79_FS_1_U82 ( .A1(u5_mult_79_n84), .A2(u5_mult_79_n40), .ZN(
        u5_mult_79_FS_1_n68) );
  NOR2_X1 u5_mult_79_FS_1_U81 ( .A1(u5_mult_79_n84), .A2(u5_mult_79_n40), .ZN(
        u5_mult_79_FS_1_n69) );
  NOR2_X1 u5_mult_79_FS_1_U80 ( .A1(u5_mult_79_FS_1_n68), .A2(
        u5_mult_79_FS_1_n69), .ZN(u5_mult_79_FS_1_n70) );
  XOR2_X1 u5_mult_79_FS_1_U79 ( .A(u5_mult_79_FS_1_n67), .B(
        u5_mult_79_FS_1_n70), .Z(u5_N36) );
  NOR2_X1 u5_mult_79_FS_1_U78 ( .A1(u5_mult_79_n89), .A2(u5_mult_79_n45), .ZN(
        u5_mult_79_FS_1_n63) );
  NAND2_X1 u5_mult_79_FS_1_U77 ( .A1(u5_mult_79_n89), .A2(u5_mult_79_n45), 
        .ZN(u5_mult_79_FS_1_n65) );
  NAND2_X1 u5_mult_79_FS_1_U76 ( .A1(u5_mult_79_FS_1_n13), .A2(
        u5_mult_79_FS_1_n65), .ZN(u5_mult_79_FS_1_n66) );
  AOI21_X1 u5_mult_79_FS_1_U75 ( .B1(u5_mult_79_FS_1_n14), .B2(
        u5_mult_79_FS_1_n67), .A(u5_mult_79_FS_1_n68), .ZN(u5_mult_79_FS_1_n64) );
  XOR2_X1 u5_mult_79_FS_1_U74 ( .A(u5_mult_79_FS_1_n66), .B(
        u5_mult_79_FS_1_n64), .Z(u5_N37) );
  OAI21_X1 u5_mult_79_FS_1_U73 ( .B1(u5_mult_79_FS_1_n63), .B2(
        u5_mult_79_FS_1_n64), .A(u5_mult_79_FS_1_n65), .ZN(u5_mult_79_FS_1_n59) );
  AND2_X1 u5_mult_79_FS_1_U72 ( .A1(u5_mult_79_n83), .A2(u5_mult_79_n39), .ZN(
        u5_mult_79_FS_1_n60) );
  NOR2_X1 u5_mult_79_FS_1_U71 ( .A1(u5_mult_79_n83), .A2(u5_mult_79_n39), .ZN(
        u5_mult_79_FS_1_n61) );
  NOR2_X1 u5_mult_79_FS_1_U70 ( .A1(u5_mult_79_FS_1_n60), .A2(
        u5_mult_79_FS_1_n61), .ZN(u5_mult_79_FS_1_n62) );
  XOR2_X1 u5_mult_79_FS_1_U69 ( .A(u5_mult_79_FS_1_n59), .B(
        u5_mult_79_FS_1_n62), .Z(u5_N38) );
  NOR2_X1 u5_mult_79_FS_1_U68 ( .A1(u5_mult_79_n88), .A2(u5_mult_79_n44), .ZN(
        u5_mult_79_FS_1_n55) );
  NAND2_X1 u5_mult_79_FS_1_U67 ( .A1(u5_mult_79_n88), .A2(u5_mult_79_n44), 
        .ZN(u5_mult_79_FS_1_n57) );
  NAND2_X1 u5_mult_79_FS_1_U66 ( .A1(u5_mult_79_FS_1_n11), .A2(
        u5_mult_79_FS_1_n57), .ZN(u5_mult_79_FS_1_n58) );
  AOI21_X1 u5_mult_79_FS_1_U65 ( .B1(u5_mult_79_FS_1_n12), .B2(
        u5_mult_79_FS_1_n59), .A(u5_mult_79_FS_1_n60), .ZN(u5_mult_79_FS_1_n56) );
  XOR2_X1 u5_mult_79_FS_1_U64 ( .A(u5_mult_79_FS_1_n58), .B(
        u5_mult_79_FS_1_n56), .Z(u5_N39) );
  OAI21_X1 u5_mult_79_FS_1_U63 ( .B1(u5_mult_79_FS_1_n55), .B2(
        u5_mult_79_FS_1_n56), .A(u5_mult_79_FS_1_n57), .ZN(u5_mult_79_FS_1_n51) );
  AND2_X1 u5_mult_79_FS_1_U62 ( .A1(u5_mult_79_n82), .A2(u5_mult_79_n38), .ZN(
        u5_mult_79_FS_1_n52) );
  NOR2_X1 u5_mult_79_FS_1_U61 ( .A1(u5_mult_79_n82), .A2(u5_mult_79_n38), .ZN(
        u5_mult_79_FS_1_n53) );
  NOR2_X1 u5_mult_79_FS_1_U60 ( .A1(u5_mult_79_FS_1_n52), .A2(
        u5_mult_79_FS_1_n53), .ZN(u5_mult_79_FS_1_n54) );
  XOR2_X1 u5_mult_79_FS_1_U59 ( .A(u5_mult_79_FS_1_n51), .B(
        u5_mult_79_FS_1_n54), .Z(u5_N40) );
  NOR2_X1 u5_mult_79_FS_1_U58 ( .A1(u5_mult_79_n87), .A2(u5_mult_79_n43), .ZN(
        u5_mult_79_FS_1_n47) );
  NAND2_X1 u5_mult_79_FS_1_U57 ( .A1(u5_mult_79_n87), .A2(u5_mult_79_n43), 
        .ZN(u5_mult_79_FS_1_n49) );
  NAND2_X1 u5_mult_79_FS_1_U56 ( .A1(u5_mult_79_FS_1_n9), .A2(
        u5_mult_79_FS_1_n49), .ZN(u5_mult_79_FS_1_n50) );
  AOI21_X1 u5_mult_79_FS_1_U55 ( .B1(u5_mult_79_FS_1_n10), .B2(
        u5_mult_79_FS_1_n51), .A(u5_mult_79_FS_1_n52), .ZN(u5_mult_79_FS_1_n48) );
  XOR2_X1 u5_mult_79_FS_1_U54 ( .A(u5_mult_79_FS_1_n50), .B(
        u5_mult_79_FS_1_n48), .Z(u5_N41) );
  OAI21_X1 u5_mult_79_FS_1_U53 ( .B1(u5_mult_79_FS_1_n47), .B2(
        u5_mult_79_FS_1_n48), .A(u5_mult_79_FS_1_n49), .ZN(u5_mult_79_FS_1_n43) );
  AND2_X1 u5_mult_79_FS_1_U52 ( .A1(u5_mult_79_n81), .A2(u5_mult_79_n37), .ZN(
        u5_mult_79_FS_1_n44) );
  NOR2_X1 u5_mult_79_FS_1_U51 ( .A1(u5_mult_79_n81), .A2(u5_mult_79_n37), .ZN(
        u5_mult_79_FS_1_n45) );
  NOR2_X1 u5_mult_79_FS_1_U50 ( .A1(u5_mult_79_FS_1_n44), .A2(
        u5_mult_79_FS_1_n45), .ZN(u5_mult_79_FS_1_n46) );
  XOR2_X1 u5_mult_79_FS_1_U49 ( .A(u5_mult_79_FS_1_n43), .B(
        u5_mult_79_FS_1_n46), .Z(u5_N42) );
  NOR2_X1 u5_mult_79_FS_1_U48 ( .A1(u5_mult_79_n86), .A2(u5_mult_79_n42), .ZN(
        u5_mult_79_FS_1_n39) );
  NAND2_X1 u5_mult_79_FS_1_U47 ( .A1(u5_mult_79_n86), .A2(u5_mult_79_n42), 
        .ZN(u5_mult_79_FS_1_n41) );
  NAND2_X1 u5_mult_79_FS_1_U46 ( .A1(u5_mult_79_FS_1_n7), .A2(
        u5_mult_79_FS_1_n41), .ZN(u5_mult_79_FS_1_n42) );
  AOI21_X1 u5_mult_79_FS_1_U45 ( .B1(u5_mult_79_FS_1_n8), .B2(
        u5_mult_79_FS_1_n43), .A(u5_mult_79_FS_1_n44), .ZN(u5_mult_79_FS_1_n40) );
  XOR2_X1 u5_mult_79_FS_1_U44 ( .A(u5_mult_79_FS_1_n42), .B(
        u5_mult_79_FS_1_n40), .Z(u5_N43) );
  OAI21_X1 u5_mult_79_FS_1_U43 ( .B1(u5_mult_79_FS_1_n39), .B2(
        u5_mult_79_FS_1_n40), .A(u5_mult_79_FS_1_n41), .ZN(u5_mult_79_FS_1_n35) );
  AND2_X1 u5_mult_79_FS_1_U42 ( .A1(u5_mult_79_n80), .A2(u5_mult_79_n36), .ZN(
        u5_mult_79_FS_1_n36) );
  NOR2_X1 u5_mult_79_FS_1_U41 ( .A1(u5_mult_79_n80), .A2(u5_mult_79_n36), .ZN(
        u5_mult_79_FS_1_n37) );
  NOR2_X1 u5_mult_79_FS_1_U40 ( .A1(u5_mult_79_FS_1_n36), .A2(
        u5_mult_79_FS_1_n37), .ZN(u5_mult_79_FS_1_n38) );
  XOR2_X1 u5_mult_79_FS_1_U39 ( .A(u5_mult_79_FS_1_n35), .B(
        u5_mult_79_FS_1_n38), .Z(u5_N44) );
  NOR2_X1 u5_mult_79_FS_1_U38 ( .A1(u5_mult_79_n85), .A2(u5_mult_79_n41), .ZN(
        u5_mult_79_FS_1_n31) );
  NAND2_X1 u5_mult_79_FS_1_U37 ( .A1(u5_mult_79_n85), .A2(u5_mult_79_n41), 
        .ZN(u5_mult_79_FS_1_n33) );
  NAND2_X1 u5_mult_79_FS_1_U36 ( .A1(u5_mult_79_FS_1_n5), .A2(
        u5_mult_79_FS_1_n33), .ZN(u5_mult_79_FS_1_n34) );
  AOI21_X1 u5_mult_79_FS_1_U35 ( .B1(u5_mult_79_FS_1_n6), .B2(
        u5_mult_79_FS_1_n35), .A(u5_mult_79_FS_1_n36), .ZN(u5_mult_79_FS_1_n32) );
  XOR2_X1 u5_mult_79_FS_1_U34 ( .A(u5_mult_79_FS_1_n34), .B(
        u5_mult_79_FS_1_n32), .Z(u5_N45) );
  OAI21_X1 u5_mult_79_FS_1_U33 ( .B1(u5_mult_79_FS_1_n31), .B2(
        u5_mult_79_FS_1_n32), .A(u5_mult_79_FS_1_n33), .ZN(u5_mult_79_FS_1_n27) );
  AND2_X1 u5_mult_79_FS_1_U32 ( .A1(u5_mult_79_n93), .A2(u5_mult_79_n46), .ZN(
        u5_mult_79_FS_1_n28) );
  NOR2_X1 u5_mult_79_FS_1_U31 ( .A1(u5_mult_79_n93), .A2(u5_mult_79_n46), .ZN(
        u5_mult_79_FS_1_n29) );
  NOR2_X1 u5_mult_79_FS_1_U30 ( .A1(u5_mult_79_FS_1_n28), .A2(
        u5_mult_79_FS_1_n29), .ZN(u5_mult_79_FS_1_n30) );
  XOR2_X1 u5_mult_79_FS_1_U29 ( .A(u5_mult_79_FS_1_n27), .B(
        u5_mult_79_FS_1_n30), .Z(u5_N46) );
  AOI21_X1 u5_mult_79_FS_1_U28 ( .B1(u5_mult_79_FS_1_n27), .B2(
        u5_mult_79_FS_1_n4), .A(u5_mult_79_FS_1_n28), .ZN(u5_mult_79_FS_1_n26)
         );
  XOR2_X1 u5_mult_79_FS_1_U27 ( .A(u5_mult_79_FS_1_n3), .B(u5_mult_79_FS_1_n26), .Z(u5_N47) );
  INV_X4 u5_mult_79_FS_1_U26 ( .A(u5_mult_79_FS_1_n110), .ZN(
        u5_mult_79_FS_1_n25) );
  INV_X4 u5_mult_79_FS_1_U25 ( .A(u5_mult_79_FS_1_n108), .ZN(
        u5_mult_79_FS_1_n24) );
  INV_X4 u5_mult_79_FS_1_U24 ( .A(u5_mult_79_FS_1_n103), .ZN(
        u5_mult_79_FS_1_n23) );
  INV_X4 u5_mult_79_FS_1_U23 ( .A(u5_mult_79_FS_1_n101), .ZN(
        u5_mult_79_FS_1_n22) );
  INV_X4 u5_mult_79_FS_1_U22 ( .A(u5_mult_79_FS_1_n95), .ZN(
        u5_mult_79_FS_1_n21) );
  INV_X4 u5_mult_79_FS_1_U21 ( .A(u5_mult_79_FS_1_n93), .ZN(
        u5_mult_79_FS_1_n20) );
  INV_X4 u5_mult_79_FS_1_U20 ( .A(u5_mult_79_FS_1_n87), .ZN(
        u5_mult_79_FS_1_n19) );
  INV_X4 u5_mult_79_FS_1_U19 ( .A(u5_mult_79_FS_1_n85), .ZN(
        u5_mult_79_FS_1_n18) );
  INV_X4 u5_mult_79_FS_1_U18 ( .A(u5_mult_79_FS_1_n79), .ZN(
        u5_mult_79_FS_1_n17) );
  INV_X4 u5_mult_79_FS_1_U17 ( .A(u5_mult_79_FS_1_n77), .ZN(
        u5_mult_79_FS_1_n16) );
  INV_X4 u5_mult_79_FS_1_U16 ( .A(u5_mult_79_FS_1_n71), .ZN(
        u5_mult_79_FS_1_n15) );
  INV_X4 u5_mult_79_FS_1_U15 ( .A(u5_mult_79_FS_1_n69), .ZN(
        u5_mult_79_FS_1_n14) );
  INV_X4 u5_mult_79_FS_1_U14 ( .A(u5_mult_79_FS_1_n63), .ZN(
        u5_mult_79_FS_1_n13) );
  INV_X4 u5_mult_79_FS_1_U13 ( .A(u5_mult_79_FS_1_n61), .ZN(
        u5_mult_79_FS_1_n12) );
  INV_X4 u5_mult_79_FS_1_U12 ( .A(u5_mult_79_FS_1_n55), .ZN(
        u5_mult_79_FS_1_n11) );
  INV_X4 u5_mult_79_FS_1_U11 ( .A(u5_mult_79_FS_1_n53), .ZN(
        u5_mult_79_FS_1_n10) );
  INV_X4 u5_mult_79_FS_1_U10 ( .A(u5_mult_79_FS_1_n47), .ZN(u5_mult_79_FS_1_n9) );
  INV_X4 u5_mult_79_FS_1_U9 ( .A(u5_mult_79_FS_1_n45), .ZN(u5_mult_79_FS_1_n8)
         );
  INV_X4 u5_mult_79_FS_1_U8 ( .A(u5_mult_79_FS_1_n39), .ZN(u5_mult_79_FS_1_n7)
         );
  INV_X4 u5_mult_79_FS_1_U7 ( .A(u5_mult_79_FS_1_n37), .ZN(u5_mult_79_FS_1_n6)
         );
  INV_X4 u5_mult_79_FS_1_U6 ( .A(u5_mult_79_FS_1_n31), .ZN(u5_mult_79_FS_1_n5)
         );
  INV_X4 u5_mult_79_FS_1_U5 ( .A(u5_mult_79_FS_1_n29), .ZN(u5_mult_79_FS_1_n4)
         );
  INV_X4 u5_mult_79_FS_1_U4 ( .A(u5_mult_79_n92), .ZN(u5_mult_79_FS_1_n3) );
  AND2_X4 u5_mult_79_FS_1_U3 ( .A1(u5_mult_79_FS_1_n1), .A2(
        u5_mult_79_FS_1_n110), .ZN(u5_N25) );
  OR2_X4 u5_mult_79_FS_1_U2 ( .A1(u5_mult_79_n79), .A2(u5_mult_79_n30), .ZN(
        u5_mult_79_FS_1_n1) );
endmodule

