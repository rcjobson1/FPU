
module fpu ( clk, rmode, fpu_op, opa, opb, out, inf, snan, qnan, ine, overflow, 
        underflow, zero, div_by_zero );
  input [1:0] rmode;
  input [2:0] fpu_op;
  input [15:0] opa;
  input [15:0] opb;
  output [15:0] out;
  input clk;
  output inf, snan, qnan, ine, overflow, underflow, zero, div_by_zero;
  wire   snan_d, opa_nan, opb_nan, opa_00, opb_00, opa_inf, opb_inf, opa_dn,
         opb_dn, sign_fasu, nan_sign_d, result_zero_sign_d, fasu_op,
         sign_fasu_r, sign_mul, sign_exe, inf_mul, sign_mul_r, sign_exe_r, N34,
         N44, N56, N65, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77,
         N96, N97, N98, N99, N100, N106, N110, N111, N112, N113, N114, N115,
         N116, fract_i2f_7_, N138, N139, N140, N141, N150, N151, N179, N180,
         N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191,
         N192, N193, N194, N195, N196, opas_r1, opas_r2, sign, N216,
         fasu_op_r1, N220, N221, N222, N223, N224, N225, N226, N227, N228,
         N229, N230, N231, N232, N233, N234, N254, N268, N278, N281, N283,
         N285, N290, N291, N292, N296, u0_N17, u0_N16, u0_expb_00, u0_expa_00,
         u0_N11, u0_N10, u0_N7, u0_N6, u0_N5, u0_N4, u0_infb_f_r, u0_infa_f_r,
         u0_expb_ff, u0_expa_ff, u1_N133, u1_fracta_eq_fractb, u1_N124,
         u1_fracta_lt_fractb, u1_N123, u1_N122, u1_add_r, u1_signa_r,
         u1_sign_d, u1_fractb_lt_fracta, u1_adj_op_out_sft_0_,
         u1_adj_op_out_sft_1_, u1_adj_op_out_sft_2_, u1_adj_op_out_sft_3_,
         u1_adj_op_out_sft_4_, u1_adj_op_out_sft_5_, u1_adj_op_out_sft_6_,
         u1_adj_op_out_sft_7_, u1_adj_op_out_sft_8_, u1_adj_op_out_sft_9_,
         u1_adj_op_out_sft_10_, u1_adj_op_out_sft_11_, u1_adj_op_out_sft_12_,
         u1_adj_op_out_sft_13_, u1_exp_diff_sft_0_, u1_exp_lt_27, u1_adj_op_9_,
         u1_N39, u1_N38, u1_N37, u1_N36, u1_N35, u1_N32, u1_exp_diff_1_,
         u1_exp_diff_2_, u1_exp_diff_3_, u1_exp_diff_4_, u1_expa_lt_expb,
         u2_N73, u2_sign_d, u2_N66, u2_exp_ovf_d_0_, u2_exp_ovf_d_1_, u2_N44,
         u2_N43, u2_N42, u2_N41, u2_N40, u2_N39, u2_N38, u2_N37, u2_N36,
         u2_N34, u2_N33, u2_N32, u2_N31, u2_exp_tmp4_0_, u2_exp_tmp4_1_,
         u2_exp_tmp4_2_, u2_exp_tmp4_3_, u2_exp_tmp4_4_, u2_exp_tmp3_1_,
         u2_exp_tmp3_2_, u2_exp_tmp3_3_, u2_exp_tmp3_4_, u2_N29, u2_N28,
         u2_N27, u2_N26, u2_N25, u2_N23, u2_N22, u2_N21, u2_N20, u2_N19,
         u2_N17, u2_N16, u2_N15, u2_N14, u2_N13, u2_N12, u2_N11, u2_N10, u2_N9,
         u2_N8, u2_N7, u2_N6, u3_N32, u3_N31, u3_N30, u3_N29, u3_N28, u3_N27,
         u3_N26, u3_N25, u3_N24, u3_N23, u3_N22, u3_N21, u3_N20, u3_N19,
         u3_N18, u3_N17, u3_N16, u3_N15, u3_N14, u3_N13, u3_N12, u3_N11,
         u3_N10, u3_N9, u3_N8, u3_N7, u3_N6, u3_N5, u3_N4, u3_N3, u5_N21,
         u5_N20, u5_N19, u5_N18, u5_N17, u5_N16, u5_N15, u5_N14, u5_N13,
         u5_N12, u5_N11, u5_N10, u5_N9, u5_N8, u5_N7, u5_N6, u5_N5, u5_N4,
         u5_N3, u5_N2, u5_N1, u5_N0, u6_N23, u6_N22, u6_N21, u6_N20, u6_N19,
         u6_N18, u6_N17, u6_N16, u6_N15, u6_N14, u6_N13, u6_N10, u6_N9, u6_N8,
         u6_N7, u6_N6, u6_N5, u6_N4, u6_N3, u6_N2, u6_N1, u6_N0, u4_N798,
         u4_N797, u4_N796, u4_N656, u4_N655, u4_N654, u4_N653, u4_N581,
         u4_N558, u4_N487, u4_div_exp1_0_, u4_div_exp1_1_, u4_div_exp1_2_,
         u4_div_exp1_3_, u4_div_exp1_4_, u4_fi_ldz_2a_0_, u4_fi_ldz_2a_1_,
         u4_fi_ldz_2a_2_, u4_fi_ldz_2a_3_, u4_fi_ldz_2a_4_, u4_ldz_all_1_,
         u4_ldz_all_2_, u4_ldz_all_3_, u4_ldz_all_4_, u4_ldz_all_5_, u4_N447,
         u4_N446, u4_N445, u4_N444, u4_exp_out_pl1_1_, u4_exp_out_pl1_2_,
         u4_exp_out_pl1_3_, u4_exp_out_pl1_4_, u4_fi_ldz_mi1_1_,
         u4_fi_ldz_mi1_2_, u4_fi_ldz_mi1_3_, u4_fi_ldz_mi1_4_,
         u4_fi_ldz_mi1_6_, u4_N433, u4_N432, u4_N431, u4_N430, u4_N429,
         u4_N428, u4_N427, u4_N426, u4_N425, u4_N424, u4_N423, u4_N422,
         u4_N421, u4_N420, u4_N419, u4_N418, u4_N417, u4_N416, u4_N415,
         u4_N414, u4_N413, u4_N412, u4_N409, u4_N408, u4_N407, u4_N406,
         u4_N405, u4_N404, u4_N403, u4_N402, u4_N401, u4_N400, u4_N399,
         u4_N398, u4_N397, u4_N396, u4_N395, u4_N394, u4_N393, u4_N392,
         u4_N391, u4_N390, u4_N389, u4_N388, u4_N386, u4_exp_in_pl1_0_,
         u4_exp_in_pl1_1_, u4_exp_in_pl1_2_, u4_exp_in_pl1_3_,
         u4_exp_in_pl1_4_, u4_exp_in_pl1_5_, u4_f2i_shft_0_, u4_f2i_shft_1_,
         u4_f2i_shft_2_, u4_f2i_shft_3_, u4_f2i_shft_4_, u4_N326,
         u4_div_shft3_0_, u4_div_shft3_1_, u4_div_shft3_2_, u4_div_shft3_3_,
         u4_div_shft3_4_, u4_exp_in_mi1_1_, u4_exp_in_mi1_2_, u4_exp_in_mi1_3_,
         u4_exp_in_mi1_4_, u4_exp_in_mi1_5_, u4_fract_out_pl1_0_,
         u4_fract_out_pl1_1_, u4_fract_out_pl1_2_, u4_fract_out_pl1_3_,
         u4_fract_out_pl1_4_, u4_fract_out_pl1_5_, u4_fract_out_pl1_6_,
         u4_fract_out_pl1_7_, u4_fract_out_pl1_8_, u4_fract_out_pl1_9_,
         u4_fract_out_pl1_10_, u4_exp_next_mi_0_, u4_exp_next_mi_1_,
         u4_exp_next_mi_2_, u4_exp_next_mi_3_, u4_exp_next_mi_4_,
         u4_exp_next_mi_5_, u4_fract_out_0_, u4_fract_out_1_, u4_fract_out_2_,
         u4_fract_out_3_, u4_fract_out_4_, u4_fract_out_5_, u4_fract_out_6_,
         u4_fract_out_7_, u4_fract_out_8_, u4_fract_out_9_, u4_exp_out_0_,
         u4_exp_out_1_, u4_exp_out_2_, u4_exp_out_3_, u4_exp_out_4_, u4_N264,
         u4_N203, u4_N152, u4_N95, n831, n842, n845, n848, n850, n851, n852,
         n872, n888, n889, n1521, n1522, n1523, u4_ldz_dif_4_, u4_ldz_dif_3_,
         u4_ldz_dif_2_, u4_ldz_dif_1_, u4_ldz_dif_0_, u4_fi_ldz_mi22_4_,
         u4_fi_ldz_mi22_3_, u4_fi_ldz_mi22_2_, u4_fi_ldz_mi22_1_,
         u2_lt_130_A_0_, u2_lt_130_A_1_, u2_lt_130_A_2_, u2_lt_130_A_3_,
         u2_gt_140_B_5_, u1_gt_234_B_0_, u1_gt_234_B_1_, u1_gt_234_B_2_,
         u1_gt_234_B_3_, u1_gt_234_B_4_, u1_gt_234_B_5_, u1_gt_234_B_6_,
         u1_gt_234_B_7_, u1_gt_234_B_8_, u1_gt_234_B_9_, u1_gt_234_B_10_,
         u1_gt_234_B_11_, u1_gt_234_B_12_, u1_gt_234_B_13_, u1_gt_234_A_0_,
         u1_gt_234_A_1_, u1_gt_234_A_2_, u1_gt_234_A_3_, u1_gt_234_A_4_,
         u1_gt_234_A_5_, u1_gt_234_A_6_, u1_gt_234_A_7_, u1_gt_234_A_8_,
         u1_gt_234_A_9_, u1_gt_234_A_10_, u1_gt_234_A_11_, u1_gt_234_A_12_,
         u1_gt_234_A_13_, u1_gt_144_B_0_, u4_sub_414_carry_2_,
         u4_sub_414_carry_3_, u4_sub_414_carry_4_, u4_sub_465_A_0_,
         u4_sub_465_A_1_, u4_sub_465_A_2_, u4_sub_465_A_3_, u4_sub_465_A_4_,
         u2_add_113_A_0_, u2_add_113_A_1_, u2_add_113_A_2_, u2_add_113_A_3_,
         u2_add_113_A_4_, u2_sub_111_carry_2_, u2_sub_111_carry_3_,
         u2_sub_111_carry_4_, u2_sub_111_carry_5_, u2_add_111_carry_2_,
         u2_add_111_carry_3_, u2_add_111_carry_4_, u2_add_111_carry_5_,
         sub_1_root_u1_sub_128_aco_CI, sub_1_root_u1_sub_128_aco_B_0_,
         sub_1_root_u1_sub_128_aco_B_1_, sub_1_root_u1_sub_128_aco_B_2_,
         sub_1_root_u1_sub_128_aco_A_0_, sub_1_root_u1_sub_128_aco_A_1_,
         sub_1_root_u1_sub_128_aco_A_2_, sub_1_root_u1_sub_128_aco_A_3_,
         sub_1_root_u1_sub_128_aco_A_4_,
         add_1_root_sub_0_root_u4_sub_469_carry_2_,
         add_1_root_sub_0_root_u4_sub_469_carry_3_,
         add_1_root_sub_0_root_u4_sub_469_carry_4_, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         u4_srl_450_n76, u4_srl_450_n75, u4_srl_450_n74, u4_srl_450_n73,
         u4_srl_450_n72, u4_srl_450_n71, u4_srl_450_n70, u4_srl_450_n69,
         u4_srl_450_n68, u4_srl_450_n67, u4_srl_450_n66, u4_srl_450_n65,
         u4_srl_450_n64, u4_srl_450_n63, u4_srl_450_n62, u4_srl_450_n61,
         u4_srl_450_n60, u4_srl_450_n59, u4_srl_450_n58, u4_srl_450_n57,
         u4_srl_450_n56, u4_srl_450_n55, u4_srl_450_n54, u4_srl_450_n53,
         u4_srl_450_n52, u4_srl_450_n51, u4_srl_450_n50, u4_srl_450_n49,
         u4_srl_450_n48, u4_srl_450_n47, u4_srl_450_n46, u4_srl_450_n45,
         u4_srl_450_n44, u4_srl_450_n43, u4_srl_450_n42, u4_srl_450_n41,
         u4_srl_450_n40, u4_srl_450_n39, u4_srl_450_n38, u4_srl_450_n37,
         u4_srl_450_n36, u4_srl_450_n35, u4_srl_450_n34, u4_srl_450_n33,
         u4_srl_450_n32, u4_srl_450_n31, u4_srl_450_n30, u4_srl_450_n29,
         u4_srl_450_n28, u4_srl_450_n27, u4_srl_450_n26, u4_srl_450_n25,
         u4_srl_450_n24, u4_srl_450_n23, u4_srl_450_n22, u4_srl_450_n21,
         u4_srl_450_n20, u4_srl_450_n19, u4_srl_450_n18, u4_srl_450_n17,
         u4_srl_450_n16, u4_srl_450_n15, u4_srl_450_n14, u4_srl_450_n13,
         u4_srl_450_n12, u4_srl_450_n11, u4_srl_450_n10, u4_srl_450_n9,
         u4_srl_450_n8, u4_srl_450_n7, u4_srl_450_n6, u4_srl_450_n5,
         u4_srl_450_n4, u4_srl_450_n3, u4_srl_450_n2, u4_srl_450_n1,
         u4_sll_451_n8, u4_sll_451_n7, u4_sll_451_n6, u4_sll_451_n5,
         u4_sll_451_n4, u4_sll_451_n3, u4_sll_451_n2, u4_sll_451_n1,
         u4_sll_451_ML_int_2__0_, u4_sll_451_ML_int_2__1_,
         u4_sll_451_ML_int_2__2_, u4_sll_451_ML_int_2__3_,
         u4_sll_451_ML_int_2__4_, u4_sll_451_ML_int_2__5_,
         u4_sll_451_ML_int_2__6_, u4_sll_451_ML_int_2__7_,
         u4_sll_451_ML_int_2__8_, u4_sll_451_ML_int_2__9_,
         u4_sll_451_ML_int_2__10_, u4_sll_451_ML_int_2__11_,
         u4_sll_451_ML_int_2__12_, u4_sll_451_ML_int_2__13_,
         u4_sll_451_ML_int_2__14_, u4_sll_451_ML_int_2__15_,
         u4_sll_451_ML_int_2__16_, u4_sll_451_ML_int_2__17_,
         u4_sll_451_ML_int_2__18_, u4_sll_451_ML_int_2__19_,
         u4_sll_451_ML_int_2__20_, u4_sll_451_ML_int_2__21_,
         u4_sll_451_ML_int_1__0_, u4_sll_451_ML_int_1__1_,
         u4_sll_451_ML_int_1__2_, u4_sll_451_ML_int_1__3_,
         u4_sll_451_ML_int_1__4_, u4_sll_451_ML_int_1__5_,
         u4_sll_451_ML_int_1__6_, u4_sll_451_ML_int_1__7_,
         u4_sll_451_ML_int_1__8_, u4_sll_451_ML_int_1__9_,
         u4_sll_451_ML_int_1__10_, u4_sll_451_ML_int_1__11_,
         u4_sll_451_ML_int_1__12_, u4_sll_451_ML_int_1__13_,
         u4_sll_451_ML_int_1__14_, u4_sll_451_ML_int_1__15_,
         u4_sll_451_ML_int_1__16_, u4_sll_451_ML_int_1__17_,
         u4_sll_451_ML_int_1__18_, u4_sll_451_ML_int_1__19_,
         u4_sll_451_ML_int_1__20_, u4_sll_451_ML_int_1__21_, u4_sll_479_n11,
         u4_sll_479_n10, u4_sll_479_n9, u4_sll_479_n8, u4_sll_479_n7,
         u4_sll_479_n6, u4_sll_479_n5, u4_sll_479_n4, u4_sll_479_n3,
         u4_sll_479_n2, u4_sll_479_n1, u4_sll_479_ML_int_4__7_,
         u4_sll_479_ML_int_4__8_, u4_sll_479_ML_int_4__9_,
         u4_sll_479_ML_int_4__10_, u4_sll_479_ML_int_4__11_,
         u4_sll_479_ML_int_4__23_, u4_sll_479_ML_int_4__24_,
         u4_sll_479_ML_int_4__25_, u4_sll_479_ML_int_4__26_,
         u4_sll_479_ML_int_4__27_, u4_sll_479_ML_int_3__0_,
         u4_sll_479_ML_int_3__1_, u4_sll_479_ML_int_3__2_,
         u4_sll_479_ML_int_3__3_, u4_sll_479_ML_int_3__7_,
         u4_sll_479_ML_int_3__8_, u4_sll_479_ML_int_3__9_,
         u4_sll_479_ML_int_3__10_, u4_sll_479_ML_int_3__11_,
         u4_sll_479_ML_int_3__15_, u4_sll_479_ML_int_3__16_,
         u4_sll_479_ML_int_3__17_, u4_sll_479_ML_int_3__18_,
         u4_sll_479_ML_int_3__19_, u4_sll_479_ML_int_3__23_,
         u4_sll_479_ML_int_3__24_, u4_sll_479_ML_int_3__25_,
         u4_sll_479_ML_int_3__26_, u4_sll_479_ML_int_3__27_,
         u4_sll_479_ML_int_2__2_, u4_sll_479_ML_int_2__3_,
         u4_sll_479_ML_int_2__4_, u4_sll_479_ML_int_2__5_,
         u4_sll_479_ML_int_2__6_, u4_sll_479_ML_int_2__7_,
         u4_sll_479_ML_int_2__8_, u4_sll_479_ML_int_2__9_,
         u4_sll_479_ML_int_2__10_, u4_sll_479_ML_int_2__11_,
         u4_sll_479_ML_int_2__12_, u4_sll_479_ML_int_2__13_,
         u4_sll_479_ML_int_2__14_, u4_sll_479_ML_int_2__15_,
         u4_sll_479_ML_int_2__16_, u4_sll_479_ML_int_2__17_,
         u4_sll_479_ML_int_2__18_, u4_sll_479_ML_int_2__19_,
         u4_sll_479_ML_int_2__20_, u4_sll_479_ML_int_2__21_,
         u4_sll_479_ML_int_2__22_, u4_sll_479_ML_int_2__23_,
         u4_sll_479_ML_int_2__24_, u4_sll_479_ML_int_2__25_,
         u4_sll_479_ML_int_2__26_, u4_sll_479_ML_int_2__27_,
         u4_sll_479_ML_int_1__0_, u4_sll_479_ML_int_1__1_,
         u4_sll_479_ML_int_1__2_, u4_sll_479_ML_int_1__3_,
         u4_sll_479_ML_int_1__4_, u4_sll_479_ML_int_1__5_,
         u4_sll_479_ML_int_1__6_, u4_sll_479_ML_int_1__7_,
         u4_sll_479_ML_int_1__8_, u4_sll_479_ML_int_1__9_,
         u4_sll_479_ML_int_1__10_, u4_sll_479_ML_int_1__11_,
         u4_sll_479_ML_int_1__12_, u4_sll_479_ML_int_1__13_,
         u4_sll_479_ML_int_1__14_, u4_sll_479_ML_int_1__15_,
         u4_sll_479_ML_int_1__16_, u4_sll_479_ML_int_1__17_,
         u4_sll_479_ML_int_1__18_, u4_sll_479_ML_int_1__19_,
         u4_sll_479_ML_int_1__20_, u4_sll_479_ML_int_1__21_,
         u4_sll_479_ML_int_1__22_, u4_sll_479_ML_int_1__23_,
         u4_sll_479_ML_int_1__24_, u4_sll_479_ML_int_1__25_,
         u4_sll_479_ML_int_1__26_, u4_sll_479_ML_int_1__27_, u4_sub_467_n7,
         u4_sub_467_n6, u4_sub_467_n5, u4_sub_467_n4, u4_sub_467_n3,
         u4_sub_467_n2, u4_sub_467_n1, u3_sub_59_n16, u3_sub_59_n15,
         u3_sub_59_n14, u3_sub_59_n13, u3_sub_59_n12, u3_sub_59_n11,
         u3_sub_59_n10, u3_sub_59_n9, u3_sub_59_n8, u3_sub_59_n7, u3_sub_59_n6,
         u3_sub_59_n5, u3_sub_59_n4, u3_sub_59_n3, u3_sub_59_n1, u3_add_59_n1,
         u1_srl_146_n47, u1_srl_146_n46, u1_srl_146_n45, u1_srl_146_n44,
         u1_srl_146_n43, u1_srl_146_n42, u1_srl_146_n41, u1_srl_146_n40,
         u1_srl_146_n39, u1_srl_146_n38, u1_srl_146_n37, u1_srl_146_n36,
         u1_srl_146_n35, u1_srl_146_n34, u1_srl_146_n33, u1_srl_146_n32,
         u1_srl_146_n31, u1_srl_146_n30, u1_srl_146_n29, u1_srl_146_n28,
         u1_srl_146_n27, u1_srl_146_n26, u1_srl_146_n25, u1_srl_146_n24,
         u1_srl_146_n23, u1_srl_146_n22, u1_srl_146_n21, u1_srl_146_n20,
         u1_srl_146_n19, u1_srl_146_n18, u1_srl_146_n17, u1_srl_146_n16,
         u1_srl_146_n15, u1_srl_146_n14, u1_srl_146_n13, u1_srl_146_n12,
         u1_srl_146_n11, u1_srl_146_n10, u1_srl_146_n9, u1_srl_146_n8,
         u1_srl_146_n7, u1_srl_146_n6, u1_srl_146_n5, u1_srl_146_n4,
         u1_srl_146_n3, u1_srl_146_n2, u1_srl_146_n1, sll_384_n11, sll_384_n10,
         sll_384_n9, sll_384_n8, sll_384_n7, sll_384_n6, sll_384_n5,
         sll_384_n4, sll_384_n3, sll_384_n2, sll_384_n1, sll_384_ML_int_3__0_,
         sll_384_ML_int_3__1_, sll_384_ML_int_3__2_, sll_384_ML_int_3__4_,
         sll_384_ML_int_3__5_, sll_384_ML_int_3__6_, sll_384_ML_int_3__7_,
         sll_384_ML_int_3__8_, sll_384_ML_int_3__9_, sll_384_ML_int_3__10_,
         sll_384_ML_int_2__2_, sll_384_ML_int_2__3_, sll_384_ML_int_2__4_,
         sll_384_ML_int_2__5_, sll_384_ML_int_2__6_, sll_384_ML_int_2__7_,
         sll_384_ML_int_2__8_, sll_384_ML_int_2__9_, sll_384_ML_int_2__10_,
         sll_384_ML_int_1__0_, sll_384_ML_int_1__1_, sll_384_ML_int_1__2_,
         sll_384_ML_int_1__3_, sll_384_ML_int_1__4_, sll_384_ML_int_1__5_,
         sll_384_ML_int_1__6_, sll_384_ML_int_1__7_, sll_384_ML_int_1__8_,
         sll_384_ML_int_1__9_, sll_384_ML_int_1__10_, u5_mult_78_n64,
         u5_mult_78_n63, u5_mult_78_n62, u5_mult_78_n61, u5_mult_78_n60,
         u5_mult_78_n59, u5_mult_78_n58, u5_mult_78_n57, u5_mult_78_n56,
         u5_mult_78_n55, u5_mult_78_n54, u5_mult_78_n53, u5_mult_78_n52,
         u5_mult_78_n51, u5_mult_78_n50, u5_mult_78_n49, u5_mult_78_n48,
         u5_mult_78_n47, u5_mult_78_n46, u5_mult_78_n45, u5_mult_78_n44,
         u5_mult_78_n43, u5_mult_78_n40, u5_mult_78_n39, u5_mult_78_n38,
         u5_mult_78_n37, u5_mult_78_n36, u5_mult_78_n35, u5_mult_78_n34,
         u5_mult_78_n33, u5_mult_78_n32, u5_mult_78_n31, u5_mult_78_n30,
         u5_mult_78_n29, u5_mult_78_n28, u5_mult_78_n27, u5_mult_78_n26,
         u5_mult_78_n25, u5_mult_78_n24, u5_mult_78_n23, u5_mult_78_n22,
         u5_mult_78_n21, u5_mult_78_n20, u5_mult_78_n19, u5_mult_78_n18,
         u5_mult_78_n17, u5_mult_78_n16, u5_mult_78_n15, u5_mult_78_n14,
         u5_mult_78_n13, u5_mult_78_n12, u5_mult_78_n11, u5_mult_78_n10,
         u5_mult_78_n9, u5_mult_78_n8, u5_mult_78_n7, u5_mult_78_n6,
         u5_mult_78_n5, u5_mult_78_n4, u5_mult_78_n3, u5_mult_78_SUMB_2__1_,
         u5_mult_78_SUMB_2__2_, u5_mult_78_SUMB_2__3_, u5_mult_78_SUMB_2__4_,
         u5_mult_78_SUMB_2__5_, u5_mult_78_SUMB_2__6_, u5_mult_78_SUMB_2__7_,
         u5_mult_78_SUMB_2__8_, u5_mult_78_SUMB_2__9_, u5_mult_78_SUMB_3__1_,
         u5_mult_78_SUMB_3__2_, u5_mult_78_SUMB_3__3_, u5_mult_78_SUMB_3__4_,
         u5_mult_78_SUMB_3__5_, u5_mult_78_SUMB_3__6_, u5_mult_78_SUMB_3__7_,
         u5_mult_78_SUMB_3__8_, u5_mult_78_SUMB_3__9_, u5_mult_78_SUMB_4__1_,
         u5_mult_78_SUMB_4__2_, u5_mult_78_SUMB_4__3_, u5_mult_78_SUMB_4__4_,
         u5_mult_78_SUMB_4__5_, u5_mult_78_SUMB_4__6_, u5_mult_78_SUMB_4__7_,
         u5_mult_78_SUMB_4__8_, u5_mult_78_SUMB_4__9_, u5_mult_78_SUMB_5__1_,
         u5_mult_78_SUMB_5__2_, u5_mult_78_SUMB_5__3_, u5_mult_78_SUMB_5__4_,
         u5_mult_78_SUMB_5__5_, u5_mult_78_SUMB_5__6_, u5_mult_78_SUMB_5__7_,
         u5_mult_78_SUMB_5__8_, u5_mult_78_SUMB_5__9_, u5_mult_78_SUMB_6__1_,
         u5_mult_78_SUMB_6__2_, u5_mult_78_SUMB_6__3_, u5_mult_78_SUMB_6__4_,
         u5_mult_78_SUMB_6__5_, u5_mult_78_SUMB_6__6_, u5_mult_78_SUMB_6__7_,
         u5_mult_78_SUMB_6__8_, u5_mult_78_SUMB_6__9_, u5_mult_78_SUMB_7__1_,
         u5_mult_78_SUMB_7__2_, u5_mult_78_SUMB_7__3_, u5_mult_78_SUMB_7__4_,
         u5_mult_78_SUMB_7__5_, u5_mult_78_SUMB_7__6_, u5_mult_78_SUMB_7__7_,
         u5_mult_78_SUMB_7__8_, u5_mult_78_SUMB_7__9_, u5_mult_78_SUMB_8__1_,
         u5_mult_78_SUMB_8__2_, u5_mult_78_SUMB_8__3_, u5_mult_78_SUMB_8__4_,
         u5_mult_78_SUMB_8__5_, u5_mult_78_SUMB_8__6_, u5_mult_78_SUMB_8__7_,
         u5_mult_78_SUMB_8__8_, u5_mult_78_SUMB_8__9_, u5_mult_78_SUMB_9__1_,
         u5_mult_78_SUMB_9__2_, u5_mult_78_SUMB_9__3_, u5_mult_78_SUMB_9__4_,
         u5_mult_78_SUMB_9__5_, u5_mult_78_SUMB_9__6_, u5_mult_78_SUMB_9__7_,
         u5_mult_78_SUMB_9__8_, u5_mult_78_SUMB_9__9_, u5_mult_78_SUMB_10__1_,
         u5_mult_78_SUMB_10__2_, u5_mult_78_SUMB_10__3_,
         u5_mult_78_SUMB_10__4_, u5_mult_78_SUMB_10__5_,
         u5_mult_78_SUMB_10__6_, u5_mult_78_SUMB_10__7_,
         u5_mult_78_SUMB_10__8_, u5_mult_78_SUMB_10__9_,
         u5_mult_78_CARRYB_2__0_, u5_mult_78_CARRYB_2__1_,
         u5_mult_78_CARRYB_2__2_, u5_mult_78_CARRYB_2__3_,
         u5_mult_78_CARRYB_2__4_, u5_mult_78_CARRYB_2__5_,
         u5_mult_78_CARRYB_2__6_, u5_mult_78_CARRYB_2__7_,
         u5_mult_78_CARRYB_2__8_, u5_mult_78_CARRYB_2__9_,
         u5_mult_78_CARRYB_3__0_, u5_mult_78_CARRYB_3__1_,
         u5_mult_78_CARRYB_3__2_, u5_mult_78_CARRYB_3__3_,
         u5_mult_78_CARRYB_3__4_, u5_mult_78_CARRYB_3__5_,
         u5_mult_78_CARRYB_3__6_, u5_mult_78_CARRYB_3__7_,
         u5_mult_78_CARRYB_3__8_, u5_mult_78_CARRYB_3__9_,
         u5_mult_78_CARRYB_4__0_, u5_mult_78_CARRYB_4__1_,
         u5_mult_78_CARRYB_4__2_, u5_mult_78_CARRYB_4__3_,
         u5_mult_78_CARRYB_4__4_, u5_mult_78_CARRYB_4__5_,
         u5_mult_78_CARRYB_4__6_, u5_mult_78_CARRYB_4__7_,
         u5_mult_78_CARRYB_4__8_, u5_mult_78_CARRYB_4__9_,
         u5_mult_78_CARRYB_5__0_, u5_mult_78_CARRYB_5__1_,
         u5_mult_78_CARRYB_5__2_, u5_mult_78_CARRYB_5__3_,
         u5_mult_78_CARRYB_5__4_, u5_mult_78_CARRYB_5__5_,
         u5_mult_78_CARRYB_5__6_, u5_mult_78_CARRYB_5__7_,
         u5_mult_78_CARRYB_5__8_, u5_mult_78_CARRYB_5__9_,
         u5_mult_78_CARRYB_6__0_, u5_mult_78_CARRYB_6__1_,
         u5_mult_78_CARRYB_6__2_, u5_mult_78_CARRYB_6__3_,
         u5_mult_78_CARRYB_6__4_, u5_mult_78_CARRYB_6__5_,
         u5_mult_78_CARRYB_6__6_, u5_mult_78_CARRYB_6__7_,
         u5_mult_78_CARRYB_6__8_, u5_mult_78_CARRYB_6__9_,
         u5_mult_78_CARRYB_7__0_, u5_mult_78_CARRYB_7__1_,
         u5_mult_78_CARRYB_7__2_, u5_mult_78_CARRYB_7__3_,
         u5_mult_78_CARRYB_7__4_, u5_mult_78_CARRYB_7__5_,
         u5_mult_78_CARRYB_7__6_, u5_mult_78_CARRYB_7__7_,
         u5_mult_78_CARRYB_7__8_, u5_mult_78_CARRYB_7__9_,
         u5_mult_78_CARRYB_8__0_, u5_mult_78_CARRYB_8__1_,
         u5_mult_78_CARRYB_8__2_, u5_mult_78_CARRYB_8__3_,
         u5_mult_78_CARRYB_8__4_, u5_mult_78_CARRYB_8__5_,
         u5_mult_78_CARRYB_8__6_, u5_mult_78_CARRYB_8__7_,
         u5_mult_78_CARRYB_8__8_, u5_mult_78_CARRYB_8__9_,
         u5_mult_78_CARRYB_9__0_, u5_mult_78_CARRYB_9__1_,
         u5_mult_78_CARRYB_9__2_, u5_mult_78_CARRYB_9__3_,
         u5_mult_78_CARRYB_9__4_, u5_mult_78_CARRYB_9__5_,
         u5_mult_78_CARRYB_9__6_, u5_mult_78_CARRYB_9__7_,
         u5_mult_78_CARRYB_9__8_, u5_mult_78_CARRYB_9__9_,
         u5_mult_78_CARRYB_10__0_, u5_mult_78_CARRYB_10__1_,
         u5_mult_78_CARRYB_10__2_, u5_mult_78_CARRYB_10__3_,
         u5_mult_78_CARRYB_10__4_, u5_mult_78_CARRYB_10__5_,
         u5_mult_78_CARRYB_10__6_, u5_mult_78_CARRYB_10__7_,
         u5_mult_78_CARRYB_10__8_, u5_mult_78_CARRYB_10__9_,
         u5_mult_78_ab_0__1_, u5_mult_78_ab_0__2_, u5_mult_78_ab_0__3_,
         u5_mult_78_ab_0__4_, u5_mult_78_ab_0__5_, u5_mult_78_ab_0__6_,
         u5_mult_78_ab_0__7_, u5_mult_78_ab_0__8_, u5_mult_78_ab_0__9_,
         u5_mult_78_ab_0__10_, u5_mult_78_ab_1__0_, u5_mult_78_ab_1__1_,
         u5_mult_78_ab_1__2_, u5_mult_78_ab_1__3_, u5_mult_78_ab_1__4_,
         u5_mult_78_ab_1__5_, u5_mult_78_ab_1__6_, u5_mult_78_ab_1__7_,
         u5_mult_78_ab_1__8_, u5_mult_78_ab_1__9_, u5_mult_78_ab_1__10_,
         u5_mult_78_ab_2__0_, u5_mult_78_ab_2__1_, u5_mult_78_ab_2__2_,
         u5_mult_78_ab_2__3_, u5_mult_78_ab_2__4_, u5_mult_78_ab_2__5_,
         u5_mult_78_ab_2__6_, u5_mult_78_ab_2__7_, u5_mult_78_ab_2__8_,
         u5_mult_78_ab_2__9_, u5_mult_78_ab_2__10_, u5_mult_78_ab_3__0_,
         u5_mult_78_ab_3__1_, u5_mult_78_ab_3__2_, u5_mult_78_ab_3__3_,
         u5_mult_78_ab_3__4_, u5_mult_78_ab_3__5_, u5_mult_78_ab_3__6_,
         u5_mult_78_ab_3__7_, u5_mult_78_ab_3__8_, u5_mult_78_ab_3__9_,
         u5_mult_78_ab_3__10_, u5_mult_78_ab_4__0_, u5_mult_78_ab_4__1_,
         u5_mult_78_ab_4__2_, u5_mult_78_ab_4__3_, u5_mult_78_ab_4__4_,
         u5_mult_78_ab_4__5_, u5_mult_78_ab_4__6_, u5_mult_78_ab_4__7_,
         u5_mult_78_ab_4__8_, u5_mult_78_ab_4__9_, u5_mult_78_ab_4__10_,
         u5_mult_78_ab_5__0_, u5_mult_78_ab_5__1_, u5_mult_78_ab_5__2_,
         u5_mult_78_ab_5__3_, u5_mult_78_ab_5__4_, u5_mult_78_ab_5__5_,
         u5_mult_78_ab_5__6_, u5_mult_78_ab_5__7_, u5_mult_78_ab_5__8_,
         u5_mult_78_ab_5__9_, u5_mult_78_ab_5__10_, u5_mult_78_ab_6__0_,
         u5_mult_78_ab_6__1_, u5_mult_78_ab_6__2_, u5_mult_78_ab_6__3_,
         u5_mult_78_ab_6__4_, u5_mult_78_ab_6__5_, u5_mult_78_ab_6__6_,
         u5_mult_78_ab_6__7_, u5_mult_78_ab_6__8_, u5_mult_78_ab_6__9_,
         u5_mult_78_ab_6__10_, u5_mult_78_ab_7__0_, u5_mult_78_ab_7__1_,
         u5_mult_78_ab_7__2_, u5_mult_78_ab_7__3_, u5_mult_78_ab_7__4_,
         u5_mult_78_ab_7__5_, u5_mult_78_ab_7__6_, u5_mult_78_ab_7__7_,
         u5_mult_78_ab_7__8_, u5_mult_78_ab_7__9_, u5_mult_78_ab_7__10_,
         u5_mult_78_ab_8__0_, u5_mult_78_ab_8__1_, u5_mult_78_ab_8__2_,
         u5_mult_78_ab_8__3_, u5_mult_78_ab_8__4_, u5_mult_78_ab_8__5_,
         u5_mult_78_ab_8__6_, u5_mult_78_ab_8__7_, u5_mult_78_ab_8__8_,
         u5_mult_78_ab_8__9_, u5_mult_78_ab_8__10_, u5_mult_78_ab_9__0_,
         u5_mult_78_ab_9__1_, u5_mult_78_ab_9__2_, u5_mult_78_ab_9__3_,
         u5_mult_78_ab_9__4_, u5_mult_78_ab_9__5_, u5_mult_78_ab_9__6_,
         u5_mult_78_ab_9__7_, u5_mult_78_ab_9__8_, u5_mult_78_ab_9__9_,
         u5_mult_78_ab_9__10_, u5_mult_78_ab_10__0_, u5_mult_78_ab_10__1_,
         u5_mult_78_ab_10__2_, u5_mult_78_ab_10__3_, u5_mult_78_ab_10__4_,
         u5_mult_78_ab_10__5_, u5_mult_78_ab_10__6_, u5_mult_78_ab_10__7_,
         u5_mult_78_ab_10__8_, u5_mult_78_ab_10__9_, u5_mult_78_ab_10__10_,
         u5_mult_78_FS_1_n44, u5_mult_78_FS_1_n43, u5_mult_78_FS_1_n42,
         u5_mult_78_FS_1_n41, u5_mult_78_FS_1_n40, u5_mult_78_FS_1_n39,
         u5_mult_78_FS_1_n38, u5_mult_78_FS_1_n37, u5_mult_78_FS_1_n36,
         u5_mult_78_FS_1_n35, u5_mult_78_FS_1_n34, u5_mult_78_FS_1_n33,
         u5_mult_78_FS_1_n32, u5_mult_78_FS_1_n31, u5_mult_78_FS_1_n30,
         u5_mult_78_FS_1_n29, u5_mult_78_FS_1_n28, u5_mult_78_FS_1_n27,
         u5_mult_78_FS_1_n26, u5_mult_78_FS_1_n25, u5_mult_78_FS_1_n24,
         u5_mult_78_FS_1_n23, u5_mult_78_FS_1_n22, u5_mult_78_FS_1_n21,
         u5_mult_78_FS_1_n20, u5_mult_78_FS_1_n19, u5_mult_78_FS_1_n18,
         u5_mult_78_FS_1_n17, u5_mult_78_FS_1_n16, u5_mult_78_FS_1_n15,
         u5_mult_78_FS_1_n14, u5_mult_78_FS_1_n13, u5_mult_78_FS_1_n12,
         u5_mult_78_FS_1_n11, u5_mult_78_FS_1_n10, u5_mult_78_FS_1_n9,
         u5_mult_78_FS_1_n8, u5_mult_78_FS_1_n7, u5_mult_78_FS_1_n6,
         u5_mult_78_FS_1_n5, u5_mult_78_FS_1_n4, u5_mult_78_FS_1_n3,
         u5_mult_78_FS_1_n1;
  wire   [15:10] opa_r;
  wire   [15:10] opb_r;
  wire   [1:0] rmode_r1;
  wire   [1:0] rmode_r2;
  wire   [1:0] rmode_r3;
  wire   [2:0] fpu_op_r1;
  wire   [2:0] fpu_op_r2;
  wire   [13:0] fracta;
  wire   [13:0] fractb;
  wire   [9:0] fracta_mul;
  wire   [1:0] exp_ovf;
  wire   [2:0] underflow_fmul_d;
  wire   [14:1] fract_out_q;
  wire   [21:2] prod;
  wire   [22:0] quo;
  wire   [22:0] remainder;
  wire   [3:0] div_opa_ldz_r1;
  wire   [3:0] div_opa_ldz_r2;
  wire   [4:1] exp_r;
  wire   [11:4] opa_r1;
  wire   [21:8] fract_denorm;
  wire   [2:1] underflow_fmul_r;
  wire   [13:0] u1_fractb_s;
  wire   [13:0] u1_fracta_s;
  wire   [4:0] u1_exp_diff2;
  wire   [4:3] u1_exp_small;
  wire   [2:0] u2_underflow_d;
  wire   [21:0] u5_prod1;
  wire   [23:0] u6_remainder;
  wire   [23:0] u6_quo1;
  wire   [4:0] u4_div_exp3;
  wire   [4:0] u4_div_exp2;
  wire   [27:23] u4_exp_f2i_1;
  wire   [4:0] u4_exp_fix_divb;
  wire   [4:0] u4_exp_fix_diva;
  wire   [4:0] u4_exp_out1_mi1;
  wire   [4:1] u4_exp_out_mi1;
  wire   [2:0] u4_shift_left;
  wire   [4:0] u4_shift_right;
  wire   [4:0] u4_div_shft4;
  wire   [4:0] u4_div_shft2;
  wire   [5:0] u4_div_scht1a;
  wire   [4:1] u4_sub_470_carry;
  wire   [4:2] u4_add_461_carry;
  wire   [4:3] u4_add_407_carry;
  wire   [4:1] u4_sub_409_carry;
  wire   [4:1] u4_add_408_carry;
  wire   [4:2] u4_sub_478_carry;
  wire   [4:1] u4_sub_493_carry;
  wire   [4:1] u4_add_486_carry;
  wire   [4:2] u4_add_463_carry;
  wire   [4:1] u4_add_491_carry;
  wire   [5:1] u4_sub_406_carry;
  wire   [4:2] u2_add_115_carry;
  wire   [4:2] u2_add_113_carry;
  wire   [4:1] u2_add_110_carry;
  wire   [5:1] u2_sub_110_carry;
  wire   [4:1] sub_1_root_u1_sub_128_aco_carry;
  wire   [20:8] sub_434_3_carry;
  wire   [10:2] sub_434_b0_carry;
  wire   [4:2] u4_sub_488_carry;
  wire   [4:1] sub_0_root_sub_0_root_u4_sub_469_carry;
  wire   [4:1] add_0_root_sub_0_root_u4_add_494_carry;
  wire   [4:1] sub_1_root_sub_0_root_u4_add_494_carry;
  wire   [9:2] u4_add_393_carry;
  wire   [5:1] u4_sub_467_carry;
  wire   [14:1] u3_sub_59_carry;
  wire   [13:2] u3_add_59_carry;

  OR2_X2 u4_C1739 ( .A1(u4_N655), .A2(u4_exp_out_0_), .ZN(u4_N656) );
  OR2_X2 u4_C1740 ( .A1(u4_N654), .A2(u4_exp_out_1_), .ZN(u4_N655) );
  OR2_X2 u4_C1741 ( .A1(u4_N653), .A2(u4_exp_out_2_), .ZN(u4_N654) );
  OR2_X2 u4_C1742 ( .A1(u4_exp_out_4_), .A2(u4_exp_out_3_), .ZN(u4_N653) );
  OR2_X2 u4_C1935 ( .A1(u4_shift_right[4]), .A2(u4_shift_right[3]), .ZN(
        u4_N386) );
  OR2_X2 u4_C2104 ( .A1(u4_N796), .A2(u4_N797), .ZN(u4_N798) );
  AND2_X2 u4_C2106 ( .A1(u4_exp_out_4_), .A2(1'b1), .ZN(u4_N797) );
  AOI22_X2 U16 ( .A1(u4_div_exp3[1]), .A2(n842), .B1(n848), .B2(
        u4_sub_465_A_1_), .ZN(n845) );
  OAI211_X2 U18 ( .C1(n850), .C2(n831), .A(n851), .B(n852), .ZN(u4_exp_out_2_)
         );
  OAI221_X2 U100 ( .B1(u4_N581), .B2(n872), .C1(n888), .C2(n1631), .A(n889), 
        .ZN(u4_shift_right[0]) );
  DFF_X2 opa_r_reg_15_ ( .D(opa[15]), .CK(clk), .Q(opa_r[15]), .QN(n1594) );
  DFF_X2 opa_r_reg_14_ ( .D(opa[14]), .CK(clk), .Q(opa_r[14]), .QN(n1577) );
  DFF_X2 opa_r_reg_13_ ( .D(opa[13]), .CK(clk), .Q(opa_r[13]), .QN(n1579) );
  DFF_X2 opa_r_reg_12_ ( .D(opa[12]), .CK(clk), .Q(opa_r[12]), .QN(n1547) );
  DFF_X2 opa_r_reg_11_ ( .D(opa[11]), .CK(clk), .Q(opa_r[11]), .QN(n1578) );
  DFF_X2 opa_r_reg_10_ ( .D(opa[10]), .CK(clk), .Q(opa_r[10]), .QN(n1580) );
  DFF_X2 opa_r_reg_9_ ( .D(opa[9]), .CK(clk), .Q(fracta_mul[9]), .QN(n1856) );
  DFF_X2 opa_r_reg_8_ ( .D(opa[8]), .CK(clk), .Q(fracta_mul[8]), .QN(n1855) );
  DFF_X2 opa_r_reg_7_ ( .D(opa[7]), .CK(clk), .Q(fracta_mul[7]), .QN(n1854) );
  DFF_X2 opa_r_reg_6_ ( .D(opa[6]), .CK(clk), .Q(fracta_mul[6]), .QN(n1853) );
  DFF_X2 opa_r_reg_5_ ( .D(opa[5]), .CK(clk), .Q(fracta_mul[5]), .QN(n1852) );
  DFF_X2 opa_r_reg_4_ ( .D(opa[4]), .CK(clk), .Q(fracta_mul[4]), .QN(n1851) );
  DFF_X2 opa_r_reg_3_ ( .D(opa[3]), .CK(clk), .Q(fracta_mul[3]), .QN(n1850) );
  DFF_X2 opa_r_reg_2_ ( .D(opa[2]), .CK(clk), .Q(fracta_mul[2]), .QN(n1849) );
  DFF_X2 opa_r_reg_1_ ( .D(opa[1]), .CK(clk), .Q(fracta_mul[1]), .QN(n1848) );
  DFF_X2 opa_r_reg_0_ ( .D(opa[0]), .CK(clk), .Q(fracta_mul[0]), .QN(n1847) );
  DFF_X2 opb_r_reg_15_ ( .D(opb[15]), .CK(clk), .Q(opb_r[15]), .QN(n1554) );
  DFF_X2 opb_r_reg_14_ ( .D(opb[14]), .CK(clk), .Q(opb_r[14]), .QN(n1582) );
  DFF_X2 opb_r_reg_13_ ( .D(opb[13]), .CK(clk), .Q(opb_r[13]), .QN(n1583) );
  DFF_X2 opb_r_reg_12_ ( .D(opb[12]), .CK(clk), .Q(opb_r[12]), .QN(n1584) );
  DFF_X2 opb_r_reg_11_ ( .D(opb[11]), .CK(clk), .Q(opb_r[11]), .QN(n1587) );
  DFF_X2 opb_r_reg_10_ ( .D(opb[10]), .CK(clk), .Q(opb_r[10]), .QN(n1588) );
  DFF_X2 opb_r_reg_9_ ( .D(opb[9]), .CK(clk), .Q(u6_N9), .QN(n1846) );
  DFF_X2 opb_r_reg_8_ ( .D(opb[8]), .CK(clk), .Q(u6_N8) );
  DFF_X2 opb_r_reg_7_ ( .D(opb[7]), .CK(clk), .Q(u6_N7), .QN(n1845) );
  DFF_X2 opb_r_reg_6_ ( .D(opb[6]), .CK(clk), .Q(u6_N6), .QN(n1844) );
  DFF_X2 opb_r_reg_5_ ( .D(opb[5]), .CK(clk), .Q(u6_N5), .QN(n1843) );
  DFF_X2 opb_r_reg_4_ ( .D(opb[4]), .CK(clk), .Q(u6_N4), .QN(n1842) );
  DFF_X2 opb_r_reg_3_ ( .D(opb[3]), .CK(clk), .Q(u6_N3), .QN(n1841) );
  DFF_X2 opb_r_reg_2_ ( .D(opb[2]), .CK(clk), .Q(u6_N2), .QN(n1840) );
  DFF_X2 opb_r_reg_1_ ( .D(opb[1]), .CK(clk), .Q(u6_N1), .QN(n1839) );
  DFF_X2 opb_r_reg_0_ ( .D(opb[0]), .CK(clk), .Q(u6_N0), .QN(n1838) );
  DFF_X2 rmode_r1_reg_1_ ( .D(rmode[1]), .CK(clk), .Q(rmode_r1[1]) );
  DFF_X2 rmode_r1_reg_0_ ( .D(rmode[0]), .CK(clk), .Q(rmode_r1[0]) );
  DFF_X2 rmode_r2_reg_1_ ( .D(rmode_r1[1]), .CK(clk), .Q(rmode_r2[1]) );
  DFF_X2 rmode_r2_reg_0_ ( .D(rmode_r1[0]), .CK(clk), .Q(rmode_r2[0]) );
  DFF_X2 rmode_r3_reg_1_ ( .D(rmode_r2[1]), .CK(clk), .Q(rmode_r3[1]), .QN(
        n1548) );
  DFF_X2 rmode_r3_reg_0_ ( .D(rmode_r2[0]), .CK(clk), .Q(rmode_r3[0]), .QN(
        n1576) );
  DFF_X2 fpu_op_r1_reg_2_ ( .D(fpu_op[2]), .CK(clk), .Q(fpu_op_r1[2]), .QN(
        n1837) );
  DFF_X2 fpu_op_r1_reg_1_ ( .D(fpu_op[1]), .CK(clk), .Q(fpu_op_r1[1]) );
  DFF_X2 fpu_op_r1_reg_0_ ( .D(fpu_op[0]), .CK(clk), .Q(fpu_op_r1[0]), .QN(
        n2702) );
  DFF_X2 fpu_op_r2_reg_2_ ( .D(fpu_op_r1[2]), .CK(clk), .Q(fpu_op_r2[2]), .QN(
        n1836) );
  DFF_X2 fpu_op_r2_reg_1_ ( .D(fpu_op_r1[1]), .CK(clk), .Q(fpu_op_r2[1]), .QN(
        n1835) );
  DFF_X2 fpu_op_r2_reg_0_ ( .D(fpu_op_r1[0]), .CK(clk), .Q(fpu_op_r2[0]), .QN(
        n1834) );
  DFF_X2 fpu_op_r3_reg_2_ ( .D(fpu_op_r2[2]), .CK(clk), .Q(n1560), .QN(n1833)
         );
  DFF_X2 fpu_op_r3_reg_1_ ( .D(fpu_op_r2[1]), .CK(clk), .QN(n1832) );
  DFF_X2 fpu_op_r3_reg_0_ ( .D(fpu_op_r2[0]), .CK(clk), .Q(n1536), .QN(n1831)
         );
  DFF_X2 div_opa_ldz_r1_reg_3_ ( .D(N34), .CK(clk), .Q(div_opa_ldz_r1[3]) );
  DFF_X2 div_opa_ldz_r1_reg_2_ ( .D(N44), .CK(clk), .Q(div_opa_ldz_r1[2]) );
  DFF_X2 div_opa_ldz_r1_reg_1_ ( .D(N56), .CK(clk), .Q(div_opa_ldz_r1[1]) );
  DFF_X2 div_opa_ldz_r1_reg_0_ ( .D(N65), .CK(clk), .Q(div_opa_ldz_r1[0]) );
  DFF_X2 div_opa_ldz_r2_reg_3_ ( .D(div_opa_ldz_r1[3]), .CK(clk), .Q(
        div_opa_ldz_r2[3]), .QN(n2475) );
  DFF_X2 div_opa_ldz_r2_reg_2_ ( .D(div_opa_ldz_r1[2]), .CK(clk), .Q(
        div_opa_ldz_r2[2]), .QN(n1830) );
  DFF_X2 div_opa_ldz_r2_reg_1_ ( .D(div_opa_ldz_r1[1]), .CK(clk), .Q(
        div_opa_ldz_r2[1]), .QN(n1829) );
  DFF_X2 div_opa_ldz_r2_reg_0_ ( .D(div_opa_ldz_r1[0]), .CK(clk), .Q(
        div_opa_ldz_r2[0]), .QN(n1828) );
  DFF_X2 opa_r1_reg_14_ ( .D(opa_r[14]), .CK(clk), .QN(n1620) );
  DFF_X2 opa_r1_reg_13_ ( .D(opa_r[13]), .CK(clk), .QN(n1621) );
  DFF_X2 opa_r1_reg_12_ ( .D(opa_r[12]), .CK(clk), .QN(n1622) );
  DFF_X2 opa_r1_reg_11_ ( .D(opa_r[11]), .CK(clk), .Q(opa_r1[11]), .QN(n1618)
         );
  DFF_X2 opa_r1_reg_10_ ( .D(opa_r[10]), .CK(clk), .Q(opa_r1[10]), .QN(n1619)
         );
  DFF_X2 opa_r1_reg_9_ ( .D(fracta_mul[9]), .CK(clk), .QN(n1614) );
  DFF_X2 opa_r1_reg_8_ ( .D(fracta_mul[8]), .CK(clk), .QN(n1615) );
  DFF_X2 opa_r1_reg_7_ ( .D(fracta_mul[7]), .CK(clk), .QN(n1616) );
  DFF_X2 opa_r1_reg_6_ ( .D(fracta_mul[6]), .CK(clk), .QN(n1617) );
  DFF_X2 opa_r1_reg_5_ ( .D(fracta_mul[5]), .CK(clk), .Q(opa_r1[5]), .QN(n1612) );
  DFF_X2 opa_r1_reg_4_ ( .D(fracta_mul[4]), .CK(clk), .Q(opa_r1[4]), .QN(n1613) );
  DFF_X2 opa_r1_reg_3_ ( .D(fracta_mul[3]), .CK(clk), .QN(n1589) );
  DFF_X2 opa_r1_reg_2_ ( .D(fracta_mul[2]), .CK(clk), .QN(n1590) );
  DFF_X2 opa_r1_reg_1_ ( .D(fracta_mul[1]), .CK(clk), .QN(n1591) );
  DFF_X2 opa_r1_reg_0_ ( .D(fracta_mul[0]), .CK(clk), .Q(N106), .QN(n1599) );
  DFF_X2 opas_r1_reg ( .D(opa_r[15]), .CK(clk), .Q(opas_r1) );
  DFF_X2 opas_r2_reg ( .D(opas_r1), .CK(clk), .Q(opas_r2), .QN(n1573) );
  DFF_X2 u0_fractb_00_reg ( .D(n2701), .CK(clk), .QN(n1827) );
  DFF_X2 u0_fracta_00_reg ( .D(n2699), .CK(clk), .QN(n1826) );
  DFF_X2 u0_expb_00_reg ( .D(n1523), .CK(clk), .Q(u0_expb_00), .QN(n1825) );
  DFF_X2 u0_opb_dn_reg ( .D(u0_expb_00), .CK(clk), .Q(opb_dn), .QN(n1538) );
  DFF_X2 u0_opb_00_reg ( .D(u0_N17), .CK(clk), .Q(opb_00), .QN(n1553) );
  DFF_X2 u0_expa_00_reg ( .D(n1522), .CK(clk), .Q(u0_expa_00), .QN(n1824) );
  DFF_X2 u0_opa_dn_reg ( .D(u0_expa_00), .CK(clk), .Q(opa_dn), .QN(n1574) );
  DFF_X2 u0_opa_00_reg ( .D(u0_N16), .CK(clk), .Q(opa_00), .QN(n1592) );
  DFF_X2 u0_opb_nan_reg ( .D(u0_N11), .CK(clk), .Q(opb_nan), .QN(n1610) );
  DFF_X2 u0_opa_nan_reg ( .D(u0_N10), .CK(clk), .Q(opa_nan), .QN(n1600) );
  DFF_X2 opa_nan_r_reg ( .D(N291), .CK(clk), .QN(n1823) );
  DFF_X2 u0_snan_r_b_reg ( .D(u0_N5), .CK(clk), .QN(n1822) );
  DFF_X2 u0_qnan_r_b_reg ( .D(u6_N9), .CK(clk), .QN(n1821) );
  DFF_X2 u0_snan_r_a_reg ( .D(u0_N4), .CK(clk), .QN(n1820) );
  DFF_X2 u0_qnan_r_a_reg ( .D(fracta_mul[9]), .CK(clk), .QN(n1819) );
  DFF_X2 u0_infb_f_r_reg ( .D(n2701), .CK(clk), .Q(u0_infb_f_r) );
  DFF_X2 u0_infa_f_r_reg ( .D(n2699), .CK(clk), .Q(u0_infa_f_r) );
  DFF_X2 u0_expb_ff_reg ( .D(n2700), .CK(clk), .Q(u0_expb_ff), .QN(n1596) );
  DFF_X2 u0_opb_inf_reg ( .D(n2714), .CK(clk), .Q(opb_inf), .QN(n1549) );
  DFF_X2 u0_expa_ff_reg ( .D(n2697), .CK(clk), .Q(u0_expa_ff), .QN(n1555) );
  DFF_X2 u0_snan_reg ( .D(n2712), .CK(clk), .Q(snan_d), .QN(n1818) );
  DFF_X2 snan_reg ( .D(snan_d), .CK(clk), .Q(snan) );
  DFF_X2 u0_qnan_reg ( .D(n2713), .CK(clk), .QN(n1817) );
  DFF_X2 u0_opa_inf_reg ( .D(n2715), .CK(clk), .Q(opa_inf), .QN(n1595) );
  DFF_X2 div_by_zero_reg ( .D(N292), .CK(clk), .Q(div_by_zero) );
  DFF_X2 u0_inf_reg ( .D(u0_N7), .CK(clk), .Q(n1597), .QN(n1816) );
  DFF_X2 u0_ind_reg ( .D(u0_N6), .CK(clk), .Q(n1598) );
  DFF_X2 u1_fasu_op_reg ( .D(n2684), .CK(clk), .Q(fasu_op), .QN(n1815) );
  DFF_X2 fasu_op_r1_reg ( .D(fasu_op), .CK(clk), .Q(fasu_op_r1) );
  DFF_X2 fasu_op_r2_reg ( .D(fasu_op_r1), .CK(clk), .QN(n1814) );
  DFF_X2 qnan_reg ( .D(N283), .CK(clk), .Q(qnan) );
  DFF_X2 u1_fracta_eq_fractb_reg ( .D(u1_N124), .CK(clk), .Q(
        u1_fracta_eq_fractb) );
  DFF_X2 u1_fracta_lt_fractb_reg ( .D(u1_N123), .CK(clk), .Q(
        u1_fracta_lt_fractb), .QN(n1609) );
  DFF_X2 u1_add_r_reg ( .D(n2702), .CK(clk), .Q(u1_add_r) );
  DFF_X2 u1_signb_r_reg ( .D(opb_r[15]), .CK(clk), .QN(n1593) );
  DFF_X2 u1_signa_r_reg ( .D(opa_r[15]), .CK(clk), .Q(u1_signa_r), .QN(n1608)
         );
  DFF_X2 u1_result_zero_sign_reg ( .D(u1_N122), .CK(clk), .Q(
        result_zero_sign_d) );
  DFF_X2 u1_nan_sign_reg ( .D(u1_N133), .CK(clk), .Q(nan_sign_d) );
  DFF_X2 u1_sign_reg ( .D(u1_sign_d), .CK(clk), .Q(sign_fasu) );
  DFF_X2 sign_fasu_r_reg ( .D(sign_fasu), .CK(clk), .Q(sign_fasu_r) );
  DFF_X2 u1_fractb_out_reg_0_ ( .D(u1_fractb_s[0]), .CK(clk), .Q(fractb[0]) );
  DFF_X2 u1_fractb_out_reg_1_ ( .D(u1_fractb_s[1]), .CK(clk), .Q(fractb[1]) );
  DFF_X2 u1_fractb_out_reg_2_ ( .D(u1_fractb_s[2]), .CK(clk), .Q(fractb[2]) );
  DFF_X2 u1_fractb_out_reg_3_ ( .D(u1_fractb_s[3]), .CK(clk), .Q(fractb[3]) );
  DFF_X2 u1_fractb_out_reg_4_ ( .D(u1_fractb_s[4]), .CK(clk), .Q(fractb[4]) );
  DFF_X2 u1_fractb_out_reg_5_ ( .D(u1_fractb_s[5]), .CK(clk), .Q(fractb[5]) );
  DFF_X2 u1_fractb_out_reg_6_ ( .D(u1_fractb_s[6]), .CK(clk), .Q(fractb[6]) );
  DFF_X2 u1_fractb_out_reg_7_ ( .D(u1_fractb_s[7]), .CK(clk), .Q(fractb[7]) );
  DFF_X2 u1_fractb_out_reg_8_ ( .D(u1_fractb_s[8]), .CK(clk), .Q(fractb[8]) );
  DFF_X2 u1_fractb_out_reg_9_ ( .D(u1_fractb_s[9]), .CK(clk), .Q(fractb[9]) );
  DFF_X2 u1_fractb_out_reg_10_ ( .D(u1_fractb_s[10]), .CK(clk), .Q(fractb[10])
         );
  DFF_X2 u1_fractb_out_reg_11_ ( .D(u1_fractb_s[11]), .CK(clk), .Q(fractb[11])
         );
  DFF_X2 u1_fractb_out_reg_12_ ( .D(u1_fractb_s[12]), .CK(clk), .Q(fractb[12])
         );
  DFF_X2 u1_fractb_out_reg_13_ ( .D(u1_fractb_s[13]), .CK(clk), .Q(fractb[13])
         );
  DFF_X2 u1_fracta_out_reg_0_ ( .D(u1_fracta_s[0]), .CK(clk), .Q(fracta[0]) );
  DFF_X2 u1_fracta_out_reg_1_ ( .D(u1_fracta_s[1]), .CK(clk), .Q(fracta[1]) );
  DFF_X2 u1_fracta_out_reg_2_ ( .D(u1_fracta_s[2]), .CK(clk), .Q(fracta[2]) );
  DFF_X2 u1_fracta_out_reg_3_ ( .D(u1_fracta_s[3]), .CK(clk), .Q(fracta[3]) );
  DFF_X2 u1_fracta_out_reg_4_ ( .D(u1_fracta_s[4]), .CK(clk), .Q(fracta[4]) );
  DFF_X2 u1_fracta_out_reg_5_ ( .D(u1_fracta_s[5]), .CK(clk), .Q(fracta[5]) );
  DFF_X2 u1_fracta_out_reg_6_ ( .D(u1_fracta_s[6]), .CK(clk), .Q(fracta[6]) );
  DFF_X2 u1_fracta_out_reg_7_ ( .D(u1_fracta_s[7]), .CK(clk), .Q(fracta[7]) );
  DFF_X2 u1_fracta_out_reg_8_ ( .D(u1_fracta_s[8]), .CK(clk), .Q(fracta[8]) );
  DFF_X2 u1_fracta_out_reg_9_ ( .D(u1_fracta_s[9]), .CK(clk), .Q(fracta[9]) );
  DFF_X2 u1_fracta_out_reg_10_ ( .D(u1_fracta_s[10]), .CK(clk), .Q(fracta[10])
         );
  DFF_X2 u1_fracta_out_reg_11_ ( .D(u1_fracta_s[11]), .CK(clk), .Q(fracta[11])
         );
  DFF_X2 u1_fracta_out_reg_12_ ( .D(u1_fracta_s[12]), .CK(clk), .Q(fracta[12])
         );
  DFF_X2 u1_fracta_out_reg_13_ ( .D(u1_fracta_s[13]), .CK(clk), .Q(fracta[13])
         );
  DFF_X2 fract_out_q_reg_0_ ( .D(n2683), .CK(clk), .QN(n1813) );
  DFF_X2 fract_out_q_reg_1_ ( .D(n2682), .CK(clk), .Q(fract_out_q[1]) );
  DFF_X2 fract_out_q_reg_2_ ( .D(n2681), .CK(clk), .Q(fract_out_q[2]) );
  DFF_X2 fract_out_q_reg_3_ ( .D(n2680), .CK(clk), .Q(fract_out_q[3]) );
  DFF_X2 fract_out_q_reg_4_ ( .D(n2679), .CK(clk), .Q(fract_out_q[4]) );
  DFF_X2 fract_out_q_reg_5_ ( .D(n2678), .CK(clk), .Q(fract_out_q[5]) );
  DFF_X2 fract_out_q_reg_6_ ( .D(n2677), .CK(clk), .Q(fract_out_q[6]) );
  DFF_X2 fract_out_q_reg_7_ ( .D(n2676), .CK(clk), .Q(fract_out_q[7]) );
  DFF_X2 fract_out_q_reg_8_ ( .D(n2675), .CK(clk), .Q(fract_out_q[8]) );
  DFF_X2 fract_out_q_reg_9_ ( .D(n2674), .CK(clk), .Q(fract_out_q[9]) );
  DFF_X2 fract_out_q_reg_10_ ( .D(n2673), .CK(clk), .Q(fract_out_q[10]) );
  DFF_X2 fract_out_q_reg_11_ ( .D(n2672), .CK(clk), .Q(fract_out_q[11]) );
  DFF_X2 fract_out_q_reg_12_ ( .D(n2671), .CK(clk), .Q(fract_out_q[12]) );
  DFF_X2 fract_out_q_reg_13_ ( .D(n2670), .CK(clk), .Q(fract_out_q[13]) );
  DFF_X2 fract_out_q_reg_14_ ( .D(n2669), .CK(clk), .Q(fract_out_q[14]) );
  DFF_X2 u1_exp_dn_out_reg_0_ ( .D(u1_N35), .CK(clk), .QN(n1812) );
  DFF_X2 u1_exp_dn_out_reg_1_ ( .D(u1_N36), .CK(clk), .QN(n1811) );
  DFF_X2 u1_exp_dn_out_reg_2_ ( .D(u1_N37), .CK(clk), .QN(n1810) );
  DFF_X2 u1_exp_dn_out_reg_3_ ( .D(u1_N38), .CK(clk), .QN(n1809) );
  DFF_X2 u1_exp_dn_out_reg_4_ ( .D(u1_N39), .CK(clk), .QN(n1808) );
  DFF_X2 u2_sign_exe_reg ( .D(u2_N73), .CK(clk), .Q(sign_exe) );
  DFF_X2 sign_exe_r_reg ( .D(sign_exe), .CK(clk), .Q(sign_exe_r), .QN(n1611)
         );
  DFF_X2 u2_sign_reg ( .D(u2_sign_d), .CK(clk), .Q(sign_mul) );
  DFF_X2 sign_mul_r_reg ( .D(sign_mul), .CK(clk), .Q(sign_mul_r) );
  DFF_X2 sign_reg ( .D(N216), .CK(clk), .Q(sign), .QN(n1581) );
  DFF_X2 fract_i2f_reg_21_ ( .D(N196), .CK(clk), .QN(n1807) );
  DFF_X2 fract_i2f_reg_20_ ( .D(N195), .CK(clk), .QN(n1806) );
  DFF_X2 fract_i2f_reg_19_ ( .D(N194), .CK(clk), .QN(n1805) );
  DFF_X2 fract_i2f_reg_18_ ( .D(N193), .CK(clk), .QN(n1804) );
  DFF_X2 fract_i2f_reg_17_ ( .D(N192), .CK(clk), .QN(n1803) );
  DFF_X2 fract_i2f_reg_16_ ( .D(N191), .CK(clk), .QN(n1802) );
  DFF_X2 fract_i2f_reg_15_ ( .D(N190), .CK(clk), .QN(n1801) );
  DFF_X2 fract_i2f_reg_14_ ( .D(N189), .CK(clk), .QN(n1800) );
  DFF_X2 fract_i2f_reg_13_ ( .D(N188), .CK(clk), .QN(n1799) );
  DFF_X2 fract_i2f_reg_12_ ( .D(N187), .CK(clk), .QN(n1798) );
  DFF_X2 fract_i2f_reg_11_ ( .D(N186), .CK(clk), .QN(n1797) );
  DFF_X2 fract_i2f_reg_10_ ( .D(N185), .CK(clk), .QN(n1796) );
  DFF_X2 fract_i2f_reg_9_ ( .D(N184), .CK(clk), .QN(n1795) );
  DFF_X2 fract_i2f_reg_8_ ( .D(N183), .CK(clk), .QN(n1794) );
  DFF_X2 fract_i2f_reg_7_ ( .D(N182), .CK(clk), .Q(fract_i2f_7_) );
  DFF_X2 fract_i2f_reg_6_ ( .D(N181), .CK(clk), .Q(n1540) );
  DFF_X2 fract_i2f_reg_5_ ( .D(N180), .CK(clk), .Q(n1541) );
  DFF_X2 fract_i2f_reg_4_ ( .D(N179), .CK(clk), .Q(n1542) );
  DFF_X2 fract_i2f_reg_3_ ( .D(n2666), .CK(clk), .Q(n1543) );
  DFF_X2 fract_i2f_reg_2_ ( .D(n2667), .CK(clk), .Q(n1539) );
  DFF_X2 fract_i2f_reg_1_ ( .D(n2668), .CK(clk), .QN(n1793) );
  DFF_X2 fract_i2f_reg_0_ ( .D(n2703), .CK(clk), .QN(n1792) );
  DFF_X2 u2_inf_reg ( .D(u2_N66), .CK(clk), .Q(inf_mul) );
  DFF_X2 inf_mul_r_reg ( .D(inf_mul), .CK(clk), .Q(n1604), .QN(n1791) );
  DFF_X2 u2_underflow_reg_0_ ( .D(u2_underflow_d[0]), .CK(clk), .Q(
        underflow_fmul_d[0]) );
  DFF_X2 underflow_fmul_r_reg_0_ ( .D(underflow_fmul_d[0]), .CK(clk), .QN(
        n1790) );
  DFF_X2 u2_underflow_reg_1_ ( .D(u2_underflow_d[1]), .CK(clk), .Q(
        underflow_fmul_d[1]) );
  DFF_X2 underflow_fmul_r_reg_1_ ( .D(underflow_fmul_d[1]), .CK(clk), .Q(
        underflow_fmul_r[1]) );
  DFF_X2 u2_underflow_reg_2_ ( .D(u2_underflow_d[2]), .CK(clk), .Q(
        underflow_fmul_d[2]) );
  DFF_X2 underflow_fmul_r_reg_2_ ( .D(underflow_fmul_d[2]), .CK(clk), .Q(
        underflow_fmul_r[2]) );
  DFF_X2 u2_exp_ovf_reg_0_ ( .D(u2_exp_ovf_d_0_), .CK(clk), .Q(exp_ovf[0]) );
  DFF_X2 exp_ovf_r_reg_0_ ( .D(exp_ovf[0]), .CK(clk), .Q(n1546), .QN(n1789) );
  DFF_X2 u2_exp_ovf_reg_1_ ( .D(u2_exp_ovf_d_1_), .CK(clk), .Q(exp_ovf[1]) );
  DFF_X2 exp_ovf_r_reg_1_ ( .D(exp_ovf[1]), .CK(clk), .Q(n1575), .QN(n1788) );
  DFF_X2 u2_exp_out_reg_0_ ( .D(u2_N40), .CK(clk), .QN(n1787) );
  DFF_X2 exp_r_reg_0_ ( .D(N96), .CK(clk), .Q(u4_div_shft2[0]), .QN(n1786) );
  DFF_X2 u2_exp_out_reg_1_ ( .D(u2_N41), .CK(clk), .QN(n1785) );
  DFF_X2 exp_r_reg_1_ ( .D(N97), .CK(clk), .Q(exp_r[1]), .QN(n1784) );
  DFF_X2 u2_exp_out_reg_2_ ( .D(u2_N42), .CK(clk), .QN(n1783) );
  DFF_X2 exp_r_reg_2_ ( .D(N98), .CK(clk), .Q(exp_r[2]), .QN(n1782) );
  DFF_X2 u2_exp_out_reg_3_ ( .D(u2_N43), .CK(clk), .QN(n1781) );
  DFF_X2 exp_r_reg_3_ ( .D(N99), .CK(clk), .Q(n1533), .QN(n1780) );
  DFF_X2 u2_exp_out_reg_4_ ( .D(u2_N44), .CK(clk), .QN(n1779) );
  DFF_X2 inf_mul2_reg ( .D(N296), .CK(clk), .QN(n1778) );
  DFF_X2 exp_r_reg_4_ ( .D(N100), .CK(clk), .Q(exp_r[4]), .QN(n1777) );
  DFF_X2 u5_prod1_reg_0_ ( .D(u5_N0), .CK(clk), .Q(u5_prod1[0]) );
  DFF_X2 u5_prod_reg_0_ ( .D(u5_prod1[0]), .CK(clk), .QN(n1544) );
  DFF_X2 u5_prod1_reg_1_ ( .D(u5_N1), .CK(clk), .Q(u5_prod1[1]) );
  DFF_X2 u5_prod_reg_1_ ( .D(u5_prod1[1]), .CK(clk), .QN(n1537) );
  DFF_X2 u5_prod1_reg_2_ ( .D(u5_N2), .CK(clk), .Q(u5_prod1[2]) );
  DFF_X2 u5_prod_reg_2_ ( .D(u5_prod1[2]), .CK(clk), .Q(prod[2]) );
  DFF_X2 u5_prod1_reg_3_ ( .D(u5_N3), .CK(clk), .Q(u5_prod1[3]) );
  DFF_X2 u5_prod_reg_3_ ( .D(u5_prod1[3]), .CK(clk), .Q(prod[3]) );
  DFF_X2 u5_prod1_reg_4_ ( .D(u5_N4), .CK(clk), .Q(u5_prod1[4]) );
  DFF_X2 u5_prod_reg_4_ ( .D(u5_prod1[4]), .CK(clk), .Q(prod[4]) );
  DFF_X2 u5_prod1_reg_5_ ( .D(u5_N5), .CK(clk), .Q(u5_prod1[5]) );
  DFF_X2 u5_prod_reg_5_ ( .D(u5_prod1[5]), .CK(clk), .Q(prod[5]) );
  DFF_X2 u5_prod1_reg_6_ ( .D(u5_N6), .CK(clk), .Q(u5_prod1[6]) );
  DFF_X2 u5_prod_reg_6_ ( .D(u5_prod1[6]), .CK(clk), .Q(prod[6]) );
  DFF_X2 u5_prod1_reg_7_ ( .D(u5_N7), .CK(clk), .Q(u5_prod1[7]) );
  DFF_X2 u5_prod_reg_7_ ( .D(u5_prod1[7]), .CK(clk), .Q(prod[7]) );
  DFF_X2 u5_prod1_reg_8_ ( .D(u5_N8), .CK(clk), .Q(u5_prod1[8]) );
  DFF_X2 u5_prod_reg_8_ ( .D(u5_prod1[8]), .CK(clk), .Q(prod[8]), .QN(n1557)
         );
  DFF_X2 u5_prod1_reg_9_ ( .D(u5_N9), .CK(clk), .Q(u5_prod1[9]) );
  DFF_X2 u5_prod_reg_9_ ( .D(u5_prod1[9]), .CK(clk), .Q(prod[9]), .QN(n1570)
         );
  DFF_X2 u5_prod1_reg_10_ ( .D(u5_N10), .CK(clk), .Q(u5_prod1[10]) );
  DFF_X2 u5_prod_reg_10_ ( .D(u5_prod1[10]), .CK(clk), .QN(n1562) );
  DFF_X2 u5_prod1_reg_11_ ( .D(u5_N11), .CK(clk), .Q(u5_prod1[11]) );
  DFF_X2 u5_prod_reg_11_ ( .D(u5_prod1[11]), .CK(clk), .Q(prod[11]), .QN(n1568) );
  DFF_X2 u5_prod1_reg_12_ ( .D(u5_N12), .CK(clk), .Q(u5_prod1[12]) );
  DFF_X2 u5_prod_reg_12_ ( .D(u5_prod1[12]), .CK(clk), .Q(prod[12]), .QN(n1571) );
  DFF_X2 u5_prod1_reg_13_ ( .D(u5_N13), .CK(clk), .Q(u5_prod1[13]) );
  DFF_X2 u5_prod_reg_13_ ( .D(u5_prod1[13]), .CK(clk), .Q(prod[13]), .QN(n1569) );
  DFF_X2 u5_prod1_reg_14_ ( .D(u5_N14), .CK(clk), .Q(u5_prod1[14]) );
  DFF_X2 u5_prod_reg_14_ ( .D(u5_prod1[14]), .CK(clk), .Q(prod[14]), .QN(n1565) );
  DFF_X2 u5_prod1_reg_15_ ( .D(u5_N15), .CK(clk), .Q(u5_prod1[15]) );
  DFF_X2 u5_prod_reg_15_ ( .D(u5_prod1[15]), .CK(clk), .Q(prod[15]), .QN(n1567) );
  DFF_X2 u5_prod1_reg_16_ ( .D(u5_N16), .CK(clk), .Q(u5_prod1[16]) );
  DFF_X2 u5_prod_reg_16_ ( .D(u5_prod1[16]), .CK(clk), .Q(prod[16]), .QN(n1566) );
  DFF_X2 u5_prod1_reg_17_ ( .D(u5_N17), .CK(clk), .Q(u5_prod1[17]) );
  DFF_X2 u5_prod_reg_17_ ( .D(u5_prod1[17]), .CK(clk), .QN(n1563) );
  DFF_X2 u5_prod1_reg_18_ ( .D(u5_N18), .CK(clk), .Q(u5_prod1[18]) );
  DFF_X2 u5_prod_reg_18_ ( .D(u5_prod1[18]), .CK(clk), .QN(n1534) );
  DFF_X2 u5_prod1_reg_19_ ( .D(u5_N19), .CK(clk), .Q(u5_prod1[19]) );
  DFF_X2 u5_prod_reg_19_ ( .D(u5_prod1[19]), .CK(clk), .QN(n1545) );
  DFF_X2 u5_prod1_reg_20_ ( .D(u5_N20), .CK(clk), .Q(u5_prod1[20]) );
  DFF_X2 u5_prod_reg_20_ ( .D(u5_prod1[20]), .CK(clk), .QN(n1561) );
  DFF_X2 u5_prod1_reg_21_ ( .D(u5_N21), .CK(clk), .Q(u5_prod1[21]) );
  DFF_X2 u5_prod_reg_21_ ( .D(u5_prod1[21]), .CK(clk), .Q(prod[21]) );
  DFF_X2 u6_remainder_reg_0_ ( .D(u6_N0), .CK(clk), .Q(u6_remainder[0]) );
  DFF_X2 u6_rem_reg_0_ ( .D(u6_remainder[0]), .CK(clk), .Q(remainder[0]) );
  DFF_X2 u6_remainder_reg_1_ ( .D(u6_N1), .CK(clk), .Q(u6_remainder[1]) );
  DFF_X2 u6_rem_reg_1_ ( .D(u6_remainder[1]), .CK(clk), .QN(n1776) );
  DFF_X2 u6_remainder_reg_2_ ( .D(u6_N2), .CK(clk), .Q(u6_remainder[2]) );
  DFF_X2 u6_rem_reg_2_ ( .D(u6_remainder[2]), .CK(clk), .QN(n1775) );
  DFF_X2 u6_remainder_reg_3_ ( .D(u6_N3), .CK(clk), .Q(u6_remainder[3]) );
  DFF_X2 u6_rem_reg_3_ ( .D(u6_remainder[3]), .CK(clk), .QN(n1774) );
  DFF_X2 u6_remainder_reg_4_ ( .D(u6_N4), .CK(clk), .Q(u6_remainder[4]) );
  DFF_X2 u6_rem_reg_4_ ( .D(u6_remainder[4]), .CK(clk), .Q(remainder[4]) );
  DFF_X2 u6_remainder_reg_5_ ( .D(u6_N5), .CK(clk), .Q(u6_remainder[5]) );
  DFF_X2 u6_rem_reg_5_ ( .D(u6_remainder[5]), .CK(clk), .Q(remainder[5]) );
  DFF_X2 u6_remainder_reg_6_ ( .D(u6_N6), .CK(clk), .Q(u6_remainder[6]) );
  DFF_X2 u6_rem_reg_6_ ( .D(u6_remainder[6]), .CK(clk), .Q(remainder[6]) );
  DFF_X2 u6_remainder_reg_7_ ( .D(u6_N7), .CK(clk), .Q(u6_remainder[7]) );
  DFF_X2 u6_rem_reg_7_ ( .D(u6_remainder[7]), .CK(clk), .QN(n1773) );
  DFF_X2 u6_remainder_reg_8_ ( .D(u6_N8), .CK(clk), .Q(u6_remainder[8]) );
  DFF_X2 u6_rem_reg_8_ ( .D(u6_remainder[8]), .CK(clk), .QN(n1772) );
  DFF_X2 u6_remainder_reg_9_ ( .D(u6_N9), .CK(clk), .Q(u6_remainder[9]) );
  DFF_X2 u6_rem_reg_9_ ( .D(u6_remainder[9]), .CK(clk), .QN(n1771) );
  DFF_X2 u6_remainder_reg_10_ ( .D(u6_N10), .CK(clk), .Q(u6_remainder[10]) );
  DFF_X2 u6_rem_reg_10_ ( .D(u6_remainder[10]), .CK(clk), .Q(remainder[10]) );
  DFF_X2 u6_remainder_reg_13_ ( .D(u6_N13), .CK(clk), .Q(u6_remainder[13]) );
  DFF_X2 u6_rem_reg_13_ ( .D(u6_remainder[13]), .CK(clk), .QN(n1770) );
  DFF_X2 u6_remainder_reg_14_ ( .D(u6_N14), .CK(clk), .Q(u6_remainder[14]) );
  DFF_X2 u6_rem_reg_14_ ( .D(u6_remainder[14]), .CK(clk), .QN(n1769) );
  DFF_X2 u6_remainder_reg_15_ ( .D(u6_N15), .CK(clk), .Q(u6_remainder[15]) );
  DFF_X2 u6_rem_reg_15_ ( .D(u6_remainder[15]), .CK(clk), .Q(remainder[15]) );
  DFF_X2 u6_remainder_reg_16_ ( .D(u6_N16), .CK(clk), .Q(u6_remainder[16]) );
  DFF_X2 u6_rem_reg_16_ ( .D(u6_remainder[16]), .CK(clk), .Q(remainder[16]) );
  DFF_X2 u6_remainder_reg_17_ ( .D(u6_N17), .CK(clk), .Q(u6_remainder[17]) );
  DFF_X2 u6_rem_reg_17_ ( .D(u6_remainder[17]), .CK(clk), .Q(remainder[17]) );
  DFF_X2 u6_remainder_reg_18_ ( .D(u6_N18), .CK(clk), .Q(u6_remainder[18]) );
  DFF_X2 u6_rem_reg_18_ ( .D(u6_remainder[18]), .CK(clk), .QN(n1768) );
  DFF_X2 u6_remainder_reg_19_ ( .D(u6_N19), .CK(clk), .Q(u6_remainder[19]) );
  DFF_X2 u6_rem_reg_19_ ( .D(u6_remainder[19]), .CK(clk), .QN(n1767) );
  DFF_X2 u6_remainder_reg_20_ ( .D(u6_N20), .CK(clk), .Q(u6_remainder[20]) );
  DFF_X2 u6_rem_reg_20_ ( .D(u6_remainder[20]), .CK(clk), .Q(remainder[20]) );
  DFF_X2 u6_remainder_reg_21_ ( .D(u6_N21), .CK(clk), .Q(u6_remainder[21]) );
  DFF_X2 u6_rem_reg_21_ ( .D(u6_remainder[21]), .CK(clk), .Q(remainder[21]) );
  DFF_X2 u6_remainder_reg_22_ ( .D(u6_N22), .CK(clk), .Q(u6_remainder[22]) );
  DFF_X2 u6_rem_reg_22_ ( .D(u6_remainder[22]), .CK(clk), .Q(remainder[22]) );
  DFF_X2 u6_remainder_reg_23_ ( .D(u6_N23), .CK(clk), .Q(u6_remainder[23]) );
  DFF_X2 u6_rem_reg_23_ ( .D(u6_remainder[23]), .CK(clk), .QN(n1766) );
  DFF_X2 u6_quo1_reg_0_ ( .D(u6_N0), .CK(clk), .Q(u6_quo1[0]) );
  DFF_X2 u6_quo_reg_0_ ( .D(u6_quo1[0]), .CK(clk), .Q(quo[0]) );
  DFF_X2 u6_quo1_reg_1_ ( .D(u6_N1), .CK(clk), .Q(u6_quo1[1]) );
  DFF_X2 u6_quo_reg_1_ ( .D(u6_quo1[1]), .CK(clk), .Q(quo[1]) );
  DFF_X2 u6_quo1_reg_2_ ( .D(u6_N2), .CK(clk), .Q(u6_quo1[2]) );
  DFF_X2 u6_quo_reg_2_ ( .D(u6_quo1[2]), .CK(clk), .Q(quo[2]), .QN(n1572) );
  DFF_X2 u6_quo1_reg_3_ ( .D(u6_N3), .CK(clk), .Q(u6_quo1[3]) );
  DFF_X2 u6_quo_reg_3_ ( .D(u6_quo1[3]), .CK(clk), .Q(quo[3]), .QN(n1558) );
  DFF_X2 u6_quo1_reg_4_ ( .D(u6_N4), .CK(clk), .Q(u6_quo1[4]) );
  DFF_X2 u6_quo_reg_4_ ( .D(u6_quo1[4]), .CK(clk), .Q(quo[4]) );
  DFF_X2 u6_quo1_reg_5_ ( .D(u6_N5), .CK(clk), .Q(u6_quo1[5]) );
  DFF_X2 u6_quo_reg_5_ ( .D(u6_quo1[5]), .CK(clk), .Q(quo[5]) );
  DFF_X2 u6_quo1_reg_6_ ( .D(u6_N6), .CK(clk), .Q(u6_quo1[6]) );
  DFF_X2 u6_quo_reg_6_ ( .D(u6_quo1[6]), .CK(clk), .Q(quo[6]) );
  DFF_X2 u6_quo1_reg_7_ ( .D(u6_N7), .CK(clk), .Q(u6_quo1[7]) );
  DFF_X2 u6_quo_reg_7_ ( .D(u6_quo1[7]), .CK(clk), .Q(quo[7]) );
  DFF_X2 u6_quo1_reg_8_ ( .D(u6_N8), .CK(clk), .Q(u6_quo1[8]) );
  DFF_X2 u6_quo_reg_8_ ( .D(u6_quo1[8]), .CK(clk), .Q(quo[8]) );
  DFF_X2 u6_quo1_reg_9_ ( .D(u6_N9), .CK(clk), .Q(u6_quo1[9]) );
  DFF_X2 u6_quo_reg_9_ ( .D(u6_quo1[9]), .CK(clk), .Q(quo[9]), .QN(n1556) );
  DFF_X2 u6_quo1_reg_10_ ( .D(u6_N10), .CK(clk), .Q(u6_quo1[10]) );
  DFF_X2 u6_quo_reg_10_ ( .D(u6_quo1[10]), .CK(clk), .Q(quo[10]) );
  DFF_X2 u6_quo1_reg_13_ ( .D(u6_N13), .CK(clk), .Q(u6_quo1[13]) );
  DFF_X2 u6_quo_reg_13_ ( .D(u6_quo1[13]), .CK(clk), .Q(quo[13]), .QN(n1564)
         );
  DFF_X2 u6_quo1_reg_14_ ( .D(u6_N14), .CK(clk), .Q(u6_quo1[14]) );
  DFF_X2 u6_quo_reg_14_ ( .D(u6_quo1[14]), .CK(clk), .Q(quo[14]) );
  DFF_X2 u6_quo1_reg_15_ ( .D(u6_N15), .CK(clk), .Q(u6_quo1[15]) );
  DFF_X2 u6_quo_reg_15_ ( .D(u6_quo1[15]), .CK(clk), .Q(quo[15]) );
  DFF_X2 u6_quo1_reg_16_ ( .D(u6_N16), .CK(clk), .Q(u6_quo1[16]) );
  DFF_X2 u6_quo_reg_16_ ( .D(u6_quo1[16]), .CK(clk), .Q(quo[16]) );
  DFF_X2 u6_quo1_reg_17_ ( .D(u6_N17), .CK(clk), .Q(u6_quo1[17]) );
  DFF_X2 u6_quo_reg_17_ ( .D(u6_quo1[17]), .CK(clk), .Q(quo[17]) );
  DFF_X2 u6_quo1_reg_18_ ( .D(u6_N18), .CK(clk), .Q(u6_quo1[18]) );
  DFF_X2 u6_quo_reg_18_ ( .D(u6_quo1[18]), .CK(clk), .Q(quo[18]) );
  DFF_X2 u6_quo1_reg_19_ ( .D(u6_N19), .CK(clk), .Q(u6_quo1[19]) );
  DFF_X2 u6_quo_reg_19_ ( .D(u6_quo1[19]), .CK(clk), .Q(quo[19]) );
  DFF_X2 u6_quo1_reg_20_ ( .D(u6_N20), .CK(clk), .Q(u6_quo1[20]) );
  DFF_X2 u6_quo_reg_20_ ( .D(u6_quo1[20]), .CK(clk), .Q(quo[20]) );
  DFF_X2 u6_quo1_reg_21_ ( .D(u6_N21), .CK(clk), .Q(u6_quo1[21]) );
  DFF_X2 u6_quo_reg_21_ ( .D(u6_quo1[21]), .CK(clk), .Q(quo[21]) );
  DFF_X2 u6_quo1_reg_22_ ( .D(u6_N22), .CK(clk), .Q(u6_quo1[22]) );
  DFF_X2 u6_quo_reg_22_ ( .D(u6_quo1[22]), .CK(clk), .Q(quo[22]) );
  DFF_X2 out_reg_10_ ( .D(N230), .CK(clk), .Q(out[10]) );
  DFF_X2 out_reg_13_ ( .D(N233), .CK(clk), .Q(out[13]) );
  DFF_X2 out_reg_14_ ( .D(N234), .CK(clk), .Q(out[14]) );
  DFF_X2 out_reg_12_ ( .D(N232), .CK(clk), .Q(out[12]) );
  DFF_X2 out_reg_11_ ( .D(N231), .CK(clk), .Q(out[11]) );
  DFF_X2 overflow_reg ( .D(N278), .CK(clk), .Q(overflow) );
  DFF_X2 out_reg_9_ ( .D(N229), .CK(clk), .Q(out[9]) );
  DFF_X2 out_reg_8_ ( .D(N228), .CK(clk), .Q(out[8]) );
  DFF_X2 out_reg_7_ ( .D(N227), .CK(clk), .Q(out[7]) );
  DFF_X2 out_reg_6_ ( .D(N226), .CK(clk), .Q(out[6]) );
  DFF_X2 out_reg_5_ ( .D(N225), .CK(clk), .Q(out[5]) );
  DFF_X2 out_reg_4_ ( .D(N224), .CK(clk), .Q(out[4]) );
  DFF_X2 out_reg_3_ ( .D(N223), .CK(clk), .Q(out[3]) );
  DFF_X2 out_reg_2_ ( .D(N222), .CK(clk), .Q(out[2]) );
  DFF_X2 out_reg_1_ ( .D(N221), .CK(clk), .Q(out[1]) );
  DFF_X2 inf_reg ( .D(N285), .CK(clk), .Q(inf) );
  DFF_X2 underflow_reg ( .D(N281), .CK(clk), .Q(underflow) );
  DFF_X2 ine_reg ( .D(N268), .CK(clk), .Q(ine) );
  DFF_X2 zero_reg ( .D(N290), .CK(clk), .Q(zero) );
  DFF_X2 out_reg_15_ ( .D(N254), .CK(clk), .Q(out[15]) );
  DFF_X2 out_reg_0_ ( .D(N220), .CK(clk), .Q(out[0]) );
  DFF_X2 u6_quo1_reg_23_ ( .D(u6_N23), .CK(clk), .Q(u6_quo1[23]) );
  DFF_X2 u6_quo_reg_23_ ( .D(u6_quo1[23]), .CK(clk), .QN(n1765) );
  FA_X1 u4_sub_470_U2_1 ( .A(exp_r[1]), .B(n1657), .CI(u4_sub_470_carry[1]), 
        .CO(u4_sub_470_carry[2]), .S(u4_exp_fix_divb[1]) );
  FA_X1 u4_sub_470_U2_2 ( .A(exp_r[2]), .B(n1676), .CI(u4_sub_470_carry[2]), 
        .CO(u4_sub_470_carry[3]), .S(u4_exp_fix_divb[2]) );
  FA_X1 u4_sub_470_U2_3 ( .A(n1533), .B(n1675), .CI(u4_sub_470_carry[3]), .CO(
        u4_sub_470_carry[4]), .S(u4_exp_fix_divb[3]) );
  FA_X1 u4_sub_470_U2_4 ( .A(exp_r[4]), .B(n1674), .CI(u4_sub_470_carry[4]), 
        .S(u4_exp_fix_divb[4]) );
  HA_X1 u4_add_461_U1_1_1 ( .A(u4_exp_out_1_), .B(u4_exp_out_0_), .CO(
        u4_add_461_carry[2]), .S(u4_exp_out_pl1_1_) );
  HA_X1 u4_add_461_U1_1_2 ( .A(u4_exp_out_2_), .B(u4_add_461_carry[2]), .CO(
        u4_add_461_carry[3]), .S(u4_exp_out_pl1_2_) );
  HA_X1 u4_add_461_U1_1_3 ( .A(u4_exp_out_3_), .B(u4_add_461_carry[3]), .CO(
        u4_add_461_carry[4]), .S(u4_exp_out_pl1_3_) );
  FA_X1 u4_sub_409_U2_1 ( .A(div_opa_ldz_r2[1]), .B(n1784), .CI(
        u4_sub_409_carry[1]), .CO(u4_sub_409_carry[2]), .S(u4_div_shft4[1]) );
  FA_X1 u4_sub_409_U2_2 ( .A(div_opa_ldz_r2[2]), .B(n1782), .CI(
        u4_sub_409_carry[2]), .CO(u4_sub_409_carry[3]), .S(u4_div_shft4[2]) );
  FA_X1 u4_sub_409_U2_3 ( .A(div_opa_ldz_r2[3]), .B(n1780), .CI(
        u4_sub_409_carry[3]), .CO(u4_sub_409_carry[4]), .S(u4_div_shft4[3]) );
  FA_X1 u4_add_408_U1_1 ( .A(div_opa_ldz_r2[1]), .B(exp_r[1]), .CI(
        u4_add_408_carry[1]), .CO(u4_add_408_carry[2]), .S(u4_div_shft3_1_) );
  FA_X1 u4_add_408_U1_2 ( .A(div_opa_ldz_r2[2]), .B(exp_r[2]), .CI(
        u4_add_408_carry[2]), .CO(u4_add_408_carry[3]), .S(u4_div_shft3_2_) );
  FA_X1 u4_add_408_U1_3 ( .A(div_opa_ldz_r2[3]), .B(n1533), .CI(
        u4_add_408_carry[3]), .CO(u4_add_408_carry[4]), .S(u4_div_shft3_3_) );
  FA_X1 u4_sub_493_U2_1 ( .A(u4_exp_in_pl1_1_), .B(n1653), .CI(
        u4_sub_493_carry[1]), .CO(u4_sub_493_carry[2]), .S(u4_div_exp2[1]) );
  FA_X1 u4_sub_493_U2_2 ( .A(u4_exp_in_pl1_2_), .B(n1654), .CI(
        u4_sub_493_carry[2]), .CO(u4_sub_493_carry[3]), .S(u4_div_exp2[2]) );
  FA_X1 u4_sub_493_U2_3 ( .A(u4_exp_in_pl1_3_), .B(n1655), .CI(
        u4_sub_493_carry[3]), .CO(u4_sub_493_carry[4]), .S(u4_div_exp2[3]) );
  FA_X1 u4_sub_493_U2_4 ( .A(u4_exp_in_pl1_4_), .B(n1656), .CI(
        u4_sub_493_carry[4]), .S(u4_div_exp2[4]) );
  FA_X1 u4_add_486_U1_1 ( .A(div_opa_ldz_r2[1]), .B(u4_N264), .CI(
        u4_add_486_carry[1]), .CO(u4_add_486_carry[2]), .S(u4_ldz_all_1_) );
  FA_X1 u4_add_486_U1_2 ( .A(div_opa_ldz_r2[2]), .B(u4_N203), .CI(
        u4_add_486_carry[2]), .CO(u4_add_486_carry[3]), .S(u4_ldz_all_2_) );
  FA_X1 u4_add_486_U1_3 ( .A(div_opa_ldz_r2[3]), .B(u4_N152), .CI(
        u4_add_486_carry[3]), .CO(u4_add_486_carry[4]), .S(u4_ldz_all_3_) );
  HA_X1 u4_add_463_U1_1_1 ( .A(exp_r[1]), .B(n1626), .CO(u4_add_463_carry[2]), 
        .S(u4_exp_in_pl1_1_) );
  HA_X1 u4_add_463_U1_1_2 ( .A(exp_r[2]), .B(u4_add_463_carry[2]), .CO(
        u4_add_463_carry[3]), .S(u4_exp_in_pl1_2_) );
  HA_X1 u4_add_463_U1_1_3 ( .A(n1533), .B(u4_add_463_carry[3]), .CO(
        u4_add_463_carry[4]), .S(u4_exp_in_pl1_3_) );
  HA_X1 u4_add_463_U1_1_4 ( .A(exp_r[4]), .B(u4_add_463_carry[4]), .CO(
        u4_exp_in_pl1_5_), .S(u4_exp_in_pl1_4_) );
  FA_X1 u4_add_491_U1_1 ( .A(u4_exp_in_mi1_1_), .B(u4_fi_ldz_2a_1_), .CI(
        u4_add_491_carry[1]), .CO(u4_add_491_carry[2]), .S(u4_div_exp1_1_) );
  FA_X1 u4_add_491_U1_2 ( .A(u4_exp_in_mi1_2_), .B(u4_fi_ldz_2a_2_), .CI(
        u4_add_491_carry[2]), .CO(u4_add_491_carry[3]), .S(u4_div_exp1_2_) );
  FA_X1 u4_add_491_U1_3 ( .A(u4_exp_in_mi1_3_), .B(u4_fi_ldz_2a_3_), .CI(
        u4_add_491_carry[3]), .CO(u4_add_491_carry[4]), .S(u4_div_exp1_3_) );
  FA_X1 u4_add_491_U1_4 ( .A(u4_exp_in_mi1_4_), .B(u4_fi_ldz_2a_4_), .CI(
        u4_add_491_carry[4]), .S(u4_div_exp1_4_) );
  FA_X1 u4_sub_406_U2_1 ( .A(exp_r[1]), .B(n1829), .CI(u4_sub_406_carry[1]), 
        .CO(u4_sub_406_carry[2]), .S(u4_div_scht1a[1]) );
  FA_X1 u4_sub_406_U2_2 ( .A(exp_r[2]), .B(n1830), .CI(u4_sub_406_carry[2]), 
        .CO(u4_sub_406_carry[3]), .S(u4_div_scht1a[2]) );
  FA_X1 u4_sub_406_U2_3 ( .A(n1533), .B(n2475), .CI(u4_sub_406_carry[3]), .CO(
        u4_sub_406_carry[4]), .S(u4_div_scht1a[3]) );
  HA_X1 u2_add_115_U1_1_1 ( .A(u2_exp_tmp4_1_), .B(u2_exp_tmp4_0_), .CO(
        u2_add_115_carry[2]), .S(u2_N31) );
  HA_X1 u2_add_115_U1_1_2 ( .A(u2_exp_tmp4_2_), .B(u2_add_115_carry[2]), .CO(
        u2_add_115_carry[3]), .S(u2_N32) );
  HA_X1 u2_add_115_U1_1_3 ( .A(u2_exp_tmp4_3_), .B(u2_add_115_carry[3]), .CO(
        u2_add_115_carry[4]), .S(u2_N33) );
  HA_X1 u2_add_113_U1_1_1 ( .A(u2_add_113_A_1_), .B(u2_add_113_A_0_), .CO(
        u2_add_113_carry[2]), .S(u2_exp_tmp3_1_) );
  HA_X1 u2_add_113_U1_1_2 ( .A(u2_add_113_A_2_), .B(u2_add_113_carry[2]), .CO(
        u2_add_113_carry[3]), .S(u2_exp_tmp3_2_) );
  HA_X1 u2_add_113_U1_1_3 ( .A(u2_add_113_A_3_), .B(u2_add_113_carry[3]), .CO(
        u2_add_113_carry[4]), .S(u2_exp_tmp3_3_) );
  FA_X1 u2_add_110_U1_1 ( .A(opa_r[11]), .B(opb_r[11]), .CI(
        u2_add_110_carry[1]), .CO(u2_add_110_carry[2]), .S(u2_N13) );
  FA_X1 u2_add_110_U1_2 ( .A(opa_r[12]), .B(opb_r[12]), .CI(
        u2_add_110_carry[2]), .CO(u2_add_110_carry[3]), .S(u2_N14) );
  FA_X1 u2_add_110_U1_3 ( .A(opa_r[13]), .B(opb_r[13]), .CI(
        u2_add_110_carry[3]), .CO(u2_add_110_carry[4]), .S(u2_N15) );
  FA_X1 u2_add_110_U1_4 ( .A(opa_r[14]), .B(opb_r[14]), .CI(
        u2_add_110_carry[4]), .CO(u2_N17), .S(u2_N16) );
  FA_X1 u2_sub_110_U2_1 ( .A(opa_r[11]), .B(n1587), .CI(u2_sub_110_carry[1]), 
        .CO(u2_sub_110_carry[2]), .S(u2_N7) );
  FA_X1 u2_sub_110_U2_2 ( .A(opa_r[12]), .B(n1584), .CI(u2_sub_110_carry[2]), 
        .CO(u2_sub_110_carry[3]), .S(u2_N8) );
  FA_X1 u2_sub_110_U2_3 ( .A(opa_r[13]), .B(n1583), .CI(u2_sub_110_carry[3]), 
        .CO(u2_sub_110_carry[4]), .S(u2_N9) );
  FA_X1 u2_sub_110_U2_4 ( .A(opa_r[14]), .B(n1582), .CI(u2_sub_110_carry[4]), 
        .CO(u2_sub_110_carry[5]), .S(u2_N10) );
  FA_X1 sub_1_root_u1_sub_128_aco_U2_0 ( .A(sub_1_root_u1_sub_128_aco_A_0_), 
        .B(n1638), .CI(n1934), .CO(sub_1_root_u1_sub_128_aco_carry[1]), .S(
        u1_exp_diff2[0]) );
  FA_X1 sub_1_root_u1_sub_128_aco_U2_1 ( .A(sub_1_root_u1_sub_128_aco_A_1_), 
        .B(n1639), .CI(sub_1_root_u1_sub_128_aco_carry[1]), .CO(
        sub_1_root_u1_sub_128_aco_carry[2]), .S(u1_exp_diff2[1]) );
  FA_X1 sub_1_root_u1_sub_128_aco_U2_2 ( .A(sub_1_root_u1_sub_128_aco_A_2_), 
        .B(n1640), .CI(sub_1_root_u1_sub_128_aco_carry[2]), .CO(
        sub_1_root_u1_sub_128_aco_carry[3]), .S(u1_exp_diff2[2]) );
  FA_X1 sub_1_root_u1_sub_128_aco_U2_3 ( .A(sub_1_root_u1_sub_128_aco_A_3_), 
        .B(n1641), .CI(sub_1_root_u1_sub_128_aco_carry[3]), .CO(
        sub_1_root_u1_sub_128_aco_carry[4]), .S(u1_exp_diff2[3]) );
  FA_X1 sub_1_root_u1_sub_128_aco_U2_4 ( .A(sub_1_root_u1_sub_128_aco_A_4_), 
        .B(n1642), .CI(sub_1_root_u1_sub_128_aco_carry[4]), .S(u1_exp_diff2[4]) );
  FA_X1 sub_0_root_sub_0_root_u4_sub_469_U2_1 ( .A(u4_fi_ldz_mi22_1_), .B(
        n2351), .CI(sub_0_root_sub_0_root_u4_sub_469_carry[1]), .CO(
        sub_0_root_sub_0_root_u4_sub_469_carry[2]), .S(u4_exp_fix_diva[1]) );
  FA_X1 sub_0_root_sub_0_root_u4_sub_469_U2_2 ( .A(u4_fi_ldz_mi22_2_), .B(
        n2362), .CI(sub_0_root_sub_0_root_u4_sub_469_carry[2]), .CO(
        sub_0_root_sub_0_root_u4_sub_469_carry[3]), .S(u4_exp_fix_diva[2]) );
  FA_X1 sub_0_root_sub_0_root_u4_sub_469_U2_3 ( .A(u4_fi_ldz_mi22_3_), .B(
        n1666), .CI(sub_0_root_sub_0_root_u4_sub_469_carry[3]), .CO(
        sub_0_root_sub_0_root_u4_sub_469_carry[4]), .S(u4_exp_fix_diva[3]) );
  FA_X1 sub_0_root_sub_0_root_u4_sub_469_U2_4 ( .A(u4_fi_ldz_mi22_4_), .B(
        n2349), .CI(sub_0_root_sub_0_root_u4_sub_469_carry[4]), .S(
        u4_exp_fix_diva[4]) );
  FA_X1 add_0_root_sub_0_root_u4_add_494_U1_1 ( .A(u4_ldz_dif_1_), .B(
        u4_fi_ldz_2a_1_), .CI(add_0_root_sub_0_root_u4_add_494_carry[1]), .CO(
        add_0_root_sub_0_root_u4_add_494_carry[2]), .S(u4_div_exp3[1]) );
  FA_X1 add_0_root_sub_0_root_u4_add_494_U1_2 ( .A(u4_ldz_dif_2_), .B(
        u4_fi_ldz_2a_2_), .CI(add_0_root_sub_0_root_u4_add_494_carry[2]), .CO(
        add_0_root_sub_0_root_u4_add_494_carry[3]), .S(u4_div_exp3[2]) );
  FA_X1 add_0_root_sub_0_root_u4_add_494_U1_3 ( .A(u4_ldz_dif_3_), .B(
        u4_fi_ldz_2a_3_), .CI(add_0_root_sub_0_root_u4_add_494_carry[3]), .CO(
        add_0_root_sub_0_root_u4_add_494_carry[4]), .S(u4_div_exp3[3]) );
  FA_X1 add_0_root_sub_0_root_u4_add_494_U1_4 ( .A(u4_ldz_dif_4_), .B(
        u4_fi_ldz_2a_4_), .CI(add_0_root_sub_0_root_u4_add_494_carry[4]), .S(
        u4_div_exp3[4]) );
  FA_X1 sub_1_root_sub_0_root_u4_add_494_U2_1 ( .A(exp_r[1]), .B(n1829), .CI(
        sub_1_root_sub_0_root_u4_add_494_carry[1]), .CO(
        sub_1_root_sub_0_root_u4_add_494_carry[2]), .S(u4_ldz_dif_1_) );
  FA_X1 sub_1_root_sub_0_root_u4_add_494_U2_2 ( .A(exp_r[2]), .B(n1830), .CI(
        sub_1_root_sub_0_root_u4_add_494_carry[2]), .CO(
        sub_1_root_sub_0_root_u4_add_494_carry[3]), .S(u4_ldz_dif_2_) );
  FA_X1 sub_1_root_sub_0_root_u4_add_494_U2_3 ( .A(n1533), .B(n2475), .CI(
        sub_1_root_sub_0_root_u4_add_494_carry[3]), .CO(
        sub_1_root_sub_0_root_u4_add_494_carry[4]), .S(u4_ldz_dif_3_) );
  NAND2_X2 U1188 ( .A1(n1770), .A2(n1769), .ZN(n2455) );
  NAND2_X2 U1189 ( .A1(n1524), .A2(n1525), .ZN(u4_sub_406_carry[5]) );
  XNOR2_X2 U1190 ( .A(exp_r[4]), .B(u4_sub_406_carry[4]), .ZN(u4_div_scht1a[4]) );
  INV_X4 U1191 ( .A(exp_r[4]), .ZN(n1524) );
  INV_X4 U1192 ( .A(u4_sub_406_carry[4]), .ZN(n1525) );
  XNOR2_X2 U1193 ( .A(exp_r[4]), .B(sub_1_root_sub_0_root_u4_add_494_carry[4]), 
        .ZN(u4_ldz_dif_4_) );
  AOI222_X1 U1194 ( .A1(quo[2]), .A2(n2487), .B1(n2065), .B2(fract_out_q[3]), 
        .C1(1'b0), .C2(n2481), .ZN(n2498) );
  AOI222_X1 U1195 ( .A1(1'b0), .A2(n2487), .B1(n2065), .B2(fract_out_q[13]), 
        .C1(quo[22]), .C2(n2481), .ZN(n2486) );
  AOI222_X1 U1196 ( .A1(quo[1]), .A2(n2487), .B1(n2065), .B2(fract_out_q[2]), 
        .C1(1'b0), .C2(n2481), .ZN(n2497) );
  AOI222_X1 U1197 ( .A1(1'b0), .A2(n2487), .B1(n2065), .B2(fract_out_q[12]), 
        .C1(quo[21]), .C2(n2481), .ZN(n2488) );
  NOR4_X1 U1198 ( .A1(n2455), .A2(remainder[0]), .A3(1'b0), .A4(remainder[10]), 
        .ZN(n2448) );
  XNOR2_X2 U1199 ( .A(n1777), .B(u4_sub_409_carry[4]), .ZN(n1526) );
  INV_X4 U1200 ( .A(n1526), .ZN(u4_div_shft4[4]) );
  XNOR2_X2 U1201 ( .A(exp_r[4]), .B(u4_add_408_carry[4]), .ZN(n1527) );
  INV_X4 U1202 ( .A(n1527), .ZN(u4_div_shft3_4_) );
  NAND2_X2 U1203 ( .A1(u4_N95), .A2(u4_add_486_carry[4]), .ZN(n1528) );
  INV_X4 U1204 ( .A(n1528), .ZN(u4_ldz_all_5_) );
  XNOR2_X2 U1205 ( .A(u4_N95), .B(u4_add_486_carry[4]), .ZN(n1529) );
  INV_X4 U1206 ( .A(n1529), .ZN(u4_ldz_all_4_) );
  INV_X4 U1207 ( .A(n1777), .ZN(n2404) );
  NAND2_X2 U1208 ( .A1(n2405), .A2(n2406), .ZN(n2403) );
  NOR3_X2 U1209 ( .A1(n2460), .A2(n2461), .A3(n2462), .ZN(n2437) );
  NOR2_X2 U1210 ( .A1(u4_N386), .A2(n2466), .ZN(n2439) );
  INV_X4 U1211 ( .A(n2483), .ZN(n2481) );
  NAND2_X2 U1212 ( .A1(n2265), .A2(n2271), .ZN(n2232) );
  NAND2_X2 U1213 ( .A1(n2265), .A2(n2266), .ZN(n2233) );
  OAI211_X2 U1214 ( .C1(n2149), .C2(n2259), .A(n2260), .B(n2200), .ZN(n2235)
         );
  INV_X4 U1215 ( .A(n1924), .ZN(n1941) );
  INV_X4 U1216 ( .A(u4_div_shft2[0]), .ZN(n1625) );
  INV_X4 U1217 ( .A(n2482), .ZN(n2484) );
  NOR2_X2 U1218 ( .A1(n2507), .A2(n1831), .ZN(n1877) );
  NAND3_X2 U1219 ( .A1(fpu_op_r1[0]), .A2(fpu_op_r1[1]), .A3(n1837), .ZN(n1924) );
  NAND2_X2 U1220 ( .A1(n2531), .A2(n2513), .ZN(n1990) );
  NAND2_X2 U1221 ( .A1(n2527), .A2(n2040), .ZN(n2519) );
  NAND2_X2 U1222 ( .A1(n2513), .A2(n2040), .ZN(n2520) );
  NAND2_X2 U1223 ( .A1(n1551), .A2(n2521), .ZN(n2514) );
  NOR2_X2 U1224 ( .A1(n2484), .A2(n1560), .ZN(n2124) );
  INV_X4 U1225 ( .A(fract_denorm[21]), .ZN(n1902) );
  INV_X4 U1226 ( .A(n2698), .ZN(n1522) );
  AND4_X4 U1227 ( .A1(n1621), .A2(n1620), .A3(n1622), .A4(n2532), .ZN(n1530)
         );
  NAND2_X2 U1228 ( .A1(n1628), .A2(n2501), .ZN(n1531) );
  INV_X4 U1229 ( .A(n1630), .ZN(n1629) );
  XNOR2_X2 U1230 ( .A(n1618), .B(sub_434_3_carry[17]), .ZN(n1532) );
  INV_X4 U1231 ( .A(n1632), .ZN(n1631) );
  OAI21_X2 U1232 ( .B1(opb_r[14]), .B2(n1577), .A(n1684), .ZN(u1_expa_lt_expb)
         );
  XNOR2_X2 U1233 ( .A(n1619), .B(sub_434_3_carry[16]), .ZN(n1535) );
  INV_X4 U1234 ( .A(n1625), .ZN(n1626) );
  INV_X4 U1235 ( .A(n1966), .ZN(n1630) );
  INV_X4 U1236 ( .A(n1623), .ZN(n1624) );
  XNOR2_X2 U1237 ( .A(n1622), .B(sub_434_3_carry[18]), .ZN(n1550) );
  NAND2_X2 U1238 ( .A1(sub_434_b0_carry[10]), .A2(n1530), .ZN(n1551) );
  NAND2_X2 U1239 ( .A1(sub_434_3_carry[20]), .A2(n1620), .ZN(n1552) );
  OAI221_X2 U1240 ( .B1(n1631), .B2(n2509), .C1(n1807), .C2(n2507), .A(n2510), 
        .ZN(fract_denorm[21]) );
  XNOR2_X2 U1241 ( .A(u4_fi_ldz_2a_0_), .B(div_opa_ldz_r2[0]), .ZN(n1559) );
  INV_X4 U1242 ( .A(n1560), .ZN(n1628) );
  NAND2_X2 U1243 ( .A1(n2395), .A2(n2396), .ZN(u4_exp_out_0_) );
  INV_X4 U1244 ( .A(n1531), .ZN(n1632) );
  OAI21_X2 U1245 ( .B1(fract_denorm[20]), .B2(n1901), .A(n1902), .ZN(
        u4_fi_ldz_2a_0_) );
  INV_X4 U1246 ( .A(u1_fractb_lt_fracta), .ZN(n1634) );
  INV_X4 U1247 ( .A(n1634), .ZN(n1633) );
  INV_X4 U1248 ( .A(n1625), .ZN(n1627) );
  XNOR2_X2 U1249 ( .A(n1614), .B(sub_434_3_carry[15]), .ZN(n1585) );
  XNOR2_X2 U1250 ( .A(n1615), .B(sub_434_3_carry[14]), .ZN(n1586) );
  XNOR2_X2 U1251 ( .A(n1616), .B(sub_434_3_carry[13]), .ZN(n1601) );
  XNOR2_X2 U1252 ( .A(n1617), .B(sub_434_3_carry[12]), .ZN(n1602) );
  XNOR2_X2 U1253 ( .A(n1612), .B(sub_434_3_carry[11]), .ZN(n1603) );
  XNOR2_X2 U1254 ( .A(n1589), .B(sub_434_b0_carry[3]), .ZN(n1605) );
  XNOR2_X2 U1255 ( .A(n1590), .B(sub_434_b0_carry[2]), .ZN(n1606) );
  XNOR2_X2 U1256 ( .A(n1591), .B(n1599), .ZN(n1607) );
  INV_X4 U1260 ( .A(u1_expa_lt_expb), .ZN(n1623) );
  NAND3_X2 U1261 ( .A1(n1580), .A2(n1578), .A3(n2037), .ZN(n2698) );
  OAI22_X2 U1262 ( .A1(n2189), .A2(n2252), .B1(n1888), .B2(n2253), .ZN(n2229)
         );
  AND3_X4 U1263 ( .A1(n2473), .A2(n1902), .A3(n2435), .ZN(u4_N152) );
  INV_X4 U1264 ( .A(n2096), .ZN(n2155) );
  AND2_X4 U1265 ( .A1(n2501), .A2(n1538), .ZN(n2487) );
  INV_X4 U1266 ( .A(n2125), .ZN(n2065) );
  XOR2_X1 U1267 ( .A(exp_r[4]), .B(add_1_root_sub_0_root_u4_sub_469_carry_4_), 
        .Z(u4_fi_ldz_mi22_4_) );
  OR2_X1 U1268 ( .A1(n1533), .A2(add_1_root_sub_0_root_u4_sub_469_carry_3_), 
        .ZN(add_1_root_sub_0_root_u4_sub_469_carry_4_) );
  XNOR2_X1 U1269 ( .A(add_1_root_sub_0_root_u4_sub_469_carry_3_), .B(n1533), 
        .ZN(u4_fi_ldz_mi22_3_) );
  AND2_X1 U1270 ( .A1(exp_r[2]), .A2(add_1_root_sub_0_root_u4_sub_469_carry_2_), .ZN(add_1_root_sub_0_root_u4_sub_469_carry_3_) );
  XOR2_X1 U1271 ( .A(exp_r[2]), .B(add_1_root_sub_0_root_u4_sub_469_carry_2_), 
        .Z(u4_fi_ldz_mi22_2_) );
  AND2_X1 U1272 ( .A1(exp_r[1]), .A2(n1627), .ZN(
        add_1_root_sub_0_root_u4_sub_469_carry_2_) );
  XOR2_X1 U1273 ( .A(n1891), .B(n1627), .Z(u4_fi_ldz_mi22_1_) );
  OR2_X1 U1274 ( .A1(u4_fi_ldz_2a_0_), .A2(n1626), .ZN(u4_sub_470_carry[1]) );
  XNOR2_X1 U1275 ( .A(n1626), .B(u4_fi_ldz_2a_0_), .ZN(u4_exp_fix_divb[0]) );
  OR2_X1 U1276 ( .A1(n1667), .A2(n1668), .ZN(
        sub_0_root_sub_0_root_u4_sub_469_carry[1]) );
  XNOR2_X1 U1277 ( .A(n1668), .B(n1667), .ZN(u4_exp_fix_diva[0]) );
  XOR2_X1 U1278 ( .A(exp_r[4]), .B(u4_add_407_carry[4]), .Z(u4_div_shft2[4])
         );
  AND2_X1 U1279 ( .A1(n1533), .A2(u4_add_407_carry[3]), .ZN(
        u4_add_407_carry[4]) );
  XOR2_X1 U1280 ( .A(n1533), .B(u4_add_407_carry[3]), .Z(u4_div_shft2[3]) );
  AND2_X1 U1281 ( .A1(exp_r[2]), .A2(n1891), .ZN(u4_add_407_carry[3]) );
  XOR2_X1 U1282 ( .A(exp_r[2]), .B(n1891), .Z(u4_div_shft2[2]) );
  XOR2_X1 U1283 ( .A(n2349), .B(u4_sub_488_carry[4]), .Z(u4_fi_ldz_2a_4_) );
  OR2_X1 U1284 ( .A1(n1666), .A2(u4_sub_488_carry[3]), .ZN(u4_sub_488_carry[4]) );
  XNOR2_X1 U1285 ( .A(u4_sub_488_carry[3]), .B(n1666), .ZN(u4_fi_ldz_2a_3_) );
  AND2_X1 U1286 ( .A1(u4_sub_488_carry[2]), .A2(n2362), .ZN(
        u4_sub_488_carry[3]) );
  XOR2_X1 U1287 ( .A(n2362), .B(u4_sub_488_carry[2]), .Z(u4_fi_ldz_2a_2_) );
  XNOR2_X1 U1288 ( .A(n2349), .B(u4_sub_478_carry[4]), .ZN(u4_N447) );
  OR2_X1 U1289 ( .A1(n1666), .A2(u4_sub_478_carry[3]), .ZN(u4_sub_478_carry[4]) );
  XNOR2_X1 U1290 ( .A(u4_sub_478_carry[3]), .B(n1666), .ZN(u4_N446) );
  OR2_X1 U1291 ( .A1(n2362), .A2(u4_sub_478_carry[2]), .ZN(u4_sub_478_carry[3]) );
  XNOR2_X1 U1292 ( .A(u4_sub_478_carry[2]), .B(n2362), .ZN(u4_N445) );
  AND2_X1 U1293 ( .A1(u4_fi_ldz_2a_0_), .A2(u4_ldz_dif_0_), .ZN(
        add_0_root_sub_0_root_u4_add_494_carry[1]) );
  XOR2_X1 U1294 ( .A(u4_fi_ldz_2a_0_), .B(u4_ldz_dif_0_), .Z(u4_div_exp3[0])
         );
  OR2_X1 U1295 ( .A1(n1828), .A2(n1626), .ZN(
        sub_1_root_sub_0_root_u4_add_494_carry[1]) );
  XNOR2_X1 U1296 ( .A(n1627), .B(n1828), .ZN(u4_ldz_dif_0_) );
  XOR2_X1 U1297 ( .A(exp_r[4]), .B(u4_sub_414_carry_4_), .Z(u4_f2i_shft_4_) );
  AND2_X1 U1298 ( .A1(u4_sub_414_carry_3_), .A2(n1533), .ZN(
        u4_sub_414_carry_4_) );
  XOR2_X1 U1299 ( .A(n1533), .B(u4_sub_414_carry_3_), .Z(u4_f2i_shft_3_) );
  AND2_X1 U1300 ( .A1(u4_sub_414_carry_2_), .A2(exp_r[2]), .ZN(
        u4_sub_414_carry_3_) );
  XOR2_X1 U1301 ( .A(exp_r[2]), .B(u4_sub_414_carry_2_), .Z(u4_f2i_shft_2_) );
  OR2_X1 U1302 ( .A1(n1891), .A2(n1627), .ZN(u4_sub_414_carry_2_) );
  XNOR2_X1 U1303 ( .A(n1627), .B(n1891), .ZN(u4_f2i_shft_1_) );
  OR2_X1 U1304 ( .A1(n2351), .A2(n1667), .ZN(u4_sub_478_carry[2]) );
  XNOR2_X1 U1305 ( .A(n1667), .B(n2351), .ZN(u4_N444) );
  OR2_X1 U1306 ( .A1(n1559), .A2(u4_exp_in_pl1_0_), .ZN(u4_sub_493_carry[1])
         );
  XNOR2_X1 U1307 ( .A(u4_exp_in_pl1_0_), .B(n1559), .ZN(u4_div_exp2[0]) );
  AND2_X1 U1308 ( .A1(u4_fi_ldz_2a_0_), .A2(div_opa_ldz_r2[0]), .ZN(
        u4_add_486_carry[1]) );
  AND2_X1 U1309 ( .A1(u4_fi_ldz_2a_0_), .A2(n1668), .ZN(u4_add_491_carry[1])
         );
  XOR2_X1 U1310 ( .A(u4_fi_ldz_2a_0_), .B(n1668), .Z(u4_div_exp1_0_) );
  OR2_X1 U1311 ( .A1(n2351), .A2(n1667), .ZN(u4_sub_488_carry[2]) );
  XNOR2_X1 U1312 ( .A(n1667), .B(n2351), .ZN(u4_fi_ldz_2a_1_) );
  OR2_X1 U1313 ( .A1(n1828), .A2(n1627), .ZN(u4_sub_406_carry[1]) );
  XNOR2_X1 U1314 ( .A(n1626), .B(n1828), .ZN(u4_div_scht1a[0]) );
  OR2_X1 U1315 ( .A1(n1668), .A2(div_opa_ldz_r2[0]), .ZN(u4_sub_409_carry[1])
         );
  XNOR2_X1 U1316 ( .A(div_opa_ldz_r2[0]), .B(n1668), .ZN(u4_div_shft4[0]) );
  AND2_X1 U1317 ( .A1(n1626), .A2(div_opa_ldz_r2[0]), .ZN(u4_add_408_carry[1])
         );
  XOR2_X1 U1318 ( .A(n1626), .B(div_opa_ldz_r2[0]), .Z(u4_div_shft3_0_) );
  XOR2_X1 U1319 ( .A(u2_gt_140_B_5_), .B(u2_add_111_carry_5_), .Z(u2_N23) );
  AND2_X1 U1320 ( .A1(u2_add_111_carry_4_), .A2(u2_exp_tmp4_4_), .ZN(
        u2_add_111_carry_5_) );
  XOR2_X1 U1321 ( .A(u2_exp_tmp4_4_), .B(u2_add_111_carry_4_), .Z(u2_N22) );
  OR2_X1 U1322 ( .A1(u2_lt_130_A_3_), .A2(u2_add_111_carry_3_), .ZN(
        u2_add_111_carry_4_) );
  XNOR2_X1 U1323 ( .A(u2_add_111_carry_3_), .B(u2_lt_130_A_3_), .ZN(u2_N21) );
  OR2_X1 U1324 ( .A1(u2_lt_130_A_2_), .A2(u2_add_111_carry_2_), .ZN(
        u2_add_111_carry_3_) );
  XNOR2_X1 U1325 ( .A(u2_add_111_carry_2_), .B(u2_lt_130_A_2_), .ZN(u2_N20) );
  OR2_X1 U1326 ( .A1(u2_lt_130_A_1_), .A2(u2_lt_130_A_0_), .ZN(
        u2_add_111_carry_2_) );
  XNOR2_X1 U1327 ( .A(u2_lt_130_A_0_), .B(u2_lt_130_A_1_), .ZN(u2_N19) );
  XNOR2_X1 U1328 ( .A(u2_gt_140_B_5_), .B(u2_sub_111_carry_5_), .ZN(u2_N29) );
  OR2_X1 U1329 ( .A1(u2_exp_tmp4_4_), .A2(u2_sub_111_carry_4_), .ZN(
        u2_sub_111_carry_5_) );
  XNOR2_X1 U1330 ( .A(u2_sub_111_carry_4_), .B(u2_exp_tmp4_4_), .ZN(u2_N28) );
  AND2_X1 U1331 ( .A1(u2_sub_111_carry_3_), .A2(u2_lt_130_A_3_), .ZN(
        u2_sub_111_carry_4_) );
  XOR2_X1 U1332 ( .A(u2_lt_130_A_3_), .B(u2_sub_111_carry_3_), .Z(u2_N27) );
  AND2_X1 U1333 ( .A1(u2_sub_111_carry_2_), .A2(u2_lt_130_A_2_), .ZN(
        u2_sub_111_carry_3_) );
  XOR2_X1 U1334 ( .A(u2_lt_130_A_2_), .B(u2_sub_111_carry_2_), .Z(u2_N26) );
  AND2_X1 U1335 ( .A1(u2_lt_130_A_0_), .A2(u2_lt_130_A_1_), .ZN(
        u2_sub_111_carry_2_) );
  XOR2_X1 U1336 ( .A(u2_lt_130_A_1_), .B(u2_lt_130_A_0_), .Z(u2_N25) );
  AND2_X1 U1337 ( .A1(opa_r[10]), .A2(opb_r[10]), .ZN(u2_add_110_carry[1]) );
  XOR2_X1 U1338 ( .A(opb_r[10]), .B(opa_r[10]), .Z(u2_N12) );
  OR2_X1 U1339 ( .A1(n1588), .A2(opa_r[10]), .ZN(u2_sub_110_carry[1]) );
  XNOR2_X1 U1340 ( .A(opa_r[10]), .B(n1588), .ZN(u2_N6) );
  XOR2_X1 U1341 ( .A(n1620), .B(sub_434_3_carry[20]), .Z(N151) );
  AND2_X1 U1342 ( .A1(sub_434_3_carry[19]), .A2(n1621), .ZN(
        sub_434_3_carry[20]) );
  XOR2_X1 U1343 ( .A(n1621), .B(sub_434_3_carry[19]), .Z(N150) );
  AND2_X1 U1344 ( .A1(sub_434_3_carry[18]), .A2(n1622), .ZN(
        sub_434_3_carry[19]) );
  AND2_X1 U1345 ( .A1(sub_434_3_carry[17]), .A2(n1618), .ZN(
        sub_434_3_carry[18]) );
  AND2_X1 U1346 ( .A1(sub_434_3_carry[16]), .A2(n1619), .ZN(
        sub_434_3_carry[17]) );
  AND2_X1 U1347 ( .A1(sub_434_3_carry[15]), .A2(n1614), .ZN(
        sub_434_3_carry[16]) );
  AND2_X1 U1348 ( .A1(sub_434_3_carry[14]), .A2(n1615), .ZN(
        sub_434_3_carry[15]) );
  AND2_X1 U1349 ( .A1(sub_434_3_carry[13]), .A2(n1616), .ZN(
        sub_434_3_carry[14]) );
  AND2_X1 U1350 ( .A1(sub_434_3_carry[12]), .A2(n1617), .ZN(
        sub_434_3_carry[13]) );
  AND2_X1 U1351 ( .A1(sub_434_3_carry[11]), .A2(n1612), .ZN(
        sub_434_3_carry[12]) );
  AND2_X1 U1352 ( .A1(sub_434_3_carry[10]), .A2(n1613), .ZN(
        sub_434_3_carry[11]) );
  XOR2_X1 U1353 ( .A(n1613), .B(sub_434_3_carry[10]), .Z(N141) );
  AND2_X1 U1354 ( .A1(sub_434_3_carry[9]), .A2(n1589), .ZN(sub_434_3_carry[10]) );
  XOR2_X1 U1355 ( .A(n1589), .B(sub_434_3_carry[9]), .Z(N140) );
  AND2_X1 U1356 ( .A1(sub_434_3_carry[8]), .A2(n1590), .ZN(sub_434_3_carry[9])
         );
  XOR2_X1 U1357 ( .A(n1590), .B(sub_434_3_carry[8]), .Z(N139) );
  AND2_X1 U1358 ( .A1(n1599), .A2(n1591), .ZN(sub_434_3_carry[8]) );
  XOR2_X1 U1359 ( .A(n1591), .B(n1599), .Z(N138) );
  XOR2_X1 U1360 ( .A(n1530), .B(sub_434_b0_carry[10]), .Z(N116) );
  AND2_X1 U1361 ( .A1(sub_434_b0_carry[9]), .A2(n1614), .ZN(
        sub_434_b0_carry[10]) );
  XOR2_X1 U1362 ( .A(n1614), .B(sub_434_b0_carry[9]), .Z(N115) );
  AND2_X1 U1363 ( .A1(sub_434_b0_carry[8]), .A2(n1615), .ZN(
        sub_434_b0_carry[9]) );
  XOR2_X1 U1364 ( .A(n1615), .B(sub_434_b0_carry[8]), .Z(N114) );
  AND2_X1 U1365 ( .A1(sub_434_b0_carry[7]), .A2(n1616), .ZN(
        sub_434_b0_carry[8]) );
  XOR2_X1 U1366 ( .A(n1616), .B(sub_434_b0_carry[7]), .Z(N113) );
  AND2_X1 U1367 ( .A1(sub_434_b0_carry[6]), .A2(n1617), .ZN(
        sub_434_b0_carry[7]) );
  XOR2_X1 U1368 ( .A(n1617), .B(sub_434_b0_carry[6]), .Z(N112) );
  AND2_X1 U1369 ( .A1(sub_434_b0_carry[5]), .A2(n1612), .ZN(
        sub_434_b0_carry[6]) );
  XOR2_X1 U1370 ( .A(n1612), .B(sub_434_b0_carry[5]), .Z(N111) );
  AND2_X1 U1371 ( .A1(sub_434_b0_carry[4]), .A2(n1613), .ZN(
        sub_434_b0_carry[5]) );
  XOR2_X1 U1372 ( .A(n1613), .B(sub_434_b0_carry[4]), .Z(N110) );
  AND2_X1 U1373 ( .A1(sub_434_b0_carry[3]), .A2(n1589), .ZN(
        sub_434_b0_carry[4]) );
  AND2_X1 U1374 ( .A1(sub_434_b0_carry[2]), .A2(n1590), .ZN(
        sub_434_b0_carry[3]) );
  AND2_X1 U1375 ( .A1(n1599), .A2(n1591), .ZN(sub_434_b0_carry[2]) );
  INV_X4 U1376 ( .A(sub_1_root_u1_sub_128_aco_B_0_), .ZN(n1638) );
  INV_X4 U1377 ( .A(sub_1_root_u1_sub_128_aco_B_1_), .ZN(n1639) );
  INV_X4 U1378 ( .A(sub_1_root_u1_sub_128_aco_B_2_), .ZN(n1640) );
  INV_X4 U1379 ( .A(u1_exp_small[3]), .ZN(n1641) );
  INV_X4 U1380 ( .A(u1_exp_small[4]), .ZN(n1642) );
  INV_X4 U1381 ( .A(u2_sub_110_carry[5]), .ZN(u2_N11) );
  XOR2_X1 U1382 ( .A(u2_add_113_carry[4]), .B(u2_add_113_A_4_), .Z(
        u2_exp_tmp3_4_) );
  INV_X4 U1383 ( .A(u2_lt_130_A_0_), .ZN(u2_exp_tmp4_0_) );
  INV_X4 U1384 ( .A(u2_lt_130_A_1_), .ZN(u2_exp_tmp4_1_) );
  INV_X4 U1385 ( .A(u2_lt_130_A_2_), .ZN(u2_exp_tmp4_2_) );
  INV_X4 U1386 ( .A(u2_lt_130_A_3_), .ZN(u2_exp_tmp4_3_) );
  XOR2_X1 U1387 ( .A(u2_add_115_carry[4]), .B(u2_exp_tmp4_4_), .Z(u2_N34) );
  NOR2_X1 U1388 ( .A1(u2_exp_tmp4_1_), .A2(u2_exp_tmp4_0_), .ZN(n1644) );
  AOI21_X1 U1389 ( .B1(u2_exp_tmp4_0_), .B2(u2_exp_tmp4_1_), .A(n1644), .ZN(
        n1643) );
  NAND2_X1 U1390 ( .A1(n1644), .A2(u2_lt_130_A_2_), .ZN(n1645) );
  OAI21_X1 U1391 ( .B1(n1644), .B2(u2_lt_130_A_2_), .A(n1645), .ZN(u2_N37) );
  XNOR2_X1 U1392 ( .A(u2_exp_tmp4_3_), .B(n1645), .ZN(u2_N38) );
  NOR2_X1 U1393 ( .A1(u2_exp_tmp4_3_), .A2(n1645), .ZN(n1646) );
  XOR2_X1 U1394 ( .A(u2_exp_tmp4_4_), .B(n1646), .Z(u2_N39) );
  INV_X4 U1395 ( .A(n1643), .ZN(u2_N36) );
  INV_X4 U1396 ( .A(u4_sub_406_carry[5]), .ZN(u4_div_scht1a[5]) );
  NOR2_X1 U1397 ( .A1(n1891), .A2(n1627), .ZN(n1648) );
  AOI21_X1 U1398 ( .B1(n1626), .B2(n1891), .A(n1648), .ZN(n1647) );
  NAND2_X1 U1399 ( .A1(n1648), .A2(n1782), .ZN(n1649) );
  OAI21_X1 U1400 ( .B1(n1648), .B2(n1782), .A(n1649), .ZN(u4_exp_in_mi1_2_) );
  XNOR2_X1 U1401 ( .A(n1533), .B(n1649), .ZN(u4_exp_in_mi1_3_) );
  NOR3_X1 U1402 ( .A1(n1533), .A2(exp_r[4]), .A3(n1649), .ZN(u4_exp_in_mi1_5_)
         );
  OAI21_X1 U1403 ( .B1(n1533), .B2(n1649), .A(exp_r[4]), .ZN(n1650) );
  NAND2_X1 U1404 ( .A1(n2179), .A2(n1650), .ZN(u4_exp_in_mi1_4_) );
  INV_X4 U1405 ( .A(n1647), .ZN(u4_exp_in_mi1_1_) );
  INV_X4 U1406 ( .A(n1626), .ZN(u4_exp_in_pl1_0_) );
  INV_X4 U1407 ( .A(u4_ldz_all_1_), .ZN(n1653) );
  INV_X4 U1408 ( .A(u4_ldz_all_2_), .ZN(n1654) );
  INV_X4 U1409 ( .A(u4_ldz_all_3_), .ZN(n1655) );
  INV_X4 U1410 ( .A(u4_ldz_all_4_), .ZN(n1656) );
  NOR2_X1 U1411 ( .A1(u4_N264), .A2(u4_fi_ldz_2a_0_), .ZN(n1658) );
  AOI21_X1 U1412 ( .B1(u4_fi_ldz_2a_0_), .B2(u4_N264), .A(n1658), .ZN(n1657)
         );
  NAND2_X1 U1413 ( .A1(n1658), .A2(n2362), .ZN(n1659) );
  OAI21_X1 U1414 ( .B1(n1658), .B2(n2362), .A(n1659), .ZN(u4_fi_ldz_mi1_2_) );
  XNOR2_X1 U1415 ( .A(u4_N152), .B(n1659), .ZN(u4_fi_ldz_mi1_3_) );
  NOR3_X1 U1416 ( .A1(u4_N152), .A2(u4_N95), .A3(n1659), .ZN(u4_fi_ldz_mi1_6_)
         );
  OAI21_X1 U1417 ( .B1(u4_N152), .B2(n1659), .A(u4_N95), .ZN(n1660) );
  NAND2_X1 U1418 ( .A1(n1661), .A2(n1660), .ZN(u4_fi_ldz_mi1_4_) );
  INV_X4 U1419 ( .A(u4_fi_ldz_mi1_6_), .ZN(n1661) );
  INV_X4 U1420 ( .A(n1657), .ZN(u4_fi_ldz_mi1_1_) );
  NOR2_X1 U1421 ( .A1(u4_sub_465_A_1_), .A2(u4_sub_465_A_0_), .ZN(n1663) );
  AOI21_X1 U1422 ( .B1(u4_sub_465_A_0_), .B2(u4_sub_465_A_1_), .A(n1663), .ZN(
        n1662) );
  NAND2_X1 U1423 ( .A1(n1663), .A2(n850), .ZN(n1664) );
  OAI21_X1 U1424 ( .B1(n1663), .B2(n850), .A(n1664), .ZN(u4_exp_out1_mi1[2])
         );
  XNOR2_X1 U1425 ( .A(u4_sub_465_A_3_), .B(n1664), .ZN(u4_exp_out1_mi1[3]) );
  NOR2_X1 U1426 ( .A1(u4_sub_465_A_3_), .A2(n1664), .ZN(n1665) );
  XOR2_X1 U1427 ( .A(u4_sub_465_A_4_), .B(n1665), .Z(u4_exp_out1_mi1[4]) );
  INV_X4 U1428 ( .A(u4_sub_465_A_0_), .ZN(u4_exp_out1_mi1[0]) );
  INV_X4 U1429 ( .A(n1662), .ZN(u4_exp_out1_mi1[1]) );
  INV_X4 U1430 ( .A(n1627), .ZN(u4_f2i_shft_0_) );
  INV_X4 U1431 ( .A(u4_N152), .ZN(n1666) );
  INV_X4 U1432 ( .A(u4_fi_ldz_2a_0_), .ZN(n1667) );
  INV_X4 U1433 ( .A(n1627), .ZN(n1668) );
  XOR2_X1 U1434 ( .A(u4_add_461_carry[4]), .B(u4_exp_out_4_), .Z(
        u4_exp_out_pl1_4_) );
  NOR2_X1 U1435 ( .A1(u4_exp_out_1_), .A2(u4_exp_out_0_), .ZN(n1670) );
  AOI21_X1 U1436 ( .B1(u4_exp_out_0_), .B2(u4_exp_out_1_), .A(n1670), .ZN(
        n1669) );
  INV_X1 U1437 ( .A(n1669), .ZN(u4_exp_out_mi1[1]) );
  NAND2_X1 U1438 ( .A1(n1670), .A2(n1867), .ZN(n1671) );
  OAI21_X1 U1439 ( .B1(n1670), .B2(n1867), .A(n1671), .ZN(u4_exp_out_mi1[2])
         );
  XNOR2_X1 U1440 ( .A(u4_exp_out_3_), .B(n1671), .ZN(u4_exp_out_mi1[3]) );
  NOR2_X1 U1441 ( .A1(u4_exp_out_3_), .A2(n1671), .ZN(n1672) );
  XOR2_X1 U1442 ( .A(u4_exp_out_4_), .B(n1672), .Z(u4_exp_out_mi1[4]) );
  INV_X4 U1443 ( .A(u4_fi_ldz_mi1_4_), .ZN(n1674) );
  INV_X4 U1444 ( .A(u4_fi_ldz_mi1_3_), .ZN(n1675) );
  INV_X4 U1445 ( .A(u4_fi_ldz_mi1_2_), .ZN(n1676) );
  AND2_X1 U1446 ( .A1(opb_r[10]), .A2(n1580), .ZN(n1677) );
  OAI22_X1 U1447 ( .A1(n1677), .A2(n1578), .B1(opb_r[11]), .B2(n1677), .ZN(
        n1678) );
  OAI21_X1 U1448 ( .B1(opa_r[14]), .B2(n1582), .A(n1678), .ZN(n1686) );
  NAND2_X1 U1449 ( .A1(opb_r[13]), .A2(n1579), .ZN(n1682) );
  NOR2_X1 U1450 ( .A1(n1580), .A2(opb_r[10]), .ZN(n1680) );
  OAI21_X1 U1451 ( .B1(n1687), .B2(n1578), .A(opb_r[11]), .ZN(n1679) );
  NAND2_X1 U1452 ( .A1(opb_r[12]), .A2(n1547), .ZN(n1685) );
  OAI211_X1 U1453 ( .C1(opa_r[11]), .C2(n1680), .A(n1679), .B(n1685), .ZN(
        n1681) );
  OAI221_X1 U1454 ( .B1(opb_r[12]), .B2(n1547), .C1(opb_r[13]), .C2(n1579), 
        .A(n1681), .ZN(n1683) );
  OAI211_X1 U1455 ( .C1(opa_r[14]), .C2(n1582), .A(n1683), .B(n1682), .ZN(
        n1684) );
  NOR4_X1 U1456 ( .A1(n1686), .A2(n1689), .A3(n1624), .A4(n1688), .ZN(u1_N32)
         );
  INV_X4 U1457 ( .A(n1680), .ZN(n1687) );
  INV_X4 U1458 ( .A(n1685), .ZN(n1688) );
  INV_X4 U1459 ( .A(n1682), .ZN(n1689) );
  AND2_X1 U1460 ( .A1(fracta_mul[0]), .A2(n1838), .ZN(n1690) );
  OAI22_X1 U1461 ( .A1(fracta_mul[1]), .A2(n1690), .B1(n1690), .B2(n1839), 
        .ZN(n1692) );
  NAND2_X1 U1462 ( .A1(fracta_mul[7]), .A2(n1845), .ZN(n1693) );
  NAND2_X1 U1463 ( .A1(fracta_mul[5]), .A2(n1843), .ZN(n1701) );
  NAND2_X1 U1464 ( .A1(fracta_mul[6]), .A2(n1844), .ZN(n1702) );
  AND2_X1 U1465 ( .A1(n1701), .A2(n1702), .ZN(n1691) );
  OR2_X1 U1466 ( .A1(n1855), .A2(u6_N8), .ZN(n1694) );
  NAND4_X1 U1467 ( .A1(n1692), .A2(n1693), .A3(n1691), .A4(n1694), .ZN(n1712)
         );
  NAND2_X1 U1468 ( .A1(fracta_mul[9]), .A2(n1846), .ZN(n1708) );
  AND2_X1 U1469 ( .A1(n1694), .A2(n1693), .ZN(n1705) );
  NAND2_X1 U1470 ( .A1(fracta_mul[4]), .A2(n1842), .ZN(n1710) );
  NAND2_X1 U1471 ( .A1(fracta_mul[3]), .A2(n1841), .ZN(n1709) );
  NOR2_X1 U1472 ( .A1(n1838), .A2(fracta_mul[0]), .ZN(n1696) );
  OAI21_X1 U1473 ( .B1(fracta_mul[1]), .B2(n1713), .A(n1839), .ZN(n1695) );
  NAND2_X1 U1474 ( .A1(fracta_mul[2]), .A2(n1840), .ZN(n1707) );
  OAI211_X1 U1475 ( .C1(n1696), .C2(n1848), .A(n1695), .B(n1707), .ZN(n1697)
         );
  OAI221_X1 U1476 ( .B1(fracta_mul[2]), .B2(n1840), .C1(fracta_mul[3]), .C2(
        n1841), .A(n1697), .ZN(n1698) );
  NAND3_X1 U1477 ( .A1(n1710), .A2(n1709), .A3(n1698), .ZN(n1699) );
  OAI221_X1 U1478 ( .B1(fracta_mul[4]), .B2(n1842), .C1(fracta_mul[5]), .C2(
        n1843), .A(n1699), .ZN(n1700) );
  NAND3_X1 U1479 ( .A1(n1702), .A2(n1701), .A3(n1700), .ZN(n1703) );
  OAI221_X1 U1480 ( .B1(fracta_mul[6]), .B2(n1844), .C1(fracta_mul[7]), .C2(
        n1845), .A(n1703), .ZN(n1704) );
  AOI22_X1 U1481 ( .A1(u6_N8), .A2(n1855), .B1(n1705), .B2(n1704), .ZN(n1706)
         );
  OAI22_X1 U1482 ( .A1(fracta_mul[9]), .A2(n1846), .B1(n1716), .B2(n1706), 
        .ZN(u1_N123) );
  NAND3_X1 U1483 ( .A1(n1708), .A2(n1717), .A3(n1707), .ZN(n1711) );
  NOR4_X1 U1484 ( .A1(n1712), .A2(n1711), .A3(n1714), .A4(n1715), .ZN(u1_N124)
         );
  INV_X4 U1485 ( .A(n1696), .ZN(n1713) );
  INV_X4 U1486 ( .A(n1709), .ZN(n1714) );
  INV_X4 U1487 ( .A(n1710), .ZN(n1715) );
  INV_X4 U1488 ( .A(n1708), .ZN(n1716) );
  INV_X4 U1489 ( .A(u1_N123), .ZN(n1717) );
  AND4_X1 U1490 ( .A1(u1_exp_diff_3_), .A2(u1_exp_diff_2_), .A3(u1_gt_144_B_0_), .A4(u1_exp_diff_1_), .ZN(n1718) );
  OR2_X1 U1491 ( .A1(n1718), .A2(u1_exp_diff_4_), .ZN(u1_exp_lt_27) );
  NOR2_X1 U1492 ( .A1(u1_gt_234_A_12_), .A2(n1751), .ZN(n1732) );
  NOR2_X1 U1493 ( .A1(n1734), .A2(u1_gt_234_A_0_), .ZN(n1719) );
  AOI21_X1 U1494 ( .B1(n1719), .B2(n1740), .A(u1_gt_234_B_1_), .ZN(n1720) );
  AOI221_X1 U1495 ( .B1(u1_gt_234_A_2_), .B2(n1735), .C1(u1_gt_234_A_1_), .C2(
        n1736), .A(n1720), .ZN(n1721) );
  AOI221_X1 U1496 ( .B1(u1_gt_234_B_3_), .B2(n1742), .C1(u1_gt_234_B_2_), .C2(
        n1741), .A(n1721), .ZN(n1722) );
  AOI221_X1 U1497 ( .B1(u1_gt_234_A_4_), .B2(n1754), .C1(u1_gt_234_A_3_), .C2(
        n1753), .A(n1722), .ZN(n1723) );
  AOI221_X1 U1498 ( .B1(u1_gt_234_B_5_), .B2(n1744), .C1(u1_gt_234_B_4_), .C2(
        n1743), .A(n1723), .ZN(n1724) );
  AOI221_X1 U1499 ( .B1(u1_gt_234_A_6_), .B2(n1756), .C1(u1_gt_234_A_5_), .C2(
        n1755), .A(n1724), .ZN(n1725) );
  AOI221_X1 U1500 ( .B1(u1_gt_234_B_7_), .B2(n1746), .C1(u1_gt_234_B_6_), .C2(
        n1745), .A(n1725), .ZN(n1726) );
  AOI221_X1 U1501 ( .B1(u1_gt_234_A_8_), .B2(n1758), .C1(u1_gt_234_A_7_), .C2(
        n1757), .A(n1726), .ZN(n1727) );
  AOI221_X1 U1502 ( .B1(u1_gt_234_B_9_), .B2(n1748), .C1(u1_gt_234_B_8_), .C2(
        n1747), .A(n1727), .ZN(n1728) );
  AOI221_X1 U1503 ( .B1(u1_gt_234_A_9_), .B2(n1759), .C1(u1_gt_234_A_10_), 
        .C2(n1749), .A(n1728), .ZN(n1729) );
  AOI221_X1 U1504 ( .B1(u1_gt_234_B_11_), .B2(n1738), .C1(u1_gt_234_B_10_), 
        .C2(n1737), .A(n1729), .ZN(n1730) );
  AOI221_X1 U1505 ( .B1(u1_gt_234_A_12_), .B2(n1751), .C1(u1_gt_234_A_11_), 
        .C2(n1750), .A(n1730), .ZN(n1731) );
  OAI22_X1 U1506 ( .A1(n1732), .A2(n1731), .B1(u1_gt_234_B_13_), .B2(n1739), 
        .ZN(n1733) );
  OAI21_X1 U1507 ( .B1(u1_gt_234_A_13_), .B2(n1752), .A(n1733), .ZN(
        u1_fractb_lt_fracta) );
  INV_X4 U1508 ( .A(u1_gt_234_B_0_), .ZN(n1734) );
  INV_X4 U1509 ( .A(u1_gt_234_B_2_), .ZN(n1735) );
  INV_X4 U1510 ( .A(n1719), .ZN(n1736) );
  INV_X4 U1511 ( .A(u1_gt_234_A_10_), .ZN(n1737) );
  INV_X4 U1512 ( .A(u1_gt_234_A_11_), .ZN(n1738) );
  INV_X4 U1513 ( .A(u1_gt_234_A_13_), .ZN(n1739) );
  INV_X4 U1514 ( .A(u1_gt_234_A_1_), .ZN(n1740) );
  INV_X4 U1515 ( .A(u1_gt_234_A_2_), .ZN(n1741) );
  INV_X4 U1516 ( .A(u1_gt_234_A_3_), .ZN(n1742) );
  INV_X4 U1517 ( .A(u1_gt_234_A_4_), .ZN(n1743) );
  INV_X4 U1518 ( .A(u1_gt_234_A_5_), .ZN(n1744) );
  INV_X4 U1519 ( .A(u1_gt_234_A_6_), .ZN(n1745) );
  INV_X4 U1520 ( .A(u1_gt_234_A_7_), .ZN(n1746) );
  INV_X4 U1521 ( .A(u1_gt_234_A_8_), .ZN(n1747) );
  INV_X4 U1522 ( .A(u1_gt_234_A_9_), .ZN(n1748) );
  INV_X4 U1523 ( .A(u1_gt_234_B_10_), .ZN(n1749) );
  INV_X4 U1524 ( .A(u1_gt_234_B_11_), .ZN(n1750) );
  INV_X4 U1525 ( .A(u1_gt_234_B_12_), .ZN(n1751) );
  INV_X4 U1526 ( .A(u1_gt_234_B_13_), .ZN(n1752) );
  INV_X4 U1527 ( .A(u1_gt_234_B_3_), .ZN(n1753) );
  INV_X4 U1528 ( .A(u1_gt_234_B_4_), .ZN(n1754) );
  INV_X4 U1529 ( .A(u1_gt_234_B_5_), .ZN(n1755) );
  INV_X4 U1530 ( .A(u1_gt_234_B_6_), .ZN(n1756) );
  INV_X4 U1531 ( .A(u1_gt_234_B_7_), .ZN(n1757) );
  INV_X4 U1532 ( .A(u1_gt_234_B_8_), .ZN(n1758) );
  INV_X4 U1533 ( .A(u1_gt_234_B_9_), .ZN(n1759) );
  OAI21_X1 U1534 ( .B1(u4_div_shft3_2_), .B2(u4_div_shft3_1_), .A(
        u4_div_shft3_3_), .ZN(n1760) );
  NAND2_X1 U1535 ( .A1(n1761), .A2(n1760), .ZN(u4_N326) );
  INV_X4 U1536 ( .A(u4_div_shft3_4_), .ZN(n1761) );
  AND4_X1 U1537 ( .A1(u4_div_exp1_0_), .A2(u4_div_exp1_1_), .A3(u4_div_exp1_3_), .A4(u4_div_exp1_2_), .ZN(n1762) );
  NOR2_X1 U1538 ( .A1(u4_div_exp1_4_), .A2(n1762), .ZN(u4_N487) );
  OAI21_X1 U1539 ( .B1(u4_ldz_all_2_), .B2(u4_ldz_all_1_), .A(u4_ldz_all_3_), 
        .ZN(n1763) );
  NOR3_X1 U1540 ( .A1(n1764), .A2(u4_ldz_all_5_), .A3(u4_ldz_all_4_), .ZN(
        u4_N558) );
  INV_X4 U1541 ( .A(n1763), .ZN(n1764) );
  OAI221_X1 U1542 ( .B1(n1631), .B2(n1857), .C1(n872), .C2(u4_N796), .A(n1858), 
        .ZN(u4_shift_right[4]) );
  NAND2_X1 U1543 ( .A1(u4_exp_in_mi1_4_), .A2(n1859), .ZN(n1858) );
  AOI222_X1 U1544 ( .A1(u4_div_shft3_4_), .A2(n1860), .B1(u4_div_shft4[4]), 
        .B2(n1861), .C1(u4_div_shft2[4]), .C2(n1862), .ZN(n1857) );
  OAI221_X1 U1545 ( .B1(n1531), .B2(n1863), .C1(n872), .C2(n1864), .A(n1865), 
        .ZN(u4_shift_right[3]) );
  NAND2_X1 U1546 ( .A1(u4_exp_in_mi1_3_), .A2(n1859), .ZN(n1865) );
  AOI222_X1 U1547 ( .A1(u4_div_shft3_3_), .A2(n1860), .B1(u4_div_shft4[3]), 
        .B2(n1861), .C1(u4_div_shft2[3]), .C2(n1862), .ZN(n1863) );
  OAI221_X1 U1548 ( .B1(n1631), .B2(n1866), .C1(n872), .C2(n1867), .A(n1868), 
        .ZN(u4_shift_right[2]) );
  NAND2_X1 U1549 ( .A1(u4_exp_in_mi1_2_), .A2(n1859), .ZN(n1868) );
  AOI222_X1 U1550 ( .A1(u4_div_shft3_2_), .A2(n1860), .B1(u4_div_shft4[2]), 
        .B2(n1861), .C1(u4_div_shft2[2]), .C2(n1862), .ZN(n1866) );
  OAI221_X1 U1551 ( .B1(n1531), .B2(n1869), .C1(n872), .C2(n1870), .A(n1871), 
        .ZN(u4_shift_right[1]) );
  NAND2_X1 U1552 ( .A1(u4_exp_in_mi1_1_), .A2(n1859), .ZN(n1871) );
  AOI222_X1 U1553 ( .A1(u4_div_shft3_1_), .A2(n1860), .B1(u4_div_shft4[1]), 
        .B2(n1861), .C1(n1784), .C2(n1862), .ZN(n1869) );
  NAND2_X1 U1554 ( .A1(n1872), .A2(n1873), .ZN(u4_shift_left[2]) );
  AOI222_X1 U1555 ( .A1(n1874), .A2(exp_r[2]), .B1(u4_div_scht1a[2]), .B2(
        n1875), .C1(n1876), .C2(div_opa_ldz_r2[2]), .ZN(n1873) );
  AOI222_X1 U1556 ( .A1(u4_f2i_shft_2_), .A2(n1877), .B1(u4_N203), .B2(n1878), 
        .C1(u4_exp_in_pl1_2_), .C2(n1879), .ZN(n1872) );
  NAND2_X1 U1557 ( .A1(n1880), .A2(n1881), .ZN(u4_shift_left[1]) );
  AOI221_X1 U1558 ( .B1(u4_div_scht1a[1]), .B2(n1875), .C1(n1876), .C2(
        div_opa_ldz_r2[1]), .A(n1882), .ZN(n1881) );
  OAI33_X1 U1559 ( .A1(n1883), .A2(n1884), .A3(n1885), .B1(n1886), .B2(n1887), 
        .B3(n1888), .ZN(n1882) );
  OAI21_X1 U1560 ( .B1(u4_exp_in_pl1_1_), .B2(n1889), .A(n1890), .ZN(n1886) );
  INV_X1 U1561 ( .A(u4_exp_in_pl1_1_), .ZN(n1883) );
  AOI222_X1 U1562 ( .A1(u4_f2i_shft_1_), .A2(n1877), .B1(n1874), .B2(n1891), 
        .C1(u4_N264), .C2(n1878), .ZN(n1880) );
  NAND2_X1 U1563 ( .A1(n1892), .A2(n1893), .ZN(u4_shift_left[0]) );
  AOI222_X1 U1564 ( .A1(n1874), .A2(n1894), .B1(u4_div_scht1a[0]), .B2(n1875), 
        .C1(n1876), .C2(div_opa_ldz_r2[0]), .ZN(n1893) );
  NOR2_X1 U1565 ( .A1(n1895), .A2(n1896), .ZN(n1876) );
  NOR2_X1 U1566 ( .A1(n1895), .A2(n1889), .ZN(n1875) );
  AOI222_X1 U1567 ( .A1(u4_f2i_shft_0_), .A2(n1877), .B1(u4_fi_ldz_2a_0_), 
        .B2(n1878), .C1(u4_exp_in_pl1_0_), .C2(n1879), .ZN(n1892) );
  INV_X1 U1568 ( .A(n1897), .ZN(u4_fract_out_9_) );
  INV_X1 U1569 ( .A(n1898), .ZN(u4_fract_out_8_) );
  INV_X1 U1570 ( .A(n1899), .ZN(u4_fract_out_7_) );
  INV_X1 U1571 ( .A(n1900), .ZN(u4_fract_out_1_) );
  AOI21_X1 U1572 ( .B1(n1903), .B2(n1904), .A(fract_denorm[19]), .ZN(n1901) );
  INV_X1 U1573 ( .A(fract_denorm[18]), .ZN(n1904) );
  OAI21_X1 U1574 ( .B1(fract_denorm[16]), .B2(n1905), .A(n1906), .ZN(n1903) );
  INV_X1 U1575 ( .A(fract_denorm[17]), .ZN(n1906) );
  AOI21_X1 U1576 ( .B1(n1907), .B2(n1908), .A(fract_denorm[15]), .ZN(n1905) );
  OAI21_X1 U1577 ( .B1(fract_denorm[12]), .B2(n1909), .A(n1910), .ZN(n1907) );
  AOI21_X1 U1578 ( .B1(n1911), .B2(n1912), .A(fract_denorm[11]), .ZN(n1909) );
  OAI21_X1 U1579 ( .B1(fract_denorm[8]), .B2(n1913), .A(n1914), .ZN(n1911) );
  AOI21_X1 U1580 ( .B1(n1915), .B2(n1916), .A(n2704), .ZN(n1913) );
  OAI21_X1 U1581 ( .B1(n2710), .B2(n1917), .A(n1918), .ZN(n1915) );
  AOI21_X1 U1582 ( .B1(n2705), .B2(n1919), .A(n2711), .ZN(n1917) );
  NOR2_X1 U1583 ( .A1(n1920), .A2(n1921), .ZN(u2_underflow_d[2]) );
  MUX2_X1 U1584 ( .A(n1922), .B(n1923), .S(n1924), .Z(n1921) );
  NAND4_X1 U1585 ( .A1(u2_N15), .A2(u2_N14), .A3(n1925), .A4(u2_N13), .ZN(
        n1923) );
  NOR2_X1 U1586 ( .A1(u2_N16), .A2(n1926), .ZN(n1925) );
  INV_X1 U1587 ( .A(u2_N12), .ZN(n1926) );
  NAND4_X1 U1588 ( .A1(u2_N9), .A2(u2_N8), .A3(n1927), .A4(u2_N7), .ZN(n1922)
         );
  NOR2_X1 U1589 ( .A1(u2_N10), .A2(n1928), .ZN(n1927) );
  INV_X1 U1590 ( .A(u2_N6), .ZN(n1928) );
  INV_X1 U1591 ( .A(n1929), .ZN(u2_underflow_d[1]) );
  AOI221_X1 U1592 ( .B1(n1522), .B2(n1930), .C1(n1523), .C2(n1931), .A(n1932), 
        .ZN(n1929) );
  AOI21_X1 U1593 ( .B1(n1577), .B2(n1582), .A(n1920), .ZN(n1932) );
  OAI22_X1 U1594 ( .A1(u6_N10), .A2(n1931), .B1(n2698), .B2(n1930), .ZN(n1920)
         );
  AND3_X1 U1595 ( .A1(n1933), .A2(n1934), .A3(n1935), .ZN(u2_underflow_d[0])
         );
  NOR2_X1 U1596 ( .A1(n1577), .A2(n1936), .ZN(u2_exp_ovf_d_0_) );
  MUX2_X1 U1597 ( .A(n1937), .B(n1924), .S(n1582), .Z(n1936) );
  NAND2_X1 U1598 ( .A1(n1938), .A2(n1924), .ZN(n1937) );
  NOR2_X1 U1599 ( .A1(n1554), .A2(n1594), .ZN(u2_N73) );
  MUX2_X1 U1600 ( .A(n1939), .B(n1940), .S(n1924), .Z(u2_N66) );
  NOR2_X1 U1601 ( .A1(n1933), .A2(n1935), .ZN(n1940) );
  INV_X1 U1602 ( .A(u2_gt_140_B_5_), .ZN(n1935) );
  MUX2_X1 U1603 ( .A(u2_N17), .B(u2_N11), .S(n1941), .Z(u2_gt_140_B_5_) );
  NOR2_X1 U1604 ( .A1(u2_exp_tmp4_4_), .A2(n1942), .ZN(n1933) );
  AND4_X1 U1605 ( .A1(u2_lt_130_A_3_), .A2(u2_lt_130_A_2_), .A3(u2_lt_130_A_0_), .A4(u2_lt_130_A_1_), .ZN(n1942) );
  MUX2_X1 U1606 ( .A(u2_N13), .B(u2_N7), .S(n1941), .Z(u2_lt_130_A_1_) );
  MUX2_X1 U1607 ( .A(u2_N12), .B(u2_N6), .S(n1941), .Z(u2_lt_130_A_0_) );
  MUX2_X1 U1608 ( .A(u2_N14), .B(u2_N8), .S(n1941), .Z(u2_lt_130_A_2_) );
  MUX2_X1 U1609 ( .A(u2_N15), .B(u2_N9), .S(n1941), .Z(u2_lt_130_A_3_) );
  MUX2_X1 U1610 ( .A(u2_N10), .B(u2_N16), .S(n1924), .Z(u2_exp_tmp4_4_) );
  NOR2_X1 U1611 ( .A1(opa_r[14]), .A2(u6_N10), .ZN(n1939) );
  OAI211_X1 U1612 ( .C1(n1943), .C2(n1944), .A(n1945), .B(n1946), .ZN(u2_N44)
         );
  AOI22_X1 U1613 ( .A1(u2_exp_tmp4_4_), .A2(n1947), .B1(u2_exp_tmp3_4_), .B2(
        n1948), .ZN(n1946) );
  AOI22_X1 U1614 ( .A1(u2_N39), .A2(n1949), .B1(u2_N34), .B2(n1950), .ZN(n1945) );
  OAI211_X1 U1615 ( .C1(n1951), .C2(n1944), .A(n1952), .B(n1953), .ZN(u2_N43)
         );
  AOI22_X1 U1616 ( .A1(u2_exp_tmp4_3_), .A2(n1947), .B1(u2_exp_tmp3_3_), .B2(
        n1948), .ZN(n1953) );
  AOI22_X1 U1617 ( .A1(u2_N38), .A2(n1949), .B1(u2_N33), .B2(n1950), .ZN(n1952) );
  INV_X1 U1618 ( .A(u2_add_113_A_3_), .ZN(n1951) );
  OAI211_X1 U1619 ( .C1(n1954), .C2(n1944), .A(n1955), .B(n1956), .ZN(u2_N42)
         );
  AOI22_X1 U1620 ( .A1(u2_exp_tmp4_2_), .A2(n1947), .B1(u2_exp_tmp3_2_), .B2(
        n1948), .ZN(n1956) );
  AOI22_X1 U1621 ( .A1(u2_N37), .A2(n1949), .B1(u2_N32), .B2(n1950), .ZN(n1955) );
  INV_X1 U1622 ( .A(u2_add_113_A_2_), .ZN(n1954) );
  OAI211_X1 U1623 ( .C1(n1957), .C2(n1944), .A(n1958), .B(n1959), .ZN(u2_N41)
         );
  AOI22_X1 U1624 ( .A1(u2_exp_tmp4_1_), .A2(n1947), .B1(u2_exp_tmp3_1_), .B2(
        n1948), .ZN(n1959) );
  AOI22_X1 U1625 ( .A1(u2_N36), .A2(n1949), .B1(u2_N31), .B2(n1950), .ZN(n1958) );
  INV_X1 U1626 ( .A(u2_add_113_A_1_), .ZN(n1957) );
  OAI211_X1 U1627 ( .C1(n1960), .C2(n1944), .A(n1961), .B(n1962), .ZN(u2_N40)
         );
  AOI22_X1 U1628 ( .A1(u2_exp_tmp4_0_), .A2(n1947), .B1(n1960), .B2(n1948), 
        .ZN(n1962) );
  NOR2_X1 U1629 ( .A1(n1934), .A2(u2_exp_ovf_d_1_), .ZN(n1948) );
  INV_X1 U1630 ( .A(n1963), .ZN(u2_exp_ovf_d_1_) );
  NOR2_X1 U1631 ( .A1(n1963), .A2(sub_1_root_u1_sub_128_aco_CI), .ZN(n1947) );
  AOI22_X1 U1632 ( .A1(u2_lt_130_A_0_), .A2(n1949), .B1(u2_lt_130_A_0_), .B2(
        n1950), .ZN(n1961) );
  AND3_X1 U1633 ( .A1(n1941), .A2(sub_1_root_u1_sub_128_aco_CI), .A3(n1938), 
        .ZN(n1950) );
  NOR3_X1 U1634 ( .A1(n1941), .A2(n1934), .A3(n1963), .ZN(n1949) );
  NAND2_X1 U1635 ( .A1(n1934), .A2(n1963), .ZN(n1944) );
  NOR2_X1 U1636 ( .A1(n1938), .A2(n1964), .ZN(n1963) );
  NOR4_X1 U1637 ( .A1(n1943), .A2(n1941), .A3(opa_r[14]), .A4(opb_r[14]), .ZN(
        n1964) );
  INV_X1 U1638 ( .A(u2_add_113_A_4_), .ZN(n1943) );
  MUX2_X1 U1639 ( .A(u2_N29), .B(u2_N23), .S(n1941), .Z(n1938) );
  INV_X1 U1640 ( .A(u2_add_113_A_0_), .ZN(n1960) );
  MUX2_X1 U1641 ( .A(opa_r[15]), .B(n1965), .S(n1633), .Z(u1_sign_d) );
  XNOR2_X1 U1642 ( .A(n1554), .B(fpu_op_r1[0]), .ZN(n1965) );
  MUX2_X1 U1643 ( .A(u1_gt_234_B_9_), .B(u1_gt_234_A_9_), .S(n1633), .Z(
        u1_fractb_s[9]) );
  MUX2_X1 U1644 ( .A(u1_gt_234_B_8_), .B(u1_gt_234_A_8_), .S(n1633), .Z(
        u1_fractb_s[8]) );
  MUX2_X1 U1645 ( .A(u1_gt_234_B_7_), .B(u1_gt_234_A_7_), .S(n1633), .Z(
        u1_fractb_s[7]) );
  MUX2_X1 U1646 ( .A(u1_gt_234_B_6_), .B(u1_gt_234_A_6_), .S(n1633), .Z(
        u1_fractb_s[6]) );
  MUX2_X1 U1647 ( .A(u1_gt_234_B_5_), .B(u1_gt_234_A_5_), .S(n1633), .Z(
        u1_fractb_s[5]) );
  MUX2_X1 U1648 ( .A(u1_gt_234_B_4_), .B(u1_gt_234_A_4_), .S(n1633), .Z(
        u1_fractb_s[4]) );
  MUX2_X1 U1649 ( .A(u1_gt_234_B_3_), .B(u1_gt_234_A_3_), .S(n1633), .Z(
        u1_fractb_s[3]) );
  MUX2_X1 U1650 ( .A(u1_gt_234_B_2_), .B(u1_gt_234_A_2_), .S(n1633), .Z(
        u1_fractb_s[2]) );
  MUX2_X1 U1651 ( .A(u1_gt_234_B_1_), .B(u1_gt_234_A_1_), .S(n1633), .Z(
        u1_fractb_s[1]) );
  MUX2_X1 U1652 ( .A(u1_gt_234_B_13_), .B(u1_gt_234_A_13_), .S(n1633), .Z(
        u1_fractb_s[13]) );
  MUX2_X1 U1653 ( .A(u1_gt_234_B_12_), .B(u1_gt_234_A_12_), .S(
        u1_fractb_lt_fracta), .Z(u1_fractb_s[12]) );
  MUX2_X1 U1654 ( .A(u1_gt_234_B_11_), .B(u1_gt_234_A_11_), .S(
        u1_fractb_lt_fracta), .Z(u1_fractb_s[11]) );
  MUX2_X1 U1655 ( .A(u1_gt_234_B_10_), .B(u1_gt_234_A_10_), .S(
        u1_fractb_lt_fracta), .Z(u1_fractb_s[10]) );
  MUX2_X1 U1656 ( .A(u1_gt_234_B_0_), .B(u1_gt_234_A_0_), .S(n1633), .Z(
        u1_fractb_s[0]) );
  MUX2_X1 U1657 ( .A(u1_gt_234_A_9_), .B(u1_gt_234_B_9_), .S(
        u1_fractb_lt_fracta), .Z(u1_fracta_s[9]) );
  MUX2_X1 U1658 ( .A(u1_gt_234_A_8_), .B(u1_gt_234_B_8_), .S(
        u1_fractb_lt_fracta), .Z(u1_fracta_s[8]) );
  MUX2_X1 U1659 ( .A(u1_gt_234_A_7_), .B(u1_gt_234_B_7_), .S(
        u1_fractb_lt_fracta), .Z(u1_fracta_s[7]) );
  MUX2_X1 U1660 ( .A(u1_gt_234_A_6_), .B(u1_gt_234_B_6_), .S(
        u1_fractb_lt_fracta), .Z(u1_fracta_s[6]) );
  MUX2_X1 U1661 ( .A(u1_gt_234_A_5_), .B(u1_gt_234_B_5_), .S(
        u1_fractb_lt_fracta), .Z(u1_fracta_s[5]) );
  MUX2_X1 U1662 ( .A(u1_gt_234_A_4_), .B(u1_gt_234_B_4_), .S(
        u1_fractb_lt_fracta), .Z(u1_fracta_s[4]) );
  MUX2_X1 U1663 ( .A(u1_gt_234_A_3_), .B(u1_gt_234_B_3_), .S(n1633), .Z(
        u1_fracta_s[3]) );
  MUX2_X1 U1664 ( .A(u1_gt_234_A_2_), .B(u1_gt_234_B_2_), .S(n1633), .Z(
        u1_fracta_s[2]) );
  MUX2_X1 U1665 ( .A(u1_gt_234_A_1_), .B(u1_gt_234_B_1_), .S(n1633), .Z(
        u1_fracta_s[1]) );
  MUX2_X1 U1666 ( .A(u1_gt_234_A_13_), .B(u1_gt_234_B_13_), .S(n1633), .Z(
        u1_fracta_s[13]) );
  MUX2_X1 U1667 ( .A(u1_gt_234_A_12_), .B(u1_gt_234_B_12_), .S(n1633), .Z(
        u1_fracta_s[12]) );
  MUX2_X1 U1668 ( .A(u1_gt_234_A_11_), .B(u1_gt_234_B_11_), .S(n1633), .Z(
        u1_fracta_s[11]) );
  MUX2_X1 U1669 ( .A(u1_gt_234_A_10_), .B(u1_gt_234_B_10_), .S(n1633), .Z(
        u1_fracta_s[10]) );
  MUX2_X1 U1670 ( .A(u1_gt_234_A_0_), .B(u1_gt_234_B_0_), .S(
        u1_fractb_lt_fracta), .Z(u1_fracta_s[0]) );
  MUX2_X1 U1671 ( .A(opb_r[14]), .B(opa_r[14]), .S(n1629), .Z(u1_exp_small[4])
         );
  MUX2_X1 U1672 ( .A(opb_r[13]), .B(opa_r[13]), .S(n1966), .Z(u1_exp_small[3])
         );
  AND2_X1 U1673 ( .A1(u1_exp_diff2[4]), .A2(n1967), .ZN(u1_exp_diff_4_) );
  INV_X1 U1674 ( .A(n1968), .ZN(u1_exp_diff_2_) );
  NOR2_X1 U1675 ( .A1(n1969), .A2(n1970), .ZN(u1_N39) );
  NOR2_X1 U1676 ( .A1(n1969), .A2(n1971), .ZN(u1_N38) );
  INV_X1 U1677 ( .A(sub_1_root_u1_sub_128_aco_A_3_), .ZN(n1971) );
  NOR2_X1 U1678 ( .A1(n1969), .A2(n1972), .ZN(u1_N37) );
  INV_X1 U1679 ( .A(sub_1_root_u1_sub_128_aco_A_2_), .ZN(n1972) );
  NOR2_X1 U1680 ( .A1(n1969), .A2(n1973), .ZN(u1_N36) );
  INV_X1 U1681 ( .A(sub_1_root_u1_sub_128_aco_A_1_), .ZN(n1973) );
  NOR2_X1 U1682 ( .A1(n1969), .A2(n1974), .ZN(u1_N35) );
  INV_X1 U1683 ( .A(sub_1_root_u1_sub_128_aco_A_0_), .ZN(n1974) );
  AND3_X1 U1684 ( .A1(n1975), .A2(u1_N124), .A3(u1_N32), .ZN(n1969) );
  OAI21_X1 U1685 ( .B1(n1976), .B2(n1593), .A(n1977), .ZN(u1_N133) );
  OAI21_X1 U1686 ( .B1(n1978), .B2(n1610), .A(u1_signa_r), .ZN(n1977) );
  NOR3_X1 U1687 ( .A1(n1600), .A2(u1_fracta_lt_fractb), .A3(
        u1_fracta_eq_fractb), .ZN(n1978) );
  AOI21_X1 U1688 ( .B1(opb_nan), .B2(n1979), .A(u1_signa_r), .ZN(n1976) );
  OAI21_X1 U1689 ( .B1(u1_fracta_eq_fractb), .B2(n1609), .A(opa_nan), .ZN(
        n1979) );
  OAI22_X1 U1690 ( .A1(n1608), .A2(n1980), .B1(n1981), .B2(n1982), .ZN(u1_N122) );
  XNOR2_X1 U1691 ( .A(n1593), .B(u1_add_r), .ZN(n1982) );
  NOR2_X1 U1692 ( .A1(n1983), .A2(u1_signa_r), .ZN(n1981) );
  NAND2_X1 U1693 ( .A1(n1984), .A2(n1985), .ZN(u0_N7) );
  NOR2_X1 U1694 ( .A1(n1985), .A2(n1984), .ZN(u0_N6) );
  NOR2_X1 U1695 ( .A1(n1986), .A2(u6_N9), .ZN(u0_N5) );
  NOR2_X1 U1696 ( .A1(n1987), .A2(fracta_mul[9]), .ZN(u0_N4) );
  NOR2_X1 U1697 ( .A1(n1825), .A2(n1827), .ZN(u0_N17) );
  NOR2_X1 U1698 ( .A1(n1824), .A2(n1826), .ZN(u0_N16) );
  NOR2_X1 U1699 ( .A1(n2701), .A2(n1988), .ZN(u0_N11) );
  NOR2_X1 U1700 ( .A1(n2699), .A2(n1989), .ZN(u0_N10) );
  MUX2_X1 U1701 ( .A(N76), .B(fracta_mul[9]), .S(n2698), .Z(u6_N22) );
  MUX2_X1 U1702 ( .A(fracta_mul[8]), .B(N75), .S(n1522), .Z(u6_N21) );
  MUX2_X1 U1703 ( .A(fracta_mul[7]), .B(N74), .S(n1522), .Z(u6_N20) );
  MUX2_X1 U1704 ( .A(fracta_mul[6]), .B(N73), .S(n1522), .Z(u6_N19) );
  MUX2_X1 U1705 ( .A(fracta_mul[5]), .B(N72), .S(n1522), .Z(u6_N18) );
  MUX2_X1 U1706 ( .A(fracta_mul[4]), .B(N71), .S(n1522), .Z(u6_N17) );
  MUX2_X1 U1707 ( .A(fracta_mul[3]), .B(N70), .S(n1522), .Z(u6_N16) );
  MUX2_X1 U1708 ( .A(fracta_mul[2]), .B(N69), .S(n1522), .Z(u6_N15) );
  MUX2_X1 U1709 ( .A(N68), .B(fracta_mul[1]), .S(n2698), .Z(u6_N14) );
  MUX2_X1 U1710 ( .A(N67), .B(fracta_mul[0]), .S(n2698), .Z(u6_N13) );
  OAI22_X1 U1711 ( .A1(n1990), .A2(n1589), .B1(n1991), .B2(n1605), .ZN(n2666)
         );
  OAI22_X1 U1712 ( .A1(n1990), .A2(n1590), .B1(n1991), .B2(n1606), .ZN(n2667)
         );
  OAI22_X1 U1713 ( .A1(n1990), .A2(n1591), .B1(n1991), .B2(n1607), .ZN(n2668)
         );
  MUX2_X1 U1714 ( .A(u2_N22), .B(u2_N28), .S(n1924), .Z(u2_add_113_A_4_) );
  MUX2_X1 U1715 ( .A(u2_N21), .B(u2_N27), .S(n1924), .Z(u2_add_113_A_3_) );
  MUX2_X1 U1716 ( .A(u2_N26), .B(u2_N20), .S(n1941), .Z(u2_add_113_A_2_) );
  MUX2_X1 U1717 ( .A(u2_N19), .B(u2_N25), .S(n1924), .Z(u2_add_113_A_1_) );
  MUX2_X1 U1718 ( .A(u2_exp_tmp4_0_), .B(u2_exp_tmp4_0_), .S(n1941), .Z(
        u2_add_113_A_0_) );
  MUX2_X1 U1719 ( .A(u3_N17), .B(u3_N32), .S(n1815), .Z(n2669) );
  MUX2_X1 U1720 ( .A(u3_N16), .B(u3_N31), .S(n1815), .Z(n2670) );
  MUX2_X1 U1721 ( .A(u3_N15), .B(u3_N30), .S(n1815), .Z(n2671) );
  MUX2_X1 U1722 ( .A(u3_N14), .B(u3_N29), .S(n1815), .Z(n2672) );
  MUX2_X1 U1723 ( .A(u3_N13), .B(u3_N28), .S(n1815), .Z(n2673) );
  MUX2_X1 U1724 ( .A(u3_N12), .B(u3_N27), .S(n1815), .Z(n2674) );
  MUX2_X1 U1725 ( .A(u3_N11), .B(u3_N26), .S(n1815), .Z(n2675) );
  MUX2_X1 U1726 ( .A(u3_N10), .B(u3_N25), .S(n1815), .Z(n2676) );
  MUX2_X1 U1727 ( .A(u3_N9), .B(u3_N24), .S(n1815), .Z(n2677) );
  MUX2_X1 U1728 ( .A(u3_N8), .B(u3_N23), .S(n1815), .Z(n2678) );
  MUX2_X1 U1729 ( .A(u3_N7), .B(u3_N22), .S(n1815), .Z(n2679) );
  MUX2_X1 U1730 ( .A(u3_N6), .B(u3_N21), .S(n1815), .Z(n2680) );
  MUX2_X1 U1731 ( .A(u3_N5), .B(u3_N20), .S(n1815), .Z(n2681) );
  MUX2_X1 U1732 ( .A(u3_N4), .B(u3_N19), .S(n1815), .Z(n2682) );
  MUX2_X1 U1733 ( .A(u3_N3), .B(u3_N18), .S(n1815), .Z(n2683) );
  MUX2_X1 U1734 ( .A(u4_exp_in_pl1_1_), .B(u4_exp_next_mi_1_), .S(n1902), .Z(
        u4_sub_465_A_1_) );
  INV_X1 U1735 ( .A(n1975), .ZN(n2684) );
  XOR2_X1 U1736 ( .A(fpu_op_r1[0]), .B(u2_sign_d), .Z(n1975) );
  XNOR2_X1 U1737 ( .A(n1594), .B(opb_r[15]), .ZN(u2_sign_d) );
  MUX2_X1 U1738 ( .A(u1_adj_op_out_sft_9_), .B(u6_N6), .S(n1966), .Z(
        u1_gt_234_B_9_) );
  MUX2_X1 U1739 ( .A(u1_adj_op_out_sft_8_), .B(u6_N5), .S(n1966), .Z(
        u1_gt_234_B_8_) );
  MUX2_X1 U1740 ( .A(u1_adj_op_out_sft_7_), .B(u6_N4), .S(n1966), .Z(
        u1_gt_234_B_7_) );
  MUX2_X1 U1741 ( .A(u1_adj_op_out_sft_6_), .B(u6_N3), .S(n1966), .Z(
        u1_gt_234_B_6_) );
  MUX2_X1 U1742 ( .A(u1_adj_op_out_sft_5_), .B(u6_N2), .S(n1966), .Z(
        u1_gt_234_B_5_) );
  MUX2_X1 U1743 ( .A(u1_adj_op_out_sft_4_), .B(u6_N1), .S(n1966), .Z(
        u1_gt_234_B_4_) );
  MUX2_X1 U1744 ( .A(u1_adj_op_out_sft_3_), .B(u6_N0), .S(n1966), .Z(
        u1_gt_234_B_3_) );
  MUX2_X1 U1745 ( .A(u1_adj_op_out_sft_13_), .B(u6_N10), .S(n1966), .Z(
        u1_gt_234_B_13_) );
  MUX2_X1 U1746 ( .A(u1_adj_op_out_sft_12_), .B(u6_N9), .S(n1966), .Z(
        u1_gt_234_B_12_) );
  MUX2_X1 U1747 ( .A(u1_adj_op_out_sft_11_), .B(u6_N8), .S(n1629), .Z(
        u1_gt_234_B_11_) );
  MUX2_X1 U1748 ( .A(u6_N7), .B(u1_adj_op_out_sft_10_), .S(n1624), .Z(
        u1_gt_234_B_10_) );
  MUX2_X1 U1749 ( .A(fracta_mul[6]), .B(u1_adj_op_out_sft_9_), .S(n1629), .Z(
        u1_gt_234_A_9_) );
  MUX2_X1 U1750 ( .A(fracta_mul[5]), .B(u1_adj_op_out_sft_8_), .S(n1629), .Z(
        u1_gt_234_A_8_) );
  MUX2_X1 U1751 ( .A(fracta_mul[4]), .B(u1_adj_op_out_sft_7_), .S(n1629), .Z(
        u1_gt_234_A_7_) );
  MUX2_X1 U1752 ( .A(fracta_mul[3]), .B(u1_adj_op_out_sft_6_), .S(n1629), .Z(
        u1_gt_234_A_6_) );
  MUX2_X1 U1753 ( .A(fracta_mul[2]), .B(u1_adj_op_out_sft_5_), .S(n1629), .Z(
        u1_gt_234_A_5_) );
  MUX2_X1 U1754 ( .A(fracta_mul[1]), .B(u1_adj_op_out_sft_4_), .S(n1629), .Z(
        u1_gt_234_A_4_) );
  MUX2_X1 U1755 ( .A(fracta_mul[0]), .B(u1_adj_op_out_sft_3_), .S(n1629), .Z(
        u1_gt_234_A_3_) );
  AND2_X1 U1756 ( .A1(u1_adj_op_out_sft_2_), .A2(n1629), .ZN(u1_gt_234_A_2_)
         );
  AND2_X1 U1757 ( .A1(u1_adj_op_out_sft_1_), .A2(n1966), .ZN(u1_gt_234_A_1_)
         );
  MUX2_X1 U1758 ( .A(n2698), .B(u1_adj_op_out_sft_13_), .S(n1629), .Z(
        u1_gt_234_A_13_) );
  MUX2_X1 U1759 ( .A(fracta_mul[9]), .B(u1_adj_op_out_sft_12_), .S(n1629), .Z(
        u1_gt_234_A_12_) );
  MUX2_X1 U1760 ( .A(fracta_mul[8]), .B(u1_adj_op_out_sft_11_), .S(n1629), .Z(
        u1_gt_234_A_11_) );
  MUX2_X1 U1761 ( .A(u1_adj_op_out_sft_10_), .B(fracta_mul[7]), .S(n1624), .Z(
        u1_gt_234_A_10_) );
  AND2_X1 U1762 ( .A1(n1992), .A2(n1629), .ZN(u1_gt_234_A_0_) );
  AND2_X1 U1763 ( .A1(u1_adj_op_out_sft_2_), .A2(n1624), .ZN(u1_gt_234_B_2_)
         );
  AND2_X1 U1764 ( .A1(u1_adj_op_out_sft_1_), .A2(n1630), .ZN(u1_gt_234_B_1_)
         );
  AND2_X1 U1765 ( .A1(n1624), .A2(n1992), .ZN(u1_gt_234_B_0_) );
  OR2_X1 U1766 ( .A1(u1_adj_op_out_sft_0_), .A2(n1993), .ZN(n1992) );
  MUX2_X1 U1767 ( .A(n1994), .B(n1995), .S(n2686), .Z(n1993) );
  MUX2_X1 U1768 ( .A(n1996), .B(n1997), .S(n2685), .Z(n1995) );
  AND2_X1 U1769 ( .A1(n1998), .A2(n1999), .ZN(n1997) );
  OAI21_X1 U1770 ( .B1(n2000), .B2(n2001), .A(n2002), .ZN(n1998) );
  OAI221_X1 U1771 ( .B1(n1999), .B2(n2003), .C1(n2000), .C2(n2004), .A(n2005), 
        .ZN(n1996) );
  AOI211_X1 U1772 ( .C1(u1_exp_diff_sft_0_), .C2(u1_adj_op_9_), .A(n2006), .B(
        n2688), .ZN(n2003) );
  INV_X1 U1773 ( .A(n2007), .ZN(n2006) );
  MUX2_X1 U1774 ( .A(fracta_mul[9]), .B(u6_N9), .S(n1624), .Z(u1_adj_op_9_) );
  NOR2_X1 U1775 ( .A1(n1999), .A2(n2008), .ZN(n1994) );
  AOI221_X1 U1776 ( .B1(n2009), .B2(n2685), .C1(u1_exp_diff_sft_0_), .C2(n2010), .A(n2011), .ZN(n2008) );
  OAI21_X1 U1777 ( .B1(n2012), .B2(n2007), .A(n2013), .ZN(n2010) );
  NOR2_X1 U1778 ( .A1(n2009), .A2(n2689), .ZN(n2007) );
  INV_X1 U1779 ( .A(n2000), .ZN(u1_exp_diff_sft_0_) );
  NAND2_X1 U1780 ( .A1(u1_gt_144_B_0_), .A2(n2014), .ZN(n2000) );
  OR3_X1 U1781 ( .A1(n2691), .A2(n2690), .A3(n2011), .ZN(n2009) );
  NAND2_X1 U1782 ( .A1(n2001), .A2(n2015), .ZN(n2011) );
  INV_X1 U1783 ( .A(n2692), .ZN(n2015) );
  NOR2_X1 U1784 ( .A1(n2016), .A2(n2693), .ZN(n2001) );
  INV_X1 U1785 ( .A(n2002), .ZN(n2016) );
  NOR3_X1 U1786 ( .A1(n2694), .A2(n2696), .A3(n2695), .ZN(n2002) );
  INV_X1 U1787 ( .A(n2012), .ZN(n2685) );
  NOR2_X1 U1788 ( .A1(u1_exp_diff_1_), .A2(u1_exp_lt_27), .ZN(n2012) );
  AND2_X1 U1789 ( .A1(u1_exp_diff2[1]), .A2(n1967), .ZN(u1_exp_diff_1_) );
  NAND2_X1 U1790 ( .A1(n1968), .A2(n2014), .ZN(n2686) );
  INV_X1 U1791 ( .A(u1_exp_lt_27), .ZN(n2014) );
  NAND2_X1 U1792 ( .A1(u1_exp_diff2[2]), .A2(n1967), .ZN(n1968) );
  INV_X1 U1793 ( .A(n1999), .ZN(n2687) );
  NOR2_X1 U1794 ( .A1(u1_exp_diff_3_), .A2(u1_exp_lt_27), .ZN(n1999) );
  AND2_X1 U1795 ( .A1(u1_exp_diff2[3]), .A2(n1967), .ZN(u1_exp_diff_3_) );
  MUX2_X1 U1796 ( .A(opa_r[12]), .B(opb_r[12]), .S(n1624), .Z(
        sub_1_root_u1_sub_128_aco_B_2_) );
  MUX2_X1 U1797 ( .A(opa_r[11]), .B(opb_r[11]), .S(n1624), .Z(
        sub_1_root_u1_sub_128_aco_B_1_) );
  AND2_X1 U1798 ( .A1(u1_exp_diff2[0]), .A2(n1967), .ZN(u1_gt_144_B_0_) );
  NAND2_X1 U1799 ( .A1(n1523), .A2(n1522), .ZN(n1967) );
  MUX2_X1 U1800 ( .A(opa_r[10]), .B(opb_r[10]), .S(u1_expa_lt_expb), .Z(
        sub_1_root_u1_sub_128_aco_B_0_) );
  MUX2_X1 U1801 ( .A(fracta_mul[8]), .B(u6_N8), .S(n1630), .Z(n2688) );
  MUX2_X1 U1802 ( .A(fracta_mul[7]), .B(u6_N7), .S(n1624), .Z(n2689) );
  MUX2_X1 U1803 ( .A(fracta_mul[6]), .B(u6_N6), .S(n1624), .Z(n2690) );
  INV_X1 U1804 ( .A(n2013), .ZN(n2691) );
  MUX2_X1 U1805 ( .A(n1843), .B(n1852), .S(n1629), .Z(n2013) );
  MUX2_X1 U1806 ( .A(u6_N4), .B(fracta_mul[4]), .S(n1629), .Z(n2692) );
  MUX2_X1 U1807 ( .A(fracta_mul[3]), .B(u6_N3), .S(n1630), .Z(n2693) );
  MUX2_X1 U1808 ( .A(fracta_mul[2]), .B(u6_N2), .S(n1624), .Z(n2694) );
  INV_X1 U1809 ( .A(n2004), .ZN(n2695) );
  MUX2_X1 U1810 ( .A(n1848), .B(n1839), .S(n1624), .Z(n2004) );
  INV_X1 U1811 ( .A(n2005), .ZN(n2696) );
  MUX2_X1 U1812 ( .A(n1838), .B(n1847), .S(n1629), .Z(n2005) );
  INV_X1 U1813 ( .A(n1970), .ZN(sub_1_root_u1_sub_128_aco_A_4_) );
  MUX2_X1 U1814 ( .A(n1577), .B(n1582), .S(n1966), .Z(n1970) );
  INV_X1 U1815 ( .A(n1624), .ZN(n1966) );
  MUX2_X1 U1816 ( .A(opb_r[13]), .B(opa_r[13]), .S(n1624), .Z(
        sub_1_root_u1_sub_128_aco_A_3_) );
  MUX2_X1 U1817 ( .A(opb_r[12]), .B(opa_r[12]), .S(n1624), .Z(
        sub_1_root_u1_sub_128_aco_A_2_) );
  MUX2_X1 U1818 ( .A(opb_r[11]), .B(opa_r[11]), .S(n1624), .Z(
        sub_1_root_u1_sub_128_aco_A_1_) );
  MUX2_X1 U1819 ( .A(opb_r[10]), .B(opa_r[10]), .S(u1_expa_lt_expb), .Z(
        sub_1_root_u1_sub_128_aco_A_0_) );
  INV_X1 U1820 ( .A(n1989), .ZN(n2697) );
  NAND4_X1 U1821 ( .A1(opa_r[13]), .A2(opa_r[14]), .A3(opa_r[12]), .A4(n2017), 
        .ZN(n1989) );
  NOR2_X1 U1822 ( .A1(n1578), .A2(n1580), .ZN(n2017) );
  INV_X1 U1823 ( .A(n1934), .ZN(sub_1_root_u1_sub_128_aco_CI) );
  NOR2_X1 U1824 ( .A1(n1522), .A2(n1523), .ZN(n1934) );
  INV_X1 U1825 ( .A(n1930), .ZN(n2699) );
  NAND2_X1 U1826 ( .A1(n1856), .A2(n1987), .ZN(n1930) );
  AND4_X1 U1827 ( .A1(n1854), .A2(n1849), .A3(n1855), .A4(n2018), .ZN(n1987)
         );
  NOR3_X1 U1828 ( .A1(fracta_mul[1]), .A2(n2019), .A3(fracta_mul[0]), .ZN(
        n2018) );
  INV_X1 U1829 ( .A(n1988), .ZN(n2700) );
  NAND4_X1 U1830 ( .A1(opb_r[13]), .A2(opb_r[14]), .A3(opb_r[12]), .A4(n2020), 
        .ZN(n1988) );
  NOR2_X1 U1831 ( .A1(n1587), .A2(n1588), .ZN(n2020) );
  INV_X1 U1832 ( .A(n1931), .ZN(n2701) );
  NAND2_X1 U1833 ( .A1(n1846), .A2(n1986), .ZN(n1931) );
  AND4_X1 U1834 ( .A1(n1842), .A2(n1841), .A3(n2021), .A4(n2022), .ZN(n1986)
         );
  NOR4_X1 U1835 ( .A1(u6_N5), .A2(u6_N6), .A3(u6_N7), .A4(u6_N8), .ZN(n2022)
         );
  NOR3_X1 U1836 ( .A1(u6_N2), .A2(u6_N0), .A3(u6_N1), .ZN(n2021) );
  OAI22_X1 U1837 ( .A1(n1990), .A2(n1599), .B1(n1991), .B2(n1599), .ZN(n2703)
         );
  INV_X1 U1838 ( .A(n2023), .ZN(n2710) );
  INV_X1 U1839 ( .A(n2024), .ZN(n2711) );
  OAI22_X1 U1840 ( .A1(n1596), .A2(n1822), .B1(n1555), .B2(n1820), .ZN(n2712)
         );
  OAI22_X1 U1841 ( .A1(n1596), .A2(n1821), .B1(n1555), .B2(n1819), .ZN(n2713)
         );
  INV_X1 U1842 ( .A(n1984), .ZN(n2714) );
  NAND2_X1 U1843 ( .A1(u0_infb_f_r), .A2(u0_expb_ff), .ZN(n1984) );
  INV_X1 U1844 ( .A(n1985), .ZN(n2715) );
  NAND2_X1 U1845 ( .A1(u0_infa_f_r), .A2(u0_expa_ff), .ZN(n1985) );
  NAND2_X1 U1846 ( .A1(n1668), .A2(n1859), .ZN(n889) );
  NOR2_X1 U1847 ( .A1(n2025), .A2(n1632), .ZN(n1859) );
  AOI222_X1 U1848 ( .A1(n1626), .A2(n1862), .B1(u4_div_shft4[0]), .B2(n1861), 
        .C1(u4_div_shft3_0_), .C2(n1860), .ZN(n888) );
  NOR2_X1 U1849 ( .A1(n2026), .A2(n1860), .ZN(n1861) );
  INV_X1 U1850 ( .A(n2027), .ZN(n1860) );
  NAND2_X1 U1851 ( .A1(n2025), .A2(n1531), .ZN(n872) );
  AOI221_X1 U1852 ( .B1(u4_exp_f2i_1[25]), .B2(n2028), .C1(u4_N445), .C2(n2029), .A(n2030), .ZN(n852) );
  NOR2_X1 U1853 ( .A1(n2031), .A2(n2032), .ZN(n2030) );
  AOI222_X1 U1854 ( .A1(u4_div_exp1_2_), .A2(opb_dn), .B1(u4_exp_out1_mi1[2]), 
        .B2(n2033), .C1(u4_div_exp2[2]), .C2(n2034), .ZN(n2031) );
  AOI21_X1 U1855 ( .B1(u4_div_exp3[2]), .B2(n842), .A(n2035), .ZN(n851) );
  INV_X1 U1856 ( .A(u4_sub_465_A_2_), .ZN(n850) );
  MUX2_X1 U1857 ( .A(u4_exp_in_pl1_2_), .B(u4_exp_next_mi_2_), .S(n1902), .Z(
        u4_sub_465_A_2_) );
  INV_X1 U1858 ( .A(u6_N10), .ZN(n1523) );
  MUX2_X1 U1859 ( .A(n2698), .B(u6_N10), .S(n1624), .Z(n1521) );
  NAND3_X1 U1860 ( .A1(n1588), .A2(n1587), .A3(n2036), .ZN(u6_N10) );
  NOR3_X1 U1861 ( .A1(opb_r[12]), .A2(opb_r[14]), .A3(opb_r[13]), .ZN(n2036)
         );
  OR2_X1 U1862 ( .A1(N77), .A2(n2698), .ZN(u6_N23) );
  NOR3_X1 U1863 ( .A1(opa_r[12]), .A2(opa_r[14]), .A3(opa_r[13]), .ZN(n2037)
         );
  OAI222_X1 U1864 ( .A1(n1809), .A2(n2038), .B1(n1781), .B2(n2039), .C1(n2040), 
        .C2(n1621), .ZN(N99) );
  OAI222_X1 U1865 ( .A1(n1810), .A2(n2038), .B1(n2041), .B2(n1622), .C1(n1835), 
        .C2(n1783), .ZN(N98) );
  OAI222_X1 U1866 ( .A1(n1811), .A2(n2038), .B1(n2041), .B2(n1618), .C1(n1835), 
        .C2(n1785), .ZN(N97) );
  OAI222_X1 U1867 ( .A1(n1812), .A2(n2038), .B1(n2041), .B2(n1619), .C1(n1835), 
        .C2(n1787), .ZN(N96) );
  OAI21_X1 U1868 ( .B1(n2042), .B2(fracta_mul[8]), .A(n1856), .ZN(N65) );
  AOI21_X1 U1869 ( .B1(n1853), .B2(n2043), .A(fracta_mul[7]), .ZN(n2042) );
  OAI21_X1 U1870 ( .B1(n2044), .B2(fracta_mul[4]), .A(n1852), .ZN(n2043) );
  AOI21_X1 U1871 ( .B1(n1849), .B2(fracta_mul[1]), .A(fracta_mul[3]), .ZN(
        n2044) );
  NOR2_X1 U1872 ( .A1(n2045), .A2(fracta_mul[9]), .ZN(N56) );
  AOI211_X1 U1873 ( .C1(n2046), .C2(n1853), .A(fracta_mul[8]), .B(
        fracta_mul[7]), .ZN(n2045) );
  AOI21_X1 U1874 ( .B1(n2047), .B2(n1851), .A(fracta_mul[5]), .ZN(n2046) );
  AOI21_X1 U1875 ( .B1(n1849), .B2(n1848), .A(fracta_mul[3]), .ZN(n2047) );
  NOR2_X1 U1876 ( .A1(n2048), .A2(n2049), .ZN(N44) );
  INV_X1 U1877 ( .A(n2019), .ZN(n2048) );
  NOR2_X1 U1878 ( .A1(n2019), .A2(n2049), .ZN(N34) );
  NAND3_X1 U1879 ( .A1(n1855), .A2(n1854), .A3(n1856), .ZN(n2049) );
  NAND4_X1 U1880 ( .A1(n1853), .A2(n1852), .A3(n1851), .A4(n1850), .ZN(n2019)
         );
  NOR4_X1 U1881 ( .A1(n2050), .A2(n1783), .A3(n1787), .A4(n1785), .ZN(N296) );
  OR2_X1 U1882 ( .A1(n1779), .A2(n1781), .ZN(n2050) );
  NOR4_X1 U1883 ( .A1(opa_inf), .A2(opa_00), .A3(n1823), .A4(n1553), .ZN(N292)
         );
  NOR3_X1 U1884 ( .A1(n2039), .A2(opa_nan), .A3(n1834), .ZN(N291) );
  OAI22_X1 U1885 ( .A1(n1887), .A2(n2051), .B1(n2052), .B2(n2053), .ZN(N290)
         );
  NOR3_X1 U1886 ( .A1(n2054), .A2(n2055), .A3(n2056), .ZN(n2052) );
  NOR4_X1 U1887 ( .A1(opb_inf), .A2(opb_00), .A3(n1631), .A4(n2057), .ZN(n2056) );
  AOI21_X1 U1888 ( .B1(n2058), .B2(n2059), .A(opa_inf), .ZN(n2054) );
  OR4_X1 U1889 ( .A1(n2060), .A2(n2057), .A3(n1885), .A4(opb_inf), .ZN(n2059)
         );
  OAI21_X1 U1890 ( .B1(n1553), .B2(n1592), .A(n2061), .ZN(n2058) );
  AOI21_X1 U1891 ( .B1(n2062), .B2(n2063), .A(n2053), .ZN(N285) );
  NAND3_X1 U1892 ( .A1(n2064), .A2(n1597), .A3(n2065), .ZN(n2063) );
  NAND2_X1 U1893 ( .A1(n1628), .A2(n2066), .ZN(n2062) );
  NAND4_X1 U1894 ( .A1(n2067), .A2(n2068), .A3(n2069), .A4(n2070), .ZN(n2066)
         );
  NAND4_X1 U1895 ( .A1(n2071), .A2(n2072), .A3(n2073), .A4(n2074), .ZN(n2069)
         );
  NOR4_X1 U1896 ( .A1(n2075), .A2(n2076), .A3(n2077), .A4(n2078), .ZN(n2074)
         );
  NOR4_X1 U1897 ( .A1(n2079), .A2(n2080), .A3(n2081), .A4(n2082), .ZN(n2073)
         );
  NAND3_X1 U1898 ( .A1(n1632), .A2(n1549), .A3(opa_inf), .ZN(n2068) );
  NAND2_X1 U1899 ( .A1(n2083), .A2(n1592), .ZN(n2067) );
  AND2_X1 U1900 ( .A1(n2084), .A2(n1628), .ZN(N283) );
  OAI33_X1 U1901 ( .A1(n2085), .A2(n1831), .A3(n2086), .B1(n2087), .B2(n2088), 
        .B3(n1604), .ZN(N281) );
  AOI221_X1 U1902 ( .B1(underflow_fmul_r[2]), .B2(n2089), .C1(
        underflow_fmul_r[1]), .C2(n2090), .A(n2091), .ZN(n2088) );
  OAI21_X1 U1903 ( .B1(n2092), .B2(n2093), .A(n1790), .ZN(n2091) );
  OR2_X1 U1904 ( .A1(n2057), .A2(n1581), .ZN(n2093) );
  OAI21_X1 U1905 ( .B1(n2094), .B2(n2095), .A(n2096), .ZN(n2092) );
  NAND4_X1 U1906 ( .A1(n1544), .A2(n1562), .A3(n2097), .A4(n2098), .ZN(n2095)
         );
  NOR4_X1 U1907 ( .A1(n2099), .A2(prod[14]), .A3(prod[16]), .A4(prod[15]), 
        .ZN(n2098) );
  NAND3_X1 U1908 ( .A1(n1534), .A2(n1545), .A3(n1563), .ZN(n2099) );
  NOR3_X1 U1909 ( .A1(prod[11]), .A2(prod[13]), .A3(prod[12]), .ZN(n2097) );
  NAND4_X1 U1910 ( .A1(n1537), .A2(n1561), .A3(n2100), .A4(n2101), .ZN(n2094)
         );
  NOR4_X1 U1911 ( .A1(n2102), .A2(prod[4]), .A3(prod[6]), .A4(prod[5]), .ZN(
        n2101) );
  OR3_X1 U1912 ( .A1(prod[8]), .A2(prod[9]), .A3(prod[7]), .ZN(n2102) );
  NOR3_X1 U1913 ( .A1(prod[21]), .A2(prod[3]), .A3(prod[2]), .ZN(n2100) );
  OAI33_X1 U1914 ( .A1(n2103), .A2(n2104), .A3(n2105), .B1(n2106), .B2(n2107), 
        .B3(n2108), .ZN(n2089) );
  NAND2_X1 U1915 ( .A1(n2109), .A2(n2110), .ZN(n2108) );
  NAND3_X1 U1916 ( .A1(n2111), .A2(n2112), .A3(n2113), .ZN(n2107) );
  NAND4_X1 U1917 ( .A1(n2114), .A2(n2115), .A3(n2116), .A4(n2117), .ZN(n2106)
         );
  NOR2_X1 U1918 ( .A1(n2080), .A2(n2081), .ZN(n2116) );
  NAND3_X1 U1919 ( .A1(n2078), .A2(n2079), .A3(n2077), .ZN(n2103) );
  INV_X1 U1920 ( .A(n2090), .ZN(n2086) );
  OAI21_X1 U1921 ( .B1(n2118), .B2(n2119), .A(n2120), .ZN(N278) );
  OR3_X1 U1922 ( .A1(n1560), .A2(n2121), .A3(n2085), .ZN(n2120) );
  AOI22_X1 U1923 ( .A1(n2122), .A2(n2123), .B1(n2124), .B2(n2060), .ZN(n2118)
         );
  OAI21_X1 U1924 ( .B1(n1560), .B2(n1536), .A(n2125), .ZN(n2123) );
  OAI221_X1 U1925 ( .B1(n2126), .B2(n2127), .C1(n1833), .C2(n2128), .A(n2129), 
        .ZN(N268) );
  NAND4_X1 U1926 ( .A1(n2130), .A2(n2124), .A3(n2131), .A4(n1592), .ZN(n2129)
         );
  NAND3_X1 U1927 ( .A1(n2070), .A2(n2057), .A3(n2132), .ZN(n2131) );
  AOI21_X1 U1928 ( .B1(n2133), .B2(n2060), .A(n2134), .ZN(n2132) );
  INV_X1 U1929 ( .A(n2126), .ZN(n2134) );
  NAND3_X1 U1930 ( .A1(n2124), .A2(n2135), .A3(n2136), .ZN(n2070) );
  NAND3_X1 U1931 ( .A1(n1595), .A2(n1549), .A3(n2137), .ZN(n2135) );
  INV_X1 U1932 ( .A(n2138), .ZN(n2128) );
  AOI22_X1 U1933 ( .A1(n2139), .A2(n2065), .B1(n2130), .B2(n1632), .ZN(n2127)
         );
  INV_X1 U1934 ( .A(n2085), .ZN(n2130) );
  NAND2_X1 U1935 ( .A1(n2139), .A2(n1553), .ZN(n2085) );
  INV_X1 U1936 ( .A(n2119), .ZN(n2139) );
  NOR3_X1 U1937 ( .A1(n2122), .A2(n2138), .A3(n2090), .ZN(n2126) );
  NAND3_X1 U1938 ( .A1(n2140), .A2(n2141), .A3(n2142), .ZN(n2090) );
  NAND3_X1 U1939 ( .A1(n2143), .A2(n2144), .A3(n2145), .ZN(n2142) );
  NAND4_X1 U1940 ( .A1(n2146), .A2(n1632), .A3(n2147), .A4(n2148), .ZN(n2141)
         );
  NOR3_X1 U1941 ( .A1(n2149), .A2(n2150), .A3(n2151), .ZN(n2148) );
  OAI22_X1 U1942 ( .A1(n2152), .A2(opb_dn), .B1(n2153), .B2(n1546), .ZN(n2147)
         );
  NAND4_X1 U1943 ( .A1(n2154), .A2(u4_N656), .A3(n1788), .A4(n2026), .ZN(n2146) );
  MUX2_X1 U1944 ( .A(n2155), .B(n2153), .S(n1789), .Z(n2154) );
  INV_X1 U1945 ( .A(n2156), .ZN(n2153) );
  OAI211_X1 U1946 ( .C1(n2157), .C2(n2158), .A(n2159), .B(n2160), .ZN(n2156)
         );
  OR4_X1 U1947 ( .A1(n2161), .A2(n1575), .A3(n2155), .A4(u4_N656), .ZN(n2160)
         );
  OAI211_X1 U1948 ( .C1(n2162), .C2(n2163), .A(n2164), .B(n2165), .ZN(n2159)
         );
  NOR3_X1 U1949 ( .A1(n1782), .A2(n1786), .A3(n1784), .ZN(n2162) );
  NOR2_X1 U1950 ( .A1(n2025), .A2(n2166), .ZN(n2158) );
  MUX2_X1 U1951 ( .A(n2167), .B(n2168), .S(n1777), .Z(n2166) );
  OAI221_X1 U1952 ( .B1(n2163), .B2(n2169), .C1(n2170), .C2(n2171), .A(n2172), 
        .ZN(n2168) );
  OAI211_X1 U1953 ( .C1(n2173), .C2(n2165), .A(n1782), .B(n1784), .ZN(n2172)
         );
  NOR4_X1 U1954 ( .A1(n2174), .A2(n1575), .A3(u4_N656), .A4(n2163), .ZN(n2173)
         );
  NAND2_X1 U1955 ( .A1(u4_N558), .A2(n2155), .ZN(n2174) );
  INV_X1 U1956 ( .A(n2165), .ZN(n2169) );
  NOR2_X1 U1957 ( .A1(n2161), .A2(n2027), .ZN(n2165) );
  NOR2_X1 U1958 ( .A1(n2175), .A2(n2170), .ZN(n2167) );
  NAND4_X1 U1959 ( .A1(n2124), .A2(n2176), .A3(n2177), .A4(n2178), .ZN(n2140)
         );
  NAND4_X1 U1960 ( .A1(n1896), .A2(n2179), .A3(n2180), .A4(n2181), .ZN(n2178)
         );
  NOR2_X1 U1961 ( .A1(n1575), .A2(n2182), .ZN(n2181) );
  INV_X1 U1962 ( .A(n2183), .ZN(n2180) );
  OAI211_X1 U1963 ( .C1(n1631), .C2(n2157), .A(n2184), .B(n2185), .ZN(n2138)
         );
  AOI222_X1 U1964 ( .A1(n2186), .A2(n2187), .B1(n1877), .B2(n2188), .C1(n2189), 
        .C2(n2177), .ZN(n2185) );
  OAI211_X1 U1965 ( .C1(n2190), .C2(n2191), .A(n2192), .B(n2152), .ZN(n2188)
         );
  INV_X1 U1966 ( .A(n2177), .ZN(n2152) );
  INV_X1 U1967 ( .A(n2121), .ZN(n2122) );
  MUX2_X1 U1968 ( .A(n2193), .B(n2194), .S(n1631), .Z(n2121) );
  NOR2_X1 U1969 ( .A1(n2195), .A2(n2196), .ZN(n2194) );
  INV_X1 U1970 ( .A(n2197), .ZN(n2196) );
  AOI211_X1 U1971 ( .C1(n2195), .C2(n2198), .A(n2199), .B(n2150), .ZN(n2193)
         );
  NAND2_X1 U1972 ( .A1(n2184), .A2(n2200), .ZN(n2199) );
  INV_X1 U1973 ( .A(n2149), .ZN(n2184) );
  OAI21_X1 U1974 ( .B1(n1777), .B2(n2155), .A(n1789), .ZN(n2198) );
  MUX2_X1 U1975 ( .A(n2201), .B(n2202), .S(n2055), .Z(N254) );
  NOR2_X1 U1976 ( .A1(n2057), .A2(n2203), .ZN(n2055) );
  NOR3_X1 U1977 ( .A1(n2053), .A2(n2204), .A3(n1573), .ZN(n2202) );
  MUX2_X1 U1978 ( .A(n2205), .B(n2206), .S(n2087), .Z(n2201) );
  NAND2_X1 U1979 ( .A1(n2207), .A2(n2124), .ZN(n2087) );
  MUX2_X1 U1980 ( .A(n2208), .B(n2209), .S(n2210), .Z(n2206) );
  NOR2_X1 U1981 ( .A1(n1531), .A2(n2053), .ZN(n2210) );
  MUX2_X1 U1982 ( .A(n2211), .B(n2212), .S(sign_mul_r), .Z(n2209) );
  OAI21_X1 U1983 ( .B1(n1553), .B2(n1592), .A(n2212), .ZN(n2211) );
  NAND3_X1 U1984 ( .A1(opa_inf), .A2(opb_inf), .A3(sign_exe_r), .ZN(n2212) );
  MUX2_X1 U1985 ( .A(nan_sign_d), .B(n2213), .S(n2214), .Z(n2208) );
  NOR2_X1 U1986 ( .A1(n2053), .A2(n1598), .ZN(n2214) );
  MUX2_X1 U1987 ( .A(result_zero_sign_d), .B(sign_fasu_r), .S(n2051), .Z(n2213) );
  OR2_X1 U1988 ( .A1(n2119), .A2(n2057), .ZN(n2051) );
  NAND4_X1 U1989 ( .A1(n2071), .A2(n2072), .A3(n2215), .A4(n2216), .ZN(n2057)
         );
  NOR4_X1 U1990 ( .A1(n2217), .A2(n2218), .A3(n2219), .A4(n2104), .ZN(n2216)
         );
  INV_X1 U1991 ( .A(n2076), .ZN(n2104) );
  NOR4_X1 U1992 ( .A1(n2105), .A2(n2080), .A3(n2081), .A4(n2082), .ZN(n2215)
         );
  INV_X1 U1993 ( .A(n2075), .ZN(n2105) );
  NOR4_X1 U1994 ( .A1(n2220), .A2(n2221), .A3(n2222), .A4(n2223), .ZN(n2072)
         );
  NOR3_X1 U1995 ( .A1(n2224), .A2(n2225), .A3(n2226), .ZN(n2071) );
  NAND2_X1 U1996 ( .A1(n1816), .A2(n2207), .ZN(n2119) );
  XOR2_X1 U1997 ( .A(sign_mul_r), .B(n2227), .Z(n2205) );
  NOR2_X1 U1998 ( .A1(n2136), .A2(n1611), .ZN(n2227) );
  NAND2_X1 U1999 ( .A1(n2228), .A2(n2076), .ZN(N234) );
  NAND2_X1 U2000 ( .A1(n2228), .A2(n2075), .ZN(N233) );
  NAND2_X1 U2001 ( .A1(n2228), .A2(n2078), .ZN(N232) );
  NAND2_X1 U2002 ( .A1(n2228), .A2(n2079), .ZN(N231) );
  NAND2_X1 U2003 ( .A1(n2228), .A2(n2077), .ZN(N230) );
  INV_X1 U2004 ( .A(n2229), .ZN(n2228) );
  OAI21_X1 U2005 ( .B1(n2230), .B2(n2229), .A(n2231), .ZN(N229) );
  INV_X1 U2006 ( .A(n2080), .ZN(n2230) );
  OAI221_X1 U2007 ( .B1(n1897), .B2(n2232), .C1(n2233), .C2(n2234), .A(n2235), 
        .ZN(n2080) );
  INV_X1 U2008 ( .A(u4_fract_out_pl1_9_), .ZN(n2234) );
  OAI21_X1 U2009 ( .B1(n2236), .B2(n2229), .A(n2231), .ZN(N228) );
  INV_X1 U2010 ( .A(n2081), .ZN(n2236) );
  OAI221_X1 U2011 ( .B1(n1898), .B2(n2232), .C1(n2233), .C2(n2237), .A(n2235), 
        .ZN(n2081) );
  INV_X1 U2012 ( .A(u4_fract_out_pl1_8_), .ZN(n2237) );
  OAI21_X1 U2013 ( .B1(n2117), .B2(n2229), .A(n2231), .ZN(N227) );
  INV_X1 U2014 ( .A(n2082), .ZN(n2117) );
  OAI221_X1 U2015 ( .B1(n1899), .B2(n2232), .C1(n2233), .C2(n2238), .A(n2235), 
        .ZN(n2082) );
  INV_X1 U2016 ( .A(u4_fract_out_pl1_7_), .ZN(n2238) );
  OAI21_X1 U2017 ( .B1(n2115), .B2(n2229), .A(n2231), .ZN(N226) );
  INV_X1 U2018 ( .A(n2220), .ZN(n2115) );
  OAI221_X1 U2019 ( .B1(n2239), .B2(n2232), .C1(n2233), .C2(n2240), .A(n2235), 
        .ZN(n2220) );
  INV_X1 U2020 ( .A(u4_fract_out_pl1_6_), .ZN(n2240) );
  NOR2_X1 U2021 ( .A1(n2114), .A2(n2229), .ZN(N225) );
  INV_X1 U2022 ( .A(n2221), .ZN(n2114) );
  OAI221_X1 U2023 ( .B1(n2241), .B2(n2232), .C1(n2233), .C2(n2242), .A(n2235), 
        .ZN(n2221) );
  INV_X1 U2024 ( .A(u4_fract_out_pl1_5_), .ZN(n2242) );
  NOR2_X1 U2025 ( .A1(n2112), .A2(n2229), .ZN(N224) );
  INV_X1 U2026 ( .A(n2222), .ZN(n2112) );
  OAI221_X1 U2027 ( .B1(n2243), .B2(n2232), .C1(n2233), .C2(n2244), .A(n2235), 
        .ZN(n2222) );
  INV_X1 U2028 ( .A(u4_fract_out_pl1_4_), .ZN(n2244) );
  NOR2_X1 U2029 ( .A1(n2111), .A2(n2229), .ZN(N223) );
  INV_X1 U2030 ( .A(n2223), .ZN(n2111) );
  OAI221_X1 U2031 ( .B1(n2245), .B2(n2232), .C1(n2233), .C2(n2246), .A(n2235), 
        .ZN(n2223) );
  INV_X1 U2032 ( .A(u4_fract_out_pl1_3_), .ZN(n2246) );
  NOR2_X1 U2033 ( .A1(n2113), .A2(n2229), .ZN(N222) );
  INV_X1 U2034 ( .A(n2225), .ZN(n2113) );
  OAI221_X1 U2035 ( .B1(n2247), .B2(n2232), .C1(n2233), .C2(n2248), .A(n2235), 
        .ZN(n2225) );
  INV_X1 U2036 ( .A(u4_fract_out_pl1_2_), .ZN(n2248) );
  NOR2_X1 U2037 ( .A1(n2110), .A2(n2229), .ZN(N221) );
  INV_X1 U2038 ( .A(n2226), .ZN(n2110) );
  OAI221_X1 U2039 ( .B1(n1900), .B2(n2232), .C1(n2233), .C2(n2249), .A(n2235), 
        .ZN(n2226) );
  INV_X1 U2040 ( .A(u4_fract_out_pl1_1_), .ZN(n2249) );
  OAI21_X1 U2041 ( .B1(n2109), .B2(n2229), .A(n2231), .ZN(N220) );
  NAND2_X1 U2042 ( .A1(n2229), .A2(n2084), .ZN(n2231) );
  OAI211_X1 U2043 ( .C1(n2136), .C2(n1885), .A(n2207), .B(n2250), .ZN(n2084)
         );
  AOI21_X1 U2044 ( .B1(n2083), .B2(opa_00), .A(n2251), .ZN(n2250) );
  INV_X1 U2045 ( .A(n2064), .ZN(n2251) );
  NAND2_X1 U2046 ( .A1(n1814), .A2(n1598), .ZN(n2064) );
  AOI22_X1 U2047 ( .A1(opb_inf), .A2(opa_00), .B1(opb_00), .B2(opa_inf), .ZN(
        n2136) );
  NAND2_X1 U2048 ( .A1(n1531), .A2(n1597), .ZN(n2253) );
  AOI211_X1 U2049 ( .C1(n2254), .C2(n2124), .A(n2255), .B(n2083), .ZN(n2252)
         );
  NOR2_X1 U2050 ( .A1(n1553), .A2(n1531), .ZN(n2083) );
  OAI21_X1 U2051 ( .B1(n1531), .B2(n1595), .A(n2207), .ZN(n2255) );
  INV_X1 U2052 ( .A(n2053), .ZN(n2207) );
  NAND2_X1 U2053 ( .A1(n1817), .A2(n1818), .ZN(n2053) );
  INV_X1 U2054 ( .A(n2137), .ZN(n2254) );
  NAND2_X1 U2055 ( .A1(n2256), .A2(n2060), .ZN(n2137) );
  NAND2_X1 U2056 ( .A1(n1791), .A2(n1778), .ZN(n2060) );
  INV_X1 U2057 ( .A(n2224), .ZN(n2109) );
  OAI221_X1 U2058 ( .B1(n2257), .B2(n2232), .C1(n2233), .C2(n2258), .A(n2235), 
        .ZN(n2224) );
  OAI21_X1 U2059 ( .B1(n2203), .B2(n2192), .A(n2261), .ZN(n2259) );
  NAND4_X1 U2060 ( .A1(n2262), .A2(n2263), .A3(n2187), .A4(n1631), .ZN(n2261)
         );
  OAI21_X1 U2061 ( .B1(n1548), .B2(n1581), .A(n2264), .ZN(n2263) );
  INV_X1 U2062 ( .A(u4_fract_out_pl1_0_), .ZN(n2258) );
  OAI22_X1 U2063 ( .A1(n2267), .A2(n2268), .B1(n2269), .B2(n1548), .ZN(n2266)
         );
  INV_X1 U2064 ( .A(n2270), .ZN(n2269) );
  OAI221_X1 U2065 ( .B1(n2272), .B2(n2268), .C1(n1548), .C2(n2270), .A(n2264), 
        .ZN(n2271) );
  AND3_X1 U2066 ( .A1(n2260), .A2(n2197), .A3(n2200), .ZN(n2265) );
  NAND4_X1 U2067 ( .A1(n2218), .A2(n2219), .A3(n2217), .A4(n2273), .ZN(n2197)
         );
  NOR4_X1 U2068 ( .A1(n1877), .A2(n2133), .A3(n2075), .A4(n2076), .ZN(n2273)
         );
  NAND2_X1 U2069 ( .A1(n2274), .A2(n2275), .ZN(n2076) );
  OAI211_X1 U2070 ( .C1(n1777), .C2(n2276), .A(n2277), .B(n2278), .ZN(n2275)
         );
  INV_X1 U2071 ( .A(n2279), .ZN(n2277) );
  NAND2_X1 U2072 ( .A1(n2274), .A2(n2280), .ZN(n2075) );
  NAND4_X1 U2073 ( .A1(n2281), .A2(n2282), .A3(n2283), .A4(n2284), .ZN(n2280)
         );
  AOI22_X1 U2074 ( .A1(u4_exp_out_pl1_3_), .A2(n2285), .B1(n2286), .B2(
        u4_exp_next_mi_3_), .ZN(n2284) );
  AOI22_X1 U2075 ( .A1(n2287), .A2(u4_exp_out_3_), .B1(u4_exp_fix_diva[3]), 
        .B2(n2288), .ZN(n2283) );
  AOI22_X1 U2076 ( .A1(u4_exp_fix_divb[3]), .A2(n2289), .B1(n2290), .B2(n2163), 
        .ZN(n2282) );
  AOI21_X1 U2077 ( .B1(u4_exp_out_mi1[3]), .B2(n2291), .A(n2292), .ZN(n2281)
         );
  INV_X1 U2078 ( .A(n2079), .ZN(n2217) );
  NAND2_X1 U2079 ( .A1(n2274), .A2(n2293), .ZN(n2079) );
  NAND4_X1 U2080 ( .A1(n2294), .A2(n2295), .A3(n2296), .A4(n2297), .ZN(n2293)
         );
  AOI22_X1 U2081 ( .A1(u4_exp_out_pl1_1_), .A2(n2285), .B1(n2286), .B2(
        u4_exp_next_mi_1_), .ZN(n2297) );
  AOI22_X1 U2082 ( .A1(n2287), .A2(u4_exp_out_1_), .B1(u4_exp_fix_diva[1]), 
        .B2(n2288), .ZN(n2296) );
  AOI22_X1 U2083 ( .A1(u4_exp_fix_divb[1]), .A2(n2289), .B1(n2290), .B2(n1891), 
        .ZN(n2295) );
  AOI21_X1 U2084 ( .B1(u4_exp_out_mi1[1]), .B2(n2291), .A(n2292), .ZN(n2294)
         );
  INV_X1 U2085 ( .A(n2077), .ZN(n2219) );
  OAI21_X1 U2086 ( .B1(n2298), .B2(n2299), .A(n2274), .ZN(n2077) );
  AOI21_X1 U2087 ( .B1(n2300), .B2(n2301), .A(n2292), .ZN(n2298) );
  AOI221_X1 U2088 ( .B1(n2302), .B2(u4_N581), .C1(n2303), .C2(n2304), .A(n2305), .ZN(n2301) );
  OAI22_X1 U2089 ( .A1(n2306), .A2(u4_N581), .B1(n2307), .B2(n2308), .ZN(n2305) );
  INV_X1 U2090 ( .A(u4_exp_next_mi_0_), .ZN(n2307) );
  MUX2_X1 U2091 ( .A(u4_exp_out_0_), .B(n2309), .S(n2310), .Z(n2304) );
  MUX2_X1 U2092 ( .A(u4_N581), .B(u4_N581), .S(n2311), .Z(n2309) );
  AOI21_X1 U2093 ( .B1(n2262), .B2(sign), .A(n1548), .ZN(n2303) );
  NOR2_X1 U2094 ( .A1(n2312), .A2(n2268), .ZN(n2302) );
  AOI222_X1 U2095 ( .A1(n2290), .A2(n1894), .B1(u4_exp_fix_diva[0]), .B2(n2288), .C1(u4_exp_fix_divb[0]), .C2(n2289), .ZN(n2300) );
  INV_X1 U2096 ( .A(n2078), .ZN(n2218) );
  NAND2_X1 U2097 ( .A1(n2274), .A2(n2313), .ZN(n2078) );
  NAND4_X1 U2098 ( .A1(n2314), .A2(n2315), .A3(n2316), .A4(n2317), .ZN(n2313)
         );
  AOI22_X1 U2099 ( .A1(u4_exp_out_pl1_2_), .A2(n2285), .B1(n2286), .B2(
        u4_exp_next_mi_2_), .ZN(n2317) );
  AOI22_X1 U2100 ( .A1(u4_exp_out_2_), .A2(n2287), .B1(u4_exp_fix_diva[2]), 
        .B2(n2288), .ZN(n2316) );
  AOI22_X1 U2101 ( .A1(u4_exp_fix_divb[2]), .A2(n2289), .B1(n2290), .B2(
        exp_r[2]), .ZN(n2315) );
  INV_X1 U2102 ( .A(n2276), .ZN(n2290) );
  NAND3_X1 U2103 ( .A1(n2133), .A2(n2318), .A3(n2195), .ZN(n2276) );
  AOI21_X1 U2104 ( .B1(u4_exp_out_mi1[2]), .B2(n2291), .A(n2292), .ZN(n2314)
         );
  INV_X1 U2105 ( .A(n2278), .ZN(n2292) );
  NOR2_X1 U2106 ( .A1(n2149), .A2(n2299), .ZN(n2278) );
  OAI211_X1 U2107 ( .C1(n2203), .C2(n2192), .A(n2319), .B(n2200), .ZN(n2299)
         );
  INV_X1 U2108 ( .A(n2151), .ZN(n2200) );
  OAI33_X1 U2109 ( .A1(n2268), .A2(n1631), .A3(n2320), .B1(n1548), .B2(sign), 
        .B3(n2321), .ZN(n2151) );
  AOI22_X1 U2110 ( .A1(n2322), .A2(n1887), .B1(n2323), .B2(n1632), .ZN(n2321)
         );
  OAI21_X1 U2111 ( .B1(n2324), .B2(n2320), .A(n2325), .ZN(n2323) );
  OR3_X1 U2112 ( .A1(n2176), .A2(n2155), .A3(n2326), .ZN(n2325) );
  AOI21_X1 U2113 ( .B1(n2327), .B2(n2176), .A(n2025), .ZN(n2324) );
  OAI21_X1 U2114 ( .B1(n1632), .B2(n2176), .A(n2328), .ZN(n2322) );
  OAI21_X1 U2115 ( .B1(n1889), .B2(n2164), .A(n2150), .ZN(n2328) );
  NAND3_X1 U2116 ( .A1(n2150), .A2(n1632), .A3(n2256), .ZN(n2319) );
  OAI221_X1 U2117 ( .B1(n2320), .B2(n2329), .C1(n2330), .C2(n1575), .A(n2331), 
        .ZN(n2149) );
  NAND3_X1 U2118 ( .A1(n1887), .A2(n2268), .A3(n2150), .ZN(n2331) );
  NOR2_X1 U2119 ( .A1(n1788), .A2(n1789), .ZN(n2150) );
  AOI21_X1 U2120 ( .B1(n2195), .B2(n2332), .A(n2333), .ZN(n2330) );
  OAI33_X1 U2121 ( .A1(n2334), .A2(n1631), .A3(n2335), .B1(n2336), .B2(n2176), 
        .B3(n2326), .ZN(n2333) );
  OAI21_X1 U2122 ( .B1(n2337), .B2(n2338), .A(n2339), .ZN(n2326) );
  AOI21_X1 U2123 ( .B1(u4_fi_ldz_2a_1_), .B2(u4_fi_ldz_2a_0_), .A(
        u4_fi_ldz_2a_2_), .ZN(n2337) );
  NAND3_X1 U2124 ( .A1(n1887), .A2(n2268), .A3(n1789), .ZN(n2336) );
  AOI211_X1 U2125 ( .C1(n2340), .C2(fract_denorm[21]), .A(n2341), .B(n2342), 
        .ZN(n2335) );
  NOR4_X1 U2126 ( .A1(n1777), .A2(n2343), .A3(n2344), .A4(n2279), .ZN(n2342)
         );
  OAI211_X1 U2127 ( .C1(u4_N796), .C2(n2345), .A(n2346), .B(n2347), .ZN(n2279)
         );
  AOI222_X1 U2128 ( .A1(u4_exp_out_mi1[4]), .A2(n2291), .B1(u4_exp_fix_diva[4]), .B2(n2288), .C1(u4_exp_fix_divb[4]), .C2(n2289), .ZN(n2347) );
  NOR3_X1 U2129 ( .A1(n2318), .A2(n2329), .A3(n2161), .ZN(n2289) );
  AND3_X1 U2130 ( .A1(n2332), .A2(n2161), .A3(n2348), .ZN(n2288) );
  NAND2_X1 U2131 ( .A1(n2349), .A2(n2350), .ZN(n2161) );
  OAI21_X1 U2132 ( .B1(u4_N203), .B2(u4_N264), .A(u4_N152), .ZN(n2350) );
  INV_X1 U2133 ( .A(n2351), .ZN(u4_N264) );
  OAI21_X1 U2134 ( .B1(n2352), .B2(n2353), .A(n1902), .ZN(n2351) );
  NOR3_X1 U2135 ( .A1(n2354), .A2(fract_denorm[18]), .A3(fract_denorm[17]), 
        .ZN(n2352) );
  AOI211_X1 U2136 ( .C1(n2355), .C2(n2356), .A(fract_denorm[16]), .B(
        fract_denorm[15]), .ZN(n2354) );
  OAI21_X1 U2137 ( .B1(n2357), .B2(n2358), .A(n2359), .ZN(n2356) );
  AOI211_X1 U2138 ( .C1(n2360), .C2(n2361), .A(n2704), .B(fract_denorm[8]), 
        .ZN(n2357) );
  OAI211_X1 U2139 ( .C1(n2705), .C2(n2706), .A(n2024), .B(n2023), .ZN(n2361)
         );
  INV_X1 U2140 ( .A(n2362), .ZN(u4_N203) );
  OAI211_X1 U2141 ( .C1(n2363), .C2(n2364), .A(n1902), .B(n2365), .ZN(n2362)
         );
  AOI211_X1 U2142 ( .C1(n2366), .C2(n2367), .A(n2368), .B(n2369), .ZN(n2363)
         );
  NAND3_X1 U2143 ( .A1(n2024), .A2(n2023), .A3(n2360), .ZN(n2367) );
  AOI22_X1 U2144 ( .A1(u4_exp_out_pl1_4_), .A2(n2285), .B1(n2286), .B2(
        u4_exp_next_mi_4_), .ZN(n2346) );
  INV_X1 U2145 ( .A(n2308), .ZN(n2286) );
  NAND3_X1 U2146 ( .A1(n2133), .A2(n1531), .A3(n2348), .ZN(n2308) );
  OAI22_X1 U2147 ( .A1(n2143), .A2(n2370), .B1(n2312), .B2(n2268), .ZN(n2285)
         );
  INV_X1 U2148 ( .A(n2256), .ZN(n2268) );
  INV_X1 U2149 ( .A(n2287), .ZN(n2345) );
  OAI21_X1 U2150 ( .B1(n2310), .B2(n1548), .A(n2306), .ZN(n2287) );
  AOI21_X1 U2151 ( .B1(n2312), .B2(n2256), .A(n2371), .ZN(n2306) );
  NOR3_X1 U2152 ( .A1(n2262), .A2(n2348), .A3(n2264), .ZN(n2371) );
  INV_X1 U2153 ( .A(n2318), .ZN(n2348) );
  NAND4_X1 U2154 ( .A1(n2372), .A2(n2373), .A3(n2374), .A4(u4_fract_out_0_), 
        .ZN(n2318) );
  INV_X1 U2155 ( .A(n2176), .ZN(n2373) );
  AND2_X1 U2156 ( .A1(n2195), .A2(n2203), .ZN(n2262) );
  NAND2_X1 U2157 ( .A1(n2272), .A2(u4_fract_out_pl1_10_), .ZN(n2312) );
  INV_X1 U2158 ( .A(n2267), .ZN(n2272) );
  OAI21_X1 U2159 ( .B1(u4_fract_out_0_), .B2(n2374), .A(n2372), .ZN(n2267) );
  INV_X1 U2160 ( .A(n2257), .ZN(u4_fract_out_0_) );
  NOR4_X1 U2161 ( .A1(n1864), .A2(n1870), .A3(u4_N581), .A4(n1867), .ZN(n2344)
         );
  INV_X1 U2162 ( .A(u4_exp_out_2_), .ZN(n1867) );
  INV_X1 U2163 ( .A(u4_exp_out_0_), .ZN(u4_N581) );
  INV_X1 U2164 ( .A(u4_exp_out_1_), .ZN(n1870) );
  AOI21_X1 U2165 ( .B1(n2320), .B2(n2375), .A(n1896), .ZN(n2341) );
  OAI21_X1 U2166 ( .B1(n2338), .B2(n2339), .A(n2195), .ZN(n2375) );
  INV_X1 U2167 ( .A(u4_fi_ldz_2a_4_), .ZN(n2339) );
  INV_X1 U2168 ( .A(u4_fi_ldz_2a_3_), .ZN(n2338) );
  OAI21_X1 U2169 ( .B1(n1789), .B2(n2176), .A(n2320), .ZN(n2340) );
  NAND3_X1 U2170 ( .A1(n2164), .A2(n1894), .A3(n2376), .ZN(n2176) );
  NAND2_X1 U2171 ( .A1(sign), .A2(rmode_r3[1]), .ZN(n2334) );
  AND4_X1 U2172 ( .A1(u4_exp_out_2_), .A2(u4_exp_out_0_), .A3(n2377), .A4(
        u4_exp_out_1_), .ZN(n2195) );
  OAI211_X1 U2173 ( .C1(n2378), .C2(n2032), .A(n2379), .B(n2380), .ZN(
        u4_exp_out_1_) );
  AOI221_X1 U2174 ( .B1(u4_N444), .B2(n2029), .C1(u4_exp_f2i_1[24]), .C2(n2028), .A(n2381), .ZN(n2380) );
  INV_X1 U2175 ( .A(n845), .ZN(n2381) );
  AOI21_X1 U2176 ( .B1(n2382), .B2(fract_denorm[21]), .A(n2035), .ZN(n2379) );
  INV_X1 U2177 ( .A(n2383), .ZN(n2382) );
  AOI222_X1 U2178 ( .A1(u4_div_exp1_1_), .A2(opb_dn), .B1(u4_div_exp2[1]), 
        .B2(n2034), .C1(u4_exp_out1_mi1[1]), .C2(n2033), .ZN(n2378) );
  NOR2_X1 U2179 ( .A1(u4_N796), .A2(n1864), .ZN(n2377) );
  INV_X1 U2180 ( .A(u4_exp_out_3_), .ZN(n1864) );
  NAND2_X1 U2181 ( .A1(n2384), .A2(n2385), .ZN(u4_exp_out_3_) );
  AOI211_X1 U2182 ( .C1(u4_N446), .C2(n2029), .A(n2035), .B(n2386), .ZN(n2385)
         );
  NOR2_X1 U2183 ( .A1(n2387), .A2(n2032), .ZN(n2386) );
  AOI222_X1 U2184 ( .A1(u4_div_exp1_3_), .A2(opb_dn), .B1(u4_div_exp2[3]), 
        .B2(n2034), .C1(u4_exp_out1_mi1[3]), .C2(n2033), .ZN(n2387) );
  AOI222_X1 U2185 ( .A1(u4_div_exp3[3]), .A2(n842), .B1(u4_exp_f2i_1[26]), 
        .B2(n2028), .C1(u4_sub_465_A_3_), .C2(n848), .ZN(n2384) );
  MUX2_X1 U2186 ( .A(u4_exp_in_pl1_3_), .B(u4_exp_next_mi_3_), .S(n1902), .Z(
        u4_sub_465_A_3_) );
  INV_X1 U2187 ( .A(u4_exp_out_4_), .ZN(u4_N796) );
  OAI211_X1 U2188 ( .C1(n831), .C2(n2388), .A(n2389), .B(n2390), .ZN(
        u4_exp_out_4_) );
  AOI221_X1 U2189 ( .B1(u4_N447), .B2(n2029), .C1(n2171), .C2(n1632), .A(n2035), .ZN(n2390) );
  NOR4_X1 U2190 ( .A1(n1573), .A2(n2144), .A3(n2391), .A4(n1877), .ZN(n2035)
         );
  INV_X1 U2191 ( .A(n2175), .ZN(n2171) );
  MUX2_X1 U2192 ( .A(n2392), .B(n2393), .S(n2394), .Z(n2175) );
  AOI222_X1 U2193 ( .A1(u4_div_exp1_4_), .A2(opb_dn), .B1(u4_div_exp2[4]), 
        .B2(n2034), .C1(u4_exp_out1_mi1[4]), .C2(n2033), .ZN(n2393) );
  INV_X1 U2194 ( .A(u4_div_exp3[4]), .ZN(n2392) );
  NAND2_X1 U2195 ( .A1(u4_exp_f2i_1[27]), .A2(n2028), .ZN(n2389) );
  INV_X1 U2196 ( .A(u4_sub_465_A_4_), .ZN(n2388) );
  MUX2_X1 U2197 ( .A(u4_exp_in_pl1_4_), .B(u4_exp_next_mi_4_), .S(n1902), .Z(
        u4_sub_465_A_4_) );
  AOI21_X1 U2198 ( .B1(u4_fi_ldz_2a_0_), .B2(n2029), .A(n2397), .ZN(n2396) );
  OAI22_X1 U2199 ( .A1(n2398), .A2(n2032), .B1(n2399), .B2(n2383), .ZN(n2397)
         );
  NAND2_X1 U2200 ( .A1(n2400), .A2(n2391), .ZN(n2383) );
  INV_X1 U2201 ( .A(fract_denorm[20]), .ZN(n2399) );
  NAND2_X1 U2202 ( .A1(n2394), .A2(n1632), .ZN(n2032) );
  AOI222_X1 U2203 ( .A1(u4_div_exp1_0_), .A2(opb_dn), .B1(u4_div_exp2[0]), 
        .B2(n2034), .C1(u4_exp_out1_mi1[0]), .C2(n2033), .ZN(n2398) );
  NOR2_X1 U2204 ( .A1(n2096), .A2(n2025), .ZN(n2033) );
  INV_X1 U2205 ( .A(n2401), .ZN(n2025) );
  INV_X1 U2206 ( .A(n2402), .ZN(n2034) );
  OAI21_X1 U2207 ( .B1(n2403), .B2(n2404), .A(opa_dn), .ZN(n2402) );
  OAI221_X1 U2208 ( .B1(n2475), .B2(n2163), .C1(n1830), .C2(exp_r[2]), .A(
        n2407), .ZN(n2406) );
  OAI221_X1 U2209 ( .B1(n1784), .B2(n2408), .C1(n1782), .C2(div_opa_ldz_r2[2]), 
        .A(n2409), .ZN(n2407) );
  OAI21_X1 U2210 ( .B1(n1891), .B2(n2410), .A(n1829), .ZN(n2409) );
  INV_X1 U2211 ( .A(n2410), .ZN(n2408) );
  NAND2_X1 U2212 ( .A1(n1786), .A2(div_opa_ldz_r2[0]), .ZN(n2410) );
  NAND2_X1 U2213 ( .A1(n2475), .A2(n2163), .ZN(n2405) );
  NOR3_X1 U2214 ( .A1(n2391), .A2(n1877), .A3(n2190), .ZN(n2029) );
  AOI222_X1 U2215 ( .A1(u4_div_exp3[0]), .A2(n842), .B1(u4_exp_f2i_1[23]), 
        .B2(n2028), .C1(u4_sub_465_A_0_), .C2(n848), .ZN(n2395) );
  INV_X1 U2216 ( .A(n831), .ZN(n848) );
  NAND4_X1 U2217 ( .A1(n2187), .A2(n1631), .A3(n2411), .A4(n2412), .ZN(n831)
         );
  AOI21_X1 U2218 ( .B1(n2183), .B2(n2124), .A(n1888), .ZN(n2412) );
  NAND3_X1 U2219 ( .A1(n2143), .A2(n2370), .A3(n1789), .ZN(n2411) );
  INV_X1 U2220 ( .A(n2311), .ZN(n2143) );
  MUX2_X1 U2221 ( .A(u4_exp_in_pl1_0_), .B(u4_exp_next_mi_0_), .S(n1902), .Z(
        u4_sub_465_A_0_) );
  AND3_X1 U2222 ( .A1(n2191), .A2(n2192), .A3(n1877), .ZN(n2028) );
  NAND2_X1 U2223 ( .A1(n2204), .A2(n2413), .ZN(n2192) );
  INV_X1 U2224 ( .A(n2414), .ZN(n2413) );
  NOR2_X1 U2225 ( .A1(n2394), .A2(n1631), .ZN(n842) );
  NAND2_X1 U2226 ( .A1(opa_dn), .A2(opb_dn), .ZN(n2394) );
  INV_X1 U2227 ( .A(n2332), .ZN(n2329) );
  NOR2_X1 U2228 ( .A1(n2264), .A2(n1531), .ZN(n2332) );
  INV_X1 U2229 ( .A(n2133), .ZN(n2264) );
  NOR2_X1 U2230 ( .A1(n1576), .A2(rmode_r3[1]), .ZN(n2133) );
  NAND3_X1 U2231 ( .A1(opb_dn), .A2(n1574), .A3(u4_N487), .ZN(n2320) );
  NOR2_X1 U2232 ( .A1(n2370), .A2(n2311), .ZN(n2291) );
  NAND2_X1 U2233 ( .A1(n2310), .A2(rmode_r3[1]), .ZN(n2370) );
  AND2_X1 U2234 ( .A1(u4_fract_out_pl1_10_), .A2(n2270), .ZN(n2310) );
  OAI21_X1 U2235 ( .B1(sign), .B2(n2415), .A(n2416), .ZN(n2270) );
  OAI211_X1 U2236 ( .C1(n2417), .C2(n2177), .A(n1576), .B(n1877), .ZN(n2416)
         );
  NAND2_X1 U2237 ( .A1(n2418), .A2(n2419), .ZN(n2177) );
  AOI211_X1 U2238 ( .C1(n2420), .C2(n2366), .A(n2164), .B(opas_r2), .ZN(n2417)
         );
  MUX2_X1 U2239 ( .A(n2421), .B(n2422), .S(n2423), .Z(n2415) );
  NAND3_X1 U2240 ( .A1(n2186), .A2(n2203), .A3(u4_N798), .ZN(n2422) );
  INV_X1 U2241 ( .A(n2424), .ZN(n2186) );
  AOI22_X1 U2242 ( .A1(n2425), .A2(n2426), .B1(n2427), .B2(n2428), .ZN(n2421)
         );
  NAND4_X1 U2243 ( .A1(n2429), .A2(n2430), .A3(n2431), .A4(n1631), .ZN(n2428)
         );
  NAND3_X1 U2244 ( .A1(n2343), .A2(n2164), .A3(n1788), .ZN(n2431) );
  NAND2_X1 U2245 ( .A1(n2183), .A2(n1789), .ZN(n2430) );
  INV_X1 U2246 ( .A(n2327), .ZN(n2429) );
  NOR2_X1 U2247 ( .A1(n1546), .A2(n1575), .ZN(n2327) );
  INV_X1 U2248 ( .A(n2432), .ZN(n2426) );
  AOI211_X1 U2249 ( .C1(n1631), .C2(n2155), .A(n2145), .B(n2427), .ZN(n2432)
         );
  OAI21_X1 U2250 ( .B1(n1531), .B2(n2157), .A(n2424), .ZN(n2427) );
  NOR2_X1 U2251 ( .A1(n2374), .A2(n2372), .ZN(n2424) );
  AOI21_X1 U2252 ( .B1(n2433), .B2(n2434), .A(n2418), .ZN(n2372) );
  AND3_X1 U2253 ( .A1(n2435), .A2(n2355), .A3(u4_N326), .ZN(n2434) );
  NOR4_X1 U2254 ( .A1(n2369), .A2(n2027), .A3(fract_denorm[10]), .A4(n1631), 
        .ZN(n2433) );
  INV_X1 U2255 ( .A(n2359), .ZN(n2369) );
  OAI21_X1 U2256 ( .B1(n1531), .B2(n2418), .A(n2419), .ZN(n2374) );
  AOI22_X1 U2257 ( .A1(n2436), .A2(n2437), .B1(n2438), .B2(n2439), .ZN(n2419)
         );
  NAND4_X1 U2258 ( .A1(n2440), .A2(n2441), .A3(n2442), .A4(n2443), .ZN(n2438)
         );
  NOR3_X1 U2259 ( .A1(u4_N396), .A2(u4_N398), .A3(u4_N397), .ZN(n2443) );
  NOR3_X1 U2260 ( .A1(u4_N393), .A2(u4_N395), .A3(u4_N394), .ZN(n2442) );
  NOR3_X1 U2261 ( .A1(u4_N390), .A2(u4_N392), .A3(u4_N391), .ZN(n2441) );
  NOR2_X1 U2262 ( .A1(u4_N389), .A2(u4_N388), .ZN(n2440) );
  NAND4_X1 U2263 ( .A1(n2444), .A2(n2445), .A3(n2446), .A4(n2447), .ZN(n2436)
         );
  NOR3_X1 U2264 ( .A1(u4_N420), .A2(u4_N422), .A3(u4_N421), .ZN(n2447) );
  NOR3_X1 U2265 ( .A1(u4_N417), .A2(u4_N419), .A3(u4_N418), .ZN(n2446) );
  NOR3_X1 U2266 ( .A1(u4_N414), .A2(u4_N416), .A3(u4_N415), .ZN(n2445) );
  NOR2_X1 U2267 ( .A1(u4_N413), .A2(u4_N412), .ZN(n2444) );
  AOI22_X1 U2268 ( .A1(u4_N399), .A2(n2439), .B1(u4_N423), .B2(n2437), .ZN(
        n2418) );
  AND4_X1 U2269 ( .A1(n2448), .A2(n2449), .A3(n2450), .A4(n2451), .ZN(n2157)
         );
  NOR4_X1 U2270 ( .A1(n2452), .A2(remainder[4]), .A3(remainder[6]), .A4(
        remainder[5]), .ZN(n2451) );
  NAND3_X1 U2271 ( .A1(n1772), .A2(n1771), .A3(n1773), .ZN(n2452) );
  NOR4_X1 U2272 ( .A1(n2453), .A2(remainder[20]), .A3(remainder[22]), .A4(
        remainder[21]), .ZN(n2450) );
  NAND3_X1 U2273 ( .A1(n1775), .A2(n1774), .A3(n1766), .ZN(n2453) );
  NOR4_X1 U2274 ( .A1(n2454), .A2(remainder[15]), .A3(remainder[17]), .A4(
        remainder[16]), .ZN(n2449) );
  NAND3_X1 U2275 ( .A1(n1767), .A2(n1776), .A3(n1768), .ZN(n2454) );
  AND4_X1 U2276 ( .A1(n2257), .A2(n1900), .A3(n2456), .A4(n2457), .ZN(n2145)
         );
  NOR3_X1 U2277 ( .A1(n2458), .A2(u4_fract_out_6_), .A3(u4_fract_out_5_), .ZN(
        n2457) );
  INV_X1 U2278 ( .A(n2241), .ZN(u4_fract_out_5_) );
  AOI22_X1 U2279 ( .A1(u4_N429), .A2(n2437), .B1(u4_N405), .B2(n2439), .ZN(
        n2241) );
  INV_X1 U2280 ( .A(n2239), .ZN(u4_fract_out_6_) );
  AOI22_X1 U2281 ( .A1(u4_N430), .A2(n2437), .B1(u4_N406), .B2(n2439), .ZN(
        n2239) );
  NAND3_X1 U2282 ( .A1(n1898), .A2(n1897), .A3(n1899), .ZN(n2458) );
  AOI22_X1 U2283 ( .A1(u4_N431), .A2(n2437), .B1(u4_N407), .B2(n2439), .ZN(
        n1899) );
  AOI22_X1 U2284 ( .A1(u4_N433), .A2(n2437), .B1(u4_N409), .B2(n2439), .ZN(
        n1897) );
  AOI22_X1 U2285 ( .A1(u4_N432), .A2(n2437), .B1(u4_N408), .B2(n2439), .ZN(
        n1898) );
  NOR3_X1 U2286 ( .A1(u4_fract_out_2_), .A2(u4_fract_out_4_), .A3(
        u4_fract_out_3_), .ZN(n2456) );
  INV_X1 U2287 ( .A(n2245), .ZN(u4_fract_out_3_) );
  AOI22_X1 U2288 ( .A1(u4_N427), .A2(n2437), .B1(u4_N403), .B2(n2439), .ZN(
        n2245) );
  INV_X1 U2289 ( .A(n2243), .ZN(u4_fract_out_4_) );
  AOI22_X1 U2290 ( .A1(u4_N428), .A2(n2437), .B1(u4_N404), .B2(n2439), .ZN(
        n2243) );
  INV_X1 U2291 ( .A(n2247), .ZN(u4_fract_out_2_) );
  AOI22_X1 U2292 ( .A1(u4_N426), .A2(n2437), .B1(u4_N402), .B2(n2439), .ZN(
        n2247) );
  AOI22_X1 U2293 ( .A1(u4_N425), .A2(n2437), .B1(u4_N401), .B2(n2439), .ZN(
        n1900) );
  NOR2_X1 U2294 ( .A1(n1788), .A2(n2190), .ZN(n2425) );
  INV_X1 U2295 ( .A(n2144), .ZN(n2190) );
  AND2_X1 U2296 ( .A1(n2260), .A2(n2459), .ZN(n2274) );
  NAND3_X1 U2297 ( .A1(n1632), .A2(n1575), .A3(n1789), .ZN(n2459) );
  AOI221_X1 U2298 ( .B1(n2124), .B2(opb_00), .C1(n1887), .C2(opa_00), .A(n2061), .ZN(n2260) );
  NOR2_X1 U2299 ( .A1(n1549), .A2(n1531), .ZN(n2061) );
  AOI22_X1 U2300 ( .A1(u4_N400), .A2(n2439), .B1(u4_N424), .B2(n2437), .ZN(
        n2257) );
  OAI221_X1 U2301 ( .B1(n1895), .B2(n2463), .C1(n2464), .C2(n2465), .A(n2466), 
        .ZN(n2462) );
  INV_X1 U2302 ( .A(n1878), .ZN(n2465) );
  OAI221_X1 U2303 ( .B1(n1631), .B2(n2467), .C1(n1885), .C2(n2468), .A(n2469), 
        .ZN(n1878) );
  MUX2_X1 U2304 ( .A(n2470), .B(n1877), .S(n1888), .Z(n2469) );
  INV_X1 U2305 ( .A(n2391), .ZN(n1888) );
  NAND2_X1 U2306 ( .A1(n2471), .A2(n2423), .ZN(n2470) );
  AOI21_X1 U2307 ( .B1(n2472), .B2(n2027), .A(u4_N656), .ZN(n2467) );
  OAI21_X1 U2308 ( .B1(n1789), .B2(n2155), .A(n2170), .ZN(n2472) );
  NAND2_X1 U2309 ( .A1(n2155), .A2(n1575), .ZN(n2170) );
  NOR2_X1 U2310 ( .A1(u4_N95), .A2(u4_N152), .ZN(n2464) );
  MUX2_X1 U2311 ( .A(n2474), .B(n2475), .S(n1889), .Z(n2463) );
  NOR2_X1 U2312 ( .A1(u4_div_scht1a[4]), .A2(u4_div_scht1a[3]), .ZN(n2474) );
  NAND3_X1 U2313 ( .A1(n1632), .A2(n2182), .A3(n2476), .ZN(n1895) );
  OAI21_X1 U2314 ( .B1(n2155), .B2(n1546), .A(n2027), .ZN(n2476) );
  OAI21_X1 U2315 ( .B1(n2477), .B2(n2203), .A(n2478), .ZN(n2461) );
  OAI21_X1 U2316 ( .B1(n2163), .B2(n2164), .A(n1874), .ZN(n2478) );
  NOR4_X1 U2317 ( .A1(n2096), .A2(n1575), .A3(n1631), .A4(u4_N656), .ZN(n1874)
         );
  INV_X1 U2318 ( .A(n1777), .ZN(n2164) );
  INV_X1 U2319 ( .A(n1877), .ZN(n2203) );
  NOR3_X1 U2320 ( .A1(n2479), .A2(u4_f2i_shft_4_), .A3(u4_f2i_shft_3_), .ZN(
        n2477) );
  INV_X1 U2321 ( .A(n2191), .ZN(n2479) );
  NAND2_X1 U2322 ( .A1(n2204), .A2(n2414), .ZN(n2191) );
  NAND4_X1 U2323 ( .A1(rmode_r3[1]), .A2(rmode_r3[0]), .A3(opas_r2), .A4(n2144), .ZN(n2414) );
  NAND2_X1 U2324 ( .A1(u4_N95), .A2(n2420), .ZN(n2144) );
  AND4_X1 U2325 ( .A1(n2024), .A2(n2023), .A3(n2360), .A4(n2480), .ZN(n2420)
         );
  NOR3_X1 U2326 ( .A1(n2707), .A2(n2705), .A3(n2706), .ZN(n2480) );
  INV_X1 U2327 ( .A(n1919), .ZN(n2706) );
  AOI222_X1 U2328 ( .A1(n2481), .A2(quo[4]), .B1(n1560), .B2(n1539), .C1(n2482), .C2(prod[2]), .ZN(n1919) );
  OAI222_X1 U2329 ( .A1(n2483), .A2(n1558), .B1(n1628), .B2(n1793), .C1(n2484), 
        .C2(n1537), .ZN(n2705) );
  OAI222_X1 U2330 ( .A1(n2483), .A2(n1572), .B1(n1628), .B2(n1792), .C1(n2484), 
        .C2(n1544), .ZN(n2707) );
  NOR2_X1 U2331 ( .A1(n2709), .A2(n2708), .ZN(n2360) );
  INV_X1 U2332 ( .A(n1916), .ZN(n2708) );
  AOI222_X1 U2333 ( .A1(n2481), .A2(quo[8]), .B1(n1560), .B2(n1540), .C1(n2482), .C2(prod[6]), .ZN(n1916) );
  INV_X1 U2334 ( .A(n1918), .ZN(n2709) );
  AOI222_X1 U2335 ( .A1(n2481), .A2(quo[7]), .B1(n1560), .B2(n1541), .C1(n2482), .C2(prod[5]), .ZN(n1918) );
  AOI222_X1 U2336 ( .A1(n2481), .A2(quo[6]), .B1(n1560), .B2(n1542), .C1(n2482), .C2(prod[4]), .ZN(n2023) );
  AOI222_X1 U2337 ( .A1(n2481), .A2(quo[5]), .B1(n1560), .B2(n1543), .C1(n2482), .C2(prod[3]), .ZN(n2024) );
  INV_X1 U2338 ( .A(n2349), .ZN(u4_N95) );
  NAND3_X1 U2339 ( .A1(n2485), .A2(n1902), .A3(n2435), .ZN(n2349) );
  NOR2_X1 U2340 ( .A1(n2364), .A2(n2353), .ZN(n2435) );
  INV_X1 U2341 ( .A(n2365), .ZN(n2353) );
  NOR2_X1 U2342 ( .A1(fract_denorm[19]), .A2(fract_denorm[20]), .ZN(n2365) );
  OAI221_X1 U2343 ( .B1(n2484), .B2(n1561), .C1(n1628), .C2(n1806), .A(n2486), 
        .ZN(fract_denorm[20]) );
  OAI221_X1 U2344 ( .B1(n2484), .B2(n1545), .C1(n1628), .C2(n1805), .A(n2488), 
        .ZN(fract_denorm[19]) );
  OR4_X1 U2345 ( .A1(fract_denorm[15]), .A2(fract_denorm[16]), .A3(
        fract_denorm[17]), .A4(fract_denorm[18]), .ZN(n2364) );
  OAI221_X1 U2346 ( .B1(n2484), .B2(n1534), .C1(n1628), .C2(n1804), .A(n2489), 
        .ZN(fract_denorm[18]) );
  AOI222_X1 U2347 ( .A1(quo[10]), .A2(n2487), .B1(n2065), .B2(fract_out_q[11]), 
        .C1(quo[20]), .C2(n2481), .ZN(n2489) );
  OAI221_X1 U2348 ( .B1(n2484), .B2(n1563), .C1(n1833), .C2(n1803), .A(n2490), 
        .ZN(fract_denorm[17]) );
  AOI222_X1 U2349 ( .A1(quo[9]), .A2(n2487), .B1(n2065), .B2(fract_out_q[10]), 
        .C1(quo[19]), .C2(n2481), .ZN(n2490) );
  OAI221_X1 U2350 ( .B1(n2484), .B2(n1566), .C1(n1833), .C2(n1802), .A(n2491), 
        .ZN(fract_denorm[16]) );
  AOI222_X1 U2351 ( .A1(quo[8]), .A2(n2487), .B1(n2065), .B2(fract_out_q[9]), 
        .C1(quo[18]), .C2(n2481), .ZN(n2491) );
  OAI221_X1 U2352 ( .B1(n2484), .B2(n1567), .C1(n1628), .C2(n1801), .A(n2492), 
        .ZN(fract_denorm[15]) );
  AOI222_X1 U2353 ( .A1(quo[7]), .A2(n2487), .B1(n2065), .B2(fract_out_q[8]), 
        .C1(quo[17]), .C2(n2481), .ZN(n2492) );
  INV_X1 U2354 ( .A(n2473), .ZN(n2485) );
  NAND3_X1 U2355 ( .A1(n2366), .A2(n2359), .A3(n2355), .ZN(n2473) );
  INV_X1 U2356 ( .A(n2368), .ZN(n2355) );
  NAND2_X1 U2357 ( .A1(n1910), .A2(n1908), .ZN(n2368) );
  INV_X1 U2358 ( .A(fract_denorm[14]), .ZN(n1908) );
  OAI221_X1 U2359 ( .B1(n2484), .B2(n1565), .C1(n1628), .C2(n1800), .A(n2493), 
        .ZN(fract_denorm[14]) );
  AOI222_X1 U2360 ( .A1(quo[6]), .A2(n2487), .B1(n2065), .B2(fract_out_q[7]), 
        .C1(quo[16]), .C2(n2481), .ZN(n2493) );
  INV_X1 U2361 ( .A(fract_denorm[13]), .ZN(n1910) );
  OAI221_X1 U2362 ( .B1(n2484), .B2(n1569), .C1(n1628), .C2(n1799), .A(n2494), 
        .ZN(fract_denorm[13]) );
  AOI222_X1 U2363 ( .A1(quo[5]), .A2(n2487), .B1(n2065), .B2(fract_out_q[6]), 
        .C1(quo[15]), .C2(n2481), .ZN(n2494) );
  NOR2_X1 U2364 ( .A1(fract_denorm[11]), .A2(fract_denorm[12]), .ZN(n2359) );
  OAI221_X1 U2365 ( .B1(n2484), .B2(n1571), .C1(n1628), .C2(n1798), .A(n2495), 
        .ZN(fract_denorm[12]) );
  AOI222_X1 U2366 ( .A1(quo[4]), .A2(n2487), .B1(n2065), .B2(fract_out_q[5]), 
        .C1(quo[14]), .C2(n2481), .ZN(n2495) );
  OAI221_X1 U2367 ( .B1(n2484), .B2(n1568), .C1(n1628), .C2(n1797), .A(n2496), 
        .ZN(fract_denorm[11]) );
  AOI222_X1 U2368 ( .A1(quo[3]), .A2(n2487), .B1(n2065), .B2(fract_out_q[4]), 
        .C1(quo[13]), .C2(n2481), .ZN(n2496) );
  NOR3_X1 U2369 ( .A1(fract_denorm[8]), .A2(n2704), .A3(n2358), .ZN(n2366) );
  NAND2_X1 U2370 ( .A1(n1912), .A2(n1914), .ZN(n2358) );
  INV_X1 U2371 ( .A(fract_denorm[9]), .ZN(n1914) );
  OAI221_X1 U2372 ( .B1(n2484), .B2(n1570), .C1(n1628), .C2(n1795), .A(n2497), 
        .ZN(fract_denorm[9]) );
  INV_X1 U2373 ( .A(fract_denorm[10]), .ZN(n1912) );
  OAI221_X1 U2374 ( .B1(n2484), .B2(n1562), .C1(n1833), .C2(n1796), .A(n2498), 
        .ZN(fract_denorm[10]) );
  OAI221_X1 U2375 ( .B1(n1813), .B2(n2125), .C1(n2483), .C2(n1556), .A(n2499), 
        .ZN(n2704) );
  AOI22_X1 U2376 ( .A1(prod[7]), .A2(n2482), .B1(n1560), .B2(fract_i2f_7_), 
        .ZN(n2499) );
  OAI221_X1 U2377 ( .B1(n2484), .B2(n1557), .C1(n1628), .C2(n1794), .A(n2500), 
        .ZN(fract_denorm[8]) );
  AOI222_X1 U2378 ( .A1(quo[0]), .A2(n2487), .B1(n2065), .B2(fract_out_q[1]), 
        .C1(quo[10]), .C2(n2481), .ZN(n2500) );
  NAND2_X1 U2379 ( .A1(opb_dn), .A2(n2501), .ZN(n2483) );
  AND2_X1 U2380 ( .A1(n1777), .A2(n2502), .ZN(n2204) );
  OAI21_X1 U2381 ( .B1(n2256), .B2(n1894), .A(n2376), .ZN(n2502) );
  NOR3_X1 U2382 ( .A1(n1782), .A2(n1784), .A3(n1780), .ZN(n2376) );
  NOR2_X1 U2383 ( .A1(rmode_r3[0]), .A2(rmode_r3[1]), .ZN(n2256) );
  INV_X1 U2384 ( .A(n2503), .ZN(n2460) );
  OAI21_X1 U2385 ( .B1(u4_exp_in_pl1_3_), .B2(u4_exp_in_pl1_4_), .A(n1879), 
        .ZN(n2503) );
  OAI21_X1 U2386 ( .B1(n1884), .B2(n1885), .A(n2504), .ZN(n1879) );
  NAND4_X1 U2387 ( .A1(n2391), .A2(n2423), .A3(n1890), .A4(n1896), .ZN(n2504)
         );
  INV_X1 U2388 ( .A(n2471), .ZN(n1890) );
  NOR2_X1 U2389 ( .A1(n2182), .A2(n2400), .ZN(n2471) );
  INV_X1 U2390 ( .A(n2187), .ZN(n2400) );
  NAND2_X1 U2391 ( .A1(n2423), .A2(n2505), .ZN(n2187) );
  OAI21_X1 U2392 ( .B1(fract_denorm[21]), .B2(n2506), .A(n1896), .ZN(n2505) );
  INV_X1 U2393 ( .A(u4_exp_next_mi_5_), .ZN(n2506) );
  INV_X1 U2394 ( .A(n1887), .ZN(n2423) );
  NAND2_X1 U2395 ( .A1(n1631), .A2(n1885), .ZN(n1887) );
  NOR2_X1 U2396 ( .A1(n1877), .A2(n2189), .ZN(n2391) );
  NOR2_X1 U2397 ( .A1(n1536), .A2(n2507), .ZN(n2189) );
  INV_X1 U2398 ( .A(n2124), .ZN(n1885) );
  INV_X1 U2399 ( .A(n2468), .ZN(n1884) );
  OAI211_X1 U2400 ( .C1(n2508), .C2(n1575), .A(n2401), .B(n2179), .ZN(n2468)
         );
  INV_X1 U2401 ( .A(u4_exp_in_mi1_5_), .ZN(n2179) );
  NAND2_X1 U2402 ( .A1(n1788), .A2(n1889), .ZN(n2401) );
  INV_X1 U2403 ( .A(n1896), .ZN(n1889) );
  NOR2_X1 U2404 ( .A1(n2183), .A2(n2182), .ZN(n2508) );
  INV_X1 U2405 ( .A(u4_N656), .ZN(n2182) );
  MUX2_X1 U2406 ( .A(u4_exp_in_pl1_5_), .B(u4_exp_next_mi_5_), .S(n1902), .Z(
        n2183) );
  AOI22_X1 U2407 ( .A1(n2065), .A2(fract_out_q[14]), .B1(prod[21]), .B2(n2124), 
        .ZN(n2510) );
  NAND2_X1 U2408 ( .A1(n1832), .A2(n1833), .ZN(n2125) );
  NAND2_X1 U2409 ( .A1(n1832), .A2(n1560), .ZN(n2507) );
  MUX2_X1 U2410 ( .A(n1564), .B(n1765), .S(opb_dn), .Z(n2509) );
  NAND2_X1 U2411 ( .A1(n2511), .A2(n2512), .ZN(n2466) );
  OAI21_X1 U2412 ( .B1(u4_exp_in_mi1_5_), .B2(n2311), .A(n1531), .ZN(n2512) );
  NOR2_X1 U2413 ( .A1(n1831), .A2(n1832), .ZN(n2501) );
  NAND2_X1 U2414 ( .A1(n2124), .A2(n1575), .ZN(n2311) );
  NOR2_X1 U2415 ( .A1(n1536), .A2(n1832), .ZN(n2482) );
  OAI21_X1 U2416 ( .B1(n1862), .B2(n1546), .A(n1788), .ZN(n2511) );
  AND2_X1 U2417 ( .A1(n2026), .A2(n2027), .ZN(n1862) );
  NAND2_X1 U2418 ( .A1(n2096), .A2(n1575), .ZN(n2027) );
  NAND3_X1 U2419 ( .A1(n1896), .A2(n2096), .A3(u4_div_scht1a[5]), .ZN(n2026)
         );
  NAND2_X1 U2420 ( .A1(n1574), .A2(n1538), .ZN(n2096) );
  NAND2_X1 U2421 ( .A1(n1777), .A2(n2343), .ZN(n1896) );
  NOR4_X1 U2422 ( .A1(n1894), .A2(n1891), .A3(exp_r[2]), .A4(n2163), .ZN(n2343) );
  INV_X1 U2423 ( .A(n1780), .ZN(n2163) );
  INV_X1 U2424 ( .A(n1784), .ZN(n1891) );
  INV_X1 U2425 ( .A(n1786), .ZN(n1894) );
  XNOR2_X1 U2426 ( .A(n2513), .B(n1983), .ZN(N216) );
  INV_X1 U2427 ( .A(n1980), .ZN(n1983) );
  NAND2_X1 U2428 ( .A1(rmode_r2[1]), .A2(rmode_r2[0]), .ZN(n1980) );
  NAND2_X1 U2429 ( .A1(n2514), .A2(n2515), .ZN(N196) );
  NAND2_X1 U2430 ( .A1(n1552), .A2(n2516), .ZN(n2515) );
  NAND2_X1 U2431 ( .A1(n2514), .A2(n2517), .ZN(N195) );
  NAND2_X1 U2432 ( .A1(N151), .A2(n2516), .ZN(n2517) );
  NAND2_X1 U2433 ( .A1(n2514), .A2(n2518), .ZN(N194) );
  NAND2_X1 U2434 ( .A1(N150), .A2(n2516), .ZN(n2518) );
  OAI221_X1 U2435 ( .B1(n2519), .B2(n1550), .C1(n2520), .C2(n1620), .A(n2514), 
        .ZN(N193) );
  OAI221_X1 U2436 ( .B1(n2519), .B2(n1532), .C1(n1621), .C2(n2520), .A(n2514), 
        .ZN(N192) );
  OAI221_X1 U2437 ( .B1(n2519), .B2(n1535), .C1(n1622), .C2(n2520), .A(n2514), 
        .ZN(N191) );
  OAI221_X1 U2438 ( .B1(n2519), .B2(n1585), .C1(n1618), .C2(n2520), .A(n2514), 
        .ZN(N190) );
  OAI221_X1 U2439 ( .B1(n2519), .B2(n1586), .C1(n1619), .C2(n2520), .A(n2514), 
        .ZN(N189) );
  OAI221_X1 U2440 ( .B1(n2519), .B2(n1601), .C1(n2520), .C2(n1614), .A(n2514), 
        .ZN(N188) );
  OAI221_X1 U2441 ( .B1(n2519), .B2(n1602), .C1(n2520), .C2(n1615), .A(n2514), 
        .ZN(N187) );
  OAI221_X1 U2442 ( .B1(n2519), .B2(n1603), .C1(n2520), .C2(n1616), .A(n2514), 
        .ZN(N186) );
  OAI221_X1 U2443 ( .B1(n1530), .B2(n1990), .C1(n2520), .C2(n1617), .A(n2522), 
        .ZN(N185) );
  AOI22_X1 U2444 ( .A1(N141), .A2(n2516), .B1(N116), .B2(n2521), .ZN(n2522) );
  OAI221_X1 U2445 ( .B1(n1990), .B2(n1614), .C1(n2520), .C2(n1612), .A(n2523), 
        .ZN(N184) );
  AOI22_X1 U2446 ( .A1(N140), .A2(n2516), .B1(N115), .B2(n2521), .ZN(n2523) );
  OAI221_X1 U2447 ( .B1(n1990), .B2(n1615), .C1(n2520), .C2(n1613), .A(n2524), 
        .ZN(N183) );
  AOI22_X1 U2448 ( .A1(N139), .A2(n2516), .B1(N114), .B2(n2521), .ZN(n2524) );
  OAI221_X1 U2449 ( .B1(n1990), .B2(n1616), .C1(n1589), .C2(n2520), .A(n2525), 
        .ZN(N182) );
  AOI22_X1 U2450 ( .A1(N138), .A2(n2516), .B1(N113), .B2(n2521), .ZN(n2525) );
  OAI221_X1 U2451 ( .B1(n1990), .B2(n1617), .C1(n1590), .C2(n2520), .A(n2526), 
        .ZN(N181) );
  AOI22_X1 U2452 ( .A1(n2516), .A2(N106), .B1(N112), .B2(n2521), .ZN(n2526) );
  INV_X1 U2453 ( .A(n2519), .ZN(n2516) );
  OAI21_X1 U2454 ( .B1(n1591), .B2(n2520), .A(n2528), .ZN(N180) );
  AOI22_X1 U2455 ( .A1(N111), .A2(n2521), .B1(opa_r1[5]), .B2(n2529), .ZN(
        n2528) );
  OAI21_X1 U2456 ( .B1(n1599), .B2(n2520), .A(n2530), .ZN(N179) );
  AOI22_X1 U2457 ( .A1(N110), .A2(n2521), .B1(opa_r1[4]), .B2(n2529), .ZN(
        n2530) );
  INV_X1 U2458 ( .A(n1990), .ZN(n2529) );
  INV_X1 U2459 ( .A(n1991), .ZN(n2521) );
  NAND2_X1 U2460 ( .A1(n2531), .A2(n2527), .ZN(n1991) );
  INV_X1 U2461 ( .A(n2527), .ZN(n2513) );
  MUX2_X1 U2462 ( .A(sign_fasu), .B(sign_mul), .S(fpu_op_r2[1]), .Z(n2527) );
  NOR2_X1 U2463 ( .A1(opa_r1[11]), .A2(opa_r1[10]), .ZN(n2532) );
  OAI222_X1 U2464 ( .A1(n1808), .A2(n2038), .B1(n1779), .B2(n2039), .C1(n2040), 
        .C2(n1620), .ZN(N100) );
  INV_X1 U2465 ( .A(n2531), .ZN(n2040) );
  NOR2_X1 U2466 ( .A1(fpu_op_r2[1]), .A2(n2041), .ZN(n2531) );
  OR2_X1 U2467 ( .A1(n1834), .A2(n1836), .ZN(n2041) );
  NAND2_X1 U2468 ( .A1(n1836), .A2(fpu_op_r2[1]), .ZN(n2039) );
  NAND2_X1 U2469 ( .A1(n1836), .A2(n1835), .ZN(n2038) );
  INV_X1 u4_add_393_U1 ( .A(u4_fract_out_0_), .ZN(u4_fract_out_pl1_0_) );
  HA_X1 u4_add_393_U1_1_1 ( .A(u4_fract_out_1_), .B(u4_fract_out_0_), .CO(
        u4_add_393_carry[2]), .S(u4_fract_out_pl1_1_) );
  HA_X1 u4_add_393_U1_1_2 ( .A(u4_fract_out_2_), .B(u4_add_393_carry[2]), .CO(
        u4_add_393_carry[3]), .S(u4_fract_out_pl1_2_) );
  HA_X1 u4_add_393_U1_1_3 ( .A(u4_fract_out_3_), .B(u4_add_393_carry[3]), .CO(
        u4_add_393_carry[4]), .S(u4_fract_out_pl1_3_) );
  HA_X1 u4_add_393_U1_1_4 ( .A(u4_fract_out_4_), .B(u4_add_393_carry[4]), .CO(
        u4_add_393_carry[5]), .S(u4_fract_out_pl1_4_) );
  HA_X1 u4_add_393_U1_1_5 ( .A(u4_fract_out_5_), .B(u4_add_393_carry[5]), .CO(
        u4_add_393_carry[6]), .S(u4_fract_out_pl1_5_) );
  HA_X1 u4_add_393_U1_1_6 ( .A(u4_fract_out_6_), .B(u4_add_393_carry[6]), .CO(
        u4_add_393_carry[7]), .S(u4_fract_out_pl1_6_) );
  HA_X1 u4_add_393_U1_1_7 ( .A(u4_fract_out_7_), .B(u4_add_393_carry[7]), .CO(
        u4_add_393_carry[8]), .S(u4_fract_out_pl1_7_) );
  HA_X1 u4_add_393_U1_1_8 ( .A(u4_fract_out_8_), .B(u4_add_393_carry[8]), .CO(
        u4_add_393_carry[9]), .S(u4_fract_out_pl1_8_) );
  HA_X1 u4_add_393_U1_1_9 ( .A(u4_fract_out_9_), .B(u4_add_393_carry[9]), .CO(
        u4_fract_out_pl1_10_), .S(u4_fract_out_pl1_9_) );
  INV_X1 u4_srl_450_U100 ( .A(u4_shift_right[0]), .ZN(u4_srl_450_n76) );
  AOI22_X1 u4_srl_450_U99 ( .A1(n2705), .A2(u4_srl_450_n6), .B1(n2707), .B2(
        u4_srl_450_n3), .ZN(u4_srl_450_n75) );
  OAI221_X1 u4_srl_450_U98 ( .B1(u4_srl_450_n39), .B2(u4_srl_450_n29), .C1(
        u4_srl_450_n7), .C2(u4_srl_450_n25), .A(u4_srl_450_n75), .ZN(
        u4_srl_450_n73) );
  AOI22_X1 u4_srl_450_U97 ( .A1(n2709), .A2(u4_srl_450_n41), .B1(n2710), .B2(
        u4_srl_450_n4), .ZN(u4_srl_450_n74) );
  OAI221_X1 u4_srl_450_U96 ( .B1(u4_srl_450_n39), .B2(u4_srl_450_n20), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n26), .A(u4_srl_450_n74), .ZN(
        u4_srl_450_n42) );
  MUX2_X1 u4_srl_450_U95 ( .A(u4_srl_450_n73), .B(u4_srl_450_n42), .S(
        u4_srl_450_n9), .Z(u4_N388) );
  AOI22_X1 u4_srl_450_U94 ( .A1(u4_srl_450_n41), .A2(fract_denorm[11]), .B1(
        u4_srl_450_n3), .B2(fract_denorm[10]), .ZN(u4_srl_450_n72) );
  OAI221_X1 u4_srl_450_U93 ( .B1(u4_srl_450_n39), .B2(u4_srl_450_n17), .C1(
        u4_srl_450_n24), .C2(u4_srl_450_n7), .A(u4_srl_450_n72), .ZN(
        u4_srl_450_n37) );
  AOI22_X1 u4_srl_450_U92 ( .A1(fract_denorm[15]), .A2(u4_srl_450_n41), .B1(
        fract_denorm[14]), .B2(u4_srl_450_n4), .ZN(u4_srl_450_n71) );
  OAI221_X1 u4_srl_450_U91 ( .B1(u4_srl_450_n39), .B2(u4_srl_450_n15), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n16), .A(u4_srl_450_n71), .ZN(
        u4_srl_450_n63) );
  MUX2_X1 u4_srl_450_U90 ( .A(u4_srl_450_n37), .B(u4_srl_450_n63), .S(
        u4_srl_450_n9), .Z(u4_N398) );
  AOI22_X1 u4_srl_450_U89 ( .A1(u4_srl_450_n41), .A2(fract_denorm[12]), .B1(
        u4_srl_450_n4), .B2(fract_denorm[11]), .ZN(u4_srl_450_n70) );
  OAI221_X1 u4_srl_450_U88 ( .B1(u4_srl_450_n39), .B2(u4_srl_450_n18), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n17), .A(u4_srl_450_n70), .ZN(
        u4_srl_450_n35) );
  AOI22_X1 u4_srl_450_U87 ( .A1(fract_denorm[16]), .A2(u4_srl_450_n6), .B1(
        fract_denorm[15]), .B2(u4_srl_450_n3), .ZN(u4_srl_450_n69) );
  OAI221_X1 u4_srl_450_U86 ( .B1(u4_srl_450_n39), .B2(u4_srl_450_n13), .C1(
        u4_srl_450_n7), .C2(u4_srl_450_n15), .A(u4_srl_450_n69), .ZN(
        u4_srl_450_n61) );
  MUX2_X1 u4_srl_450_U85 ( .A(u4_srl_450_n35), .B(u4_srl_450_n61), .S(
        u4_srl_450_n9), .Z(u4_N399) );
  AOI22_X1 u4_srl_450_U84 ( .A1(fract_denorm[13]), .A2(u4_srl_450_n6), .B1(
        u4_srl_450_n4), .B2(fract_denorm[12]), .ZN(u4_srl_450_n68) );
  OAI221_X1 u4_srl_450_U83 ( .B1(u4_srl_450_n39), .B2(u4_srl_450_n14), .C1(
        u4_srl_450_n7), .C2(u4_srl_450_n18), .A(u4_srl_450_n68), .ZN(
        u4_srl_450_n33) );
  AOI22_X1 u4_srl_450_U82 ( .A1(fract_denorm[17]), .A2(u4_srl_450_n41), .B1(
        fract_denorm[16]), .B2(u4_srl_450_n3), .ZN(u4_srl_450_n67) );
  OAI221_X1 u4_srl_450_U81 ( .B1(u4_srl_450_n39), .B2(u4_srl_450_n11), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n13), .A(u4_srl_450_n67), .ZN(
        u4_srl_450_n59) );
  MUX2_X1 u4_srl_450_U80 ( .A(u4_srl_450_n33), .B(u4_srl_450_n59), .S(
        u4_srl_450_n9), .Z(u4_N400) );
  AOI22_X1 u4_srl_450_U79 ( .A1(fract_denorm[14]), .A2(u4_srl_450_n41), .B1(
        fract_denorm[13]), .B2(u4_srl_450_n4), .ZN(u4_srl_450_n66) );
  OAI221_X1 u4_srl_450_U78 ( .B1(u4_srl_450_n39), .B2(u4_srl_450_n16), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n14), .A(u4_srl_450_n66), .ZN(
        u4_srl_450_n31) );
  AOI22_X1 u4_srl_450_U77 ( .A1(fract_denorm[18]), .A2(u4_srl_450_n6), .B1(
        fract_denorm[17]), .B2(u4_srl_450_n4), .ZN(u4_srl_450_n65) );
  OAI221_X1 u4_srl_450_U76 ( .B1(u4_srl_450_n39), .B2(u4_srl_450_n12), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n11), .A(u4_srl_450_n65), .ZN(
        u4_srl_450_n57) );
  MUX2_X1 u4_srl_450_U75 ( .A(u4_srl_450_n31), .B(u4_srl_450_n57), .S(
        u4_srl_450_n9), .Z(u4_N401) );
  AOI22_X1 u4_srl_450_U74 ( .A1(fract_denorm[19]), .A2(u4_srl_450_n6), .B1(
        fract_denorm[18]), .B2(u4_srl_450_n3), .ZN(u4_srl_450_n64) );
  OAI221_X1 u4_srl_450_U73 ( .B1(u4_srl_450_n39), .B2(u4_srl_450_n10), .C1(
        u4_srl_450_n7), .C2(u4_srl_450_n12), .A(u4_srl_450_n64), .ZN(
        u4_srl_450_n56) );
  MUX2_X1 u4_srl_450_U72 ( .A(u4_srl_450_n63), .B(u4_srl_450_n56), .S(
        u4_srl_450_n9), .Z(u4_N402) );
  AOI222_X1 u4_srl_450_U71 ( .A1(u4_srl_450_n6), .A2(fract_denorm[20]), .B1(
        u4_srl_450_n1), .B2(fract_denorm[21]), .C1(u4_srl_450_n3), .C2(
        fract_denorm[19]), .ZN(u4_srl_450_n54) );
  INV_X1 u4_srl_450_U70 ( .A(u4_srl_450_n54), .ZN(u4_srl_450_n62) );
  MUX2_X1 u4_srl_450_U69 ( .A(u4_srl_450_n61), .B(u4_srl_450_n62), .S(
        u4_srl_450_n9), .Z(u4_N403) );
  AOI22_X1 u4_srl_450_U68 ( .A1(u4_srl_450_n3), .A2(fract_denorm[20]), .B1(
        u4_srl_450_n6), .B2(fract_denorm[21]), .ZN(u4_srl_450_n50) );
  INV_X1 u4_srl_450_U67 ( .A(u4_srl_450_n50), .ZN(u4_srl_450_n60) );
  MUX2_X1 u4_srl_450_U66 ( .A(u4_srl_450_n59), .B(u4_srl_450_n60), .S(
        u4_srl_450_n9), .Z(u4_N404) );
  NOR2_X1 u4_srl_450_U65 ( .A1(u4_srl_450_n2), .A2(u4_srl_450_n10), .ZN(
        u4_srl_450_n58) );
  MUX2_X1 u4_srl_450_U64 ( .A(u4_srl_450_n57), .B(u4_srl_450_n58), .S(
        u4_srl_450_n9), .Z(u4_N405) );
  INV_X1 u4_srl_450_U63 ( .A(u4_srl_450_n56), .ZN(u4_srl_450_n55) );
  NOR2_X1 u4_srl_450_U62 ( .A1(u4_srl_450_n9), .A2(u4_srl_450_n55), .ZN(
        u4_N406) );
  NOR2_X1 u4_srl_450_U61 ( .A1(u4_srl_450_n9), .A2(u4_srl_450_n54), .ZN(
        u4_N407) );
  AOI22_X1 u4_srl_450_U60 ( .A1(n2706), .A2(u4_srl_450_n41), .B1(n2705), .B2(
        u4_srl_450_n3), .ZN(u4_srl_450_n53) );
  OAI221_X1 u4_srl_450_U59 ( .B1(u4_srl_450_n39), .B2(u4_srl_450_n28), .C1(
        u4_srl_450_n7), .C2(u4_srl_450_n29), .A(u4_srl_450_n53), .ZN(
        u4_srl_450_n51) );
  AOI22_X1 u4_srl_450_U58 ( .A1(n2708), .A2(u4_srl_450_n41), .B1(n2709), .B2(
        u4_srl_450_n4), .ZN(u4_srl_450_n52) );
  OAI221_X1 u4_srl_450_U57 ( .B1(u4_srl_450_n39), .B2(u4_srl_450_n21), .C1(
        u4_srl_450_n7), .C2(u4_srl_450_n20), .A(u4_srl_450_n52), .ZN(
        u4_srl_450_n38) );
  MUX2_X1 u4_srl_450_U56 ( .A(u4_srl_450_n51), .B(u4_srl_450_n38), .S(
        u4_srl_450_n9), .Z(u4_N389) );
  NOR2_X1 u4_srl_450_U55 ( .A1(u4_srl_450_n9), .A2(u4_srl_450_n50), .ZN(
        u4_N408) );
  NOR3_X1 u4_srl_450_U54 ( .A1(u4_srl_450_n10), .A2(u4_srl_450_n9), .A3(
        u4_srl_450_n2), .ZN(u4_N409) );
  AOI22_X1 u4_srl_450_U53 ( .A1(n2711), .A2(u4_srl_450_n6), .B1(n2706), .B2(
        u4_srl_450_n4), .ZN(u4_srl_450_n49) );
  OAI221_X1 u4_srl_450_U52 ( .B1(u4_srl_450_n39), .B2(u4_srl_450_n27), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n28), .A(u4_srl_450_n49), .ZN(
        u4_srl_450_n47) );
  AOI22_X1 u4_srl_450_U51 ( .A1(n2704), .A2(u4_srl_450_n6), .B1(n2708), .B2(
        u4_srl_450_n3), .ZN(u4_srl_450_n48) );
  OAI221_X1 u4_srl_450_U50 ( .B1(u4_srl_450_n39), .B2(u4_srl_450_n22), .C1(
        u4_srl_450_n7), .C2(u4_srl_450_n21), .A(u4_srl_450_n48), .ZN(
        u4_srl_450_n36) );
  MUX2_X1 u4_srl_450_U49 ( .A(u4_srl_450_n47), .B(u4_srl_450_n36), .S(
        u4_srl_450_n9), .Z(u4_N390) );
  AOI22_X1 u4_srl_450_U48 ( .A1(n2710), .A2(u4_srl_450_n41), .B1(n2711), .B2(
        u4_srl_450_n3), .ZN(u4_srl_450_n46) );
  OAI221_X1 u4_srl_450_U47 ( .B1(u4_srl_450_n39), .B2(u4_srl_450_n26), .C1(
        u4_srl_450_n7), .C2(u4_srl_450_n27), .A(u4_srl_450_n46), .ZN(
        u4_srl_450_n44) );
  AOI22_X1 u4_srl_450_U46 ( .A1(fract_denorm[8]), .A2(u4_srl_450_n41), .B1(
        n2704), .B2(u4_srl_450_n4), .ZN(u4_srl_450_n45) );
  OAI221_X1 u4_srl_450_U45 ( .B1(u4_srl_450_n39), .B2(u4_srl_450_n19), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n22), .A(u4_srl_450_n45), .ZN(
        u4_srl_450_n34) );
  MUX2_X1 u4_srl_450_U44 ( .A(u4_srl_450_n44), .B(u4_srl_450_n34), .S(
        u4_srl_450_n9), .Z(u4_N391) );
  AOI22_X1 u4_srl_450_U43 ( .A1(fract_denorm[9]), .A2(u4_srl_450_n6), .B1(
        fract_denorm[8]), .B2(u4_srl_450_n4), .ZN(u4_srl_450_n43) );
  OAI221_X1 u4_srl_450_U42 ( .B1(u4_srl_450_n39), .B2(u4_srl_450_n23), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n19), .A(u4_srl_450_n43), .ZN(
        u4_srl_450_n32) );
  MUX2_X1 u4_srl_450_U41 ( .A(u4_srl_450_n42), .B(u4_srl_450_n32), .S(
        u4_srl_450_n9), .Z(u4_N392) );
  AOI22_X1 u4_srl_450_U40 ( .A1(fract_denorm[10]), .A2(u4_srl_450_n6), .B1(
        fract_denorm[9]), .B2(u4_srl_450_n3), .ZN(u4_srl_450_n40) );
  OAI221_X1 u4_srl_450_U39 ( .B1(u4_srl_450_n39), .B2(u4_srl_450_n24), .C1(
        u4_srl_450_n8), .C2(u4_srl_450_n23), .A(u4_srl_450_n40), .ZN(
        u4_srl_450_n30) );
  MUX2_X1 u4_srl_450_U38 ( .A(u4_srl_450_n38), .B(u4_srl_450_n30), .S(
        u4_srl_450_n9), .Z(u4_N393) );
  MUX2_X1 u4_srl_450_U37 ( .A(u4_srl_450_n36), .B(u4_srl_450_n37), .S(
        u4_srl_450_n9), .Z(u4_N394) );
  MUX2_X1 u4_srl_450_U36 ( .A(u4_srl_450_n34), .B(u4_srl_450_n35), .S(
        u4_srl_450_n9), .Z(u4_N395) );
  MUX2_X1 u4_srl_450_U35 ( .A(u4_srl_450_n32), .B(u4_srl_450_n33), .S(
        u4_srl_450_n9), .Z(u4_N396) );
  MUX2_X1 u4_srl_450_U34 ( .A(u4_srl_450_n30), .B(u4_srl_450_n31), .S(
        u4_srl_450_n9), .Z(u4_N397) );
  INV_X4 u4_srl_450_U33 ( .A(n2711), .ZN(u4_srl_450_n29) );
  INV_X4 u4_srl_450_U32 ( .A(n2710), .ZN(u4_srl_450_n28) );
  INV_X4 u4_srl_450_U31 ( .A(n2709), .ZN(u4_srl_450_n27) );
  INV_X4 u4_srl_450_U30 ( .A(n2708), .ZN(u4_srl_450_n26) );
  INV_X4 u4_srl_450_U29 ( .A(n2706), .ZN(u4_srl_450_n25) );
  INV_X4 u4_srl_450_U28 ( .A(fract_denorm[12]), .ZN(u4_srl_450_n24) );
  INV_X4 u4_srl_450_U27 ( .A(fract_denorm[11]), .ZN(u4_srl_450_n23) );
  INV_X4 u4_srl_450_U26 ( .A(fract_denorm[9]), .ZN(u4_srl_450_n22) );
  INV_X4 u4_srl_450_U25 ( .A(fract_denorm[8]), .ZN(u4_srl_450_n21) );
  INV_X4 u4_srl_450_U24 ( .A(n2704), .ZN(u4_srl_450_n20) );
  INV_X4 u4_srl_450_U23 ( .A(fract_denorm[10]), .ZN(u4_srl_450_n19) );
  INV_X4 u4_srl_450_U22 ( .A(fract_denorm[14]), .ZN(u4_srl_450_n18) );
  INV_X4 u4_srl_450_U21 ( .A(fract_denorm[13]), .ZN(u4_srl_450_n17) );
  INV_X4 u4_srl_450_U20 ( .A(fract_denorm[16]), .ZN(u4_srl_450_n16) );
  INV_X4 u4_srl_450_U19 ( .A(fract_denorm[17]), .ZN(u4_srl_450_n15) );
  INV_X4 u4_srl_450_U18 ( .A(fract_denorm[15]), .ZN(u4_srl_450_n14) );
  INV_X4 u4_srl_450_U17 ( .A(fract_denorm[18]), .ZN(u4_srl_450_n13) );
  INV_X4 u4_srl_450_U16 ( .A(fract_denorm[20]), .ZN(u4_srl_450_n12) );
  INV_X4 u4_srl_450_U15 ( .A(fract_denorm[19]), .ZN(u4_srl_450_n11) );
  INV_X4 u4_srl_450_U14 ( .A(fract_denorm[21]), .ZN(u4_srl_450_n10) );
  NOR2_X2 u4_srl_450_U13 ( .A1(u4_srl_450_n76), .A2(u4_shift_right[1]), .ZN(
        u4_srl_450_n41) );
  INV_X4 u4_srl_450_U12 ( .A(u4_srl_450_n41), .ZN(u4_srl_450_n5) );
  INV_X4 u4_srl_450_U11 ( .A(u4_srl_450_n1), .ZN(u4_srl_450_n7) );
  INV_X4 u4_srl_450_U10 ( .A(u4_srl_450_n1), .ZN(u4_srl_450_n8) );
  INV_X4 u4_srl_450_U9 ( .A(u4_srl_450_n2), .ZN(u4_srl_450_n4) );
  OR2_X4 u4_srl_450_U8 ( .A1(u4_shift_right[0]), .A2(u4_shift_right[1]), .ZN(
        u4_srl_450_n2) );
  AND2_X4 u4_srl_450_U7 ( .A1(u4_shift_right[1]), .A2(u4_srl_450_n76), .ZN(
        u4_srl_450_n1) );
  BUF_X4 u4_srl_450_U6 ( .A(u4_shift_right[2]), .Z(u4_srl_450_n9) );
  INV_X4 u4_srl_450_U5 ( .A(u4_srl_450_n2), .ZN(u4_srl_450_n3) );
  INV_X4 u4_srl_450_U4 ( .A(u4_srl_450_n5), .ZN(u4_srl_450_n6) );
  NAND2_X2 u4_srl_450_U3 ( .A1(u4_shift_right[1]), .A2(u4_shift_right[0]), 
        .ZN(u4_srl_450_n39) );
  AND2_X1 u4_sll_451_U17 ( .A1(n2707), .A2(u4_sll_451_n1), .ZN(
        u4_sll_451_ML_int_1__0_) );
  NAND2_X1 u4_sll_451_U16 ( .A1(u4_sll_451_ML_int_1__0_), .A2(u4_sll_451_n3), 
        .ZN(u4_sll_451_n8) );
  INV_X1 u4_sll_451_U15 ( .A(u4_sll_451_n8), .ZN(u4_sll_451_ML_int_2__0_) );
  NAND2_X1 u4_sll_451_U14 ( .A1(u4_sll_451_ML_int_1__1_), .A2(u4_sll_451_n3), 
        .ZN(u4_sll_451_n7) );
  INV_X1 u4_sll_451_U13 ( .A(u4_sll_451_n7), .ZN(u4_sll_451_ML_int_2__1_) );
  NOR2_X1 u4_sll_451_U12 ( .A1(u4_sll_451_n6), .A2(u4_sll_451_n8), .ZN(u4_N412) );
  NOR2_X1 u4_sll_451_U11 ( .A1(u4_sll_451_n6), .A2(u4_sll_451_n7), .ZN(u4_N413) );
  AND2_X1 u4_sll_451_U10 ( .A1(u4_sll_451_ML_int_2__2_), .A2(u4_sll_451_n5), 
        .ZN(u4_N414) );
  AND2_X1 u4_sll_451_U9 ( .A1(u4_sll_451_ML_int_2__3_), .A2(u4_sll_451_n5), 
        .ZN(u4_N415) );
  INV_X4 u4_sll_451_U8 ( .A(u4_shift_left[0]), .ZN(u4_sll_451_n1) );
  INV_X4 u4_sll_451_U7 ( .A(u4_sll_451_n1), .ZN(u4_sll_451_n2) );
  INV_X4 u4_sll_451_U6 ( .A(u4_shift_left[2]), .ZN(u4_sll_451_n5) );
  INV_X4 u4_sll_451_U5 ( .A(u4_sll_451_n5), .ZN(u4_sll_451_n6) );
  INV_X4 u4_sll_451_U4 ( .A(u4_shift_left[1]), .ZN(u4_sll_451_n3) );
  INV_X4 u4_sll_451_U3 ( .A(u4_sll_451_n3), .ZN(u4_sll_451_n4) );
  MUX2_X2 u4_sll_451_M1_0_1 ( .A(n2705), .B(n2707), .S(u4_shift_left[0]), .Z(
        u4_sll_451_ML_int_1__1_) );
  MUX2_X2 u4_sll_451_M1_0_2 ( .A(n2706), .B(n2705), .S(u4_shift_left[0]), .Z(
        u4_sll_451_ML_int_1__2_) );
  MUX2_X2 u4_sll_451_M1_0_3 ( .A(n2711), .B(n2706), .S(u4_sll_451_n2), .Z(
        u4_sll_451_ML_int_1__3_) );
  MUX2_X2 u4_sll_451_M1_0_4 ( .A(n2710), .B(n2711), .S(u4_sll_451_n2), .Z(
        u4_sll_451_ML_int_1__4_) );
  MUX2_X2 u4_sll_451_M1_0_5 ( .A(n2709), .B(n2710), .S(u4_sll_451_n2), .Z(
        u4_sll_451_ML_int_1__5_) );
  MUX2_X2 u4_sll_451_M1_0_6 ( .A(n2708), .B(n2709), .S(u4_shift_left[0]), .Z(
        u4_sll_451_ML_int_1__6_) );
  MUX2_X2 u4_sll_451_M1_0_7 ( .A(n2704), .B(n2708), .S(u4_shift_left[0]), .Z(
        u4_sll_451_ML_int_1__7_) );
  MUX2_X2 u4_sll_451_M1_0_8 ( .A(fract_denorm[8]), .B(n2704), .S(
        u4_shift_left[0]), .Z(u4_sll_451_ML_int_1__8_) );
  MUX2_X2 u4_sll_451_M1_0_9 ( .A(fract_denorm[9]), .B(fract_denorm[8]), .S(
        u4_shift_left[0]), .Z(u4_sll_451_ML_int_1__9_) );
  MUX2_X2 u4_sll_451_M1_0_10 ( .A(fract_denorm[10]), .B(fract_denorm[9]), .S(
        u4_shift_left[0]), .Z(u4_sll_451_ML_int_1__10_) );
  MUX2_X2 u4_sll_451_M1_0_11 ( .A(fract_denorm[11]), .B(fract_denorm[10]), .S(
        u4_shift_left[0]), .Z(u4_sll_451_ML_int_1__11_) );
  MUX2_X2 u4_sll_451_M1_0_12 ( .A(fract_denorm[12]), .B(fract_denorm[11]), .S(
        u4_sll_451_n2), .Z(u4_sll_451_ML_int_1__12_) );
  MUX2_X2 u4_sll_451_M1_0_13 ( .A(fract_denorm[13]), .B(fract_denorm[12]), .S(
        u4_sll_451_n2), .Z(u4_sll_451_ML_int_1__13_) );
  MUX2_X2 u4_sll_451_M1_0_14 ( .A(fract_denorm[14]), .B(fract_denorm[13]), .S(
        u4_sll_451_n2), .Z(u4_sll_451_ML_int_1__14_) );
  MUX2_X2 u4_sll_451_M1_0_15 ( .A(fract_denorm[15]), .B(fract_denorm[14]), .S(
        u4_sll_451_n2), .Z(u4_sll_451_ML_int_1__15_) );
  MUX2_X2 u4_sll_451_M1_0_16 ( .A(fract_denorm[16]), .B(fract_denorm[15]), .S(
        u4_sll_451_n2), .Z(u4_sll_451_ML_int_1__16_) );
  MUX2_X2 u4_sll_451_M1_0_17 ( .A(fract_denorm[17]), .B(fract_denorm[16]), .S(
        u4_sll_451_n2), .Z(u4_sll_451_ML_int_1__17_) );
  MUX2_X2 u4_sll_451_M1_0_18 ( .A(fract_denorm[18]), .B(fract_denorm[17]), .S(
        u4_sll_451_n2), .Z(u4_sll_451_ML_int_1__18_) );
  MUX2_X2 u4_sll_451_M1_0_19 ( .A(fract_denorm[19]), .B(fract_denorm[18]), .S(
        u4_sll_451_n2), .Z(u4_sll_451_ML_int_1__19_) );
  MUX2_X2 u4_sll_451_M1_0_20 ( .A(fract_denorm[20]), .B(fract_denorm[19]), .S(
        u4_sll_451_n2), .Z(u4_sll_451_ML_int_1__20_) );
  MUX2_X2 u4_sll_451_M1_0_21 ( .A(fract_denorm[21]), .B(fract_denorm[20]), .S(
        u4_sll_451_n2), .Z(u4_sll_451_ML_int_1__21_) );
  MUX2_X2 u4_sll_451_M1_1_2 ( .A(u4_sll_451_ML_int_1__2_), .B(
        u4_sll_451_ML_int_1__0_), .S(u4_sll_451_n4), .Z(
        u4_sll_451_ML_int_2__2_) );
  MUX2_X2 u4_sll_451_M1_1_3 ( .A(u4_sll_451_ML_int_1__3_), .B(
        u4_sll_451_ML_int_1__1_), .S(u4_sll_451_n4), .Z(
        u4_sll_451_ML_int_2__3_) );
  MUX2_X2 u4_sll_451_M1_1_4 ( .A(u4_sll_451_ML_int_1__4_), .B(
        u4_sll_451_ML_int_1__2_), .S(u4_sll_451_n4), .Z(
        u4_sll_451_ML_int_2__4_) );
  MUX2_X2 u4_sll_451_M1_1_5 ( .A(u4_sll_451_ML_int_1__5_), .B(
        u4_sll_451_ML_int_1__3_), .S(u4_sll_451_n4), .Z(
        u4_sll_451_ML_int_2__5_) );
  MUX2_X2 u4_sll_451_M1_1_6 ( .A(u4_sll_451_ML_int_1__6_), .B(
        u4_sll_451_ML_int_1__4_), .S(u4_sll_451_n4), .Z(
        u4_sll_451_ML_int_2__6_) );
  MUX2_X2 u4_sll_451_M1_1_7 ( .A(u4_sll_451_ML_int_1__7_), .B(
        u4_sll_451_ML_int_1__5_), .S(u4_sll_451_n4), .Z(
        u4_sll_451_ML_int_2__7_) );
  MUX2_X2 u4_sll_451_M1_1_8 ( .A(u4_sll_451_ML_int_1__8_), .B(
        u4_sll_451_ML_int_1__6_), .S(u4_sll_451_n4), .Z(
        u4_sll_451_ML_int_2__8_) );
  MUX2_X2 u4_sll_451_M1_1_9 ( .A(u4_sll_451_ML_int_1__9_), .B(
        u4_sll_451_ML_int_1__7_), .S(u4_sll_451_n4), .Z(
        u4_sll_451_ML_int_2__9_) );
  MUX2_X2 u4_sll_451_M1_1_10 ( .A(u4_sll_451_ML_int_1__10_), .B(
        u4_sll_451_ML_int_1__8_), .S(u4_sll_451_n4), .Z(
        u4_sll_451_ML_int_2__10_) );
  MUX2_X2 u4_sll_451_M1_1_11 ( .A(u4_sll_451_ML_int_1__11_), .B(
        u4_sll_451_ML_int_1__9_), .S(u4_sll_451_n4), .Z(
        u4_sll_451_ML_int_2__11_) );
  MUX2_X2 u4_sll_451_M1_1_12 ( .A(u4_sll_451_ML_int_1__12_), .B(
        u4_sll_451_ML_int_1__10_), .S(u4_sll_451_n4), .Z(
        u4_sll_451_ML_int_2__12_) );
  MUX2_X2 u4_sll_451_M1_1_13 ( .A(u4_sll_451_ML_int_1__13_), .B(
        u4_sll_451_ML_int_1__11_), .S(u4_sll_451_n4), .Z(
        u4_sll_451_ML_int_2__13_) );
  MUX2_X2 u4_sll_451_M1_1_14 ( .A(u4_sll_451_ML_int_1__14_), .B(
        u4_sll_451_ML_int_1__12_), .S(u4_sll_451_n4), .Z(
        u4_sll_451_ML_int_2__14_) );
  MUX2_X2 u4_sll_451_M1_1_15 ( .A(u4_sll_451_ML_int_1__15_), .B(
        u4_sll_451_ML_int_1__13_), .S(u4_sll_451_n4), .Z(
        u4_sll_451_ML_int_2__15_) );
  MUX2_X2 u4_sll_451_M1_1_16 ( .A(u4_sll_451_ML_int_1__16_), .B(
        u4_sll_451_ML_int_1__14_), .S(u4_sll_451_n4), .Z(
        u4_sll_451_ML_int_2__16_) );
  MUX2_X2 u4_sll_451_M1_1_17 ( .A(u4_sll_451_ML_int_1__17_), .B(
        u4_sll_451_ML_int_1__15_), .S(u4_sll_451_n4), .Z(
        u4_sll_451_ML_int_2__17_) );
  MUX2_X2 u4_sll_451_M1_1_18 ( .A(u4_sll_451_ML_int_1__18_), .B(
        u4_sll_451_ML_int_1__16_), .S(u4_sll_451_n4), .Z(
        u4_sll_451_ML_int_2__18_) );
  MUX2_X2 u4_sll_451_M1_1_19 ( .A(u4_sll_451_ML_int_1__19_), .B(
        u4_sll_451_ML_int_1__17_), .S(u4_sll_451_n4), .Z(
        u4_sll_451_ML_int_2__19_) );
  MUX2_X2 u4_sll_451_M1_1_20 ( .A(u4_sll_451_ML_int_1__20_), .B(
        u4_sll_451_ML_int_1__18_), .S(u4_sll_451_n4), .Z(
        u4_sll_451_ML_int_2__20_) );
  MUX2_X2 u4_sll_451_M1_1_21 ( .A(u4_sll_451_ML_int_1__21_), .B(
        u4_sll_451_ML_int_1__19_), .S(u4_sll_451_n4), .Z(
        u4_sll_451_ML_int_2__21_) );
  MUX2_X2 u4_sll_451_M1_2_4 ( .A(u4_sll_451_ML_int_2__4_), .B(
        u4_sll_451_ML_int_2__0_), .S(u4_sll_451_n6), .Z(u4_N416) );
  MUX2_X2 u4_sll_451_M1_2_5 ( .A(u4_sll_451_ML_int_2__5_), .B(
        u4_sll_451_ML_int_2__1_), .S(u4_sll_451_n6), .Z(u4_N417) );
  MUX2_X2 u4_sll_451_M1_2_6 ( .A(u4_sll_451_ML_int_2__6_), .B(
        u4_sll_451_ML_int_2__2_), .S(u4_sll_451_n6), .Z(u4_N418) );
  MUX2_X2 u4_sll_451_M1_2_7 ( .A(u4_sll_451_ML_int_2__7_), .B(
        u4_sll_451_ML_int_2__3_), .S(u4_sll_451_n6), .Z(u4_N419) );
  MUX2_X2 u4_sll_451_M1_2_8 ( .A(u4_sll_451_ML_int_2__8_), .B(
        u4_sll_451_ML_int_2__4_), .S(u4_sll_451_n6), .Z(u4_N420) );
  MUX2_X2 u4_sll_451_M1_2_9 ( .A(u4_sll_451_ML_int_2__9_), .B(
        u4_sll_451_ML_int_2__5_), .S(u4_sll_451_n6), .Z(u4_N421) );
  MUX2_X2 u4_sll_451_M1_2_10 ( .A(u4_sll_451_ML_int_2__10_), .B(
        u4_sll_451_ML_int_2__6_), .S(u4_sll_451_n6), .Z(u4_N422) );
  MUX2_X2 u4_sll_451_M1_2_11 ( .A(u4_sll_451_ML_int_2__11_), .B(
        u4_sll_451_ML_int_2__7_), .S(u4_sll_451_n6), .Z(u4_N423) );
  MUX2_X2 u4_sll_451_M1_2_12 ( .A(u4_sll_451_ML_int_2__12_), .B(
        u4_sll_451_ML_int_2__8_), .S(u4_sll_451_n6), .Z(u4_N424) );
  MUX2_X2 u4_sll_451_M1_2_13 ( .A(u4_sll_451_ML_int_2__13_), .B(
        u4_sll_451_ML_int_2__9_), .S(u4_sll_451_n6), .Z(u4_N425) );
  MUX2_X2 u4_sll_451_M1_2_14 ( .A(u4_sll_451_ML_int_2__14_), .B(
        u4_sll_451_ML_int_2__10_), .S(u4_sll_451_n6), .Z(u4_N426) );
  MUX2_X2 u4_sll_451_M1_2_15 ( .A(u4_sll_451_ML_int_2__15_), .B(
        u4_sll_451_ML_int_2__11_), .S(u4_sll_451_n6), .Z(u4_N427) );
  MUX2_X2 u4_sll_451_M1_2_16 ( .A(u4_sll_451_ML_int_2__16_), .B(
        u4_sll_451_ML_int_2__12_), .S(u4_sll_451_n6), .Z(u4_N428) );
  MUX2_X2 u4_sll_451_M1_2_17 ( .A(u4_sll_451_ML_int_2__17_), .B(
        u4_sll_451_ML_int_2__13_), .S(u4_sll_451_n6), .Z(u4_N429) );
  MUX2_X2 u4_sll_451_M1_2_18 ( .A(u4_sll_451_ML_int_2__18_), .B(
        u4_sll_451_ML_int_2__14_), .S(u4_sll_451_n6), .Z(u4_N430) );
  MUX2_X2 u4_sll_451_M1_2_19 ( .A(u4_sll_451_ML_int_2__19_), .B(
        u4_sll_451_ML_int_2__15_), .S(u4_sll_451_n6), .Z(u4_N431) );
  MUX2_X2 u4_sll_451_M1_2_20 ( .A(u4_sll_451_ML_int_2__20_), .B(
        u4_sll_451_ML_int_2__16_), .S(u4_sll_451_n6), .Z(u4_N432) );
  MUX2_X2 u4_sll_451_M1_2_21 ( .A(u4_sll_451_ML_int_2__21_), .B(
        u4_sll_451_ML_int_2__17_), .S(u4_sll_451_n6), .Z(u4_N433) );
  AND2_X1 u4_sll_479_U19 ( .A1(n2707), .A2(u4_sll_479_n8), .ZN(
        u4_sll_479_ML_int_1__0_) );
  NOR2_X1 u4_sll_479_U18 ( .A1(u4_sll_479_n2), .A2(u4_sll_479_n1), .ZN(
        u4_sll_479_n11) );
  AND2_X1 u4_sll_479_U17 ( .A1(u4_sll_479_n11), .A2(u4_sll_479_ML_int_1__0_), 
        .ZN(u4_sll_479_ML_int_3__0_) );
  AND2_X1 u4_sll_479_U16 ( .A1(u4_sll_479_ML_int_1__1_), .A2(u4_sll_479_n11), 
        .ZN(u4_sll_479_ML_int_3__1_) );
  AND2_X1 u4_sll_479_U15 ( .A1(u4_sll_479_ML_int_2__2_), .A2(u4_sll_479_n10), 
        .ZN(u4_sll_479_ML_int_3__2_) );
  AND2_X1 u4_sll_479_U14 ( .A1(u4_sll_479_ML_int_2__3_), .A2(u4_sll_479_n10), 
        .ZN(u4_sll_479_ML_int_3__3_) );
  AND2_X1 u4_sll_479_U13 ( .A1(u4_sll_479_ML_int_3__7_), .A2(u4_sll_479_n9), 
        .ZN(u4_sll_479_ML_int_4__7_) );
  INV_X4 u4_sll_479_U12 ( .A(u4_sll_479_n1), .ZN(u4_sll_479_n10) );
  INV_X4 u4_sll_479_U11 ( .A(u4_f2i_shft_3_), .ZN(u4_sll_479_n9) );
  INV_X4 u4_sll_479_U10 ( .A(u4_sll_479_n4), .ZN(u4_sll_479_n3) );
  INV_X4 u4_sll_479_U9 ( .A(u4_sll_479_n4), .ZN(u4_sll_479_n2) );
  INV_X4 u4_sll_479_U8 ( .A(u4_f2i_shft_1_), .ZN(u4_sll_479_n4) );
  INV_X4 u4_sll_479_U7 ( .A(u4_sll_479_n5), .ZN(u4_sll_479_n8) );
  INV_X4 u4_sll_479_U6 ( .A(u4_sll_479_n6), .ZN(u4_sll_479_n5) );
  INV_X4 u4_sll_479_U5 ( .A(u4_sll_479_n8), .ZN(u4_sll_479_n7) );
  INV_X4 u4_sll_479_U4 ( .A(u4_f2i_shft_0_), .ZN(u4_sll_479_n6) );
  BUF_X4 u4_sll_479_U3 ( .A(u4_f2i_shft_2_), .Z(u4_sll_479_n1) );
  MUX2_X2 u4_sll_479_M1_0_1 ( .A(n2705), .B(n2707), .S(u4_sll_479_n7), .Z(
        u4_sll_479_ML_int_1__1_) );
  MUX2_X2 u4_sll_479_M1_0_2 ( .A(n2706), .B(n2705), .S(u4_sll_479_n7), .Z(
        u4_sll_479_ML_int_1__2_) );
  MUX2_X2 u4_sll_479_M1_0_3 ( .A(n2711), .B(n2706), .S(u4_sll_479_n7), .Z(
        u4_sll_479_ML_int_1__3_) );
  MUX2_X2 u4_sll_479_M1_0_4 ( .A(n2710), .B(n2711), .S(u4_sll_479_n7), .Z(
        u4_sll_479_ML_int_1__4_) );
  MUX2_X2 u4_sll_479_M1_0_5 ( .A(n2709), .B(n2710), .S(u4_sll_479_n7), .Z(
        u4_sll_479_ML_int_1__5_) );
  MUX2_X2 u4_sll_479_M1_0_6 ( .A(n2708), .B(n2709), .S(u4_sll_479_n7), .Z(
        u4_sll_479_ML_int_1__6_) );
  MUX2_X2 u4_sll_479_M1_0_7 ( .A(n2704), .B(n2708), .S(u4_sll_479_n7), .Z(
        u4_sll_479_ML_int_1__7_) );
  MUX2_X2 u4_sll_479_M1_0_8 ( .A(fract_denorm[8]), .B(n2704), .S(u4_sll_479_n7), .Z(u4_sll_479_ML_int_1__8_) );
  MUX2_X2 u4_sll_479_M1_0_9 ( .A(fract_denorm[9]), .B(fract_denorm[8]), .S(
        u4_sll_479_n7), .Z(u4_sll_479_ML_int_1__9_) );
  MUX2_X2 u4_sll_479_M1_0_10 ( .A(fract_denorm[10]), .B(fract_denorm[9]), .S(
        u4_sll_479_n7), .Z(u4_sll_479_ML_int_1__10_) );
  MUX2_X2 u4_sll_479_M1_0_11 ( .A(fract_denorm[11]), .B(fract_denorm[10]), .S(
        u4_sll_479_n7), .Z(u4_sll_479_ML_int_1__11_) );
  MUX2_X2 u4_sll_479_M1_0_12 ( .A(fract_denorm[12]), .B(fract_denorm[11]), .S(
        u4_f2i_shft_0_), .Z(u4_sll_479_ML_int_1__12_) );
  MUX2_X2 u4_sll_479_M1_0_13 ( .A(fract_denorm[13]), .B(fract_denorm[12]), .S(
        u4_sll_479_n7), .Z(u4_sll_479_ML_int_1__13_) );
  MUX2_X2 u4_sll_479_M1_0_14 ( .A(fract_denorm[14]), .B(fract_denorm[13]), .S(
        u4_f2i_shft_0_), .Z(u4_sll_479_ML_int_1__14_) );
  MUX2_X2 u4_sll_479_M1_0_15 ( .A(fract_denorm[15]), .B(fract_denorm[14]), .S(
        u4_sll_479_n7), .Z(u4_sll_479_ML_int_1__15_) );
  MUX2_X2 u4_sll_479_M1_0_16 ( .A(fract_denorm[16]), .B(fract_denorm[15]), .S(
        u4_f2i_shft_0_), .Z(u4_sll_479_ML_int_1__16_) );
  MUX2_X2 u4_sll_479_M1_0_17 ( .A(fract_denorm[17]), .B(fract_denorm[16]), .S(
        u4_sll_479_n5), .Z(u4_sll_479_ML_int_1__17_) );
  MUX2_X2 u4_sll_479_M1_0_18 ( .A(fract_denorm[18]), .B(fract_denorm[17]), .S(
        u4_f2i_shft_0_), .Z(u4_sll_479_ML_int_1__18_) );
  MUX2_X2 u4_sll_479_M1_0_19 ( .A(fract_denorm[19]), .B(fract_denorm[18]), .S(
        u4_sll_479_n7), .Z(u4_sll_479_ML_int_1__19_) );
  MUX2_X2 u4_sll_479_M1_0_20 ( .A(fract_denorm[20]), .B(fract_denorm[19]), .S(
        u4_f2i_shft_0_), .Z(u4_sll_479_ML_int_1__20_) );
  MUX2_X2 u4_sll_479_M1_0_21 ( .A(fract_denorm[21]), .B(fract_denorm[20]), .S(
        u4_sll_479_n7), .Z(u4_sll_479_ML_int_1__21_) );
  MUX2_X2 u4_sll_479_M1_0_22 ( .A(fract_denorm[21]), .B(fract_denorm[21]), .S(
        u4_f2i_shft_0_), .Z(u4_sll_479_ML_int_1__22_) );
  MUX2_X2 u4_sll_479_M1_0_23 ( .A(fract_denorm[21]), .B(fract_denorm[21]), .S(
        u4_sll_479_n7), .Z(u4_sll_479_ML_int_1__23_) );
  MUX2_X2 u4_sll_479_M1_0_24 ( .A(fract_denorm[21]), .B(fract_denorm[21]), .S(
        u4_f2i_shft_0_), .Z(u4_sll_479_ML_int_1__24_) );
  MUX2_X2 u4_sll_479_M1_0_25 ( .A(fract_denorm[21]), .B(fract_denorm[21]), .S(
        u4_f2i_shft_0_), .Z(u4_sll_479_ML_int_1__25_) );
  MUX2_X2 u4_sll_479_M1_0_26 ( .A(fract_denorm[21]), .B(fract_denorm[21]), .S(
        u4_f2i_shft_0_), .Z(u4_sll_479_ML_int_1__26_) );
  MUX2_X2 u4_sll_479_M1_0_27 ( .A(fract_denorm[21]), .B(fract_denorm[21]), .S(
        u4_f2i_shft_0_), .Z(u4_sll_479_ML_int_1__27_) );
  MUX2_X2 u4_sll_479_M1_1_2 ( .A(u4_sll_479_ML_int_1__2_), .B(
        u4_sll_479_ML_int_1__0_), .S(u4_f2i_shft_1_), .Z(
        u4_sll_479_ML_int_2__2_) );
  MUX2_X2 u4_sll_479_M1_1_3 ( .A(u4_sll_479_ML_int_1__3_), .B(
        u4_sll_479_ML_int_1__1_), .S(u4_f2i_shft_1_), .Z(
        u4_sll_479_ML_int_2__3_) );
  MUX2_X2 u4_sll_479_M1_1_4 ( .A(u4_sll_479_ML_int_1__4_), .B(
        u4_sll_479_ML_int_1__2_), .S(u4_sll_479_n3), .Z(
        u4_sll_479_ML_int_2__4_) );
  MUX2_X2 u4_sll_479_M1_1_5 ( .A(u4_sll_479_ML_int_1__5_), .B(
        u4_sll_479_ML_int_1__3_), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_2__5_) );
  MUX2_X2 u4_sll_479_M1_1_6 ( .A(u4_sll_479_ML_int_1__6_), .B(
        u4_sll_479_ML_int_1__4_), .S(u4_sll_479_n3), .Z(
        u4_sll_479_ML_int_2__6_) );
  MUX2_X2 u4_sll_479_M1_1_7 ( .A(u4_sll_479_ML_int_1__7_), .B(
        u4_sll_479_ML_int_1__5_), .S(u4_sll_479_n3), .Z(
        u4_sll_479_ML_int_2__7_) );
  MUX2_X2 u4_sll_479_M1_1_8 ( .A(u4_sll_479_ML_int_1__8_), .B(
        u4_sll_479_ML_int_1__6_), .S(u4_sll_479_n3), .Z(
        u4_sll_479_ML_int_2__8_) );
  MUX2_X2 u4_sll_479_M1_1_9 ( .A(u4_sll_479_ML_int_1__9_), .B(
        u4_sll_479_ML_int_1__7_), .S(u4_sll_479_n3), .Z(
        u4_sll_479_ML_int_2__9_) );
  MUX2_X2 u4_sll_479_M1_1_10 ( .A(u4_sll_479_ML_int_1__10_), .B(
        u4_sll_479_ML_int_1__8_), .S(u4_sll_479_n3), .Z(
        u4_sll_479_ML_int_2__10_) );
  MUX2_X2 u4_sll_479_M1_1_11 ( .A(u4_sll_479_ML_int_1__11_), .B(
        u4_sll_479_ML_int_1__9_), .S(u4_sll_479_n3), .Z(
        u4_sll_479_ML_int_2__11_) );
  MUX2_X2 u4_sll_479_M1_1_12 ( .A(u4_sll_479_ML_int_1__12_), .B(
        u4_sll_479_ML_int_1__10_), .S(u4_sll_479_n3), .Z(
        u4_sll_479_ML_int_2__12_) );
  MUX2_X2 u4_sll_479_M1_1_13 ( .A(u4_sll_479_ML_int_1__13_), .B(
        u4_sll_479_ML_int_1__11_), .S(u4_sll_479_n3), .Z(
        u4_sll_479_ML_int_2__13_) );
  MUX2_X2 u4_sll_479_M1_1_14 ( .A(u4_sll_479_ML_int_1__14_), .B(
        u4_sll_479_ML_int_1__12_), .S(u4_sll_479_n3), .Z(
        u4_sll_479_ML_int_2__14_) );
  MUX2_X2 u4_sll_479_M1_1_15 ( .A(u4_sll_479_ML_int_1__15_), .B(
        u4_sll_479_ML_int_1__13_), .S(u4_sll_479_n3), .Z(
        u4_sll_479_ML_int_2__15_) );
  MUX2_X2 u4_sll_479_M1_1_16 ( .A(u4_sll_479_ML_int_1__16_), .B(
        u4_sll_479_ML_int_1__14_), .S(u4_sll_479_n3), .Z(
        u4_sll_479_ML_int_2__16_) );
  MUX2_X2 u4_sll_479_M1_1_17 ( .A(u4_sll_479_ML_int_1__17_), .B(
        u4_sll_479_ML_int_1__15_), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_2__17_) );
  MUX2_X2 u4_sll_479_M1_1_18 ( .A(u4_sll_479_ML_int_1__18_), .B(
        u4_sll_479_ML_int_1__16_), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_2__18_) );
  MUX2_X2 u4_sll_479_M1_1_19 ( .A(u4_sll_479_ML_int_1__19_), .B(
        u4_sll_479_ML_int_1__17_), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_2__19_) );
  MUX2_X2 u4_sll_479_M1_1_20 ( .A(u4_sll_479_ML_int_1__20_), .B(
        u4_sll_479_ML_int_1__18_), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_2__20_) );
  MUX2_X2 u4_sll_479_M1_1_21 ( .A(u4_sll_479_ML_int_1__21_), .B(
        u4_sll_479_ML_int_1__19_), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_2__21_) );
  MUX2_X2 u4_sll_479_M1_1_22 ( .A(u4_sll_479_ML_int_1__22_), .B(
        u4_sll_479_ML_int_1__20_), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_2__22_) );
  MUX2_X2 u4_sll_479_M1_1_23 ( .A(u4_sll_479_ML_int_1__23_), .B(
        u4_sll_479_ML_int_1__21_), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_2__23_) );
  MUX2_X2 u4_sll_479_M1_1_24 ( .A(u4_sll_479_ML_int_1__24_), .B(
        u4_sll_479_ML_int_1__22_), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_2__24_) );
  MUX2_X2 u4_sll_479_M1_1_25 ( .A(u4_sll_479_ML_int_1__25_), .B(
        u4_sll_479_ML_int_1__23_), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_2__25_) );
  MUX2_X2 u4_sll_479_M1_1_26 ( .A(u4_sll_479_ML_int_1__26_), .B(
        u4_sll_479_ML_int_1__24_), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_2__26_) );
  MUX2_X2 u4_sll_479_M1_1_27 ( .A(u4_sll_479_ML_int_1__27_), .B(
        u4_sll_479_ML_int_1__25_), .S(u4_sll_479_n2), .Z(
        u4_sll_479_ML_int_2__27_) );
  MUX2_X2 u4_sll_479_M1_2_7 ( .A(u4_sll_479_ML_int_2__7_), .B(
        u4_sll_479_ML_int_2__3_), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_3__7_) );
  MUX2_X2 u4_sll_479_M1_2_8 ( .A(u4_sll_479_ML_int_2__8_), .B(
        u4_sll_479_ML_int_2__4_), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_3__8_) );
  MUX2_X2 u4_sll_479_M1_2_9 ( .A(u4_sll_479_ML_int_2__9_), .B(
        u4_sll_479_ML_int_2__5_), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_3__9_) );
  MUX2_X2 u4_sll_479_M1_2_10 ( .A(u4_sll_479_ML_int_2__10_), .B(
        u4_sll_479_ML_int_2__6_), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_3__10_) );
  MUX2_X2 u4_sll_479_M1_2_11 ( .A(u4_sll_479_ML_int_2__11_), .B(
        u4_sll_479_ML_int_2__7_), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_3__11_) );
  MUX2_X2 u4_sll_479_M1_2_15 ( .A(u4_sll_479_ML_int_2__15_), .B(
        u4_sll_479_ML_int_2__11_), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_3__15_) );
  MUX2_X2 u4_sll_479_M1_2_16 ( .A(u4_sll_479_ML_int_2__16_), .B(
        u4_sll_479_ML_int_2__12_), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_3__16_) );
  MUX2_X2 u4_sll_479_M1_2_17 ( .A(u4_sll_479_ML_int_2__17_), .B(
        u4_sll_479_ML_int_2__13_), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_3__17_) );
  MUX2_X2 u4_sll_479_M1_2_18 ( .A(u4_sll_479_ML_int_2__18_), .B(
        u4_sll_479_ML_int_2__14_), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_3__18_) );
  MUX2_X2 u4_sll_479_M1_2_19 ( .A(u4_sll_479_ML_int_2__19_), .B(
        u4_sll_479_ML_int_2__15_), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_3__19_) );
  MUX2_X2 u4_sll_479_M1_2_23 ( .A(u4_sll_479_ML_int_2__23_), .B(
        u4_sll_479_ML_int_2__19_), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_3__23_) );
  MUX2_X2 u4_sll_479_M1_2_24 ( .A(u4_sll_479_ML_int_2__24_), .B(
        u4_sll_479_ML_int_2__20_), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_3__24_) );
  MUX2_X2 u4_sll_479_M1_2_25 ( .A(u4_sll_479_ML_int_2__25_), .B(
        u4_sll_479_ML_int_2__21_), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_3__25_) );
  MUX2_X2 u4_sll_479_M1_2_26 ( .A(u4_sll_479_ML_int_2__26_), .B(
        u4_sll_479_ML_int_2__22_), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_3__26_) );
  MUX2_X2 u4_sll_479_M1_2_27 ( .A(u4_sll_479_ML_int_2__27_), .B(
        u4_sll_479_ML_int_2__23_), .S(u4_sll_479_n1), .Z(
        u4_sll_479_ML_int_3__27_) );
  MUX2_X2 u4_sll_479_M1_3_8 ( .A(u4_sll_479_ML_int_3__8_), .B(
        u4_sll_479_ML_int_3__0_), .S(u4_f2i_shft_3_), .Z(
        u4_sll_479_ML_int_4__8_) );
  MUX2_X2 u4_sll_479_M1_3_9 ( .A(u4_sll_479_ML_int_3__9_), .B(
        u4_sll_479_ML_int_3__1_), .S(u4_f2i_shft_3_), .Z(
        u4_sll_479_ML_int_4__9_) );
  MUX2_X2 u4_sll_479_M1_3_10 ( .A(u4_sll_479_ML_int_3__10_), .B(
        u4_sll_479_ML_int_3__2_), .S(u4_f2i_shft_3_), .Z(
        u4_sll_479_ML_int_4__10_) );
  MUX2_X2 u4_sll_479_M1_3_11 ( .A(u4_sll_479_ML_int_3__11_), .B(
        u4_sll_479_ML_int_3__3_), .S(u4_f2i_shft_3_), .Z(
        u4_sll_479_ML_int_4__11_) );
  MUX2_X2 u4_sll_479_M1_3_23 ( .A(u4_sll_479_ML_int_3__23_), .B(
        u4_sll_479_ML_int_3__15_), .S(u4_f2i_shft_3_), .Z(
        u4_sll_479_ML_int_4__23_) );
  MUX2_X2 u4_sll_479_M1_3_24 ( .A(u4_sll_479_ML_int_3__24_), .B(
        u4_sll_479_ML_int_3__16_), .S(u4_f2i_shft_3_), .Z(
        u4_sll_479_ML_int_4__24_) );
  MUX2_X2 u4_sll_479_M1_3_25 ( .A(u4_sll_479_ML_int_3__25_), .B(
        u4_sll_479_ML_int_3__17_), .S(u4_f2i_shft_3_), .Z(
        u4_sll_479_ML_int_4__25_) );
  MUX2_X2 u4_sll_479_M1_3_26 ( .A(u4_sll_479_ML_int_3__26_), .B(
        u4_sll_479_ML_int_3__18_), .S(u4_f2i_shft_3_), .Z(
        u4_sll_479_ML_int_4__26_) );
  MUX2_X2 u4_sll_479_M1_3_27 ( .A(u4_sll_479_ML_int_3__27_), .B(
        u4_sll_479_ML_int_3__19_), .S(u4_f2i_shft_3_), .Z(
        u4_sll_479_ML_int_4__27_) );
  MUX2_X2 u4_sll_479_M1_4_23 ( .A(u4_sll_479_ML_int_4__23_), .B(
        u4_sll_479_ML_int_4__7_), .S(u4_f2i_shft_4_), .Z(u4_exp_f2i_1[23]) );
  MUX2_X2 u4_sll_479_M1_4_24 ( .A(u4_sll_479_ML_int_4__24_), .B(
        u4_sll_479_ML_int_4__8_), .S(u4_f2i_shft_4_), .Z(u4_exp_f2i_1[24]) );
  MUX2_X2 u4_sll_479_M1_4_25 ( .A(u4_sll_479_ML_int_4__25_), .B(
        u4_sll_479_ML_int_4__9_), .S(u4_f2i_shft_4_), .Z(u4_exp_f2i_1[25]) );
  MUX2_X2 u4_sll_479_M1_4_26 ( .A(u4_sll_479_ML_int_4__26_), .B(
        u4_sll_479_ML_int_4__10_), .S(u4_f2i_shft_4_), .Z(u4_exp_f2i_1[26]) );
  MUX2_X2 u4_sll_479_M1_4_27 ( .A(u4_sll_479_ML_int_4__27_), .B(
        u4_sll_479_ML_int_4__11_), .S(u4_f2i_shft_4_), .Z(u4_exp_f2i_1[27]) );
  INV_X4 u4_sub_467_U9 ( .A(n1667), .ZN(u4_sub_467_n7) );
  INV_X4 u4_sub_467_U8 ( .A(u4_fi_ldz_mi1_4_), .ZN(u4_sub_467_n6) );
  INV_X4 u4_sub_467_U7 ( .A(u4_fi_ldz_mi1_6_), .ZN(u4_sub_467_n5) );
  INV_X4 u4_sub_467_U6 ( .A(u4_fi_ldz_mi1_3_), .ZN(u4_sub_467_n4) );
  INV_X4 u4_sub_467_U5 ( .A(u4_fi_ldz_mi1_2_), .ZN(u4_sub_467_n3) );
  INV_X4 u4_sub_467_U4 ( .A(u4_fi_ldz_mi1_1_), .ZN(u4_sub_467_n2) );
  INV_X4 u4_sub_467_U3 ( .A(u4_exp_in_pl1_0_), .ZN(u4_sub_467_n1) );
  XNOR2_X2 u4_sub_467_U2 ( .A(u4_sub_467_n7), .B(u4_exp_in_pl1_0_), .ZN(
        u4_exp_next_mi_0_) );
  NAND2_X2 u4_sub_467_U1 ( .A1(n1667), .A2(u4_sub_467_n1), .ZN(
        u4_sub_467_carry[1]) );
  FA_X1 u4_sub_467_U2_1 ( .A(u4_exp_in_pl1_1_), .B(u4_sub_467_n2), .CI(
        u4_sub_467_carry[1]), .CO(u4_sub_467_carry[2]), .S(u4_exp_next_mi_1_)
         );
  FA_X1 u4_sub_467_U2_2 ( .A(u4_exp_in_pl1_2_), .B(u4_sub_467_n3), .CI(
        u4_sub_467_carry[2]), .CO(u4_sub_467_carry[3]), .S(u4_exp_next_mi_2_)
         );
  FA_X1 u4_sub_467_U2_3 ( .A(u4_exp_in_pl1_3_), .B(u4_sub_467_n4), .CI(
        u4_sub_467_carry[3]), .CO(u4_sub_467_carry[4]), .S(u4_exp_next_mi_3_)
         );
  FA_X1 u4_sub_467_U2_4 ( .A(u4_exp_in_pl1_4_), .B(u4_sub_467_n6), .CI(
        u4_sub_467_carry[4]), .CO(u4_sub_467_carry[5]), .S(u4_exp_next_mi_4_)
         );
  FA_X1 u4_sub_467_U2_5 ( .A(u4_exp_in_pl1_5_), .B(u4_sub_467_n5), .CI(
        u4_sub_467_carry[5]), .S(u4_exp_next_mi_5_) );
  INV_X4 u3_sub_59_U18 ( .A(fractb[13]), .ZN(u3_sub_59_n16) );
  INV_X4 u3_sub_59_U17 ( .A(fractb[12]), .ZN(u3_sub_59_n15) );
  INV_X4 u3_sub_59_U16 ( .A(fractb[11]), .ZN(u3_sub_59_n14) );
  INV_X4 u3_sub_59_U15 ( .A(fractb[10]), .ZN(u3_sub_59_n13) );
  INV_X4 u3_sub_59_U14 ( .A(fractb[9]), .ZN(u3_sub_59_n12) );
  INV_X4 u3_sub_59_U13 ( .A(fractb[8]), .ZN(u3_sub_59_n11) );
  INV_X4 u3_sub_59_U12 ( .A(fractb[7]), .ZN(u3_sub_59_n10) );
  INV_X4 u3_sub_59_U11 ( .A(fractb[6]), .ZN(u3_sub_59_n9) );
  INV_X4 u3_sub_59_U10 ( .A(fractb[5]), .ZN(u3_sub_59_n8) );
  INV_X4 u3_sub_59_U9 ( .A(fractb[4]), .ZN(u3_sub_59_n7) );
  INV_X4 u3_sub_59_U8 ( .A(fractb[3]), .ZN(u3_sub_59_n6) );
  INV_X4 u3_sub_59_U7 ( .A(fractb[2]), .ZN(u3_sub_59_n5) );
  INV_X4 u3_sub_59_U6 ( .A(fractb[1]), .ZN(u3_sub_59_n4) );
  INV_X4 u3_sub_59_U5 ( .A(fractb[0]), .ZN(u3_sub_59_n3) );
  INV_X4 u3_sub_59_U4 ( .A(u3_sub_59_carry[14]), .ZN(u3_N32) );
  INV_X4 u3_sub_59_U3 ( .A(fracta[0]), .ZN(u3_sub_59_n1) );
  XNOR2_X2 u3_sub_59_U2 ( .A(u3_sub_59_n3), .B(fracta[0]), .ZN(u3_N18) );
  NAND2_X2 u3_sub_59_U1 ( .A1(fractb[0]), .A2(u3_sub_59_n1), .ZN(
        u3_sub_59_carry[1]) );
  FA_X1 u3_sub_59_U2_1 ( .A(fracta[1]), .B(u3_sub_59_n4), .CI(
        u3_sub_59_carry[1]), .CO(u3_sub_59_carry[2]), .S(u3_N19) );
  FA_X1 u3_sub_59_U2_2 ( .A(fracta[2]), .B(u3_sub_59_n5), .CI(
        u3_sub_59_carry[2]), .CO(u3_sub_59_carry[3]), .S(u3_N20) );
  FA_X1 u3_sub_59_U2_3 ( .A(fracta[3]), .B(u3_sub_59_n6), .CI(
        u3_sub_59_carry[3]), .CO(u3_sub_59_carry[4]), .S(u3_N21) );
  FA_X1 u3_sub_59_U2_4 ( .A(fracta[4]), .B(u3_sub_59_n7), .CI(
        u3_sub_59_carry[4]), .CO(u3_sub_59_carry[5]), .S(u3_N22) );
  FA_X1 u3_sub_59_U2_5 ( .A(fracta[5]), .B(u3_sub_59_n8), .CI(
        u3_sub_59_carry[5]), .CO(u3_sub_59_carry[6]), .S(u3_N23) );
  FA_X1 u3_sub_59_U2_6 ( .A(fracta[6]), .B(u3_sub_59_n9), .CI(
        u3_sub_59_carry[6]), .CO(u3_sub_59_carry[7]), .S(u3_N24) );
  FA_X1 u3_sub_59_U2_7 ( .A(fracta[7]), .B(u3_sub_59_n10), .CI(
        u3_sub_59_carry[7]), .CO(u3_sub_59_carry[8]), .S(u3_N25) );
  FA_X1 u3_sub_59_U2_8 ( .A(fracta[8]), .B(u3_sub_59_n11), .CI(
        u3_sub_59_carry[8]), .CO(u3_sub_59_carry[9]), .S(u3_N26) );
  FA_X1 u3_sub_59_U2_9 ( .A(fracta[9]), .B(u3_sub_59_n12), .CI(
        u3_sub_59_carry[9]), .CO(u3_sub_59_carry[10]), .S(u3_N27) );
  FA_X1 u3_sub_59_U2_10 ( .A(fracta[10]), .B(u3_sub_59_n13), .CI(
        u3_sub_59_carry[10]), .CO(u3_sub_59_carry[11]), .S(u3_N28) );
  FA_X1 u3_sub_59_U2_11 ( .A(fracta[11]), .B(u3_sub_59_n14), .CI(
        u3_sub_59_carry[11]), .CO(u3_sub_59_carry[12]), .S(u3_N29) );
  FA_X1 u3_sub_59_U2_12 ( .A(fracta[12]), .B(u3_sub_59_n15), .CI(
        u3_sub_59_carry[12]), .CO(u3_sub_59_carry[13]), .S(u3_N30) );
  FA_X1 u3_sub_59_U2_13 ( .A(fracta[13]), .B(u3_sub_59_n16), .CI(
        u3_sub_59_carry[13]), .CO(u3_sub_59_carry[14]), .S(u3_N31) );
  XOR2_X2 u3_add_59_U2 ( .A(fractb[0]), .B(fracta[0]), .Z(u3_N3) );
  AND2_X4 u3_add_59_U1 ( .A1(fractb[0]), .A2(fracta[0]), .ZN(u3_add_59_n1) );
  FA_X1 u3_add_59_U1_1 ( .A(fracta[1]), .B(fractb[1]), .CI(u3_add_59_n1), .CO(
        u3_add_59_carry[2]), .S(u3_N4) );
  FA_X1 u3_add_59_U1_2 ( .A(fracta[2]), .B(fractb[2]), .CI(u3_add_59_carry[2]), 
        .CO(u3_add_59_carry[3]), .S(u3_N5) );
  FA_X1 u3_add_59_U1_3 ( .A(fracta[3]), .B(fractb[3]), .CI(u3_add_59_carry[3]), 
        .CO(u3_add_59_carry[4]), .S(u3_N6) );
  FA_X1 u3_add_59_U1_4 ( .A(fracta[4]), .B(fractb[4]), .CI(u3_add_59_carry[4]), 
        .CO(u3_add_59_carry[5]), .S(u3_N7) );
  FA_X1 u3_add_59_U1_5 ( .A(fracta[5]), .B(fractb[5]), .CI(u3_add_59_carry[5]), 
        .CO(u3_add_59_carry[6]), .S(u3_N8) );
  FA_X1 u3_add_59_U1_6 ( .A(fracta[6]), .B(fractb[6]), .CI(u3_add_59_carry[6]), 
        .CO(u3_add_59_carry[7]), .S(u3_N9) );
  FA_X1 u3_add_59_U1_7 ( .A(fracta[7]), .B(fractb[7]), .CI(u3_add_59_carry[7]), 
        .CO(u3_add_59_carry[8]), .S(u3_N10) );
  FA_X1 u3_add_59_U1_8 ( .A(fracta[8]), .B(fractb[8]), .CI(u3_add_59_carry[8]), 
        .CO(u3_add_59_carry[9]), .S(u3_N11) );
  FA_X1 u3_add_59_U1_9 ( .A(fracta[9]), .B(fractb[9]), .CI(u3_add_59_carry[9]), 
        .CO(u3_add_59_carry[10]), .S(u3_N12) );
  FA_X1 u3_add_59_U1_10 ( .A(fracta[10]), .B(fractb[10]), .CI(
        u3_add_59_carry[10]), .CO(u3_add_59_carry[11]), .S(u3_N13) );
  FA_X1 u3_add_59_U1_11 ( .A(fracta[11]), .B(fractb[11]), .CI(
        u3_add_59_carry[11]), .CO(u3_add_59_carry[12]), .S(u3_N14) );
  FA_X1 u3_add_59_U1_12 ( .A(fracta[12]), .B(fractb[12]), .CI(
        u3_add_59_carry[12]), .CO(u3_add_59_carry[13]), .S(u3_N15) );
  FA_X1 u3_add_59_U1_13 ( .A(fracta[13]), .B(fractb[13]), .CI(
        u3_add_59_carry[13]), .CO(u3_N17), .S(u3_N16) );
  NAND2_X1 u1_srl_146_U63 ( .A1(n2687), .A2(u1_srl_146_n13), .ZN(
        u1_srl_146_n27) );
  NAND2_X1 u1_srl_146_U62 ( .A1(u1_exp_diff_sft_0_), .A2(n2685), .ZN(
        u1_srl_146_n45) );
  AOI22_X1 u1_srl_146_U61 ( .A1(n2689), .A2(u1_srl_146_n34), .B1(u1_srl_146_n9), .B2(n2688), .ZN(u1_srl_146_n47) );
  AOI221_X1 u1_srl_146_U60 ( .B1(u1_srl_146_n31), .B2(n2690), .C1(
        u1_srl_146_n32), .C2(n2691), .A(u1_srl_146_n1), .ZN(u1_srl_146_n17) );
  AOI22_X1 u1_srl_146_U59 ( .A1(n2693), .A2(u1_srl_146_n34), .B1(n2692), .B2(
        u1_srl_146_n9), .ZN(u1_srl_146_n46) );
  AOI221_X1 u1_srl_146_U58 ( .B1(u1_srl_146_n31), .B2(n2694), .C1(
        u1_srl_146_n32), .C2(n2695), .A(u1_srl_146_n2), .ZN(u1_srl_146_n29) );
  AOI22_X1 u1_srl_146_U57 ( .A1(u1_adj_op_9_), .A2(u1_srl_146_n32), .B1(
        u1_srl_146_n31), .B2(n1521), .ZN(u1_srl_146_n19) );
  OAI33_X1 u1_srl_146_U56 ( .A1(u1_srl_146_n14), .A2(u1_srl_146_n19), .A3(
        u1_srl_146_n13), .B1(u1_srl_146_n15), .B2(u1_srl_146_n45), .B3(
        u1_srl_146_n18), .ZN(u1_srl_146_n44) );
  OAI221_X1 u1_srl_146_U55 ( .B1(u1_srl_146_n27), .B2(u1_srl_146_n17), .C1(
        u1_srl_146_n20), .C2(u1_srl_146_n29), .A(u1_srl_146_n10), .ZN(
        u1_adj_op_out_sft_0_) );
  AOI22_X1 u1_srl_146_U54 ( .A1(u1_adj_op_9_), .A2(u1_srl_146_n34), .B1(n1521), 
        .B2(u1_srl_146_n9), .ZN(u1_srl_146_n43) );
  AOI221_X1 u1_srl_146_U53 ( .B1(n2688), .B2(u1_srl_146_n31), .C1(n2689), .C2(
        u1_srl_146_n32), .A(u1_srl_146_n3), .ZN(u1_srl_146_n24) );
  NOR2_X1 u1_srl_146_U52 ( .A1(u1_srl_146_n24), .A2(u1_srl_146_n18), .ZN(
        u1_adj_op_out_sft_10_) );
  AOI222_X1 u1_srl_146_U51 ( .A1(u1_adj_op_9_), .A2(u1_srl_146_n31), .B1(
        u1_srl_146_n34), .B2(n1521), .C1(n2688), .C2(u1_srl_146_n32), .ZN(
        u1_srl_146_n22) );
  NOR2_X1 u1_srl_146_U50 ( .A1(u1_srl_146_n22), .A2(u1_srl_146_n18), .ZN(
        u1_adj_op_out_sft_11_) );
  NOR2_X1 u1_srl_146_U49 ( .A1(u1_srl_146_n19), .A2(u1_srl_146_n18), .ZN(
        u1_adj_op_out_sft_12_) );
  NAND2_X1 u1_srl_146_U48 ( .A1(n1521), .A2(u1_srl_146_n32), .ZN(
        u1_srl_146_n26) );
  NOR2_X1 u1_srl_146_U47 ( .A1(u1_srl_146_n26), .A2(u1_srl_146_n18), .ZN(
        u1_adj_op_out_sft_13_) );
  AOI22_X1 u1_srl_146_U46 ( .A1(n2692), .A2(u1_srl_146_n34), .B1(n2691), .B2(
        u1_srl_146_n9), .ZN(u1_srl_146_n42) );
  AOI221_X1 u1_srl_146_U45 ( .B1(u1_srl_146_n31), .B2(n2693), .C1(
        u1_srl_146_n32), .C2(n2694), .A(u1_srl_146_n4), .ZN(u1_srl_146_n28) );
  AOI22_X1 u1_srl_146_U44 ( .A1(n2688), .A2(u1_srl_146_n34), .B1(u1_adj_op_9_), 
        .B2(u1_srl_146_n9), .ZN(u1_srl_146_n41) );
  AOI221_X1 u1_srl_146_U43 ( .B1(u1_srl_146_n31), .B2(n2689), .C1(
        u1_srl_146_n32), .C2(n2690), .A(u1_srl_146_n5), .ZN(u1_srl_146_n25) );
  MUX2_X1 u1_srl_146_U42 ( .A(u1_srl_146_n25), .B(u1_srl_146_n26), .S(n2686), 
        .Z(u1_srl_146_n16) );
  MUX2_X1 u1_srl_146_U41 ( .A(n2696), .B(n2695), .S(u1_exp_diff_sft_0_), .Z(
        u1_srl_146_n40) );
  NAND3_X1 u1_srl_146_U40 ( .A1(u1_srl_146_n12), .A2(n2685), .A3(
        u1_srl_146_n40), .ZN(u1_srl_146_n39) );
  OAI221_X1 u1_srl_146_U39 ( .B1(u1_srl_146_n28), .B2(u1_srl_146_n20), .C1(
        u1_srl_146_n16), .C2(u1_srl_146_n14), .A(u1_srl_146_n39), .ZN(
        u1_adj_op_out_sft_1_) );
  MUX2_X1 u1_srl_146_U38 ( .A(n2695), .B(n2694), .S(u1_exp_diff_sft_0_), .Z(
        u1_srl_146_n38) );
  AOI22_X1 u1_srl_146_U37 ( .A1(n2696), .A2(u1_srl_146_n31), .B1(
        u1_srl_146_n38), .B2(n2685), .ZN(u1_srl_146_n36) );
  AOI22_X1 u1_srl_146_U36 ( .A1(n2691), .A2(u1_srl_146_n34), .B1(n2690), .B2(
        u1_srl_146_n9), .ZN(u1_srl_146_n37) );
  AOI221_X1 u1_srl_146_U35 ( .B1(u1_srl_146_n31), .B2(n2692), .C1(
        u1_srl_146_n32), .C2(n2693), .A(u1_srl_146_n6), .ZN(u1_srl_146_n23) );
  OAI222_X1 u1_srl_146_U34 ( .A1(u1_srl_146_n24), .A2(u1_srl_146_n27), .B1(
        u1_srl_146_n36), .B2(u1_srl_146_n18), .C1(u1_srl_146_n23), .C2(
        u1_srl_146_n20), .ZN(u1_adj_op_out_sft_2_) );
  AOI22_X1 u1_srl_146_U33 ( .A1(n2690), .A2(u1_srl_146_n34), .B1(n2689), .B2(
        u1_srl_146_n9), .ZN(u1_srl_146_n35) );
  AOI221_X1 u1_srl_146_U32 ( .B1(u1_srl_146_n31), .B2(n2691), .C1(
        u1_srl_146_n32), .C2(n2692), .A(u1_srl_146_n7), .ZN(u1_srl_146_n21) );
  AOI22_X1 u1_srl_146_U31 ( .A1(u1_srl_146_n9), .A2(n2693), .B1(u1_srl_146_n34), .B2(n2694), .ZN(u1_srl_146_n33) );
  AOI221_X1 u1_srl_146_U30 ( .B1(n2695), .B2(u1_srl_146_n31), .C1(n2696), .C2(
        u1_srl_146_n32), .A(u1_srl_146_n8), .ZN(u1_srl_146_n30) );
  OAI222_X1 u1_srl_146_U29 ( .A1(u1_srl_146_n21), .A2(u1_srl_146_n20), .B1(
        u1_srl_146_n22), .B2(u1_srl_146_n27), .C1(u1_srl_146_n30), .C2(
        u1_srl_146_n18), .ZN(u1_adj_op_out_sft_3_) );
  OAI222_X1 u1_srl_146_U28 ( .A1(u1_srl_146_n17), .A2(u1_srl_146_n20), .B1(
        u1_srl_146_n19), .B2(u1_srl_146_n27), .C1(u1_srl_146_n29), .C2(
        u1_srl_146_n18), .ZN(u1_adj_op_out_sft_4_) );
  OAI222_X1 u1_srl_146_U27 ( .A1(u1_srl_146_n25), .A2(u1_srl_146_n20), .B1(
        u1_srl_146_n26), .B2(u1_srl_146_n27), .C1(u1_srl_146_n28), .C2(
        u1_srl_146_n18), .ZN(u1_adj_op_out_sft_5_) );
  OAI22_X1 u1_srl_146_U26 ( .A1(u1_srl_146_n23), .A2(u1_srl_146_n18), .B1(
        u1_srl_146_n24), .B2(u1_srl_146_n20), .ZN(u1_adj_op_out_sft_6_) );
  OAI22_X1 u1_srl_146_U25 ( .A1(u1_srl_146_n21), .A2(u1_srl_146_n18), .B1(
        u1_srl_146_n22), .B2(u1_srl_146_n20), .ZN(u1_adj_op_out_sft_7_) );
  OAI22_X1 u1_srl_146_U24 ( .A1(u1_srl_146_n17), .A2(u1_srl_146_n18), .B1(
        u1_srl_146_n19), .B2(u1_srl_146_n20), .ZN(u1_adj_op_out_sft_8_) );
  NOR2_X1 u1_srl_146_U23 ( .A1(n2687), .A2(u1_srl_146_n16), .ZN(
        u1_adj_op_out_sft_9_) );
  INV_X4 u1_srl_146_U22 ( .A(n2696), .ZN(u1_srl_146_n15) );
  INV_X4 u1_srl_146_U21 ( .A(n2687), .ZN(u1_srl_146_n14) );
  INV_X4 u1_srl_146_U20 ( .A(n2686), .ZN(u1_srl_146_n13) );
  INV_X4 u1_srl_146_U19 ( .A(u1_srl_146_n18), .ZN(u1_srl_146_n12) );
  INV_X4 u1_srl_146_U18 ( .A(u1_exp_diff_sft_0_), .ZN(u1_srl_146_n11) );
  INV_X4 u1_srl_146_U17 ( .A(u1_srl_146_n44), .ZN(u1_srl_146_n10) );
  INV_X4 u1_srl_146_U16 ( .A(u1_srl_146_n45), .ZN(u1_srl_146_n9) );
  INV_X4 u1_srl_146_U15 ( .A(u1_srl_146_n33), .ZN(u1_srl_146_n8) );
  INV_X4 u1_srl_146_U14 ( .A(u1_srl_146_n35), .ZN(u1_srl_146_n7) );
  INV_X4 u1_srl_146_U13 ( .A(u1_srl_146_n37), .ZN(u1_srl_146_n6) );
  INV_X4 u1_srl_146_U12 ( .A(u1_srl_146_n41), .ZN(u1_srl_146_n5) );
  INV_X4 u1_srl_146_U11 ( .A(u1_srl_146_n42), .ZN(u1_srl_146_n4) );
  INV_X4 u1_srl_146_U10 ( .A(u1_srl_146_n43), .ZN(u1_srl_146_n3) );
  INV_X4 u1_srl_146_U9 ( .A(u1_srl_146_n46), .ZN(u1_srl_146_n2) );
  INV_X4 u1_srl_146_U8 ( .A(u1_srl_146_n47), .ZN(u1_srl_146_n1) );
  AND2_X4 u1_srl_146_U7 ( .A1(n2685), .A2(u1_srl_146_n11), .ZN(u1_srl_146_n34)
         );
  NAND2_X2 u1_srl_146_U6 ( .A1(n2686), .A2(u1_srl_146_n14), .ZN(u1_srl_146_n20) );
  NAND2_X2 u1_srl_146_U5 ( .A1(u1_srl_146_n13), .A2(u1_srl_146_n14), .ZN(
        u1_srl_146_n18) );
  NOR2_X2 u1_srl_146_U4 ( .A1(u1_srl_146_n11), .A2(n2685), .ZN(u1_srl_146_n31)
         );
  NOR2_X2 u1_srl_146_U3 ( .A1(u1_exp_diff_sft_0_), .A2(n2685), .ZN(
        u1_srl_146_n32) );
  AND2_X1 sll_384_U25 ( .A1(fracta_mul[0]), .A2(sll_384_n3), .ZN(
        sll_384_ML_int_1__0_) );
  NAND2_X1 sll_384_U24 ( .A1(sll_384_ML_int_1__0_), .A2(sll_384_n8), .ZN(
        sll_384_n11) );
  NAND2_X1 sll_384_U23 ( .A1(sll_384_ML_int_1__1_), .A2(sll_384_n8), .ZN(
        sll_384_n10) );
  NOR2_X1 sll_384_U22 ( .A1(N44), .A2(sll_384_n11), .ZN(sll_384_ML_int_3__0_)
         );
  NOR2_X1 sll_384_U21 ( .A1(N44), .A2(sll_384_n10), .ZN(sll_384_ML_int_3__1_)
         );
  NOR2_X1 sll_384_U20 ( .A1(N44), .A2(sll_384_n2), .ZN(sll_384_ML_int_3__2_)
         );
  NAND2_X1 sll_384_U19 ( .A1(sll_384_n7), .A2(sll_384_n6), .ZN(sll_384_n9) );
  NOR2_X1 sll_384_U18 ( .A1(sll_384_n9), .A2(sll_384_n11), .ZN(N67) );
  NOR2_X1 sll_384_U17 ( .A1(sll_384_n9), .A2(sll_384_n10), .ZN(N68) );
  NOR2_X1 sll_384_U16 ( .A1(sll_384_n9), .A2(sll_384_n2), .ZN(N69) );
  NOR2_X1 sll_384_U15 ( .A1(sll_384_n5), .A2(sll_384_n9), .ZN(N70) );
  AND2_X1 sll_384_U14 ( .A1(sll_384_ML_int_3__4_), .A2(sll_384_n6), .ZN(N71)
         );
  AND2_X1 sll_384_U13 ( .A1(sll_384_ML_int_3__5_), .A2(sll_384_n6), .ZN(N72)
         );
  AND2_X1 sll_384_U12 ( .A1(sll_384_ML_int_3__6_), .A2(sll_384_n6), .ZN(N73)
         );
  AND2_X1 sll_384_U11 ( .A1(sll_384_ML_int_3__7_), .A2(sll_384_n6), .ZN(N74)
         );
  INV_X4 sll_384_U10 ( .A(N56), .ZN(sll_384_n8) );
  INV_X4 sll_384_U9 ( .A(N44), .ZN(sll_384_n7) );
  INV_X4 sll_384_U8 ( .A(N34), .ZN(sll_384_n6) );
  INV_X4 sll_384_U7 ( .A(sll_384_ML_int_2__3_), .ZN(sll_384_n5) );
  INV_X4 sll_384_U6 ( .A(sll_384_n10), .ZN(sll_384_n4) );
  INV_X4 sll_384_U5 ( .A(N65), .ZN(sll_384_n3) );
  INV_X4 sll_384_U4 ( .A(sll_384_ML_int_2__2_), .ZN(sll_384_n2) );
  INV_X4 sll_384_U3 ( .A(sll_384_n11), .ZN(sll_384_n1) );
  MUX2_X2 sll_384_M1_0_1 ( .A(fracta_mul[1]), .B(fracta_mul[0]), .S(N65), .Z(
        sll_384_ML_int_1__1_) );
  MUX2_X2 sll_384_M1_0_2 ( .A(fracta_mul[2]), .B(fracta_mul[1]), .S(N65), .Z(
        sll_384_ML_int_1__2_) );
  MUX2_X2 sll_384_M1_0_3 ( .A(fracta_mul[3]), .B(fracta_mul[2]), .S(N65), .Z(
        sll_384_ML_int_1__3_) );
  MUX2_X2 sll_384_M1_0_4 ( .A(fracta_mul[4]), .B(fracta_mul[3]), .S(N65), .Z(
        sll_384_ML_int_1__4_) );
  MUX2_X2 sll_384_M1_0_5 ( .A(fracta_mul[5]), .B(fracta_mul[4]), .S(N65), .Z(
        sll_384_ML_int_1__5_) );
  MUX2_X2 sll_384_M1_0_6 ( .A(fracta_mul[6]), .B(fracta_mul[5]), .S(N65), .Z(
        sll_384_ML_int_1__6_) );
  MUX2_X2 sll_384_M1_0_7 ( .A(fracta_mul[7]), .B(fracta_mul[6]), .S(N65), .Z(
        sll_384_ML_int_1__7_) );
  MUX2_X2 sll_384_M1_0_8 ( .A(fracta_mul[8]), .B(fracta_mul[7]), .S(N65), .Z(
        sll_384_ML_int_1__8_) );
  MUX2_X2 sll_384_M1_0_9 ( .A(fracta_mul[9]), .B(fracta_mul[8]), .S(N65), .Z(
        sll_384_ML_int_1__9_) );
  MUX2_X2 sll_384_M1_0_10 ( .A(n2698), .B(fracta_mul[9]), .S(N65), .Z(
        sll_384_ML_int_1__10_) );
  MUX2_X2 sll_384_M1_1_2 ( .A(sll_384_ML_int_1__2_), .B(sll_384_ML_int_1__0_), 
        .S(N56), .Z(sll_384_ML_int_2__2_) );
  MUX2_X2 sll_384_M1_1_3 ( .A(sll_384_ML_int_1__3_), .B(sll_384_ML_int_1__1_), 
        .S(N56), .Z(sll_384_ML_int_2__3_) );
  MUX2_X2 sll_384_M1_1_4 ( .A(sll_384_ML_int_1__4_), .B(sll_384_ML_int_1__2_), 
        .S(N56), .Z(sll_384_ML_int_2__4_) );
  MUX2_X2 sll_384_M1_1_5 ( .A(sll_384_ML_int_1__5_), .B(sll_384_ML_int_1__3_), 
        .S(N56), .Z(sll_384_ML_int_2__5_) );
  MUX2_X2 sll_384_M1_1_6 ( .A(sll_384_ML_int_1__6_), .B(sll_384_ML_int_1__4_), 
        .S(N56), .Z(sll_384_ML_int_2__6_) );
  MUX2_X2 sll_384_M1_1_7 ( .A(sll_384_ML_int_1__7_), .B(sll_384_ML_int_1__5_), 
        .S(N56), .Z(sll_384_ML_int_2__7_) );
  MUX2_X2 sll_384_M1_1_8 ( .A(sll_384_ML_int_1__8_), .B(sll_384_ML_int_1__6_), 
        .S(N56), .Z(sll_384_ML_int_2__8_) );
  MUX2_X2 sll_384_M1_1_9 ( .A(sll_384_ML_int_1__9_), .B(sll_384_ML_int_1__7_), 
        .S(N56), .Z(sll_384_ML_int_2__9_) );
  MUX2_X2 sll_384_M1_1_10 ( .A(sll_384_ML_int_1__10_), .B(sll_384_ML_int_1__8_), .S(N56), .Z(sll_384_ML_int_2__10_) );
  MUX2_X2 sll_384_M1_2_4 ( .A(sll_384_ML_int_2__4_), .B(sll_384_n1), .S(N44), 
        .Z(sll_384_ML_int_3__4_) );
  MUX2_X2 sll_384_M1_2_5 ( .A(sll_384_ML_int_2__5_), .B(sll_384_n4), .S(N44), 
        .Z(sll_384_ML_int_3__5_) );
  MUX2_X2 sll_384_M1_2_6 ( .A(sll_384_ML_int_2__6_), .B(sll_384_ML_int_2__2_), 
        .S(N44), .Z(sll_384_ML_int_3__6_) );
  MUX2_X2 sll_384_M1_2_7 ( .A(sll_384_ML_int_2__7_), .B(sll_384_ML_int_2__3_), 
        .S(N44), .Z(sll_384_ML_int_3__7_) );
  MUX2_X2 sll_384_M1_2_8 ( .A(sll_384_ML_int_2__8_), .B(sll_384_ML_int_2__4_), 
        .S(N44), .Z(sll_384_ML_int_3__8_) );
  MUX2_X2 sll_384_M1_2_9 ( .A(sll_384_ML_int_2__9_), .B(sll_384_ML_int_2__5_), 
        .S(N44), .Z(sll_384_ML_int_3__9_) );
  MUX2_X2 sll_384_M1_2_10 ( .A(sll_384_ML_int_2__10_), .B(sll_384_ML_int_2__6_), .S(N44), .Z(sll_384_ML_int_3__10_) );
  MUX2_X2 sll_384_M1_3_8 ( .A(sll_384_ML_int_3__8_), .B(sll_384_ML_int_3__0_), 
        .S(N34), .Z(N75) );
  MUX2_X2 sll_384_M1_3_9 ( .A(sll_384_ML_int_3__9_), .B(sll_384_ML_int_3__1_), 
        .S(N34), .Z(N76) );
  MUX2_X2 sll_384_M1_3_10 ( .A(sll_384_ML_int_3__10_), .B(sll_384_ML_int_3__2_), .S(N34), .Z(N77) );
  NOR2_X1 u5_mult_78_U185 ( .A1(u5_mult_78_n64), .A2(u5_mult_78_n53), .ZN(
        u5_N0) );
  NOR2_X1 u5_mult_78_U184 ( .A1(u5_mult_78_n54), .A2(u5_mult_78_n53), .ZN(
        u5_mult_78_ab_0__10_) );
  NOR2_X1 u5_mult_78_U183 ( .A1(u5_mult_78_n63), .A2(u5_mult_78_n53), .ZN(
        u5_mult_78_ab_0__1_) );
  NOR2_X1 u5_mult_78_U182 ( .A1(u5_mult_78_n62), .A2(u5_mult_78_n53), .ZN(
        u5_mult_78_ab_0__2_) );
  NOR2_X1 u5_mult_78_U181 ( .A1(u5_mult_78_n61), .A2(u5_mult_78_n53), .ZN(
        u5_mult_78_ab_0__3_) );
  NOR2_X1 u5_mult_78_U180 ( .A1(u5_mult_78_n60), .A2(u5_mult_78_n53), .ZN(
        u5_mult_78_ab_0__4_) );
  NOR2_X1 u5_mult_78_U179 ( .A1(u5_mult_78_n59), .A2(u5_mult_78_n53), .ZN(
        u5_mult_78_ab_0__5_) );
  NOR2_X1 u5_mult_78_U178 ( .A1(u5_mult_78_n58), .A2(u5_mult_78_n53), .ZN(
        u5_mult_78_ab_0__6_) );
  NOR2_X1 u5_mult_78_U177 ( .A1(u5_mult_78_n57), .A2(u5_mult_78_n53), .ZN(
        u5_mult_78_ab_0__7_) );
  NOR2_X1 u5_mult_78_U176 ( .A1(u5_mult_78_n56), .A2(u5_mult_78_n53), .ZN(
        u5_mult_78_ab_0__8_) );
  NOR2_X1 u5_mult_78_U175 ( .A1(u5_mult_78_n55), .A2(u5_mult_78_n53), .ZN(
        u5_mult_78_ab_0__9_) );
  NOR2_X1 u5_mult_78_U174 ( .A1(u5_mult_78_n64), .A2(u5_mult_78_n43), .ZN(
        u5_mult_78_ab_10__0_) );
  NOR2_X1 u5_mult_78_U173 ( .A1(u5_mult_78_n54), .A2(u5_mult_78_n43), .ZN(
        u5_mult_78_ab_10__10_) );
  NOR2_X1 u5_mult_78_U172 ( .A1(u5_mult_78_n63), .A2(u5_mult_78_n43), .ZN(
        u5_mult_78_ab_10__1_) );
  NOR2_X1 u5_mult_78_U171 ( .A1(u5_mult_78_n62), .A2(u5_mult_78_n43), .ZN(
        u5_mult_78_ab_10__2_) );
  NOR2_X1 u5_mult_78_U170 ( .A1(u5_mult_78_n61), .A2(u5_mult_78_n43), .ZN(
        u5_mult_78_ab_10__3_) );
  NOR2_X1 u5_mult_78_U169 ( .A1(u5_mult_78_n60), .A2(u5_mult_78_n43), .ZN(
        u5_mult_78_ab_10__4_) );
  NOR2_X1 u5_mult_78_U168 ( .A1(u5_mult_78_n59), .A2(u5_mult_78_n43), .ZN(
        u5_mult_78_ab_10__5_) );
  NOR2_X1 u5_mult_78_U167 ( .A1(u5_mult_78_n58), .A2(u5_mult_78_n43), .ZN(
        u5_mult_78_ab_10__6_) );
  NOR2_X1 u5_mult_78_U166 ( .A1(u5_mult_78_n57), .A2(u5_mult_78_n43), .ZN(
        u5_mult_78_ab_10__7_) );
  NOR2_X1 u5_mult_78_U165 ( .A1(u5_mult_78_n56), .A2(u5_mult_78_n43), .ZN(
        u5_mult_78_ab_10__8_) );
  NOR2_X1 u5_mult_78_U164 ( .A1(u5_mult_78_n55), .A2(u5_mult_78_n43), .ZN(
        u5_mult_78_ab_10__9_) );
  NOR2_X1 u5_mult_78_U163 ( .A1(u5_mult_78_n64), .A2(u5_mult_78_n52), .ZN(
        u5_mult_78_ab_1__0_) );
  NOR2_X1 u5_mult_78_U162 ( .A1(u5_mult_78_n54), .A2(u5_mult_78_n52), .ZN(
        u5_mult_78_ab_1__10_) );
  NOR2_X1 u5_mult_78_U161 ( .A1(u5_mult_78_n63), .A2(u5_mult_78_n52), .ZN(
        u5_mult_78_ab_1__1_) );
  NOR2_X1 u5_mult_78_U160 ( .A1(u5_mult_78_n62), .A2(u5_mult_78_n52), .ZN(
        u5_mult_78_ab_1__2_) );
  NOR2_X1 u5_mult_78_U159 ( .A1(u5_mult_78_n61), .A2(u5_mult_78_n52), .ZN(
        u5_mult_78_ab_1__3_) );
  NOR2_X1 u5_mult_78_U158 ( .A1(u5_mult_78_n60), .A2(u5_mult_78_n52), .ZN(
        u5_mult_78_ab_1__4_) );
  NOR2_X1 u5_mult_78_U157 ( .A1(u5_mult_78_n59), .A2(u5_mult_78_n52), .ZN(
        u5_mult_78_ab_1__5_) );
  NOR2_X1 u5_mult_78_U156 ( .A1(u5_mult_78_n58), .A2(u5_mult_78_n52), .ZN(
        u5_mult_78_ab_1__6_) );
  NOR2_X1 u5_mult_78_U155 ( .A1(u5_mult_78_n57), .A2(u5_mult_78_n52), .ZN(
        u5_mult_78_ab_1__7_) );
  NOR2_X1 u5_mult_78_U154 ( .A1(u5_mult_78_n56), .A2(u5_mult_78_n52), .ZN(
        u5_mult_78_ab_1__8_) );
  NOR2_X1 u5_mult_78_U153 ( .A1(u5_mult_78_n55), .A2(u5_mult_78_n52), .ZN(
        u5_mult_78_ab_1__9_) );
  NOR2_X1 u5_mult_78_U152 ( .A1(u5_mult_78_n64), .A2(u5_mult_78_n51), .ZN(
        u5_mult_78_ab_2__0_) );
  NOR2_X1 u5_mult_78_U151 ( .A1(u5_mult_78_n54), .A2(u5_mult_78_n51), .ZN(
        u5_mult_78_ab_2__10_) );
  NOR2_X1 u5_mult_78_U150 ( .A1(u5_mult_78_n63), .A2(u5_mult_78_n51), .ZN(
        u5_mult_78_ab_2__1_) );
  NOR2_X1 u5_mult_78_U149 ( .A1(u5_mult_78_n62), .A2(u5_mult_78_n51), .ZN(
        u5_mult_78_ab_2__2_) );
  NOR2_X1 u5_mult_78_U148 ( .A1(u5_mult_78_n61), .A2(u5_mult_78_n51), .ZN(
        u5_mult_78_ab_2__3_) );
  NOR2_X1 u5_mult_78_U147 ( .A1(u5_mult_78_n60), .A2(u5_mult_78_n51), .ZN(
        u5_mult_78_ab_2__4_) );
  NOR2_X1 u5_mult_78_U146 ( .A1(u5_mult_78_n59), .A2(u5_mult_78_n51), .ZN(
        u5_mult_78_ab_2__5_) );
  NOR2_X1 u5_mult_78_U145 ( .A1(u5_mult_78_n58), .A2(u5_mult_78_n51), .ZN(
        u5_mult_78_ab_2__6_) );
  NOR2_X1 u5_mult_78_U144 ( .A1(u5_mult_78_n57), .A2(u5_mult_78_n51), .ZN(
        u5_mult_78_ab_2__7_) );
  NOR2_X1 u5_mult_78_U143 ( .A1(u5_mult_78_n56), .A2(u5_mult_78_n51), .ZN(
        u5_mult_78_ab_2__8_) );
  NOR2_X1 u5_mult_78_U142 ( .A1(u5_mult_78_n55), .A2(u5_mult_78_n51), .ZN(
        u5_mult_78_ab_2__9_) );
  NOR2_X1 u5_mult_78_U141 ( .A1(u5_mult_78_n64), .A2(u5_mult_78_n50), .ZN(
        u5_mult_78_ab_3__0_) );
  NOR2_X1 u5_mult_78_U140 ( .A1(u5_mult_78_n54), .A2(u5_mult_78_n50), .ZN(
        u5_mult_78_ab_3__10_) );
  NOR2_X1 u5_mult_78_U139 ( .A1(u5_mult_78_n63), .A2(u5_mult_78_n50), .ZN(
        u5_mult_78_ab_3__1_) );
  NOR2_X1 u5_mult_78_U138 ( .A1(u5_mult_78_n62), .A2(u5_mult_78_n50), .ZN(
        u5_mult_78_ab_3__2_) );
  NOR2_X1 u5_mult_78_U137 ( .A1(u5_mult_78_n61), .A2(u5_mult_78_n50), .ZN(
        u5_mult_78_ab_3__3_) );
  NOR2_X1 u5_mult_78_U136 ( .A1(u5_mult_78_n60), .A2(u5_mult_78_n50), .ZN(
        u5_mult_78_ab_3__4_) );
  NOR2_X1 u5_mult_78_U135 ( .A1(u5_mult_78_n59), .A2(u5_mult_78_n50), .ZN(
        u5_mult_78_ab_3__5_) );
  NOR2_X1 u5_mult_78_U134 ( .A1(u5_mult_78_n58), .A2(u5_mult_78_n50), .ZN(
        u5_mult_78_ab_3__6_) );
  NOR2_X1 u5_mult_78_U133 ( .A1(u5_mult_78_n57), .A2(u5_mult_78_n50), .ZN(
        u5_mult_78_ab_3__7_) );
  NOR2_X1 u5_mult_78_U132 ( .A1(u5_mult_78_n56), .A2(u5_mult_78_n50), .ZN(
        u5_mult_78_ab_3__8_) );
  NOR2_X1 u5_mult_78_U131 ( .A1(u5_mult_78_n55), .A2(u5_mult_78_n50), .ZN(
        u5_mult_78_ab_3__9_) );
  NOR2_X1 u5_mult_78_U130 ( .A1(u5_mult_78_n64), .A2(u5_mult_78_n49), .ZN(
        u5_mult_78_ab_4__0_) );
  NOR2_X1 u5_mult_78_U129 ( .A1(u5_mult_78_n54), .A2(u5_mult_78_n49), .ZN(
        u5_mult_78_ab_4__10_) );
  NOR2_X1 u5_mult_78_U128 ( .A1(u5_mult_78_n63), .A2(u5_mult_78_n49), .ZN(
        u5_mult_78_ab_4__1_) );
  NOR2_X1 u5_mult_78_U127 ( .A1(u5_mult_78_n62), .A2(u5_mult_78_n49), .ZN(
        u5_mult_78_ab_4__2_) );
  NOR2_X1 u5_mult_78_U126 ( .A1(u5_mult_78_n61), .A2(u5_mult_78_n49), .ZN(
        u5_mult_78_ab_4__3_) );
  NOR2_X1 u5_mult_78_U125 ( .A1(u5_mult_78_n60), .A2(u5_mult_78_n49), .ZN(
        u5_mult_78_ab_4__4_) );
  NOR2_X1 u5_mult_78_U124 ( .A1(u5_mult_78_n59), .A2(u5_mult_78_n49), .ZN(
        u5_mult_78_ab_4__5_) );
  NOR2_X1 u5_mult_78_U123 ( .A1(u5_mult_78_n58), .A2(u5_mult_78_n49), .ZN(
        u5_mult_78_ab_4__6_) );
  NOR2_X1 u5_mult_78_U122 ( .A1(u5_mult_78_n57), .A2(u5_mult_78_n49), .ZN(
        u5_mult_78_ab_4__7_) );
  NOR2_X1 u5_mult_78_U121 ( .A1(u5_mult_78_n56), .A2(u5_mult_78_n49), .ZN(
        u5_mult_78_ab_4__8_) );
  NOR2_X1 u5_mult_78_U120 ( .A1(u5_mult_78_n55), .A2(u5_mult_78_n49), .ZN(
        u5_mult_78_ab_4__9_) );
  NOR2_X1 u5_mult_78_U119 ( .A1(u5_mult_78_n64), .A2(u5_mult_78_n48), .ZN(
        u5_mult_78_ab_5__0_) );
  NOR2_X1 u5_mult_78_U118 ( .A1(u5_mult_78_n54), .A2(u5_mult_78_n48), .ZN(
        u5_mult_78_ab_5__10_) );
  NOR2_X1 u5_mult_78_U117 ( .A1(u5_mult_78_n63), .A2(u5_mult_78_n48), .ZN(
        u5_mult_78_ab_5__1_) );
  NOR2_X1 u5_mult_78_U116 ( .A1(u5_mult_78_n62), .A2(u5_mult_78_n48), .ZN(
        u5_mult_78_ab_5__2_) );
  NOR2_X1 u5_mult_78_U115 ( .A1(u5_mult_78_n61), .A2(u5_mult_78_n48), .ZN(
        u5_mult_78_ab_5__3_) );
  NOR2_X1 u5_mult_78_U114 ( .A1(u5_mult_78_n60), .A2(u5_mult_78_n48), .ZN(
        u5_mult_78_ab_5__4_) );
  NOR2_X1 u5_mult_78_U113 ( .A1(u5_mult_78_n59), .A2(u5_mult_78_n48), .ZN(
        u5_mult_78_ab_5__5_) );
  NOR2_X1 u5_mult_78_U112 ( .A1(u5_mult_78_n58), .A2(u5_mult_78_n48), .ZN(
        u5_mult_78_ab_5__6_) );
  NOR2_X1 u5_mult_78_U111 ( .A1(u5_mult_78_n57), .A2(u5_mult_78_n48), .ZN(
        u5_mult_78_ab_5__7_) );
  NOR2_X1 u5_mult_78_U110 ( .A1(u5_mult_78_n56), .A2(u5_mult_78_n48), .ZN(
        u5_mult_78_ab_5__8_) );
  NOR2_X1 u5_mult_78_U109 ( .A1(u5_mult_78_n55), .A2(u5_mult_78_n48), .ZN(
        u5_mult_78_ab_5__9_) );
  NOR2_X1 u5_mult_78_U108 ( .A1(u5_mult_78_n64), .A2(u5_mult_78_n47), .ZN(
        u5_mult_78_ab_6__0_) );
  NOR2_X1 u5_mult_78_U107 ( .A1(u5_mult_78_n54), .A2(u5_mult_78_n47), .ZN(
        u5_mult_78_ab_6__10_) );
  NOR2_X1 u5_mult_78_U106 ( .A1(u5_mult_78_n63), .A2(u5_mult_78_n47), .ZN(
        u5_mult_78_ab_6__1_) );
  NOR2_X1 u5_mult_78_U105 ( .A1(u5_mult_78_n62), .A2(u5_mult_78_n47), .ZN(
        u5_mult_78_ab_6__2_) );
  NOR2_X1 u5_mult_78_U104 ( .A1(u5_mult_78_n61), .A2(u5_mult_78_n47), .ZN(
        u5_mult_78_ab_6__3_) );
  NOR2_X1 u5_mult_78_U103 ( .A1(u5_mult_78_n60), .A2(u5_mult_78_n47), .ZN(
        u5_mult_78_ab_6__4_) );
  NOR2_X1 u5_mult_78_U102 ( .A1(u5_mult_78_n59), .A2(u5_mult_78_n47), .ZN(
        u5_mult_78_ab_6__5_) );
  NOR2_X1 u5_mult_78_U101 ( .A1(u5_mult_78_n58), .A2(u5_mult_78_n47), .ZN(
        u5_mult_78_ab_6__6_) );
  NOR2_X1 u5_mult_78_U100 ( .A1(u5_mult_78_n57), .A2(u5_mult_78_n47), .ZN(
        u5_mult_78_ab_6__7_) );
  NOR2_X1 u5_mult_78_U99 ( .A1(u5_mult_78_n56), .A2(u5_mult_78_n47), .ZN(
        u5_mult_78_ab_6__8_) );
  NOR2_X1 u5_mult_78_U98 ( .A1(u5_mult_78_n55), .A2(u5_mult_78_n47), .ZN(
        u5_mult_78_ab_6__9_) );
  NOR2_X1 u5_mult_78_U97 ( .A1(u5_mult_78_n64), .A2(u5_mult_78_n46), .ZN(
        u5_mult_78_ab_7__0_) );
  NOR2_X1 u5_mult_78_U96 ( .A1(u5_mult_78_n54), .A2(u5_mult_78_n46), .ZN(
        u5_mult_78_ab_7__10_) );
  NOR2_X1 u5_mult_78_U95 ( .A1(u5_mult_78_n63), .A2(u5_mult_78_n46), .ZN(
        u5_mult_78_ab_7__1_) );
  NOR2_X1 u5_mult_78_U94 ( .A1(u5_mult_78_n62), .A2(u5_mult_78_n46), .ZN(
        u5_mult_78_ab_7__2_) );
  NOR2_X1 u5_mult_78_U93 ( .A1(u5_mult_78_n61), .A2(u5_mult_78_n46), .ZN(
        u5_mult_78_ab_7__3_) );
  NOR2_X1 u5_mult_78_U92 ( .A1(u5_mult_78_n60), .A2(u5_mult_78_n46), .ZN(
        u5_mult_78_ab_7__4_) );
  NOR2_X1 u5_mult_78_U91 ( .A1(u5_mult_78_n59), .A2(u5_mult_78_n46), .ZN(
        u5_mult_78_ab_7__5_) );
  NOR2_X1 u5_mult_78_U90 ( .A1(u5_mult_78_n58), .A2(u5_mult_78_n46), .ZN(
        u5_mult_78_ab_7__6_) );
  NOR2_X1 u5_mult_78_U89 ( .A1(u5_mult_78_n57), .A2(u5_mult_78_n46), .ZN(
        u5_mult_78_ab_7__7_) );
  NOR2_X1 u5_mult_78_U88 ( .A1(u5_mult_78_n56), .A2(u5_mult_78_n46), .ZN(
        u5_mult_78_ab_7__8_) );
  NOR2_X1 u5_mult_78_U87 ( .A1(u5_mult_78_n55), .A2(u5_mult_78_n46), .ZN(
        u5_mult_78_ab_7__9_) );
  NOR2_X1 u5_mult_78_U86 ( .A1(u5_mult_78_n64), .A2(u5_mult_78_n45), .ZN(
        u5_mult_78_ab_8__0_) );
  NOR2_X1 u5_mult_78_U85 ( .A1(u5_mult_78_n54), .A2(u5_mult_78_n45), .ZN(
        u5_mult_78_ab_8__10_) );
  NOR2_X1 u5_mult_78_U84 ( .A1(u5_mult_78_n63), .A2(u5_mult_78_n45), .ZN(
        u5_mult_78_ab_8__1_) );
  NOR2_X1 u5_mult_78_U83 ( .A1(u5_mult_78_n62), .A2(u5_mult_78_n45), .ZN(
        u5_mult_78_ab_8__2_) );
  NOR2_X1 u5_mult_78_U82 ( .A1(u5_mult_78_n61), .A2(u5_mult_78_n45), .ZN(
        u5_mult_78_ab_8__3_) );
  NOR2_X1 u5_mult_78_U81 ( .A1(u5_mult_78_n60), .A2(u5_mult_78_n45), .ZN(
        u5_mult_78_ab_8__4_) );
  NOR2_X1 u5_mult_78_U80 ( .A1(u5_mult_78_n59), .A2(u5_mult_78_n45), .ZN(
        u5_mult_78_ab_8__5_) );
  NOR2_X1 u5_mult_78_U79 ( .A1(u5_mult_78_n58), .A2(u5_mult_78_n45), .ZN(
        u5_mult_78_ab_8__6_) );
  NOR2_X1 u5_mult_78_U78 ( .A1(u5_mult_78_n57), .A2(u5_mult_78_n45), .ZN(
        u5_mult_78_ab_8__7_) );
  NOR2_X1 u5_mult_78_U77 ( .A1(u5_mult_78_n56), .A2(u5_mult_78_n45), .ZN(
        u5_mult_78_ab_8__8_) );
  NOR2_X1 u5_mult_78_U76 ( .A1(u5_mult_78_n55), .A2(u5_mult_78_n45), .ZN(
        u5_mult_78_ab_8__9_) );
  NOR2_X1 u5_mult_78_U75 ( .A1(u5_mult_78_n44), .A2(u5_mult_78_n64), .ZN(
        u5_mult_78_ab_9__0_) );
  NOR2_X1 u5_mult_78_U74 ( .A1(u5_mult_78_n44), .A2(u5_mult_78_n54), .ZN(
        u5_mult_78_ab_9__10_) );
  NOR2_X1 u5_mult_78_U73 ( .A1(u5_mult_78_n44), .A2(u5_mult_78_n63), .ZN(
        u5_mult_78_ab_9__1_) );
  NOR2_X1 u5_mult_78_U72 ( .A1(u5_mult_78_n44), .A2(u5_mult_78_n62), .ZN(
        u5_mult_78_ab_9__2_) );
  NOR2_X1 u5_mult_78_U71 ( .A1(u5_mult_78_n44), .A2(u5_mult_78_n61), .ZN(
        u5_mult_78_ab_9__3_) );
  NOR2_X1 u5_mult_78_U70 ( .A1(u5_mult_78_n44), .A2(u5_mult_78_n60), .ZN(
        u5_mult_78_ab_9__4_) );
  NOR2_X1 u5_mult_78_U69 ( .A1(u5_mult_78_n44), .A2(u5_mult_78_n59), .ZN(
        u5_mult_78_ab_9__5_) );
  NOR2_X1 u5_mult_78_U68 ( .A1(u5_mult_78_n44), .A2(u5_mult_78_n58), .ZN(
        u5_mult_78_ab_9__6_) );
  NOR2_X1 u5_mult_78_U67 ( .A1(u5_mult_78_n44), .A2(u5_mult_78_n57), .ZN(
        u5_mult_78_ab_9__7_) );
  NOR2_X1 u5_mult_78_U66 ( .A1(u5_mult_78_n44), .A2(u5_mult_78_n56), .ZN(
        u5_mult_78_ab_9__8_) );
  NOR2_X1 u5_mult_78_U65 ( .A1(u5_mult_78_n44), .A2(u5_mult_78_n55), .ZN(
        u5_mult_78_ab_9__9_) );
  XOR2_X2 u5_mult_78_U63 ( .A(u5_mult_78_ab_1__0_), .B(u5_mult_78_ab_0__1_), 
        .Z(u5_N1) );
  XOR2_X2 u5_mult_78_U62 ( .A(u5_mult_78_CARRYB_10__0_), .B(
        u5_mult_78_SUMB_10__1_), .Z(u5_N11) );
  AND2_X4 u5_mult_78_U61 ( .A1(u5_mult_78_SUMB_10__1_), .A2(
        u5_mult_78_CARRYB_10__0_), .ZN(u5_mult_78_n40) );
  AND2_X4 u5_mult_78_U60 ( .A1(u5_mult_78_SUMB_10__3_), .A2(
        u5_mult_78_CARRYB_10__2_), .ZN(u5_mult_78_n39) );
  AND2_X4 u5_mult_78_U59 ( .A1(u5_mult_78_SUMB_10__5_), .A2(
        u5_mult_78_CARRYB_10__4_), .ZN(u5_mult_78_n38) );
  AND2_X4 u5_mult_78_U58 ( .A1(u5_mult_78_SUMB_10__7_), .A2(
        u5_mult_78_CARRYB_10__6_), .ZN(u5_mult_78_n37) );
  AND2_X4 u5_mult_78_U57 ( .A1(u5_mult_78_SUMB_10__9_), .A2(
        u5_mult_78_CARRYB_10__8_), .ZN(u5_mult_78_n36) );
  AND2_X4 u5_mult_78_U56 ( .A1(u5_mult_78_SUMB_10__2_), .A2(
        u5_mult_78_CARRYB_10__1_), .ZN(u5_mult_78_n35) );
  AND2_X4 u5_mult_78_U55 ( .A1(u5_mult_78_SUMB_10__4_), .A2(
        u5_mult_78_CARRYB_10__3_), .ZN(u5_mult_78_n34) );
  AND2_X4 u5_mult_78_U54 ( .A1(u5_mult_78_SUMB_10__6_), .A2(
        u5_mult_78_CARRYB_10__5_), .ZN(u5_mult_78_n33) );
  AND2_X4 u5_mult_78_U53 ( .A1(u5_mult_78_SUMB_10__8_), .A2(
        u5_mult_78_CARRYB_10__7_), .ZN(u5_mult_78_n32) );
  AND2_X4 u5_mult_78_U52 ( .A1(u5_mult_78_ab_10__10_), .A2(
        u5_mult_78_CARRYB_10__9_), .ZN(u5_mult_78_n31) );
  XOR2_X2 u5_mult_78_U51 ( .A(u5_mult_78_ab_1__1_), .B(u5_mult_78_ab_0__2_), 
        .Z(u5_mult_78_n30) );
  XOR2_X2 u5_mult_78_U50 ( .A(u5_mult_78_ab_1__2_), .B(u5_mult_78_ab_0__3_), 
        .Z(u5_mult_78_n29) );
  XOR2_X2 u5_mult_78_U49 ( .A(u5_mult_78_ab_1__3_), .B(u5_mult_78_ab_0__4_), 
        .Z(u5_mult_78_n28) );
  XOR2_X2 u5_mult_78_U48 ( .A(u5_mult_78_ab_1__4_), .B(u5_mult_78_ab_0__5_), 
        .Z(u5_mult_78_n27) );
  XOR2_X2 u5_mult_78_U47 ( .A(u5_mult_78_ab_1__5_), .B(u5_mult_78_ab_0__6_), 
        .Z(u5_mult_78_n26) );
  XOR2_X2 u5_mult_78_U46 ( .A(u5_mult_78_ab_1__6_), .B(u5_mult_78_ab_0__7_), 
        .Z(u5_mult_78_n25) );
  XOR2_X2 u5_mult_78_U45 ( .A(u5_mult_78_ab_1__7_), .B(u5_mult_78_ab_0__8_), 
        .Z(u5_mult_78_n24) );
  XOR2_X2 u5_mult_78_U44 ( .A(u5_mult_78_ab_1__8_), .B(u5_mult_78_ab_0__9_), 
        .Z(u5_mult_78_n23) );
  XOR2_X2 u5_mult_78_U43 ( .A(u5_mult_78_ab_1__9_), .B(u5_mult_78_ab_0__10_), 
        .Z(u5_mult_78_n22) );
  AND2_X4 u5_mult_78_U42 ( .A1(u5_mult_78_ab_0__10_), .A2(u5_mult_78_ab_1__9_), 
        .ZN(u5_mult_78_n21) );
  XOR2_X2 u5_mult_78_U41 ( .A(u5_mult_78_CARRYB_10__3_), .B(
        u5_mult_78_SUMB_10__4_), .Z(u5_mult_78_n20) );
  XOR2_X2 u5_mult_78_U40 ( .A(u5_mult_78_CARRYB_10__5_), .B(
        u5_mult_78_SUMB_10__6_), .Z(u5_mult_78_n19) );
  XOR2_X2 u5_mult_78_U39 ( .A(u5_mult_78_CARRYB_10__7_), .B(
        u5_mult_78_SUMB_10__8_), .Z(u5_mult_78_n18) );
  XOR2_X2 u5_mult_78_U38 ( .A(u5_mult_78_CARRYB_10__1_), .B(
        u5_mult_78_SUMB_10__2_), .Z(u5_mult_78_n17) );
  XOR2_X2 u5_mult_78_U37 ( .A(u5_mult_78_CARRYB_10__2_), .B(
        u5_mult_78_SUMB_10__3_), .Z(u5_mult_78_n16) );
  XOR2_X2 u5_mult_78_U36 ( .A(u5_mult_78_CARRYB_10__4_), .B(
        u5_mult_78_SUMB_10__5_), .Z(u5_mult_78_n15) );
  XOR2_X2 u5_mult_78_U35 ( .A(u5_mult_78_CARRYB_10__6_), .B(
        u5_mult_78_SUMB_10__7_), .Z(u5_mult_78_n14) );
  XOR2_X2 u5_mult_78_U34 ( .A(u5_mult_78_CARRYB_10__8_), .B(
        u5_mult_78_SUMB_10__9_), .Z(u5_mult_78_n13) );
  XOR2_X2 u5_mult_78_U33 ( .A(u5_mult_78_CARRYB_10__9_), .B(
        u5_mult_78_ab_10__10_), .Z(u5_mult_78_n12) );
  AND2_X4 u5_mult_78_U32 ( .A1(u5_mult_78_ab_0__1_), .A2(u5_mult_78_ab_1__0_), 
        .ZN(u5_mult_78_n11) );
  AND2_X4 u5_mult_78_U31 ( .A1(u5_mult_78_ab_0__2_), .A2(u5_mult_78_ab_1__1_), 
        .ZN(u5_mult_78_n10) );
  AND2_X4 u5_mult_78_U30 ( .A1(u5_mult_78_ab_0__3_), .A2(u5_mult_78_ab_1__2_), 
        .ZN(u5_mult_78_n9) );
  AND2_X4 u5_mult_78_U29 ( .A1(u5_mult_78_ab_0__4_), .A2(u5_mult_78_ab_1__3_), 
        .ZN(u5_mult_78_n8) );
  AND2_X4 u5_mult_78_U28 ( .A1(u5_mult_78_ab_0__5_), .A2(u5_mult_78_ab_1__4_), 
        .ZN(u5_mult_78_n7) );
  AND2_X4 u5_mult_78_U27 ( .A1(u5_mult_78_ab_0__6_), .A2(u5_mult_78_ab_1__5_), 
        .ZN(u5_mult_78_n6) );
  AND2_X4 u5_mult_78_U26 ( .A1(u5_mult_78_ab_0__7_), .A2(u5_mult_78_ab_1__6_), 
        .ZN(u5_mult_78_n5) );
  AND2_X4 u5_mult_78_U25 ( .A1(u5_mult_78_ab_0__8_), .A2(u5_mult_78_ab_1__7_), 
        .ZN(u5_mult_78_n4) );
  AND2_X4 u5_mult_78_U24 ( .A1(u5_mult_78_ab_0__9_), .A2(u5_mult_78_ab_1__8_), 
        .ZN(u5_mult_78_n3) );
  INV_X4 u5_mult_78_U23 ( .A(u6_N0), .ZN(u5_mult_78_n64) );
  INV_X4 u5_mult_78_U22 ( .A(fracta_mul[0]), .ZN(u5_mult_78_n53) );
  INV_X4 u5_mult_78_U21 ( .A(fracta_mul[2]), .ZN(u5_mult_78_n51) );
  INV_X4 u5_mult_78_U20 ( .A(fracta_mul[3]), .ZN(u5_mult_78_n50) );
  INV_X4 u5_mult_78_U19 ( .A(fracta_mul[4]), .ZN(u5_mult_78_n49) );
  INV_X4 u5_mult_78_U18 ( .A(fracta_mul[5]), .ZN(u5_mult_78_n48) );
  INV_X4 u5_mult_78_U17 ( .A(fracta_mul[6]), .ZN(u5_mult_78_n47) );
  INV_X4 u5_mult_78_U16 ( .A(fracta_mul[7]), .ZN(u5_mult_78_n46) );
  INV_X4 u5_mult_78_U15 ( .A(fracta_mul[8]), .ZN(u5_mult_78_n45) );
  INV_X4 u5_mult_78_U14 ( .A(fracta_mul[9]), .ZN(u5_mult_78_n44) );
  INV_X4 u5_mult_78_U13 ( .A(n2698), .ZN(u5_mult_78_n43) );
  INV_X4 u5_mult_78_U12 ( .A(u6_N1), .ZN(u5_mult_78_n63) );
  INV_X4 u5_mult_78_U11 ( .A(fracta_mul[1]), .ZN(u5_mult_78_n52) );
  INV_X4 u5_mult_78_U10 ( .A(u6_N2), .ZN(u5_mult_78_n62) );
  INV_X4 u5_mult_78_U9 ( .A(u6_N10), .ZN(u5_mult_78_n54) );
  INV_X4 u5_mult_78_U8 ( .A(u6_N9), .ZN(u5_mult_78_n55) );
  INV_X4 u5_mult_78_U7 ( .A(u6_N3), .ZN(u5_mult_78_n61) );
  INV_X4 u5_mult_78_U6 ( .A(u6_N4), .ZN(u5_mult_78_n60) );
  INV_X4 u5_mult_78_U5 ( .A(u6_N5), .ZN(u5_mult_78_n59) );
  INV_X4 u5_mult_78_U4 ( .A(u6_N6), .ZN(u5_mult_78_n58) );
  INV_X4 u5_mult_78_U3 ( .A(u6_N7), .ZN(u5_mult_78_n57) );
  INV_X4 u5_mult_78_U2 ( .A(u6_N8), .ZN(u5_mult_78_n56) );
  FA_X1 u5_mult_78_S3_2_9 ( .A(u5_mult_78_ab_2__9_), .B(u5_mult_78_n21), .CI(
        u5_mult_78_ab_1__10_), .CO(u5_mult_78_CARRYB_2__9_), .S(
        u5_mult_78_SUMB_2__9_) );
  FA_X1 u5_mult_78_S2_2_8 ( .A(u5_mult_78_ab_2__8_), .B(u5_mult_78_n3), .CI(
        u5_mult_78_n22), .CO(u5_mult_78_CARRYB_2__8_), .S(
        u5_mult_78_SUMB_2__8_) );
  FA_X1 u5_mult_78_S2_2_7 ( .A(u5_mult_78_ab_2__7_), .B(u5_mult_78_n4), .CI(
        u5_mult_78_n23), .CO(u5_mult_78_CARRYB_2__7_), .S(
        u5_mult_78_SUMB_2__7_) );
  FA_X1 u5_mult_78_S2_2_6 ( .A(u5_mult_78_ab_2__6_), .B(u5_mult_78_n5), .CI(
        u5_mult_78_n24), .CO(u5_mult_78_CARRYB_2__6_), .S(
        u5_mult_78_SUMB_2__6_) );
  FA_X1 u5_mult_78_S2_2_5 ( .A(u5_mult_78_ab_2__5_), .B(u5_mult_78_n6), .CI(
        u5_mult_78_n25), .CO(u5_mult_78_CARRYB_2__5_), .S(
        u5_mult_78_SUMB_2__5_) );
  FA_X1 u5_mult_78_S2_2_4 ( .A(u5_mult_78_ab_2__4_), .B(u5_mult_78_n7), .CI(
        u5_mult_78_n26), .CO(u5_mult_78_CARRYB_2__4_), .S(
        u5_mult_78_SUMB_2__4_) );
  FA_X1 u5_mult_78_S2_2_3 ( .A(u5_mult_78_ab_2__3_), .B(u5_mult_78_n8), .CI(
        u5_mult_78_n27), .CO(u5_mult_78_CARRYB_2__3_), .S(
        u5_mult_78_SUMB_2__3_) );
  FA_X1 u5_mult_78_S2_2_2 ( .A(u5_mult_78_ab_2__2_), .B(u5_mult_78_n9), .CI(
        u5_mult_78_n28), .CO(u5_mult_78_CARRYB_2__2_), .S(
        u5_mult_78_SUMB_2__2_) );
  FA_X1 u5_mult_78_S2_2_1 ( .A(u5_mult_78_ab_2__1_), .B(u5_mult_78_n10), .CI(
        u5_mult_78_n29), .CO(u5_mult_78_CARRYB_2__1_), .S(
        u5_mult_78_SUMB_2__1_) );
  FA_X1 u5_mult_78_S1_2_0 ( .A(u5_mult_78_ab_2__0_), .B(u5_mult_78_n11), .CI(
        u5_mult_78_n30), .CO(u5_mult_78_CARRYB_2__0_), .S(u5_N2) );
  FA_X1 u5_mult_78_S3_3_9 ( .A(u5_mult_78_ab_3__9_), .B(
        u5_mult_78_CARRYB_2__9_), .CI(u5_mult_78_ab_2__10_), .CO(
        u5_mult_78_CARRYB_3__9_), .S(u5_mult_78_SUMB_3__9_) );
  FA_X1 u5_mult_78_S2_3_8 ( .A(u5_mult_78_ab_3__8_), .B(
        u5_mult_78_CARRYB_2__8_), .CI(u5_mult_78_SUMB_2__9_), .CO(
        u5_mult_78_CARRYB_3__8_), .S(u5_mult_78_SUMB_3__8_) );
  FA_X1 u5_mult_78_S2_3_7 ( .A(u5_mult_78_ab_3__7_), .B(
        u5_mult_78_CARRYB_2__7_), .CI(u5_mult_78_SUMB_2__8_), .CO(
        u5_mult_78_CARRYB_3__7_), .S(u5_mult_78_SUMB_3__7_) );
  FA_X1 u5_mult_78_S2_3_6 ( .A(u5_mult_78_ab_3__6_), .B(
        u5_mult_78_CARRYB_2__6_), .CI(u5_mult_78_SUMB_2__7_), .CO(
        u5_mult_78_CARRYB_3__6_), .S(u5_mult_78_SUMB_3__6_) );
  FA_X1 u5_mult_78_S2_3_5 ( .A(u5_mult_78_ab_3__5_), .B(
        u5_mult_78_CARRYB_2__5_), .CI(u5_mult_78_SUMB_2__6_), .CO(
        u5_mult_78_CARRYB_3__5_), .S(u5_mult_78_SUMB_3__5_) );
  FA_X1 u5_mult_78_S2_3_4 ( .A(u5_mult_78_ab_3__4_), .B(
        u5_mult_78_CARRYB_2__4_), .CI(u5_mult_78_SUMB_2__5_), .CO(
        u5_mult_78_CARRYB_3__4_), .S(u5_mult_78_SUMB_3__4_) );
  FA_X1 u5_mult_78_S2_3_3 ( .A(u5_mult_78_ab_3__3_), .B(
        u5_mult_78_CARRYB_2__3_), .CI(u5_mult_78_SUMB_2__4_), .CO(
        u5_mult_78_CARRYB_3__3_), .S(u5_mult_78_SUMB_3__3_) );
  FA_X1 u5_mult_78_S2_3_2 ( .A(u5_mult_78_ab_3__2_), .B(
        u5_mult_78_CARRYB_2__2_), .CI(u5_mult_78_SUMB_2__3_), .CO(
        u5_mult_78_CARRYB_3__2_), .S(u5_mult_78_SUMB_3__2_) );
  FA_X1 u5_mult_78_S2_3_1 ( .A(u5_mult_78_ab_3__1_), .B(
        u5_mult_78_CARRYB_2__1_), .CI(u5_mult_78_SUMB_2__2_), .CO(
        u5_mult_78_CARRYB_3__1_), .S(u5_mult_78_SUMB_3__1_) );
  FA_X1 u5_mult_78_S1_3_0 ( .A(u5_mult_78_ab_3__0_), .B(
        u5_mult_78_CARRYB_2__0_), .CI(u5_mult_78_SUMB_2__1_), .CO(
        u5_mult_78_CARRYB_3__0_), .S(u5_N3) );
  FA_X1 u5_mult_78_S3_4_9 ( .A(u5_mult_78_ab_4__9_), .B(
        u5_mult_78_CARRYB_3__9_), .CI(u5_mult_78_ab_3__10_), .CO(
        u5_mult_78_CARRYB_4__9_), .S(u5_mult_78_SUMB_4__9_) );
  FA_X1 u5_mult_78_S2_4_8 ( .A(u5_mult_78_ab_4__8_), .B(
        u5_mult_78_CARRYB_3__8_), .CI(u5_mult_78_SUMB_3__9_), .CO(
        u5_mult_78_CARRYB_4__8_), .S(u5_mult_78_SUMB_4__8_) );
  FA_X1 u5_mult_78_S2_4_7 ( .A(u5_mult_78_ab_4__7_), .B(
        u5_mult_78_CARRYB_3__7_), .CI(u5_mult_78_SUMB_3__8_), .CO(
        u5_mult_78_CARRYB_4__7_), .S(u5_mult_78_SUMB_4__7_) );
  FA_X1 u5_mult_78_S2_4_6 ( .A(u5_mult_78_ab_4__6_), .B(
        u5_mult_78_CARRYB_3__6_), .CI(u5_mult_78_SUMB_3__7_), .CO(
        u5_mult_78_CARRYB_4__6_), .S(u5_mult_78_SUMB_4__6_) );
  FA_X1 u5_mult_78_S2_4_5 ( .A(u5_mult_78_ab_4__5_), .B(
        u5_mult_78_CARRYB_3__5_), .CI(u5_mult_78_SUMB_3__6_), .CO(
        u5_mult_78_CARRYB_4__5_), .S(u5_mult_78_SUMB_4__5_) );
  FA_X1 u5_mult_78_S2_4_4 ( .A(u5_mult_78_ab_4__4_), .B(
        u5_mult_78_CARRYB_3__4_), .CI(u5_mult_78_SUMB_3__5_), .CO(
        u5_mult_78_CARRYB_4__4_), .S(u5_mult_78_SUMB_4__4_) );
  FA_X1 u5_mult_78_S2_4_3 ( .A(u5_mult_78_ab_4__3_), .B(
        u5_mult_78_CARRYB_3__3_), .CI(u5_mult_78_SUMB_3__4_), .CO(
        u5_mult_78_CARRYB_4__3_), .S(u5_mult_78_SUMB_4__3_) );
  FA_X1 u5_mult_78_S2_4_2 ( .A(u5_mult_78_ab_4__2_), .B(
        u5_mult_78_CARRYB_3__2_), .CI(u5_mult_78_SUMB_3__3_), .CO(
        u5_mult_78_CARRYB_4__2_), .S(u5_mult_78_SUMB_4__2_) );
  FA_X1 u5_mult_78_S2_4_1 ( .A(u5_mult_78_ab_4__1_), .B(
        u5_mult_78_CARRYB_3__1_), .CI(u5_mult_78_SUMB_3__2_), .CO(
        u5_mult_78_CARRYB_4__1_), .S(u5_mult_78_SUMB_4__1_) );
  FA_X1 u5_mult_78_S1_4_0 ( .A(u5_mult_78_ab_4__0_), .B(
        u5_mult_78_CARRYB_3__0_), .CI(u5_mult_78_SUMB_3__1_), .CO(
        u5_mult_78_CARRYB_4__0_), .S(u5_N4) );
  FA_X1 u5_mult_78_S3_5_9 ( .A(u5_mult_78_ab_5__9_), .B(
        u5_mult_78_CARRYB_4__9_), .CI(u5_mult_78_ab_4__10_), .CO(
        u5_mult_78_CARRYB_5__9_), .S(u5_mult_78_SUMB_5__9_) );
  FA_X1 u5_mult_78_S2_5_8 ( .A(u5_mult_78_ab_5__8_), .B(
        u5_mult_78_CARRYB_4__8_), .CI(u5_mult_78_SUMB_4__9_), .CO(
        u5_mult_78_CARRYB_5__8_), .S(u5_mult_78_SUMB_5__8_) );
  FA_X1 u5_mult_78_S2_5_7 ( .A(u5_mult_78_ab_5__7_), .B(
        u5_mult_78_CARRYB_4__7_), .CI(u5_mult_78_SUMB_4__8_), .CO(
        u5_mult_78_CARRYB_5__7_), .S(u5_mult_78_SUMB_5__7_) );
  FA_X1 u5_mult_78_S2_5_6 ( .A(u5_mult_78_ab_5__6_), .B(
        u5_mult_78_CARRYB_4__6_), .CI(u5_mult_78_SUMB_4__7_), .CO(
        u5_mult_78_CARRYB_5__6_), .S(u5_mult_78_SUMB_5__6_) );
  FA_X1 u5_mult_78_S2_5_5 ( .A(u5_mult_78_ab_5__5_), .B(
        u5_mult_78_CARRYB_4__5_), .CI(u5_mult_78_SUMB_4__6_), .CO(
        u5_mult_78_CARRYB_5__5_), .S(u5_mult_78_SUMB_5__5_) );
  FA_X1 u5_mult_78_S2_5_4 ( .A(u5_mult_78_ab_5__4_), .B(
        u5_mult_78_CARRYB_4__4_), .CI(u5_mult_78_SUMB_4__5_), .CO(
        u5_mult_78_CARRYB_5__4_), .S(u5_mult_78_SUMB_5__4_) );
  FA_X1 u5_mult_78_S2_5_3 ( .A(u5_mult_78_ab_5__3_), .B(
        u5_mult_78_CARRYB_4__3_), .CI(u5_mult_78_SUMB_4__4_), .CO(
        u5_mult_78_CARRYB_5__3_), .S(u5_mult_78_SUMB_5__3_) );
  FA_X1 u5_mult_78_S2_5_2 ( .A(u5_mult_78_ab_5__2_), .B(
        u5_mult_78_CARRYB_4__2_), .CI(u5_mult_78_SUMB_4__3_), .CO(
        u5_mult_78_CARRYB_5__2_), .S(u5_mult_78_SUMB_5__2_) );
  FA_X1 u5_mult_78_S2_5_1 ( .A(u5_mult_78_ab_5__1_), .B(
        u5_mult_78_CARRYB_4__1_), .CI(u5_mult_78_SUMB_4__2_), .CO(
        u5_mult_78_CARRYB_5__1_), .S(u5_mult_78_SUMB_5__1_) );
  FA_X1 u5_mult_78_S1_5_0 ( .A(u5_mult_78_ab_5__0_), .B(
        u5_mult_78_CARRYB_4__0_), .CI(u5_mult_78_SUMB_4__1_), .CO(
        u5_mult_78_CARRYB_5__0_), .S(u5_N5) );
  FA_X1 u5_mult_78_S3_6_9 ( .A(u5_mult_78_ab_6__9_), .B(
        u5_mult_78_CARRYB_5__9_), .CI(u5_mult_78_ab_5__10_), .CO(
        u5_mult_78_CARRYB_6__9_), .S(u5_mult_78_SUMB_6__9_) );
  FA_X1 u5_mult_78_S2_6_8 ( .A(u5_mult_78_ab_6__8_), .B(
        u5_mult_78_CARRYB_5__8_), .CI(u5_mult_78_SUMB_5__9_), .CO(
        u5_mult_78_CARRYB_6__8_), .S(u5_mult_78_SUMB_6__8_) );
  FA_X1 u5_mult_78_S2_6_7 ( .A(u5_mult_78_ab_6__7_), .B(
        u5_mult_78_CARRYB_5__7_), .CI(u5_mult_78_SUMB_5__8_), .CO(
        u5_mult_78_CARRYB_6__7_), .S(u5_mult_78_SUMB_6__7_) );
  FA_X1 u5_mult_78_S2_6_6 ( .A(u5_mult_78_ab_6__6_), .B(
        u5_mult_78_CARRYB_5__6_), .CI(u5_mult_78_SUMB_5__7_), .CO(
        u5_mult_78_CARRYB_6__6_), .S(u5_mult_78_SUMB_6__6_) );
  FA_X1 u5_mult_78_S2_6_5 ( .A(u5_mult_78_ab_6__5_), .B(
        u5_mult_78_CARRYB_5__5_), .CI(u5_mult_78_SUMB_5__6_), .CO(
        u5_mult_78_CARRYB_6__5_), .S(u5_mult_78_SUMB_6__5_) );
  FA_X1 u5_mult_78_S2_6_4 ( .A(u5_mult_78_ab_6__4_), .B(
        u5_mult_78_CARRYB_5__4_), .CI(u5_mult_78_SUMB_5__5_), .CO(
        u5_mult_78_CARRYB_6__4_), .S(u5_mult_78_SUMB_6__4_) );
  FA_X1 u5_mult_78_S2_6_3 ( .A(u5_mult_78_ab_6__3_), .B(
        u5_mult_78_CARRYB_5__3_), .CI(u5_mult_78_SUMB_5__4_), .CO(
        u5_mult_78_CARRYB_6__3_), .S(u5_mult_78_SUMB_6__3_) );
  FA_X1 u5_mult_78_S2_6_2 ( .A(u5_mult_78_ab_6__2_), .B(
        u5_mult_78_CARRYB_5__2_), .CI(u5_mult_78_SUMB_5__3_), .CO(
        u5_mult_78_CARRYB_6__2_), .S(u5_mult_78_SUMB_6__2_) );
  FA_X1 u5_mult_78_S2_6_1 ( .A(u5_mult_78_ab_6__1_), .B(
        u5_mult_78_CARRYB_5__1_), .CI(u5_mult_78_SUMB_5__2_), .CO(
        u5_mult_78_CARRYB_6__1_), .S(u5_mult_78_SUMB_6__1_) );
  FA_X1 u5_mult_78_S1_6_0 ( .A(u5_mult_78_ab_6__0_), .B(
        u5_mult_78_CARRYB_5__0_), .CI(u5_mult_78_SUMB_5__1_), .CO(
        u5_mult_78_CARRYB_6__0_), .S(u5_N6) );
  FA_X1 u5_mult_78_S3_7_9 ( .A(u5_mult_78_ab_7__9_), .B(
        u5_mult_78_CARRYB_6__9_), .CI(u5_mult_78_ab_6__10_), .CO(
        u5_mult_78_CARRYB_7__9_), .S(u5_mult_78_SUMB_7__9_) );
  FA_X1 u5_mult_78_S2_7_8 ( .A(u5_mult_78_ab_7__8_), .B(
        u5_mult_78_CARRYB_6__8_), .CI(u5_mult_78_SUMB_6__9_), .CO(
        u5_mult_78_CARRYB_7__8_), .S(u5_mult_78_SUMB_7__8_) );
  FA_X1 u5_mult_78_S2_7_7 ( .A(u5_mult_78_ab_7__7_), .B(
        u5_mult_78_CARRYB_6__7_), .CI(u5_mult_78_SUMB_6__8_), .CO(
        u5_mult_78_CARRYB_7__7_), .S(u5_mult_78_SUMB_7__7_) );
  FA_X1 u5_mult_78_S2_7_6 ( .A(u5_mult_78_ab_7__6_), .B(
        u5_mult_78_CARRYB_6__6_), .CI(u5_mult_78_SUMB_6__7_), .CO(
        u5_mult_78_CARRYB_7__6_), .S(u5_mult_78_SUMB_7__6_) );
  FA_X1 u5_mult_78_S2_7_5 ( .A(u5_mult_78_ab_7__5_), .B(
        u5_mult_78_CARRYB_6__5_), .CI(u5_mult_78_SUMB_6__6_), .CO(
        u5_mult_78_CARRYB_7__5_), .S(u5_mult_78_SUMB_7__5_) );
  FA_X1 u5_mult_78_S2_7_4 ( .A(u5_mult_78_ab_7__4_), .B(
        u5_mult_78_CARRYB_6__4_), .CI(u5_mult_78_SUMB_6__5_), .CO(
        u5_mult_78_CARRYB_7__4_), .S(u5_mult_78_SUMB_7__4_) );
  FA_X1 u5_mult_78_S2_7_3 ( .A(u5_mult_78_ab_7__3_), .B(
        u5_mult_78_CARRYB_6__3_), .CI(u5_mult_78_SUMB_6__4_), .CO(
        u5_mult_78_CARRYB_7__3_), .S(u5_mult_78_SUMB_7__3_) );
  FA_X1 u5_mult_78_S2_7_2 ( .A(u5_mult_78_ab_7__2_), .B(
        u5_mult_78_CARRYB_6__2_), .CI(u5_mult_78_SUMB_6__3_), .CO(
        u5_mult_78_CARRYB_7__2_), .S(u5_mult_78_SUMB_7__2_) );
  FA_X1 u5_mult_78_S2_7_1 ( .A(u5_mult_78_ab_7__1_), .B(
        u5_mult_78_CARRYB_6__1_), .CI(u5_mult_78_SUMB_6__2_), .CO(
        u5_mult_78_CARRYB_7__1_), .S(u5_mult_78_SUMB_7__1_) );
  FA_X1 u5_mult_78_S1_7_0 ( .A(u5_mult_78_ab_7__0_), .B(
        u5_mult_78_CARRYB_6__0_), .CI(u5_mult_78_SUMB_6__1_), .CO(
        u5_mult_78_CARRYB_7__0_), .S(u5_N7) );
  FA_X1 u5_mult_78_S3_8_9 ( .A(u5_mult_78_ab_8__9_), .B(
        u5_mult_78_CARRYB_7__9_), .CI(u5_mult_78_ab_7__10_), .CO(
        u5_mult_78_CARRYB_8__9_), .S(u5_mult_78_SUMB_8__9_) );
  FA_X1 u5_mult_78_S2_8_8 ( .A(u5_mult_78_ab_8__8_), .B(
        u5_mult_78_CARRYB_7__8_), .CI(u5_mult_78_SUMB_7__9_), .CO(
        u5_mult_78_CARRYB_8__8_), .S(u5_mult_78_SUMB_8__8_) );
  FA_X1 u5_mult_78_S2_8_7 ( .A(u5_mult_78_ab_8__7_), .B(
        u5_mult_78_CARRYB_7__7_), .CI(u5_mult_78_SUMB_7__8_), .CO(
        u5_mult_78_CARRYB_8__7_), .S(u5_mult_78_SUMB_8__7_) );
  FA_X1 u5_mult_78_S2_8_6 ( .A(u5_mult_78_ab_8__6_), .B(
        u5_mult_78_CARRYB_7__6_), .CI(u5_mult_78_SUMB_7__7_), .CO(
        u5_mult_78_CARRYB_8__6_), .S(u5_mult_78_SUMB_8__6_) );
  FA_X1 u5_mult_78_S2_8_5 ( .A(u5_mult_78_ab_8__5_), .B(
        u5_mult_78_CARRYB_7__5_), .CI(u5_mult_78_SUMB_7__6_), .CO(
        u5_mult_78_CARRYB_8__5_), .S(u5_mult_78_SUMB_8__5_) );
  FA_X1 u5_mult_78_S2_8_4 ( .A(u5_mult_78_ab_8__4_), .B(
        u5_mult_78_CARRYB_7__4_), .CI(u5_mult_78_SUMB_7__5_), .CO(
        u5_mult_78_CARRYB_8__4_), .S(u5_mult_78_SUMB_8__4_) );
  FA_X1 u5_mult_78_S2_8_3 ( .A(u5_mult_78_ab_8__3_), .B(
        u5_mult_78_CARRYB_7__3_), .CI(u5_mult_78_SUMB_7__4_), .CO(
        u5_mult_78_CARRYB_8__3_), .S(u5_mult_78_SUMB_8__3_) );
  FA_X1 u5_mult_78_S2_8_2 ( .A(u5_mult_78_ab_8__2_), .B(
        u5_mult_78_CARRYB_7__2_), .CI(u5_mult_78_SUMB_7__3_), .CO(
        u5_mult_78_CARRYB_8__2_), .S(u5_mult_78_SUMB_8__2_) );
  FA_X1 u5_mult_78_S2_8_1 ( .A(u5_mult_78_ab_8__1_), .B(
        u5_mult_78_CARRYB_7__1_), .CI(u5_mult_78_SUMB_7__2_), .CO(
        u5_mult_78_CARRYB_8__1_), .S(u5_mult_78_SUMB_8__1_) );
  FA_X1 u5_mult_78_S1_8_0 ( .A(u5_mult_78_ab_8__0_), .B(
        u5_mult_78_CARRYB_7__0_), .CI(u5_mult_78_SUMB_7__1_), .CO(
        u5_mult_78_CARRYB_8__0_), .S(u5_N8) );
  FA_X1 u5_mult_78_S3_9_9 ( .A(u5_mult_78_ab_9__9_), .B(
        u5_mult_78_CARRYB_8__9_), .CI(u5_mult_78_ab_8__10_), .CO(
        u5_mult_78_CARRYB_9__9_), .S(u5_mult_78_SUMB_9__9_) );
  FA_X1 u5_mult_78_S2_9_8 ( .A(u5_mult_78_ab_9__8_), .B(
        u5_mult_78_CARRYB_8__8_), .CI(u5_mult_78_SUMB_8__9_), .CO(
        u5_mult_78_CARRYB_9__8_), .S(u5_mult_78_SUMB_9__8_) );
  FA_X1 u5_mult_78_S2_9_7 ( .A(u5_mult_78_ab_9__7_), .B(
        u5_mult_78_CARRYB_8__7_), .CI(u5_mult_78_SUMB_8__8_), .CO(
        u5_mult_78_CARRYB_9__7_), .S(u5_mult_78_SUMB_9__7_) );
  FA_X1 u5_mult_78_S2_9_6 ( .A(u5_mult_78_ab_9__6_), .B(
        u5_mult_78_CARRYB_8__6_), .CI(u5_mult_78_SUMB_8__7_), .CO(
        u5_mult_78_CARRYB_9__6_), .S(u5_mult_78_SUMB_9__6_) );
  FA_X1 u5_mult_78_S2_9_5 ( .A(u5_mult_78_ab_9__5_), .B(
        u5_mult_78_CARRYB_8__5_), .CI(u5_mult_78_SUMB_8__6_), .CO(
        u5_mult_78_CARRYB_9__5_), .S(u5_mult_78_SUMB_9__5_) );
  FA_X1 u5_mult_78_S2_9_4 ( .A(u5_mult_78_ab_9__4_), .B(
        u5_mult_78_CARRYB_8__4_), .CI(u5_mult_78_SUMB_8__5_), .CO(
        u5_mult_78_CARRYB_9__4_), .S(u5_mult_78_SUMB_9__4_) );
  FA_X1 u5_mult_78_S2_9_3 ( .A(u5_mult_78_ab_9__3_), .B(
        u5_mult_78_CARRYB_8__3_), .CI(u5_mult_78_SUMB_8__4_), .CO(
        u5_mult_78_CARRYB_9__3_), .S(u5_mult_78_SUMB_9__3_) );
  FA_X1 u5_mult_78_S2_9_2 ( .A(u5_mult_78_ab_9__2_), .B(
        u5_mult_78_CARRYB_8__2_), .CI(u5_mult_78_SUMB_8__3_), .CO(
        u5_mult_78_CARRYB_9__2_), .S(u5_mult_78_SUMB_9__2_) );
  FA_X1 u5_mult_78_S2_9_1 ( .A(u5_mult_78_ab_9__1_), .B(
        u5_mult_78_CARRYB_8__1_), .CI(u5_mult_78_SUMB_8__2_), .CO(
        u5_mult_78_CARRYB_9__1_), .S(u5_mult_78_SUMB_9__1_) );
  FA_X1 u5_mult_78_S1_9_0 ( .A(u5_mult_78_ab_9__0_), .B(
        u5_mult_78_CARRYB_8__0_), .CI(u5_mult_78_SUMB_8__1_), .CO(
        u5_mult_78_CARRYB_9__0_), .S(u5_N9) );
  FA_X1 u5_mult_78_S5_9 ( .A(u5_mult_78_ab_10__9_), .B(u5_mult_78_CARRYB_9__9_), .CI(u5_mult_78_ab_9__10_), .CO(u5_mult_78_CARRYB_10__9_), .S(
        u5_mult_78_SUMB_10__9_) );
  FA_X1 u5_mult_78_S4_8 ( .A(u5_mult_78_ab_10__8_), .B(u5_mult_78_CARRYB_9__8_), .CI(u5_mult_78_SUMB_9__9_), .CO(u5_mult_78_CARRYB_10__8_), .S(
        u5_mult_78_SUMB_10__8_) );
  FA_X1 u5_mult_78_S4_7 ( .A(u5_mult_78_ab_10__7_), .B(u5_mult_78_CARRYB_9__7_), .CI(u5_mult_78_SUMB_9__8_), .CO(u5_mult_78_CARRYB_10__7_), .S(
        u5_mult_78_SUMB_10__7_) );
  FA_X1 u5_mult_78_S4_6 ( .A(u5_mult_78_ab_10__6_), .B(u5_mult_78_CARRYB_9__6_), .CI(u5_mult_78_SUMB_9__7_), .CO(u5_mult_78_CARRYB_10__6_), .S(
        u5_mult_78_SUMB_10__6_) );
  FA_X1 u5_mult_78_S4_5 ( .A(u5_mult_78_ab_10__5_), .B(u5_mult_78_CARRYB_9__5_), .CI(u5_mult_78_SUMB_9__6_), .CO(u5_mult_78_CARRYB_10__5_), .S(
        u5_mult_78_SUMB_10__5_) );
  FA_X1 u5_mult_78_S4_4 ( .A(u5_mult_78_ab_10__4_), .B(u5_mult_78_CARRYB_9__4_), .CI(u5_mult_78_SUMB_9__5_), .CO(u5_mult_78_CARRYB_10__4_), .S(
        u5_mult_78_SUMB_10__4_) );
  FA_X1 u5_mult_78_S4_3 ( .A(u5_mult_78_ab_10__3_), .B(u5_mult_78_CARRYB_9__3_), .CI(u5_mult_78_SUMB_9__4_), .CO(u5_mult_78_CARRYB_10__3_), .S(
        u5_mult_78_SUMB_10__3_) );
  FA_X1 u5_mult_78_S4_2 ( .A(u5_mult_78_ab_10__2_), .B(u5_mult_78_CARRYB_9__2_), .CI(u5_mult_78_SUMB_9__3_), .CO(u5_mult_78_CARRYB_10__2_), .S(
        u5_mult_78_SUMB_10__2_) );
  FA_X1 u5_mult_78_S4_1 ( .A(u5_mult_78_ab_10__1_), .B(u5_mult_78_CARRYB_9__1_), .CI(u5_mult_78_SUMB_9__2_), .CO(u5_mult_78_CARRYB_10__1_), .S(
        u5_mult_78_SUMB_10__1_) );
  FA_X1 u5_mult_78_S4_0 ( .A(u5_mult_78_ab_10__0_), .B(u5_mult_78_CARRYB_9__0_), .CI(u5_mult_78_SUMB_9__1_), .CO(u5_mult_78_CARRYB_10__0_), .S(u5_N10) );
  NAND2_X1 u5_mult_78_FS_1_U54 ( .A1(u5_mult_78_n40), .A2(u5_mult_78_n17), 
        .ZN(u5_mult_78_FS_1_n44) );
  AND2_X1 u5_mult_78_FS_1_U53 ( .A1(u5_mult_78_n35), .A2(u5_mult_78_n16), .ZN(
        u5_mult_78_FS_1_n41) );
  NOR2_X1 u5_mult_78_FS_1_U52 ( .A1(u5_mult_78_n35), .A2(u5_mult_78_n16), .ZN(
        u5_mult_78_FS_1_n42) );
  NOR2_X1 u5_mult_78_FS_1_U51 ( .A1(u5_mult_78_FS_1_n41), .A2(
        u5_mult_78_FS_1_n42), .ZN(u5_mult_78_FS_1_n43) );
  XOR2_X1 u5_mult_78_FS_1_U50 ( .A(u5_mult_78_FS_1_n11), .B(
        u5_mult_78_FS_1_n43), .Z(u5_N13) );
  NOR2_X1 u5_mult_78_FS_1_U49 ( .A1(u5_mult_78_n39), .A2(u5_mult_78_n20), .ZN(
        u5_mult_78_FS_1_n37) );
  NAND2_X1 u5_mult_78_FS_1_U48 ( .A1(u5_mult_78_n39), .A2(u5_mult_78_n20), 
        .ZN(u5_mult_78_FS_1_n39) );
  NAND2_X1 u5_mult_78_FS_1_U47 ( .A1(u5_mult_78_FS_1_n9), .A2(
        u5_mult_78_FS_1_n39), .ZN(u5_mult_78_FS_1_n40) );
  AOI21_X1 u5_mult_78_FS_1_U46 ( .B1(u5_mult_78_FS_1_n10), .B2(
        u5_mult_78_FS_1_n11), .A(u5_mult_78_FS_1_n41), .ZN(u5_mult_78_FS_1_n38) );
  XOR2_X1 u5_mult_78_FS_1_U45 ( .A(u5_mult_78_FS_1_n40), .B(
        u5_mult_78_FS_1_n38), .Z(u5_N14) );
  OAI21_X1 u5_mult_78_FS_1_U44 ( .B1(u5_mult_78_FS_1_n37), .B2(
        u5_mult_78_FS_1_n38), .A(u5_mult_78_FS_1_n39), .ZN(u5_mult_78_FS_1_n33) );
  AND2_X1 u5_mult_78_FS_1_U43 ( .A1(u5_mult_78_n34), .A2(u5_mult_78_n15), .ZN(
        u5_mult_78_FS_1_n34) );
  NOR2_X1 u5_mult_78_FS_1_U42 ( .A1(u5_mult_78_n34), .A2(u5_mult_78_n15), .ZN(
        u5_mult_78_FS_1_n35) );
  NOR2_X1 u5_mult_78_FS_1_U41 ( .A1(u5_mult_78_FS_1_n34), .A2(
        u5_mult_78_FS_1_n35), .ZN(u5_mult_78_FS_1_n36) );
  XOR2_X1 u5_mult_78_FS_1_U40 ( .A(u5_mult_78_FS_1_n33), .B(
        u5_mult_78_FS_1_n36), .Z(u5_N15) );
  NOR2_X1 u5_mult_78_FS_1_U39 ( .A1(u5_mult_78_n38), .A2(u5_mult_78_n19), .ZN(
        u5_mult_78_FS_1_n29) );
  NAND2_X1 u5_mult_78_FS_1_U38 ( .A1(u5_mult_78_n38), .A2(u5_mult_78_n19), 
        .ZN(u5_mult_78_FS_1_n31) );
  NAND2_X1 u5_mult_78_FS_1_U37 ( .A1(u5_mult_78_FS_1_n7), .A2(
        u5_mult_78_FS_1_n31), .ZN(u5_mult_78_FS_1_n32) );
  AOI21_X1 u5_mult_78_FS_1_U36 ( .B1(u5_mult_78_FS_1_n8), .B2(
        u5_mult_78_FS_1_n33), .A(u5_mult_78_FS_1_n34), .ZN(u5_mult_78_FS_1_n30) );
  XOR2_X1 u5_mult_78_FS_1_U35 ( .A(u5_mult_78_FS_1_n32), .B(
        u5_mult_78_FS_1_n30), .Z(u5_N16) );
  OAI21_X1 u5_mult_78_FS_1_U34 ( .B1(u5_mult_78_FS_1_n29), .B2(
        u5_mult_78_FS_1_n30), .A(u5_mult_78_FS_1_n31), .ZN(u5_mult_78_FS_1_n25) );
  AND2_X1 u5_mult_78_FS_1_U33 ( .A1(u5_mult_78_n33), .A2(u5_mult_78_n14), .ZN(
        u5_mult_78_FS_1_n26) );
  NOR2_X1 u5_mult_78_FS_1_U32 ( .A1(u5_mult_78_n33), .A2(u5_mult_78_n14), .ZN(
        u5_mult_78_FS_1_n27) );
  NOR2_X1 u5_mult_78_FS_1_U31 ( .A1(u5_mult_78_FS_1_n26), .A2(
        u5_mult_78_FS_1_n27), .ZN(u5_mult_78_FS_1_n28) );
  XOR2_X1 u5_mult_78_FS_1_U30 ( .A(u5_mult_78_FS_1_n25), .B(
        u5_mult_78_FS_1_n28), .Z(u5_N17) );
  NOR2_X1 u5_mult_78_FS_1_U29 ( .A1(u5_mult_78_n37), .A2(u5_mult_78_n18), .ZN(
        u5_mult_78_FS_1_n21) );
  NAND2_X1 u5_mult_78_FS_1_U28 ( .A1(u5_mult_78_n37), .A2(u5_mult_78_n18), 
        .ZN(u5_mult_78_FS_1_n23) );
  NAND2_X1 u5_mult_78_FS_1_U27 ( .A1(u5_mult_78_FS_1_n5), .A2(
        u5_mult_78_FS_1_n23), .ZN(u5_mult_78_FS_1_n24) );
  AOI21_X1 u5_mult_78_FS_1_U26 ( .B1(u5_mult_78_FS_1_n6), .B2(
        u5_mult_78_FS_1_n25), .A(u5_mult_78_FS_1_n26), .ZN(u5_mult_78_FS_1_n22) );
  XOR2_X1 u5_mult_78_FS_1_U25 ( .A(u5_mult_78_FS_1_n24), .B(
        u5_mult_78_FS_1_n22), .Z(u5_N18) );
  OAI21_X1 u5_mult_78_FS_1_U24 ( .B1(u5_mult_78_FS_1_n21), .B2(
        u5_mult_78_FS_1_n22), .A(u5_mult_78_FS_1_n23), .ZN(u5_mult_78_FS_1_n17) );
  AND2_X1 u5_mult_78_FS_1_U23 ( .A1(u5_mult_78_n32), .A2(u5_mult_78_n13), .ZN(
        u5_mult_78_FS_1_n18) );
  NOR2_X1 u5_mult_78_FS_1_U22 ( .A1(u5_mult_78_n32), .A2(u5_mult_78_n13), .ZN(
        u5_mult_78_FS_1_n19) );
  NOR2_X1 u5_mult_78_FS_1_U21 ( .A1(u5_mult_78_FS_1_n18), .A2(
        u5_mult_78_FS_1_n19), .ZN(u5_mult_78_FS_1_n20) );
  XOR2_X1 u5_mult_78_FS_1_U20 ( .A(u5_mult_78_FS_1_n17), .B(
        u5_mult_78_FS_1_n20), .Z(u5_N19) );
  NOR2_X1 u5_mult_78_FS_1_U19 ( .A1(u5_mult_78_n36), .A2(u5_mult_78_n12), .ZN(
        u5_mult_78_FS_1_n13) );
  NAND2_X1 u5_mult_78_FS_1_U18 ( .A1(u5_mult_78_n36), .A2(u5_mult_78_n12), 
        .ZN(u5_mult_78_FS_1_n15) );
  NAND2_X1 u5_mult_78_FS_1_U17 ( .A1(u5_mult_78_FS_1_n3), .A2(
        u5_mult_78_FS_1_n15), .ZN(u5_mult_78_FS_1_n16) );
  AOI21_X1 u5_mult_78_FS_1_U16 ( .B1(u5_mult_78_FS_1_n4), .B2(
        u5_mult_78_FS_1_n17), .A(u5_mult_78_FS_1_n18), .ZN(u5_mult_78_FS_1_n14) );
  XOR2_X1 u5_mult_78_FS_1_U15 ( .A(u5_mult_78_FS_1_n16), .B(
        u5_mult_78_FS_1_n14), .Z(u5_N20) );
  OAI21_X1 u5_mult_78_FS_1_U14 ( .B1(u5_mult_78_FS_1_n13), .B2(
        u5_mult_78_FS_1_n14), .A(u5_mult_78_FS_1_n15), .ZN(u5_mult_78_FS_1_n12) );
  XOR2_X1 u5_mult_78_FS_1_U13 ( .A(u5_mult_78_FS_1_n12), .B(u5_mult_78_n31), 
        .Z(u5_N21) );
  INV_X4 u5_mult_78_FS_1_U12 ( .A(u5_mult_78_FS_1_n44), .ZN(
        u5_mult_78_FS_1_n11) );
  INV_X4 u5_mult_78_FS_1_U11 ( .A(u5_mult_78_FS_1_n42), .ZN(
        u5_mult_78_FS_1_n10) );
  INV_X4 u5_mult_78_FS_1_U10 ( .A(u5_mult_78_FS_1_n37), .ZN(u5_mult_78_FS_1_n9) );
  INV_X4 u5_mult_78_FS_1_U9 ( .A(u5_mult_78_FS_1_n35), .ZN(u5_mult_78_FS_1_n8)
         );
  INV_X4 u5_mult_78_FS_1_U8 ( .A(u5_mult_78_FS_1_n29), .ZN(u5_mult_78_FS_1_n7)
         );
  INV_X4 u5_mult_78_FS_1_U7 ( .A(u5_mult_78_FS_1_n27), .ZN(u5_mult_78_FS_1_n6)
         );
  INV_X4 u5_mult_78_FS_1_U6 ( .A(u5_mult_78_FS_1_n21), .ZN(u5_mult_78_FS_1_n5)
         );
  INV_X4 u5_mult_78_FS_1_U5 ( .A(u5_mult_78_FS_1_n19), .ZN(u5_mult_78_FS_1_n4)
         );
  INV_X4 u5_mult_78_FS_1_U4 ( .A(u5_mult_78_FS_1_n13), .ZN(u5_mult_78_FS_1_n3)
         );
  AND2_X4 u5_mult_78_FS_1_U3 ( .A1(u5_mult_78_FS_1_n1), .A2(
        u5_mult_78_FS_1_n44), .ZN(u5_N12) );
  OR2_X4 u5_mult_78_FS_1_U2 ( .A1(u5_mult_78_n40), .A2(u5_mult_78_n17), .ZN(
        u5_mult_78_FS_1_n1) );
endmodule

