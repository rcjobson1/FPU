
module fpu ( clk, rmode, fpu_op, opa, opb, out, inf, snan, qnan, ine, overflow, 
        underflow, zero, div_by_zero );
  input [1:0] rmode;
  input [2:0] fpu_op;
  input [31:0] opa;
  input [31:0] opb;
  output [31:0] out;
  input clk;
  output inf, snan, qnan, ine, overflow, underflow, zero, div_by_zero;
  wire   fpu_op_r3_1_, inf_d, ind_d, snan_d, opa_nan, opb_nan, opa_00, opb_00,
         opa_inf, opb_inf, opa_dn, sign_fasu, result_zero_sign_d, sign_fasu_r,
         sign_mul, sign_exe, inf_mul, sign_mul_r, sign_exe_r, exp_ovf_r_0_,
         N107, N141, N170, N172, N173, N174, N175, N176, N177, N178, N179,
         N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190,
         N191, N192, N193, N194, N195, N214, N215, N216, N217, N218, N219,
         N220, N221, N224, N227, N228, N229, N230, N231, N232, N233, N234,
         N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245,
         N246, N247, N248, N249, N250, N251, N298, N299, N300, N301, N302,
         N303, N304, N305, N306, N307, N308, N309, N310, N311, N312, N313,
         N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324,
         N325, N391, N392, N393, N394, N395, N396, N397, N398, N399, N400,
         N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, N411,
         N412, N413, N414, N415, N416, N417, N418, N419, N420, N421, opas_r1,
         opas_r2, sign, N441, fasu_op_r1, N445, N446, N447, N448, N449, N450,
         N451, N452, N453, N454, N455, N456, N457, N458, N459, N460, N461,
         N462, N463, N464, N465, N466, N467, N468, N469, N470, N471, N473,
         N475, N495, N509, N519, N522, N524, N526, N531, N532, opa_nan_r, N533,
         N540, u0_N17, u0_N16, u0_fractb_00, u0_fracta_00, u0_expb_00,
         u0_expa_00, u0_N11, u0_N10, u0_N7, u0_N6, u0_snan_r_b, u0_N5,
         u0_qnan_r_b, u0_snan_r_a, u0_N4, u0_qnan_r_a, u0_infb_f_r,
         u0_infa_f_r, u0_expb_ff, u0_expa_ff, u1_N140, u1_fracta_eq_fractb,
         u1_N131, u1_fracta_lt_fractb, u1_N130, u1_N129, u1_add_r, u1_signa_r,
         u1_sign_d, u1_adj_op_out_sft_0_, u1_adj_op_out_sft_1_,
         u1_adj_op_out_sft_2_, u1_adj_op_out_sft_3_, u1_adj_op_out_sft_4_,
         u1_adj_op_out_sft_5_, u1_adj_op_out_sft_6_, u1_adj_op_out_sft_7_,
         u1_adj_op_out_sft_8_, u1_adj_op_out_sft_9_, u1_adj_op_out_sft_10_,
         u1_adj_op_out_sft_11_, u1_adj_op_out_sft_12_, u1_adj_op_out_sft_13_,
         u1_adj_op_out_sft_14_, u1_adj_op_out_sft_15_, u1_adj_op_out_sft_16_,
         u1_adj_op_out_sft_17_, u1_adj_op_out_sft_18_, u1_adj_op_out_sft_19_,
         u1_adj_op_out_sft_20_, u1_adj_op_out_sft_21_, u1_adj_op_out_sft_22_,
         u1_adj_op_out_sft_23_, u1_adj_op_out_sft_24_, u1_adj_op_out_sft_25_,
         u1_adj_op_out_sft_26_, u1_exp_diff_sft_4_, u1_adj_op_10_,
         u1_adj_op_17_, u1_adj_op_18_, u1_adj_op_19_, u1_adj_op_20_,
         u1_adj_op_22_, u1_N44, u1_N43, u1_N42, u1_N41, u1_N40, u1_N39, u1_N38,
         u1_N37, u2_N124, u2_N97, u2_sign_d, u2_N90, u2_exp_ovf_d_0_,
         u2_exp_ovf_d_1_, u2_N65, u2_N64, u2_N63, u2_N62, u2_N61, u2_N60,
         u2_N59, u2_N58, u2_N49, u2_N48, u2_N47, u2_N46, u2_N45, u2_N44,
         u2_N43, u2_N42, u2_exp_tmp4_0_, u2_exp_tmp4_1_, u2_exp_tmp4_2_,
         u2_exp_tmp4_3_, u2_exp_tmp4_4_, u2_exp_tmp4_5_, u2_exp_tmp4_6_,
         u2_exp_tmp4_7_, u2_exp_tmp3_0_, u2_exp_tmp3_1_, u2_exp_tmp3_2_,
         u2_exp_tmp3_3_, u2_exp_tmp3_4_, u2_exp_tmp3_5_, u2_exp_tmp3_6_,
         u2_exp_tmp3_7_, u2_N23, u2_N22, u2_N21, u2_N20, u2_N19, u2_N18,
         u2_N17, u2_N16, u2_N15, u2_N14, u2_N13, u2_N12, u2_N11, u2_N10, u2_N9,
         u2_N8, u2_N7, u2_N6, u3_N58, u3_N57, u3_N56, u3_N55, u3_N54, u3_N53,
         u3_N52, u3_N51, u3_N50, u3_N49, u3_N48, u3_N47, u3_N46, u3_N45,
         u3_N44, u3_N43, u3_N42, u3_N41, u3_N40, u3_N39, u3_N38, u3_N37,
         u3_N36, u3_N35, u3_N34, u3_N33, u3_N32, u3_N31, u3_N30, u3_N29,
         u3_N28, u3_N27, u3_N26, u3_N25, u3_N24, u3_N23, u3_N22, u3_N21,
         u3_N20, u3_N19, u3_N18, u3_N17, u3_N16, u3_N15, u3_N14, u3_N13,
         u3_N12, u3_N11, u3_N10, u3_N9, u3_N8, u3_N7, u3_N6, u3_N5, u3_N4,
         u3_N3, u5_N47, u5_N46, u5_N45, u5_N44, u5_N43, u5_N42, u5_N41, u5_N40,
         u5_N39, u5_N38, u5_N37, u5_N36, u5_N35, u5_N34, u5_N33, u5_N32,
         u5_N31, u5_N30, u5_N29, u5_N28, u5_N27, u5_N26, u5_N25, u5_N24,
         u5_N23, u5_N22, u5_N21, u5_N20, u5_N19, u5_N18, u5_N17, u5_N16,
         u5_N15, u5_N14, u5_N13, u5_N12, u5_N11, u5_N10, u5_N9, u5_N8, u5_N7,
         u5_N6, u5_N5, u5_N4, u5_N3, u5_N2, u5_N1, u5_N0, u6_N49, u6_N48,
         u6_N47, u6_N46, u6_N45, u6_N44, u6_N43, u6_N42, u6_N41, u6_N40,
         u6_N39, u6_N38, u6_N37, u6_N36, u6_N35, u6_N34, u6_N33, u6_N32,
         u6_N31, u6_N30, u6_N29, u6_N28, u6_N27, u6_N26, u6_N23, u6_N22,
         u6_N18, u6_N17, u6_N15, u6_N13, u6_N10, u6_N9, u6_N8, u6_N7, u6_N6,
         u6_N5, u6_N4, u6_N3, u6_N2, u6_N1, u6_N0, u4_N1977, u4_N1733,
         u4_N1600, u4_N1598, u4_div_exp2_0_, u4_div_exp2_1_, u4_div_exp2_2_,
         u4_div_exp2_3_, u4_div_exp2_4_, u4_div_exp2_5_, u4_div_exp2_6_,
         u4_div_exp2_7_, u4_div_exp1_0_, u4_div_exp1_1_, u4_div_exp1_2_,
         u4_div_exp1_3_, u4_div_exp1_4_, u4_div_exp1_5_, u4_div_exp1_6_,
         u4_div_exp1_7_, u4_div_exp1_8_, u4_fi_ldz_2a_3_, u4_fi_ldz_2a_4_,
         u4_fi_ldz_2a_5_, u4_fi_ldz_2a_6_, u4_ldz_all_0_, u4_ldz_all_1_,
         u4_ldz_all_2_, u4_ldz_all_3_, u4_ldz_all_5_, u4_ldz_all_6_,
         u4_exp_out_pl1_0_, u4_exp_out_pl1_1_, u4_exp_out_pl1_2_,
         u4_exp_out_pl1_3_, u4_exp_out_pl1_4_, u4_exp_out_pl1_5_,
         u4_exp_out_pl1_6_, u4_exp_out_pl1_7_, u4_fi_ldz_mi1_1_,
         u4_fi_ldz_mi1_2_, u4_fi_ldz_mi1_3_, u4_fi_ldz_mi1_4_,
         u4_fi_ldz_mi1_5_, u4_N1455, u4_N1454, u4_N1453, u4_N1452, u4_N1451,
         u4_N1450, u4_N1449, u4_N1448, u4_N1447, u4_N1446, u4_N1445, u4_N1444,
         u4_N1443, u4_N1442, u4_N1441, u4_N1440, u4_N1439, u4_N1438, u4_N1437,
         u4_N1436, u4_N1435, u4_N1434, u4_N1433, u4_N1432, u4_N1431, u4_N1430,
         u4_N1429, u4_N1428, u4_N1427, u4_N1426, u4_N1425, u4_N1424, u4_N1423,
         u4_N1422, u4_N1421, u4_N1420, u4_N1419, u4_N1418, u4_N1417, u4_N1416,
         u4_N1415, u4_N1414, u4_N1413, u4_N1412, u4_N1411, u4_N1410, u4_N1409,
         u4_N1408, u4_N1405, u4_N1404, u4_N1403, u4_N1402, u4_N1401, u4_N1400,
         u4_N1399, u4_N1398, u4_N1397, u4_N1396, u4_N1395, u4_N1394, u4_N1393,
         u4_N1392, u4_N1391, u4_N1390, u4_N1389, u4_N1388, u4_N1387, u4_N1386,
         u4_N1385, u4_N1384, u4_N1383, u4_N1382, u4_N1381, u4_N1380, u4_N1379,
         u4_N1378, u4_N1377, u4_N1376, u4_N1375, u4_N1374, u4_N1373, u4_N1372,
         u4_N1371, u4_N1370, u4_N1369, u4_N1368, u4_N1367, u4_N1366, u4_N1365,
         u4_N1364, u4_N1363, u4_N1362, u4_N1361, u4_N1360, u4_N1359, u4_N1358,
         u4_exp_in_pl1_0_, u4_exp_in_pl1_1_, u4_exp_in_pl1_2_,
         u4_exp_in_pl1_3_, u4_exp_in_pl1_4_, u4_exp_in_pl1_5_,
         u4_exp_in_pl1_6_, u4_exp_in_pl1_7_, u4_exp_in_pl1_8_, u4_f2i_shft_2_,
         u4_f2i_shft_3_, u4_f2i_shft_4_, u4_f2i_shft_5_, u4_f2i_shft_6_,
         u4_f2i_shft_7_, u4_div_shft3_0_, u4_div_shft3_1_, u4_div_shft3_2_,
         u4_div_shft3_3_, u4_div_shft3_4_, u4_div_shft3_5_, u4_div_shft3_6_,
         u4_div_shft3_7_, u4_exp_in_mi1_1_, u4_exp_in_mi1_2_, u4_exp_in_mi1_4_,
         u4_exp_in_mi1_5_, u4_exp_in_mi1_6_, u4_exp_in_mi1_7_,
         u4_fract_out_pl1_0_, u4_fract_out_pl1_1_, u4_fract_out_pl1_2_,
         u4_fract_out_pl1_3_, u4_fract_out_pl1_4_, u4_fract_out_pl1_5_,
         u4_fract_out_pl1_6_, u4_fract_out_pl1_7_, u4_fract_out_pl1_8_,
         u4_fract_out_pl1_9_, u4_fract_out_pl1_10_, u4_fract_out_pl1_11_,
         u4_fract_out_pl1_12_, u4_fract_out_pl1_13_, u4_fract_out_pl1_14_,
         u4_fract_out_pl1_15_, u4_fract_out_pl1_16_, u4_fract_out_pl1_17_,
         u4_fract_out_pl1_18_, u4_fract_out_pl1_19_, u4_fract_out_pl1_20_,
         u4_fract_out_pl1_21_, u4_fract_out_pl1_22_, u4_fract_out_pl1_23_,
         u4_exp_next_mi_0_, u4_exp_next_mi_1_, u4_exp_next_mi_2_,
         u4_exp_next_mi_3_, u4_exp_next_mi_4_, u4_exp_next_mi_5_,
         u4_exp_next_mi_6_, u4_exp_next_mi_7_, u4_exp_next_mi_8_,
         u4_fract_out_0_, u4_fract_out_1_, u4_fract_out_2_, u4_fract_out_3_,
         u4_fract_out_4_, u4_fract_out_5_, u4_fract_out_6_, u4_fract_out_7_,
         u4_fract_out_8_, u4_fract_out_9_, u4_fract_out_10_, u4_fract_out_11_,
         u4_fract_out_12_, u4_fract_out_13_, u4_fract_out_14_,
         u4_fract_out_15_, u4_fract_out_16_, u4_fract_out_17_,
         u4_fract_out_18_, u4_fract_out_19_, u4_fract_out_20_,
         u4_fract_out_21_, u4_fract_out_22_, u4_exp_out_1_, u4_exp_out_2_,
         u4_exp_out_4_, u4_exp_out_6_, n1371, n1373, n1416, n1451, n1452,
         n1453, n1454, n1456, n1457, n1458, n1459, n1460, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1735,
         n1742, n1743, n1744, n1745, n1746, n1749, n1751, n1752, n1753, n1754,
         n1756, n1821, n1822, n1823, n1889, n1890, n1892, n1893, n1895, n1896,
         n1898, n1900, n1901, n1903, n2051, n2058, n2060, n2065, n2069, n2076,
         n2083, n2087, n2091, n2093, n2245, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2278, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2437, n2443, n2444, n2445, n2448,
         n2449, n2450, n2451, n2452, n2453, n2459, u4_ldz_dif_7_,
         u4_ldz_dif_6_, u4_ldz_dif_5_, u4_ldz_dif_4_, u4_ldz_dif_3_,
         u4_ldz_dif_2_, u4_ldz_dif_1_, u4_ldz_dif_0_, net17652, net17653,
         net17654, net17655, net17656, net17657, net17659, net17682, net17683,
         net17684, net17685, net17686, net17690, net17692, net17693, net17694,
         net17695, net22501, net23043, net23097, net23104, net23180, net23182,
         net28939, net33106, net48876, net82010, net82011, net82013, net82014,
         net82023, net82024, net82029, net82030, net82034, net82035, net82036,
         net82039, net82040, net82753, net82757, net82762, net82764, net82767,
         net82776, net82778, net82781, net82782, net82784, net82792, net82807,
         net82826, net82829, net82850, net82853, net82856, net82873, net82876,
         net82891, net82893, net82902, net82911, net82918, net82925, net82927,
         net82929, net82931, net82932, net82934, net82938, net82940, net82950,
         net82951, net82952, net82957, net82965, net82988, net82991, net82997,
         net83007, net83009, net83016, net83017, net83018, net83019, net83020,
         net83030, net83036, net83041, net83042, net83044, net83045, net83057,
         net83059, net83061, net83064, net83066, net83068, net83070, net83074,
         net83090, net83109, net83113, net83115, net83119, net83120, net83126,
         net83168, net83197, net83198, net83214, net83220, net83233, net83234,
         net83247, net83248, net83254, net83262, net83263, net83264, net83271,
         net83274, net83275, net83276, net83278, net83279, net83282, net83288,
         net83292, net83294, net83295, net83297, net83300, net83305, net83312,
         net83316, net83326, net83327, net83328, net83329, net83338, net83342,
         net83344, net83348, net83349, net83350, net83356, net83357, net83358,
         net83359, net83367, net83368, net83369, net83370, net83371, net83373,
         net83375, net83381, net83383, net83384, net83385, net83393, net83396,
         net83404, net83408, net83409, net83415, net83416, net83417, net83422,
         net83428, net83430, net83431, net83433, net83434, net83435, net83446,
         net83463, net83468, net83474, net83487, net83492, net83495, net83497,
         net83498, net83499, net83500, net83507, net83510, net83514, net83518,
         net83525, net83526, net83527, net83532, net83534, net83535, net83555,
         net83556, net83562, net83563, net83565, net83567, net83568, net83569,
         net83579, net83580, net83591, net83593, net83596, net83599, net83606,
         net83616, net83620, net83621, net83622, net83624, net83630, net83632,
         net83633, net83634, net83636, net83638, net83642, net83660, net83713,
         net83714, net83715, net83721, net83724, net83725, net83727, net83735,
         net83736, net83738, net83744, net83745, net83747, net83749, net83750,
         net83751, net83752, net83753, net83754, net83756, net83757, net83759,
         net83761, net83762, net83766, net83767, net83770, net83771, net83773,
         net83775, net83776, net83791, net83796, net83797, net83799, net83807,
         net83811, net83823, net83824, net83828, net83836, net83837, net83841,
         net83842, net83846, net83851, net83854, net83857, net83858, net83862,
         net83863, net83864, net83865, net83868, net83869, net83870, net83878,
         net83886, net83887, net83888, net83902, net83903, net83918, net83919,
         net83921, net83924, net83925, net83926, net83927, net83928, net83932,
         net83933, net83941, net83943, net83948, net83953, net83957, net83959,
         net83963, net83965, net83971, net83977, net83991, net83995, net84000,
         net84002, net84003, net84013, net84014, net84015, net84016, net84018,
         net84030, net84032, net84035, net84043, net84054, net84067, net84075,
         net84083, net84091, net84092, net84100, net84101, net84115, net84116,
         net84117, net84121, net84124, net84128, net84131, net84132, net84135,
         net84138, net84139, net84140, net84141, net84142, net84143, net84149,
         net84150, net84151, net84158, net84166, net84167, net84172, net84178,
         net84181, net84182, net84183, net84185, net84188, net84189, net84191,
         net84201, net84204, net84205, net84207, net84224, net84225, net84231,
         net84237, net84238, net84242, net84257, net84261, net84262, net84272,
         net84273, net84275, net84284, net84285, net84286, net84293, net84298,
         net84301, net84302, net84306, net84311, net84312, net84314, net84321,
         net84323, net84324, net84341, net84343, net84345, net84347, net84348,
         net84349, net84350, net84351, net84353, net84355, net84363, net84364,
         net84370, net84375, net84376, net84377, net84382, net84385, net84387,
         net84396, net84397, net84400, net84411, net84435, net84436, net84443,
         net84444, net84450, net84455, net84490, net84496, net84557, net84559,
         net84568, net84605, net84736, net84737, net84738, net85121, net85117,
         net85115, net85111, net85145, net85143, net85139, net85135, net85133,
         net85131, net85149, net85167, net85165, net85159, net85157, net85179,
         net85175, net85377, net85393, net85391, net85901, net85905, net85929,
         net85933, net85932, net85937, net85976, net85975, net85989, net85988,
         net85987, net85986, net85985, net86001, net85999, net85998, net85997,
         net86012, net86015, net86014, net86013, net86028, net86032, net86040,
         net86045, net86236, net86235, net86257, net86295, net86294, net86309,
         net86315, net86401, net86418, net86478, net86486, net86497, net86532,
         net86531, net86571, net90897, net90945, net91297, net91406, net91498,
         net91595, net91594, net91733, net91817, net92015, net92028, net92065,
         net92365, net92392, net92566, net92573, net92599, net92624, net92622,
         net92661, net92690, net92738, net92781, net92895, net93218, net93364,
         net93404, net93422, net93507, net93671, net93695, net93714, net93777,
         net93776, net93902, net93937, net94004, net94019, net94138, net94146,
         net94305, net94374, net94373, net94442, net94516, net94515, net94514,
         net94513, net94566, net94587, net94595, net94614, net94692, net94701,
         net94703, net94725, net94811, net94825, net94834, net94896, net94933,
         net94948, net94966, net94976, net95019, net95070, net95118, net95132,
         net95137, net95136, net95138, net95148, net95173, net95178, net95236,
         net95242, net95279, net95297, net95357, net95365, net95431, net95473,
         net95479, net95504, net95525, net95549, net95574, net95605, net95614,
         net93655, net85177, net84451, net84362, net84361, net84239, net84202,
         net83635, net83625, net82037, net83123, net83121, net83117, net84118,
         net82993, net83043, net83038, net84495, net84271, net84270, net84258,
         net84236, net93455, net85399, net85397, net26607, net95353, net93416,
         net84354, net84305, net84283, net84282, net84280, net84235, net84171,
         net86481, net83343, net84356, net84300, net84281, net83458, net83405,
         net83403, net83402, net86234, net83730, net83723, n2085, net83325,
         net83039, net86496, net83166, n1461, net85990, net83345, net83196,
         net82780, net85928, net84049, net84048, net84046, net84044, net84017,
         net83958, net83445, net83418, net83319, net82012, net83826, net83818,
         net83817, net83816, net83665, net92408, net92066, net85904, net83639,
         net83602, net83601, net83421, net82038, net92626, net86570, net84548,
         net84547, net84546, net84180, net83722, fract_denorm_46_, net84102,
         net84080, net83114, net83052, net82852, u4_N1640, net83444, net83443,
         net83442, net83441, net83440, net83439, net83438, net83437, net83436,
         net83410, net83259, net83667, net83605, net82939, net85183, net84042,
         net83787, net83785, net83778, net83005, net83800, net83731, net82999,
         n1450, u4_exp_out_3_, net84082, net83994, net83993, net83803,
         net83802, net83801, net83726, net83668, net82953, n2067, net95102,
         net93036, net83788, net94620, net86044, net83931, net83930, net83929,
         net83834, net83832, net83831, net83827, net83374, u4_N1976, net83783,
         net83780, net83779, net83777, u4_exp_out_5_, net84079, net84036,
         net83808, net85141, net85119, net84556, u4_N1732, net92816, net92815,
         net91838, net91045, net91044, net90736, net83974, net83973, net83972,
         net83781, net93471, net86027, net85169, net85163, net85125, net84077,
         net84076, net82998, net82916, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2518, n2519, n2520, n2521, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2768, n2769, n2770,
         n2771, n2772, n2773, n2776, n2777, n2779, n2780, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2948, n2949, n2950, n2951, n2952, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3015, n3016, n3017, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, u4_sub_472_n9, u4_sub_472_n8,
         u4_sub_472_n7, u4_sub_472_n6, u4_sub_472_n5, u4_sub_472_n4,
         u4_sub_472_n3, u4_sub_472_n2, u4_sub_472_n1, u4_sub_472_carry_1_,
         u4_sub_472_carry_2_, u4_sub_472_carry_3_, u4_sub_472_carry_4_,
         u4_sub_472_carry_5_, u4_sub_472_carry_6_, u4_sub_472_carry_7_,
         u4_sub_471_n8, u4_sub_471_n7, u4_sub_471_n6, u4_sub_471_n5,
         u4_sub_471_n4, u4_sub_471_n3, u4_sub_471_n2, u4_sub_471_n1,
         u4_sll_453_n267, u4_sll_453_n266, u4_sll_453_n265, u4_sll_453_n264,
         u4_sll_453_n263, u4_sll_453_n262, u4_sll_453_n261, u4_sll_453_n260,
         u4_sll_453_n259, u4_sll_453_n258, u4_sll_453_n257, u4_sll_453_n256,
         u4_sll_453_n255, u4_sll_453_n254, u4_sll_453_n253, u4_sll_453_n252,
         u4_sll_453_n251, u4_sll_453_n250, u4_sll_453_n249, u4_sll_453_n248,
         u4_sll_453_n247, u4_sll_453_n246, u4_sll_453_n245, u4_sll_453_n244,
         u4_sll_453_n243, u4_sll_453_n242, u4_sll_453_n241, u4_sll_453_n240,
         u4_sll_453_n239, u4_sll_453_n238, u4_sll_453_n237, u4_sll_453_n236,
         u4_sll_453_n235, u4_sll_453_n234, u4_sll_453_n233, u4_sll_453_n232,
         u4_sll_453_n231, u4_sll_453_n230, u4_sll_453_n229, u4_sll_453_n228,
         u4_sll_453_n227, u4_sll_453_n226, u4_sll_453_n225, u4_sll_453_n224,
         u4_sll_453_n223, u4_sll_453_n222, u4_sll_453_n221, u4_sll_453_n220,
         u4_sll_453_n219, u4_sll_453_n218, u4_sll_453_n217, u4_sll_453_n216,
         u4_sll_453_n215, u4_sll_453_n214, u4_sll_453_n213, u4_sll_453_n212,
         u4_sll_453_n211, u4_sll_453_n210, u4_sll_453_n209, u4_sll_453_n208,
         u4_sll_453_n207, u4_sll_453_n206, u4_sll_453_n205, u4_sll_453_n204,
         u4_sll_453_n203, u4_sll_453_n202, u4_sll_453_n201, u4_sll_453_n200,
         u4_sll_453_n199, u4_sll_453_n198, u4_sll_453_n197, u4_sll_453_n196,
         u4_sll_453_n195, u4_sll_453_n194, u4_sll_453_n193, u4_sll_453_n192,
         u4_sll_453_n191, u4_sll_453_n190, u4_sll_453_n189, u4_sll_453_n188,
         u4_sll_453_n187, u4_sll_453_n186, u4_sll_453_n185, u4_sll_453_n184,
         u4_sll_453_n183, u4_sll_453_n182, u4_sll_453_n181, u4_sll_453_n180,
         u4_sll_453_n179, u4_sll_453_n178, u4_sll_453_n177, u4_sll_453_n176,
         u4_sll_453_n175, u4_sll_453_n174, u4_sll_453_n173, u4_sll_453_n172,
         u4_sll_453_n171, u4_sll_453_n170, u4_sll_453_n169, u4_sll_453_n168,
         u4_sll_453_n167, u4_sll_453_n166, u4_sll_453_n165, u4_sll_453_n164,
         u4_sll_453_n163, u4_sll_453_n162, u4_sll_453_n161, u4_sll_453_n160,
         u4_sll_453_n159, u4_sll_453_n158, u4_sll_453_n157, u4_sll_453_n156,
         u4_sll_453_n155, u4_sll_453_n154, u4_sll_453_n153, u4_sll_453_n152,
         u4_sll_453_n151, u4_sll_453_n150, u4_sll_453_n149, u4_sll_453_n148,
         u4_sll_453_n147, u4_sll_453_n146, u4_sll_453_n145, u4_sll_453_n144,
         u4_sll_453_n143, u4_sll_453_n142, u4_sll_453_n141, u4_sll_453_n140,
         u4_sll_453_n139, u4_sll_453_n138, u4_sll_453_n137, u4_sll_453_n136,
         u4_sll_453_n135, u4_sll_453_n134, u4_sll_453_n133, u4_sll_453_n132,
         u4_sll_453_n131, u4_sll_453_n130, u4_sll_453_n129, u4_sll_453_n128,
         u4_sll_453_n127, u4_sll_453_n126, u4_sll_453_n125, u4_sll_453_n124,
         u4_sll_453_n123, u4_sll_453_n122, u4_sll_453_n121, u4_sll_453_n120,
         u4_sll_453_n119, u4_sll_453_n118, u4_sll_453_n117, u4_sll_453_n116,
         u4_sll_453_n115, u4_sll_453_n114, u4_sll_453_n113, u4_sll_453_n112,
         u4_sll_453_n111, u4_sll_453_n110, u4_sll_453_n109, u4_sll_453_n108,
         u4_sll_453_n107, u4_sll_453_n106, u4_sll_453_n105, u4_sll_453_n104,
         u4_sll_453_n103, u4_sll_453_n102, u4_sll_453_n101, u4_sll_453_n100,
         u4_sll_453_n99, u4_sll_453_n98, u4_sll_453_n97, u4_sll_453_n96,
         u4_sll_453_n95, u4_sll_453_n94, u4_sll_453_n93, u4_sll_453_n92,
         u4_sll_453_n91, u4_sll_453_n90, u4_sll_453_n89, u4_sll_453_n88,
         u4_sll_453_n87, u4_sll_453_n86, u4_sll_453_n85, u4_sll_453_n84,
         u4_sll_453_n83, u4_sll_453_n82, u4_sll_453_n81, u4_sll_453_n80,
         u4_sll_453_n79, u4_sll_453_n78, u4_sll_453_n77, u4_sll_453_n76,
         u4_sll_453_n75, u4_sll_453_n74, u4_sll_453_n73, u4_sll_453_n72,
         u4_sll_453_n71, u4_sll_453_n70, u4_sll_453_n69, u4_sll_453_n68,
         u4_sll_453_n67, u4_sll_453_n66, u4_sll_453_n65, u4_sll_453_n64,
         u4_sll_453_n63, u4_sll_453_n62, u4_sll_453_n61, u4_sll_453_n60,
         u4_sll_453_n59, u4_sll_453_n58, u4_sll_453_n57, u4_sll_453_n56,
         u4_sll_453_n55, u4_sll_453_n54, u4_sll_453_n53, u4_sll_453_n52,
         u4_sll_453_n51, u4_sll_453_n50, u4_sll_453_n49, u4_sll_453_n48,
         u4_sll_453_n47, u4_sll_453_n46, u4_sll_453_n45, u4_sll_453_n44,
         u4_sll_453_n43, u4_sll_453_n42, u4_sll_453_n41, u4_sll_453_n40,
         u4_sll_453_n39, u4_sll_453_n38, u4_sll_453_n37, u4_sll_453_n36,
         u4_sll_453_n35, u4_sll_453_n34, u4_sll_453_n33, u4_sll_453_n32,
         u4_sll_453_n31, u4_sll_453_n30, u4_sll_453_n29, u4_sll_453_n28,
         u4_sll_453_n27, u4_sll_453_n26, u4_sll_453_n25, u4_sll_453_n24,
         u4_sll_453_n23, u4_sll_453_n22, u4_sll_453_n21, u4_sll_453_n20,
         u4_sll_453_n19, u4_sll_453_n18, u4_sll_453_n17, u4_sll_453_n16,
         u4_sll_453_n15, u4_sll_453_n14, u4_sll_453_n13, u4_sll_453_n12,
         u4_sll_453_n11, u4_sll_453_n10, u4_sll_453_n9, u4_sll_453_n8,
         u4_sll_453_n7, u4_sll_453_n6, u4_sll_453_n5, u4_sll_453_n4,
         u4_sll_453_n3, u4_sll_453_n2, u4_sll_453_n1, u4_sll_453_ML_int_2__30_,
         u4_sll_453_ML_int_3__34_, u4_sll_453_ML_int_4__18_,
         u4_sll_453_ML_int_4__34_, u4_sll_453_ML_int_5__34_,
         u4_sll_453_net85299, u4_sll_453_net85319, u4_sll_453_net85349,
         u4_sll_453_net85351, u4_sll_453_ML_int_1__8_,
         u4_sll_453_ML_int_2__10_, u4_sll_453_net85269, u4_sll_453_net85271,
         u4_sll_453_ML_int_2__6_, u4_sll_453_ML_int_3__10_,
         u4_sll_453_net85267, u4_sll_453_net85275, u4_sll_453_ML_int_5__2_,
         u4_sll_453_net12807, u4_sll_453_net85337, u4_sll_453_net85347,
         u4_sll_453_net85365, u4_sll_453_ML_int_3__18_, u4_sll_453_net95318,
         u4_sll_453_net94330, u4_sll_453_net94297, u4_sll_453_net94228,
         u4_sll_453_net94113, u4_sll_453_net94050, u4_sll_453_net93991,
         u4_sll_453_net93929, u4_sll_453_net93930, u4_sll_453_net93876,
         u4_sll_453_net93857, u4_sll_453_net93725, u4_sll_453_net93728,
         u4_sll_453_net93710, u4_sll_453_net93645, u4_sll_453_net93630,
         u4_sll_453_net93631, u4_sll_453_net93359, u4_sll_453_net93284,
         u4_sll_453_net93219, u4_sll_453_net93122, u4_sll_453_net93041,
         u4_sll_453_net92631, u4_sll_453_net92610, u4_sll_453_net92613,
         u4_sll_453_net91550, u4_sll_453_net86373, u4_sll_453_net86374,
         u4_sll_453_net85353, u4_sll_453_net85355, u4_sll_453_net85333,
         u4_sll_453_net85339, u4_sll_453_net85341, u4_sll_453_net85343,
         u4_sll_453_net85301, u4_sll_453_net85303, u4_sll_453_net85313,
         u4_sll_453_net85315, u4_sll_453_net85321, u4_sll_453_net85273,
         u4_sll_453_net85285, u4_sll_453_net85287, u4_sll_453_net85289,
         u4_sll_453_net85257, u4_sll_453_net85259, u4_sll_453_net85261,
         u4_sll_453_net85263, u4_sll_453_net85265, u4_sll_453_net85229,
         u4_sll_453_net85231, u4_sll_453_net85237, u4_sll_453_ML_int_5__0_,
         u4_sll_453_ML_int_5__1_, u4_sll_453_ML_int_5__3_,
         u4_sll_453_ML_int_5__4_, u4_sll_453_ML_int_5__5_,
         u4_sll_453_ML_int_5__6_, u4_sll_453_ML_int_5__7_,
         u4_sll_453_ML_int_5__8_, u4_sll_453_ML_int_5__9_,
         u4_sll_453_ML_int_5__10_, u4_sll_453_ML_int_5__11_,
         u4_sll_453_ML_int_5__12_, u4_sll_453_ML_int_5__13_,
         u4_sll_453_ML_int_5__14_, u4_sll_453_ML_int_5__15_,
         u4_sll_453_ML_int_5__16_, u4_sll_453_ML_int_5__17_,
         u4_sll_453_ML_int_5__18_, u4_sll_453_ML_int_5__19_,
         u4_sll_453_ML_int_5__20_, u4_sll_453_ML_int_5__21_,
         u4_sll_453_ML_int_5__22_, u4_sll_453_ML_int_5__23_,
         u4_sll_453_ML_int_5__24_, u4_sll_453_ML_int_5__25_,
         u4_sll_453_ML_int_5__26_, u4_sll_453_ML_int_5__27_,
         u4_sll_453_ML_int_5__28_, u4_sll_453_ML_int_5__29_,
         u4_sll_453_ML_int_5__30_, u4_sll_453_ML_int_5__31_,
         u4_sll_453_ML_int_5__32_, u4_sll_453_ML_int_5__33_,
         u4_sll_453_ML_int_5__35_, u4_sll_453_ML_int_5__36_,
         u4_sll_453_ML_int_5__37_, u4_sll_453_ML_int_5__38_,
         u4_sll_453_ML_int_5__39_, u4_sll_453_ML_int_5__40_,
         u4_sll_453_ML_int_5__41_, u4_sll_453_ML_int_5__42_,
         u4_sll_453_ML_int_5__43_, u4_sll_453_ML_int_5__44_,
         u4_sll_453_ML_int_5__45_, u4_sll_453_ML_int_5__46_,
         u4_sll_453_ML_int_5__47_, u4_sll_453_ML_int_4__0_,
         u4_sll_453_ML_int_4__1_, u4_sll_453_ML_int_4__2_,
         u4_sll_453_ML_int_4__3_, u4_sll_453_ML_int_4__4_,
         u4_sll_453_ML_int_4__5_, u4_sll_453_ML_int_4__6_,
         u4_sll_453_ML_int_4__7_, u4_sll_453_ML_int_4__8_,
         u4_sll_453_ML_int_4__9_, u4_sll_453_ML_int_4__10_,
         u4_sll_453_ML_int_4__11_, u4_sll_453_ML_int_4__12_,
         u4_sll_453_ML_int_4__13_, u4_sll_453_ML_int_4__14_,
         u4_sll_453_ML_int_4__15_, u4_sll_453_ML_int_4__16_,
         u4_sll_453_ML_int_4__17_, u4_sll_453_ML_int_4__19_,
         u4_sll_453_ML_int_4__20_, u4_sll_453_ML_int_4__21_,
         u4_sll_453_ML_int_4__22_, u4_sll_453_ML_int_4__23_,
         u4_sll_453_ML_int_4__24_, u4_sll_453_ML_int_4__25_,
         u4_sll_453_ML_int_4__26_, u4_sll_453_ML_int_4__27_,
         u4_sll_453_ML_int_4__28_, u4_sll_453_ML_int_4__29_,
         u4_sll_453_ML_int_4__30_, u4_sll_453_ML_int_4__31_,
         u4_sll_453_ML_int_4__32_, u4_sll_453_ML_int_4__33_,
         u4_sll_453_ML_int_4__35_, u4_sll_453_ML_int_4__36_,
         u4_sll_453_ML_int_4__37_, u4_sll_453_ML_int_4__38_,
         u4_sll_453_ML_int_4__39_, u4_sll_453_ML_int_4__40_,
         u4_sll_453_ML_int_4__41_, u4_sll_453_ML_int_4__42_,
         u4_sll_453_ML_int_4__43_, u4_sll_453_ML_int_4__44_,
         u4_sll_453_ML_int_4__45_, u4_sll_453_ML_int_4__46_,
         u4_sll_453_ML_int_4__47_, u4_sll_453_ML_int_3__0_,
         u4_sll_453_ML_int_3__1_, u4_sll_453_ML_int_3__2_,
         u4_sll_453_ML_int_3__3_, u4_sll_453_ML_int_3__4_,
         u4_sll_453_ML_int_3__5_, u4_sll_453_ML_int_3__6_,
         u4_sll_453_ML_int_3__7_, u4_sll_453_ML_int_3__8_,
         u4_sll_453_ML_int_3__9_, u4_sll_453_ML_int_3__11_,
         u4_sll_453_ML_int_3__12_, u4_sll_453_ML_int_3__13_,
         u4_sll_453_ML_int_3__14_, u4_sll_453_ML_int_3__15_,
         u4_sll_453_ML_int_3__16_, u4_sll_453_ML_int_3__17_,
         u4_sll_453_ML_int_3__19_, u4_sll_453_ML_int_3__20_,
         u4_sll_453_ML_int_3__21_, u4_sll_453_ML_int_3__22_,
         u4_sll_453_ML_int_3__23_, u4_sll_453_ML_int_3__24_,
         u4_sll_453_ML_int_3__25_, u4_sll_453_ML_int_3__26_,
         u4_sll_453_ML_int_3__27_, u4_sll_453_ML_int_3__28_,
         u4_sll_453_ML_int_3__29_, u4_sll_453_ML_int_3__30_,
         u4_sll_453_ML_int_3__31_, u4_sll_453_ML_int_3__32_,
         u4_sll_453_ML_int_3__33_, u4_sll_453_ML_int_3__35_,
         u4_sll_453_ML_int_3__36_, u4_sll_453_ML_int_3__37_,
         u4_sll_453_ML_int_3__38_, u4_sll_453_ML_int_3__39_,
         u4_sll_453_ML_int_3__40_, u4_sll_453_ML_int_3__41_,
         u4_sll_453_ML_int_3__42_, u4_sll_453_ML_int_3__43_,
         u4_sll_453_ML_int_3__44_, u4_sll_453_ML_int_3__45_,
         u4_sll_453_ML_int_3__46_, u4_sll_453_ML_int_3__47_,
         u4_sll_453_ML_int_2__0_, u4_sll_453_ML_int_2__1_,
         u4_sll_453_ML_int_2__2_, u4_sll_453_ML_int_2__3_,
         u4_sll_453_ML_int_2__4_, u4_sll_453_ML_int_2__5_,
         u4_sll_453_ML_int_2__7_, u4_sll_453_ML_int_2__8_,
         u4_sll_453_ML_int_2__9_, u4_sll_453_ML_int_2__11_,
         u4_sll_453_ML_int_2__12_, u4_sll_453_ML_int_2__13_,
         u4_sll_453_ML_int_2__14_, u4_sll_453_ML_int_2__15_,
         u4_sll_453_ML_int_2__16_, u4_sll_453_ML_int_2__17_,
         u4_sll_453_ML_int_2__18_, u4_sll_453_ML_int_2__19_,
         u4_sll_453_ML_int_2__20_, u4_sll_453_ML_int_2__21_,
         u4_sll_453_ML_int_2__22_, u4_sll_453_ML_int_2__23_,
         u4_sll_453_ML_int_2__24_, u4_sll_453_ML_int_2__25_,
         u4_sll_453_ML_int_2__26_, u4_sll_453_ML_int_2__27_,
         u4_sll_453_ML_int_2__28_, u4_sll_453_ML_int_2__29_,
         u4_sll_453_ML_int_2__31_, u4_sll_453_ML_int_2__32_,
         u4_sll_453_ML_int_2__33_, u4_sll_453_ML_int_2__34_,
         u4_sll_453_ML_int_2__35_, u4_sll_453_ML_int_2__36_,
         u4_sll_453_ML_int_2__37_, u4_sll_453_ML_int_2__38_,
         u4_sll_453_ML_int_2__39_, u4_sll_453_ML_int_2__40_,
         u4_sll_453_ML_int_2__41_, u4_sll_453_ML_int_2__42_,
         u4_sll_453_ML_int_2__43_, u4_sll_453_ML_int_2__44_,
         u4_sll_453_ML_int_2__45_, u4_sll_453_ML_int_2__46_,
         u4_sll_453_ML_int_2__47_, u4_sll_453_ML_int_1__0_,
         u4_sll_453_ML_int_1__1_, u4_sll_453_ML_int_1__2_,
         u4_sll_453_ML_int_1__3_, u4_sll_453_ML_int_1__4_,
         u4_sll_453_ML_int_1__5_, u4_sll_453_ML_int_1__6_,
         u4_sll_453_ML_int_1__7_, u4_sll_453_ML_int_1__9_,
         u4_sll_453_ML_int_1__10_, u4_sll_453_ML_int_1__11_,
         u4_sll_453_ML_int_1__12_, u4_sll_453_ML_int_1__13_,
         u4_sll_453_ML_int_1__14_, u4_sll_453_ML_int_1__15_,
         u4_sll_453_ML_int_1__16_, u4_sll_453_ML_int_1__17_,
         u4_sll_453_ML_int_1__18_, u4_sll_453_ML_int_1__19_,
         u4_sll_453_ML_int_1__20_, u4_sll_453_ML_int_1__21_,
         u4_sll_453_ML_int_1__22_, u4_sll_453_ML_int_1__23_,
         u4_sll_453_ML_int_1__24_, u4_sll_453_ML_int_1__25_,
         u4_sll_453_ML_int_1__26_, u4_sll_453_ML_int_1__27_,
         u4_sll_453_ML_int_1__28_, u4_sll_453_ML_int_1__29_,
         u4_sll_453_ML_int_1__30_, u4_sll_453_ML_int_1__31_,
         u4_sll_453_ML_int_1__32_, u4_sll_453_ML_int_1__33_,
         u4_sll_453_ML_int_1__34_, u4_sll_453_ML_int_1__35_,
         u4_sll_453_ML_int_1__36_, u4_sll_453_ML_int_1__37_,
         u4_sll_453_ML_int_1__38_, u4_sll_453_ML_int_1__39_,
         u4_sll_453_ML_int_1__40_, u4_sll_453_ML_int_1__41_,
         u4_sll_453_ML_int_1__42_, u4_sll_453_ML_int_1__43_,
         u4_sll_453_ML_int_1__44_, u4_sll_453_ML_int_1__45_,
         u4_sll_453_ML_int_1__46_, u4_sll_453_ML_int_1__47_, u4_srl_452_n309,
         u4_srl_452_n308, u4_srl_452_n307, u4_srl_452_n306, u4_srl_452_n305,
         u4_srl_452_n304, u4_srl_452_n303, u4_srl_452_n302, u4_srl_452_n301,
         u4_srl_452_n300, u4_srl_452_n299, u4_srl_452_n298, u4_srl_452_n297,
         u4_srl_452_n296, u4_srl_452_n295, u4_srl_452_n294, u4_srl_452_n293,
         u4_srl_452_n292, u4_srl_452_n291, u4_srl_452_n290, u4_srl_452_n289,
         u4_srl_452_n288, u4_srl_452_n287, u4_srl_452_n286, u4_srl_452_n285,
         u4_srl_452_n284, u4_srl_452_n283, u4_srl_452_n282, u4_srl_452_n281,
         u4_srl_452_n280, u4_srl_452_n279, u4_srl_452_n278, u4_srl_452_n277,
         u4_srl_452_n276, u4_srl_452_n275, u4_srl_452_n274, u4_srl_452_n273,
         u4_srl_452_n272, u4_srl_452_n271, u4_srl_452_n270, u4_srl_452_n269,
         u4_srl_452_n268, u4_srl_452_n267, u4_srl_452_n266, u4_srl_452_n265,
         u4_srl_452_n264, u4_srl_452_n263, u4_srl_452_n262, u4_srl_452_n261,
         u4_srl_452_n260, u4_srl_452_n259, u4_srl_452_n258, u4_srl_452_n257,
         u4_srl_452_n256, u4_srl_452_n255, u4_srl_452_n254, u4_srl_452_n253,
         u4_srl_452_n252, u4_srl_452_n251, u4_srl_452_n250, u4_srl_452_n249,
         u4_srl_452_n248, u4_srl_452_n247, u4_srl_452_n246, u4_srl_452_n245,
         u4_srl_452_n244, u4_srl_452_n243, u4_srl_452_n242, u4_srl_452_n241,
         u4_srl_452_n240, u4_srl_452_n239, u4_srl_452_n238, u4_srl_452_n237,
         u4_srl_452_n236, u4_srl_452_n235, u4_srl_452_n234, u4_srl_452_n233,
         u4_srl_452_n232, u4_srl_452_n231, u4_srl_452_n230, u4_srl_452_n229,
         u4_srl_452_n228, u4_srl_452_n227, u4_srl_452_n226, u4_srl_452_n225,
         u4_srl_452_n224, u4_srl_452_n223, u4_srl_452_n222, u4_srl_452_n221,
         u4_srl_452_n220, u4_srl_452_n219, u4_srl_452_n218, u4_srl_452_n217,
         u4_srl_452_n216, u4_srl_452_n215, u4_srl_452_n214, u4_srl_452_n213,
         u4_srl_452_n212, u4_srl_452_n211, u4_srl_452_n210, u4_srl_452_n209,
         u4_srl_452_n208, u4_srl_452_n207, u4_srl_452_n206, u4_srl_452_n205,
         u4_srl_452_n204, u4_srl_452_n203, u4_srl_452_n202, u4_srl_452_n201,
         u4_srl_452_n200, u4_srl_452_n199, u4_srl_452_n198, u4_srl_452_n197,
         u4_srl_452_n196, u4_srl_452_n195, u4_srl_452_n194, u4_srl_452_n193,
         u4_srl_452_n192, u4_srl_452_n191, u4_srl_452_n190, u4_srl_452_n189,
         u4_srl_452_n188, u4_srl_452_n187, u4_srl_452_n186, u4_srl_452_n185,
         u4_srl_452_n184, u4_srl_452_n183, u4_srl_452_n182, u4_srl_452_n181,
         u4_srl_452_n180, u4_srl_452_n179, u4_srl_452_n178, u4_srl_452_n177,
         u4_srl_452_n176, u4_srl_452_n175, u4_srl_452_n174, u4_srl_452_n173,
         u4_srl_452_n172, u4_srl_452_n171, u4_srl_452_n170, u4_srl_452_n169,
         u4_srl_452_n168, u4_srl_452_n167, u4_srl_452_n166, u4_srl_452_n165,
         u4_srl_452_n164, u4_srl_452_n163, u4_srl_452_n162, u4_srl_452_n161,
         u4_srl_452_n160, u4_srl_452_n159, u4_srl_452_n158, u4_srl_452_n157,
         u4_srl_452_n156, u4_srl_452_n155, u4_srl_452_n154, u4_srl_452_n153,
         u4_srl_452_n152, u4_srl_452_n151, u4_srl_452_n150, u4_srl_452_n149,
         u4_srl_452_n148, u4_srl_452_n147, u4_srl_452_n146, u4_srl_452_n145,
         u4_srl_452_n144, u4_srl_452_n143, u4_srl_452_n142, u4_srl_452_n141,
         u4_srl_452_n140, u4_srl_452_n139, u4_srl_452_n138, u4_srl_452_n137,
         u4_srl_452_n136, u4_srl_452_n135, u4_srl_452_n134, u4_srl_452_n133,
         u4_srl_452_n132, u4_srl_452_n131, u4_srl_452_n130, u4_srl_452_n129,
         u4_srl_452_n128, u4_srl_452_n127, u4_srl_452_n126, u4_srl_452_n125,
         u4_srl_452_n124, u4_srl_452_n123, u4_srl_452_n122, u4_srl_452_n121,
         u4_srl_452_n120, u4_srl_452_n119, u4_srl_452_n118, u4_srl_452_n117,
         u4_srl_452_n116, u4_srl_452_n115, u4_srl_452_n114, u4_srl_452_n113,
         u4_srl_452_n112, u4_srl_452_n111, u4_srl_452_n110, u4_srl_452_n109,
         u4_srl_452_n108, u4_srl_452_n107, u4_srl_452_n106, u4_srl_452_n105,
         u4_srl_452_n104, u4_srl_452_n103, u4_srl_452_n102, u4_srl_452_n101,
         u4_srl_452_n100, u4_srl_452_n99, u4_srl_452_n98, u4_srl_452_n97,
         u4_srl_452_n96, u4_srl_452_n95, u4_srl_452_n94, u4_srl_452_n93,
         u4_srl_452_n92, u4_srl_452_n91, u4_srl_452_n90, u4_srl_452_n89,
         u4_srl_452_n88, u4_srl_452_n87, u4_srl_452_n86, u4_srl_452_n85,
         u4_srl_452_n84, u4_srl_452_n83, u4_srl_452_n82, u4_srl_452_n81,
         u4_srl_452_n80, u4_srl_452_n79, u4_srl_452_n78, u4_srl_452_n77,
         u4_srl_452_n76, u4_srl_452_n75, u4_srl_452_n74, u4_srl_452_n73,
         u4_srl_452_n72, u4_srl_452_n71, u4_srl_452_n70, u4_srl_452_n69,
         u4_srl_452_n68, u4_srl_452_n67, u4_srl_452_n66, u4_srl_452_n65,
         u4_srl_452_n64, u4_srl_452_n63, u4_srl_452_n62, u4_srl_452_n61,
         u4_srl_452_n60, u4_srl_452_n59, u4_srl_452_n58, u4_srl_452_n57,
         u4_srl_452_n56, u4_srl_452_n55, u4_srl_452_n54, u4_srl_452_n53,
         u4_srl_452_n52, u4_srl_452_n51, u4_srl_452_n50, u4_srl_452_n49,
         u4_srl_452_n48, u4_srl_452_n47, u4_srl_452_n46, u4_srl_452_n45,
         u4_srl_452_n44, u4_srl_452_n43, u4_srl_452_n42, u4_srl_452_n41,
         u4_srl_452_n40, u4_srl_452_n39, u4_srl_452_n38, u4_srl_452_n37,
         u4_srl_452_n36, u4_srl_452_n35, u4_srl_452_n34, u4_srl_452_n33,
         u4_srl_452_n32, u4_srl_452_n31, u4_srl_452_n30, u4_srl_452_n29,
         u4_srl_452_n28, u4_srl_452_n27, u4_srl_452_n26, u4_srl_452_n25,
         u4_srl_452_n24, u4_srl_452_n23, u4_srl_452_n22, u4_srl_452_n21,
         u4_srl_452_n20, u4_srl_452_n19, u4_srl_452_n18, u4_srl_452_n17,
         u4_srl_452_n16, u4_srl_452_n15, u4_srl_452_n14, u4_srl_452_n13,
         u4_srl_452_n12, u4_srl_452_n11, u4_srl_452_n10, u4_srl_452_n9,
         u4_srl_452_n8, u4_srl_452_n7, u4_srl_452_n6, u4_srl_452_n5,
         u4_srl_452_n4, u4_srl_452_n3, u4_srl_452_n2, u4_srl_452_n1,
         u4_sll_481_n95, u4_sll_481_n94, u4_sll_481_n93, u4_sll_481_n92,
         u4_sll_481_n91, u4_sll_481_n90, u4_sll_481_n89, u4_sll_481_n88,
         u4_sll_481_n87, u4_sll_481_n86, u4_sll_481_n85, u4_sll_481_n84,
         u4_sll_481_n83, u4_sll_481_n82, u4_sll_481_n81, u4_sll_481_n80,
         u4_sll_481_n79, u4_sll_481_n78, u4_sll_481_n77, u4_sll_481_n76,
         u4_sll_481_n75, u4_sll_481_n74, u4_sll_481_n73, u4_sll_481_n72,
         u4_sll_481_n71, u4_sll_481_n70, u4_sll_481_n69, u4_sll_481_n68,
         u4_sll_481_n67, u4_sll_481_n66, u4_sll_481_n65, u4_sll_481_n64,
         u4_sll_481_n63, u4_sll_481_n62, u4_sll_481_n61, u4_sll_481_n60,
         u4_sll_481_n59, u4_sll_481_n58, u4_sll_481_n57, u4_sll_481_n56,
         u4_sll_481_n55, u4_sll_481_n54, u4_sll_481_n53, u4_sll_481_n52,
         u4_sll_481_n51, u4_sll_481_n50, u4_sll_481_n49, u4_sll_481_n48,
         u4_sll_481_n47, u4_sll_481_n46, u4_sll_481_n45, u4_sll_481_n44,
         u4_sll_481_n43, u4_sll_481_n42, u4_sll_481_n41, u4_sll_481_n40,
         u4_sll_481_n39, u4_sll_481_n38, u4_sll_481_n37, u4_sll_481_n36,
         u4_sll_481_n35, u4_sll_481_n34, u4_sll_481_n33, u4_sll_481_n32,
         u4_sll_481_n31, u4_sll_481_n30, u4_sll_481_n29, u4_sll_481_n28,
         u4_sll_481_n27, u4_sll_481_n26, u4_sll_481_n25, u4_sll_481_n24,
         u4_sll_481_n23, u4_sll_481_n22, u4_sll_481_n21, u4_sll_481_n20,
         u4_sll_481_n19, u4_sll_481_n18, u4_sll_481_n17, u4_sll_481_n16,
         u4_sll_481_n15, u4_sll_481_n14, u4_sll_481_n13, u4_sll_481_n12,
         u4_sll_481_n11, u4_sll_481_n10, u4_sll_481_n9, u4_sll_481_n8,
         u4_sll_481_n7, u4_sll_481_n6, u4_sll_481_n5, u4_sll_481_n4,
         u4_sll_481_n3, u4_sll_481_n2, u4_sll_481_n1, u4_sll_481_ML_int_6__49_,
         u4_sll_481_ML_int_6__50_, u4_sll_481_ML_int_6__51_,
         u4_sll_481_ML_int_6__52_, u4_sll_481_ML_int_6__53_,
         u4_sll_481_ML_int_6__54_, u4_sll_481_ML_int_6__55_,
         u4_sll_481_ML_int_6__56_, u4_sll_481_ML_int_5__17_,
         u4_sll_481_ML_int_5__18_, u4_sll_481_ML_int_5__19_,
         u4_sll_481_ML_int_5__20_, u4_sll_481_ML_int_5__21_,
         u4_sll_481_ML_int_5__22_, u4_sll_481_ML_int_5__23_,
         u4_sll_481_ML_int_5__24_, u4_sll_481_ML_int_5__49_,
         u4_sll_481_ML_int_5__50_, u4_sll_481_ML_int_5__51_,
         u4_sll_481_ML_int_5__52_, u4_sll_481_ML_int_5__53_,
         u4_sll_481_ML_int_5__54_, u4_sll_481_ML_int_5__55_,
         u4_sll_481_ML_int_5__56_, u4_sll_481_ML_int_4__1_,
         u4_sll_481_ML_int_4__2_, u4_sll_481_ML_int_4__3_,
         u4_sll_481_ML_int_4__4_, u4_sll_481_ML_int_4__5_,
         u4_sll_481_ML_int_4__6_, u4_sll_481_ML_int_4__7_,
         u4_sll_481_ML_int_4__8_, u4_sll_481_ML_int_4__17_,
         u4_sll_481_ML_int_4__18_, u4_sll_481_ML_int_4__19_,
         u4_sll_481_ML_int_4__20_, u4_sll_481_ML_int_4__21_,
         u4_sll_481_ML_int_4__22_, u4_sll_481_ML_int_4__23_,
         u4_sll_481_ML_int_4__24_, u4_sll_481_ML_int_4__33_,
         u4_sll_481_ML_int_4__34_, u4_sll_481_ML_int_4__35_,
         u4_sll_481_ML_int_4__36_, u4_sll_481_ML_int_4__37_,
         u4_sll_481_ML_int_4__38_, u4_sll_481_ML_int_4__39_,
         u4_sll_481_ML_int_4__40_, u4_sll_481_ML_int_4__49_,
         u4_sll_481_ML_int_4__50_, u4_sll_481_ML_int_4__51_,
         u4_sll_481_ML_int_4__52_, u4_sll_481_ML_int_4__53_,
         u4_sll_481_ML_int_4__54_, u4_sll_481_ML_int_4__55_,
         u4_sll_481_ML_int_4__56_, u4_sll_481_ML_int_3__0_,
         u4_sll_481_ML_int_3__4_, u4_sll_481_ML_int_3__5_,
         u4_sll_481_ML_int_3__6_, u4_sll_481_ML_int_3__7_,
         u4_sll_481_ML_int_3__8_, u4_sll_481_ML_int_3__9_,
         u4_sll_481_ML_int_3__10_, u4_sll_481_ML_int_3__11_,
         u4_sll_481_ML_int_3__12_, u4_sll_481_ML_int_3__13_,
         u4_sll_481_ML_int_3__14_, u4_sll_481_ML_int_3__15_,
         u4_sll_481_ML_int_3__16_, u4_sll_481_ML_int_3__17_,
         u4_sll_481_ML_int_3__18_, u4_sll_481_ML_int_3__19_,
         u4_sll_481_ML_int_3__20_, u4_sll_481_ML_int_3__21_,
         u4_sll_481_ML_int_3__22_, u4_sll_481_ML_int_3__23_,
         u4_sll_481_ML_int_3__24_, u4_sll_481_ML_int_3__25_,
         u4_sll_481_ML_int_3__26_, u4_sll_481_ML_int_3__27_,
         u4_sll_481_ML_int_3__28_, u4_sll_481_ML_int_3__29_,
         u4_sll_481_ML_int_3__30_, u4_sll_481_ML_int_3__31_,
         u4_sll_481_ML_int_3__32_, u4_sll_481_ML_int_3__33_,
         u4_sll_481_ML_int_3__34_, u4_sll_481_ML_int_3__35_,
         u4_sll_481_ML_int_3__36_, u4_sll_481_ML_int_3__37_,
         u4_sll_481_ML_int_3__38_, u4_sll_481_ML_int_3__39_,
         u4_sll_481_ML_int_3__40_, u4_sll_481_ML_int_3__41_,
         u4_sll_481_ML_int_3__42_, u4_sll_481_ML_int_3__43_,
         u4_sll_481_ML_int_3__44_, u4_sll_481_ML_int_3__45_,
         u4_sll_481_ML_int_3__46_, u4_sll_481_ML_int_3__47_,
         u4_sll_481_ML_int_3__48_, u4_sll_481_ML_int_3__49_,
         u4_sll_481_ML_int_3__50_, u4_sll_481_ML_int_3__51_,
         u4_sll_481_ML_int_3__52_, u4_sll_481_ML_int_3__53_,
         u4_sll_481_ML_int_3__54_, u4_sll_481_ML_int_3__55_,
         u4_sll_481_ML_int_3__56_, u4_sll_481_ML_int_2__1_,
         u4_sll_481_ML_int_2__2_, u4_sll_481_ML_int_2__3_,
         u4_sll_481_ML_int_2__4_, u4_sll_481_ML_int_2__5_,
         u4_sll_481_ML_int_2__6_, u4_sll_481_ML_int_2__8_,
         u4_sll_481_ML_int_2__9_, u4_sll_481_ML_int_2__10_,
         u4_sll_481_ML_int_2__11_, u4_sll_481_ML_int_2__12_,
         u4_sll_481_ML_int_2__13_, u4_sll_481_ML_int_2__14_,
         u4_sll_481_ML_int_2__15_, u4_sll_481_ML_int_2__16_,
         u4_sll_481_ML_int_2__17_, u4_sll_481_ML_int_2__18_,
         u4_sll_481_ML_int_2__19_, u4_sll_481_ML_int_2__20_,
         u4_sll_481_ML_int_2__21_, u4_sll_481_ML_int_2__22_,
         u4_sll_481_ML_int_2__23_, u4_sll_481_ML_int_2__24_,
         u4_sll_481_ML_int_2__25_, u4_sll_481_ML_int_2__26_,
         u4_sll_481_ML_int_2__27_, u4_sll_481_ML_int_2__28_,
         u4_sll_481_ML_int_2__29_, u4_sll_481_ML_int_2__30_,
         u4_sll_481_ML_int_2__31_, u4_sll_481_ML_int_2__32_,
         u4_sll_481_ML_int_2__33_, u4_sll_481_ML_int_2__34_,
         u4_sll_481_ML_int_2__35_, u4_sll_481_ML_int_2__36_,
         u4_sll_481_ML_int_2__37_, u4_sll_481_ML_int_2__38_,
         u4_sll_481_ML_int_2__39_, u4_sll_481_ML_int_2__40_,
         u4_sll_481_ML_int_2__41_, u4_sll_481_ML_int_2__42_,
         u4_sll_481_ML_int_2__43_, u4_sll_481_ML_int_2__44_,
         u4_sll_481_ML_int_2__45_, u4_sll_481_ML_int_2__46_,
         u4_sll_481_ML_int_2__47_, u4_sll_481_ML_int_2__48_,
         u4_sll_481_ML_int_2__49_, u4_sll_481_ML_int_2__50_,
         u4_sll_481_ML_int_2__51_, u4_sll_481_ML_int_2__52_,
         u4_sll_481_ML_int_2__53_, u4_sll_481_ML_int_2__54_,
         u4_sll_481_ML_int_2__55_, u4_sll_481_ML_int_2__56_,
         u4_sll_481_ML_int_1__0_, u4_sll_481_ML_int_1__1_,
         u4_sll_481_ML_int_1__2_, u4_sll_481_ML_int_1__3_,
         u4_sll_481_ML_int_1__4_, u4_sll_481_ML_int_1__5_,
         u4_sll_481_ML_int_1__6_, u4_sll_481_ML_int_1__7_,
         u4_sll_481_ML_int_1__8_, u4_sll_481_ML_int_1__9_,
         u4_sll_481_ML_int_1__10_, u4_sll_481_ML_int_1__11_,
         u4_sll_481_ML_int_1__12_, u4_sll_481_ML_int_1__13_,
         u4_sll_481_ML_int_1__14_, u4_sll_481_ML_int_1__15_,
         u4_sll_481_ML_int_1__16_, u4_sll_481_ML_int_1__17_,
         u4_sll_481_ML_int_1__18_, u4_sll_481_ML_int_1__19_,
         u4_sll_481_ML_int_1__20_, u4_sll_481_ML_int_1__21_,
         u4_sll_481_ML_int_1__22_, u4_sll_481_ML_int_1__23_,
         u4_sll_481_ML_int_1__24_, u4_sll_481_ML_int_1__25_,
         u4_sll_481_ML_int_1__26_, u4_sll_481_ML_int_1__27_,
         u4_sll_481_ML_int_1__28_, u4_sll_481_ML_int_1__29_,
         u4_sll_481_ML_int_1__30_, u4_sll_481_ML_int_1__31_,
         u4_sll_481_ML_int_1__32_, u4_sll_481_ML_int_1__33_,
         u4_sll_481_ML_int_1__34_, u4_sll_481_ML_int_1__35_,
         u4_sll_481_ML_int_1__36_, u4_sll_481_ML_int_1__37_,
         u4_sll_481_ML_int_1__38_, u4_sll_481_ML_int_1__39_,
         u4_sll_481_ML_int_1__40_, u4_sll_481_ML_int_1__41_,
         u4_sll_481_ML_int_1__42_, u4_sll_481_ML_int_1__43_,
         u4_sll_481_ML_int_1__44_, u4_sll_481_ML_int_1__45_,
         u4_sll_481_ML_int_1__46_, u4_sll_481_ML_int_1__47_,
         u4_sll_481_ML_int_1__49_, u4_sll_481_ML_int_1__51_,
         u4_sll_481_ML_int_1__52_, u4_sll_481_ML_int_1__53_,
         u4_sll_481_ML_int_1__54_, u4_sll_481_ML_int_1__55_,
         u4_sll_481_MR_int_1__55_, u4_sll_481_SHMAG_4_, u4_sll_481_SHMAG_5_,
         u4_sll_481_temp_int_SH_0_, u4_sll_481_temp_int_SH_1_,
         u4_sll_481_temp_int_SH_3_, u4_sub_411_n15, u4_sub_411_n14,
         u4_sub_411_n13, u4_sub_411_n12, u4_sub_411_n11, u4_sub_411_n10,
         u4_sub_411_n9, u4_sub_411_n8, u4_sub_411_n7, u4_sub_411_n6,
         u4_sub_411_n5, u4_sub_411_n4, u4_sub_411_carry_1_,
         u4_sub_411_carry_2_, u4_sub_411_carry_3_, u4_sub_411_carry_4_,
         u4_sub_411_carry_5_, u4_sub_411_carry_6_, u4_sub_411_carry_7_,
         u4_add_410_n7, u4_add_410_n6, u4_add_410_n5, u4_add_410_n4,
         u4_add_410_n3, u4_add_410_n2, u4_add_410_carry_1_,
         u4_add_410_carry_2_, u4_add_410_carry_3_, u4_add_410_carry_4_,
         u4_add_410_carry_5_, u4_add_410_carry_6_, u4_add_410_carry_7_,
         u3_sub_60_n30, u3_sub_60_n29, u3_sub_60_n28, u3_sub_60_n27,
         u3_sub_60_n26, u3_sub_60_n25, u3_sub_60_n24, u3_sub_60_n23,
         u3_sub_60_n22, u3_sub_60_n21, u3_sub_60_n20, u3_sub_60_n19,
         u3_sub_60_n18, u3_sub_60_n17, u3_sub_60_n16, u3_sub_60_n15,
         u3_sub_60_n14, u3_sub_60_n13, u3_sub_60_n12, u3_sub_60_n11,
         u3_sub_60_n10, u3_sub_60_n9, u3_sub_60_n8, u3_sub_60_n7, u3_sub_60_n6,
         u3_sub_60_n5, u3_sub_60_n4, u3_sub_60_n2, u3_sub_60_n1, u3_add_60_n3,
         u3_add_60_n2, u3_add_60_n1, u2_add_112_n2, u2_sub_112_n11,
         u2_sub_112_n10, u2_sub_112_n9, u2_sub_112_n8, u2_sub_112_n7,
         u2_sub_112_n6, u2_sub_112_n5, u2_sub_112_n4, u2_sub_112_n2,
         u2_sub_112_n1, u1_srl_148_n147, u1_srl_148_n146, u1_srl_148_n145,
         u1_srl_148_n144, u1_srl_148_n143, u1_srl_148_n142, u1_srl_148_n141,
         u1_srl_148_n140, u1_srl_148_n139, u1_srl_148_n138, u1_srl_148_n137,
         u1_srl_148_n136, u1_srl_148_n135, u1_srl_148_n134, u1_srl_148_n133,
         u1_srl_148_n132, u1_srl_148_n131, u1_srl_148_n130, u1_srl_148_n129,
         u1_srl_148_n128, u1_srl_148_n127, u1_srl_148_n126, u1_srl_148_n125,
         u1_srl_148_n124, u1_srl_148_n123, u1_srl_148_n122, u1_srl_148_n121,
         u1_srl_148_n120, u1_srl_148_n119, u1_srl_148_n118, u1_srl_148_n117,
         u1_srl_148_n116, u1_srl_148_n115, u1_srl_148_n114, u1_srl_148_n113,
         u1_srl_148_n112, u1_srl_148_n111, u1_srl_148_n110, u1_srl_148_n109,
         u1_srl_148_n108, u1_srl_148_n107, u1_srl_148_n106, u1_srl_148_n105,
         u1_srl_148_n104, u1_srl_148_n103, u1_srl_148_n102, u1_srl_148_n101,
         u1_srl_148_n100, u1_srl_148_n99, u1_srl_148_n98, u1_srl_148_n97,
         u1_srl_148_n96, u1_srl_148_n95, u1_srl_148_n94, u1_srl_148_n93,
         u1_srl_148_n92, u1_srl_148_n91, u1_srl_148_n90, u1_srl_148_n89,
         u1_srl_148_n88, u1_srl_148_n87, u1_srl_148_n86, u1_srl_148_n85,
         u1_srl_148_n84, u1_srl_148_n83, u1_srl_148_n82, u1_srl_148_n81,
         u1_srl_148_n80, u1_srl_148_n79, u1_srl_148_n78, u1_srl_148_n77,
         u1_srl_148_n76, u1_srl_148_n75, u1_srl_148_n74, u1_srl_148_n73,
         u1_srl_148_n72, u1_srl_148_n71, u1_srl_148_n70, u1_srl_148_n69,
         u1_srl_148_n68, u1_srl_148_n67, u1_srl_148_n66, u1_srl_148_n65,
         u1_srl_148_n64, u1_srl_148_n63, u1_srl_148_n62, u1_srl_148_n61,
         u1_srl_148_n60, u1_srl_148_n59, u1_srl_148_n58, u1_srl_148_n57,
         u1_srl_148_n56, u1_srl_148_n55, u1_srl_148_n54, u1_srl_148_n53,
         u1_srl_148_n52, u1_srl_148_n51, u1_srl_148_n50, u1_srl_148_n49,
         u1_srl_148_n48, u1_srl_148_n47, u1_srl_148_n46, u1_srl_148_n45,
         u1_srl_148_n44, u1_srl_148_n43, u1_srl_148_n42, u1_srl_148_n41,
         u1_srl_148_n40, u1_srl_148_n39, u1_srl_148_n38, u1_srl_148_n37,
         u1_srl_148_n36, u1_srl_148_n35, u1_srl_148_n34, u1_srl_148_n33,
         u1_srl_148_n32, u1_srl_148_n31, u1_srl_148_n30, u1_srl_148_n29,
         u1_srl_148_n28, u1_srl_148_n27, u1_srl_148_n26, u1_srl_148_n25,
         u1_srl_148_n24, u1_srl_148_n23, u1_srl_148_n22, u1_srl_148_n21,
         u1_srl_148_n20, u1_srl_148_n19, u1_srl_148_n18, u1_srl_148_n17,
         u1_srl_148_n16, u1_srl_148_n14, u1_srl_148_n12, u1_srl_148_n11,
         u1_srl_148_n10, u1_srl_148_n9, u1_srl_148_n8, u1_srl_148_n7,
         u1_srl_148_n6, u1_srl_148_n5, u1_srl_148_n4, u1_srl_148_n3,
         u1_srl_148_n2, u1_srl_148_n1, sub_434_3_n84, sub_434_3_n83,
         sub_434_3_n82, sub_434_3_n81, sub_434_3_n80, sub_434_3_n79,
         sub_434_3_n78, sub_434_3_n77, sub_434_3_n76, sub_434_3_n75,
         sub_434_3_n74, sub_434_3_n73, sub_434_3_n72, sub_434_3_n71,
         sub_434_3_n70, sub_434_3_n69, sub_434_3_n68, sub_434_3_n67,
         sub_434_3_n66, sub_434_3_n65, sub_434_3_n64, sub_434_3_n63,
         sub_434_3_n62, sub_434_3_n61, sub_434_3_n60, sub_434_3_n59,
         sub_434_3_n58, sub_434_3_n57, sub_434_3_n56, sub_434_3_n55,
         sub_434_3_n54, sub_434_3_n53, sub_434_3_n52, sub_434_3_n51,
         sub_434_3_n50, sub_434_3_n49, sub_434_3_n48, sub_434_3_n47,
         sub_434_3_n46, sub_434_3_n45, sub_434_3_n44, sub_434_3_n43,
         sub_434_3_n42, sub_434_3_n41, sub_434_3_n40, sub_434_3_n39,
         sub_434_3_n38, sub_434_3_n37, sub_434_3_n36, sub_434_3_n35,
         sub_434_3_n34, sub_434_3_n33, sub_434_3_n32, sub_434_3_n31,
         sub_434_3_n30, sub_434_3_n29, sub_434_3_n28, sub_434_3_n27,
         sub_434_3_n26, sub_434_3_n25, sub_434_3_carry_21_,
         sub_434_3_carry_22_, sub_434_3_carry_23_, sub_434_3_carry_24_,
         sub_434_3_carry_25_, sub_434_3_carry_26_, sub_434_3_carry_27_,
         sub_434_3_carry_28_, sub_434_3_carry_29_, sub_434_3_carry_30_,
         sub_434_3_carry_31_, sub_434_3_carry_32_, sub_434_3_carry_33_,
         sub_434_3_carry_34_, sub_434_3_carry_35_, sub_434_3_carry_36_,
         sub_434_3_carry_37_, sub_434_3_carry_38_, sub_434_3_carry_39_,
         sub_434_3_carry_40_, sub_434_3_carry_41_, sub_434_3_carry_42_,
         sub_434_3_carry_43_, sub_434_3_carry_44_, sub_434_3_carry_45_,
         sub_434_3_carry_46_, sub_434_3_carry_47_, sub_434_b0_n70,
         sub_434_b0_n69, sub_434_b0_n68, sub_434_b0_n67, sub_434_b0_n66,
         sub_434_b0_n65, sub_434_b0_n64, sub_434_b0_n63, sub_434_b0_n62,
         sub_434_b0_n61, sub_434_b0_n60, sub_434_b0_n59, sub_434_b0_n58,
         sub_434_b0_n57, sub_434_b0_n56, sub_434_b0_n55, sub_434_b0_n54,
         sub_434_b0_n53, sub_434_b0_n52, sub_434_b0_n51, sub_434_b0_n50,
         sub_434_b0_n49, sub_434_b0_n48, sub_434_b0_n47, sub_434_b0_n46,
         sub_434_b0_n45, sub_434_b0_n44, sub_434_b0_n43, sub_434_b0_n42,
         sub_434_b0_n41, sub_434_b0_n40, sub_434_b0_n39, sub_434_b0_n38,
         sub_434_b0_n37, sub_434_b0_n12, sub_434_b0_n11, sub_434_b0_n10,
         sub_434_b0_n9, sub_434_b0_n8, sub_434_b0_n7, sub_434_b0_n6,
         sub_434_b0_n5, sub_434_b0_n4, sub_434_b0_n3, sub_434_b0_n2,
         sub_434_b0_n1, sub_434_b0_carry_3_, sub_434_b0_carry_5_,
         sub_434_b0_carry_8_, sub_434_b0_carry_10_, sub_434_b0_carry_12_,
         sub_434_b0_carry_14_, sub_434_b0_carry_16_, sub_434_b0_carry_18_,
         sub_434_b0_carry_20_, sub_434_b0_carry_22_, sll_384_n24, sll_384_n23,
         sll_384_n22, sll_384_n21, sll_384_n20, sll_384_n19, sll_384_n18,
         sll_384_n17, sll_384_n16, sll_384_n15, sll_384_n14, sll_384_n13,
         sll_384_n12, sll_384_n11, sll_384_n10, sll_384_n9, sll_384_n8,
         sll_384_n7, sll_384_n6, sll_384_n5, sll_384_n4, sll_384_n3,
         sll_384_n2, sll_384_n1, sll_384_ML_int_4__8_, sll_384_ML_int_4__9_,
         sll_384_ML_int_4__10_, sll_384_ML_int_4__11_, sll_384_ML_int_4__12_,
         sll_384_ML_int_4__13_, sll_384_ML_int_4__14_, sll_384_ML_int_4__15_,
         sll_384_ML_int_4__16_, sll_384_ML_int_4__17_, sll_384_ML_int_4__18_,
         sll_384_ML_int_4__19_, sll_384_ML_int_4__20_, sll_384_ML_int_4__21_,
         sll_384_ML_int_4__22_, sll_384_ML_int_4__23_, sll_384_ML_int_3__0_,
         sll_384_ML_int_3__1_, sll_384_ML_int_3__2_, sll_384_ML_int_3__3_,
         sll_384_ML_int_3__4_, sll_384_ML_int_3__5_, sll_384_ML_int_3__6_,
         sll_384_ML_int_3__7_, sll_384_ML_int_3__8_, sll_384_ML_int_3__9_,
         sll_384_ML_int_3__10_, sll_384_ML_int_3__11_, sll_384_ML_int_3__12_,
         sll_384_ML_int_3__13_, sll_384_ML_int_3__14_, sll_384_ML_int_3__15_,
         sll_384_ML_int_3__16_, sll_384_ML_int_3__17_, sll_384_ML_int_3__18_,
         sll_384_ML_int_3__19_, sll_384_ML_int_3__20_, sll_384_ML_int_3__21_,
         sll_384_ML_int_3__22_, sll_384_ML_int_3__23_, sll_384_ML_int_2__0_,
         sll_384_ML_int_2__1_, sll_384_ML_int_2__2_, sll_384_ML_int_2__3_,
         sll_384_ML_int_2__4_, sll_384_ML_int_2__5_, sll_384_ML_int_2__6_,
         sll_384_ML_int_2__7_, sll_384_ML_int_2__8_, sll_384_ML_int_2__9_,
         sll_384_ML_int_2__10_, sll_384_ML_int_2__11_, sll_384_ML_int_2__12_,
         sll_384_ML_int_2__13_, sll_384_ML_int_2__14_, sll_384_ML_int_2__15_,
         sll_384_ML_int_2__16_, sll_384_ML_int_2__17_, sll_384_ML_int_2__18_,
         sll_384_ML_int_2__19_, sll_384_ML_int_2__20_, sll_384_ML_int_2__21_,
         sll_384_ML_int_2__22_, sll_384_ML_int_2__23_, sll_384_ML_int_1__0_,
         sll_384_ML_int_1__1_, sll_384_ML_int_1__2_, sll_384_ML_int_1__3_,
         sll_384_ML_int_1__4_, sll_384_ML_int_1__5_, sll_384_ML_int_1__6_,
         sll_384_ML_int_1__7_, sll_384_ML_int_1__8_, sll_384_ML_int_1__9_,
         sll_384_ML_int_1__10_, sll_384_ML_int_1__11_, sll_384_ML_int_1__12_,
         sll_384_ML_int_1__13_, sll_384_ML_int_1__14_, sll_384_ML_int_1__15_,
         sll_384_ML_int_1__16_, sll_384_ML_int_1__17_, sll_384_ML_int_1__18_,
         sll_384_ML_int_1__19_, sll_384_ML_int_1__20_, sll_384_ML_int_1__21_,
         sll_384_ML_int_1__22_, sll_384_ML_int_1__23_, r473_n81, r473_n80,
         r473_n79, r473_n78, r473_n77, r473_n76, r473_n75, r473_n74, r473_n73,
         r473_n72, r473_n71, r473_n70, r473_n69, r473_n68, r473_n67, r473_n66,
         r473_n65, r473_n64, r473_n63, r473_n62, r473_n61, r473_n60, r473_n59,
         r473_n58, r473_n57, r473_n56, r473_n55, r473_n54, r473_n53, r473_n52,
         r473_n51, r473_n50, r473_n49, r473_n48, r473_n47, r473_n46, r473_n45,
         r473_n44, r473_n43, r473_n42, r473_n41, r473_n40, r473_n39, r473_n38,
         r473_n37, r473_n36, r473_n35, r473_n34, r473_n33, r473_n32, r473_n31,
         r473_n30, r473_n29, r473_n28, r473_n27, r473_n26, r473_n25, r473_n24,
         r473_n23, r473_n22, r473_n21, r473_n20, r473_n19, r473_n18, r473_n17,
         r473_n16, r473_n15, r473_n14, r473_n13, r473_n12, r473_n11, r473_n10,
         r473_n9, r473_n8, r473_n7, r473_n6, r473_n5, r473_n4, r473_n3,
         r473_n2, sub_1_root_sub_0_root_u4_add_496_n10,
         sub_1_root_sub_0_root_u4_add_496_n9,
         sub_1_root_sub_0_root_u4_add_496_n8,
         sub_1_root_sub_0_root_u4_add_496_n7,
         sub_1_root_sub_0_root_u4_add_496_n6,
         sub_1_root_sub_0_root_u4_add_496_n5,
         sub_1_root_sub_0_root_u4_add_496_n4,
         sub_1_root_sub_0_root_u4_add_496_n3,
         sub_1_root_sub_0_root_u4_add_496_n2,
         sub_1_root_sub_0_root_u4_add_496_n1,
         sub_1_root_sub_0_root_u4_add_496_carry_1_,
         sub_1_root_sub_0_root_u4_add_496_carry_2_,
         sub_1_root_sub_0_root_u4_add_496_carry_3_,
         sub_1_root_sub_0_root_u4_add_496_carry_4_,
         sub_1_root_sub_0_root_u4_add_496_carry_5_,
         sub_1_root_sub_0_root_u4_add_496_carry_6_,
         sub_1_root_sub_0_root_u4_add_496_carry_7_, u5_mult_79_n1882,
         u5_mult_79_n1881, u5_mult_79_n1880, u5_mult_79_n1879,
         u5_mult_79_n1878, u5_mult_79_n1877, u5_mult_79_n1876,
         u5_mult_79_n1875, u5_mult_79_n1874, u5_mult_79_n1873,
         u5_mult_79_n1872, u5_mult_79_n1871, u5_mult_79_n1870,
         u5_mult_79_n1869, u5_mult_79_n1868, u5_mult_79_n1867,
         u5_mult_79_n1866, u5_mult_79_n1865, u5_mult_79_n1864,
         u5_mult_79_n1863, u5_mult_79_n1862, u5_mult_79_n1861,
         u5_mult_79_n1860, u5_mult_79_n1859, u5_mult_79_n1858,
         u5_mult_79_n1857, u5_mult_79_n1856, u5_mult_79_n1855,
         u5_mult_79_n1854, u5_mult_79_n1853, u5_mult_79_n1852,
         u5_mult_79_n1851, u5_mult_79_n1850, u5_mult_79_n1849,
         u5_mult_79_n1848, u5_mult_79_n1847, u5_mult_79_n1846,
         u5_mult_79_n1845, u5_mult_79_n1844, u5_mult_79_n1843,
         u5_mult_79_n1842, u5_mult_79_n1841, u5_mult_79_n1840,
         u5_mult_79_n1839, u5_mult_79_n1838, u5_mult_79_n1837,
         u5_mult_79_n1836, u5_mult_79_n1835, u5_mult_79_n1834,
         u5_mult_79_n1833, u5_mult_79_n1832, u5_mult_79_n1831,
         u5_mult_79_n1830, u5_mult_79_n1829, u5_mult_79_n1828,
         u5_mult_79_n1827, u5_mult_79_n1826, u5_mult_79_n1825,
         u5_mult_79_n1824, u5_mult_79_n1823, u5_mult_79_n1822,
         u5_mult_79_n1821, u5_mult_79_n1820, u5_mult_79_n1819,
         u5_mult_79_n1818, u5_mult_79_n1817, u5_mult_79_n1816,
         u5_mult_79_n1815, u5_mult_79_n1814, u5_mult_79_n1813,
         u5_mult_79_n1812, u5_mult_79_n1811, u5_mult_79_n1810,
         u5_mult_79_n1809, u5_mult_79_n1808, u5_mult_79_n1807,
         u5_mult_79_n1806, u5_mult_79_n1805, u5_mult_79_n1804,
         u5_mult_79_n1803, u5_mult_79_n1802, u5_mult_79_n1801,
         u5_mult_79_n1800, u5_mult_79_n1799, u5_mult_79_n1798,
         u5_mult_79_n1797, u5_mult_79_n1796, u5_mult_79_n1795,
         u5_mult_79_n1794, u5_mult_79_n1793, u5_mult_79_n1792,
         u5_mult_79_n1791, u5_mult_79_n1790, u5_mult_79_n1789,
         u5_mult_79_n1788, u5_mult_79_n1787, u5_mult_79_n1786,
         u5_mult_79_n1785, u5_mult_79_n1784, u5_mult_79_n1783,
         u5_mult_79_n1782, u5_mult_79_n1781, u5_mult_79_n1780,
         u5_mult_79_n1779, u5_mult_79_n1778, u5_mult_79_n1777,
         u5_mult_79_n1776, u5_mult_79_n1775, u5_mult_79_n1774,
         u5_mult_79_n1773, u5_mult_79_n1772, u5_mult_79_n1771,
         u5_mult_79_n1770, u5_mult_79_n1769, u5_mult_79_n1768,
         u5_mult_79_n1767, u5_mult_79_n1766, u5_mult_79_n1765,
         u5_mult_79_n1764, u5_mult_79_n1763, u5_mult_79_n1762,
         u5_mult_79_n1761, u5_mult_79_n1760, u5_mult_79_n1759,
         u5_mult_79_n1758, u5_mult_79_n1757, u5_mult_79_n1756,
         u5_mult_79_n1755, u5_mult_79_n1754, u5_mult_79_n1753,
         u5_mult_79_n1752, u5_mult_79_n1751, u5_mult_79_n1750,
         u5_mult_79_n1749, u5_mult_79_n1748, u5_mult_79_n1747,
         u5_mult_79_n1746, u5_mult_79_n1745, u5_mult_79_n1744,
         u5_mult_79_n1743, u5_mult_79_n1742, u5_mult_79_n1741,
         u5_mult_79_n1740, u5_mult_79_n1739, u5_mult_79_n1738,
         u5_mult_79_n1737, u5_mult_79_n1736, u5_mult_79_n1735,
         u5_mult_79_n1734, u5_mult_79_n1733, u5_mult_79_n1732,
         u5_mult_79_n1731, u5_mult_79_n1730, u5_mult_79_n1729,
         u5_mult_79_n1728, u5_mult_79_n1727, u5_mult_79_n1726,
         u5_mult_79_n1725, u5_mult_79_n1724, u5_mult_79_n1723,
         u5_mult_79_n1722, u5_mult_79_n1721, u5_mult_79_n1720,
         u5_mult_79_n1719, u5_mult_79_n1718, u5_mult_79_n1717,
         u5_mult_79_n1716, u5_mult_79_n1715, u5_mult_79_n1714,
         u5_mult_79_n1713, u5_mult_79_n1712, u5_mult_79_n1711,
         u5_mult_79_n1710, u5_mult_79_n1709, u5_mult_79_n1708,
         u5_mult_79_n1707, u5_mult_79_n1706, u5_mult_79_n1705,
         u5_mult_79_n1704, u5_mult_79_n1703, u5_mult_79_n1702,
         u5_mult_79_n1701, u5_mult_79_n1700, u5_mult_79_n1699,
         u5_mult_79_n1698, u5_mult_79_n1697, u5_mult_79_n1696,
         u5_mult_79_n1695, u5_mult_79_n1694, u5_mult_79_n1693,
         u5_mult_79_n1692, u5_mult_79_n1691, u5_mult_79_n1690,
         u5_mult_79_n1689, u5_mult_79_n1688, u5_mult_79_n1687,
         u5_mult_79_n1686, u5_mult_79_n1685, u5_mult_79_n1684,
         u5_mult_79_n1683, u5_mult_79_n1682, u5_mult_79_n1681,
         u5_mult_79_n1680, u5_mult_79_n1679, u5_mult_79_n1678,
         u5_mult_79_n1677, u5_mult_79_n1676, u5_mult_79_n1675,
         u5_mult_79_n1674, u5_mult_79_n1673, u5_mult_79_n1672,
         u5_mult_79_n1671, u5_mult_79_n1670, u5_mult_79_n1669,
         u5_mult_79_n1668, u5_mult_79_n1667, u5_mult_79_n1666,
         u5_mult_79_n1665, u5_mult_79_n1664, u5_mult_79_n1663,
         u5_mult_79_n1662, u5_mult_79_n1661, u5_mult_79_n1660,
         u5_mult_79_n1659, u5_mult_79_n1658, u5_mult_79_n1657,
         u5_mult_79_n1656, u5_mult_79_n1655, u5_mult_79_n1654,
         u5_mult_79_n1653, u5_mult_79_n1652, u5_mult_79_n1651,
         u5_mult_79_n1650, u5_mult_79_n1649, u5_mult_79_n1648,
         u5_mult_79_n1647, u5_mult_79_n1646, u5_mult_79_n1645,
         u5_mult_79_n1644, u5_mult_79_n1643, u5_mult_79_n1642,
         u5_mult_79_n1641, u5_mult_79_n1640, u5_mult_79_n1639,
         u5_mult_79_n1638, u5_mult_79_n1637, u5_mult_79_n1636,
         u5_mult_79_n1635, u5_mult_79_n1634, u5_mult_79_n1633,
         u5_mult_79_n1632, u5_mult_79_n1631, u5_mult_79_n1630,
         u5_mult_79_n1629, u5_mult_79_n1628, u5_mult_79_n1627,
         u5_mult_79_n1626, u5_mult_79_n1625, u5_mult_79_n1624,
         u5_mult_79_n1623, u5_mult_79_n1622, u5_mult_79_n1621,
         u5_mult_79_n1620, u5_mult_79_n1619, u5_mult_79_n1618,
         u5_mult_79_n1617, u5_mult_79_n1616, u5_mult_79_n1615,
         u5_mult_79_n1614, u5_mult_79_n1613, u5_mult_79_n1612,
         u5_mult_79_n1611, u5_mult_79_n1610, u5_mult_79_n1609,
         u5_mult_79_n1608, u5_mult_79_n1607, u5_mult_79_n1606,
         u5_mult_79_n1605, u5_mult_79_n1604, u5_mult_79_n1603,
         u5_mult_79_n1602, u5_mult_79_n1601, u5_mult_79_n1600,
         u5_mult_79_n1599, u5_mult_79_n1598, u5_mult_79_n1597,
         u5_mult_79_n1596, u5_mult_79_n1595, u5_mult_79_n1594,
         u5_mult_79_n1593, u5_mult_79_n1592, u5_mult_79_n1591,
         u5_mult_79_n1590, u5_mult_79_n1589, u5_mult_79_n1588,
         u5_mult_79_n1587, u5_mult_79_n1586, u5_mult_79_n1585,
         u5_mult_79_n1584, u5_mult_79_n1583, u5_mult_79_n1582,
         u5_mult_79_n1581, u5_mult_79_n1580, u5_mult_79_n1579,
         u5_mult_79_n1578, u5_mult_79_n1577, u5_mult_79_n1576,
         u5_mult_79_n1575, u5_mult_79_n1574, u5_mult_79_n1573,
         u5_mult_79_n1572, u5_mult_79_n1571, u5_mult_79_n1570,
         u5_mult_79_n1569, u5_mult_79_n1568, u5_mult_79_n1567,
         u5_mult_79_n1566, u5_mult_79_n1565, u5_mult_79_n1564,
         u5_mult_79_n1563, u5_mult_79_n1562, u5_mult_79_n1561,
         u5_mult_79_n1560, u5_mult_79_n1559, u5_mult_79_n1558,
         u5_mult_79_n1557, u5_mult_79_n1556, u5_mult_79_n1555,
         u5_mult_79_n1554, u5_mult_79_n1553, u5_mult_79_n1552,
         u5_mult_79_n1551, u5_mult_79_n1550, u5_mult_79_n1549,
         u5_mult_79_n1548, u5_mult_79_n1547, u5_mult_79_n1546,
         u5_mult_79_n1545, u5_mult_79_n1544, u5_mult_79_n1543,
         u5_mult_79_n1542, u5_mult_79_n1541, u5_mult_79_n1540,
         u5_mult_79_n1539, u5_mult_79_n1538, u5_mult_79_n1537,
         u5_mult_79_n1536, u5_mult_79_n1535, u5_mult_79_n1534,
         u5_mult_79_n1533, u5_mult_79_n1532, u5_mult_79_n1531,
         u5_mult_79_n1530, u5_mult_79_n1529, u5_mult_79_n1528,
         u5_mult_79_n1527, u5_mult_79_n1526, u5_mult_79_n1525,
         u5_mult_79_n1524, u5_mult_79_n1523, u5_mult_79_n1522,
         u5_mult_79_n1521, u5_mult_79_n1520, u5_mult_79_n1519,
         u5_mult_79_n1518, u5_mult_79_n1517, u5_mult_79_n1516,
         u5_mult_79_n1515, u5_mult_79_n1514, u5_mult_79_n1513,
         u5_mult_79_n1512, u5_mult_79_n1511, u5_mult_79_n1510,
         u5_mult_79_n1509, u5_mult_79_n1508, u5_mult_79_n1507,
         u5_mult_79_n1506, u5_mult_79_n1505, u5_mult_79_n1504,
         u5_mult_79_n1503, u5_mult_79_n1502, u5_mult_79_n1501,
         u5_mult_79_n1500, u5_mult_79_n1499, u5_mult_79_n1498,
         u5_mult_79_n1497, u5_mult_79_n1496, u5_mult_79_n1495,
         u5_mult_79_n1494, u5_mult_79_n1493, u5_mult_79_n1492,
         u5_mult_79_n1491, u5_mult_79_n1490, u5_mult_79_n1489,
         u5_mult_79_n1488, u5_mult_79_n1487, u5_mult_79_n1486,
         u5_mult_79_n1485, u5_mult_79_n1484, u5_mult_79_n1483,
         u5_mult_79_n1482, u5_mult_79_n1481, u5_mult_79_n1480,
         u5_mult_79_n1479, u5_mult_79_n1478, u5_mult_79_n1477,
         u5_mult_79_n1476, u5_mult_79_n1475, u5_mult_79_n1474,
         u5_mult_79_n1473, u5_mult_79_n1472, u5_mult_79_n1471,
         u5_mult_79_n1470, u5_mult_79_n1469, u5_mult_79_n1468,
         u5_mult_79_n1467, u5_mult_79_n1466, u5_mult_79_n1465,
         u5_mult_79_n1464, u5_mult_79_n1463, u5_mult_79_n1462,
         u5_mult_79_n1461, u5_mult_79_n1460, u5_mult_79_n1459,
         u5_mult_79_n1458, u5_mult_79_n1457, u5_mult_79_n1456,
         u5_mult_79_n1455, u5_mult_79_n1454, u5_mult_79_n1453,
         u5_mult_79_n1452, u5_mult_79_n1451, u5_mult_79_n1450,
         u5_mult_79_n1449, u5_mult_79_n1448, u5_mult_79_n1447,
         u5_mult_79_n1446, u5_mult_79_n1445, u5_mult_79_n1444,
         u5_mult_79_n1443, u5_mult_79_n1442, u5_mult_79_n1441,
         u5_mult_79_n1440, u5_mult_79_n1439, u5_mult_79_n1438,
         u5_mult_79_n1437, u5_mult_79_n1436, u5_mult_79_n1435,
         u5_mult_79_n1434, u5_mult_79_n1433, u5_mult_79_n1432,
         u5_mult_79_n1431, u5_mult_79_n1430, u5_mult_79_n1429,
         u5_mult_79_n1428, u5_mult_79_n1427, u5_mult_79_n1426,
         u5_mult_79_n1425, u5_mult_79_n1424, u5_mult_79_n1423,
         u5_mult_79_n1422, u5_mult_79_n1421, u5_mult_79_n1420,
         u5_mult_79_n1419, u5_mult_79_n1418, u5_mult_79_n1417,
         u5_mult_79_n1416, u5_mult_79_n1415, u5_mult_79_n1414,
         u5_mult_79_n1413, u5_mult_79_n1412, u5_mult_79_n1411,
         u5_mult_79_n1410, u5_mult_79_n1409, u5_mult_79_n1408,
         u5_mult_79_n1407, u5_mult_79_n1406, u5_mult_79_n1405,
         u5_mult_79_n1404, u5_mult_79_n1403, u5_mult_79_n1402,
         u5_mult_79_n1401, u5_mult_79_n1400, u5_mult_79_n1399,
         u5_mult_79_n1398, u5_mult_79_n1397, u5_mult_79_n1396,
         u5_mult_79_n1395, u5_mult_79_n1394, u5_mult_79_n1393,
         u5_mult_79_n1392, u5_mult_79_n1391, u5_mult_79_n1390,
         u5_mult_79_n1389, u5_mult_79_n1388, u5_mult_79_n1387,
         u5_mult_79_n1386, u5_mult_79_n1385, u5_mult_79_n1384,
         u5_mult_79_n1383, u5_mult_79_n1382, u5_mult_79_n1381,
         u5_mult_79_n1380, u5_mult_79_n1379, u5_mult_79_n1378,
         u5_mult_79_n1377, u5_mult_79_n1376, u5_mult_79_n1375,
         u5_mult_79_n1374, u5_mult_79_n1373, u5_mult_79_n1372,
         u5_mult_79_n1371, u5_mult_79_n1370, u5_mult_79_n1369,
         u5_mult_79_n1368, u5_mult_79_n1367, u5_mult_79_n1366,
         u5_mult_79_n1365, u5_mult_79_n1364, u5_mult_79_n1363,
         u5_mult_79_n1362, u5_mult_79_n1361, u5_mult_79_n1360,
         u5_mult_79_n1359, u5_mult_79_n1358, u5_mult_79_n1357,
         u5_mult_79_n1356, u5_mult_79_n1355, u5_mult_79_n1354,
         u5_mult_79_n1353, u5_mult_79_n1352, u5_mult_79_n1351,
         u5_mult_79_n1350, u5_mult_79_n1349, u5_mult_79_n1348,
         u5_mult_79_n1347, u5_mult_79_n1346, u5_mult_79_n1345,
         u5_mult_79_n1344, u5_mult_79_n1343, u5_mult_79_n1342,
         u5_mult_79_n1341, u5_mult_79_n1340, u5_mult_79_n1339,
         u5_mult_79_n1338, u5_mult_79_n1337, u5_mult_79_n1336,
         u5_mult_79_n1335, u5_mult_79_n1334, u5_mult_79_n1333,
         u5_mult_79_n1332, u5_mult_79_n1331, u5_mult_79_n1330,
         u5_mult_79_n1329, u5_mult_79_n1328, u5_mult_79_n1327,
         u5_mult_79_n1326, u5_mult_79_n1325, u5_mult_79_n1324,
         u5_mult_79_n1323, u5_mult_79_n1322, u5_mult_79_n1321,
         u5_mult_79_n1320, u5_mult_79_n1319, u5_mult_79_n1318,
         u5_mult_79_n1317, u5_mult_79_n1316, u5_mult_79_n1315,
         u5_mult_79_n1314, u5_mult_79_n1313, u5_mult_79_n1312,
         u5_mult_79_n1311, u5_mult_79_n1310, u5_mult_79_n1309,
         u5_mult_79_n1308, u5_mult_79_n1307, u5_mult_79_n1306,
         u5_mult_79_n1305, u5_mult_79_n1304, u5_mult_79_n1303,
         u5_mult_79_n1302, u5_mult_79_n1301, u5_mult_79_n1300,
         u5_mult_79_n1299, u5_mult_79_n1298, u5_mult_79_n1297,
         u5_mult_79_n1296, u5_mult_79_n1295, u5_mult_79_n1294,
         u5_mult_79_n1293, u5_mult_79_n1292, u5_mult_79_n1291,
         u5_mult_79_n1290, u5_mult_79_n1289, u5_mult_79_n1288,
         u5_mult_79_n1287, u5_mult_79_n1286, u5_mult_79_n1285,
         u5_mult_79_n1284, u5_mult_79_n1283, u5_mult_79_n1282,
         u5_mult_79_n1281, u5_mult_79_n1280, u5_mult_79_n1279,
         u5_mult_79_n1278, u5_mult_79_n1277, u5_mult_79_n1276,
         u5_mult_79_n1275, u5_mult_79_n1274, u5_mult_79_n1273,
         u5_mult_79_n1272, u5_mult_79_n1271, u5_mult_79_n1270,
         u5_mult_79_n1269, u5_mult_79_n1268, u5_mult_79_n1267,
         u5_mult_79_n1266, u5_mult_79_n1265, u5_mult_79_n1264,
         u5_mult_79_n1263, u5_mult_79_n1262, u5_mult_79_n1261,
         u5_mult_79_n1260, u5_mult_79_n1259, u5_mult_79_n1258,
         u5_mult_79_n1257, u5_mult_79_n1256, u5_mult_79_n1255,
         u5_mult_79_n1254, u5_mult_79_n1253, u5_mult_79_n1252,
         u5_mult_79_n1251, u5_mult_79_n1250, u5_mult_79_n1249,
         u5_mult_79_n1248, u5_mult_79_n1247, u5_mult_79_n1246,
         u5_mult_79_n1245, u5_mult_79_n1244, u5_mult_79_n1243,
         u5_mult_79_n1242, u5_mult_79_n1241, u5_mult_79_n1240,
         u5_mult_79_n1239, u5_mult_79_n1238, u5_mult_79_n1237,
         u5_mult_79_n1236, u5_mult_79_n1235, u5_mult_79_n1234,
         u5_mult_79_n1233, u5_mult_79_n1232, u5_mult_79_n1231,
         u5_mult_79_n1230, u5_mult_79_n1229, u5_mult_79_n1228,
         u5_mult_79_n1227, u5_mult_79_n1226, u5_mult_79_n1225,
         u5_mult_79_n1224, u5_mult_79_n1223, u5_mult_79_n1222,
         u5_mult_79_n1221, u5_mult_79_n1220, u5_mult_79_n1219,
         u5_mult_79_n1218, u5_mult_79_n1217, u5_mult_79_n1216,
         u5_mult_79_n1215, u5_mult_79_n1214, u5_mult_79_n1213,
         u5_mult_79_n1212, u5_mult_79_n1211, u5_mult_79_n1210,
         u5_mult_79_n1209, u5_mult_79_n1208, u5_mult_79_n1207,
         u5_mult_79_n1206, u5_mult_79_n1205, u5_mult_79_n1204,
         u5_mult_79_n1203, u5_mult_79_n1202, u5_mult_79_n1201,
         u5_mult_79_n1200, u5_mult_79_n1199, u5_mult_79_n1198,
         u5_mult_79_n1197, u5_mult_79_n1196, u5_mult_79_n1195,
         u5_mult_79_n1194, u5_mult_79_n1193, u5_mult_79_n1192,
         u5_mult_79_n1191, u5_mult_79_n1190, u5_mult_79_n1189,
         u5_mult_79_n1188, u5_mult_79_n1187, u5_mult_79_n1186,
         u5_mult_79_n1185, u5_mult_79_n1184, u5_mult_79_n1183,
         u5_mult_79_n1182, u5_mult_79_n1181, u5_mult_79_n1180,
         u5_mult_79_n1179, u5_mult_79_n1178, u5_mult_79_n1177,
         u5_mult_79_n1176, u5_mult_79_n1175, u5_mult_79_n1174,
         u5_mult_79_n1173, u5_mult_79_n1172, u5_mult_79_n1171,
         u5_mult_79_n1170, u5_mult_79_n1169, u5_mult_79_n1168,
         u5_mult_79_n1167, u5_mult_79_n1166, u5_mult_79_n1165,
         u5_mult_79_n1164, u5_mult_79_n1163, u5_mult_79_n1162,
         u5_mult_79_n1161, u5_mult_79_n1160, u5_mult_79_n1159,
         u5_mult_79_n1158, u5_mult_79_n1157, u5_mult_79_n1156,
         u5_mult_79_n1155, u5_mult_79_n1154, u5_mult_79_n1153,
         u5_mult_79_n1152, u5_mult_79_n1151, u5_mult_79_n1150,
         u5_mult_79_n1149, u5_mult_79_n1148, u5_mult_79_n1147,
         u5_mult_79_n1146, u5_mult_79_n1145, u5_mult_79_n1144,
         u5_mult_79_n1143, u5_mult_79_n1142, u5_mult_79_n1141,
         u5_mult_79_n1140, u5_mult_79_n1139, u5_mult_79_n1138,
         u5_mult_79_n1137, u5_mult_79_n1136, u5_mult_79_n1135,
         u5_mult_79_n1134, u5_mult_79_n1133, u5_mult_79_n1132,
         u5_mult_79_n1131, u5_mult_79_n1130, u5_mult_79_n1129,
         u5_mult_79_n1128, u5_mult_79_n1127, u5_mult_79_n1126,
         u5_mult_79_n1125, u5_mult_79_n1124, u5_mult_79_n1123,
         u5_mult_79_n1122, u5_mult_79_n1121, u5_mult_79_n1120,
         u5_mult_79_n1119, u5_mult_79_n1118, u5_mult_79_n1117,
         u5_mult_79_n1116, u5_mult_79_n1115, u5_mult_79_n1114,
         u5_mult_79_n1113, u5_mult_79_n1112, u5_mult_79_n1111,
         u5_mult_79_n1110, u5_mult_79_n1109, u5_mult_79_n1108,
         u5_mult_79_n1107, u5_mult_79_n1106, u5_mult_79_n1105,
         u5_mult_79_n1104, u5_mult_79_n1103, u5_mult_79_n1102,
         u5_mult_79_n1101, u5_mult_79_n1100, u5_mult_79_n1099,
         u5_mult_79_n1098, u5_mult_79_n1097, u5_mult_79_n1096,
         u5_mult_79_n1095, u5_mult_79_n1094, u5_mult_79_n1093,
         u5_mult_79_n1092, u5_mult_79_n1091, u5_mult_79_n1090,
         u5_mult_79_n1089, u5_mult_79_n1088, u5_mult_79_n1087,
         u5_mult_79_n1086, u5_mult_79_n1085, u5_mult_79_n1084,
         u5_mult_79_n1083, u5_mult_79_n1082, u5_mult_79_n1081,
         u5_mult_79_n1080, u5_mult_79_n1079, u5_mult_79_n1078,
         u5_mult_79_n1077, u5_mult_79_n1076, u5_mult_79_n1075,
         u5_mult_79_n1074, u5_mult_79_n1073, u5_mult_79_n1072,
         u5_mult_79_n1071, u5_mult_79_n1070, u5_mult_79_n1069,
         u5_mult_79_n1068, u5_mult_79_n1067, u5_mult_79_n1066,
         u5_mult_79_n1065, u5_mult_79_n1064, u5_mult_79_n1063,
         u5_mult_79_n1062, u5_mult_79_n1061, u5_mult_79_n1060,
         u5_mult_79_n1059, u5_mult_79_n1058, u5_mult_79_n1057,
         u5_mult_79_n1056, u5_mult_79_n1055, u5_mult_79_n1054,
         u5_mult_79_n1053, u5_mult_79_n1052, u5_mult_79_n1051,
         u5_mult_79_n1050, u5_mult_79_n1049, u5_mult_79_n1048,
         u5_mult_79_n1047, u5_mult_79_n1046, u5_mult_79_n1045,
         u5_mult_79_n1044, u5_mult_79_n1043, u5_mult_79_n1042,
         u5_mult_79_n1041, u5_mult_79_n1040, u5_mult_79_n1039,
         u5_mult_79_n1038, u5_mult_79_n1037, u5_mult_79_n1036,
         u5_mult_79_n1035, u5_mult_79_n1034, u5_mult_79_n1033,
         u5_mult_79_n1032, u5_mult_79_n1031, u5_mult_79_n1030,
         u5_mult_79_n1029, u5_mult_79_n1028, u5_mult_79_n1027,
         u5_mult_79_n1026, u5_mult_79_n1025, u5_mult_79_n1024,
         u5_mult_79_n1023, u5_mult_79_n1022, u5_mult_79_n1021,
         u5_mult_79_n1020, u5_mult_79_n1019, u5_mult_79_n1018,
         u5_mult_79_n1017, u5_mult_79_n1016, u5_mult_79_n1015,
         u5_mult_79_n1014, u5_mult_79_n1013, u5_mult_79_n1012,
         u5_mult_79_n1011, u5_mult_79_n1010, u5_mult_79_n1009,
         u5_mult_79_n1008, u5_mult_79_n1007, u5_mult_79_n1006,
         u5_mult_79_n1005, u5_mult_79_n1004, u5_mult_79_n1003,
         u5_mult_79_n1002, u5_mult_79_n1001, u5_mult_79_n1000, u5_mult_79_n999,
         u5_mult_79_n998, u5_mult_79_n997, u5_mult_79_n996, u5_mult_79_n995,
         u5_mult_79_n994, u5_mult_79_n993, u5_mult_79_n992, u5_mult_79_n991,
         u5_mult_79_n990, u5_mult_79_n989, u5_mult_79_n988, u5_mult_79_n987,
         u5_mult_79_n986, u5_mult_79_n985, u5_mult_79_n984, u5_mult_79_n983,
         u5_mult_79_n982, u5_mult_79_n981, u5_mult_79_n980, u5_mult_79_n979,
         u5_mult_79_n978, u5_mult_79_n977, u5_mult_79_n976, u5_mult_79_n975,
         u5_mult_79_n974, u5_mult_79_n973, u5_mult_79_n972, u5_mult_79_n971,
         u5_mult_79_n970, u5_mult_79_n969, u5_mult_79_n968, u5_mult_79_n967,
         u5_mult_79_n966, u5_mult_79_n965, u5_mult_79_n964, u5_mult_79_n963,
         u5_mult_79_n962, u5_mult_79_n961, u5_mult_79_n960, u5_mult_79_n959,
         u5_mult_79_n958, u5_mult_79_n957, u5_mult_79_n956, u5_mult_79_n955,
         u5_mult_79_n954, u5_mult_79_n953, u5_mult_79_n952, u5_mult_79_n951,
         u5_mult_79_n950, u5_mult_79_n949, u5_mult_79_n948, u5_mult_79_n947,
         u5_mult_79_n946, u5_mult_79_n945, u5_mult_79_n944, u5_mult_79_n943,
         u5_mult_79_n942, u5_mult_79_n941, u5_mult_79_n940, u5_mult_79_n939,
         u5_mult_79_n938, u5_mult_79_n937, u5_mult_79_n936, u5_mult_79_n935,
         u5_mult_79_n934, u5_mult_79_n933, u5_mult_79_n932, u5_mult_79_n931,
         u5_mult_79_n930, u5_mult_79_n929, u5_mult_79_n928, u5_mult_79_n927,
         u5_mult_79_n926, u5_mult_79_n925, u5_mult_79_n924, u5_mult_79_n923,
         u5_mult_79_n922, u5_mult_79_n921, u5_mult_79_n920, u5_mult_79_n919,
         u5_mult_79_n918, u5_mult_79_n917, u5_mult_79_n916, u5_mult_79_n915,
         u5_mult_79_n914, u5_mult_79_n913, u5_mult_79_n912, u5_mult_79_n911,
         u5_mult_79_n910, u5_mult_79_n909, u5_mult_79_n908, u5_mult_79_n907,
         u5_mult_79_n906, u5_mult_79_n905, u5_mult_79_n904, u5_mult_79_n903,
         u5_mult_79_n902, u5_mult_79_n901, u5_mult_79_n900, u5_mult_79_n899,
         u5_mult_79_n898, u5_mult_79_n897, u5_mult_79_n896, u5_mult_79_n895,
         u5_mult_79_n894, u5_mult_79_n893, u5_mult_79_n892, u5_mult_79_n891,
         u5_mult_79_n890, u5_mult_79_n889, u5_mult_79_n888, u5_mult_79_n887,
         u5_mult_79_n886, u5_mult_79_n885, u5_mult_79_n884, u5_mult_79_n883,
         u5_mult_79_n882, u5_mult_79_n881, u5_mult_79_n880, u5_mult_79_n879,
         u5_mult_79_n878, u5_mult_79_n877, u5_mult_79_n876, u5_mult_79_n875,
         u5_mult_79_n874, u5_mult_79_n873, u5_mult_79_n872, u5_mult_79_n871,
         u5_mult_79_n870, u5_mult_79_n869, u5_mult_79_n868, u5_mult_79_n867,
         u5_mult_79_n866, u5_mult_79_n865, u5_mult_79_n864, u5_mult_79_n863,
         u5_mult_79_n862, u5_mult_79_n861, u5_mult_79_n860, u5_mult_79_n859,
         u5_mult_79_n858, u5_mult_79_n857, u5_mult_79_n856, u5_mult_79_n855,
         u5_mult_79_n854, u5_mult_79_n853, u5_mult_79_n852, u5_mult_79_n851,
         u5_mult_79_n850, u5_mult_79_n849, u5_mult_79_n848, u5_mult_79_n847,
         u5_mult_79_n846, u5_mult_79_n845, u5_mult_79_n844, u5_mult_79_n843,
         u5_mult_79_n842, u5_mult_79_n841, u5_mult_79_n840, u5_mult_79_n839,
         u5_mult_79_n838, u5_mult_79_n837, u5_mult_79_n836, u5_mult_79_n835,
         u5_mult_79_n834, u5_mult_79_n833, u5_mult_79_n832, u5_mult_79_n831,
         u5_mult_79_n830, u5_mult_79_n829, u5_mult_79_n828, u5_mult_79_n827,
         u5_mult_79_n826, u5_mult_79_n825, u5_mult_79_n824, u5_mult_79_n823,
         u5_mult_79_n822, u5_mult_79_n821, u5_mult_79_n820, u5_mult_79_n819,
         u5_mult_79_n818, u5_mult_79_n817, u5_mult_79_n816, u5_mult_79_n815,
         u5_mult_79_n814, u5_mult_79_n813, u5_mult_79_n812, u5_mult_79_n811,
         u5_mult_79_n810, u5_mult_79_n809, u5_mult_79_n808, u5_mult_79_n807,
         u5_mult_79_n806, u5_mult_79_n805, u5_mult_79_n804, u5_mult_79_n803,
         u5_mult_79_n802, u5_mult_79_n801, u5_mult_79_n800, u5_mult_79_n799,
         u5_mult_79_n798, u5_mult_79_n797, u5_mult_79_n796, u5_mult_79_n795,
         u5_mult_79_n794, u5_mult_79_n793, u5_mult_79_n792, u5_mult_79_n791,
         u5_mult_79_n790, u5_mult_79_n789, u5_mult_79_n788, u5_mult_79_n787,
         u5_mult_79_n786, u5_mult_79_n785, u5_mult_79_n784, u5_mult_79_n783,
         u5_mult_79_n782, u5_mult_79_n781, u5_mult_79_n780, u5_mult_79_n779,
         u5_mult_79_n778, u5_mult_79_n777, u5_mult_79_n776, u5_mult_79_n775,
         u5_mult_79_n774, u5_mult_79_n773, u5_mult_79_n772, u5_mult_79_n771,
         u5_mult_79_n770, u5_mult_79_n769, u5_mult_79_n768, u5_mult_79_n767,
         u5_mult_79_n766, u5_mult_79_n765, u5_mult_79_n764, u5_mult_79_n763,
         u5_mult_79_n762, u5_mult_79_n761, u5_mult_79_n760, u5_mult_79_n759,
         u5_mult_79_n758, u5_mult_79_n757, u5_mult_79_n756, u5_mult_79_n755,
         u5_mult_79_n754, u5_mult_79_n753, u5_mult_79_n752, u5_mult_79_n751,
         u5_mult_79_n750, u5_mult_79_n749, u5_mult_79_n748, u5_mult_79_n747,
         u5_mult_79_n746, u5_mult_79_n745, u5_mult_79_n744, u5_mult_79_n743,
         u5_mult_79_n742, u5_mult_79_n741, u5_mult_79_n740, u5_mult_79_n739,
         u5_mult_79_n738, u5_mult_79_n737, u5_mult_79_n736, u5_mult_79_n735,
         u5_mult_79_n734, u5_mult_79_n733, u5_mult_79_n732, u5_mult_79_n731,
         u5_mult_79_n730, u5_mult_79_n729, u5_mult_79_n728, u5_mult_79_n727,
         u5_mult_79_n726, u5_mult_79_n725, u5_mult_79_n724, u5_mult_79_n723,
         u5_mult_79_n722, u5_mult_79_n721, u5_mult_79_n720, u5_mult_79_n719,
         u5_mult_79_n718, u5_mult_79_n717, u5_mult_79_n716, u5_mult_79_n715,
         u5_mult_79_n714, u5_mult_79_n713, u5_mult_79_n712, u5_mult_79_n711,
         u5_mult_79_n710, u5_mult_79_n709, u5_mult_79_n708, u5_mult_79_n707,
         u5_mult_79_n706, u5_mult_79_n705, u5_mult_79_n704, u5_mult_79_n703,
         u5_mult_79_n702, u5_mult_79_n701, u5_mult_79_n700, u5_mult_79_n699,
         u5_mult_79_n698, u5_mult_79_n697, u5_mult_79_n696, u5_mult_79_n695,
         u5_mult_79_n694, u5_mult_79_n693, u5_mult_79_n692, u5_mult_79_n691,
         u5_mult_79_n690, u5_mult_79_n689, u5_mult_79_n688, u5_mult_79_n687,
         u5_mult_79_n686, u5_mult_79_n685, u5_mult_79_n684, u5_mult_79_n683,
         u5_mult_79_n682, u5_mult_79_n681, u5_mult_79_n680, u5_mult_79_n679,
         u5_mult_79_n678, u5_mult_79_n677, u5_mult_79_n676, u5_mult_79_n675,
         u5_mult_79_n674, u5_mult_79_n673, u5_mult_79_n672, u5_mult_79_n671,
         u5_mult_79_n670, u5_mult_79_n669, u5_mult_79_n668, u5_mult_79_n667,
         u5_mult_79_n666, u5_mult_79_n665, u5_mult_79_n664, u5_mult_79_n663,
         u5_mult_79_n662, u5_mult_79_n661, u5_mult_79_n660, u5_mult_79_n659,
         u5_mult_79_n658, u5_mult_79_n657, u5_mult_79_n656, u5_mult_79_n655,
         u5_mult_79_n654, u5_mult_79_n653, u5_mult_79_n652, u5_mult_79_n651,
         u5_mult_79_n650, u5_mult_79_n649, u5_mult_79_n648, u5_mult_79_n647,
         u5_mult_79_n646, u5_mult_79_n645, u5_mult_79_n644, u5_mult_79_n643,
         u5_mult_79_n642, u5_mult_79_n641, u5_mult_79_n640, u5_mult_79_n639,
         u5_mult_79_n638, u5_mult_79_n637, u5_mult_79_n636, u5_mult_79_n635,
         u5_mult_79_n634, u5_mult_79_n633, u5_mult_79_n632, u5_mult_79_n631,
         u5_mult_79_n630, u5_mult_79_n629, u5_mult_79_n628, u5_mult_79_n627,
         u5_mult_79_n626, u5_mult_79_n625, u5_mult_79_n624, u5_mult_79_n623,
         u5_mult_79_n622, u5_mult_79_n621, u5_mult_79_n620, u5_mult_79_n619,
         u5_mult_79_n618, u5_mult_79_n617, u5_mult_79_n616, u5_mult_79_n615,
         u5_mult_79_n614, u5_mult_79_n613, u5_mult_79_n612, u5_mult_79_n611,
         u5_mult_79_n610, u5_mult_79_n609, u5_mult_79_n608, u5_mult_79_n607,
         u5_mult_79_n606, u5_mult_79_n605, u5_mult_79_n604, u5_mult_79_n603,
         u5_mult_79_n602, u5_mult_79_n601, u5_mult_79_n600, u5_mult_79_n599,
         u5_mult_79_n598, u5_mult_79_n597, u5_mult_79_n596, u5_mult_79_n595,
         u5_mult_79_n594, u5_mult_79_n593, u5_mult_79_n592, u5_mult_79_n591,
         u5_mult_79_n590, u5_mult_79_n589, u5_mult_79_n588, u5_mult_79_n587,
         u5_mult_79_n586, u5_mult_79_n585, u5_mult_79_n584, u5_mult_79_n583,
         u5_mult_79_n582, u5_mult_79_n581, u5_mult_79_n580, u5_mult_79_n579,
         u5_mult_79_n578, u5_mult_79_n577, u5_mult_79_n576, u5_mult_79_n575,
         u5_mult_79_n574, u5_mult_79_n573, u5_mult_79_n572, u5_mult_79_n571,
         u5_mult_79_n570, u5_mult_79_n569, u5_mult_79_n568, u5_mult_79_n567,
         u5_mult_79_n566, u5_mult_79_n565, u5_mult_79_n564, u5_mult_79_n563,
         u5_mult_79_n562, u5_mult_79_n561, u5_mult_79_n560, u5_mult_79_n559,
         u5_mult_79_n558, u5_mult_79_n557, u5_mult_79_n556, u5_mult_79_n555,
         u5_mult_79_n554, u5_mult_79_n553, u5_mult_79_n552, u5_mult_79_n551,
         u5_mult_79_n550, u5_mult_79_n549, u5_mult_79_n548, u5_mult_79_n547,
         u5_mult_79_n546, u5_mult_79_n545, u5_mult_79_n544, u5_mult_79_n543,
         u5_mult_79_n542, u5_mult_79_n541, u5_mult_79_n540, u5_mult_79_n539,
         u5_mult_79_n538, u5_mult_79_n537, u5_mult_79_n536, u5_mult_79_n535,
         u5_mult_79_n534, u5_mult_79_n533, u5_mult_79_n532, u5_mult_79_n531,
         u5_mult_79_n530, u5_mult_79_n529, u5_mult_79_n528, u5_mult_79_n527,
         u5_mult_79_n526, u5_mult_79_n525, u5_mult_79_n524, u5_mult_79_n523,
         u5_mult_79_n522, u5_mult_79_n521, u5_mult_79_n520, u5_mult_79_n519,
         u5_mult_79_n518, u5_mult_79_n517, u5_mult_79_n516, u5_mult_79_n515,
         u5_mult_79_n514, u5_mult_79_n513, u5_mult_79_n512, u5_mult_79_n511,
         u5_mult_79_n510, u5_mult_79_n509, u5_mult_79_n508, u5_mult_79_n507,
         u5_mult_79_n506, u5_mult_79_n505, u5_mult_79_n504, u5_mult_79_n503,
         u5_mult_79_n502, u5_mult_79_n501, u5_mult_79_n500, u5_mult_79_n499,
         u5_mult_79_n498, u5_mult_79_n497, u5_mult_79_n496, u5_mult_79_n495,
         u5_mult_79_n494, u5_mult_79_n493, u5_mult_79_n492, u5_mult_79_n491,
         u5_mult_79_n490, u5_mult_79_n489, u5_mult_79_n488, u5_mult_79_n487,
         u5_mult_79_n486, u5_mult_79_n485, u5_mult_79_n484, u5_mult_79_n483,
         u5_mult_79_n482, u5_mult_79_n481, u5_mult_79_n480, u5_mult_79_n479,
         u5_mult_79_n478, u5_mult_79_n477, u5_mult_79_n476, u5_mult_79_n475,
         u5_mult_79_n474, u5_mult_79_n473, u5_mult_79_n472, u5_mult_79_n471,
         u5_mult_79_n470, u5_mult_79_n469, u5_mult_79_n468, u5_mult_79_n467,
         u5_mult_79_n466, u5_mult_79_n465, u5_mult_79_n464, u5_mult_79_n463,
         u5_mult_79_n462, u5_mult_79_n461, u5_mult_79_n460, u5_mult_79_n459,
         u5_mult_79_n458, u5_mult_79_n457, u5_mult_79_n456, u5_mult_79_n455,
         u5_mult_79_n454, u5_mult_79_n453, u5_mult_79_n452, u5_mult_79_n451,
         u5_mult_79_n450, u5_mult_79_n449, u5_mult_79_n448, u5_mult_79_n447,
         u5_mult_79_n446, u5_mult_79_n445, u5_mult_79_n444, u5_mult_79_n443,
         u5_mult_79_n442, u5_mult_79_n441, u5_mult_79_n440, u5_mult_79_n439,
         u5_mult_79_n438, u5_mult_79_n437, u5_mult_79_n436, u5_mult_79_n435,
         u5_mult_79_n434, u5_mult_79_n433, u5_mult_79_n432, u5_mult_79_n431,
         u5_mult_79_n430, u5_mult_79_n429, u5_mult_79_n428, u5_mult_79_n427,
         u5_mult_79_n426, u5_mult_79_n425, u5_mult_79_n424, u5_mult_79_n423,
         u5_mult_79_n422, u5_mult_79_n421, u5_mult_79_n420, u5_mult_79_n419,
         u5_mult_79_n418, u5_mult_79_n417, u5_mult_79_n416, u5_mult_79_n415,
         u5_mult_79_n414, u5_mult_79_n413, u5_mult_79_n412, u5_mult_79_n411,
         u5_mult_79_n410, u5_mult_79_n409, u5_mult_79_n408, u5_mult_79_n407,
         u5_mult_79_n406, u5_mult_79_n405, u5_mult_79_n404, u5_mult_79_n403,
         u5_mult_79_n402, u5_mult_79_n401, u5_mult_79_n400, u5_mult_79_n399,
         u5_mult_79_n398, u5_mult_79_n397, u5_mult_79_n396, u5_mult_79_n395,
         u5_mult_79_n394, u5_mult_79_n393, u5_mult_79_n392, u5_mult_79_n391,
         u5_mult_79_n390, u5_mult_79_n389, u5_mult_79_n388, u5_mult_79_n387,
         u5_mult_79_n386, u5_mult_79_n385, u5_mult_79_n384, u5_mult_79_n383,
         u5_mult_79_n382, u5_mult_79_n381, u5_mult_79_n380, u5_mult_79_n379,
         u5_mult_79_n378, u5_mult_79_n377, u5_mult_79_n376, u5_mult_79_n375,
         u5_mult_79_n374, u5_mult_79_n373, u5_mult_79_n372, u5_mult_79_n371,
         u5_mult_79_n370, u5_mult_79_n369, u5_mult_79_n368, u5_mult_79_n367,
         u5_mult_79_n366, u5_mult_79_n365, u5_mult_79_n364, u5_mult_79_n363,
         u5_mult_79_n362, u5_mult_79_n361, u5_mult_79_n360, u5_mult_79_n359,
         u5_mult_79_n358, u5_mult_79_n357, u5_mult_79_n356, u5_mult_79_n355,
         u5_mult_79_n354, u5_mult_79_n353, u5_mult_79_n352, u5_mult_79_n351,
         u5_mult_79_n350, u5_mult_79_n349, u5_mult_79_n348, u5_mult_79_n347,
         u5_mult_79_n346, u5_mult_79_n345, u5_mult_79_n344, u5_mult_79_n343,
         u5_mult_79_n342, u5_mult_79_n341, u5_mult_79_n340, u5_mult_79_n339,
         u5_mult_79_n338, u5_mult_79_n337, u5_mult_79_n336, u5_mult_79_n335,
         u5_mult_79_n334, u5_mult_79_n333, u5_mult_79_n332, u5_mult_79_n331,
         u5_mult_79_n330, u5_mult_79_n329, u5_mult_79_n328, u5_mult_79_n327,
         u5_mult_79_n326, u5_mult_79_n325, u5_mult_79_n324, u5_mult_79_n323,
         u5_mult_79_n322, u5_mult_79_n321, u5_mult_79_n320, u5_mult_79_n319,
         u5_mult_79_n318, u5_mult_79_n317, u5_mult_79_n316, u5_mult_79_n315,
         u5_mult_79_n314, u5_mult_79_n313, u5_mult_79_n312, u5_mult_79_n311,
         u5_mult_79_n310, u5_mult_79_n309, u5_mult_79_n308, u5_mult_79_n307,
         u5_mult_79_n306, u5_mult_79_n305, u5_mult_79_n304, u5_mult_79_n303,
         u5_mult_79_n302, u5_mult_79_n301, u5_mult_79_n300, u5_mult_79_n299,
         u5_mult_79_n298, u5_mult_79_n297, u5_mult_79_n296, u5_mult_79_n295,
         u5_mult_79_n294, u5_mult_79_n293, u5_mult_79_n292, u5_mult_79_n291,
         u5_mult_79_n290, u5_mult_79_n289, u5_mult_79_n288, u5_mult_79_n287,
         u5_mult_79_n286, u5_mult_79_n285, u5_mult_79_n284, u5_mult_79_n283,
         u5_mult_79_n282, u5_mult_79_n281, u5_mult_79_n280, u5_mult_79_n279,
         u5_mult_79_n278, u5_mult_79_n277, u5_mult_79_n276, u5_mult_79_n275,
         u5_mult_79_n274, u5_mult_79_n273, u5_mult_79_n272, u5_mult_79_n271,
         u5_mult_79_n270, u5_mult_79_n269, u5_mult_79_n268, u5_mult_79_n267,
         u5_mult_79_n266, u5_mult_79_n265, u5_mult_79_n264, u5_mult_79_n263,
         u5_mult_79_n262, u5_mult_79_n261, u5_mult_79_n260, u5_mult_79_n259,
         u5_mult_79_n258, u5_mult_79_n257, u5_mult_79_n256, u5_mult_79_n255,
         u5_mult_79_n254, u5_mult_79_n253, u5_mult_79_n252, u5_mult_79_n251,
         u5_mult_79_n250, u5_mult_79_n249, u5_mult_79_n248, u5_mult_79_n247,
         u5_mult_79_n245, u5_mult_79_n244, u5_mult_79_n243, u5_mult_79_n242,
         u5_mult_79_n241, u5_mult_79_n240, u5_mult_79_n239, u5_mult_79_n238,
         u5_mult_79_n237, u5_mult_79_n236, u5_mult_79_n235, u5_mult_79_n234,
         u5_mult_79_n233, u5_mult_79_n232, u5_mult_79_n231, u5_mult_79_n230,
         u5_mult_79_n229, u5_mult_79_n228, u5_mult_79_n227, u5_mult_79_n226,
         u5_mult_79_n225, u5_mult_79_n224, u5_mult_79_n223, u5_mult_79_n222,
         u5_mult_79_n221, u5_mult_79_n220, u5_mult_79_n219, u5_mult_79_n218,
         u5_mult_79_n217, u5_mult_79_n216, u5_mult_79_n215, u5_mult_79_n214,
         u5_mult_79_n213, u5_mult_79_n212, u5_mult_79_n211, u5_mult_79_n210,
         u5_mult_79_n209, u5_mult_79_n208, u5_mult_79_n207, u5_mult_79_n206,
         u5_mult_79_n205, u5_mult_79_n204, u5_mult_79_n203, u5_mult_79_n202,
         u5_mult_79_n201, u5_mult_79_n200, u5_mult_79_n199, u5_mult_79_n198,
         u5_mult_79_n197, u5_mult_79_n196, u5_mult_79_n195, u5_mult_79_n194,
         u5_mult_79_n193, u5_mult_79_n192, u5_mult_79_n191, u5_mult_79_n190,
         u5_mult_79_n189, u5_mult_79_n188, u5_mult_79_n187, u5_mult_79_n186,
         u5_mult_79_n185, u5_mult_79_n184, u5_mult_79_n183, u5_mult_79_n182,
         u5_mult_79_n181, u5_mult_79_n180, u5_mult_79_n179, u5_mult_79_n178,
         u5_mult_79_n177, u5_mult_79_n176, u5_mult_79_n175, u5_mult_79_n174,
         u5_mult_79_n173, u5_mult_79_n172, u5_mult_79_n171, u5_mult_79_n170,
         u5_mult_79_n169, u5_mult_79_n168, u5_mult_79_n167, u5_mult_79_n166,
         u5_mult_79_n165, u5_mult_79_n164, u5_mult_79_n163, u5_mult_79_n162,
         u5_mult_79_n161, u5_mult_79_n160, u5_mult_79_n159, u5_mult_79_n158,
         u5_mult_79_n157, u5_mult_79_n156, u5_mult_79_n155, u5_mult_79_n154,
         u5_mult_79_n153, u5_mult_79_n152, u5_mult_79_n151, u5_mult_79_n150,
         u5_mult_79_n149, u5_mult_79_n148, u5_mult_79_n147, u5_mult_79_n146,
         u5_mult_79_n145, u5_mult_79_n144, u5_mult_79_n143, u5_mult_79_n142,
         u5_mult_79_n141, u5_mult_79_n140, u5_mult_79_n139, u5_mult_79_n138,
         u5_mult_79_n137, u5_mult_79_n136, u5_mult_79_n135, u5_mult_79_n134,
         u5_mult_79_n133, u5_mult_79_n132, u5_mult_79_n131, u5_mult_79_n130,
         u5_mult_79_n129, u5_mult_79_n128, u5_mult_79_n127, u5_mult_79_n126,
         u5_mult_79_n125, u5_mult_79_n124, u5_mult_79_n123, u5_mult_79_n122,
         u5_mult_79_n121, u5_mult_79_n120, u5_mult_79_n119, u5_mult_79_n118,
         u5_mult_79_n117, u5_mult_79_n116, u5_mult_79_n115, u5_mult_79_n114,
         u5_mult_79_n113, u5_mult_79_n112, u5_mult_79_n111, u5_mult_79_n110,
         u5_mult_79_n109, u5_mult_79_n108, u5_mult_79_n107, u5_mult_79_n106,
         u5_mult_79_n105, u5_mult_79_n104, u5_mult_79_n103, u5_mult_79_n102,
         u5_mult_79_n101, u5_mult_79_n100, u5_mult_79_n99, u5_mult_79_n98,
         u5_mult_79_n96, u5_mult_79_n95, u5_mult_79_n94, u5_mult_79_n93,
         u5_mult_79_n92, u5_mult_79_n91, u5_mult_79_n90, u5_mult_79_n89,
         u5_mult_79_n88, u5_mult_79_n87, u5_mult_79_n86, u5_mult_79_n85,
         u5_mult_79_n84, u5_mult_79_n83, u5_mult_79_n82, u5_mult_79_n81,
         u5_mult_79_n80, u5_mult_79_n79, u5_mult_79_n78, u5_mult_79_n77,
         u5_mult_79_n76, u5_mult_79_n75, u5_mult_79_n74, u5_mult_79_n73,
         u5_mult_79_n72, u5_mult_79_n71, u5_mult_79_n70, u5_mult_79_n69,
         u5_mult_79_n68, u5_mult_79_n67, u5_mult_79_n66, u5_mult_79_n65,
         u5_mult_79_n64, u5_mult_79_n63, u5_mult_79_n62, u5_mult_79_n61,
         u5_mult_79_n60, u5_mult_79_n59, u5_mult_79_n58, u5_mult_79_n57,
         u5_mult_79_n56, u5_mult_79_n55, u5_mult_79_n54, u5_mult_79_n53,
         u5_mult_79_n52, u5_mult_79_n51, u5_mult_79_n50, u5_mult_79_n49,
         u5_mult_79_n48, u5_mult_79_n47, u5_mult_79_n46, u5_mult_79_n45,
         u5_mult_79_n44, u5_mult_79_n43, u5_mult_79_n42, u5_mult_79_n41,
         u5_mult_79_n40, u5_mult_79_n39, u5_mult_79_n38, u5_mult_79_n37,
         u5_mult_79_n36, u5_mult_79_n35, u5_mult_79_n34, u5_mult_79_n33,
         u5_mult_79_n32, u5_mult_79_n31, u5_mult_79_n30, u5_mult_79_n29,
         u5_mult_79_n28, u5_mult_79_n27, u5_mult_79_n26, u5_mult_79_n25,
         u5_mult_79_n24, u5_mult_79_n23, u5_mult_79_n22, u5_mult_79_n21,
         u5_mult_79_n20, u5_mult_79_n19, u5_mult_79_n18, u5_mult_79_n17,
         u5_mult_79_n16, u5_mult_79_n15, u5_mult_79_n14, u5_mult_79_n13,
         u5_mult_79_n12, u5_mult_79_n11, u5_mult_79_n10, u5_mult_79_n9,
         u5_mult_79_n8, u5_mult_79_n7, u5_mult_79_n6, u5_mult_79_n5,
         u5_mult_79_n4, u5_mult_79_n3, u5_mult_79_SUMB_1__1_,
         u5_mult_79_SUMB_1__2_, u5_mult_79_SUMB_1__3_, u5_mult_79_SUMB_1__4_,
         u5_mult_79_SUMB_1__5_, u5_mult_79_SUMB_1__6_, u5_mult_79_SUMB_1__7_,
         u5_mult_79_SUMB_1__8_, u5_mult_79_SUMB_1__9_, u5_mult_79_SUMB_1__10_,
         u5_mult_79_SUMB_1__11_, u5_mult_79_SUMB_1__12_,
         u5_mult_79_SUMB_1__13_, u5_mult_79_SUMB_1__14_,
         u5_mult_79_SUMB_1__15_, u5_mult_79_SUMB_1__16_,
         u5_mult_79_SUMB_1__17_, u5_mult_79_SUMB_1__18_,
         u5_mult_79_SUMB_1__19_, u5_mult_79_SUMB_1__20_,
         u5_mult_79_SUMB_1__21_, u5_mult_79_SUMB_1__22_, u5_mult_79_SUMB_2__1_,
         u5_mult_79_SUMB_2__2_, u5_mult_79_SUMB_2__3_, u5_mult_79_SUMB_2__4_,
         u5_mult_79_SUMB_2__5_, u5_mult_79_SUMB_2__6_, u5_mult_79_SUMB_2__7_,
         u5_mult_79_SUMB_2__8_, u5_mult_79_SUMB_2__9_, u5_mult_79_SUMB_2__10_,
         u5_mult_79_SUMB_2__11_, u5_mult_79_SUMB_2__12_,
         u5_mult_79_SUMB_2__13_, u5_mult_79_SUMB_2__14_,
         u5_mult_79_SUMB_2__15_, u5_mult_79_SUMB_2__16_,
         u5_mult_79_SUMB_2__17_, u5_mult_79_SUMB_2__18_,
         u5_mult_79_SUMB_2__19_, u5_mult_79_SUMB_2__20_,
         u5_mult_79_SUMB_2__21_, u5_mult_79_SUMB_2__22_, u5_mult_79_SUMB_3__1_,
         u5_mult_79_SUMB_3__2_, u5_mult_79_SUMB_3__3_, u5_mult_79_SUMB_3__4_,
         u5_mult_79_SUMB_3__5_, u5_mult_79_SUMB_3__6_, u5_mult_79_SUMB_3__7_,
         u5_mult_79_SUMB_3__8_, u5_mult_79_SUMB_3__9_, u5_mult_79_SUMB_3__10_,
         u5_mult_79_SUMB_3__11_, u5_mult_79_SUMB_3__12_,
         u5_mult_79_SUMB_3__13_, u5_mult_79_SUMB_3__14_,
         u5_mult_79_SUMB_3__15_, u5_mult_79_SUMB_3__16_,
         u5_mult_79_SUMB_3__17_, u5_mult_79_SUMB_3__18_,
         u5_mult_79_SUMB_3__19_, u5_mult_79_SUMB_3__20_,
         u5_mult_79_SUMB_3__21_, u5_mult_79_SUMB_3__22_, u5_mult_79_SUMB_4__1_,
         u5_mult_79_SUMB_4__2_, u5_mult_79_SUMB_4__3_, u5_mult_79_SUMB_4__4_,
         u5_mult_79_SUMB_4__5_, u5_mult_79_SUMB_4__6_, u5_mult_79_SUMB_4__7_,
         u5_mult_79_SUMB_4__8_, u5_mult_79_SUMB_4__9_, u5_mult_79_SUMB_4__10_,
         u5_mult_79_SUMB_4__11_, u5_mult_79_SUMB_4__12_,
         u5_mult_79_SUMB_4__13_, u5_mult_79_SUMB_4__14_,
         u5_mult_79_SUMB_4__15_, u5_mult_79_SUMB_4__16_,
         u5_mult_79_SUMB_4__17_, u5_mult_79_SUMB_4__18_,
         u5_mult_79_SUMB_4__19_, u5_mult_79_SUMB_4__20_,
         u5_mult_79_SUMB_4__21_, u5_mult_79_SUMB_4__22_, u5_mult_79_SUMB_5__1_,
         u5_mult_79_SUMB_5__2_, u5_mult_79_SUMB_5__3_, u5_mult_79_SUMB_5__4_,
         u5_mult_79_SUMB_5__5_, u5_mult_79_SUMB_5__6_, u5_mult_79_SUMB_5__7_,
         u5_mult_79_SUMB_5__8_, u5_mult_79_SUMB_5__9_, u5_mult_79_SUMB_5__10_,
         u5_mult_79_SUMB_5__11_, u5_mult_79_SUMB_5__12_,
         u5_mult_79_SUMB_5__13_, u5_mult_79_SUMB_5__14_,
         u5_mult_79_SUMB_5__15_, u5_mult_79_SUMB_5__16_,
         u5_mult_79_SUMB_5__17_, u5_mult_79_SUMB_5__19_,
         u5_mult_79_SUMB_5__20_, u5_mult_79_SUMB_5__21_,
         u5_mult_79_SUMB_5__22_, u5_mult_79_SUMB_6__1_, u5_mult_79_SUMB_6__2_,
         u5_mult_79_SUMB_6__3_, u5_mult_79_SUMB_6__4_, u5_mult_79_SUMB_6__5_,
         u5_mult_79_SUMB_6__6_, u5_mult_79_SUMB_6__7_, u5_mult_79_SUMB_6__8_,
         u5_mult_79_SUMB_6__9_, u5_mult_79_SUMB_6__10_, u5_mult_79_SUMB_6__11_,
         u5_mult_79_SUMB_6__12_, u5_mult_79_SUMB_6__13_,
         u5_mult_79_SUMB_6__14_, u5_mult_79_SUMB_6__15_,
         u5_mult_79_SUMB_6__16_, u5_mult_79_SUMB_6__17_,
         u5_mult_79_SUMB_6__18_, u5_mult_79_SUMB_6__19_,
         u5_mult_79_SUMB_6__20_, u5_mult_79_SUMB_6__21_,
         u5_mult_79_SUMB_6__22_, u5_mult_79_SUMB_7__1_, u5_mult_79_SUMB_7__2_,
         u5_mult_79_SUMB_7__3_, u5_mult_79_SUMB_7__4_, u5_mult_79_SUMB_7__5_,
         u5_mult_79_SUMB_7__6_, u5_mult_79_SUMB_7__7_, u5_mult_79_SUMB_7__8_,
         u5_mult_79_SUMB_7__9_, u5_mult_79_SUMB_7__10_, u5_mult_79_SUMB_7__11_,
         u5_mult_79_SUMB_7__12_, u5_mult_79_SUMB_7__13_,
         u5_mult_79_SUMB_7__14_, u5_mult_79_SUMB_7__15_,
         u5_mult_79_SUMB_7__16_, u5_mult_79_SUMB_7__17_,
         u5_mult_79_SUMB_7__18_, u5_mult_79_SUMB_7__19_,
         u5_mult_79_SUMB_7__20_, u5_mult_79_SUMB_7__21_,
         u5_mult_79_SUMB_7__22_, u5_mult_79_SUMB_8__1_, u5_mult_79_SUMB_8__2_,
         u5_mult_79_SUMB_8__3_, u5_mult_79_SUMB_8__4_, u5_mult_79_SUMB_8__5_,
         u5_mult_79_SUMB_8__6_, u5_mult_79_SUMB_8__7_, u5_mult_79_SUMB_8__8_,
         u5_mult_79_SUMB_8__9_, u5_mult_79_SUMB_8__10_, u5_mult_79_SUMB_8__11_,
         u5_mult_79_SUMB_8__12_, u5_mult_79_SUMB_8__13_,
         u5_mult_79_SUMB_8__14_, u5_mult_79_SUMB_8__15_,
         u5_mult_79_SUMB_8__16_, u5_mult_79_SUMB_8__17_,
         u5_mult_79_SUMB_8__18_, u5_mult_79_SUMB_8__19_,
         u5_mult_79_SUMB_8__20_, u5_mult_79_SUMB_8__21_,
         u5_mult_79_SUMB_8__22_, u5_mult_79_SUMB_9__1_, u5_mult_79_SUMB_9__2_,
         u5_mult_79_SUMB_9__3_, u5_mult_79_SUMB_9__4_, u5_mult_79_SUMB_9__5_,
         u5_mult_79_SUMB_9__6_, u5_mult_79_SUMB_9__7_, u5_mult_79_SUMB_9__8_,
         u5_mult_79_SUMB_9__9_, u5_mult_79_SUMB_9__10_, u5_mult_79_SUMB_9__11_,
         u5_mult_79_SUMB_9__12_, u5_mult_79_SUMB_9__13_,
         u5_mult_79_SUMB_9__14_, u5_mult_79_SUMB_9__15_,
         u5_mult_79_SUMB_9__16_, u5_mult_79_SUMB_9__17_,
         u5_mult_79_SUMB_9__18_, u5_mult_79_SUMB_9__19_,
         u5_mult_79_SUMB_9__20_, u5_mult_79_SUMB_9__21_,
         u5_mult_79_SUMB_9__22_, u5_mult_79_SUMB_10__1_,
         u5_mult_79_SUMB_10__2_, u5_mult_79_SUMB_10__3_,
         u5_mult_79_SUMB_10__4_, u5_mult_79_SUMB_10__5_,
         u5_mult_79_SUMB_10__6_, u5_mult_79_SUMB_10__7_,
         u5_mult_79_SUMB_10__8_, u5_mult_79_SUMB_10__9_,
         u5_mult_79_SUMB_10__10_, u5_mult_79_SUMB_10__11_,
         u5_mult_79_SUMB_10__12_, u5_mult_79_SUMB_10__13_,
         u5_mult_79_SUMB_10__14_, u5_mult_79_SUMB_10__15_,
         u5_mult_79_SUMB_10__16_, u5_mult_79_SUMB_10__17_,
         u5_mult_79_SUMB_10__18_, u5_mult_79_SUMB_10__19_,
         u5_mult_79_SUMB_10__20_, u5_mult_79_SUMB_10__21_,
         u5_mult_79_SUMB_10__22_, u5_mult_79_SUMB_11__1_,
         u5_mult_79_SUMB_11__2_, u5_mult_79_SUMB_11__3_,
         u5_mult_79_SUMB_11__4_, u5_mult_79_SUMB_11__5_,
         u5_mult_79_SUMB_11__6_, u5_mult_79_SUMB_11__7_,
         u5_mult_79_SUMB_11__8_, u5_mult_79_SUMB_11__9_,
         u5_mult_79_SUMB_11__10_, u5_mult_79_SUMB_11__11_,
         u5_mult_79_SUMB_11__12_, u5_mult_79_SUMB_11__13_,
         u5_mult_79_SUMB_11__14_, u5_mult_79_SUMB_11__15_,
         u5_mult_79_SUMB_11__16_, u5_mult_79_SUMB_11__17_,
         u5_mult_79_SUMB_11__18_, u5_mult_79_SUMB_11__19_,
         u5_mult_79_SUMB_11__20_, u5_mult_79_SUMB_11__21_,
         u5_mult_79_SUMB_11__22_, u5_mult_79_SUMB_12__1_,
         u5_mult_79_SUMB_12__2_, u5_mult_79_SUMB_12__3_,
         u5_mult_79_SUMB_12__4_, u5_mult_79_SUMB_12__5_,
         u5_mult_79_SUMB_12__6_, u5_mult_79_SUMB_12__7_,
         u5_mult_79_SUMB_12__8_, u5_mult_79_SUMB_12__9_,
         u5_mult_79_SUMB_12__10_, u5_mult_79_SUMB_12__11_,
         u5_mult_79_SUMB_12__12_, u5_mult_79_SUMB_12__13_,
         u5_mult_79_SUMB_12__14_, u5_mult_79_SUMB_12__15_,
         u5_mult_79_SUMB_12__16_, u5_mult_79_SUMB_12__17_,
         u5_mult_79_SUMB_12__18_, u5_mult_79_SUMB_12__19_,
         u5_mult_79_SUMB_12__20_, u5_mult_79_SUMB_12__21_,
         u5_mult_79_SUMB_12__22_, u5_mult_79_SUMB_13__1_,
         u5_mult_79_SUMB_13__2_, u5_mult_79_SUMB_13__3_,
         u5_mult_79_SUMB_13__4_, u5_mult_79_SUMB_13__5_,
         u5_mult_79_SUMB_13__6_, u5_mult_79_SUMB_13__7_,
         u5_mult_79_SUMB_13__8_, u5_mult_79_SUMB_13__9_,
         u5_mult_79_SUMB_13__10_, u5_mult_79_SUMB_13__11_,
         u5_mult_79_SUMB_13__12_, u5_mult_79_SUMB_13__14_,
         u5_mult_79_SUMB_13__15_, u5_mult_79_SUMB_13__16_,
         u5_mult_79_SUMB_13__17_, u5_mult_79_SUMB_13__18_,
         u5_mult_79_SUMB_13__19_, u5_mult_79_SUMB_13__20_,
         u5_mult_79_SUMB_13__21_, u5_mult_79_SUMB_13__22_,
         u5_mult_79_SUMB_14__1_, u5_mult_79_SUMB_14__2_,
         u5_mult_79_SUMB_14__3_, u5_mult_79_SUMB_14__4_,
         u5_mult_79_SUMB_14__5_, u5_mult_79_SUMB_14__6_,
         u5_mult_79_SUMB_14__7_, u5_mult_79_SUMB_14__8_,
         u5_mult_79_SUMB_14__9_, u5_mult_79_SUMB_14__10_,
         u5_mult_79_SUMB_14__11_, u5_mult_79_SUMB_14__12_,
         u5_mult_79_SUMB_14__13_, u5_mult_79_SUMB_14__14_,
         u5_mult_79_SUMB_14__15_, u5_mult_79_SUMB_14__16_,
         u5_mult_79_SUMB_14__17_, u5_mult_79_SUMB_14__18_,
         u5_mult_79_SUMB_14__19_, u5_mult_79_SUMB_14__20_,
         u5_mult_79_SUMB_14__21_, u5_mult_79_SUMB_14__22_,
         u5_mult_79_SUMB_15__1_, u5_mult_79_SUMB_15__2_,
         u5_mult_79_SUMB_15__3_, u5_mult_79_SUMB_15__4_,
         u5_mult_79_SUMB_15__5_, u5_mult_79_SUMB_15__6_,
         u5_mult_79_SUMB_15__7_, u5_mult_79_SUMB_15__8_,
         u5_mult_79_SUMB_15__9_, u5_mult_79_SUMB_15__10_,
         u5_mult_79_SUMB_15__11_, u5_mult_79_SUMB_15__12_,
         u5_mult_79_SUMB_15__13_, u5_mult_79_SUMB_15__14_,
         u5_mult_79_SUMB_15__15_, u5_mult_79_SUMB_15__16_,
         u5_mult_79_SUMB_15__17_, u5_mult_79_SUMB_15__18_,
         u5_mult_79_SUMB_15__19_, u5_mult_79_SUMB_15__20_,
         u5_mult_79_SUMB_15__21_, u5_mult_79_SUMB_15__22_,
         u5_mult_79_SUMB_16__1_, u5_mult_79_SUMB_16__2_,
         u5_mult_79_SUMB_16__3_, u5_mult_79_SUMB_16__4_,
         u5_mult_79_SUMB_16__5_, u5_mult_79_SUMB_16__6_,
         u5_mult_79_SUMB_16__7_, u5_mult_79_SUMB_16__9_,
         u5_mult_79_SUMB_16__10_, u5_mult_79_SUMB_16__11_,
         u5_mult_79_SUMB_16__13_, u5_mult_79_SUMB_16__14_,
         u5_mult_79_SUMB_16__15_, u5_mult_79_SUMB_16__16_,
         u5_mult_79_SUMB_16__17_, u5_mult_79_SUMB_16__18_,
         u5_mult_79_SUMB_16__19_, u5_mult_79_SUMB_16__20_,
         u5_mult_79_SUMB_16__21_, u5_mult_79_SUMB_16__22_,
         u5_mult_79_SUMB_17__1_, u5_mult_79_SUMB_17__2_,
         u5_mult_79_SUMB_17__3_, u5_mult_79_SUMB_17__4_,
         u5_mult_79_SUMB_17__5_, u5_mult_79_SUMB_17__6_,
         u5_mult_79_SUMB_17__7_, u5_mult_79_SUMB_17__8_,
         u5_mult_79_SUMB_17__9_, u5_mult_79_SUMB_17__10_,
         u5_mult_79_SUMB_17__11_, u5_mult_79_SUMB_17__12_,
         u5_mult_79_SUMB_17__13_, u5_mult_79_SUMB_17__14_,
         u5_mult_79_SUMB_17__15_, u5_mult_79_SUMB_17__16_,
         u5_mult_79_SUMB_17__17_, u5_mult_79_SUMB_17__18_,
         u5_mult_79_SUMB_17__19_, u5_mult_79_SUMB_17__20_,
         u5_mult_79_SUMB_17__21_, u5_mult_79_SUMB_17__22_,
         u5_mult_79_SUMB_18__1_, u5_mult_79_SUMB_18__2_,
         u5_mult_79_SUMB_18__3_, u5_mult_79_SUMB_18__4_,
         u5_mult_79_SUMB_18__5_, u5_mult_79_SUMB_18__6_,
         u5_mult_79_SUMB_18__7_, u5_mult_79_SUMB_18__8_,
         u5_mult_79_SUMB_18__9_, u5_mult_79_SUMB_18__10_,
         u5_mult_79_SUMB_18__11_, u5_mult_79_SUMB_18__12_,
         u5_mult_79_SUMB_18__13_, u5_mult_79_SUMB_18__14_,
         u5_mult_79_SUMB_18__15_, u5_mult_79_SUMB_18__16_,
         u5_mult_79_SUMB_18__17_, u5_mult_79_SUMB_18__18_,
         u5_mult_79_SUMB_18__19_, u5_mult_79_SUMB_18__20_,
         u5_mult_79_SUMB_18__21_, u5_mult_79_SUMB_18__22_,
         u5_mult_79_SUMB_19__1_, u5_mult_79_SUMB_19__2_,
         u5_mult_79_SUMB_19__3_, u5_mult_79_SUMB_19__4_,
         u5_mult_79_SUMB_19__5_, u5_mult_79_SUMB_19__6_,
         u5_mult_79_SUMB_19__7_, u5_mult_79_SUMB_19__8_,
         u5_mult_79_SUMB_19__9_, u5_mult_79_SUMB_19__10_,
         u5_mult_79_SUMB_19__11_, u5_mult_79_SUMB_19__12_,
         u5_mult_79_SUMB_19__13_, u5_mult_79_SUMB_19__14_,
         u5_mult_79_SUMB_19__15_, u5_mult_79_SUMB_19__16_,
         u5_mult_79_SUMB_19__17_, u5_mult_79_SUMB_19__18_,
         u5_mult_79_SUMB_19__19_, u5_mult_79_SUMB_19__20_,
         u5_mult_79_SUMB_19__21_, u5_mult_79_SUMB_19__22_,
         u5_mult_79_SUMB_20__1_, u5_mult_79_SUMB_20__2_,
         u5_mult_79_SUMB_20__3_, u5_mult_79_SUMB_20__4_,
         u5_mult_79_SUMB_20__5_, u5_mult_79_SUMB_20__6_,
         u5_mult_79_SUMB_20__7_, u5_mult_79_SUMB_20__8_,
         u5_mult_79_SUMB_20__9_, u5_mult_79_SUMB_20__10_,
         u5_mult_79_SUMB_20__11_, u5_mult_79_SUMB_20__12_,
         u5_mult_79_SUMB_20__13_, u5_mult_79_SUMB_20__14_,
         u5_mult_79_SUMB_20__15_, u5_mult_79_SUMB_20__16_,
         u5_mult_79_SUMB_20__17_, u5_mult_79_SUMB_20__18_,
         u5_mult_79_SUMB_20__19_, u5_mult_79_SUMB_20__20_,
         u5_mult_79_SUMB_20__21_, u5_mult_79_SUMB_20__22_,
         u5_mult_79_SUMB_21__1_, u5_mult_79_SUMB_21__2_,
         u5_mult_79_SUMB_21__4_, u5_mult_79_SUMB_21__5_,
         u5_mult_79_SUMB_21__6_, u5_mult_79_SUMB_21__7_,
         u5_mult_79_SUMB_21__8_, u5_mult_79_SUMB_21__9_,
         u5_mult_79_SUMB_21__10_, u5_mult_79_SUMB_21__11_,
         u5_mult_79_SUMB_21__12_, u5_mult_79_SUMB_21__13_,
         u5_mult_79_SUMB_21__14_, u5_mult_79_SUMB_21__15_,
         u5_mult_79_SUMB_21__16_, u5_mult_79_SUMB_21__17_,
         u5_mult_79_SUMB_21__18_, u5_mult_79_SUMB_21__19_,
         u5_mult_79_SUMB_21__20_, u5_mult_79_SUMB_21__21_,
         u5_mult_79_SUMB_21__22_, u5_mult_79_SUMB_22__1_,
         u5_mult_79_SUMB_22__2_, u5_mult_79_SUMB_22__3_,
         u5_mult_79_SUMB_22__4_, u5_mult_79_SUMB_22__5_,
         u5_mult_79_SUMB_22__6_, u5_mult_79_SUMB_22__7_,
         u5_mult_79_SUMB_22__8_, u5_mult_79_SUMB_22__9_,
         u5_mult_79_SUMB_22__10_, u5_mult_79_SUMB_22__11_,
         u5_mult_79_SUMB_22__12_, u5_mult_79_SUMB_22__13_,
         u5_mult_79_SUMB_22__14_, u5_mult_79_SUMB_22__15_,
         u5_mult_79_SUMB_22__16_, u5_mult_79_SUMB_22__17_,
         u5_mult_79_SUMB_22__18_, u5_mult_79_SUMB_22__19_,
         u5_mult_79_SUMB_22__20_, u5_mult_79_SUMB_22__21_,
         u5_mult_79_SUMB_22__22_, u5_mult_79_SUMB_23__1_,
         u5_mult_79_SUMB_23__2_, u5_mult_79_SUMB_23__3_,
         u5_mult_79_SUMB_23__4_, u5_mult_79_SUMB_23__5_,
         u5_mult_79_SUMB_23__6_, u5_mult_79_SUMB_23__7_,
         u5_mult_79_SUMB_23__8_, u5_mult_79_SUMB_23__9_,
         u5_mult_79_SUMB_23__10_, u5_mult_79_SUMB_23__11_,
         u5_mult_79_SUMB_23__12_, u5_mult_79_SUMB_23__13_,
         u5_mult_79_SUMB_23__14_, u5_mult_79_SUMB_23__15_,
         u5_mult_79_SUMB_23__16_, u5_mult_79_SUMB_23__17_,
         u5_mult_79_SUMB_23__18_, u5_mult_79_SUMB_23__19_,
         u5_mult_79_SUMB_23__20_, u5_mult_79_SUMB_23__21_,
         u5_mult_79_SUMB_23__22_, u5_mult_79_CARRYB_1__0_,
         u5_mult_79_CARRYB_1__1_, u5_mult_79_CARRYB_1__2_,
         u5_mult_79_CARRYB_1__3_, u5_mult_79_CARRYB_1__4_,
         u5_mult_79_CARRYB_1__5_, u5_mult_79_CARRYB_1__6_,
         u5_mult_79_CARRYB_1__7_, u5_mult_79_CARRYB_1__8_,
         u5_mult_79_CARRYB_1__10_, u5_mult_79_CARRYB_1__11_,
         u5_mult_79_CARRYB_1__12_, u5_mult_79_CARRYB_1__13_,
         u5_mult_79_CARRYB_1__14_, u5_mult_79_CARRYB_1__15_,
         u5_mult_79_CARRYB_1__16_, u5_mult_79_CARRYB_1__18_,
         u5_mult_79_CARRYB_1__19_, u5_mult_79_CARRYB_1__20_,
         u5_mult_79_CARRYB_1__21_, u5_mult_79_CARRYB_1__22_,
         u5_mult_79_CARRYB_2__0_, u5_mult_79_CARRYB_2__1_,
         u5_mult_79_CARRYB_2__2_, u5_mult_79_CARRYB_2__3_,
         u5_mult_79_CARRYB_2__4_, u5_mult_79_CARRYB_2__5_,
         u5_mult_79_CARRYB_2__6_, u5_mult_79_CARRYB_2__7_,
         u5_mult_79_CARRYB_2__8_, u5_mult_79_CARRYB_2__9_,
         u5_mult_79_CARRYB_2__10_, u5_mult_79_CARRYB_2__11_,
         u5_mult_79_CARRYB_2__12_, u5_mult_79_CARRYB_2__13_,
         u5_mult_79_CARRYB_2__14_, u5_mult_79_CARRYB_2__15_,
         u5_mult_79_CARRYB_2__16_, u5_mult_79_CARRYB_2__17_,
         u5_mult_79_CARRYB_2__18_, u5_mult_79_CARRYB_2__19_,
         u5_mult_79_CARRYB_2__20_, u5_mult_79_CARRYB_2__21_,
         u5_mult_79_CARRYB_2__22_, u5_mult_79_CARRYB_3__0_,
         u5_mult_79_CARRYB_3__1_, u5_mult_79_CARRYB_3__2_,
         u5_mult_79_CARRYB_3__3_, u5_mult_79_CARRYB_3__4_,
         u5_mult_79_CARRYB_3__5_, u5_mult_79_CARRYB_3__6_,
         u5_mult_79_CARRYB_3__7_, u5_mult_79_CARRYB_3__8_,
         u5_mult_79_CARRYB_3__9_, u5_mult_79_CARRYB_3__10_,
         u5_mult_79_CARRYB_3__11_, u5_mult_79_CARRYB_3__12_,
         u5_mult_79_CARRYB_3__13_, u5_mult_79_CARRYB_3__14_,
         u5_mult_79_CARRYB_3__15_, u5_mult_79_CARRYB_3__16_,
         u5_mult_79_CARRYB_3__17_, u5_mult_79_CARRYB_3__18_,
         u5_mult_79_CARRYB_3__19_, u5_mult_79_CARRYB_3__20_,
         u5_mult_79_CARRYB_3__21_, u5_mult_79_CARRYB_3__22_,
         u5_mult_79_CARRYB_4__0_, u5_mult_79_CARRYB_4__1_,
         u5_mult_79_CARRYB_4__2_, u5_mult_79_CARRYB_4__3_,
         u5_mult_79_CARRYB_4__4_, u5_mult_79_CARRYB_4__5_,
         u5_mult_79_CARRYB_4__6_, u5_mult_79_CARRYB_4__7_,
         u5_mult_79_CARRYB_4__8_, u5_mult_79_CARRYB_4__9_,
         u5_mult_79_CARRYB_4__10_, u5_mult_79_CARRYB_4__11_,
         u5_mult_79_CARRYB_4__12_, u5_mult_79_CARRYB_4__13_,
         u5_mult_79_CARRYB_4__14_, u5_mult_79_CARRYB_4__15_,
         u5_mult_79_CARRYB_4__16_, u5_mult_79_CARRYB_4__17_,
         u5_mult_79_CARRYB_4__18_, u5_mult_79_CARRYB_4__19_,
         u5_mult_79_CARRYB_4__20_, u5_mult_79_CARRYB_4__21_,
         u5_mult_79_CARRYB_4__22_, u5_mult_79_CARRYB_5__0_,
         u5_mult_79_CARRYB_5__1_, u5_mult_79_CARRYB_5__2_,
         u5_mult_79_CARRYB_5__3_, u5_mult_79_CARRYB_5__4_,
         u5_mult_79_CARRYB_5__5_, u5_mult_79_CARRYB_5__6_,
         u5_mult_79_CARRYB_5__7_, u5_mult_79_CARRYB_5__8_,
         u5_mult_79_CARRYB_5__9_, u5_mult_79_CARRYB_5__10_,
         u5_mult_79_CARRYB_5__11_, u5_mult_79_CARRYB_5__12_,
         u5_mult_79_CARRYB_5__13_, u5_mult_79_CARRYB_5__14_,
         u5_mult_79_CARRYB_5__15_, u5_mult_79_CARRYB_5__16_,
         u5_mult_79_CARRYB_5__17_, u5_mult_79_CARRYB_5__18_,
         u5_mult_79_CARRYB_5__19_, u5_mult_79_CARRYB_5__20_,
         u5_mult_79_CARRYB_5__21_, u5_mult_79_CARRYB_5__22_,
         u5_mult_79_CARRYB_6__0_, u5_mult_79_CARRYB_6__1_,
         u5_mult_79_CARRYB_6__2_, u5_mult_79_CARRYB_6__3_,
         u5_mult_79_CARRYB_6__4_, u5_mult_79_CARRYB_6__5_,
         u5_mult_79_CARRYB_6__6_, u5_mult_79_CARRYB_6__7_,
         u5_mult_79_CARRYB_6__8_, u5_mult_79_CARRYB_6__9_,
         u5_mult_79_CARRYB_6__10_, u5_mult_79_CARRYB_6__11_,
         u5_mult_79_CARRYB_6__12_, u5_mult_79_CARRYB_6__13_,
         u5_mult_79_CARRYB_6__14_, u5_mult_79_CARRYB_6__15_,
         u5_mult_79_CARRYB_6__16_, u5_mult_79_CARRYB_6__17_,
         u5_mult_79_CARRYB_6__18_, u5_mult_79_CARRYB_6__19_,
         u5_mult_79_CARRYB_6__20_, u5_mult_79_CARRYB_6__21_,
         u5_mult_79_CARRYB_6__22_, u5_mult_79_CARRYB_7__0_,
         u5_mult_79_CARRYB_7__1_, u5_mult_79_CARRYB_7__2_,
         u5_mult_79_CARRYB_7__3_, u5_mult_79_CARRYB_7__4_,
         u5_mult_79_CARRYB_7__5_, u5_mult_79_CARRYB_7__6_,
         u5_mult_79_CARRYB_7__7_, u5_mult_79_CARRYB_7__8_,
         u5_mult_79_CARRYB_7__9_, u5_mult_79_CARRYB_7__10_,
         u5_mult_79_CARRYB_7__11_, u5_mult_79_CARRYB_7__12_,
         u5_mult_79_CARRYB_7__13_, u5_mult_79_CARRYB_7__14_,
         u5_mult_79_CARRYB_7__15_, u5_mult_79_CARRYB_7__16_,
         u5_mult_79_CARRYB_7__17_, u5_mult_79_CARRYB_7__18_,
         u5_mult_79_CARRYB_7__19_, u5_mult_79_CARRYB_7__20_,
         u5_mult_79_CARRYB_7__21_, u5_mult_79_CARRYB_7__22_,
         u5_mult_79_CARRYB_8__0_, u5_mult_79_CARRYB_8__1_,
         u5_mult_79_CARRYB_8__2_, u5_mult_79_CARRYB_8__3_,
         u5_mult_79_CARRYB_8__4_, u5_mult_79_CARRYB_8__5_,
         u5_mult_79_CARRYB_8__6_, u5_mult_79_CARRYB_8__7_,
         u5_mult_79_CARRYB_8__8_, u5_mult_79_CARRYB_8__9_,
         u5_mult_79_CARRYB_8__10_, u5_mult_79_CARRYB_8__11_,
         u5_mult_79_CARRYB_8__12_, u5_mult_79_CARRYB_8__13_,
         u5_mult_79_CARRYB_8__14_, u5_mult_79_CARRYB_8__15_,
         u5_mult_79_CARRYB_8__16_, u5_mult_79_CARRYB_8__17_,
         u5_mult_79_CARRYB_8__18_, u5_mult_79_CARRYB_8__19_,
         u5_mult_79_CARRYB_8__20_, u5_mult_79_CARRYB_8__21_,
         u5_mult_79_CARRYB_8__22_, u5_mult_79_CARRYB_9__0_,
         u5_mult_79_CARRYB_9__1_, u5_mult_79_CARRYB_9__2_,
         u5_mult_79_CARRYB_9__3_, u5_mult_79_CARRYB_9__4_,
         u5_mult_79_CARRYB_9__5_, u5_mult_79_CARRYB_9__6_,
         u5_mult_79_CARRYB_9__7_, u5_mult_79_CARRYB_9__8_,
         u5_mult_79_CARRYB_9__9_, u5_mult_79_CARRYB_9__10_,
         u5_mult_79_CARRYB_9__11_, u5_mult_79_CARRYB_9__12_,
         u5_mult_79_CARRYB_9__13_, u5_mult_79_CARRYB_9__14_,
         u5_mult_79_CARRYB_9__15_, u5_mult_79_CARRYB_9__16_,
         u5_mult_79_CARRYB_9__17_, u5_mult_79_CARRYB_9__18_,
         u5_mult_79_CARRYB_9__19_, u5_mult_79_CARRYB_9__20_,
         u5_mult_79_CARRYB_9__21_, u5_mult_79_CARRYB_9__22_,
         u5_mult_79_CARRYB_10__0_, u5_mult_79_CARRYB_10__1_,
         u5_mult_79_CARRYB_10__2_, u5_mult_79_CARRYB_10__3_,
         u5_mult_79_CARRYB_10__4_, u5_mult_79_CARRYB_10__5_,
         u5_mult_79_CARRYB_10__6_, u5_mult_79_CARRYB_10__7_,
         u5_mult_79_CARRYB_10__8_, u5_mult_79_CARRYB_10__9_,
         u5_mult_79_CARRYB_10__10_, u5_mult_79_CARRYB_10__11_,
         u5_mult_79_CARRYB_10__12_, u5_mult_79_CARRYB_10__13_,
         u5_mult_79_CARRYB_10__14_, u5_mult_79_CARRYB_10__15_,
         u5_mult_79_CARRYB_10__16_, u5_mult_79_CARRYB_10__17_,
         u5_mult_79_CARRYB_10__18_, u5_mult_79_CARRYB_10__19_,
         u5_mult_79_CARRYB_10__20_, u5_mult_79_CARRYB_10__21_,
         u5_mult_79_CARRYB_10__22_, u5_mult_79_CARRYB_11__0_,
         u5_mult_79_CARRYB_11__1_, u5_mult_79_CARRYB_11__2_,
         u5_mult_79_CARRYB_11__3_, u5_mult_79_CARRYB_11__4_,
         u5_mult_79_CARRYB_11__5_, u5_mult_79_CARRYB_11__6_,
         u5_mult_79_CARRYB_11__7_, u5_mult_79_CARRYB_11__8_,
         u5_mult_79_CARRYB_11__9_, u5_mult_79_CARRYB_11__10_,
         u5_mult_79_CARRYB_11__11_, u5_mult_79_CARRYB_11__12_,
         u5_mult_79_CARRYB_11__13_, u5_mult_79_CARRYB_11__14_,
         u5_mult_79_CARRYB_11__15_, u5_mult_79_CARRYB_11__16_,
         u5_mult_79_CARRYB_11__17_, u5_mult_79_CARRYB_11__18_,
         u5_mult_79_CARRYB_11__19_, u5_mult_79_CARRYB_11__20_,
         u5_mult_79_CARRYB_11__21_, u5_mult_79_CARRYB_11__22_,
         u5_mult_79_CARRYB_12__0_, u5_mult_79_CARRYB_12__1_,
         u5_mult_79_CARRYB_12__2_, u5_mult_79_CARRYB_12__3_,
         u5_mult_79_CARRYB_12__4_, u5_mult_79_CARRYB_12__5_,
         u5_mult_79_CARRYB_12__6_, u5_mult_79_CARRYB_12__7_,
         u5_mult_79_CARRYB_12__8_, u5_mult_79_CARRYB_12__9_,
         u5_mult_79_CARRYB_12__10_, u5_mult_79_CARRYB_12__11_,
         u5_mult_79_CARRYB_12__12_, u5_mult_79_CARRYB_12__13_,
         u5_mult_79_CARRYB_12__14_, u5_mult_79_CARRYB_12__15_,
         u5_mult_79_CARRYB_12__16_, u5_mult_79_CARRYB_12__17_,
         u5_mult_79_CARRYB_12__18_, u5_mult_79_CARRYB_12__19_,
         u5_mult_79_CARRYB_12__20_, u5_mult_79_CARRYB_12__21_,
         u5_mult_79_CARRYB_12__22_, u5_mult_79_CARRYB_13__0_,
         u5_mult_79_CARRYB_13__1_, u5_mult_79_CARRYB_13__2_,
         u5_mult_79_CARRYB_13__3_, u5_mult_79_CARRYB_13__4_,
         u5_mult_79_CARRYB_13__5_, u5_mult_79_CARRYB_13__6_,
         u5_mult_79_CARRYB_13__7_, u5_mult_79_CARRYB_13__8_,
         u5_mult_79_CARRYB_13__9_, u5_mult_79_CARRYB_13__10_,
         u5_mult_79_CARRYB_13__11_, u5_mult_79_CARRYB_13__12_,
         u5_mult_79_CARRYB_13__13_, u5_mult_79_CARRYB_13__14_,
         u5_mult_79_CARRYB_13__15_, u5_mult_79_CARRYB_13__16_,
         u5_mult_79_CARRYB_13__17_, u5_mult_79_CARRYB_13__18_,
         u5_mult_79_CARRYB_13__19_, u5_mult_79_CARRYB_13__20_,
         u5_mult_79_CARRYB_13__21_, u5_mult_79_CARRYB_13__22_,
         u5_mult_79_CARRYB_14__0_, u5_mult_79_CARRYB_14__1_,
         u5_mult_79_CARRYB_14__2_, u5_mult_79_CARRYB_14__3_,
         u5_mult_79_CARRYB_14__4_, u5_mult_79_CARRYB_14__5_,
         u5_mult_79_CARRYB_14__6_, u5_mult_79_CARRYB_14__7_,
         u5_mult_79_CARRYB_14__8_, u5_mult_79_CARRYB_14__9_,
         u5_mult_79_CARRYB_14__10_, u5_mult_79_CARRYB_14__11_,
         u5_mult_79_CARRYB_14__12_, u5_mult_79_CARRYB_14__13_,
         u5_mult_79_CARRYB_14__14_, u5_mult_79_CARRYB_14__15_,
         u5_mult_79_CARRYB_14__16_, u5_mult_79_CARRYB_14__17_,
         u5_mult_79_CARRYB_14__18_, u5_mult_79_CARRYB_14__19_,
         u5_mult_79_CARRYB_14__20_, u5_mult_79_CARRYB_14__21_,
         u5_mult_79_CARRYB_14__22_, u5_mult_79_CARRYB_15__0_,
         u5_mult_79_CARRYB_15__1_, u5_mult_79_CARRYB_15__2_,
         u5_mult_79_CARRYB_15__3_, u5_mult_79_CARRYB_15__4_,
         u5_mult_79_CARRYB_15__5_, u5_mult_79_CARRYB_15__6_,
         u5_mult_79_CARRYB_15__7_, u5_mult_79_CARRYB_15__8_,
         u5_mult_79_CARRYB_15__9_, u5_mult_79_CARRYB_15__10_,
         u5_mult_79_CARRYB_15__11_, u5_mult_79_CARRYB_15__12_,
         u5_mult_79_CARRYB_15__13_, u5_mult_79_CARRYB_15__14_,
         u5_mult_79_CARRYB_15__15_, u5_mult_79_CARRYB_15__16_,
         u5_mult_79_CARRYB_15__17_, u5_mult_79_CARRYB_15__18_,
         u5_mult_79_CARRYB_15__19_, u5_mult_79_CARRYB_15__20_,
         u5_mult_79_CARRYB_15__21_, u5_mult_79_CARRYB_15__22_,
         u5_mult_79_CARRYB_16__0_, u5_mult_79_CARRYB_16__1_,
         u5_mult_79_CARRYB_16__2_, u5_mult_79_CARRYB_16__3_,
         u5_mult_79_CARRYB_16__4_, u5_mult_79_CARRYB_16__5_,
         u5_mult_79_CARRYB_16__6_, u5_mult_79_CARRYB_16__7_,
         u5_mult_79_CARRYB_16__8_, u5_mult_79_CARRYB_16__9_,
         u5_mult_79_CARRYB_16__10_, u5_mult_79_CARRYB_16__11_,
         u5_mult_79_CARRYB_16__12_, u5_mult_79_CARRYB_16__13_,
         u5_mult_79_CARRYB_16__14_, u5_mult_79_CARRYB_16__15_,
         u5_mult_79_CARRYB_16__16_, u5_mult_79_CARRYB_16__17_,
         u5_mult_79_CARRYB_16__18_, u5_mult_79_CARRYB_16__19_,
         u5_mult_79_CARRYB_16__20_, u5_mult_79_CARRYB_16__21_,
         u5_mult_79_CARRYB_16__22_, u5_mult_79_CARRYB_17__0_,
         u5_mult_79_CARRYB_17__1_, u5_mult_79_CARRYB_17__2_,
         u5_mult_79_CARRYB_17__3_, u5_mult_79_CARRYB_17__4_,
         u5_mult_79_CARRYB_17__5_, u5_mult_79_CARRYB_17__6_,
         u5_mult_79_CARRYB_17__7_, u5_mult_79_CARRYB_17__8_,
         u5_mult_79_CARRYB_17__9_, u5_mult_79_CARRYB_17__10_,
         u5_mult_79_CARRYB_17__11_, u5_mult_79_CARRYB_17__12_,
         u5_mult_79_CARRYB_17__13_, u5_mult_79_CARRYB_17__14_,
         u5_mult_79_CARRYB_17__15_, u5_mult_79_CARRYB_17__16_,
         u5_mult_79_CARRYB_17__17_, u5_mult_79_CARRYB_17__18_,
         u5_mult_79_CARRYB_17__19_, u5_mult_79_CARRYB_17__20_,
         u5_mult_79_CARRYB_17__21_, u5_mult_79_CARRYB_17__22_,
         u5_mult_79_CARRYB_18__0_, u5_mult_79_CARRYB_18__1_,
         u5_mult_79_CARRYB_18__2_, u5_mult_79_CARRYB_18__3_,
         u5_mult_79_CARRYB_18__4_, u5_mult_79_CARRYB_18__5_,
         u5_mult_79_CARRYB_18__6_, u5_mult_79_CARRYB_18__7_,
         u5_mult_79_CARRYB_18__8_, u5_mult_79_CARRYB_18__9_,
         u5_mult_79_CARRYB_18__10_, u5_mult_79_CARRYB_18__11_,
         u5_mult_79_CARRYB_18__12_, u5_mult_79_CARRYB_18__13_,
         u5_mult_79_CARRYB_18__14_, u5_mult_79_CARRYB_18__15_,
         u5_mult_79_CARRYB_18__16_, u5_mult_79_CARRYB_18__17_,
         u5_mult_79_CARRYB_18__18_, u5_mult_79_CARRYB_18__19_,
         u5_mult_79_CARRYB_18__20_, u5_mult_79_CARRYB_18__21_,
         u5_mult_79_CARRYB_18__22_, u5_mult_79_CARRYB_19__0_,
         u5_mult_79_CARRYB_19__1_, u5_mult_79_CARRYB_19__2_,
         u5_mult_79_CARRYB_19__3_, u5_mult_79_CARRYB_19__4_,
         u5_mult_79_CARRYB_19__5_, u5_mult_79_CARRYB_19__6_,
         u5_mult_79_CARRYB_19__7_, u5_mult_79_CARRYB_19__8_,
         u5_mult_79_CARRYB_19__9_, u5_mult_79_CARRYB_19__10_,
         u5_mult_79_CARRYB_19__11_, u5_mult_79_CARRYB_19__12_,
         u5_mult_79_CARRYB_19__13_, u5_mult_79_CARRYB_19__14_,
         u5_mult_79_CARRYB_19__15_, u5_mult_79_CARRYB_19__16_,
         u5_mult_79_CARRYB_19__17_, u5_mult_79_CARRYB_19__18_,
         u5_mult_79_CARRYB_19__19_, u5_mult_79_CARRYB_19__20_,
         u5_mult_79_CARRYB_19__21_, u5_mult_79_CARRYB_19__22_,
         u5_mult_79_CARRYB_20__0_, u5_mult_79_CARRYB_20__1_,
         u5_mult_79_CARRYB_20__2_, u5_mult_79_CARRYB_20__3_,
         u5_mult_79_CARRYB_20__4_, u5_mult_79_CARRYB_20__5_,
         u5_mult_79_CARRYB_20__6_, u5_mult_79_CARRYB_20__7_,
         u5_mult_79_CARRYB_20__8_, u5_mult_79_CARRYB_20__9_,
         u5_mult_79_CARRYB_20__10_, u5_mult_79_CARRYB_20__11_,
         u5_mult_79_CARRYB_20__12_, u5_mult_79_CARRYB_20__13_,
         u5_mult_79_CARRYB_20__14_, u5_mult_79_CARRYB_20__15_,
         u5_mult_79_CARRYB_20__16_, u5_mult_79_CARRYB_20__17_,
         u5_mult_79_CARRYB_20__18_, u5_mult_79_CARRYB_20__19_,
         u5_mult_79_CARRYB_20__20_, u5_mult_79_CARRYB_20__21_,
         u5_mult_79_CARRYB_20__22_, u5_mult_79_CARRYB_21__0_,
         u5_mult_79_CARRYB_21__1_, u5_mult_79_CARRYB_21__2_,
         u5_mult_79_CARRYB_21__3_, u5_mult_79_CARRYB_21__4_,
         u5_mult_79_CARRYB_21__5_, u5_mult_79_CARRYB_21__6_,
         u5_mult_79_CARRYB_21__7_, u5_mult_79_CARRYB_21__8_,
         u5_mult_79_CARRYB_21__9_, u5_mult_79_CARRYB_21__10_,
         u5_mult_79_CARRYB_21__11_, u5_mult_79_CARRYB_21__12_,
         u5_mult_79_CARRYB_21__13_, u5_mult_79_CARRYB_21__14_,
         u5_mult_79_CARRYB_21__15_, u5_mult_79_CARRYB_21__16_,
         u5_mult_79_CARRYB_21__17_, u5_mult_79_CARRYB_21__18_,
         u5_mult_79_CARRYB_21__19_, u5_mult_79_CARRYB_21__20_,
         u5_mult_79_CARRYB_21__21_, u5_mult_79_CARRYB_21__22_,
         u5_mult_79_CARRYB_22__0_, u5_mult_79_CARRYB_22__1_,
         u5_mult_79_CARRYB_22__2_, u5_mult_79_CARRYB_22__3_,
         u5_mult_79_CARRYB_22__4_, u5_mult_79_CARRYB_22__5_,
         u5_mult_79_CARRYB_22__6_, u5_mult_79_CARRYB_22__7_,
         u5_mult_79_CARRYB_22__8_, u5_mult_79_CARRYB_22__9_,
         u5_mult_79_CARRYB_22__10_, u5_mult_79_CARRYB_22__11_,
         u5_mult_79_CARRYB_22__12_, u5_mult_79_CARRYB_22__13_,
         u5_mult_79_CARRYB_22__14_, u5_mult_79_CARRYB_22__15_,
         u5_mult_79_CARRYB_22__16_, u5_mult_79_CARRYB_22__17_,
         u5_mult_79_CARRYB_22__18_, u5_mult_79_CARRYB_22__19_,
         u5_mult_79_CARRYB_22__20_, u5_mult_79_CARRYB_22__21_,
         u5_mult_79_CARRYB_22__22_, u5_mult_79_CARRYB_23__0_,
         u5_mult_79_CARRYB_23__1_, u5_mult_79_CARRYB_23__2_,
         u5_mult_79_CARRYB_23__3_, u5_mult_79_CARRYB_23__4_,
         u5_mult_79_CARRYB_23__5_, u5_mult_79_CARRYB_23__6_,
         u5_mult_79_CARRYB_23__7_, u5_mult_79_CARRYB_23__8_,
         u5_mult_79_CARRYB_23__9_, u5_mult_79_CARRYB_23__10_,
         u5_mult_79_CARRYB_23__11_, u5_mult_79_CARRYB_23__12_,
         u5_mult_79_CARRYB_23__13_, u5_mult_79_CARRYB_23__14_,
         u5_mult_79_CARRYB_23__15_, u5_mult_79_CARRYB_23__16_,
         u5_mult_79_CARRYB_23__17_, u5_mult_79_CARRYB_23__18_,
         u5_mult_79_CARRYB_23__19_, u5_mult_79_CARRYB_23__20_,
         u5_mult_79_CARRYB_23__21_, u5_mult_79_CARRYB_23__22_,
         u5_mult_79_ab_0__1_, u5_mult_79_ab_0__2_, u5_mult_79_ab_0__3_,
         u5_mult_79_ab_0__4_, u5_mult_79_ab_0__5_, u5_mult_79_ab_0__6_,
         u5_mult_79_ab_0__7_, u5_mult_79_ab_0__8_, u5_mult_79_ab_0__9_,
         u5_mult_79_ab_0__10_, u5_mult_79_ab_0__11_, u5_mult_79_ab_0__12_,
         u5_mult_79_ab_0__13_, u5_mult_79_ab_0__14_, u5_mult_79_ab_0__15_,
         u5_mult_79_ab_0__16_, u5_mult_79_ab_0__17_, u5_mult_79_ab_0__18_,
         u5_mult_79_ab_0__19_, u5_mult_79_ab_0__20_, u5_mult_79_ab_0__21_,
         u5_mult_79_ab_0__22_, u5_mult_79_ab_1__0_, u5_mult_79_ab_1__1_,
         u5_mult_79_ab_1__2_, u5_mult_79_ab_1__3_, u5_mult_79_ab_1__4_,
         u5_mult_79_ab_1__5_, u5_mult_79_ab_1__6_, u5_mult_79_ab_1__7_,
         u5_mult_79_ab_1__8_, u5_mult_79_ab_1__9_, u5_mult_79_ab_1__10_,
         u5_mult_79_ab_1__11_, u5_mult_79_ab_1__12_, u5_mult_79_ab_1__13_,
         u5_mult_79_ab_1__14_, u5_mult_79_ab_1__15_, u5_mult_79_ab_1__16_,
         u5_mult_79_ab_1__17_, u5_mult_79_ab_1__18_, u5_mult_79_ab_1__19_,
         u5_mult_79_ab_1__20_, u5_mult_79_ab_1__21_, u5_mult_79_ab_1__22_,
         u5_mult_79_ab_1__23_, u5_mult_79_ab_2__0_, u5_mult_79_ab_2__1_,
         u5_mult_79_ab_2__2_, u5_mult_79_ab_2__3_, u5_mult_79_ab_2__4_,
         u5_mult_79_ab_2__5_, u5_mult_79_ab_2__6_, u5_mult_79_ab_2__7_,
         u5_mult_79_ab_2__8_, u5_mult_79_ab_2__9_, u5_mult_79_ab_2__10_,
         u5_mult_79_ab_2__11_, u5_mult_79_ab_2__12_, u5_mult_79_ab_2__13_,
         u5_mult_79_ab_2__14_, u5_mult_79_ab_2__15_, u5_mult_79_ab_2__16_,
         u5_mult_79_ab_2__17_, u5_mult_79_ab_2__18_, u5_mult_79_ab_2__19_,
         u5_mult_79_ab_2__20_, u5_mult_79_ab_2__21_, u5_mult_79_ab_2__22_,
         u5_mult_79_ab_2__23_, u5_mult_79_ab_3__0_, u5_mult_79_ab_3__1_,
         u5_mult_79_ab_3__2_, u5_mult_79_ab_3__3_, u5_mult_79_ab_3__4_,
         u5_mult_79_ab_3__5_, u5_mult_79_ab_3__6_, u5_mult_79_ab_3__7_,
         u5_mult_79_ab_3__8_, u5_mult_79_ab_3__9_, u5_mult_79_ab_3__10_,
         u5_mult_79_ab_3__11_, u5_mult_79_ab_3__12_, u5_mult_79_ab_3__13_,
         u5_mult_79_ab_3__14_, u5_mult_79_ab_3__15_, u5_mult_79_ab_3__16_,
         u5_mult_79_ab_3__17_, u5_mult_79_ab_3__18_, u5_mult_79_ab_3__19_,
         u5_mult_79_ab_3__20_, u5_mult_79_ab_3__21_, u5_mult_79_ab_3__22_,
         u5_mult_79_ab_3__23_, u5_mult_79_ab_4__0_, u5_mult_79_ab_4__1_,
         u5_mult_79_ab_4__2_, u5_mult_79_ab_4__3_, u5_mult_79_ab_4__4_,
         u5_mult_79_ab_4__5_, u5_mult_79_ab_4__6_, u5_mult_79_ab_4__7_,
         u5_mult_79_ab_4__8_, u5_mult_79_ab_4__9_, u5_mult_79_ab_4__10_,
         u5_mult_79_ab_4__11_, u5_mult_79_ab_4__12_, u5_mult_79_ab_4__13_,
         u5_mult_79_ab_4__14_, u5_mult_79_ab_4__15_, u5_mult_79_ab_4__16_,
         u5_mult_79_ab_4__17_, u5_mult_79_ab_4__18_, u5_mult_79_ab_4__19_,
         u5_mult_79_ab_4__20_, u5_mult_79_ab_4__21_, u5_mult_79_ab_4__22_,
         u5_mult_79_ab_4__23_, u5_mult_79_ab_5__0_, u5_mult_79_ab_5__1_,
         u5_mult_79_ab_5__2_, u5_mult_79_ab_5__3_, u5_mult_79_ab_5__4_,
         u5_mult_79_ab_5__5_, u5_mult_79_ab_5__6_, u5_mult_79_ab_5__7_,
         u5_mult_79_ab_5__8_, u5_mult_79_ab_5__9_, u5_mult_79_ab_5__10_,
         u5_mult_79_ab_5__11_, u5_mult_79_ab_5__12_, u5_mult_79_ab_5__13_,
         u5_mult_79_ab_5__14_, u5_mult_79_ab_5__15_, u5_mult_79_ab_5__16_,
         u5_mult_79_ab_5__17_, u5_mult_79_ab_5__18_, u5_mult_79_ab_5__19_,
         u5_mult_79_ab_5__20_, u5_mult_79_ab_5__21_, u5_mult_79_ab_5__22_,
         u5_mult_79_ab_5__23_, u5_mult_79_ab_6__0_, u5_mult_79_ab_6__1_,
         u5_mult_79_ab_6__2_, u5_mult_79_ab_6__3_, u5_mult_79_ab_6__4_,
         u5_mult_79_ab_6__5_, u5_mult_79_ab_6__6_, u5_mult_79_ab_6__7_,
         u5_mult_79_ab_6__8_, u5_mult_79_ab_6__9_, u5_mult_79_ab_6__10_,
         u5_mult_79_ab_6__11_, u5_mult_79_ab_6__12_, u5_mult_79_ab_6__13_,
         u5_mult_79_ab_6__14_, u5_mult_79_ab_6__15_, u5_mult_79_ab_6__16_,
         u5_mult_79_ab_6__17_, u5_mult_79_ab_6__18_, u5_mult_79_ab_6__19_,
         u5_mult_79_ab_6__20_, u5_mult_79_ab_6__21_, u5_mult_79_ab_6__22_,
         u5_mult_79_ab_6__23_, u5_mult_79_ab_7__0_, u5_mult_79_ab_7__1_,
         u5_mult_79_ab_7__2_, u5_mult_79_ab_7__3_, u5_mult_79_ab_7__4_,
         u5_mult_79_ab_7__5_, u5_mult_79_ab_7__6_, u5_mult_79_ab_7__7_,
         u5_mult_79_ab_7__8_, u5_mult_79_ab_7__9_, u5_mult_79_ab_7__10_,
         u5_mult_79_ab_7__11_, u5_mult_79_ab_7__12_, u5_mult_79_ab_7__13_,
         u5_mult_79_ab_7__14_, u5_mult_79_ab_7__15_, u5_mult_79_ab_7__16_,
         u5_mult_79_ab_7__17_, u5_mult_79_ab_7__18_, u5_mult_79_ab_7__19_,
         u5_mult_79_ab_7__20_, u5_mult_79_ab_7__21_, u5_mult_79_ab_7__22_,
         u5_mult_79_ab_7__23_, u5_mult_79_ab_8__0_, u5_mult_79_ab_8__1_,
         u5_mult_79_ab_8__2_, u5_mult_79_ab_8__3_, u5_mult_79_ab_8__4_,
         u5_mult_79_ab_8__5_, u5_mult_79_ab_8__6_, u5_mult_79_ab_8__7_,
         u5_mult_79_ab_8__8_, u5_mult_79_ab_8__9_, u5_mult_79_ab_8__10_,
         u5_mult_79_ab_8__11_, u5_mult_79_ab_8__12_, u5_mult_79_ab_8__13_,
         u5_mult_79_ab_8__14_, u5_mult_79_ab_8__15_, u5_mult_79_ab_8__16_,
         u5_mult_79_ab_8__17_, u5_mult_79_ab_8__18_, u5_mult_79_ab_8__19_,
         u5_mult_79_ab_8__20_, u5_mult_79_ab_8__21_, u5_mult_79_ab_8__22_,
         u5_mult_79_ab_8__23_, u5_mult_79_ab_9__0_, u5_mult_79_ab_9__1_,
         u5_mult_79_ab_9__2_, u5_mult_79_ab_9__3_, u5_mult_79_ab_9__4_,
         u5_mult_79_ab_9__5_, u5_mult_79_ab_9__6_, u5_mult_79_ab_9__7_,
         u5_mult_79_ab_9__8_, u5_mult_79_ab_9__9_, u5_mult_79_ab_9__10_,
         u5_mult_79_ab_9__11_, u5_mult_79_ab_9__12_, u5_mult_79_ab_9__13_,
         u5_mult_79_ab_9__14_, u5_mult_79_ab_9__15_, u5_mult_79_ab_9__16_,
         u5_mult_79_ab_9__17_, u5_mult_79_ab_9__18_, u5_mult_79_ab_9__19_,
         u5_mult_79_ab_9__20_, u5_mult_79_ab_9__21_, u5_mult_79_ab_9__22_,
         u5_mult_79_ab_9__23_, u5_mult_79_ab_10__0_, u5_mult_79_ab_10__1_,
         u5_mult_79_ab_10__2_, u5_mult_79_ab_10__3_, u5_mult_79_ab_10__4_,
         u5_mult_79_ab_10__5_, u5_mult_79_ab_10__6_, u5_mult_79_ab_10__7_,
         u5_mult_79_ab_10__8_, u5_mult_79_ab_10__9_, u5_mult_79_ab_10__10_,
         u5_mult_79_ab_10__11_, u5_mult_79_ab_10__12_, u5_mult_79_ab_10__13_,
         u5_mult_79_ab_10__14_, u5_mult_79_ab_10__15_, u5_mult_79_ab_10__16_,
         u5_mult_79_ab_10__17_, u5_mult_79_ab_10__18_, u5_mult_79_ab_10__19_,
         u5_mult_79_ab_10__20_, u5_mult_79_ab_10__21_, u5_mult_79_ab_10__22_,
         u5_mult_79_ab_10__23_, u5_mult_79_ab_11__0_, u5_mult_79_ab_11__1_,
         u5_mult_79_ab_11__2_, u5_mult_79_ab_11__3_, u5_mult_79_ab_11__4_,
         u5_mult_79_ab_11__5_, u5_mult_79_ab_11__6_, u5_mult_79_ab_11__7_,
         u5_mult_79_ab_11__8_, u5_mult_79_ab_11__9_, u5_mult_79_ab_11__10_,
         u5_mult_79_ab_11__11_, u5_mult_79_ab_11__12_, u5_mult_79_ab_11__13_,
         u5_mult_79_ab_11__14_, u5_mult_79_ab_11__15_, u5_mult_79_ab_11__16_,
         u5_mult_79_ab_11__17_, u5_mult_79_ab_11__18_, u5_mult_79_ab_11__19_,
         u5_mult_79_ab_11__20_, u5_mult_79_ab_11__21_, u5_mult_79_ab_11__22_,
         u5_mult_79_ab_11__23_, u5_mult_79_ab_12__0_, u5_mult_79_ab_12__1_,
         u5_mult_79_ab_12__2_, u5_mult_79_ab_12__3_, u5_mult_79_ab_12__4_,
         u5_mult_79_ab_12__5_, u5_mult_79_ab_12__6_, u5_mult_79_ab_12__7_,
         u5_mult_79_ab_12__8_, u5_mult_79_ab_12__9_, u5_mult_79_ab_12__10_,
         u5_mult_79_ab_12__11_, u5_mult_79_ab_12__12_, u5_mult_79_ab_12__13_,
         u5_mult_79_ab_12__14_, u5_mult_79_ab_12__15_, u5_mult_79_ab_12__16_,
         u5_mult_79_ab_12__17_, u5_mult_79_ab_12__18_, u5_mult_79_ab_12__19_,
         u5_mult_79_ab_12__20_, u5_mult_79_ab_12__21_, u5_mult_79_ab_12__22_,
         u5_mult_79_ab_12__23_, u5_mult_79_ab_13__0_, u5_mult_79_ab_13__1_,
         u5_mult_79_ab_13__2_, u5_mult_79_ab_13__3_, u5_mult_79_ab_13__4_,
         u5_mult_79_ab_13__5_, u5_mult_79_ab_13__6_, u5_mult_79_ab_13__7_,
         u5_mult_79_ab_13__8_, u5_mult_79_ab_13__9_, u5_mult_79_ab_13__10_,
         u5_mult_79_ab_13__11_, u5_mult_79_ab_13__12_, u5_mult_79_ab_13__13_,
         u5_mult_79_ab_13__14_, u5_mult_79_ab_13__15_, u5_mult_79_ab_13__16_,
         u5_mult_79_ab_13__17_, u5_mult_79_ab_13__18_, u5_mult_79_ab_13__19_,
         u5_mult_79_ab_13__20_, u5_mult_79_ab_13__21_, u5_mult_79_ab_13__22_,
         u5_mult_79_ab_13__23_, u5_mult_79_ab_14__0_, u5_mult_79_ab_14__1_,
         u5_mult_79_ab_14__2_, u5_mult_79_ab_14__3_, u5_mult_79_ab_14__4_,
         u5_mult_79_ab_14__5_, u5_mult_79_ab_14__6_, u5_mult_79_ab_14__7_,
         u5_mult_79_ab_14__8_, u5_mult_79_ab_14__9_, u5_mult_79_ab_14__10_,
         u5_mult_79_ab_14__11_, u5_mult_79_ab_14__12_, u5_mult_79_ab_14__13_,
         u5_mult_79_ab_14__14_, u5_mult_79_ab_14__15_, u5_mult_79_ab_14__16_,
         u5_mult_79_ab_14__17_, u5_mult_79_ab_14__18_, u5_mult_79_ab_14__19_,
         u5_mult_79_ab_14__20_, u5_mult_79_ab_14__21_, u5_mult_79_ab_14__22_,
         u5_mult_79_ab_14__23_, u5_mult_79_ab_15__0_, u5_mult_79_ab_15__1_,
         u5_mult_79_ab_15__2_, u5_mult_79_ab_15__3_, u5_mult_79_ab_15__4_,
         u5_mult_79_ab_15__5_, u5_mult_79_ab_15__6_, u5_mult_79_ab_15__7_,
         u5_mult_79_ab_15__8_, u5_mult_79_ab_15__9_, u5_mult_79_ab_15__10_,
         u5_mult_79_ab_15__11_, u5_mult_79_ab_15__12_, u5_mult_79_ab_15__13_,
         u5_mult_79_ab_15__14_, u5_mult_79_ab_15__15_, u5_mult_79_ab_15__16_,
         u5_mult_79_ab_15__17_, u5_mult_79_ab_15__18_, u5_mult_79_ab_15__19_,
         u5_mult_79_ab_15__20_, u5_mult_79_ab_15__21_, u5_mult_79_ab_15__22_,
         u5_mult_79_ab_15__23_, u5_mult_79_ab_16__0_, u5_mult_79_ab_16__1_,
         u5_mult_79_ab_16__2_, u5_mult_79_ab_16__3_, u5_mult_79_ab_16__4_,
         u5_mult_79_ab_16__5_, u5_mult_79_ab_16__6_, u5_mult_79_ab_16__7_,
         u5_mult_79_ab_16__8_, u5_mult_79_ab_16__9_, u5_mult_79_ab_16__10_,
         u5_mult_79_ab_16__11_, u5_mult_79_ab_16__12_, u5_mult_79_ab_16__13_,
         u5_mult_79_ab_16__14_, u5_mult_79_ab_16__15_, u5_mult_79_ab_16__16_,
         u5_mult_79_ab_16__17_, u5_mult_79_ab_16__18_, u5_mult_79_ab_16__19_,
         u5_mult_79_ab_16__20_, u5_mult_79_ab_16__21_, u5_mult_79_ab_16__22_,
         u5_mult_79_ab_16__23_, u5_mult_79_ab_17__0_, u5_mult_79_ab_17__1_,
         u5_mult_79_ab_17__2_, u5_mult_79_ab_17__3_, u5_mult_79_ab_17__4_,
         u5_mult_79_ab_17__5_, u5_mult_79_ab_17__6_, u5_mult_79_ab_17__7_,
         u5_mult_79_ab_17__8_, u5_mult_79_ab_17__9_, u5_mult_79_ab_17__10_,
         u5_mult_79_ab_17__11_, u5_mult_79_ab_17__12_, u5_mult_79_ab_17__13_,
         u5_mult_79_ab_17__14_, u5_mult_79_ab_17__15_, u5_mult_79_ab_17__16_,
         u5_mult_79_ab_17__17_, u5_mult_79_ab_17__18_, u5_mult_79_ab_17__19_,
         u5_mult_79_ab_17__20_, u5_mult_79_ab_17__21_, u5_mult_79_ab_17__22_,
         u5_mult_79_ab_17__23_, u5_mult_79_ab_18__0_, u5_mult_79_ab_18__1_,
         u5_mult_79_ab_18__2_, u5_mult_79_ab_18__3_, u5_mult_79_ab_18__4_,
         u5_mult_79_ab_18__5_, u5_mult_79_ab_18__6_, u5_mult_79_ab_18__7_,
         u5_mult_79_ab_18__8_, u5_mult_79_ab_18__9_, u5_mult_79_ab_18__10_,
         u5_mult_79_ab_18__11_, u5_mult_79_ab_18__12_, u5_mult_79_ab_18__13_,
         u5_mult_79_ab_18__14_, u5_mult_79_ab_18__15_, u5_mult_79_ab_18__16_,
         u5_mult_79_ab_18__17_, u5_mult_79_ab_18__18_, u5_mult_79_ab_18__19_,
         u5_mult_79_ab_18__20_, u5_mult_79_ab_18__21_, u5_mult_79_ab_18__22_,
         u5_mult_79_ab_18__23_, u5_mult_79_ab_19__0_, u5_mult_79_ab_19__1_,
         u5_mult_79_ab_19__2_, u5_mult_79_ab_19__3_, u5_mult_79_ab_19__4_,
         u5_mult_79_ab_19__5_, u5_mult_79_ab_19__6_, u5_mult_79_ab_19__7_,
         u5_mult_79_ab_19__8_, u5_mult_79_ab_19__9_, u5_mult_79_ab_19__10_,
         u5_mult_79_ab_19__11_, u5_mult_79_ab_19__12_, u5_mult_79_ab_19__13_,
         u5_mult_79_ab_19__14_, u5_mult_79_ab_19__15_, u5_mult_79_ab_19__16_,
         u5_mult_79_ab_19__17_, u5_mult_79_ab_19__18_, u5_mult_79_ab_19__19_,
         u5_mult_79_ab_19__20_, u5_mult_79_ab_19__21_, u5_mult_79_ab_19__22_,
         u5_mult_79_ab_19__23_, u5_mult_79_ab_20__0_, u5_mult_79_ab_20__1_,
         u5_mult_79_ab_20__2_, u5_mult_79_ab_20__3_, u5_mult_79_ab_20__4_,
         u5_mult_79_ab_20__5_, u5_mult_79_ab_20__6_, u5_mult_79_ab_20__7_,
         u5_mult_79_ab_20__8_, u5_mult_79_ab_20__9_, u5_mult_79_ab_20__10_,
         u5_mult_79_ab_20__11_, u5_mult_79_ab_20__12_, u5_mult_79_ab_20__13_,
         u5_mult_79_ab_20__14_, u5_mult_79_ab_20__15_, u5_mult_79_ab_20__16_,
         u5_mult_79_ab_20__17_, u5_mult_79_ab_20__18_, u5_mult_79_ab_20__19_,
         u5_mult_79_ab_20__20_, u5_mult_79_ab_20__21_, u5_mult_79_ab_20__22_,
         u5_mult_79_ab_20__23_, u5_mult_79_ab_21__0_, u5_mult_79_ab_21__1_,
         u5_mult_79_ab_21__2_, u5_mult_79_ab_21__3_, u5_mult_79_ab_21__4_,
         u5_mult_79_ab_21__5_, u5_mult_79_ab_21__6_, u5_mult_79_ab_21__7_,
         u5_mult_79_ab_21__8_, u5_mult_79_ab_21__9_, u5_mult_79_ab_21__10_,
         u5_mult_79_ab_21__11_, u5_mult_79_ab_21__12_, u5_mult_79_ab_21__13_,
         u5_mult_79_ab_21__14_, u5_mult_79_ab_21__15_, u5_mult_79_ab_21__16_,
         u5_mult_79_ab_21__17_, u5_mult_79_ab_21__18_, u5_mult_79_ab_21__19_,
         u5_mult_79_ab_21__20_, u5_mult_79_ab_21__21_, u5_mult_79_ab_21__22_,
         u5_mult_79_ab_21__23_, u5_mult_79_ab_22__0_, u5_mult_79_ab_22__1_,
         u5_mult_79_ab_22__2_, u5_mult_79_ab_22__3_, u5_mult_79_ab_22__4_,
         u5_mult_79_ab_22__5_, u5_mult_79_ab_22__6_, u5_mult_79_ab_22__7_,
         u5_mult_79_ab_22__8_, u5_mult_79_ab_22__9_, u5_mult_79_ab_22__10_,
         u5_mult_79_ab_22__11_, u5_mult_79_ab_22__12_, u5_mult_79_ab_22__13_,
         u5_mult_79_ab_22__14_, u5_mult_79_ab_22__15_, u5_mult_79_ab_22__16_,
         u5_mult_79_ab_22__17_, u5_mult_79_ab_22__18_, u5_mult_79_ab_22__19_,
         u5_mult_79_ab_22__20_, u5_mult_79_ab_22__21_, u5_mult_79_ab_22__22_,
         u5_mult_79_ab_22__23_, u5_mult_79_ab_23__0_, u5_mult_79_ab_23__1_,
         u5_mult_79_ab_23__2_, u5_mult_79_ab_23__3_, u5_mult_79_ab_23__4_,
         u5_mult_79_ab_23__5_, u5_mult_79_ab_23__6_, u5_mult_79_ab_23__7_,
         u5_mult_79_ab_23__8_, u5_mult_79_ab_23__9_, u5_mult_79_ab_23__10_,
         u5_mult_79_ab_23__11_, u5_mult_79_ab_23__12_, u5_mult_79_ab_23__13_,
         u5_mult_79_ab_23__14_, u5_mult_79_ab_23__15_, u5_mult_79_ab_23__16_,
         u5_mult_79_ab_23__17_, u5_mult_79_ab_23__18_, u5_mult_79_ab_23__19_,
         u5_mult_79_ab_23__20_, u5_mult_79_ab_23__21_, u5_mult_79_ab_23__22_,
         u5_mult_79_ab_23__23_, u5_mult_79_FS_1_n285, u5_mult_79_FS_1_n284,
         u5_mult_79_FS_1_n283, u5_mult_79_FS_1_n282, u5_mult_79_FS_1_n281,
         u5_mult_79_FS_1_n280, u5_mult_79_FS_1_n279, u5_mult_79_FS_1_n278,
         u5_mult_79_FS_1_n277, u5_mult_79_FS_1_n276, u5_mult_79_FS_1_n275,
         u5_mult_79_FS_1_n274, u5_mult_79_FS_1_n273, u5_mult_79_FS_1_n272,
         u5_mult_79_FS_1_n271, u5_mult_79_FS_1_n270, u5_mult_79_FS_1_n269,
         u5_mult_79_FS_1_n268, u5_mult_79_FS_1_n267, u5_mult_79_FS_1_n266,
         u5_mult_79_FS_1_n265, u5_mult_79_FS_1_n264, u5_mult_79_FS_1_n263,
         u5_mult_79_FS_1_n262, u5_mult_79_FS_1_n261, u5_mult_79_FS_1_n260,
         u5_mult_79_FS_1_n259, u5_mult_79_FS_1_n258, u5_mult_79_FS_1_n257,
         u5_mult_79_FS_1_n256, u5_mult_79_FS_1_n255, u5_mult_79_FS_1_n254,
         u5_mult_79_FS_1_n253, u5_mult_79_FS_1_n252, u5_mult_79_FS_1_n251,
         u5_mult_79_FS_1_n250, u5_mult_79_FS_1_n249, u5_mult_79_FS_1_n248,
         u5_mult_79_FS_1_n247, u5_mult_79_FS_1_n246, u5_mult_79_FS_1_n245,
         u5_mult_79_FS_1_n244, u5_mult_79_FS_1_n243, u5_mult_79_FS_1_n242,
         u5_mult_79_FS_1_n241, u5_mult_79_FS_1_n240, u5_mult_79_FS_1_n239,
         u5_mult_79_FS_1_n238, u5_mult_79_FS_1_n237, u5_mult_79_FS_1_n236,
         u5_mult_79_FS_1_n235, u5_mult_79_FS_1_n234, u5_mult_79_FS_1_n233,
         u5_mult_79_FS_1_n232, u5_mult_79_FS_1_n231, u5_mult_79_FS_1_n230,
         u5_mult_79_FS_1_n229, u5_mult_79_FS_1_n228, u5_mult_79_FS_1_n227,
         u5_mult_79_FS_1_n226, u5_mult_79_FS_1_n225, u5_mult_79_FS_1_n224,
         u5_mult_79_FS_1_n223, u5_mult_79_FS_1_n222, u5_mult_79_FS_1_n221,
         u5_mult_79_FS_1_n220, u5_mult_79_FS_1_n219, u5_mult_79_FS_1_n218,
         u5_mult_79_FS_1_n217, u5_mult_79_FS_1_n216, u5_mult_79_FS_1_n215,
         u5_mult_79_FS_1_n214, u5_mult_79_FS_1_n213, u5_mult_79_FS_1_n212,
         u5_mult_79_FS_1_n211, u5_mult_79_FS_1_n210, u5_mult_79_FS_1_n209,
         u5_mult_79_FS_1_n208, u5_mult_79_FS_1_n207, u5_mult_79_FS_1_n206,
         u5_mult_79_FS_1_n205, u5_mult_79_FS_1_n204, u5_mult_79_FS_1_n203,
         u5_mult_79_FS_1_n202, u5_mult_79_FS_1_n201, u5_mult_79_FS_1_n200,
         u5_mult_79_FS_1_n199, u5_mult_79_FS_1_n198, u5_mult_79_FS_1_n197,
         u5_mult_79_FS_1_n196, u5_mult_79_FS_1_n195, u5_mult_79_FS_1_n194,
         u5_mult_79_FS_1_n193, u5_mult_79_FS_1_n192, u5_mult_79_FS_1_n191,
         u5_mult_79_FS_1_n190, u5_mult_79_FS_1_n189, u5_mult_79_FS_1_n188,
         u5_mult_79_FS_1_n187, u5_mult_79_FS_1_n186, u5_mult_79_FS_1_n185,
         u5_mult_79_FS_1_n184, u5_mult_79_FS_1_n183, u5_mult_79_FS_1_n182,
         u5_mult_79_FS_1_n181, u5_mult_79_FS_1_n180, u5_mult_79_FS_1_n179,
         u5_mult_79_FS_1_n178, u5_mult_79_FS_1_n177, u5_mult_79_FS_1_n176,
         u5_mult_79_FS_1_n175, u5_mult_79_FS_1_n174, u5_mult_79_FS_1_n173,
         u5_mult_79_FS_1_n172, u5_mult_79_FS_1_n171, u5_mult_79_FS_1_n170,
         u5_mult_79_FS_1_n169, u5_mult_79_FS_1_n168, u5_mult_79_FS_1_n167,
         u5_mult_79_FS_1_n166, u5_mult_79_FS_1_n165, u5_mult_79_FS_1_n164,
         u5_mult_79_FS_1_n163, u5_mult_79_FS_1_n162, u5_mult_79_FS_1_n161,
         u5_mult_79_FS_1_n160, u5_mult_79_FS_1_n159, u5_mult_79_FS_1_n158,
         u5_mult_79_FS_1_n157, u5_mult_79_FS_1_n156, u5_mult_79_FS_1_n155,
         u5_mult_79_FS_1_n154, u5_mult_79_FS_1_n153, u5_mult_79_FS_1_n152,
         u5_mult_79_FS_1_n151, u5_mult_79_FS_1_n150, u5_mult_79_FS_1_n149,
         u5_mult_79_FS_1_n148, u5_mult_79_FS_1_n147, u5_mult_79_FS_1_n146,
         u5_mult_79_FS_1_n145, u5_mult_79_FS_1_n144, u5_mult_79_FS_1_n143,
         u5_mult_79_FS_1_n142, u5_mult_79_FS_1_n141, u5_mult_79_FS_1_n140,
         u5_mult_79_FS_1_n139, u5_mult_79_FS_1_n138, u5_mult_79_FS_1_n137,
         u5_mult_79_FS_1_n136, u5_mult_79_FS_1_n135, u5_mult_79_FS_1_n134,
         u5_mult_79_FS_1_n133, u5_mult_79_FS_1_n132, u5_mult_79_FS_1_n131,
         u5_mult_79_FS_1_n130, u5_mult_79_FS_1_n129, u5_mult_79_FS_1_n128,
         u5_mult_79_FS_1_n127, u5_mult_79_FS_1_n126, u5_mult_79_FS_1_n125,
         u5_mult_79_FS_1_n124, u5_mult_79_FS_1_n123, u5_mult_79_FS_1_n122,
         u5_mult_79_FS_1_n121, u5_mult_79_FS_1_n120, u5_mult_79_FS_1_n119,
         u5_mult_79_FS_1_n118, u5_mult_79_FS_1_n117, u5_mult_79_FS_1_n116,
         u5_mult_79_FS_1_n115, u5_mult_79_FS_1_n114, u5_mult_79_FS_1_n113,
         u5_mult_79_FS_1_n112, u5_mult_79_FS_1_n111, u5_mult_79_FS_1_n110,
         u5_mult_79_FS_1_n109, u5_mult_79_FS_1_n108, u5_mult_79_FS_1_n107,
         u5_mult_79_FS_1_n106, u5_mult_79_FS_1_n105, u5_mult_79_FS_1_n104,
         u5_mult_79_FS_1_n103, u5_mult_79_FS_1_n102, u5_mult_79_FS_1_n101,
         u5_mult_79_FS_1_n100, u5_mult_79_FS_1_n99, u5_mult_79_FS_1_n98,
         u5_mult_79_FS_1_n97, u5_mult_79_FS_1_n96, u5_mult_79_FS_1_n95,
         u5_mult_79_FS_1_n94, u5_mult_79_FS_1_n93, u5_mult_79_FS_1_n92,
         u5_mult_79_FS_1_n91, u5_mult_79_FS_1_n90, u5_mult_79_FS_1_n89,
         u5_mult_79_FS_1_n88, u5_mult_79_FS_1_n87, u5_mult_79_FS_1_n86,
         u5_mult_79_FS_1_n85, u5_mult_79_FS_1_n84, u5_mult_79_FS_1_n83,
         u5_mult_79_FS_1_n82, u5_mult_79_FS_1_n81, u5_mult_79_FS_1_n80,
         u5_mult_79_FS_1_n79, u5_mult_79_FS_1_n78, u5_mult_79_FS_1_n77,
         u5_mult_79_FS_1_n76, u5_mult_79_FS_1_n75, u5_mult_79_FS_1_n74,
         u5_mult_79_FS_1_n73, u5_mult_79_FS_1_n72, u5_mult_79_FS_1_n71,
         u5_mult_79_FS_1_n70, u5_mult_79_FS_1_n69, u5_mult_79_FS_1_n68,
         u5_mult_79_FS_1_n67, u5_mult_79_FS_1_n66, u5_mult_79_FS_1_n65,
         u5_mult_79_FS_1_n64, u5_mult_79_FS_1_n63, u5_mult_79_FS_1_n62,
         u5_mult_79_FS_1_n61, u5_mult_79_FS_1_n60, u5_mult_79_FS_1_n59,
         u5_mult_79_FS_1_n58, u5_mult_79_FS_1_n57, u5_mult_79_FS_1_n56,
         u5_mult_79_FS_1_n55, u5_mult_79_FS_1_n54, u5_mult_79_FS_1_n53,
         u5_mult_79_FS_1_n52, u5_mult_79_FS_1_n51, u5_mult_79_FS_1_n50,
         u5_mult_79_FS_1_n49, u5_mult_79_FS_1_n48, u5_mult_79_FS_1_n47,
         u5_mult_79_FS_1_n46, u5_mult_79_FS_1_n45, u5_mult_79_FS_1_n44,
         u5_mult_79_FS_1_n43, u5_mult_79_FS_1_n42, u5_mult_79_FS_1_n41,
         u5_mult_79_FS_1_n40, u5_mult_79_FS_1_n39, u5_mult_79_FS_1_n38,
         u5_mult_79_FS_1_n37, u5_mult_79_FS_1_n36, u5_mult_79_FS_1_n35,
         u5_mult_79_FS_1_n34, u5_mult_79_FS_1_n33, u5_mult_79_FS_1_n32,
         u5_mult_79_FS_1_n31, u5_mult_79_FS_1_n30, u5_mult_79_FS_1_n29,
         u5_mult_79_FS_1_n28, u5_mult_79_FS_1_n27, u5_mult_79_FS_1_n26,
         u5_mult_79_FS_1_n25, u5_mult_79_FS_1_n24, u5_mult_79_FS_1_n23,
         u5_mult_79_FS_1_n22, u5_mult_79_FS_1_n21, u5_mult_79_FS_1_n20,
         u5_mult_79_FS_1_n19, u5_mult_79_FS_1_n18, u5_mult_79_FS_1_n17,
         u5_mult_79_FS_1_n16, u5_mult_79_FS_1_n15, u5_mult_79_FS_1_n14,
         u5_mult_79_FS_1_n13, u5_mult_79_FS_1_n12, u5_mult_79_FS_1_n11,
         u5_mult_79_FS_1_n10, u5_mult_79_FS_1_n9, u5_mult_79_FS_1_n8,
         u5_mult_79_FS_1_n7, u5_mult_79_FS_1_n6, u5_mult_79_FS_1_n5,
         u5_mult_79_FS_1_n4, u5_mult_79_FS_1_n3, u5_mult_79_FS_1_n2,
         u5_mult_79_FS_1_n1, u4_add_395_n68, u4_add_395_n67, u4_add_395_n66,
         u4_add_395_n65, u4_add_395_n64, u4_add_395_n63, u4_add_395_n62,
         u4_add_395_n61, u4_add_395_n60, u4_add_395_n59, u4_add_395_n58,
         u4_add_395_n57, u4_add_395_n56, u4_add_395_n55, u4_add_395_n54,
         u4_add_395_n53, u4_add_395_n52, u4_add_395_n51, u4_add_395_n50,
         u4_add_395_n49, u4_add_395_n48, u4_add_395_n47, u4_add_395_n46,
         u4_add_395_n45, u4_add_395_n44, u4_add_395_n43, u4_add_395_n42,
         u4_add_395_n41, u4_add_395_n40, u4_add_395_n39, u4_add_395_n38,
         u4_add_395_n37, u4_add_395_n36, u4_add_395_n35, u4_add_395_n34,
         u4_add_395_n33, u4_add_395_n32, u4_add_395_n31, u4_add_395_n30,
         u4_add_395_n29, u4_add_395_n28, u4_add_395_n27, u4_add_395_n26,
         u4_add_395_n25, u4_add_395_n24, u4_add_395_n23, u4_add_395_n22,
         u4_add_395_n21, u4_add_395_n20, u4_add_395_n19, u4_add_395_n18,
         u4_add_395_n17, u4_add_395_n16, u4_add_395_n15, u4_add_395_n14,
         u4_add_395_n13, u4_add_395_n12, u4_add_395_n11, u4_add_395_n10,
         u4_add_395_n9, u4_add_395_n8, u4_add_395_n7, u4_add_395_n5,
         u4_add_395_n3, u4_add_395_n2, u4_add_395_n1, u4_sub_495_n35,
         u4_sub_495_n34, u4_sub_495_n33, u4_sub_495_n32, u4_sub_495_n31,
         u4_sub_495_n30, u4_sub_495_n29, u4_sub_495_n28, u4_sub_495_n27,
         u4_sub_495_n26, u4_sub_495_n25, u4_sub_495_n24, u4_sub_495_n23,
         u4_sub_495_n22, u4_sub_495_n21, u4_sub_495_n20, u4_sub_495_n19,
         u4_sub_495_n18, u4_sub_495_n17, u4_sub_495_n16, u4_sub_495_n15,
         u4_sub_495_n14, u4_sub_495_n13, u4_sub_495_n12, u4_sub_495_n11,
         u4_sub_495_n10, u4_sub_495_n9, u4_sub_495_n8, u4_sub_495_n7,
         u4_sub_495_n6, u4_sub_495_n5, u4_sub_495_n4, u4_sub_495_n3,
         u4_sub_495_n2, u4_sub_495_n1, u4_sub_495_net32049,
         u4_sub_495_net32012, u4_sub_495_net32015, u4_sub_495_net32016,
         u4_sub_495_net32019, u4_sub_495_net32021, u4_sub_495_net32024,
         u4_sub_495_net32030, u4_sub_495_net32039, u4_sub_495_net32040,
         u4_sub_495_net32048, u4_sub_495_net32031, u4_sub_495_net32036,
         u4_sub_495_net32042, u4_sub_495_net32043, u4_sub_495_net32046,
         u4_sub_495_net32047, u4_sub_495_net32052, u4_sub_495_net32025,
         u4_sub_495_net32027, u4_sub_495_net32013, u4_sub_495_net95073,
         u4_sub_495_net94054, u4_sub_495_net91261, u4_sub_495_net32017,
         u4_sub_495_net32018, u4_sub_495_net32028, u4_sub_495_net32029,
         u4_sub_495_net32035, u4_sub_495_net32044, u4_sub_495_net32045,
         u4_sub_495_net32050, u4_sub_495_net32051, u4_sub_495_net32054,
         u4_sub_495_net32055, u4_add_463_n14, u4_add_463_n13, u4_add_463_n12,
         u4_add_463_n11, u4_add_463_n10, u4_add_463_n9, u4_add_463_n8,
         u4_add_463_n7, u4_add_463_n6, u4_add_463_n5, u4_add_463_n4,
         u4_add_463_n3, u4_add_463_n1, u4_add_493_n72, u4_add_493_n71,
         u4_add_493_n70, u4_add_493_n69, u4_add_493_n68, u4_add_493_n67,
         u4_add_493_n66, u4_add_493_n65, u4_add_493_n64, u4_add_493_n63,
         u4_add_493_n62, u4_add_493_n61, u4_add_493_n60, u4_add_493_n59,
         u4_add_493_n58, u4_add_493_n57, u4_add_493_n56, u4_add_493_n55,
         u4_add_493_n54, u4_add_493_n53, u4_add_493_n52, u4_add_493_n51,
         u4_add_493_n50, u4_add_493_n49, u4_add_493_n48, u4_add_493_n47,
         u4_add_493_n46, u4_add_493_n45, u4_add_493_n44, u4_add_493_n43,
         u4_add_493_n42, u4_add_493_n41, u4_add_493_n40, u4_add_493_n39,
         u4_add_493_n38, u4_add_493_n37, u4_add_493_n36, u4_add_493_n35,
         u4_add_493_n34, u4_add_493_n33, u4_add_493_n32, u4_add_493_n31,
         u4_add_493_n30, u4_add_493_n29, u4_add_493_n28, u4_add_493_n27,
         u4_add_493_n26, u4_add_493_n25, u4_add_493_n24, u4_add_493_n23,
         u4_add_493_n22, u4_add_493_n21, u4_add_493_n20, u4_add_493_n19,
         u4_add_493_n18, u4_add_493_n17, u4_add_493_n16, u4_add_493_n15,
         u4_add_493_n14, u4_add_493_n13, u4_add_493_n12, u4_add_493_n11,
         u4_add_493_n10, u4_add_493_n9, u4_add_493_n8, u4_add_493_n7,
         u4_add_493_n6, u4_add_493_n5, u4_add_493_n4, u4_add_493_n3,
         u4_add_493_n2, u4_add_493_n1, add_0_root_sub_0_root_u4_add_496_n66,
         add_0_root_sub_0_root_u4_add_496_n65,
         add_0_root_sub_0_root_u4_add_496_n64,
         add_0_root_sub_0_root_u4_add_496_n63,
         add_0_root_sub_0_root_u4_add_496_n62,
         add_0_root_sub_0_root_u4_add_496_n61,
         add_0_root_sub_0_root_u4_add_496_n60,
         add_0_root_sub_0_root_u4_add_496_n59,
         add_0_root_sub_0_root_u4_add_496_n58,
         add_0_root_sub_0_root_u4_add_496_n57,
         add_0_root_sub_0_root_u4_add_496_n56,
         add_0_root_sub_0_root_u4_add_496_n55,
         add_0_root_sub_0_root_u4_add_496_n54,
         add_0_root_sub_0_root_u4_add_496_n53,
         add_0_root_sub_0_root_u4_add_496_n52,
         add_0_root_sub_0_root_u4_add_496_n51,
         add_0_root_sub_0_root_u4_add_496_n50,
         add_0_root_sub_0_root_u4_add_496_n49,
         add_0_root_sub_0_root_u4_add_496_n48,
         add_0_root_sub_0_root_u4_add_496_n47,
         add_0_root_sub_0_root_u4_add_496_n46,
         add_0_root_sub_0_root_u4_add_496_n45,
         add_0_root_sub_0_root_u4_add_496_n44,
         add_0_root_sub_0_root_u4_add_496_n43,
         add_0_root_sub_0_root_u4_add_496_n42,
         add_0_root_sub_0_root_u4_add_496_n41,
         add_0_root_sub_0_root_u4_add_496_n40,
         add_0_root_sub_0_root_u4_add_496_n39,
         add_0_root_sub_0_root_u4_add_496_n38,
         add_0_root_sub_0_root_u4_add_496_n37,
         add_0_root_sub_0_root_u4_add_496_n36,
         add_0_root_sub_0_root_u4_add_496_n35,
         add_0_root_sub_0_root_u4_add_496_n34,
         add_0_root_sub_0_root_u4_add_496_n33,
         add_0_root_sub_0_root_u4_add_496_n32,
         add_0_root_sub_0_root_u4_add_496_n31,
         add_0_root_sub_0_root_u4_add_496_n30,
         add_0_root_sub_0_root_u4_add_496_n29,
         add_0_root_sub_0_root_u4_add_496_n28,
         add_0_root_sub_0_root_u4_add_496_n27,
         add_0_root_sub_0_root_u4_add_496_n26,
         add_0_root_sub_0_root_u4_add_496_n25,
         add_0_root_sub_0_root_u4_add_496_n24,
         add_0_root_sub_0_root_u4_add_496_n23,
         add_0_root_sub_0_root_u4_add_496_n22,
         add_0_root_sub_0_root_u4_add_496_n21,
         add_0_root_sub_0_root_u4_add_496_n20,
         add_0_root_sub_0_root_u4_add_496_n19,
         add_0_root_sub_0_root_u4_add_496_n18,
         add_0_root_sub_0_root_u4_add_496_n17,
         add_0_root_sub_0_root_u4_add_496_n16,
         add_0_root_sub_0_root_u4_add_496_n15,
         add_0_root_sub_0_root_u4_add_496_n14,
         add_0_root_sub_0_root_u4_add_496_n13,
         add_0_root_sub_0_root_u4_add_496_n12,
         add_0_root_sub_0_root_u4_add_496_n11,
         add_0_root_sub_0_root_u4_add_496_n10,
         add_0_root_sub_0_root_u4_add_496_n9,
         add_0_root_sub_0_root_u4_add_496_n8,
         add_0_root_sub_0_root_u4_add_496_n7,
         add_0_root_sub_0_root_u4_add_496_n6,
         add_0_root_sub_0_root_u4_add_496_n5,
         add_0_root_sub_0_root_u4_add_496_n4,
         add_0_root_sub_0_root_u4_add_496_n3,
         add_0_root_sub_0_root_u4_add_496_n2,
         add_0_root_sub_0_root_u4_add_496_n1, u4_add_465_n12, u4_add_465_n11,
         u4_add_465_n10, u4_add_465_n9, u4_add_465_n8, u4_add_465_n7,
         u4_add_465_n6, u4_add_465_n5, u4_add_465_n4, u4_add_465_n3,
         u4_add_465_n2, u4_add_465_n1, sub_1_root_u1_sub_130_aco_n99,
         sub_1_root_u1_sub_130_aco_n98, sub_1_root_u1_sub_130_aco_n97,
         sub_1_root_u1_sub_130_aco_n96, sub_1_root_u1_sub_130_aco_n95,
         sub_1_root_u1_sub_130_aco_n94, sub_1_root_u1_sub_130_aco_n93,
         sub_1_root_u1_sub_130_aco_n92, sub_1_root_u1_sub_130_aco_n91,
         sub_1_root_u1_sub_130_aco_n90, sub_1_root_u1_sub_130_aco_n89,
         sub_1_root_u1_sub_130_aco_n88, sub_1_root_u1_sub_130_aco_n87,
         sub_1_root_u1_sub_130_aco_n86, sub_1_root_u1_sub_130_aco_n85,
         sub_1_root_u1_sub_130_aco_n84, sub_1_root_u1_sub_130_aco_n83,
         sub_1_root_u1_sub_130_aco_n82, sub_1_root_u1_sub_130_aco_n81,
         sub_1_root_u1_sub_130_aco_n80, sub_1_root_u1_sub_130_aco_n79,
         sub_1_root_u1_sub_130_aco_n78, sub_1_root_u1_sub_130_aco_n77,
         sub_1_root_u1_sub_130_aco_n76, sub_1_root_u1_sub_130_aco_n75,
         sub_1_root_u1_sub_130_aco_n74, sub_1_root_u1_sub_130_aco_n73,
         sub_1_root_u1_sub_130_aco_n72, sub_1_root_u1_sub_130_aco_n71,
         sub_1_root_u1_sub_130_aco_n70, sub_1_root_u1_sub_130_aco_n69,
         sub_1_root_u1_sub_130_aco_n68, sub_1_root_u1_sub_130_aco_n67,
         sub_1_root_u1_sub_130_aco_n66, sub_1_root_u1_sub_130_aco_n65,
         sub_1_root_u1_sub_130_aco_n64, sub_1_root_u1_sub_130_aco_n63,
         sub_1_root_u1_sub_130_aco_n62, sub_1_root_u1_sub_130_aco_n61,
         sub_1_root_u1_sub_130_aco_n60, sub_1_root_u1_sub_130_aco_n59,
         sub_1_root_u1_sub_130_aco_n58, sub_1_root_u1_sub_130_aco_n57,
         sub_1_root_u1_sub_130_aco_n56, sub_1_root_u1_sub_130_aco_n55,
         sub_1_root_u1_sub_130_aco_n54, sub_1_root_u1_sub_130_aco_n53,
         sub_1_root_u1_sub_130_aco_n52, sub_1_root_u1_sub_130_aco_n51,
         sub_1_root_u1_sub_130_aco_n50, sub_1_root_u1_sub_130_aco_n49,
         sub_1_root_u1_sub_130_aco_n48, sub_1_root_u1_sub_130_aco_n47,
         sub_1_root_u1_sub_130_aco_n46, sub_1_root_u1_sub_130_aco_n45,
         sub_1_root_u1_sub_130_aco_n44, sub_1_root_u1_sub_130_aco_n43,
         sub_1_root_u1_sub_130_aco_n42, sub_1_root_u1_sub_130_aco_n41,
         sub_1_root_u1_sub_130_aco_n40, sub_1_root_u1_sub_130_aco_n39,
         sub_1_root_u1_sub_130_aco_n38, sub_1_root_u1_sub_130_aco_n37,
         sub_1_root_u1_sub_130_aco_n36, sub_1_root_u1_sub_130_aco_n35,
         sub_1_root_u1_sub_130_aco_n34, sub_1_root_u1_sub_130_aco_n33,
         sub_1_root_u1_sub_130_aco_n32, sub_1_root_u1_sub_130_aco_n31,
         sub_1_root_u1_sub_130_aco_n30, sub_1_root_u1_sub_130_aco_n29,
         sub_1_root_u1_sub_130_aco_n28, sub_1_root_u1_sub_130_aco_n27,
         sub_1_root_u1_sub_130_aco_n26, sub_1_root_u1_sub_130_aco_n25,
         sub_1_root_u1_sub_130_aco_n24, sub_1_root_u1_sub_130_aco_n23,
         sub_1_root_u1_sub_130_aco_n22, sub_1_root_u1_sub_130_aco_n21,
         sub_1_root_u1_sub_130_aco_n20, sub_1_root_u1_sub_130_aco_n19,
         sub_1_root_u1_sub_130_aco_n18, sub_1_root_u1_sub_130_aco_n17,
         sub_1_root_u1_sub_130_aco_n16, sub_1_root_u1_sub_130_aco_n15,
         sub_1_root_u1_sub_130_aco_n14, sub_1_root_u1_sub_130_aco_n13,
         sub_1_root_u1_sub_130_aco_n12, sub_1_root_u1_sub_130_aco_n11,
         sub_1_root_u1_sub_130_aco_n10, sub_1_root_u1_sub_130_aco_n9,
         sub_1_root_u1_sub_130_aco_n8, sub_1_root_u1_sub_130_aco_n7,
         sub_1_root_u1_sub_130_aco_n6, sub_1_root_u1_sub_130_aco_n5,
         sub_1_root_u1_sub_130_aco_n4, sub_1_root_u1_sub_130_aco_n3,
         sub_1_root_u1_sub_130_aco_n2, sub_1_root_u1_sub_130_aco_n1,
         u4_sub_469_n62, u4_sub_469_n61, u4_sub_469_n60, u4_sub_469_n59,
         u4_sub_469_n58, u4_sub_469_n57, u4_sub_469_n56, u4_sub_469_n55,
         u4_sub_469_n54, u4_sub_469_n53, u4_sub_469_n52, u4_sub_469_n51,
         u4_sub_469_n50, u4_sub_469_n49, u4_sub_469_n48, u4_sub_469_n47,
         u4_sub_469_n46, u4_sub_469_n45, u4_sub_469_n44, u4_sub_469_n43,
         u4_sub_469_n42, u4_sub_469_n41, u4_sub_469_n40, u4_sub_469_n39,
         u4_sub_469_n38, u4_sub_469_n37, u4_sub_469_n36, u4_sub_469_n35,
         u4_sub_469_n34, u4_sub_469_n33, u4_sub_469_n32, u4_sub_469_n31,
         u4_sub_469_n30, u4_sub_469_n29, u4_sub_469_n28, u4_sub_469_n27,
         u4_sub_469_n26, u4_sub_469_n25, u4_sub_469_n24, u4_sub_469_n23,
         u4_sub_469_n22, u4_sub_469_n21, u4_sub_469_n20, u4_sub_469_n19,
         u4_sub_469_n18, u4_sub_469_n17, u4_sub_469_n16, u4_sub_469_n15,
         u4_sub_469_n14, u4_sub_469_n13, u4_sub_469_n12, u4_sub_469_n11,
         u4_sub_469_n10, u4_sub_469_n9, u4_sub_469_n8, u4_sub_469_n7,
         u4_sub_469_n6, u4_sub_469_n5, u4_sub_469_n4, u4_sub_469_n2,
         u4_sub_469_n1;
  wire   [31:23] opa_r;
  wire   [31:23] opb_r;
  wire   [1:0] rmode_r1;
  wire   [1:0] rmode_r2;
  wire   [1:0] rmode_r3;
  wire   [2:0] fpu_op_r1;
  wire   [2:0] fpu_op_r2;
  wire   [26:0] fracta;
  wire   [26:0] fractb;
  wire   [7:0] exp_fasu;
  wire   [22:0] fracta_mul;
  wire   [7:0] exp_mul;
  wire   [1:0] exp_ovf;
  wire   [2:0] underflow_fmul_d;
  wire   [27:0] fract_out_q;
  wire   [47:0] prod;
  wire   [49:0] quo;
  wire   [49:0] remainder;
  wire   [4:0] div_opa_ldz_r1;
  wire   [4:0] div_opa_ldz_r2;
  wire   [6:3] exp_r;
  wire   [30:1] opa_r1;
  wire   [47:0] fract_i2f;
  wire   [45:21] fract_denorm;
  wire   [1:0] underflow_fmul_r;
  wire   [26:0] u1_fractb_s;
  wire   [26:0] u1_fracta_s;
  wire   [7:0] u1_exp_diff2;
  wire   [7:0] u1_exp_small;
  wire   [2:1] u2_underflow_d;
  wire   [47:0] u5_prod1;
  wire   [49:0] u6_remainder;
  wire   [49:0] u6_quo1;
  wire   [7:0] u4_div_exp3;
  wire   [56:49] u4_exp_f2i_1;
  wire   [7:0] u4_exp_fix_divb;
  wire   [7:0] u4_exp_fix_diva;
  wire   [6:2] u4_fi_ldz_mi22;
  wire   [5:0] u4_shift_left;
  wire   [7:0] u4_shift_right;
  wire   [7:0] u4_div_shft4;
  wire   [7:1] u4_sub_471_carry;
  wire   [27:1] u3_sub_60_carry;
  wire   [26:1] u3_add_60_carry;
  wire   [7:2] u2_add_117_carry;
  wire   [7:2] u2_add_115_carry;
  wire   [7:1] u2_add_112_carry;
  wire   [8:1] u2_sub_112_carry;
  wire   [44:25] u5_mult_79_CLA_SUM;
  wire   [45:24] u5_mult_79_CLA_CARRY;

  NOR2_X4 U16 ( .A1(net85393), .A2(n4759), .ZN(n1371) );
  NOR2_X4 U34 ( .A1(n4759), .A2(net23180), .ZN(n1373) );
  AND2_X2 U258 ( .A1(opb_r[31]), .A2(opa_r[31]), .ZN(u2_N97) );
  AOI221_X2 U500 ( .B1(opb_nan), .B2(n1725), .C1(n1726), .C2(
        u1_fracta_lt_fractb), .A(u1_signa_r), .ZN(n1722) );
  NAND2_X2 U502 ( .A1(opa_nan), .A2(opb_nan), .ZN(n1725) );
  OAI22_X2 U503 ( .A1(n2750), .A2(n1727), .B1(n1728), .B2(n1729), .ZN(u1_N129)
         );
  XNOR2_X2 U504 ( .A(n2748), .B(u1_add_r), .ZN(n1729) );
  AND2_X2 U505 ( .A1(n1727), .A2(n2750), .ZN(n1728) );
  AOI22_X2 U506 ( .A1(u0_snan_r_a), .A2(u0_expa_ff), .B1(u0_snan_r_b), .B2(
        u0_expb_ff), .ZN(n1730) );
  AOI22_X2 U507 ( .A1(u0_qnan_r_a), .A2(u0_expa_ff), .B1(u0_qnan_r_b), .B2(
        u0_expb_ff), .ZN(n1731) );
  NAND2_X2 U508 ( .A1(n1732), .A2(n1733), .ZN(u0_N7) );
  AND2_X2 U512 ( .A1(u0_fractb_00), .A2(u0_expb_00), .ZN(u0_N17) );
  AND2_X2 U513 ( .A1(u0_fracta_00), .A2(u0_expa_00), .ZN(u0_N16) );
  NAND2_X2 U514 ( .A1(u0_infb_f_r), .A2(u0_expb_ff), .ZN(n1732) );
  NAND2_X2 U515 ( .A1(u0_infa_f_r), .A2(u0_expa_ff), .ZN(n1733) );
  AND4_X2 U526 ( .A1(n1742), .A2(n1743), .A3(n1744), .A4(n1745), .ZN(n1735) );
  NOR4_X2 U527 ( .A1(fracta_mul[8]), .A2(fracta_mul[6]), .A3(fracta_mul[5]), 
        .A4(fracta_mul[4]), .ZN(n1745) );
  NOR4_X2 U529 ( .A1(fracta_mul[18]), .A2(fracta_mul[16]), .A3(fracta_mul[14]), 
        .A4(fracta_mul[12]), .ZN(n1743) );
  NOR4_X2 U538 ( .A1(n1754), .A2(n3049), .A3(u6_N3), .A4(u6_N2), .ZN(n1751) );
  OR2_X2 U543 ( .A1(u6_N0), .A2(u6_N10), .ZN(n1756) );
  NAND4_X2 U603 ( .A1(exp_mul[7]), .A2(exp_mul[6]), .A3(exp_mul[5]), .A4(
        exp_mul[4]), .ZN(n1822) );
  NAND4_X2 U604 ( .A1(exp_mul[3]), .A2(exp_mul[2]), .A3(exp_mul[1]), .A4(
        exp_mul[0]), .ZN(n1821) );
  AND4_X2 U605 ( .A1(opb_00), .A2(opa_nan_r), .A3(n2753), .A4(n2594), .ZN(N533) );
  NOR4_X2 U633 ( .A1(n1893), .A2(prod[26]), .A3(prod[28]), .A4(prod[27]), .ZN(
        n1892) );
  OR3_X2 U634 ( .A1(prod[2]), .A2(prod[30]), .A3(prod[29]), .ZN(n1893) );
  NOR4_X2 U637 ( .A1(n1895), .A2(prod[15]), .A3(prod[17]), .A4(prod[16]), .ZN(
        n1890) );
  OR3_X2 U638 ( .A1(prod[19]), .A2(prod[1]), .A3(prod[18]), .ZN(n1895) );
  NOR4_X2 U639 ( .A1(n1896), .A2(prod[0]), .A3(prod[11]), .A4(prod[10]), .ZN(
        n1889) );
  OR3_X2 U640 ( .A1(prod[13]), .A2(prod[14]), .A3(prod[12]), .ZN(n1896) );
  NOR4_X2 U642 ( .A1(n1901), .A2(prod[4]), .A3(prod[6]), .A4(prod[5]), .ZN(
        n1900) );
  OR3_X2 U643 ( .A1(prod[8]), .A2(prod[9]), .A3(prod[7]), .ZN(n1901) );
  NOR4_X2 U646 ( .A1(n1903), .A2(prod[37]), .A3(prod[39]), .A4(prod[38]), .ZN(
        n1898) );
  OR3_X2 U647 ( .A1(prod[40]), .A2(prod[41]), .A3(prod[3]), .ZN(n1903) );
  OR3_X2 U771 ( .A1(fracta_mul[13]), .A2(fracta_mul[15]), .A3(fracta_mul[14]), 
        .ZN(n2051) );
  AOI22_X2 U1017 ( .A1(u4_N1389), .A2(net85377), .B1(u4_N1439), .B2(n2794), 
        .ZN(n2083) );
  NOR3_X4 U1074 ( .A1(u4_N1361), .A2(u4_N1363), .A3(u4_N1362), .ZN(n2261) );
  XNOR2_X2 U1329 ( .A(n1727), .B(n5322), .ZN(N441) );
  NAND2_X2 U1330 ( .A1(rmode_r2[1]), .A2(rmode_r2[0]), .ZN(n1727) );
  OAI221_X2 U1395 ( .B1(n5321), .B2(n2616), .C1(n2759), .C2(n1823), .A(n2425), 
        .ZN(N221) );
  NAND2_X2 U1396 ( .A1(exp_fasu[7]), .A2(n2426), .ZN(n2425) );
  OAI221_X2 U1397 ( .B1(n5321), .B2(n2617), .C1(n2761), .C2(n1823), .A(n2427), 
        .ZN(N220) );
  NAND2_X2 U1398 ( .A1(exp_fasu[6]), .A2(n2426), .ZN(n2427) );
  OAI221_X2 U1399 ( .B1(n5321), .B2(n2612), .C1(n2757), .C2(n1823), .A(n2428), 
        .ZN(N219) );
  NAND2_X2 U1400 ( .A1(exp_fasu[5]), .A2(n2426), .ZN(n2428) );
  OAI221_X2 U1401 ( .B1(n5321), .B2(n2615), .C1(n2755), .C2(n1823), .A(n2429), 
        .ZN(N218) );
  NAND2_X2 U1402 ( .A1(exp_fasu[4]), .A2(n2426), .ZN(n2429) );
  OAI221_X2 U1403 ( .B1(n5321), .B2(n2611), .C1(n2758), .C2(n1823), .A(n2430), 
        .ZN(N217) );
  NAND2_X2 U1404 ( .A1(exp_fasu[3]), .A2(n2426), .ZN(n2430) );
  OR2_X2 U1405 ( .A1(n2567), .A2(fpu_op_r2[2]), .ZN(n1823) );
  OAI221_X2 U1407 ( .B1(n2431), .B2(n2614), .C1(n2760), .C2(n2567), .A(n2432), 
        .ZN(N216) );
  NAND2_X2 U1408 ( .A1(exp_fasu[2]), .A2(n2426), .ZN(n2432) );
  OAI221_X2 U1409 ( .B1(n2431), .B2(n2610), .C1(n2756), .C2(n2567), .A(n2433), 
        .ZN(N215) );
  NAND2_X2 U1410 ( .A1(exp_fasu[1]), .A2(n2426), .ZN(n2433) );
  OAI221_X2 U1411 ( .B1(n2431), .B2(n2613), .C1(n2754), .C2(n2567), .A(n2434), 
        .ZN(N214) );
  NAND2_X2 U1412 ( .A1(exp_fasu[0]), .A2(n2426), .ZN(n2434) );
  NOR4_X2 U1425 ( .A1(fracta_mul[15]), .A2(fracta_mul[17]), .A3(fracta_mul[19]), .A4(fracta_mul[21]), .ZN(n2437) );
  OAI211_X2 U1429 ( .C1(n2449), .C2(n2450), .A(n2687), .B(n2696), .ZN(n2448)
         );
  OR3_X2 U1431 ( .A1(fracta_mul[6]), .A2(fracta_mul[7]), .A3(fracta_mul[11]), 
        .ZN(n2452) );
  OR2_X2 U1432 ( .A1(fracta_mul[12]), .A2(fracta_mul[13]), .ZN(n2449) );
  OAI33_X1 U1932 ( .A1(n2451), .A2(fracta_mul[11]), .A3(fracta_mul[10]), .B1(
        n2452), .B2(fracta_mul[10]), .B3(n2453), .ZN(n2450) );
  DFF_X2 opa_r_reg_31_ ( .D(opa[31]), .CK(clk), .Q(opa_r[31]) );
  DFF_X2 opa_r_reg_30_ ( .D(opa[30]), .CK(clk), .Q(opa_r[30]), .QN(n2566) );
  DFF_X2 opa_r_reg_29_ ( .D(opa[29]), .CK(clk), .Q(opa_r[29]), .QN(n2653) );
  DFF_X2 opa_r_reg_28_ ( .D(opa[28]), .CK(clk), .Q(opa_r[28]), .QN(n2582) );
  DFF_X2 opa_r_reg_27_ ( .D(opa[27]), .CK(clk), .Q(opa_r[27]), .QN(n2657) );
  DFF_X2 opa_r_reg_26_ ( .D(opa[26]), .CK(clk), .Q(opa_r[26]), .QN(n2764) );
  DFF_X2 opa_r_reg_25_ ( .D(opa[25]), .CK(clk), .Q(opa_r[25]), .QN(n2765) );
  DFF_X2 opa_r_reg_24_ ( .D(opa[24]), .CK(clk), .Q(opa_r[24]), .QN(n2763) );
  DFF_X2 opa_r_reg_23_ ( .D(opa[23]), .CK(clk), .Q(opa_r[23]), .QN(n2655) );
  DFF_X2 opa_r_reg_22_ ( .D(opa[22]), .CK(clk), .Q(fracta_mul[22]), .QN(n2591)
         );
  DFF_X2 opa_r_reg_21_ ( .D(opa[21]), .CK(clk), .Q(fracta_mul[21]), .QN(n2599)
         );
  DFF_X2 opa_r_reg_20_ ( .D(opa[20]), .CK(clk), .Q(fracta_mul[20]), .QN(n2683)
         );
  DFF_X2 opa_r_reg_19_ ( .D(opa[19]), .CK(clk), .Q(fracta_mul[19]), .QN(n2592)
         );
  DFF_X2 opa_r_reg_18_ ( .D(opa[18]), .CK(clk), .Q(fracta_mul[18]), .QN(n2677)
         );
  DFF_X2 opa_r_reg_17_ ( .D(opa[17]), .CK(clk), .Q(fracta_mul[17]), .QN(n2590)
         );
  DFF_X2 opa_r_reg_16_ ( .D(opa[16]), .CK(clk), .Q(fracta_mul[16]), .QN(n2675)
         );
  DFF_X2 opa_r_reg_15_ ( .D(opa[15]), .CK(clk), .Q(fracta_mul[15]), .QN(n2696)
         );
  DFF_X2 opa_r_reg_14_ ( .D(opa[14]), .CK(clk), .Q(fracta_mul[14]), .QN(n2687)
         );
  DFF_X2 opa_r_reg_13_ ( .D(opa[13]), .CK(clk), .Q(fracta_mul[13]), .QN(n2678)
         );
  DFF_X2 opa_r_reg_12_ ( .D(opa[12]), .CK(clk), .Q(fracta_mul[12]), .QN(n2692)
         );
  DFF_X2 opa_r_reg_11_ ( .D(opa[11]), .CK(clk), .Q(fracta_mul[11]), .QN(n2697)
         );
  DFF_X2 opa_r_reg_10_ ( .D(opa[10]), .CK(clk), .Q(fracta_mul[10]), .QN(n2593)
         );
  DFF_X2 opa_r_reg_9_ ( .D(opa[9]), .CK(clk), .Q(fracta_mul[9]), .QN(n2681) );
  DFF_X2 opa_r_reg_8_ ( .D(opa[8]), .CK(clk), .Q(fracta_mul[8]), .QN(n2695) );
  DFF_X2 opa_r_reg_7_ ( .D(opa[7]), .CK(clk), .Q(fracta_mul[7]), .QN(n2689) );
  DFF_X2 opa_r_reg_6_ ( .D(opa[6]), .CK(clk), .Q(fracta_mul[6]), .QN(n2685) );
  DFF_X2 opa_r_reg_5_ ( .D(opa[5]), .CK(clk), .Q(fracta_mul[5]), .QN(n2596) );
  DFF_X2 opa_r_reg_4_ ( .D(opa[4]), .CK(clk), .Q(fracta_mul[4]), .QN(n2690) );
  DFF_X2 opa_r_reg_3_ ( .D(opa[3]), .CK(clk), .Q(fracta_mul[3]), .QN(n2598) );
  DFF_X2 opa_r_reg_2_ ( .D(opa[2]), .CK(clk), .Q(fracta_mul[2]), .QN(n2999) );
  DFF_X2 opa_r_reg_1_ ( .D(opa[1]), .CK(clk), .Q(n2586), .QN(n3033) );
  DFF_X2 opa_r_reg_0_ ( .D(opa[0]), .CK(clk), .Q(fracta_mul[0]), .QN(n3053) );
  DFF_X2 opb_r_reg_31_ ( .D(opb[31]), .CK(clk), .Q(opb_r[31]) );
  DFF_X2 opb_r_reg_29_ ( .D(opb[29]), .CK(clk), .Q(opb_r[29]), .QN(n3060) );
  DFF_X2 opb_r_reg_28_ ( .D(opb[28]), .CK(clk), .Q(opb_r[28]), .QN(n3063) );
  DFF_X2 opb_r_reg_27_ ( .D(opb[27]), .CK(clk), .Q(opb_r[27]), .QN(n3064) );
  DFF_X2 opb_r_reg_26_ ( .D(opb[26]), .CK(clk), .Q(opb_r[26]), .QN(n3061) );
  DFF_X2 opb_r_reg_25_ ( .D(opb[25]), .CK(clk), .Q(opb_r[25]), .QN(n3062) );
  DFF_X2 opb_r_reg_24_ ( .D(opb[24]), .CK(clk), .Q(opb_r[24]), .QN(n3058) );
  DFF_X2 opb_r_reg_23_ ( .D(opb[23]), .CK(clk), .Q(opb_r[23]), .QN(n3059) );
  DFF_X2 opb_r_reg_18_ ( .D(opb[18]), .CK(clk), .Q(u6_N18), .QN(n3034) );
  DFF_X2 opb_r_reg_17_ ( .D(opb[17]), .CK(clk), .Q(u6_N17), .QN(n3031) );
  DFF_X2 opb_r_reg_15_ ( .D(opb[15]), .CK(clk), .Q(u6_N15), .QN(n2941) );
  DFF_X2 opb_r_reg_13_ ( .D(opb[13]), .CK(clk), .Q(u6_N13), .QN(n3004) );
  DFF_X2 opb_r_reg_10_ ( .D(opb[10]), .CK(clk), .Q(u6_N10), .QN(n2943) );
  DFF_X2 opb_r_reg_9_ ( .D(opb[9]), .CK(clk), .Q(u6_N9), .QN(n2922) );
  DFF_X2 opb_r_reg_8_ ( .D(opb[8]), .CK(clk), .Q(u6_N8), .QN(n2920) );
  DFF_X2 opb_r_reg_7_ ( .D(opb[7]), .CK(clk), .Q(u6_N7), .QN(n2768) );
  DFF_X2 opb_r_reg_6_ ( .D(opb[6]), .CK(clk), .Q(u6_N6), .QN(n2589) );
  DFF_X2 opb_r_reg_5_ ( .D(opb[5]), .CK(clk), .Q(u6_N5), .QN(n2706) );
  DFF_X2 opb_r_reg_4_ ( .D(opb[4]), .CK(clk), .Q(u6_N4), .QN(n2705) );
  DFF_X2 opb_r_reg_3_ ( .D(opb[3]), .CK(clk), .Q(u6_N3), .QN(n2703) );
  DFF_X2 opb_r_reg_2_ ( .D(opb[2]), .CK(clk), .Q(u6_N2), .QN(n2702) );
  DFF_X2 opb_r_reg_1_ ( .D(opb[1]), .CK(clk), .Q(u6_N1), .QN(n2701) );
  DFF_X2 opb_r_reg_0_ ( .D(opb[0]), .CK(clk), .Q(u6_N0), .QN(n2708) );
  DFF_X2 rmode_r1_reg_1_ ( .D(rmode[1]), .CK(clk), .Q(rmode_r1[1]) );
  DFF_X2 rmode_r1_reg_0_ ( .D(rmode[0]), .CK(clk), .Q(rmode_r1[0]) );
  DFF_X2 rmode_r2_reg_1_ ( .D(rmode_r1[1]), .CK(clk), .Q(rmode_r2[1]) );
  DFF_X2 rmode_r2_reg_0_ ( .D(rmode_r1[0]), .CK(clk), .Q(rmode_r2[0]) );
  DFF_X2 rmode_r3_reg_1_ ( .D(rmode_r2[1]), .CK(clk), .Q(rmode_r3[1]), .QN(
        n2578) );
  DFF_X2 rmode_r3_reg_0_ ( .D(rmode_r2[0]), .CK(clk), .Q(rmode_r3[0]), .QN(
        n2660) );
  DFF_X2 fpu_op_r1_reg_2_ ( .D(fpu_op[2]), .CK(clk), .Q(fpu_op_r1[2]), .QN(
        n2711) );
  DFF_X2 fpu_op_r1_reg_1_ ( .D(fpu_op[1]), .CK(clk), .Q(fpu_op_r1[1]) );
  DFF_X2 fpu_op_r1_reg_0_ ( .D(fpu_op[0]), .CK(clk), .Q(fpu_op_r1[0]), .QN(
        n2700) );
  DFF_X2 fpu_op_r2_reg_2_ ( .D(fpu_op_r1[2]), .CK(clk), .Q(fpu_op_r2[2]) );
  DFF_X2 fpu_op_r2_reg_1_ ( .D(fpu_op_r1[1]), .CK(clk), .Q(fpu_op_r2[1]), .QN(
        n2567) );
  DFF_X2 fpu_op_r2_reg_0_ ( .D(fpu_op_r1[0]), .CK(clk), .Q(fpu_op_r2[0]), .QN(
        n2752) );
  DFF_X2 fpu_op_r3_reg_2_ ( .D(fpu_op_r2[2]), .CK(clk), .Q(net90945), .QN(
        net86257) );
  DFF_X2 fpu_op_r3_reg_1_ ( .D(fpu_op_r2[1]), .CK(clk), .Q(fpu_op_r3_1_), .QN(
        net86236) );
  DFF_X2 div_opa_ldz_r1_reg_4_ ( .D(n2587), .CK(clk), .Q(div_opa_ldz_r1[4]) );
  DFF_X2 div_opa_ldz_r1_reg_3_ ( .D(n2597), .CK(clk), .Q(div_opa_ldz_r1[3]) );
  DFF_X2 div_opa_ldz_r1_reg_2_ ( .D(N107), .CK(clk), .Q(div_opa_ldz_r1[2]) );
  DFF_X2 div_opa_ldz_r1_reg_1_ ( .D(N141), .CK(clk), .Q(div_opa_ldz_r1[1]) );
  DFF_X2 div_opa_ldz_r1_reg_0_ ( .D(N170), .CK(clk), .Q(div_opa_ldz_r1[0]) );
  DFF_X2 div_opa_ldz_r2_reg_4_ ( .D(div_opa_ldz_r1[4]), .CK(clk), .Q(
        div_opa_ldz_r2[4]), .QN(n2688) );
  DFF_X2 div_opa_ldz_r2_reg_3_ ( .D(div_opa_ldz_r1[3]), .CK(clk), .Q(
        div_opa_ldz_r2[3]), .QN(n2694) );
  DFF_X2 div_opa_ldz_r2_reg_2_ ( .D(div_opa_ldz_r1[2]), .CK(clk), .Q(
        div_opa_ldz_r2[2]), .QN(n2691) );
  DFF_X2 div_opa_ldz_r2_reg_1_ ( .D(div_opa_ldz_r1[1]), .CK(clk), .Q(
        div_opa_ldz_r2[1]), .QN(n2654) );
  DFF_X2 div_opa_ldz_r2_reg_0_ ( .D(div_opa_ldz_r1[0]), .CK(clk), .Q(
        div_opa_ldz_r2[0]), .QN(n2581) );
  DFF_X2 opa_r1_reg_30_ ( .D(opa_r[30]), .CK(clk), .Q(opa_r1[30]), .QN(n2616)
         );
  DFF_X2 opa_r1_reg_29_ ( .D(opa_r[29]), .CK(clk), .Q(opa_r1[29]), .QN(n2617)
         );
  DFF_X2 opa_r1_reg_28_ ( .D(opa_r[28]), .CK(clk), .Q(opa_r1[28]), .QN(n2612)
         );
  DFF_X2 opa_r1_reg_27_ ( .D(opa_r[27]), .CK(clk), .Q(opa_r1[27]), .QN(n2615)
         );
  DFF_X2 opa_r1_reg_26_ ( .D(opa_r[26]), .CK(clk), .Q(opa_r1[26]), .QN(n2611)
         );
  DFF_X2 opa_r1_reg_25_ ( .D(opa_r[25]), .CK(clk), .Q(opa_r1[25]), .QN(n2614)
         );
  DFF_X2 opa_r1_reg_24_ ( .D(opa_r[24]), .CK(clk), .Q(opa_r1[24]), .QN(n2610)
         );
  DFF_X2 opa_r1_reg_23_ ( .D(opa_r[23]), .CK(clk), .Q(opa_r1[23]), .QN(n2613)
         );
  DFF_X2 opa_r1_reg_22_ ( .D(fracta_mul[22]), .CK(clk), .Q(opa_r1[22]) );
  DFF_X2 opa_r1_reg_21_ ( .D(fracta_mul[21]), .CK(clk), .Q(opa_r1[21]) );
  DFF_X2 opa_r1_reg_20_ ( .D(fracta_mul[20]), .CK(clk), .Q(opa_r1[20]) );
  DFF_X2 opa_r1_reg_19_ ( .D(fracta_mul[19]), .CK(clk), .Q(opa_r1[19]) );
  DFF_X2 opa_r1_reg_18_ ( .D(fracta_mul[18]), .CK(clk), .Q(opa_r1[18]) );
  DFF_X2 opa_r1_reg_17_ ( .D(fracta_mul[17]), .CK(clk), .Q(opa_r1[17]) );
  DFF_X2 opa_r1_reg_16_ ( .D(fracta_mul[16]), .CK(clk), .Q(opa_r1[16]) );
  DFF_X2 opa_r1_reg_15_ ( .D(fracta_mul[15]), .CK(clk), .Q(opa_r1[15]) );
  DFF_X2 opa_r1_reg_14_ ( .D(fracta_mul[14]), .CK(clk), .Q(opa_r1[14]) );
  DFF_X2 opa_r1_reg_13_ ( .D(fracta_mul[13]), .CK(clk), .Q(opa_r1[13]) );
  DFF_X2 opa_r1_reg_12_ ( .D(fracta_mul[12]), .CK(clk), .Q(opa_r1[12]) );
  DFF_X2 opa_r1_reg_11_ ( .D(fracta_mul[11]), .CK(clk), .Q(opa_r1[11]) );
  DFF_X2 opa_r1_reg_10_ ( .D(fracta_mul[10]), .CK(clk), .Q(opa_r1[10]) );
  DFF_X2 opa_r1_reg_9_ ( .D(fracta_mul[9]), .CK(clk), .Q(opa_r1[9]) );
  DFF_X2 opa_r1_reg_8_ ( .D(fracta_mul[8]), .CK(clk), .Q(opa_r1[8]) );
  DFF_X2 opa_r1_reg_7_ ( .D(fracta_mul[7]), .CK(clk), .Q(opa_r1[7]) );
  DFF_X2 opa_r1_reg_6_ ( .D(fracta_mul[6]), .CK(clk), .Q(opa_r1[6]) );
  DFF_X2 opa_r1_reg_5_ ( .D(fracta_mul[5]), .CK(clk), .Q(opa_r1[5]) );
  DFF_X2 opa_r1_reg_4_ ( .D(fracta_mul[4]), .CK(clk), .Q(opa_r1[4]) );
  DFF_X2 opa_r1_reg_3_ ( .D(fracta_mul[3]), .CK(clk), .Q(opa_r1[3]) );
  DFF_X2 opa_r1_reg_2_ ( .D(fracta_mul[2]), .CK(clk), .Q(opa_r1[2]) );
  DFF_X2 opa_r1_reg_1_ ( .D(n2586), .CK(clk), .Q(opa_r1[1]) );
  DFF_X2 opa_r1_reg_0_ ( .D(fracta_mul[0]), .CK(clk), .Q(N227), .QN(n2749) );
  DFF_X2 opas_r1_reg ( .D(opa_r[31]), .CK(clk), .Q(opas_r1) );
  DFF_X2 opas_r2_reg ( .D(opas_r1), .CK(clk), .Q(opas_r2), .QN(n2577) );
  DFF_X2 u0_fractb_00_reg ( .D(n4763), .CK(clk), .Q(u0_fractb_00) );
  DFF_X2 u0_fracta_00_reg ( .D(n4762), .CK(clk), .Q(u0_fracta_00) );
  DFF_X2 u0_expb_00_reg ( .D(n4765), .CK(clk), .Q(u0_expb_00) );
  DFF_X2 u0_opb_dn_reg ( .D(u0_expb_00), .CK(clk), .Q(net94019), .QN(net86235)
         );
  DFF_X2 u0_opb_00_reg ( .D(u0_N17), .CK(clk), .Q(opb_00), .QN(n2698) );
  DFF_X2 u0_expa_00_reg ( .D(n3093), .CK(clk), .Q(u0_expa_00) );
  DFF_X2 u0_opa_dn_reg ( .D(u0_expa_00), .CK(clk), .Q(opa_dn), .QN(n2584) );
  DFF_X2 u0_opa_00_reg ( .D(u0_N16), .CK(clk), .Q(opa_00), .QN(n2753) );
  DFF_X2 u0_opb_nan_reg ( .D(u0_N11), .CK(clk), .Q(opb_nan), .QN(n2751) );
  DFF_X2 u0_opa_nan_reg ( .D(u0_N10), .CK(clk), .Q(opa_nan) );
  DFF_X2 opa_nan_r_reg ( .D(N532), .CK(clk), .Q(opa_nan_r) );
  DFF_X2 u0_snan_r_b_reg ( .D(u0_N5), .CK(clk), .Q(u0_snan_r_b) );
  DFF_X2 u0_qnan_r_b_reg ( .D(u6_N22), .CK(clk), .Q(u0_qnan_r_b) );
  DFF_X2 u0_snan_r_a_reg ( .D(u0_N4), .CK(clk), .Q(u0_snan_r_a) );
  DFF_X2 u0_qnan_r_a_reg ( .D(fracta_mul[22]), .CK(clk), .Q(u0_qnan_r_a) );
  DFF_X2 u0_infb_f_r_reg ( .D(n4763), .CK(clk), .Q(u0_infb_f_r) );
  DFF_X2 u0_infa_f_r_reg ( .D(n4762), .CK(clk), .Q(u0_infa_f_r) );
  DFF_X2 u0_expb_ff_reg ( .D(n4760), .CK(clk), .Q(u0_expb_ff) );
  DFF_X2 u0_opb_inf_reg ( .D(n5329), .CK(clk), .Q(opb_inf), .QN(n2707) );
  DFF_X2 u0_expa_ff_reg ( .D(n4761), .CK(clk), .Q(u0_expa_ff) );
  DFF_X2 u0_snan_reg ( .D(n5327), .CK(clk), .Q(snan_d), .QN(n2607) );
  DFF_X2 snan_reg ( .D(snan_d), .CK(clk), .Q(snan) );
  DFF_X2 u0_qnan_reg ( .D(n5328), .CK(clk), .QN(n2736) );
  DFF_X2 u0_opa_inf_reg ( .D(n5330), .CK(clk), .Q(opa_inf), .QN(n2594) );
  DFF_X2 div_by_zero_reg ( .D(N533), .CK(clk), .Q(div_by_zero) );
  DFF_X2 u0_inf_reg ( .D(u0_N7), .CK(clk), .Q(inf_d), .QN(n2709) );
  DFF_X2 u0_ind_reg ( .D(u0_N6), .CK(clk), .Q(ind_d), .QN(n2731) );
  DFF_X2 u1_fasu_op_reg ( .D(n5287), .CK(clk), .Q(n2570), .QN(n2609) );
  DFF_X2 fasu_op_r1_reg ( .D(n3095), .CK(clk), .Q(fasu_op_r1) );
  DFF_X2 fasu_op_r2_reg ( .D(fasu_op_r1), .CK(clk), .QN(n2738) );
  DFF_X2 qnan_reg ( .D(N524), .CK(clk), .Q(qnan) );
  DFF_X2 u1_fracta_eq_fractb_reg ( .D(u1_N131), .CK(clk), .Q(
        u1_fracta_eq_fractb) );
  DFF_X2 u1_fracta_lt_fractb_reg ( .D(u1_N130), .CK(clk), .Q(
        u1_fracta_lt_fractb) );
  DFF_X2 u1_add_r_reg ( .D(n2700), .CK(clk), .Q(u1_add_r) );
  DFF_X2 u1_signb_r_reg ( .D(opb_r[31]), .CK(clk), .QN(n2748) );
  DFF_X2 u1_signa_r_reg ( .D(opa_r[31]), .CK(clk), .Q(u1_signa_r), .QN(n2750)
         );
  DFF_X2 u1_result_zero_sign_reg ( .D(u1_N129), .CK(clk), .Q(
        result_zero_sign_d) );
  DFF_X2 u1_nan_sign_reg ( .D(u1_N140), .CK(clk), .QN(n2728) );
  DFF_X2 sign_fasu_r_reg ( .D(sign_fasu), .CK(clk), .Q(sign_fasu_r) );
  DFF_X2 u1_fractb_out_reg_0_ ( .D(u1_fractb_s[0]), .CK(clk), .Q(fractb[0]) );
  DFF_X2 u1_fractb_out_reg_1_ ( .D(u1_fractb_s[1]), .CK(clk), .Q(fractb[1]) );
  DFF_X2 u1_fractb_out_reg_2_ ( .D(u1_fractb_s[2]), .CK(clk), .Q(fractb[2]) );
  DFF_X2 u1_fractb_out_reg_3_ ( .D(u1_fractb_s[3]), .CK(clk), .Q(fractb[3]) );
  DFF_X2 u1_fractb_out_reg_4_ ( .D(u1_fractb_s[4]), .CK(clk), .Q(fractb[4]) );
  DFF_X2 u1_fractb_out_reg_5_ ( .D(u1_fractb_s[5]), .CK(clk), .Q(fractb[5]) );
  DFF_X2 u1_fractb_out_reg_6_ ( .D(u1_fractb_s[6]), .CK(clk), .Q(fractb[6]) );
  DFF_X2 u1_fractb_out_reg_7_ ( .D(u1_fractb_s[7]), .CK(clk), .Q(fractb[7]) );
  DFF_X2 u1_fractb_out_reg_8_ ( .D(u1_fractb_s[8]), .CK(clk), .Q(fractb[8]) );
  DFF_X2 u1_fractb_out_reg_9_ ( .D(u1_fractb_s[9]), .CK(clk), .Q(fractb[9]) );
  DFF_X2 u1_fractb_out_reg_10_ ( .D(u1_fractb_s[10]), .CK(clk), .Q(fractb[10])
         );
  DFF_X2 u1_fractb_out_reg_11_ ( .D(u1_fractb_s[11]), .CK(clk), .Q(fractb[11])
         );
  DFF_X2 u1_fractb_out_reg_12_ ( .D(u1_fractb_s[12]), .CK(clk), .Q(fractb[12])
         );
  DFF_X2 u1_fractb_out_reg_13_ ( .D(u1_fractb_s[13]), .CK(clk), .Q(fractb[13])
         );
  DFF_X2 u1_fractb_out_reg_14_ ( .D(u1_fractb_s[14]), .CK(clk), .Q(fractb[14])
         );
  DFF_X2 u1_fractb_out_reg_15_ ( .D(u1_fractb_s[15]), .CK(clk), .Q(fractb[15])
         );
  DFF_X2 u1_fractb_out_reg_16_ ( .D(u1_fractb_s[16]), .CK(clk), .Q(fractb[16])
         );
  DFF_X2 u1_fractb_out_reg_17_ ( .D(u1_fractb_s[17]), .CK(clk), .Q(fractb[17])
         );
  DFF_X2 u1_fractb_out_reg_18_ ( .D(u1_fractb_s[18]), .CK(clk), .Q(fractb[18])
         );
  DFF_X2 u1_fractb_out_reg_19_ ( .D(u1_fractb_s[19]), .CK(clk), .Q(fractb[19])
         );
  DFF_X2 u1_fractb_out_reg_20_ ( .D(u1_fractb_s[20]), .CK(clk), .Q(fractb[20])
         );
  DFF_X2 u1_fractb_out_reg_21_ ( .D(u1_fractb_s[21]), .CK(clk), .Q(fractb[21])
         );
  DFF_X2 u1_fractb_out_reg_22_ ( .D(u1_fractb_s[22]), .CK(clk), .Q(fractb[22])
         );
  DFF_X2 u1_fractb_out_reg_23_ ( .D(u1_fractb_s[23]), .CK(clk), .Q(fractb[23])
         );
  DFF_X2 u1_fractb_out_reg_24_ ( .D(u1_fractb_s[24]), .CK(clk), .Q(fractb[24])
         );
  DFF_X2 u1_fractb_out_reg_25_ ( .D(u1_fractb_s[25]), .CK(clk), .Q(fractb[25])
         );
  DFF_X2 u1_fractb_out_reg_26_ ( .D(u1_fractb_s[26]), .CK(clk), .Q(fractb[26])
         );
  DFF_X2 u1_fracta_out_reg_0_ ( .D(u1_fracta_s[0]), .CK(clk), .Q(fracta[0]) );
  DFF_X2 u1_fracta_out_reg_1_ ( .D(u1_fracta_s[1]), .CK(clk), .Q(fracta[1]) );
  DFF_X2 u1_fracta_out_reg_2_ ( .D(u1_fracta_s[2]), .CK(clk), .Q(fracta[2]) );
  DFF_X2 u1_fracta_out_reg_3_ ( .D(u1_fracta_s[3]), .CK(clk), .Q(fracta[3]) );
  DFF_X2 u1_fracta_out_reg_4_ ( .D(u1_fracta_s[4]), .CK(clk), .Q(fracta[4]) );
  DFF_X2 u1_fracta_out_reg_5_ ( .D(u1_fracta_s[5]), .CK(clk), .Q(fracta[5]) );
  DFF_X2 u1_fracta_out_reg_6_ ( .D(u1_fracta_s[6]), .CK(clk), .Q(fracta[6]) );
  DFF_X2 u1_fracta_out_reg_7_ ( .D(u1_fracta_s[7]), .CK(clk), .Q(fracta[7]) );
  DFF_X2 u1_fracta_out_reg_8_ ( .D(u1_fracta_s[8]), .CK(clk), .Q(fracta[8]) );
  DFF_X2 u1_fracta_out_reg_9_ ( .D(u1_fracta_s[9]), .CK(clk), .Q(fracta[9]) );
  DFF_X2 u1_fracta_out_reg_10_ ( .D(u1_fracta_s[10]), .CK(clk), .Q(fracta[10])
         );
  DFF_X2 u1_fracta_out_reg_11_ ( .D(u1_fracta_s[11]), .CK(clk), .Q(fracta[11])
         );
  DFF_X2 u1_fracta_out_reg_12_ ( .D(u1_fracta_s[12]), .CK(clk), .Q(fracta[12])
         );
  DFF_X2 u1_fracta_out_reg_13_ ( .D(u1_fracta_s[13]), .CK(clk), .Q(fracta[13])
         );
  DFF_X2 u1_fracta_out_reg_14_ ( .D(u1_fracta_s[14]), .CK(clk), .Q(fracta[14])
         );
  DFF_X2 u1_fracta_out_reg_15_ ( .D(u1_fracta_s[15]), .CK(clk), .Q(fracta[15])
         );
  DFF_X2 u1_fracta_out_reg_16_ ( .D(u1_fracta_s[16]), .CK(clk), .Q(fracta[16])
         );
  DFF_X2 u1_fracta_out_reg_17_ ( .D(u1_fracta_s[17]), .CK(clk), .Q(fracta[17])
         );
  DFF_X2 u1_fracta_out_reg_18_ ( .D(u1_fracta_s[18]), .CK(clk), .Q(fracta[18])
         );
  DFF_X2 u1_fracta_out_reg_19_ ( .D(u1_fracta_s[19]), .CK(clk), .Q(fracta[19])
         );
  DFF_X2 u1_fracta_out_reg_20_ ( .D(u1_fracta_s[20]), .CK(clk), .Q(fracta[20])
         );
  DFF_X2 u1_fracta_out_reg_21_ ( .D(u1_fracta_s[21]), .CK(clk), .Q(fracta[21])
         );
  DFF_X2 u1_fracta_out_reg_22_ ( .D(u1_fracta_s[22]), .CK(clk), .Q(fracta[22])
         );
  DFF_X2 u1_fracta_out_reg_23_ ( .D(u1_fracta_s[23]), .CK(clk), .Q(fracta[23])
         );
  DFF_X2 u1_fracta_out_reg_24_ ( .D(u1_fracta_s[24]), .CK(clk), .Q(fracta[24])
         );
  DFF_X2 u1_fracta_out_reg_25_ ( .D(u1_fracta_s[25]), .CK(clk), .Q(fracta[25])
         );
  DFF_X2 u1_fracta_out_reg_26_ ( .D(u1_fracta_s[26]), .CK(clk), .Q(fracta[26])
         );
  DFF_X2 fract_out_q_reg_0_ ( .D(n5286), .CK(clk), .Q(fract_out_q[0]) );
  DFF_X2 fract_out_q_reg_1_ ( .D(n5285), .CK(clk), .Q(fract_out_q[1]) );
  DFF_X2 fract_out_q_reg_2_ ( .D(n5284), .CK(clk), .Q(fract_out_q[2]) );
  DFF_X2 fract_out_q_reg_3_ ( .D(n5283), .CK(clk), .QN(n2636) );
  DFF_X2 fract_out_q_reg_4_ ( .D(n5282), .CK(clk), .QN(n2635) );
  DFF_X2 fract_out_q_reg_5_ ( .D(n5281), .CK(clk), .Q(fract_out_q[5]) );
  DFF_X2 fract_out_q_reg_6_ ( .D(n5280), .CK(clk), .Q(fract_out_q[6]) );
  DFF_X2 fract_out_q_reg_7_ ( .D(n5279), .CK(clk), .Q(fract_out_q[7]) );
  DFF_X2 fract_out_q_reg_8_ ( .D(n5278), .CK(clk), .Q(fract_out_q[8]) );
  DFF_X2 fract_out_q_reg_9_ ( .D(n5277), .CK(clk), .QN(n2633) );
  DFF_X2 fract_out_q_reg_10_ ( .D(n5276), .CK(clk), .QN(n2646) );
  DFF_X2 fract_out_q_reg_11_ ( .D(n5275), .CK(clk), .Q(fract_out_q[11]) );
  DFF_X2 fract_out_q_reg_12_ ( .D(n5274), .CK(clk), .Q(fract_out_q[12]) );
  DFF_X2 fract_out_q_reg_13_ ( .D(n5273), .CK(clk), .Q(fract_out_q[13]) );
  DFF_X2 fract_out_q_reg_14_ ( .D(n5272), .CK(clk), .Q(fract_out_q[14]) );
  DFF_X2 fract_out_q_reg_15_ ( .D(n5271), .CK(clk), .QN(n2634) );
  DFF_X2 fract_out_q_reg_16_ ( .D(n5270), .CK(clk), .QN(n2629) );
  DFF_X2 fract_out_q_reg_17_ ( .D(n5269), .CK(clk), .QN(n2628) );
  DFF_X2 fract_out_q_reg_18_ ( .D(n5268), .CK(clk), .QN(n2647) );
  DFF_X2 fract_out_q_reg_21_ ( .D(n5265), .CK(clk), .Q(fract_out_q[21]) );
  DFF_X2 fract_out_q_reg_22_ ( .D(n5264), .CK(clk), .QN(n2630) );
  DFF_X2 fract_out_q_reg_23_ ( .D(n5263), .CK(clk), .QN(n2631) );
  DFF_X2 fract_out_q_reg_24_ ( .D(n5262), .CK(clk), .QN(n2627) );
  DFF_X2 fract_out_q_reg_25_ ( .D(n5261), .CK(clk), .QN(n2632) );
  DFF_X2 fract_out_q_reg_26_ ( .D(n5260), .CK(clk), .Q(fract_out_q[26]) );
  DFF_X2 fract_out_q_reg_27_ ( .D(n5259), .CK(clk), .Q(fract_out_q[27]) );
  DFF_X2 u1_exp_dn_out_reg_0_ ( .D(u1_N37), .CK(clk), .Q(exp_fasu[0]) );
  DFF_X2 u1_exp_dn_out_reg_1_ ( .D(u1_N38), .CK(clk), .Q(exp_fasu[1]) );
  DFF_X2 u1_exp_dn_out_reg_2_ ( .D(u1_N39), .CK(clk), .Q(exp_fasu[2]) );
  DFF_X2 u1_exp_dn_out_reg_3_ ( .D(u1_N40), .CK(clk), .Q(exp_fasu[3]) );
  DFF_X2 u1_exp_dn_out_reg_4_ ( .D(u1_N41), .CK(clk), .Q(exp_fasu[4]) );
  DFF_X2 u1_exp_dn_out_reg_5_ ( .D(u1_N42), .CK(clk), .Q(exp_fasu[5]) );
  DFF_X2 u1_exp_dn_out_reg_6_ ( .D(u1_N43), .CK(clk), .Q(exp_fasu[6]) );
  DFF_X2 u1_exp_dn_out_reg_7_ ( .D(u1_N44), .CK(clk), .Q(exp_fasu[7]) );
  DFF_X2 u2_sign_exe_reg ( .D(u2_N97), .CK(clk), .Q(sign_exe) );
  DFF_X2 sign_exe_r_reg ( .D(sign_exe), .CK(clk), .Q(sign_exe_r) );
  DFF_X2 u2_sign_reg ( .D(u2_sign_d), .CK(clk), .Q(sign_mul), .QN(n2734) );
  DFF_X2 sign_mul_r_reg ( .D(sign_mul), .CK(clk), .Q(sign_mul_r) );
  DFF_X2 sign_reg ( .D(N441), .CK(clk), .Q(sign), .QN(n2676) );
  DFF_X2 fract_i2f_reg_47_ ( .D(N421), .CK(clk), .Q(fract_i2f[47]) );
  DFF_X2 fract_i2f_reg_46_ ( .D(N420), .CK(clk), .Q(fract_i2f[46]) );
  DFF_X2 fract_i2f_reg_45_ ( .D(N419), .CK(clk), .Q(fract_i2f[45]) );
  DFF_X2 fract_i2f_reg_44_ ( .D(N418), .CK(clk), .Q(fract_i2f[44]) );
  DFF_X2 fract_i2f_reg_43_ ( .D(N417), .CK(clk), .Q(fract_i2f[43]) );
  DFF_X2 fract_i2f_reg_42_ ( .D(N416), .CK(clk), .Q(fract_i2f[42]) );
  DFF_X2 fract_i2f_reg_41_ ( .D(N415), .CK(clk), .Q(fract_i2f[41]) );
  DFF_X2 fract_i2f_reg_40_ ( .D(N414), .CK(clk), .Q(fract_i2f[40]) );
  DFF_X2 fract_i2f_reg_39_ ( .D(N413), .CK(clk), .Q(fract_i2f[39]) );
  DFF_X2 fract_i2f_reg_38_ ( .D(N412), .CK(clk), .Q(fract_i2f[38]) );
  DFF_X2 fract_i2f_reg_37_ ( .D(N411), .CK(clk), .Q(fract_i2f[37]) );
  DFF_X2 fract_i2f_reg_36_ ( .D(N410), .CK(clk), .Q(fract_i2f[36]) );
  DFF_X2 fract_i2f_reg_35_ ( .D(N409), .CK(clk), .Q(fract_i2f[35]) );
  DFF_X2 fract_i2f_reg_34_ ( .D(N408), .CK(clk), .Q(fract_i2f[34]) );
  DFF_X2 fract_i2f_reg_33_ ( .D(N407), .CK(clk), .Q(fract_i2f[33]) );
  DFF_X2 fract_i2f_reg_32_ ( .D(N406), .CK(clk), .Q(fract_i2f[32]) );
  DFF_X2 fract_i2f_reg_31_ ( .D(N405), .CK(clk), .Q(fract_i2f[31]) );
  DFF_X2 fract_i2f_reg_30_ ( .D(N404), .CK(clk), .Q(fract_i2f[30]) );
  DFF_X2 fract_i2f_reg_29_ ( .D(N403), .CK(clk), .QN(n3045) );
  DFF_X2 fract_i2f_reg_28_ ( .D(N402), .CK(clk), .Q(fract_i2f[28]) );
  DFF_X2 fract_i2f_reg_27_ ( .D(N401), .CK(clk), .Q(fract_i2f[27]) );
  DFF_X2 fract_i2f_reg_26_ ( .D(N400), .CK(clk), .Q(fract_i2f[26]) );
  DFF_X2 fract_i2f_reg_25_ ( .D(N399), .CK(clk), .Q(fract_i2f[25]) );
  DFF_X2 fract_i2f_reg_24_ ( .D(N398), .CK(clk), .Q(fract_i2f[24]) );
  DFF_X2 fract_i2f_reg_23_ ( .D(N397), .CK(clk), .Q(fract_i2f[23]) );
  DFF_X2 fract_i2f_reg_22_ ( .D(N396), .CK(clk), .Q(fract_i2f[22]) );
  DFF_X2 fract_i2f_reg_21_ ( .D(N395), .CK(clk), .Q(fract_i2f[21]) );
  DFF_X2 fract_i2f_reg_20_ ( .D(N394), .CK(clk), .Q(fract_i2f[20]) );
  DFF_X2 fract_i2f_reg_19_ ( .D(N393), .CK(clk), .Q(fract_i2f[19]) );
  DFF_X2 fract_i2f_reg_18_ ( .D(N392), .CK(clk), .Q(fract_i2f[18]) );
  DFF_X2 fract_i2f_reg_17_ ( .D(N391), .CK(clk), .Q(fract_i2f[17]) );
  DFF_X2 fract_i2f_reg_16_ ( .D(n5237), .CK(clk), .Q(fract_i2f[16]) );
  DFF_X2 fract_i2f_reg_15_ ( .D(n5238), .CK(clk), .Q(fract_i2f[15]) );
  DFF_X2 fract_i2f_reg_14_ ( .D(n5239), .CK(clk), .Q(fract_i2f[14]) );
  DFF_X2 fract_i2f_reg_13_ ( .D(n5240), .CK(clk), .Q(fract_i2f[13]) );
  DFF_X2 fract_i2f_reg_12_ ( .D(n5241), .CK(clk), .Q(fract_i2f[12]) );
  DFF_X2 fract_i2f_reg_11_ ( .D(n5242), .CK(clk), .Q(fract_i2f[11]) );
  DFF_X2 fract_i2f_reg_10_ ( .D(n5243), .CK(clk), .Q(fract_i2f[10]) );
  DFF_X2 fract_i2f_reg_9_ ( .D(n5244), .CK(clk), .Q(fract_i2f[9]) );
  DFF_X2 fract_i2f_reg_8_ ( .D(n5245), .CK(clk), .Q(fract_i2f[8]) );
  DFF_X2 fract_i2f_reg_7_ ( .D(n5246), .CK(clk), .Q(fract_i2f[7]) );
  DFF_X2 fract_i2f_reg_6_ ( .D(n5247), .CK(clk), .Q(fract_i2f[6]) );
  DFF_X2 fract_i2f_reg_5_ ( .D(n5248), .CK(clk), .Q(fract_i2f[5]) );
  DFF_X2 fract_i2f_reg_4_ ( .D(n5249), .CK(clk), .Q(fract_i2f[4]) );
  DFF_X2 fract_i2f_reg_3_ ( .D(n5250), .CK(clk), .Q(fract_i2f[3]) );
  DFF_X2 fract_i2f_reg_2_ ( .D(n5251), .CK(clk), .Q(fract_i2f[2]) );
  DFF_X2 fract_i2f_reg_1_ ( .D(n5252), .CK(clk), .Q(fract_i2f[1]) );
  DFF_X2 fract_i2f_reg_0_ ( .D(n5320), .CK(clk), .Q(fract_i2f[0]) );
  DFF_X2 u2_inf_reg ( .D(u2_N90), .CK(clk), .Q(inf_mul) );
  DFF_X2 inf_mul_r_reg ( .D(inf_mul), .CK(clk), .QN(n2605) );
  DFF_X2 u2_underflow_reg_0_ ( .D(n2739), .CK(clk), .Q(underflow_fmul_d[0]) );
  DFF_X2 underflow_fmul_r_reg_0_ ( .D(underflow_fmul_d[0]), .CK(clk), .Q(
        underflow_fmul_r[0]) );
  DFF_X2 u2_underflow_reg_1_ ( .D(u2_underflow_d[1]), .CK(clk), .Q(
        underflow_fmul_d[1]) );
  DFF_X2 underflow_fmul_r_reg_1_ ( .D(underflow_fmul_d[1]), .CK(clk), .Q(
        underflow_fmul_r[1]) );
  DFF_X2 u2_underflow_reg_2_ ( .D(u2_underflow_d[2]), .CK(clk), .Q(
        underflow_fmul_d[2]) );
  DFF_X2 underflow_fmul_r_reg_2_ ( .D(underflow_fmul_d[2]), .CK(clk), .QN(
        n2762) );
  DFF_X2 u2_exp_ovf_reg_0_ ( .D(u2_exp_ovf_d_0_), .CK(clk), .Q(exp_ovf[0]) );
  DFF_X2 exp_ovf_r_reg_0_ ( .D(exp_ovf[0]), .CK(clk), .Q(exp_ovf_r_0_), .QN(
        n2674) );
  DFF_X2 u2_exp_ovf_reg_1_ ( .D(u2_exp_ovf_d_1_), .CK(clk), .Q(exp_ovf[1]) );
  DFF_X2 exp_ovf_r_reg_1_ ( .D(exp_ovf[1]), .CK(clk), .QN(n2747) );
  DFF_X2 exp_r_reg_0_ ( .D(N214), .CK(clk), .QN(net92065) );
  DFF_X2 exp_r_reg_1_ ( .D(N215), .CK(clk), .QN(n2956) );
  DFF_X2 exp_r_reg_2_ ( .D(N216), .CK(clk), .QN(n2916) );
  DFF_X2 exp_r_reg_3_ ( .D(N217), .CK(clk), .Q(exp_r[3]), .QN(n2579) );
  DFF_X2 exp_r_reg_4_ ( .D(N218), .CK(clk), .Q(exp_r[4]), .QN(n2908) );
  DFF_X2 exp_r_reg_5_ ( .D(N219), .CK(clk), .Q(exp_r[5]), .QN(net95297) );
  DFF_X2 exp_r_reg_6_ ( .D(N220), .CK(clk), .Q(exp_r[6]), .QN(n2618) );
  DFF_X2 exp_r_reg_7_ ( .D(N221), .CK(clk), .QN(n2668) );
  DFF_X2 inf_mul2_reg ( .D(N540), .CK(clk), .QN(n2737) );
  DFF_X2 u5_prod1_reg_0_ ( .D(u5_N0), .CK(clk), .Q(u5_prod1[0]) );
  DFF_X2 u5_prod_reg_0_ ( .D(u5_prod1[0]), .CK(clk), .Q(prod[0]) );
  DFF_X2 u5_prod1_reg_1_ ( .D(u5_N1), .CK(clk), .Q(u5_prod1[1]) );
  DFF_X2 u5_prod_reg_1_ ( .D(u5_prod1[1]), .CK(clk), .Q(prod[1]) );
  DFF_X2 u5_prod1_reg_2_ ( .D(u5_N2), .CK(clk), .Q(u5_prod1[2]) );
  DFF_X2 u5_prod_reg_2_ ( .D(u5_prod1[2]), .CK(clk), .Q(prod[2]) );
  DFF_X2 u5_prod1_reg_3_ ( .D(u5_N3), .CK(clk), .Q(u5_prod1[3]) );
  DFF_X2 u5_prod_reg_3_ ( .D(u5_prod1[3]), .CK(clk), .Q(prod[3]) );
  DFF_X2 u5_prod1_reg_4_ ( .D(u5_N4), .CK(clk), .Q(u5_prod1[4]) );
  DFF_X2 u5_prod_reg_4_ ( .D(u5_prod1[4]), .CK(clk), .Q(prod[4]) );
  DFF_X2 u5_prod1_reg_5_ ( .D(u5_N5), .CK(clk), .Q(u5_prod1[5]) );
  DFF_X2 u5_prod_reg_5_ ( .D(u5_prod1[5]), .CK(clk), .Q(prod[5]) );
  DFF_X2 u5_prod1_reg_6_ ( .D(u5_N6), .CK(clk), .Q(u5_prod1[6]) );
  DFF_X2 u5_prod_reg_6_ ( .D(u5_prod1[6]), .CK(clk), .Q(prod[6]) );
  DFF_X2 u5_prod1_reg_7_ ( .D(u5_N7), .CK(clk), .Q(u5_prod1[7]) );
  DFF_X2 u5_prod_reg_7_ ( .D(u5_prod1[7]), .CK(clk), .Q(prod[7]) );
  DFF_X2 u5_prod1_reg_8_ ( .D(u5_N8), .CK(clk), .Q(u5_prod1[8]) );
  DFF_X2 u5_prod_reg_8_ ( .D(u5_prod1[8]), .CK(clk), .Q(prod[8]) );
  DFF_X2 u5_prod1_reg_9_ ( .D(u5_N9), .CK(clk), .Q(u5_prod1[9]) );
  DFF_X2 u5_prod_reg_9_ ( .D(u5_prod1[9]), .CK(clk), .Q(prod[9]) );
  DFF_X2 u5_prod1_reg_10_ ( .D(u5_N10), .CK(clk), .Q(u5_prod1[10]) );
  DFF_X2 u5_prod_reg_10_ ( .D(u5_prod1[10]), .CK(clk), .Q(prod[10]) );
  DFF_X2 u5_prod1_reg_11_ ( .D(u5_N11), .CK(clk), .Q(u5_prod1[11]) );
  DFF_X2 u5_prod_reg_11_ ( .D(u5_prod1[11]), .CK(clk), .Q(prod[11]) );
  DFF_X2 u5_prod1_reg_12_ ( .D(u5_N12), .CK(clk), .Q(u5_prod1[12]) );
  DFF_X2 u5_prod_reg_12_ ( .D(u5_prod1[12]), .CK(clk), .Q(prod[12]) );
  DFF_X2 u5_prod1_reg_13_ ( .D(u5_N13), .CK(clk), .Q(u5_prod1[13]) );
  DFF_X2 u5_prod_reg_13_ ( .D(u5_prod1[13]), .CK(clk), .Q(prod[13]) );
  DFF_X2 u5_prod1_reg_14_ ( .D(u5_N14), .CK(clk), .Q(u5_prod1[14]) );
  DFF_X2 u5_prod_reg_14_ ( .D(u5_prod1[14]), .CK(clk), .Q(prod[14]) );
  DFF_X2 u5_prod1_reg_15_ ( .D(u5_N15), .CK(clk), .Q(u5_prod1[15]) );
  DFF_X2 u5_prod_reg_15_ ( .D(u5_prod1[15]), .CK(clk), .Q(prod[15]) );
  DFF_X2 u5_prod1_reg_16_ ( .D(u5_N16), .CK(clk), .Q(u5_prod1[16]) );
  DFF_X2 u5_prod_reg_16_ ( .D(u5_prod1[16]), .CK(clk), .Q(prod[16]) );
  DFF_X2 u5_prod1_reg_17_ ( .D(u5_N17), .CK(clk), .Q(u5_prod1[17]) );
  DFF_X2 u5_prod_reg_17_ ( .D(u5_prod1[17]), .CK(clk), .Q(prod[17]) );
  DFF_X2 u5_prod1_reg_18_ ( .D(u5_N18), .CK(clk), .Q(u5_prod1[18]) );
  DFF_X2 u5_prod_reg_18_ ( .D(u5_prod1[18]), .CK(clk), .Q(prod[18]) );
  DFF_X2 u5_prod_reg_19_ ( .D(u5_prod1[19]), .CK(clk), .Q(prod[19]) );
  DFF_X2 u5_prod_reg_20_ ( .D(u5_prod1[20]), .CK(clk), .Q(prod[20]) );
  DFF_X2 u5_prod_reg_21_ ( .D(u5_prod1[21]), .CK(clk), .Q(prod[21]) );
  DFF_X2 u5_prod1_reg_22_ ( .D(u5_N22), .CK(clk), .Q(u5_prod1[22]) );
  DFF_X2 u5_prod1_reg_23_ ( .D(u5_N23), .CK(clk), .Q(u5_prod1[23]) );
  DFF_X2 u5_prod_reg_23_ ( .D(u5_prod1[23]), .CK(clk), .Q(prod[23]) );
  DFF_X2 u5_prod1_reg_24_ ( .D(u5_N24), .CK(clk), .Q(u5_prod1[24]) );
  DFF_X2 u5_prod_reg_24_ ( .D(u5_prod1[24]), .CK(clk), .Q(prod[24]), .QN(n2642) );
  DFF_X2 u5_prod1_reg_26_ ( .D(u5_N26), .CK(clk), .Q(u5_prod1[26]) );
  DFF_X2 u5_prod_reg_26_ ( .D(u5_prod1[26]), .CK(clk), .Q(prod[26]) );
  DFF_X2 u5_prod1_reg_27_ ( .D(u5_N27), .CK(clk), .Q(u5_prod1[27]) );
  DFF_X2 u5_prod_reg_27_ ( .D(u5_prod1[27]), .CK(clk), .Q(prod[27]) );
  DFF_X2 u5_prod1_reg_28_ ( .D(u5_N28), .CK(clk), .Q(u5_prod1[28]) );
  DFF_X2 u5_prod_reg_28_ ( .D(u5_prod1[28]), .CK(clk), .Q(prod[28]) );
  DFF_X2 u5_prod1_reg_29_ ( .D(u5_N29), .CK(clk), .Q(u5_prod1[29]) );
  DFF_X2 u5_prod_reg_29_ ( .D(u5_prod1[29]), .CK(clk), .Q(prod[29]), .QN(n3070) );
  DFF_X2 u5_prod_reg_30_ ( .D(u5_prod1[30]), .CK(clk), .Q(prod[30]) );
  DFF_X2 u5_prod1_reg_31_ ( .D(u5_N31), .CK(clk), .Q(u5_prod1[31]) );
  DFF_X2 u5_prod1_reg_32_ ( .D(u5_N32), .CK(clk), .Q(u5_prod1[32]) );
  DFF_X2 u5_prod1_reg_33_ ( .D(u5_N33), .CK(clk), .Q(u5_prod1[33]) );
  DFF_X2 u5_prod1_reg_34_ ( .D(u5_N34), .CK(clk), .Q(u5_prod1[34]) );
  DFF_X2 u5_prod_reg_36_ ( .D(u5_prod1[36]), .CK(clk), .Q(prod[36]), .QN(n2625) );
  DFF_X2 u5_prod_reg_37_ ( .D(u5_prod1[37]), .CK(clk), .Q(prod[37]) );
  DFF_X2 u5_prod_reg_38_ ( .D(u5_prod1[38]), .CK(clk), .Q(prod[38]) );
  DFF_X2 u5_prod_reg_39_ ( .D(u5_prod1[39]), .CK(clk), .Q(prod[39]) );
  DFF_X2 u5_prod_reg_40_ ( .D(u5_prod1[40]), .CK(clk), .Q(prod[40]) );
  DFF_X2 u5_prod_reg_41_ ( .D(u5_prod1[41]), .CK(clk), .Q(prod[41]) );
  DFF_X2 u5_prod_reg_42_ ( .D(u5_prod1[42]), .CK(clk), .Q(prod[42]) );
  DFF_X2 u5_prod_reg_43_ ( .D(u5_prod1[43]), .CK(clk), .Q(prod[43]) );
  DFF_X2 u5_prod_reg_44_ ( .D(u5_prod1[44]), .CK(clk), .Q(prod[44]) );
  DFF_X2 u5_prod_reg_45_ ( .D(u5_prod1[45]), .CK(clk), .Q(prod[45]) );
  DFF_X2 u5_prod_reg_46_ ( .D(u5_prod1[46]), .CK(clk), .Q(prod[46]) );
  DFF_X2 u6_remainder_reg_0_ ( .D(u6_N0), .CK(clk), .Q(u6_remainder[0]) );
  DFF_X2 u6_rem_reg_0_ ( .D(u6_remainder[0]), .CK(clk), .Q(remainder[0]) );
  DFF_X2 u6_remainder_reg_1_ ( .D(u6_N1), .CK(clk), .Q(u6_remainder[1]) );
  DFF_X2 u6_rem_reg_1_ ( .D(u6_remainder[1]), .CK(clk), .Q(remainder[1]) );
  DFF_X2 u6_remainder_reg_2_ ( .D(u6_N2), .CK(clk), .Q(u6_remainder[2]) );
  DFF_X2 u6_rem_reg_2_ ( .D(u6_remainder[2]), .CK(clk), .Q(remainder[2]) );
  DFF_X2 u6_remainder_reg_3_ ( .D(u6_N3), .CK(clk), .Q(u6_remainder[3]) );
  DFF_X2 u6_rem_reg_3_ ( .D(u6_remainder[3]), .CK(clk), .Q(remainder[3]) );
  DFF_X2 u6_remainder_reg_4_ ( .D(u6_N4), .CK(clk), .Q(u6_remainder[4]) );
  DFF_X2 u6_rem_reg_4_ ( .D(u6_remainder[4]), .CK(clk), .Q(remainder[4]) );
  DFF_X2 u6_remainder_reg_5_ ( .D(u6_N5), .CK(clk), .Q(u6_remainder[5]) );
  DFF_X2 u6_rem_reg_5_ ( .D(u6_remainder[5]), .CK(clk), .Q(remainder[5]) );
  DFF_X2 u6_remainder_reg_6_ ( .D(u6_N6), .CK(clk), .Q(u6_remainder[6]) );
  DFF_X2 u6_rem_reg_6_ ( .D(u6_remainder[6]), .CK(clk), .QN(n2732) );
  DFF_X2 u6_remainder_reg_7_ ( .D(u6_N7), .CK(clk), .Q(u6_remainder[7]) );
  DFF_X2 u6_rem_reg_7_ ( .D(u6_remainder[7]), .CK(clk), .Q(remainder[7]) );
  DFF_X2 u6_remainder_reg_8_ ( .D(u6_N8), .CK(clk), .Q(u6_remainder[8]) );
  DFF_X2 u6_rem_reg_8_ ( .D(u6_remainder[8]), .CK(clk), .Q(remainder[8]) );
  DFF_X2 u6_remainder_reg_9_ ( .D(u6_N9), .CK(clk), .Q(u6_remainder[9]) );
  DFF_X2 u6_rem_reg_9_ ( .D(u6_remainder[9]), .CK(clk), .Q(remainder[9]) );
  DFF_X2 u6_remainder_reg_10_ ( .D(u6_N10), .CK(clk), .Q(u6_remainder[10]) );
  DFF_X2 u6_rem_reg_10_ ( .D(u6_remainder[10]), .CK(clk), .Q(remainder[10]) );
  DFF_X2 u6_remainder_reg_11_ ( .D(n2982), .CK(clk), .Q(u6_remainder[11]) );
  DFF_X2 u6_rem_reg_11_ ( .D(u6_remainder[11]), .CK(clk), .Q(remainder[11]) );
  DFF_X2 u6_remainder_reg_12_ ( .D(n2986), .CK(clk), .Q(u6_remainder[12]) );
  DFF_X2 u6_rem_reg_12_ ( .D(u6_remainder[12]), .CK(clk), .Q(remainder[12]) );
  DFF_X2 u6_remainder_reg_13_ ( .D(u6_N13), .CK(clk), .Q(u6_remainder[13]) );
  DFF_X2 u6_rem_reg_13_ ( .D(u6_remainder[13]), .CK(clk), .Q(remainder[13]) );
  DFF_X2 u6_remainder_reg_14_ ( .D(n2672), .CK(clk), .Q(u6_remainder[14]) );
  DFF_X2 u6_rem_reg_14_ ( .D(u6_remainder[14]), .CK(clk), .Q(remainder[14]) );
  DFF_X2 u6_remainder_reg_15_ ( .D(u6_N15), .CK(clk), .Q(u6_remainder[15]) );
  DFF_X2 u6_rem_reg_15_ ( .D(u6_remainder[15]), .CK(clk), .Q(remainder[15]) );
  DFF_X2 u6_remainder_reg_16_ ( .D(n2963), .CK(clk), .Q(u6_remainder[16]) );
  DFF_X2 u6_rem_reg_16_ ( .D(u6_remainder[16]), .CK(clk), .Q(remainder[16]) );
  DFF_X2 u6_remainder_reg_17_ ( .D(u6_N17), .CK(clk), .Q(u6_remainder[17]) );
  DFF_X2 u6_rem_reg_17_ ( .D(u6_remainder[17]), .CK(clk), .Q(remainder[17]) );
  DFF_X2 u6_remainder_reg_18_ ( .D(u6_N18), .CK(clk), .Q(u6_remainder[18]) );
  DFF_X2 u6_rem_reg_18_ ( .D(u6_remainder[18]), .CK(clk), .Q(remainder[18]) );
  DFF_X2 u6_remainder_reg_19_ ( .D(n2968), .CK(clk), .Q(u6_remainder[19]) );
  DFF_X2 u6_rem_reg_19_ ( .D(u6_remainder[19]), .CK(clk), .Q(remainder[19]) );
  DFF_X2 u6_remainder_reg_20_ ( .D(n3040), .CK(clk), .Q(u6_remainder[20]) );
  DFF_X2 u6_rem_reg_20_ ( .D(u6_remainder[20]), .CK(clk), .Q(remainder[20]) );
  DFF_X2 u6_remainder_reg_21_ ( .D(n3049), .CK(clk), .Q(u6_remainder[21]) );
  DFF_X2 u6_rem_reg_21_ ( .D(u6_remainder[21]), .CK(clk), .Q(remainder[21]) );
  DFF_X2 u6_remainder_reg_22_ ( .D(u6_N22), .CK(clk), .Q(u6_remainder[22]) );
  DFF_X2 u6_rem_reg_22_ ( .D(u6_remainder[22]), .CK(clk), .Q(remainder[22]) );
  DFF_X2 u6_remainder_reg_23_ ( .D(n2930), .CK(clk), .Q(u6_remainder[23]) );
  DFF_X2 u6_rem_reg_23_ ( .D(u6_remainder[23]), .CK(clk), .Q(remainder[23]) );
  DFF_X2 u6_remainder_reg_26_ ( .D(u6_N26), .CK(clk), .Q(u6_remainder[26]) );
  DFF_X2 u6_rem_reg_26_ ( .D(u6_remainder[26]), .CK(clk), .Q(remainder[26]) );
  DFF_X2 u6_remainder_reg_27_ ( .D(u6_N27), .CK(clk), .Q(u6_remainder[27]) );
  DFF_X2 u6_rem_reg_27_ ( .D(u6_remainder[27]), .CK(clk), .Q(remainder[27]) );
  DFF_X2 u6_remainder_reg_28_ ( .D(u6_N28), .CK(clk), .Q(u6_remainder[28]) );
  DFF_X2 u6_rem_reg_28_ ( .D(u6_remainder[28]), .CK(clk), .Q(remainder[28]) );
  DFF_X2 u6_remainder_reg_29_ ( .D(u6_N29), .CK(clk), .Q(u6_remainder[29]) );
  DFF_X2 u6_rem_reg_29_ ( .D(u6_remainder[29]), .CK(clk), .Q(remainder[29]) );
  DFF_X2 u6_remainder_reg_30_ ( .D(u6_N30), .CK(clk), .Q(u6_remainder[30]) );
  DFF_X2 u6_rem_reg_30_ ( .D(u6_remainder[30]), .CK(clk), .Q(remainder[30]) );
  DFF_X2 u6_remainder_reg_31_ ( .D(u6_N31), .CK(clk), .Q(u6_remainder[31]) );
  DFF_X2 u6_rem_reg_31_ ( .D(u6_remainder[31]), .CK(clk), .QN(n2733) );
  DFF_X2 u6_remainder_reg_32_ ( .D(u6_N32), .CK(clk), .Q(u6_remainder[32]) );
  DFF_X2 u6_rem_reg_32_ ( .D(u6_remainder[32]), .CK(clk), .Q(remainder[32]) );
  DFF_X2 u6_remainder_reg_33_ ( .D(u6_N33), .CK(clk), .Q(u6_remainder[33]) );
  DFF_X2 u6_rem_reg_33_ ( .D(u6_remainder[33]), .CK(clk), .Q(remainder[33]) );
  DFF_X2 u6_remainder_reg_34_ ( .D(u6_N34), .CK(clk), .Q(u6_remainder[34]) );
  DFF_X2 u6_rem_reg_34_ ( .D(u6_remainder[34]), .CK(clk), .Q(remainder[34]) );
  DFF_X2 u6_remainder_reg_35_ ( .D(u6_N35), .CK(clk), .Q(u6_remainder[35]) );
  DFF_X2 u6_rem_reg_35_ ( .D(u6_remainder[35]), .CK(clk), .Q(remainder[35]) );
  DFF_X2 u6_remainder_reg_36_ ( .D(u6_N36), .CK(clk), .Q(u6_remainder[36]) );
  DFF_X2 u6_rem_reg_36_ ( .D(u6_remainder[36]), .CK(clk), .Q(remainder[36]) );
  DFF_X2 u6_remainder_reg_37_ ( .D(u6_N37), .CK(clk), .Q(u6_remainder[37]) );
  DFF_X2 u6_rem_reg_37_ ( .D(u6_remainder[37]), .CK(clk), .Q(remainder[37]) );
  DFF_X2 u6_remainder_reg_38_ ( .D(u6_N38), .CK(clk), .Q(u6_remainder[38]) );
  DFF_X2 u6_rem_reg_38_ ( .D(u6_remainder[38]), .CK(clk), .Q(remainder[38]) );
  DFF_X2 u6_remainder_reg_39_ ( .D(u6_N39), .CK(clk), .Q(u6_remainder[39]) );
  DFF_X2 u6_rem_reg_39_ ( .D(u6_remainder[39]), .CK(clk), .Q(remainder[39]) );
  DFF_X2 u6_remainder_reg_40_ ( .D(u6_N40), .CK(clk), .Q(u6_remainder[40]) );
  DFF_X2 u6_rem_reg_40_ ( .D(u6_remainder[40]), .CK(clk), .Q(remainder[40]) );
  DFF_X2 u6_remainder_reg_41_ ( .D(u6_N41), .CK(clk), .Q(u6_remainder[41]) );
  DFF_X2 u6_rem_reg_41_ ( .D(u6_remainder[41]), .CK(clk), .Q(remainder[41]) );
  DFF_X2 u6_remainder_reg_42_ ( .D(u6_N42), .CK(clk), .Q(u6_remainder[42]) );
  DFF_X2 u6_rem_reg_42_ ( .D(u6_remainder[42]), .CK(clk), .Q(remainder[42]) );
  DFF_X2 u6_remainder_reg_43_ ( .D(u6_N43), .CK(clk), .Q(u6_remainder[43]) );
  DFF_X2 u6_rem_reg_43_ ( .D(u6_remainder[43]), .CK(clk), .Q(remainder[43]) );
  DFF_X2 u6_remainder_reg_44_ ( .D(u6_N44), .CK(clk), .Q(u6_remainder[44]) );
  DFF_X2 u6_rem_reg_44_ ( .D(u6_remainder[44]), .CK(clk), .Q(remainder[44]) );
  DFF_X2 u6_remainder_reg_45_ ( .D(u6_N45), .CK(clk), .Q(u6_remainder[45]) );
  DFF_X2 u6_rem_reg_45_ ( .D(u6_remainder[45]), .CK(clk), .Q(remainder[45]) );
  DFF_X2 u6_remainder_reg_46_ ( .D(u6_N46), .CK(clk), .Q(u6_remainder[46]) );
  DFF_X2 u6_rem_reg_46_ ( .D(u6_remainder[46]), .CK(clk), .Q(remainder[46]) );
  DFF_X2 u6_remainder_reg_47_ ( .D(u6_N47), .CK(clk), .Q(u6_remainder[47]) );
  DFF_X2 u6_rem_reg_47_ ( .D(u6_remainder[47]), .CK(clk), .Q(remainder[47]) );
  DFF_X2 u6_remainder_reg_48_ ( .D(u6_N48), .CK(clk), .Q(u6_remainder[48]) );
  DFF_X2 u6_rem_reg_48_ ( .D(u6_remainder[48]), .CK(clk), .Q(remainder[48]) );
  DFF_X2 u6_remainder_reg_49_ ( .D(u6_N49), .CK(clk), .Q(u6_remainder[49]) );
  DFF_X2 u6_rem_reg_49_ ( .D(u6_remainder[49]), .CK(clk), .Q(remainder[49]) );
  DFF_X2 u6_quo1_reg_0_ ( .D(u6_N0), .CK(clk), .Q(u6_quo1[0]) );
  DFF_X2 u6_quo_reg_0_ ( .D(u6_quo1[0]), .CK(clk), .Q(quo[0]) );
  DFF_X2 u6_quo1_reg_1_ ( .D(u6_N1), .CK(clk), .Q(u6_quo1[1]) );
  DFF_X2 u6_quo_reg_1_ ( .D(u6_quo1[1]), .CK(clk), .Q(quo[1]) );
  DFF_X2 u6_quo1_reg_2_ ( .D(u6_N2), .CK(clk), .Q(u6_quo1[2]) );
  DFF_X2 u6_quo_reg_2_ ( .D(u6_quo1[2]), .CK(clk), .Q(quo[2]), .QN(n2650) );
  DFF_X2 u6_quo1_reg_3_ ( .D(u6_N3), .CK(clk), .Q(u6_quo1[3]) );
  DFF_X2 u6_quo_reg_3_ ( .D(u6_quo1[3]), .CK(clk), .Q(quo[3]) );
  DFF_X2 u6_quo1_reg_4_ ( .D(u6_N4), .CK(clk), .Q(u6_quo1[4]) );
  DFF_X2 u6_quo_reg_4_ ( .D(u6_quo1[4]), .CK(clk), .Q(quo[4]) );
  DFF_X2 u6_quo1_reg_5_ ( .D(u6_N5), .CK(clk), .Q(u6_quo1[5]) );
  DFF_X2 u6_quo_reg_5_ ( .D(u6_quo1[5]), .CK(clk), .Q(quo[5]) );
  DFF_X2 u6_quo1_reg_6_ ( .D(u6_N6), .CK(clk), .Q(u6_quo1[6]) );
  DFF_X2 u6_quo_reg_6_ ( .D(u6_quo1[6]), .CK(clk), .Q(quo[6]) );
  DFF_X2 u6_quo1_reg_7_ ( .D(u6_N7), .CK(clk), .Q(u6_quo1[7]) );
  DFF_X2 u6_quo_reg_7_ ( .D(u6_quo1[7]), .CK(clk), .Q(quo[7]) );
  DFF_X2 u6_quo1_reg_8_ ( .D(u6_N8), .CK(clk), .Q(u6_quo1[8]) );
  DFF_X2 u6_quo_reg_8_ ( .D(u6_quo1[8]), .CK(clk), .Q(quo[8]) );
  DFF_X2 u6_quo1_reg_9_ ( .D(u6_N9), .CK(clk), .Q(u6_quo1[9]) );
  DFF_X2 u6_quo_reg_9_ ( .D(u6_quo1[9]), .CK(clk), .Q(quo[9]) );
  DFF_X2 u6_quo1_reg_10_ ( .D(u6_N10), .CK(clk), .Q(u6_quo1[10]) );
  DFF_X2 u6_quo_reg_10_ ( .D(u6_quo1[10]), .CK(clk), .Q(quo[10]) );
  DFF_X2 u6_quo1_reg_11_ ( .D(n2982), .CK(clk), .Q(u6_quo1[11]) );
  DFF_X2 u6_quo_reg_11_ ( .D(u6_quo1[11]), .CK(clk), .Q(quo[11]) );
  DFF_X2 u6_quo1_reg_12_ ( .D(n2986), .CK(clk), .Q(u6_quo1[12]) );
  DFF_X2 u6_quo_reg_12_ ( .D(u6_quo1[12]), .CK(clk), .Q(quo[12]) );
  DFF_X2 u6_quo1_reg_13_ ( .D(u6_N13), .CK(clk), .Q(u6_quo1[13]) );
  DFF_X2 u6_quo_reg_13_ ( .D(u6_quo1[13]), .CK(clk), .Q(quo[13]), .QN(n2639)
         );
  DFF_X2 u6_quo1_reg_14_ ( .D(n2672), .CK(clk), .Q(u6_quo1[14]) );
  DFF_X2 u6_quo_reg_14_ ( .D(u6_quo1[14]), .CK(clk), .Q(quo[14]) );
  DFF_X2 u6_quo1_reg_15_ ( .D(u6_N15), .CK(clk), .Q(u6_quo1[15]) );
  DFF_X2 u6_quo_reg_15_ ( .D(u6_quo1[15]), .CK(clk), .Q(quo[15]) );
  DFF_X2 u6_quo1_reg_16_ ( .D(n2963), .CK(clk), .Q(u6_quo1[16]) );
  DFF_X2 u6_quo_reg_16_ ( .D(u6_quo1[16]), .CK(clk), .Q(quo[16]) );
  DFF_X2 u6_quo1_reg_17_ ( .D(u6_N17), .CK(clk), .Q(u6_quo1[17]) );
  DFF_X2 u6_quo_reg_17_ ( .D(u6_quo1[17]), .CK(clk), .Q(quo[17]) );
  DFF_X2 u6_quo1_reg_18_ ( .D(u6_N18), .CK(clk), .Q(u6_quo1[18]) );
  DFF_X2 u6_quo_reg_18_ ( .D(u6_quo1[18]), .CK(clk), .Q(quo[18]) );
  DFF_X2 u6_quo1_reg_19_ ( .D(n2968), .CK(clk), .Q(u6_quo1[19]) );
  DFF_X2 u6_quo_reg_19_ ( .D(u6_quo1[19]), .CK(clk), .Q(quo[19]) );
  DFF_X2 u6_quo1_reg_20_ ( .D(n3040), .CK(clk), .Q(u6_quo1[20]) );
  DFF_X2 u6_quo_reg_20_ ( .D(u6_quo1[20]), .CK(clk), .Q(quo[20]) );
  DFF_X2 u6_quo1_reg_21_ ( .D(n3049), .CK(clk), .Q(u6_quo1[21]) );
  DFF_X2 u6_quo_reg_21_ ( .D(u6_quo1[21]), .CK(clk), .Q(quo[21]) );
  DFF_X2 u6_quo1_reg_22_ ( .D(u6_N22), .CK(clk), .Q(u6_quo1[22]) );
  DFF_X2 u6_quo_reg_22_ ( .D(u6_quo1[22]), .CK(clk), .Q(quo[22]), .QN(n2648)
         );
  DFF_X2 u6_quo1_reg_23_ ( .D(n2930), .CK(clk), .Q(u6_quo1[23]) );
  DFF_X2 u6_quo1_reg_26_ ( .D(u6_N26), .CK(clk), .Q(u6_quo1[26]) );
  DFF_X2 u6_quo_reg_26_ ( .D(u6_quo1[26]), .CK(clk), .Q(quo[26]) );
  DFF_X2 u6_quo1_reg_27_ ( .D(u6_N27), .CK(clk), .Q(u6_quo1[27]) );
  DFF_X2 u6_quo_reg_27_ ( .D(u6_quo1[27]), .CK(clk), .Q(quo[27]) );
  DFF_X2 u6_quo1_reg_28_ ( .D(u6_N28), .CK(clk), .Q(u6_quo1[28]) );
  DFF_X2 u6_quo_reg_28_ ( .D(u6_quo1[28]), .CK(clk), .QN(n2651) );
  DFF_X2 u6_quo1_reg_29_ ( .D(u6_N29), .CK(clk), .Q(u6_quo1[29]) );
  DFF_X2 u6_quo_reg_29_ ( .D(u6_quo1[29]), .CK(clk), .Q(quo[29]) );
  DFF_X2 u6_quo1_reg_30_ ( .D(u6_N30), .CK(clk), .Q(u6_quo1[30]) );
  DFF_X2 u6_quo_reg_30_ ( .D(u6_quo1[30]), .CK(clk), .Q(quo[30]) );
  DFF_X2 u6_quo1_reg_31_ ( .D(u6_N31), .CK(clk), .Q(u6_quo1[31]) );
  DFF_X2 u6_quo_reg_31_ ( .D(u6_quo1[31]), .CK(clk), .Q(quo[31]) );
  DFF_X2 u6_quo1_reg_32_ ( .D(u6_N32), .CK(clk), .Q(u6_quo1[32]) );
  DFF_X2 u6_quo_reg_32_ ( .D(u6_quo1[32]), .CK(clk), .Q(quo[32]) );
  DFF_X2 u6_quo1_reg_33_ ( .D(u6_N33), .CK(clk), .Q(u6_quo1[33]) );
  DFF_X2 u6_quo_reg_33_ ( .D(u6_quo1[33]), .CK(clk), .Q(quo[33]) );
  DFF_X2 u6_quo1_reg_34_ ( .D(u6_N34), .CK(clk), .Q(u6_quo1[34]) );
  DFF_X2 u6_quo_reg_34_ ( .D(u6_quo1[34]), .CK(clk), .Q(quo[34]) );
  DFF_X2 u6_quo1_reg_35_ ( .D(u6_N35), .CK(clk), .Q(u6_quo1[35]) );
  DFF_X2 u6_quo_reg_35_ ( .D(u6_quo1[35]), .CK(clk), .Q(quo[35]) );
  DFF_X2 u6_quo1_reg_36_ ( .D(u6_N36), .CK(clk), .Q(u6_quo1[36]) );
  DFF_X2 u6_quo_reg_36_ ( .D(u6_quo1[36]), .CK(clk), .Q(quo[36]) );
  DFF_X2 u6_quo1_reg_37_ ( .D(u6_N37), .CK(clk), .Q(u6_quo1[37]) );
  DFF_X2 u6_quo_reg_37_ ( .D(u6_quo1[37]), .CK(clk), .Q(quo[37]) );
  DFF_X2 u6_quo1_reg_38_ ( .D(u6_N38), .CK(clk), .Q(u6_quo1[38]) );
  DFF_X2 u6_quo_reg_38_ ( .D(u6_quo1[38]), .CK(clk), .Q(quo[38]) );
  DFF_X2 u6_quo1_reg_39_ ( .D(u6_N39), .CK(clk), .Q(u6_quo1[39]) );
  DFF_X2 u6_quo_reg_39_ ( .D(u6_quo1[39]), .CK(clk), .Q(quo[39]) );
  DFF_X2 u6_quo1_reg_40_ ( .D(u6_N40), .CK(clk), .Q(u6_quo1[40]) );
  DFF_X2 u6_quo_reg_40_ ( .D(u6_quo1[40]), .CK(clk), .Q(quo[40]) );
  DFF_X2 u6_quo1_reg_41_ ( .D(u6_N41), .CK(clk), .Q(u6_quo1[41]) );
  DFF_X2 u6_quo_reg_41_ ( .D(u6_quo1[41]), .CK(clk), .Q(quo[41]) );
  DFF_X2 u6_quo1_reg_42_ ( .D(u6_N42), .CK(clk), .Q(u6_quo1[42]) );
  DFF_X2 u6_quo_reg_42_ ( .D(u6_quo1[42]), .CK(clk), .Q(quo[42]) );
  DFF_X2 u6_quo1_reg_43_ ( .D(u6_N43), .CK(clk), .Q(u6_quo1[43]) );
  DFF_X2 u6_quo_reg_43_ ( .D(u6_quo1[43]), .CK(clk), .Q(quo[43]) );
  DFF_X2 u6_quo1_reg_44_ ( .D(u6_N44), .CK(clk), .Q(u6_quo1[44]) );
  DFF_X2 u6_quo_reg_44_ ( .D(u6_quo1[44]), .CK(clk), .Q(quo[44]) );
  DFF_X2 u6_quo1_reg_45_ ( .D(u6_N45), .CK(clk), .Q(u6_quo1[45]) );
  DFF_X2 u6_quo_reg_45_ ( .D(u6_quo1[45]), .CK(clk), .Q(quo[45]) );
  DFF_X2 u6_quo1_reg_46_ ( .D(u6_N46), .CK(clk), .Q(u6_quo1[46]) );
  DFF_X2 u6_quo_reg_46_ ( .D(u6_quo1[46]), .CK(clk), .Q(quo[46]) );
  DFF_X2 u6_quo1_reg_47_ ( .D(u6_N47), .CK(clk), .Q(u6_quo1[47]) );
  DFF_X2 u6_quo_reg_47_ ( .D(u6_quo1[47]), .CK(clk), .Q(quo[47]) );
  DFF_X2 u6_quo1_reg_48_ ( .D(u6_N48), .CK(clk), .Q(u6_quo1[48]) );
  DFF_X2 u6_quo_reg_48_ ( .D(u6_quo1[48]), .CK(clk), .QN(n2649) );
  DFF_X2 out_reg_23_ ( .D(N468), .CK(clk), .Q(out[23]) );
  DFF_X2 out_reg_29_ ( .D(n2520), .CK(clk), .Q(out[29]) );
  DFF_X2 out_reg_30_ ( .D(N475), .CK(clk), .Q(out[30]) );
  DFF_X2 out_reg_24_ ( .D(N469), .CK(clk), .Q(out[24]) );
  DFF_X2 out_reg_25_ ( .D(N470), .CK(clk), .Q(out[25]) );
  DFF_X2 out_reg_26_ ( .D(N471), .CK(clk), .Q(out[26]) );
  DFF_X2 out_reg_22_ ( .D(N467), .CK(clk), .Q(out[22]) );
  DFF_X2 out_reg_21_ ( .D(N466), .CK(clk), .Q(out[21]) );
  DFF_X2 out_reg_20_ ( .D(N465), .CK(clk), .Q(out[20]) );
  DFF_X2 out_reg_19_ ( .D(N464), .CK(clk), .Q(out[19]) );
  DFF_X2 out_reg_18_ ( .D(N463), .CK(clk), .Q(out[18]) );
  DFF_X2 out_reg_17_ ( .D(N462), .CK(clk), .Q(out[17]) );
  DFF_X2 out_reg_16_ ( .D(N461), .CK(clk), .Q(out[16]) );
  DFF_X2 out_reg_15_ ( .D(N460), .CK(clk), .Q(out[15]) );
  DFF_X2 out_reg_14_ ( .D(N459), .CK(clk), .Q(out[14]) );
  DFF_X2 out_reg_13_ ( .D(N458), .CK(clk), .Q(out[13]) );
  DFF_X2 out_reg_12_ ( .D(N457), .CK(clk), .Q(out[12]) );
  DFF_X2 out_reg_11_ ( .D(N456), .CK(clk), .Q(out[11]) );
  DFF_X2 out_reg_10_ ( .D(N455), .CK(clk), .Q(out[10]) );
  DFF_X2 out_reg_9_ ( .D(N454), .CK(clk), .Q(out[9]) );
  DFF_X2 out_reg_8_ ( .D(N453), .CK(clk), .Q(out[8]) );
  DFF_X2 out_reg_7_ ( .D(N452), .CK(clk), .Q(out[7]) );
  DFF_X2 out_reg_6_ ( .D(N451), .CK(clk), .Q(out[6]) );
  DFF_X2 out_reg_5_ ( .D(N450), .CK(clk), .Q(out[5]) );
  DFF_X2 out_reg_4_ ( .D(N449), .CK(clk), .Q(out[4]) );
  DFF_X2 out_reg_3_ ( .D(N448), .CK(clk), .Q(out[3]) );
  DFF_X2 out_reg_2_ ( .D(N447), .CK(clk), .Q(out[2]) );
  DFF_X2 out_reg_1_ ( .D(N446), .CK(clk), .Q(out[1]) );
  DFF_X2 ine_reg ( .D(N509), .CK(clk), .Q(ine) );
  DFF_X2 out_reg_0_ ( .D(N445), .CK(clk), .Q(out[0]) );
  DFF_X2 u6_quo1_reg_49_ ( .D(u6_N49), .CK(clk), .Q(u6_quo1[49]) );
  DFF_X1 u5_prod1_reg_38_ ( .D(u5_N38), .CK(clk), .Q(u5_prod1[38]) );
  DFF_X2 opb_r_reg_30_ ( .D(opb[30]), .CK(clk), .Q(opb_r[30]), .QN(n2996) );
  DFF_X1 underflow_reg ( .D(N522), .CK(clk), .Q(underflow) );
  DFF_X2 fpu_op_r3_reg_0_ ( .D(fpu_op_r2[0]), .CK(clk), .Q(net91406), .QN(
        net86294) );
  DFF_X2 fract_out_q_reg_20_ ( .D(n5266), .CK(clk), .QN(n3043) );
  DFF_X2 fract_out_q_reg_19_ ( .D(n5267), .CK(clk), .QN(n3042) );
  DFF_X1 u5_prod1_reg_39_ ( .D(u5_N39), .CK(clk), .Q(u5_prod1[39]) );
  DFF_X1 u5_prod1_reg_42_ ( .D(u5_N42), .CK(clk), .Q(u5_prod1[42]) );
  DFF_X1 u5_prod1_reg_40_ ( .D(u5_N40), .CK(clk), .Q(u5_prod1[40]) );
  DFF_X1 u5_prod1_reg_41_ ( .D(u5_N41), .CK(clk), .Q(u5_prod1[41]) );
  DFF_X1 u5_prod1_reg_46_ ( .D(u5_N46), .CK(clk), .Q(u5_prod1[46]) );
  DFF_X1 u5_prod1_reg_36_ ( .D(u5_N36), .CK(clk), .Q(u5_prod1[36]) );
  DFF_X1 u5_prod1_reg_43_ ( .D(u5_N43), .CK(clk), .Q(u5_prod1[43]) );
  DFF_X1 u5_prod1_reg_44_ ( .D(u5_N44), .CK(clk), .Q(u5_prod1[44]) );
  DFF_X1 u5_prod1_reg_45_ ( .D(u5_N45), .CK(clk), .Q(u5_prod1[45]) );
  DFF_X2 opb_r_reg_22_ ( .D(opb[22]), .CK(clk), .Q(u6_N22), .QN(n3002) );
  DFF_X1 u5_prod1_reg_37_ ( .D(u5_N37), .CK(clk), .Q(u5_prod1[37]) );
  DFF_X1 u5_prod1_reg_35_ ( .D(u5_N35), .CK(clk), .Q(u5_prod1[35]) );
  DFF_X1 zero_reg ( .D(N531), .CK(clk), .Q(zero) );
  DFF_X1 out_reg_31_ ( .D(N495), .CK(clk), .Q(out[31]) );
  DFF_X1 u6_quo_reg_49_ ( .D(u6_quo1[49]), .CK(clk), .Q(quo[49]) );
  DFF_X1 inf_reg ( .D(N526), .CK(clk), .Q(inf) );
  DFF_X1 u5_prod1_reg_47_ ( .D(u5_N47), .CK(clk), .Q(u5_prod1[47]) );
  DFF_X1 u5_prod1_reg_30_ ( .D(u5_N30), .CK(clk), .Q(u5_prod1[30]) );
  DFF_X1 overflow_reg ( .D(N519), .CK(clk), .Q(overflow) );
  DFF_X2 opb_r_reg_11_ ( .D(opb[11]), .CK(clk), .QN(n2772) );
  DFF_X2 opb_r_reg_12_ ( .D(opb[12]), .CK(clk), .QN(n2771) );
  DFF_X2 opb_r_reg_14_ ( .D(opb[14]), .CK(clk), .Q(n2672), .QN(n2770) );
  DFF_X1 out_reg_28_ ( .D(N473), .CK(clk), .Q(out[28]) );
  DFF_X1 u5_prod1_reg_20_ ( .D(u5_N20), .CK(clk), .Q(u5_prod1[20]) );
  DFF_X1 u2_exp_out_reg_6_ ( .D(u2_N64), .CK(clk), .Q(exp_mul[6]), .QN(n2761)
         );
  DFF_X1 u2_exp_out_reg_2_ ( .D(u2_N60), .CK(clk), .Q(exp_mul[2]), .QN(n2760)
         );
  DFF_X1 u2_exp_out_reg_7_ ( .D(u2_N65), .CK(clk), .Q(exp_mul[7]), .QN(n2759)
         );
  DFF_X1 u2_exp_out_reg_3_ ( .D(u2_N61), .CK(clk), .Q(exp_mul[3]), .QN(n2758)
         );
  DFF_X1 u2_exp_out_reg_5_ ( .D(u2_N63), .CK(clk), .Q(exp_mul[5]), .QN(n2757)
         );
  DFF_X1 u2_exp_out_reg_1_ ( .D(u2_N59), .CK(clk), .Q(exp_mul[1]), .QN(n2756)
         );
  DFF_X1 u2_exp_out_reg_4_ ( .D(u2_N62), .CK(clk), .Q(exp_mul[4]), .QN(n2755)
         );
  DFF_X1 u2_exp_out_reg_0_ ( .D(u2_N58), .CK(clk), .Q(exp_mul[0]), .QN(n2754)
         );
  DFF_X1 u5_prod_reg_47_ ( .D(u5_prod1[47]), .CK(clk), .Q(prod[47]), .QN(n2730) );
  DFF_X1 u5_prod_reg_31_ ( .D(u5_prod1[31]), .CK(clk), .Q(prod[31]), .QN(n2717) );
  DFF_X1 u5_prod_reg_34_ ( .D(u5_prod1[34]), .CK(clk), .Q(prod[34]), .QN(n2713) );
  DFF_X1 u5_prod_reg_22_ ( .D(u5_prod1[22]), .CK(clk), .Q(prod[22]), .QN(n2712) );
  DFF_X2 u6_quo_reg_23_ ( .D(u6_quo1[23]), .CK(clk), .QN(n3026) );
  DFF_X1 u1_sign_reg ( .D(u1_sign_d), .CK(clk), .Q(sign_fasu), .QN(n2608) );
  DFF_X1 u5_prod_reg_32_ ( .D(u5_prod1[32]), .CK(clk), .Q(prod[32]), .QN(n2602) );
  DFF_X1 u5_prod_reg_35_ ( .D(u5_prod1[35]), .CK(clk), .Q(prod[35]), .QN(n2601) );
  DFF_X2 opb_r_reg_21_ ( .D(opb[21]), .CK(clk), .QN(n2693) );
  DFF_X2 opb_r_reg_19_ ( .D(opb[19]), .CK(clk), .QN(n2679) );
  DFF_X2 opb_r_reg_16_ ( .D(opb[16]), .CK(clk), .QN(n2680) );
  DFF_X2 opb_r_reg_20_ ( .D(opb[20]), .CK(clk), .QN(n2682) );
  DFF_X1 u5_prod_reg_33_ ( .D(u5_prod1[33]), .CK(clk), .Q(prod[33]), .QN(n2569) );
  DFF_X1 u5_prod_reg_25_ ( .D(u5_prod1[25]), .CK(clk), .Q(prod[25]), .QN(n2568) );
  DFF_X1 u5_prod1_reg_25_ ( .D(u5_N25), .CK(clk), .Q(u5_prod1[25]) );
  DFF_X1 out_reg_27_ ( .D(n2518), .CK(clk), .Q(out[27]) );
  DFF_X1 u5_prod1_reg_21_ ( .D(u5_N21), .CK(clk), .Q(u5_prod1[21]) );
  DFF_X1 u5_prod1_reg_19_ ( .D(u5_N19), .CK(clk), .Q(u5_prod1[19]) );
  NAND2_X2 U1933 ( .A1(n2810), .A2(net86234), .ZN(net84548) );
  AOI22_X4 U1934 ( .A1(1'b0), .A2(net85133), .B1(prod[23]), .B2(n2936), .ZN(
        n3170) );
  INV_X4 U1935 ( .A(n3234), .ZN(n3235) );
  INV_X4 U1936 ( .A(n3201), .ZN(n3202) );
  INV_X4 U1937 ( .A(remainder[26]), .ZN(n3637) );
  NOR2_X4 U1938 ( .A1(remainder[23]), .A2(remainder[22]), .ZN(n3617) );
  INV_X2 U1939 ( .A(n4076), .ZN(n2460) );
  INV_X4 U1940 ( .A(n4076), .ZN(n3918) );
  NAND2_X2 U1941 ( .A1(net83415), .A2(net92622), .ZN(n2990) );
  BUF_X16 U1942 ( .A(n2892), .Z(n2461) );
  AOI211_X2 U1943 ( .C1(n4099), .C2(net85989), .A(net82757), .B(net85976), 
        .ZN(N461) );
  BUF_X16 U1944 ( .A(n2998), .Z(n2462) );
  INV_X4 U1945 ( .A(n2467), .ZN(n2463) );
  INV_X4 U1946 ( .A(net92626), .ZN(n2467) );
  NAND2_X2 U1947 ( .A1(n3843), .A2(n3054), .ZN(n2464) );
  INV_X8 U1948 ( .A(n4034), .ZN(n2997) );
  NAND3_X2 U1949 ( .A1(n3753), .A2(n3752), .A3(n3751), .ZN(n2465) );
  INV_X8 U1950 ( .A(n3796), .ZN(n3800) );
  OAI22_X4 U1951 ( .A1(n3057), .A2(n2658), .B1(net83326), .B2(net83327), .ZN(
        n3803) );
  INV_X2 U1952 ( .A(net95614), .ZN(net82891) );
  NAND2_X1 U1953 ( .A1(net83297), .A2(n3844), .ZN(net82957) );
  INV_X8 U1954 ( .A(n4108), .ZN(n3919) );
  OAI22_X4 U1955 ( .A1(net86014), .A2(n2624), .B1(net86001), .B2(n3867), .ZN(
        n4108) );
  AND3_X2 U1956 ( .A1(n4044), .A2(net91733), .A3(net82876), .ZN(n4057) );
  NAND2_X1 U1957 ( .A1(n3917), .A2(n3921), .ZN(n2466) );
  NAND2_X4 U1958 ( .A1(net86497), .A2(n2992), .ZN(n3873) );
  INV_X2 U1959 ( .A(n3054), .ZN(n4074) );
  NOR3_X2 U1960 ( .A1(n4039), .A2(n4074), .A3(n4038), .ZN(n4040) );
  INV_X4 U1961 ( .A(n4095), .ZN(n2549) );
  INV_X4 U1962 ( .A(n4107), .ZN(n3868) );
  NAND4_X4 U1963 ( .A1(net83119), .A2(net83120), .A3(net83117), .A4(net95549), 
        .ZN(n2475) );
  INV_X4 U1964 ( .A(n2478), .ZN(n3920) );
  INV_X8 U1965 ( .A(n4098), .ZN(n4024) );
  INV_X1 U1966 ( .A(net95549), .ZN(net94976) );
  NAND2_X2 U1967 ( .A1(n3895), .A2(u4_fract_out_21_), .ZN(n3865) );
  INV_X1 U1968 ( .A(net83441), .ZN(n2468) );
  INV_X2 U1969 ( .A(n3741), .ZN(n3742) );
  CLKBUF_X3 U1970 ( .A(u4_div_exp2_7_), .Z(net93036) );
  INV_X16 U1971 ( .A(net23043), .ZN(n2469) );
  INV_X16 U1972 ( .A(net83754), .ZN(net23043) );
  INV_X1 U1973 ( .A(n2924), .ZN(n2970) );
  NOR2_X2 U1974 ( .A1(n3495), .A2(net95173), .ZN(n3477) );
  NAND2_X2 U1975 ( .A1(div_opa_ldz_r2[2]), .A2(net83754), .ZN(net84132) );
  OAI211_X2 U1976 ( .C1(net94513), .C2(net86028), .A(net83991), .B(n2795), 
        .ZN(u4_exp_out_3_) );
  INV_X2 U1977 ( .A(net94513), .ZN(net83018) );
  OR2_X2 U1978 ( .A1(n3473), .A2(net94004), .ZN(n2470) );
  NAND2_X2 U1979 ( .A1(n3394), .A2(net91297), .ZN(n3405) );
  CLKBUF_X2 U1980 ( .A(n3431), .Z(n2471) );
  INV_X4 U1981 ( .A(n3207), .ZN(n2472) );
  INV_X4 U1982 ( .A(n2472), .ZN(n2473) );
  AOI22_X4 U1983 ( .A1(fract_i2f[33]), .A2(net85115), .B1(prod[33]), .B2(n2936), .ZN(n3207) );
  BUF_X8 U1984 ( .A(n3612), .Z(n2474) );
  NAND2_X4 U1985 ( .A1(n2513), .A2(n3672), .ZN(n3675) );
  NAND3_X2 U1986 ( .A1(n3672), .A2(n2901), .A3(n3671), .ZN(n3673) );
  NAND4_X4 U1987 ( .A1(quo[38]), .A2(net85175), .A3(net85159), .A4(net85135), 
        .ZN(n3251) );
  NAND2_X2 U1988 ( .A1(n4118), .A2(n4121), .ZN(n3927) );
  NOR2_X4 U1989 ( .A1(n4063), .A2(net85976), .ZN(n4068) );
  OAI21_X4 U1990 ( .B1(n3655), .B2(n3656), .A(n2794), .ZN(n3672) );
  NOR2_X2 U1991 ( .A1(n2485), .A2(n2505), .ZN(n2780) );
  INV_X4 U1992 ( .A(net82902), .ZN(net82781) );
  INV_X4 U1993 ( .A(n4100), .ZN(n4026) );
  NAND2_X4 U1994 ( .A1(net83057), .A2(n2834), .ZN(n2833) );
  BUF_X32 U1995 ( .A(u4_exp_out_6_), .Z(n2476) );
  OAI21_X4 U1996 ( .B1(n3655), .B2(n3656), .A(n2794), .ZN(n2477) );
  NAND4_X4 U1997 ( .A1(n3654), .A2(n3653), .A3(n3652), .A4(n3651), .ZN(n3655)
         );
  OAI22_X4 U1998 ( .A1(net85999), .A2(n3888), .B1(n3887), .B2(net86015), .ZN(
        n2478) );
  OAI22_X2 U1999 ( .A1(net85999), .A2(n3888), .B1(n3887), .B2(net86015), .ZN(
        n4095) );
  INV_X1 U2000 ( .A(n4028), .ZN(n2479) );
  INV_X8 U2001 ( .A(n4103), .ZN(n4028) );
  NAND3_X4 U2002 ( .A1(n3843), .A2(net82826), .A3(net85986), .ZN(n4039) );
  CLKBUF_X2 U2003 ( .A(u4_fract_out_9_), .Z(n2480) );
  INV_X2 U2004 ( .A(fract_denorm[37]), .ZN(net84355) );
  BUF_X32 U2005 ( .A(n2975), .Z(n2481) );
  INV_X1 U2006 ( .A(fract_denorm[34]), .ZN(n2482) );
  NAND3_X4 U2007 ( .A1(n3255), .A2(n3257), .A3(n3256), .ZN(n2483) );
  NAND3_X2 U2008 ( .A1(n3255), .A2(n3257), .A3(n3256), .ZN(fract_denorm[35])
         );
  NAND3_X2 U2009 ( .A1(n3728), .A2(n3727), .A3(n3726), .ZN(n3729) );
  NOR2_X1 U2010 ( .A1(n2505), .A2(n1452), .ZN(n3056) );
  NAND2_X2 U2011 ( .A1(net86497), .A2(u4_fract_out_18_), .ZN(n3863) );
  BUF_X32 U2012 ( .A(net82953), .Z(n2484) );
  NOR2_X1 U2013 ( .A1(net83126), .A2(n3883), .ZN(n3884) );
  NOR2_X1 U2014 ( .A1(net83126), .A2(n3841), .ZN(n3842) );
  NAND2_X1 U2015 ( .A1(net86497), .A2(u4_fract_out_19_), .ZN(n3861) );
  INV_X1 U2016 ( .A(n1457), .ZN(u4_fract_out_18_) );
  NAND2_X4 U2017 ( .A1(n1457), .A2(n1459), .ZN(n2491) );
  INV_X2 U2018 ( .A(n1450), .ZN(u4_fract_out_9_) );
  INV_X1 U2019 ( .A(u4_fract_out_15_), .ZN(n2485) );
  INV_X2 U2020 ( .A(n2058), .ZN(u4_fract_out_21_) );
  NAND2_X2 U2021 ( .A1(net84132), .A2(n2488), .ZN(n2875) );
  NAND3_X2 U2022 ( .A1(net84171), .A2(net84349), .A3(net84350), .ZN(net84293)
         );
  INV_X1 U2023 ( .A(net23043), .ZN(net95431) );
  AOI21_X2 U2024 ( .B1(net93422), .B2(net84382), .A(n3344), .ZN(n3368) );
  OR2_X2 U2025 ( .A1(n3502), .A2(n2906), .ZN(net94516) );
  INV_X8 U2026 ( .A(u4_div_exp2_6_), .ZN(net83767) );
  NAND2_X2 U2027 ( .A1(n2486), .A2(n2487), .ZN(n2488) );
  INV_X1 U2028 ( .A(div_opa_ldz_r2[2]), .ZN(n2486) );
  INV_X4 U2029 ( .A(net83754), .ZN(n2487) );
  INV_X8 U2030 ( .A(net93776), .ZN(net93777) );
  INV_X4 U2031 ( .A(net84270), .ZN(n2489) );
  INV_X4 U2032 ( .A(n2489), .ZN(n2490) );
  NOR2_X4 U2033 ( .A1(net84271), .A2(net94138), .ZN(net84270) );
  NOR2_X2 U2034 ( .A1(net83771), .A2(net95136), .ZN(net83770) );
  BUF_X32 U2035 ( .A(n4001), .Z(n2903) );
  NAND2_X2 U2036 ( .A1(net83446), .A2(n2662), .ZN(net83416) );
  NOR3_X2 U2037 ( .A1(n3411), .A2(n3410), .A3(n3409), .ZN(net84204) );
  NAND2_X2 U2038 ( .A1(n2492), .A2(n2093), .ZN(n3603) );
  INV_X4 U2039 ( .A(n2491), .ZN(n2492) );
  NOR2_X2 U2040 ( .A1(net85111), .A2(n2634), .ZN(n2493) );
  NOR2_X2 U2041 ( .A1(net92028), .A2(n2494), .ZN(n3253) );
  INV_X4 U2042 ( .A(n2493), .ZN(n2494) );
  BUF_X32 U2043 ( .A(net83020), .Z(n2495) );
  NAND2_X4 U2044 ( .A1(n2666), .A2(n3395), .ZN(net84238) );
  INV_X4 U2045 ( .A(net83931), .ZN(net83930) );
  INV_X8 U2046 ( .A(net84121), .ZN(net84128) );
  INV_X8 U2047 ( .A(net83864), .ZN(n2791) );
  NAND3_X4 U2048 ( .A1(n3242), .A2(n3241), .A3(n3240), .ZN(fract_denorm[42])
         );
  NAND3_X2 U2049 ( .A1(n3242), .A2(n3241), .A3(n3240), .ZN(net94305) );
  NAND2_X4 U2050 ( .A1(n3601), .A2(n3600), .ZN(net83738) );
  NAND2_X2 U2051 ( .A1(n3471), .A2(n2496), .ZN(n2497) );
  NAND2_X1 U2052 ( .A1(n3472), .A2(net93695), .ZN(n2498) );
  NAND2_X2 U2053 ( .A1(n2497), .A2(n2498), .ZN(n3476) );
  INV_X1 U2054 ( .A(net93695), .ZN(n2496) );
  INV_X1 U2055 ( .A(u4_fi_ldz_mi1_1_), .ZN(n2499) );
  INV_X2 U2056 ( .A(n2499), .ZN(n2500) );
  INV_X2 U2057 ( .A(u4_exp_in_pl1_5_), .ZN(n3472) );
  INV_X16 U2058 ( .A(net85393), .ZN(net93695) );
  OAI221_X4 U2059 ( .B1(net83766), .B2(net83750), .C1(net83767), .C2(net95102), 
        .A(n3590), .ZN(n3955) );
  INV_X4 U2060 ( .A(u4_exp_next_mi_5_), .ZN(n3471) );
  NAND2_X2 U2061 ( .A1(n4069), .A2(net85121), .ZN(n4073) );
  NAND3_X1 U2062 ( .A1(n3895), .A2(net86013), .A3(u4_fract_out_pl1_5_), .ZN(
        n3857) );
  NAND2_X4 U2063 ( .A1(n2558), .A2(n2559), .ZN(n3752) );
  NAND2_X2 U2064 ( .A1(net83518), .A2(rmode_r3[1]), .ZN(n2502) );
  BUF_X8 U2065 ( .A(net83499), .Z(n2501) );
  AOI211_X2 U2066 ( .C1(n4096), .C2(net85988), .A(net82757), .B(net85976), 
        .ZN(N459) );
  INV_X4 U2067 ( .A(n1452), .ZN(u4_fract_out_7_) );
  NAND2_X2 U2068 ( .A1(sign), .A2(net82853), .ZN(n2503) );
  NAND2_X1 U2069 ( .A1(n2504), .A2(net95525), .ZN(net82850) );
  INV_X4 U2070 ( .A(n2503), .ZN(n2504) );
  NAND2_X1 U2071 ( .A1(n2463), .A2(net83422), .ZN(net83418) );
  INV_X8 U2072 ( .A(net86481), .ZN(n2505) );
  INV_X4 U2073 ( .A(net86481), .ZN(net86496) );
  INV_X4 U2074 ( .A(net83279), .ZN(net83274) );
  AND2_X2 U2075 ( .A1(n3796), .A2(n3821), .ZN(n2525) );
  NAND4_X2 U2076 ( .A1(net83842), .A2(n3579), .A3(n3580), .A4(n3578), .ZN(
        u4_shift_left[1]) );
  INV_X4 U2077 ( .A(n2779), .ZN(n2964) );
  INV_X8 U2078 ( .A(n3999), .ZN(n3684) );
  NOR2_X4 U2079 ( .A1(n3731), .A2(n3825), .ZN(n3754) );
  NAND2_X1 U2080 ( .A1(n3825), .A2(net83271), .ZN(n3826) );
  INV_X8 U2081 ( .A(n1453), .ZN(u4_fract_out_3_) );
  NOR2_X2 U2082 ( .A1(n2906), .A2(n2926), .ZN(n3494) );
  INV_X2 U2083 ( .A(n2470), .ZN(n2906) );
  NOR2_X1 U2084 ( .A1(net83474), .A2(net85901), .ZN(n2506) );
  NOR2_X4 U2085 ( .A1(u4_N1733), .A2(n2507), .ZN(net82998) );
  INV_X4 U2086 ( .A(n2506), .ZN(n2507) );
  INV_X8 U2087 ( .A(net84324), .ZN(net94138) );
  NAND3_X1 U2088 ( .A1(n3210), .A2(n3211), .A3(n3212), .ZN(n2552) );
  INV_X8 U2089 ( .A(n2747), .ZN(net85901) );
  CLKBUF_X3 U2090 ( .A(net82998), .Z(net94933) );
  INV_X8 U2091 ( .A(u4_div_exp2_4_), .ZN(net84017) );
  NAND2_X4 U2092 ( .A1(n2861), .A2(net95353), .ZN(n2866) );
  NAND3_X2 U2093 ( .A1(net17694), .A2(net84280), .A3(n2557), .ZN(n2861) );
  NOR2_X4 U2094 ( .A1(net85143), .A2(n2556), .ZN(n3246) );
  INV_X8 U2095 ( .A(n2555), .ZN(n2556) );
  INV_X8 U2096 ( .A(n3475), .ZN(n2976) );
  NAND2_X4 U2097 ( .A1(n1450), .A2(n1452), .ZN(net83731) );
  NAND2_X2 U2098 ( .A1(n3737), .A2(n2508), .ZN(n2509) );
  NAND2_X1 U2099 ( .A1(n3808), .A2(net83507), .ZN(n2510) );
  NAND2_X2 U2100 ( .A1(n2509), .A2(n2510), .ZN(n3738) );
  INV_X1 U2101 ( .A(net83507), .ZN(n2508) );
  INV_X2 U2102 ( .A(net83526), .ZN(n2511) );
  NAND2_X1 U2103 ( .A1(net86028), .A2(n3659), .ZN(n2512) );
  INV_X4 U2104 ( .A(n2512), .ZN(n2513) );
  INV_X1 U2105 ( .A(n3736), .ZN(n3737) );
  INV_X4 U2106 ( .A(u4_exp_out_1_), .ZN(net83507) );
  NAND3_X2 U2107 ( .A1(n3738), .A2(n3739), .A3(n2972), .ZN(n3828) );
  INV_X16 U2108 ( .A(net86027), .ZN(net86028) );
  BUF_X4 U2109 ( .A(n2278), .Z(n2901) );
  BUF_X32 U2110 ( .A(u4_fract_out_10_), .Z(n2514) );
  INV_X8 U2111 ( .A(n4553), .ZN(n5290) );
  INV_X16 U2112 ( .A(n4726), .ZN(n3079) );
  INV_X2 U2113 ( .A(opb_r[24]), .ZN(n4473) );
  NAND2_X1 U2114 ( .A1(opb_r[24]), .A2(opb_r[23]), .ZN(n4738) );
  NAND2_X2 U2115 ( .A1(n4121), .A2(n2519), .ZN(n2518) );
  INV_X32 U2116 ( .A(net82757), .ZN(n2519) );
  NAND2_X2 U2117 ( .A1(n3950), .A2(n2521), .ZN(n2520) );
  INV_X32 U2118 ( .A(net82757), .ZN(n2521) );
  INV_X2 U2119 ( .A(n2589), .ZN(n2523) );
  AOI211_X4 U2120 ( .C1(n4093), .C2(net85989), .A(net82757), .B(net85976), 
        .ZN(N457) );
  AOI211_X4 U2121 ( .C1(net82792), .C2(net85990), .A(net82757), .B(net85976), 
        .ZN(N462) );
  AOI211_X4 U2122 ( .C1(n4102), .C2(net85989), .A(net82757), .B(net85976), 
        .ZN(N463) );
  AOI211_X4 U2123 ( .C1(n4104), .C2(net85989), .A(net82757), .B(net85976), 
        .ZN(N464) );
  AOI211_X4 U2124 ( .C1(n4106), .C2(net85989), .A(net82757), .B(net85976), 
        .ZN(N465) );
  AOI211_X4 U2125 ( .C1(net82784), .C2(net85990), .A(net82757), .B(net85976), 
        .ZN(N466) );
  AOI211_X4 U2126 ( .C1(n4086), .C2(net85988), .A(net82757), .B(net85976), 
        .ZN(N452) );
  AOI211_X4 U2127 ( .C1(n4092), .C2(net85988), .A(net82757), .B(net85976), 
        .ZN(N456) );
  AOI211_X4 U2128 ( .C1(n4094), .C2(net85988), .A(net82757), .B(net85976), 
        .ZN(N458) );
  AOI211_X4 U2129 ( .C1(n4077), .C2(net85987), .A(net82757), .B(net85976), 
        .ZN(N447) );
  AOI211_X4 U2130 ( .C1(n4088), .C2(net85987), .A(net82757), .B(net85976), 
        .ZN(N453) );
  AOI211_X4 U2131 ( .C1(n4090), .C2(net85987), .A(net82757), .B(net85976), 
        .ZN(N454) );
  AOI211_X4 U2132 ( .C1(n4091), .C2(net85987), .A(net82757), .B(net85976), 
        .ZN(N455) );
  AOI211_X4 U2133 ( .C1(n4075), .C2(net85986), .A(net82757), .B(net85976), 
        .ZN(N446) );
  AOI211_X4 U2134 ( .C1(n4079), .C2(net85986), .A(net82757), .B(net85976), 
        .ZN(N448) );
  AOI211_X4 U2135 ( .C1(n4081), .C2(net85986), .A(net82757), .B(net85976), 
        .ZN(N449) );
  AOI211_X4 U2136 ( .C1(n4083), .C2(net85986), .A(net82757), .B(net85976), 
        .ZN(N450) );
  NOR3_X4 U2137 ( .A1(n3800), .A2(n2524), .A3(n3799), .ZN(n3057) );
  INV_X32 U2138 ( .A(n3802), .ZN(n2524) );
  OAI21_X2 U2139 ( .B1(net82931), .B2(n3793), .A(n3790), .ZN(n3799) );
  INV_X2 U2140 ( .A(n3919), .ZN(n2893) );
  NAND2_X4 U2141 ( .A1(n4007), .A2(n3817), .ZN(net83349) );
  INV_X2 U2142 ( .A(n2693), .ZN(n2526) );
  INV_X2 U2143 ( .A(n4122), .ZN(n3846) );
  NAND2_X2 U2144 ( .A1(net82753), .A2(n4122), .ZN(N468) );
  OAI21_X2 U2145 ( .B1(n4023), .B2(n4113), .A(n4022), .ZN(N509) );
  OAI211_X2 U2146 ( .C1(n4068), .C2(n2911), .A(n4066), .B(n4065), .ZN(n4069)
         );
  INV_X8 U2147 ( .A(net85163), .ZN(net85157) );
  INV_X2 U2148 ( .A(net84385), .ZN(net92690) );
  NAND2_X4 U2149 ( .A1(n2842), .A2(net83278), .ZN(net86481) );
  NOR2_X2 U2150 ( .A1(n3229), .A2(net85175), .ZN(n3209) );
  AND3_X4 U2151 ( .A1(prod[41]), .A2(net85133), .A3(net85165), .ZN(n2527) );
  NOR2_X2 U2152 ( .A1(net94019), .A2(net85163), .ZN(net86295) );
  AND2_X2 U2153 ( .A1(n4753), .A2(n4752), .ZN(n2528) );
  AND2_X2 U2154 ( .A1(n4753), .A2(n3514), .ZN(n2529) );
  INV_X8 U2155 ( .A(net26607), .ZN(net85399) );
  OR2_X1 U2156 ( .A1(net86571), .A2(fract_denorm[45]), .ZN(n2530) );
  NOR2_X4 U2157 ( .A1(net85157), .A2(net85143), .ZN(n3238) );
  INV_X16 U2158 ( .A(fract_denorm[28]), .ZN(n3021) );
  NOR2_X4 U2159 ( .A1(net85145), .A2(net85157), .ZN(n3174) );
  INV_X8 U2160 ( .A(net92573), .ZN(net84321) );
  AND2_X2 U2161 ( .A1(net83744), .A2(net94614), .ZN(n2531) );
  INV_X8 U2162 ( .A(net84298), .ZN(net84377) );
  OR2_X1 U2163 ( .A1(net83660), .A2(net83041), .ZN(n2532) );
  INV_X8 U2164 ( .A(net94566), .ZN(net83487) );
  INV_X8 U2165 ( .A(net83796), .ZN(net23182) );
  NAND2_X4 U2166 ( .A1(net83797), .A2(n2670), .ZN(net83796) );
  AND2_X4 U2167 ( .A1(net83854), .A2(n3573), .ZN(n2533) );
  OR2_X1 U2168 ( .A1(n2745), .A2(net94725), .ZN(n2534) );
  INV_X2 U2169 ( .A(net83282), .ZN(net83271) );
  AOI21_X2 U2170 ( .B1(n3822), .B2(n3821), .A(n3824), .ZN(net83282) );
  INV_X4 U2171 ( .A(n3677), .ZN(n3998) );
  NAND2_X4 U2172 ( .A1(n3674), .A2(n3673), .ZN(net83565) );
  INV_X4 U2173 ( .A(u4_fract_out_22_), .ZN(n3016) );
  AND2_X2 U2174 ( .A1(net86497), .A2(u4_fract_out_5_), .ZN(n2535) );
  NAND2_X4 U2175 ( .A1(net94703), .A2(net83278), .ZN(n3895) );
  INV_X8 U2176 ( .A(net85997), .ZN(net85998) );
  INV_X16 U2177 ( .A(net86013), .ZN(net86015) );
  OR2_X2 U2178 ( .A1(n3733), .A2(net83514), .ZN(n2536) );
  AOI22_X4 U2179 ( .A1(net92566), .A2(n3884), .B1(n3056), .B2(net85997), .ZN(
        n2898) );
  OR2_X2 U2180 ( .A1(net83126), .A2(n3864), .ZN(n2537) );
  OR2_X2 U2181 ( .A1(net83126), .A2(n3860), .ZN(n2538) );
  OAI22_X4 U2182 ( .A1(net92365), .A2(net86015), .B1(net85998), .B2(net83166), 
        .ZN(net95614) );
  BUF_X16 U2183 ( .A(n1454), .Z(n2952) );
  NOR2_X1 U2184 ( .A1(n3715), .A2(n3714), .ZN(n3716) );
  AOI21_X4 U2185 ( .B1(n3608), .B2(n3430), .A(n3429), .ZN(n3433) );
  NAND2_X4 U2186 ( .A1(u4_N1455), .A2(n2794), .ZN(n2539) );
  BUF_X8 U2187 ( .A(net84356), .Z(n2540) );
  NAND2_X2 U2188 ( .A1(n3895), .A2(u4_fract_out_4_), .ZN(n3852) );
  OAI21_X4 U2189 ( .B1(net83562), .B2(net83563), .A(net83234), .ZN(net83498)
         );
  NAND2_X2 U2190 ( .A1(n3732), .A2(n2541), .ZN(n2542) );
  NAND2_X1 U2191 ( .A1(net83368), .A2(net83518), .ZN(n2543) );
  NAND2_X2 U2192 ( .A1(n2542), .A2(n2543), .ZN(n3733) );
  INV_X1 U2193 ( .A(net83518), .ZN(n2541) );
  NAND2_X2 U2194 ( .A1(net85997), .A2(n2535), .ZN(n2544) );
  NAND2_X4 U2195 ( .A1(n2544), .A2(n3857), .ZN(n4082) );
  NAND2_X1 U2196 ( .A1(u4_exp_out_pl1_0_), .A2(net82040), .ZN(n3732) );
  INV_X1 U2197 ( .A(net48876), .ZN(net83368) );
  NAND4_X4 U2198 ( .A1(n3754), .A2(net83329), .A3(n3828), .A4(n2536), .ZN(
        n2910) );
  AOI21_X2 U2199 ( .B1(net83807), .B2(net83808), .A(net86032), .ZN(net83800)
         );
  INV_X4 U2200 ( .A(net84257), .ZN(net84341) );
  INV_X1 U2201 ( .A(fract_denorm[27]), .ZN(n2545) );
  INV_X2 U2202 ( .A(n2545), .ZN(n2546) );
  AOI22_X2 U2203 ( .A1(net84556), .A2(fract_out_q[26]), .B1(fract_i2f[46]), 
        .B2(net90945), .ZN(net84546) );
  INV_X1 U2204 ( .A(n3021), .ZN(n2547) );
  NOR3_X2 U2205 ( .A1(n3043), .A2(net92028), .A3(net90945), .ZN(n3214) );
  NAND2_X2 U2206 ( .A1(n3895), .A2(u4_fract_out_13_), .ZN(n2912) );
  AOI22_X4 U2207 ( .A1(n3174), .A2(prod[37]), .B1(fract_i2f[37]), .B2(net85115), .ZN(n3270) );
  NAND2_X2 U2208 ( .A1(n2549), .A2(n2779), .ZN(n2896) );
  INV_X4 U2209 ( .A(n3606), .ZN(n3024) );
  NOR3_X4 U2210 ( .A1(n2627), .A2(net92028), .A3(net85111), .ZN(n3243) );
  INV_X4 U2211 ( .A(net85119), .ZN(net85117) );
  INV_X4 U2212 ( .A(net83445), .ZN(net83444) );
  INV_X8 U2213 ( .A(n4024), .ZN(n2892) );
  OR2_X4 U2214 ( .A1(n5324), .A2(n5325), .ZN(n2548) );
  NAND3_X2 U2215 ( .A1(n3169), .A2(n3170), .A3(n3168), .ZN(n3068) );
  INV_X4 U2216 ( .A(n2964), .ZN(n2958) );
  CLKBUF_X3 U2217 ( .A(net83771), .Z(n2561) );
  NAND4_X1 U2218 ( .A1(n4035), .A2(net95549), .A3(n3917), .A4(net86418), .ZN(
        n3925) );
  INV_X1 U2219 ( .A(n3917), .ZN(n2895) );
  INV_X8 U2220 ( .A(net83811), .ZN(net83854) );
  NAND2_X4 U2221 ( .A1(n3541), .A2(net86045), .ZN(net83811) );
  INV_X8 U2222 ( .A(n3532), .ZN(n3541) );
  NOR3_X4 U2223 ( .A1(u4_N1431), .A2(u4_N1430), .A3(u4_N1429), .ZN(n3654) );
  INV_X2 U2224 ( .A(n1459), .ZN(u4_fract_out_13_) );
  INV_X2 U2225 ( .A(u4_fract_out_pl1_22_), .ZN(n3866) );
  BUF_X32 U2226 ( .A(u4_fract_out_20_), .Z(n2550) );
  INV_X32 U2227 ( .A(net86013), .ZN(net86014) );
  NAND3_X1 U2228 ( .A1(n2536), .A2(net83305), .A3(n3812), .ZN(n3813) );
  INV_X8 U2229 ( .A(n2060), .ZN(u4_fract_out_20_) );
  NAND2_X4 U2230 ( .A1(net83036), .A2(n3688), .ZN(n3715) );
  OAI22_X4 U2231 ( .A1(net86001), .A2(n3882), .B1(net86014), .B2(net86478), 
        .ZN(n4089) );
  NAND2_X4 U2232 ( .A1(quo[26]), .A2(net92028), .ZN(n3158) );
  INV_X4 U2233 ( .A(fract_denorm[24]), .ZN(n3334) );
  NAND2_X2 U2234 ( .A1(net83715), .A2(net84324), .ZN(n3391) );
  INV_X8 U2235 ( .A(net86257), .ZN(net85125) );
  INV_X16 U2236 ( .A(net85125), .ZN(net85121) );
  NAND2_X2 U2237 ( .A1(net85139), .A2(net85159), .ZN(n3229) );
  NAND3_X2 U2238 ( .A1(n3210), .A2(n3211), .A3(n3212), .ZN(n2551) );
  NAND3_X2 U2239 ( .A1(n3210), .A2(n3211), .A3(n3212), .ZN(fract_denorm[39])
         );
  INV_X1 U2240 ( .A(n2481), .ZN(n2553) );
  INV_X2 U2241 ( .A(n2553), .ZN(n2554) );
  NOR2_X4 U2242 ( .A1(net85157), .A2(n2625), .ZN(n2555) );
  XNOR2_X1 U2243 ( .A(n3027), .B(net85933), .ZN(n3585) );
  NOR2_X2 U2244 ( .A1(n3045), .A2(net85121), .ZN(n3044) );
  NOR2_X4 U2245 ( .A1(n3371), .A2(n3370), .ZN(n3407) );
  INV_X1 U2246 ( .A(fract_denorm[36]), .ZN(net84351) );
  NOR2_X4 U2247 ( .A1(net33106), .A2(n2654), .ZN(n2877) );
  INV_X4 U2248 ( .A(net84281), .ZN(n2557) );
  INV_X8 U2249 ( .A(net84281), .ZN(net84201) );
  NAND2_X2 U2250 ( .A1(n3747), .A2(net94566), .ZN(n2558) );
  NAND2_X1 U2251 ( .A1(n3746), .A2(net83487), .ZN(n2559) );
  NOR2_X4 U2252 ( .A1(net93714), .A2(n2532), .ZN(n3644) );
  NAND3_X2 U2253 ( .A1(n3753), .A2(n3752), .A3(n3751), .ZN(net83329) );
  AOI211_X2 U2254 ( .C1(n3743), .C2(n2621), .A(net83492), .B(n3742), .ZN(n3747) );
  AOI211_X2 U2255 ( .C1(net82036), .C2(n2674), .A(n3643), .B(n3763), .ZN(
        net83660) );
  AND2_X2 U2256 ( .A1(net95019), .A2(u4_fract_out_3_), .ZN(n2560) );
  NAND2_X2 U2257 ( .A1(n3895), .A2(n2480), .ZN(n3882) );
  INV_X16 U2258 ( .A(net85997), .ZN(net86001) );
  NAND2_X1 U2259 ( .A1(net48876), .A2(net83446), .ZN(n3718) );
  NAND3_X4 U2260 ( .A1(n4001), .A2(n3675), .A3(n2669), .ZN(n3661) );
  NAND2_X4 U2261 ( .A1(n4001), .A2(n3675), .ZN(n3999) );
  OAI21_X2 U2262 ( .B1(n3658), .B2(n3657), .A(net85377), .ZN(n3659) );
  NAND2_X2 U2263 ( .A1(n3736), .A2(u4_exp_out_2_), .ZN(n3719) );
  NAND2_X4 U2264 ( .A1(n3677), .A2(n3676), .ZN(net83563) );
  NAND2_X2 U2265 ( .A1(n3999), .A2(n2093), .ZN(n3676) );
  NOR2_X1 U2266 ( .A1(net82782), .A2(n4082), .ZN(n4083) );
  INV_X4 U2267 ( .A(n2087), .ZN(u4_fract_out_4_) );
  NOR2_X1 U2268 ( .A1(n3376), .A2(n3447), .ZN(n3377) );
  OR2_X1 U2269 ( .A1(n2552), .A2(fract_denorm[40]), .ZN(n2955) );
  NAND4_X4 U2270 ( .A1(quo[47]), .A2(net85175), .A3(net92028), .A4(net85159), 
        .ZN(n3236) );
  NAND2_X4 U2271 ( .A1(net83929), .A2(net83834), .ZN(n2790) );
  NAND2_X1 U2272 ( .A1(net84356), .A2(n2856), .ZN(n2562) );
  AOI22_X4 U2273 ( .A1(n3258), .A2(prod[45]), .B1(fract_i2f[45]), .B2(net85115), .ZN(n3237) );
  NOR2_X2 U2274 ( .A1(net85145), .A2(net85159), .ZN(n3258) );
  NOR3_X2 U2275 ( .A1(net93364), .A2(net85143), .A3(n3070), .ZN(n3069) );
  INV_X1 U2276 ( .A(n2540), .ZN(n2563) );
  INV_X16 U2277 ( .A(fract_denorm[43]), .ZN(net84180) );
  INV_X8 U2278 ( .A(net86014), .ZN(net92566) );
  NAND4_X4 U2279 ( .A1(net83723), .A2(net83724), .A3(net83725), .A4(net83726), 
        .ZN(net82953) );
  INV_X4 U2280 ( .A(net82038), .ZN(net83601) );
  NAND2_X1 U2281 ( .A1(sign_fasu_r), .A2(n2833), .ZN(n2989) );
  INV_X4 U2282 ( .A(net84312), .ZN(net84311) );
  INV_X4 U2283 ( .A(n3447), .ZN(n3355) );
  INV_X8 U2284 ( .A(fpu_op_r3_1_), .ZN(net90897) );
  NAND2_X2 U2285 ( .A1(net85135), .A2(net85159), .ZN(n3252) );
  NOR3_X2 U2286 ( .A1(n2633), .A2(net85111), .A3(net85135), .ZN(n3186) );
  NAND2_X1 U2287 ( .A1(net85135), .A2(net85121), .ZN(n3282) );
  AOI22_X2 U2288 ( .A1(n3199), .A2(fract_out_q[2]), .B1(fract_i2f[22]), .B2(
        net85115), .ZN(n3204) );
  NAND3_X4 U2289 ( .A1(quo[0]), .A2(net85133), .A3(n3284), .ZN(n3195) );
  AND4_X4 U2290 ( .A1(n3228), .A2(n3227), .A3(n3226), .A4(n3225), .ZN(n2564)
         );
  INV_X4 U2291 ( .A(n2564), .ZN(fract_denorm[32]) );
  NOR2_X2 U2292 ( .A1(n3252), .A2(net85175), .ZN(n3254) );
  INV_X1 U2293 ( .A(n3475), .ZN(n3495) );
  INV_X16 U2294 ( .A(net85169), .ZN(net85163) );
  INV_X8 U2295 ( .A(n2851), .ZN(n2856) );
  NAND2_X2 U2296 ( .A1(net85143), .A2(net85121), .ZN(n4109) );
  AOI22_X4 U2297 ( .A1(u4_exp_f2i_1[55]), .A2(n2652), .B1(n1373), .B2(net83776), .ZN(n3593) );
  INV_X8 U2298 ( .A(net86294), .ZN(net85169) );
  INV_X32 U2299 ( .A(net85163), .ZN(net85159) );
  NOR2_X2 U2300 ( .A1(n3477), .A2(n2561), .ZN(n3481) );
  NAND2_X4 U2301 ( .A1(n2791), .A2(div_opa_ldz_r2[0]), .ZN(n2788) );
  NOR3_X4 U2302 ( .A1(n3927), .A2(n3930), .A3(n4119), .ZN(n3847) );
  AND2_X2 U2303 ( .A1(net95019), .A2(u4_fract_out_3_), .ZN(n3052) );
  NOR4_X2 U2304 ( .A1(n3925), .A2(n3924), .A3(n3923), .A4(n3922), .ZN(net83057) );
  OAI21_X2 U2305 ( .B1(n3980), .B2(n3979), .A(n2534), .ZN(n3981) );
  AOI211_X2 U2306 ( .C1(net83417), .C2(net83418), .A(n2511), .B(net95504), 
        .ZN(net83415) );
  INV_X4 U2307 ( .A(net84003), .ZN(net94515) );
  INV_X4 U2308 ( .A(net84002), .ZN(net94514) );
  NAND4_X2 U2309 ( .A1(n4034), .A2(n4026), .A3(n3921), .A4(n4025), .ZN(n3922)
         );
  NOR2_X1 U2310 ( .A1(net85933), .A2(net84738), .ZN(n3134) );
  OAI21_X2 U2311 ( .B1(n3466), .B2(n4747), .A(net82029), .ZN(n3900) );
  INV_X4 U2312 ( .A(n2668), .ZN(net85937) );
  NOR2_X1 U2313 ( .A1(net83862), .A2(n3734), .ZN(net83858) );
  NOR2_X2 U2314 ( .A1(net83381), .A2(n3781), .ZN(n3782) );
  NOR3_X2 U2315 ( .A1(u4_N1408), .A2(u4_N1409), .A3(u4_N1410), .ZN(n3647) );
  NOR2_X2 U2316 ( .A1(n4119), .A2(net83064), .ZN(n3931) );
  AOI21_X2 U2317 ( .B1(n3967), .B2(n3966), .A(n3965), .ZN(n3987) );
  OAI21_X2 U2318 ( .B1(n3985), .B2(n3984), .A(n3983), .ZN(n3986) );
  OAI21_X1 U2319 ( .B1(net83030), .B2(n3765), .A(n3764), .ZN(n3766) );
  NOR2_X1 U2320 ( .A1(exp_ovf_r_0_), .A2(net82856), .ZN(n3529) );
  OAI21_X1 U2321 ( .B1(exp_ovf_r_0_), .B2(n4006), .A(net82929), .ZN(n4008) );
  NAND2_X2 U2322 ( .A1(n1373), .A2(net94004), .ZN(net83991) );
  OAI21_X2 U2323 ( .B1(net83994), .B2(net83783), .A(net83995), .ZN(net83993)
         );
  OAI21_X1 U2324 ( .B1(net83773), .B2(net84079), .A(net83744), .ZN(n2785) );
  AOI22_X2 U2325 ( .A1(u4_exp_f2i_1[54]), .A2(n2652), .B1(n1373), .B2(n2787), 
        .ZN(net84036) );
  OAI21_X1 U2326 ( .B1(net83773), .B2(net84079), .A(net83744), .ZN(n3592) );
  INV_X16 U2327 ( .A(net85937), .ZN(net82029) );
  OAI21_X2 U2328 ( .B1(n2578), .B2(net83396), .A(n2879), .ZN(n2878) );
  NOR2_X2 U2329 ( .A1(net83036), .A2(n2880), .ZN(n2879) );
  NOR2_X1 U2330 ( .A1(fracta_mul[9]), .A2(fracta_mul[8]), .ZN(n2451) );
  INV_X4 U2331 ( .A(exp_r[6]), .ZN(net85932) );
  AOI21_X2 U2332 ( .B1(net83780), .B2(net83775), .A(net83781), .ZN(net83779)
         );
  AOI22_X2 U2333 ( .A1(u4_exp_f2i_1[56]), .A2(n2652), .B1(n1373), .B2(net93671), .ZN(net83777) );
  INV_X8 U2334 ( .A(n4288), .ZN(n4318) );
  NOR2_X1 U2335 ( .A1(n4706), .A2(n4664), .ZN(n4520) );
  NOR2_X2 U2336 ( .A1(n4665), .A2(n4708), .ZN(n4521) );
  NOR2_X2 U2337 ( .A1(n4515), .A2(n4514), .ZN(n4611) );
  NOR2_X1 U2338 ( .A1(n4690), .A2(n4658), .ZN(n4507) );
  NOR2_X1 U2339 ( .A1(n4659), .A2(n4692), .ZN(n4508) );
  NAND2_X2 U2340 ( .A1(n3015), .A2(fract_denorm[25]), .ZN(n3388) );
  NOR2_X1 U2341 ( .A1(div_opa_ldz_r2[4]), .A2(net86532), .ZN(n3454) );
  OAI21_X2 U2342 ( .B1(net85901), .B2(net83385), .A(net86028), .ZN(n3643) );
  NOR2_X1 U2343 ( .A1(n3088), .A2(n3085), .ZN(n3972) );
  NOR2_X1 U2344 ( .A1(n4766), .A2(n3961), .ZN(net83009) );
  NAND3_X2 U2345 ( .A1(n3762), .A2(u4_div_exp1_6_), .A3(n3761), .ZN(n3781) );
  AOI211_X2 U2346 ( .C1(net86027), .C2(net83736), .A(n2531), .B(net83738), 
        .ZN(net95357) );
  NOR3_X2 U2347 ( .A1(n3998), .A2(net83356), .A3(n3646), .ZN(n3645) );
  NOR2_X2 U2348 ( .A1(n2821), .A2(n2822), .ZN(net84049) );
  NAND3_X2 U2349 ( .A1(n2823), .A2(net83918), .A3(n2824), .ZN(net84044) );
  NOR2_X1 U2350 ( .A1(net85929), .A2(net84054), .ZN(n2824) );
  INV_X4 U2351 ( .A(net83802), .ZN(net83846) );
  NOR2_X2 U2352 ( .A1(n4501), .A2(n4500), .ZN(n4639) );
  OAI21_X1 U2353 ( .B1(n4541), .B2(n4555), .A(n4540), .ZN(n4542) );
  AOI211_X2 U2354 ( .C1(n5289), .C2(n5292), .A(n5293), .B(n4550), .ZN(n4541)
         );
  NOR2_X1 U2355 ( .A1(n5291), .A2(n4544), .ZN(n4547) );
  NAND3_X2 U2356 ( .A1(n3133), .A2(n2908), .A3(n2579), .ZN(net84736) );
  AOI22_X2 U2357 ( .A1(n3238), .A2(prod[42]), .B1(fract_i2f[42]), .B2(net85115), .ZN(n3242) );
  NOR2_X1 U2358 ( .A1(rmode_r3[0]), .A2(net86032), .ZN(n3674) );
  NAND3_X1 U2359 ( .A1(n3670), .A2(net82029), .A3(n2577), .ZN(n3671) );
  AOI211_X2 U2360 ( .C1(net83854), .C2(n3544), .A(n3543), .B(n3542), .ZN(n3547) );
  NOR3_X1 U2361 ( .A1(prod[36]), .A2(prod[42]), .A3(prod[43]), .ZN(n4045) );
  NOR3_X1 U2362 ( .A1(prod[44]), .A2(prod[46]), .A3(prod[45]), .ZN(net82873)
         );
  NAND3_X2 U2363 ( .A1(n4050), .A2(n2712), .A3(n4049), .ZN(n4053) );
  NOR2_X1 U2364 ( .A1(prod[23]), .A2(prod[24]), .ZN(n4050) );
  NOR2_X1 U2365 ( .A1(prod[21]), .A2(prod[20]), .ZN(n4049) );
  NAND3_X2 U2366 ( .A1(n2601), .A2(n2713), .A3(n2569), .ZN(n4051) );
  INV_X4 U2367 ( .A(net83292), .ZN(net93937) );
  AOI21_X2 U2368 ( .B1(net83220), .B2(n2841), .A(net83294), .ZN(net83292) );
  OAI21_X2 U2369 ( .B1(net83278), .B2(net83295), .A(n3818), .ZN(net83294) );
  NOR2_X1 U2370 ( .A1(net82856), .A2(net83367), .ZN(n2845) );
  NOR2_X1 U2371 ( .A1(exp_ovf_r_0_), .A2(net83234), .ZN(n3787) );
  NOR2_X1 U2372 ( .A1(net83041), .A2(net83367), .ZN(n3786) );
  NOR2_X1 U2373 ( .A1(n4645), .A2(n4676), .ZN(n4495) );
  NOR2_X1 U2374 ( .A1(n5288), .A2(n4555), .ZN(n4556) );
  AOI21_X1 U2375 ( .B1(n4554), .B2(n4553), .A(n2715), .ZN(n4557) );
  NOR2_X2 U2376 ( .A1(n4441), .A2(n4440), .ZN(n4445) );
  AOI222_X1 U2377 ( .A1(n4753), .A2(n3734), .B1(u4_div_shft4[1]), .B2(n4755), 
        .C1(u4_div_shft3_1_), .C2(n4754), .ZN(n3520) );
  NOR2_X2 U2378 ( .A1(n4749), .A2(n3504), .ZN(n3505) );
  OAI21_X2 U2379 ( .B1(n3136), .B2(n2908), .A(net84736), .ZN(u4_exp_in_mi1_4_)
         );
  NOR2_X1 U2380 ( .A1(n3088), .A2(n3137), .ZN(n3136) );
  AOI21_X2 U2381 ( .B1(n3487), .B2(n3467), .A(n2668), .ZN(n3469) );
  NOR2_X2 U2382 ( .A1(net85933), .A2(net85929), .ZN(n3467) );
  AOI22_X2 U2383 ( .A1(n3174), .A2(prod[35]), .B1(fract_i2f[35]), .B2(net85115), .ZN(n3257) );
  NAND3_X1 U2384 ( .A1(quo[33]), .A2(net84450), .A3(net85131), .ZN(n3222) );
  NOR2_X2 U2385 ( .A1(n4214), .A2(n4220), .ZN(n4208) );
  NOR2_X2 U2386 ( .A1(n4265), .A2(n4186), .ZN(n4221) );
  NAND4_X2 U2387 ( .A1(n4067), .A2(n3995), .A3(n3994), .A4(n3993), .ZN(n3996)
         );
  NOR2_X2 U2388 ( .A1(net83126), .A2(n3889), .ZN(n3890) );
  NOR2_X2 U2389 ( .A1(opa_r1[23]), .A2(opa_r1[24]), .ZN(n4321) );
  NAND3_X1 U2390 ( .A1(u1_N131), .A2(n3076), .A3(n2600), .ZN(n4464) );
  NOR2_X1 U2391 ( .A1(n4749), .A2(n4748), .ZN(n4750) );
  AOI21_X2 U2392 ( .B1(net82952), .B2(net86045), .A(net86027), .ZN(n3587) );
  AOI21_X2 U2393 ( .B1(n3586), .B2(n2674), .A(net85901), .ZN(n3588) );
  NAND2_X2 U2394 ( .A1(n4010), .A2(net86028), .ZN(n2950) );
  NOR2_X1 U2395 ( .A1(n2577), .A2(net82829), .ZN(n3901) );
  NAND2_X2 U2396 ( .A1(n2989), .A2(net92661), .ZN(n3936) );
  AOI22_X2 U2397 ( .A1(n3856), .A2(net86013), .B1(n3052), .B2(net85997), .ZN(
        n2904) );
  NAND2_X2 U2398 ( .A1(n3895), .A2(u4_fract_out_pl1_13_), .ZN(n2913) );
  OAI21_X1 U2399 ( .B1(n3840), .B2(n3839), .A(net83233), .ZN(net82753) );
  NAND3_X2 U2400 ( .A1(fpu_op_r1[1]), .A2(fpu_op_r1[0]), .A3(n2711), .ZN(n4288) );
  NOR2_X1 U2401 ( .A1(u2_N13), .A2(n4296), .ZN(n4300) );
  NOR2_X2 U2402 ( .A1(n4298), .A2(n4297), .ZN(n4299) );
  NOR2_X1 U2403 ( .A1(u2_N22), .A2(n4290), .ZN(n4294) );
  NOR2_X2 U2404 ( .A1(n4292), .A2(n4291), .ZN(n4293) );
  INV_X4 U2405 ( .A(n4328), .ZN(n4389) );
  NOR2_X2 U2406 ( .A1(u1_fracta_eq_fractb), .A2(n1725), .ZN(n1726) );
  NAND3_X2 U2407 ( .A1(n3837), .A2(n3836), .A3(n3835), .ZN(n4728) );
  AOI21_X1 U2408 ( .B1(n3834), .B2(net82035), .A(n3833), .ZN(n3835) );
  AOI211_X1 U2409 ( .C1(n4524), .C2(n2598), .A(fracta_mul[5]), .B(
        fracta_mul[4]), .ZN(n2453) );
  NAND3_X2 U2410 ( .A1(n2593), .A2(n2699), .A3(n3112), .ZN(n3116) );
  NOR2_X1 U2411 ( .A1(fracta_mul[13]), .A2(n3113), .ZN(n3115) );
  INV_X16 U2412 ( .A(net85399), .ZN(net85397) );
  NAND3_X2 U2413 ( .A1(n4276), .A2(n4275), .A3(n4274), .ZN(u2_N59) );
  NAND3_X2 U2414 ( .A1(n4253), .A2(n4252), .A3(n4251), .ZN(u2_N63) );
  NAND3_X2 U2415 ( .A1(n4263), .A2(n4262), .A3(n4261), .ZN(u2_N61) );
  NAND3_X2 U2416 ( .A1(n2719), .A2(n4241), .A3(n4240), .ZN(u2_N65) );
  AOI222_X1 U2417 ( .A1(u2_exp_tmp3_7_), .A2(n4278), .B1(u2_N49), .B2(n4242), 
        .C1(n4279), .C2(n5253), .ZN(n4240) );
  OAI21_X2 U2418 ( .B1(n4267), .B2(n4266), .A(n4273), .ZN(n4269) );
  NAND2_X2 U2419 ( .A1(net90736), .A2(net91838), .ZN(u4_N1732) );
  NOR2_X2 U2420 ( .A1(n4570), .A2(n4716), .ZN(n4571) );
  NOR2_X2 U2421 ( .A1(n4705), .A2(n4600), .ZN(n4594) );
  NOR2_X2 U2422 ( .A1(n4521), .A2(n4520), .ZN(n4596) );
  NOR2_X2 U2423 ( .A1(n4698), .A2(n4661), .ZN(n4514) );
  NOR2_X2 U2424 ( .A1(n4662), .A2(n4700), .ZN(n4515) );
  OAI21_X1 U2425 ( .B1(div_opa_ldz_r2[0]), .B2(net22501), .A(net83841), .ZN(
        n2818) );
  NOR2_X2 U2426 ( .A1(n4508), .A2(n4507), .ZN(n4625) );
  AOI21_X2 U2427 ( .B1(net83886), .B2(net83888), .A(n2827), .ZN(n2826) );
  NOR2_X1 U2428 ( .A1(n3008), .A2(n3428), .ZN(n3429) );
  NOR2_X1 U2429 ( .A1(n3576), .A2(net86032), .ZN(n3577) );
  INV_X4 U2430 ( .A(net83823), .ZN(n2812) );
  NOR3_X2 U2431 ( .A1(u4_N1417), .A2(u4_N1418), .A3(u4_N1419), .ZN(n3650) );
  NOR3_X2 U2432 ( .A1(u4_N1414), .A2(u4_N1415), .A3(u4_N1416), .ZN(n3649) );
  NOR3_X2 U2433 ( .A1(u4_N1411), .A2(u4_N1412), .A3(u4_N1413), .ZN(n3648) );
  NOR2_X2 U2434 ( .A1(n3734), .A2(net83434), .ZN(n3735) );
  NAND3_X1 U2435 ( .A1(net85937), .A2(net83665), .A3(n2618), .ZN(net83385) );
  NOR2_X2 U2436 ( .A1(n4682), .A2(n4655), .ZN(n4500) );
  NOR2_X2 U2437 ( .A1(n4656), .A2(n4684), .ZN(n4501) );
  NAND3_X2 U2438 ( .A1(net85165), .A2(net85133), .A3(prod[30]), .ZN(n3180) );
  NOR2_X2 U2439 ( .A1(u4_div_exp1_8_), .A2(n3782), .ZN(n3784) );
  NOR2_X2 U2440 ( .A1(n3401), .A2(n3400), .ZN(n3415) );
  NOR2_X1 U2441 ( .A1(net17684), .A2(net84207), .ZN(n3416) );
  NOR2_X2 U2442 ( .A1(net83625), .A2(net83635), .ZN(n2886) );
  AOI21_X2 U2443 ( .B1(n3977), .B2(n3976), .A(n3975), .ZN(n3984) );
  NOR2_X1 U2444 ( .A1(n3985), .A2(net82029), .ZN(n3959) );
  OAI21_X1 U2445 ( .B1(net83009), .B2(net82988), .A(net82999), .ZN(net83007)
         );
  NOR3_X2 U2446 ( .A1(remainder[18]), .A2(remainder[17]), .A3(remainder[16]), 
        .ZN(n3619) );
  NOR3_X2 U2447 ( .A1(remainder[15]), .A2(remainder[14]), .A3(remainder[13]), 
        .ZN(n3620) );
  NOR2_X2 U2448 ( .A1(remainder[28]), .A2(remainder[27]), .ZN(n3636) );
  NOR2_X2 U2449 ( .A1(remainder[1]), .A2(remainder[0]), .ZN(n3625) );
  NOR2_X2 U2450 ( .A1(remainder[3]), .A2(remainder[2]), .ZN(n3624) );
  NOR2_X1 U2451 ( .A1(net85901), .A2(exp_ovf_r_0_), .ZN(n3763) );
  NAND2_X2 U2452 ( .A1(n3744), .A2(net83446), .ZN(n3741) );
  NAND3_X1 U2453 ( .A1(n2659), .A2(n3702), .A3(n3701), .ZN(n3703) );
  NOR2_X1 U2454 ( .A1(net86028), .A2(net83357), .ZN(n3767) );
  NOR2_X1 U2455 ( .A1(net83316), .A2(n3805), .ZN(n3806) );
  NAND2_X2 U2456 ( .A1(n2660), .A2(n2578), .ZN(net83357) );
  NOR2_X1 U2457 ( .A1(opb_r[26]), .A2(n2764), .ZN(n4440) );
  NOR2_X1 U2458 ( .A1(net82856), .A2(net82029), .ZN(n4006) );
  OAI21_X2 U2459 ( .B1(n2583), .B2(net86532), .A(net83775), .ZN(net84014) );
  NOR2_X2 U2460 ( .A1(net83233), .A2(n2577), .ZN(net84015) );
  NOR2_X2 U2461 ( .A1(net83428), .A2(n3709), .ZN(n3710) );
  NOR2_X2 U2462 ( .A1(net83428), .A2(n2807), .ZN(n2803) );
  NOR2_X2 U2463 ( .A1(net82029), .A2(net83434), .ZN(n2804) );
  NOR2_X2 U2464 ( .A1(net83431), .A2(n3694), .ZN(n3698) );
  NOR2_X2 U2465 ( .A1(net83428), .A2(n3691), .ZN(n3699) );
  NAND3_X1 U2466 ( .A1(n3817), .A2(net83297), .A3(n3816), .ZN(net83295) );
  INV_X8 U2467 ( .A(net83357), .ZN(net83234) );
  NAND3_X2 U2468 ( .A1(n4217), .A2(n4214), .A3(n4218), .ZN(n4212) );
  NOR2_X2 U2469 ( .A1(n4315), .A2(n4288), .ZN(n4237) );
  NAND3_X2 U2470 ( .A1(n4264), .A2(n4281), .A3(n4265), .ZN(n4226) );
  INV_X4 U2471 ( .A(net83965), .ZN(net83963) );
  NAND3_X2 U2472 ( .A1(n3547), .A2(n3546), .A3(n3545), .ZN(u4_shift_left[4])
         );
  NOR2_X2 U2473 ( .A1(net83773), .A2(net83783), .ZN(net83780) );
  NOR2_X2 U2474 ( .A1(n2684), .A2(n3909), .ZN(n3912) );
  NOR2_X2 U2475 ( .A1(n3910), .A2(n2728), .ZN(n3911) );
  NAND3_X2 U2476 ( .A1(opb_inf), .A2(opa_inf), .A3(sign_exe_r), .ZN(n3903) );
  INV_X4 U2477 ( .A(net84043), .ZN(net83749) );
  NOR3_X2 U2478 ( .A1(n4053), .A2(n4052), .A3(n4051), .ZN(n4054) );
  NAND3_X2 U2479 ( .A1(n2717), .A2(n2602), .A3(n2568), .ZN(n4052) );
  NOR2_X1 U2480 ( .A1(net85901), .A2(net82036), .ZN(n3948) );
  NOR2_X2 U2481 ( .A1(net83036), .A2(n2704), .ZN(n2829) );
  OAI21_X1 U2482 ( .B1(n2843), .B2(n2844), .A(net83356), .ZN(net83405) );
  NOR2_X1 U2483 ( .A1(net86027), .A2(net83408), .ZN(n2844) );
  NOR2_X1 U2484 ( .A1(net83409), .A2(net82925), .ZN(n2843) );
  NAND3_X1 U2485 ( .A1(net86027), .A2(net85901), .A3(n2674), .ZN(net83325) );
  NOR2_X1 U2486 ( .A1(net83113), .A2(n2709), .ZN(n3838) );
  NOR2_X1 U2487 ( .A1(n4231), .A2(n4193), .ZN(n4195) );
  NOR2_X1 U2488 ( .A1(n4675), .A2(n4650), .ZN(n4651) );
  AOI21_X2 U2489 ( .B1(n4560), .B2(n4559), .A(u1_exp_diff_sft_4_), .ZN(n4561)
         );
  INV_X4 U2490 ( .A(n4452), .ZN(n4453) );
  NOR3_X1 U2491 ( .A1(n1746), .A2(fracta_mul[10]), .A3(fracta_mul[0]), .ZN(
        n1742) );
  NAND3_X2 U2492 ( .A1(n2437), .A2(n2697), .A3(n2444), .ZN(n1746) );
  NOR3_X1 U2493 ( .A1(fracta_mul[13]), .A2(fracta_mul[9]), .A3(fracta_mul[7]), 
        .ZN(n2444) );
  NAND3_X2 U2494 ( .A1(n3508), .A2(n3507), .A3(n3506), .ZN(u4_shift_right[3])
         );
  OAI21_X2 U2495 ( .B1(net84737), .B2(net82988), .A(net84738), .ZN(
        u4_exp_in_mi1_5_) );
  NOR2_X2 U2496 ( .A1(n4749), .A2(n3488), .ZN(n3489) );
  NOR2_X2 U2497 ( .A1(n4749), .A2(n3498), .ZN(n3499) );
  OAI21_X1 U2498 ( .B1(u2_exp_tmp4_5_), .B2(n4208), .A(n4207), .ZN(n4209) );
  OAI21_X1 U2499 ( .B1(u2_exp_tmp4_3_), .B2(n4221), .A(n4220), .ZN(n4222) );
  NOR2_X1 U2500 ( .A1(n4265), .A2(n4264), .ZN(n4267) );
  NOR3_X2 U2501 ( .A1(net83045), .A2(n3941), .A3(opa_inf), .ZN(net83044) );
  AOI21_X2 U2502 ( .B1(n3940), .B2(n3939), .A(opb_inf), .ZN(net83042) );
  NAND3_X1 U2503 ( .A1(n2594), .A2(n4110), .A3(net82035), .ZN(n3939) );
  NOR2_X1 U2504 ( .A1(net83924), .A2(net83761), .ZN(n3534) );
  NAND3_X2 U2505 ( .A1(n4005), .A2(net82934), .A3(n4004), .ZN(n4019) );
  INV_X4 U2506 ( .A(n2898), .ZN(n4085) );
  NOR2_X2 U2507 ( .A1(fpu_op_r2[1]), .A2(fpu_op_r2[2]), .ZN(n2426) );
  INV_X4 U2508 ( .A(n4329), .ZN(n4384) );
  NOR2_X2 U2509 ( .A1(opa_r1[29]), .A2(opa_r1[30]), .ZN(n4324) );
  NOR2_X2 U2510 ( .A1(opa_r1[27]), .A2(opa_r1[28]), .ZN(n4323) );
  NOR2_X2 U2511 ( .A1(opa_r1[25]), .A2(opa_r1[26]), .ZN(n4322) );
  INV_X8 U2512 ( .A(n3073), .ZN(n3074) );
  NAND3_X1 U2513 ( .A1(n4456), .A2(n4455), .A3(n4454), .ZN(n4463) );
  NOR2_X2 U2514 ( .A1(n4305), .A2(n4304), .ZN(n4308) );
  NOR3_X1 U2515 ( .A1(n4730), .A2(n2566), .A3(n2653), .ZN(n4733) );
  NOR3_X1 U2516 ( .A1(n4731), .A2(n2764), .A3(n2765), .ZN(n4732) );
  NOR3_X1 U2517 ( .A1(n4738), .A2(n4737), .A3(n4736), .ZN(n4739) );
  NOR3_X1 U2518 ( .A1(n4735), .A2(n4734), .A3(n3065), .ZN(n4740) );
  AOI21_X1 U2519 ( .B1(n2690), .B2(n5319), .A(fracta_mul[5]), .ZN(n2443) );
  AOI21_X1 U2520 ( .B1(n3125), .B2(n2692), .A(fracta_mul[13]), .ZN(n3127) );
  OAI21_X1 U2521 ( .B1(n2695), .B2(fracta_mul[9]), .A(n2593), .ZN(n3124) );
  OAI21_X1 U2522 ( .B1(fracta_mul[19]), .B2(n3128), .A(n2683), .ZN(n3129) );
  AOI21_X1 U2523 ( .B1(fracta_mul[16]), .B2(n2590), .A(fracta_mul[18]), .ZN(
        n3128) );
  NOR2_X1 U2524 ( .A1(fracta_mul[10]), .A2(n3111), .ZN(n3105) );
  NOR2_X1 U2525 ( .A1(n2051), .A2(fracta_mul[12]), .ZN(n3104) );
  NOR2_X1 U2526 ( .A1(fracta_mul[16]), .A2(fracta_mul[19]), .ZN(n3107) );
  OAI21_X2 U2527 ( .B1(u4_exp_in_pl1_7_), .B2(u4_exp_in_pl1_6_), .A(n3582), 
        .ZN(n3583) );
  AOI21_X2 U2528 ( .B1(net85933), .B2(n3581), .A(net85937), .ZN(n3584) );
  NOR2_X1 U2529 ( .A1(exp_ovf_r_0_), .A2(net82040), .ZN(net82039) );
  NOR2_X2 U2530 ( .A1(n2684), .A2(n3933), .ZN(n3934) );
  NOR2_X1 U2531 ( .A1(net82782), .A2(n4078), .ZN(n4079) );
  NOR2_X1 U2532 ( .A1(net82782), .A2(n4085), .ZN(n4086) );
  INV_X4 U2533 ( .A(n2776), .ZN(net82778) );
  OAI21_X2 U2534 ( .B1(n2777), .B2(net85985), .A(net85975), .ZN(n2776) );
  NOR2_X2 U2535 ( .A1(n1821), .A2(n1822), .ZN(N540) );
  NOR2_X1 U2536 ( .A1(n4289), .A2(n2566), .ZN(u2_exp_ovf_d_0_) );
  NOR2_X2 U2537 ( .A1(n4309), .A2(n4312), .ZN(u2_underflow_d[2]) );
  NOR2_X1 U2538 ( .A1(n4476), .A2(n4465), .ZN(u1_N44) );
  NOR2_X1 U2539 ( .A1(n4476), .A2(n4466), .ZN(u1_N43) );
  NOR2_X1 U2540 ( .A1(n4476), .A2(n4468), .ZN(u1_N42) );
  NOR2_X1 U2541 ( .A1(n4476), .A2(n4470), .ZN(u1_N41) );
  NOR2_X1 U2542 ( .A1(n4476), .A2(n4471), .ZN(u1_N40) );
  NOR2_X1 U2543 ( .A1(n4476), .A2(n4472), .ZN(u1_N39) );
  NOR2_X1 U2544 ( .A1(n4476), .A2(n4474), .ZN(u1_N38) );
  NOR2_X1 U2545 ( .A1(n4477), .A2(n4476), .ZN(u1_N37) );
  OAI21_X2 U2546 ( .B1(n1722), .B2(n2748), .A(n1723), .ZN(u1_N140) );
  OAI21_X2 U2547 ( .B1(n1724), .B2(n2751), .A(u1_signa_r), .ZN(n1723) );
  NOR3_X2 U2548 ( .A1(n1725), .A2(u1_fracta_lt_fractb), .A3(
        u1_fracta_eq_fractb), .ZN(n1724) );
  NOR2_X1 U2549 ( .A1(net85115), .A2(n4729), .ZN(N524) );
  NOR2_X2 U2550 ( .A1(n1733), .A2(n1732), .ZN(u0_N6) );
  NOR2_X1 U2551 ( .A1(fracta_mul[22]), .A2(n1735), .ZN(u0_N4) );
  NOR3_X2 U2552 ( .A1(n2752), .A2(opa_nan), .A3(n1823), .ZN(N532) );
  NOR2_X2 U2553 ( .A1(n4762), .A2(n4743), .ZN(u0_N10) );
  NOR2_X2 U2554 ( .A1(n4763), .A2(n4744), .ZN(u0_N11) );
  NAND3_X2 U2555 ( .A1(n2435), .A2(n3131), .A3(n3130), .ZN(N170) );
  AOI21_X1 U2556 ( .B1(n2599), .B2(n3129), .A(fracta_mul[22]), .ZN(n3130) );
  OAI21_X2 U2557 ( .B1(n3127), .B2(n3126), .A(n2437), .ZN(n3131) );
  OAI21_X1 U2558 ( .B1(n2443), .B2(fracta_mul[6]), .A(n5318), .ZN(n2435) );
  NOR2_X1 U2559 ( .A1(n3123), .A2(fracta_mul[22]), .ZN(N141) );
  NOR2_X1 U2560 ( .A1(fracta_mul[19]), .A2(fracta_mul[18]), .ZN(n3122) );
  AOI21_X2 U2561 ( .B1(n3119), .B2(n3118), .A(n3117), .ZN(N107) );
  NAND3_X2 U2562 ( .A1(n3116), .A2(n3115), .A3(n3114), .ZN(n3118) );
  NOR2_X1 U2563 ( .A1(fracta_mul[15]), .A2(fracta_mul[14]), .ZN(n3114) );
  NOR2_X1 U2564 ( .A1(net86027), .A2(net82034), .ZN(n4745) );
  NOR3_X2 U2565 ( .A1(u4_N1370), .A2(u4_N1372), .A3(u4_N1371), .ZN(n2264) );
  NOR3_X2 U2566 ( .A1(u4_N1373), .A2(u4_N1375), .A3(u4_N1374), .ZN(n2265) );
  NOR3_X2 U2567 ( .A1(u4_N1376), .A2(u4_N1378), .A3(u4_N1377), .ZN(n2266) );
  NOR3_X2 U2568 ( .A1(u4_N1379), .A2(u4_N1381), .A3(u4_N1380), .ZN(n2267) );
  NOR3_X2 U2569 ( .A1(u4_N1358), .A2(u4_N1360), .A3(u4_N1359), .ZN(n2260) );
  NOR3_X2 U2570 ( .A1(u4_N1364), .A2(u4_N1366), .A3(u4_N1365), .ZN(n2262) );
  NOR3_X2 U2571 ( .A1(u4_N1367), .A2(u4_N1369), .A3(u4_N1368), .ZN(n2263) );
  AND2_X4 U2572 ( .A1(n4362), .A2(n5321), .ZN(n2565) );
  INV_X4 U2573 ( .A(n4277), .ZN(n4242) );
  INV_X1 U2574 ( .A(opb_r[30]), .ZN(n3065) );
  INV_X16 U2575 ( .A(net85125), .ZN(net85119) );
  INV_X16 U2576 ( .A(net82826), .ZN(net82782) );
  INV_X8 U2577 ( .A(n2917), .ZN(n3479) );
  INV_X8 U2578 ( .A(net82916), .ZN(net86027) );
  INV_X2 U2579 ( .A(n4277), .ZN(n4249) );
  INV_X4 U2580 ( .A(n4109), .ZN(n3150) );
  INV_X4 U2581 ( .A(n4109), .ZN(n4071) );
  AND3_X4 U2582 ( .A1(net84300), .A2(net84231), .A3(net92895), .ZN(n2571) );
  OR2_X4 U2583 ( .A1(net83282), .A2(net94374), .ZN(n2572) );
  OR2_X4 U2584 ( .A1(net83282), .A2(n3827), .ZN(n2573) );
  OR2_X1 U2585 ( .A1(net83282), .A2(n3823), .ZN(n2574) );
  AND2_X2 U2586 ( .A1(n3795), .A2(net83328), .ZN(n2575) );
  OR2_X1 U2587 ( .A1(net83282), .A2(net83262), .ZN(n2576) );
  INV_X4 U2588 ( .A(net83416), .ZN(net83441) );
  AND2_X4 U2589 ( .A1(net84080), .A2(net85159), .ZN(n2580) );
  AND2_X4 U2590 ( .A1(net84082), .A2(n2798), .ZN(n2583) );
  AND2_X4 U2591 ( .A1(net83596), .A2(net83487), .ZN(n2585) );
  AND2_X4 U2592 ( .A1(n3109), .A2(n2723), .ZN(n2587) );
  AND2_X4 U2593 ( .A1(n5321), .A2(n5322), .ZN(n2588) );
  AND3_X4 U2594 ( .A1(n2883), .A2(net83248), .A3(net83045), .ZN(n2595) );
  AND2_X4 U2595 ( .A1(n2723), .A2(n3110), .ZN(n2597) );
  XOR2_X2 U2596 ( .A(n4439), .B(n2700), .Z(n2600) );
  AND2_X2 U2597 ( .A1(net86027), .A2(n3978), .ZN(n2603) );
  AND3_X4 U2598 ( .A1(n4308), .A2(n4307), .A3(n4306), .ZN(n2604) );
  AND2_X2 U2599 ( .A1(u4_div_shft3_4_), .A2(n2741), .ZN(n2606) );
  OR2_X2 U2600 ( .A1(net83126), .A2(n3858), .ZN(n2619) );
  AND2_X4 U2601 ( .A1(fract_i2f[41]), .A2(net85115), .ZN(n2620) );
  OR2_X2 U2602 ( .A1(rmode_r3[1]), .A2(net83497), .ZN(n2621) );
  AND2_X2 U2603 ( .A1(net17692), .A2(net84202), .ZN(n2622) );
  AND2_X2 U2604 ( .A1(fract_i2f[30]), .A2(net85115), .ZN(n2623) );
  OR2_X2 U2605 ( .A1(net83126), .A2(n3866), .ZN(n2624) );
  AND2_X2 U2606 ( .A1(u4_exp_fix_divb[3]), .A2(net95605), .ZN(n2626) );
  OR2_X2 U2607 ( .A1(net83061), .A2(n2835), .ZN(n2637) );
  AND2_X4 U2608 ( .A1(n3184), .A2(n3185), .ZN(n2638) );
  OR2_X2 U2609 ( .A1(net83126), .A2(n3853), .ZN(n2640) );
  OR2_X2 U2610 ( .A1(net83126), .A2(n3777), .ZN(n2641) );
  AND2_X2 U2611 ( .A1(fract_i2f[26]), .A2(net85115), .ZN(n2643) );
  OR2_X2 U2612 ( .A1(net83126), .A2(n3862), .ZN(n2644) );
  AND3_X4 U2613 ( .A1(n3776), .A2(n3774), .A3(n3775), .ZN(n2645) );
  AND3_X4 U2614 ( .A1(net83113), .A2(net83808), .A3(net83350), .ZN(n2652) );
  INV_X16 U2615 ( .A(net86044), .ZN(net86045) );
  INV_X16 U2616 ( .A(net83374), .ZN(net86044) );
  XOR2_X2 U2617 ( .A(n3137), .B(n2579), .Z(n2656) );
  AND2_X4 U2618 ( .A1(n3802), .A2(n3801), .ZN(n2658) );
  AND2_X2 U2619 ( .A1(net95138), .A2(net86032), .ZN(n2659) );
  INV_X4 U2620 ( .A(n2908), .ZN(n3085) );
  AND2_X2 U2621 ( .A1(n3465), .A2(n3088), .ZN(n2661) );
  AND2_X4 U2622 ( .A1(net83535), .A2(net83534), .ZN(n2662) );
  AND2_X2 U2623 ( .A1(net83878), .A2(n2798), .ZN(n2663) );
  AND2_X2 U2624 ( .A1(n4664), .A2(n4706), .ZN(n2664) );
  AND2_X2 U2625 ( .A1(net85115), .A2(n4019), .ZN(n2665) );
  AND2_X2 U2626 ( .A1(n2981), .A2(n3396), .ZN(n2666) );
  OR2_X2 U2627 ( .A1(net83316), .A2(net83510), .ZN(n2667) );
  INV_X16 U2628 ( .A(net85928), .ZN(net85929) );
  INV_X8 U2629 ( .A(net85929), .ZN(net82988) );
  AND2_X2 U2630 ( .A1(net83642), .A2(n3660), .ZN(n2669) );
  NOR2_X2 U2631 ( .A1(u4_shift_right[7]), .A2(u4_shift_right[6]), .ZN(n2670)
         );
  AND2_X2 U2632 ( .A1(net83963), .A2(n3599), .ZN(n2671) );
  AND2_X4 U2633 ( .A1(n2595), .A2(net83325), .ZN(n2673) );
  NAND2_X2 U2634 ( .A1(u2_N124), .A2(n2930), .ZN(n5317) );
  INV_X4 U2635 ( .A(net82753), .ZN(net82757) );
  AND2_X2 U2636 ( .A1(net83070), .A2(net82035), .ZN(n2684) );
  AND2_X4 U2637 ( .A1(n2595), .A2(net83297), .ZN(n2686) );
  INV_X2 U2638 ( .A(n4277), .ZN(n4254) );
  OR4_X4 U2639 ( .A1(fracta_mul[7]), .A2(fracta_mul[6]), .A3(fracta_mul[5]), 
        .A4(fracta_mul[4]), .ZN(n2699) );
  AND2_X2 U2640 ( .A1(sign), .A2(rmode_r3[1]), .ZN(n2704) );
  OR2_X4 U2641 ( .A1(u4_fi_ldz_2a_6_), .A2(net86045), .ZN(n2710) );
  OR2_X2 U2642 ( .A1(net86027), .A2(net83474), .ZN(n2714) );
  AND3_X4 U2643 ( .A1(n4554), .A2(n4538), .A3(n4537), .ZN(n2715) );
  XOR2_X2 U2644 ( .A(n4318), .B(n4230), .Z(n2716) );
  NOR2_X2 U2645 ( .A1(net83350), .A2(net86032), .ZN(n4003) );
  OR2_X4 U2646 ( .A1(n2802), .A2(net83358), .ZN(n2718) );
  OR2_X4 U2647 ( .A1(n4231), .A2(n4243), .ZN(n2719) );
  AND2_X2 U2648 ( .A1(n3077), .A2(u1_adj_op_out_sft_2_), .ZN(n2720) );
  AND2_X2 U2649 ( .A1(n3078), .A2(u1_adj_op_out_sft_1_), .ZN(n2721) );
  AND3_X4 U2650 ( .A1(n4532), .A2(n4540), .A3(n4531), .ZN(n2722) );
  AND4_X4 U2651 ( .A1(n3108), .A2(n2590), .A3(n2677), .A4(n3107), .ZN(n2723)
         );
  AND2_X2 U2652 ( .A1(n4661), .A2(n4698), .ZN(n2724) );
  AND2_X2 U2653 ( .A1(n4658), .A2(n4690), .ZN(n2725) );
  AND2_X2 U2654 ( .A1(n4655), .A2(n4682), .ZN(n2726) );
  AND2_X2 U2655 ( .A1(u4_div_shft3_2_), .A2(n3611), .ZN(n2727) );
  INV_X4 U2656 ( .A(net85985), .ZN(net85990) );
  OR2_X1 U2657 ( .A1(n3089), .A2(n3091), .ZN(n2729) );
  OR2_X4 U2658 ( .A1(opa_inf), .A2(opb_00), .ZN(n2735) );
  AND3_X4 U2659 ( .A1(n4316), .A2(n4315), .A3(n4317), .ZN(n2739) );
  OR2_X4 U2660 ( .A1(net82856), .A2(n2674), .ZN(n2740) );
  OR2_X4 U2661 ( .A1(u4_div_shft3_3_), .A2(n2727), .ZN(n2741) );
  AND2_X4 U2662 ( .A1(n3915), .A2(n3914), .ZN(n2742) );
  AND2_X4 U2663 ( .A1(n4014), .A2(n4065), .ZN(n2743) );
  OR2_X4 U2664 ( .A1(n4265), .A2(n4288), .ZN(n2744) );
  OR2_X4 U2665 ( .A1(net85901), .A2(net82856), .ZN(n2745) );
  INV_X2 U2666 ( .A(n3692), .ZN(n3982) );
  AND2_X4 U2667 ( .A1(n2605), .A2(n2684), .ZN(n2746) );
  INV_X1 U2668 ( .A(n4764), .ZN(n3094) );
  INV_X1 U2669 ( .A(u2_N124), .ZN(n4764) );
  INV_X4 U2670 ( .A(n3094), .ZN(n3092) );
  INV_X4 U2671 ( .A(n3094), .ZN(n3093) );
  INV_X16 U2672 ( .A(net85904), .ZN(net85905) );
  INV_X4 U2673 ( .A(n2609), .ZN(n3095) );
  INV_X8 U2674 ( .A(n4487), .ZN(n4489) );
  NAND3_X1 U2675 ( .A1(u1_exp_diff2[2]), .A2(n4488), .A3(n4487), .ZN(n4544) );
  OAI21_X2 U2676 ( .B1(u1_exp_diff2[3]), .B2(n4489), .A(n4488), .ZN(n4555) );
  NAND3_X2 U2677 ( .A1(u1_exp_diff2[3]), .A2(u1_exp_diff2[2]), .A3(
        u1_exp_diff2[4]), .ZN(n4482) );
  AOI21_X1 U2678 ( .B1(n5290), .B2(n4550), .A(n5296), .ZN(n4552) );
  INV_X8 U2679 ( .A(n4555), .ZN(n5291) );
  INV_X8 U2680 ( .A(n4551), .ZN(n5289) );
  NOR2_X2 U2681 ( .A1(n4532), .A2(n4551), .ZN(n4543) );
  OAI21_X2 U2682 ( .B1(n4545), .B2(n4551), .A(n2722), .ZN(n4546) );
  NOR2_X2 U2683 ( .A1(n4552), .A2(n4551), .ZN(n4558) );
  OAI211_X1 U2684 ( .C1(opa_r[23]), .C2(n4475), .A(n4458), .B(n4457), .ZN(
        n4462) );
  NOR2_X2 U2685 ( .A1(opa_r[23]), .A2(opa_r[24]), .ZN(n3100) );
  NOR2_X2 U2686 ( .A1(opa_r[27]), .A2(opa_r[28]), .ZN(n3102) );
  NAND2_X1 U2687 ( .A1(opa_r[27]), .A2(opa_r[28]), .ZN(n4730) );
  NAND2_X1 U2688 ( .A1(opa_r[23]), .A2(opa_r[24]), .ZN(n4731) );
  NOR2_X2 U2689 ( .A1(opa_r[25]), .A2(opa_r[26]), .ZN(n3101) );
  OAI21_X4 U2690 ( .B1(opb_r[30]), .B2(n2566), .A(n4453), .ZN(n4672) );
  OAI211_X4 U2691 ( .C1(n4649), .C2(n4648), .A(n4647), .B(n4646), .ZN(n4652)
         );
  OAI211_X4 U2692 ( .C1(n4591), .C2(n4590), .A(n4589), .B(n4588), .ZN(n4595)
         );
  OAI211_X4 U2693 ( .C1(n4606), .C2(n4605), .A(n4604), .B(n4603), .ZN(n4610)
         );
  OAI211_X4 U2694 ( .C1(n4621), .C2(n4620), .A(n4619), .B(n4618), .ZN(n4624)
         );
  OAI211_X4 U2695 ( .C1(n4635), .C2(n4634), .A(n4633), .B(n4632), .ZN(n4638)
         );
  INV_X8 U2696 ( .A(n4672), .ZN(n4670) );
  NAND2_X1 U2697 ( .A1(n4562), .A2(n4672), .ZN(n4671) );
  NOR2_X2 U2698 ( .A1(n4673), .A2(n4672), .ZN(n4725) );
  NOR2_X2 U2699 ( .A1(n4120), .A2(n3950), .ZN(n3951) );
  NOR2_X2 U2700 ( .A1(n4121), .A2(n4120), .ZN(n3831) );
  INV_X4 U2701 ( .A(n2768), .ZN(n2769) );
  NOR4_X1 U2702 ( .A1(n1753), .A2(u6_N4), .A3(u6_N6), .A4(u6_N5), .ZN(n1752)
         );
  AOI21_X2 U2703 ( .B1(n4115), .B2(n4112), .A(n4111), .ZN(n4117) );
  AND2_X2 U2704 ( .A1(n4039), .A2(net85975), .ZN(n2773) );
  OAI21_X2 U2705 ( .B1(n4117), .B2(net82767), .A(n4116), .ZN(N519) );
  NOR3_X2 U2706 ( .A1(net82957), .A2(net86028), .A3(n4002), .ZN(n3993) );
  AOI21_X2 U2707 ( .B1(n4003), .B2(net82029), .A(n4002), .ZN(n4004) );
  OR2_X2 U2708 ( .A1(net82782), .A2(n2893), .ZN(n2777) );
  INV_X16 U2709 ( .A(net82781), .ZN(net85975) );
  NAND2_X1 U2710 ( .A1(n2949), .A2(net82902), .ZN(n4010) );
  INV_X4 U2711 ( .A(net85976), .ZN(net91733) );
  AOI211_X2 U2712 ( .C1(n4084), .C2(net85987), .A(net82757), .B(net85976), 
        .ZN(N451) );
  INV_X1 U2713 ( .A(u6_N7), .ZN(n4517) );
  NOR2_X2 U2714 ( .A1(net82762), .A2(n2831), .ZN(n3954) );
  INV_X4 U2715 ( .A(net84150), .ZN(net84286) );
  NAND2_X2 U2716 ( .A1(n3402), .A2(n3397), .ZN(net84150) );
  AOI22_X4 U2717 ( .A1(n2780), .A2(net85997), .B1(n3890), .B2(net86013), .ZN(
        n2779) );
  OR2_X2 U2718 ( .A1(net83126), .A2(net83168), .ZN(net92365) );
  OAI21_X2 U2719 ( .B1(net83068), .B2(n3815), .A(net93937), .ZN(n2954) );
  AND2_X4 U2720 ( .A1(net82998), .A2(net86027), .ZN(net93471) );
  INV_X1 U2721 ( .A(net93471), .ZN(net83802) );
  MUX2_X2 U2722 ( .A(net93471), .B(n2580), .S(net22501), .Z(net92408) );
  NAND2_X1 U2723 ( .A1(net84076), .A2(net85121), .ZN(net82916) );
  INV_X1 U2724 ( .A(net84077), .ZN(net84076) );
  OAI21_X4 U2725 ( .B1(net83930), .B2(net82998), .A(net83233), .ZN(net83832)
         );
  NAND2_X4 U2726 ( .A1(net85135), .A2(net85159), .ZN(net84077) );
  NOR2_X2 U2727 ( .A1(net84077), .A2(net85175), .ZN(net84568) );
  NOR2_X1 U2728 ( .A1(net85115), .A2(net84077), .ZN(net84496) );
  INV_X8 U2729 ( .A(net85169), .ZN(net85167) );
  INV_X4 U2730 ( .A(net85169), .ZN(net85165) );
  INV_X16 U2731 ( .A(net85141), .ZN(net85135) );
  OR2_X4 U2732 ( .A1(u4_N1732), .A2(net48876), .ZN(u4_N1733) );
  NOR2_X4 U2733 ( .A1(u4_exp_out_2_), .A2(u4_exp_out_1_), .ZN(net91838) );
  NOR2_X4 U2734 ( .A1(net92815), .A2(net92816), .ZN(net90736) );
  NAND2_X4 U2735 ( .A1(n2783), .A2(n2784), .ZN(net92816) );
  INV_X4 U2736 ( .A(u4_exp_out_3_), .ZN(n2784) );
  INV_X8 U2737 ( .A(u4_exp_out_4_), .ZN(n2783) );
  NAND2_X4 U2738 ( .A1(net91045), .A2(net91044), .ZN(net92815) );
  INV_X8 U2739 ( .A(u4_exp_out_5_), .ZN(net91044) );
  NOR2_X4 U2740 ( .A1(u4_N1976), .A2(u4_exp_out_6_), .ZN(net91045) );
  NAND3_X4 U2741 ( .A1(net83971), .A2(net83972), .A3(net83973), .ZN(
        u4_exp_out_2_) );
  AOI21_X2 U2742 ( .B1(net83974), .B2(net83744), .A(net83781), .ZN(net83973)
         );
  INV_X4 U2743 ( .A(net83995), .ZN(net83781) );
  AOI21_X4 U2744 ( .B1(net84014), .B2(net83744), .A(net83781), .ZN(net84013)
         );
  AOI221_X2 U2745 ( .B1(n1373), .B2(net83963), .C1(u4_exp_f2i_1[50]), .C2(
        n2652), .A(net83781), .ZN(net83953) );
  OAI21_X1 U2746 ( .B1(n2782), .B2(n2469), .A(net83580), .ZN(net83974) );
  INV_X2 U2747 ( .A(net84083), .ZN(n2782) );
  NAND2_X1 U2748 ( .A1(n2782), .A2(n2469), .ZN(net83580) );
  NAND2_X2 U2749 ( .A1(net86027), .A2(net83017), .ZN(net83972) );
  NOR2_X4 U2750 ( .A1(net92028), .A2(net85115), .ZN(net84556) );
  INV_X32 U2751 ( .A(net85119), .ZN(net85115) );
  INV_X16 U2752 ( .A(net85141), .ZN(net92028) );
  INV_X16 U2753 ( .A(net85149), .ZN(net85141) );
  INV_X8 U2754 ( .A(net86236), .ZN(net85149) );
  NOR2_X2 U2755 ( .A1(net86235), .A2(net86236), .ZN(net86234) );
  NAND3_X4 U2756 ( .A1(net84036), .A2(n2786), .A3(n2785), .ZN(u4_exp_out_5_)
         );
  BUF_X32 U2757 ( .A(u4_exp_out_5_), .Z(net94896) );
  INV_X4 U2758 ( .A(net83775), .ZN(net84079) );
  NAND2_X4 U2759 ( .A1(net83020), .A2(net86027), .ZN(n2786) );
  INV_X1 U2760 ( .A(net95173), .ZN(n2787) );
  INV_X4 U2761 ( .A(net82940), .ZN(net83808) );
  INV_X4 U2762 ( .A(net86032), .ZN(net83113) );
  INV_X16 U2763 ( .A(n2580), .ZN(net86032) );
  NAND3_X4 U2764 ( .A1(net83778), .A2(net83777), .A3(net83779), .ZN(u4_N1976)
         );
  BUF_X32 U2765 ( .A(u4_N1976), .Z(net95138) );
  INV_X4 U2766 ( .A(net83744), .ZN(net83783) );
  OAI21_X2 U2767 ( .B1(net86532), .B2(net93218), .A(net83773), .ZN(net84138)
         );
  NAND2_X1 U2768 ( .A1(net83773), .A2(net84124), .ZN(net82991) );
  NAND3_X4 U2769 ( .A1(net83828), .A2(n2789), .A3(n2788), .ZN(net83827) );
  NOR2_X4 U2770 ( .A1(net83827), .A2(net83826), .ZN(net83816) );
  NAND2_X1 U2771 ( .A1(n2791), .A2(div_opa_ldz_r2[1]), .ZN(net83863) );
  OAI211_X2 U2772 ( .C1(net94620), .C2(net83831), .A(n2790), .B(net94614), 
        .ZN(n2789) );
  INV_X1 U2773 ( .A(net83836), .ZN(net83834) );
  INV_X2 U2774 ( .A(net83834), .ZN(net95473) );
  INV_X8 U2775 ( .A(net83832), .ZN(net83929) );
  INV_X2 U2776 ( .A(net83929), .ZN(net94620) );
  OAI21_X1 U2777 ( .B1(net83927), .B2(net83928), .A(net83929), .ZN(net83868)
         );
  NOR2_X4 U2778 ( .A1(net83932), .A2(net86028), .ZN(net83931) );
  NOR3_X2 U2779 ( .A1(net83837), .A2(net82965), .A3(net86044), .ZN(net83831)
         );
  NAND2_X4 U2780 ( .A1(net83665), .A2(net82999), .ZN(net83374) );
  INV_X4 U2781 ( .A(net84054), .ZN(net82999) );
  NAND2_X1 U2782 ( .A1(net94933), .A2(net82999), .ZN(net82997) );
  OAI21_X1 U2783 ( .B1(net82999), .B2(net83802), .A(net83803), .ZN(net83801)
         );
  NAND2_X4 U2784 ( .A1(net83788), .A2(net93036), .ZN(n2792) );
  OAI211_X4 U2785 ( .C1(net83785), .C2(net83750), .A(n2792), .B(net83787), 
        .ZN(net83005) );
  INV_X8 U2786 ( .A(net95102), .ZN(net83788) );
  AOI221_X4 U2787 ( .B1(net94516), .B2(net83747), .C1(net83788), .C2(net94514), 
        .A(net94515), .ZN(net94513) );
  INV_X1 U2788 ( .A(net83788), .ZN(net95178) );
  NAND4_X4 U2789 ( .A1(u4_div_exp2_7_), .A2(u4_div_exp2_6_), .A3(net84048), 
        .A4(net84049), .ZN(n2793) );
  NAND3_X4 U2790 ( .A1(n2793), .A2(net84044), .A3(net84046), .ZN(net95102) );
  OAI221_X2 U2791 ( .B1(net84016), .B2(net83750), .C1(net83753), .C2(net84017), 
        .A(net84018), .ZN(net83019) );
  OAI221_X2 U2792 ( .B1(net83957), .B2(net83750), .C1(net83753), .C2(net83958), 
        .A(net83959), .ZN(net83016) );
  NAND3_X4 U2793 ( .A1(n2793), .A2(net84044), .A3(net84046), .ZN(net83753) );
  NAND3_X4 U2794 ( .A1(net82953), .A2(n2714), .A3(net93714), .ZN(net83668) );
  NAND2_X4 U2795 ( .A1(net83668), .A2(net83667), .ZN(net83605) );
  NOR3_X4 U2796 ( .A1(net83727), .A2(u4_fract_out_15_), .A3(u4_fract_out_16_), 
        .ZN(net83726) );
  INV_X8 U2797 ( .A(n2067), .ZN(u4_fract_out_15_) );
  AOI22_X4 U2798 ( .A1(u4_N1398), .A2(net85377), .B1(u4_N1448), .B2(n2794), 
        .ZN(n2067) );
  NOR3_X4 U2799 ( .A1(net83799), .A2(net83800), .A3(net83801), .ZN(n2794) );
  INV_X4 U2800 ( .A(net83797), .ZN(net83803) );
  OAI221_X1 U2801 ( .B1(net86032), .B2(net83941), .C1(net82988), .C2(net83802), 
        .A(net83943), .ZN(net83921) );
  BUF_X32 U2802 ( .A(u4_exp_out_3_), .Z(net94566) );
  AOI21_X4 U2803 ( .B1(u4_exp_f2i_1[52]), .B2(n2652), .A(net83993), .ZN(n2795)
         );
  NOR2_X4 U2804 ( .A1(n2583), .A2(n2796), .ZN(net83994) );
  INV_X4 U2805 ( .A(n2797), .ZN(n2796) );
  NAND2_X1 U2806 ( .A1(net83580), .A2(net83762), .ZN(n2797) );
  INV_X8 U2807 ( .A(u4_fi_ldz_2a_3_), .ZN(net83762) );
  NAND2_X2 U2808 ( .A1(n2583), .A2(net86532), .ZN(net83775) );
  INV_X1 U2809 ( .A(net83762), .ZN(n2798) );
  NAND3_X1 U2810 ( .A1(net93902), .A2(n2798), .A3(n2469), .ZN(net83756) );
  INV_X1 U2811 ( .A(net83580), .ZN(net84082) );
  NOR3_X4 U2812 ( .A1(u4_fract_out_20_), .A2(net83731), .A3(net83730), .ZN(
        net83723) );
  AOI22_X4 U2813 ( .A1(u4_N1392), .A2(net85377), .B1(u4_N1442), .B2(n2794), 
        .ZN(n1450) );
  NAND2_X4 U2814 ( .A1(net83005), .A2(net86027), .ZN(net83778) );
  BUF_X32 U2815 ( .A(net83005), .Z(net94825) );
  AOI22_X4 U2816 ( .A1(u4_div_exp1_7_), .A2(net83752), .B1(u4_div_exp3[7]), 
        .B2(net83749), .ZN(net83787) );
  INV_X4 U2817 ( .A(net84042), .ZN(net83752) );
  NAND2_X1 U2818 ( .A1(net85175), .A2(net84043), .ZN(net84042) );
  INV_X16 U2819 ( .A(net85179), .ZN(net85175) );
  INV_X16 U2820 ( .A(net85183), .ZN(net85179) );
  INV_X4 U2821 ( .A(net86235), .ZN(net85183) );
  XNOR2_X2 U2822 ( .A(n2799), .B(net93671), .ZN(net83785) );
  INV_X8 U2823 ( .A(n2801), .ZN(n2799) );
  NOR2_X4 U2824 ( .A1(n2799), .A2(net83770), .ZN(net83766) );
  NAND2_X4 U2825 ( .A1(net83771), .A2(n2800), .ZN(n2801) );
  MUX2_X2 U2826 ( .A(net83430), .B(net83791), .S(net93455), .Z(n2800) );
  INV_X4 U2827 ( .A(net85393), .ZN(net93455) );
  INV_X8 U2828 ( .A(net83605), .ZN(net83639) );
  NOR2_X4 U2829 ( .A1(net83041), .A2(n2718), .ZN(net83667) );
  NAND3_X1 U2830 ( .A1(net83356), .A2(n2718), .A3(net83660), .ZN(net83642) );
  INV_X4 U2831 ( .A(net85901), .ZN(net83358) );
  INV_X4 U2832 ( .A(net82939), .ZN(n2802) );
  NOR2_X4 U2833 ( .A1(n2802), .A2(net83233), .ZN(net83744) );
  NAND2_X2 U2834 ( .A1(n2802), .A2(net84015), .ZN(net83995) );
  INV_X8 U2835 ( .A(net83356), .ZN(net83041) );
  NAND2_X2 U2836 ( .A1(net84100), .A2(net83633), .ZN(net82939) );
  NAND3_X2 U2837 ( .A1(net82951), .A2(net82952), .A3(net82939), .ZN(net82950)
         );
  NAND4_X2 U2838 ( .A1(rmode_r3[1]), .A2(rmode_r3[0]), .A3(net82939), .A4(
        opas_r2), .ZN(net84091) );
  NAND4_X2 U2839 ( .A1(net82938), .A2(net82939), .A3(net82029), .A4(net82940), 
        .ZN(net82934) );
  NAND2_X4 U2840 ( .A1(net83259), .A2(net83262), .ZN(net83410) );
  INV_X8 U2841 ( .A(net83410), .ZN(net83402) );
  NAND3_X4 U2842 ( .A1(net83437), .A2(net83436), .A3(net83438), .ZN(net83259)
         );
  NOR3_X4 U2843 ( .A1(net83259), .A2(net83383), .A3(net83384), .ZN(net83279)
         );
  INV_X1 U2844 ( .A(net83259), .ZN(net94373) );
  AOI22_X2 U2845 ( .A1(net83435), .A2(u4_exp_out_pl1_7_), .B1(
        u4_exp_fix_divb[7]), .B2(net95605), .ZN(net83438) );
  NOR3_X4 U2846 ( .A1(n2803), .A2(n2804), .A3(n2805), .ZN(net83436) );
  NOR2_X1 U2847 ( .A1(net83316), .A2(n2806), .ZN(n2805) );
  INV_X1 U2848 ( .A(u4_exp_next_mi_7_), .ZN(n2806) );
  INV_X4 U2849 ( .A(u4_exp_fix_diva[7]), .ZN(n2807) );
  MUX2_X2 U2850 ( .A(net83439), .B(net83440), .S(u4_N1640), .Z(net83437) );
  INV_X1 U2851 ( .A(net95138), .ZN(u4_N1640) );
  OAI221_X1 U2852 ( .B1(net82011), .B2(net82023), .C1(u4_N1640), .C2(net82013), 
        .A(net82024), .ZN(u4_shift_right[7]) );
  OR2_X1 U2853 ( .A1(u4_N1640), .A2(net95138), .ZN(u4_N1977) );
  NAND2_X2 U2854 ( .A1(net83441), .A2(net83442), .ZN(net83440) );
  INV_X1 U2855 ( .A(n2476), .ZN(net83442) );
  NOR3_X4 U2856 ( .A1(net83443), .A2(net83319), .A3(net83444), .ZN(net83439)
         );
  OAI211_X4 U2857 ( .C1(net92626), .C2(net82012), .A(n2808), .B(net83422), 
        .ZN(net83443) );
  NAND2_X4 U2858 ( .A1(net83446), .A2(net94896), .ZN(n2808) );
  INV_X16 U2859 ( .A(net83421), .ZN(net83446) );
  INV_X8 U2860 ( .A(net83446), .ZN(net92626) );
  NAND2_X4 U2861 ( .A1(net82852), .A2(net83113), .ZN(net83052) );
  INV_X8 U2862 ( .A(net83052), .ZN(net83043) );
  INV_X4 U2863 ( .A(net84102), .ZN(net84080) );
  NAND2_X2 U2864 ( .A1(net84080), .A2(net86309), .ZN(net83233) );
  NAND2_X1 U2865 ( .A1(net85115), .A2(net85145), .ZN(net84102) );
  INV_X16 U2866 ( .A(net85149), .ZN(net85145) );
  NOR3_X4 U2867 ( .A1(net83114), .A2(n2475), .A3(net83115), .ZN(net82852) );
  NAND3_X4 U2868 ( .A1(net83198), .A2(net83197), .A3(net83196), .ZN(net83114)
         );
  NOR3_X4 U2869 ( .A1(net83114), .A2(n2475), .A3(net83115), .ZN(net95525) );
  NAND3_X4 U2870 ( .A1(net84387), .A2(n2809), .A3(net84180), .ZN(net83722) );
  NOR2_X4 U2871 ( .A1(net83721), .A2(net83722), .ZN(net84370) );
  INV_X8 U2872 ( .A(net83722), .ZN(net84324) );
  NAND3_X1 U2873 ( .A1(net84180), .A2(net84225), .A3(net94305), .ZN(net84224)
         );
  OAI21_X1 U2874 ( .B1(fract_denorm[44]), .B2(net84180), .A(net84181), .ZN(
        net84178) );
  AOI211_X2 U2875 ( .C1(net84306), .C2(net84180), .A(net85391), .B(
        fract_denorm[45]), .ZN(net84301) );
  NOR2_X4 U2876 ( .A1(fract_denorm[44]), .A2(net86571), .ZN(n2809) );
  INV_X16 U2877 ( .A(net86570), .ZN(net86571) );
  INV_X4 U2878 ( .A(fract_denorm_46_), .ZN(net86570) );
  NAND3_X2 U2879 ( .A1(net84546), .A2(net84547), .A3(net84548), .ZN(
        fract_denorm_46_) );
  NOR2_X2 U2880 ( .A1(net85167), .A2(n2649), .ZN(n2810) );
  NAND3_X2 U2881 ( .A1(net85165), .A2(net85133), .A3(prod[46]), .ZN(net84547)
         );
  INV_X16 U2882 ( .A(net85143), .ZN(net85133) );
  INV_X16 U2883 ( .A(net85149), .ZN(net85143) );
  NAND3_X4 U2884 ( .A1(net83602), .A2(net83601), .A3(n2676), .ZN(net83421) );
  INV_X1 U2885 ( .A(net83601), .ZN(net95279) );
  NAND2_X2 U2886 ( .A1(rmode_r3[1]), .A2(n2676), .ZN(net83343) );
  OAI21_X4 U2887 ( .B1(n2676), .B2(net83348), .A(rmode_r3[1]), .ZN(net83514)
         );
  OAI21_X2 U2888 ( .B1(net83639), .B2(net83606), .A(n2676), .ZN(net83569) );
  NOR2_X4 U2889 ( .A1(n2811), .A2(net82040), .ZN(net83602) );
  NAND2_X4 U2890 ( .A1(u4_fract_out_pl1_23_), .A2(rmode_r3[1]), .ZN(net82038)
         );
  NOR2_X1 U2891 ( .A1(net82038), .A2(net83569), .ZN(net83568) );
  NOR2_X1 U2892 ( .A1(net82038), .A2(net83565), .ZN(net83567) );
  NAND2_X2 U2893 ( .A1(sign), .A2(net83565), .ZN(net83500) );
  NOR2_X4 U2894 ( .A1(net83639), .A2(net83606), .ZN(n2811) );
  NAND2_X2 U2895 ( .A1(net83565), .A2(n2811), .ZN(net83499) );
  INV_X4 U2896 ( .A(net92408), .ZN(net83828) );
  INV_X8 U2897 ( .A(net92066), .ZN(net85904) );
  INV_X4 U2898 ( .A(net92065), .ZN(net92066) );
  NAND3_X4 U2899 ( .A1(net83816), .A2(net83817), .A3(net83818), .ZN(
        u4_shift_left[0]) );
  OAI221_X4 U2900 ( .B1(net82035), .B2(n2812), .C1(n2813), .C2(n2814), .A(
        u4_exp_in_pl1_0_), .ZN(net83818) );
  NAND3_X4 U2901 ( .A1(n2815), .A2(net86045), .A3(net83823), .ZN(n2814) );
  INV_X4 U2902 ( .A(net84738), .ZN(net83665) );
  INV_X4 U2903 ( .A(n2819), .ZN(n2815) );
  NAND3_X4 U2904 ( .A1(net82035), .A2(net86045), .A3(n2815), .ZN(net83870) );
  NOR2_X1 U2905 ( .A1(net85901), .A2(u4_N1733), .ZN(n2819) );
  NOR2_X4 U2906 ( .A1(net85901), .A2(net83824), .ZN(n2813) );
  INV_X8 U2907 ( .A(net82776), .ZN(net82035) );
  OAI211_X2 U2908 ( .C1(net85901), .C2(net83824), .A(n2816), .B(net94614), 
        .ZN(net83817) );
  INV_X4 U2909 ( .A(net83870), .ZN(n2816) );
  OAI221_X2 U2910 ( .B1(net83868), .B2(n2816), .C1(net95242), .C2(net83869), 
        .A(net93902), .ZN(net83842) );
  NOR2_X4 U2911 ( .A1(n2817), .A2(net83811), .ZN(net83826) );
  INV_X4 U2912 ( .A(n2818), .ZN(n2817) );
  INV_X4 U2913 ( .A(net85905), .ZN(net22501) );
  INV_X1 U2914 ( .A(n2476), .ZN(net82012) );
  INV_X1 U2915 ( .A(net82012), .ZN(net92622) );
  NAND2_X1 U2916 ( .A1(net82012), .A2(n2468), .ZN(net92624) );
  OAI221_X2 U2917 ( .B1(net82010), .B2(net82011), .C1(net82012), .C2(net82013), 
        .A(net82014), .ZN(u4_shift_right[6]) );
  NAND2_X4 U2918 ( .A1(net83498), .A2(net83495), .ZN(net83319) );
  INV_X8 U2919 ( .A(net83319), .ZN(net83526) );
  NAND2_X1 U2920 ( .A1(net83319), .A2(net48876), .ZN(net83305) );
  NAND2_X2 U2921 ( .A1(net83527), .A2(net83446), .ZN(net83445) );
  NAND3_X1 U2922 ( .A1(net83422), .A2(net83526), .A3(net83445), .ZN(net83525)
         );
  NAND2_X4 U2923 ( .A1(net83518), .A2(rmode_r3[1]), .ZN(net83422) );
  NAND2_X2 U2924 ( .A1(u4_div_exp2_1_), .A2(u4_div_exp2_0_), .ZN(n2822) );
  NAND2_X2 U2925 ( .A1(u4_div_exp2_3_), .A2(u4_div_exp2_2_), .ZN(n2821) );
  NOR2_X4 U2926 ( .A1(net84017), .A2(n2820), .ZN(net84048) );
  INV_X4 U2927 ( .A(u4_div_exp2_5_), .ZN(n2820) );
  OAI221_X1 U2928 ( .B1(net84016), .B2(net83750), .C1(net84017), .C2(net95178), 
        .A(net84018), .ZN(net95148) );
  INV_X8 U2929 ( .A(exp_r[5]), .ZN(net85928) );
  NAND2_X2 U2930 ( .A1(net84737), .A2(net85928), .ZN(net84738) );
  OAI21_X4 U2931 ( .B1(n2825), .B2(n2826), .A(net83919), .ZN(n2823) );
  NAND2_X2 U2932 ( .A1(net83887), .A2(net83902), .ZN(n2827) );
  INV_X4 U2933 ( .A(net83903), .ZN(n2825) );
  NOR2_X4 U2934 ( .A1(net83749), .A2(n2584), .ZN(net84046) );
  NAND2_X2 U2935 ( .A1(n2584), .A2(net85179), .ZN(net83474) );
  INV_X4 U2936 ( .A(u4_div_exp2_1_), .ZN(net83958) );
  NAND3_X4 U2937 ( .A1(net84559), .A2(net84557), .A3(n2828), .ZN(
        fract_denorm[44]) );
  NAND4_X2 U2938 ( .A1(quo[46]), .A2(net85175), .A3(net85135), .A4(net85159), 
        .ZN(n2828) );
  NOR3_X4 U2939 ( .A1(net82782), .A2(net83074), .A3(net85985), .ZN(net83196)
         );
  INV_X8 U2940 ( .A(net82780), .ZN(net85985) );
  NAND4_X4 U2941 ( .A1(net83344), .A2(n2595), .A3(net86028), .A4(net83345), 
        .ZN(net82780) );
  NOR2_X2 U2942 ( .A1(net23180), .A2(n2829), .ZN(net83345) );
  NAND2_X2 U2943 ( .A1(n2704), .A2(net86027), .ZN(net83359) );
  INV_X4 U2944 ( .A(net83300), .ZN(net83036) );
  INV_X8 U2945 ( .A(net82932), .ZN(net23180) );
  NAND3_X2 U2946 ( .A1(net23180), .A2(net86571), .A3(net83735), .ZN(net83593)
         );
  NAND3_X4 U2947 ( .A1(net82927), .A2(n2595), .A3(net83349), .ZN(net82826) );
  NAND2_X2 U2948 ( .A1(net86497), .A2(u4_fract_out_11_), .ZN(net83166) );
  INV_X4 U2949 ( .A(n1461), .ZN(u4_fract_out_11_) );
  INV_X16 U2950 ( .A(n2505), .ZN(net86497) );
  INV_X4 U2951 ( .A(net86496), .ZN(net95019) );
  AOI22_X4 U2952 ( .A1(u4_N1394), .A2(net85377), .B1(u4_N1444), .B2(n2794), 
        .ZN(n1461) );
  NAND3_X2 U2953 ( .A1(n1451), .A2(n1461), .A3(n1460), .ZN(net83727) );
  NAND2_X4 U2954 ( .A1(n2830), .A2(net83593), .ZN(net48876) );
  AOI211_X4 U2955 ( .C1(net86027), .C2(net83736), .A(n2531), .B(net83738), 
        .ZN(n2830) );
  OAI21_X2 U2956 ( .B1(net83038), .B2(net82829), .A(net83039), .ZN(N531) );
  NAND2_X2 U2957 ( .A1(net83041), .A2(n2839), .ZN(net83039) );
  INV_X2 U2958 ( .A(n2838), .ZN(n2839) );
  INV_X1 U2959 ( .A(n2832), .ZN(n2838) );
  INV_X4 U2960 ( .A(n2833), .ZN(n2832) );
  NAND2_X2 U2961 ( .A1(result_zero_sign_d), .A2(n2832), .ZN(net92661) );
  NOR2_X4 U2962 ( .A1(net83059), .A2(n2637), .ZN(n2834) );
  NAND2_X1 U2963 ( .A1(n2836), .A2(net83068), .ZN(n2835) );
  NOR2_X4 U2964 ( .A1(n2837), .A2(net82767), .ZN(n2836) );
  INV_X8 U2965 ( .A(n2831), .ZN(n2837) );
  NOR2_X2 U2966 ( .A1(net83064), .A2(n2837), .ZN(net83214) );
  NAND2_X4 U2967 ( .A1(net83066), .A2(n2837), .ZN(net83254) );
  OAI21_X4 U2968 ( .B1(net86486), .B2(net83263), .A(n2673), .ZN(n2831) );
  NAND3_X2 U2969 ( .A1(n2087), .A2(n2083), .A3(n2085), .ZN(net83730) );
  AOI22_X4 U2970 ( .A1(u4_N1388), .A2(net85377), .B1(u4_N1438), .B2(n2794), 
        .ZN(n2085) );
  INV_X4 U2971 ( .A(n2085), .ZN(u4_fract_out_5_) );
  INV_X4 U2972 ( .A(net86234), .ZN(net84490) );
  OAI21_X4 U2973 ( .B1(net83402), .B2(net83403), .A(n2841), .ZN(n2842) );
  NAND2_X4 U2974 ( .A1(n2842), .A2(net83278), .ZN(net86012) );
  INV_X4 U2975 ( .A(n2840), .ZN(n2841) );
  OAI21_X2 U2976 ( .B1(net83402), .B2(net83403), .A(n2841), .ZN(net94703) );
  OAI21_X4 U2977 ( .B1(n2845), .B2(net83458), .A(net86027), .ZN(net83403) );
  OAI21_X4 U2978 ( .B1(net83403), .B2(net83404), .A(net83405), .ZN(n2840) );
  INV_X4 U2979 ( .A(net83403), .ZN(net83276) );
  INV_X4 U2980 ( .A(net83404), .ZN(net83458) );
  NOR2_X1 U2981 ( .A1(n2840), .A2(n2465), .ZN(net83326) );
  OAI21_X4 U2982 ( .B1(net83276), .B2(n2840), .A(net83278), .ZN(net83275) );
  INV_X4 U2983 ( .A(net84030), .ZN(net83409) );
  NAND2_X4 U2984 ( .A1(n2856), .A2(net84356), .ZN(net84281) );
  OR4_X4 U2985 ( .A1(n2562), .A2(net17692), .A3(net17654), .A4(net84282), .ZN(
        net95353) );
  INV_X8 U2986 ( .A(n2848), .ZN(net84356) );
  NAND3_X1 U2987 ( .A1(net84189), .A2(net84188), .A3(net84356), .ZN(net84185)
         );
  OAI211_X2 U2988 ( .C1(net17654), .C2(net17692), .A(n2856), .B(net84356), 
        .ZN(net84345) );
  NAND4_X4 U2989 ( .A1(net84300), .A2(n2855), .A3(net84324), .A4(n2850), .ZN(
        n2848) );
  NOR2_X1 U2990 ( .A1(net84375), .A2(n2563), .ZN(net84343) );
  NOR2_X4 U2991 ( .A1(n2848), .A2(net84298), .ZN(net91297) );
  NOR2_X4 U2992 ( .A1(net17686), .A2(fract_denorm[33]), .ZN(n2850) );
  NOR2_X4 U2993 ( .A1(net84323), .A2(net84272), .ZN(n2855) );
  INV_X4 U2994 ( .A(net83721), .ZN(net84300) );
  INV_X1 U2995 ( .A(net84300), .ZN(net92015) );
  NAND3_X2 U2996 ( .A1(net84171), .A2(net84300), .A3(fract_denorm[33]), .ZN(
        net84262) );
  NAND3_X2 U2997 ( .A1(n2853), .A2(n2852), .A3(net91817), .ZN(n2851) );
  NOR2_X4 U2998 ( .A1(net84312), .A2(net83630), .ZN(n2852) );
  NOR3_X4 U2999 ( .A1(net95365), .A2(n2849), .A3(net84191), .ZN(n2853) );
  NAND2_X4 U3000 ( .A1(n2847), .A2(n2846), .ZN(n2849) );
  INV_X8 U3001 ( .A(net17656), .ZN(n2846) );
  AND2_X2 U3002 ( .A1(n2847), .A2(n2846), .ZN(net92738) );
  NAND2_X2 U3003 ( .A1(net83622), .A2(n2846), .ZN(net83621) );
  INV_X8 U3004 ( .A(n2854), .ZN(n2847) );
  NAND2_X1 U3005 ( .A1(n2847), .A2(net83638), .ZN(net83634) );
  NAND4_X2 U3006 ( .A1(net84321), .A2(net17656), .A3(n2847), .A4(net84204), 
        .ZN(net84151) );
  NAND2_X4 U3007 ( .A1(net84411), .A2(net84207), .ZN(n2854) );
  INV_X8 U3008 ( .A(net17685), .ZN(net84207) );
  NAND2_X1 U3009 ( .A1(u4_fract_out_pl1_9_), .A2(net86012), .ZN(net86478) );
  INV_X4 U3010 ( .A(net83343), .ZN(net83278) );
  NAND2_X2 U3011 ( .A1(net83342), .A2(net83343), .ZN(net83328) );
  NAND3_X4 U3012 ( .A1(n2857), .A2(net93416), .A3(n2858), .ZN(net83754) );
  NAND2_X2 U3013 ( .A1(n2859), .A2(net17683), .ZN(n2858) );
  INV_X2 U3014 ( .A(net84275), .ZN(n2859) );
  INV_X8 U3015 ( .A(net84235), .ZN(net93416) );
  NAND4_X2 U3016 ( .A1(net84140), .A2(net93416), .A3(net84143), .A4(net84142), 
        .ZN(net84135) );
  NAND4_X4 U3017 ( .A1(net84236), .A2(net84239), .A3(net84238), .A4(net84237), 
        .ZN(net84235) );
  NOR2_X4 U3018 ( .A1(n2860), .A2(n2866), .ZN(n2857) );
  INV_X4 U3019 ( .A(net17693), .ZN(net84282) );
  NAND2_X2 U3020 ( .A1(net84282), .A2(net83625), .ZN(net84382) );
  NAND3_X4 U3021 ( .A1(net84282), .A2(net84362), .A3(net84202), .ZN(net83635)
         );
  INV_X2 U3022 ( .A(net84242), .ZN(net84280) );
  NAND3_X1 U3023 ( .A1(net84280), .A2(net93422), .A3(net83632), .ZN(net84101)
         );
  NAND3_X2 U3024 ( .A1(net84285), .A2(net84286), .A3(n2865), .ZN(n2860) );
  INV_X4 U3025 ( .A(n2864), .ZN(n2865) );
  NAND2_X2 U3026 ( .A1(net84284), .A2(net84283), .ZN(n2864) );
  AOI21_X4 U3027 ( .B1(net84301), .B2(net84302), .A(n2862), .ZN(net84283) );
  INV_X4 U3028 ( .A(n2863), .ZN(n2862) );
  NAND3_X2 U3029 ( .A1(fract_denorm[36]), .A2(net84305), .A3(net84171), .ZN(
        n2863) );
  INV_X8 U3030 ( .A(net84353), .ZN(net84171) );
  NAND3_X1 U3031 ( .A1(net84171), .A2(net84172), .A3(fract_denorm[37]), .ZN(
        net84167) );
  INV_X4 U3032 ( .A(net84354), .ZN(net84305) );
  NAND2_X4 U3033 ( .A1(net84305), .A2(net84351), .ZN(net84273) );
  NOR2_X1 U3034 ( .A1(net84305), .A2(net84353), .ZN(net84347) );
  NAND2_X2 U3035 ( .A1(net84172), .A2(net84355), .ZN(net84354) );
  INV_X1 U3036 ( .A(u4_exp_out_4_), .ZN(net83596) );
  AOI22_X2 U3037 ( .A1(u4_exp_out_pl1_4_), .A2(net83435), .B1(net83556), .B2(
        u4_exp_out_4_), .ZN(net83555) );
  NAND2_X1 U3038 ( .A1(opa_dn), .A2(net85175), .ZN(net84043) );
  NOR2_X1 U3039 ( .A1(opa_dn), .A2(net85179), .ZN(net83463) );
  MUX2_X2 U3040 ( .A(net95574), .B(net83791), .S(net93455), .Z(net95137) );
  MUX2_X2 U3041 ( .A(net83430), .B(net83791), .S(net93455), .Z(net95136) );
  MUX2_X2 U3042 ( .A(net83510), .B(net83865), .S(net93455), .Z(net83965) );
  INV_X32 U3043 ( .A(net85397), .ZN(net85393) );
  MUX2_X2 U3044 ( .A(u4_exp_next_mi_3_), .B(u4_exp_in_pl1_3_), .S(net85397), 
        .Z(net94004) );
  NAND2_X2 U3045 ( .A1(net84495), .A2(net84400), .ZN(net26607) );
  NOR2_X4 U3046 ( .A1(n2867), .A2(n2868), .ZN(net84236) );
  NAND4_X2 U3047 ( .A1(net84236), .A2(net84239), .A3(net84237), .A4(net84238), 
        .ZN(net95070) );
  AOI211_X4 U3048 ( .C1(n2869), .C2(net84314), .A(net84166), .B(net84257), 
        .ZN(n2868) );
  NAND2_X2 U3049 ( .A1(net17657), .A2(net84258), .ZN(n2869) );
  INV_X2 U3050 ( .A(net17683), .ZN(net84258) );
  NAND4_X4 U3051 ( .A1(net84261), .A2(net84262), .A3(n2870), .A4(n2871), .ZN(
        n2867) );
  NAND2_X2 U3052 ( .A1(n2872), .A2(net28939), .ZN(n2871) );
  INV_X4 U3053 ( .A(n2874), .ZN(n2872) );
  NAND2_X4 U3054 ( .A1(n2872), .A2(net83714), .ZN(net84183) );
  NAND2_X2 U3055 ( .A1(net84324), .A2(net85399), .ZN(n2874) );
  OAI221_X1 U3056 ( .B1(net85393), .B2(net83369), .C1(net83370), .C2(net82931), 
        .A(net83371), .ZN(net83288) );
  NAND2_X4 U3057 ( .A1(u4_exp_next_mi_8_), .A2(net85393), .ZN(net83836) );
  NAND2_X2 U3058 ( .A1(net86045), .A2(net85393), .ZN(net83373) );
  INV_X4 U3059 ( .A(net84397), .ZN(net84495) );
  NAND2_X2 U3060 ( .A1(n2873), .A2(n2490), .ZN(n2870) );
  INV_X1 U3061 ( .A(n2483), .ZN(net84271) );
  INV_X2 U3062 ( .A(net84271), .ZN(net94442) );
  NOR2_X1 U3063 ( .A1(net92690), .A2(net84273), .ZN(n2873) );
  XNOR2_X2 U3064 ( .A(net84118), .B(n2875), .ZN(net82993) );
  AOI211_X4 U3065 ( .C1(net83042), .C2(net94587), .A(net83044), .B(net83043), 
        .ZN(net83038) );
  INV_X2 U3066 ( .A(net83043), .ZN(net92392) );
  NAND2_X1 U3067 ( .A1(net83109), .A2(net83043), .ZN(net83090) );
  INV_X8 U3068 ( .A(net82993), .ZN(u4_ldz_all_2_) );
  NOR2_X4 U3069 ( .A1(n2876), .A2(n2877), .ZN(net84118) );
  OAI21_X4 U3070 ( .B1(net84118), .B2(net84131), .A(net84132), .ZN(net84121)
         );
  XNOR2_X2 U3071 ( .A(net33106), .B(n2654), .ZN(net84116) );
  AOI21_X4 U3072 ( .B1(net33106), .B2(n2654), .A(net84117), .ZN(n2876) );
  NAND2_X2 U3073 ( .A1(net83858), .A2(n2654), .ZN(net83857) );
  INV_X16 U3074 ( .A(net83757), .ZN(net33106) );
  NOR3_X2 U3075 ( .A1(net94966), .A2(net95614), .A3(net82807), .ZN(net83117)
         );
  INV_X16 U3076 ( .A(net83121), .ZN(net85997) );
  NAND3_X4 U3077 ( .A1(n2878), .A2(net83393), .A3(n2686), .ZN(net83121) );
  NAND3_X4 U3078 ( .A1(net83393), .A2(n2882), .A3(n2686), .ZN(net83123) );
  NAND2_X2 U3079 ( .A1(net83356), .A2(opa_00), .ZN(n2883) );
  NOR2_X4 U3080 ( .A1(n2881), .A2(net83357), .ZN(n2880) );
  INV_X4 U3081 ( .A(net83563), .ZN(n2881) );
  NAND2_X2 U3082 ( .A1(n2881), .A2(net83234), .ZN(n2884) );
  OAI21_X4 U3083 ( .B1(net82037), .B2(n2578), .A(n2884), .ZN(n2882) );
  NAND2_X2 U3084 ( .A1(rmode_r3[0]), .A2(n2578), .ZN(net83300) );
  INV_X16 U3085 ( .A(net83123), .ZN(net86013) );
  INV_X4 U3086 ( .A(net83396), .ZN(net82037) );
  OAI21_X1 U3087 ( .B1(net82037), .B2(net95279), .A(net82039), .ZN(net82030)
         );
  AOI22_X4 U3088 ( .A1(n2557), .A2(n2885), .B1(net84201), .B2(n2886), .ZN(
        net84239) );
  INV_X4 U3089 ( .A(net17653), .ZN(net83625) );
  NAND2_X1 U3090 ( .A1(net83624), .A2(net83625), .ZN(net83620) );
  NAND2_X2 U3091 ( .A1(net84361), .A2(net83625), .ZN(net84242) );
  NOR3_X4 U3092 ( .A1(net84242), .A2(n2887), .A3(net17694), .ZN(n2885) );
  INV_X4 U3093 ( .A(net17695), .ZN(n2887) );
  NAND2_X2 U3094 ( .A1(n2887), .A2(net84364), .ZN(net84363) );
  INV_X4 U3095 ( .A(net83635), .ZN(net84361) );
  NOR3_X4 U3096 ( .A1(net83634), .A2(net83635), .A3(net83636), .ZN(net83616)
         );
  INV_X4 U3097 ( .A(net17654), .ZN(net84202) );
  INV_X4 U3098 ( .A(net17692), .ZN(net84362) );
  NAND3_X2 U3099 ( .A1(net84435), .A2(net84436), .A3(n2888), .ZN(net17653) );
  NAND2_X1 U3100 ( .A1(quo[5]), .A2(net86315), .ZN(n2888) );
  INV_X8 U3101 ( .A(n2890), .ZN(net86315) );
  NAND2_X4 U3102 ( .A1(n2889), .A2(net92028), .ZN(n2890) );
  INV_X8 U3103 ( .A(net84451), .ZN(n2889) );
  INV_X16 U3104 ( .A(n2889), .ZN(net86040) );
  AOI22_X2 U3105 ( .A1(u4_div_exp2_0_), .A2(net83751), .B1(u4_div_exp1_0_), 
        .B2(net83752), .ZN(net83745) );
  INV_X4 U3106 ( .A(u4_div_exp2_3_), .ZN(net84002) );
  INV_X4 U3107 ( .A(u4_div_exp2_2_), .ZN(net83977) );
  NAND3_X4 U3108 ( .A1(net84443), .A2(net84444), .A3(n2891), .ZN(net17686) );
  NAND2_X1 U3109 ( .A1(quo[15]), .A2(net86315), .ZN(n2891) );
  NAND2_X4 U3110 ( .A1(net85177), .A2(net93655), .ZN(net84451) );
  INV_X8 U3111 ( .A(net85167), .ZN(net93655) );
  INV_X8 U3112 ( .A(net85179), .ZN(net85177) );
  NOR3_X2 U3113 ( .A1(n3186), .A2(n3069), .A3(n3044), .ZN(n3187) );
  NAND2_X2 U3114 ( .A1(net86497), .A2(u4_fract_out_2_), .ZN(n3854) );
  NAND2_X2 U3115 ( .A1(net86315), .A2(quo[11]), .ZN(n3300) );
  NOR2_X2 U3116 ( .A1(net85145), .A2(net85157), .ZN(n3154) );
  NAND3_X1 U3117 ( .A1(n2585), .A2(n2502), .A3(n3745), .ZN(net83417) );
  NOR2_X2 U3118 ( .A1(net82782), .A2(n4107), .ZN(net82784) );
  INV_X8 U3119 ( .A(n4089), .ZN(n3921) );
  INV_X8 U3120 ( .A(n3779), .ZN(n3843) );
  NAND3_X1 U3121 ( .A1(net83526), .A2(n3741), .A3(n2502), .ZN(net83556) );
  NOR2_X2 U3122 ( .A1(n3692), .A2(n3690), .ZN(net95605) );
  INV_X8 U3123 ( .A(net95605), .ZN(net83431) );
  NAND2_X4 U3124 ( .A1(n3689), .A2(n3695), .ZN(n3690) );
  NAND3_X1 U3125 ( .A1(n3997), .A2(n3996), .A3(net82950), .ZN(n2933) );
  NAND2_X1 U3126 ( .A1(n4060), .A2(n2933), .ZN(n4061) );
  AOI21_X2 U3127 ( .B1(underflow_fmul_r[1]), .B2(n2933), .A(
        underflow_fmul_r[0]), .ZN(n4056) );
  OAI211_X1 U3128 ( .C1(n3789), .C2(n3788), .A(n3787), .B(n3786), .ZN(n3790)
         );
  BUF_X8 U3129 ( .A(net83430), .Z(net95574) );
  INV_X1 U3130 ( .A(fract_denorm[40]), .ZN(n3606) );
  INV_X2 U3131 ( .A(net83498), .ZN(net83497) );
  AOI22_X4 U3132 ( .A1(n2894), .A2(net94595), .B1(n3876), .B2(net86013), .ZN(
        net95549) );
  AND2_X2 U3133 ( .A1(net86497), .A2(u4_fract_out_12_), .ZN(n2894) );
  INV_X4 U3134 ( .A(net85999), .ZN(net94595) );
  NOR2_X1 U3135 ( .A1(net83126), .A2(n3875), .ZN(n3876) );
  INV_X4 U3136 ( .A(n2938), .ZN(n2998) );
  NOR2_X2 U3137 ( .A1(net82782), .A2(n4074), .ZN(n4075) );
  INV_X4 U3138 ( .A(n4035), .ZN(n2897) );
  AND2_X2 U3139 ( .A1(net83446), .A2(net94896), .ZN(net95504) );
  NOR2_X2 U3140 ( .A1(n3391), .A2(n2985), .ZN(n3383) );
  NOR2_X4 U3141 ( .A1(fract_denorm[21]), .A2(fract_denorm[22]), .ZN(net95479)
         );
  AOI22_X4 U3142 ( .A1(u4_N1387), .A2(net85377), .B1(u4_N1437), .B2(n2794), 
        .ZN(n2087) );
  NOR2_X4 U3143 ( .A1(n3259), .A2(net85175), .ZN(n3261) );
  NOR3_X4 U3144 ( .A1(n4032), .A2(n4100), .A3(n2892), .ZN(net83120) );
  NAND2_X2 U3145 ( .A1(n2622), .A2(net84201), .ZN(n2995) );
  INV_X4 U3146 ( .A(n3382), .ZN(n3392) );
  OAI21_X2 U3147 ( .B1(n3403), .B2(n2530), .A(net85393), .ZN(n3404) );
  NAND3_X2 U3148 ( .A1(n2909), .A2(n3350), .A3(n3335), .ZN(net95365) );
  CLKBUF_X2 U3149 ( .A(n3402), .Z(n2899) );
  NAND2_X2 U3150 ( .A1(net84140), .A2(net84141), .ZN(net94614) );
  NAND2_X2 U3151 ( .A1(n2946), .A2(n3399), .ZN(n3424) );
  OAI21_X2 U3152 ( .B1(n3425), .B2(net84185), .A(n3424), .ZN(n3436) );
  NAND3_X2 U3153 ( .A1(n3431), .A2(n2564), .A3(fract_denorm[31]), .ZN(n3432)
         );
  INV_X2 U3154 ( .A(n3397), .ZN(n3401) );
  XNOR2_X2 U3155 ( .A(net94614), .B(n2581), .ZN(u4_ldz_all_0_) );
  CLKBUF_X3 U3156 ( .A(u4_fract_out_0_), .Z(n2900) );
  NAND2_X4 U3157 ( .A1(net83745), .A2(n3598), .ZN(net83736) );
  INV_X4 U3158 ( .A(net85929), .ZN(net91498) );
  INV_X2 U3159 ( .A(u4_fract_out_pl1_21_), .ZN(n3864) );
  INV_X4 U3160 ( .A(net83926), .ZN(net95242) );
  INV_X4 U3161 ( .A(net83868), .ZN(net83926) );
  NOR2_X2 U3162 ( .A1(net83126), .A2(n3855), .ZN(n3856) );
  NOR2_X2 U3163 ( .A1(net83126), .A2(n3849), .ZN(n3850) );
  INV_X2 U3164 ( .A(net82891), .ZN(net95236) );
  INV_X2 U3165 ( .A(n4118), .ZN(n3832) );
  NAND2_X2 U3166 ( .A1(n3895), .A2(u4_fract_out_14_), .ZN(n3888) );
  INV_X16 U3167 ( .A(net86012), .ZN(net83126) );
  OAI21_X2 U3168 ( .B1(net83579), .B2(net83580), .A(n3755), .ZN(n3692) );
  OAI21_X1 U3169 ( .B1(net83487), .B2(net83596), .A(net83527), .ZN(n3687) );
  NOR2_X1 U3170 ( .A1(net83535), .A2(net83596), .ZN(n3679) );
  MUX2_X2 U3171 ( .A(n3471), .B(n3472), .S(net93695), .Z(net95173) );
  NOR2_X2 U3172 ( .A1(n3495), .A2(n3494), .ZN(net84016) );
  INV_X1 U3173 ( .A(u4_ldz_all_6_), .ZN(net95132) );
  INV_X1 U3174 ( .A(net83624), .ZN(net95118) );
  INV_X1 U3175 ( .A(n3471), .ZN(n2905) );
  NAND2_X2 U3176 ( .A1(n3355), .A2(n3444), .ZN(n3358) );
  XNOR2_X2 U3177 ( .A(net84128), .B(n3457), .ZN(n2907) );
  INV_X4 U3178 ( .A(n2907), .ZN(u4_ldz_all_3_) );
  AOI22_X2 U3179 ( .A1(fract_out_q[5]), .A2(n4071), .B1(quo[4]), .B2(n3072), 
        .ZN(n3171) );
  MUX2_X2 U3180 ( .A(n3696), .B(n3474), .S(net93695), .Z(n3493) );
  INV_X4 U3181 ( .A(net84273), .ZN(net84350) );
  NOR2_X4 U3182 ( .A1(net17683), .A2(net17657), .ZN(n2909) );
  INV_X4 U3183 ( .A(n2909), .ZN(n3663) );
  NAND3_X1 U3184 ( .A1(net83713), .A2(net83714), .A3(net83715), .ZN(n3614) );
  OAI22_X4 U3185 ( .A1(net86001), .A2(n2912), .B1(n2913), .B2(net86014), .ZN(
        net94966) );
  INV_X8 U3186 ( .A(n4082), .ZN(n4035) );
  NAND4_X1 U3187 ( .A1(n3954), .A2(n3953), .A3(n3952), .A4(n3951), .ZN(n2911)
         );
  NOR2_X2 U3188 ( .A1(net86401), .A2(n4118), .ZN(n3953) );
  INV_X4 U3189 ( .A(net94966), .ZN(net86418) );
  CLKBUF_X3 U3190 ( .A(n3422), .Z(n2959) );
  INV_X4 U3191 ( .A(net83507), .ZN(net94948) );
  AOI22_X2 U3192 ( .A1(u4_exp_fix_diva[1]), .A2(net83312), .B1(
        u4_exp_fix_divb[1]), .B2(net95605), .ZN(n3739) );
  NAND2_X4 U3193 ( .A1(n3947), .A2(net95473), .ZN(n3527) );
  NOR2_X1 U3194 ( .A1(n3091), .A2(net85905), .ZN(n2914) );
  BUF_X32 U3195 ( .A(u4_ldz_all_1_), .Z(n2915) );
  INV_X4 U3196 ( .A(n2916), .ZN(n2917) );
  INV_X16 U3197 ( .A(net86040), .ZN(net84605) );
  INV_X4 U3198 ( .A(net95070), .ZN(net84141) );
  INV_X1 U3199 ( .A(u4_ldz_all_3_), .ZN(n2918) );
  INV_X2 U3200 ( .A(n2918), .ZN(n2919) );
  NAND2_X1 U3201 ( .A1(net83525), .A2(net94896), .ZN(n3728) );
  NOR3_X2 U3202 ( .A1(n3958), .A2(n3957), .A3(n3956), .ZN(n3960) );
  INV_X4 U3203 ( .A(n2920), .ZN(n2921) );
  INV_X4 U3204 ( .A(n2922), .ZN(n2923) );
  XNOR2_X2 U3205 ( .A(n3452), .B(n3455), .ZN(n2924) );
  NOR2_X1 U3206 ( .A1(n2914), .A2(n3479), .ZN(n2925) );
  INV_X1 U3207 ( .A(u4_ldz_all_2_), .ZN(net94834) );
  INV_X2 U3208 ( .A(u6_N8), .ZN(n4592) );
  OR3_X1 U3209 ( .A1(u6_N8), .A2(u6_N9), .A3(u6_N7), .ZN(n1753) );
  MUX2_X2 U3210 ( .A(n3474), .B(n3696), .S(net85393), .Z(n2926) );
  INV_X1 U3211 ( .A(n4071), .ZN(n2927) );
  BUF_X32 U3212 ( .A(n3955), .Z(n2928) );
  INV_X2 U3213 ( .A(n2929), .ZN(net94811) );
  AND2_X2 U3214 ( .A1(net83041), .A2(net83928), .ZN(n2929) );
  NOR3_X4 U3215 ( .A1(n2628), .A2(net85111), .A3(net85135), .ZN(n3266) );
  BUF_X32 U3216 ( .A(u6_N23), .Z(n2930) );
  INV_X2 U3217 ( .A(net82965), .ZN(net94725) );
  INV_X2 U3218 ( .A(u4_N1733), .ZN(net82965) );
  OAI21_X2 U3219 ( .B1(net83567), .B2(net83568), .A(net82040), .ZN(n3700) );
  INV_X4 U3220 ( .A(n2931), .ZN(n3804) );
  AOI21_X2 U3221 ( .B1(n2931), .B2(u4_exp_out_pl1_0_), .A(n3806), .ZN(n3811)
         );
  NOR3_X2 U3222 ( .A1(net83357), .A2(net83562), .A3(net83563), .ZN(n2931) );
  INV_X1 U3223 ( .A(net82893), .ZN(net94701) );
  INV_X1 U3224 ( .A(n2460), .ZN(n2932) );
  NOR2_X4 U3225 ( .A1(n4122), .A2(n4121), .ZN(n3952) );
  NOR2_X1 U3226 ( .A1(net82782), .A2(net94701), .ZN(n4091) );
  NOR2_X1 U3227 ( .A1(net82782), .A2(n2932), .ZN(n4077) );
  INV_X2 U3228 ( .A(net83562), .ZN(net94692) );
  NOR2_X2 U3229 ( .A1(net82782), .A2(net95236), .ZN(n4092) );
  BUF_X32 U3230 ( .A(u4_exp_next_mi_2_), .Z(n2934) );
  INV_X16 U3231 ( .A(n3517), .ZN(n2935) );
  INV_X32 U3232 ( .A(n2935), .ZN(n2936) );
  INV_X4 U3233 ( .A(n3139), .ZN(n3517) );
  INV_X1 U3234 ( .A(n3021), .ZN(n2937) );
  AOI22_X4 U3235 ( .A1(net94595), .A2(n2939), .B1(n2940), .B2(net86013), .ZN(
        n2938) );
  AND2_X2 U3236 ( .A1(net95019), .A2(u4_fract_out_6_), .ZN(n2939) );
  NOR2_X1 U3237 ( .A1(net83126), .A2(n3877), .ZN(n2940) );
  INV_X2 U3238 ( .A(net82918), .ZN(net94587) );
  INV_X2 U3239 ( .A(net95525), .ZN(net82918) );
  INV_X2 U3240 ( .A(net93776), .ZN(net94146) );
  INV_X4 U3241 ( .A(n2941), .ZN(n2942) );
  INV_X4 U3242 ( .A(n2943), .ZN(n2944) );
  NAND2_X4 U3243 ( .A1(net82856), .A2(n3764), .ZN(net83750) );
  NOR2_X4 U3244 ( .A1(n3213), .A2(net85175), .ZN(n3215) );
  NOR2_X2 U3245 ( .A1(n2547), .A2(n3612), .ZN(n3348) );
  INV_X8 U3246 ( .A(fract_denorm[31]), .ZN(n3338) );
  AOI21_X4 U3247 ( .B1(n3267), .B2(net92028), .A(n3266), .ZN(n3268) );
  INV_X4 U3248 ( .A(n3897), .ZN(n3898) );
  NAND2_X2 U3249 ( .A1(net92392), .A2(n2742), .ZN(n3916) );
  NAND2_X4 U3250 ( .A1(n2645), .A2(n3773), .ZN(net83262) );
  NAND2_X1 U3251 ( .A1(net83041), .A2(n3646), .ZN(n3660) );
  NAND3_X2 U3252 ( .A1(n2477), .A2(n3659), .A3(n2901), .ZN(n4001) );
  NAND2_X1 U3253 ( .A1(net83433), .A2(net85933), .ZN(n3775) );
  NOR3_X2 U3254 ( .A1(n3772), .A2(n3771), .A3(n3770), .ZN(n3774) );
  INV_X2 U3255 ( .A(net94373), .ZN(net94374) );
  NAND2_X2 U3256 ( .A1(n3398), .A2(net84377), .ZN(n2945) );
  INV_X2 U3257 ( .A(n2945), .ZN(n2946) );
  NAND3_X2 U3258 ( .A1(net23043), .A2(net83762), .A3(net84139), .ZN(n3449) );
  INV_X4 U3259 ( .A(n3388), .ZN(n3371) );
  NOR2_X4 U3260 ( .A1(n3008), .A2(n3006), .ZN(n3369) );
  INV_X16 U3261 ( .A(n3007), .ZN(n3008) );
  NAND4_X2 U3262 ( .A1(n3954), .A2(n3953), .A3(n3952), .A4(n3951), .ZN(n4067)
         );
  NAND3_X2 U3263 ( .A1(net84376), .A2(net83630), .A3(net84377), .ZN(net84375)
         );
  NAND2_X4 U3264 ( .A1(n3423), .A2(net84188), .ZN(net83630) );
  NAND2_X2 U3265 ( .A1(u4_fract_out_22_), .A2(net86497), .ZN(n3867) );
  NAND4_X2 U3266 ( .A1(quo[40]), .A2(net85175), .A3(net92028), .A4(net85159), 
        .ZN(n3263) );
  NAND2_X4 U3267 ( .A1(net85135), .A2(net85159), .ZN(n3259) );
  INV_X1 U3268 ( .A(n2465), .ZN(net83342) );
  INV_X16 U3269 ( .A(net85997), .ZN(net85999) );
  NOR2_X2 U3270 ( .A1(n2464), .A2(n3927), .ZN(n3928) );
  NOR2_X2 U3271 ( .A1(net85115), .A2(net85139), .ZN(n3199) );
  INV_X4 U3272 ( .A(n3892), .ZN(n3893) );
  NOR3_X2 U3273 ( .A1(n4033), .A2(net94966), .A3(n2896), .ZN(n4042) );
  INV_X8 U3274 ( .A(n4029), .ZN(n3869) );
  NAND2_X4 U3275 ( .A1(n3929), .A2(n3928), .ZN(net83059) );
  NAND2_X2 U3276 ( .A1(net92028), .A2(net85159), .ZN(n3274) );
  NOR3_X4 U3277 ( .A1(n4015), .A2(n2927), .A3(net82767), .ZN(n4021) );
  NAND3_X4 U3278 ( .A1(n2910), .A2(net83278), .A3(net83276), .ZN(net83393) );
  NOR2_X1 U3279 ( .A1(net83282), .A2(n3828), .ZN(net83264) );
  NOR2_X2 U3280 ( .A1(n3926), .A2(n3020), .ZN(n3929) );
  NAND2_X2 U3281 ( .A1(n4058), .A2(n2746), .ZN(n4062) );
  OAI22_X4 U3282 ( .A1(n2640), .A2(net86014), .B1(net85999), .B2(n3854), .ZN(
        n4076) );
  NOR2_X1 U3283 ( .A1(net82782), .A2(n2479), .ZN(n4104) );
  INV_X4 U3284 ( .A(n4020), .ZN(n4015) );
  AOI22_X4 U3285 ( .A1(u4_N1384), .A2(net85377), .B1(u4_N1434), .B2(n2794), 
        .ZN(n2091) );
  MUX2_X2 U3286 ( .A(u4_exp_next_mi_2_), .B(u4_exp_in_pl1_2_), .S(net93695), 
        .Z(n2948) );
  INV_X4 U3287 ( .A(n2948), .ZN(n3509) );
  INV_X2 U3288 ( .A(n2934), .ZN(n3708) );
  INV_X2 U3289 ( .A(u4_exp_in_pl1_2_), .ZN(n3558) );
  NAND2_X4 U3290 ( .A1(n3375), .A2(n3360), .ZN(net84312) );
  NOR3_X4 U3291 ( .A1(n2629), .A2(net85111), .A3(net85135), .ZN(n3247) );
  NAND2_X1 U3292 ( .A1(net83383), .A2(net95138), .ZN(net82931) );
  OR2_X1 U3293 ( .A1(n2929), .A2(net82931), .ZN(n2949) );
  NAND2_X2 U3294 ( .A1(n4009), .A2(net86027), .ZN(n2951) );
  NAND2_X4 U3295 ( .A1(n2950), .A2(n2951), .ZN(n4115) );
  OAI21_X2 U3296 ( .B1(n2545), .B2(n2974), .A(n3388), .ZN(n3390) );
  NOR3_X4 U3297 ( .A1(n2630), .A2(net92028), .A3(net85111), .ZN(n3239) );
  NAND2_X4 U3298 ( .A1(n2983), .A2(n3509), .ZN(n3473) );
  INV_X1 U3299 ( .A(u6_N15), .ZN(n4504) );
  INV_X4 U3300 ( .A(net94004), .ZN(net84000) );
  NAND3_X2 U3301 ( .A1(n2938), .A2(net82893), .A3(n2898), .ZN(n3926) );
  INV_X1 U3302 ( .A(n3402), .ZN(n3408) );
  INV_X8 U3303 ( .A(n3715), .ZN(n3807) );
  INV_X1 U3304 ( .A(net33106), .ZN(net93902) );
  NOR3_X4 U3305 ( .A1(n2897), .A2(n4038), .A3(n2997), .ZN(net83198) );
  INV_X4 U3306 ( .A(n2956), .ZN(n2957) );
  NOR2_X1 U3307 ( .A1(net82782), .A2(n4095), .ZN(n4096) );
  NOR3_X1 U3308 ( .A1(n2729), .A2(u4_ldz_all_5_), .A3(net82997), .ZN(n3977) );
  INV_X1 U3309 ( .A(n3091), .ZN(n3734) );
  INV_X4 U3310 ( .A(net84135), .ZN(net93776) );
  NAND2_X2 U3311 ( .A1(n3354), .A2(net84201), .ZN(n3444) );
  NOR3_X4 U3312 ( .A1(n3800), .A2(n3820), .A3(n3799), .ZN(n3814) );
  AOI22_X1 U3313 ( .A1(net22501), .A2(net23097), .B1(net23104), .B2(net48876), 
        .ZN(n1416) );
  NOR2_X4 U3314 ( .A1(n3677), .A2(n2603), .ZN(net93714) );
  NOR2_X2 U3315 ( .A1(net83316), .A2(n3708), .ZN(n3711) );
  INV_X4 U3316 ( .A(n3452), .ZN(n3456) );
  NAND2_X2 U3317 ( .A1(net84124), .A2(net83761), .ZN(n2965) );
  NOR2_X1 U3318 ( .A1(net83636), .A2(net83622), .ZN(n2960) );
  NOR2_X4 U3319 ( .A1(n3419), .A2(n2961), .ZN(n3384) );
  INV_X4 U3320 ( .A(n2960), .ZN(n2961) );
  OAI221_X2 U3321 ( .B1(n3513), .B2(net83750), .C1(net83977), .C2(net83753), 
        .A(n3512), .ZN(net83017) );
  NOR2_X2 U3322 ( .A1(div_opa_ldz_r2[2]), .A2(net83754), .ZN(net84131) );
  MUX2_X2 U3323 ( .A(u4_exp_next_mi_7_), .B(u4_exp_in_pl1_7_), .S(net93695), 
        .Z(net93671) );
  NAND3_X2 U3324 ( .A1(n3170), .A2(n3169), .A3(n3168), .ZN(fract_denorm[23])
         );
  INV_X1 U3325 ( .A(n2925), .ZN(n3138) );
  NAND2_X2 U3326 ( .A1(net84151), .A2(n3444), .ZN(n3412) );
  NOR3_X2 U3327 ( .A1(net85139), .A2(net85111), .A3(n2646), .ZN(n3181) );
  NAND2_X4 U3328 ( .A1(n3693), .A2(n3692), .ZN(net83428) );
  INV_X4 U3329 ( .A(n2680), .ZN(n2962) );
  INV_X1 U3330 ( .A(n2680), .ZN(n2963) );
  INV_X2 U3331 ( .A(u4_ldz_all_0_), .ZN(n3969) );
  NOR2_X2 U3332 ( .A1(net83126), .A2(n3891), .ZN(n3892) );
  INV_X4 U3333 ( .A(n3879), .ZN(n3880) );
  NOR2_X4 U3334 ( .A1(net83126), .A2(n3878), .ZN(n3879) );
  INV_X4 U3335 ( .A(n4105), .ZN(n4027) );
  NOR2_X2 U3336 ( .A1(n4105), .A2(n4107), .ZN(n3019) );
  INV_X8 U3337 ( .A(n4087), .ZN(n3917) );
  NAND2_X2 U3338 ( .A1(net83636), .A2(net84205), .ZN(n3353) );
  NAND2_X4 U3339 ( .A1(net93507), .A2(net83773), .ZN(n2966) );
  NAND2_X4 U3340 ( .A1(n2965), .A2(n2966), .ZN(u4_ldz_all_5_) );
  INV_X4 U3341 ( .A(net84124), .ZN(net93507) );
  NAND3_X2 U3342 ( .A1(n3380), .A2(n3398), .A3(n3379), .ZN(net83761) );
  AOI21_X1 U3343 ( .B1(n3948), .B2(n3947), .A(net83030), .ZN(n3949) );
  NOR2_X4 U3344 ( .A1(n4109), .A2(n2635), .ZN(n3160) );
  NOR2_X2 U3345 ( .A1(n2691), .A2(net83864), .ZN(n3559) );
  NOR2_X2 U3346 ( .A1(n2694), .A2(net83864), .ZN(n3551) );
  NOR2_X2 U3347 ( .A1(n2688), .A2(net83864), .ZN(n3542) );
  AOI21_X1 U3348 ( .B1(n3533), .B2(n3581), .A(net83811), .ZN(n3535) );
  AOI211_X1 U3349 ( .C1(net83854), .C2(n3561), .A(n3560), .B(n3559), .ZN(n3567) );
  NOR3_X2 U3350 ( .A1(net83921), .A2(n3535), .A3(n3534), .ZN(n3536) );
  NOR2_X2 U3351 ( .A1(n4103), .A2(n4101), .ZN(n3870) );
  INV_X1 U3352 ( .A(u6_N10), .ZN(n4509) );
  NAND3_X2 U3353 ( .A1(n4015), .A2(net82918), .A3(n2743), .ZN(n4018) );
  INV_X2 U3354 ( .A(u4_exp_next_mi_8_), .ZN(net83948) );
  INV_X8 U3355 ( .A(net84067), .ZN(net83771) );
  NAND2_X1 U3356 ( .A1(n3562), .A2(net83823), .ZN(n3582) );
  NOR2_X1 U3357 ( .A1(net83823), .A2(n3558), .ZN(n3560) );
  NAND3_X1 U3358 ( .A1(n3170), .A2(n3169), .A3(n3168), .ZN(n3067) );
  CLKBUF_X3 U3359 ( .A(n2557), .Z(net93422) );
  NAND2_X1 U3360 ( .A1(prod[14]), .A2(n2936), .ZN(n3311) );
  NAND2_X2 U3361 ( .A1(prod[11]), .A2(n2936), .ZN(n3308) );
  NAND2_X1 U3362 ( .A1(prod[6]), .A2(n2936), .ZN(n3326) );
  NAND2_X1 U3363 ( .A1(prod[5]), .A2(n2936), .ZN(n3323) );
  NOR2_X1 U3364 ( .A1(n4110), .A2(net82776), .ZN(n4111) );
  NOR2_X1 U3365 ( .A1(opa_00), .A2(net82776), .ZN(n4017) );
  NOR2_X1 U3366 ( .A1(net82776), .A2(n3943), .ZN(n3946) );
  OAI21_X1 U3367 ( .B1(net82776), .B2(n3944), .A(net83070), .ZN(n3839) );
  NOR2_X1 U3368 ( .A1(net82776), .A2(net83865), .ZN(n3569) );
  NAND3_X2 U3369 ( .A1(n3442), .A2(n3441), .A3(n3440), .ZN(net17652) );
  NAND3_X2 U3370 ( .A1(n3329), .A2(n3328), .A3(n3327), .ZN(net17695) );
  NAND3_X2 U3371 ( .A1(n3332), .A2(n3331), .A3(n3330), .ZN(net17694) );
  NAND3_X2 U3372 ( .A1(n3320), .A2(n3319), .A3(n3318), .ZN(net17693) );
  NAND3_X2 U3373 ( .A1(n3323), .A2(n3322), .A3(n3321), .ZN(net17692) );
  INV_X2 U3374 ( .A(net83713), .ZN(net93404) );
  INV_X2 U3375 ( .A(n3384), .ZN(n3364) );
  NOR3_X4 U3376 ( .A1(n2631), .A2(net92028), .A3(net85111), .ZN(n3230) );
  XNOR2_X1 U3377 ( .A(n3460), .B(net91498), .ZN(net83941) );
  INV_X4 U3378 ( .A(net85165), .ZN(net93364) );
  NOR2_X4 U3379 ( .A1(n3046), .A2(n3243), .ZN(net84559) );
  AOI22_X4 U3380 ( .A1(u4_N1385), .A2(net23182), .B1(u4_N1435), .B2(n2794), 
        .ZN(n1454) );
  AOI21_X2 U3381 ( .B1(net84182), .B2(n2955), .A(n3376), .ZN(n3366) );
  INV_X4 U3382 ( .A(net83759), .ZN(net86531) );
  INV_X16 U3383 ( .A(net86531), .ZN(net86532) );
  NAND3_X2 U3384 ( .A1(net85165), .A2(net85133), .A3(prod[21]), .ZN(n3197) );
  NAND2_X4 U3385 ( .A1(n3350), .A2(net83622), .ZN(n3409) );
  NAND3_X2 U3386 ( .A1(net83762), .A2(net84139), .A3(net23043), .ZN(net93218)
         );
  INV_X2 U3387 ( .A(u4_div_exp1_7_), .ZN(net83381) );
  NAND2_X1 U3388 ( .A1(n3381), .A2(net83761), .ZN(u4_fi_ldz_2a_6_) );
  NAND2_X1 U3389 ( .A1(net83761), .A2(n3381), .ZN(u4_fi_ldz_2a_5_) );
  AOI21_X1 U3390 ( .B1(net83846), .B2(n3091), .A(n3577), .ZN(n3578) );
  XOR2_X1 U3391 ( .A(n3089), .B(n3091), .Z(n3514) );
  XOR2_X1 U3392 ( .A(div_opa_ldz_r2[1]), .B(n3091), .Z(n3570) );
  NAND2_X1 U3393 ( .A1(n3091), .A2(n3089), .ZN(n3503) );
  INV_X4 U3394 ( .A(n2679), .ZN(n2967) );
  INV_X1 U3395 ( .A(n2679), .ZN(n2968) );
  INV_X16 U3396 ( .A(n3090), .ZN(n3091) );
  INV_X1 U3397 ( .A(fract_denorm[45]), .ZN(net84181) );
  AND2_X4 U3398 ( .A1(n3063), .A2(n3064), .ZN(n3097) );
  NOR3_X2 U3399 ( .A1(n3447), .A2(n3446), .A3(n3445), .ZN(net84143) );
  AOI22_X4 U3400 ( .A1(n1371), .A2(n2929), .B1(net86027), .B2(net83016), .ZN(
        n3518) );
  AOI21_X2 U3401 ( .B1(u4_exp_out_pl1_1_), .B2(net83435), .A(n3735), .ZN(n3740) );
  NOR3_X2 U3402 ( .A1(n4037), .A2(n4085), .A3(n2466), .ZN(n4041) );
  NOR2_X4 U3403 ( .A1(net84347), .A2(net84348), .ZN(n3357) );
  AOI22_X4 U3404 ( .A1(u4_N1386), .A2(net23182), .B1(u4_N1436), .B2(n2794), 
        .ZN(n1453) );
  INV_X2 U3405 ( .A(u6_N9), .ZN(n4597) );
  NAND2_X4 U3406 ( .A1(n4758), .A2(div_opa_ldz_r2[0]), .ZN(net84117) );
  INV_X4 U3407 ( .A(n2770), .ZN(n2969) );
  INV_X8 U3408 ( .A(n2771), .ZN(n2986) );
  NAND2_X1 U3409 ( .A1(fract_i2f[3]), .A2(net85115), .ZN(net84436) );
  INV_X8 U3410 ( .A(n2772), .ZN(n2982) );
  NAND2_X2 U3411 ( .A1(n2667), .A2(n3740), .ZN(n2971) );
  INV_X4 U3412 ( .A(n2971), .ZN(n2972) );
  NAND2_X4 U3413 ( .A1(n3843), .A2(n3054), .ZN(net83074) );
  INV_X2 U3414 ( .A(n2974), .ZN(n2973) );
  INV_X2 U3415 ( .A(n3345), .ZN(n3346) );
  INV_X8 U3416 ( .A(n3411), .ZN(n3398) );
  NAND3_X2 U3417 ( .A1(net85165), .A2(net85133), .A3(prod[22]), .ZN(n3203) );
  NAND3_X2 U3418 ( .A1(n3273), .A2(n3272), .A3(n3271), .ZN(n3278) );
  NAND3_X2 U3419 ( .A1(prod[20]), .A2(net85165), .A3(net85131), .ZN(n3192) );
  INV_X1 U3420 ( .A(n3375), .ZN(n2974) );
  NOR2_X2 U3421 ( .A1(n3846), .A2(net83066), .ZN(n3848) );
  NAND2_X4 U3422 ( .A1(n3051), .A2(n3918), .ZN(n4038) );
  NAND2_X1 U3423 ( .A1(n2925), .A2(n3088), .ZN(n3461) );
  NAND2_X1 U3424 ( .A1(n2914), .A2(n3479), .ZN(n3137) );
  XNOR2_X1 U3425 ( .A(n3087), .B(n2925), .ZN(n3463) );
  INV_X1 U3426 ( .A(n2914), .ZN(n3961) );
  INV_X4 U3427 ( .A(n4059), .ZN(n4013) );
  NOR2_X1 U3428 ( .A1(fract_denorm[27]), .A2(n3373), .ZN(n3374) );
  NAND2_X1 U3429 ( .A1(net82753), .A2(n4118), .ZN(N471) );
  NOR3_X4 U3430 ( .A1(n2998), .A2(n4085), .A3(n4036), .ZN(net83119) );
  INV_X4 U3431 ( .A(net84323), .ZN(net83713) );
  NOR2_X4 U3432 ( .A1(net17659), .A2(net17682), .ZN(n3335) );
  NOR2_X4 U3433 ( .A1(fract_denorm[35]), .A2(fract_denorm[36]), .ZN(n2975) );
  NOR2_X1 U3434 ( .A1(n3970), .A2(n2919), .ZN(n3971) );
  NAND2_X2 U3435 ( .A1(quo[39]), .A2(net94019), .ZN(n3265) );
  NAND2_X2 U3436 ( .A1(net83757), .A2(n4758), .ZN(net84083) );
  NOR2_X1 U3437 ( .A1(net84323), .A2(net84272), .ZN(net92895) );
  NAND2_X1 U3438 ( .A1(u4_exp_out_2_), .A2(net94948), .ZN(n3713) );
  NOR2_X2 U3439 ( .A1(fract_denorm[26]), .A2(fract_denorm[27]), .ZN(n3009) );
  NOR2_X2 U3440 ( .A1(n3974), .A2(n3973), .ZN(n3976) );
  NAND2_X1 U3441 ( .A1(n3027), .A2(net92781), .ZN(n2977) );
  NAND2_X4 U3442 ( .A1(n3458), .A2(net85937), .ZN(n2978) );
  NAND2_X4 U3443 ( .A1(n2977), .A2(n2978), .ZN(n3459) );
  INV_X1 U3444 ( .A(net85937), .ZN(net92781) );
  INV_X2 U3445 ( .A(n2548), .ZN(n2979) );
  NAND3_X2 U3446 ( .A1(n3302), .A2(n3301), .A3(n3300), .ZN(n2980) );
  NAND3_X2 U3447 ( .A1(n3302), .A2(n3301), .A3(n3300), .ZN(n2981) );
  NAND3_X2 U3448 ( .A1(n3302), .A2(n3301), .A3(n3300), .ZN(n5325) );
  NOR2_X4 U3449 ( .A1(n3333), .A2(n3612), .ZN(net91817) );
  NOR2_X4 U3450 ( .A1(net83963), .A2(n3599), .ZN(n2983) );
  NOR3_X4 U3451 ( .A1(n3664), .A2(net83630), .A3(n3663), .ZN(n3669) );
  INV_X1 U3452 ( .A(n2672), .ZN(n4502) );
  NAND3_X2 U3453 ( .A1(n3383), .A2(n2571), .A3(n3392), .ZN(net84284) );
  INV_X1 U3454 ( .A(n3666), .ZN(n2984) );
  INV_X4 U3455 ( .A(n2984), .ZN(n2985) );
  INV_X8 U3456 ( .A(n5326), .ZN(n3666) );
  INV_X8 U3457 ( .A(net17655), .ZN(net83624) );
  NOR2_X1 U3458 ( .A1(net82782), .A2(net94966), .ZN(n4094) );
  NAND2_X2 U3459 ( .A1(n3386), .A2(n3422), .ZN(n3387) );
  INV_X4 U3460 ( .A(net84272), .ZN(net84385) );
  INV_X1 U3461 ( .A(n2982), .ZN(n4511) );
  INV_X1 U3462 ( .A(net83527), .ZN(net83534) );
  INV_X1 U3463 ( .A(n2986), .ZN(n4607) );
  AND2_X4 U3464 ( .A1(n3058), .A2(n3059), .ZN(n3099) );
  INV_X1 U3465 ( .A(n2915), .ZN(n3968) );
  INV_X4 U3466 ( .A(u4_exp_next_mi_6_), .ZN(net83430) );
  OAI21_X2 U3467 ( .B1(n2469), .B2(net94146), .A(u4_fi_ldz_2a_3_), .ZN(n3448)
         );
  NAND2_X4 U3468 ( .A1(n2990), .A2(net92624), .ZN(n3773) );
  INV_X1 U3469 ( .A(n2514), .ZN(n2991) );
  INV_X2 U3470 ( .A(n2991), .ZN(n2992) );
  NOR3_X2 U3471 ( .A1(u4_N1420), .A2(u4_N1421), .A3(u4_N1422), .ZN(n3651) );
  AOI211_X2 U3472 ( .C1(n4097), .C2(net85988), .A(net82757), .B(net85976), 
        .ZN(N460) );
  INV_X2 U3473 ( .A(net84376), .ZN(net92599) );
  INV_X2 U3474 ( .A(net84191), .ZN(net84376) );
  NAND3_X4 U3475 ( .A1(quo[1]), .A2(net85133), .A3(n3284), .ZN(n3200) );
  NAND3_X2 U3476 ( .A1(net84370), .A2(n3349), .A3(net83713), .ZN(net84166) );
  NOR2_X2 U3477 ( .A1(net84231), .A2(net84166), .ZN(n3399) );
  NOR3_X1 U3478 ( .A1(fract_denorm[27]), .A2(fract_denorm[25]), .A3(
        fract_denorm[26]), .ZN(n3347) );
  AOI22_X4 U3479 ( .A1(fract_i2f[25]), .A2(net85115), .B1(prod[25]), .B2(n2936), .ZN(n3173) );
  NAND2_X1 U3480 ( .A1(n2936), .A2(net85121), .ZN(net82776) );
  NAND2_X1 U3481 ( .A1(prod[0]), .A2(n2936), .ZN(n3442) );
  NAND2_X1 U3482 ( .A1(prod[1]), .A2(n2936), .ZN(n3329) );
  NAND2_X1 U3483 ( .A1(prod[2]), .A2(n2936), .ZN(n3332) );
  NAND2_X1 U3484 ( .A1(prod[3]), .A2(n2936), .ZN(net84435) );
  NAND2_X1 U3485 ( .A1(prod[4]), .A2(n2936), .ZN(n3320) );
  NAND2_X1 U3486 ( .A1(prod[13]), .A2(n2936), .ZN(net84443) );
  NAND2_X2 U3487 ( .A1(prod[12]), .A2(n2936), .ZN(n3305) );
  INV_X4 U3488 ( .A(fract_denorm[23]), .ZN(net83638) );
  NAND2_X2 U3489 ( .A1(net83500), .A2(u4_fract_out_pl1_23_), .ZN(n2993) );
  NAND2_X4 U3490 ( .A1(net83499), .A2(n2994), .ZN(net83518) );
  INV_X4 U3491 ( .A(n2993), .ZN(n2994) );
  NAND3_X4 U3492 ( .A1(net84370), .A2(n3349), .A3(net83713), .ZN(net92573) );
  NOR2_X2 U3493 ( .A1(net83126), .A2(n3871), .ZN(n3872) );
  NAND2_X2 U3494 ( .A1(net86027), .A2(net83932), .ZN(n3532) );
  NAND2_X2 U3495 ( .A1(net86045), .A2(u4_N1733), .ZN(n3526) );
  INV_X1 U3496 ( .A(net94896), .ZN(net83535) );
  NAND3_X2 U3497 ( .A1(n3348), .A2(n3369), .A3(n3347), .ZN(n3362) );
  AND2_X2 U3498 ( .A1(n3417), .A2(n2995), .ZN(n3439) );
  NAND3_X2 U3499 ( .A1(quo[34]), .A2(net84605), .A3(net85133), .ZN(n3227) );
  INV_X4 U3500 ( .A(net86040), .ZN(net84455) );
  NOR2_X1 U3501 ( .A1(net85901), .A2(net82965), .ZN(n3988) );
  OAI21_X1 U3502 ( .B1(net82036), .B2(net82965), .A(net83358), .ZN(n3525) );
  NOR2_X4 U3503 ( .A1(n3025), .A2(n3026), .ZN(n3046) );
  NAND2_X2 U3504 ( .A1(net86295), .A2(fpu_op_r3_1_), .ZN(n3025) );
  NOR2_X4 U3505 ( .A1(u4_N1733), .A2(n3531), .ZN(net83932) );
  AND2_X2 U3506 ( .A1(n2996), .A2(n3060), .ZN(n3096) );
  NOR3_X2 U3507 ( .A1(n4031), .A2(n4030), .A3(n4029), .ZN(n4043) );
  NAND2_X4 U3508 ( .A1(n3868), .A2(n3919), .ZN(n4029) );
  INV_X4 U3509 ( .A(n2999), .ZN(n3000) );
  NAND3_X2 U3510 ( .A1(net83068), .A2(n3844), .A3(net83220), .ZN(n3845) );
  NAND3_X2 U3511 ( .A1(n4011), .A2(n4013), .A3(n4012), .ZN(n4020) );
  INV_X1 U3512 ( .A(n3921), .ZN(n3001) );
  NOR2_X2 U3513 ( .A1(net82782), .A2(n4105), .ZN(n4106) );
  NAND3_X1 U3514 ( .A1(n4026), .A2(n4025), .A3(n4024), .ZN(n4031) );
  INV_X4 U3515 ( .A(n3872), .ZN(n3874) );
  INV_X4 U3516 ( .A(n3002), .ZN(n3003) );
  AOI21_X1 U3517 ( .B1(n4055), .B2(n4054), .A(net82856), .ZN(net82853) );
  NAND4_X1 U3518 ( .A1(net92028), .A2(net85159), .A3(net85179), .A4(quo[8]), 
        .ZN(n3188) );
  NOR2_X1 U3519 ( .A1(net86309), .A2(n4113), .ZN(n4060) );
  NAND2_X4 U3520 ( .A1(n2638), .A2(n3183), .ZN(fract_denorm[30]) );
  NAND4_X1 U3521 ( .A1(fpu_op_r3_1_), .A2(net85159), .A3(net85179), .A4(quo[9]), .ZN(n3184) );
  NOR3_X2 U3522 ( .A1(n3182), .A2(n2623), .A3(n3181), .ZN(n3183) );
  INV_X16 U3523 ( .A(n3479), .ZN(n3089) );
  INV_X8 U3524 ( .A(fract_denorm[38]), .ZN(net84172) );
  INV_X1 U3525 ( .A(n2551), .ZN(n3607) );
  NAND2_X2 U3526 ( .A1(quo[3]), .A2(n3072), .ZN(n3163) );
  NOR2_X2 U3527 ( .A1(net86040), .A2(n3158), .ZN(n3159) );
  NOR2_X1 U3528 ( .A1(net90897), .A2(net85159), .ZN(n3219) );
  NOR2_X1 U3529 ( .A1(net82782), .A2(n4100), .ZN(net82792) );
  NOR2_X1 U3530 ( .A1(net82782), .A2(net94976), .ZN(n4093) );
  NAND2_X4 U3531 ( .A1(n3661), .A2(n3662), .ZN(net83606) );
  NAND2_X2 U3532 ( .A1(net86497), .A2(u4_fract_out_8_), .ZN(n3881) );
  NAND2_X2 U3533 ( .A1(net86497), .A2(n2900), .ZN(n3778) );
  INV_X4 U3534 ( .A(n3004), .ZN(n3005) );
  NOR2_X1 U3535 ( .A1(net82782), .A2(n2895), .ZN(n4088) );
  OAI211_X2 U3536 ( .C1(n4057), .C2(n2762), .A(net82850), .B(n4056), .ZN(n4058) );
  NAND2_X2 U3537 ( .A1(net86497), .A2(u4_fract_out_16_), .ZN(n3899) );
  NOR3_X4 U3538 ( .A1(n2632), .A2(net92028), .A3(net85111), .ZN(n3234) );
  NAND2_X2 U3539 ( .A1(net85149), .A2(net85167), .ZN(n3139) );
  INV_X8 U3540 ( .A(n3428), .ZN(n3006) );
  INV_X4 U3541 ( .A(net84293), .ZN(net84348) );
  NAND2_X4 U3542 ( .A1(net84324), .A2(net84385), .ZN(net84353) );
  INV_X8 U3543 ( .A(fract_denorm[30]), .ZN(n3007) );
  CLKBUF_X2 U3544 ( .A(n3606), .Z(n3029) );
  AND3_X2 U3545 ( .A1(fract_out_q[8]), .A2(net85121), .A3(net85145), .ZN(n3175) );
  INV_X16 U3546 ( .A(net85121), .ZN(net85111) );
  NAND2_X1 U3547 ( .A1(net23104), .A2(net94566), .ZN(n3508) );
  NAND2_X4 U3548 ( .A1(net91817), .A2(net84311), .ZN(n3411) );
  NAND4_X2 U3549 ( .A1(n3393), .A2(n2571), .A3(n2985), .A4(n3392), .ZN(
        net84237) );
  INV_X1 U3550 ( .A(fract_denorm[21]), .ZN(n3418) );
  NOR2_X2 U3551 ( .A1(fract_denorm[24]), .A2(net83638), .ZN(n3430) );
  INV_X8 U3552 ( .A(net85141), .ZN(net85139) );
  INV_X8 U3553 ( .A(n3244), .ZN(n3284) );
  NAND3_X2 U3554 ( .A1(fract_i2f[47]), .A2(net85145), .A3(net85111), .ZN(n3279) );
  NOR2_X2 U3555 ( .A1(net84490), .A2(n3287), .ZN(n3339) );
  NOR3_X2 U3556 ( .A1(n2647), .A2(net85111), .A3(net85135), .ZN(n3260) );
  NOR2_X1 U3557 ( .A1(net85115), .A2(net92028), .ZN(n3194) );
  NOR3_X2 U3558 ( .A1(n3042), .A2(net85139), .A3(net90945), .ZN(n3208) );
  NOR2_X1 U3559 ( .A1(n3418), .A2(fract_denorm[22]), .ZN(n3421) );
  NAND4_X2 U3560 ( .A1(net92028), .A2(net85159), .A3(net85179), .A4(quo[15]), 
        .ZN(n3250) );
  NOR4_X1 U3561 ( .A1(n3615), .A2(n3614), .A3(n3613), .A4(n2474), .ZN(n3616)
         );
  AND2_X2 U3562 ( .A1(net85139), .A2(net86295), .ZN(n3176) );
  NOR2_X4 U3563 ( .A1(fract_denorm[26]), .A2(fract_denorm[27]), .ZN(n3010) );
  INV_X4 U3564 ( .A(n3010), .ZN(n3333) );
  INV_X2 U3565 ( .A(fract_denorm[26]), .ZN(n3373) );
  NOR2_X1 U3566 ( .A1(n2983), .A2(n2671), .ZN(net83957) );
  AND2_X4 U3567 ( .A1(n3375), .A2(n3009), .ZN(n3015) );
  INV_X4 U3568 ( .A(n3405), .ZN(n3395) );
  INV_X8 U3569 ( .A(fract_denorm[25]), .ZN(n3360) );
  INV_X16 U3570 ( .A(net85145), .ZN(net85131) );
  INV_X2 U3571 ( .A(n3016), .ZN(n3017) );
  NOR4_X1 U3572 ( .A1(n1756), .A2(n2982), .A3(u6_N13), .A4(n2986), .ZN(n1749)
         );
  INV_X4 U3573 ( .A(n3019), .ZN(n3020) );
  OAI22_X4 U3574 ( .A1(net86014), .A2(n2537), .B1(n3865), .B2(net85998), .ZN(
        n4107) );
  OAI22_X4 U3575 ( .A1(net86015), .A2(n2619), .B1(n3859), .B2(net85998), .ZN(
        n4105) );
  INV_X4 U3576 ( .A(n1451), .ZN(u4_fract_out_8_) );
  NOR2_X1 U3577 ( .A1(net82782), .A2(n4101), .ZN(n4102) );
  INV_X2 U3578 ( .A(n4044), .ZN(n4063) );
  NAND3_X2 U3579 ( .A1(n2058), .A2(n2091), .A3(n2069), .ZN(n3602) );
  NOR3_X4 U3580 ( .A1(u4_N1426), .A2(u4_N1427), .A3(u4_N1428), .ZN(n3653) );
  NAND3_X1 U3581 ( .A1(net82035), .A2(n2903), .A3(n3949), .ZN(n3997) );
  INV_X1 U3582 ( .A(fract_denorm[45]), .ZN(net91594) );
  INV_X2 U3583 ( .A(net91594), .ZN(net91595) );
  NOR2_X4 U3584 ( .A1(fract_denorm[39]), .A2(fract_denorm[40]), .ZN(n3022) );
  INV_X1 U3585 ( .A(n3607), .ZN(n3023) );
  INV_X2 U3586 ( .A(net86040), .ZN(net84450) );
  NOR3_X2 U3587 ( .A1(n2639), .A2(n3274), .A3(net85175), .ZN(n3277) );
  NAND4_X2 U3588 ( .A1(net85135), .A2(net93364), .A3(quo[30]), .A4(net85175), 
        .ZN(n3178) );
  NAND2_X2 U3589 ( .A1(quo[16]), .A2(net86315), .ZN(n3309) );
  NAND2_X4 U3590 ( .A1(n3541), .A2(net86044), .ZN(net83864) );
  OAI211_X4 U3591 ( .C1(net84314), .C2(net84275), .A(n3364), .B(n3365), .ZN(
        n3376) );
  NOR2_X4 U3592 ( .A1(n3460), .A2(net95297), .ZN(n3027) );
  INV_X1 U3593 ( .A(fract_denorm[44]), .ZN(net84225) );
  AOI22_X4 U3594 ( .A1(u4_N1396), .A2(net85377), .B1(u4_N1446), .B2(n2794), 
        .ZN(n1459) );
  NOR2_X2 U3595 ( .A1(net85905), .A2(net83234), .ZN(n3466) );
  INV_X1 U3596 ( .A(n2981), .ZN(n3406) );
  INV_X1 U3597 ( .A(net95137), .ZN(net83776) );
  AOI22_X4 U3598 ( .A1(u4_N1397), .A2(net85377), .B1(u4_N1447), .B2(n2794), 
        .ZN(n2069) );
  NOR2_X1 U3599 ( .A1(u4_f2i_shft_6_), .A2(u4_f2i_shft_7_), .ZN(net83807) );
  NAND3_X1 U3600 ( .A1(net84182), .A2(n3029), .A3(n2552), .ZN(n3427) );
  INV_X8 U3601 ( .A(n3356), .ZN(fract_denorm[34]) );
  NAND4_X2 U3602 ( .A1(quo[16]), .A2(net85179), .A3(net85135), .A4(net85157), 
        .ZN(n3269) );
  INV_X1 U3603 ( .A(n3424), .ZN(n3400) );
  NAND3_X1 U3604 ( .A1(net84204), .A2(net84205), .A3(n3416), .ZN(n3417) );
  INV_X4 U3605 ( .A(net84400), .ZN(net84396) );
  INV_X1 U3606 ( .A(n5324), .ZN(n3396) );
  NAND2_X4 U3607 ( .A1(n3666), .A2(net83624), .ZN(n3336) );
  NOR2_X2 U3608 ( .A1(net83316), .A2(n3696), .ZN(n3697) );
  INV_X1 U3609 ( .A(n3473), .ZN(n3511) );
  INV_X1 U3610 ( .A(n2926), .ZN(n3492) );
  NOR2_X1 U3611 ( .A1(u6_N15), .A2(n2672), .ZN(n4307) );
  NOR2_X1 U3612 ( .A1(net83316), .A2(net95574), .ZN(n3771) );
  INV_X4 U3613 ( .A(n3053), .ZN(n3030) );
  INV_X4 U3614 ( .A(n3031), .ZN(n3032) );
  INV_X8 U3615 ( .A(n2682), .ZN(n3039) );
  INV_X4 U3616 ( .A(n3034), .ZN(n3035) );
  INV_X1 U3617 ( .A(u6_N17), .ZN(n4626) );
  OAI221_X2 U3618 ( .B1(n3481), .B2(net83750), .C1(n2820), .C2(net83753), .A(
        n3480), .ZN(net83020) );
  NAND2_X4 U3619 ( .A1(n3027), .A2(net85933), .ZN(n3458) );
  XNOR2_X1 U3620 ( .A(n3089), .B(n2914), .ZN(u4_f2i_shft_2_) );
  INV_X1 U3621 ( .A(n2682), .ZN(n3040) );
  NOR2_X1 U3622 ( .A1(fract_denorm[44]), .A2(net94305), .ZN(net84306) );
  OAI21_X1 U3623 ( .B1(n2970), .B2(n3971), .A(net95132), .ZN(n3974) );
  INV_X1 U3624 ( .A(net84117), .ZN(net84115) );
  NOR2_X4 U3625 ( .A1(n3473), .A2(net94004), .ZN(n3041) );
  NAND2_X1 U3626 ( .A1(fract_i2f[34]), .A2(net85115), .ZN(n3272) );
  NAND2_X1 U3627 ( .A1(fract_i2f[17]), .A2(net85115), .ZN(n3147) );
  INV_X1 U3628 ( .A(u6_N18), .ZN(n4496) );
  AOI22_X4 U3629 ( .A1(n3238), .A2(prod[44]), .B1(fract_i2f[44]), .B2(net85115), .ZN(net84557) );
  NAND3_X1 U3630 ( .A1(fract_out_q[21]), .A2(net85121), .A3(net85145), .ZN(
        n3286) );
  NAND3_X1 U3631 ( .A1(fract_out_q[27]), .A2(net85143), .A3(net85121), .ZN(
        n3280) );
  NAND3_X1 U3632 ( .A1(net85121), .A2(net85145), .A3(fract_out_q[11]), .ZN(
        n3220) );
  NAND3_X1 U3633 ( .A1(net85121), .A2(net85143), .A3(fract_out_q[12]), .ZN(
        n3225) );
  NAND3_X1 U3634 ( .A1(fract_out_q[14]), .A2(net85121), .A3(net85143), .ZN(
        n3273) );
  INV_X8 U3635 ( .A(fract_denorm[29]), .ZN(n3428) );
  INV_X8 U3636 ( .A(n1456), .ZN(u4_fract_out_19_) );
  AOI22_X4 U3637 ( .A1(u4_N1402), .A2(net85377), .B1(u4_N1452), .B2(n2794), 
        .ZN(n1456) );
  NAND2_X2 U3638 ( .A1(net84377), .A2(n3398), .ZN(n3382) );
  OR2_X1 U3639 ( .A1(u6_N1), .A2(n3040), .ZN(n1754) );
  NOR2_X4 U3640 ( .A1(n5324), .A2(n5325), .ZN(n3048) );
  NAND4_X2 U3641 ( .A1(n3378), .A2(net84101), .A3(n2899), .A4(n3377), .ZN(
        net83759) );
  NOR4_X1 U3642 ( .A1(n2968), .A2(u6_N18), .A3(u6_N17), .A4(n2963), .ZN(n4306)
         );
  NAND2_X1 U3643 ( .A1(net83744), .A2(n2500), .ZN(n3519) );
  OAI22_X4 U3644 ( .A1(net86015), .A2(n2641), .B1(net86001), .B2(n3778), .ZN(
        n3779) );
  OR3_X2 U3645 ( .A1(n3026), .A2(net84490), .A3(net85167), .ZN(n3071) );
  NOR2_X1 U3646 ( .A1(n3265), .A2(net85167), .ZN(n3267) );
  NOR2_X1 U3647 ( .A1(n3511), .A2(net84000), .ZN(n3502) );
  NAND2_X1 U3648 ( .A1(u4_fi_ldz_2a_3_), .A2(net86532), .ZN(n3381) );
  NAND2_X1 U3649 ( .A1(div_opa_ldz_r2[3]), .A2(u4_fi_ldz_2a_3_), .ZN(n3450) );
  NAND3_X2 U3650 ( .A1(net85165), .A2(net85133), .A3(prod[34]), .ZN(n3271) );
  NAND3_X2 U3651 ( .A1(prod[17]), .A2(net85165), .A3(net85131), .ZN(n3148) );
  INV_X1 U3652 ( .A(net83753), .ZN(net83751) );
  INV_X8 U3653 ( .A(n3336), .ZN(n3386) );
  INV_X8 U3654 ( .A(n3389), .ZN(n3375) );
  NOR2_X2 U3655 ( .A1(net83632), .A2(net84242), .ZN(n3354) );
  NAND3_X2 U3656 ( .A1(n3326), .A2(n3325), .A3(n3324), .ZN(net17654) );
  AOI22_X4 U3657 ( .A1(n3154), .A2(prod[39]), .B1(fract_i2f[39]), .B2(net85115), .ZN(n3212) );
  NOR2_X1 U3658 ( .A1(net17686), .A2(net17682), .ZN(n3665) );
  INV_X2 U3659 ( .A(net17686), .ZN(net84231) );
  NAND2_X1 U3660 ( .A1(net84377), .A2(n2959), .ZN(n3425) );
  NOR3_X1 U3661 ( .A1(n3604), .A2(net92015), .A3(net94138), .ZN(n3605) );
  OAI21_X1 U3662 ( .B1(net83714), .B2(net94138), .A(net84224), .ZN(n3403) );
  NOR2_X2 U3663 ( .A1(net85143), .A2(n3275), .ZN(n3276) );
  NAND3_X2 U3664 ( .A1(quo[36]), .A2(net85175), .A3(net85157), .ZN(n3275) );
  OAI22_X4 U3665 ( .A1(net86015), .A2(n3874), .B1(net86001), .B2(n3873), .ZN(
        net82807) );
  NAND3_X2 U3666 ( .A1(prod[18]), .A2(net85165), .A3(net85131), .ZN(n3145) );
  NAND4_X1 U3667 ( .A1(n3680), .A2(net94566), .A3(n3679), .A4(n2476), .ZN(
        n3789) );
  NOR2_X1 U3668 ( .A1(n2983), .A2(n3509), .ZN(n3510) );
  INV_X8 U3670 ( .A(n4101), .ZN(n4025) );
  INV_X1 U3671 ( .A(net93364), .ZN(net86309) );
  NAND4_X1 U3672 ( .A1(net85179), .A2(quo[10]), .A3(net85157), .A4(net85131), 
        .ZN(n3221) );
  NAND4_X1 U3673 ( .A1(net85179), .A2(quo[11]), .A3(net85157), .A4(net85131), 
        .ZN(n3226) );
  AOI22_X4 U3674 ( .A1(fract_out_q[0]), .A2(n4071), .B1(fract_i2f[20]), .B2(
        net85115), .ZN(n3191) );
  NOR4_X4 U3675 ( .A1(net84396), .A2(net84397), .A3(n3340), .A4(n3339), .ZN(
        n3343) );
  OAI211_X4 U3676 ( .C1(n3282), .C2(n3281), .A(n3280), .B(n3279), .ZN(net84397) );
  AOI22_X4 U3677 ( .A1(net92566), .A2(n3842), .B1(n3055), .B2(net85997), .ZN(
        n3054) );
  INV_X1 U3678 ( .A(n2904), .ZN(n4078) );
  INV_X8 U3679 ( .A(n1460), .ZN(u4_fract_out_12_) );
  AOI22_X4 U3680 ( .A1(u4_N1395), .A2(net85377), .B1(u4_N1445), .B2(n2794), 
        .ZN(n1460) );
  AOI22_X4 U3681 ( .A1(u4_N1383), .A2(net85377), .B1(u4_N1433), .B2(n2794), 
        .ZN(n2093) );
  AOI22_X4 U3682 ( .A1(u4_N1401), .A2(net85377), .B1(u4_N1451), .B2(n2794), 
        .ZN(n1457) );
  NAND3_X2 U3683 ( .A1(n3725), .A2(n3724), .A3(n3723), .ZN(n3730) );
  INV_X1 U3684 ( .A(n2693), .ZN(n3049) );
  AOI21_X1 U3685 ( .B1(n2905), .B2(net83532), .A(net83441), .ZN(n3724) );
  OAI21_X1 U3686 ( .B1(n3985), .B2(net94825), .A(n3963), .ZN(n3964) );
  OAI21_X1 U3687 ( .B1(n3960), .B2(n3959), .A(net94825), .ZN(n3967) );
  NOR2_X2 U3688 ( .A1(n3408), .A2(n3443), .ZN(n3414) );
  NOR3_X1 U3689 ( .A1(net94834), .A2(n3969), .A3(n3968), .ZN(n3970) );
  NAND2_X4 U3690 ( .A1(net83041), .A2(net83928), .ZN(net82932) );
  NAND2_X4 U3691 ( .A1(net83836), .A2(net86045), .ZN(net83928) );
  INV_X4 U3692 ( .A(n3033), .ZN(n3050) );
  NAND3_X1 U3693 ( .A1(net95148), .A2(n2928), .A3(n2495), .ZN(n3958) );
  NOR2_X4 U3694 ( .A1(n2665), .A2(n4021), .ZN(n4022) );
  OAI22_X4 U3695 ( .A1(net85998), .A2(n3861), .B1(n2538), .B2(net86014), .ZN(
        n4103) );
  OAI22_X4 U3696 ( .A1(net85998), .A2(n3852), .B1(net86015), .B2(n3851), .ZN(
        n4080) );
  NOR4_X1 U3697 ( .A1(fracta_mul[3]), .A2(fracta_mul[2]), .A3(fracta_mul[20]), 
        .A4(n2586), .ZN(n1744) );
  INV_X1 U3698 ( .A(n2586), .ZN(n4523) );
  OAI21_X4 U3699 ( .B1(net83274), .B2(n3824), .A(net83275), .ZN(net86486) );
  OAI21_X2 U3700 ( .B1(n3795), .B2(net94703), .A(net83278), .ZN(n3844) );
  NAND3_X2 U3701 ( .A1(n3706), .A2(n3705), .A3(net83555), .ZN(n3823) );
  AOI22_X4 U3702 ( .A1(n3856), .A2(net86013), .B1(n2560), .B2(net85997), .ZN(
        n3051) );
  AOI21_X2 U3703 ( .B1(n4073), .B2(n4072), .A(net82829), .ZN(N526) );
  NOR2_X1 U3704 ( .A1(n3930), .A2(net83066), .ZN(n3932) );
  INV_X1 U3705 ( .A(net83066), .ZN(net86401) );
  NAND3_X2 U3706 ( .A1(net83214), .A2(n3848), .A3(n3847), .ZN(net82876) );
  NOR2_X1 U3707 ( .A1(u6_N22), .A2(n2604), .ZN(u0_N5) );
  INV_X1 U3708 ( .A(u6_N22), .ZN(n4491) );
  OAI22_X4 U3709 ( .A1(net85999), .A2(n3899), .B1(n3898), .B2(net86014), .ZN(
        n4098) );
  NOR2_X4 U3710 ( .A1(net83279), .A2(net83288), .ZN(n3796) );
  NAND4_X4 U3711 ( .A1(n3816), .A2(n3817), .A3(net83297), .A4(n3798), .ZN(
        n3820) );
  INV_X2 U3712 ( .A(n3820), .ZN(n3802) );
  AND2_X2 U3713 ( .A1(net86481), .A2(u4_fract_out_1_), .ZN(n3055) );
  NAND2_X4 U3714 ( .A1(n3920), .A2(n2779), .ZN(n4032) );
  INV_X8 U3715 ( .A(n4080), .ZN(n4034) );
  NOR2_X2 U3716 ( .A1(net82782), .A2(n2997), .ZN(n4081) );
  AOI21_X1 U3717 ( .B1(n4524), .B2(n2586), .A(fracta_mul[3]), .ZN(n2445) );
  NAND2_X4 U3718 ( .A1(n3845), .A2(n2673), .ZN(n4122) );
  NAND2_X4 U3719 ( .A1(n3804), .A2(n3700), .ZN(net83435) );
  NOR2_X1 U3720 ( .A1(net82782), .A2(n2462), .ZN(n4084) );
  INV_X8 U3721 ( .A(net82764), .ZN(net83066) );
  NOR2_X1 U3722 ( .A1(net82782), .A2(n2461), .ZN(n4099) );
  NAND4_X4 U3723 ( .A1(n3832), .A2(n3830), .A3(n2954), .A4(n3831), .ZN(
        net82902) );
  NAND3_X2 U3724 ( .A1(net82891), .A2(net95549), .A3(net82893), .ZN(n4033) );
  NAND2_X1 U3725 ( .A1(n3895), .A2(u4_fract_out_17_), .ZN(n3894) );
  AOI22_X4 U3726 ( .A1(u4_N1403), .A2(net85377), .B1(u4_N1453), .B2(n2794), 
        .ZN(n2060) );
  INV_X1 U3727 ( .A(n2484), .ZN(net82951) );
  INV_X8 U3728 ( .A(n1458), .ZN(u4_fract_out_17_) );
  AOI22_X4 U3729 ( .A1(u4_N1400), .A2(net85377), .B1(u4_N1450), .B2(n2794), 
        .ZN(n1458) );
  AOI22_X4 U3730 ( .A1(u4_N1404), .A2(net85377), .B1(u4_N1454), .B2(n2794), 
        .ZN(n2058) );
  OAI22_X4 U3731 ( .A1(n2644), .A2(net86015), .B1(n3863), .B2(net85999), .ZN(
        n4101) );
  AOI22_X4 U3732 ( .A1(u4_N1391), .A2(net85377), .B1(u4_N1441), .B2(n2794), 
        .ZN(n1451) );
  INV_X2 U3733 ( .A(u4_fract_out_pl1_23_), .ZN(net83562) );
  OAI22_X4 U3734 ( .A1(n3894), .A2(net85998), .B1(n3893), .B2(net86014), .ZN(
        n4100) );
  AND2_X2 U3735 ( .A1(n3061), .A2(n3062), .ZN(n3098) );
  AOI21_X1 U3736 ( .B1(n3687), .B2(n2467), .A(n3686), .ZN(n3706) );
  AOI21_X1 U3737 ( .B1(n3717), .B2(n2467), .A(n3716), .ZN(n3720) );
  NAND2_X1 U3738 ( .A1(n3745), .A2(n2467), .ZN(n3746) );
  NAND2_X1 U3739 ( .A1(net83368), .A2(n2467), .ZN(n3808) );
  AOI22_X4 U3740 ( .A1(u4_N1390), .A2(net85377), .B1(u4_N1440), .B2(n2794), 
        .ZN(n1452) );
  NOR2_X1 U3741 ( .A1(opb_r[25]), .A2(n2765), .ZN(n4441) );
  NAND2_X1 U3742 ( .A1(opb_r[27]), .A2(n2657), .ZN(n4460) );
  INV_X1 U3743 ( .A(n2930), .ZN(n4765) );
  INV_X8 U3744 ( .A(n2076), .ZN(u4_fract_out_10_) );
  AOI22_X4 U3745 ( .A1(u4_N1393), .A2(net85377), .B1(u4_N1443), .B2(n2794), 
        .ZN(n2076) );
  NAND3_X1 U3746 ( .A1(n1454), .A2(n1453), .A3(n3016), .ZN(n2245) );
  NAND2_X4 U3747 ( .A1(n2539), .A2(n3589), .ZN(u4_fract_out_22_) );
  AOI22_X4 U3748 ( .A1(u4_N1399), .A2(net85377), .B1(u4_N1449), .B2(n2794), 
        .ZN(n2065) );
  INV_X8 U3749 ( .A(n2065), .ZN(u4_fract_out_16_) );
  NOR3_X2 U3750 ( .A1(net85145), .A2(net85159), .A3(n2642), .ZN(n3161) );
  NOR2_X1 U3751 ( .A1(n3341), .A2(n3340), .ZN(n3290) );
  NAND3_X2 U3752 ( .A1(n3290), .A2(n3289), .A3(n3288), .ZN(net28939) );
  NAND2_X4 U3753 ( .A1(n3010), .A2(n3375), .ZN(n3359) );
  NAND2_X1 U3754 ( .A1(net86315), .A2(quo[2]), .ZN(n3441) );
  NAND2_X1 U3755 ( .A1(quo[3]), .A2(net86315), .ZN(n3327) );
  NAND2_X1 U3756 ( .A1(quo[4]), .A2(net86315), .ZN(n3330) );
  NAND2_X1 U3757 ( .A1(quo[6]), .A2(net86315), .ZN(n3318) );
  NAND2_X1 U3758 ( .A1(quo[7]), .A2(net86315), .ZN(n3321) );
  NAND2_X1 U3759 ( .A1(quo[8]), .A2(net86315), .ZN(n3324) );
  NOR2_X1 U3760 ( .A1(net85145), .A2(n2650), .ZN(n3167) );
  NOR2_X1 U3761 ( .A1(net90897), .A2(net85159), .ZN(n3224) );
  NAND3_X1 U3762 ( .A1(n2979), .A2(n2985), .A3(n3665), .ZN(n3667) );
  NAND3_X2 U3763 ( .A1(n3427), .A2(net85393), .A3(n3426), .ZN(n3435) );
  INV_X2 U3764 ( .A(net86571), .ZN(net84302) );
  AOI22_X4 U3765 ( .A1(n3174), .A2(prod[40]), .B1(fract_i2f[40]), .B2(net85115), .ZN(n3218) );
  AND2_X4 U3766 ( .A1(n3195), .A2(n3071), .ZN(n3196) );
  INV_X8 U3767 ( .A(n2957), .ZN(n3090) );
  NOR2_X2 U3768 ( .A1(n3511), .A2(n3510), .ZN(n3513) );
  NOR3_X2 U3769 ( .A1(n3443), .A2(net84149), .A3(net84150), .ZN(net84142) );
  NAND2_X4 U3770 ( .A1(n3363), .A2(net84205), .ZN(n3419) );
  NAND2_X4 U3771 ( .A1(n3346), .A2(net92738), .ZN(net84298) );
  NAND4_X4 U3772 ( .A1(n3096), .A2(n3098), .A3(n3097), .A4(n3099), .ZN(u6_N23)
         );
  NAND4_X1 U3773 ( .A1(n3608), .A2(n3607), .A3(n3605), .A4(n3029), .ZN(n3615)
         );
  NOR2_X1 U3774 ( .A1(n2482), .A2(n2483), .ZN(net84349) );
  NAND2_X4 U3775 ( .A1(net85135), .A2(net85159), .ZN(n3213) );
  NAND2_X4 U3776 ( .A1(n3283), .A2(net84496), .ZN(net84400) );
  NOR2_X4 U3777 ( .A1(n3244), .A2(net90897), .ZN(n3072) );
  NOR3_X1 U3778 ( .A1(n3006), .A2(n3008), .A3(n3021), .ZN(n3385) );
  NAND3_X2 U3779 ( .A1(quo[20]), .A2(net85133), .A3(n3284), .ZN(n3285) );
  NAND2_X4 U3780 ( .A1(net93218), .A2(n3448), .ZN(u4_fi_ldz_mi1_3_) );
  NAND2_X4 U3781 ( .A1(n3338), .A2(n2564), .ZN(net84323) );
  NAND2_X1 U3782 ( .A1(opb_r[28]), .A2(opb_r[27]), .ZN(n4735) );
  OAI22_X1 U3783 ( .A1(opb_r[28]), .A2(n2582), .B1(opb_r[27]), .B2(n2657), 
        .ZN(n4446) );
  AOI22_X4 U3784 ( .A1(u4_N1382), .A2(net85377), .B1(u4_N1432), .B2(n2794), 
        .ZN(n2278) );
  NAND3_X1 U3785 ( .A1(n2903), .A2(net85179), .A3(n3990), .ZN(n3991) );
  AOI22_X4 U3786 ( .A1(fract_out_q[6]), .A2(n3150), .B1(n3072), .B2(quo[5]), 
        .ZN(n3151) );
  NAND2_X1 U3787 ( .A1(quo[43]), .A2(net85159), .ZN(n3287) );
  NAND4_X4 U3788 ( .A1(n3223), .A2(n3222), .A3(n3221), .A4(n3220), .ZN(
        fract_denorm[31]) );
  AOI22_X4 U3789 ( .A1(fract_out_q[7]), .A2(n3150), .B1(n3072), .B2(quo[6]), 
        .ZN(n3155) );
  NOR2_X1 U3790 ( .A1(net86040), .A2(n2648), .ZN(n3190) );
  NOR3_X1 U3791 ( .A1(net86040), .A2(net85143), .A3(n2651), .ZN(n3149) );
  OAI21_X1 U3792 ( .B1(net85111), .B2(net93364), .A(n2927), .ZN(n4112) );
  OAI21_X1 U3793 ( .B1(net23043), .B2(net33106), .A(net83762), .ZN(n3596) );
  NOR2_X1 U3794 ( .A1(opa_r[30]), .A2(opb_r[30]), .ZN(n4313) );
  OAI22_X1 U3795 ( .A1(u2_N124), .A2(n4741), .B1(n2930), .B2(n4742), .ZN(n4312) );
  NOR2_X1 U3796 ( .A1(opa_r[30]), .A2(n2930), .ZN(n4319) );
  NOR2_X1 U3797 ( .A1(opa_r[30]), .A2(opb_r[30]), .ZN(n4465) );
  NAND2_X1 U3798 ( .A1(opb_r[30]), .A2(n2566), .ZN(n4455) );
  INV_X1 U3799 ( .A(n3419), .ZN(n3420) );
  NAND2_X4 U3800 ( .A1(n2976), .A2(n3476), .ZN(net84067) );
  AOI22_X1 U3801 ( .A1(net84321), .A2(n3372), .B1(n2471), .B2(net93404), .ZN(
        n3378) );
  NOR2_X1 U3802 ( .A1(n3391), .A2(net83624), .ZN(n3393) );
  NOR3_X2 U3803 ( .A1(n3391), .A2(net92690), .A3(net83721), .ZN(n3431) );
  NOR2_X1 U3804 ( .A1(net92573), .A2(n3409), .ZN(n3379) );
  NAND2_X4 U3805 ( .A1(net83638), .A2(n3334), .ZN(n3612) );
  INV_X8 U3806 ( .A(net84158), .ZN(net84140) );
  NAND3_X1 U3807 ( .A1(n2545), .A2(n3021), .A3(n3407), .ZN(n3372) );
  NAND2_X4 U3808 ( .A1(n3955), .A2(net86027), .ZN(n3591) );
  NAND2_X4 U3809 ( .A1(net86315), .A2(quo[12]), .ZN(n3297) );
  INV_X1 U3810 ( .A(n3444), .ZN(n3446) );
  INV_X8 U3811 ( .A(net92573), .ZN(net84205) );
  NAND2_X4 U3812 ( .A1(n3459), .A2(net84054), .ZN(u4_f2i_shft_7_) );
  NAND2_X4 U3813 ( .A1(net94146), .A2(net84083), .ZN(u4_fi_ldz_mi1_1_) );
  NOR2_X1 U3814 ( .A1(n2554), .A2(net84353), .ZN(n3344) );
  NAND2_X1 U3815 ( .A1(net95138), .A2(net83368), .ZN(n3788) );
  XNOR2_X1 U3816 ( .A(net95431), .B(net33106), .ZN(u4_fi_ldz_mi22[2]) );
  NAND2_X1 U3817 ( .A1(net83878), .A2(n2469), .ZN(n3566) );
  NAND2_X4 U3818 ( .A1(n3422), .A2(n3351), .ZN(net84257) );
  NAND2_X4 U3819 ( .A1(net91406), .A2(net85179), .ZN(n3244) );
  NAND2_X4 U3820 ( .A1(n3048), .A2(n3386), .ZN(net84191) );
  NAND3_X2 U3821 ( .A1(n2909), .A2(net95479), .A3(n3335), .ZN(n3345) );
  NAND3_X2 U3822 ( .A1(n3394), .A2(n5324), .A3(net91297), .ZN(n3397) );
  NOR2_X1 U3823 ( .A1(net82782), .A2(n2964), .ZN(n4097) );
  NAND3_X1 U3824 ( .A1(net84205), .A2(n2474), .A3(n3608), .ZN(n3365) );
  AOI211_X2 U3825 ( .C1(n3385), .C2(net84205), .A(net84348), .B(n3384), .ZN(
        net84285) );
  NAND2_X1 U3826 ( .A1(net84341), .A2(net84205), .ZN(net84275) );
  NAND3_X2 U3827 ( .A1(net84205), .A2(n2973), .A3(n3374), .ZN(n3402) );
  NAND3_X1 U3828 ( .A1(n4115), .A2(net85121), .A3(n4114), .ZN(n4116) );
  NAND2_X1 U3829 ( .A1(n3999), .A2(n3998), .ZN(n4000) );
  NAND3_X1 U3830 ( .A1(n3807), .A2(net85905), .A3(net82929), .ZN(n3809) );
  AOI22_X1 U3831 ( .A1(u4_exp_next_mi_3_), .A2(net83532), .B1(
        u4_exp_fix_diva[3]), .B2(net83312), .ZN(n3753) );
  NAND3_X1 U3832 ( .A1(net85929), .A2(net82929), .A3(n3807), .ZN(n3727) );
  NAND3_X1 U3833 ( .A1(n3088), .A2(net82929), .A3(n3807), .ZN(n3748) );
  NAND3_X1 U3834 ( .A1(n3085), .A2(net82929), .A3(n3807), .ZN(n3685) );
  NAND2_X1 U3835 ( .A1(net82929), .A2(n3807), .ZN(net83434) );
  NAND2_X4 U3836 ( .A1(n3807), .A2(n3703), .ZN(net83495) );
  OAI21_X1 U3837 ( .B1(u4_fi_ldz_2a_3_), .B2(net86532), .A(n3381), .ZN(
        u4_fi_ldz_2a_4_) );
  NOR2_X1 U3838 ( .A1(div_opa_ldz_r2[3]), .A2(u4_fi_ldz_2a_3_), .ZN(n3451) );
  XNOR2_X1 U3839 ( .A(u4_fi_ldz_2a_3_), .B(div_opa_ldz_r2[3]), .ZN(n3457) );
  NAND2_X4 U3840 ( .A1(net84140), .A2(net84141), .ZN(n4758) );
  OAI22_X4 U3841 ( .A1(net86001), .A2(n3881), .B1(n3880), .B2(net86014), .ZN(
        n4087) );
  NAND2_X4 U3842 ( .A1(n3041), .A2(n3493), .ZN(n3475) );
  NAND2_X4 U3843 ( .A1(n3917), .A2(n3921), .ZN(n4036) );
  NOR2_X1 U3844 ( .A1(net82782), .A2(n3001), .ZN(n4090) );
  AOI221_X1 U3845 ( .B1(n2903), .B2(net82034), .C1(n4000), .C2(net94811), .A(
        n2603), .ZN(n4005) );
  NAND2_X1 U3846 ( .A1(net86497), .A2(n2550), .ZN(n3859) );
  NAND4_X1 U3847 ( .A1(net83498), .A2(n2501), .A3(net83500), .A4(net94692), 
        .ZN(n3743) );
  AOI21_X1 U3848 ( .B1(net94725), .B2(net94811), .A(net83837), .ZN(n3575) );
  NAND2_X1 U3849 ( .A1(net83933), .A2(net94725), .ZN(net83927) );
  NOR2_X1 U3850 ( .A1(n3423), .A2(net92599), .ZN(net84189) );
  INV_X8 U3851 ( .A(net85985), .ZN(net85986) );
  INV_X8 U3852 ( .A(net85985), .ZN(net85987) );
  INV_X8 U3853 ( .A(net85985), .ZN(net85988) );
  INV_X8 U3854 ( .A(net85985), .ZN(net85989) );
  INV_X32 U3855 ( .A(net85975), .ZN(net85976) );
  INV_X8 U3856 ( .A(n4436), .ZN(n3073) );
  NAND2_X4 U3857 ( .A1(N251), .A2(n4389), .ZN(n4436) );
  INV_X32 U3858 ( .A(n4670), .ZN(n3075) );
  INV_X32 U3859 ( .A(n3075), .ZN(n3076) );
  INV_X32 U3860 ( .A(n3075), .ZN(n3077) );
  INV_X32 U3861 ( .A(n3075), .ZN(n3078) );
  INV_X16 U3862 ( .A(n3079), .ZN(n3080) );
  INV_X16 U3863 ( .A(n3079), .ZN(n3081) );
  INV_X16 U3864 ( .A(n3079), .ZN(n3082) );
  INV_X16 U3865 ( .A(n3079), .ZN(n3083) );
  INV_X16 U3866 ( .A(n3079), .ZN(n3084) );
  INV_X32 U3867 ( .A(net85932), .ZN(net85933) );
  INV_X8 U3868 ( .A(exp_r[3]), .ZN(n3086) );
  INV_X8 U3869 ( .A(n3086), .ZN(n3087) );
  INV_X8 U3870 ( .A(n3086), .ZN(n3088) );
  INV_X32 U3871 ( .A(net85393), .ZN(net85391) );
  INV_X32 U3872 ( .A(net83796), .ZN(net85377) );
  NOR2_X4 U3873 ( .A1(opa_r[29]), .A2(opa_r[30]), .ZN(n3103) );
  NAND4_X2 U3874 ( .A1(n3103), .A2(n3102), .A3(n3101), .A4(n3100), .ZN(u2_N124) );
  NAND2_X2 U3875 ( .A1(n2697), .A2(n2451), .ZN(n3111) );
  NAND2_X2 U3876 ( .A1(n3105), .A2(n3104), .ZN(n3110) );
  INV_X4 U3877 ( .A(n3110), .ZN(n3109) );
  NAND2_X2 U3878 ( .A1(n2599), .A2(n2683), .ZN(n3120) );
  INV_X4 U3879 ( .A(n3120), .ZN(n3106) );
  NAND2_X2 U3880 ( .A1(n3106), .A2(n2591), .ZN(n3117) );
  INV_X4 U3881 ( .A(n3117), .ZN(n3108) );
  NOR4_X2 U3882 ( .A1(fracta_mul[16]), .A2(fracta_mul[17]), .A3(fracta_mul[19]), .A4(fracta_mul[18]), .ZN(n3119) );
  INV_X4 U3883 ( .A(n3111), .ZN(n3112) );
  INV_X4 U3884 ( .A(n2692), .ZN(n3113) );
  NAND3_X4 U3885 ( .A1(n2590), .A2(n2675), .A3(n2448), .ZN(n3121) );
  AOI21_X4 U3886 ( .B1(n3122), .B2(n3121), .A(n3120), .ZN(n3123) );
  NAND2_X2 U3887 ( .A1(n2697), .A2(n3124), .ZN(n3125) );
  INV_X4 U3888 ( .A(n2687), .ZN(n3126) );
  INV_X4 U3889 ( .A(N195), .ZN(n3132) );
  NAND2_X2 U3890 ( .A1(n3132), .A2(n3092), .ZN(u6_N49) );
  NOR2_X4 U3891 ( .A1(n3091), .A2(net85905), .ZN(n3464) );
  INV_X4 U3892 ( .A(n3137), .ZN(n3133) );
  INV_X4 U3893 ( .A(net84736), .ZN(net84737) );
  NAND2_X2 U3894 ( .A1(net82029), .A2(n2618), .ZN(net84054) );
  NAND2_X2 U3895 ( .A1(n3134), .A2(net86045), .ZN(n3135) );
  NAND2_X2 U3896 ( .A1(net86045), .A2(net82029), .ZN(net84030) );
  NAND2_X2 U3897 ( .A1(n3135), .A2(net84030), .ZN(net82023) );
  INV_X4 U3898 ( .A(net82023), .ZN(u4_exp_in_mi1_7_) );
  XNOR2_X2 U3899 ( .A(net84738), .B(n2618), .ZN(net82010) );
  INV_X4 U3900 ( .A(net82010), .ZN(u4_exp_in_mi1_6_) );
  NOR2_X4 U3901 ( .A1(n3464), .A2(n3479), .ZN(n3462) );
  NAND2_X2 U3902 ( .A1(n3138), .A2(n3137), .ZN(u4_exp_in_mi1_2_) );
  OAI21_X4 U3903 ( .B1(net22501), .B2(n3734), .A(n3961), .ZN(u4_exp_in_mi1_1_)
         );
  NAND2_X2 U3904 ( .A1(prod[19]), .A2(n2936), .ZN(n3142) );
  NAND2_X2 U3905 ( .A1(fract_i2f[19]), .A2(net85117), .ZN(n3141) );
  NAND3_X4 U3906 ( .A1(quo[21]), .A2(net84605), .A3(net85131), .ZN(n3140) );
  NAND3_X4 U3907 ( .A1(n3142), .A2(n3141), .A3(n3140), .ZN(net17682) );
  NAND2_X2 U3908 ( .A1(fract_i2f[18]), .A2(net85117), .ZN(n3144) );
  NAND3_X4 U3909 ( .A1(quo[20]), .A2(net84605), .A3(net85131), .ZN(n3143) );
  NAND3_X4 U3910 ( .A1(n3145), .A2(n3144), .A3(n3143), .ZN(net17683) );
  NAND3_X4 U3911 ( .A1(quo[19]), .A2(net84605), .A3(net85131), .ZN(n3146) );
  NAND3_X4 U3912 ( .A1(n3148), .A2(n3147), .A3(n3146), .ZN(net17657) );
  NOR2_X4 U3913 ( .A1(n3149), .A2(n2643), .ZN(n3153) );
  NAND2_X2 U3914 ( .A1(prod[26]), .A2(n2936), .ZN(n3152) );
  NAND3_X4 U3915 ( .A1(n3153), .A2(n3152), .A3(n3151), .ZN(fract_denorm[26])
         );
  AOI22_X2 U3916 ( .A1(n3154), .A2(prod[27]), .B1(fract_i2f[27]), .B2(net85115), .ZN(n3157) );
  NAND3_X4 U3917 ( .A1(quo[29]), .A2(net85133), .A3(net84455), .ZN(n3156) );
  NAND3_X4 U3918 ( .A1(n3157), .A2(n3156), .A3(n3155), .ZN(fract_denorm[27])
         );
  NAND2_X2 U3919 ( .A1(fract_i2f[24]), .A2(net85115), .ZN(n3164) );
  NOR3_X4 U3920 ( .A1(n3159), .A2(n3161), .A3(n3160), .ZN(n3162) );
  NAND3_X4 U3921 ( .A1(n3164), .A2(n3163), .A3(n3162), .ZN(fract_denorm[24])
         );
  NAND2_X2 U3922 ( .A1(fract_i2f[23]), .A2(net85115), .ZN(n3169) );
  NOR2_X4 U3923 ( .A1(net85117), .A2(n2636), .ZN(n3166) );
  AOI22_X2 U3924 ( .A1(n3167), .A2(n3284), .B1(n3166), .B2(net85143), .ZN(
        n3168) );
  NAND3_X4 U3925 ( .A1(quo[27]), .A2(net85133), .A3(net84605), .ZN(n3172) );
  NAND3_X4 U3926 ( .A1(n3173), .A2(n3172), .A3(n3171), .ZN(fract_denorm[25])
         );
  AOI22_X2 U3927 ( .A1(n3174), .A2(prod[28]), .B1(fract_i2f[28]), .B2(net85115), .ZN(n3179) );
  AOI21_X4 U3928 ( .B1(n3176), .B2(quo[7]), .A(n3175), .ZN(n3177) );
  NAND3_X4 U3929 ( .A1(n3177), .A2(n3179), .A3(n3178), .ZN(fract_denorm[28])
         );
  NAND4_X2 U3930 ( .A1(quo[32]), .A2(net85175), .A3(net85159), .A4(net92028), 
        .ZN(n3185) );
  INV_X4 U3931 ( .A(n3180), .ZN(n3182) );
  NAND4_X2 U3932 ( .A1(quo[31]), .A2(net85175), .A3(net85159), .A4(net85135), 
        .ZN(n3189) );
  NAND3_X4 U3933 ( .A1(n3189), .A2(n3188), .A3(n3187), .ZN(fract_denorm[29])
         );
  NAND2_X2 U3934 ( .A1(n3190), .A2(net85133), .ZN(n3193) );
  NAND3_X4 U3935 ( .A1(n3193), .A2(n3192), .A3(n3191), .ZN(net17659) );
  AOI22_X2 U3936 ( .A1(n3194), .A2(fract_out_q[1]), .B1(fract_i2f[21]), .B2(
        net85115), .ZN(n3198) );
  NAND3_X4 U3937 ( .A1(n3198), .A2(n3197), .A3(n3196), .ZN(fract_denorm[21])
         );
  INV_X4 U3938 ( .A(n3200), .ZN(n3201) );
  NAND3_X4 U3939 ( .A1(n3202), .A2(n3203), .A3(n3204), .ZN(fract_denorm[22])
         );
  NAND3_X4 U3940 ( .A1(quo[35]), .A2(net84605), .A3(net85131), .ZN(n3206) );
  AOI22_X2 U3941 ( .A1(fract_out_q[13]), .A2(n3150), .B1(quo[12]), .B2(n3072), 
        .ZN(n3205) );
  NAND3_X4 U3942 ( .A1(n2473), .A2(n3206), .A3(n3205), .ZN(fract_denorm[33])
         );
  NAND4_X2 U3943 ( .A1(quo[41]), .A2(net85175), .A3(net92028), .A4(net85159), 
        .ZN(n3211) );
  AOI21_X4 U3944 ( .B1(n3209), .B2(quo[18]), .A(n3208), .ZN(n3210) );
  NAND4_X2 U3945 ( .A1(quo[42]), .A2(net85175), .A3(net92028), .A4(net85159), 
        .ZN(n3217) );
  AOI21_X4 U3946 ( .B1(n3215), .B2(quo[19]), .A(n3214), .ZN(n3216) );
  NAND3_X4 U3947 ( .A1(n3216), .A2(n3217), .A3(n3218), .ZN(fract_denorm[40])
         );
  AOI22_X2 U3948 ( .A1(n3219), .A2(prod[31]), .B1(fract_i2f[31]), .B2(net85115), .ZN(n3223) );
  AOI22_X2 U3949 ( .A1(n3224), .A2(prod[32]), .B1(fract_i2f[32]), .B2(net85115), .ZN(n3228) );
  AOI22_X2 U3950 ( .A1(n3238), .A2(prod[43]), .B1(fract_i2f[43]), .B2(net85115), .ZN(n3233) );
  NAND4_X2 U3951 ( .A1(quo[45]), .A2(net85175), .A3(net85131), .A4(net85159), 
        .ZN(n3232) );
  AOI21_X4 U3952 ( .B1(n3261), .B2(quo[22]), .A(n3230), .ZN(n3231) );
  NAND3_X4 U3953 ( .A1(n3233), .A2(n3232), .A3(n3231), .ZN(fract_denorm[43])
         );
  NAND3_X4 U3954 ( .A1(n3235), .A2(n3236), .A3(n3237), .ZN(fract_denorm[45])
         );
  NAND4_X2 U3955 ( .A1(quo[44]), .A2(net85175), .A3(net85133), .A4(net85159), 
        .ZN(n3241) );
  AOI21_X4 U3956 ( .B1(net84568), .B2(quo[21]), .A(n3239), .ZN(n3240) );
  NAND2_X2 U3957 ( .A1(fract_i2f[36]), .A2(net85115), .ZN(n3245) );
  INV_X4 U3958 ( .A(n3245), .ZN(n3248) );
  NOR3_X4 U3959 ( .A1(n3248), .A2(n3247), .A3(n3246), .ZN(n3249) );
  NAND3_X4 U3960 ( .A1(n3251), .A2(n3250), .A3(n3249), .ZN(fract_denorm[36])
         );
  NAND4_X2 U3961 ( .A1(quo[37]), .A2(net85175), .A3(net85135), .A4(net85159), 
        .ZN(n3256) );
  AOI21_X4 U3962 ( .B1(n3254), .B2(quo[14]), .A(n3253), .ZN(n3255) );
  AOI22_X2 U3963 ( .A1(n3258), .A2(prod[38]), .B1(fract_i2f[38]), .B2(net85115), .ZN(n3264) );
  AOI21_X4 U3964 ( .B1(n3261), .B2(quo[17]), .A(n3260), .ZN(n3262) );
  NAND3_X4 U3965 ( .A1(n3262), .A2(n3263), .A3(n3264), .ZN(fract_denorm[38])
         );
  NAND3_X4 U3966 ( .A1(n3270), .A2(n3269), .A3(n3268), .ZN(fract_denorm[37])
         );
  NOR3_X4 U3967 ( .A1(n3278), .A2(n3277), .A3(n3276), .ZN(n3356) );
  NAND2_X2 U3968 ( .A1(prod[47]), .A2(net85167), .ZN(n3281) );
  MUX2_X2 U3969 ( .A(quo[26]), .B(quo[49]), .S(net94019), .Z(n3283) );
  INV_X4 U3970 ( .A(n3285), .ZN(n3340) );
  INV_X4 U3971 ( .A(n3286), .ZN(n3341) );
  INV_X4 U3972 ( .A(n3339), .ZN(n3289) );
  NOR2_X4 U3973 ( .A1(n2620), .A2(n2527), .ZN(n3288) );
  NAND2_X2 U3974 ( .A1(prod[7]), .A2(n2936), .ZN(n3293) );
  NAND2_X2 U3975 ( .A1(fract_i2f[7]), .A2(net85115), .ZN(n3292) );
  NAND2_X2 U3976 ( .A1(quo[9]), .A2(net86315), .ZN(n3291) );
  NAND3_X4 U3977 ( .A1(n3293), .A2(n3292), .A3(n3291), .ZN(n5323) );
  NAND2_X2 U3978 ( .A1(prod[8]), .A2(n2936), .ZN(n3296) );
  NAND2_X2 U3979 ( .A1(fract_i2f[8]), .A2(net85115), .ZN(n3295) );
  NAND2_X2 U3980 ( .A1(quo[10]), .A2(net86315), .ZN(n3294) );
  NAND3_X4 U3981 ( .A1(n3296), .A2(n3295), .A3(n3294), .ZN(net17690) );
  NAND2_X2 U3982 ( .A1(prod[10]), .A2(n2936), .ZN(n3299) );
  NAND2_X2 U3983 ( .A1(fract_i2f[10]), .A2(net85115), .ZN(n3298) );
  NAND3_X4 U3984 ( .A1(n3299), .A2(n3298), .A3(n3297), .ZN(n5324) );
  NAND2_X2 U3985 ( .A1(prod[9]), .A2(n2936), .ZN(n3302) );
  NAND2_X2 U3986 ( .A1(fract_i2f[9]), .A2(net85115), .ZN(n3301) );
  NAND2_X2 U3987 ( .A1(fract_i2f[12]), .A2(net85115), .ZN(n3304) );
  NAND3_X4 U3988 ( .A1(quo[14]), .A2(net84605), .A3(net85131), .ZN(n3303) );
  NAND3_X4 U3989 ( .A1(n3305), .A2(n3304), .A3(n3303), .ZN(n5326) );
  NAND2_X2 U3990 ( .A1(fract_i2f[11]), .A2(net85115), .ZN(n3307) );
  NAND3_X4 U3991 ( .A1(quo[13]), .A2(net84605), .A3(net85131), .ZN(n3306) );
  NAND3_X4 U3992 ( .A1(n3308), .A2(n3307), .A3(n3306), .ZN(net17655) );
  NAND2_X2 U3993 ( .A1(fract_i2f[14]), .A2(net85115), .ZN(n3310) );
  NAND3_X4 U3994 ( .A1(n3311), .A2(n3310), .A3(n3309), .ZN(net17656) );
  NAND2_X2 U3995 ( .A1(prod[16]), .A2(n2936), .ZN(n3314) );
  NAND2_X2 U3996 ( .A1(fract_i2f[16]), .A2(net85115), .ZN(n3313) );
  NAND3_X4 U3997 ( .A1(quo[18]), .A2(net84605), .A3(net85131), .ZN(n3312) );
  NAND3_X4 U3998 ( .A1(n3314), .A2(n3313), .A3(n3312), .ZN(net17684) );
  NAND2_X2 U3999 ( .A1(prod[15]), .A2(n2936), .ZN(n3317) );
  NAND2_X2 U4000 ( .A1(fract_i2f[15]), .A2(net85115), .ZN(n3316) );
  NAND3_X4 U4001 ( .A1(quo[17]), .A2(net84455), .A3(net85131), .ZN(n3315) );
  NAND3_X4 U4002 ( .A1(n3317), .A2(n3316), .A3(n3315), .ZN(net17685) );
  NAND2_X2 U4003 ( .A1(fract_i2f[13]), .A2(net85115), .ZN(net84444) );
  NAND2_X2 U4004 ( .A1(fract_i2f[4]), .A2(net85115), .ZN(n3319) );
  NAND2_X2 U4005 ( .A1(fract_i2f[5]), .A2(net85117), .ZN(n3322) );
  NAND2_X2 U4006 ( .A1(fract_i2f[6]), .A2(net85117), .ZN(n3325) );
  NAND2_X2 U4007 ( .A1(fract_i2f[1]), .A2(net85117), .ZN(n3328) );
  NAND2_X2 U4008 ( .A1(fract_i2f[2]), .A2(net85117), .ZN(n3331) );
  NAND3_X4 U4009 ( .A1(n3021), .A2(n3007), .A3(n3428), .ZN(n3389) );
  INV_X4 U4010 ( .A(n5323), .ZN(n3423) );
  INV_X4 U4011 ( .A(net17690), .ZN(net84188) );
  NOR2_X4 U4012 ( .A1(fract_denorm[21]), .A2(fract_denorm[22]), .ZN(n3350) );
  INV_X4 U4013 ( .A(net17684), .ZN(net84411) );
  NOR2_X4 U4014 ( .A1(fract_denorm[34]), .A2(fract_denorm[37]), .ZN(n3337) );
  NAND3_X4 U4015 ( .A1(n3337), .A2(n2975), .A3(net84172), .ZN(net83721) );
  NOR3_X4 U4016 ( .A1(n2620), .A2(n3341), .A3(n2527), .ZN(n3342) );
  NAND3_X4 U4017 ( .A1(n3343), .A2(n3022), .A3(n3342), .ZN(net84272) );
  NOR2_X4 U4018 ( .A1(fract_denorm[42]), .A2(fract_denorm[45]), .ZN(net84387)
         );
  NOR3_X4 U4019 ( .A1(n3359), .A2(fract_denorm[25]), .A3(n3612), .ZN(n3422) );
  INV_X4 U4020 ( .A(net95479), .ZN(net83636) );
  NOR2_X4 U4021 ( .A1(net84272), .A2(fract_denorm[33]), .ZN(n3349) );
  INV_X4 U4022 ( .A(net17682), .ZN(net84314) );
  INV_X4 U4023 ( .A(net17659), .ZN(net83622) );
  INV_X4 U4024 ( .A(n3409), .ZN(n3351) );
  NAND4_X2 U4025 ( .A1(net84341), .A2(net84321), .A3(net84314), .A4(n3663), 
        .ZN(n3352) );
  OAI21_X4 U4026 ( .B1(n3353), .B2(n3362), .A(n3352), .ZN(n3447) );
  INV_X4 U4027 ( .A(net17694), .ZN(net84364) );
  INV_X4 U4028 ( .A(net84363), .ZN(net83632) );
  NAND3_X4 U4029 ( .A1(net84345), .A2(net84262), .A3(n3357), .ZN(n3445) );
  AOI211_X4 U4030 ( .C1(net84343), .C2(n2959), .A(n3445), .B(n3358), .ZN(n3367) );
  INV_X4 U4031 ( .A(net28939), .ZN(net83714) );
  NAND2_X2 U4032 ( .A1(n3360), .A2(n3015), .ZN(n3361) );
  INV_X4 U4033 ( .A(n3361), .ZN(n3608) );
  INV_X4 U4034 ( .A(n3362), .ZN(n3363) );
  NAND3_X4 U4035 ( .A1(n3367), .A2(n3368), .A3(n3366), .ZN(u4_fi_ldz_2a_3_) );
  INV_X4 U4036 ( .A(n3369), .ZN(n3370) );
  INV_X4 U4037 ( .A(fract_denorm[33]), .ZN(net83715) );
  NAND2_X2 U4038 ( .A1(n2909), .A2(net84314), .ZN(n3410) );
  INV_X4 U4039 ( .A(n3410), .ZN(n3380) );
  INV_X4 U4040 ( .A(n3387), .ZN(n3394) );
  NAND2_X2 U4041 ( .A1(net84321), .A2(n3390), .ZN(net84261) );
  OAI221_X2 U4042 ( .B1(n3407), .B2(net92573), .C1(n3405), .C2(n3406), .A(
        n3404), .ZN(n3443) );
  NOR3_X4 U4043 ( .A1(n3412), .A2(n3447), .A3(n3445), .ZN(n3413) );
  NAND3_X4 U4044 ( .A1(n3415), .A2(n3414), .A3(n3413), .ZN(net83757) );
  NAND2_X2 U4045 ( .A1(n3421), .A2(n3420), .ZN(n3438) );
  INV_X4 U4046 ( .A(net84183), .ZN(net84182) );
  NAND2_X2 U4047 ( .A1(net84178), .A2(net84302), .ZN(n3426) );
  OAI211_X2 U4048 ( .C1(net92573), .C2(n3433), .A(n3432), .B(net84167), .ZN(
        n3434) );
  NOR3_X4 U4049 ( .A1(n3436), .A2(n3434), .A3(n3435), .ZN(n3437) );
  NAND3_X4 U4050 ( .A1(n3437), .A2(n3439), .A3(n3438), .ZN(net84158) );
  INV_X4 U4051 ( .A(n4758), .ZN(n4757) );
  NAND2_X2 U4052 ( .A1(fract_i2f[0]), .A2(net85117), .ZN(n3440) );
  INV_X4 U4054 ( .A(net84151), .ZN(net84149) );
  INV_X4 U4055 ( .A(net93777), .ZN(net84139) );
  INV_X4 U4056 ( .A(net84138), .ZN(u4_fi_ldz_mi1_5_) );
  XNOR2_X2 U4057 ( .A(n3449), .B(net86532), .ZN(u4_fi_ldz_mi1_4_) );
  XNOR2_X2 U4058 ( .A(net93777), .B(net83754), .ZN(u4_fi_ldz_mi1_2_) );
  OAI21_X4 U4059 ( .B1(net84128), .B2(n3451), .A(n3450), .ZN(n3452) );
  NAND2_X2 U4060 ( .A1(div_opa_ldz_r2[4]), .A2(net86532), .ZN(n3453) );
  OAI21_X4 U4061 ( .B1(n3456), .B2(n3454), .A(n3453), .ZN(net84124) );
  INV_X4 U4062 ( .A(net82991), .ZN(u4_ldz_all_6_) );
  XNOR2_X2 U4063 ( .A(div_opa_ldz_r2[4]), .B(net86532), .ZN(n3455) );
  XNOR2_X2 U4064 ( .A(net84116), .B(net84115), .ZN(u4_ldz_all_1_) );
  NAND3_X4 U4065 ( .A1(n3462), .A2(exp_r[4]), .A3(n3087), .ZN(n3460) );
  INV_X4 U4066 ( .A(n3585), .ZN(u4_f2i_shft_6_) );
  INV_X4 U4067 ( .A(net83941), .ZN(u4_f2i_shft_5_) );
  XNOR2_X2 U4068 ( .A(n3085), .B(n3461), .ZN(u4_f2i_shft_4_) );
  INV_X4 U4069 ( .A(n3463), .ZN(u4_f2i_shft_3_) );
  INV_X4 U4070 ( .A(net84101), .ZN(net84100) );
  INV_X4 U4071 ( .A(net17652), .ZN(net83633) );
  INV_X4 U4072 ( .A(net84091), .ZN(net84092) );
  INV_X4 U4073 ( .A(n3503), .ZN(n3465) );
  NAND2_X2 U4074 ( .A1(n2661), .A2(n3085), .ZN(n3487) );
  NOR2_X4 U4075 ( .A1(n3487), .A2(net82988), .ZN(n4751) );
  NAND2_X2 U4076 ( .A1(net85933), .A2(n4751), .ZN(n4747) );
  NAND2_X2 U4077 ( .A1(n3469), .A2(opas_r2), .ZN(n3468) );
  OAI21_X4 U4078 ( .B1(net84092), .B2(n3900), .A(n3468), .ZN(net82940) );
  INV_X4 U4079 ( .A(n3900), .ZN(n3470) );
  AOI22_X2 U4080 ( .A1(net84092), .A2(n3470), .B1(n3469), .B2(n2577), .ZN(
        net83350) );
  INV_X4 U4081 ( .A(u4_exp_in_pl1_1_), .ZN(net83865) );
  INV_X4 U4082 ( .A(u4_exp_next_mi_1_), .ZN(net83510) );
  INV_X4 U4083 ( .A(u4_exp_in_pl1_0_), .ZN(net84075) );
  INV_X4 U4084 ( .A(u4_exp_next_mi_0_), .ZN(n3805) );
  MUX2_X2 U4085 ( .A(net84075), .B(n3805), .S(net85393), .Z(n3597) );
  INV_X4 U4086 ( .A(u4_exp_in_pl1_4_), .ZN(n3474) );
  INV_X4 U4087 ( .A(u4_exp_next_mi_4_), .ZN(n3696) );
  INV_X4 U4088 ( .A(net83474), .ZN(net82856) );
  NAND2_X2 U4089 ( .A1(net86044), .A2(net83358), .ZN(n3764) );
  NAND2_X2 U4090 ( .A1(n3088), .A2(n2694), .ZN(net83903) );
  NAND2_X2 U4091 ( .A1(div_opa_ldz_r2[0]), .A2(net22501), .ZN(net83841) );
  INV_X4 U4092 ( .A(net83841), .ZN(net83862) );
  NAND2_X2 U4093 ( .A1(net83862), .A2(n3734), .ZN(n3478) );
  AOI21_X4 U4094 ( .B1(n3478), .B2(n2654), .A(net83858), .ZN(net83886) );
  NAND2_X2 U4095 ( .A1(n3089), .A2(n2691), .ZN(net83888) );
  NAND2_X2 U4096 ( .A1(div_opa_ldz_r2[2]), .A2(n3479), .ZN(net83887) );
  NAND2_X2 U4097 ( .A1(div_opa_ldz_r2[3]), .A2(n2579), .ZN(net83902) );
  NAND2_X2 U4098 ( .A1(div_opa_ldz_r2[4]), .A2(n2908), .ZN(net83919) );
  NAND2_X2 U4099 ( .A1(n3085), .A2(n2688), .ZN(net83918) );
  AOI22_X2 U4100 ( .A1(u4_div_exp1_5_), .A2(net83752), .B1(u4_div_exp3[5]), 
        .B2(net83749), .ZN(n3480) );
  INV_X4 U4101 ( .A(u4_exp_in_mi1_5_), .ZN(n3491) );
  NAND2_X2 U4102 ( .A1(n3764), .A2(net86028), .ZN(net82011) );
  INV_X4 U4103 ( .A(n3764), .ZN(n3975) );
  NAND2_X2 U4104 ( .A1(n3975), .A2(net86028), .ZN(net82013) );
  NOR2_X4 U4105 ( .A1(net82856), .A2(net83358), .ZN(n3530) );
  NAND2_X2 U4106 ( .A1(n3530), .A2(net86027), .ZN(n3604) );
  INV_X4 U4107 ( .A(n3604), .ZN(n4754) );
  INV_X4 U4108 ( .A(net83919), .ZN(net84032) );
  INV_X4 U4109 ( .A(net83887), .ZN(net84035) );
  OAI21_X4 U4110 ( .B1(net84035), .B2(net83886), .A(net83888), .ZN(n3548) );
  NAND2_X2 U4111 ( .A1(n3548), .A2(net83902), .ZN(n3482) );
  NAND2_X2 U4112 ( .A1(n3482), .A2(net83903), .ZN(n3483) );
  INV_X4 U4113 ( .A(n3483), .ZN(n3537) );
  OAI21_X4 U4114 ( .B1(net84032), .B2(n3537), .A(net83918), .ZN(n3528) );
  INV_X4 U4115 ( .A(n3528), .ZN(n3484) );
  NAND2_X2 U4116 ( .A1(n3484), .A2(net82988), .ZN(n3581) );
  INV_X4 U4117 ( .A(n3581), .ZN(n3485) );
  NAND4_X2 U4118 ( .A1(n3485), .A2(n2618), .A3(net83409), .A4(net83474), .ZN(
        n3989) );
  NOR3_X4 U4119 ( .A1(n3530), .A2(n3989), .A3(net86028), .ZN(n4755) );
  INV_X4 U4120 ( .A(n3530), .ZN(n3979) );
  NAND2_X2 U4121 ( .A1(n3989), .A2(n3979), .ZN(n3586) );
  INV_X4 U4122 ( .A(n3586), .ZN(n3486) );
  NAND2_X2 U4123 ( .A1(n3486), .A2(net86027), .ZN(n4749) );
  XNOR2_X2 U4124 ( .A(n3487), .B(net82988), .ZN(n3488) );
  AOI221_X2 U4125 ( .B1(u4_div_shft3_5_), .B2(n4754), .C1(u4_div_shft4[5]), 
        .C2(n4755), .A(n3489), .ZN(n3490) );
  OAI221_X2 U4126 ( .B1(n3491), .B2(net82011), .C1(net83535), .C2(net82013), 
        .A(n3490), .ZN(u4_shift_right[5]) );
  AOI22_X2 U4127 ( .A1(u4_exp_f2i_1[53]), .A2(n2652), .B1(n1373), .B2(n3492), 
        .ZN(n3497) );
  AOI22_X2 U4128 ( .A1(u4_div_exp1_4_), .A2(net83752), .B1(u4_div_exp3[4]), 
        .B2(net83749), .ZN(net84018) );
  NAND2_X2 U4129 ( .A1(net86027), .A2(net83019), .ZN(n3496) );
  NAND3_X4 U4130 ( .A1(n3497), .A2(n3496), .A3(net84013), .ZN(u4_exp_out_4_)
         );
  INV_X4 U4131 ( .A(u4_exp_in_mi1_4_), .ZN(n3501) );
  XNOR2_X2 U4132 ( .A(n3085), .B(n2661), .ZN(n3498) );
  AOI221_X2 U4133 ( .B1(u4_div_shft4[4]), .B2(n4755), .C1(u4_div_shft3_4_), 
        .C2(n4754), .A(n3499), .ZN(n3500) );
  OAI221_X2 U4134 ( .B1(n3501), .B2(net82011), .C1(net83596), .C2(net82013), 
        .A(n3500), .ZN(u4_shift_right[4]) );
  AOI22_X2 U4135 ( .A1(u4_div_exp1_3_), .A2(net83752), .B1(u4_div_exp3[3]), 
        .B2(net83749), .ZN(net84003) );
  INV_X4 U4136 ( .A(net82013), .ZN(net23104) );
  INV_X4 U4137 ( .A(net82011), .ZN(net23097) );
  NAND2_X2 U4138 ( .A1(n2656), .A2(net23097), .ZN(n3507) );
  XNOR2_X2 U4139 ( .A(n3503), .B(n2579), .ZN(n3504) );
  AOI221_X2 U4140 ( .B1(u4_div_shft3_3_), .B2(n4754), .C1(u4_div_shft4[3]), 
        .C2(n4755), .A(n3505), .ZN(n3506) );
  AOI22_X2 U4141 ( .A1(u4_exp_f2i_1[51]), .A2(n2652), .B1(n1373), .B2(n2948), 
        .ZN(net83971) );
  AOI22_X2 U4142 ( .A1(u4_div_exp1_2_), .A2(net83752), .B1(u4_div_exp3[2]), 
        .B2(net83749), .ZN(n3512) );
  INV_X4 U4143 ( .A(u4_exp_in_mi1_2_), .ZN(n3516) );
  INV_X4 U4144 ( .A(u4_exp_out_2_), .ZN(net83599) );
  INV_X4 U4145 ( .A(n4749), .ZN(n4753) );
  AOI221_X2 U4146 ( .B1(u4_div_shft4[2]), .B2(n4755), .C1(u4_div_shft3_2_), 
        .C2(n4754), .A(n2529), .ZN(n3515) );
  OAI221_X2 U4147 ( .B1(n3516), .B2(net82011), .C1(net83599), .C2(net82013), 
        .A(n3515), .ZN(u4_shift_right[2]) );
  NAND2_X2 U4148 ( .A1(net82776), .A2(net86028), .ZN(net83356) );
  INV_X4 U4149 ( .A(n3597), .ZN(n3599) );
  AOI22_X2 U4150 ( .A1(u4_div_exp1_1_), .A2(net83752), .B1(u4_div_exp3[1]), 
        .B2(net83749), .ZN(net83959) );
  NAND3_X4 U4151 ( .A1(n3518), .A2(n3519), .A3(net83953), .ZN(u4_exp_out_1_)
         );
  INV_X4 U4152 ( .A(u4_exp_in_mi1_1_), .ZN(n3576) );
  OAI221_X2 U4153 ( .B1(n3576), .B2(net82011), .C1(net83507), .C2(net82013), 
        .A(n3520), .ZN(u4_shift_right[1]) );
  NAND2_X2 U4154 ( .A1(n4753), .A2(net85905), .ZN(n3523) );
  NAND2_X2 U4155 ( .A1(u4_div_shft3_0_), .A2(n4754), .ZN(n3522) );
  NAND2_X2 U4156 ( .A1(u4_div_shft4[0]), .A2(n4755), .ZN(n3521) );
  NAND4_X2 U4157 ( .A1(n3523), .A2(n3522), .A3(n3521), .A4(n1416), .ZN(
        u4_shift_right[0]) );
  INV_X4 U4158 ( .A(u4_exp_in_pl1_8_), .ZN(n3524) );
  MUX2_X2 U4159 ( .A(n3524), .B(net83948), .S(net85393), .Z(net83824) );
  INV_X4 U4160 ( .A(net83824), .ZN(net82036) );
  NAND2_X2 U4161 ( .A1(n3525), .A2(net86045), .ZN(n3568) );
  NAND2_X2 U4162 ( .A1(net82035), .A2(n3568), .ZN(n3562) );
  NAND2_X2 U4163 ( .A1(net86032), .A2(net83233), .ZN(net82034) );
  INV_X4 U4164 ( .A(net82034), .ZN(net83735) );
  NAND2_X2 U4165 ( .A1(net83735), .A2(net83041), .ZN(net83837) );
  INV_X4 U4166 ( .A(net83837), .ZN(net83933) );
  INV_X4 U4167 ( .A(n3526), .ZN(n3947) );
  NAND3_X4 U4168 ( .A1(net83933), .A2(n3527), .A3(net86045), .ZN(net83823) );
  NAND2_X2 U4169 ( .A1(u4_exp_in_pl1_5_), .A2(n3582), .ZN(net83943) );
  NAND2_X2 U4170 ( .A1(net85929), .A2(n3528), .ZN(n3533) );
  NOR2_X4 U4171 ( .A1(n3530), .A2(n3529), .ZN(n3531) );
  NAND2_X2 U4172 ( .A1(net82036), .A2(net83358), .ZN(net83869) );
  INV_X4 U4173 ( .A(net83869), .ZN(net83925) );
  OAI21_X4 U4174 ( .B1(net83925), .B2(net83870), .A(net83926), .ZN(net83878)
         );
  INV_X4 U4175 ( .A(net83878), .ZN(net83924) );
  INV_X4 U4176 ( .A(n3536), .ZN(u4_shift_left[5]) );
  NAND2_X2 U4177 ( .A1(net83918), .A2(net83919), .ZN(n3539) );
  XNOR2_X2 U4178 ( .A(div_opa_ldz_r2[4]), .B(n3085), .ZN(n3538) );
  MUX2_X2 U4179 ( .A(n3539), .B(n3538), .S(n3537), .Z(n3544) );
  NAND2_X2 U4180 ( .A1(net83878), .A2(net86532), .ZN(n3540) );
  INV_X4 U4181 ( .A(n3540), .ZN(n3543) );
  NAND2_X2 U4182 ( .A1(u4_f2i_shft_4_), .A2(net83113), .ZN(n3546) );
  AOI22_X2 U4183 ( .A1(net83846), .A2(n3085), .B1(u4_exp_in_pl1_4_), .B2(n3582), .ZN(n3545) );
  XNOR2_X2 U4184 ( .A(div_opa_ldz_r2[3]), .B(n3087), .ZN(n3550) );
  NAND2_X2 U4185 ( .A1(net83902), .A2(net83903), .ZN(n3549) );
  MUX2_X2 U4186 ( .A(n3550), .B(n3549), .S(n3548), .Z(n3552) );
  AOI211_X4 U4187 ( .C1(net83854), .C2(n3552), .A(n2663), .B(n3551), .ZN(n3555) );
  NAND2_X2 U4188 ( .A1(u4_f2i_shft_3_), .A2(net83113), .ZN(n3554) );
  AOI22_X2 U4189 ( .A1(net83846), .A2(n3088), .B1(u4_exp_in_pl1_3_), .B2(n3582), .ZN(n3553) );
  NAND3_X4 U4190 ( .A1(n3555), .A2(n3554), .A3(n3553), .ZN(u4_shift_left[3])
         );
  NAND2_X2 U4191 ( .A1(net83887), .A2(net83888), .ZN(n3557) );
  XNOR2_X2 U4192 ( .A(div_opa_ldz_r2[2]), .B(n3089), .ZN(n3556) );
  MUX2_X2 U4193 ( .A(n3557), .B(n3556), .S(net83886), .Z(n3561) );
  INV_X4 U4194 ( .A(n3562), .ZN(n3563) );
  NAND2_X2 U4195 ( .A1(n3563), .A2(u4_exp_in_pl1_2_), .ZN(n3565) );
  AOI22_X2 U4196 ( .A1(u4_f2i_shft_2_), .A2(net82938), .B1(net83846), .B2(
        n3089), .ZN(n3564) );
  NAND4_X2 U4197 ( .A1(n3567), .A2(n3566), .A3(n3565), .A4(n3564), .ZN(
        u4_shift_left[2]) );
  NAND2_X2 U4198 ( .A1(n3569), .A2(n3568), .ZN(n3580) );
  NAND2_X2 U4199 ( .A1(net86045), .A2(net83865), .ZN(n3574) );
  INV_X4 U4200 ( .A(net83863), .ZN(net83851) );
  NAND2_X2 U4201 ( .A1(div_opa_ldz_r2[1]), .A2(n3734), .ZN(n3571) );
  MUX2_X2 U4202 ( .A(n3571), .B(n3570), .S(net83862), .Z(n3572) );
  NAND2_X2 U4203 ( .A1(n3572), .A2(net83857), .ZN(n3573) );
  AOI211_X4 U4204 ( .C1(n3575), .C2(n3574), .A(net83851), .B(n2533), .ZN(n3579) );
  OAI21_X4 U4205 ( .B1(net83811), .B2(n3584), .A(n3583), .ZN(net83799) );
  NAND2_X2 U4206 ( .A1(net82035), .A2(net85901), .ZN(net82040) );
  INV_X4 U4207 ( .A(net82040), .ZN(net82952) );
  NOR2_X4 U4208 ( .A1(n3588), .A2(n3587), .ZN(net83797) );
  NAND2_X2 U4209 ( .A1(u4_N1405), .A2(net85377), .ZN(n3589) );
  INV_X4 U4210 ( .A(n2069), .ZN(u4_fract_out_14_) );
  INV_X4 U4211 ( .A(n2083), .ZN(u4_fract_out_6_) );
  INV_X4 U4212 ( .A(n2952), .ZN(u4_fract_out_2_) );
  INV_X4 U4213 ( .A(n2091), .ZN(u4_fract_out_1_) );
  INV_X4 U4214 ( .A(n2093), .ZN(u4_fract_out_0_) );
  INV_X4 U4215 ( .A(u4_exp_in_pl1_6_), .ZN(net83791) );
  INV_X4 U4216 ( .A(net83761), .ZN(net83773) );
  AOI22_X2 U4217 ( .A1(u4_div_exp1_6_), .A2(net83752), .B1(u4_div_exp3[6]), 
        .B2(net83749), .ZN(n3590) );
  NAND3_X4 U4218 ( .A1(n3591), .A2(n3593), .A3(n3592), .ZN(u4_exp_out_6_) );
  INV_X4 U4219 ( .A(net86532), .ZN(net83579) );
  INV_X4 U4220 ( .A(n3596), .ZN(n3595) );
  OAI21_X4 U4221 ( .B1(net83579), .B2(n3595), .A(net83761), .ZN(n3594) );
  INV_X4 U4222 ( .A(n3594), .ZN(u4_fi_ldz_mi22[6]) );
  XNOR2_X2 U4223 ( .A(n3595), .B(net86532), .ZN(u4_fi_ldz_mi22[4]) );
  NAND2_X2 U4224 ( .A1(n3596), .A2(net83756), .ZN(u4_fi_ldz_mi22[3]) );
  INV_X4 U4225 ( .A(net83750), .ZN(net83747) );
  AOI22_X2 U4226 ( .A1(net83747), .A2(n3597), .B1(u4_div_exp3[0]), .B2(
        net83749), .ZN(n3598) );
  NAND2_X2 U4227 ( .A1(n1373), .A2(n3599), .ZN(n3601) );
  NAND2_X2 U4228 ( .A1(u4_exp_f2i_1[49]), .A2(n2652), .ZN(n3600) );
  NAND2_X2 U4229 ( .A1(net95357), .A2(net83593), .ZN(n4756) );
  NOR3_X4 U4230 ( .A1(n3602), .A2(u4_fract_out_19_), .A3(u4_fract_out_17_), 
        .ZN(net83724) );
  NOR3_X4 U4231 ( .A1(n3603), .A2(u4_fract_out_10_), .A3(n2245), .ZN(net83725)
         );
  INV_X4 U4232 ( .A(u4_div_shft3_1_), .ZN(n3610) );
  INV_X4 U4233 ( .A(u4_div_shft3_0_), .ZN(n3609) );
  NOR2_X4 U4234 ( .A1(n3610), .A2(n3609), .ZN(n3611) );
  NOR4_X2 U4235 ( .A1(u4_div_shft3_7_), .A2(u4_div_shft3_6_), .A3(
        u4_div_shft3_5_), .A4(n2606), .ZN(n3613) );
  NOR2_X4 U4236 ( .A1(n2278), .A2(n3616), .ZN(n3677) );
  NOR3_X4 U4237 ( .A1(remainder[21]), .A2(remainder[20]), .A3(remainder[19]), 
        .ZN(n3618) );
  NAND4_X2 U4238 ( .A1(n3620), .A2(n3619), .A3(n3618), .A4(n3617), .ZN(n3628)
         );
  NOR3_X4 U4239 ( .A1(remainder[9]), .A2(remainder[8]), .A3(remainder[7]), 
        .ZN(n3622) );
  NOR3_X4 U4240 ( .A1(remainder[12]), .A2(remainder[11]), .A3(remainder[10]), 
        .ZN(n3621) );
  NAND2_X2 U4241 ( .A1(n3622), .A2(n3621), .ZN(n3627) );
  NOR2_X4 U4242 ( .A1(remainder[5]), .A2(remainder[4]), .ZN(n3623) );
  NAND4_X2 U4243 ( .A1(n3625), .A2(n3624), .A3(n3623), .A4(n2732), .ZN(n3626)
         );
  NOR3_X4 U4244 ( .A1(n3628), .A2(n3627), .A3(n3626), .ZN(n3642) );
  NOR3_X4 U4245 ( .A1(remainder[40]), .A2(remainder[39]), .A3(remainder[38]), 
        .ZN(n3632) );
  NOR3_X4 U4246 ( .A1(remainder[43]), .A2(remainder[42]), .A3(remainder[41]), 
        .ZN(n3631) );
  NOR3_X4 U4247 ( .A1(remainder[46]), .A2(remainder[45]), .A3(remainder[44]), 
        .ZN(n3630) );
  NOR3_X4 U4248 ( .A1(remainder[49]), .A2(remainder[48]), .A3(remainder[47]), 
        .ZN(n3629) );
  NAND4_X2 U4249 ( .A1(n3632), .A2(n3631), .A3(n3630), .A4(n3629), .ZN(n3640)
         );
  NOR3_X4 U4250 ( .A1(remainder[34]), .A2(remainder[33]), .A3(remainder[32]), 
        .ZN(n3634) );
  NOR3_X4 U4251 ( .A1(remainder[37]), .A2(remainder[36]), .A3(remainder[35]), 
        .ZN(n3633) );
  NAND2_X2 U4252 ( .A1(n3634), .A2(n3633), .ZN(n3639) );
  NOR2_X4 U4253 ( .A1(remainder[30]), .A2(remainder[29]), .ZN(n3635) );
  NAND4_X2 U4254 ( .A1(n3637), .A2(n3636), .A3(n3635), .A4(n2733), .ZN(n3638)
         );
  NOR3_X4 U4255 ( .A1(n3640), .A2(n3639), .A3(n3638), .ZN(n3641) );
  NAND2_X2 U4256 ( .A1(n3642), .A2(n3641), .ZN(n3978) );
  NAND2_X2 U4257 ( .A1(u4_N1977), .A2(net86032), .ZN(n3646) );
  NOR2_X4 U4258 ( .A1(n3645), .A2(n3644), .ZN(n3662) );
  NAND4_X2 U4259 ( .A1(n3650), .A2(n3649), .A3(n3648), .A4(n3647), .ZN(n3656)
         );
  NOR3_X4 U4260 ( .A1(u4_N1424), .A2(u4_N1423), .A3(u4_N1425), .ZN(n3652) );
  NAND4_X2 U4261 ( .A1(n2264), .A2(n2265), .A3(n2266), .A4(n2267), .ZN(n3658)
         );
  NAND4_X2 U4262 ( .A1(n2260), .A2(n2261), .A3(n2262), .A4(n2263), .ZN(n3657)
         );
  NAND2_X2 U4263 ( .A1(net83632), .A2(net83633), .ZN(n3664) );
  NOR3_X4 U4264 ( .A1(n3667), .A2(net83620), .A3(net83621), .ZN(n3668) );
  NAND3_X4 U4265 ( .A1(net83616), .A2(n3669), .A3(n3668), .ZN(n3670) );
  NAND2_X2 U4266 ( .A1(net83569), .A2(net83565), .ZN(net83396) );
  NAND2_X2 U4267 ( .A1(net83599), .A2(net83507), .ZN(n3678) );
  INV_X4 U4268 ( .A(n3678), .ZN(n3704) );
  NAND2_X2 U4269 ( .A1(n2585), .A2(n3745), .ZN(net83527) );
  INV_X4 U4270 ( .A(n3713), .ZN(n3680) );
  INV_X4 U4271 ( .A(n3789), .ZN(n3702) );
  NAND2_X2 U4272 ( .A1(net95357), .A2(net83593), .ZN(n3701) );
  NAND2_X2 U4273 ( .A1(n3702), .A2(n3701), .ZN(net83591) );
  INV_X4 U4274 ( .A(net83591), .ZN(net83383) );
  INV_X4 U4275 ( .A(net82931), .ZN(net82929) );
  INV_X4 U4276 ( .A(n4747), .ZN(n3681) );
  NAND2_X2 U4277 ( .A1(n3681), .A2(net85905), .ZN(n3962) );
  INV_X4 U4278 ( .A(n3962), .ZN(n3682) );
  NAND2_X2 U4279 ( .A1(n3682), .A2(net85937), .ZN(net83408) );
  NOR2_X4 U4280 ( .A1(n3998), .A2(net83408), .ZN(n3683) );
  NAND3_X4 U4281 ( .A1(n3684), .A2(n2900), .A3(n3683), .ZN(n3688) );
  INV_X4 U4282 ( .A(n3685), .ZN(n3686) );
  NAND2_X2 U4283 ( .A1(net83036), .A2(net86027), .ZN(n3793) );
  INV_X4 U4284 ( .A(n3793), .ZN(n3689) );
  INV_X4 U4285 ( .A(n3688), .ZN(n3695) );
  INV_X4 U4286 ( .A(n3690), .ZN(n3693) );
  INV_X4 U4287 ( .A(u4_fi_ldz_2a_6_), .ZN(n3755) );
  INV_X4 U4288 ( .A(u4_exp_fix_diva[4]), .ZN(n3691) );
  INV_X4 U4289 ( .A(u4_exp_fix_divb[4]), .ZN(n3694) );
  NAND3_X4 U4290 ( .A1(n3695), .A2(net83036), .A3(net86028), .ZN(net83316) );
  NOR3_X4 U4291 ( .A1(n3699), .A2(n3698), .A3(n3697), .ZN(n3705) );
  NAND2_X2 U4292 ( .A1(n3704), .A2(net83368), .ZN(n3744) );
  INV_X4 U4293 ( .A(u4_exp_fix_divb[2]), .ZN(n3707) );
  NOR2_X4 U4294 ( .A1(net83431), .A2(n3707), .ZN(n3712) );
  INV_X4 U4295 ( .A(u4_exp_fix_diva[2]), .ZN(n3709) );
  NOR3_X4 U4296 ( .A1(n3712), .A2(n3711), .A3(n3710), .ZN(n3722) );
  NAND2_X2 U4297 ( .A1(u4_exp_out_pl1_2_), .A2(net83435), .ZN(n3721) );
  NAND2_X2 U4298 ( .A1(n3744), .A2(n3713), .ZN(n3717) );
  NAND2_X2 U4299 ( .A1(net82929), .A2(n3089), .ZN(n3714) );
  NAND3_X2 U4300 ( .A1(n3718), .A2(n2502), .A3(net83526), .ZN(n3736) );
  NAND4_X2 U4301 ( .A1(n3722), .A2(n3721), .A3(n3720), .A4(n3719), .ZN(n3827)
         );
  NAND2_X2 U4302 ( .A1(n3823), .A2(n3827), .ZN(n3731) );
  NAND2_X2 U4303 ( .A1(u4_exp_fix_diva[5]), .A2(net83312), .ZN(n3725) );
  INV_X4 U4304 ( .A(net83316), .ZN(net83532) );
  NAND2_X2 U4305 ( .A1(u4_exp_fix_divb[5]), .A2(net95605), .ZN(n3723) );
  NAND2_X2 U4306 ( .A1(u4_exp_out_pl1_5_), .A2(net83435), .ZN(n3726) );
  NOR2_X4 U4307 ( .A1(n3730), .A2(n3729), .ZN(n3825) );
  NAND2_X2 U4308 ( .A1(net83383), .A2(n2659), .ZN(net83348) );
  INV_X4 U4309 ( .A(net83428), .ZN(net83312) );
  INV_X4 U4310 ( .A(net83495), .ZN(net83492) );
  INV_X4 U4311 ( .A(n3744), .ZN(n3745) );
  NAND2_X2 U4312 ( .A1(u4_exp_out_pl1_3_), .A2(net83435), .ZN(n3749) );
  NAND2_X2 U4313 ( .A1(n3749), .A2(n3748), .ZN(n3750) );
  NOR2_X4 U4314 ( .A1(n2626), .A2(n3750), .ZN(n3751) );
  INV_X4 U4315 ( .A(net83408), .ZN(net83030) );
  NAND2_X2 U4316 ( .A1(net83030), .A2(n3755), .ZN(net83367) );
  INV_X4 U4317 ( .A(u4_div_exp1_5_), .ZN(n3757) );
  INV_X4 U4318 ( .A(u4_div_exp1_4_), .ZN(n3756) );
  NOR2_X4 U4319 ( .A1(n3757), .A2(n3756), .ZN(n3762) );
  INV_X4 U4320 ( .A(u4_div_exp1_3_), .ZN(n3760) );
  INV_X4 U4321 ( .A(u4_div_exp1_2_), .ZN(n3759) );
  INV_X4 U4322 ( .A(u4_div_exp1_0_), .ZN(net83468) );
  INV_X4 U4323 ( .A(u4_div_exp1_1_), .ZN(n3758) );
  NOR4_X2 U4324 ( .A1(n3760), .A2(n3759), .A3(net83468), .A4(n3758), .ZN(n3761) );
  NAND3_X4 U4325 ( .A1(n3781), .A2(net83381), .A3(net83463), .ZN(n3792) );
  INV_X4 U4326 ( .A(n3792), .ZN(n3785) );
  INV_X4 U4327 ( .A(n3763), .ZN(n3765) );
  NAND2_X2 U4328 ( .A1(n3785), .A2(n3766), .ZN(net83404) );
  NAND2_X2 U4329 ( .A1(opb_00), .A2(net82035), .ZN(net83248) );
  NAND2_X2 U4330 ( .A1(opb_inf), .A2(net86027), .ZN(net83045) );
  NAND2_X2 U4331 ( .A1(n3767), .A2(n3785), .ZN(net83297) );
  NAND2_X2 U4332 ( .A1(u4_exp_out_pl1_6_), .A2(net83435), .ZN(n3776) );
  INV_X4 U4333 ( .A(net83434), .ZN(net83433) );
  INV_X4 U4334 ( .A(u4_exp_fix_divb[6]), .ZN(n3768) );
  NOR2_X4 U4335 ( .A1(net83431), .A2(n3768), .ZN(n3772) );
  INV_X4 U4336 ( .A(u4_exp_fix_diva[6]), .ZN(n3769) );
  NOR2_X4 U4337 ( .A1(net83428), .A2(n3769), .ZN(n3770) );
  NAND2_X2 U4338 ( .A1(exp_ovf_r_0_), .A2(net85901), .ZN(net82925) );
  INV_X4 U4339 ( .A(u4_fract_out_pl1_0_), .ZN(n3777) );
  NAND2_X2 U4340 ( .A1(n2910), .A2(net83276), .ZN(n3780) );
  INV_X4 U4341 ( .A(n3780), .ZN(n3795) );
  INV_X4 U4342 ( .A(net82957), .ZN(net82927) );
  NAND2_X2 U4343 ( .A1(net85937), .A2(net83385), .ZN(net83384) );
  NAND2_X2 U4344 ( .A1(exp_ovf_r_0_), .A2(net83030), .ZN(net83369) );
  INV_X4 U4345 ( .A(n4006), .ZN(n3783) );
  OAI21_X4 U4346 ( .B1(n3784), .B2(n3783), .A(n2710), .ZN(net83375) );
  INV_X4 U4347 ( .A(net83375), .ZN(net83370) );
  NAND2_X2 U4348 ( .A1(n3785), .A2(net83373), .ZN(net83371) );
  INV_X4 U4349 ( .A(n3799), .ZN(n3821) );
  NAND2_X2 U4350 ( .A1(n3821), .A2(net83359), .ZN(n3819) );
  NAND2_X2 U4351 ( .A1(n3819), .A2(net83358), .ZN(n3801) );
  INV_X4 U4352 ( .A(net82925), .ZN(net83338) );
  NAND3_X2 U4353 ( .A1(net83338), .A2(net83356), .A3(net83357), .ZN(n3791) );
  OAI21_X4 U4354 ( .B1(n3793), .B2(n3792), .A(n3791), .ZN(n3794) );
  INV_X4 U4355 ( .A(n3794), .ZN(n3798) );
  OAI21_X4 U4356 ( .B1(n2525), .B2(n3801), .A(n3798), .ZN(n4002) );
  INV_X4 U4357 ( .A(n4002), .ZN(n4007) );
  INV_X4 U4358 ( .A(n4003), .ZN(n3817) );
  INV_X4 U4359 ( .A(net83348), .ZN(net83344) );
  NAND2_X2 U4360 ( .A1(net83338), .A2(net83234), .ZN(n3995) );
  INV_X4 U4361 ( .A(n3995), .ZN(n3797) );
  NAND2_X2 U4362 ( .A1(n3797), .A2(net86027), .ZN(n3816) );
  INV_X4 U4363 ( .A(net83328), .ZN(net83327) );
  OAI21_X4 U4364 ( .B1(n3803), .B2(n2575), .A(n2673), .ZN(n4118) );
  AOI22_X2 U4365 ( .A1(u4_exp_fix_diva[0]), .A2(net83312), .B1(
        u4_exp_fix_divb[0]), .B2(net95605), .ZN(n3810) );
  AND4_X2 U4366 ( .A1(n3811), .A2(n3810), .A3(n3809), .A4(n3808), .ZN(n3812)
         );
  OAI21_X4 U4367 ( .B1(n3814), .B2(n2658), .A(n3813), .ZN(net83068) );
  NAND2_X2 U4368 ( .A1(net83300), .A2(net86032), .ZN(n3815) );
  INV_X4 U4369 ( .A(n3815), .ZN(n3818) );
  INV_X4 U4370 ( .A(net83295), .ZN(net83220) );
  NOR2_X4 U4371 ( .A1(net83288), .A2(n3820), .ZN(n3822) );
  OAI22_X2 U4372 ( .A1(n2747), .A2(n3820), .B1(n3820), .B2(n3819), .ZN(n3824)
         );
  OAI21_X4 U4373 ( .B1(net83274), .B2(n3824), .A(net83275), .ZN(n3829) );
  OAI21_X4 U4374 ( .B1(net86486), .B2(n2574), .A(n2673), .ZN(n4121) );
  OAI21_X4 U4375 ( .B1(n3829), .B2(n3826), .A(n2673), .ZN(n4120) );
  OAI21_X4 U4376 ( .B1(n3829), .B2(n2573), .A(n2673), .ZN(net82764) );
  INV_X4 U4377 ( .A(net83264), .ZN(net83263) );
  OAI21_X4 U4378 ( .B1(net86486), .B2(n2576), .A(n2673), .ZN(n3950) );
  OAI21_X4 U4379 ( .B1(n3829), .B2(n2572), .A(n2673), .ZN(net82762) );
  NOR3_X4 U4380 ( .A1(net83254), .A2(n3950), .A3(net82762), .ZN(n3830) );
  NAND2_X2 U4381 ( .A1(opb_00), .A2(opa_00), .ZN(n3902) );
  INV_X4 U4382 ( .A(n3902), .ZN(n3941) );
  NAND2_X2 U4383 ( .A1(n3941), .A2(net86027), .ZN(n3837) );
  INV_X4 U4384 ( .A(net83248), .ZN(net83247) );
  NAND2_X2 U4385 ( .A1(net83247), .A2(opa_inf), .ZN(n3836) );
  NAND2_X2 U4386 ( .A1(opb_inf), .A2(opa_00), .ZN(n3906) );
  INV_X4 U4387 ( .A(n3906), .ZN(n3834) );
  NAND2_X2 U4388 ( .A1(n2736), .A2(n2607), .ZN(net82829) );
  INV_X4 U4389 ( .A(net82829), .ZN(net83070) );
  NAND2_X2 U4390 ( .A1(ind_d), .A2(n2738), .ZN(n4070) );
  NAND2_X2 U4391 ( .A1(net83070), .A2(n4070), .ZN(n3833) );
  MUX2_X2 U4392 ( .A(n3838), .B(n2735), .S(net86027), .Z(n3840) );
  NAND2_X2 U4393 ( .A1(n2737), .A2(n2605), .ZN(n3942) );
  NAND2_X2 U4394 ( .A1(net83234), .A2(n3942), .ZN(n3944) );
  MUX2_X2 U4395 ( .A(n2773), .B(n4728), .S(net82757), .Z(N445) );
  INV_X4 U4396 ( .A(u4_fract_out_pl1_1_), .ZN(n3841) );
  INV_X4 U4397 ( .A(net82762), .ZN(net83064) );
  INV_X4 U4398 ( .A(n4120), .ZN(n3930) );
  INV_X4 U4399 ( .A(n3950), .ZN(n4119) );
  INV_X4 U4400 ( .A(net82876), .ZN(net83197) );
  INV_X4 U4401 ( .A(u4_fract_out_pl1_4_), .ZN(n3849) );
  INV_X4 U4402 ( .A(n3850), .ZN(n3851) );
  INV_X4 U4403 ( .A(u4_fract_out_pl1_2_), .ZN(n3853) );
  INV_X4 U4404 ( .A(u4_fract_out_pl1_3_), .ZN(n3855) );
  INV_X4 U4405 ( .A(u4_fract_out_pl1_20_), .ZN(n3858) );
  INV_X4 U4406 ( .A(u4_fract_out_pl1_19_), .ZN(n3860) );
  INV_X4 U4407 ( .A(u4_fract_out_pl1_18_), .ZN(n3862) );
  NAND3_X4 U4408 ( .A1(n4027), .A2(n3870), .A3(n3869), .ZN(net83115) );
  INV_X4 U4409 ( .A(u4_fract_out_pl1_11_), .ZN(net83168) );
  INV_X4 U4410 ( .A(u4_fract_out_pl1_10_), .ZN(n3871) );
  INV_X4 U4411 ( .A(u4_fract_out_pl1_12_), .ZN(n3875) );
  INV_X4 U4412 ( .A(u4_fract_out_pl1_6_), .ZN(n3877) );
  INV_X4 U4413 ( .A(u4_fract_out_pl1_8_), .ZN(n3878) );
  INV_X4 U4414 ( .A(u4_fract_out_pl1_7_), .ZN(n3883) );
  INV_X4 U4415 ( .A(u4_fract_out_pl1_14_), .ZN(n3885) );
  NOR2_X4 U4416 ( .A1(net83126), .A2(n3885), .ZN(n3886) );
  INV_X4 U4417 ( .A(n3886), .ZN(n3887) );
  INV_X4 U4418 ( .A(u4_fract_out_pl1_15_), .ZN(n3889) );
  INV_X4 U4419 ( .A(u4_fract_out_pl1_17_), .ZN(n3891) );
  INV_X4 U4420 ( .A(u4_fract_out_pl1_16_), .ZN(n3896) );
  NOR2_X4 U4421 ( .A1(net83126), .A2(n3896), .ZN(n3897) );
  NAND2_X2 U4422 ( .A1(n3901), .A2(n3900), .ZN(net83109) );
  NAND2_X2 U4423 ( .A1(net83070), .A2(net86027), .ZN(n3935) );
  INV_X4 U4424 ( .A(n3935), .ZN(n3909) );
  NAND2_X2 U4425 ( .A1(n3903), .A2(n3902), .ZN(n3904) );
  MUX2_X2 U4426 ( .A(n3904), .B(n3903), .S(sign_mul_r), .Z(n3905) );
  NAND2_X2 U4427 ( .A1(n3909), .A2(n3905), .ZN(n3915) );
  NAND2_X2 U4428 ( .A1(opb_00), .A2(opa_inf), .ZN(n3907) );
  NAND2_X2 U4429 ( .A1(n3907), .A2(n3906), .ZN(n3943) );
  NAND2_X2 U4430 ( .A1(sign_exe_r), .A2(n3943), .ZN(n3908) );
  XNOR2_X2 U4431 ( .A(sign_mul_r), .B(n3908), .ZN(n3913) );
  NAND2_X2 U4432 ( .A1(net83070), .A2(n2731), .ZN(n3933) );
  INV_X4 U4433 ( .A(n3933), .ZN(n3910) );
  AOI22_X2 U4434 ( .A1(n3913), .A2(n2684), .B1(n3912), .B2(n3911), .ZN(n3914)
         );
  NAND2_X2 U4435 ( .A1(n3916), .A2(net83090), .ZN(n3938) );
  NAND4_X2 U4436 ( .A1(n2958), .A2(n3919), .A3(n2460), .A4(n2549), .ZN(n3924)
         );
  NAND4_X2 U4437 ( .A1(net82891), .A2(n4028), .A3(n4024), .A4(n2904), .ZN(
        n3923) );
  INV_X4 U4438 ( .A(net82807), .ZN(net82893) );
  NAND2_X2 U4439 ( .A1(net83070), .A2(n2709), .ZN(net82767) );
  NAND2_X2 U4440 ( .A1(n3932), .A2(n3931), .ZN(net83061) );
  NAND4_X2 U4441 ( .A1(n3936), .A2(net92392), .A3(n3935), .A4(n3934), .ZN(
        n3937) );
  NAND2_X2 U4442 ( .A1(n3938), .A2(n3937), .ZN(N495) );
  NAND2_X2 U4443 ( .A1(net86027), .A2(n2698), .ZN(n3940) );
  INV_X4 U4444 ( .A(n3942), .ZN(n4110) );
  NAND2_X2 U4445 ( .A1(net83036), .A2(n3942), .ZN(n4014) );
  NAND3_X2 U4446 ( .A1(n3944), .A2(n2594), .A3(n2707), .ZN(n3945) );
  NAND2_X2 U4447 ( .A1(n3946), .A2(n3945), .ZN(n4065) );
  NAND2_X2 U4448 ( .A1(net83017), .A2(net83018), .ZN(n3957) );
  NAND2_X2 U4449 ( .A1(net86044), .A2(net83016), .ZN(n3956) );
  INV_X4 U4450 ( .A(n3978), .ZN(n3985) );
  NAND2_X2 U4451 ( .A1(net83007), .A2(n3962), .ZN(n3963) );
  NAND2_X2 U4452 ( .A1(n3964), .A2(net82029), .ZN(n3966) );
  NAND2_X2 U4453 ( .A1(net82856), .A2(net85901), .ZN(n3965) );
  NAND2_X2 U4454 ( .A1(n3972), .A2(net82988), .ZN(n3973) );
  AOI21_X2 U4455 ( .B1(u4_N1600), .B2(n3978), .A(u4_N1598), .ZN(n3980) );
  NAND2_X2 U4456 ( .A1(n3982), .A2(n3981), .ZN(n3983) );
  OAI21_X4 U4457 ( .B1(n3987), .B2(n3986), .A(n2674), .ZN(n3992) );
  NAND3_X2 U4458 ( .A1(n2740), .A2(n3989), .A3(n3988), .ZN(n3990) );
  NAND2_X2 U4459 ( .A1(n3992), .A2(n3991), .ZN(n3994) );
  NAND3_X2 U4460 ( .A1(n3996), .A2(n3997), .A3(net82950), .ZN(n4059) );
  INV_X4 U4461 ( .A(net86032), .ZN(net82938) );
  INV_X4 U4462 ( .A(n4019), .ZN(n4012) );
  NAND4_X2 U4463 ( .A1(n4008), .A2(net82925), .A3(n4007), .A4(net82927), .ZN(
        n4009) );
  INV_X4 U4464 ( .A(n4115), .ZN(n4011) );
  NOR2_X4 U4465 ( .A1(n4015), .A2(net86028), .ZN(n4016) );
  AOI21_X4 U4466 ( .B1(n4018), .B2(n4017), .A(n4016), .ZN(n4023) );
  INV_X4 U4467 ( .A(net82767), .ZN(net82911) );
  NAND2_X2 U4468 ( .A1(net82911), .A2(n2698), .ZN(n4113) );
  NAND2_X2 U4469 ( .A1(n4028), .A2(n4027), .ZN(n4030) );
  NAND3_X4 U4470 ( .A1(n4035), .A2(n2938), .A3(n4034), .ZN(n4037) );
  NAND4_X2 U4471 ( .A1(n4043), .A2(n4042), .A3(n4041), .A4(n4040), .ZN(n4044)
         );
  NAND2_X2 U4472 ( .A1(net82873), .A2(n4045), .ZN(n4048) );
  NAND3_X2 U4473 ( .A1(n1898), .A2(n1900), .A3(n2730), .ZN(n4047) );
  NAND3_X2 U4474 ( .A1(n1890), .A2(n1892), .A3(n1889), .ZN(n4046) );
  NOR3_X2 U4475 ( .A1(n4048), .A2(n4047), .A3(n4046), .ZN(n4055) );
  NAND2_X2 U4476 ( .A1(n4062), .A2(n4061), .ZN(N522) );
  OAI22_X2 U4477 ( .A1(opa_00), .A2(n2698), .B1(opb_inf), .B2(n2594), .ZN(
        n4064) );
  NAND2_X2 U4478 ( .A1(net86027), .A2(n4064), .ZN(n4066) );
  NAND3_X2 U4479 ( .A1(inf_d), .A2(n4071), .A3(n4070), .ZN(n4072) );
  MUX2_X2 U4480 ( .A(net82778), .B(n4728), .S(net82757), .Z(N467) );
  INV_X4 U4481 ( .A(n4113), .ZN(n4114) );
  NAND2_X2 U4482 ( .A1(net82753), .A2(net82764), .ZN(N470) );
  NAND2_X2 U4483 ( .A1(net82753), .A2(n2831), .ZN(N469) );
  NAND2_X2 U4484 ( .A1(net82753), .A2(net82762), .ZN(N475) );
  NAND2_X2 U4485 ( .A1(net82753), .A2(n4120), .ZN(N473) );
  INV_X4 U4486 ( .A(N194), .ZN(n4123) );
  MUX2_X2 U4487 ( .A(n2591), .B(n4123), .S(n3092), .Z(n4124) );
  INV_X4 U4488 ( .A(n4124), .ZN(u6_N48) );
  INV_X4 U4489 ( .A(N193), .ZN(n4125) );
  MUX2_X2 U4490 ( .A(n2599), .B(n4125), .S(n3092), .Z(n4126) );
  INV_X4 U4491 ( .A(n4126), .ZN(u6_N47) );
  INV_X4 U4492 ( .A(N192), .ZN(n4127) );
  MUX2_X2 U4493 ( .A(n2683), .B(n4127), .S(n3092), .Z(n4128) );
  INV_X4 U4494 ( .A(n4128), .ZN(u6_N46) );
  INV_X4 U4495 ( .A(N191), .ZN(n4129) );
  MUX2_X2 U4496 ( .A(n2592), .B(n4129), .S(n3092), .Z(n4130) );
  INV_X4 U4497 ( .A(n4130), .ZN(u6_N45) );
  INV_X4 U4498 ( .A(N190), .ZN(n4131) );
  MUX2_X2 U4499 ( .A(n2677), .B(n4131), .S(n3092), .Z(n4132) );
  INV_X4 U4500 ( .A(n4132), .ZN(u6_N44) );
  INV_X4 U4501 ( .A(N189), .ZN(n4133) );
  MUX2_X2 U4502 ( .A(n2590), .B(n4133), .S(n3093), .Z(n4134) );
  INV_X4 U4503 ( .A(n4134), .ZN(u6_N43) );
  INV_X4 U4504 ( .A(N188), .ZN(n4135) );
  MUX2_X2 U4505 ( .A(n2675), .B(n4135), .S(n3092), .Z(n4136) );
  INV_X4 U4506 ( .A(n4136), .ZN(u6_N42) );
  INV_X4 U4507 ( .A(N187), .ZN(n4137) );
  MUX2_X2 U4508 ( .A(n2696), .B(n4137), .S(n3092), .Z(n4138) );
  INV_X4 U4509 ( .A(n4138), .ZN(u6_N41) );
  INV_X4 U4510 ( .A(N186), .ZN(n4139) );
  MUX2_X2 U4511 ( .A(n2687), .B(n4139), .S(n3092), .Z(n4140) );
  INV_X4 U4512 ( .A(n4140), .ZN(u6_N40) );
  INV_X4 U4513 ( .A(N185), .ZN(n4141) );
  MUX2_X2 U4514 ( .A(n2678), .B(n4141), .S(n3092), .Z(n4142) );
  INV_X4 U4515 ( .A(n4142), .ZN(u6_N39) );
  INV_X4 U4516 ( .A(N184), .ZN(n4143) );
  MUX2_X2 U4517 ( .A(n2692), .B(n4143), .S(n3092), .Z(n4144) );
  INV_X4 U4518 ( .A(n4144), .ZN(u6_N38) );
  INV_X4 U4519 ( .A(N183), .ZN(n4145) );
  MUX2_X2 U4520 ( .A(n2697), .B(n4145), .S(n3092), .Z(n4146) );
  INV_X4 U4521 ( .A(n4146), .ZN(u6_N37) );
  INV_X4 U4522 ( .A(N182), .ZN(n4147) );
  MUX2_X2 U4523 ( .A(n2593), .B(n4147), .S(n3093), .Z(n4148) );
  INV_X4 U4524 ( .A(n4148), .ZN(u6_N36) );
  INV_X4 U4525 ( .A(N181), .ZN(n4149) );
  MUX2_X2 U4526 ( .A(n2681), .B(n4149), .S(n3093), .Z(n4150) );
  INV_X4 U4527 ( .A(n4150), .ZN(u6_N35) );
  INV_X4 U4528 ( .A(N180), .ZN(n4151) );
  MUX2_X2 U4529 ( .A(n2695), .B(n4151), .S(n3093), .Z(n4152) );
  INV_X4 U4530 ( .A(n4152), .ZN(u6_N34) );
  INV_X4 U4531 ( .A(N179), .ZN(n4153) );
  MUX2_X2 U4532 ( .A(n2689), .B(n4153), .S(n3093), .Z(n4154) );
  INV_X4 U4533 ( .A(n4154), .ZN(u6_N33) );
  INV_X4 U4534 ( .A(N178), .ZN(n4155) );
  MUX2_X2 U4535 ( .A(n2685), .B(n4155), .S(n3093), .Z(n4156) );
  INV_X4 U4536 ( .A(n4156), .ZN(u6_N32) );
  INV_X4 U4537 ( .A(N177), .ZN(n4157) );
  MUX2_X2 U4538 ( .A(n2596), .B(n4157), .S(n3093), .Z(n4158) );
  INV_X4 U4539 ( .A(n4158), .ZN(u6_N31) );
  INV_X4 U4540 ( .A(N176), .ZN(n4159) );
  MUX2_X2 U4541 ( .A(n2690), .B(n4159), .S(n3093), .Z(n4160) );
  INV_X4 U4542 ( .A(n4160), .ZN(u6_N30) );
  INV_X4 U4543 ( .A(N175), .ZN(n4161) );
  MUX2_X2 U4544 ( .A(n2598), .B(n4161), .S(n3093), .Z(n4162) );
  INV_X4 U4545 ( .A(n4162), .ZN(u6_N29) );
  INV_X4 U4546 ( .A(fracta_mul[2]), .ZN(n4524) );
  INV_X4 U4547 ( .A(N174), .ZN(n4163) );
  MUX2_X2 U4548 ( .A(n4524), .B(n4163), .S(n3093), .Z(n4164) );
  INV_X4 U4549 ( .A(n4164), .ZN(u6_N28) );
  INV_X4 U4550 ( .A(N173), .ZN(n4165) );
  MUX2_X2 U4551 ( .A(n4523), .B(n4165), .S(n3093), .Z(n4166) );
  INV_X4 U4552 ( .A(n4166), .ZN(u6_N27) );
  INV_X4 U4553 ( .A(fracta_mul[0]), .ZN(n4530) );
  INV_X4 U4554 ( .A(N172), .ZN(n4167) );
  MUX2_X2 U4555 ( .A(n4530), .B(n4167), .S(n3092), .Z(n4168) );
  INV_X4 U4556 ( .A(n4168), .ZN(u6_N26) );
  INV_X4 U4557 ( .A(u2_N22), .ZN(n4170) );
  INV_X4 U4558 ( .A(u2_N13), .ZN(n4169) );
  MUX2_X2 U4559 ( .A(n4170), .B(n4169), .S(n4318), .Z(n4231) );
  INV_X4 U4560 ( .A(n4231), .ZN(u2_exp_tmp4_7_) );
  INV_X4 U4561 ( .A(u2_N16), .ZN(n4172) );
  INV_X4 U4562 ( .A(u2_N7), .ZN(n4171) );
  MUX2_X2 U4563 ( .A(n4172), .B(n4171), .S(n4318), .Z(u2_exp_tmp4_1_) );
  INV_X4 U4564 ( .A(u2_exp_tmp4_1_), .ZN(n4264) );
  INV_X4 U4565 ( .A(u2_N15), .ZN(n4174) );
  INV_X4 U4566 ( .A(u2_N6), .ZN(n4173) );
  MUX2_X2 U4567 ( .A(n4174), .B(n4173), .S(n4318), .Z(u2_exp_tmp4_0_) );
  INV_X4 U4568 ( .A(u2_exp_tmp4_0_), .ZN(n4281) );
  INV_X4 U4569 ( .A(u2_N17), .ZN(n4176) );
  INV_X4 U4570 ( .A(u2_N8), .ZN(n4175) );
  MUX2_X2 U4571 ( .A(n4176), .B(n4175), .S(n4318), .Z(u2_exp_tmp4_2_) );
  INV_X4 U4572 ( .A(u2_exp_tmp4_2_), .ZN(n4265) );
  INV_X4 U4573 ( .A(n4226), .ZN(n4217) );
  INV_X4 U4574 ( .A(u2_N19), .ZN(n4178) );
  INV_X4 U4575 ( .A(u2_N10), .ZN(n4177) );
  MUX2_X2 U4576 ( .A(n4178), .B(n4177), .S(n4318), .Z(u2_exp_tmp4_4_) );
  INV_X4 U4577 ( .A(u2_exp_tmp4_4_), .ZN(n4214) );
  INV_X4 U4578 ( .A(u2_N18), .ZN(n4180) );
  INV_X4 U4579 ( .A(u2_N9), .ZN(n4179) );
  MUX2_X2 U4580 ( .A(n4180), .B(n4179), .S(n4318), .Z(u2_exp_tmp4_3_) );
  INV_X4 U4581 ( .A(u2_exp_tmp4_3_), .ZN(n4218) );
  INV_X4 U4582 ( .A(n4212), .ZN(n4204) );
  INV_X4 U4583 ( .A(u2_N20), .ZN(n4182) );
  INV_X4 U4584 ( .A(u2_N11), .ZN(n4181) );
  MUX2_X2 U4585 ( .A(n4182), .B(n4181), .S(n4318), .Z(u2_exp_tmp4_5_) );
  INV_X4 U4586 ( .A(u2_exp_tmp4_5_), .ZN(n4205) );
  NAND2_X2 U4587 ( .A1(n4204), .A2(n4205), .ZN(n4199) );
  INV_X4 U4588 ( .A(n4199), .ZN(n4183) );
  INV_X4 U4589 ( .A(u2_N21), .ZN(n4290) );
  INV_X4 U4590 ( .A(u2_N12), .ZN(n4296) );
  MUX2_X2 U4591 ( .A(n4290), .B(n4296), .S(n4318), .Z(u2_exp_tmp4_6_) );
  INV_X4 U4592 ( .A(u2_exp_tmp4_6_), .ZN(n4201) );
  NAND2_X2 U4593 ( .A1(n4183), .A2(n4201), .ZN(n4232) );
  INV_X4 U4594 ( .A(n4232), .ZN(n4184) );
  NAND2_X2 U4595 ( .A1(n4184), .A2(u2_exp_tmp4_7_), .ZN(n4185) );
  NAND2_X2 U4596 ( .A1(n4231), .A2(n4232), .ZN(n4314) );
  NAND2_X2 U4597 ( .A1(n4185), .A2(n4314), .ZN(n4190) );
  NAND2_X2 U4598 ( .A1(u2_exp_tmp4_1_), .A2(u2_exp_tmp4_0_), .ZN(n4186) );
  INV_X4 U4599 ( .A(n4221), .ZN(n4187) );
  NOR2_X4 U4600 ( .A1(n4218), .A2(n4187), .ZN(n4219) );
  INV_X4 U4601 ( .A(n4208), .ZN(n4188) );
  NOR2_X4 U4602 ( .A1(n4205), .A2(n4188), .ZN(n4206) );
  NOR2_X4 U4603 ( .A1(n4201), .A2(n4207), .ZN(n4193) );
  XNOR2_X2 U4604 ( .A(u2_exp_tmp4_7_), .B(n4193), .ZN(n4189) );
  MUX2_X2 U4605 ( .A(n4190), .B(n4189), .S(n4318), .Z(n5253) );
  NAND4_X2 U4606 ( .A1(n4288), .A2(n3065), .A3(n2566), .A4(n5253), .ZN(n4198)
         );
  INV_X4 U4607 ( .A(u2_N23), .ZN(n4192) );
  INV_X4 U4608 ( .A(u2_N14), .ZN(n4191) );
  MUX2_X2 U4609 ( .A(n4192), .B(n4191), .S(n4318), .Z(n4317) );
  XNOR2_X2 U4610 ( .A(n4317), .B(n4314), .ZN(n4197) );
  INV_X4 U4611 ( .A(n4317), .ZN(n4194) );
  XNOR2_X2 U4612 ( .A(n4195), .B(n4194), .ZN(n4196) );
  MUX2_X2 U4613 ( .A(n4197), .B(n4196), .S(n4318), .Z(n4236) );
  NAND2_X2 U4614 ( .A1(n4198), .A2(n4236), .ZN(u2_exp_ovf_d_1_) );
  NAND2_X2 U4615 ( .A1(u2_exp_tmp4_6_), .A2(n4199), .ZN(n4200) );
  NAND2_X2 U4616 ( .A1(n4200), .A2(n4232), .ZN(n4244) );
  XNOR2_X2 U4617 ( .A(n4201), .B(n4206), .ZN(n4202) );
  MUX2_X2 U4618 ( .A(n4244), .B(n4202), .S(n4318), .Z(n4203) );
  INV_X4 U4619 ( .A(n4203), .ZN(n5254) );
  XNOR2_X2 U4620 ( .A(n4205), .B(n4204), .ZN(n4250) );
  INV_X4 U4621 ( .A(n4250), .ZN(n4210) );
  INV_X4 U4622 ( .A(n4206), .ZN(n4207) );
  MUX2_X2 U4623 ( .A(n4210), .B(n4209), .S(n4318), .Z(n5255) );
  NAND2_X2 U4624 ( .A1(n4217), .A2(n4218), .ZN(n4211) );
  NAND2_X2 U4625 ( .A1(u2_exp_tmp4_4_), .A2(n4211), .ZN(n4213) );
  NAND2_X2 U4626 ( .A1(n4213), .A2(n4212), .ZN(n4255) );
  XNOR2_X2 U4627 ( .A(n4214), .B(n4219), .ZN(n4215) );
  MUX2_X2 U4628 ( .A(n4255), .B(n4215), .S(n4318), .Z(n4216) );
  INV_X4 U4629 ( .A(n4216), .ZN(n5256) );
  XNOR2_X2 U4630 ( .A(n4218), .B(n4217), .ZN(n4260) );
  INV_X4 U4631 ( .A(n4260), .ZN(n4223) );
  INV_X4 U4632 ( .A(n4219), .ZN(n4220) );
  MUX2_X2 U4633 ( .A(n4223), .B(n4222), .S(n4318), .Z(n5257) );
  NAND2_X2 U4634 ( .A1(n4318), .A2(n4265), .ZN(n4224) );
  MUX2_X2 U4635 ( .A(n4224), .B(n4265), .S(n4281), .Z(n4225) );
  MUX2_X2 U4636 ( .A(n4225), .B(n2744), .S(n4264), .Z(n4228) );
  OAI21_X4 U4637 ( .B1(n4265), .B2(n4281), .A(n4226), .ZN(n4266) );
  NAND2_X2 U4638 ( .A1(n4266), .A2(n4288), .ZN(n4227) );
  NAND2_X2 U4639 ( .A1(n4228), .A2(n4227), .ZN(n4229) );
  INV_X4 U4640 ( .A(n4229), .ZN(n5258) );
  XNOR2_X2 U4641 ( .A(n4281), .B(n4264), .ZN(n4272) );
  INV_X4 U4642 ( .A(n4272), .ZN(n4230) );
  INV_X4 U4643 ( .A(n5317), .ZN(n4315) );
  NAND2_X2 U4644 ( .A1(u2_exp_ovf_d_1_), .A2(n4315), .ZN(n4243) );
  NAND3_X4 U4645 ( .A1(n5317), .A2(n4288), .A3(u2_exp_ovf_d_1_), .ZN(n4282) );
  INV_X4 U4646 ( .A(n4282), .ZN(n4234) );
  XNOR2_X2 U4647 ( .A(u2_exp_tmp4_7_), .B(n4232), .ZN(n4233) );
  NAND2_X2 U4648 ( .A1(n4234), .A2(n4233), .ZN(n4241) );
  INV_X4 U4649 ( .A(u2_exp_ovf_d_1_), .ZN(n4238) );
  NAND2_X2 U4650 ( .A1(n5317), .A2(n4238), .ZN(n4235) );
  INV_X4 U4651 ( .A(n4235), .ZN(n4278) );
  INV_X4 U4652 ( .A(n4236), .ZN(n4286) );
  NAND2_X2 U4653 ( .A1(n4237), .A2(n4286), .ZN(n4277) );
  NAND2_X2 U4654 ( .A1(n4315), .A2(n4238), .ZN(n4239) );
  INV_X4 U4655 ( .A(n4239), .ZN(n4279) );
  AOI22_X2 U4656 ( .A1(u2_N48), .A2(n4242), .B1(u2_exp_tmp3_6_), .B2(n4278), 
        .ZN(n4248) );
  INV_X4 U4657 ( .A(n4243), .ZN(n4280) );
  NAND2_X2 U4658 ( .A1(n4280), .A2(u2_exp_tmp4_6_), .ZN(n4247) );
  INV_X4 U4659 ( .A(n4282), .ZN(n4273) );
  NAND2_X2 U4660 ( .A1(n4273), .A2(n4244), .ZN(n4246) );
  NAND2_X2 U4661 ( .A1(n5254), .A2(n4279), .ZN(n4245) );
  NAND4_X2 U4662 ( .A1(n4248), .A2(n4247), .A3(n4246), .A4(n4245), .ZN(u2_N64)
         );
  AOI22_X2 U4663 ( .A1(u2_N47), .A2(n4249), .B1(n5255), .B2(n4279), .ZN(n4253)
         );
  NAND2_X2 U4664 ( .A1(u2_exp_tmp3_5_), .A2(n4278), .ZN(n4252) );
  AOI22_X2 U4665 ( .A1(n4280), .A2(u2_exp_tmp4_5_), .B1(n4273), .B2(n4250), 
        .ZN(n4251) );
  AOI22_X2 U4666 ( .A1(u2_N46), .A2(n4254), .B1(u2_exp_tmp3_4_), .B2(n4278), 
        .ZN(n4259) );
  NAND2_X2 U4667 ( .A1(n4280), .A2(u2_exp_tmp4_4_), .ZN(n4258) );
  NAND2_X2 U4668 ( .A1(n4273), .A2(n4255), .ZN(n4257) );
  NAND2_X2 U4669 ( .A1(n4279), .A2(n5256), .ZN(n4256) );
  NAND4_X2 U4670 ( .A1(n4259), .A2(n4258), .A3(n4257), .A4(n4256), .ZN(u2_N62)
         );
  AOI22_X2 U4671 ( .A1(u2_N45), .A2(n4254), .B1(n5257), .B2(n4279), .ZN(n4263)
         );
  NAND2_X2 U4672 ( .A1(u2_exp_tmp3_3_), .A2(n4278), .ZN(n4262) );
  AOI22_X2 U4673 ( .A1(n4280), .A2(u2_exp_tmp4_3_), .B1(n4273), .B2(n4260), 
        .ZN(n4261) );
  AOI22_X2 U4674 ( .A1(u2_N44), .A2(n4249), .B1(u2_exp_tmp3_2_), .B2(n4278), 
        .ZN(n4271) );
  NAND2_X2 U4675 ( .A1(n4280), .A2(u2_exp_tmp4_2_), .ZN(n4270) );
  NAND2_X2 U4676 ( .A1(n5258), .A2(n4279), .ZN(n4268) );
  NAND4_X2 U4677 ( .A1(n4271), .A2(n4270), .A3(n4269), .A4(n4268), .ZN(u2_N60)
         );
  AOI22_X2 U4678 ( .A1(u2_N43), .A2(n4242), .B1(n4279), .B2(n2716), .ZN(n4276)
         );
  NAND2_X2 U4679 ( .A1(u2_exp_tmp3_1_), .A2(n4278), .ZN(n4275) );
  AOI22_X2 U4680 ( .A1(n4280), .A2(u2_exp_tmp4_1_), .B1(n4273), .B2(n4272), 
        .ZN(n4274) );
  AOI22_X2 U4681 ( .A1(u2_N42), .A2(n4254), .B1(u2_exp_tmp3_0_), .B2(n4278), 
        .ZN(n4285) );
  NOR2_X4 U4682 ( .A1(n4280), .A2(n4279), .ZN(n4283) );
  MUX2_X2 U4683 ( .A(n4283), .B(n4282), .S(n4281), .Z(n4284) );
  NAND2_X2 U4684 ( .A1(n4285), .A2(n4284), .ZN(u2_N58) );
  NAND2_X2 U4685 ( .A1(n4286), .A2(n4288), .ZN(n4287) );
  MUX2_X2 U4686 ( .A(n4288), .B(n4287), .S(opb_r[30]), .Z(n4289) );
  AND2_X2 U4687 ( .A1(u2_N20), .A2(u2_N19), .ZN(n4295) );
  NAND2_X2 U4688 ( .A1(u2_N18), .A2(u2_N17), .ZN(n4292) );
  NAND2_X2 U4689 ( .A1(u2_N16), .A2(u2_N15), .ZN(n4291) );
  NAND3_X2 U4690 ( .A1(n4295), .A2(n4294), .A3(n4293), .ZN(n4303) );
  AND2_X2 U4691 ( .A1(u2_N11), .A2(u2_N10), .ZN(n4301) );
  NAND2_X2 U4692 ( .A1(u2_N9), .A2(u2_N8), .ZN(n4298) );
  NAND2_X2 U4693 ( .A1(u2_N7), .A2(u2_N6), .ZN(n4297) );
  NAND3_X2 U4694 ( .A1(n4301), .A2(n4300), .A3(n4299), .ZN(n4302) );
  MUX2_X2 U4695 ( .A(n4303), .B(n4302), .S(n4318), .Z(n4309) );
  NAND2_X2 U4696 ( .A1(n1735), .A2(n2591), .ZN(n4741) );
  NAND2_X2 U4697 ( .A1(n1751), .A2(n1752), .ZN(n4305) );
  INV_X4 U4698 ( .A(n1749), .ZN(n4304) );
  NAND2_X2 U4699 ( .A1(n2604), .A2(n4491), .ZN(n4742) );
  NAND2_X2 U4700 ( .A1(n4742), .A2(n4765), .ZN(n4311) );
  NAND2_X2 U4701 ( .A1(n4741), .A2(n3093), .ZN(n4310) );
  OAI211_X2 U4702 ( .C1(n4313), .C2(n4312), .A(n4311), .B(n4310), .ZN(
        u2_underflow_d[1]) );
  INV_X4 U4703 ( .A(n4314), .ZN(n4316) );
  NOR2_X4 U4704 ( .A1(n4317), .A2(n4316), .ZN(n4320) );
  MUX2_X2 U4705 ( .A(n4320), .B(n4319), .S(n4318), .Z(u2_N90) );
  NAND4_X2 U4706 ( .A1(n4324), .A2(n4323), .A3(n4322), .A4(n4321), .ZN(N224)
         );
  NAND2_X2 U4707 ( .A1(fpu_op_r2[0]), .A2(fpu_op_r2[2]), .ZN(n2431) );
  INV_X4 U4708 ( .A(n2431), .ZN(n4325) );
  NAND2_X2 U4709 ( .A1(n4325), .A2(n2567), .ZN(n5321) );
  MUX2_X2 U4710 ( .A(n2608), .B(n2734), .S(fpu_op_r2[1]), .Z(n4362) );
  INV_X4 U4711 ( .A(n4362), .ZN(n5322) );
  INV_X4 U4712 ( .A(n5321), .ZN(n4326) );
  NAND2_X2 U4713 ( .A1(n5322), .A2(n4326), .ZN(n4328) );
  INV_X4 U4714 ( .A(N227), .ZN(n4327) );
  NAND2_X2 U4715 ( .A1(n4362), .A2(n4326), .ZN(n4329) );
  OAI22_X2 U4716 ( .A1(n4328), .A2(n4327), .B1(n4329), .B2(n2749), .ZN(n5320)
         );
  NAND2_X2 U4717 ( .A1(N228), .A2(n4389), .ZN(n4331) );
  NAND2_X2 U4718 ( .A1(opa_r1[1]), .A2(n4384), .ZN(n4330) );
  NAND2_X2 U4719 ( .A1(n4331), .A2(n4330), .ZN(n5252) );
  NAND2_X2 U4720 ( .A1(N229), .A2(n4389), .ZN(n4333) );
  NAND2_X2 U4721 ( .A1(opa_r1[2]), .A2(n4384), .ZN(n4332) );
  NAND2_X2 U4722 ( .A1(n4333), .A2(n4332), .ZN(n5251) );
  NAND2_X2 U4723 ( .A1(N230), .A2(n4389), .ZN(n4335) );
  NAND2_X2 U4724 ( .A1(opa_r1[3]), .A2(n4384), .ZN(n4334) );
  NAND2_X2 U4725 ( .A1(n4335), .A2(n4334), .ZN(n5250) );
  NAND2_X2 U4726 ( .A1(N231), .A2(n4389), .ZN(n4337) );
  NAND2_X2 U4727 ( .A1(opa_r1[4]), .A2(n4384), .ZN(n4336) );
  NAND2_X2 U4728 ( .A1(n4337), .A2(n4336), .ZN(n5249) );
  NAND2_X2 U4729 ( .A1(N232), .A2(n4389), .ZN(n4339) );
  NAND2_X2 U4730 ( .A1(opa_r1[5]), .A2(n4384), .ZN(n4338) );
  NAND2_X2 U4731 ( .A1(n4339), .A2(n4338), .ZN(n5248) );
  NAND2_X2 U4732 ( .A1(N233), .A2(n4389), .ZN(n4341) );
  NAND2_X2 U4733 ( .A1(n4384), .A2(opa_r1[6]), .ZN(n4340) );
  NAND2_X2 U4734 ( .A1(n4341), .A2(n4340), .ZN(n5247) );
  NAND2_X2 U4735 ( .A1(N234), .A2(n4389), .ZN(n4343) );
  NAND2_X2 U4736 ( .A1(n4384), .A2(opa_r1[7]), .ZN(n4342) );
  NAND2_X2 U4737 ( .A1(n4343), .A2(n4342), .ZN(n5246) );
  NAND2_X2 U4738 ( .A1(N235), .A2(n4389), .ZN(n4345) );
  NAND2_X2 U4739 ( .A1(n4384), .A2(opa_r1[8]), .ZN(n4344) );
  NAND2_X2 U4740 ( .A1(n4345), .A2(n4344), .ZN(n5245) );
  NAND2_X2 U4741 ( .A1(N236), .A2(n4389), .ZN(n4347) );
  NAND2_X2 U4742 ( .A1(n4384), .A2(opa_r1[9]), .ZN(n4346) );
  NAND2_X2 U4743 ( .A1(n4347), .A2(n4346), .ZN(n5244) );
  NAND2_X2 U4744 ( .A1(N237), .A2(n4389), .ZN(n4349) );
  NAND2_X2 U4745 ( .A1(n4384), .A2(opa_r1[10]), .ZN(n4348) );
  NAND2_X2 U4746 ( .A1(n4349), .A2(n4348), .ZN(n5243) );
  NAND2_X2 U4747 ( .A1(N238), .A2(n4389), .ZN(n4351) );
  NAND2_X2 U4748 ( .A1(n4384), .A2(opa_r1[11]), .ZN(n4350) );
  NAND2_X2 U4749 ( .A1(n4351), .A2(n4350), .ZN(n5242) );
  NAND2_X2 U4750 ( .A1(N239), .A2(n4389), .ZN(n4353) );
  NAND2_X2 U4751 ( .A1(n4384), .A2(opa_r1[12]), .ZN(n4352) );
  NAND2_X2 U4752 ( .A1(n4353), .A2(n4352), .ZN(n5241) );
  NAND2_X2 U4753 ( .A1(N240), .A2(n4389), .ZN(n4355) );
  NAND2_X2 U4754 ( .A1(n4384), .A2(opa_r1[13]), .ZN(n4354) );
  NAND2_X2 U4755 ( .A1(n4355), .A2(n4354), .ZN(n5240) );
  NAND2_X2 U4756 ( .A1(N241), .A2(n4389), .ZN(n4357) );
  NAND2_X2 U4757 ( .A1(n4384), .A2(opa_r1[14]), .ZN(n4356) );
  NAND2_X2 U4758 ( .A1(n4357), .A2(n4356), .ZN(n5239) );
  NAND2_X2 U4759 ( .A1(N242), .A2(n4389), .ZN(n4359) );
  NAND2_X2 U4760 ( .A1(n4384), .A2(opa_r1[15]), .ZN(n4358) );
  NAND2_X2 U4761 ( .A1(n4359), .A2(n4358), .ZN(n5238) );
  NAND2_X2 U4762 ( .A1(N243), .A2(n4389), .ZN(n4361) );
  NAND2_X2 U4763 ( .A1(n4384), .A2(opa_r1[16]), .ZN(n4360) );
  NAND2_X2 U4764 ( .A1(n4361), .A2(n4360), .ZN(n5237) );
  NAND2_X2 U4765 ( .A1(N244), .A2(n4389), .ZN(n4365) );
  NAND2_X2 U4766 ( .A1(N227), .A2(n2565), .ZN(n4364) );
  NAND2_X2 U4767 ( .A1(n4384), .A2(opa_r1[17]), .ZN(n4363) );
  NAND3_X2 U4768 ( .A1(n4365), .A2(n4364), .A3(n4363), .ZN(N391) );
  NAND2_X2 U4769 ( .A1(N245), .A2(n4389), .ZN(n4368) );
  NAND2_X2 U4770 ( .A1(opa_r1[1]), .A2(n2565), .ZN(n4367) );
  NAND2_X2 U4771 ( .A1(n4384), .A2(opa_r1[18]), .ZN(n4366) );
  NAND3_X2 U4772 ( .A1(n4368), .A2(n4367), .A3(n4366), .ZN(N392) );
  NAND2_X2 U4773 ( .A1(n4384), .A2(opa_r1[19]), .ZN(n4371) );
  NAND2_X2 U4774 ( .A1(N246), .A2(n4389), .ZN(n4370) );
  AOI22_X2 U4775 ( .A1(N227), .A2(n2588), .B1(opa_r1[2]), .B2(n2565), .ZN(
        n4369) );
  NAND3_X2 U4776 ( .A1(n4371), .A2(n4370), .A3(n4369), .ZN(N393) );
  NAND2_X2 U4777 ( .A1(N298), .A2(n2588), .ZN(n4375) );
  NAND2_X2 U4778 ( .A1(opa_r1[3]), .A2(n2565), .ZN(n4374) );
  NAND2_X2 U4779 ( .A1(N247), .A2(n4389), .ZN(n4373) );
  NAND2_X2 U4780 ( .A1(n4384), .A2(opa_r1[20]), .ZN(n4372) );
  NAND4_X2 U4781 ( .A1(n4375), .A2(n4374), .A3(n4373), .A4(n4372), .ZN(N394)
         );
  NAND2_X2 U4782 ( .A1(N299), .A2(n2588), .ZN(n4379) );
  NAND2_X2 U4783 ( .A1(opa_r1[4]), .A2(n2565), .ZN(n4378) );
  NAND2_X2 U4784 ( .A1(N248), .A2(n4389), .ZN(n4377) );
  NAND2_X2 U4785 ( .A1(n4384), .A2(opa_r1[21]), .ZN(n4376) );
  NAND4_X2 U4786 ( .A1(n4379), .A2(n4378), .A3(n4377), .A4(n4376), .ZN(N395)
         );
  NAND2_X2 U4787 ( .A1(N300), .A2(n2588), .ZN(n4383) );
  NAND2_X2 U4788 ( .A1(opa_r1[5]), .A2(n2565), .ZN(n4382) );
  NAND2_X2 U4789 ( .A1(N249), .A2(n4389), .ZN(n4381) );
  NAND2_X2 U4790 ( .A1(n4384), .A2(opa_r1[22]), .ZN(n4380) );
  NAND4_X2 U4791 ( .A1(n4383), .A2(n4382), .A3(n4381), .A4(n4380), .ZN(N396)
         );
  NAND2_X2 U4792 ( .A1(N301), .A2(n2588), .ZN(n4388) );
  NAND2_X2 U4793 ( .A1(opa_r1[6]), .A2(n2565), .ZN(n4387) );
  NAND2_X2 U4794 ( .A1(N250), .A2(n4389), .ZN(n4386) );
  NAND2_X2 U4795 ( .A1(n4384), .A2(N224), .ZN(n4385) );
  NAND4_X2 U4796 ( .A1(n4388), .A2(n4387), .A3(n4386), .A4(n4385), .ZN(N397)
         );
  NAND2_X2 U4797 ( .A1(N302), .A2(n2588), .ZN(n4391) );
  NAND2_X2 U4798 ( .A1(opa_r1[7]), .A2(n2565), .ZN(n4390) );
  NAND3_X2 U4799 ( .A1(n4391), .A2(n4436), .A3(n4390), .ZN(N398) );
  NAND2_X2 U4800 ( .A1(N303), .A2(n2588), .ZN(n4393) );
  NAND2_X2 U4801 ( .A1(opa_r1[8]), .A2(n2565), .ZN(n4392) );
  NAND3_X2 U4802 ( .A1(n4393), .A2(n3074), .A3(n4392), .ZN(N399) );
  NAND2_X2 U4803 ( .A1(N304), .A2(n2588), .ZN(n4395) );
  NAND2_X2 U4804 ( .A1(opa_r1[9]), .A2(n2565), .ZN(n4394) );
  NAND3_X2 U4805 ( .A1(n4395), .A2(n4436), .A3(n4394), .ZN(N400) );
  NAND2_X2 U4806 ( .A1(N305), .A2(n2588), .ZN(n4397) );
  NAND2_X2 U4807 ( .A1(opa_r1[10]), .A2(n2565), .ZN(n4396) );
  NAND3_X2 U4808 ( .A1(n4397), .A2(n3074), .A3(n4396), .ZN(N401) );
  NAND2_X2 U4809 ( .A1(N306), .A2(n2588), .ZN(n4399) );
  NAND2_X2 U4810 ( .A1(opa_r1[11]), .A2(n2565), .ZN(n4398) );
  NAND3_X2 U4811 ( .A1(n4399), .A2(n4436), .A3(n4398), .ZN(N402) );
  NAND2_X2 U4812 ( .A1(N307), .A2(n2588), .ZN(n4401) );
  NAND2_X2 U4813 ( .A1(opa_r1[12]), .A2(n2565), .ZN(n4400) );
  NAND3_X2 U4814 ( .A1(n4401), .A2(n3074), .A3(n4400), .ZN(N403) );
  NAND2_X2 U4815 ( .A1(N308), .A2(n2588), .ZN(n4403) );
  NAND2_X2 U4816 ( .A1(opa_r1[13]), .A2(n2565), .ZN(n4402) );
  NAND3_X2 U4817 ( .A1(n4403), .A2(n4436), .A3(n4402), .ZN(N404) );
  NAND2_X2 U4818 ( .A1(N309), .A2(n2588), .ZN(n4405) );
  NAND2_X2 U4819 ( .A1(opa_r1[14]), .A2(n2565), .ZN(n4404) );
  NAND3_X2 U4820 ( .A1(n4405), .A2(n3074), .A3(n4404), .ZN(N405) );
  NAND2_X2 U4821 ( .A1(N310), .A2(n2588), .ZN(n4407) );
  NAND2_X2 U4822 ( .A1(opa_r1[15]), .A2(n2565), .ZN(n4406) );
  NAND3_X2 U4823 ( .A1(n4407), .A2(n4436), .A3(n4406), .ZN(N406) );
  NAND2_X2 U4824 ( .A1(N311), .A2(n2588), .ZN(n4409) );
  NAND2_X2 U4825 ( .A1(opa_r1[16]), .A2(n2565), .ZN(n4408) );
  NAND3_X2 U4826 ( .A1(n4409), .A2(n3074), .A3(n4408), .ZN(N407) );
  NAND2_X2 U4827 ( .A1(N312), .A2(n2588), .ZN(n4411) );
  NAND2_X2 U4828 ( .A1(opa_r1[17]), .A2(n2565), .ZN(n4410) );
  NAND3_X2 U4829 ( .A1(n4411), .A2(n4436), .A3(n4410), .ZN(N408) );
  NAND2_X2 U4830 ( .A1(N313), .A2(n2588), .ZN(n4413) );
  NAND2_X2 U4831 ( .A1(opa_r1[18]), .A2(n2565), .ZN(n4412) );
  NAND3_X2 U4832 ( .A1(n4413), .A2(n3074), .A3(n4412), .ZN(N409) );
  NAND2_X2 U4833 ( .A1(N314), .A2(n2588), .ZN(n4415) );
  NAND2_X2 U4834 ( .A1(opa_r1[19]), .A2(n2565), .ZN(n4414) );
  NAND3_X2 U4835 ( .A1(n4415), .A2(n4436), .A3(n4414), .ZN(N410) );
  NAND2_X2 U4836 ( .A1(N315), .A2(n2588), .ZN(n4417) );
  NAND2_X2 U4837 ( .A1(opa_r1[20]), .A2(n2565), .ZN(n4416) );
  NAND3_X2 U4838 ( .A1(n4417), .A2(n3074), .A3(n4416), .ZN(N411) );
  NAND2_X2 U4839 ( .A1(N316), .A2(n2588), .ZN(n4419) );
  NAND2_X2 U4840 ( .A1(opa_r1[21]), .A2(n2565), .ZN(n4418) );
  NAND3_X2 U4841 ( .A1(n4419), .A2(n4436), .A3(n4418), .ZN(N412) );
  NAND2_X2 U4842 ( .A1(N317), .A2(n2588), .ZN(n4421) );
  NAND2_X2 U4843 ( .A1(opa_r1[22]), .A2(n2565), .ZN(n4420) );
  NAND3_X2 U4844 ( .A1(n4421), .A2(n3074), .A3(n4420), .ZN(N413) );
  NAND2_X2 U4845 ( .A1(N318), .A2(n2588), .ZN(n4423) );
  NAND2_X2 U4846 ( .A1(n2565), .A2(opa_r1[23]), .ZN(n4422) );
  NAND3_X2 U4847 ( .A1(n4423), .A2(n4436), .A3(n4422), .ZN(N414) );
  NAND2_X2 U4848 ( .A1(N319), .A2(n2588), .ZN(n4425) );
  NAND2_X2 U4849 ( .A1(n2565), .A2(opa_r1[24]), .ZN(n4424) );
  NAND3_X2 U4850 ( .A1(n4425), .A2(n3074), .A3(n4424), .ZN(N415) );
  NAND2_X2 U4851 ( .A1(N320), .A2(n2588), .ZN(n4427) );
  NAND2_X2 U4852 ( .A1(n2565), .A2(opa_r1[25]), .ZN(n4426) );
  NAND3_X2 U4853 ( .A1(n4427), .A2(n4436), .A3(n4426), .ZN(N416) );
  NAND2_X2 U4854 ( .A1(N321), .A2(n2588), .ZN(n4429) );
  NAND2_X2 U4855 ( .A1(n2565), .A2(opa_r1[26]), .ZN(n4428) );
  NAND3_X2 U4856 ( .A1(n4429), .A2(n3074), .A3(n4428), .ZN(N417) );
  NAND2_X2 U4857 ( .A1(N322), .A2(n2588), .ZN(n4431) );
  NAND2_X2 U4858 ( .A1(n2565), .A2(opa_r1[27]), .ZN(n4430) );
  NAND3_X2 U4859 ( .A1(n4431), .A2(n4436), .A3(n4430), .ZN(N418) );
  NAND2_X2 U4860 ( .A1(N323), .A2(n2588), .ZN(n4433) );
  NAND2_X2 U4861 ( .A1(n2565), .A2(opa_r1[28]), .ZN(n4432) );
  NAND3_X2 U4862 ( .A1(n4433), .A2(n3074), .A3(n4432), .ZN(N419) );
  NAND2_X2 U4863 ( .A1(N324), .A2(n2588), .ZN(n4435) );
  NAND2_X2 U4864 ( .A1(n2565), .A2(opa_r1[29]), .ZN(n4434) );
  NAND3_X2 U4865 ( .A1(n4435), .A2(n4436), .A3(n4434), .ZN(N420) );
  NAND2_X2 U4866 ( .A1(n2565), .A2(opa_r1[30]), .ZN(n4438) );
  NAND2_X2 U4867 ( .A1(N325), .A2(n2588), .ZN(n4437) );
  NAND3_X2 U4868 ( .A1(n4438), .A2(n4437), .A3(n3074), .ZN(N421) );
  XNOR2_X2 U4869 ( .A(opb_r[31]), .B(opa_r[31]), .ZN(n4439) );
  INV_X4 U4870 ( .A(n4439), .ZN(u2_sign_d) );
  INV_X4 U4871 ( .A(n4465), .ZN(n5309) );
  NAND2_X2 U4872 ( .A1(opb_r[24]), .A2(n2763), .ZN(n4459) );
  OAI22_X2 U4873 ( .A1(opb_r[23]), .A2(n2655), .B1(opb_r[24]), .B2(n2763), 
        .ZN(n4442) );
  NAND2_X2 U4874 ( .A1(opb_r[25]), .A2(n2765), .ZN(n4456) );
  NAND3_X2 U4875 ( .A1(n4459), .A2(n4442), .A3(n4456), .ZN(n4444) );
  NAND2_X2 U4876 ( .A1(opb_r[26]), .A2(n2764), .ZN(n4454) );
  NAND2_X2 U4877 ( .A1(n4460), .A2(n4454), .ZN(n4443) );
  AOI21_X4 U4878 ( .B1(n4445), .B2(n4444), .A(n4443), .ZN(n4447) );
  NAND2_X2 U4879 ( .A1(opb_r[28]), .A2(n2582), .ZN(n4457) );
  OAI21_X4 U4880 ( .B1(n4447), .B2(n4446), .A(n4457), .ZN(n4451) );
  INV_X4 U4881 ( .A(opb_r[29]), .ZN(n4734) );
  NAND2_X2 U4882 ( .A1(opa_r[29]), .A2(n4734), .ZN(n4450) );
  INV_X4 U4883 ( .A(n4455), .ZN(n4449) );
  NAND2_X2 U4884 ( .A1(opb_r[29]), .A2(n2653), .ZN(n4458) );
  INV_X4 U4885 ( .A(n4458), .ZN(n4448) );
  AOI211_X4 U4886 ( .C1(n4451), .C2(n4450), .A(n4449), .B(n4448), .ZN(n4452)
         );
  INV_X4 U4887 ( .A(opb_r[23]), .ZN(n4475) );
  NAND2_X2 U4888 ( .A1(n4460), .A2(n4459), .ZN(n4461) );
  NOR4_X2 U4889 ( .A1(n4464), .A2(n4463), .A3(n4462), .A4(n4461), .ZN(n4476)
         );
  MUX2_X2 U4890 ( .A(n2653), .B(n4734), .S(n3077), .Z(n4466) );
  INV_X4 U4891 ( .A(n4466), .ZN(n5310) );
  INV_X4 U4892 ( .A(opb_r[28]), .ZN(n4467) );
  MUX2_X2 U4893 ( .A(n2582), .B(n4467), .S(n3078), .Z(n4468) );
  INV_X4 U4894 ( .A(n4468), .ZN(n5311) );
  INV_X4 U4895 ( .A(opb_r[27]), .ZN(n4469) );
  MUX2_X2 U4896 ( .A(n2657), .B(n4469), .S(n3077), .Z(n4470) );
  INV_X4 U4897 ( .A(n4470), .ZN(n5312) );
  INV_X4 U4898 ( .A(opb_r[26]), .ZN(n4736) );
  MUX2_X2 U4899 ( .A(n2764), .B(n4736), .S(n3078), .Z(n4471) );
  INV_X4 U4900 ( .A(n4471), .ZN(n5313) );
  INV_X4 U4901 ( .A(opb_r[25]), .ZN(n4737) );
  MUX2_X2 U4902 ( .A(n2765), .B(n4737), .S(n3076), .Z(n4472) );
  INV_X4 U4903 ( .A(n4472), .ZN(n5314) );
  MUX2_X2 U4904 ( .A(n2763), .B(n4473), .S(n3077), .Z(n4474) );
  INV_X4 U4905 ( .A(n4474), .ZN(n5315) );
  MUX2_X2 U4906 ( .A(n2655), .B(n4475), .S(n3078), .Z(n4477) );
  INV_X4 U4907 ( .A(n4477), .ZN(n5316) );
  MUX2_X2 U4908 ( .A(u3_N58), .B(u3_N30), .S(n3095), .Z(n5259) );
  MUX2_X2 U4909 ( .A(u3_N57), .B(u3_N29), .S(n3095), .Z(n5260) );
  MUX2_X2 U4910 ( .A(u3_N56), .B(u3_N28), .S(n3095), .Z(n5261) );
  MUX2_X2 U4911 ( .A(u3_N55), .B(u3_N27), .S(n3095), .Z(n5262) );
  MUX2_X2 U4912 ( .A(u3_N54), .B(u3_N26), .S(n3095), .Z(n5263) );
  MUX2_X2 U4913 ( .A(u3_N53), .B(u3_N25), .S(n3095), .Z(n5264) );
  MUX2_X2 U4914 ( .A(u3_N52), .B(u3_N24), .S(n3095), .Z(n5265) );
  MUX2_X2 U4915 ( .A(u3_N51), .B(u3_N23), .S(n3095), .Z(n5266) );
  MUX2_X2 U4916 ( .A(u3_N50), .B(u3_N22), .S(n3095), .Z(n5267) );
  MUX2_X2 U4917 ( .A(u3_N49), .B(u3_N21), .S(n3095), .Z(n5268) );
  MUX2_X2 U4918 ( .A(u3_N48), .B(u3_N20), .S(n3095), .Z(n5269) );
  MUX2_X2 U4919 ( .A(u3_N47), .B(u3_N19), .S(n2570), .Z(n5270) );
  MUX2_X2 U4920 ( .A(u3_N46), .B(u3_N18), .S(n3095), .Z(n5271) );
  MUX2_X2 U4921 ( .A(u3_N45), .B(u3_N17), .S(n3095), .Z(n5272) );
  MUX2_X2 U4922 ( .A(u3_N44), .B(u3_N16), .S(n2570), .Z(n5273) );
  MUX2_X2 U4923 ( .A(u3_N43), .B(u3_N15), .S(n3095), .Z(n5274) );
  MUX2_X2 U4924 ( .A(u3_N42), .B(u3_N14), .S(n2570), .Z(n5275) );
  MUX2_X2 U4925 ( .A(u3_N41), .B(u3_N13), .S(n2570), .Z(n5276) );
  MUX2_X2 U4926 ( .A(u3_N40), .B(u3_N12), .S(n2570), .Z(n5277) );
  MUX2_X2 U4927 ( .A(u3_N39), .B(u3_N11), .S(n2570), .Z(n5278) );
  MUX2_X2 U4928 ( .A(u3_N38), .B(u3_N10), .S(n2570), .Z(n5279) );
  MUX2_X2 U4929 ( .A(u3_N37), .B(u3_N9), .S(n2570), .Z(n5280) );
  MUX2_X2 U4930 ( .A(u3_N36), .B(u3_N8), .S(n3095), .Z(n5281) );
  MUX2_X2 U4931 ( .A(u3_N35), .B(u3_N7), .S(n2570), .Z(n5282) );
  MUX2_X2 U4932 ( .A(u3_N34), .B(u3_N6), .S(n3095), .Z(n5283) );
  MUX2_X2 U4933 ( .A(u3_N33), .B(u3_N5), .S(n2570), .Z(n5284) );
  MUX2_X2 U4934 ( .A(u3_N32), .B(u3_N4), .S(n3095), .Z(n5285) );
  MUX2_X2 U4935 ( .A(u3_N31), .B(u3_N3), .S(n2570), .Z(n5286) );
  MUX2_X2 U4936 ( .A(n2930), .B(u2_N124), .S(n3076), .Z(n2459) );
  MUX2_X2 U4937 ( .A(u6_N22), .B(fracta_mul[22]), .S(n3077), .Z(u1_adj_op_22_)
         );
  MUX2_X2 U4938 ( .A(n3049), .B(fracta_mul[21]), .S(n3078), .Z(n5300) );
  MUX2_X2 U4939 ( .A(n3040), .B(fracta_mul[20]), .S(n3076), .Z(u1_adj_op_20_)
         );
  MUX2_X2 U4940 ( .A(n2968), .B(fracta_mul[19]), .S(n3077), .Z(u1_adj_op_19_)
         );
  MUX2_X2 U4941 ( .A(u6_N18), .B(fracta_mul[18]), .S(n3078), .Z(u1_adj_op_18_)
         );
  MUX2_X2 U4942 ( .A(u6_N17), .B(fracta_mul[17]), .S(n3076), .Z(u1_adj_op_17_)
         );
  MUX2_X2 U4943 ( .A(n2963), .B(fracta_mul[16]), .S(n3077), .Z(n5302) );
  MUX2_X2 U4944 ( .A(u6_N15), .B(fracta_mul[15]), .S(n3078), .Z(n5303) );
  MUX2_X2 U4945 ( .A(n2672), .B(fracta_mul[14]), .S(n3076), .Z(n5304) );
  MUX2_X2 U4946 ( .A(u6_N13), .B(fracta_mul[13]), .S(n3077), .Z(n5305) );
  MUX2_X2 U4947 ( .A(n2986), .B(fracta_mul[12]), .S(n3078), .Z(n5306) );
  MUX2_X2 U4948 ( .A(n2982), .B(fracta_mul[11]), .S(n3076), .Z(n5307) );
  MUX2_X2 U4949 ( .A(u6_N10), .B(fracta_mul[10]), .S(n3077), .Z(u1_adj_op_10_)
         );
  MUX2_X2 U4950 ( .A(n4597), .B(n2681), .S(n3078), .Z(n4478) );
  INV_X4 U4951 ( .A(n4478), .ZN(n5292) );
  MUX2_X2 U4952 ( .A(n4592), .B(n2695), .S(n3076), .Z(n4479) );
  INV_X4 U4953 ( .A(n4479), .ZN(n5293) );
  MUX2_X2 U4954 ( .A(n4517), .B(n2689), .S(n3077), .Z(n4539) );
  INV_X4 U4955 ( .A(n4539), .ZN(n5294) );
  MUX2_X2 U4956 ( .A(n2589), .B(n2685), .S(n3078), .Z(n4538) );
  INV_X4 U4957 ( .A(n4538), .ZN(n5295) );
  MUX2_X2 U4958 ( .A(n2706), .B(n2596), .S(n3077), .Z(n4537) );
  INV_X4 U4959 ( .A(n4537), .ZN(n5296) );
  MUX2_X2 U4960 ( .A(n2705), .B(n2690), .S(n3078), .Z(n4535) );
  INV_X4 U4961 ( .A(n4535), .ZN(n5297) );
  MUX2_X2 U4962 ( .A(n2703), .B(n2598), .S(n3076), .Z(n4533) );
  INV_X4 U4963 ( .A(n4533), .ZN(n5298) );
  MUX2_X2 U4964 ( .A(n2702), .B(n4524), .S(n3077), .Z(n4531) );
  INV_X4 U4965 ( .A(n4531), .ZN(n5299) );
  MUX2_X2 U4966 ( .A(n2701), .B(n4523), .S(n3078), .Z(n4532) );
  INV_X4 U4967 ( .A(n4532), .ZN(n5301) );
  MUX2_X2 U4968 ( .A(n2708), .B(n4530), .S(n3076), .Z(n4540) );
  INV_X4 U4969 ( .A(n4540), .ZN(n5308) );
  MUX2_X2 U4970 ( .A(opb_r[30]), .B(opa_r[30]), .S(n3076), .Z(u1_exp_small[7])
         );
  MUX2_X2 U4971 ( .A(opb_r[29]), .B(opa_r[29]), .S(n3077), .Z(u1_exp_small[6])
         );
  MUX2_X2 U4972 ( .A(opb_r[28]), .B(opa_r[28]), .S(n3078), .Z(u1_exp_small[5])
         );
  MUX2_X2 U4973 ( .A(opb_r[27]), .B(opa_r[27]), .S(n3076), .Z(u1_exp_small[4])
         );
  MUX2_X2 U4974 ( .A(opb_r[26]), .B(opa_r[26]), .S(n3077), .Z(u1_exp_small[3])
         );
  MUX2_X2 U4975 ( .A(opb_r[25]), .B(opa_r[25]), .S(n3078), .Z(u1_exp_small[2])
         );
  MUX2_X2 U4976 ( .A(opb_r[24]), .B(opa_r[24]), .S(n3076), .Z(u1_exp_small[1])
         );
  MUX2_X2 U4977 ( .A(opb_r[23]), .B(opa_r[23]), .S(n3077), .Z(u1_exp_small[0])
         );
  NAND2_X2 U4978 ( .A1(n4765), .A2(n4764), .ZN(n4488) );
  INV_X4 U4979 ( .A(n4488), .ZN(n4486) );
  INV_X4 U4980 ( .A(u1_exp_diff2[4]), .ZN(n4485) );
  NOR2_X4 U4981 ( .A1(u1_exp_diff2[7]), .A2(u1_exp_diff2[6]), .ZN(n4480) );
  INV_X4 U4982 ( .A(n4480), .ZN(n4484) );
  INV_X4 U4983 ( .A(u1_exp_diff2[5]), .ZN(n4481) );
  NAND2_X2 U4984 ( .A1(n4482), .A2(n4481), .ZN(n4483) );
  OAI21_X4 U4985 ( .B1(n4484), .B2(n4483), .A(n4488), .ZN(n4487) );
  OAI21_X4 U4986 ( .B1(n4486), .B2(n4485), .A(n4487), .ZN(u1_exp_diff_sft_4_)
         );
  INV_X4 U4987 ( .A(n4544), .ZN(n5288) );
  OAI21_X4 U4988 ( .B1(u1_exp_diff2[1]), .B2(n4489), .A(n4488), .ZN(n4553) );
  OAI21_X4 U4989 ( .B1(u1_exp_diff2[0]), .B2(n4489), .A(n4488), .ZN(n4551) );
  INV_X4 U4990 ( .A(u1_adj_op_out_sft_26_), .ZN(n4490) );
  MUX2_X2 U4991 ( .A(n4490), .B(n4765), .S(n3078), .Z(n4650) );
  NAND2_X2 U4992 ( .A1(n4490), .A2(n3076), .ZN(n4675) );
  INV_X4 U4993 ( .A(n4675), .ZN(n4493) );
  NAND2_X2 U4994 ( .A1(n4650), .A2(n4493), .ZN(u1_fracta_s[26]) );
  INV_X4 U4995 ( .A(u1_adj_op_out_sft_25_), .ZN(n4492) );
  MUX2_X2 U4996 ( .A(n4492), .B(n4491), .S(n3076), .Z(n4644) );
  INV_X4 U4997 ( .A(n4644), .ZN(n4676) );
  MUX2_X2 U4998 ( .A(n2591), .B(n4492), .S(n3077), .Z(n4645) );
  INV_X4 U4999 ( .A(n4645), .ZN(n4677) );
  INV_X4 U5000 ( .A(n4650), .ZN(n4674) );
  NOR2_X4 U5001 ( .A1(n4674), .A2(n4493), .ZN(n4494) );
  NOR2_X4 U5002 ( .A1(n4495), .A2(n4494), .ZN(n4653) );
  INV_X4 U5003 ( .A(u1_adj_op_out_sft_21_), .ZN(n4497) );
  MUX2_X2 U5004 ( .A(n2677), .B(n4497), .S(n3078), .Z(n4656) );
  MUX2_X2 U5005 ( .A(n4497), .B(n4496), .S(n3076), .Z(n4631) );
  INV_X4 U5006 ( .A(n4631), .ZN(n4684) );
  INV_X4 U5007 ( .A(u1_adj_op_out_sft_22_), .ZN(n4499) );
  MUX2_X2 U5008 ( .A(n4499), .B(n2679), .S(n3077), .Z(n4498) );
  INV_X4 U5009 ( .A(n4498), .ZN(n4682) );
  MUX2_X2 U5010 ( .A(n2592), .B(n4499), .S(n3078), .Z(n4655) );
  INV_X4 U5011 ( .A(u1_adj_op_out_sft_17_), .ZN(n4503) );
  MUX2_X2 U5012 ( .A(n2687), .B(n4503), .S(n3076), .Z(n4659) );
  MUX2_X2 U5013 ( .A(n4503), .B(n4502), .S(n3077), .Z(n4617) );
  INV_X4 U5014 ( .A(n4617), .ZN(n4692) );
  INV_X4 U5015 ( .A(u1_adj_op_out_sft_18_), .ZN(n4506) );
  MUX2_X2 U5016 ( .A(n4506), .B(n4504), .S(n3078), .Z(n4505) );
  INV_X4 U5017 ( .A(n4505), .ZN(n4690) );
  MUX2_X2 U5018 ( .A(n2696), .B(n4506), .S(n3076), .Z(n4658) );
  INV_X4 U5019 ( .A(u1_adj_op_out_sft_13_), .ZN(n4510) );
  MUX2_X2 U5020 ( .A(n2593), .B(n4510), .S(n3077), .Z(n4662) );
  MUX2_X2 U5021 ( .A(n4510), .B(n4509), .S(n3078), .Z(n4602) );
  INV_X4 U5022 ( .A(n4602), .ZN(n4700) );
  INV_X4 U5023 ( .A(u1_adj_op_out_sft_14_), .ZN(n4513) );
  MUX2_X2 U5024 ( .A(n4513), .B(n4511), .S(n3076), .Z(n4512) );
  INV_X4 U5025 ( .A(n4512), .ZN(n4698) );
  MUX2_X2 U5026 ( .A(n2697), .B(n4513), .S(n3077), .Z(n4661) );
  INV_X4 U5027 ( .A(u1_adj_op_out_sft_9_), .ZN(n4516) );
  MUX2_X2 U5028 ( .A(n2685), .B(n4516), .S(n3078), .Z(n4665) );
  MUX2_X2 U5029 ( .A(n4516), .B(n2589), .S(n3076), .Z(n4587) );
  INV_X4 U5030 ( .A(n4587), .ZN(n4708) );
  INV_X4 U5031 ( .A(u1_adj_op_out_sft_10_), .ZN(n4519) );
  MUX2_X2 U5032 ( .A(n4519), .B(n4517), .S(n3077), .Z(n4518) );
  INV_X4 U5033 ( .A(n4518), .ZN(n4706) );
  MUX2_X2 U5034 ( .A(n2689), .B(n4519), .S(n3078), .Z(n4664) );
  INV_X4 U5035 ( .A(u1_adj_op_out_sft_4_), .ZN(n4522) );
  MUX2_X2 U5036 ( .A(n4522), .B(n2701), .S(n3076), .Z(n4667) );
  MUX2_X2 U5037 ( .A(n4523), .B(n4522), .S(n3077), .Z(n4528) );
  INV_X4 U5038 ( .A(n4528), .ZN(n4719) );
  NOR2_X4 U5039 ( .A1(n4667), .A2(n4719), .ZN(n4527) );
  INV_X4 U5040 ( .A(u1_adj_op_out_sft_5_), .ZN(n4525) );
  MUX2_X2 U5041 ( .A(n4524), .B(n4525), .S(n3078), .Z(n4570) );
  INV_X4 U5042 ( .A(n4570), .ZN(n4717) );
  MUX2_X2 U5043 ( .A(n4525), .B(n2702), .S(n3076), .Z(n4569) );
  NOR2_X4 U5044 ( .A1(n4717), .A2(n4569), .ZN(n4526) );
  NOR2_X4 U5045 ( .A1(n4527), .A2(n4526), .ZN(n4573) );
  NAND2_X2 U5046 ( .A1(n4719), .A2(n4667), .ZN(n4568) );
  INV_X4 U5047 ( .A(u1_adj_op_out_sft_3_), .ZN(n4529) );
  MUX2_X2 U5048 ( .A(n4529), .B(n2708), .S(n3077), .Z(n4565) );
  INV_X4 U5049 ( .A(n4565), .ZN(n4720) );
  MUX2_X2 U5050 ( .A(n4530), .B(n4529), .S(n3078), .Z(n4564) );
  NAND2_X2 U5051 ( .A1(n4720), .A2(n4564), .ZN(n4563) );
  NAND2_X2 U5052 ( .A1(u1_adj_op_out_sft_2_), .A2(n4672), .ZN(n4668) );
  NAND2_X2 U5053 ( .A1(u1_adj_op_out_sft_1_), .A2(n4672), .ZN(n4669) );
  NAND2_X2 U5054 ( .A1(n2722), .A2(n4533), .ZN(n4534) );
  INV_X4 U5055 ( .A(n4534), .ZN(n4545) );
  NAND2_X2 U5056 ( .A1(n4545), .A2(n4535), .ZN(n4536) );
  INV_X4 U5057 ( .A(n4536), .ZN(n4554) );
  NAND2_X2 U5058 ( .A1(n2715), .A2(n4539), .ZN(n4550) );
  OAI21_X4 U5059 ( .B1(n4543), .B2(n4542), .A(n5288), .ZN(n4549) );
  NAND2_X2 U5060 ( .A1(n4547), .A2(n4546), .ZN(n4548) );
  MUX2_X2 U5061 ( .A(n4549), .B(n4548), .S(n5290), .Z(n4560) );
  OAI21_X4 U5062 ( .B1(n4558), .B2(n4557), .A(n4556), .ZN(n4559) );
  NOR2_X4 U5063 ( .A1(u1_adj_op_out_sft_0_), .A2(n4561), .ZN(n4673) );
  INV_X4 U5064 ( .A(n4673), .ZN(n4562) );
  NAND4_X2 U5065 ( .A1(n4563), .A2(n4668), .A3(n4669), .A4(n4671), .ZN(n4567)
         );
  INV_X4 U5066 ( .A(n4564), .ZN(n4721) );
  NAND2_X2 U5067 ( .A1(n4565), .A2(n4721), .ZN(n4566) );
  NAND3_X4 U5068 ( .A1(n4568), .A2(n4567), .A3(n4566), .ZN(n4572) );
  INV_X4 U5069 ( .A(n4569), .ZN(n4716) );
  AOI21_X4 U5070 ( .B1(n4573), .B2(n4572), .A(n4571), .ZN(n4582) );
  INV_X4 U5071 ( .A(u1_adj_op_out_sft_6_), .ZN(n4574) );
  MUX2_X2 U5072 ( .A(n2598), .B(n4574), .S(n3076), .Z(n4576) );
  INV_X4 U5073 ( .A(n4576), .ZN(n4715) );
  MUX2_X2 U5074 ( .A(n4574), .B(n2703), .S(n3077), .Z(n4575) );
  NAND2_X2 U5075 ( .A1(n4715), .A2(n4575), .ZN(n4581) );
  INV_X4 U5076 ( .A(n4575), .ZN(n4714) );
  NAND2_X2 U5077 ( .A1(n4576), .A2(n4714), .ZN(n4577) );
  INV_X4 U5078 ( .A(n4577), .ZN(n4580) );
  INV_X4 U5079 ( .A(u1_adj_op_out_sft_7_), .ZN(n4578) );
  MUX2_X2 U5080 ( .A(n2690), .B(n4578), .S(n3078), .Z(n4586) );
  INV_X4 U5081 ( .A(n4586), .ZN(n4713) );
  MUX2_X2 U5082 ( .A(n4578), .B(n2705), .S(n3076), .Z(n4585) );
  NOR2_X4 U5083 ( .A1(n4713), .A2(n4585), .ZN(n4579) );
  AOI211_X4 U5084 ( .C1(n4582), .C2(n4581), .A(n4580), .B(n4579), .ZN(n4591)
         );
  INV_X4 U5085 ( .A(u1_adj_op_out_sft_8_), .ZN(n4584) );
  MUX2_X2 U5086 ( .A(n4584), .B(n2706), .S(n3077), .Z(n4583) );
  INV_X4 U5087 ( .A(n4583), .ZN(n4710) );
  MUX2_X2 U5088 ( .A(n2596), .B(n4584), .S(n3078), .Z(n4666) );
  INV_X4 U5089 ( .A(n4585), .ZN(n4712) );
  OAI22_X2 U5090 ( .A1(n4710), .A2(n4666), .B1(n4586), .B2(n4712), .ZN(n4590)
         );
  NAND2_X2 U5091 ( .A1(n4708), .A2(n4665), .ZN(n4589) );
  NAND2_X2 U5092 ( .A1(n4666), .A2(n4710), .ZN(n4588) );
  INV_X4 U5093 ( .A(u1_adj_op_out_sft_11_), .ZN(n4593) );
  MUX2_X2 U5094 ( .A(n2695), .B(n4593), .S(n3076), .Z(n4601) );
  INV_X4 U5095 ( .A(n4601), .ZN(n4705) );
  MUX2_X2 U5096 ( .A(n4593), .B(n4592), .S(n3077), .Z(n4600) );
  AOI211_X4 U5097 ( .C1(n4596), .C2(n4595), .A(n2664), .B(n4594), .ZN(n4606)
         );
  INV_X4 U5098 ( .A(u1_adj_op_out_sft_12_), .ZN(n4599) );
  MUX2_X2 U5099 ( .A(n4599), .B(n4597), .S(n3078), .Z(n4598) );
  INV_X4 U5100 ( .A(n4598), .ZN(n4702) );
  MUX2_X2 U5101 ( .A(n2681), .B(n4599), .S(n3076), .Z(n4663) );
  INV_X4 U5102 ( .A(n4600), .ZN(n4704) );
  OAI22_X2 U5103 ( .A1(n4702), .A2(n4663), .B1(n4601), .B2(n4704), .ZN(n4605)
         );
  NAND2_X2 U5104 ( .A1(n4700), .A2(n4662), .ZN(n4604) );
  NAND2_X2 U5105 ( .A1(n4663), .A2(n4702), .ZN(n4603) );
  INV_X4 U5106 ( .A(u1_adj_op_out_sft_15_), .ZN(n4608) );
  MUX2_X2 U5107 ( .A(n2692), .B(n4608), .S(n3077), .Z(n4616) );
  INV_X4 U5108 ( .A(n4616), .ZN(n4697) );
  MUX2_X2 U5109 ( .A(n4608), .B(n4607), .S(n3078), .Z(n4615) );
  NOR2_X4 U5110 ( .A1(n4697), .A2(n4615), .ZN(n4609) );
  AOI211_X4 U5111 ( .C1(n4611), .C2(n4610), .A(n2724), .B(n4609), .ZN(n4621)
         );
  INV_X4 U5112 ( .A(u1_adj_op_out_sft_16_), .ZN(n4614) );
  INV_X4 U5113 ( .A(u6_N13), .ZN(n4612) );
  MUX2_X2 U5114 ( .A(n4614), .B(n4612), .S(n3076), .Z(n4613) );
  INV_X4 U5115 ( .A(n4613), .ZN(n4694) );
  MUX2_X2 U5116 ( .A(n2678), .B(n4614), .S(n3077), .Z(n4660) );
  INV_X4 U5117 ( .A(n4615), .ZN(n4696) );
  OAI22_X2 U5118 ( .A1(n4694), .A2(n4660), .B1(n4616), .B2(n4696), .ZN(n4620)
         );
  NAND2_X2 U5119 ( .A1(n4692), .A2(n4659), .ZN(n4619) );
  NAND2_X2 U5120 ( .A1(n4660), .A2(n4694), .ZN(n4618) );
  INV_X4 U5121 ( .A(u1_adj_op_out_sft_19_), .ZN(n4622) );
  MUX2_X2 U5122 ( .A(n2675), .B(n4622), .S(n3078), .Z(n4630) );
  INV_X4 U5123 ( .A(n4630), .ZN(n4689) );
  MUX2_X2 U5124 ( .A(n4622), .B(n2680), .S(n3076), .Z(n4629) );
  NOR2_X4 U5125 ( .A1(n4689), .A2(n4629), .ZN(n4623) );
  AOI211_X4 U5126 ( .C1(n4625), .C2(n4624), .A(n2725), .B(n4623), .ZN(n4635)
         );
  INV_X4 U5127 ( .A(u1_adj_op_out_sft_20_), .ZN(n4628) );
  MUX2_X2 U5128 ( .A(n4628), .B(n4626), .S(n3077), .Z(n4627) );
  INV_X4 U5129 ( .A(n4627), .ZN(n4686) );
  MUX2_X2 U5130 ( .A(n2590), .B(n4628), .S(n3078), .Z(n4657) );
  INV_X4 U5131 ( .A(n4629), .ZN(n4688) );
  OAI22_X2 U5132 ( .A1(n4686), .A2(n4657), .B1(n4630), .B2(n4688), .ZN(n4634)
         );
  NAND2_X2 U5133 ( .A1(n4684), .A2(n4656), .ZN(n4633) );
  NAND2_X2 U5134 ( .A1(n4657), .A2(n4686), .ZN(n4632) );
  INV_X4 U5135 ( .A(u1_adj_op_out_sft_23_), .ZN(n4636) );
  MUX2_X2 U5136 ( .A(n2683), .B(n4636), .S(n3076), .Z(n4643) );
  INV_X4 U5137 ( .A(n4643), .ZN(n4681) );
  MUX2_X2 U5138 ( .A(n4636), .B(n2682), .S(n3077), .Z(n4642) );
  NOR2_X4 U5139 ( .A1(n4681), .A2(n4642), .ZN(n4637) );
  AOI211_X4 U5140 ( .C1(n4639), .C2(n4638), .A(n2726), .B(n4637), .ZN(n4649)
         );
  INV_X4 U5141 ( .A(u1_adj_op_out_sft_24_), .ZN(n4641) );
  MUX2_X2 U5142 ( .A(n4641), .B(n2693), .S(n3078), .Z(n4640) );
  INV_X4 U5143 ( .A(n4640), .ZN(n4678) );
  MUX2_X2 U5144 ( .A(n2599), .B(n4641), .S(n3076), .Z(n4654) );
  INV_X4 U5145 ( .A(n4642), .ZN(n4680) );
  OAI22_X2 U5146 ( .A1(n4678), .A2(n4654), .B1(n4643), .B2(n4680), .ZN(n4648)
         );
  NAND2_X2 U5147 ( .A1(n4676), .A2(n4645), .ZN(n4647) );
  NAND2_X2 U5148 ( .A1(n4654), .A2(n4678), .ZN(n4646) );
  AOI21_X4 U5149 ( .B1(n4653), .B2(n4652), .A(n4651), .ZN(n4726) );
  MUX2_X2 U5150 ( .A(n4676), .B(n4677), .S(n3080), .Z(u1_fracta_s[25]) );
  INV_X4 U5151 ( .A(n4654), .ZN(n4679) );
  MUX2_X2 U5152 ( .A(n4678), .B(n4679), .S(n3081), .Z(u1_fracta_s[24]) );
  MUX2_X2 U5153 ( .A(n4680), .B(n4681), .S(n3082), .Z(u1_fracta_s[23]) );
  INV_X4 U5154 ( .A(n4655), .ZN(n4683) );
  MUX2_X2 U5155 ( .A(n4682), .B(n4683), .S(n3083), .Z(u1_fracta_s[22]) );
  INV_X4 U5156 ( .A(n4656), .ZN(n4685) );
  MUX2_X2 U5157 ( .A(n4684), .B(n4685), .S(n3084), .Z(u1_fracta_s[21]) );
  INV_X4 U5158 ( .A(n4657), .ZN(n4687) );
  MUX2_X2 U5159 ( .A(n4686), .B(n4687), .S(n3084), .Z(u1_fracta_s[20]) );
  MUX2_X2 U5160 ( .A(n4688), .B(n4689), .S(n3080), .Z(u1_fracta_s[19]) );
  INV_X4 U5161 ( .A(n4658), .ZN(n4691) );
  MUX2_X2 U5162 ( .A(n4690), .B(n4691), .S(n3081), .Z(u1_fracta_s[18]) );
  INV_X4 U5163 ( .A(n4659), .ZN(n4693) );
  MUX2_X2 U5164 ( .A(n4692), .B(n4693), .S(n3082), .Z(u1_fracta_s[17]) );
  INV_X4 U5165 ( .A(n4660), .ZN(n4695) );
  MUX2_X2 U5166 ( .A(n4694), .B(n4695), .S(n3080), .Z(u1_fracta_s[16]) );
  MUX2_X2 U5167 ( .A(n4696), .B(n4697), .S(n3083), .Z(u1_fracta_s[15]) );
  INV_X4 U5168 ( .A(n4661), .ZN(n4699) );
  MUX2_X2 U5169 ( .A(n4698), .B(n4699), .S(n3084), .Z(u1_fracta_s[14]) );
  INV_X4 U5170 ( .A(n4662), .ZN(n4701) );
  MUX2_X2 U5171 ( .A(n4700), .B(n4701), .S(n3080), .Z(u1_fracta_s[13]) );
  INV_X4 U5172 ( .A(n4663), .ZN(n4703) );
  MUX2_X2 U5173 ( .A(n4702), .B(n4703), .S(n3081), .Z(u1_fracta_s[12]) );
  MUX2_X2 U5174 ( .A(n4704), .B(n4705), .S(n3081), .Z(u1_fracta_s[11]) );
  INV_X4 U5175 ( .A(n4664), .ZN(n4707) );
  MUX2_X2 U5176 ( .A(n4706), .B(n4707), .S(n3082), .Z(u1_fracta_s[10]) );
  INV_X4 U5177 ( .A(n4665), .ZN(n4709) );
  MUX2_X2 U5178 ( .A(n4708), .B(n4709), .S(n3083), .Z(u1_fracta_s[9]) );
  INV_X4 U5179 ( .A(n4666), .ZN(n4711) );
  MUX2_X2 U5180 ( .A(n4710), .B(n4711), .S(n3084), .Z(u1_fracta_s[8]) );
  MUX2_X2 U5181 ( .A(n4712), .B(n4713), .S(n3080), .Z(u1_fracta_s[7]) );
  MUX2_X2 U5182 ( .A(n4714), .B(n4715), .S(n3082), .Z(u1_fracta_s[6]) );
  MUX2_X2 U5183 ( .A(n4716), .B(n4717), .S(n3081), .Z(u1_fracta_s[5]) );
  INV_X4 U5184 ( .A(n4667), .ZN(n4718) );
  MUX2_X2 U5185 ( .A(n4718), .B(n4719), .S(n3082), .Z(u1_fracta_s[4]) );
  MUX2_X2 U5186 ( .A(n4720), .B(n4721), .S(n3083), .Z(u1_fracta_s[3]) );
  INV_X4 U5187 ( .A(n4668), .ZN(n4722) );
  MUX2_X2 U5188 ( .A(n4722), .B(n2720), .S(n3084), .Z(u1_fracta_s[2]) );
  INV_X4 U5189 ( .A(n4669), .ZN(n4723) );
  MUX2_X2 U5190 ( .A(n4723), .B(n2721), .S(n3083), .Z(u1_fracta_s[1]) );
  INV_X4 U5191 ( .A(n4671), .ZN(n4724) );
  MUX2_X2 U5192 ( .A(n4724), .B(n4725), .S(n3080), .Z(u1_fracta_s[0]) );
  MUX2_X2 U5193 ( .A(n4675), .B(n4674), .S(n3081), .Z(u1_fractb_s[26]) );
  MUX2_X2 U5194 ( .A(n4677), .B(n4676), .S(n3082), .Z(u1_fractb_s[25]) );
  MUX2_X2 U5195 ( .A(n4679), .B(n4678), .S(n3083), .Z(u1_fractb_s[24]) );
  MUX2_X2 U5196 ( .A(n4681), .B(n4680), .S(n3084), .Z(u1_fractb_s[23]) );
  MUX2_X2 U5197 ( .A(n4683), .B(n4682), .S(n3084), .Z(u1_fractb_s[22]) );
  MUX2_X2 U5198 ( .A(n4685), .B(n4684), .S(n3080), .Z(u1_fractb_s[21]) );
  MUX2_X2 U5199 ( .A(n4687), .B(n4686), .S(n3081), .Z(u1_fractb_s[20]) );
  MUX2_X2 U5200 ( .A(n4689), .B(n4688), .S(n3082), .Z(u1_fractb_s[19]) );
  MUX2_X2 U5201 ( .A(n4691), .B(n4690), .S(n3080), .Z(u1_fractb_s[18]) );
  MUX2_X2 U5202 ( .A(n4693), .B(n4692), .S(n3083), .Z(u1_fractb_s[17]) );
  MUX2_X2 U5203 ( .A(n4695), .B(n4694), .S(n3084), .Z(u1_fractb_s[16]) );
  MUX2_X2 U5204 ( .A(n4697), .B(n4696), .S(n3080), .Z(u1_fractb_s[15]) );
  MUX2_X2 U5205 ( .A(n4699), .B(n4698), .S(n3081), .Z(u1_fractb_s[14]) );
  MUX2_X2 U5206 ( .A(n4701), .B(n4700), .S(n3081), .Z(u1_fractb_s[13]) );
  MUX2_X2 U5207 ( .A(n4703), .B(n4702), .S(n3082), .Z(u1_fractb_s[12]) );
  MUX2_X2 U5208 ( .A(n4705), .B(n4704), .S(n3083), .Z(u1_fractb_s[11]) );
  MUX2_X2 U5209 ( .A(n4707), .B(n4706), .S(n3084), .Z(u1_fractb_s[10]) );
  MUX2_X2 U5210 ( .A(n4709), .B(n4708), .S(n3080), .Z(u1_fractb_s[9]) );
  MUX2_X2 U5211 ( .A(n4711), .B(n4710), .S(n3082), .Z(u1_fractb_s[8]) );
  MUX2_X2 U5212 ( .A(n4713), .B(n4712), .S(n3081), .Z(u1_fractb_s[7]) );
  MUX2_X2 U5213 ( .A(n4715), .B(n4714), .S(n3082), .Z(u1_fractb_s[6]) );
  MUX2_X2 U5214 ( .A(n4717), .B(n4716), .S(n3083), .Z(u1_fractb_s[5]) );
  MUX2_X2 U5215 ( .A(n4719), .B(n4718), .S(n3084), .Z(u1_fractb_s[4]) );
  MUX2_X2 U5216 ( .A(n4721), .B(n4720), .S(n3083), .Z(u1_fractb_s[3]) );
  MUX2_X2 U5217 ( .A(n2720), .B(n4722), .S(n3080), .Z(u1_fractb_s[2]) );
  MUX2_X2 U5218 ( .A(n2721), .B(n4723), .S(n3081), .Z(u1_fractb_s[1]) );
  MUX2_X2 U5219 ( .A(n4725), .B(n4724), .S(n3082), .Z(u1_fractb_s[0]) );
  XOR2_X2 U5220 ( .A(opb_r[31]), .B(fpu_op_r1[0]), .Z(n4727) );
  MUX2_X2 U5221 ( .A(n4727), .B(opa_r[31]), .S(n3083), .Z(u1_sign_d) );
  INV_X4 U5222 ( .A(n4728), .ZN(n4729) );
  NAND2_X2 U5223 ( .A1(n4733), .A2(n4732), .ZN(n4743) );
  INV_X4 U5224 ( .A(n4743), .ZN(n4761) );
  NAND2_X2 U5225 ( .A1(n4740), .A2(n4739), .ZN(n4744) );
  INV_X4 U5226 ( .A(n4744), .ZN(n4760) );
  INV_X4 U5227 ( .A(n4741), .ZN(n4762) );
  INV_X4 U5228 ( .A(n4742), .ZN(n4763) );
  NAND2_X2 U5229 ( .A1(net82035), .A2(net82036), .ZN(n4746) );
  NAND3_X2 U5230 ( .A1(net82030), .A2(n4746), .A3(n4745), .ZN(n4759) );
  XNOR2_X2 U5231 ( .A(n4747), .B(net82029), .ZN(n4748) );
  AOI221_X2 U5232 ( .B1(u4_div_shft3_7_), .B2(n4754), .C1(u4_div_shft4[7]), 
        .C2(n4755), .A(n4750), .ZN(net82024) );
  XNOR2_X2 U5233 ( .A(n4751), .B(n2618), .ZN(n4752) );
  AOI221_X2 U5234 ( .B1(u4_div_shft4[6]), .B2(n4755), .C1(u4_div_shft3_6_), 
        .C2(n4754), .A(n2528), .ZN(net82014) );
  OR3_X1 U5235 ( .A1(n3085), .A2(n3087), .A3(n3089), .ZN(n4766) );
  AND3_X1 U5236 ( .A1(n3091), .A2(net85905), .A3(n3089), .ZN(n4767) );
  OAI21_X1 U5237 ( .B1(n3087), .B2(n4767), .A(n3085), .ZN(n4768) );
  NOR4_X1 U5238 ( .A1(net85937), .A2(net85933), .A3(net85929), .A4(n4769), 
        .ZN(u4_N1600) );
  INV_X4 U5239 ( .A(n4768), .ZN(n4769) );
  AND3_X1 U5240 ( .A1(n3091), .A2(net85905), .A3(n3089), .ZN(n4770) );
  OAI21_X1 U5241 ( .B1(n4770), .B2(n3088), .A(n3085), .ZN(n4771) );
  OR4_X1 U5242 ( .A1(net85929), .A2(n4772), .A3(net85937), .A4(net85933), .ZN(
        u4_N1598) );
  INV_X4 U5243 ( .A(n4771), .ZN(n4772) );
  INV_X4 U5244 ( .A(n2600), .ZN(n5287) );
  INV_X4 U5245 ( .A(n1746), .ZN(n5318) );
  INV_X4 U5246 ( .A(n2445), .ZN(n5319) );
  INV_X4 U5247 ( .A(n1730), .ZN(n5327) );
  INV_X4 U5248 ( .A(n1731), .ZN(n5328) );
  INV_X4 U5249 ( .A(n1732), .ZN(n5329) );
  INV_X4 U5250 ( .A(n1733), .ZN(n5330) );
  INV_X4 u4_sub_472_U14 ( .A(u4_fi_ldz_mi1_5_), .ZN(u4_sub_472_n7) );
  INV_X1 u4_sub_472_U13 ( .A(u4_fi_ldz_mi1_2_), .ZN(u4_sub_472_n4) );
  INV_X1 u4_sub_472_U12 ( .A(n4757), .ZN(u4_sub_472_n9) );
  INV_X4 u4_sub_472_U11 ( .A(u4_sub_472_carry_6_), .ZN(u4_sub_472_n3) );
  INV_X4 u4_sub_472_U10 ( .A(net85933), .ZN(u4_sub_472_n2) );
  XNOR2_X2 u4_sub_472_U9 ( .A(net85933), .B(u4_sub_472_carry_6_), .ZN(
        u4_exp_fix_divb[6]) );
  NAND2_X2 u4_sub_472_U8 ( .A1(u4_sub_472_n2), .A2(u4_sub_472_n3), .ZN(
        u4_sub_472_carry_7_) );
  INV_X4 u4_sub_472_U7 ( .A(net85905), .ZN(u4_sub_472_n1) );
  NAND2_X2 u4_sub_472_U6 ( .A1(n4757), .A2(u4_sub_472_n1), .ZN(
        u4_sub_472_carry_1_) );
  XNOR2_X2 u4_sub_472_U5 ( .A(net85937), .B(u4_sub_472_carry_7_), .ZN(
        u4_exp_fix_divb[7]) );
  INV_X1 u4_sub_472_U4 ( .A(u4_fi_ldz_mi1_4_), .ZN(u4_sub_472_n6) );
  INV_X1 u4_sub_472_U3 ( .A(n2500), .ZN(u4_sub_472_n8) );
  INV_X1 u4_sub_472_U2 ( .A(u4_fi_ldz_mi1_3_), .ZN(u4_sub_472_n5) );
  XNOR2_X1 u4_sub_472_U1 ( .A(u4_sub_472_n9), .B(net85905), .ZN(
        u4_exp_fix_divb[0]) );
  FA_X1 u4_sub_472_U2_1 ( .A(n3091), .B(u4_sub_472_n8), .CI(
        u4_sub_472_carry_1_), .CO(u4_sub_472_carry_2_), .S(u4_exp_fix_divb[1])
         );
  FA_X1 u4_sub_472_U2_2 ( .A(n3089), .B(u4_sub_472_n4), .CI(
        u4_sub_472_carry_2_), .CO(u4_sub_472_carry_3_), .S(u4_exp_fix_divb[2])
         );
  FA_X1 u4_sub_472_U2_3 ( .A(n3088), .B(u4_sub_472_n5), .CI(
        u4_sub_472_carry_3_), .CO(u4_sub_472_carry_4_), .S(u4_exp_fix_divb[3])
         );
  FA_X1 u4_sub_472_U2_4 ( .A(n3085), .B(u4_sub_472_n6), .CI(
        u4_sub_472_carry_4_), .CO(u4_sub_472_carry_5_), .S(u4_exp_fix_divb[4])
         );
  FA_X1 u4_sub_472_U2_5 ( .A(net85929), .B(u4_sub_472_n7), .CI(
        u4_sub_472_carry_5_), .CO(u4_sub_472_carry_6_), .S(u4_exp_fix_divb[5])
         );
  INV_X4 u4_sub_471_U11 ( .A(u4_fi_ldz_mi22[2]), .ZN(u4_sub_471_n6) );
  INV_X4 u4_sub_471_U10 ( .A(u4_fi_ldz_mi22[3]), .ZN(u4_sub_471_n5) );
  INV_X4 u4_sub_471_U9 ( .A(u4_fi_ldz_mi22[4]), .ZN(u4_sub_471_n4) );
  INV_X4 u4_sub_471_U8 ( .A(u4_fi_ldz_mi22[6]), .ZN(u4_sub_471_n3) );
  INV_X1 u4_sub_471_U7 ( .A(net94614), .ZN(u4_sub_471_n8) );
  INV_X4 u4_sub_471_U6 ( .A(net85905), .ZN(u4_sub_471_n2) );
  INV_X4 u4_sub_471_U5 ( .A(u4_sub_471_n8), .ZN(u4_sub_471_n1) );
  NAND2_X2 u4_sub_471_U4 ( .A1(u4_sub_471_n1), .A2(u4_sub_471_n2), .ZN(
        u4_sub_471_carry[1]) );
  XNOR2_X2 u4_sub_471_U3 ( .A(net85937), .B(u4_sub_471_carry[7]), .ZN(
        u4_exp_fix_diva[7]) );
  INV_X1 u4_sub_471_U2 ( .A(net33106), .ZN(u4_sub_471_n7) );
  XNOR2_X1 u4_sub_471_U1 ( .A(u4_sub_471_n8), .B(net85905), .ZN(
        u4_exp_fix_diva[0]) );
  FA_X1 u4_sub_471_U2_1 ( .A(n3091), .B(u4_sub_471_n7), .CI(
        u4_sub_471_carry[1]), .CO(u4_sub_471_carry[2]), .S(u4_exp_fix_diva[1])
         );
  FA_X1 u4_sub_471_U2_2 ( .A(n3089), .B(u4_sub_471_n6), .CI(
        u4_sub_471_carry[2]), .CO(u4_sub_471_carry[3]), .S(u4_exp_fix_diva[2])
         );
  FA_X1 u4_sub_471_U2_3 ( .A(n3088), .B(u4_sub_471_n5), .CI(
        u4_sub_471_carry[3]), .CO(u4_sub_471_carry[4]), .S(u4_exp_fix_diva[3])
         );
  FA_X1 u4_sub_471_U2_4 ( .A(n3085), .B(u4_sub_471_n4), .CI(
        u4_sub_471_carry[4]), .CO(u4_sub_471_carry[5]), .S(u4_exp_fix_diva[4])
         );
  FA_X1 u4_sub_471_U2_5 ( .A(net85929), .B(u4_sub_471_n3), .CI(
        u4_sub_471_carry[5]), .CO(u4_sub_471_carry[6]), .S(u4_exp_fix_diva[5])
         );
  FA_X1 u4_sub_471_U2_6 ( .A(net85933), .B(u4_sub_471_n3), .CI(
        u4_sub_471_carry[6]), .CO(u4_sub_471_carry[7]), .S(u4_exp_fix_diva[6])
         );
  AND2_X1 u4_sll_453_U509 ( .A1(u4_sll_453_ML_int_1__0_), .A2(
        u4_sll_453_net94113), .ZN(u4_sll_453_ML_int_2__0_) );
  AND2_X1 u4_sll_453_U508 ( .A1(u4_sll_453_ML_int_2__0_), .A2(
        u4_sll_453_net85273), .ZN(u4_sll_453_ML_int_3__0_) );
  AND2_X1 u4_sll_453_U507 ( .A1(u4_sll_453_ML_int_3__0_), .A2(
        u4_sll_453_net85301), .ZN(u4_sll_453_ML_int_4__0_) );
  AND2_X1 u4_sll_453_U506 ( .A1(u4_sll_453_ML_int_3__1_), .A2(
        u4_sll_453_net85303), .ZN(u4_sll_453_ML_int_4__1_) );
  AND2_X1 u4_sll_453_U505 ( .A1(u4_sll_453_ML_int_3__2_), .A2(
        u4_sll_453_net85321), .ZN(u4_sll_453_ML_int_4__2_) );
  AND2_X1 u4_sll_453_U504 ( .A1(u4_sll_453_ML_int_3__3_), .A2(
        u4_sll_453_net85321), .ZN(u4_sll_453_ML_int_4__3_) );
  NAND2_X1 u4_sll_453_U503 ( .A1(u4_sll_453_ML_int_4__0_), .A2(
        u4_sll_453_net85333), .ZN(u4_sll_453_n267) );
  INV_X1 u4_sll_453_U502 ( .A(u4_sll_453_n267), .ZN(u4_sll_453_ML_int_5__0_)
         );
  NAND2_X1 u4_sll_453_U501 ( .A1(u4_sll_453_ML_int_4__10_), .A2(
        u4_sll_453_net85333), .ZN(u4_sll_453_n266) );
  INV_X1 u4_sll_453_U500 ( .A(u4_sll_453_n266), .ZN(u4_sll_453_ML_int_5__10_)
         );
  NAND2_X1 u4_sll_453_U499 ( .A1(u4_sll_453_n179), .A2(u4_sll_453_net85333), 
        .ZN(u4_sll_453_n264) );
  INV_X1 u4_sll_453_U498 ( .A(u4_sll_453_n264), .ZN(u4_sll_453_ML_int_5__12_)
         );
  INV_X1 u4_sll_453_U497 ( .A(u4_sll_453_n262), .ZN(u4_sll_453_ML_int_5__14_)
         );
  NAND2_X1 u4_sll_453_U496 ( .A1(u4_sll_453_ML_int_4__1_), .A2(
        u4_sll_453_net85347), .ZN(u4_sll_453_n260) );
  INV_X1 u4_sll_453_U495 ( .A(u4_sll_453_n260), .ZN(u4_sll_453_ML_int_5__1_)
         );
  NAND2_X1 u4_sll_453_U494 ( .A1(u4_sll_453_ML_int_4__3_), .A2(
        u4_sll_453_net85347), .ZN(u4_sll_453_n259) );
  INV_X1 u4_sll_453_U493 ( .A(u4_sll_453_n259), .ZN(u4_sll_453_ML_int_5__3_)
         );
  NAND2_X1 u4_sll_453_U492 ( .A1(u4_sll_453_ML_int_4__4_), .A2(
        u4_sll_453_net85347), .ZN(u4_sll_453_n258) );
  INV_X1 u4_sll_453_U491 ( .A(u4_sll_453_n258), .ZN(u4_sll_453_ML_int_5__4_)
         );
  NAND2_X1 u4_sll_453_U490 ( .A1(u4_sll_453_ML_int_4__5_), .A2(
        u4_sll_453_net85347), .ZN(u4_sll_453_n257) );
  INV_X1 u4_sll_453_U489 ( .A(u4_sll_453_n257), .ZN(u4_sll_453_ML_int_5__5_)
         );
  NAND2_X1 u4_sll_453_U488 ( .A1(u4_sll_453_ML_int_4__6_), .A2(
        u4_sll_453_net85347), .ZN(u4_sll_453_n256) );
  INV_X1 u4_sll_453_U487 ( .A(u4_sll_453_n256), .ZN(u4_sll_453_ML_int_5__6_)
         );
  NAND2_X1 u4_sll_453_U486 ( .A1(u4_sll_453_ML_int_4__7_), .A2(
        u4_sll_453_net85347), .ZN(u4_sll_453_n255) );
  INV_X1 u4_sll_453_U485 ( .A(u4_sll_453_n255), .ZN(u4_sll_453_ML_int_5__7_)
         );
  NAND2_X1 u4_sll_453_U484 ( .A1(u4_sll_453_ML_int_4__8_), .A2(
        u4_sll_453_net94330), .ZN(u4_sll_453_n254) );
  INV_X1 u4_sll_453_U483 ( .A(u4_sll_453_n254), .ZN(u4_sll_453_ML_int_5__8_)
         );
  NAND2_X1 u4_sll_453_U482 ( .A1(u4_sll_453_ML_int_4__9_), .A2(
        u4_sll_453_net85347), .ZN(u4_sll_453_n253) );
  INV_X1 u4_sll_453_U481 ( .A(u4_sll_453_n253), .ZN(u4_sll_453_ML_int_5__9_)
         );
  NOR2_X1 u4_sll_453_U480 ( .A1(u4_sll_453_net85353), .A2(u4_sll_453_n267), 
        .ZN(u4_N1408) );
  NOR2_X1 u4_sll_453_U479 ( .A1(u4_sll_453_net85355), .A2(u4_sll_453_n266), 
        .ZN(u4_N1418) );
  NOR2_X1 u4_sll_453_U478 ( .A1(u4_sll_453_net85355), .A2(u4_sll_453_n265), 
        .ZN(u4_N1419) );
  NOR2_X1 u4_sll_453_U477 ( .A1(u4_sll_453_net85355), .A2(u4_sll_453_n264), 
        .ZN(u4_N1420) );
  NOR2_X1 u4_sll_453_U476 ( .A1(u4_sll_453_net85355), .A2(u4_sll_453_n263), 
        .ZN(u4_N1421) );
  NOR2_X1 u4_sll_453_U475 ( .A1(u4_sll_453_net85355), .A2(u4_sll_453_n262), 
        .ZN(u4_N1422) );
  NOR2_X1 u4_sll_453_U474 ( .A1(u4_sll_453_net85355), .A2(u4_sll_453_n260), 
        .ZN(u4_N1409) );
  NOR2_X1 u4_sll_453_U473 ( .A1(u4_sll_453_net85355), .A2(u4_sll_453_n259), 
        .ZN(u4_N1411) );
  NOR2_X1 u4_sll_453_U472 ( .A1(u4_sll_453_net85355), .A2(u4_sll_453_n258), 
        .ZN(u4_N1412) );
  NOR2_X1 u4_sll_453_U471 ( .A1(u4_sll_453_net85355), .A2(u4_sll_453_n257), 
        .ZN(u4_N1413) );
  NOR2_X1 u4_sll_453_U470 ( .A1(u4_sll_453_net85355), .A2(u4_sll_453_n256), 
        .ZN(u4_N1414) );
  NOR2_X1 u4_sll_453_U469 ( .A1(u4_sll_453_net85355), .A2(u4_sll_453_n255), 
        .ZN(u4_N1415) );
  NOR2_X1 u4_sll_453_U468 ( .A1(u4_sll_453_net85355), .A2(u4_sll_453_n254), 
        .ZN(u4_N1416) );
  NOR2_X1 u4_sll_453_U467 ( .A1(u4_sll_453_net85355), .A2(u4_sll_453_n253), 
        .ZN(u4_N1417) );
  AND2_X2 u4_sll_453_U466 ( .A1(u4_sll_453_ML_int_5__17_), .A2(
        u4_sll_453_net93876), .ZN(u4_N1425) );
  MUX2_X2 u4_sll_453_U465 ( .A(u4_sll_453_ML_int_2__18_), .B(
        u4_sll_453_ML_int_2__22_), .S(u4_sll_453_net85299), .Z(
        u4_sll_453_ML_int_3__22_) );
  MUX2_X2 u4_sll_453_U464 ( .A(u4_sll_453_ML_int_1__7_), .B(u4_sll_453_n237), 
        .S(u4_sll_453_net85265), .Z(u4_sll_453_ML_int_2__9_) );
  NAND2_X2 u4_sll_453_U463 ( .A1(u4_sll_453_n248), .A2(u4_sll_453_n249), .ZN(
        u4_sll_453_ML_int_1__20_) );
  NAND2_X1 u4_sll_453_U462 ( .A1(net17682), .A2(u4_sll_453_net94297), .ZN(
        u4_sll_453_n249) );
  NAND2_X2 u4_sll_453_U461 ( .A1(u4_sll_453_n246), .A2(u4_sll_453_n247), .ZN(
        u4_N1449) );
  NAND2_X1 u4_sll_453_U460 ( .A1(u4_sll_453_ML_int_5__9_), .A2(
        u4_sll_453_net85353), .ZN(u4_sll_453_n247) );
  NAND2_X2 u4_sll_453_U459 ( .A1(u4_sll_453_n244), .A2(u4_sll_453_n245), .ZN(
        u4_sll_453_ML_int_3__20_) );
  AND2_X2 u4_sll_453_U458 ( .A1(u4_sll_453_ML_int_5__20_), .A2(
        u4_sll_453_net93041), .ZN(u4_N1428) );
  INV_X4 u4_sll_453_U457 ( .A(u4_sll_453_net85285), .ZN(u4_sll_453_net85273)
         );
  MUX2_X2 u4_sll_453_U456 ( .A(u4_sll_453_ML_int_2__4_), .B(
        u4_sll_453_ML_int_2__8_), .S(u4_sll_453_net85273), .Z(
        u4_sll_453_ML_int_3__8_) );
  NAND2_X2 u4_sll_453_U455 ( .A1(u4_sll_453_n242), .A2(u4_sll_453_n243), .ZN(
        u4_N1450) );
  NAND2_X1 u4_sll_453_U454 ( .A1(u4_sll_453_ML_int_5__10_), .A2(
        u4_sll_453_net85353), .ZN(u4_sll_453_n243) );
  NAND2_X2 u4_sll_453_U453 ( .A1(u4_sll_453_n240), .A2(u4_sll_453_n241), .ZN(
        u4_sll_453_ML_int_1__12_) );
  NAND2_X1 u4_sll_453_U452 ( .A1(n5326), .A2(u4_sll_453_net92610), .ZN(
        u4_sll_453_n240) );
  MUX2_X2 u4_sll_453_U451 ( .A(u4_sll_453_ML_int_2__9_), .B(u4_sll_453_n238), 
        .S(u4_sll_453_n83), .Z(u4_sll_453_n239) );
  AND2_X2 u4_sll_453_U450 ( .A1(u4_sll_453_ML_int_5__23_), .A2(
        u4_sll_453_net93645), .ZN(u4_N1431) );
  AND2_X2 u4_sll_453_U449 ( .A1(u4_sll_453_ML_int_5__16_), .A2(
        u4_sll_453_net93728), .ZN(u4_N1424) );
  AND2_X2 u4_sll_453_U448 ( .A1(u4_sll_453_ML_int_5__24_), .A2(
        u4_sll_453_net93728), .ZN(u4_N1432) );
  MUX2_X2 u4_sll_453_U447 ( .A(u4_sll_453_ML_int_1__45_), .B(
        u4_sll_453_ML_int_1__47_), .S(u4_sll_453_net85265), .Z(
        u4_sll_453_ML_int_2__47_) );
  AND2_X2 u4_sll_453_U446 ( .A1(u4_sll_453_ML_int_5__29_), .A2(u4_sll_453_n109), .ZN(u4_N1437) );
  INV_X1 u4_sll_453_U445 ( .A(u4_sll_453_net85353), .ZN(u4_sll_453_net92613)
         );
  NAND2_X1 u4_sll_453_U444 ( .A1(u4_sll_453_ML_int_5__8_), .A2(
        u4_sll_453_net85353), .ZN(u4_sll_453_n236) );
  NAND2_X2 u4_sll_453_U443 ( .A1(u4_sll_453_n233), .A2(u4_sll_453_n234), .ZN(
        u4_sll_453_ML_int_1__30_) );
  NAND2_X1 u4_sll_453_U442 ( .A1(n3008), .A2(u4_sll_453_net92610), .ZN(
        u4_sll_453_n233) );
  NAND2_X2 u4_sll_453_U441 ( .A1(u4_sll_453_net92631), .A2(u4_sll_453_n232), 
        .ZN(u4_sll_453_ML_int_1__17_) );
  MUX2_X2 u4_sll_453_U440 ( .A(u4_sll_453_ML_int_1__15_), .B(
        u4_sll_453_ML_int_1__17_), .S(u4_sll_453_net85265), .Z(
        u4_sll_453_ML_int_2__17_) );
  INV_X1 u4_sll_453_U439 ( .A(u4_sll_453_net85355), .ZN(u4_sll_453_net93041)
         );
  NAND2_X2 u4_sll_453_U438 ( .A1(u4_sll_453_n230), .A2(u4_sll_453_n231), .ZN(
        u4_N1443) );
  NAND2_X1 u4_sll_453_U437 ( .A1(u4_sll_453_ML_int_5__3_), .A2(
        u4_sll_453_net85355), .ZN(u4_sll_453_n231) );
  NAND2_X2 u4_sll_453_U436 ( .A1(u4_sll_453_ML_int_5__35_), .A2(
        u4_sll_453_net93041), .ZN(u4_sll_453_n230) );
  INV_X1 u4_sll_453_U435 ( .A(u4_sll_453_net85341), .ZN(u4_sll_453_net93122)
         );
  NAND2_X2 u4_sll_453_U434 ( .A1(u4_sll_453_n228), .A2(u4_sll_453_n229), .ZN(
        u4_sll_453_ML_int_5__36_) );
  NAND2_X1 u4_sll_453_U433 ( .A1(u4_sll_453_ML_int_4__20_), .A2(
        u4_sll_453_net85341), .ZN(u4_sll_453_n229) );
  NAND2_X2 u4_sll_453_U432 ( .A1(u4_sll_453_ML_int_4__36_), .A2(
        u4_sll_453_net93122), .ZN(u4_sll_453_n228) );
  NAND2_X2 u4_sll_453_U431 ( .A1(u4_sll_453_n227), .A2(u4_sll_453_n226), .ZN(
        u4_sll_453_ML_int_5__47_) );
  NAND2_X2 u4_sll_453_U430 ( .A1(u4_sll_453_ML_int_4__47_), .A2(
        u4_sll_453_net85333), .ZN(u4_sll_453_n227) );
  INV_X1 u4_sll_453_U429 ( .A(u4_sll_453_net85341), .ZN(u4_sll_453_net93219)
         );
  NAND2_X2 u4_sll_453_U428 ( .A1(u4_sll_453_n224), .A2(u4_sll_453_n225), .ZN(
        u4_sll_453_ML_int_5__39_) );
  NAND2_X1 u4_sll_453_U427 ( .A1(u4_sll_453_ML_int_4__23_), .A2(
        u4_sll_453_net85341), .ZN(u4_sll_453_n225) );
  NAND2_X2 u4_sll_453_U426 ( .A1(u4_sll_453_ML_int_4__39_), .A2(
        u4_sll_453_net93219), .ZN(u4_sll_453_n224) );
  NAND2_X2 u4_sll_453_U425 ( .A1(u4_sll_453_n223), .A2(u4_sll_453_net93284), 
        .ZN(u4_sll_453_ML_int_3__19_) );
  NAND2_X1 u4_sll_453_U424 ( .A1(u4_sll_453_ML_int_2__15_), .A2(
        u4_sll_453_net85287), .ZN(u4_sll_453_n223) );
  INV_X2 u4_sll_453_U423 ( .A(u4_sll_453_net85315), .ZN(u4_sll_453_net93359)
         );
  NAND2_X1 u4_sll_453_U422 ( .A1(u4_sll_453_ML_int_3__9_), .A2(
        u4_sll_453_net85315), .ZN(u4_sll_453_n222) );
  NAND2_X1 u4_sll_453_U421 ( .A1(u4_sll_453_ML_int_3__17_), .A2(
        u4_sll_453_net93359), .ZN(u4_sll_453_n221) );
  AND2_X2 u4_sll_453_U420 ( .A1(u4_sll_453_ML_int_5__27_), .A2(
        u4_sll_453_net85365), .ZN(u4_N1435) );
  NAND2_X2 u4_sll_453_U419 ( .A1(u4_sll_453_net93630), .A2(u4_sll_453_net93631), .ZN(u4_sll_453_n237) );
  INV_X1 u4_sll_453_U418 ( .A(u4_sll_453_net85353), .ZN(u4_sll_453_net93645)
         );
  NAND2_X1 u4_sll_453_U417 ( .A1(u4_sll_453_ML_int_5__5_), .A2(
        u4_sll_453_net85353), .ZN(u4_sll_453_n220) );
  NAND2_X2 u4_sll_453_U416 ( .A1(u4_sll_453_n217), .A2(u4_sll_453_n218), .ZN(
        u4_sll_453_ML_int_3__29_) );
  NAND2_X1 u4_sll_453_U415 ( .A1(u4_sll_453_ML_int_2__25_), .A2(
        u4_sll_453_net85289), .ZN(u4_sll_453_n218) );
  MUX2_X2 u4_sll_453_U414 ( .A(u4_sll_453_ML_int_1__19_), .B(
        u4_sll_453_ML_int_1__21_), .S(u4_sll_453_net93710), .Z(
        u4_sll_453_ML_int_2__21_) );
  INV_X1 u4_sll_453_U413 ( .A(u4_sll_453_net85353), .ZN(u4_sll_453_net93728)
         );
  NAND2_X2 u4_sll_453_U412 ( .A1(u4_sll_453_n215), .A2(u4_sll_453_n216), .ZN(
        u4_N1446) );
  NAND2_X1 u4_sll_453_U411 ( .A1(u4_sll_453_ML_int_5__6_), .A2(
        u4_sll_453_net85353), .ZN(u4_sll_453_n216) );
  NAND2_X2 u4_sll_453_U410 ( .A1(u4_sll_453_n213), .A2(u4_sll_453_n214), .ZN(
        u4_sll_453_ML_int_3__14_) );
  NAND2_X1 u4_sll_453_U409 ( .A1(u4_sll_453_ML_int_2__10_), .A2(
        u4_sll_453_net85287), .ZN(u4_sll_453_n214) );
  NAND2_X1 u4_sll_453_U408 ( .A1(u4_sll_453_ML_int_2__14_), .A2(
        u4_sll_453_net93725), .ZN(u4_sll_453_n213) );
  AND2_X2 u4_sll_453_U407 ( .A1(u4_sll_453_ML_int_5__31_), .A2(
        u4_sll_453_net93876), .ZN(u4_N1439) );
  INV_X1 u4_sll_453_U406 ( .A(u4_sll_453_net85343), .ZN(u4_sll_453_net93857)
         );
  NAND2_X2 u4_sll_453_U405 ( .A1(u4_sll_453_n211), .A2(u4_sll_453_n212), .ZN(
        u4_sll_453_ML_int_5__43_) );
  NAND2_X2 u4_sll_453_U404 ( .A1(u4_sll_453_ML_int_4__43_), .A2(
        u4_sll_453_net93857), .ZN(u4_sll_453_n211) );
  NAND2_X4 u4_sll_453_U403 ( .A1(u4_sll_453_n209), .A2(u4_sll_453_n210), .ZN(
        u4_N1452) );
  NAND2_X2 u4_sll_453_U402 ( .A1(u4_sll_453_ML_int_5__12_), .A2(
        u4_sll_453_net85353), .ZN(u4_sll_453_n210) );
  NAND2_X4 u4_sll_453_U401 ( .A1(u4_sll_453_ML_int_5__44_), .A2(
        u4_sll_453_net93876), .ZN(u4_sll_453_n209) );
  NAND2_X2 u4_sll_453_U400 ( .A1(u4_sll_453_n207), .A2(u4_sll_453_n208), .ZN(
        u4_sll_453_ML_int_3__28_) );
  CLKBUF_X2 u4_sll_453_U399 ( .A(u4_sll_453_ML_int_3__15_), .Z(u4_sll_453_n252) );
  NAND2_X2 u4_sll_453_U398 ( .A1(u4_sll_453_n205), .A2(u4_sll_453_n206), .ZN(
        u4_sll_453_ML_int_3__15_) );
  NAND2_X2 u4_sll_453_U397 ( .A1(u4_sll_453_ML_int_2__15_), .A2(
        u4_sll_453_net93725), .ZN(u4_sll_453_n205) );
  NAND2_X2 u4_sll_453_U396 ( .A1(u4_sll_453_n203), .A2(u4_sll_453_n204), .ZN(
        u4_sll_453_ML_int_5__33_) );
  NAND2_X1 u4_sll_453_U395 ( .A1(u4_sll_453_ML_int_4__17_), .A2(
        u4_sll_453_net85341), .ZN(u4_sll_453_n204) );
  NAND2_X2 u4_sll_453_U394 ( .A1(u4_sll_453_ML_int_4__33_), .A2(
        u4_sll_453_n163), .ZN(u4_sll_453_n203) );
  NAND2_X1 u4_sll_453_U393 ( .A1(net17692), .A2(u4_sll_453_net94297), .ZN(
        u4_sll_453_n202) );
  NAND2_X1 u4_sll_453_U392 ( .A1(net17654), .A2(u4_sll_453_n61), .ZN(
        u4_sll_453_n201) );
  NAND2_X2 u4_sll_453_U391 ( .A1(u4_sll_453_net93929), .A2(u4_sll_453_net93930), .ZN(u4_sll_453_ML_int_2__8_) );
  NAND2_X2 u4_sll_453_U390 ( .A1(u4_sll_453_n199), .A2(u4_sll_453_n200), .ZN(
        u4_sll_453_ML_int_2__22_) );
  NAND2_X1 u4_sll_453_U389 ( .A1(u4_sll_453_ML_int_1__20_), .A2(
        u4_sll_453_net85259), .ZN(u4_sll_453_n200) );
  NAND2_X2 u4_sll_453_U388 ( .A1(u4_sll_453_ML_int_1__22_), .A2(
        u4_sll_453_net94113), .ZN(u4_sll_453_n199) );
  INV_X1 u4_sll_453_U387 ( .A(u4_sll_453_net85343), .ZN(u4_sll_453_net93991)
         );
  NAND2_X2 u4_sll_453_U386 ( .A1(u4_sll_453_n197), .A2(u4_sll_453_n198), .ZN(
        u4_sll_453_ML_int_5__45_) );
  NAND2_X2 u4_sll_453_U385 ( .A1(u4_sll_453_ML_int_4__45_), .A2(
        u4_sll_453_net93991), .ZN(u4_sll_453_n197) );
  INV_X4 u4_sll_453_U384 ( .A(u4_sll_453_n194), .ZN(u4_sll_453_ML_int_3__32_)
         );
  MUX2_X2 u4_sll_453_U383 ( .A(u4_sll_453_n196), .B(u4_sll_453_n195), .S(
        u4_sll_453_net85289), .Z(u4_sll_453_n194) );
  AND2_X2 u4_sll_453_U382 ( .A1(u4_sll_453_ML_int_2__2_), .A2(u4_sll_453_n90), 
        .ZN(u4_sll_453_ML_int_3__2_) );
  NAND2_X2 u4_sll_453_U381 ( .A1(u4_sll_453_n193), .A2(u4_sll_453_net94050), 
        .ZN(u4_sll_453_ML_int_2__5_) );
  NAND2_X2 u4_sll_453_U380 ( .A1(u4_sll_453_ML_int_1__3_), .A2(
        u4_sll_453_net85263), .ZN(u4_sll_453_n193) );
  NAND2_X2 u4_sll_453_U379 ( .A1(u4_sll_453_n191), .A2(u4_sll_453_n192), .ZN(
        u4_sll_453_ML_int_3__11_) );
  NAND2_X1 u4_sll_453_U378 ( .A1(u4_sll_453_ML_int_2__7_), .A2(
        u4_sll_453_net85287), .ZN(u4_sll_453_n192) );
  NAND2_X2 u4_sll_453_U377 ( .A1(u4_sll_453_ML_int_2__11_), .A2(
        u4_sll_453_net93725), .ZN(u4_sll_453_n191) );
  NAND2_X2 u4_sll_453_U376 ( .A1(u4_sll_453_n189), .A2(u4_sll_453_n190), .ZN(
        u4_sll_453_ML_int_2__7_) );
  NAND2_X1 u4_sll_453_U375 ( .A1(u4_sll_453_ML_int_1__5_), .A2(
        u4_sll_453_net85257), .ZN(u4_sll_453_n190) );
  MUX2_X2 u4_sll_453_U374 ( .A(u4_sll_453_ML_int_2__20_), .B(
        u4_sll_453_ML_int_2__24_), .S(u4_sll_453_net85299), .Z(
        u4_sll_453_ML_int_3__24_) );
  NAND2_X2 u4_sll_453_U373 ( .A1(u4_sll_453_n221), .A2(u4_sll_453_n222), .ZN(
        u4_sll_453_ML_int_4__17_) );
  NAND2_X2 u4_sll_453_U372 ( .A1(u4_sll_453_n187), .A2(u4_sll_453_n188), .ZN(
        u4_sll_453_ML_int_5__32_) );
  NAND2_X1 u4_sll_453_U371 ( .A1(u4_sll_453_ML_int_4__16_), .A2(
        u4_sll_453_net85341), .ZN(u4_sll_453_n188) );
  NAND2_X2 u4_sll_453_U370 ( .A1(u4_sll_453_ML_int_4__32_), .A2(
        u4_sll_453_net94330), .ZN(u4_sll_453_n187) );
  AND2_X2 u4_sll_453_U369 ( .A1(u4_sll_453_ML_int_5__21_), .A2(
        u4_sll_453_net93876), .ZN(u4_N1429) );
  AND2_X2 u4_sll_453_U368 ( .A1(u4_sll_453_ML_int_5__26_), .A2(u4_sll_453_n109), .ZN(u4_N1434) );
  AND2_X2 u4_sll_453_U367 ( .A1(u4_sll_453_ML_int_2__3_), .A2(u4_sll_453_n90), 
        .ZN(u4_sll_453_ML_int_3__3_) );
  AND2_X2 u4_sll_453_U366 ( .A1(u4_sll_453_ML_int_1__1_), .A2(
        u4_sll_453_net94113), .ZN(u4_sll_453_ML_int_2__1_) );
  AND2_X2 u4_sll_453_U365 ( .A1(u4_sll_453_ML_int_3__7_), .A2(
        u4_sll_453_net85321), .ZN(u4_sll_453_ML_int_4__7_) );
  INV_X1 u4_sll_453_U364 ( .A(u4_sll_453_net85315), .ZN(u4_sll_453_net94228)
         );
  NAND2_X2 u4_sll_453_U363 ( .A1(u4_sll_453_n185), .A2(u4_sll_453_n186), .ZN(
        u4_sll_453_ML_int_4__24_) );
  AND2_X2 u4_sll_453_U362 ( .A1(u4_sll_453_ML_int_3__5_), .A2(
        u4_sll_453_net85321), .ZN(u4_sll_453_ML_int_4__5_) );
  NAND2_X2 u4_sll_453_U361 ( .A1(u4_sll_453_n183), .A2(u4_sll_453_n184), .ZN(
        u4_sll_453_ML_int_5__21_) );
  NAND2_X1 u4_sll_453_U360 ( .A1(u4_sll_453_ML_int_4__5_), .A2(
        u4_sll_453_net85339), .ZN(u4_sll_453_n184) );
  NAND2_X1 u4_sll_453_U359 ( .A1(u4_sll_453_ML_int_4__21_), .A2(
        u4_sll_453_net94330), .ZN(u4_sll_453_n183) );
  AND2_X4 u4_sll_453_U358 ( .A1(u4_sll_453_ML_int_5__18_), .A2(u4_sll_453_n109), .ZN(u4_N1426) );
  NAND2_X2 u4_sll_453_U357 ( .A1(u4_sll_453_n181), .A2(u4_sll_453_n182), .ZN(
        u4_sll_453_ML_int_5__31_) );
  INV_X4 u4_sll_453_U356 ( .A(u4_sll_453_ML_int_2__32_), .ZN(u4_sll_453_n196)
         );
  INV_X4 u4_sll_453_U355 ( .A(u4_sll_453_net85237), .ZN(u4_sll_453_net85229)
         );
  MUX2_X2 u4_sll_453_U354 ( .A(u4_sll_453_n238), .B(u4_sll_453_ML_int_2__17_), 
        .S(u4_sll_453_net85275), .Z(u4_sll_453_ML_int_3__17_) );
  INV_X4 u4_sll_453_U353 ( .A(u4_sll_453_n261), .ZN(u4_sll_453_ML_int_5__15_)
         );
  INV_X1 u4_sll_453_U352 ( .A(u4_sll_453_ML_int_5__15_), .ZN(u4_sll_453_n180)
         );
  AND2_X2 u4_sll_453_U351 ( .A1(u4_sll_453_ML_int_5__30_), .A2(u4_sll_453_n109), .ZN(u4_N1438) );
  MUX2_X2 u4_sll_453_U350 ( .A(u4_sll_453_ML_int_3__30_), .B(u4_sll_453_n177), 
        .S(u4_sll_453_net85315), .Z(u4_sll_453_n178) );
  INV_X2 u4_sll_453_U349 ( .A(u4_sll_453_ML_int_2__28_), .ZN(u4_sll_453_n195)
         );
  NAND2_X2 u4_sll_453_U348 ( .A1(u4_sll_453_ML_int_2__28_), .A2(
        u4_sll_453_net93725), .ZN(u4_sll_453_n207) );
  AND2_X2 u4_sll_453_U347 ( .A1(u4_sll_453_ML_int_5__25_), .A2(
        u4_sll_453_net92613), .ZN(u4_N1433) );
  MUX2_X2 u4_sll_453_U346 ( .A(u4_sll_453_ML_int_2__18_), .B(
        u4_sll_453_ML_int_2__22_), .S(u4_sll_453_net85299), .Z(u4_sll_453_n177) );
  INV_X32 u4_sll_453_U345 ( .A(u4_sll_453_net85265), .ZN(u4_sll_453_net85259)
         );
  MUX2_X2 u4_sll_453_U344 ( .A(u4_sll_453_ML_int_1__18_), .B(u4_sll_453_n1), 
        .S(u4_sll_453_net85259), .Z(u4_sll_453_n175) );
  NOR2_X1 u4_sll_453_U343 ( .A1(u4_sll_453_net85355), .A2(u4_sll_453_net12807), 
        .ZN(u4_N1410) );
  NAND2_X1 u4_sll_453_U342 ( .A1(u4_sll_453_ML_int_4__2_), .A2(
        u4_sll_453_net85347), .ZN(u4_sll_453_net12807) );
  INV_X1 u4_sll_453_U341 ( .A(u4_sll_453_net12807), .ZN(
        u4_sll_453_ML_int_5__2_) );
  INV_X32 u4_sll_453_U340 ( .A(u4_sll_453_net85365), .ZN(u4_sll_453_net85355)
         );
  NAND2_X2 u4_sll_453_U339 ( .A1(u4_sll_453_ML_int_1__6_), .A2(
        u4_sll_453_net85263), .ZN(u4_sll_453_net93929) );
  NAND2_X1 u4_sll_453_U338 ( .A1(u4_sll_453_ML_int_1__5_), .A2(
        u4_sll_453_net85267), .ZN(u4_sll_453_net94050) );
  AND2_X1 u4_sll_453_U337 ( .A1(u4_sll_453_ML_int_2__1_), .A2(
        u4_sll_453_net85275), .ZN(u4_sll_453_ML_int_3__1_) );
  NAND2_X1 u4_sll_453_U336 ( .A1(u4_sll_453_ML_int_2__19_), .A2(
        u4_sll_453_net85275), .ZN(u4_sll_453_net93284) );
  INV_X8 u4_sll_453_U335 ( .A(u4_sll_453_net85237), .ZN(u4_sll_453_net85231)
         );
  NAND2_X1 u4_sll_453_U334 ( .A1(net17657), .A2(u4_sll_453_net92610), .ZN(
        u4_sll_453_net92631) );
  NAND2_X1 u4_sll_453_U333 ( .A1(net17690), .A2(u4_sll_453_net92610), .ZN(
        u4_sll_453_n173) );
  NAND2_X1 u4_sll_453_U332 ( .A1(n5323), .A2(u4_sll_453_net86374), .ZN(
        u4_sll_453_n174) );
  NAND2_X1 u4_sll_453_U331 ( .A1(u4_sll_453_ML_int_1__8_), .A2(
        u4_sll_453_net85265), .ZN(u4_sll_453_net93930) );
  NAND2_X2 u4_sll_453_U330 ( .A1(u4_sll_453_n173), .A2(u4_sll_453_n174), .ZN(
        u4_sll_453_ML_int_1__8_) );
  INV_X32 u4_sll_453_U329 ( .A(u4_sll_453_net85269), .ZN(u4_sll_453_net85265)
         );
  INV_X32 u4_sll_453_U328 ( .A(u4_sll_453_net85265), .ZN(u4_sll_453_net85261)
         );
  MUX2_X2 u4_sll_453_U327 ( .A(u4_sll_453_ML_int_1__28_), .B(
        u4_sll_453_ML_int_1__30_), .S(u4_sll_453_net85265), .Z(
        u4_sll_453_ML_int_2__30_) );
  INV_X32 u4_sll_453_U326 ( .A(u4_sll_453_net85319), .ZN(u4_sll_453_net85315)
         );
  INV_X32 u4_sll_453_U325 ( .A(u4_sll_453_net85319), .ZN(u4_sll_453_net85313)
         );
  MUX2_X2 u4_sll_453_U324 ( .A(u4_sll_453_ML_int_3__21_), .B(
        u4_sll_453_ML_int_3__29_), .S(u4_sll_453_net85319), .Z(
        u4_sll_453_ML_int_4__29_) );
  NAND2_X1 u4_sll_453_U323 ( .A1(n2981), .A2(u4_sll_453_n104), .ZN(
        u4_sll_453_net93630) );
  INV_X16 u4_sll_453_U322 ( .A(u4_shift_left[0]), .ZN(u4_sll_453_net85237) );
  MUX2_X2 u4_sll_453_U321 ( .A(n5324), .B(n2981), .S(u4_sll_453_net85229), .Z(
        u4_sll_453_n172) );
  INV_X16 u4_sll_453_U320 ( .A(u4_sll_453_net85351), .ZN(u4_sll_453_net85339)
         );
  INV_X4 u4_sll_453_U319 ( .A(u4_sll_453_net85257), .ZN(u4_sll_453_net94113)
         );
  INV_X1 u4_sll_453_U318 ( .A(u4_sll_453_net85313), .ZN(u4_sll_453_net85301)
         );
  INV_X1 u4_sll_453_U317 ( .A(u4_sll_453_net85313), .ZN(u4_sll_453_net85303)
         );
  INV_X1 u4_sll_453_U316 ( .A(u4_sll_453_net85313), .ZN(u4_sll_453_net91550)
         );
  INV_X8 u4_sll_453_U315 ( .A(u4_shift_left[3]), .ZN(u4_sll_453_net85321) );
  INV_X16 u4_sll_453_U314 ( .A(u4_sll_453_net85299), .ZN(u4_sll_453_net85285)
         );
  INV_X16 u4_sll_453_U313 ( .A(u4_shift_left[3]), .ZN(u4_sll_453_net85319) );
  INV_X32 u4_sll_453_U312 ( .A(u4_sll_453_net85237), .ZN(u4_sll_453_net86373)
         );
  MUX2_X2 u4_sll_453_U311 ( .A(u4_sll_453_ML_int_1__13_), .B(
        u4_sll_453_ML_int_1__15_), .S(u4_sll_453_n171), .Z(
        u4_sll_453_ML_int_2__15_) );
  INV_X2 u4_sll_453_U310 ( .A(u4_sll_453_n263), .ZN(u4_sll_453_ML_int_5__13_)
         );
  NAND2_X2 u4_sll_453_U309 ( .A1(u4_sll_453_n169), .A2(u4_sll_453_n170), .ZN(
        u4_sll_453_ML_int_3__25_) );
  NAND2_X2 u4_sll_453_U308 ( .A1(u4_sll_453_ML_int_2__21_), .A2(
        u4_sll_453_net85287), .ZN(u4_sll_453_n170) );
  NAND2_X2 u4_sll_453_U307 ( .A1(u4_sll_453_ML_int_2__25_), .A2(u4_sll_453_n90), .ZN(u4_sll_453_n169) );
  INV_X1 u4_sll_453_U306 ( .A(u4_sll_453_net85315), .ZN(u4_sll_453_n166) );
  NAND2_X2 u4_sll_453_U305 ( .A1(u4_sll_453_n167), .A2(u4_sll_453_n168), .ZN(
        u4_sll_453_ML_int_4__25_) );
  NAND2_X1 u4_sll_453_U304 ( .A1(u4_sll_453_ML_int_3__17_), .A2(
        u4_sll_453_net85315), .ZN(u4_sll_453_n168) );
  NAND2_X2 u4_sll_453_U303 ( .A1(u4_sll_453_ML_int_3__25_), .A2(
        u4_sll_453_n166), .ZN(u4_sll_453_n167) );
  NAND2_X2 u4_sll_453_U302 ( .A1(u4_sll_453_n164), .A2(u4_sll_453_n165), .ZN(
        u4_sll_453_ML_int_5__41_) );
  NAND2_X2 u4_sll_453_U301 ( .A1(u4_sll_453_ML_int_4__25_), .A2(
        u4_sll_453_net85343), .ZN(u4_sll_453_n165) );
  NAND2_X2 u4_sll_453_U300 ( .A1(u4_sll_453_ML_int_4__41_), .A2(
        u4_sll_453_n163), .ZN(u4_sll_453_n164) );
  INV_X1 u4_sll_453_U299 ( .A(u4_sll_453_net94297), .ZN(u4_sll_453_n160) );
  NAND2_X2 u4_sll_453_U298 ( .A1(u4_sll_453_n161), .A2(u4_sll_453_n162), .ZN(
        u4_sll_453_ML_int_1__19_) );
  NAND2_X1 u4_sll_453_U297 ( .A1(net17683), .A2(u4_sll_453_net86374), .ZN(
        u4_sll_453_n162) );
  NAND2_X1 u4_sll_453_U296 ( .A1(net17682), .A2(u4_sll_453_n160), .ZN(
        u4_sll_453_n161) );
  NAND2_X2 u4_sll_453_U295 ( .A1(u4_sll_453_n158), .A2(u4_sll_453_n159), .ZN(
        u4_sll_453_ML_int_3__23_) );
  NAND2_X1 u4_sll_453_U294 ( .A1(u4_sll_453_ML_int_2__19_), .A2(
        u4_sll_453_net85287), .ZN(u4_sll_453_n159) );
  NAND2_X2 u4_sll_453_U293 ( .A1(u4_sll_453_ML_int_2__11_), .A2(
        u4_sll_453_net85287), .ZN(u4_sll_453_n206) );
  NAND2_X2 u4_sll_453_U292 ( .A1(u4_sll_453_ML_int_4__31_), .A2(
        u4_sll_453_n163), .ZN(u4_sll_453_n181) );
  NAND2_X2 u4_sll_453_U291 ( .A1(u4_sll_453_n156), .A2(u4_sll_453_n157), .ZN(
        u4_sll_453_ML_int_3__31_) );
  NAND2_X1 u4_sll_453_U290 ( .A1(u4_sll_453_ML_int_2__27_), .A2(
        u4_sll_453_net85289), .ZN(u4_sll_453_n157) );
  INV_X1 u4_sll_453_U289 ( .A(u4_sll_453_net85315), .ZN(u4_sll_453_n153) );
  NAND2_X4 u4_sll_453_U288 ( .A1(u4_sll_453_n154), .A2(u4_sll_453_n155), .ZN(
        u4_sll_453_ML_int_4__31_) );
  NAND2_X1 u4_sll_453_U287 ( .A1(u4_sll_453_ML_int_3__23_), .A2(
        u4_sll_453_net85315), .ZN(u4_sll_453_n155) );
  NAND2_X4 u4_sll_453_U286 ( .A1(u4_sll_453_ML_int_3__31_), .A2(
        u4_sll_453_n153), .ZN(u4_sll_453_n154) );
  MUX2_X1 u4_sll_453_U285 ( .A(u4_sll_453_ML_int_3__12_), .B(
        u4_sll_453_ML_int_3__4_), .S(u4_sll_453_net85313), .Z(u4_sll_453_n179)
         );
  AND2_X2 u4_sll_453_U284 ( .A1(u4_sll_453_ML_int_3__4_), .A2(
        u4_sll_453_net85321), .ZN(u4_sll_453_ML_int_4__4_) );
  INV_X1 u4_sll_453_U283 ( .A(u4_sll_453_net85275), .ZN(u4_sll_453_n150) );
  NAND2_X2 u4_sll_453_U282 ( .A1(u4_sll_453_n151), .A2(u4_sll_453_n152), .ZN(
        u4_sll_453_ML_int_3__10_) );
  NAND2_X1 u4_sll_453_U281 ( .A1(u4_sll_453_ML_int_2__10_), .A2(
        u4_sll_453_net85275), .ZN(u4_sll_453_n152) );
  NAND2_X2 u4_sll_453_U280 ( .A1(u4_sll_453_ML_int_2__6_), .A2(u4_sll_453_n150), .ZN(u4_sll_453_n151) );
  NAND2_X2 u4_sll_453_U279 ( .A1(u4_sll_453_n172), .A2(u4_sll_453_net85265), 
        .ZN(u4_sll_453_n149) );
  NAND2_X4 u4_sll_453_U278 ( .A1(u4_sll_453_ML_int_1__8_), .A2(
        u4_sll_453_net85263), .ZN(u4_sll_453_n148) );
  NAND2_X2 u4_sll_453_U277 ( .A1(u4_sll_453_n145), .A2(u4_sll_453_n146), .ZN(
        u4_sll_453_n238) );
  NAND2_X1 u4_sll_453_U276 ( .A1(u4_sll_453_ML_int_1__11_), .A2(
        u4_sll_453_net85259), .ZN(u4_sll_453_n146) );
  NAND2_X1 u4_sll_453_U275 ( .A1(u4_sll_453_ML_int_1__13_), .A2(
        u4_sll_453_n137), .ZN(u4_sll_453_n145) );
  INV_X4 u4_sll_453_U274 ( .A(u4_sll_453_net85351), .ZN(u4_sll_453_n142) );
  NAND2_X2 u4_sll_453_U273 ( .A1(u4_sll_453_n144), .A2(u4_sll_453_n143), .ZN(
        u4_sll_453_ML_int_5__34_) );
  NAND2_X2 u4_sll_453_U272 ( .A1(u4_sll_453_ML_int_4__34_), .A2(
        u4_sll_453_net85351), .ZN(u4_sll_453_n144) );
  NAND2_X2 u4_sll_453_U271 ( .A1(u4_sll_453_ML_int_4__18_), .A2(
        u4_sll_453_n142), .ZN(u4_sll_453_n143) );
  NAND2_X2 u4_sll_453_U270 ( .A1(u4_sll_453_ML_int_2__23_), .A2(
        u4_sll_453_net93725), .ZN(u4_sll_453_n158) );
  NAND2_X2 u4_sll_453_U269 ( .A1(u4_sll_453_n140), .A2(u4_sll_453_n141), .ZN(
        u4_sll_453_ML_int_1__21_) );
  NAND2_X1 u4_sll_453_U268 ( .A1(net17659), .A2(u4_sll_453_net85231), .ZN(
        u4_sll_453_n141) );
  NAND2_X1 u4_sll_453_U267 ( .A1(fract_denorm[21]), .A2(u4_sll_453_n104), .ZN(
        u4_sll_453_n140) );
  NAND2_X2 u4_sll_453_U266 ( .A1(u4_sll_453_ML_int_1__21_), .A2(
        u4_sll_453_net85259), .ZN(u4_sll_453_n139) );
  NAND2_X2 u4_sll_453_U265 ( .A1(u4_sll_453_ML_int_1__23_), .A2(
        u4_sll_453_n137), .ZN(u4_sll_453_n138) );
  NAND2_X2 u4_sll_453_U264 ( .A1(u4_sll_453_ML_int_4__15_), .A2(
        u4_sll_453_net85341), .ZN(u4_sll_453_n182) );
  NAND2_X2 u4_sll_453_U263 ( .A1(u4_sll_453_ML_int_4__15_), .A2(
        u4_sll_453_net85347), .ZN(u4_sll_453_n261) );
  INV_X1 u4_sll_453_U262 ( .A(u4_sll_453_net85315), .ZN(u4_sll_453_net95318)
         );
  NAND2_X4 u4_sll_453_U261 ( .A1(u4_sll_453_n135), .A2(u4_sll_453_n136), .ZN(
        u4_sll_453_ML_int_4__15_) );
  NAND2_X2 u4_sll_453_U260 ( .A1(u4_sll_453_n252), .A2(u4_sll_453_net95318), 
        .ZN(u4_sll_453_n136) );
  NAND2_X2 u4_sll_453_U259 ( .A1(u4_sll_453_ML_int_3__7_), .A2(u4_sll_453_n134), .ZN(u4_sll_453_n135) );
  NAND2_X2 u4_sll_453_U258 ( .A1(u4_sll_453_ML_int_5__15_), .A2(
        u4_sll_453_net85353), .ZN(u4_sll_453_n133) );
  NAND2_X4 u4_sll_453_U257 ( .A1(u4_sll_453_ML_int_5__47_), .A2(
        u4_sll_453_n109), .ZN(u4_sll_453_n132) );
  NAND2_X4 u4_sll_453_U256 ( .A1(u4_sll_453_n219), .A2(u4_sll_453_n220), .ZN(
        u4_N1445) );
  INV_X1 u4_sll_453_U255 ( .A(u4_sll_453_n112), .ZN(u4_sll_453_n129) );
  NAND2_X2 u4_sll_453_U254 ( .A1(u4_sll_453_n130), .A2(u4_sll_453_n131), .ZN(
        u4_sll_453_ML_int_3__13_) );
  NAND2_X1 u4_sll_453_U253 ( .A1(u4_sll_453_ML_int_2__13_), .A2(
        u4_sll_453_net93725), .ZN(u4_sll_453_n131) );
  NAND2_X1 u4_sll_453_U252 ( .A1(u4_sll_453_ML_int_2__9_), .A2(u4_sll_453_n129), .ZN(u4_sll_453_n130) );
  NAND2_X2 u4_sll_453_U251 ( .A1(u4_sll_453_ML_int_2__20_), .A2(
        u4_sll_453_n112), .ZN(u4_sll_453_n244) );
  AND2_X2 u4_sll_453_U250 ( .A1(u4_sll_453_ML_int_3__6_), .A2(
        u4_sll_453_net85321), .ZN(u4_sll_453_ML_int_4__6_) );
  AND2_X2 u4_sll_453_U249 ( .A1(net17652), .A2(u4_sll_453_net92610), .ZN(
        u4_sll_453_ML_int_1__0_) );
  NAND2_X4 u4_sll_453_U248 ( .A1(u4_sll_453_ML_int_5__46_), .A2(
        u4_sll_453_n109), .ZN(u4_sll_453_n250) );
  NAND2_X2 u4_sll_453_U247 ( .A1(u4_sll_453_ML_int_5__14_), .A2(
        u4_sll_453_net85353), .ZN(u4_sll_453_n251) );
  NAND2_X4 u4_sll_453_U246 ( .A1(u4_sll_453_n250), .A2(u4_sll_453_n251), .ZN(
        u4_N1454) );
  NAND2_X2 u4_sll_453_U245 ( .A1(u4_sll_453_n127), .A2(u4_sll_453_n128), .ZN(
        u4_sll_453_ML_int_5__30_) );
  NAND2_X2 u4_sll_453_U244 ( .A1(u4_sll_453_ML_int_4__14_), .A2(
        u4_sll_453_net85341), .ZN(u4_sll_453_n128) );
  NAND2_X2 u4_sll_453_U243 ( .A1(u4_sll_453_n178), .A2(u4_sll_453_net94330), 
        .ZN(u4_sll_453_n127) );
  NAND2_X4 u4_sll_453_U242 ( .A1(u4_sll_453_n235), .A2(u4_sll_453_n236), .ZN(
        u4_N1448) );
  NAND2_X4 u4_sll_453_U241 ( .A1(u4_sll_453_ML_int_5__40_), .A2(
        u4_sll_453_net92613), .ZN(u4_sll_453_n235) );
  NAND2_X1 u4_sll_453_U240 ( .A1(u4_sll_453_ML_int_5__42_), .A2(
        u4_sll_453_n109), .ZN(u4_sll_453_n242) );
  INV_X32 u4_sll_453_U239 ( .A(u4_sll_453_net85351), .ZN(u4_sll_453_net85343)
         );
  INV_X1 u4_sll_453_U238 ( .A(u4_sll_453_net85315), .ZN(u4_sll_453_n124) );
  NAND2_X2 u4_sll_453_U237 ( .A1(u4_sll_453_n125), .A2(u4_sll_453_n126), .ZN(
        u4_sll_453_ML_int_4__26_) );
  NAND2_X2 u4_sll_453_U236 ( .A1(u4_sll_453_ML_int_3__18_), .A2(
        u4_sll_453_net85315), .ZN(u4_sll_453_n126) );
  INV_X1 u4_sll_453_U235 ( .A(u4_sll_453_net85343), .ZN(u4_sll_453_n121) );
  NAND2_X2 u4_sll_453_U234 ( .A1(u4_sll_453_n122), .A2(u4_sll_453_n123), .ZN(
        u4_sll_453_ML_int_5__42_) );
  NAND2_X2 u4_sll_453_U233 ( .A1(u4_sll_453_ML_int_4__26_), .A2(
        u4_sll_453_net85343), .ZN(u4_sll_453_n123) );
  NAND2_X2 u4_sll_453_U232 ( .A1(u4_sll_453_ML_int_4__42_), .A2(
        u4_sll_453_n121), .ZN(u4_sll_453_n122) );
  MUX2_X2 u4_sll_453_U231 ( .A(u4_sll_453_ML_int_4__40_), .B(
        u4_sll_453_ML_int_4__24_), .S(u4_sll_453_net85349), .Z(
        u4_sll_453_ML_int_5__40_) );
  AND2_X2 u4_sll_453_U230 ( .A1(u4_sll_453_ML_int_5__19_), .A2(
        u4_sll_453_net93645), .ZN(u4_N1427) );
  MUX2_X2 u4_sll_453_U229 ( .A(u4_sll_453_ML_int_2__43_), .B(
        u4_sll_453_ML_int_2__47_), .S(u4_sll_453_net85299), .Z(
        u4_sll_453_ML_int_3__47_) );
  MUX2_X2 u4_sll_453_U228 ( .A(u4_sll_453_ML_int_2__37_), .B(
        u4_sll_453_ML_int_2__33_), .S(u4_sll_453_net85289), .Z(u4_sll_453_n119) );
  INV_X32 u4_sll_453_U227 ( .A(u4_sll_453_net85313), .ZN(u4_sll_453_n118) );
  MUX2_X2 u4_sll_453_U226 ( .A(u4_sll_453_ML_int_3__4_), .B(
        u4_sll_453_ML_int_3__12_), .S(u4_sll_453_n118), .Z(
        u4_sll_453_ML_int_4__12_) );
  AND2_X2 u4_sll_453_U225 ( .A1(u4_sll_453_ML_int_5__22_), .A2(
        u4_sll_453_net93041), .ZN(u4_N1430) );
  INV_X32 u4_sll_453_U224 ( .A(u4_sll_453_net85313), .ZN(u4_sll_453_n117) );
  MUX2_X2 u4_sll_453_U223 ( .A(u4_sll_453_ML_int_3__30_), .B(
        u4_sll_453_ML_int_3__38_), .S(u4_sll_453_n117), .Z(
        u4_sll_453_ML_int_4__38_) );
  NAND2_X2 u4_sll_453_U222 ( .A1(u4_sll_453_n116), .A2(u4_sll_453_n115), .ZN(
        u4_sll_453_ML_int_1__16_) );
  NAND2_X1 u4_sll_453_U221 ( .A1(net17684), .A2(u4_sll_453_n104), .ZN(
        u4_sll_453_n115) );
  NAND2_X2 u4_sll_453_U220 ( .A1(u4_sll_453_n113), .A2(u4_sll_453_n114), .ZN(
        u4_sll_453_ML_int_3__12_) );
  NAND2_X1 u4_sll_453_U219 ( .A1(u4_sll_453_ML_int_2__8_), .A2(
        u4_sll_453_net85287), .ZN(u4_sll_453_n114) );
  NAND2_X2 u4_sll_453_U218 ( .A1(u4_sll_453_ML_int_2__24_), .A2(
        u4_sll_453_net85289), .ZN(u4_sll_453_n208) );
  BUF_X4 u4_sll_453_U217 ( .A(u4_sll_453_ML_int_1__24_), .Z(u4_sll_453_n176)
         );
  INV_X4 u4_sll_453_U216 ( .A(u4_sll_453_net85355), .ZN(u4_sll_453_n109) );
  NAND2_X4 u4_sll_453_U215 ( .A1(u4_sll_453_n110), .A2(u4_sll_453_n111), .ZN(
        u4_N1440) );
  NAND2_X1 u4_sll_453_U214 ( .A1(u4_sll_453_ML_int_5__0_), .A2(
        u4_sll_453_net85355), .ZN(u4_sll_453_n111) );
  NAND2_X4 u4_sll_453_U213 ( .A1(u4_sll_453_ML_int_5__32_), .A2(
        u4_sll_453_n109), .ZN(u4_sll_453_n110) );
  NAND2_X4 u4_sll_453_U212 ( .A1(u4_sll_453_n107), .A2(u4_sll_453_n108), .ZN(
        u4_sll_453_ML_int_2__24_) );
  NAND2_X1 u4_sll_453_U211 ( .A1(u4_sll_453_ML_int_1__22_), .A2(
        u4_sll_453_net85259), .ZN(u4_sll_453_n108) );
  NAND2_X4 u4_sll_453_U210 ( .A1(u4_sll_453_n176), .A2(u4_sll_453_n137), .ZN(
        u4_sll_453_n107) );
  NAND2_X2 u4_sll_453_U209 ( .A1(u4_sll_453_n106), .A2(u4_sll_453_n105), .ZN(
        u4_sll_453_ML_int_1__24_) );
  NAND2_X1 u4_sll_453_U208 ( .A1(fract_denorm[24]), .A2(u4_sll_453_n104), .ZN(
        u4_sll_453_n105) );
  NAND2_X2 u4_sll_453_U207 ( .A1(net17684), .A2(u4_sll_453_net86374), .ZN(
        u4_sll_453_n232) );
  INV_X16 u4_sll_453_U206 ( .A(u4_sll_453_net85237), .ZN(u4_sll_453_net86374)
         );
  NAND2_X2 u4_sll_453_U205 ( .A1(n3006), .A2(u4_sll_453_net94297), .ZN(
        u4_sll_453_n234) );
  AND2_X4 u4_sll_453_U204 ( .A1(u4_sll_453_ML_int_5__28_), .A2(
        u4_sll_453_net85365), .ZN(u4_N1436) );
  INV_X1 u4_sll_453_U203 ( .A(u4_sll_453_net85341), .ZN(u4_sll_453_n147) );
  INV_X4 u4_sll_453_U202 ( .A(u4_sll_453_n147), .ZN(u4_sll_453_n101) );
  NAND2_X2 u4_sll_453_U201 ( .A1(u4_sll_453_n102), .A2(u4_sll_453_n103), .ZN(
        u4_sll_453_ML_int_5__28_) );
  NAND2_X1 u4_sll_453_U200 ( .A1(u4_sll_453_ML_int_4__28_), .A2(
        u4_sll_453_n147), .ZN(u4_sll_453_n103) );
  NAND2_X2 u4_sll_453_U199 ( .A1(u4_sll_453_ML_int_4__12_), .A2(
        u4_sll_453_n101), .ZN(u4_sll_453_n102) );
  NAND2_X2 u4_sll_453_U198 ( .A1(u4_sll_453_ML_int_4__27_), .A2(
        u4_sll_453_net85343), .ZN(u4_sll_453_n212) );
  INV_X1 u4_sll_453_U197 ( .A(u4_sll_453_net85315), .ZN(u4_sll_453_n98) );
  NAND2_X2 u4_sll_453_U196 ( .A1(u4_sll_453_n99), .A2(u4_sll_453_n100), .ZN(
        u4_sll_453_ML_int_4__27_) );
  NAND2_X1 u4_sll_453_U195 ( .A1(u4_sll_453_ML_int_3__19_), .A2(
        u4_sll_453_net85315), .ZN(u4_sll_453_n100) );
  INV_X1 u4_sll_453_U194 ( .A(u4_sll_453_net85261), .ZN(u4_sll_453_n95) );
  NAND2_X2 u4_sll_453_U193 ( .A1(u4_sll_453_n96), .A2(u4_sll_453_n97), .ZN(
        u4_sll_453_ML_int_2__34_) );
  NAND2_X1 u4_sll_453_U192 ( .A1(u4_sll_453_ML_int_1__32_), .A2(
        u4_sll_453_net85261), .ZN(u4_sll_453_n97) );
  INV_X1 u4_sll_453_U191 ( .A(u4_sll_453_net85313), .ZN(u4_sll_453_n120) );
  NAND2_X2 u4_sll_453_U190 ( .A1(u4_sll_453_n93), .A2(u4_sll_453_n94), .ZN(
        u4_sll_453_ML_int_4__43_) );
  NAND2_X2 u4_sll_453_U189 ( .A1(u4_sll_453_ML_int_3__43_), .A2(
        u4_sll_453_n120), .ZN(u4_sll_453_n94) );
  NAND2_X2 u4_sll_453_U188 ( .A1(u4_sll_453_n91), .A2(u4_sll_453_n92), .ZN(
        u4_sll_453_ML_int_3__36_) );
  NAND2_X1 u4_sll_453_U187 ( .A1(u4_sll_453_ML_int_2__32_), .A2(
        u4_sll_453_net85289), .ZN(u4_sll_453_n92) );
  NAND2_X2 u4_sll_453_U186 ( .A1(u4_sll_453_n88), .A2(u4_sll_453_n89), .ZN(
        u4_sll_453_ML_int_1__4_) );
  NAND2_X1 u4_sll_453_U185 ( .A1(net17693), .A2(u4_sll_453_net92610), .ZN(
        u4_sll_453_n88) );
  NAND2_X2 u4_sll_453_U184 ( .A1(u4_sll_453_n86), .A2(u4_sll_453_n87), .ZN(
        u4_sll_453_ML_int_3__21_) );
  NAND2_X1 u4_sll_453_U183 ( .A1(u4_sll_453_ML_int_2__17_), .A2(
        u4_sll_453_net85287), .ZN(u4_sll_453_n87) );
  NAND2_X1 u4_sll_453_U182 ( .A1(u4_sll_453_ML_int_2__21_), .A2(u4_sll_453_n90), .ZN(u4_sll_453_n86) );
  NAND2_X2 u4_sll_453_U181 ( .A1(u4_sll_453_n84), .A2(u4_sll_453_n85), .ZN(
        u4_sll_453_ML_int_1__15_) );
  NAND2_X1 u4_sll_453_U180 ( .A1(net17656), .A2(u4_sll_453_net85231), .ZN(
        u4_sll_453_n85) );
  NAND2_X1 u4_sll_453_U179 ( .A1(net17685), .A2(u4_sll_453_n160), .ZN(
        u4_sll_453_n84) );
  NAND2_X4 u4_sll_453_U178 ( .A1(u4_sll_453_ML_int_4__31_), .A2(
        u4_sll_453_net85339), .ZN(u4_sll_453_n226) );
  NAND2_X2 u4_sll_453_U177 ( .A1(net17690), .A2(u4_sll_453_net86374), .ZN(
        u4_sll_453_net93631) );
  NAND2_X1 u4_sll_453_U176 ( .A1(u4_sll_453_ML_int_1__7_), .A2(
        u4_sll_453_net94113), .ZN(u4_sll_453_n189) );
  INV_X4 u4_sll_453_U175 ( .A(u4_sll_453_net85259), .ZN(u4_sll_453_n171) );
  MUX2_X2 u4_sll_453_U174 ( .A(u4_sll_453_ML_int_1__35_), .B(
        u4_sll_453_ML_int_1__37_), .S(u4_sll_453_n171), .Z(
        u4_sll_453_ML_int_2__37_) );
  INV_X16 u4_sll_453_U173 ( .A(u4_sll_453_net85337), .ZN(u4_sll_453_net85333)
         );
  MUX2_X2 u4_sll_453_U172 ( .A(u4_sll_453_ML_int_4__9_), .B(
        u4_sll_453_ML_int_4__25_), .S(u4_sll_453_net85333), .Z(
        u4_sll_453_ML_int_5__25_) );
  MUX2_X2 u4_sll_453_U171 ( .A(u4_sll_453_ML_int_2__35_), .B(
        u4_sll_453_ML_int_2__39_), .S(u4_sll_453_n83), .Z(
        u4_sll_453_ML_int_3__39_) );
  NAND2_X2 u4_sll_453_U170 ( .A1(u4_sll_453_n148), .A2(u4_sll_453_n149), .ZN(
        u4_sll_453_ML_int_2__10_) );
  INV_X4 u4_sll_453_U169 ( .A(u4_sll_453_net85287), .ZN(u4_sll_453_net93725)
         );
  INV_X4 u4_sll_453_U168 ( .A(u4_sll_453_net85287), .ZN(u4_sll_453_n112) );
  INV_X2 u4_sll_453_U167 ( .A(u4_sll_453_net85285), .ZN(u4_sll_453_net85275)
         );
  INV_X4 u4_sll_453_U166 ( .A(u4_sll_453_net85289), .ZN(u4_sll_453_n83) );
  INV_X8 u4_sll_453_U165 ( .A(u4_shift_left[2]), .ZN(u4_sll_453_net85299) );
  INV_X8 u4_sll_453_U164 ( .A(u4_sll_453_net85289), .ZN(u4_sll_453_n90) );
  INV_X16 u4_sll_453_U163 ( .A(u4_sll_453_net85299), .ZN(u4_sll_453_net85289)
         );
  INV_X16 u4_sll_453_U162 ( .A(u4_shift_left[5]), .ZN(u4_sll_453_net85365) );
  INV_X16 u4_sll_453_U161 ( .A(u4_sll_453_net85365), .ZN(u4_sll_453_net85353)
         );
  INV_X4 u4_sll_453_U160 ( .A(u4_sll_453_net85353), .ZN(u4_sll_453_net93876)
         );
  INV_X16 u4_sll_453_U159 ( .A(u4_shift_left[4]), .ZN(u4_sll_453_net85351) );
  INV_X8 u4_sll_453_U158 ( .A(u4_sll_453_net85351), .ZN(u4_sll_453_net85349)
         );
  INV_X4 u4_sll_453_U157 ( .A(u4_sll_453_net85339), .ZN(u4_sll_453_net94330)
         );
  INV_X2 u4_sll_453_U156 ( .A(u4_sll_453_net85349), .ZN(u4_sll_453_net85347)
         );
  INV_X2 u4_sll_453_U155 ( .A(u4_sll_453_net85347), .ZN(u4_sll_453_net85337)
         );
  INV_X4 u4_sll_453_U154 ( .A(u4_sll_453_net85343), .ZN(u4_sll_453_n163) );
  INV_X2 u4_sll_453_U153 ( .A(u4_sll_453_net95318), .ZN(u4_sll_453_n134) );
  INV_X8 u4_sll_453_U152 ( .A(u4_sll_453_net85259), .ZN(u4_sll_453_n137) );
  NAND2_X2 u4_sll_453_U151 ( .A1(u4_sll_453_ML_int_5__37_), .A2(
        u4_sll_453_net93645), .ZN(u4_sll_453_n219) );
  INV_X32 u4_sll_453_U150 ( .A(u4_sll_453_net85351), .ZN(u4_sll_453_net85341)
         );
  INV_X1 u4_sll_453_U149 ( .A(u4_sll_453_net85341), .ZN(u4_sll_453_n80) );
  NAND2_X2 u4_sll_453_U148 ( .A1(u4_sll_453_n81), .A2(u4_sll_453_n82), .ZN(
        u4_sll_453_ML_int_5__37_) );
  NAND2_X1 u4_sll_453_U147 ( .A1(u4_sll_453_ML_int_4__21_), .A2(
        u4_sll_453_net85341), .ZN(u4_sll_453_n82) );
  NAND2_X2 u4_sll_453_U146 ( .A1(u4_sll_453_ML_int_4__37_), .A2(u4_sll_453_n80), .ZN(u4_sll_453_n81) );
  INV_X1 u4_sll_453_U145 ( .A(u4_sll_453_net85341), .ZN(u4_sll_453_n77) );
  NAND2_X2 u4_sll_453_U144 ( .A1(u4_sll_453_n78), .A2(u4_sll_453_n79), .ZN(
        u4_sll_453_ML_int_5__29_) );
  NAND2_X1 u4_sll_453_U143 ( .A1(u4_sll_453_ML_int_4__13_), .A2(
        u4_sll_453_net85341), .ZN(u4_sll_453_n79) );
  NAND2_X2 u4_sll_453_U142 ( .A1(u4_sll_453_ML_int_4__29_), .A2(u4_sll_453_n77), .ZN(u4_sll_453_n78) );
  NAND2_X2 u4_sll_453_U141 ( .A1(u4_sll_453_ML_int_2__29_), .A2(
        u4_sll_453_net93725), .ZN(u4_sll_453_n217) );
  NAND2_X2 u4_sll_453_U140 ( .A1(u4_sll_453_n75), .A2(u4_sll_453_n76), .ZN(
        u4_sll_453_ML_int_2__29_) );
  NAND2_X2 u4_sll_453_U139 ( .A1(u4_sll_453_ML_int_1__29_), .A2(u4_sll_453_n74), .ZN(u4_sll_453_n75) );
  INV_X1 u4_sll_453_U138 ( .A(u4_sll_453_net85313), .ZN(u4_sll_453_n71) );
  NAND2_X2 u4_sll_453_U137 ( .A1(u4_sll_453_n72), .A2(u4_sll_453_n73), .ZN(
        u4_sll_453_ML_int_4__33_) );
  NAND2_X1 u4_sll_453_U136 ( .A1(u4_sll_453_ML_int_3__25_), .A2(
        u4_sll_453_net85313), .ZN(u4_sll_453_n73) );
  NAND2_X2 u4_sll_453_U135 ( .A1(u4_sll_453_ML_int_3__33_), .A2(u4_sll_453_n71), .ZN(u4_sll_453_n72) );
  NAND2_X2 u4_sll_453_U134 ( .A1(u4_sll_453_ML_int_3__27_), .A2(u4_sll_453_n98), .ZN(u4_sll_453_n99) );
  INV_X32 u4_sll_453_U133 ( .A(u4_sll_453_net85299), .ZN(u4_sll_453_net85287)
         );
  NAND2_X4 u4_sll_453_U132 ( .A1(u4_sll_453_n138), .A2(u4_sll_453_n139), .ZN(
        u4_sll_453_ML_int_2__23_) );
  INV_X1 u4_sll_453_U131 ( .A(u4_sll_453_net85265), .ZN(u4_sll_453_n68) );
  NAND2_X2 u4_sll_453_U130 ( .A1(u4_sll_453_n69), .A2(u4_sll_453_n70), .ZN(
        u4_sll_453_ML_int_2__27_) );
  NAND2_X1 u4_sll_453_U129 ( .A1(u4_sll_453_ML_int_1__27_), .A2(
        u4_sll_453_net85265), .ZN(u4_sll_453_n70) );
  NAND2_X2 u4_sll_453_U128 ( .A1(u4_sll_453_ML_int_1__25_), .A2(u4_sll_453_n68), .ZN(u4_sll_453_n69) );
  INV_X1 u4_sll_453_U127 ( .A(u4_sll_453_net85287), .ZN(u4_sll_453_n65) );
  NAND2_X4 u4_sll_453_U126 ( .A1(u4_sll_453_n66), .A2(u4_sll_453_n67), .ZN(
        u4_sll_453_ML_int_3__27_) );
  NAND2_X2 u4_sll_453_U125 ( .A1(u4_sll_453_ML_int_2__23_), .A2(
        u4_sll_453_net85287), .ZN(u4_sll_453_n67) );
  NAND2_X2 u4_sll_453_U124 ( .A1(u4_sll_453_ML_int_2__27_), .A2(u4_sll_453_n65), .ZN(u4_sll_453_n66) );
  INV_X32 u4_sll_453_U123 ( .A(u4_sll_453_net85341), .ZN(u4_sll_453_n64) );
  MUX2_X2 u4_sll_453_U122 ( .A(u4_sll_453_ML_int_4__11_), .B(
        u4_sll_453_ML_int_4__27_), .S(u4_sll_453_n64), .Z(
        u4_sll_453_ML_int_5__27_) );
  NAND2_X2 u4_sll_453_U121 ( .A1(u4_sll_453_ML_int_1__34_), .A2(u4_sll_453_n95), .ZN(u4_sll_453_n96) );
  NAND2_X2 u4_sll_453_U120 ( .A1(u4_sll_453_ML_int_2__36_), .A2(u4_sll_453_n90), .ZN(u4_sll_453_n91) );
  INV_X1 u4_sll_453_U119 ( .A(u4_sll_453_net94297), .ZN(u4_sll_453_n61) );
  NAND2_X2 u4_sll_453_U118 ( .A1(u4_sll_453_n62), .A2(u4_sll_453_n63), .ZN(
        u4_sll_453_ML_int_1__34_) );
  NAND2_X2 u4_sll_453_U117 ( .A1(fract_denorm[34]), .A2(u4_sll_453_n61), .ZN(
        u4_sll_453_n62) );
  NAND2_X2 u4_sll_453_U116 ( .A1(u4_sll_453_n59), .A2(u4_sll_453_n60), .ZN(
        u4_sll_453_ML_int_2__36_) );
  NAND2_X1 u4_sll_453_U115 ( .A1(u4_sll_453_ML_int_1__34_), .A2(
        u4_sll_453_net85261), .ZN(u4_sll_453_n60) );
  INV_X2 u4_sll_453_U114 ( .A(u4_sll_453_net85229), .ZN(u4_sll_453_n55) );
  NAND2_X2 u4_sll_453_U113 ( .A1(net17695), .A2(u4_sll_453_net86374), .ZN(
        u4_sll_453_n57) );
  NAND2_X1 u4_sll_453_U112 ( .A1(net17694), .A2(u4_sll_453_n55), .ZN(
        u4_sll_453_n56) );
  INV_X2 u4_sll_453_U111 ( .A(u4_sll_453_net85267), .ZN(u4_sll_453_n52) );
  NAND2_X4 u4_sll_453_U110 ( .A1(u4_sll_453_n53), .A2(u4_sll_453_n54), .ZN(
        u4_sll_453_ML_int_2__4_) );
  NAND2_X2 u4_sll_453_U109 ( .A1(u4_sll_453_ML_int_1__4_), .A2(
        u4_sll_453_net85267), .ZN(u4_sll_453_n54) );
  NAND2_X4 u4_sll_453_U108 ( .A1(u4_sll_453_ML_int_1__2_), .A2(u4_sll_453_n52), 
        .ZN(u4_sll_453_n53) );
  INV_X1 u4_sll_453_U107 ( .A(u4_sll_453_net85229), .ZN(u4_sll_453_n49) );
  NAND2_X2 u4_sll_453_U106 ( .A1(u4_sll_453_n50), .A2(u4_sll_453_n51), .ZN(
        u4_sll_453_ML_int_1__26_) );
  NAND2_X1 u4_sll_453_U105 ( .A1(fract_denorm[25]), .A2(u4_sll_453_net86374), 
        .ZN(u4_sll_453_n51) );
  NAND2_X1 u4_sll_453_U104 ( .A1(fract_denorm[26]), .A2(u4_sll_453_n49), .ZN(
        u4_sll_453_n50) );
  INV_X1 u4_sll_453_U103 ( .A(u4_sll_453_net85315), .ZN(u4_sll_453_n46) );
  NAND2_X2 u4_sll_453_U102 ( .A1(u4_sll_453_n47), .A2(u4_sll_453_n48), .ZN(
        u4_sll_453_ML_int_4__30_) );
  NAND2_X1 u4_sll_453_U101 ( .A1(u4_sll_453_ML_int_3__22_), .A2(
        u4_sll_453_net85315), .ZN(u4_sll_453_n48) );
  NAND2_X1 u4_sll_453_U100 ( .A1(u4_sll_453_ML_int_3__30_), .A2(u4_sll_453_n46), .ZN(u4_sll_453_n47) );
  INV_X4 u4_sll_453_U99 ( .A(u4_sll_453_net85353), .ZN(u4_sll_453_n43) );
  NAND2_X4 u4_sll_453_U98 ( .A1(u4_sll_453_n44), .A2(u4_sll_453_n45), .ZN(
        u4_N1447) );
  NAND2_X2 u4_sll_453_U97 ( .A1(u4_sll_453_ML_int_5__7_), .A2(
        u4_sll_453_net85353), .ZN(u4_sll_453_n45) );
  NAND2_X4 u4_sll_453_U96 ( .A1(u4_sll_453_ML_int_5__39_), .A2(u4_sll_453_n43), 
        .ZN(u4_sll_453_n44) );
  INV_X1 u4_sll_453_U95 ( .A(u4_sll_453_net85229), .ZN(u4_sll_453_n40) );
  NAND2_X2 u4_sll_453_U94 ( .A1(u4_sll_453_n42), .A2(u4_sll_453_n41), .ZN(
        u4_sll_453_ML_int_1__39_) );
  NAND2_X1 u4_sll_453_U93 ( .A1(n2552), .A2(u4_sll_453_n40), .ZN(
        u4_sll_453_n41) );
  NAND2_X2 u4_sll_453_U92 ( .A1(u4_sll_453_ML_int_4__11_), .A2(
        u4_sll_453_net85333), .ZN(u4_sll_453_n265) );
  INV_X2 u4_sll_453_U91 ( .A(u4_sll_453_n265), .ZN(u4_sll_453_ML_int_5__11_)
         );
  NAND2_X1 u4_sll_453_U90 ( .A1(u4_sll_453_ML_int_1__36_), .A2(u4_sll_453_n58), 
        .ZN(u4_sll_453_n59) );
  NOR2_X2 u4_sll_453_U89 ( .A1(u4_sll_453_net85355), .A2(u4_sll_453_n180), 
        .ZN(u4_N1423) );
  INV_X1 u4_sll_453_U88 ( .A(u4_sll_453_net85289), .ZN(u4_sll_453_n37) );
  NAND2_X2 u4_sll_453_U87 ( .A1(u4_sll_453_n38), .A2(u4_sll_453_n39), .ZN(
        u4_sll_453_ML_int_3__37_) );
  NAND2_X1 u4_sll_453_U86 ( .A1(u4_sll_453_ML_int_2__33_), .A2(
        u4_sll_453_net85289), .ZN(u4_sll_453_n39) );
  NAND2_X1 u4_sll_453_U85 ( .A1(u4_sll_453_ML_int_2__37_), .A2(u4_sll_453_n37), 
        .ZN(u4_sll_453_n38) );
  INV_X1 u4_sll_453_U84 ( .A(u4_sll_453_net85229), .ZN(u4_sll_453_n34) );
  NAND2_X2 u4_sll_453_U83 ( .A1(u4_sll_453_n35), .A2(u4_sll_453_n36), .ZN(
        u4_sll_453_ML_int_1__18_) );
  NAND2_X1 u4_sll_453_U82 ( .A1(net17683), .A2(u4_sll_453_n34), .ZN(
        u4_sll_453_n35) );
  INV_X1 u4_sll_453_U81 ( .A(u4_sll_453_net85289), .ZN(u4_sll_453_n31) );
  NAND2_X2 u4_sll_453_U80 ( .A1(u4_sll_453_n32), .A2(u4_sll_453_n33), .ZN(
        u4_sll_453_ML_int_3__38_) );
  NAND2_X1 u4_sll_453_U79 ( .A1(u4_sll_453_ML_int_2__34_), .A2(
        u4_sll_453_net85289), .ZN(u4_sll_453_n33) );
  NAND2_X1 u4_sll_453_U78 ( .A1(u4_sll_453_ML_int_2__38_), .A2(u4_sll_453_n31), 
        .ZN(u4_sll_453_n32) );
  INV_X1 u4_sll_453_U77 ( .A(u4_sll_453_net85341), .ZN(u4_sll_453_n28) );
  NAND2_X2 u4_sll_453_U76 ( .A1(u4_sll_453_n29), .A2(u4_sll_453_n30), .ZN(
        u4_sll_453_ML_int_5__38_) );
  NAND2_X1 u4_sll_453_U75 ( .A1(u4_sll_453_ML_int_4__22_), .A2(
        u4_sll_453_net85341), .ZN(u4_sll_453_n30) );
  NAND2_X2 u4_sll_453_U74 ( .A1(u4_sll_453_ML_int_4__38_), .A2(u4_sll_453_n28), 
        .ZN(u4_sll_453_n29) );
  INV_X1 u4_sll_453_U73 ( .A(u4_sll_453_net85261), .ZN(u4_sll_453_n58) );
  INV_X1 u4_sll_453_U72 ( .A(u4_sll_453_net85261), .ZN(u4_sll_453_n74) );
  NAND2_X1 u4_sll_453_U71 ( .A1(u4_sll_453_ML_int_1__27_), .A2(
        u4_sll_453_net85261), .ZN(u4_sll_453_n76) );
  NAND2_X2 u4_sll_453_U70 ( .A1(u4_sll_453_ML_int_3__35_), .A2(u4_sll_453_n134), .ZN(u4_sll_453_n93) );
  NAND2_X2 u4_sll_453_U69 ( .A1(u4_sll_453_n90), .A2(u4_sll_453_ML_int_2__31_), 
        .ZN(u4_sll_453_n156) );
  INV_X1 u4_sll_453_U68 ( .A(u4_sll_453_net85289), .ZN(u4_sll_453_n25) );
  NAND2_X2 u4_sll_453_U67 ( .A1(u4_sll_453_n26), .A2(u4_sll_453_n27), .ZN(
        u4_sll_453_ML_int_3__35_) );
  NAND2_X1 u4_sll_453_U66 ( .A1(u4_sll_453_ML_int_2__31_), .A2(
        u4_sll_453_net85289), .ZN(u4_sll_453_n27) );
  NAND2_X2 u4_sll_453_U65 ( .A1(u4_sll_453_ML_int_2__35_), .A2(u4_sll_453_n25), 
        .ZN(u4_sll_453_n26) );
  INV_X1 u4_sll_453_U64 ( .A(u4_sll_453_net85265), .ZN(u4_sll_453_n22) );
  NAND2_X2 u4_sll_453_U63 ( .A1(u4_sll_453_n23), .A2(u4_sll_453_n24), .ZN(
        u4_sll_453_ML_int_2__31_) );
  NAND2_X1 u4_sll_453_U62 ( .A1(u4_sll_453_ML_int_1__31_), .A2(
        u4_sll_453_net85265), .ZN(u4_sll_453_n24) );
  NAND2_X2 u4_sll_453_U61 ( .A1(u4_sll_453_ML_int_1__29_), .A2(u4_sll_453_n22), 
        .ZN(u4_sll_453_n23) );
  INV_X1 u4_sll_453_U60 ( .A(u4_sll_453_net85315), .ZN(u4_sll_453_n19) );
  NAND2_X4 u4_sll_453_U59 ( .A1(u4_sll_453_n20), .A2(u4_sll_453_n21), .ZN(
        u4_sll_453_ML_int_4__18_) );
  NAND2_X1 u4_sll_453_U58 ( .A1(u4_sll_453_ML_int_3__10_), .A2(
        u4_sll_453_net85315), .ZN(u4_sll_453_n21) );
  NAND2_X2 u4_sll_453_U57 ( .A1(u4_sll_453_ML_int_3__18_), .A2(u4_sll_453_n19), 
        .ZN(u4_sll_453_n20) );
  INV_X4 u4_sll_453_U56 ( .A(u4_sll_453_net85269), .ZN(u4_sll_453_net85267) );
  INV_X1 u4_sll_453_U55 ( .A(u4_sll_453_net85313), .ZN(u4_sll_453_n16) );
  NAND2_X2 u4_sll_453_U54 ( .A1(u4_sll_453_n17), .A2(u4_sll_453_n18), .ZN(
        u4_sll_453_ML_int_4__44_) );
  NAND2_X1 u4_sll_453_U53 ( .A1(u4_sll_453_ML_int_3__36_), .A2(
        u4_sll_453_net85313), .ZN(u4_sll_453_n18) );
  NAND2_X2 u4_sll_453_U52 ( .A1(u4_sll_453_ML_int_3__44_), .A2(u4_sll_453_n16), 
        .ZN(u4_sll_453_n17) );
  MUX2_X2 u4_sll_453_U51 ( .A(n3024), .B(n2552), .S(u4_sll_453_net86374), .Z(
        u4_sll_453_n15) );
  INV_X8 u4_sll_453_U50 ( .A(u4_sll_453_net85237), .ZN(u4_sll_453_net94297) );
  INV_X1 u4_sll_453_U49 ( .A(u4_sll_453_net85313), .ZN(u4_sll_453_n12) );
  NAND2_X2 u4_sll_453_U48 ( .A1(u4_sll_453_n13), .A2(u4_sll_453_n14), .ZN(
        u4_sll_453_ML_int_4__11_) );
  NAND2_X1 u4_sll_453_U47 ( .A1(u4_sll_453_ML_int_3__3_), .A2(
        u4_sll_453_net85313), .ZN(u4_sll_453_n14) );
  NAND2_X1 u4_sll_453_U46 ( .A1(u4_sll_453_ML_int_3__11_), .A2(u4_sll_453_n12), 
        .ZN(u4_sll_453_n13) );
  INV_X4 u4_sll_453_U45 ( .A(u4_sll_453_net94297), .ZN(u4_sll_453_net92610) );
  NAND2_X2 u4_sll_453_U44 ( .A1(n3068), .A2(u4_sll_453_net86374), .ZN(
        u4_sll_453_n106) );
  NAND2_X2 u4_sll_453_U43 ( .A1(u4_sll_453_ML_int_3__16_), .A2(
        u4_sll_453_net85315), .ZN(u4_sll_453_n186) );
  NAND2_X2 u4_sll_453_U42 ( .A1(u4_sll_453_ML_int_2__12_), .A2(u4_sll_453_n112), .ZN(u4_sll_453_n113) );
  INV_X1 u4_sll_453_U41 ( .A(u4_sll_453_net85287), .ZN(u4_sll_453_n9) );
  NAND2_X2 u4_sll_453_U40 ( .A1(u4_sll_453_n10), .A2(u4_sll_453_n11), .ZN(
        u4_sll_453_ML_int_3__16_) );
  NAND2_X1 u4_sll_453_U39 ( .A1(u4_sll_453_ML_int_2__12_), .A2(
        u4_sll_453_net85287), .ZN(u4_sll_453_n11) );
  NAND2_X1 u4_sll_453_U38 ( .A1(u4_sll_453_ML_int_2__16_), .A2(u4_sll_453_n9), 
        .ZN(u4_sll_453_n10) );
  INV_X1 u4_sll_453_U37 ( .A(u4_sll_453_net85265), .ZN(u4_sll_453_n6) );
  NAND2_X2 u4_sll_453_U36 ( .A1(u4_sll_453_n7), .A2(u4_sll_453_n8), .ZN(
        u4_sll_453_ML_int_2__12_) );
  NAND2_X1 u4_sll_453_U35 ( .A1(u4_sll_453_ML_int_1__12_), .A2(
        u4_sll_453_net85265), .ZN(u4_sll_453_n8) );
  NAND2_X2 u4_sll_453_U34 ( .A1(u4_sll_453_ML_int_1__10_), .A2(u4_sll_453_n6), 
        .ZN(u4_sll_453_n7) );
  INV_X32 u4_sll_453_U33 ( .A(u4_sll_453_net85289), .ZN(u4_sll_453_n5) );
  MUX2_X2 u4_sll_453_U32 ( .A(u4_sll_453_ML_int_2__30_), .B(
        u4_sll_453_ML_int_2__34_), .S(u4_sll_453_n5), .Z(
        u4_sll_453_ML_int_3__34_) );
  NAND2_X4 u4_sll_453_U31 ( .A1(u4_sll_453_n132), .A2(u4_sll_453_n133), .ZN(
        u4_N1455) );
  NAND2_X2 u4_sll_453_U30 ( .A1(u4_sll_453_ML_int_5__38_), .A2(
        u4_sll_453_net93728), .ZN(u4_sll_453_n215) );
  NAND2_X2 u4_sll_453_U29 ( .A1(u4_sll_453_ML_int_4__13_), .A2(u4_sll_453_n163), .ZN(u4_sll_453_n263) );
  NAND2_X1 u4_sll_453_U28 ( .A1(u4_sll_453_ML_int_3__26_), .A2(u4_sll_453_n124), .ZN(u4_sll_453_n125) );
  INV_X4 u4_sll_453_U27 ( .A(u4_sll_453_net91550), .ZN(u4_sll_453_n2) );
  NAND2_X2 u4_sll_453_U26 ( .A1(u4_sll_453_n3), .A2(u4_sll_453_n4), .ZN(
        u4_sll_453_ML_int_4__47_) );
  NAND2_X2 u4_sll_453_U25 ( .A1(u4_sll_453_ML_int_3__47_), .A2(
        u4_sll_453_net91550), .ZN(u4_sll_453_n4) );
  NAND2_X2 u4_sll_453_U24 ( .A1(u4_sll_453_ML_int_3__39_), .A2(u4_sll_453_n2), 
        .ZN(u4_sll_453_n3) );
  NAND2_X2 u4_sll_453_U23 ( .A1(u4_sll_453_ML_int_4__14_), .A2(
        u4_sll_453_net85347), .ZN(u4_sll_453_n262) );
  NAND2_X2 u4_sll_453_U22 ( .A1(net17653), .A2(u4_sll_453_net94297), .ZN(
        u4_sll_453_n89) );
  NAND2_X2 u4_sll_453_U21 ( .A1(u4_sll_453_ML_int_5__41_), .A2(u4_sll_453_n109), .ZN(u4_sll_453_n246) );
  INV_X4 u4_sll_453_U20 ( .A(u4_shift_left[1]), .ZN(u4_sll_453_net85271) );
  NAND2_X4 u4_sll_453_U19 ( .A1(net17685), .A2(u4_sll_453_net85231), .ZN(
        u4_sll_453_n116) );
  NAND2_X2 u4_sll_453_U18 ( .A1(u4_sll_453_ML_int_3__24_), .A2(
        u4_sll_453_net94228), .ZN(u4_sll_453_n185) );
  NAND2_X2 u4_sll_453_U17 ( .A1(u4_sll_453_ML_int_2__16_), .A2(
        u4_sll_453_net85287), .ZN(u4_sll_453_n245) );
  INV_X4 u4_sll_453_U16 ( .A(u4_sll_453_net85259), .ZN(u4_sll_453_net93710) );
  INV_X8 u4_sll_453_U15 ( .A(u4_sll_453_net85267), .ZN(u4_sll_453_net85257) );
  INV_X8 u4_sll_453_U14 ( .A(u4_sll_453_net85265), .ZN(u4_sll_453_net85263) );
  INV_X16 u4_sll_453_U13 ( .A(u4_sll_453_net85271), .ZN(u4_sll_453_net85269)
         );
  NAND2_X2 u4_sll_453_U12 ( .A1(u4_sll_453_ML_int_4__29_), .A2(
        u4_sll_453_net85343), .ZN(u4_sll_453_n198) );
  NAND2_X1 u4_sll_453_U11 ( .A1(net17655), .A2(u4_sll_453_net86374), .ZN(
        u4_sll_453_n241) );
  NAND2_X2 u4_sll_453_U10 ( .A1(net17657), .A2(u4_sll_453_net85231), .ZN(
        u4_sll_453_n36) );
  NAND2_X2 u4_sll_453_U9 ( .A1(u4_sll_453_n201), .A2(u4_sll_453_n202), .ZN(
        u4_sll_453_ML_int_1__6_) );
  NAND2_X1 u4_sll_453_U8 ( .A1(net17659), .A2(u4_sll_453_net92610), .ZN(
        u4_sll_453_n248) );
  NAND2_X2 u4_sll_453_U7 ( .A1(u4_sll_453_n56), .A2(u4_sll_453_n57), .ZN(
        u4_sll_453_ML_int_1__2_) );
  NAND2_X2 u4_sll_453_U6 ( .A1(fract_denorm[38]), .A2(u4_sll_453_net85231), 
        .ZN(u4_sll_453_n42) );
  INV_X4 u4_sll_453_U5 ( .A(u4_sll_453_net85231), .ZN(u4_sll_453_n104) );
  NAND2_X1 u4_sll_453_U4 ( .A1(fract_denorm[33]), .A2(u4_sll_453_net85231), 
        .ZN(u4_sll_453_n63) );
  NAND2_X2 u4_sll_453_U3 ( .A1(u4_sll_453_n116), .A2(u4_sll_453_n115), .ZN(
        u4_sll_453_n1) );
  MUX2_X2 u4_sll_453_M1_0_9 ( .A(n2981), .B(net17690), .S(u4_sll_453_net86373), 
        .Z(u4_sll_453_ML_int_1__9_) );
  MUX2_X2 u4_sll_453_M1_3_34 ( .A(u4_sll_453_ML_int_3__34_), .B(
        u4_sll_453_ML_int_3__26_), .S(u4_sll_453_net85313), .Z(
        u4_sll_453_ML_int_4__34_) );
  MUX2_X2 u4_sll_453_M1_0_11 ( .A(net17655), .B(n5324), .S(u4_sll_453_net86373), .Z(u4_sll_453_ML_int_1__11_) );
  MUX2_X2 u4_sll_453_M1_0_10 ( .A(n5324), .B(n2981), .S(u4_sll_453_net85229), 
        .Z(u4_sll_453_ML_int_1__10_) );
  MUX2_X2 u4_sll_453_M1_5_34 ( .A(u4_sll_453_ML_int_5__34_), .B(
        u4_sll_453_ML_int_5__2_), .S(u4_sll_453_net85355), .Z(u4_N1442) );
  MUX2_X2 u4_sll_453_M1_4_18 ( .A(u4_sll_453_ML_int_4__18_), .B(
        u4_sll_453_ML_int_4__2_), .S(u4_sll_453_net85339), .Z(
        u4_sll_453_ML_int_5__18_) );
  MUX2_X2 u4_sll_453_M1_3_42 ( .A(u4_sll_453_ML_int_3__42_), .B(
        u4_sll_453_ML_int_3__34_), .S(u4_sll_453_net85313), .Z(
        u4_sll_453_ML_int_4__42_) );
  MUX2_X2 u4_sll_453_M1_0_7 ( .A(n5323), .B(net17654), .S(u4_sll_453_net86373), 
        .Z(u4_sll_453_ML_int_1__7_) );
  MUX2_X2 u4_sll_453_M1_1_6 ( .A(u4_sll_453_ML_int_1__6_), .B(
        u4_sll_453_ML_int_1__4_), .S(u4_sll_453_net85257), .Z(
        u4_sll_453_ML_int_2__6_) );
  MUX2_X2 u4_sll_453_M1_2_6 ( .A(u4_sll_453_ML_int_2__6_), .B(
        u4_sll_453_ML_int_2__2_), .S(u4_sll_453_net85285), .Z(
        u4_sll_453_ML_int_3__6_) );
  MUX2_X2 u4_sll_453_M1_2_18 ( .A(u4_sll_453_n175), .B(
        u4_sll_453_ML_int_2__14_), .S(u4_sll_453_net85287), .Z(
        u4_sll_453_ML_int_3__18_) );
  MUX2_X2 u4_sll_453_M1_1_13 ( .A(u4_sll_453_ML_int_1__13_), .B(
        u4_sll_453_ML_int_1__11_), .S(u4_sll_453_net85259), .Z(
        u4_sll_453_ML_int_2__13_) );
  MUX2_X1 u4_sll_453_M1_4_24 ( .A(u4_sll_453_ML_int_4__24_), .B(
        u4_sll_453_ML_int_4__8_), .S(u4_sll_453_net85341), .Z(
        u4_sll_453_ML_int_5__24_) );
  MUX2_X2 u4_sll_453_M1_0_1 ( .A(net17695), .B(net17652), .S(
        u4_sll_453_net86374), .Z(u4_sll_453_ML_int_1__1_) );
  MUX2_X2 u4_sll_453_M1_0_3 ( .A(net17653), .B(net17694), .S(
        u4_sll_453_net85231), .Z(u4_sll_453_ML_int_1__3_) );
  MUX2_X2 u4_sll_453_M1_0_5 ( .A(net17692), .B(net17693), .S(
        u4_sll_453_net86374), .Z(u4_sll_453_ML_int_1__5_) );
  MUX2_X2 u4_sll_453_M1_0_13 ( .A(net17686), .B(n5326), .S(u4_sll_453_net86374), .Z(u4_sll_453_ML_int_1__13_) );
  MUX2_X2 u4_sll_453_M1_0_14 ( .A(net17656), .B(net17686), .S(
        u4_sll_453_net86374), .Z(u4_sll_453_ML_int_1__14_) );
  MUX2_X2 u4_sll_453_M1_0_22 ( .A(fract_denorm[22]), .B(fract_denorm[21]), .S(
        u4_sll_453_net85231), .Z(u4_sll_453_ML_int_1__22_) );
  MUX2_X2 u4_sll_453_M1_0_23 ( .A(n3068), .B(fract_denorm[22]), .S(
        u4_sll_453_net85231), .Z(u4_sll_453_ML_int_1__23_) );
  MUX2_X2 u4_sll_453_M1_0_25 ( .A(fract_denorm[25]), .B(fract_denorm[24]), .S(
        u4_sll_453_net94297), .Z(u4_sll_453_ML_int_1__25_) );
  MUX2_X2 u4_sll_453_M1_0_27 ( .A(n2546), .B(fract_denorm[26]), .S(
        u4_sll_453_net85229), .Z(u4_sll_453_ML_int_1__27_) );
  MUX2_X2 u4_sll_453_M1_0_28 ( .A(n2937), .B(n2546), .S(u4_sll_453_net86373), 
        .Z(u4_sll_453_ML_int_1__28_) );
  MUX2_X2 u4_sll_453_M1_0_29 ( .A(n3006), .B(n2937), .S(u4_sll_453_net85229), 
        .Z(u4_sll_453_ML_int_1__29_) );
  MUX2_X2 u4_sll_453_M1_0_31 ( .A(fract_denorm[31]), .B(n3008), .S(
        u4_sll_453_net86373), .Z(u4_sll_453_ML_int_1__31_) );
  MUX2_X2 u4_sll_453_M1_0_32 ( .A(fract_denorm[32]), .B(fract_denorm[31]), .S(
        u4_sll_453_net94297), .Z(u4_sll_453_ML_int_1__32_) );
  MUX2_X2 u4_sll_453_M1_0_33 ( .A(fract_denorm[33]), .B(fract_denorm[32]), .S(
        u4_sll_453_net86374), .Z(u4_sll_453_ML_int_1__33_) );
  MUX2_X2 u4_sll_453_M1_0_35 ( .A(net94442), .B(fract_denorm[34]), .S(
        u4_sll_453_net94297), .Z(u4_sll_453_ML_int_1__35_) );
  MUX2_X2 u4_sll_453_M1_0_36 ( .A(fract_denorm[36]), .B(net94442), .S(
        u4_sll_453_net86373), .Z(u4_sll_453_ML_int_1__36_) );
  MUX2_X2 u4_sll_453_M1_0_37 ( .A(fract_denorm[37]), .B(fract_denorm[36]), .S(
        u4_sll_453_net86373), .Z(u4_sll_453_ML_int_1__37_) );
  MUX2_X2 u4_sll_453_M1_0_38 ( .A(fract_denorm[38]), .B(fract_denorm[37]), .S(
        u4_sll_453_net86373), .Z(u4_sll_453_ML_int_1__38_) );
  MUX2_X2 u4_sll_453_M1_0_40 ( .A(n3024), .B(n2552), .S(u4_sll_453_net86373), 
        .Z(u4_sll_453_ML_int_1__40_) );
  MUX2_X2 u4_sll_453_M1_0_41 ( .A(net28939), .B(n3024), .S(u4_sll_453_net86373), .Z(u4_sll_453_ML_int_1__41_) );
  MUX2_X2 u4_sll_453_M1_0_42 ( .A(net94305), .B(net28939), .S(
        u4_sll_453_net86373), .Z(u4_sll_453_ML_int_1__42_) );
  MUX2_X2 u4_sll_453_M1_0_43 ( .A(fract_denorm[43]), .B(net94305), .S(
        u4_sll_453_net94297), .Z(u4_sll_453_ML_int_1__43_) );
  MUX2_X2 u4_sll_453_M1_0_44 ( .A(fract_denorm[44]), .B(fract_denorm[43]), .S(
        u4_sll_453_net94297), .Z(u4_sll_453_ML_int_1__44_) );
  MUX2_X2 u4_sll_453_M1_0_45 ( .A(net91595), .B(fract_denorm[44]), .S(
        u4_sll_453_net85229), .Z(u4_sll_453_ML_int_1__45_) );
  MUX2_X2 u4_sll_453_M1_0_46 ( .A(net86571), .B(net91595), .S(
        u4_sll_453_net85229), .Z(u4_sll_453_ML_int_1__46_) );
  MUX2_X2 u4_sll_453_M1_0_47 ( .A(net85391), .B(net86571), .S(
        u4_sll_453_net85229), .Z(u4_sll_453_ML_int_1__47_) );
  MUX2_X2 u4_sll_453_M1_1_2 ( .A(u4_sll_453_ML_int_1__2_), .B(
        u4_sll_453_ML_int_1__0_), .S(u4_sll_453_net85257), .Z(
        u4_sll_453_ML_int_2__2_) );
  MUX2_X2 u4_sll_453_M1_1_3 ( .A(u4_sll_453_ML_int_1__3_), .B(
        u4_sll_453_ML_int_1__1_), .S(u4_sll_453_net85257), .Z(
        u4_sll_453_ML_int_2__3_) );
  MUX2_X2 u4_sll_453_M1_1_11 ( .A(u4_sll_453_ML_int_1__11_), .B(
        u4_sll_453_ML_int_1__9_), .S(u4_sll_453_net85259), .Z(
        u4_sll_453_ML_int_2__11_) );
  MUX2_X2 u4_sll_453_M1_1_14 ( .A(u4_sll_453_ML_int_1__14_), .B(
        u4_sll_453_ML_int_1__12_), .S(u4_sll_453_net85259), .Z(
        u4_sll_453_ML_int_2__14_) );
  MUX2_X2 u4_sll_453_M1_1_16 ( .A(u4_sll_453_n1), .B(u4_sll_453_ML_int_1__14_), 
        .S(u4_sll_453_net85259), .Z(u4_sll_453_ML_int_2__16_) );
  MUX2_X2 u4_sll_453_M1_1_18 ( .A(u4_sll_453_ML_int_1__18_), .B(
        u4_sll_453_ML_int_1__16_), .S(u4_sll_453_net85259), .Z(
        u4_sll_453_ML_int_2__18_) );
  MUX2_X2 u4_sll_453_M1_1_19 ( .A(u4_sll_453_ML_int_1__19_), .B(
        u4_sll_453_ML_int_1__17_), .S(u4_sll_453_net85259), .Z(
        u4_sll_453_ML_int_2__19_) );
  MUX2_X2 u4_sll_453_M1_1_20 ( .A(u4_sll_453_ML_int_1__20_), .B(
        u4_sll_453_ML_int_1__18_), .S(u4_sll_453_net85259), .Z(
        u4_sll_453_ML_int_2__20_) );
  MUX2_X2 u4_sll_453_M1_1_25 ( .A(u4_sll_453_ML_int_1__25_), .B(
        u4_sll_453_ML_int_1__23_), .S(u4_sll_453_net85259), .Z(
        u4_sll_453_ML_int_2__25_) );
  MUX2_X2 u4_sll_453_M1_1_26 ( .A(u4_sll_453_ML_int_1__26_), .B(
        u4_sll_453_ML_int_1__24_), .S(u4_sll_453_net85261), .Z(
        u4_sll_453_ML_int_2__26_) );
  MUX2_X2 u4_sll_453_M1_1_28 ( .A(u4_sll_453_ML_int_1__28_), .B(
        u4_sll_453_ML_int_1__26_), .S(u4_sll_453_net85261), .Z(
        u4_sll_453_ML_int_2__28_) );
  MUX2_X2 u4_sll_453_M1_1_32 ( .A(u4_sll_453_ML_int_1__32_), .B(
        u4_sll_453_ML_int_1__30_), .S(u4_sll_453_net85261), .Z(
        u4_sll_453_ML_int_2__32_) );
  MUX2_X2 u4_sll_453_M1_1_33 ( .A(u4_sll_453_ML_int_1__33_), .B(
        u4_sll_453_ML_int_1__31_), .S(u4_sll_453_net85261), .Z(
        u4_sll_453_ML_int_2__33_) );
  MUX2_X2 u4_sll_453_M1_1_35 ( .A(u4_sll_453_ML_int_1__35_), .B(
        u4_sll_453_ML_int_1__33_), .S(u4_sll_453_net85261), .Z(
        u4_sll_453_ML_int_2__35_) );
  MUX2_X2 u4_sll_453_M1_1_38 ( .A(u4_sll_453_ML_int_1__38_), .B(
        u4_sll_453_ML_int_1__36_), .S(u4_sll_453_net85261), .Z(
        u4_sll_453_ML_int_2__38_) );
  MUX2_X2 u4_sll_453_M1_1_39 ( .A(u4_sll_453_ML_int_1__39_), .B(
        u4_sll_453_ML_int_1__37_), .S(u4_sll_453_net85261), .Z(
        u4_sll_453_ML_int_2__39_) );
  MUX2_X2 u4_sll_453_M1_1_40 ( .A(u4_sll_453_n15), .B(u4_sll_453_ML_int_1__38_), .S(u4_sll_453_net85261), .Z(u4_sll_453_ML_int_2__40_) );
  MUX2_X2 u4_sll_453_M1_1_41 ( .A(u4_sll_453_ML_int_1__41_), .B(
        u4_sll_453_ML_int_1__39_), .S(u4_sll_453_net85261), .Z(
        u4_sll_453_ML_int_2__41_) );
  MUX2_X2 u4_sll_453_M1_1_42 ( .A(u4_sll_453_ML_int_1__42_), .B(
        u4_sll_453_ML_int_1__40_), .S(u4_sll_453_net85261), .Z(
        u4_sll_453_ML_int_2__42_) );
  MUX2_X2 u4_sll_453_M1_1_43 ( .A(u4_sll_453_ML_int_1__43_), .B(
        u4_sll_453_ML_int_1__41_), .S(u4_sll_453_net85261), .Z(
        u4_sll_453_ML_int_2__43_) );
  MUX2_X2 u4_sll_453_M1_1_44 ( .A(u4_sll_453_ML_int_1__44_), .B(
        u4_sll_453_ML_int_1__42_), .S(u4_sll_453_net85263), .Z(
        u4_sll_453_ML_int_2__44_) );
  MUX2_X2 u4_sll_453_M1_1_45 ( .A(u4_sll_453_ML_int_1__45_), .B(
        u4_sll_453_ML_int_1__43_), .S(u4_sll_453_net85263), .Z(
        u4_sll_453_ML_int_2__45_) );
  MUX2_X2 u4_sll_453_M1_1_46 ( .A(u4_sll_453_ML_int_1__46_), .B(
        u4_sll_453_ML_int_1__44_), .S(u4_sll_453_net85263), .Z(
        u4_sll_453_ML_int_2__46_) );
  MUX2_X2 u4_sll_453_M1_2_4 ( .A(u4_sll_453_ML_int_2__4_), .B(
        u4_sll_453_ML_int_2__0_), .S(u4_sll_453_net85285), .Z(
        u4_sll_453_ML_int_3__4_) );
  MUX2_X2 u4_sll_453_M1_2_5 ( .A(u4_sll_453_ML_int_2__5_), .B(
        u4_sll_453_ML_int_2__1_), .S(u4_sll_453_net85285), .Z(
        u4_sll_453_ML_int_3__5_) );
  MUX2_X2 u4_sll_453_M1_2_7 ( .A(u4_sll_453_ML_int_2__7_), .B(
        u4_sll_453_ML_int_2__3_), .S(u4_sll_453_net85285), .Z(
        u4_sll_453_ML_int_3__7_) );
  MUX2_X2 u4_sll_453_M1_2_9 ( .A(u4_sll_453_ML_int_2__9_), .B(
        u4_sll_453_ML_int_2__5_), .S(u4_sll_453_net85285), .Z(
        u4_sll_453_ML_int_3__9_) );
  MUX2_X2 u4_sll_453_M1_2_26 ( .A(u4_sll_453_ML_int_2__26_), .B(
        u4_sll_453_ML_int_2__22_), .S(u4_sll_453_net85287), .Z(
        u4_sll_453_ML_int_3__26_) );
  MUX2_X2 u4_sll_453_M1_2_30 ( .A(u4_sll_453_ML_int_2__30_), .B(
        u4_sll_453_ML_int_2__26_), .S(u4_sll_453_net85289), .Z(
        u4_sll_453_ML_int_3__30_) );
  MUX2_X2 u4_sll_453_M1_2_33 ( .A(u4_sll_453_ML_int_2__33_), .B(
        u4_sll_453_ML_int_2__29_), .S(u4_sll_453_net85289), .Z(
        u4_sll_453_ML_int_3__33_) );
  MUX2_X2 u4_sll_453_M1_2_40 ( .A(u4_sll_453_ML_int_2__40_), .B(
        u4_sll_453_ML_int_2__36_), .S(u4_sll_453_net85289), .Z(
        u4_sll_453_ML_int_3__40_) );
  MUX2_X2 u4_sll_453_M1_2_41 ( .A(u4_sll_453_ML_int_2__41_), .B(
        u4_sll_453_ML_int_2__37_), .S(u4_sll_453_net85289), .Z(
        u4_sll_453_ML_int_3__41_) );
  MUX2_X2 u4_sll_453_M1_2_42 ( .A(u4_sll_453_ML_int_2__42_), .B(
        u4_sll_453_ML_int_2__38_), .S(u4_sll_453_net85289), .Z(
        u4_sll_453_ML_int_3__42_) );
  MUX2_X2 u4_sll_453_M1_2_43 ( .A(u4_sll_453_ML_int_2__43_), .B(
        u4_sll_453_ML_int_2__39_), .S(u4_sll_453_net85289), .Z(
        u4_sll_453_ML_int_3__43_) );
  MUX2_X2 u4_sll_453_M1_2_44 ( .A(u4_sll_453_ML_int_2__44_), .B(
        u4_sll_453_ML_int_2__40_), .S(u4_sll_453_net85289), .Z(
        u4_sll_453_ML_int_3__44_) );
  MUX2_X2 u4_sll_453_M1_2_45 ( .A(u4_sll_453_ML_int_2__45_), .B(
        u4_sll_453_ML_int_2__41_), .S(u4_sll_453_net85289), .Z(
        u4_sll_453_ML_int_3__45_) );
  MUX2_X2 u4_sll_453_M1_2_46 ( .A(u4_sll_453_ML_int_2__46_), .B(
        u4_sll_453_ML_int_2__42_), .S(u4_sll_453_net85289), .Z(
        u4_sll_453_ML_int_3__46_) );
  MUX2_X2 u4_sll_453_M1_3_8 ( .A(u4_sll_453_ML_int_3__8_), .B(
        u4_sll_453_ML_int_3__0_), .S(u4_sll_453_net85313), .Z(
        u4_sll_453_ML_int_4__8_) );
  MUX2_X2 u4_sll_453_M1_3_9 ( .A(u4_sll_453_ML_int_3__9_), .B(
        u4_sll_453_ML_int_3__1_), .S(u4_sll_453_net85313), .Z(
        u4_sll_453_ML_int_4__9_) );
  MUX2_X2 u4_sll_453_M1_3_10 ( .A(u4_sll_453_ML_int_3__10_), .B(
        u4_sll_453_ML_int_3__2_), .S(u4_sll_453_net85313), .Z(
        u4_sll_453_ML_int_4__10_) );
  MUX2_X2 u4_sll_453_M1_3_13 ( .A(u4_sll_453_n239), .B(u4_sll_453_ML_int_3__5_), .S(u4_sll_453_net85313), .Z(u4_sll_453_ML_int_4__13_) );
  MUX2_X2 u4_sll_453_M1_3_14 ( .A(u4_sll_453_ML_int_3__14_), .B(
        u4_sll_453_ML_int_3__6_), .S(u4_sll_453_net85315), .Z(
        u4_sll_453_ML_int_4__14_) );
  MUX2_X2 u4_sll_453_M1_3_16 ( .A(u4_sll_453_ML_int_3__16_), .B(
        u4_sll_453_ML_int_3__8_), .S(u4_sll_453_net85315), .Z(
        u4_sll_453_ML_int_4__16_) );
  MUX2_X2 u4_sll_453_M1_3_19 ( .A(u4_sll_453_ML_int_3__19_), .B(
        u4_sll_453_ML_int_3__11_), .S(u4_sll_453_net85315), .Z(
        u4_sll_453_ML_int_4__19_) );
  MUX2_X2 u4_sll_453_M1_3_20 ( .A(u4_sll_453_ML_int_3__20_), .B(
        u4_sll_453_ML_int_3__12_), .S(u4_sll_453_net85315), .Z(
        u4_sll_453_ML_int_4__20_) );
  MUX2_X2 u4_sll_453_M1_3_21 ( .A(u4_sll_453_ML_int_3__21_), .B(
        u4_sll_453_ML_int_3__13_), .S(u4_sll_453_net85315), .Z(
        u4_sll_453_ML_int_4__21_) );
  MUX2_X2 u4_sll_453_M1_3_22 ( .A(u4_sll_453_n177), .B(
        u4_sll_453_ML_int_3__14_), .S(u4_sll_453_net85315), .Z(
        u4_sll_453_ML_int_4__22_) );
  MUX2_X2 u4_sll_453_M1_3_23 ( .A(u4_sll_453_ML_int_3__23_), .B(
        u4_sll_453_ML_int_3__15_), .S(u4_sll_453_net85315), .Z(
        u4_sll_453_ML_int_4__23_) );
  MUX2_X2 u4_sll_453_M1_3_28 ( .A(u4_sll_453_ML_int_3__28_), .B(
        u4_sll_453_ML_int_3__20_), .S(u4_sll_453_net85315), .Z(
        u4_sll_453_ML_int_4__28_) );
  MUX2_X2 u4_sll_453_M1_3_32 ( .A(u4_sll_453_ML_int_3__32_), .B(
        u4_sll_453_ML_int_3__24_), .S(u4_sll_453_net85313), .Z(
        u4_sll_453_ML_int_4__32_) );
  MUX2_X2 u4_sll_453_M1_3_35 ( .A(u4_sll_453_ML_int_3__35_), .B(
        u4_sll_453_ML_int_3__27_), .S(u4_sll_453_net85313), .Z(
        u4_sll_453_ML_int_4__35_) );
  MUX2_X2 u4_sll_453_M1_3_36 ( .A(u4_sll_453_ML_int_3__36_), .B(
        u4_sll_453_ML_int_3__28_), .S(u4_sll_453_net85313), .Z(
        u4_sll_453_ML_int_4__36_) );
  MUX2_X2 u4_sll_453_M1_3_37 ( .A(u4_sll_453_n119), .B(
        u4_sll_453_ML_int_3__29_), .S(u4_sll_453_net85313), .Z(
        u4_sll_453_ML_int_4__37_) );
  MUX2_X2 u4_sll_453_M1_3_39 ( .A(u4_sll_453_ML_int_3__39_), .B(
        u4_sll_453_ML_int_3__31_), .S(u4_sll_453_net85313), .Z(
        u4_sll_453_ML_int_4__39_) );
  MUX2_X2 u4_sll_453_M1_3_40 ( .A(u4_sll_453_ML_int_3__40_), .B(
        u4_sll_453_ML_int_3__32_), .S(u4_sll_453_net85313), .Z(
        u4_sll_453_ML_int_4__40_) );
  MUX2_X2 u4_sll_453_M1_3_41 ( .A(u4_sll_453_ML_int_3__41_), .B(
        u4_sll_453_ML_int_3__33_), .S(u4_sll_453_net85313), .Z(
        u4_sll_453_ML_int_4__41_) );
  MUX2_X2 u4_sll_453_M1_3_45 ( .A(u4_sll_453_ML_int_3__45_), .B(
        u4_sll_453_ML_int_3__37_), .S(u4_sll_453_net85313), .Z(
        u4_sll_453_ML_int_4__45_) );
  MUX2_X2 u4_sll_453_M1_3_46 ( .A(u4_sll_453_ML_int_3__46_), .B(
        u4_sll_453_ML_int_3__38_), .S(u4_sll_453_net85313), .Z(
        u4_sll_453_ML_int_4__46_) );
  MUX2_X2 u4_sll_453_M1_4_16 ( .A(u4_sll_453_ML_int_4__16_), .B(
        u4_sll_453_ML_int_4__0_), .S(u4_sll_453_net85339), .Z(
        u4_sll_453_ML_int_5__16_) );
  MUX2_X2 u4_sll_453_M1_4_17 ( .A(u4_sll_453_ML_int_4__17_), .B(
        u4_sll_453_ML_int_4__1_), .S(u4_sll_453_net85339), .Z(
        u4_sll_453_ML_int_5__17_) );
  MUX2_X2 u4_sll_453_M1_4_19 ( .A(u4_sll_453_ML_int_4__19_), .B(
        u4_sll_453_ML_int_4__3_), .S(u4_sll_453_net85339), .Z(
        u4_sll_453_ML_int_5__19_) );
  MUX2_X2 u4_sll_453_M1_4_20 ( .A(u4_sll_453_ML_int_4__20_), .B(
        u4_sll_453_ML_int_4__4_), .S(u4_sll_453_net85339), .Z(
        u4_sll_453_ML_int_5__20_) );
  MUX2_X2 u4_sll_453_M1_4_22 ( .A(u4_sll_453_ML_int_4__22_), .B(
        u4_sll_453_ML_int_4__6_), .S(u4_sll_453_net85341), .Z(
        u4_sll_453_ML_int_5__22_) );
  MUX2_X2 u4_sll_453_M1_4_23 ( .A(u4_sll_453_ML_int_4__23_), .B(
        u4_sll_453_ML_int_4__7_), .S(u4_sll_453_net85341), .Z(
        u4_sll_453_ML_int_5__23_) );
  MUX2_X2 u4_sll_453_M1_4_26 ( .A(u4_sll_453_ML_int_4__26_), .B(
        u4_sll_453_ML_int_4__10_), .S(u4_sll_453_net85341), .Z(
        u4_sll_453_ML_int_5__26_) );
  MUX2_X2 u4_sll_453_M1_4_35 ( .A(u4_sll_453_ML_int_4__35_), .B(
        u4_sll_453_ML_int_4__19_), .S(u4_sll_453_net85341), .Z(
        u4_sll_453_ML_int_5__35_) );
  MUX2_X2 u4_sll_453_M1_4_44 ( .A(u4_sll_453_ML_int_4__44_), .B(
        u4_sll_453_ML_int_4__28_), .S(u4_sll_453_net85343), .Z(
        u4_sll_453_ML_int_5__44_) );
  MUX2_X2 u4_sll_453_M1_4_46 ( .A(u4_sll_453_ML_int_4__46_), .B(
        u4_sll_453_ML_int_4__30_), .S(u4_sll_453_net85343), .Z(
        u4_sll_453_ML_int_5__46_) );
  MUX2_X2 u4_sll_453_M1_5_33 ( .A(u4_sll_453_ML_int_5__33_), .B(
        u4_sll_453_ML_int_5__1_), .S(u4_sll_453_net85355), .Z(u4_N1441) );
  MUX2_X2 u4_sll_453_M1_5_36 ( .A(u4_sll_453_ML_int_5__36_), .B(
        u4_sll_453_ML_int_5__4_), .S(u4_sll_453_net85355), .Z(u4_N1444) );
  MUX2_X2 u4_sll_453_M1_5_43 ( .A(u4_sll_453_ML_int_5__43_), .B(
        u4_sll_453_ML_int_5__11_), .S(u4_sll_453_net85353), .Z(u4_N1451) );
  MUX2_X2 u4_sll_453_M1_5_45 ( .A(u4_sll_453_ML_int_5__45_), .B(
        u4_sll_453_ML_int_5__13_), .S(u4_sll_453_net85353), .Z(u4_N1453) );
  INV_X1 u4_srl_452_U359 ( .A(u4_shift_right[2]), .ZN(u4_srl_452_n306) );
  INV_X1 u4_srl_452_U358 ( .A(u4_shift_right[3]), .ZN(u4_srl_452_n259) );
  NAND2_X1 u4_srl_452_U357 ( .A1(u4_srl_452_n306), .A2(u4_srl_452_n259), .ZN(
        u4_srl_452_n279) );
  NOR2_X1 u4_srl_452_U356 ( .A1(u4_srl_452_n279), .A2(u4_shift_right[4]), .ZN(
        u4_srl_452_n135) );
  AOI22_X1 u4_srl_452_U355 ( .A1(net17695), .A2(u4_srl_452_n19), .B1(net17652), 
        .B2(u4_srl_452_n22), .ZN(u4_srl_452_n308) );
  OAI221_X1 u4_srl_452_U354 ( .B1(u4_srl_452_n13), .B2(u4_srl_452_n71), .C1(
        u4_srl_452_n144), .C2(u4_srl_452_n27), .A(u4_srl_452_n308), .ZN(
        u4_srl_452_n294) );
  AOI22_X1 u4_srl_452_U353 ( .A1(n2980), .A2(u4_srl_452_n20), .B1(net17690), 
        .B2(u4_srl_452_n23), .ZN(u4_srl_452_n307) );
  OAI221_X1 u4_srl_452_U352 ( .B1(u4_srl_452_n13), .B2(u4_srl_452_n69), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n32), .A(u4_srl_452_n307), .ZN(
        u4_srl_452_n93) );
  AOI22_X1 u4_srl_452_U351 ( .A1(net17686), .A2(u4_srl_452_n20), .B1(n5326), 
        .B2(u4_srl_452_n23), .ZN(u4_srl_452_n305) );
  OAI221_X1 u4_srl_452_U350 ( .B1(u4_srl_452_n13), .B2(u4_srl_452_n36), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n68), .A(u4_srl_452_n305), .ZN(
        u4_srl_452_n89) );
  AOI22_X1 u4_srl_452_U349 ( .A1(net17692), .A2(u4_srl_452_n20), .B1(net17693), 
        .B2(u4_srl_452_n23), .ZN(u4_srl_452_n304) );
  OAI221_X1 u4_srl_452_U348 ( .B1(u4_srl_452_n13), .B2(u4_srl_452_n30), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n70), .A(u4_srl_452_n304), .ZN(
        u4_srl_452_n123) );
  NAND2_X1 u4_srl_452_U347 ( .A1(u4_shift_right[2]), .A2(u4_srl_452_n259), 
        .ZN(u4_srl_452_n276) );
  AOI222_X1 u4_srl_452_U346 ( .A1(u4_srl_452_n93), .A2(u4_srl_452_n141), .B1(
        u4_srl_452_n89), .B2(u4_srl_452_n142), .C1(u4_srl_452_n123), .C2(
        u4_srl_452_n10), .ZN(u4_srl_452_n297) );
  AOI22_X1 u4_srl_452_U345 ( .A1(n3006), .A2(u4_srl_452_n20), .B1(
        fract_denorm[28]), .B2(u4_srl_452_n23), .ZN(u4_srl_452_n303) );
  OAI221_X1 u4_srl_452_U344 ( .B1(u4_srl_452_n13), .B2(u4_srl_452_n57), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n47), .A(u4_srl_452_n303), .ZN(
        u4_srl_452_n178) );
  AOI22_X1 u4_srl_452_U343 ( .A1(fract_denorm[25]), .A2(u4_srl_452_n20), .B1(
        u4_srl_452_n22), .B2(fract_denorm[24]), .ZN(u4_srl_452_n302) );
  OAI221_X1 u4_srl_452_U342 ( .B1(u4_srl_452_n13), .B2(u4_srl_452_n45), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n44), .A(u4_srl_452_n302), .ZN(
        u4_srl_452_n179) );
  AOI22_X1 u4_srl_452_U341 ( .A1(fract_denorm[21]), .A2(u4_srl_452_n20), .B1(
        net17659), .B2(u4_srl_452_n23), .ZN(u4_srl_452_n301) );
  OAI221_X1 u4_srl_452_U340 ( .B1(u4_srl_452_n13), .B2(u4_srl_452_n49), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n41), .A(u4_srl_452_n301), .ZN(
        u4_srl_452_n90) );
  AOI22_X1 u4_srl_452_U339 ( .A1(net17657), .A2(u4_srl_452_n20), .B1(net17684), 
        .B2(u4_srl_452_n23), .ZN(u4_srl_452_n300) );
  OAI221_X1 u4_srl_452_U338 ( .B1(u4_srl_452_n13), .B2(u4_srl_452_n39), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n38), .A(u4_srl_452_n300), .ZN(
        u4_srl_452_n91) );
  AOI22_X1 u4_srl_452_U337 ( .A1(u4_srl_452_n143), .A2(u4_srl_452_n90), .B1(
        u4_srl_452_n164), .B2(u4_srl_452_n91), .ZN(u4_srl_452_n299) );
  INV_X1 u4_srl_452_U336 ( .A(u4_srl_452_n299), .ZN(u4_srl_452_n298) );
  AOI221_X1 u4_srl_452_U335 ( .B1(u4_srl_452_n178), .B2(u4_srl_452_n142), .C1(
        u4_srl_452_n179), .C2(u4_srl_452_n141), .A(u4_srl_452_n298), .ZN(
        u4_srl_452_n230) );
  MUX2_X1 u4_srl_452_U334 ( .A(u4_srl_452_n297), .B(u4_srl_452_n230), .S(
        u4_shift_right[4]), .Z(u4_srl_452_n296) );
  INV_X1 u4_srl_452_U333 ( .A(u4_srl_452_n296), .ZN(u4_srl_452_n295) );
  AOI21_X1 u4_srl_452_U332 ( .B1(u4_srl_452_n135), .B2(u4_srl_452_n294), .A(
        u4_srl_452_n295), .ZN(u4_srl_452_n288) );
  AOI22_X1 u4_srl_452_U331 ( .A1(fract_denorm[37]), .A2(u4_srl_452_n20), .B1(
        fract_denorm[36]), .B2(u4_srl_452_n23), .ZN(u4_srl_452_n293) );
  OAI221_X1 u4_srl_452_U330 ( .B1(u4_srl_452_n13), .B2(u4_srl_452_n58), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n55), .A(u4_srl_452_n293), .ZN(
        u4_srl_452_n206) );
  AOI22_X1 u4_srl_452_U329 ( .A1(fract_denorm[33]), .A2(u4_srl_452_n20), .B1(
        fract_denorm[32]), .B2(u4_srl_452_n23), .ZN(u4_srl_452_n292) );
  OAI221_X1 u4_srl_452_U328 ( .B1(u4_srl_452_n13), .B2(u4_srl_452_n53), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n52), .A(u4_srl_452_n292), .ZN(
        u4_srl_452_n183) );
  AOI22_X1 u4_srl_452_U327 ( .A1(fract_denorm[45]), .A2(u4_srl_452_n20), .B1(
        fract_denorm[44]), .B2(u4_srl_452_n23), .ZN(u4_srl_452_n291) );
  OAI221_X1 u4_srl_452_U326 ( .B1(u4_srl_452_n13), .B2(u4_srl_452_n26), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n62), .A(u4_srl_452_n291), .ZN(
        u4_srl_452_n177) );
  INV_X1 u4_srl_452_U325 ( .A(u4_srl_452_n177), .ZN(u4_srl_452_n129) );
  AOI22_X1 u4_srl_452_U324 ( .A1(net28939), .A2(u4_srl_452_n20), .B1(n3024), 
        .B2(u4_srl_452_n23), .ZN(u4_srl_452_n290) );
  OAI221_X1 u4_srl_452_U323 ( .B1(u4_srl_452_n13), .B2(u4_srl_452_n63), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n65), .A(u4_srl_452_n290), .ZN(
        u4_srl_452_n176) );
  INV_X1 u4_srl_452_U322 ( .A(u4_srl_452_n176), .ZN(u4_srl_452_n254) );
  OAI22_X1 u4_srl_452_U321 ( .A1(u4_srl_452_n172), .A2(u4_srl_452_n129), .B1(
        u4_srl_452_n174), .B2(u4_srl_452_n254), .ZN(u4_srl_452_n289) );
  AOI221_X1 u4_srl_452_U320 ( .B1(u4_srl_452_n206), .B2(u4_srl_452_n143), .C1(
        u4_srl_452_n183), .C2(u4_srl_452_n164), .A(u4_srl_452_n289), .ZN(
        u4_srl_452_n150) );
  INV_X1 u4_srl_452_U319 ( .A(u4_shift_right[4]), .ZN(u4_srl_452_n280) );
  NAND2_X1 u4_srl_452_U318 ( .A1(u4_shift_right[5]), .A2(u4_srl_452_n280), 
        .ZN(u4_srl_452_n134) );
  OAI22_X1 u4_srl_452_U317 ( .A1(u4_shift_right[5]), .A2(u4_srl_452_n288), 
        .B1(u4_srl_452_n150), .B2(u4_srl_452_n134), .ZN(u4_N1358) );
  AOI22_X1 u4_srl_452_U316 ( .A1(fract_denorm[31]), .A2(u4_srl_452_n20), .B1(
        n3008), .B2(u4_srl_452_n24), .ZN(u4_srl_452_n287) );
  OAI221_X1 u4_srl_452_U315 ( .B1(u4_srl_452_n13), .B2(u4_srl_452_n51), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n50), .A(u4_srl_452_n287), .ZN(
        u4_srl_452_n201) );
  AOI22_X1 u4_srl_452_U314 ( .A1(fract_denorm[27]), .A2(u4_srl_452_n20), .B1(
        fract_denorm[26]), .B2(u4_srl_452_n24), .ZN(u4_srl_452_n286) );
  OAI221_X1 u4_srl_452_U313 ( .B1(u4_srl_452_n13), .B2(u4_srl_452_n46), .C1(
        u4_srl_452_n16), .C2(u4_srl_452_n48), .A(u4_srl_452_n286), .ZN(
        u4_srl_452_n196) );
  AOI22_X1 u4_srl_452_U312 ( .A1(n2551), .A2(u4_srl_452_n20), .B1(
        fract_denorm[38]), .B2(u4_srl_452_n24), .ZN(u4_srl_452_n285) );
  OAI221_X1 u4_srl_452_U311 ( .B1(u4_srl_452_n13), .B2(u4_srl_452_n60), .C1(
        u4_srl_452_n16), .C2(u4_srl_452_n59), .A(u4_srl_452_n285), .ZN(
        u4_srl_452_n195) );
  INV_X1 u4_srl_452_U310 ( .A(u4_srl_452_n195), .ZN(u4_srl_452_n239) );
  AOI22_X1 u4_srl_452_U309 ( .A1(n2483), .A2(u4_srl_452_n19), .B1(
        fract_denorm[34]), .B2(u4_srl_452_n24), .ZN(u4_srl_452_n284) );
  OAI221_X1 u4_srl_452_U308 ( .B1(u4_srl_452_n13), .B2(u4_srl_452_n54), .C1(
        u4_srl_452_n16), .C2(u4_srl_452_n56), .A(u4_srl_452_n284), .ZN(
        u4_srl_452_n221) );
  INV_X1 u4_srl_452_U307 ( .A(u4_srl_452_n221), .ZN(u4_srl_452_n199) );
  OAI22_X1 u4_srl_452_U306 ( .A1(u4_srl_452_n172), .A2(u4_srl_452_n239), .B1(
        u4_srl_452_n174), .B2(u4_srl_452_n199), .ZN(u4_srl_452_n283) );
  AOI221_X1 u4_srl_452_U305 ( .B1(u4_srl_452_n201), .B2(u4_srl_452_n143), .C1(
        u4_srl_452_n196), .C2(u4_srl_452_n164), .A(u4_srl_452_n283), .ZN(
        u4_srl_452_n166) );
  INV_X1 u4_srl_452_U304 ( .A(u4_shift_right[5]), .ZN(u4_srl_452_n281) );
  INV_X1 u4_srl_452_U303 ( .A(u4_srl_452_n134), .ZN(u4_srl_452_n81) );
  AOI22_X1 u4_srl_452_U302 ( .A1(fract_denorm[43]), .A2(u4_srl_452_n20), .B1(
        net94305), .B2(u4_srl_452_n24), .ZN(u4_srl_452_n282) );
  OAI221_X1 u4_srl_452_U301 ( .B1(u4_srl_452_n13), .B2(u4_srl_452_n61), .C1(
        u4_srl_452_n16), .C2(u4_srl_452_n64), .A(u4_srl_452_n282), .ZN(
        u4_srl_452_n193) );
  AOI22_X1 u4_srl_452_U300 ( .A1(u4_srl_452_n23), .A2(net86571), .B1(
        u4_srl_452_n19), .B2(net85391), .ZN(u4_srl_452_n127) );
  INV_X1 u4_srl_452_U299 ( .A(u4_srl_452_n127), .ZN(u4_srl_452_n194) );
  AOI22_X1 u4_srl_452_U298 ( .A1(u4_srl_452_n193), .A2(u4_srl_452_n164), .B1(
        u4_srl_452_n194), .B2(u4_srl_452_n10), .ZN(u4_srl_452_n131) );
  INV_X1 u4_srl_452_U297 ( .A(u4_srl_452_n131), .ZN(u4_srl_452_n277) );
  AOI22_X1 u4_srl_452_U296 ( .A1(net17655), .A2(u4_srl_452_n20), .B1(n5324), 
        .B2(u4_srl_452_n24), .ZN(u4_srl_452_n278) );
  OAI221_X1 u4_srl_452_U295 ( .B1(u4_srl_452_n13), .B2(u4_srl_452_n35), .C1(
        u4_srl_452_n16), .C2(u4_srl_452_n34), .A(u4_srl_452_n278), .ZN(
        u4_srl_452_n107) );
  AOI22_X1 u4_srl_452_U294 ( .A1(u4_srl_452_n81), .A2(u4_srl_452_n277), .B1(
        u4_srl_452_n83), .B2(u4_srl_452_n107), .ZN(u4_srl_452_n271) );
  AOI22_X1 u4_srl_452_U293 ( .A1(net17685), .A2(u4_srl_452_n19), .B1(net17656), 
        .B2(u4_srl_452_n24), .ZN(u4_srl_452_n275) );
  OAI221_X1 u4_srl_452_U292 ( .B1(u4_srl_452_n13), .B2(u4_srl_452_n67), .C1(
        u4_srl_452_n16), .C2(u4_srl_452_n37), .A(u4_srl_452_n275), .ZN(
        u4_srl_452_n109) );
  AOI22_X1 u4_srl_452_U291 ( .A1(u4_srl_452_n19), .A2(n3067), .B1(
        u4_srl_452_n22), .B2(fract_denorm[22]), .ZN(u4_srl_452_n274) );
  OAI221_X1 u4_srl_452_U290 ( .B1(u4_srl_452_n13), .B2(u4_srl_452_n43), .C1(
        u4_srl_452_n42), .C2(u4_srl_452_n17), .A(u4_srl_452_n274), .ZN(
        u4_srl_452_n197) );
  AOI22_X1 u4_srl_452_U289 ( .A1(net17682), .A2(u4_srl_452_n20), .B1(net17683), 
        .B2(u4_srl_452_n24), .ZN(u4_srl_452_n273) );
  OAI221_X1 u4_srl_452_U288 ( .B1(u4_srl_452_n13), .B2(u4_srl_452_n40), .C1(
        u4_srl_452_n16), .C2(u4_srl_452_n66), .A(u4_srl_452_n273), .ZN(
        u4_srl_452_n108) );
  AOI222_X1 u4_srl_452_U287 ( .A1(u4_srl_452_n75), .A2(u4_srl_452_n109), .B1(
        u4_srl_452_n77), .B2(u4_srl_452_n197), .C1(u4_srl_452_n79), .C2(
        u4_srl_452_n108), .ZN(u4_srl_452_n272) );
  OAI211_X1 u4_srl_452_U286 ( .C1(u4_srl_452_n166), .C2(u4_srl_452_n6), .A(
        u4_srl_452_n271), .B(u4_srl_452_n272), .ZN(u4_N1368) );
  AOI22_X1 u4_srl_452_U285 ( .A1(fract_denorm[32]), .A2(u4_srl_452_n20), .B1(
        fract_denorm[31]), .B2(u4_srl_452_n24), .ZN(u4_srl_452_n270) );
  OAI221_X1 u4_srl_452_U284 ( .B1(u4_srl_452_n13), .B2(u4_srl_452_n52), .C1(
        u4_srl_452_n16), .C2(u4_srl_452_n51), .A(u4_srl_452_n270), .ZN(
        u4_srl_452_n192) );
  AOI22_X1 u4_srl_452_U283 ( .A1(fract_denorm[28]), .A2(u4_srl_452_n20), .B1(
        fract_denorm[27]), .B2(u4_srl_452_n24), .ZN(u4_srl_452_n269) );
  OAI221_X1 u4_srl_452_U282 ( .B1(u4_srl_452_n14), .B2(u4_srl_452_n47), .C1(
        u4_srl_452_n16), .C2(u4_srl_452_n46), .A(u4_srl_452_n269), .ZN(
        u4_srl_452_n187) );
  AOI22_X1 u4_srl_452_U281 ( .A1(n3024), .A2(u4_srl_452_n19), .B1(n2551), .B2(
        u4_srl_452_n24), .ZN(u4_srl_452_n268) );
  OAI221_X1 u4_srl_452_U280 ( .B1(u4_srl_452_n14), .B2(u4_srl_452_n65), .C1(
        u4_srl_452_n16), .C2(u4_srl_452_n60), .A(u4_srl_452_n268), .ZN(
        u4_srl_452_n186) );
  AOI22_X1 u4_srl_452_U279 ( .A1(fract_denorm[36]), .A2(u4_srl_452_n20), .B1(
        n2483), .B2(u4_srl_452_n23), .ZN(u4_srl_452_n267) );
  OAI221_X1 u4_srl_452_U278 ( .B1(u4_srl_452_n14), .B2(u4_srl_452_n55), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n54), .A(u4_srl_452_n267), .ZN(
        u4_srl_452_n191) );
  AOI22_X1 u4_srl_452_U277 ( .A1(u4_srl_452_n142), .A2(u4_srl_452_n186), .B1(
        u4_srl_452_n141), .B2(u4_srl_452_n191), .ZN(u4_srl_452_n266) );
  INV_X1 u4_srl_452_U276 ( .A(u4_srl_452_n266), .ZN(u4_srl_452_n265) );
  AOI221_X1 u4_srl_452_U275 ( .B1(u4_srl_452_n192), .B2(u4_srl_452_n10), .C1(
        u4_srl_452_n187), .C2(u4_srl_452_n164), .A(u4_srl_452_n265), .ZN(
        u4_srl_452_n165) );
  INV_X1 u4_srl_452_U274 ( .A(u4_srl_452_n165), .ZN(u4_srl_452_n262) );
  AOI22_X1 u4_srl_452_U273 ( .A1(net17684), .A2(u4_srl_452_n19), .B1(net17685), 
        .B2(u4_srl_452_n23), .ZN(u4_srl_452_n264) );
  OAI221_X1 u4_srl_452_U272 ( .B1(u4_srl_452_n14), .B2(u4_srl_452_n38), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n67), .A(u4_srl_452_n264), .ZN(
        u4_srl_452_n100) );
  AOI22_X1 u4_srl_452_U271 ( .A1(n5326), .A2(u4_srl_452_n19), .B1(net17655), 
        .B2(u4_srl_452_n23), .ZN(u4_srl_452_n263) );
  OAI221_X1 u4_srl_452_U270 ( .B1(u4_srl_452_n14), .B2(u4_srl_452_n68), .C1(
        u4_srl_452_n16), .C2(u4_srl_452_n35), .A(u4_srl_452_n263), .ZN(
        u4_srl_452_n98) );
  AOI222_X1 u4_srl_452_U269 ( .A1(u4_srl_452_n3), .A2(u4_srl_452_n262), .B1(
        u4_srl_452_n75), .B2(u4_srl_452_n100), .C1(u4_srl_452_n83), .C2(
        u4_srl_452_n98), .ZN(u4_srl_452_n255) );
  AOI22_X1 u4_srl_452_U268 ( .A1(net17659), .A2(u4_srl_452_n20), .B1(net17682), 
        .B2(u4_srl_452_n23), .ZN(u4_srl_452_n261) );
  OAI221_X1 u4_srl_452_U267 ( .B1(u4_srl_452_n14), .B2(u4_srl_452_n41), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n40), .A(u4_srl_452_n261), .ZN(
        u4_srl_452_n99) );
  AOI22_X1 u4_srl_452_U266 ( .A1(fract_denorm[44]), .A2(u4_srl_452_n19), .B1(
        fract_denorm[43]), .B2(u4_srl_452_n23), .ZN(u4_srl_452_n260) );
  OAI221_X1 u4_srl_452_U265 ( .B1(u4_srl_452_n14), .B2(u4_srl_452_n62), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n61), .A(u4_srl_452_n260), .ZN(
        u4_srl_452_n184) );
  NAND2_X1 u4_srl_452_U264 ( .A1(net85391), .A2(u4_srl_452_n23), .ZN(
        u4_srl_452_n126) );
  INV_X1 u4_srl_452_U263 ( .A(u4_srl_452_n126), .ZN(u4_srl_452_n185) );
  MUX2_X1 u4_srl_452_U262 ( .A(u4_srl_452_n184), .B(u4_srl_452_n185), .S(
        u4_shift_right[2]), .Z(u4_srl_452_n218) );
  NAND2_X1 u4_srl_452_U261 ( .A1(u4_srl_452_n218), .A2(u4_srl_452_n259), .ZN(
        u4_srl_452_n130) );
  INV_X1 u4_srl_452_U260 ( .A(u4_srl_452_n130), .ZN(u4_srl_452_n257) );
  AOI22_X1 u4_srl_452_U259 ( .A1(u4_srl_452_n19), .A2(fract_denorm[24]), .B1(
        u4_srl_452_n22), .B2(n3067), .ZN(u4_srl_452_n258) );
  OAI221_X1 u4_srl_452_U258 ( .B1(u4_srl_452_n14), .B2(u4_srl_452_n44), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n43), .A(u4_srl_452_n258), .ZN(
        u4_srl_452_n188) );
  AOI222_X1 u4_srl_452_U257 ( .A1(u4_srl_452_n79), .A2(u4_srl_452_n99), .B1(
        u4_srl_452_n257), .B2(u4_srl_452_n81), .C1(u4_srl_452_n77), .C2(
        u4_srl_452_n188), .ZN(u4_srl_452_n256) );
  NAND2_X1 u4_srl_452_U256 ( .A1(u4_srl_452_n255), .A2(u4_srl_452_n256), .ZN(
        u4_N1369) );
  INV_X1 u4_srl_452_U255 ( .A(u4_srl_452_n206), .ZN(u4_srl_452_n181) );
  OAI22_X1 u4_srl_452_U254 ( .A1(u4_srl_452_n172), .A2(u4_srl_452_n254), .B1(
        u4_srl_452_n174), .B2(u4_srl_452_n181), .ZN(u4_srl_452_n253) );
  AOI221_X1 u4_srl_452_U253 ( .B1(u4_srl_452_n183), .B2(u4_srl_452_n10), .C1(
        u4_srl_452_n178), .C2(u4_srl_452_n164), .A(u4_srl_452_n253), .ZN(
        u4_srl_452_n163) );
  AOI22_X1 u4_srl_452_U252 ( .A1(u4_srl_452_n75), .A2(u4_srl_452_n91), .B1(
        u4_srl_452_n83), .B2(u4_srl_452_n89), .ZN(u4_srl_452_n251) );
  AND2_X1 u4_srl_452_U251 ( .A1(u4_srl_452_n135), .A2(u4_shift_right[5]), .ZN(
        u4_srl_452_n233) );
  AOI222_X1 u4_srl_452_U250 ( .A1(u4_srl_452_n79), .A2(u4_srl_452_n90), .B1(
        u4_srl_452_n233), .B2(u4_srl_452_n177), .C1(u4_srl_452_n77), .C2(
        u4_srl_452_n179), .ZN(u4_srl_452_n252) );
  OAI211_X1 u4_srl_452_U249 ( .C1(u4_srl_452_n163), .C2(u4_srl_452_n6), .A(
        u4_srl_452_n251), .B(u4_srl_452_n252), .ZN(u4_N1370) );
  AOI22_X1 u4_srl_452_U248 ( .A1(fract_denorm[34]), .A2(u4_srl_452_n146), .B1(
        fract_denorm[33]), .B2(u4_srl_452_n23), .ZN(u4_srl_452_n250) );
  OAI221_X1 u4_srl_452_U247 ( .B1(u4_srl_452_n14), .B2(u4_srl_452_n56), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n53), .A(u4_srl_452_n250), .ZN(
        u4_srl_452_n205) );
  AOI22_X1 u4_srl_452_U246 ( .A1(n3008), .A2(u4_srl_452_n20), .B1(n3006), .B2(
        u4_srl_452_n23), .ZN(u4_srl_452_n249) );
  OAI221_X1 u4_srl_452_U245 ( .B1(u4_srl_452_n14), .B2(u4_srl_452_n50), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n57), .A(u4_srl_452_n249), .ZN(
        u4_srl_452_n169) );
  AOI22_X1 u4_srl_452_U244 ( .A1(net94305), .A2(u4_srl_452_n19), .B1(net28939), 
        .B2(u4_srl_452_n23), .ZN(u4_srl_452_n248) );
  OAI221_X1 u4_srl_452_U243 ( .B1(u4_srl_452_n14), .B2(u4_srl_452_n64), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n63), .A(u4_srl_452_n248), .ZN(
        u4_srl_452_n167) );
  INV_X1 u4_srl_452_U242 ( .A(u4_srl_452_n167), .ZN(u4_srl_452_n227) );
  AOI22_X1 u4_srl_452_U241 ( .A1(fract_denorm[38]), .A2(u4_srl_452_n20), .B1(
        fract_denorm[37]), .B2(u4_srl_452_n23), .ZN(u4_srl_452_n247) );
  OAI221_X1 u4_srl_452_U240 ( .B1(u4_srl_452_n14), .B2(u4_srl_452_n59), .C1(
        u4_srl_452_n16), .C2(u4_srl_452_n58), .A(u4_srl_452_n247), .ZN(
        u4_srl_452_n202) );
  INV_X1 u4_srl_452_U239 ( .A(u4_srl_452_n202), .ZN(u4_srl_452_n173) );
  OAI22_X1 u4_srl_452_U238 ( .A1(u4_srl_452_n172), .A2(u4_srl_452_n227), .B1(
        u4_srl_452_n174), .B2(u4_srl_452_n173), .ZN(u4_srl_452_n246) );
  AOI221_X1 u4_srl_452_U237 ( .B1(u4_srl_452_n205), .B2(u4_srl_452_n143), .C1(
        u4_srl_452_n169), .C2(u4_srl_452_n164), .A(u4_srl_452_n246), .ZN(
        u4_srl_452_n162) );
  AOI22_X1 u4_srl_452_U236 ( .A1(net17683), .A2(u4_srl_452_n19), .B1(net17657), 
        .B2(u4_srl_452_n23), .ZN(u4_srl_452_n245) );
  OAI221_X1 u4_srl_452_U235 ( .B1(u4_srl_452_n14), .B2(u4_srl_452_n66), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n39), .A(u4_srl_452_n245), .ZN(
        u4_srl_452_n80) );
  AOI22_X1 u4_srl_452_U234 ( .A1(net17656), .A2(u4_srl_452_n19), .B1(net17686), 
        .B2(u4_srl_452_n23), .ZN(u4_srl_452_n244) );
  OAI221_X1 u4_srl_452_U233 ( .B1(u4_srl_452_n14), .B2(u4_srl_452_n37), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n36), .A(u4_srl_452_n244), .ZN(
        u4_srl_452_n76) );
  AOI22_X1 u4_srl_452_U232 ( .A1(u4_srl_452_n75), .A2(u4_srl_452_n80), .B1(
        u4_srl_452_n83), .B2(u4_srl_452_n76), .ZN(u4_srl_452_n240) );
  AOI22_X1 u4_srl_452_U231 ( .A1(fract_denorm[22]), .A2(u4_srl_452_n20), .B1(
        fract_denorm[21]), .B2(u4_srl_452_n23), .ZN(u4_srl_452_n243) );
  OAI221_X1 u4_srl_452_U230 ( .B1(u4_srl_452_n14), .B2(u4_srl_452_n42), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n49), .A(u4_srl_452_n243), .ZN(
        u4_srl_452_n78) );
  AOI222_X1 u4_srl_452_U229 ( .A1(u4_srl_452_n19), .A2(net86571), .B1(
        u4_srl_452_n18), .B2(net85391), .C1(u4_srl_452_n22), .C2(
        fract_denorm[45]), .ZN(u4_srl_452_n128) );
  INV_X1 u4_srl_452_U228 ( .A(u4_srl_452_n128), .ZN(u4_srl_452_n168) );
  AOI22_X1 u4_srl_452_U227 ( .A1(fract_denorm[26]), .A2(u4_srl_452_n19), .B1(
        fract_denorm[25]), .B2(u4_srl_452_n22), .ZN(u4_srl_452_n242) );
  OAI221_X1 u4_srl_452_U226 ( .B1(u4_srl_452_n12), .B2(u4_srl_452_n48), .C1(
        u4_srl_452_n144), .C2(u4_srl_452_n45), .A(u4_srl_452_n242), .ZN(
        u4_srl_452_n170) );
  AOI222_X1 u4_srl_452_U225 ( .A1(u4_srl_452_n79), .A2(u4_srl_452_n78), .B1(
        u4_srl_452_n233), .B2(u4_srl_452_n168), .C1(u4_srl_452_n77), .C2(
        u4_srl_452_n170), .ZN(u4_srl_452_n241) );
  OAI211_X1 u4_srl_452_U224 ( .C1(u4_srl_452_n162), .C2(u4_srl_452_n6), .A(
        u4_srl_452_n240), .B(u4_srl_452_n241), .ZN(u4_N1371) );
  INV_X1 u4_srl_452_U223 ( .A(u4_srl_452_n193), .ZN(u4_srl_452_n223) );
  OAI22_X1 u4_srl_452_U222 ( .A1(u4_srl_452_n172), .A2(u4_srl_452_n223), .B1(
        u4_srl_452_n174), .B2(u4_srl_452_n239), .ZN(u4_srl_452_n238) );
  AOI221_X1 u4_srl_452_U221 ( .B1(u4_srl_452_n221), .B2(u4_srl_452_n143), .C1(
        u4_srl_452_n201), .C2(u4_srl_452_n164), .A(u4_srl_452_n238), .ZN(
        u4_srl_452_n153) );
  AOI22_X1 u4_srl_452_U220 ( .A1(u4_srl_452_n75), .A2(u4_srl_452_n108), .B1(
        u4_srl_452_n83), .B2(u4_srl_452_n109), .ZN(u4_srl_452_n236) );
  AOI222_X1 u4_srl_452_U219 ( .A1(u4_srl_452_n79), .A2(u4_srl_452_n197), .B1(
        u4_srl_452_n233), .B2(u4_srl_452_n194), .C1(u4_srl_452_n77), .C2(
        u4_srl_452_n196), .ZN(u4_srl_452_n237) );
  OAI211_X1 u4_srl_452_U218 ( .C1(u4_srl_452_n153), .C2(u4_srl_452_n6), .A(
        u4_srl_452_n236), .B(u4_srl_452_n237), .ZN(u4_N1372) );
  AOI22_X1 u4_srl_452_U217 ( .A1(u4_srl_452_n142), .A2(u4_srl_452_n184), .B1(
        u4_srl_452_n141), .B2(u4_srl_452_n186), .ZN(u4_srl_452_n235) );
  INV_X1 u4_srl_452_U216 ( .A(u4_srl_452_n235), .ZN(u4_srl_452_n234) );
  AOI221_X1 u4_srl_452_U215 ( .B1(u4_srl_452_n191), .B2(u4_srl_452_n10), .C1(
        u4_srl_452_n192), .C2(u4_srl_452_n164), .A(u4_srl_452_n234), .ZN(
        u4_srl_452_n151) );
  AOI22_X1 u4_srl_452_U214 ( .A1(u4_srl_452_n75), .A2(u4_srl_452_n99), .B1(
        u4_srl_452_n83), .B2(u4_srl_452_n100), .ZN(u4_srl_452_n231) );
  AOI222_X1 u4_srl_452_U213 ( .A1(u4_srl_452_n79), .A2(u4_srl_452_n188), .B1(
        u4_srl_452_n233), .B2(u4_srl_452_n185), .C1(u4_srl_452_n77), .C2(
        u4_srl_452_n187), .ZN(u4_srl_452_n232) );
  OAI211_X1 u4_srl_452_U212 ( .C1(u4_srl_452_n151), .C2(u4_srl_452_n6), .A(
        u4_srl_452_n231), .B(u4_srl_452_n232), .ZN(u4_N1373) );
  OAI22_X1 u4_srl_452_U211 ( .A1(u4_srl_452_n230), .A2(u4_srl_452_n9), .B1(
        u4_srl_452_n150), .B2(u4_srl_452_n6), .ZN(u4_N1374) );
  AOI22_X1 u4_srl_452_U210 ( .A1(u4_srl_452_n142), .A2(u4_srl_452_n169), .B1(
        u4_srl_452_n141), .B2(u4_srl_452_n170), .ZN(u4_srl_452_n229) );
  INV_X1 u4_srl_452_U209 ( .A(u4_srl_452_n229), .ZN(u4_srl_452_n228) );
  AOI221_X1 u4_srl_452_U208 ( .B1(u4_srl_452_n78), .B2(u4_srl_452_n10), .C1(
        u4_srl_452_n80), .C2(u4_srl_452_n164), .A(u4_srl_452_n228), .ZN(
        u4_srl_452_n214) );
  OAI22_X1 u4_srl_452_U207 ( .A1(u4_srl_452_n172), .A2(u4_srl_452_n128), .B1(
        u4_srl_452_n174), .B2(u4_srl_452_n227), .ZN(u4_srl_452_n226) );
  AOI221_X1 u4_srl_452_U206 ( .B1(u4_srl_452_n202), .B2(u4_srl_452_n10), .C1(
        u4_srl_452_n205), .C2(u4_srl_452_n164), .A(u4_srl_452_n226), .ZN(
        u4_srl_452_n149) );
  OAI22_X1 u4_srl_452_U205 ( .A1(u4_srl_452_n214), .A2(u4_srl_452_n9), .B1(
        u4_srl_452_n149), .B2(u4_srl_452_n6), .ZN(u4_N1375) );
  AOI22_X1 u4_srl_452_U204 ( .A1(u4_srl_452_n142), .A2(u4_srl_452_n201), .B1(
        u4_srl_452_n141), .B2(u4_srl_452_n196), .ZN(u4_srl_452_n225) );
  INV_X1 u4_srl_452_U203 ( .A(u4_srl_452_n225), .ZN(u4_srl_452_n224) );
  AOI221_X1 u4_srl_452_U202 ( .B1(u4_srl_452_n197), .B2(u4_srl_452_n10), .C1(
        u4_srl_452_n108), .C2(u4_srl_452_n164), .A(u4_srl_452_n224), .ZN(
        u4_srl_452_n159) );
  OAI22_X1 u4_srl_452_U201 ( .A1(u4_srl_452_n172), .A2(u4_srl_452_n127), .B1(
        u4_srl_452_n174), .B2(u4_srl_452_n223), .ZN(u4_srl_452_n222) );
  AOI221_X1 u4_srl_452_U200 ( .B1(u4_srl_452_n195), .B2(u4_srl_452_n10), .C1(
        u4_srl_452_n221), .C2(u4_srl_452_n164), .A(u4_srl_452_n222), .ZN(
        u4_srl_452_n148) );
  OAI22_X1 u4_srl_452_U199 ( .A1(u4_srl_452_n159), .A2(u4_srl_452_n9), .B1(
        u4_srl_452_n148), .B2(u4_srl_452_n6), .ZN(u4_N1376) );
  AOI22_X1 u4_srl_452_U198 ( .A1(u4_srl_452_n142), .A2(u4_srl_452_n192), .B1(
        u4_srl_452_n141), .B2(u4_srl_452_n187), .ZN(u4_srl_452_n220) );
  INV_X1 u4_srl_452_U197 ( .A(u4_srl_452_n220), .ZN(u4_srl_452_n219) );
  AOI221_X1 u4_srl_452_U196 ( .B1(u4_srl_452_n188), .B2(u4_srl_452_n10), .C1(
        u4_srl_452_n99), .C2(u4_srl_452_n164), .A(u4_srl_452_n219), .ZN(
        u4_srl_452_n140) );
  AOI222_X1 u4_srl_452_U195 ( .A1(u4_srl_452_n191), .A2(u4_srl_452_n164), .B1(
        u4_srl_452_n186), .B2(u4_srl_452_n143), .C1(u4_srl_452_n218), .C2(
        u4_shift_right[3]), .ZN(u4_srl_452_n133) );
  OAI22_X1 u4_srl_452_U194 ( .A1(u4_srl_452_n140), .A2(u4_srl_452_n9), .B1(
        u4_srl_452_n133), .B2(u4_srl_452_n6), .ZN(u4_N1377) );
  AOI22_X1 u4_srl_452_U193 ( .A1(net17694), .A2(u4_srl_452_n19), .B1(net17695), 
        .B2(u4_srl_452_n22), .ZN(u4_srl_452_n217) );
  OAI221_X1 u4_srl_452_U192 ( .B1(u4_srl_452_n14), .B2(u4_srl_452_n28), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n71), .A(u4_srl_452_n217), .ZN(
        u4_srl_452_n210) );
  AOI22_X1 u4_srl_452_U191 ( .A1(n5324), .A2(u4_srl_452_n19), .B1(n2980), .B2(
        u4_srl_452_n22), .ZN(u4_srl_452_n216) );
  OAI221_X1 u4_srl_452_U190 ( .B1(u4_srl_452_n14), .B2(u4_srl_452_n34), .C1(
        u4_srl_452_n16), .C2(u4_srl_452_n69), .A(u4_srl_452_n216), .ZN(
        u4_srl_452_n84) );
  AOI22_X1 u4_srl_452_U189 ( .A1(net17654), .A2(u4_srl_452_n19), .B1(net17692), 
        .B2(u4_srl_452_n22), .ZN(u4_srl_452_n215) );
  OAI221_X1 u4_srl_452_U188 ( .B1(u4_srl_452_n14), .B2(u4_srl_452_n31), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n30), .A(u4_srl_452_n215), .ZN(
        u4_srl_452_n117) );
  AOI222_X1 u4_srl_452_U187 ( .A1(u4_srl_452_n84), .A2(u4_srl_452_n141), .B1(
        u4_srl_452_n76), .B2(u4_srl_452_n142), .C1(u4_srl_452_n117), .C2(
        u4_srl_452_n10), .ZN(u4_srl_452_n213) );
  MUX2_X1 u4_srl_452_U186 ( .A(u4_srl_452_n213), .B(u4_srl_452_n214), .S(
        u4_shift_right[4]), .Z(u4_srl_452_n212) );
  INV_X1 u4_srl_452_U185 ( .A(u4_srl_452_n212), .ZN(u4_srl_452_n211) );
  AOI21_X1 u4_srl_452_U184 ( .B1(u4_srl_452_n135), .B2(u4_srl_452_n210), .A(
        u4_srl_452_n211), .ZN(u4_srl_452_n209) );
  OAI22_X1 u4_srl_452_U183 ( .A1(u4_shift_right[5]), .A2(u4_srl_452_n209), 
        .B1(u4_srl_452_n149), .B2(u4_srl_452_n134), .ZN(u4_N1359) );
  AOI22_X1 u4_srl_452_U182 ( .A1(u4_srl_452_n142), .A2(u4_srl_452_n183), .B1(
        u4_srl_452_n141), .B2(u4_srl_452_n178), .ZN(u4_srl_452_n208) );
  INV_X1 u4_srl_452_U181 ( .A(u4_srl_452_n208), .ZN(u4_srl_452_n207) );
  AOI221_X1 u4_srl_452_U180 ( .B1(u4_srl_452_n179), .B2(u4_srl_452_n10), .C1(
        u4_srl_452_n90), .C2(u4_srl_452_n164), .A(u4_srl_452_n207), .ZN(
        u4_srl_452_n119) );
  AOI222_X1 u4_srl_452_U179 ( .A1(u4_srl_452_n176), .A2(u4_srl_452_n10), .B1(
        u4_srl_452_n177), .B2(u4_srl_452_n141), .C1(u4_srl_452_n206), .C2(
        u4_srl_452_n164), .ZN(u4_srl_452_n124) );
  OAI22_X1 u4_srl_452_U178 ( .A1(u4_srl_452_n119), .A2(u4_srl_452_n8), .B1(
        u4_srl_452_n124), .B2(u4_srl_452_n6), .ZN(u4_N1378) );
  INV_X1 u4_srl_452_U177 ( .A(u4_srl_452_n205), .ZN(u4_srl_452_n175) );
  INV_X1 u4_srl_452_U176 ( .A(u4_srl_452_n169), .ZN(u4_srl_452_n204) );
  OAI22_X1 u4_srl_452_U175 ( .A1(u4_srl_452_n172), .A2(u4_srl_452_n175), .B1(
        u4_srl_452_n174), .B2(u4_srl_452_n204), .ZN(u4_srl_452_n203) );
  AOI221_X1 u4_srl_452_U174 ( .B1(u4_srl_452_n170), .B2(u4_srl_452_n10), .C1(
        u4_srl_452_n78), .C2(u4_srl_452_n164), .A(u4_srl_452_n203), .ZN(
        u4_srl_452_n113) );
  AOI222_X1 u4_srl_452_U173 ( .A1(u4_srl_452_n167), .A2(u4_srl_452_n10), .B1(
        u4_srl_452_n168), .B2(u4_srl_452_n141), .C1(u4_srl_452_n202), .C2(
        u4_srl_452_n164), .ZN(u4_srl_452_n118) );
  OAI22_X1 u4_srl_452_U172 ( .A1(u4_srl_452_n113), .A2(u4_srl_452_n9), .B1(
        u4_srl_452_n118), .B2(u4_srl_452_n6), .ZN(u4_N1379) );
  INV_X1 u4_srl_452_U171 ( .A(u4_srl_452_n201), .ZN(u4_srl_452_n200) );
  OAI22_X1 u4_srl_452_U170 ( .A1(u4_srl_452_n172), .A2(u4_srl_452_n199), .B1(
        u4_srl_452_n174), .B2(u4_srl_452_n200), .ZN(u4_srl_452_n198) );
  AOI221_X1 u4_srl_452_U169 ( .B1(u4_srl_452_n196), .B2(u4_srl_452_n10), .C1(
        u4_srl_452_n197), .C2(u4_srl_452_n164), .A(u4_srl_452_n198), .ZN(
        u4_srl_452_n104) );
  AOI222_X1 u4_srl_452_U168 ( .A1(u4_srl_452_n193), .A2(u4_srl_452_n10), .B1(
        u4_srl_452_n194), .B2(u4_srl_452_n141), .C1(u4_srl_452_n195), .C2(
        u4_srl_452_n164), .ZN(u4_srl_452_n112) );
  OAI22_X1 u4_srl_452_U167 ( .A1(u4_srl_452_n104), .A2(u4_srl_452_n8), .B1(
        u4_srl_452_n112), .B2(u4_srl_452_n7), .ZN(u4_N1380) );
  AOI22_X1 u4_srl_452_U166 ( .A1(u4_srl_452_n142), .A2(u4_srl_452_n191), .B1(
        u4_srl_452_n141), .B2(u4_srl_452_n192), .ZN(u4_srl_452_n190) );
  INV_X1 u4_srl_452_U165 ( .A(u4_srl_452_n190), .ZN(u4_srl_452_n189) );
  AOI221_X1 u4_srl_452_U164 ( .B1(u4_srl_452_n187), .B2(u4_srl_452_n10), .C1(
        u4_srl_452_n188), .C2(u4_srl_452_n164), .A(u4_srl_452_n189), .ZN(
        u4_srl_452_n95) );
  AOI222_X1 u4_srl_452_U163 ( .A1(u4_srl_452_n184), .A2(u4_srl_452_n10), .B1(
        u4_srl_452_n141), .B2(u4_srl_452_n185), .C1(u4_srl_452_n186), .C2(
        u4_srl_452_n164), .ZN(u4_srl_452_n103) );
  OAI22_X1 u4_srl_452_U162 ( .A1(u4_srl_452_n95), .A2(u4_srl_452_n8), .B1(
        u4_srl_452_n103), .B2(u4_srl_452_n6), .ZN(u4_N1381) );
  INV_X1 u4_srl_452_U161 ( .A(u4_srl_452_n183), .ZN(u4_srl_452_n182) );
  OAI22_X1 u4_srl_452_U160 ( .A1(u4_srl_452_n172), .A2(u4_srl_452_n181), .B1(
        u4_srl_452_n174), .B2(u4_srl_452_n182), .ZN(u4_srl_452_n180) );
  AOI221_X1 u4_srl_452_U159 ( .B1(u4_srl_452_n178), .B2(u4_srl_452_n10), .C1(
        u4_srl_452_n179), .C2(u4_srl_452_n164), .A(u4_srl_452_n180), .ZN(
        u4_srl_452_n86) );
  AOI22_X1 u4_srl_452_U158 ( .A1(u4_srl_452_n176), .A2(u4_srl_452_n164), .B1(
        u4_srl_452_n177), .B2(u4_srl_452_n10), .ZN(u4_srl_452_n94) );
  OAI22_X1 u4_srl_452_U157 ( .A1(u4_srl_452_n86), .A2(u4_srl_452_n8), .B1(
        u4_srl_452_n94), .B2(u4_srl_452_n6), .ZN(u4_N1382) );
  OAI22_X1 u4_srl_452_U156 ( .A1(u4_srl_452_n172), .A2(u4_srl_452_n173), .B1(
        u4_srl_452_n174), .B2(u4_srl_452_n175), .ZN(u4_srl_452_n171) );
  AOI221_X1 u4_srl_452_U155 ( .B1(u4_srl_452_n169), .B2(u4_srl_452_n10), .C1(
        u4_srl_452_n170), .C2(u4_srl_452_n164), .A(u4_srl_452_n171), .ZN(
        u4_srl_452_n72) );
  AOI22_X1 u4_srl_452_U154 ( .A1(u4_srl_452_n167), .A2(u4_srl_452_n164), .B1(
        u4_srl_452_n168), .B2(u4_srl_452_n143), .ZN(u4_srl_452_n85) );
  OAI22_X1 u4_srl_452_U153 ( .A1(u4_srl_452_n72), .A2(u4_srl_452_n8), .B1(
        u4_srl_452_n85), .B2(u4_srl_452_n6), .ZN(u4_N1383) );
  OAI22_X1 u4_srl_452_U152 ( .A1(u4_srl_452_n166), .A2(u4_srl_452_n8), .B1(
        u4_srl_452_n131), .B2(u4_srl_452_n6), .ZN(u4_N1384) );
  OAI22_X1 u4_srl_452_U151 ( .A1(u4_srl_452_n165), .A2(u4_srl_452_n8), .B1(
        u4_srl_452_n7), .B2(u4_srl_452_n130), .ZN(u4_N1385) );
  NAND2_X1 u4_srl_452_U150 ( .A1(u4_srl_452_n3), .A2(u4_srl_452_n164), .ZN(
        u4_srl_452_n152) );
  OAI22_X1 u4_srl_452_U149 ( .A1(u4_srl_452_n163), .A2(u4_srl_452_n8), .B1(
        u4_srl_452_n129), .B2(u4_srl_452_n152), .ZN(u4_N1386) );
  OAI22_X1 u4_srl_452_U148 ( .A1(u4_srl_452_n162), .A2(u4_srl_452_n8), .B1(
        u4_srl_452_n128), .B2(u4_srl_452_n152), .ZN(u4_N1387) );
  AOI22_X1 u4_srl_452_U147 ( .A1(net17653), .A2(u4_srl_452_n19), .B1(net17694), 
        .B2(u4_srl_452_n22), .ZN(u4_srl_452_n161) );
  OAI221_X1 u4_srl_452_U146 ( .B1(u4_srl_452_n14), .B2(u4_srl_452_n29), .C1(
        u4_srl_452_n144), .C2(u4_srl_452_n28), .A(u4_srl_452_n161), .ZN(
        u4_srl_452_n155) );
  AOI22_X1 u4_srl_452_U145 ( .A1(n5323), .A2(u4_srl_452_n19), .B1(net17654), 
        .B2(u4_srl_452_n22), .ZN(u4_srl_452_n160) );
  OAI221_X1 u4_srl_452_U144 ( .B1(u4_srl_452_n14), .B2(u4_srl_452_n33), .C1(
        u4_srl_452_n17), .C2(u4_srl_452_n31), .A(u4_srl_452_n160), .ZN(
        u4_srl_452_n111) );
  AOI222_X1 u4_srl_452_U143 ( .A1(u4_srl_452_n107), .A2(u4_srl_452_n141), .B1(
        u4_srl_452_n109), .B2(u4_srl_452_n142), .C1(u4_srl_452_n111), .C2(
        u4_srl_452_n10), .ZN(u4_srl_452_n158) );
  MUX2_X1 u4_srl_452_U142 ( .A(u4_srl_452_n158), .B(u4_srl_452_n159), .S(
        u4_shift_right[4]), .Z(u4_srl_452_n157) );
  INV_X1 u4_srl_452_U141 ( .A(u4_srl_452_n157), .ZN(u4_srl_452_n156) );
  AOI21_X1 u4_srl_452_U140 ( .B1(u4_srl_452_n135), .B2(u4_srl_452_n155), .A(
        u4_srl_452_n156), .ZN(u4_srl_452_n154) );
  OAI22_X1 u4_srl_452_U139 ( .A1(u4_shift_right[5]), .A2(u4_srl_452_n154), 
        .B1(u4_srl_452_n148), .B2(u4_srl_452_n134), .ZN(u4_N1360) );
  OAI22_X1 u4_srl_452_U138 ( .A1(u4_srl_452_n153), .A2(u4_srl_452_n8), .B1(
        u4_srl_452_n127), .B2(u4_srl_452_n152), .ZN(u4_N1388) );
  OAI22_X1 u4_srl_452_U137 ( .A1(u4_srl_452_n151), .A2(u4_srl_452_n8), .B1(
        u4_srl_452_n126), .B2(u4_srl_452_n152), .ZN(u4_N1389) );
  NOR2_X1 u4_srl_452_U136 ( .A1(u4_srl_452_n150), .A2(u4_srl_452_n9), .ZN(
        u4_N1390) );
  NOR2_X1 u4_srl_452_U135 ( .A1(u4_srl_452_n149), .A2(u4_srl_452_n9), .ZN(
        u4_N1391) );
  NOR2_X1 u4_srl_452_U134 ( .A1(u4_srl_452_n148), .A2(u4_srl_452_n8), .ZN(
        u4_N1392) );
  NOR2_X1 u4_srl_452_U133 ( .A1(u4_srl_452_n133), .A2(u4_srl_452_n8), .ZN(
        u4_N1393) );
  NOR2_X1 u4_srl_452_U132 ( .A1(u4_srl_452_n124), .A2(u4_srl_452_n8), .ZN(
        u4_N1394) );
  NOR2_X1 u4_srl_452_U131 ( .A1(u4_srl_452_n118), .A2(u4_srl_452_n8), .ZN(
        u4_N1395) );
  NOR2_X1 u4_srl_452_U130 ( .A1(u4_srl_452_n112), .A2(u4_srl_452_n8), .ZN(
        u4_N1396) );
  NOR2_X1 u4_srl_452_U129 ( .A1(u4_srl_452_n103), .A2(u4_srl_452_n8), .ZN(
        u4_N1397) );
  AOI22_X1 u4_srl_452_U128 ( .A1(net17693), .A2(u4_srl_452_n19), .B1(net17653), 
        .B2(u4_srl_452_n22), .ZN(u4_srl_452_n147) );
  OAI221_X1 u4_srl_452_U127 ( .B1(u4_srl_452_n14), .B2(u4_srl_452_n70), .C1(
        u4_srl_452_n144), .C2(u4_srl_452_n29), .A(u4_srl_452_n147), .ZN(
        u4_srl_452_n136) );
  AOI22_X1 u4_srl_452_U126 ( .A1(net17690), .A2(u4_srl_452_n19), .B1(n5323), 
        .B2(u4_srl_452_n24), .ZN(u4_srl_452_n145) );
  OAI221_X1 u4_srl_452_U125 ( .B1(u4_srl_452_n13), .B2(u4_srl_452_n32), .C1(
        u4_srl_452_n16), .C2(u4_srl_452_n33), .A(u4_srl_452_n145), .ZN(
        u4_srl_452_n102) );
  AOI222_X1 u4_srl_452_U124 ( .A1(u4_srl_452_n98), .A2(u4_srl_452_n141), .B1(
        u4_srl_452_n100), .B2(u4_srl_452_n142), .C1(u4_srl_452_n102), .C2(
        u4_srl_452_n10), .ZN(u4_srl_452_n139) );
  MUX2_X1 u4_srl_452_U123 ( .A(u4_srl_452_n139), .B(u4_srl_452_n140), .S(
        u4_shift_right[4]), .Z(u4_srl_452_n138) );
  INV_X1 u4_srl_452_U122 ( .A(u4_srl_452_n138), .ZN(u4_srl_452_n137) );
  AOI21_X1 u4_srl_452_U121 ( .B1(u4_srl_452_n135), .B2(u4_srl_452_n136), .A(
        u4_srl_452_n137), .ZN(u4_srl_452_n132) );
  OAI22_X1 u4_srl_452_U120 ( .A1(u4_shift_right[5]), .A2(u4_srl_452_n132), 
        .B1(u4_srl_452_n133), .B2(u4_srl_452_n134), .ZN(u4_N1361) );
  NOR2_X1 u4_srl_452_U119 ( .A1(u4_srl_452_n94), .A2(u4_srl_452_n8), .ZN(
        u4_N1398) );
  NOR2_X1 u4_srl_452_U118 ( .A1(u4_srl_452_n85), .A2(u4_srl_452_n8), .ZN(
        u4_N1399) );
  NOR2_X1 u4_srl_452_U117 ( .A1(u4_srl_452_n131), .A2(u4_srl_452_n8), .ZN(
        u4_N1400) );
  NOR2_X1 u4_srl_452_U116 ( .A1(u4_srl_452_n9), .A2(u4_srl_452_n130), .ZN(
        u4_N1401) );
  INV_X1 u4_srl_452_U115 ( .A(u4_srl_452_n83), .ZN(u4_srl_452_n125) );
  NOR2_X1 u4_srl_452_U114 ( .A1(u4_srl_452_n129), .A2(u4_srl_452_n125), .ZN(
        u4_N1402) );
  NOR2_X1 u4_srl_452_U113 ( .A1(u4_srl_452_n128), .A2(u4_srl_452_n125), .ZN(
        u4_N1403) );
  NOR2_X1 u4_srl_452_U112 ( .A1(u4_srl_452_n127), .A2(u4_srl_452_n125), .ZN(
        u4_N1404) );
  NOR2_X1 u4_srl_452_U111 ( .A1(u4_srl_452_n125), .A2(u4_srl_452_n126), .ZN(
        u4_N1405) );
  INV_X1 u4_srl_452_U110 ( .A(u4_srl_452_n124), .ZN(u4_srl_452_n122) );
  AOI22_X1 u4_srl_452_U109 ( .A1(u4_srl_452_n81), .A2(u4_srl_452_n122), .B1(
        u4_srl_452_n83), .B2(u4_srl_452_n123), .ZN(u4_srl_452_n120) );
  AOI222_X1 u4_srl_452_U108 ( .A1(u4_srl_452_n75), .A2(u4_srl_452_n93), .B1(
        u4_srl_452_n77), .B2(u4_srl_452_n91), .C1(u4_srl_452_n79), .C2(
        u4_srl_452_n89), .ZN(u4_srl_452_n121) );
  OAI211_X1 u4_srl_452_U107 ( .C1(u4_srl_452_n119), .C2(u4_srl_452_n6), .A(
        u4_srl_452_n120), .B(u4_srl_452_n121), .ZN(u4_N1362) );
  INV_X1 u4_srl_452_U106 ( .A(u4_srl_452_n118), .ZN(u4_srl_452_n116) );
  AOI22_X1 u4_srl_452_U105 ( .A1(u4_srl_452_n81), .A2(u4_srl_452_n116), .B1(
        u4_srl_452_n83), .B2(u4_srl_452_n117), .ZN(u4_srl_452_n114) );
  AOI222_X1 u4_srl_452_U104 ( .A1(u4_srl_452_n75), .A2(u4_srl_452_n84), .B1(
        u4_srl_452_n77), .B2(u4_srl_452_n80), .C1(u4_srl_452_n79), .C2(
        u4_srl_452_n76), .ZN(u4_srl_452_n115) );
  OAI211_X1 u4_srl_452_U103 ( .C1(u4_srl_452_n113), .C2(u4_srl_452_n6), .A(
        u4_srl_452_n114), .B(u4_srl_452_n115), .ZN(u4_N1363) );
  INV_X1 u4_srl_452_U102 ( .A(u4_srl_452_n112), .ZN(u4_srl_452_n110) );
  AOI22_X1 u4_srl_452_U101 ( .A1(u4_srl_452_n81), .A2(u4_srl_452_n110), .B1(
        u4_srl_452_n83), .B2(u4_srl_452_n111), .ZN(u4_srl_452_n105) );
  AOI222_X1 u4_srl_452_U100 ( .A1(u4_srl_452_n75), .A2(u4_srl_452_n107), .B1(
        u4_srl_452_n77), .B2(u4_srl_452_n108), .C1(u4_srl_452_n79), .C2(
        u4_srl_452_n109), .ZN(u4_srl_452_n106) );
  OAI211_X1 u4_srl_452_U99 ( .C1(u4_srl_452_n104), .C2(u4_srl_452_n6), .A(
        u4_srl_452_n105), .B(u4_srl_452_n106), .ZN(u4_N1364) );
  INV_X1 u4_srl_452_U98 ( .A(u4_srl_452_n103), .ZN(u4_srl_452_n101) );
  AOI22_X1 u4_srl_452_U97 ( .A1(u4_srl_452_n81), .A2(u4_srl_452_n101), .B1(
        u4_srl_452_n83), .B2(u4_srl_452_n102), .ZN(u4_srl_452_n96) );
  AOI222_X1 u4_srl_452_U96 ( .A1(u4_srl_452_n75), .A2(u4_srl_452_n98), .B1(
        u4_srl_452_n77), .B2(u4_srl_452_n99), .C1(u4_srl_452_n79), .C2(
        u4_srl_452_n100), .ZN(u4_srl_452_n97) );
  OAI211_X1 u4_srl_452_U95 ( .C1(u4_srl_452_n95), .C2(u4_srl_452_n6), .A(
        u4_srl_452_n96), .B(u4_srl_452_n97), .ZN(u4_N1365) );
  INV_X1 u4_srl_452_U94 ( .A(u4_srl_452_n94), .ZN(u4_srl_452_n92) );
  AOI22_X1 u4_srl_452_U93 ( .A1(u4_srl_452_n81), .A2(u4_srl_452_n92), .B1(
        u4_srl_452_n83), .B2(u4_srl_452_n93), .ZN(u4_srl_452_n87) );
  AOI222_X1 u4_srl_452_U92 ( .A1(u4_srl_452_n75), .A2(u4_srl_452_n89), .B1(
        u4_srl_452_n77), .B2(u4_srl_452_n90), .C1(u4_srl_452_n79), .C2(
        u4_srl_452_n91), .ZN(u4_srl_452_n88) );
  OAI211_X1 u4_srl_452_U91 ( .C1(u4_srl_452_n86), .C2(u4_srl_452_n6), .A(
        u4_srl_452_n87), .B(u4_srl_452_n88), .ZN(u4_N1366) );
  INV_X1 u4_srl_452_U90 ( .A(u4_srl_452_n85), .ZN(u4_srl_452_n82) );
  AOI22_X1 u4_srl_452_U89 ( .A1(u4_srl_452_n81), .A2(u4_srl_452_n82), .B1(
        u4_srl_452_n83), .B2(u4_srl_452_n84), .ZN(u4_srl_452_n73) );
  AOI222_X1 u4_srl_452_U88 ( .A1(u4_srl_452_n75), .A2(u4_srl_452_n76), .B1(
        u4_srl_452_n77), .B2(u4_srl_452_n78), .C1(u4_srl_452_n79), .C2(
        u4_srl_452_n80), .ZN(u4_srl_452_n74) );
  OAI211_X1 u4_srl_452_U87 ( .C1(u4_srl_452_n72), .C2(u4_srl_452_n6), .A(
        u4_srl_452_n73), .B(u4_srl_452_n74), .ZN(u4_N1367) );
  INV_X4 u4_srl_452_U86 ( .A(net17653), .ZN(u4_srl_452_n71) );
  INV_X4 u4_srl_452_U85 ( .A(net17656), .ZN(u4_srl_452_n68) );
  INV_X4 u4_srl_452_U84 ( .A(net17657), .ZN(u4_srl_452_n67) );
  INV_X4 u4_srl_452_U83 ( .A(net17659), .ZN(u4_srl_452_n66) );
  INV_X4 u4_srl_452_U82 ( .A(net86571), .ZN(u4_srl_452_n62) );
  INV_X4 u4_srl_452_U81 ( .A(net28939), .ZN(u4_srl_452_n60) );
  INV_X4 u4_srl_452_U80 ( .A(fract_denorm[37]), .ZN(u4_srl_452_n54) );
  INV_X4 u4_srl_452_U79 ( .A(fract_denorm[33]), .ZN(u4_srl_452_n51) );
  INV_X4 u4_srl_452_U78 ( .A(fract_denorm[26]), .ZN(u4_srl_452_n44) );
  INV_X4 u4_srl_452_U77 ( .A(fract_denorm[25]), .ZN(u4_srl_452_n43) );
  INV_X4 u4_srl_452_U76 ( .A(fract_denorm[24]), .ZN(u4_srl_452_n42) );
  INV_X4 u4_srl_452_U75 ( .A(net17682), .ZN(u4_srl_452_n39) );
  INV_X4 u4_srl_452_U74 ( .A(net17683), .ZN(u4_srl_452_n38) );
  INV_X4 u4_srl_452_U73 ( .A(net17684), .ZN(u4_srl_452_n37) );
  INV_X4 u4_srl_452_U72 ( .A(net17690), .ZN(u4_srl_452_n31) );
  INV_X4 u4_srl_452_U71 ( .A(n5323), .ZN(u4_srl_452_n30) );
  INV_X4 u4_srl_452_U70 ( .A(net17692), .ZN(u4_srl_452_n29) );
  INV_X4 u4_srl_452_U69 ( .A(net17693), .ZN(u4_srl_452_n28) );
  INV_X4 u4_srl_452_U68 ( .A(net17694), .ZN(u4_srl_452_n27) );
  NAND2_X4 u4_srl_452_U67 ( .A1(u4_shift_right[3]), .A2(u4_srl_452_n306), .ZN(
        u4_srl_452_n174) );
  INV_X16 u4_srl_452_U66 ( .A(u4_srl_452_n174), .ZN(u4_srl_452_n141) );
  NAND2_X4 u4_srl_452_U65 ( .A1(u4_shift_right[3]), .A2(u4_shift_right[2]), 
        .ZN(u4_srl_452_n172) );
  INV_X16 u4_srl_452_U64 ( .A(u4_srl_452_n172), .ZN(u4_srl_452_n142) );
  NOR2_X4 u4_srl_452_U63 ( .A1(u4_srl_452_n279), .A2(u4_srl_452_n8), .ZN(
        u4_srl_452_n83) );
  NOR2_X4 u4_srl_452_U62 ( .A1(u4_srl_452_n276), .A2(u4_srl_452_n9), .ZN(
        u4_srl_452_n75) );
  NOR2_X4 u4_srl_452_U61 ( .A1(u4_srl_452_n9), .A2(u4_srl_452_n172), .ZN(
        u4_srl_452_n77) );
  NOR2_X4 u4_srl_452_U60 ( .A1(u4_srl_452_n174), .A2(u4_srl_452_n9), .ZN(
        u4_srl_452_n79) );
  INV_X1 u4_srl_452_U59 ( .A(n2551), .ZN(u4_srl_452_n58) );
  INV_X1 u4_srl_452_U58 ( .A(n3067), .ZN(u4_srl_452_n49) );
  INV_X1 u4_srl_452_U57 ( .A(n3024), .ZN(u4_srl_452_n59) );
  INV_X1 u4_srl_452_U56 ( .A(fract_denorm[32]), .ZN(u4_srl_452_n50) );
  INV_X1 u4_srl_452_U55 ( .A(n2980), .ZN(u4_srl_452_n33) );
  INV_X1 u4_srl_452_U54 ( .A(n2483), .ZN(u4_srl_452_n53) );
  INV_X2 u4_srl_452_U53 ( .A(net17686), .ZN(u4_srl_452_n35) );
  INV_X2 u4_srl_452_U52 ( .A(net17654), .ZN(u4_srl_452_n70) );
  INV_X1 u4_srl_452_U51 ( .A(fract_denorm[44]), .ZN(u4_srl_452_n64) );
  INV_X2 u4_srl_452_U50 ( .A(net17685), .ZN(u4_srl_452_n36) );
  INV_X1 u4_srl_452_U49 ( .A(n3008), .ZN(u4_srl_452_n47) );
  INV_X2 u4_srl_452_U48 ( .A(fract_denorm[21]), .ZN(u4_srl_452_n40) );
  INV_X2 u4_srl_452_U47 ( .A(n3006), .ZN(u4_srl_452_n46) );
  INV_X1 u4_srl_452_U46 ( .A(net94305), .ZN(u4_srl_452_n65) );
  INV_X1 u4_srl_452_U45 ( .A(fract_denorm[22]), .ZN(u4_srl_452_n41) );
  INV_X1 u4_srl_452_U44 ( .A(n5326), .ZN(u4_srl_452_n34) );
  INV_X2 u4_srl_452_U43 ( .A(fract_denorm[27]), .ZN(u4_srl_452_n45) );
  INV_X1 u4_srl_452_U42 ( .A(fract_denorm[28]), .ZN(u4_srl_452_n48) );
  INV_X2 u4_srl_452_U41 ( .A(fract_denorm[34]), .ZN(u4_srl_452_n52) );
  INV_X4 u4_srl_452_U40 ( .A(u4_shift_right[0]), .ZN(u4_srl_452_n309) );
  INV_X1 u4_srl_452_U39 ( .A(net85391), .ZN(u4_srl_452_n26) );
  INV_X1 u4_srl_452_U38 ( .A(u4_srl_452_n3), .ZN(u4_srl_452_n7) );
  INV_X4 u4_srl_452_U37 ( .A(u4_srl_452_n1), .ZN(u4_srl_452_n8) );
  INV_X16 u4_srl_452_U36 ( .A(u4_srl_452_n23), .ZN(u4_srl_452_n25) );
  INV_X4 u4_srl_452_U35 ( .A(u4_srl_452_n11), .ZN(u4_srl_452_n10) );
  INV_X4 u4_srl_452_U34 ( .A(u4_srl_452_n143), .ZN(u4_srl_452_n11) );
  AND2_X4 u4_srl_452_U33 ( .A1(u4_shift_right[1]), .A2(u4_shift_right[0]), 
        .ZN(u4_srl_452_n4) );
  INV_X8 u4_srl_452_U32 ( .A(u4_srl_452_n15), .ZN(u4_srl_452_n14) );
  INV_X8 u4_srl_452_U31 ( .A(u4_srl_452_n4), .ZN(u4_srl_452_n12) );
  NOR2_X2 u4_srl_452_U30 ( .A1(u4_srl_452_n309), .A2(u4_shift_right[1]), .ZN(
        u4_srl_452_n146) );
  INV_X4 u4_srl_452_U29 ( .A(u4_srl_452_n276), .ZN(u4_srl_452_n143) );
  AND2_X4 u4_srl_452_U28 ( .A1(u4_shift_right[4]), .A2(u4_srl_452_n281), .ZN(
        u4_srl_452_n3) );
  INV_X4 u4_srl_452_U27 ( .A(u4_srl_452_n21), .ZN(u4_srl_452_n19) );
  INV_X4 u4_srl_452_U26 ( .A(u4_srl_452_n21), .ZN(u4_srl_452_n20) );
  INV_X4 u4_srl_452_U25 ( .A(u4_srl_452_n146), .ZN(u4_srl_452_n21) );
  INV_X16 u4_srl_452_U24 ( .A(u4_srl_452_n15), .ZN(u4_srl_452_n13) );
  INV_X8 u4_srl_452_U23 ( .A(u4_srl_452_n3), .ZN(u4_srl_452_n6) );
  INV_X4 u4_srl_452_U22 ( .A(u4_srl_452_n1), .ZN(u4_srl_452_n9) );
  INV_X16 u4_srl_452_U21 ( .A(u4_srl_452_n25), .ZN(u4_srl_452_n22) );
  INV_X8 u4_srl_452_U20 ( .A(u4_srl_452_n18), .ZN(u4_srl_452_n16) );
  INV_X16 u4_srl_452_U19 ( .A(u4_srl_452_n25), .ZN(u4_srl_452_n24) );
  INV_X4 u4_srl_452_U18 ( .A(u4_srl_452_n144), .ZN(u4_srl_452_n18) );
  INV_X4 u4_srl_452_U17 ( .A(u4_shift_right[1]), .ZN(u4_srl_452_n5) );
  INV_X2 u4_srl_452_U16 ( .A(n5324), .ZN(u4_srl_452_n32) );
  INV_X2 u4_srl_452_U15 ( .A(fract_denorm[45]), .ZN(u4_srl_452_n61) );
  INV_X1 u4_srl_452_U14 ( .A(fract_denorm[31]), .ZN(u4_srl_452_n57) );
  INV_X1 u4_srl_452_U13 ( .A(fract_denorm[43]), .ZN(u4_srl_452_n63) );
  INV_X8 u4_srl_452_U12 ( .A(u4_srl_452_n12), .ZN(u4_srl_452_n15) );
  NAND2_X1 u4_srl_452_U11 ( .A1(u4_shift_right[1]), .A2(u4_srl_452_n309), .ZN(
        u4_srl_452_n144) );
  INV_X16 u4_srl_452_U10 ( .A(u4_srl_452_n18), .ZN(u4_srl_452_n17) );
  NAND2_X2 u4_srl_452_U9 ( .A1(u4_srl_452_n309), .A2(u4_srl_452_n5), .ZN(
        u4_srl_452_n2) );
  INV_X8 u4_srl_452_U8 ( .A(u4_srl_452_n2), .ZN(u4_srl_452_n23) );
  AND2_X4 u4_srl_452_U7 ( .A1(u4_srl_452_n280), .A2(u4_srl_452_n281), .ZN(
        u4_srl_452_n1) );
  INV_X16 u4_srl_452_U6 ( .A(u4_srl_452_n279), .ZN(u4_srl_452_n164) );
  INV_X2 u4_srl_452_U5 ( .A(fract_denorm[38]), .ZN(u4_srl_452_n55) );
  INV_X1 u4_srl_452_U4 ( .A(fract_denorm[36]), .ZN(u4_srl_452_n56) );
  INV_X2 u4_srl_452_U3 ( .A(net17655), .ZN(u4_srl_452_n69) );
  AND2_X1 u4_sll_481_U150 ( .A1(net17652), .A2(u4_sll_481_n33), .ZN(
        u4_sll_481_ML_int_1__0_) );
  AND2_X1 u4_sll_481_U149 ( .A1(net85391), .A2(u4_sll_481_n58), .ZN(
        u4_sll_481_MR_int_1__55_) );
  NAND2_X1 u4_sll_481_U148 ( .A1(u4_exp_in_mi1_1_), .A2(u4_sll_481_n88), .ZN(
        u4_sll_481_n94) );
  NAND2_X1 u4_sll_481_U147 ( .A1(u4_sll_481_ML_int_1__0_), .A2(u4_sll_481_n67), 
        .ZN(u4_sll_481_n92) );
  AND2_X1 u4_sll_481_U146 ( .A1(u4_sll_481_ML_int_1__1_), .A2(u4_sll_481_n67), 
        .ZN(u4_sll_481_ML_int_2__1_) );
  NAND2_X1 u4_sll_481_U145 ( .A1(u4_f2i_shft_2_), .A2(u4_sll_481_n88), .ZN(
        u4_sll_481_n93) );
  NOR2_X1 u4_sll_481_U144 ( .A1(u4_sll_481_n74), .A2(u4_sll_481_n92), .ZN(
        u4_sll_481_ML_int_3__0_) );
  NAND2_X1 u4_sll_481_U143 ( .A1(u4_f2i_shft_3_), .A2(u4_sll_481_n88), .ZN(
        u4_sll_481_n91) );
  NOR2_X1 u4_sll_481_U142 ( .A1(u4_sll_481_n75), .A2(u4_sll_481_n80), .ZN(
        u4_sll_481_n90) );
  AND2_X1 u4_sll_481_U141 ( .A1(u4_sll_481_n90), .A2(u4_sll_481_ML_int_2__1_), 
        .ZN(u4_sll_481_ML_int_4__1_) );
  AND2_X1 u4_sll_481_U140 ( .A1(u4_sll_481_ML_int_2__2_), .A2(u4_sll_481_n90), 
        .ZN(u4_sll_481_ML_int_4__2_) );
  AND2_X1 u4_sll_481_U139 ( .A1(u4_sll_481_ML_int_2__3_), .A2(u4_sll_481_n90), 
        .ZN(u4_sll_481_ML_int_4__3_) );
  AND2_X1 u4_sll_481_U138 ( .A1(u4_sll_481_ML_int_3__4_), .A2(u4_sll_481_n82), 
        .ZN(u4_sll_481_ML_int_4__4_) );
  AND2_X1 u4_sll_481_U137 ( .A1(u4_sll_481_ML_int_3__5_), .A2(u4_sll_481_n82), 
        .ZN(u4_sll_481_ML_int_4__5_) );
  AND2_X1 u4_sll_481_U136 ( .A1(u4_sll_481_ML_int_3__6_), .A2(u4_sll_481_n82), 
        .ZN(u4_sll_481_ML_int_4__6_) );
  AND2_X1 u4_sll_481_U135 ( .A1(u4_sll_481_ML_int_3__7_), .A2(u4_sll_481_n82), 
        .ZN(u4_sll_481_ML_int_4__7_) );
  OAI21_X1 u4_sll_481_U134 ( .B1(u4_f2i_shft_4_), .B2(u4_sll_481_n86), .A(
        u4_sll_481_n88), .ZN(u4_sll_481_SHMAG_4_) );
  OAI21_X1 u4_sll_481_U133 ( .B1(u4_f2i_shft_5_), .B2(u4_sll_481_n86), .A(
        u4_sll_481_n88), .ZN(u4_sll_481_SHMAG_5_) );
  INV_X4 u4_sll_481_U132 ( .A(u4_sll_481_n89), .ZN(u4_sll_481_n86) );
  INV_X4 u4_sll_481_U131 ( .A(u4_sll_481_SHMAG_4_), .ZN(u4_sll_481_n84) );
  INV_X4 u4_sll_481_U130 ( .A(u4_sll_481_n92), .ZN(u4_sll_481_n83) );
  INV_X32 u4_sll_481_U129 ( .A(u4_sll_481_n82), .ZN(u4_sll_481_n80) );
  INV_X32 u4_sll_481_U128 ( .A(u4_sll_481_n79), .ZN(u4_sll_481_n77) );
  INV_X32 u4_sll_481_U127 ( .A(u4_sll_481_n79), .ZN(u4_sll_481_n76) );
  INV_X32 u4_sll_481_U126 ( .A(u4_sll_481_n79), .ZN(u4_sll_481_n74) );
  INV_X16 u4_sll_481_U125 ( .A(u4_sll_481_n71), .ZN(u4_sll_481_n70) );
  INV_X16 u4_sll_481_U124 ( .A(u4_sll_481_n71), .ZN(u4_sll_481_n69) );
  INV_X16 u4_sll_481_U123 ( .A(u4_sll_481_n71), .ZN(u4_sll_481_n68) );
  INV_X16 u4_sll_481_U122 ( .A(u4_sll_481_n71), .ZN(u4_sll_481_n67) );
  INV_X32 u4_sll_481_U121 ( .A(u4_sll_481_n70), .ZN(u4_sll_481_n65) );
  NAND2_X4 u4_sll_481_U120 ( .A1(u4_sll_481_n89), .A2(u4_sll_481_n95), .ZN(
        u4_sll_481_temp_int_SH_0_) );
  INV_X8 u4_sll_481_U119 ( .A(u4_sll_481_n57), .ZN(u4_sll_481_n60) );
  INV_X16 u4_sll_481_U118 ( .A(u4_sll_481_n57), .ZN(u4_sll_481_n58) );
  INV_X16 u4_sll_481_U117 ( .A(u4_sll_481_temp_int_SH_0_), .ZN(u4_sll_481_n57)
         );
  INV_X4 u4_sll_481_U116 ( .A(u4_sll_481_temp_int_SH_1_), .ZN(u4_sll_481_n72)
         );
  AND2_X2 u4_sll_481_U115 ( .A1(u4_sll_481_ML_int_6__56_), .A2(u4_sll_481_n1), 
        .ZN(u4_exp_f2i_1[56]) );
  NAND2_X4 u4_sll_481_U114 ( .A1(net22501), .A2(u4_sll_481_n88), .ZN(
        u4_sll_481_n95) );
  MUX2_X2 u4_sll_481_U113 ( .A(u4_sll_481_ML_int_4__39_), .B(
        u4_sll_481_ML_int_4__55_), .S(u4_sll_481_SHMAG_4_), .Z(
        u4_sll_481_ML_int_5__55_) );
  NAND2_X2 u4_sll_481_U112 ( .A1(u4_sll_481_n89), .A2(u4_sll_481_n94), .ZN(
        u4_sll_481_temp_int_SH_1_) );
  MUX2_X1 u4_sll_481_U111 ( .A(u4_sll_481_ML_int_3__32_), .B(
        u4_sll_481_ML_int_3__40_), .S(u4_sll_481_n54), .Z(
        u4_sll_481_ML_int_4__40_) );
  MUX2_X2 u4_sll_481_U110 ( .A(u4_sll_481_ML_int_1__38_), .B(
        u4_sll_481_ML_int_1__40_), .S(u4_sll_481_n70), .Z(
        u4_sll_481_ML_int_2__40_) );
  AND2_X2 u4_sll_481_U109 ( .A1(u4_sll_481_ML_int_6__55_), .A2(u4_sll_481_n1), 
        .ZN(u4_exp_f2i_1[55]) );
  AND2_X2 u4_sll_481_U108 ( .A1(u4_sll_481_ML_int_6__54_), .A2(u4_sll_481_n1), 
        .ZN(u4_exp_f2i_1[54]) );
  AND2_X2 u4_sll_481_U107 ( .A1(u4_sll_481_ML_int_6__53_), .A2(u4_sll_481_n1), 
        .ZN(u4_exp_f2i_1[53]) );
  AND2_X2 u4_sll_481_U106 ( .A1(u4_sll_481_ML_int_6__51_), .A2(u4_sll_481_n1), 
        .ZN(u4_exp_f2i_1[51]) );
  AND2_X2 u4_sll_481_U105 ( .A1(u4_sll_481_ML_int_6__52_), .A2(u4_sll_481_n1), 
        .ZN(u4_exp_f2i_1[52]) );
  AND2_X2 u4_sll_481_U104 ( .A1(u4_sll_481_ML_int_6__50_), .A2(u4_sll_481_n1), 
        .ZN(u4_exp_f2i_1[50]) );
  AND2_X2 u4_sll_481_U103 ( .A1(u4_sll_481_ML_int_6__49_), .A2(u4_sll_481_n1), 
        .ZN(u4_exp_f2i_1[49]) );
  NOR2_X4 u4_sll_481_U102 ( .A1(u4_sll_481_n87), .A2(u4_f2i_shft_6_), .ZN(
        u4_sll_481_n53) );
  INV_X1 u4_sll_481_U101 ( .A(u4_sll_481_n84), .ZN(u4_sll_481_n50) );
  NAND2_X2 u4_sll_481_U100 ( .A1(u4_sll_481_n51), .A2(u4_sll_481_n52), .ZN(
        u4_sll_481_ML_int_5__56_) );
  NAND2_X1 u4_sll_481_U99 ( .A1(u4_sll_481_ML_int_4__40_), .A2(u4_sll_481_n84), 
        .ZN(u4_sll_481_n52) );
  NAND2_X2 u4_sll_481_U98 ( .A1(u4_sll_481_ML_int_4__56_), .A2(u4_sll_481_n50), 
        .ZN(u4_sll_481_n51) );
  NAND2_X2 u4_sll_481_U97 ( .A1(u4_sll_481_n48), .A2(u4_sll_481_n49), .ZN(
        u4_sll_481_ML_int_2__4_) );
  NAND2_X2 u4_sll_481_U96 ( .A1(u4_sll_481_ML_int_1__2_), .A2(u4_sll_481_n63), 
        .ZN(u4_sll_481_n49) );
  NAND2_X2 u4_sll_481_U95 ( .A1(u4_sll_481_ML_int_1__4_), .A2(u4_sll_481_n30), 
        .ZN(u4_sll_481_n48) );
  NAND2_X2 u4_sll_481_U94 ( .A1(u4_f2i_shft_6_), .A2(u4_sll_481_n87), .ZN(
        u4_sll_481_n89) );
  INV_X16 u4_sll_481_U93 ( .A(u4_sll_481_n67), .ZN(u4_sll_481_n63) );
  NAND2_X2 u4_sll_481_U92 ( .A1(u4_sll_481_n46), .A2(u4_sll_481_n47), .ZN(
        u4_sll_481_ML_int_2__11_) );
  NAND2_X1 u4_sll_481_U91 ( .A1(u4_sll_481_ML_int_1__9_), .A2(u4_sll_481_n63), 
        .ZN(u4_sll_481_n47) );
  NAND2_X1 u4_sll_481_U90 ( .A1(u4_sll_481_ML_int_1__11_), .A2(u4_sll_481_n24), 
        .ZN(u4_sll_481_n46) );
  NAND2_X2 u4_sll_481_U89 ( .A1(u4_sll_481_n44), .A2(u4_sll_481_n45), .ZN(
        u4_sll_481_ML_int_1__10_) );
  NAND2_X1 u4_sll_481_U88 ( .A1(n2980), .A2(u4_sll_481_n62), .ZN(
        u4_sll_481_n45) );
  NAND2_X1 u4_sll_481_U87 ( .A1(n5324), .A2(u4_sll_481_n43), .ZN(
        u4_sll_481_n44) );
  INV_X1 u4_sll_481_U86 ( .A(u4_sll_481_n77), .ZN(u4_sll_481_n40) );
  NAND2_X2 u4_sll_481_U85 ( .A1(u4_sll_481_n41), .A2(u4_sll_481_n42), .ZN(
        u4_sll_481_ML_int_3__16_) );
  NAND2_X1 u4_sll_481_U84 ( .A1(u4_sll_481_ML_int_2__12_), .A2(u4_sll_481_n77), 
        .ZN(u4_sll_481_n42) );
  NAND2_X1 u4_sll_481_U83 ( .A1(u4_sll_481_ML_int_2__16_), .A2(u4_sll_481_n40), 
        .ZN(u4_sll_481_n41) );
  INV_X16 u4_sll_481_U82 ( .A(u4_sll_481_n68), .ZN(u4_sll_481_n66) );
  NAND2_X2 u4_sll_481_U81 ( .A1(u4_sll_481_n38), .A2(u4_sll_481_n39), .ZN(
        u4_sll_481_ML_int_2__47_) );
  NAND2_X1 u4_sll_481_U80 ( .A1(u4_sll_481_ML_int_1__45_), .A2(u4_sll_481_n66), 
        .ZN(u4_sll_481_n39) );
  NAND2_X2 u4_sll_481_U79 ( .A1(u4_sll_481_ML_int_1__47_), .A2(u4_sll_481_n30), 
        .ZN(u4_sll_481_n38) );
  NAND2_X2 u4_sll_481_U78 ( .A1(u4_sll_481_n36), .A2(u4_sll_481_n37), .ZN(
        u4_sll_481_ML_int_3__47_) );
  NAND2_X2 u4_sll_481_U77 ( .A1(u4_sll_481_ML_int_2__47_), .A2(u4_sll_481_n6), 
        .ZN(u4_sll_481_n37) );
  NAND2_X1 u4_sll_481_U76 ( .A1(u4_sll_481_ML_int_2__43_), .A2(u4_sll_481_n75), 
        .ZN(u4_sll_481_n36) );
  INV_X1 u4_sll_481_U75 ( .A(u4_sll_481_n60), .ZN(u4_sll_481_n33) );
  NAND2_X2 u4_sll_481_U74 ( .A1(u4_sll_481_n34), .A2(u4_sll_481_n35), .ZN(
        u4_sll_481_ML_int_1__24_) );
  NAND2_X2 u4_sll_481_U73 ( .A1(n3067), .A2(u4_sll_481_n55), .ZN(
        u4_sll_481_n35) );
  NAND2_X1 u4_sll_481_U72 ( .A1(fract_denorm[24]), .A2(u4_sll_481_n33), .ZN(
        u4_sll_481_n34) );
  INV_X1 u4_sll_481_U71 ( .A(u4_sll_481_n64), .ZN(u4_sll_481_n30) );
  NAND2_X2 u4_sll_481_U70 ( .A1(u4_sll_481_n31), .A2(u4_sll_481_n32), .ZN(
        u4_sll_481_ML_int_2__26_) );
  NAND2_X2 u4_sll_481_U69 ( .A1(u4_sll_481_ML_int_1__24_), .A2(u4_sll_481_n64), 
        .ZN(u4_sll_481_n32) );
  NAND2_X1 u4_sll_481_U68 ( .A1(u4_sll_481_ML_int_1__26_), .A2(u4_sll_481_n30), 
        .ZN(u4_sll_481_n31) );
  MUX2_X2 u4_sll_481_U67 ( .A(u4_sll_481_ML_int_2__36_), .B(
        u4_sll_481_ML_int_2__40_), .S(u4_sll_481_n28), .Z(
        u4_sll_481_ML_int_3__40_) );
  INV_X1 u4_sll_481_U66 ( .A(u4_sll_481_n77), .ZN(u4_sll_481_n27) );
  NAND2_X2 u4_sll_481_U65 ( .A1(u4_sll_481_n25), .A2(u4_sll_481_n26), .ZN(
        u4_sll_481_ML_int_2__13_) );
  NAND2_X2 u4_sll_481_U64 ( .A1(u4_sll_481_ML_int_1__11_), .A2(u4_sll_481_n65), 
        .ZN(u4_sll_481_n26) );
  NAND2_X2 u4_sll_481_U63 ( .A1(u4_sll_481_ML_int_1__13_), .A2(u4_sll_481_n24), 
        .ZN(u4_sll_481_n25) );
  NAND2_X2 u4_sll_481_U62 ( .A1(u4_sll_481_n22), .A2(u4_sll_481_n23), .ZN(
        u4_sll_481_ML_int_3__13_) );
  NAND2_X2 u4_sll_481_U61 ( .A1(u4_sll_481_ML_int_2__13_), .A2(u4_sll_481_n27), 
        .ZN(u4_sll_481_n23) );
  NAND2_X1 u4_sll_481_U60 ( .A1(u4_sll_481_ML_int_2__9_), .A2(u4_sll_481_n21), 
        .ZN(u4_sll_481_n22) );
  NAND2_X2 u4_sll_481_U59 ( .A1(u4_sll_481_n19), .A2(u4_sll_481_n20), .ZN(
        u4_sll_481_ML_int_6__52_) );
  NAND2_X1 u4_sll_481_U58 ( .A1(u4_sll_481_ML_int_5__20_), .A2(u4_sll_481_n85), 
        .ZN(u4_sll_481_n20) );
  NAND2_X2 u4_sll_481_U57 ( .A1(u4_sll_481_ML_int_5__52_), .A2(u4_sll_481_n9), 
        .ZN(u4_sll_481_n19) );
  NAND2_X2 u4_sll_481_U56 ( .A1(u4_sll_481_n17), .A2(u4_sll_481_n18), .ZN(
        u4_sll_481_ML_int_3__29_) );
  NAND2_X1 u4_sll_481_U55 ( .A1(u4_sll_481_ML_int_2__29_), .A2(u4_sll_481_n28), 
        .ZN(u4_sll_481_n18) );
  NAND2_X1 u4_sll_481_U54 ( .A1(u4_sll_481_ML_int_2__25_), .A2(u4_sll_481_n21), 
        .ZN(u4_sll_481_n17) );
  NAND2_X2 u4_sll_481_U53 ( .A1(u4_sll_481_n15), .A2(u4_sll_481_n16), .ZN(
        u4_sll_481_ML_int_6__53_) );
  NAND2_X1 u4_sll_481_U52 ( .A1(u4_sll_481_ML_int_5__21_), .A2(u4_sll_481_n85), 
        .ZN(u4_sll_481_n16) );
  NAND2_X2 u4_sll_481_U51 ( .A1(u4_sll_481_ML_int_5__53_), .A2(u4_sll_481_n9), 
        .ZN(u4_sll_481_n15) );
  MUX2_X1 u4_sll_481_U50 ( .A(u4_sll_481_ML_int_3__26_), .B(
        u4_sll_481_ML_int_3__34_), .S(u4_sll_481_n54), .Z(
        u4_sll_481_ML_int_4__34_) );
  INV_X16 u4_sll_481_U49 ( .A(u4_sll_481_n82), .ZN(u4_sll_481_n81) );
  MUX2_X2 u4_sll_481_U48 ( .A(u4_sll_481_ML_int_3__10_), .B(
        u4_sll_481_ML_int_3__18_), .S(u4_sll_481_n82), .Z(
        u4_sll_481_ML_int_4__18_) );
  CLKBUF_X3 u4_sll_481_U47 ( .A(u4_sll_481_ML_int_1__7_), .Z(u4_sll_481_n29)
         );
  MUX2_X2 u4_sll_481_U46 ( .A(u4_sll_481_n29), .B(u4_sll_481_ML_int_1__5_), 
        .S(u4_sll_481_n63), .Z(u4_sll_481_n14) );
  MUX2_X2 u4_sll_481_U45 ( .A(u4_sll_481_ML_int_1__8_), .B(
        u4_sll_481_ML_int_1__10_), .S(u4_sll_481_n67), .Z(
        u4_sll_481_ML_int_2__10_) );
  NAND2_X2 u4_sll_481_U44 ( .A1(u4_sll_481_n12), .A2(u4_sll_481_n13), .ZN(
        u4_sll_481_ML_int_6__51_) );
  NAND2_X1 u4_sll_481_U43 ( .A1(u4_sll_481_ML_int_5__19_), .A2(u4_sll_481_n85), 
        .ZN(u4_sll_481_n13) );
  NAND2_X2 u4_sll_481_U42 ( .A1(u4_sll_481_ML_int_5__51_), .A2(u4_sll_481_n9), 
        .ZN(u4_sll_481_n12) );
  INV_X8 u4_sll_481_U41 ( .A(u4_sll_481_n57), .ZN(u4_sll_481_n62) );
  NAND2_X2 u4_sll_481_U40 ( .A1(u4_sll_481_n10), .A2(u4_sll_481_n11), .ZN(
        u4_sll_481_ML_int_6__50_) );
  NAND2_X1 u4_sll_481_U39 ( .A1(u4_sll_481_ML_int_5__18_), .A2(u4_sll_481_n85), 
        .ZN(u4_sll_481_n11) );
  NAND2_X2 u4_sll_481_U38 ( .A1(u4_sll_481_ML_int_5__50_), .A2(u4_sll_481_n9), 
        .ZN(u4_sll_481_n10) );
  MUX2_X1 u4_sll_481_U37 ( .A(u4_sll_481_ML_int_3__25_), .B(
        u4_sll_481_ML_int_3__33_), .S(u4_sll_481_n82), .Z(
        u4_sll_481_ML_int_4__33_) );
  NAND2_X2 u4_sll_481_U36 ( .A1(u4_sll_481_n7), .A2(u4_sll_481_n8), .ZN(
        u4_sll_481_ML_int_1__17_) );
  NAND2_X1 u4_sll_481_U35 ( .A1(net17684), .A2(u4_sll_481_n61), .ZN(
        u4_sll_481_n8) );
  NAND2_X1 u4_sll_481_U34 ( .A1(net17657), .A2(u4_sll_481_n43), .ZN(
        u4_sll_481_n7) );
  INV_X2 u4_sll_481_U33 ( .A(u4_sll_481_n81), .ZN(u4_sll_481_n54) );
  INV_X4 u4_sll_481_U32 ( .A(u4_sll_481_n65), .ZN(u4_sll_481_n24) );
  INV_X4 u4_sll_481_U31 ( .A(u4_sll_481_SHMAG_5_), .ZN(u4_sll_481_n85) );
  INV_X4 u4_sll_481_U30 ( .A(u4_sll_481_n76), .ZN(u4_sll_481_n28) );
  INV_X16 u4_sll_481_U29 ( .A(u4_sll_481_n73), .ZN(u4_sll_481_n79) );
  INV_X8 u4_sll_481_U28 ( .A(u4_sll_481_n6), .ZN(u4_sll_481_n73) );
  INV_X2 u4_sll_481_U27 ( .A(u4_sll_481_n85), .ZN(u4_sll_481_n9) );
  INV_X8 u4_sll_481_U26 ( .A(u4_sll_481_temp_int_SH_3_), .ZN(u4_sll_481_n82)
         );
  AND2_X4 u4_sll_481_U25 ( .A1(u4_sll_481_n89), .A2(u4_sll_481_n93), .ZN(
        u4_sll_481_n6) );
  INV_X2 u4_sll_481_U24 ( .A(u4_sll_481_n27), .ZN(u4_sll_481_n21) );
  INV_X16 u4_sll_481_U23 ( .A(u4_sll_481_n79), .ZN(u4_sll_481_n75) );
  NAND2_X2 u4_sll_481_U22 ( .A1(u4_sll_481_n89), .A2(u4_sll_481_n91), .ZN(
        u4_sll_481_temp_int_SH_3_) );
  INV_X16 u4_sll_481_U21 ( .A(u4_sll_481_n72), .ZN(u4_sll_481_n71) );
  INV_X8 u4_sll_481_U20 ( .A(u4_sll_481_n57), .ZN(u4_sll_481_n61) );
  INV_X16 u4_sll_481_U19 ( .A(u4_sll_481_n53), .ZN(u4_sll_481_n88) );
  INV_X32 u4_sll_481_U18 ( .A(u4_sll_481_n66), .ZN(u4_sll_481_n5) );
  MUX2_X2 u4_sll_481_U17 ( .A(u4_sll_481_ML_int_1__49_), .B(
        u4_sll_481_ML_int_1__51_), .S(u4_sll_481_n5), .Z(
        u4_sll_481_ML_int_2__51_) );
  INV_X2 u4_sll_481_U16 ( .A(u4_sll_481_n57), .ZN(u4_sll_481_n59) );
  INV_X32 u4_sll_481_U15 ( .A(u4_sll_481_n69), .ZN(u4_sll_481_n64) );
  MUX2_X2 u4_sll_481_U14 ( .A(u4_sll_481_ML_int_1__25_), .B(
        u4_sll_481_ML_int_1__27_), .S(u4_sll_481_n69), .Z(
        u4_sll_481_ML_int_2__27_) );
  INV_X1 u4_sll_481_U13 ( .A(u4_sll_481_n76), .ZN(u4_sll_481_n2) );
  NAND2_X2 u4_sll_481_U12 ( .A1(u4_sll_481_n3), .A2(u4_sll_481_n4), .ZN(
        u4_sll_481_ML_int_3__31_) );
  NAND2_X1 u4_sll_481_U11 ( .A1(u4_sll_481_ML_int_2__27_), .A2(u4_sll_481_n76), 
        .ZN(u4_sll_481_n4) );
  NAND2_X1 u4_sll_481_U10 ( .A1(u4_sll_481_ML_int_2__31_), .A2(u4_sll_481_n2), 
        .ZN(u4_sll_481_n3) );
  INV_X16 u4_sll_481_U9 ( .A(u4_sll_481_n79), .ZN(u4_sll_481_n78) );
  MUX2_X2 u4_sll_481_U8 ( .A(u4_sll_481_ML_int_2__5_), .B(
        u4_sll_481_ML_int_2__9_), .S(u4_sll_481_n79), .Z(
        u4_sll_481_ML_int_3__9_) );
  INV_X32 u4_sll_481_U7 ( .A(u4_sll_481_n57), .ZN(u4_sll_481_n55) );
  INV_X1 u4_sll_481_U6 ( .A(u4_sll_481_n62), .ZN(u4_sll_481_n43) );
  INV_X16 u4_sll_481_U5 ( .A(u4_sll_481_n57), .ZN(u4_sll_481_n56) );
  INV_X8 u4_sll_481_U4 ( .A(u4_f2i_shft_7_), .ZN(u4_sll_481_n87) );
  BUF_X32 u4_sll_481_U3 ( .A(u4_sll_481_n87), .Z(u4_sll_481_n1) );
  MUX2_X2 u4_sll_481_M1_2_15 ( .A(u4_sll_481_ML_int_2__15_), .B(
        u4_sll_481_ML_int_2__11_), .S(u4_sll_481_n77), .Z(
        u4_sll_481_ML_int_3__15_) );
  MUX2_X1 u4_sll_481_M1_2_33 ( .A(u4_sll_481_ML_int_2__33_), .B(
        u4_sll_481_ML_int_2__29_), .S(u4_sll_481_n76), .Z(
        u4_sll_481_ML_int_3__33_) );
  MUX2_X1 u4_sll_481_M1_5_49 ( .A(u4_sll_481_ML_int_5__49_), .B(
        u4_sll_481_ML_int_5__17_), .S(u4_sll_481_n85), .Z(
        u4_sll_481_ML_int_6__49_) );
  MUX2_X1 u4_sll_481_M1_2_11 ( .A(u4_sll_481_ML_int_2__11_), .B(u4_sll_481_n14), .S(u4_sll_481_n78), .Z(u4_sll_481_ML_int_3__11_) );
  MUX2_X1 u4_sll_481_M1_2_10 ( .A(u4_sll_481_ML_int_2__10_), .B(
        u4_sll_481_ML_int_2__6_), .S(u4_sll_481_n78), .Z(
        u4_sll_481_ML_int_3__10_) );
  MUX2_X1 u4_sll_481_M1_2_26 ( .A(u4_sll_481_ML_int_2__26_), .B(
        u4_sll_481_ML_int_2__22_), .S(u4_sll_481_n76), .Z(
        u4_sll_481_ML_int_3__26_) );
  MUX2_X1 u4_sll_481_M1_2_25 ( .A(u4_sll_481_ML_int_2__25_), .B(
        u4_sll_481_ML_int_2__21_), .S(u4_sll_481_n76), .Z(
        u4_sll_481_ML_int_3__25_) );
  MUX2_X1 u4_sll_481_M1_3_37 ( .A(u4_sll_481_ML_int_3__37_), .B(
        u4_sll_481_ML_int_3__29_), .S(u4_sll_481_n80), .Z(
        u4_sll_481_ML_int_4__37_) );
  MUX2_X2 u4_sll_481_M1_3_55 ( .A(u4_sll_481_ML_int_3__55_), .B(
        u4_sll_481_ML_int_3__47_), .S(u4_sll_481_n81), .Z(
        u4_sll_481_ML_int_4__55_) );
  MUX2_X1 u4_sll_481_M1_2_44 ( .A(u4_sll_481_ML_int_2__44_), .B(
        u4_sll_481_ML_int_2__40_), .S(u4_sll_481_n75), .Z(
        u4_sll_481_ML_int_3__44_) );
  MUX2_X2 u4_sll_481_M1_5_55 ( .A(u4_sll_481_ML_int_5__55_), .B(
        u4_sll_481_ML_int_5__23_), .S(u4_sll_481_n85), .Z(
        u4_sll_481_ML_int_6__55_) );
  MUX2_X1 u4_sll_481_M1_5_56 ( .A(u4_sll_481_ML_int_5__56_), .B(
        u4_sll_481_ML_int_5__24_), .S(u4_sll_481_n85), .Z(
        u4_sll_481_ML_int_6__56_) );
  MUX2_X2 u4_sll_481_M1_3_39 ( .A(u4_sll_481_ML_int_3__39_), .B(
        u4_sll_481_ML_int_3__31_), .S(u4_sll_481_n81), .Z(
        u4_sll_481_ML_int_4__39_) );
  MUX2_X1 u4_sll_481_M1_2_32 ( .A(u4_sll_481_ML_int_2__32_), .B(
        u4_sll_481_ML_int_2__28_), .S(u4_sll_481_n76), .Z(
        u4_sll_481_ML_int_3__32_) );
  MUX2_X2 u4_sll_481_M1_0_1 ( .A(net17695), .B(net17652), .S(u4_sll_481_n60), 
        .Z(u4_sll_481_ML_int_1__1_) );
  MUX2_X2 u4_sll_481_M1_0_2 ( .A(net17694), .B(net17695), .S(u4_sll_481_n55), 
        .Z(u4_sll_481_ML_int_1__2_) );
  MUX2_X2 u4_sll_481_M1_0_3 ( .A(net17653), .B(net17694), .S(u4_sll_481_n61), 
        .Z(u4_sll_481_ML_int_1__3_) );
  MUX2_X2 u4_sll_481_M1_0_4 ( .A(net17693), .B(net17653), .S(u4_sll_481_n58), 
        .Z(u4_sll_481_ML_int_1__4_) );
  MUX2_X2 u4_sll_481_M1_0_5 ( .A(net17692), .B(net17693), .S(u4_sll_481_n55), 
        .Z(u4_sll_481_ML_int_1__5_) );
  MUX2_X2 u4_sll_481_M1_0_6 ( .A(net17654), .B(net17692), .S(u4_sll_481_n56), 
        .Z(u4_sll_481_ML_int_1__6_) );
  MUX2_X2 u4_sll_481_M1_0_7 ( .A(n5323), .B(net17654), .S(u4_sll_481_n58), .Z(
        u4_sll_481_ML_int_1__7_) );
  MUX2_X2 u4_sll_481_M1_0_8 ( .A(net17690), .B(n5323), .S(u4_sll_481_n62), .Z(
        u4_sll_481_ML_int_1__8_) );
  MUX2_X2 u4_sll_481_M1_0_9 ( .A(n2980), .B(net17690), .S(u4_sll_481_n62), .Z(
        u4_sll_481_ML_int_1__9_) );
  MUX2_X2 u4_sll_481_M1_0_11 ( .A(net95118), .B(n5324), .S(u4_sll_481_n55), 
        .Z(u4_sll_481_ML_int_1__11_) );
  MUX2_X2 u4_sll_481_M1_0_12 ( .A(n5326), .B(net95118), .S(u4_sll_481_n55), 
        .Z(u4_sll_481_ML_int_1__12_) );
  MUX2_X2 u4_sll_481_M1_0_13 ( .A(net17686), .B(n5326), .S(u4_sll_481_n56), 
        .Z(u4_sll_481_ML_int_1__13_) );
  MUX2_X2 u4_sll_481_M1_0_14 ( .A(net17656), .B(net17686), .S(u4_sll_481_n62), 
        .Z(u4_sll_481_ML_int_1__14_) );
  MUX2_X2 u4_sll_481_M1_0_15 ( .A(net17685), .B(net17656), .S(u4_sll_481_n55), 
        .Z(u4_sll_481_ML_int_1__15_) );
  MUX2_X2 u4_sll_481_M1_0_16 ( .A(net17684), .B(net17685), .S(u4_sll_481_n55), 
        .Z(u4_sll_481_ML_int_1__16_) );
  MUX2_X2 u4_sll_481_M1_0_18 ( .A(net17683), .B(net17657), .S(u4_sll_481_n56), 
        .Z(u4_sll_481_ML_int_1__18_) );
  MUX2_X2 u4_sll_481_M1_0_19 ( .A(net17682), .B(net17683), .S(u4_sll_481_n60), 
        .Z(u4_sll_481_ML_int_1__19_) );
  MUX2_X2 u4_sll_481_M1_0_20 ( .A(net17659), .B(net17682), .S(u4_sll_481_n61), 
        .Z(u4_sll_481_ML_int_1__20_) );
  MUX2_X2 u4_sll_481_M1_0_21 ( .A(fract_denorm[21]), .B(net17659), .S(
        u4_sll_481_n58), .Z(u4_sll_481_ML_int_1__21_) );
  MUX2_X2 u4_sll_481_M1_0_22 ( .A(fract_denorm[22]), .B(fract_denorm[21]), .S(
        u4_sll_481_n55), .Z(u4_sll_481_ML_int_1__22_) );
  MUX2_X2 u4_sll_481_M1_0_23 ( .A(n3067), .B(fract_denorm[22]), .S(
        u4_sll_481_n62), .Z(u4_sll_481_ML_int_1__23_) );
  MUX2_X2 u4_sll_481_M1_0_25 ( .A(fract_denorm[25]), .B(fract_denorm[24]), .S(
        u4_sll_481_n58), .Z(u4_sll_481_ML_int_1__25_) );
  MUX2_X2 u4_sll_481_M1_0_26 ( .A(fract_denorm[26]), .B(fract_denorm[25]), .S(
        u4_sll_481_n55), .Z(u4_sll_481_ML_int_1__26_) );
  MUX2_X2 u4_sll_481_M1_0_27 ( .A(fract_denorm[27]), .B(fract_denorm[26]), .S(
        u4_sll_481_n56), .Z(u4_sll_481_ML_int_1__27_) );
  MUX2_X2 u4_sll_481_M1_0_28 ( .A(fract_denorm[28]), .B(fract_denorm[27]), .S(
        u4_sll_481_n60), .Z(u4_sll_481_ML_int_1__28_) );
  MUX2_X2 u4_sll_481_M1_0_29 ( .A(n3006), .B(fract_denorm[28]), .S(
        u4_sll_481_n58), .Z(u4_sll_481_ML_int_1__29_) );
  MUX2_X2 u4_sll_481_M1_0_30 ( .A(n3008), .B(n3006), .S(u4_sll_481_n58), .Z(
        u4_sll_481_ML_int_1__30_) );
  MUX2_X2 u4_sll_481_M1_0_31 ( .A(fract_denorm[31]), .B(n3008), .S(
        u4_sll_481_n59), .Z(u4_sll_481_ML_int_1__31_) );
  MUX2_X2 u4_sll_481_M1_0_32 ( .A(fract_denorm[32]), .B(fract_denorm[31]), .S(
        u4_sll_481_n55), .Z(u4_sll_481_ML_int_1__32_) );
  MUX2_X2 u4_sll_481_M1_0_33 ( .A(fract_denorm[33]), .B(fract_denorm[32]), .S(
        u4_sll_481_n55), .Z(u4_sll_481_ML_int_1__33_) );
  MUX2_X2 u4_sll_481_M1_0_34 ( .A(fract_denorm[34]), .B(fract_denorm[33]), .S(
        u4_sll_481_n55), .Z(u4_sll_481_ML_int_1__34_) );
  MUX2_X2 u4_sll_481_M1_0_35 ( .A(n2483), .B(fract_denorm[34]), .S(
        u4_sll_481_n58), .Z(u4_sll_481_ML_int_1__35_) );
  MUX2_X2 u4_sll_481_M1_0_36 ( .A(fract_denorm[36]), .B(n2483), .S(
        u4_sll_481_n55), .Z(u4_sll_481_ML_int_1__36_) );
  MUX2_X2 u4_sll_481_M1_0_37 ( .A(fract_denorm[37]), .B(fract_denorm[36]), .S(
        u4_sll_481_n58), .Z(u4_sll_481_ML_int_1__37_) );
  MUX2_X2 u4_sll_481_M1_0_38 ( .A(fract_denorm[38]), .B(fract_denorm[37]), .S(
        u4_sll_481_n55), .Z(u4_sll_481_ML_int_1__38_) );
  MUX2_X2 u4_sll_481_M1_0_39 ( .A(n3023), .B(fract_denorm[38]), .S(
        u4_sll_481_n60), .Z(u4_sll_481_ML_int_1__39_) );
  MUX2_X2 u4_sll_481_M1_0_40 ( .A(n3024), .B(n3023), .S(u4_sll_481_n58), .Z(
        u4_sll_481_ML_int_1__40_) );
  MUX2_X2 u4_sll_481_M1_0_41 ( .A(net28939), .B(n3024), .S(u4_sll_481_n61), 
        .Z(u4_sll_481_ML_int_1__41_) );
  MUX2_X2 u4_sll_481_M1_0_42 ( .A(net94305), .B(net28939), .S(u4_sll_481_n58), 
        .Z(u4_sll_481_ML_int_1__42_) );
  MUX2_X2 u4_sll_481_M1_0_43 ( .A(fract_denorm[43]), .B(net94305), .S(
        u4_sll_481_n55), .Z(u4_sll_481_ML_int_1__43_) );
  MUX2_X2 u4_sll_481_M1_0_44 ( .A(fract_denorm[44]), .B(fract_denorm[43]), .S(
        u4_sll_481_n55), .Z(u4_sll_481_ML_int_1__44_) );
  MUX2_X2 u4_sll_481_M1_0_45 ( .A(fract_denorm[45]), .B(fract_denorm[44]), .S(
        u4_sll_481_n60), .Z(u4_sll_481_ML_int_1__45_) );
  MUX2_X2 u4_sll_481_M1_0_46 ( .A(net86571), .B(fract_denorm[45]), .S(
        u4_sll_481_n58), .Z(u4_sll_481_ML_int_1__46_) );
  MUX2_X2 u4_sll_481_M1_0_47 ( .A(net85391), .B(net86571), .S(u4_sll_481_n55), 
        .Z(u4_sll_481_ML_int_1__47_) );
  MUX2_X2 u4_sll_481_M1_0_49 ( .A(net85391), .B(net85391), .S(u4_sll_481_n61), 
        .Z(u4_sll_481_ML_int_1__49_) );
  MUX2_X2 u4_sll_481_M1_0_51 ( .A(net85391), .B(net85391), .S(u4_sll_481_n56), 
        .Z(u4_sll_481_ML_int_1__51_) );
  MUX2_X2 u4_sll_481_M1_0_52 ( .A(net85391), .B(net85391), .S(u4_sll_481_n61), 
        .Z(u4_sll_481_ML_int_1__52_) );
  MUX2_X2 u4_sll_481_M1_0_53 ( .A(net85391), .B(net85391), .S(u4_sll_481_n55), 
        .Z(u4_sll_481_ML_int_1__53_) );
  MUX2_X2 u4_sll_481_M1_0_54 ( .A(net85391), .B(net85391), .S(u4_sll_481_n55), 
        .Z(u4_sll_481_ML_int_1__54_) );
  MUX2_X2 u4_sll_481_M1_0_55 ( .A(net85391), .B(net85391), .S(u4_sll_481_n55), 
        .Z(u4_sll_481_ML_int_1__55_) );
  MUX2_X2 u4_sll_481_M1_1_2 ( .A(u4_sll_481_ML_int_1__2_), .B(
        u4_sll_481_ML_int_1__0_), .S(u4_sll_481_n63), .Z(
        u4_sll_481_ML_int_2__2_) );
  MUX2_X2 u4_sll_481_M1_1_3 ( .A(u4_sll_481_ML_int_1__3_), .B(
        u4_sll_481_ML_int_1__1_), .S(u4_sll_481_n63), .Z(
        u4_sll_481_ML_int_2__3_) );
  MUX2_X2 u4_sll_481_M1_1_5 ( .A(u4_sll_481_ML_int_1__5_), .B(
        u4_sll_481_ML_int_1__3_), .S(u4_sll_481_n63), .Z(
        u4_sll_481_ML_int_2__5_) );
  MUX2_X2 u4_sll_481_M1_1_6 ( .A(u4_sll_481_ML_int_1__6_), .B(
        u4_sll_481_ML_int_1__4_), .S(u4_sll_481_n63), .Z(
        u4_sll_481_ML_int_2__6_) );
  MUX2_X2 u4_sll_481_M1_1_8 ( .A(u4_sll_481_ML_int_1__8_), .B(
        u4_sll_481_ML_int_1__6_), .S(u4_sll_481_n63), .Z(
        u4_sll_481_ML_int_2__8_) );
  MUX2_X2 u4_sll_481_M1_1_9 ( .A(u4_sll_481_ML_int_1__9_), .B(
        u4_sll_481_ML_int_1__7_), .S(u4_sll_481_n63), .Z(
        u4_sll_481_ML_int_2__9_) );
  MUX2_X2 u4_sll_481_M1_1_12 ( .A(u4_sll_481_ML_int_1__12_), .B(
        u4_sll_481_ML_int_1__10_), .S(u4_sll_481_n63), .Z(
        u4_sll_481_ML_int_2__12_) );
  MUX2_X2 u4_sll_481_M1_1_14 ( .A(u4_sll_481_ML_int_1__14_), .B(
        u4_sll_481_ML_int_1__12_), .S(u4_sll_481_n66), .Z(
        u4_sll_481_ML_int_2__14_) );
  MUX2_X2 u4_sll_481_M1_1_15 ( .A(u4_sll_481_ML_int_1__15_), .B(
        u4_sll_481_ML_int_1__13_), .S(u4_sll_481_n65), .Z(
        u4_sll_481_ML_int_2__15_) );
  MUX2_X2 u4_sll_481_M1_1_16 ( .A(u4_sll_481_ML_int_1__16_), .B(
        u4_sll_481_ML_int_1__14_), .S(u4_sll_481_n66), .Z(
        u4_sll_481_ML_int_2__16_) );
  MUX2_X2 u4_sll_481_M1_1_17 ( .A(u4_sll_481_ML_int_1__17_), .B(
        u4_sll_481_ML_int_1__15_), .S(u4_sll_481_n65), .Z(
        u4_sll_481_ML_int_2__17_) );
  MUX2_X2 u4_sll_481_M1_1_18 ( .A(u4_sll_481_ML_int_1__18_), .B(
        u4_sll_481_ML_int_1__16_), .S(u4_sll_481_n65), .Z(
        u4_sll_481_ML_int_2__18_) );
  MUX2_X2 u4_sll_481_M1_1_19 ( .A(u4_sll_481_ML_int_1__19_), .B(
        u4_sll_481_ML_int_1__17_), .S(u4_sll_481_n65), .Z(
        u4_sll_481_ML_int_2__19_) );
  MUX2_X2 u4_sll_481_M1_1_20 ( .A(u4_sll_481_ML_int_1__20_), .B(
        u4_sll_481_ML_int_1__18_), .S(u4_sll_481_n65), .Z(
        u4_sll_481_ML_int_2__20_) );
  MUX2_X2 u4_sll_481_M1_1_21 ( .A(u4_sll_481_ML_int_1__21_), .B(
        u4_sll_481_ML_int_1__19_), .S(u4_sll_481_n65), .Z(
        u4_sll_481_ML_int_2__21_) );
  MUX2_X2 u4_sll_481_M1_1_22 ( .A(u4_sll_481_ML_int_1__22_), .B(
        u4_sll_481_ML_int_1__20_), .S(u4_sll_481_n65), .Z(
        u4_sll_481_ML_int_2__22_) );
  MUX2_X2 u4_sll_481_M1_1_23 ( .A(u4_sll_481_ML_int_1__23_), .B(
        u4_sll_481_ML_int_1__21_), .S(u4_sll_481_n65), .Z(
        u4_sll_481_ML_int_2__23_) );
  MUX2_X2 u4_sll_481_M1_1_24 ( .A(u4_sll_481_ML_int_1__24_), .B(
        u4_sll_481_ML_int_1__22_), .S(u4_sll_481_n64), .Z(
        u4_sll_481_ML_int_2__24_) );
  MUX2_X2 u4_sll_481_M1_1_25 ( .A(u4_sll_481_ML_int_1__25_), .B(
        u4_sll_481_ML_int_1__23_), .S(u4_sll_481_n64), .Z(
        u4_sll_481_ML_int_2__25_) );
  MUX2_X2 u4_sll_481_M1_1_28 ( .A(u4_sll_481_ML_int_1__28_), .B(
        u4_sll_481_ML_int_1__26_), .S(u4_sll_481_n64), .Z(
        u4_sll_481_ML_int_2__28_) );
  MUX2_X2 u4_sll_481_M1_1_29 ( .A(u4_sll_481_ML_int_1__29_), .B(
        u4_sll_481_ML_int_1__27_), .S(u4_sll_481_n64), .Z(
        u4_sll_481_ML_int_2__29_) );
  MUX2_X2 u4_sll_481_M1_1_30 ( .A(u4_sll_481_ML_int_1__30_), .B(
        u4_sll_481_ML_int_1__28_), .S(u4_sll_481_n64), .Z(
        u4_sll_481_ML_int_2__30_) );
  MUX2_X2 u4_sll_481_M1_1_31 ( .A(u4_sll_481_ML_int_1__31_), .B(
        u4_sll_481_ML_int_1__29_), .S(u4_sll_481_n64), .Z(
        u4_sll_481_ML_int_2__31_) );
  MUX2_X2 u4_sll_481_M1_1_32 ( .A(u4_sll_481_ML_int_1__32_), .B(
        u4_sll_481_ML_int_1__30_), .S(u4_sll_481_n64), .Z(
        u4_sll_481_ML_int_2__32_) );
  MUX2_X2 u4_sll_481_M1_1_33 ( .A(u4_sll_481_ML_int_1__33_), .B(
        u4_sll_481_ML_int_1__31_), .S(u4_sll_481_n64), .Z(
        u4_sll_481_ML_int_2__33_) );
  MUX2_X2 u4_sll_481_M1_1_34 ( .A(u4_sll_481_ML_int_1__34_), .B(
        u4_sll_481_ML_int_1__32_), .S(u4_sll_481_n64), .Z(
        u4_sll_481_ML_int_2__34_) );
  MUX2_X2 u4_sll_481_M1_1_35 ( .A(u4_sll_481_ML_int_1__35_), .B(
        u4_sll_481_ML_int_1__33_), .S(u4_sll_481_n65), .Z(
        u4_sll_481_ML_int_2__35_) );
  MUX2_X2 u4_sll_481_M1_1_36 ( .A(u4_sll_481_ML_int_1__36_), .B(
        u4_sll_481_ML_int_1__34_), .S(u4_sll_481_n65), .Z(
        u4_sll_481_ML_int_2__36_) );
  MUX2_X2 u4_sll_481_M1_1_37 ( .A(u4_sll_481_ML_int_1__37_), .B(
        u4_sll_481_ML_int_1__35_), .S(u4_sll_481_n65), .Z(
        u4_sll_481_ML_int_2__37_) );
  MUX2_X2 u4_sll_481_M1_1_38 ( .A(u4_sll_481_ML_int_1__38_), .B(
        u4_sll_481_ML_int_1__36_), .S(u4_sll_481_n65), .Z(
        u4_sll_481_ML_int_2__38_) );
  MUX2_X2 u4_sll_481_M1_1_39 ( .A(u4_sll_481_ML_int_1__39_), .B(
        u4_sll_481_ML_int_1__37_), .S(u4_sll_481_n65), .Z(
        u4_sll_481_ML_int_2__39_) );
  MUX2_X2 u4_sll_481_M1_1_41 ( .A(u4_sll_481_ML_int_1__41_), .B(
        u4_sll_481_ML_int_1__39_), .S(u4_sll_481_n65), .Z(
        u4_sll_481_ML_int_2__41_) );
  MUX2_X2 u4_sll_481_M1_1_42 ( .A(u4_sll_481_ML_int_1__42_), .B(
        u4_sll_481_ML_int_1__40_), .S(u4_sll_481_n65), .Z(
        u4_sll_481_ML_int_2__42_) );
  MUX2_X2 u4_sll_481_M1_1_43 ( .A(u4_sll_481_ML_int_1__43_), .B(
        u4_sll_481_ML_int_1__41_), .S(u4_sll_481_n65), .Z(
        u4_sll_481_ML_int_2__43_) );
  MUX2_X2 u4_sll_481_M1_1_44 ( .A(u4_sll_481_ML_int_1__44_), .B(
        u4_sll_481_ML_int_1__42_), .S(u4_sll_481_n65), .Z(
        u4_sll_481_ML_int_2__44_) );
  MUX2_X2 u4_sll_481_M1_1_45 ( .A(u4_sll_481_ML_int_1__45_), .B(
        u4_sll_481_ML_int_1__43_), .S(u4_sll_481_n65), .Z(
        u4_sll_481_ML_int_2__45_) );
  MUX2_X2 u4_sll_481_M1_1_46 ( .A(u4_sll_481_ML_int_1__46_), .B(
        u4_sll_481_ML_int_1__44_), .S(u4_sll_481_n66), .Z(
        u4_sll_481_ML_int_2__46_) );
  MUX2_X2 u4_sll_481_M1_1_48 ( .A(u4_sll_481_ML_int_1__54_), .B(
        u4_sll_481_ML_int_1__46_), .S(u4_sll_481_n66), .Z(
        u4_sll_481_ML_int_2__48_) );
  MUX2_X2 u4_sll_481_M1_1_49 ( .A(u4_sll_481_ML_int_1__49_), .B(
        u4_sll_481_ML_int_1__47_), .S(u4_sll_481_n66), .Z(
        u4_sll_481_ML_int_2__49_) );
  MUX2_X2 u4_sll_481_M1_1_50 ( .A(u4_sll_481_ML_int_1__52_), .B(
        u4_sll_481_ML_int_1__55_), .S(u4_sll_481_n66), .Z(
        u4_sll_481_ML_int_2__50_) );
  MUX2_X2 u4_sll_481_M1_1_52 ( .A(u4_sll_481_ML_int_1__52_), .B(
        u4_sll_481_ML_int_1__54_), .S(u4_sll_481_n66), .Z(
        u4_sll_481_ML_int_2__52_) );
  MUX2_X2 u4_sll_481_M1_1_53 ( .A(u4_sll_481_ML_int_1__53_), .B(
        u4_sll_481_ML_int_1__55_), .S(u4_sll_481_n66), .Z(
        u4_sll_481_ML_int_2__53_) );
  MUX2_X2 u4_sll_481_M1_1_54 ( .A(u4_sll_481_ML_int_1__54_), .B(
        u4_sll_481_ML_int_1__52_), .S(u4_sll_481_n66), .Z(
        u4_sll_481_ML_int_2__54_) );
  MUX2_X2 u4_sll_481_M1_1_55 ( .A(u4_sll_481_ML_int_1__55_), .B(
        u4_sll_481_ML_int_1__53_), .S(u4_sll_481_n66), .Z(
        u4_sll_481_ML_int_2__55_) );
  MUX2_X2 u4_sll_481_M1_1_56 ( .A(u4_sll_481_MR_int_1__55_), .B(
        u4_sll_481_ML_int_1__54_), .S(u4_sll_481_n66), .Z(
        u4_sll_481_ML_int_2__56_) );
  MUX2_X2 u4_sll_481_M1_2_4 ( .A(u4_sll_481_ML_int_2__4_), .B(u4_sll_481_n83), 
        .S(u4_sll_481_n78), .Z(u4_sll_481_ML_int_3__4_) );
  MUX2_X2 u4_sll_481_M1_2_5 ( .A(u4_sll_481_ML_int_2__5_), .B(
        u4_sll_481_ML_int_2__1_), .S(u4_sll_481_n78), .Z(
        u4_sll_481_ML_int_3__5_) );
  MUX2_X2 u4_sll_481_M1_2_6 ( .A(u4_sll_481_ML_int_2__6_), .B(
        u4_sll_481_ML_int_2__2_), .S(u4_sll_481_n78), .Z(
        u4_sll_481_ML_int_3__6_) );
  MUX2_X2 u4_sll_481_M1_2_7 ( .A(u4_sll_481_n14), .B(u4_sll_481_ML_int_2__3_), 
        .S(u4_sll_481_n78), .Z(u4_sll_481_ML_int_3__7_) );
  MUX2_X2 u4_sll_481_M1_2_8 ( .A(u4_sll_481_ML_int_2__8_), .B(
        u4_sll_481_ML_int_2__4_), .S(u4_sll_481_n78), .Z(
        u4_sll_481_ML_int_3__8_) );
  MUX2_X2 u4_sll_481_M1_2_12 ( .A(u4_sll_481_ML_int_2__12_), .B(
        u4_sll_481_ML_int_2__8_), .S(u4_sll_481_n78), .Z(
        u4_sll_481_ML_int_3__12_) );
  MUX2_X2 u4_sll_481_M1_2_14 ( .A(u4_sll_481_ML_int_2__14_), .B(
        u4_sll_481_ML_int_2__10_), .S(u4_sll_481_n77), .Z(
        u4_sll_481_ML_int_3__14_) );
  MUX2_X2 u4_sll_481_M1_2_17 ( .A(u4_sll_481_ML_int_2__17_), .B(
        u4_sll_481_ML_int_2__13_), .S(u4_sll_481_n77), .Z(
        u4_sll_481_ML_int_3__17_) );
  MUX2_X2 u4_sll_481_M1_2_18 ( .A(u4_sll_481_ML_int_2__18_), .B(
        u4_sll_481_ML_int_2__14_), .S(u4_sll_481_n77), .Z(
        u4_sll_481_ML_int_3__18_) );
  MUX2_X2 u4_sll_481_M1_2_19 ( .A(u4_sll_481_ML_int_2__19_), .B(
        u4_sll_481_ML_int_2__15_), .S(u4_sll_481_n77), .Z(
        u4_sll_481_ML_int_3__19_) );
  MUX2_X2 u4_sll_481_M1_2_20 ( .A(u4_sll_481_ML_int_2__20_), .B(
        u4_sll_481_ML_int_2__16_), .S(u4_sll_481_n77), .Z(
        u4_sll_481_ML_int_3__20_) );
  MUX2_X2 u4_sll_481_M1_2_21 ( .A(u4_sll_481_ML_int_2__21_), .B(
        u4_sll_481_ML_int_2__17_), .S(u4_sll_481_n77), .Z(
        u4_sll_481_ML_int_3__21_) );
  MUX2_X2 u4_sll_481_M1_2_22 ( .A(u4_sll_481_ML_int_2__22_), .B(
        u4_sll_481_ML_int_2__18_), .S(u4_sll_481_n77), .Z(
        u4_sll_481_ML_int_3__22_) );
  MUX2_X2 u4_sll_481_M1_2_23 ( .A(u4_sll_481_ML_int_2__23_), .B(
        u4_sll_481_ML_int_2__19_), .S(u4_sll_481_n77), .Z(
        u4_sll_481_ML_int_3__23_) );
  MUX2_X2 u4_sll_481_M1_2_24 ( .A(u4_sll_481_ML_int_2__24_), .B(
        u4_sll_481_ML_int_2__20_), .S(u4_sll_481_n76), .Z(
        u4_sll_481_ML_int_3__24_) );
  MUX2_X2 u4_sll_481_M1_2_27 ( .A(u4_sll_481_ML_int_2__27_), .B(
        u4_sll_481_ML_int_2__23_), .S(u4_sll_481_n76), .Z(
        u4_sll_481_ML_int_3__27_) );
  MUX2_X2 u4_sll_481_M1_2_28 ( .A(u4_sll_481_ML_int_2__28_), .B(
        u4_sll_481_ML_int_2__24_), .S(u4_sll_481_n76), .Z(
        u4_sll_481_ML_int_3__28_) );
  MUX2_X2 u4_sll_481_M1_2_30 ( .A(u4_sll_481_ML_int_2__30_), .B(
        u4_sll_481_ML_int_2__26_), .S(u4_sll_481_n76), .Z(
        u4_sll_481_ML_int_3__30_) );
  MUX2_X2 u4_sll_481_M1_2_34 ( .A(u4_sll_481_ML_int_2__34_), .B(
        u4_sll_481_ML_int_2__30_), .S(u4_sll_481_n76), .Z(
        u4_sll_481_ML_int_3__34_) );
  MUX2_X2 u4_sll_481_M1_2_35 ( .A(u4_sll_481_ML_int_2__35_), .B(
        u4_sll_481_ML_int_2__31_), .S(u4_sll_481_n75), .Z(
        u4_sll_481_ML_int_3__35_) );
  MUX2_X2 u4_sll_481_M1_2_36 ( .A(u4_sll_481_ML_int_2__36_), .B(
        u4_sll_481_ML_int_2__32_), .S(u4_sll_481_n75), .Z(
        u4_sll_481_ML_int_3__36_) );
  MUX2_X2 u4_sll_481_M1_2_37 ( .A(u4_sll_481_ML_int_2__37_), .B(
        u4_sll_481_ML_int_2__33_), .S(u4_sll_481_n75), .Z(
        u4_sll_481_ML_int_3__37_) );
  MUX2_X2 u4_sll_481_M1_2_38 ( .A(u4_sll_481_ML_int_2__38_), .B(
        u4_sll_481_ML_int_2__34_), .S(u4_sll_481_n75), .Z(
        u4_sll_481_ML_int_3__38_) );
  MUX2_X2 u4_sll_481_M1_2_39 ( .A(u4_sll_481_ML_int_2__39_), .B(
        u4_sll_481_ML_int_2__35_), .S(u4_sll_481_n75), .Z(
        u4_sll_481_ML_int_3__39_) );
  MUX2_X2 u4_sll_481_M1_2_41 ( .A(u4_sll_481_ML_int_2__41_), .B(
        u4_sll_481_ML_int_2__37_), .S(u4_sll_481_n75), .Z(
        u4_sll_481_ML_int_3__41_) );
  MUX2_X2 u4_sll_481_M1_2_42 ( .A(u4_sll_481_ML_int_2__42_), .B(
        u4_sll_481_ML_int_2__38_), .S(u4_sll_481_n75), .Z(
        u4_sll_481_ML_int_3__42_) );
  MUX2_X2 u4_sll_481_M1_2_43 ( .A(u4_sll_481_ML_int_2__43_), .B(
        u4_sll_481_ML_int_2__39_), .S(u4_sll_481_n75), .Z(
        u4_sll_481_ML_int_3__43_) );
  MUX2_X2 u4_sll_481_M1_2_45 ( .A(u4_sll_481_ML_int_2__45_), .B(
        u4_sll_481_ML_int_2__41_), .S(u4_sll_481_n75), .Z(
        u4_sll_481_ML_int_3__45_) );
  MUX2_X2 u4_sll_481_M1_2_46 ( .A(u4_sll_481_ML_int_2__46_), .B(
        u4_sll_481_ML_int_2__42_), .S(u4_sll_481_n74), .Z(
        u4_sll_481_ML_int_3__46_) );
  MUX2_X2 u4_sll_481_M1_2_48 ( .A(u4_sll_481_ML_int_2__48_), .B(
        u4_sll_481_ML_int_2__44_), .S(u4_sll_481_n74), .Z(
        u4_sll_481_ML_int_3__48_) );
  MUX2_X2 u4_sll_481_M1_2_49 ( .A(u4_sll_481_ML_int_2__49_), .B(
        u4_sll_481_ML_int_2__45_), .S(u4_sll_481_n74), .Z(
        u4_sll_481_ML_int_3__49_) );
  MUX2_X2 u4_sll_481_M1_2_50 ( .A(u4_sll_481_ML_int_2__50_), .B(
        u4_sll_481_ML_int_2__46_), .S(u4_sll_481_n74), .Z(
        u4_sll_481_ML_int_3__50_) );
  MUX2_X2 u4_sll_481_M1_2_51 ( .A(u4_sll_481_ML_int_2__51_), .B(
        u4_sll_481_ML_int_2__47_), .S(u4_sll_481_n74), .Z(
        u4_sll_481_ML_int_3__51_) );
  MUX2_X2 u4_sll_481_M1_2_52 ( .A(u4_sll_481_ML_int_2__52_), .B(
        u4_sll_481_ML_int_2__48_), .S(u4_sll_481_n74), .Z(
        u4_sll_481_ML_int_3__52_) );
  MUX2_X2 u4_sll_481_M1_2_53 ( .A(u4_sll_481_ML_int_2__53_), .B(
        u4_sll_481_ML_int_2__49_), .S(u4_sll_481_n74), .Z(
        u4_sll_481_ML_int_3__53_) );
  MUX2_X2 u4_sll_481_M1_2_54 ( .A(u4_sll_481_ML_int_2__54_), .B(
        u4_sll_481_ML_int_2__50_), .S(u4_sll_481_n74), .Z(
        u4_sll_481_ML_int_3__54_) );
  MUX2_X2 u4_sll_481_M1_2_55 ( .A(u4_sll_481_ML_int_2__55_), .B(
        u4_sll_481_ML_int_2__51_), .S(u4_sll_481_n74), .Z(
        u4_sll_481_ML_int_3__55_) );
  MUX2_X2 u4_sll_481_M1_2_56 ( .A(u4_sll_481_ML_int_2__56_), .B(
        u4_sll_481_ML_int_2__52_), .S(u4_sll_481_n74), .Z(
        u4_sll_481_ML_int_3__56_) );
  MUX2_X2 u4_sll_481_M1_3_8 ( .A(u4_sll_481_ML_int_3__8_), .B(
        u4_sll_481_ML_int_3__0_), .S(u4_sll_481_n81), .Z(
        u4_sll_481_ML_int_4__8_) );
  MUX2_X2 u4_sll_481_M1_3_17 ( .A(u4_sll_481_ML_int_3__17_), .B(
        u4_sll_481_ML_int_3__9_), .S(u4_sll_481_n81), .Z(
        u4_sll_481_ML_int_4__17_) );
  MUX2_X2 u4_sll_481_M1_3_19 ( .A(u4_sll_481_ML_int_3__19_), .B(
        u4_sll_481_ML_int_3__11_), .S(u4_sll_481_n80), .Z(
        u4_sll_481_ML_int_4__19_) );
  MUX2_X2 u4_sll_481_M1_3_20 ( .A(u4_sll_481_ML_int_3__20_), .B(
        u4_sll_481_ML_int_3__12_), .S(u4_sll_481_n80), .Z(
        u4_sll_481_ML_int_4__20_) );
  MUX2_X2 u4_sll_481_M1_3_21 ( .A(u4_sll_481_ML_int_3__21_), .B(
        u4_sll_481_ML_int_3__13_), .S(u4_sll_481_n80), .Z(
        u4_sll_481_ML_int_4__21_) );
  MUX2_X2 u4_sll_481_M1_3_22 ( .A(u4_sll_481_ML_int_3__22_), .B(
        u4_sll_481_ML_int_3__14_), .S(u4_sll_481_n80), .Z(
        u4_sll_481_ML_int_4__22_) );
  MUX2_X2 u4_sll_481_M1_3_23 ( .A(u4_sll_481_ML_int_3__23_), .B(
        u4_sll_481_ML_int_3__15_), .S(u4_sll_481_n80), .Z(
        u4_sll_481_ML_int_4__23_) );
  MUX2_X2 u4_sll_481_M1_3_24 ( .A(u4_sll_481_ML_int_3__24_), .B(
        u4_sll_481_ML_int_3__16_), .S(u4_sll_481_n80), .Z(
        u4_sll_481_ML_int_4__24_) );
  MUX2_X2 u4_sll_481_M1_3_35 ( .A(u4_sll_481_ML_int_3__35_), .B(
        u4_sll_481_ML_int_3__27_), .S(u4_sll_481_n80), .Z(
        u4_sll_481_ML_int_4__35_) );
  MUX2_X2 u4_sll_481_M1_3_36 ( .A(u4_sll_481_ML_int_3__36_), .B(
        u4_sll_481_ML_int_3__28_), .S(u4_sll_481_n80), .Z(
        u4_sll_481_ML_int_4__36_) );
  MUX2_X2 u4_sll_481_M1_3_38 ( .A(u4_sll_481_ML_int_3__38_), .B(
        u4_sll_481_ML_int_3__30_), .S(u4_sll_481_n81), .Z(
        u4_sll_481_ML_int_4__38_) );
  MUX2_X2 u4_sll_481_M1_3_49 ( .A(u4_sll_481_ML_int_3__49_), .B(
        u4_sll_481_ML_int_3__41_), .S(u4_sll_481_n80), .Z(
        u4_sll_481_ML_int_4__49_) );
  MUX2_X2 u4_sll_481_M1_3_50 ( .A(u4_sll_481_ML_int_3__50_), .B(
        u4_sll_481_ML_int_3__42_), .S(u4_sll_481_n81), .Z(
        u4_sll_481_ML_int_4__50_) );
  MUX2_X2 u4_sll_481_M1_3_51 ( .A(u4_sll_481_ML_int_3__51_), .B(
        u4_sll_481_ML_int_3__43_), .S(u4_sll_481_n80), .Z(
        u4_sll_481_ML_int_4__51_) );
  MUX2_X2 u4_sll_481_M1_3_52 ( .A(u4_sll_481_ML_int_3__52_), .B(
        u4_sll_481_ML_int_3__44_), .S(u4_sll_481_n80), .Z(
        u4_sll_481_ML_int_4__52_) );
  MUX2_X2 u4_sll_481_M1_3_53 ( .A(u4_sll_481_ML_int_3__53_), .B(
        u4_sll_481_ML_int_3__45_), .S(u4_sll_481_n81), .Z(
        u4_sll_481_ML_int_4__53_) );
  MUX2_X2 u4_sll_481_M1_3_54 ( .A(u4_sll_481_ML_int_3__54_), .B(
        u4_sll_481_ML_int_3__46_), .S(u4_sll_481_n80), .Z(
        u4_sll_481_ML_int_4__54_) );
  MUX2_X2 u4_sll_481_M1_3_56 ( .A(u4_sll_481_ML_int_3__56_), .B(
        u4_sll_481_ML_int_3__48_), .S(u4_sll_481_n80), .Z(
        u4_sll_481_ML_int_4__56_) );
  MUX2_X2 u4_sll_481_M1_4_17 ( .A(u4_sll_481_ML_int_4__17_), .B(
        u4_sll_481_ML_int_4__1_), .S(u4_sll_481_n84), .Z(
        u4_sll_481_ML_int_5__17_) );
  MUX2_X2 u4_sll_481_M1_4_18 ( .A(u4_sll_481_ML_int_4__18_), .B(
        u4_sll_481_ML_int_4__2_), .S(u4_sll_481_n84), .Z(
        u4_sll_481_ML_int_5__18_) );
  MUX2_X2 u4_sll_481_M1_4_19 ( .A(u4_sll_481_ML_int_4__19_), .B(
        u4_sll_481_ML_int_4__3_), .S(u4_sll_481_n84), .Z(
        u4_sll_481_ML_int_5__19_) );
  MUX2_X2 u4_sll_481_M1_4_20 ( .A(u4_sll_481_ML_int_4__20_), .B(
        u4_sll_481_ML_int_4__4_), .S(u4_sll_481_n84), .Z(
        u4_sll_481_ML_int_5__20_) );
  MUX2_X2 u4_sll_481_M1_4_21 ( .A(u4_sll_481_ML_int_4__21_), .B(
        u4_sll_481_ML_int_4__5_), .S(u4_sll_481_n84), .Z(
        u4_sll_481_ML_int_5__21_) );
  MUX2_X2 u4_sll_481_M1_4_22 ( .A(u4_sll_481_ML_int_4__22_), .B(
        u4_sll_481_ML_int_4__6_), .S(u4_sll_481_n84), .Z(
        u4_sll_481_ML_int_5__22_) );
  MUX2_X2 u4_sll_481_M1_4_23 ( .A(u4_sll_481_ML_int_4__23_), .B(
        u4_sll_481_ML_int_4__7_), .S(u4_sll_481_n84), .Z(
        u4_sll_481_ML_int_5__23_) );
  MUX2_X2 u4_sll_481_M1_4_24 ( .A(u4_sll_481_ML_int_4__24_), .B(
        u4_sll_481_ML_int_4__8_), .S(u4_sll_481_n84), .Z(
        u4_sll_481_ML_int_5__24_) );
  MUX2_X2 u4_sll_481_M1_4_49 ( .A(u4_sll_481_ML_int_4__49_), .B(
        u4_sll_481_ML_int_4__33_), .S(u4_sll_481_n84), .Z(
        u4_sll_481_ML_int_5__49_) );
  MUX2_X2 u4_sll_481_M1_4_50 ( .A(u4_sll_481_ML_int_4__50_), .B(
        u4_sll_481_ML_int_4__34_), .S(u4_sll_481_n84), .Z(
        u4_sll_481_ML_int_5__50_) );
  MUX2_X2 u4_sll_481_M1_4_51 ( .A(u4_sll_481_ML_int_4__51_), .B(
        u4_sll_481_ML_int_4__35_), .S(u4_sll_481_n84), .Z(
        u4_sll_481_ML_int_5__51_) );
  MUX2_X2 u4_sll_481_M1_4_52 ( .A(u4_sll_481_ML_int_4__52_), .B(
        u4_sll_481_ML_int_4__36_), .S(u4_sll_481_n84), .Z(
        u4_sll_481_ML_int_5__52_) );
  MUX2_X2 u4_sll_481_M1_4_53 ( .A(u4_sll_481_ML_int_4__53_), .B(
        u4_sll_481_ML_int_4__37_), .S(u4_sll_481_n84), .Z(
        u4_sll_481_ML_int_5__53_) );
  MUX2_X2 u4_sll_481_M1_4_54 ( .A(u4_sll_481_ML_int_4__54_), .B(
        u4_sll_481_ML_int_4__38_), .S(u4_sll_481_n84), .Z(
        u4_sll_481_ML_int_5__54_) );
  MUX2_X2 u4_sll_481_M1_5_54 ( .A(u4_sll_481_ML_int_5__54_), .B(
        u4_sll_481_ML_int_5__22_), .S(u4_sll_481_n85), .Z(
        u4_sll_481_ML_int_6__54_) );
  INV_X4 u4_sub_411_U19 ( .A(net85937), .ZN(u4_sub_411_n15) );
  INV_X4 u4_sub_411_U18 ( .A(net85933), .ZN(u4_sub_411_n14) );
  INV_X4 u4_sub_411_U17 ( .A(net85929), .ZN(u4_sub_411_n13) );
  INV_X4 u4_sub_411_U16 ( .A(n3085), .ZN(u4_sub_411_n12) );
  INV_X4 u4_sub_411_U15 ( .A(n3088), .ZN(u4_sub_411_n11) );
  INV_X4 u4_sub_411_U14 ( .A(n3089), .ZN(u4_sub_411_n10) );
  INV_X4 u4_sub_411_U13 ( .A(net85905), .ZN(u4_sub_411_n8) );
  INV_X4 u4_sub_411_U12 ( .A(u4_sub_411_n7), .ZN(u4_sub_411_carry_6_) );
  NAND2_X2 u4_sub_411_U11 ( .A1(u4_sub_411_n13), .A2(u4_sub_411_carry_5_), 
        .ZN(u4_sub_411_n7) );
  INV_X4 u4_sub_411_U10 ( .A(u4_sub_411_n6), .ZN(u4_sub_411_carry_7_) );
  NAND2_X2 u4_sub_411_U9 ( .A1(u4_sub_411_n14), .A2(u4_sub_411_carry_6_), .ZN(
        u4_sub_411_n6) );
  INV_X4 u4_sub_411_U8 ( .A(div_opa_ldz_r2[0]), .ZN(u4_sub_411_n5) );
  INV_X4 u4_sub_411_U7 ( .A(u4_sub_411_n8), .ZN(u4_sub_411_n4) );
  XNOR2_X2 u4_sub_411_U6 ( .A(u4_sub_411_n8), .B(div_opa_ldz_r2[0]), .ZN(
        u4_div_shft4[0]) );
  NAND2_X2 u4_sub_411_U5 ( .A1(u4_sub_411_n4), .A2(u4_sub_411_n5), .ZN(
        u4_sub_411_carry_1_) );
  INV_X1 u4_sub_411_U4 ( .A(n3091), .ZN(u4_sub_411_n9) );
  XOR2_X1 u4_sub_411_U3 ( .A(u4_sub_411_n15), .B(u4_sub_411_carry_7_), .Z(
        u4_div_shft4[7]) );
  XOR2_X1 u4_sub_411_U2 ( .A(u4_sub_411_n14), .B(u4_sub_411_carry_6_), .Z(
        u4_div_shft4[6]) );
  XOR2_X1 u4_sub_411_U1 ( .A(u4_sub_411_n13), .B(u4_sub_411_carry_5_), .Z(
        u4_div_shft4[5]) );
  FA_X1 u4_sub_411_U2_1 ( .A(div_opa_ldz_r2[1]), .B(u4_sub_411_n9), .CI(
        u4_sub_411_carry_1_), .CO(u4_sub_411_carry_2_), .S(u4_div_shft4[1]) );
  FA_X1 u4_sub_411_U2_2 ( .A(div_opa_ldz_r2[2]), .B(u4_sub_411_n10), .CI(
        u4_sub_411_carry_2_), .CO(u4_sub_411_carry_3_), .S(u4_div_shft4[2]) );
  FA_X1 u4_sub_411_U2_3 ( .A(div_opa_ldz_r2[3]), .B(u4_sub_411_n11), .CI(
        u4_sub_411_carry_3_), .CO(u4_sub_411_carry_4_), .S(u4_div_shft4[3]) );
  FA_X1 u4_sub_411_U2_4 ( .A(div_opa_ldz_r2[4]), .B(u4_sub_411_n12), .CI(
        u4_sub_411_carry_4_), .CO(u4_sub_411_carry_5_), .S(u4_div_shft4[4]) );
  INV_X4 u4_add_410_U13 ( .A(u4_add_410_n7), .ZN(u4_div_shft3_0_) );
  INV_X4 u4_add_410_U12 ( .A(u4_add_410_n6), .ZN(u4_add_410_carry_1_) );
  NAND2_X2 u4_add_410_U11 ( .A1(net85905), .A2(div_opa_ldz_r2[0]), .ZN(
        u4_add_410_n6) );
  INV_X4 u4_add_410_U10 ( .A(u4_add_410_n5), .ZN(u4_add_410_carry_6_) );
  NAND2_X2 u4_add_410_U9 ( .A1(net85929), .A2(u4_add_410_carry_5_), .ZN(
        u4_add_410_n5) );
  INV_X4 u4_add_410_U8 ( .A(u4_add_410_n4), .ZN(u4_div_shft3_6_) );
  XNOR2_X2 u4_add_410_U7 ( .A(net85933), .B(u4_add_410_carry_6_), .ZN(
        u4_add_410_n4) );
  INV_X4 u4_add_410_U6 ( .A(u4_add_410_n3), .ZN(u4_add_410_carry_7_) );
  NAND2_X2 u4_add_410_U5 ( .A1(net85933), .A2(u4_add_410_carry_6_), .ZN(
        u4_add_410_n3) );
  INV_X4 u4_add_410_U4 ( .A(u4_add_410_n2), .ZN(u4_div_shft3_7_) );
  XNOR2_X2 u4_add_410_U3 ( .A(net85937), .B(u4_add_410_carry_7_), .ZN(
        u4_add_410_n2) );
  XNOR2_X1 u4_add_410_U2 ( .A(net85905), .B(div_opa_ldz_r2[0]), .ZN(
        u4_add_410_n7) );
  XOR2_X1 u4_add_410_U1 ( .A(net85929), .B(u4_add_410_carry_5_), .Z(
        u4_div_shft3_5_) );
  FA_X1 u4_add_410_U1_1 ( .A(div_opa_ldz_r2[1]), .B(n3091), .CI(
        u4_add_410_carry_1_), .CO(u4_add_410_carry_2_), .S(u4_div_shft3_1_) );
  FA_X1 u4_add_410_U1_2 ( .A(div_opa_ldz_r2[2]), .B(n3089), .CI(
        u4_add_410_carry_2_), .CO(u4_add_410_carry_3_), .S(u4_div_shft3_2_) );
  FA_X1 u4_add_410_U1_3 ( .A(div_opa_ldz_r2[3]), .B(n3087), .CI(
        u4_add_410_carry_3_), .CO(u4_add_410_carry_4_), .S(u4_div_shft3_3_) );
  FA_X1 u4_add_410_U1_4 ( .A(div_opa_ldz_r2[4]), .B(n3085), .CI(
        u4_add_410_carry_4_), .CO(u4_add_410_carry_5_), .S(u4_div_shft3_4_) );
  INV_X4 u3_sub_60_U32 ( .A(fractb[26]), .ZN(u3_sub_60_n30) );
  INV_X4 u3_sub_60_U31 ( .A(fractb[25]), .ZN(u3_sub_60_n29) );
  INV_X4 u3_sub_60_U30 ( .A(fractb[24]), .ZN(u3_sub_60_n28) );
  INV_X4 u3_sub_60_U29 ( .A(fractb[23]), .ZN(u3_sub_60_n27) );
  INV_X4 u3_sub_60_U28 ( .A(fractb[22]), .ZN(u3_sub_60_n26) );
  INV_X4 u3_sub_60_U27 ( .A(fractb[21]), .ZN(u3_sub_60_n25) );
  INV_X4 u3_sub_60_U26 ( .A(fractb[20]), .ZN(u3_sub_60_n24) );
  INV_X4 u3_sub_60_U25 ( .A(fractb[19]), .ZN(u3_sub_60_n23) );
  INV_X4 u3_sub_60_U24 ( .A(fractb[18]), .ZN(u3_sub_60_n22) );
  INV_X4 u3_sub_60_U23 ( .A(fractb[17]), .ZN(u3_sub_60_n21) );
  INV_X4 u3_sub_60_U22 ( .A(fractb[16]), .ZN(u3_sub_60_n20) );
  INV_X4 u3_sub_60_U21 ( .A(fractb[15]), .ZN(u3_sub_60_n19) );
  INV_X4 u3_sub_60_U20 ( .A(fractb[14]), .ZN(u3_sub_60_n18) );
  INV_X4 u3_sub_60_U19 ( .A(fractb[13]), .ZN(u3_sub_60_n17) );
  INV_X4 u3_sub_60_U18 ( .A(fractb[12]), .ZN(u3_sub_60_n16) );
  INV_X4 u3_sub_60_U17 ( .A(fractb[11]), .ZN(u3_sub_60_n15) );
  INV_X4 u3_sub_60_U16 ( .A(fractb[10]), .ZN(u3_sub_60_n14) );
  INV_X4 u3_sub_60_U15 ( .A(fractb[9]), .ZN(u3_sub_60_n13) );
  INV_X4 u3_sub_60_U14 ( .A(fractb[8]), .ZN(u3_sub_60_n12) );
  INV_X4 u3_sub_60_U13 ( .A(fractb[7]), .ZN(u3_sub_60_n11) );
  INV_X4 u3_sub_60_U12 ( .A(fractb[6]), .ZN(u3_sub_60_n10) );
  INV_X4 u3_sub_60_U11 ( .A(fractb[5]), .ZN(u3_sub_60_n9) );
  INV_X4 u3_sub_60_U10 ( .A(fractb[4]), .ZN(u3_sub_60_n8) );
  INV_X4 u3_sub_60_U9 ( .A(fractb[3]), .ZN(u3_sub_60_n7) );
  INV_X4 u3_sub_60_U8 ( .A(fractb[2]), .ZN(u3_sub_60_n6) );
  INV_X4 u3_sub_60_U7 ( .A(fractb[1]), .ZN(u3_sub_60_n5) );
  INV_X4 u3_sub_60_U6 ( .A(u3_sub_60_carry[27]), .ZN(u3_N58) );
  INV_X4 u3_sub_60_U5 ( .A(u3_sub_60_n4), .ZN(u3_sub_60_n1) );
  NAND2_X2 u3_sub_60_U4 ( .A1(u3_sub_60_n1), .A2(u3_sub_60_n2), .ZN(
        u3_sub_60_carry[1]) );
  XNOR2_X1 u3_sub_60_U3 ( .A(u3_sub_60_n4), .B(fracta[0]), .ZN(u3_N31) );
  INV_X2 u3_sub_60_U2 ( .A(fracta[0]), .ZN(u3_sub_60_n2) );
  INV_X1 u3_sub_60_U1 ( .A(fractb[0]), .ZN(u3_sub_60_n4) );
  FA_X1 u3_sub_60_U2_1 ( .A(fracta[1]), .B(u3_sub_60_n5), .CI(
        u3_sub_60_carry[1]), .CO(u3_sub_60_carry[2]), .S(u3_N32) );
  FA_X1 u3_sub_60_U2_2 ( .A(fracta[2]), .B(u3_sub_60_n6), .CI(
        u3_sub_60_carry[2]), .CO(u3_sub_60_carry[3]), .S(u3_N33) );
  FA_X1 u3_sub_60_U2_3 ( .A(fracta[3]), .B(u3_sub_60_n7), .CI(
        u3_sub_60_carry[3]), .CO(u3_sub_60_carry[4]), .S(u3_N34) );
  FA_X1 u3_sub_60_U2_4 ( .A(fracta[4]), .B(u3_sub_60_n8), .CI(
        u3_sub_60_carry[4]), .CO(u3_sub_60_carry[5]), .S(u3_N35) );
  FA_X1 u3_sub_60_U2_5 ( .A(fracta[5]), .B(u3_sub_60_n9), .CI(
        u3_sub_60_carry[5]), .CO(u3_sub_60_carry[6]), .S(u3_N36) );
  FA_X1 u3_sub_60_U2_6 ( .A(fracta[6]), .B(u3_sub_60_n10), .CI(
        u3_sub_60_carry[6]), .CO(u3_sub_60_carry[7]), .S(u3_N37) );
  FA_X1 u3_sub_60_U2_7 ( .A(fracta[7]), .B(u3_sub_60_n11), .CI(
        u3_sub_60_carry[7]), .CO(u3_sub_60_carry[8]), .S(u3_N38) );
  FA_X1 u3_sub_60_U2_8 ( .A(fracta[8]), .B(u3_sub_60_n12), .CI(
        u3_sub_60_carry[8]), .CO(u3_sub_60_carry[9]), .S(u3_N39) );
  FA_X1 u3_sub_60_U2_9 ( .A(fracta[9]), .B(u3_sub_60_n13), .CI(
        u3_sub_60_carry[9]), .CO(u3_sub_60_carry[10]), .S(u3_N40) );
  FA_X1 u3_sub_60_U2_10 ( .A(fracta[10]), .B(u3_sub_60_n14), .CI(
        u3_sub_60_carry[10]), .CO(u3_sub_60_carry[11]), .S(u3_N41) );
  FA_X1 u3_sub_60_U2_11 ( .A(fracta[11]), .B(u3_sub_60_n15), .CI(
        u3_sub_60_carry[11]), .CO(u3_sub_60_carry[12]), .S(u3_N42) );
  FA_X1 u3_sub_60_U2_12 ( .A(fracta[12]), .B(u3_sub_60_n16), .CI(
        u3_sub_60_carry[12]), .CO(u3_sub_60_carry[13]), .S(u3_N43) );
  FA_X1 u3_sub_60_U2_13 ( .A(fracta[13]), .B(u3_sub_60_n17), .CI(
        u3_sub_60_carry[13]), .CO(u3_sub_60_carry[14]), .S(u3_N44) );
  FA_X1 u3_sub_60_U2_14 ( .A(fracta[14]), .B(u3_sub_60_n18), .CI(
        u3_sub_60_carry[14]), .CO(u3_sub_60_carry[15]), .S(u3_N45) );
  FA_X1 u3_sub_60_U2_15 ( .A(fracta[15]), .B(u3_sub_60_n19), .CI(
        u3_sub_60_carry[15]), .CO(u3_sub_60_carry[16]), .S(u3_N46) );
  FA_X1 u3_sub_60_U2_16 ( .A(fracta[16]), .B(u3_sub_60_n20), .CI(
        u3_sub_60_carry[16]), .CO(u3_sub_60_carry[17]), .S(u3_N47) );
  FA_X1 u3_sub_60_U2_17 ( .A(fracta[17]), .B(u3_sub_60_n21), .CI(
        u3_sub_60_carry[17]), .CO(u3_sub_60_carry[18]), .S(u3_N48) );
  FA_X1 u3_sub_60_U2_18 ( .A(fracta[18]), .B(u3_sub_60_n22), .CI(
        u3_sub_60_carry[18]), .CO(u3_sub_60_carry[19]), .S(u3_N49) );
  FA_X1 u3_sub_60_U2_19 ( .A(fracta[19]), .B(u3_sub_60_n23), .CI(
        u3_sub_60_carry[19]), .CO(u3_sub_60_carry[20]), .S(u3_N50) );
  FA_X1 u3_sub_60_U2_20 ( .A(fracta[20]), .B(u3_sub_60_n24), .CI(
        u3_sub_60_carry[20]), .CO(u3_sub_60_carry[21]), .S(u3_N51) );
  FA_X1 u3_sub_60_U2_21 ( .A(fracta[21]), .B(u3_sub_60_n25), .CI(
        u3_sub_60_carry[21]), .CO(u3_sub_60_carry[22]), .S(u3_N52) );
  FA_X1 u3_sub_60_U2_22 ( .A(fracta[22]), .B(u3_sub_60_n26), .CI(
        u3_sub_60_carry[22]), .CO(u3_sub_60_carry[23]), .S(u3_N53) );
  FA_X1 u3_sub_60_U2_23 ( .A(fracta[23]), .B(u3_sub_60_n27), .CI(
        u3_sub_60_carry[23]), .CO(u3_sub_60_carry[24]), .S(u3_N54) );
  FA_X1 u3_sub_60_U2_24 ( .A(fracta[24]), .B(u3_sub_60_n28), .CI(
        u3_sub_60_carry[24]), .CO(u3_sub_60_carry[25]), .S(u3_N55) );
  FA_X1 u3_sub_60_U2_25 ( .A(fracta[25]), .B(u3_sub_60_n29), .CI(
        u3_sub_60_carry[25]), .CO(u3_sub_60_carry[26]), .S(u3_N56) );
  FA_X1 u3_sub_60_U2_26 ( .A(fracta[26]), .B(u3_sub_60_n30), .CI(
        u3_sub_60_carry[26]), .CO(u3_sub_60_carry[27]), .S(u3_N57) );
  INV_X4 u3_add_60_U5 ( .A(u3_add_60_n3), .ZN(u3_N3) );
  INV_X4 u3_add_60_U4 ( .A(u3_add_60_n2), .ZN(u3_add_60_carry[1]) );
  XNOR2_X1 u3_add_60_U3 ( .A(fractb[0]), .B(u3_add_60_n1), .ZN(u3_add_60_n3)
         );
  BUF_X32 u3_add_60_U2 ( .A(fracta[0]), .Z(u3_add_60_n1) );
  NAND2_X4 u3_add_60_U1 ( .A1(fracta[0]), .A2(fractb[0]), .ZN(u3_add_60_n2) );
  FA_X1 u3_add_60_U1_1 ( .A(fracta[1]), .B(fractb[1]), .CI(u3_add_60_carry[1]), 
        .CO(u3_add_60_carry[2]), .S(u3_N4) );
  FA_X1 u3_add_60_U1_2 ( .A(fracta[2]), .B(fractb[2]), .CI(u3_add_60_carry[2]), 
        .CO(u3_add_60_carry[3]), .S(u3_N5) );
  FA_X1 u3_add_60_U1_3 ( .A(fracta[3]), .B(fractb[3]), .CI(u3_add_60_carry[3]), 
        .CO(u3_add_60_carry[4]), .S(u3_N6) );
  FA_X1 u3_add_60_U1_4 ( .A(fracta[4]), .B(fractb[4]), .CI(u3_add_60_carry[4]), 
        .CO(u3_add_60_carry[5]), .S(u3_N7) );
  FA_X1 u3_add_60_U1_5 ( .A(fracta[5]), .B(fractb[5]), .CI(u3_add_60_carry[5]), 
        .CO(u3_add_60_carry[6]), .S(u3_N8) );
  FA_X1 u3_add_60_U1_6 ( .A(fracta[6]), .B(fractb[6]), .CI(u3_add_60_carry[6]), 
        .CO(u3_add_60_carry[7]), .S(u3_N9) );
  FA_X1 u3_add_60_U1_7 ( .A(fracta[7]), .B(fractb[7]), .CI(u3_add_60_carry[7]), 
        .CO(u3_add_60_carry[8]), .S(u3_N10) );
  FA_X1 u3_add_60_U1_8 ( .A(fracta[8]), .B(fractb[8]), .CI(u3_add_60_carry[8]), 
        .CO(u3_add_60_carry[9]), .S(u3_N11) );
  FA_X1 u3_add_60_U1_9 ( .A(fracta[9]), .B(fractb[9]), .CI(u3_add_60_carry[9]), 
        .CO(u3_add_60_carry[10]), .S(u3_N12) );
  FA_X1 u3_add_60_U1_10 ( .A(fracta[10]), .B(fractb[10]), .CI(
        u3_add_60_carry[10]), .CO(u3_add_60_carry[11]), .S(u3_N13) );
  FA_X1 u3_add_60_U1_11 ( .A(fracta[11]), .B(fractb[11]), .CI(
        u3_add_60_carry[11]), .CO(u3_add_60_carry[12]), .S(u3_N14) );
  FA_X1 u3_add_60_U1_12 ( .A(fracta[12]), .B(fractb[12]), .CI(
        u3_add_60_carry[12]), .CO(u3_add_60_carry[13]), .S(u3_N15) );
  FA_X1 u3_add_60_U1_13 ( .A(fracta[13]), .B(fractb[13]), .CI(
        u3_add_60_carry[13]), .CO(u3_add_60_carry[14]), .S(u3_N16) );
  FA_X1 u3_add_60_U1_14 ( .A(fracta[14]), .B(fractb[14]), .CI(
        u3_add_60_carry[14]), .CO(u3_add_60_carry[15]), .S(u3_N17) );
  FA_X1 u3_add_60_U1_15 ( .A(fracta[15]), .B(fractb[15]), .CI(
        u3_add_60_carry[15]), .CO(u3_add_60_carry[16]), .S(u3_N18) );
  FA_X1 u3_add_60_U1_16 ( .A(fracta[16]), .B(fractb[16]), .CI(
        u3_add_60_carry[16]), .CO(u3_add_60_carry[17]), .S(u3_N19) );
  FA_X1 u3_add_60_U1_17 ( .A(fracta[17]), .B(fractb[17]), .CI(
        u3_add_60_carry[17]), .CO(u3_add_60_carry[18]), .S(u3_N20) );
  FA_X1 u3_add_60_U1_18 ( .A(fracta[18]), .B(fractb[18]), .CI(
        u3_add_60_carry[18]), .CO(u3_add_60_carry[19]), .S(u3_N21) );
  FA_X1 u3_add_60_U1_19 ( .A(fracta[19]), .B(fractb[19]), .CI(
        u3_add_60_carry[19]), .CO(u3_add_60_carry[20]), .S(u3_N22) );
  FA_X1 u3_add_60_U1_20 ( .A(fracta[20]), .B(fractb[20]), .CI(
        u3_add_60_carry[20]), .CO(u3_add_60_carry[21]), .S(u3_N23) );
  FA_X1 u3_add_60_U1_21 ( .A(fracta[21]), .B(fractb[21]), .CI(
        u3_add_60_carry[21]), .CO(u3_add_60_carry[22]), .S(u3_N24) );
  FA_X1 u3_add_60_U1_22 ( .A(fracta[22]), .B(fractb[22]), .CI(
        u3_add_60_carry[22]), .CO(u3_add_60_carry[23]), .S(u3_N25) );
  FA_X1 u3_add_60_U1_23 ( .A(fracta[23]), .B(fractb[23]), .CI(
        u3_add_60_carry[23]), .CO(u3_add_60_carry[24]), .S(u3_N26) );
  FA_X1 u3_add_60_U1_24 ( .A(fracta[24]), .B(fractb[24]), .CI(
        u3_add_60_carry[24]), .CO(u3_add_60_carry[25]), .S(u3_N27) );
  FA_X1 u3_add_60_U1_25 ( .A(fracta[25]), .B(fractb[25]), .CI(
        u3_add_60_carry[25]), .CO(u3_add_60_carry[26]), .S(u3_N28) );
  FA_X1 u3_add_60_U1_26 ( .A(fracta[26]), .B(fractb[26]), .CI(
        u3_add_60_carry[26]), .CO(u3_N30), .S(u3_N29) );
  XOR2_X1 u2_add_117_U2 ( .A(u2_add_117_carry[7]), .B(u2_exp_tmp4_7_), .Z(
        u2_N49) );
  INV_X4 u2_add_117_U1 ( .A(u2_exp_tmp4_0_), .ZN(u2_N42) );
  HA_X1 u2_add_117_U1_1_1 ( .A(u2_exp_tmp4_1_), .B(u2_exp_tmp4_0_), .CO(
        u2_add_117_carry[2]), .S(u2_N43) );
  HA_X1 u2_add_117_U1_1_2 ( .A(u2_exp_tmp4_2_), .B(u2_add_117_carry[2]), .CO(
        u2_add_117_carry[3]), .S(u2_N44) );
  HA_X1 u2_add_117_U1_1_3 ( .A(u2_exp_tmp4_3_), .B(u2_add_117_carry[3]), .CO(
        u2_add_117_carry[4]), .S(u2_N45) );
  HA_X1 u2_add_117_U1_1_4 ( .A(u2_exp_tmp4_4_), .B(u2_add_117_carry[4]), .CO(
        u2_add_117_carry[5]), .S(u2_N46) );
  HA_X1 u2_add_117_U1_1_5 ( .A(u2_exp_tmp4_5_), .B(u2_add_117_carry[5]), .CO(
        u2_add_117_carry[6]), .S(u2_N47) );
  HA_X1 u2_add_117_U1_1_6 ( .A(u2_exp_tmp4_6_), .B(u2_add_117_carry[6]), .CO(
        u2_add_117_carry[7]), .S(u2_N48) );
  XOR2_X1 u2_add_115_U2 ( .A(u2_add_115_carry[7]), .B(n5253), .Z(
        u2_exp_tmp3_7_) );
  INV_X4 u2_add_115_U1 ( .A(u2_exp_tmp4_0_), .ZN(u2_exp_tmp3_0_) );
  HA_X1 u2_add_115_U1_1_1 ( .A(n2716), .B(u2_exp_tmp4_0_), .CO(
        u2_add_115_carry[2]), .S(u2_exp_tmp3_1_) );
  HA_X1 u2_add_115_U1_1_2 ( .A(n5258), .B(u2_add_115_carry[2]), .CO(
        u2_add_115_carry[3]), .S(u2_exp_tmp3_2_) );
  HA_X1 u2_add_115_U1_1_3 ( .A(n5257), .B(u2_add_115_carry[3]), .CO(
        u2_add_115_carry[4]), .S(u2_exp_tmp3_3_) );
  HA_X1 u2_add_115_U1_1_4 ( .A(n5256), .B(u2_add_115_carry[4]), .CO(
        u2_add_115_carry[5]), .S(u2_exp_tmp3_4_) );
  HA_X1 u2_add_115_U1_1_5 ( .A(n5255), .B(u2_add_115_carry[5]), .CO(
        u2_add_115_carry[6]), .S(u2_exp_tmp3_5_) );
  HA_X1 u2_add_115_U1_1_6 ( .A(n5254), .B(u2_add_115_carry[6]), .CO(
        u2_add_115_carry[7]), .S(u2_exp_tmp3_6_) );
  INV_X4 u2_add_112_U3 ( .A(u2_add_112_n2), .ZN(u2_add_112_carry[1]) );
  NAND2_X2 u2_add_112_U2 ( .A1(opb_r[23]), .A2(opa_r[23]), .ZN(u2_add_112_n2)
         );
  XOR2_X1 u2_add_112_U1 ( .A(opb_r[23]), .B(opa_r[23]), .Z(u2_N15) );
  FA_X1 u2_add_112_U1_1 ( .A(opa_r[24]), .B(opb_r[24]), .CI(
        u2_add_112_carry[1]), .CO(u2_add_112_carry[2]), .S(u2_N16) );
  FA_X1 u2_add_112_U1_2 ( .A(opa_r[25]), .B(opb_r[25]), .CI(
        u2_add_112_carry[2]), .CO(u2_add_112_carry[3]), .S(u2_N17) );
  FA_X1 u2_add_112_U1_3 ( .A(opa_r[26]), .B(opb_r[26]), .CI(
        u2_add_112_carry[3]), .CO(u2_add_112_carry[4]), .S(u2_N18) );
  FA_X1 u2_add_112_U1_4 ( .A(opa_r[27]), .B(opb_r[27]), .CI(
        u2_add_112_carry[4]), .CO(u2_add_112_carry[5]), .S(u2_N19) );
  FA_X1 u2_add_112_U1_5 ( .A(opa_r[28]), .B(opb_r[28]), .CI(
        u2_add_112_carry[5]), .CO(u2_add_112_carry[6]), .S(u2_N20) );
  FA_X1 u2_add_112_U1_6 ( .A(opa_r[29]), .B(opb_r[29]), .CI(
        u2_add_112_carry[6]), .CO(u2_add_112_carry[7]), .S(u2_N21) );
  FA_X1 u2_add_112_U1_7 ( .A(opa_r[30]), .B(opb_r[30]), .CI(
        u2_add_112_carry[7]), .CO(u2_N23), .S(u2_N22) );
  INV_X4 u2_sub_112_U13 ( .A(opb_r[23]), .ZN(u2_sub_112_n11) );
  INV_X4 u2_sub_112_U12 ( .A(opb_r[25]), .ZN(u2_sub_112_n9) );
  INV_X4 u2_sub_112_U11 ( .A(opb_r[26]), .ZN(u2_sub_112_n8) );
  INV_X4 u2_sub_112_U10 ( .A(opb_r[28]), .ZN(u2_sub_112_n6) );
  INV_X4 u2_sub_112_U9 ( .A(opb_r[29]), .ZN(u2_sub_112_n5) );
  INV_X4 u2_sub_112_U8 ( .A(u2_sub_112_carry[8]), .ZN(u2_N14) );
  INV_X2 u2_sub_112_U7 ( .A(opb_r[27]), .ZN(u2_sub_112_n7) );
  INV_X1 u2_sub_112_U6 ( .A(opb_r[30]), .ZN(u2_sub_112_n4) );
  INV_X4 u2_sub_112_U5 ( .A(u2_sub_112_n11), .ZN(u2_sub_112_n1) );
  NAND2_X2 u2_sub_112_U4 ( .A1(u2_sub_112_n1), .A2(u2_sub_112_n2), .ZN(
        u2_sub_112_carry[1]) );
  XNOR2_X1 u2_sub_112_U3 ( .A(u2_sub_112_n11), .B(opa_r[23]), .ZN(u2_N6) );
  INV_X2 u2_sub_112_U2 ( .A(opa_r[23]), .ZN(u2_sub_112_n2) );
  INV_X2 u2_sub_112_U1 ( .A(opb_r[24]), .ZN(u2_sub_112_n10) );
  FA_X1 u2_sub_112_U2_1 ( .A(opa_r[24]), .B(u2_sub_112_n10), .CI(
        u2_sub_112_carry[1]), .CO(u2_sub_112_carry[2]), .S(u2_N7) );
  FA_X1 u2_sub_112_U2_2 ( .A(opa_r[25]), .B(u2_sub_112_n9), .CI(
        u2_sub_112_carry[2]), .CO(u2_sub_112_carry[3]), .S(u2_N8) );
  FA_X1 u2_sub_112_U2_3 ( .A(opa_r[26]), .B(u2_sub_112_n8), .CI(
        u2_sub_112_carry[3]), .CO(u2_sub_112_carry[4]), .S(u2_N9) );
  FA_X1 u2_sub_112_U2_4 ( .A(opa_r[27]), .B(u2_sub_112_n7), .CI(
        u2_sub_112_carry[4]), .CO(u2_sub_112_carry[5]), .S(u2_N10) );
  FA_X1 u2_sub_112_U2_5 ( .A(opa_r[28]), .B(u2_sub_112_n6), .CI(
        u2_sub_112_carry[5]), .CO(u2_sub_112_carry[6]), .S(u2_N11) );
  FA_X1 u2_sub_112_U2_6 ( .A(opa_r[29]), .B(u2_sub_112_n5), .CI(
        u2_sub_112_carry[6]), .CO(u2_sub_112_carry[7]), .S(u2_N12) );
  FA_X1 u2_sub_112_U2_7 ( .A(opa_r[30]), .B(u2_sub_112_n4), .CI(
        u2_sub_112_carry[7]), .CO(u2_sub_112_carry[8]), .S(u2_N13) );
  AOI22_X1 u1_srl_148_U174 ( .A1(n5297), .A2(u1_srl_148_n6), .B1(n5301), .B2(
        u1_srl_148_n3), .ZN(u1_srl_148_n147) );
  OAI221_X1 u1_srl_148_U173 ( .B1(u1_srl_148_n7), .B2(u1_srl_148_n46), .C1(
        u1_srl_148_n10), .C2(u1_srl_148_n45), .A(u1_srl_148_n147), .ZN(
        u1_srl_148_n146) );
  AOI22_X1 u1_srl_148_U172 ( .A1(u1_srl_148_n99), .A2(u1_adj_op_20_), .B1(
        u1_adj_op_17_), .B2(u1_srl_148_n4), .ZN(u1_srl_148_n145) );
  AND2_X1 u1_srl_148_U171 ( .A1(n5291), .A2(u1_srl_148_n20), .ZN(
        u1_srl_148_n119) );
  AOI222_X1 u1_srl_148_U170 ( .A1(u1_srl_148_n76), .A2(u1_srl_148_n111), .B1(
        u1_srl_148_n75), .B2(u1_srl_148_n119), .C1(u1_srl_148_n74), .C2(
        u1_srl_148_n110), .ZN(u1_srl_148_n120) );
  NAND2_X1 u1_srl_148_U169 ( .A1(n5291), .A2(u1_srl_148_n18), .ZN(
        u1_srl_148_n122) );
  AOI22_X1 u1_srl_148_U168 ( .A1(n5293), .A2(u1_srl_148_n99), .B1(n5296), .B2(
        u1_srl_148_n3), .ZN(u1_srl_148_n143) );
  OAI221_X1 u1_srl_148_U167 ( .B1(u1_srl_148_n8), .B2(u1_srl_148_n42), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n41), .A(u1_srl_148_n143), .ZN(
        u1_srl_148_n77) );
  AOI22_X1 u1_srl_148_U166 ( .A1(n5306), .A2(u1_srl_148_n5), .B1(n5292), .B2(
        u1_srl_148_n4), .ZN(u1_srl_148_n142) );
  NOR3_X1 u1_srl_148_U165 ( .A1(u1_srl_148_n61), .A2(u1_srl_148_n36), .A3(
        u1_srl_148_n64), .ZN(u1_srl_148_n141) );
  AOI221_X1 u1_srl_148_U164 ( .B1(u1_srl_148_n66), .B2(u1_srl_148_n77), .C1(
        u1_srl_148_n70), .C2(u1_srl_148_n92), .A(u1_srl_148_n141), .ZN(
        u1_srl_148_n140) );
  OAI221_X1 u1_srl_148_U163 ( .B1(u1_srl_148_n21), .B2(u1_srl_148_n63), .C1(
        u1_srl_148_n120), .C2(u1_srl_148_n18), .A(u1_srl_148_n140), .ZN(
        u1_adj_op_out_sft_0_) );
  AOI22_X1 u1_srl_148_U162 ( .A1(n5304), .A2(u1_srl_148_n6), .B1(n5307), .B2(
        u1_srl_148_n100), .ZN(u1_srl_148_n139) );
  OAI221_X1 u1_srl_148_U161 ( .B1(u1_srl_148_n8), .B2(u1_srl_148_n58), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n57), .A(u1_srl_148_n139), .ZN(
        u1_srl_148_n84) );
  AOI22_X1 u1_srl_148_U160 ( .A1(u1_adj_op_10_), .A2(u1_srl_148_n99), .B1(
        n5294), .B2(u1_srl_148_n3), .ZN(u1_srl_148_n138) );
  OAI221_X1 u1_srl_148_U159 ( .B1(u1_srl_148_n8), .B2(u1_srl_148_n40), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n39), .A(u1_srl_148_n138), .ZN(
        u1_srl_148_n105) );
  AOI22_X1 u1_srl_148_U158 ( .A1(u1_adj_op_18_), .A2(u1_srl_148_n5), .B1(n5303), .B2(u1_srl_148_n4), .ZN(u1_srl_148_n137) );
  OAI221_X1 u1_srl_148_U157 ( .B1(u1_srl_148_n8), .B2(u1_srl_148_n54), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n53), .A(u1_srl_148_n137), .ZN(
        u1_srl_148_n86) );
  NOR2_X1 u1_srl_148_U156 ( .A1(u1_srl_148_n22), .A2(u1_srl_148_n62), .ZN(
        u1_srl_148_n109) );
  AOI222_X1 u1_srl_148_U155 ( .A1(u1_srl_148_n66), .A2(u1_srl_148_n86), .B1(
        u1_srl_148_n109), .B2(u1_srl_148_n68), .C1(u1_srl_148_n70), .C2(
        u1_srl_148_n2), .ZN(u1_srl_148_n135) );
  OAI221_X1 u1_srl_148_U154 ( .B1(u1_srl_148_n26), .B2(u1_srl_148_n63), .C1(
        u1_srl_148_n27), .C2(u1_srl_148_n64), .A(u1_srl_148_n135), .ZN(
        u1_adj_op_out_sft_10_) );
  AOI22_X1 u1_srl_148_U153 ( .A1(u1_srl_148_n6), .A2(n2459), .B1(u1_adj_op_20_), .B2(u1_srl_148_n3), .ZN(u1_srl_148_n134) );
  AOI22_X1 u1_srl_148_U152 ( .A1(u1_srl_148_n99), .A2(u1_adj_op_19_), .B1(
        n5302), .B2(u1_srl_148_n4), .ZN(u1_srl_148_n133) );
  AOI22_X1 u1_srl_148_U151 ( .A1(n5303), .A2(u1_srl_148_n6), .B1(n5306), .B2(
        u1_srl_148_n100), .ZN(u1_srl_148_n132) );
  AOI22_X1 u1_srl_148_U150 ( .A1(n5307), .A2(u1_srl_148_n99), .B1(n5293), .B2(
        u1_srl_148_n3), .ZN(u1_srl_148_n131) );
  AOI22_X1 u1_srl_148_U149 ( .A1(u1_srl_148_n16), .A2(u1_srl_148_n79), .B1(
        u1_srl_148_n17), .B2(u1_srl_148_n82), .ZN(u1_srl_148_n130) );
  AOI221_X1 u1_srl_148_U148 ( .B1(u1_srl_148_n80), .B2(u1_srl_148_n70), .C1(
        u1_srl_148_n81), .C2(u1_srl_148_n66), .A(u1_srl_148_n14), .ZN(
        u1_srl_148_n129) );
  AOI22_X1 u1_srl_148_U147 ( .A1(u1_srl_148_n70), .A2(u1_srl_148_n75), .B1(
        u1_srl_148_n66), .B2(u1_srl_148_n76), .ZN(u1_srl_148_n128) );
  OAI221_X1 u1_srl_148_U146 ( .B1(u1_srl_148_n23), .B2(u1_srl_148_n63), .C1(
        u1_srl_148_n25), .C2(u1_srl_148_n64), .A(u1_srl_148_n128), .ZN(
        u1_adj_op_out_sft_12_) );
  AOI22_X1 u1_srl_148_U145 ( .A1(u1_adj_op_17_), .A2(u1_srl_148_n5), .B1(n5304), .B2(u1_srl_148_n4), .ZN(u1_srl_148_n127) );
  AOI22_X1 u1_srl_148_U144 ( .A1(n5305), .A2(u1_srl_148_n6), .B1(u1_adj_op_10_), .B2(u1_srl_148_n100), .ZN(u1_srl_148_n126) );
  AOI22_X1 u1_srl_148_U143 ( .A1(n5300), .A2(u1_srl_148_n99), .B1(
        u1_adj_op_18_), .B2(u1_srl_148_n3), .ZN(u1_srl_148_n125) );
  AOI22_X1 u1_srl_148_U142 ( .A1(u1_srl_148_n70), .A2(u1_srl_148_n69), .B1(
        u1_srl_148_n66), .B2(u1_srl_148_n71), .ZN(u1_srl_148_n124) );
  OAI221_X1 u1_srl_148_U141 ( .B1(u1_srl_148_n30), .B2(u1_srl_148_n63), .C1(
        u1_srl_148_n31), .C2(u1_srl_148_n64), .A(u1_srl_148_n124), .ZN(
        u1_adj_op_out_sft_13_) );
  OAI222_X1 u1_srl_148_U140 ( .A1(u1_srl_148_n28), .A2(u1_srl_148_n63), .B1(
        u1_srl_148_n19), .B2(u1_srl_148_n122), .C1(u1_srl_148_n26), .C2(
        u1_srl_148_n64), .ZN(u1_adj_op_out_sft_14_) );
  AOI222_X1 u1_srl_148_U139 ( .A1(u1_srl_148_n81), .A2(u1_srl_148_n16), .B1(
        u1_srl_148_n80), .B2(u1_srl_148_n66), .C1(u1_srl_148_n79), .C2(
        u1_srl_148_n17), .ZN(u1_srl_148_n121) );
  NOR2_X1 u1_srl_148_U138 ( .A1(u1_exp_diff_sft_4_), .A2(u1_srl_148_n120), 
        .ZN(u1_adj_op_out_sft_16_) );
  AOI222_X1 u1_srl_148_U137 ( .A1(u1_srl_148_n71), .A2(u1_srl_148_n111), .B1(
        u1_srl_148_n69), .B2(u1_srl_148_n119), .C1(u1_srl_148_n67), .C2(
        u1_srl_148_n110), .ZN(u1_srl_148_n112) );
  NOR2_X1 u1_srl_148_U136 ( .A1(u1_exp_diff_sft_4_), .A2(u1_srl_148_n112), 
        .ZN(u1_adj_op_out_sft_17_) );
  AOI222_X1 u1_srl_148_U135 ( .A1(u1_srl_148_n2), .A2(u1_srl_148_n111), .B1(
        u1_srl_148_n109), .B2(u1_srl_148_n119), .C1(u1_srl_148_n86), .C2(
        u1_srl_148_n110), .ZN(u1_srl_148_n103) );
  NOR2_X1 u1_srl_148_U134 ( .A1(u1_exp_diff_sft_4_), .A2(u1_srl_148_n103), 
        .ZN(u1_adj_op_out_sft_18_) );
  NOR2_X1 u1_srl_148_U133 ( .A1(u1_exp_diff_sft_4_), .A2(u1_srl_148_n93), .ZN(
        u1_adj_op_out_sft_19_) );
  AOI22_X1 u1_srl_148_U132 ( .A1(n5296), .A2(u1_srl_148_n5), .B1(n5299), .B2(
        u1_srl_148_n4), .ZN(u1_srl_148_n117) );
  OAI221_X1 u1_srl_148_U131 ( .B1(u1_srl_148_n7), .B2(u1_srl_148_n45), .C1(
        u1_srl_148_n10), .C2(u1_srl_148_n44), .A(u1_srl_148_n117), .ZN(
        u1_srl_148_n116) );
  AOI22_X1 u1_srl_148_U130 ( .A1(n5292), .A2(u1_srl_148_n6), .B1(n5295), .B2(
        u1_srl_148_n100), .ZN(u1_srl_148_n115) );
  OAI22_X1 u1_srl_148_U129 ( .A1(u1_srl_148_n36), .A2(u1_srl_148_n50), .B1(
        u1_srl_148_n10), .B2(u1_srl_148_n61), .ZN(u1_srl_148_n114) );
  AOI222_X1 u1_srl_148_U128 ( .A1(u1_srl_148_n66), .A2(u1_srl_148_n72), .B1(
        u1_srl_148_n17), .B2(u1_srl_148_n114), .C1(u1_srl_148_n70), .C2(
        u1_srl_148_n89), .ZN(u1_srl_148_n113) );
  OAI221_X1 u1_srl_148_U127 ( .B1(u1_srl_148_n32), .B2(u1_srl_148_n63), .C1(
        u1_srl_148_n112), .C2(u1_srl_148_n18), .A(u1_srl_148_n113), .ZN(
        u1_adj_op_out_sft_1_) );
  AOI22_X1 u1_srl_148_U126 ( .A1(u1_srl_148_n76), .A2(u1_srl_148_n110), .B1(
        u1_srl_148_n75), .B2(u1_srl_148_n111), .ZN(u1_srl_148_n90) );
  NOR2_X1 u1_srl_148_U125 ( .A1(u1_exp_diff_sft_4_), .A2(u1_srl_148_n90), .ZN(
        u1_adj_op_out_sft_20_) );
  AOI22_X1 u1_srl_148_U124 ( .A1(u1_srl_148_n71), .A2(u1_srl_148_n110), .B1(
        u1_srl_148_n69), .B2(u1_srl_148_n111), .ZN(u1_srl_148_n87) );
  NOR2_X1 u1_srl_148_U123 ( .A1(u1_exp_diff_sft_4_), .A2(u1_srl_148_n87), .ZN(
        u1_adj_op_out_sft_21_) );
  NOR3_X1 u1_srl_148_U122 ( .A1(u1_srl_148_n19), .A2(u1_exp_diff_sft_4_), .A3(
        n5291), .ZN(u1_adj_op_out_sft_22_) );
  AND2_X1 u1_srl_148_U121 ( .A1(u1_srl_148_n75), .A2(u1_srl_148_n17), .ZN(
        u1_adj_op_out_sft_24_) );
  AND2_X1 u1_srl_148_U120 ( .A1(u1_srl_148_n69), .A2(u1_srl_148_n17), .ZN(
        u1_adj_op_out_sft_25_) );
  AND2_X1 u1_srl_148_U119 ( .A1(u1_srl_148_n17), .A2(u1_srl_148_n109), .ZN(
        u1_adj_op_out_sft_26_) );
  AOI22_X1 u1_srl_148_U118 ( .A1(n5295), .A2(u1_srl_148_n99), .B1(n5298), .B2(
        u1_srl_148_n3), .ZN(u1_srl_148_n108) );
  OAI221_X1 u1_srl_148_U117 ( .B1(u1_srl_148_n7), .B2(u1_srl_148_n44), .C1(
        u1_srl_148_n10), .C2(u1_srl_148_n43), .A(u1_srl_148_n108), .ZN(
        u1_srl_148_n107) );
  OAI222_X1 u1_srl_148_U116 ( .A1(u1_srl_148_n11), .A2(u1_srl_148_n50), .B1(
        u1_srl_148_n7), .B2(u1_srl_148_n61), .C1(u1_srl_148_n36), .C2(
        u1_srl_148_n46), .ZN(u1_srl_148_n106) );
  AOI222_X1 u1_srl_148_U115 ( .A1(u1_srl_148_n66), .A2(u1_srl_148_n105), .B1(
        u1_srl_148_n17), .B2(u1_srl_148_n106), .C1(u1_srl_148_n70), .C2(
        u1_srl_148_n84), .ZN(u1_srl_148_n104) );
  OAI221_X1 u1_srl_148_U114 ( .B1(u1_srl_148_n34), .B2(u1_srl_148_n63), .C1(
        u1_srl_148_n103), .C2(u1_srl_148_n18), .A(u1_srl_148_n104), .ZN(
        u1_adj_op_out_sft_2_) );
  AOI22_X1 u1_srl_148_U113 ( .A1(n5294), .A2(u1_srl_148_n5), .B1(n5297), .B2(
        u1_srl_148_n4), .ZN(u1_srl_148_n102) );
  OAI221_X1 u1_srl_148_U112 ( .B1(u1_srl_148_n7), .B2(u1_srl_148_n43), .C1(
        u1_srl_148_n10), .C2(u1_srl_148_n42), .A(u1_srl_148_n102), .ZN(
        u1_srl_148_n101) );
  AOI22_X1 u1_srl_148_U111 ( .A1(n5298), .A2(u1_srl_148_n6), .B1(n5308), .B2(
        u1_srl_148_n100), .ZN(u1_srl_148_n98) );
  OAI221_X1 u1_srl_148_U110 ( .B1(u1_srl_148_n8), .B2(u1_srl_148_n50), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n46), .A(u1_srl_148_n98), .ZN(
        u1_srl_148_n95) );
  AOI222_X1 u1_srl_148_U109 ( .A1(u1_srl_148_n66), .A2(u1_srl_148_n82), .B1(
        u1_srl_148_n17), .B2(u1_srl_148_n95), .C1(u1_srl_148_n70), .C2(
        u1_srl_148_n79), .ZN(u1_srl_148_n94) );
  OAI221_X1 u1_srl_148_U108 ( .B1(u1_srl_148_n35), .B2(u1_srl_148_n63), .C1(
        u1_srl_148_n93), .C2(u1_srl_148_n18), .A(u1_srl_148_n94), .ZN(
        u1_adj_op_out_sft_3_) );
  AOI222_X1 u1_srl_148_U107 ( .A1(u1_srl_148_n16), .A2(u1_srl_148_n77), .B1(
        u1_srl_148_n70), .B2(u1_srl_148_n74), .C1(u1_srl_148_n66), .C2(
        u1_srl_148_n92), .ZN(u1_srl_148_n91) );
  OAI221_X1 u1_srl_148_U106 ( .B1(u1_srl_148_n21), .B2(u1_srl_148_n64), .C1(
        u1_srl_148_n90), .C2(u1_srl_148_n18), .A(u1_srl_148_n91), .ZN(
        u1_adj_op_out_sft_4_) );
  AOI222_X1 u1_srl_148_U105 ( .A1(u1_srl_148_n16), .A2(u1_srl_148_n72), .B1(
        u1_srl_148_n70), .B2(u1_srl_148_n67), .C1(u1_srl_148_n66), .C2(
        u1_srl_148_n89), .ZN(u1_srl_148_n88) );
  OAI221_X1 u1_srl_148_U104 ( .B1(u1_srl_148_n32), .B2(u1_srl_148_n64), .C1(
        u1_srl_148_n87), .C2(u1_srl_148_n18), .A(u1_srl_148_n88), .ZN(
        u1_adj_op_out_sft_5_) );
  AOI222_X1 u1_srl_148_U103 ( .A1(u1_srl_148_n66), .A2(u1_srl_148_n79), .B1(
        u1_srl_148_n68), .B2(u1_srl_148_n80), .C1(u1_srl_148_n70), .C2(
        u1_srl_148_n81), .ZN(u1_srl_148_n78) );
  OAI221_X1 u1_srl_148_U102 ( .B1(u1_srl_148_n29), .B2(u1_srl_148_n63), .C1(
        u1_srl_148_n35), .C2(u1_srl_148_n64), .A(u1_srl_148_n78), .ZN(
        u1_adj_op_out_sft_7_) );
  AOI222_X1 u1_srl_148_U101 ( .A1(u1_srl_148_n66), .A2(u1_srl_148_n74), .B1(
        u1_srl_148_n68), .B2(u1_srl_148_n75), .C1(u1_srl_148_n70), .C2(
        u1_srl_148_n76), .ZN(u1_srl_148_n73) );
  OAI221_X1 u1_srl_148_U100 ( .B1(u1_srl_148_n25), .B2(u1_srl_148_n63), .C1(
        u1_srl_148_n24), .C2(u1_srl_148_n64), .A(u1_srl_148_n73), .ZN(
        u1_adj_op_out_sft_8_) );
  AOI222_X1 u1_srl_148_U99 ( .A1(u1_srl_148_n66), .A2(u1_srl_148_n67), .B1(
        u1_srl_148_n68), .B2(u1_srl_148_n69), .C1(u1_srl_148_n70), .C2(
        u1_srl_148_n71), .ZN(u1_srl_148_n65) );
  OAI221_X1 u1_srl_148_U98 ( .B1(u1_srl_148_n31), .B2(u1_srl_148_n63), .C1(
        u1_srl_148_n33), .C2(u1_srl_148_n64), .A(u1_srl_148_n65), .ZN(
        u1_adj_op_out_sft_9_) );
  INV_X4 u1_srl_148_U97 ( .A(n2459), .ZN(u1_srl_148_n62) );
  INV_X4 u1_srl_148_U96 ( .A(n5308), .ZN(u1_srl_148_n61) );
  INV_X4 u1_srl_148_U95 ( .A(u1_adj_op_10_), .ZN(u1_srl_148_n60) );
  INV_X4 u1_srl_148_U94 ( .A(n5307), .ZN(u1_srl_148_n59) );
  INV_X4 u1_srl_148_U93 ( .A(n5306), .ZN(u1_srl_148_n58) );
  INV_X4 u1_srl_148_U92 ( .A(n5305), .ZN(u1_srl_148_n57) );
  INV_X4 u1_srl_148_U91 ( .A(n5304), .ZN(u1_srl_148_n56) );
  INV_X4 u1_srl_148_U90 ( .A(n5303), .ZN(u1_srl_148_n55) );
  INV_X4 u1_srl_148_U89 ( .A(n5302), .ZN(u1_srl_148_n54) );
  INV_X4 u1_srl_148_U88 ( .A(u1_adj_op_17_), .ZN(u1_srl_148_n53) );
  INV_X4 u1_srl_148_U87 ( .A(u1_adj_op_18_), .ZN(u1_srl_148_n52) );
  INV_X4 u1_srl_148_U86 ( .A(u1_adj_op_19_), .ZN(u1_srl_148_n51) );
  INV_X4 u1_srl_148_U85 ( .A(n5301), .ZN(u1_srl_148_n50) );
  INV_X4 u1_srl_148_U84 ( .A(u1_adj_op_20_), .ZN(u1_srl_148_n49) );
  INV_X4 u1_srl_148_U83 ( .A(n5300), .ZN(u1_srl_148_n48) );
  INV_X4 u1_srl_148_U82 ( .A(u1_adj_op_22_), .ZN(u1_srl_148_n47) );
  INV_X4 u1_srl_148_U81 ( .A(n5299), .ZN(u1_srl_148_n46) );
  INV_X4 u1_srl_148_U80 ( .A(n5298), .ZN(u1_srl_148_n45) );
  INV_X4 u1_srl_148_U79 ( .A(n5297), .ZN(u1_srl_148_n44) );
  INV_X4 u1_srl_148_U78 ( .A(n5296), .ZN(u1_srl_148_n43) );
  INV_X4 u1_srl_148_U77 ( .A(n5295), .ZN(u1_srl_148_n42) );
  INV_X4 u1_srl_148_U76 ( .A(n5294), .ZN(u1_srl_148_n41) );
  INV_X4 u1_srl_148_U75 ( .A(n5293), .ZN(u1_srl_148_n40) );
  INV_X4 u1_srl_148_U74 ( .A(n5292), .ZN(u1_srl_148_n39) );
  INV_X4 u1_srl_148_U73 ( .A(u1_srl_148_n5), .ZN(u1_srl_148_n36) );
  INV_X4 u1_srl_148_U72 ( .A(u1_srl_148_n101), .ZN(u1_srl_148_n35) );
  INV_X4 u1_srl_148_U71 ( .A(u1_srl_148_n107), .ZN(u1_srl_148_n34) );
  INV_X4 u1_srl_148_U70 ( .A(u1_srl_148_n72), .ZN(u1_srl_148_n33) );
  INV_X4 u1_srl_148_U69 ( .A(u1_srl_148_n116), .ZN(u1_srl_148_n32) );
  INV_X4 u1_srl_148_U68 ( .A(u1_srl_148_n89), .ZN(u1_srl_148_n31) );
  INV_X4 u1_srl_148_U67 ( .A(u1_srl_148_n67), .ZN(u1_srl_148_n30) );
  INV_X4 u1_srl_148_U66 ( .A(u1_srl_148_n82), .ZN(u1_srl_148_n29) );
  INV_X4 u1_srl_148_U65 ( .A(u1_srl_148_n86), .ZN(u1_srl_148_n28) );
  INV_X4 u1_srl_148_U64 ( .A(u1_srl_148_n105), .ZN(u1_srl_148_n27) );
  INV_X4 u1_srl_148_U63 ( .A(u1_srl_148_n84), .ZN(u1_srl_148_n26) );
  INV_X4 u1_srl_148_U62 ( .A(u1_srl_148_n92), .ZN(u1_srl_148_n25) );
  INV_X4 u1_srl_148_U61 ( .A(u1_srl_148_n77), .ZN(u1_srl_148_n24) );
  INV_X4 u1_srl_148_U60 ( .A(u1_srl_148_n74), .ZN(u1_srl_148_n23) );
  INV_X4 u1_srl_148_U59 ( .A(u1_srl_148_n3), .ZN(u1_srl_148_n22) );
  INV_X4 u1_srl_148_U58 ( .A(u1_srl_148_n146), .ZN(u1_srl_148_n21) );
  INV_X4 u1_srl_148_U57 ( .A(n5288), .ZN(u1_srl_148_n20) );
  INV_X4 u1_srl_148_U56 ( .A(u1_srl_148_n123), .ZN(u1_srl_148_n19) );
  INV_X4 u1_srl_148_U55 ( .A(u1_srl_148_n63), .ZN(u1_srl_148_n16) );
  INV_X4 u1_srl_148_U54 ( .A(u1_srl_148_n121), .ZN(u1_adj_op_out_sft_15_) );
  INV_X4 u1_srl_148_U53 ( .A(u1_srl_148_n130), .ZN(u1_srl_148_n14) );
  INV_X4 u1_srl_148_U52 ( .A(u1_srl_148_n129), .ZN(u1_adj_op_out_sft_11_) );
  NOR2_X4 u1_srl_148_U51 ( .A1(u1_srl_148_n38), .A2(u1_srl_148_n37), .ZN(
        u1_srl_148_n99) );
  NOR2_X4 u1_srl_148_U50 ( .A1(u1_srl_148_n38), .A2(u1_srl_148_n37), .ZN(
        u1_srl_148_n6) );
  NOR2_X4 u1_srl_148_U49 ( .A1(u1_srl_148_n38), .A2(u1_srl_148_n37), .ZN(
        u1_srl_148_n5) );
  NOR2_X4 u1_srl_148_U48 ( .A1(n5289), .A2(n5290), .ZN(u1_srl_148_n100) );
  NOR2_X4 u1_srl_148_U47 ( .A1(n5289), .A2(n5290), .ZN(u1_srl_148_n3) );
  NAND2_X4 u1_srl_148_U46 ( .A1(u1_srl_148_n111), .A2(u1_srl_148_n18), .ZN(
        u1_srl_148_n63) );
  NOR2_X4 u1_srl_148_U45 ( .A1(u1_srl_148_n122), .A2(n5288), .ZN(
        u1_srl_148_n66) );
  NOR2_X4 u1_srl_148_U44 ( .A1(u1_srl_148_n20), .A2(u1_srl_148_n122), .ZN(
        u1_srl_148_n70) );
  NAND2_X4 u1_srl_148_U43 ( .A1(u1_srl_148_n110), .A2(u1_srl_148_n18), .ZN(
        u1_srl_148_n64) );
  INV_X8 u1_srl_148_U42 ( .A(u1_exp_diff_sft_4_), .ZN(u1_srl_148_n18) );
  INV_X8 u1_srl_148_U41 ( .A(u1_srl_148_n64), .ZN(u1_srl_148_n17) );
  INV_X8 u1_srl_148_U40 ( .A(u1_srl_148_n96), .ZN(u1_srl_148_n9) );
  MUX2_X2 u1_srl_148_U39 ( .A(u1_srl_148_n109), .B(u1_srl_148_n118), .S(
        u1_srl_148_n20), .Z(u1_srl_148_n123) );
  INV_X8 u1_srl_148_U38 ( .A(u1_srl_148_n97), .ZN(u1_srl_148_n12) );
  OAI221_X2 u1_srl_148_U37 ( .B1(u1_srl_148_n27), .B2(u1_srl_148_n63), .C1(
        u1_srl_148_n34), .C2(u1_srl_148_n64), .A(u1_srl_148_n83), .ZN(
        u1_adj_op_out_sft_6_) );
  AND2_X2 u1_srl_148_U36 ( .A1(u1_srl_148_n80), .A2(u1_srl_148_n17), .ZN(
        u1_adj_op_out_sft_23_) );
  AOI222_X2 u1_srl_148_U35 ( .A1(u1_srl_148_n66), .A2(u1_srl_148_n84), .B1(
        u1_srl_148_n85), .B2(u1_exp_diff_sft_4_), .C1(u1_srl_148_n70), .C2(
        u1_srl_148_n86), .ZN(u1_srl_148_n83) );
  INV_X16 u1_srl_148_U34 ( .A(u1_srl_148_n9), .ZN(u1_srl_148_n8) );
  OAI222_X2 u1_srl_148_U33 ( .A1(u1_srl_148_n62), .A2(u1_srl_148_n10), .B1(
        u1_srl_148_n8), .B2(u1_srl_148_n47), .C1(u1_srl_148_n22), .C2(
        u1_srl_148_n48), .ZN(u1_srl_148_n75) );
  OAI221_X2 u1_srl_148_U32 ( .B1(u1_srl_148_n8), .B2(u1_srl_148_n48), .C1(
        u1_srl_148_n47), .C2(u1_srl_148_n10), .A(u1_srl_148_n134), .ZN(
        u1_srl_148_n80) );
  AOI22_X1 u1_srl_148_U31 ( .A1(u1_srl_148_n81), .A2(u1_srl_148_n110), .B1(
        u1_srl_148_n80), .B2(u1_srl_148_n111), .ZN(u1_srl_148_n93) );
  OAI221_X4 u1_srl_148_U30 ( .B1(u1_srl_148_n7), .B2(u1_srl_148_n55), .C1(
        u1_srl_148_n10), .C2(u1_srl_148_n54), .A(u1_srl_148_n127), .ZN(
        u1_srl_148_n67) );
  INV_X8 u1_srl_148_U29 ( .A(u1_srl_148_n9), .ZN(u1_srl_148_n7) );
  OAI221_X2 u1_srl_148_U28 ( .B1(u1_srl_148_n7), .B2(u1_srl_148_n57), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n56), .A(u1_srl_148_n132), .ZN(
        u1_srl_148_n79) );
  AOI22_X2 u1_srl_148_U27 ( .A1(u1_srl_148_n5), .A2(u1_adj_op_22_), .B1(
        u1_adj_op_19_), .B2(u1_srl_148_n100), .ZN(u1_srl_148_n136) );
  INV_X16 u1_srl_148_U26 ( .A(u1_srl_148_n12), .ZN(u1_srl_148_n11) );
  OAI221_X2 u1_srl_148_U25 ( .B1(u1_srl_148_n7), .B2(u1_srl_148_n59), .C1(
        u1_srl_148_n10), .C2(u1_srl_148_n58), .A(u1_srl_148_n126), .ZN(
        u1_srl_148_n89) );
  AOI22_X2 u1_srl_148_U24 ( .A1(n5302), .A2(u1_srl_148_n6), .B1(n5305), .B2(
        u1_srl_148_n100), .ZN(u1_srl_148_n144) );
  OAI221_X2 u1_srl_148_U23 ( .B1(u1_srl_148_n8), .B2(u1_srl_148_n56), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n55), .A(u1_srl_148_n144), .ZN(
        u1_srl_148_n74) );
  NOR2_X4 u1_srl_148_U22 ( .A1(n5288), .A2(n5291), .ZN(u1_srl_148_n110) );
  AND2_X4 u1_srl_148_U21 ( .A1(u1_exp_diff_sft_4_), .A2(u1_srl_148_n110), .ZN(
        u1_srl_148_n68) );
  OAI221_X2 u1_srl_148_U20 ( .B1(u1_srl_148_n7), .B2(u1_srl_148_n53), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n52), .A(u1_srl_148_n133), .ZN(
        u1_srl_148_n81) );
  OAI221_X2 u1_srl_148_U19 ( .B1(u1_srl_148_n7), .B2(u1_srl_148_n51), .C1(
        u1_srl_148_n10), .C2(u1_srl_148_n49), .A(u1_srl_148_n125), .ZN(
        u1_srl_148_n71) );
  OAI221_X2 u1_srl_148_U18 ( .B1(u1_srl_148_n8), .B2(u1_srl_148_n60), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n59), .A(u1_srl_148_n142), .ZN(
        u1_srl_148_n92) );
  OAI221_X2 u1_srl_148_U17 ( .B1(u1_srl_148_n8), .B2(u1_srl_148_n49), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n48), .A(u1_srl_148_n136), .ZN(
        u1_srl_148_n118) );
  INV_X2 u1_srl_148_U16 ( .A(u1_srl_148_n1), .ZN(u1_srl_148_n2) );
  NOR2_X2 u1_srl_148_U15 ( .A1(n5291), .A2(u1_srl_148_n19), .ZN(u1_srl_148_n85) );
  OAI22_X4 u1_srl_148_U14 ( .A1(u1_srl_148_n22), .A2(u1_srl_148_n47), .B1(
        u1_srl_148_n7), .B2(u1_srl_148_n62), .ZN(u1_srl_148_n69) );
  INV_X8 u1_srl_148_U13 ( .A(u1_srl_148_n12), .ZN(u1_srl_148_n10) );
  NOR2_X4 u1_srl_148_U12 ( .A1(u1_srl_148_n20), .A2(n5291), .ZN(
        u1_srl_148_n111) );
  OAI221_X2 u1_srl_148_U11 ( .B1(u1_srl_148_n7), .B2(u1_srl_148_n39), .C1(
        u1_srl_148_n11), .C2(u1_srl_148_n60), .A(u1_srl_148_n131), .ZN(
        u1_srl_148_n82) );
  NAND2_X2 u1_srl_148_U10 ( .A1(n5289), .A2(u1_srl_148_n38), .ZN(
        u1_srl_148_n96) );
  OAI221_X2 u1_srl_148_U9 ( .B1(u1_srl_148_n7), .B2(u1_srl_148_n41), .C1(
        u1_srl_148_n10), .C2(u1_srl_148_n40), .A(u1_srl_148_n115), .ZN(
        u1_srl_148_n72) );
  INV_X8 u1_srl_148_U8 ( .A(n5289), .ZN(u1_srl_148_n37) );
  NAND2_X2 u1_srl_148_U7 ( .A1(n5290), .A2(u1_srl_148_n37), .ZN(u1_srl_148_n97) );
  INV_X4 u1_srl_148_U6 ( .A(n5290), .ZN(u1_srl_148_n38) );
  NOR2_X2 u1_srl_148_U5 ( .A1(n5289), .A2(n5290), .ZN(u1_srl_148_n4) );
  OAI221_X2 u1_srl_148_U4 ( .B1(u1_srl_148_n8), .B2(u1_srl_148_n52), .C1(
        u1_srl_148_n51), .C2(u1_srl_148_n10), .A(u1_srl_148_n145), .ZN(
        u1_srl_148_n76) );
  INV_X2 u1_srl_148_U3 ( .A(u1_srl_148_n118), .ZN(u1_srl_148_n1) );
  INV_X4 sub_434_3_U115 ( .A(N227), .ZN(sub_434_3_n84) );
  INV_X4 sub_434_3_U114 ( .A(opa_r1[1]), .ZN(sub_434_3_n83) );
  INV_X4 sub_434_3_U113 ( .A(opa_r1[2]), .ZN(sub_434_3_n82) );
  INV_X4 sub_434_3_U112 ( .A(opa_r1[3]), .ZN(sub_434_3_n81) );
  INV_X4 sub_434_3_U111 ( .A(opa_r1[4]), .ZN(sub_434_3_n80) );
  INV_X4 sub_434_3_U110 ( .A(opa_r1[5]), .ZN(sub_434_3_n79) );
  INV_X4 sub_434_3_U109 ( .A(opa_r1[6]), .ZN(sub_434_3_n78) );
  INV_X4 sub_434_3_U108 ( .A(opa_r1[7]), .ZN(sub_434_3_n77) );
  INV_X4 sub_434_3_U107 ( .A(opa_r1[8]), .ZN(sub_434_3_n76) );
  INV_X4 sub_434_3_U106 ( .A(opa_r1[9]), .ZN(sub_434_3_n75) );
  INV_X4 sub_434_3_U105 ( .A(opa_r1[10]), .ZN(sub_434_3_n74) );
  INV_X4 sub_434_3_U104 ( .A(opa_r1[11]), .ZN(sub_434_3_n73) );
  INV_X4 sub_434_3_U103 ( .A(opa_r1[12]), .ZN(sub_434_3_n72) );
  INV_X4 sub_434_3_U102 ( .A(opa_r1[13]), .ZN(sub_434_3_n71) );
  INV_X4 sub_434_3_U101 ( .A(opa_r1[14]), .ZN(sub_434_3_n70) );
  INV_X4 sub_434_3_U100 ( .A(opa_r1[15]), .ZN(sub_434_3_n69) );
  INV_X4 sub_434_3_U99 ( .A(opa_r1[16]), .ZN(sub_434_3_n68) );
  INV_X4 sub_434_3_U98 ( .A(opa_r1[17]), .ZN(sub_434_3_n67) );
  INV_X4 sub_434_3_U97 ( .A(opa_r1[18]), .ZN(sub_434_3_n66) );
  INV_X4 sub_434_3_U96 ( .A(opa_r1[19]), .ZN(sub_434_3_n65) );
  INV_X4 sub_434_3_U95 ( .A(opa_r1[20]), .ZN(sub_434_3_n64) );
  INV_X4 sub_434_3_U94 ( .A(opa_r1[21]), .ZN(sub_434_3_n63) );
  INV_X4 sub_434_3_U93 ( .A(opa_r1[22]), .ZN(sub_434_3_n62) );
  INV_X4 sub_434_3_U92 ( .A(opa_r1[23]), .ZN(sub_434_3_n61) );
  INV_X4 sub_434_3_U91 ( .A(opa_r1[24]), .ZN(sub_434_3_n60) );
  INV_X4 sub_434_3_U90 ( .A(opa_r1[25]), .ZN(sub_434_3_n59) );
  INV_X4 sub_434_3_U89 ( .A(opa_r1[26]), .ZN(sub_434_3_n58) );
  INV_X4 sub_434_3_U88 ( .A(opa_r1[27]), .ZN(sub_434_3_n57) );
  INV_X4 sub_434_3_U87 ( .A(opa_r1[28]), .ZN(sub_434_3_n56) );
  INV_X4 sub_434_3_U86 ( .A(sub_434_3_n55), .ZN(sub_434_3_carry_21_) );
  NAND2_X2 sub_434_3_U85 ( .A1(sub_434_3_n83), .A2(sub_434_3_n84), .ZN(
        sub_434_3_n55) );
  INV_X4 sub_434_3_U84 ( .A(sub_434_3_n54), .ZN(sub_434_3_carry_22_) );
  NAND2_X2 sub_434_3_U83 ( .A1(sub_434_3_n82), .A2(sub_434_3_carry_21_), .ZN(
        sub_434_3_n54) );
  INV_X4 sub_434_3_U82 ( .A(sub_434_3_n53), .ZN(sub_434_3_carry_23_) );
  NAND2_X2 sub_434_3_U81 ( .A1(sub_434_3_n81), .A2(sub_434_3_carry_22_), .ZN(
        sub_434_3_n53) );
  INV_X4 sub_434_3_U80 ( .A(sub_434_3_n52), .ZN(sub_434_3_carry_24_) );
  NAND2_X2 sub_434_3_U79 ( .A1(sub_434_3_n80), .A2(sub_434_3_carry_23_), .ZN(
        sub_434_3_n52) );
  INV_X4 sub_434_3_U78 ( .A(sub_434_3_n51), .ZN(sub_434_3_carry_25_) );
  NAND2_X2 sub_434_3_U77 ( .A1(sub_434_3_n79), .A2(sub_434_3_carry_24_), .ZN(
        sub_434_3_n51) );
  INV_X4 sub_434_3_U76 ( .A(sub_434_3_n50), .ZN(sub_434_3_carry_26_) );
  NAND2_X2 sub_434_3_U75 ( .A1(sub_434_3_n78), .A2(sub_434_3_carry_25_), .ZN(
        sub_434_3_n50) );
  INV_X4 sub_434_3_U74 ( .A(sub_434_3_n49), .ZN(sub_434_3_carry_27_) );
  NAND2_X2 sub_434_3_U73 ( .A1(sub_434_3_n77), .A2(sub_434_3_carry_26_), .ZN(
        sub_434_3_n49) );
  INV_X4 sub_434_3_U72 ( .A(sub_434_3_n48), .ZN(sub_434_3_carry_28_) );
  NAND2_X2 sub_434_3_U71 ( .A1(sub_434_3_n76), .A2(sub_434_3_carry_27_), .ZN(
        sub_434_3_n48) );
  INV_X4 sub_434_3_U70 ( .A(sub_434_3_n47), .ZN(sub_434_3_carry_29_) );
  NAND2_X2 sub_434_3_U69 ( .A1(sub_434_3_n75), .A2(sub_434_3_carry_28_), .ZN(
        sub_434_3_n47) );
  INV_X4 sub_434_3_U68 ( .A(sub_434_3_n46), .ZN(sub_434_3_carry_30_) );
  NAND2_X2 sub_434_3_U67 ( .A1(sub_434_3_n74), .A2(sub_434_3_carry_29_), .ZN(
        sub_434_3_n46) );
  INV_X4 sub_434_3_U66 ( .A(sub_434_3_n45), .ZN(sub_434_3_carry_31_) );
  NAND2_X2 sub_434_3_U65 ( .A1(sub_434_3_n73), .A2(sub_434_3_carry_30_), .ZN(
        sub_434_3_n45) );
  INV_X4 sub_434_3_U64 ( .A(sub_434_3_n44), .ZN(sub_434_3_carry_32_) );
  NAND2_X2 sub_434_3_U63 ( .A1(sub_434_3_n72), .A2(sub_434_3_carry_31_), .ZN(
        sub_434_3_n44) );
  INV_X4 sub_434_3_U62 ( .A(sub_434_3_n43), .ZN(sub_434_3_carry_33_) );
  NAND2_X2 sub_434_3_U61 ( .A1(sub_434_3_n71), .A2(sub_434_3_carry_32_), .ZN(
        sub_434_3_n43) );
  INV_X4 sub_434_3_U60 ( .A(sub_434_3_n42), .ZN(sub_434_3_carry_34_) );
  NAND2_X2 sub_434_3_U59 ( .A1(sub_434_3_n70), .A2(sub_434_3_carry_33_), .ZN(
        sub_434_3_n42) );
  INV_X4 sub_434_3_U58 ( .A(sub_434_3_n41), .ZN(sub_434_3_carry_35_) );
  NAND2_X2 sub_434_3_U57 ( .A1(sub_434_3_n69), .A2(sub_434_3_carry_34_), .ZN(
        sub_434_3_n41) );
  INV_X4 sub_434_3_U56 ( .A(sub_434_3_n40), .ZN(sub_434_3_carry_36_) );
  NAND2_X2 sub_434_3_U55 ( .A1(sub_434_3_n68), .A2(sub_434_3_carry_35_), .ZN(
        sub_434_3_n40) );
  INV_X4 sub_434_3_U54 ( .A(sub_434_3_n39), .ZN(sub_434_3_carry_37_) );
  NAND2_X2 sub_434_3_U53 ( .A1(sub_434_3_n67), .A2(sub_434_3_carry_36_), .ZN(
        sub_434_3_n39) );
  INV_X4 sub_434_3_U52 ( .A(sub_434_3_n38), .ZN(sub_434_3_carry_38_) );
  NAND2_X2 sub_434_3_U51 ( .A1(sub_434_3_n66), .A2(sub_434_3_carry_37_), .ZN(
        sub_434_3_n38) );
  INV_X4 sub_434_3_U50 ( .A(sub_434_3_n37), .ZN(sub_434_3_carry_39_) );
  NAND2_X2 sub_434_3_U49 ( .A1(sub_434_3_n65), .A2(sub_434_3_carry_38_), .ZN(
        sub_434_3_n37) );
  INV_X4 sub_434_3_U48 ( .A(sub_434_3_n36), .ZN(sub_434_3_carry_40_) );
  NAND2_X2 sub_434_3_U47 ( .A1(sub_434_3_n64), .A2(sub_434_3_carry_39_), .ZN(
        sub_434_3_n36) );
  INV_X4 sub_434_3_U46 ( .A(sub_434_3_n35), .ZN(sub_434_3_carry_41_) );
  NAND2_X2 sub_434_3_U45 ( .A1(sub_434_3_n63), .A2(sub_434_3_carry_40_), .ZN(
        sub_434_3_n35) );
  INV_X4 sub_434_3_U44 ( .A(sub_434_3_n34), .ZN(sub_434_3_carry_42_) );
  NAND2_X2 sub_434_3_U43 ( .A1(sub_434_3_n62), .A2(sub_434_3_carry_41_), .ZN(
        sub_434_3_n34) );
  INV_X4 sub_434_3_U42 ( .A(sub_434_3_n33), .ZN(sub_434_3_carry_43_) );
  NAND2_X2 sub_434_3_U41 ( .A1(sub_434_3_n61), .A2(sub_434_3_carry_42_), .ZN(
        sub_434_3_n33) );
  INV_X4 sub_434_3_U40 ( .A(sub_434_3_n32), .ZN(sub_434_3_carry_44_) );
  NAND2_X2 sub_434_3_U39 ( .A1(sub_434_3_n60), .A2(sub_434_3_carry_43_), .ZN(
        sub_434_3_n32) );
  INV_X4 sub_434_3_U38 ( .A(sub_434_3_n31), .ZN(N322) );
  XNOR2_X2 sub_434_3_U37 ( .A(sub_434_3_n59), .B(sub_434_3_carry_44_), .ZN(
        sub_434_3_n31) );
  INV_X4 sub_434_3_U36 ( .A(sub_434_3_n30), .ZN(sub_434_3_carry_45_) );
  NAND2_X2 sub_434_3_U35 ( .A1(sub_434_3_n59), .A2(sub_434_3_carry_44_), .ZN(
        sub_434_3_n30) );
  INV_X4 sub_434_3_U34 ( .A(sub_434_3_n29), .ZN(N323) );
  XNOR2_X2 sub_434_3_U33 ( .A(sub_434_3_n58), .B(sub_434_3_carry_45_), .ZN(
        sub_434_3_n29) );
  INV_X4 sub_434_3_U32 ( .A(sub_434_3_n28), .ZN(sub_434_3_carry_46_) );
  NAND2_X2 sub_434_3_U31 ( .A1(sub_434_3_n58), .A2(sub_434_3_carry_45_), .ZN(
        sub_434_3_n28) );
  INV_X4 sub_434_3_U30 ( .A(sub_434_3_n27), .ZN(N324) );
  XNOR2_X2 sub_434_3_U29 ( .A(sub_434_3_n57), .B(sub_434_3_carry_46_), .ZN(
        sub_434_3_n27) );
  INV_X4 sub_434_3_U28 ( .A(sub_434_3_n26), .ZN(sub_434_3_carry_47_) );
  NAND2_X2 sub_434_3_U27 ( .A1(sub_434_3_n57), .A2(sub_434_3_carry_46_), .ZN(
        sub_434_3_n26) );
  INV_X4 sub_434_3_U26 ( .A(sub_434_3_n25), .ZN(N325) );
  XNOR2_X2 sub_434_3_U25 ( .A(sub_434_3_n56), .B(sub_434_3_carry_47_), .ZN(
        sub_434_3_n25) );
  XOR2_X1 sub_434_3_U24 ( .A(sub_434_3_n60), .B(sub_434_3_carry_43_), .Z(N321)
         );
  XOR2_X1 sub_434_3_U23 ( .A(sub_434_3_n61), .B(sub_434_3_carry_42_), .Z(N320)
         );
  XOR2_X1 sub_434_3_U22 ( .A(sub_434_3_n62), .B(sub_434_3_carry_41_), .Z(N319)
         );
  XOR2_X1 sub_434_3_U21 ( .A(sub_434_3_n63), .B(sub_434_3_carry_40_), .Z(N318)
         );
  XOR2_X1 sub_434_3_U20 ( .A(sub_434_3_n64), .B(sub_434_3_carry_39_), .Z(N317)
         );
  XOR2_X1 sub_434_3_U19 ( .A(sub_434_3_n65), .B(sub_434_3_carry_38_), .Z(N316)
         );
  XOR2_X1 sub_434_3_U18 ( .A(sub_434_3_n66), .B(sub_434_3_carry_37_), .Z(N315)
         );
  XOR2_X1 sub_434_3_U17 ( .A(sub_434_3_n67), .B(sub_434_3_carry_36_), .Z(N314)
         );
  XOR2_X1 sub_434_3_U16 ( .A(sub_434_3_n68), .B(sub_434_3_carry_35_), .Z(N313)
         );
  XOR2_X1 sub_434_3_U15 ( .A(sub_434_3_n69), .B(sub_434_3_carry_34_), .Z(N312)
         );
  XOR2_X1 sub_434_3_U14 ( .A(sub_434_3_n70), .B(sub_434_3_carry_33_), .Z(N311)
         );
  XOR2_X1 sub_434_3_U13 ( .A(sub_434_3_n71), .B(sub_434_3_carry_32_), .Z(N310)
         );
  XOR2_X1 sub_434_3_U12 ( .A(sub_434_3_n72), .B(sub_434_3_carry_31_), .Z(N309)
         );
  XOR2_X1 sub_434_3_U11 ( .A(sub_434_3_n73), .B(sub_434_3_carry_30_), .Z(N308)
         );
  XOR2_X1 sub_434_3_U10 ( .A(sub_434_3_n74), .B(sub_434_3_carry_29_), .Z(N307)
         );
  XOR2_X1 sub_434_3_U9 ( .A(sub_434_3_n75), .B(sub_434_3_carry_28_), .Z(N306)
         );
  XOR2_X1 sub_434_3_U8 ( .A(sub_434_3_n76), .B(sub_434_3_carry_27_), .Z(N305)
         );
  XOR2_X1 sub_434_3_U7 ( .A(sub_434_3_n77), .B(sub_434_3_carry_26_), .Z(N304)
         );
  XOR2_X1 sub_434_3_U6 ( .A(sub_434_3_n78), .B(sub_434_3_carry_25_), .Z(N303)
         );
  XOR2_X1 sub_434_3_U5 ( .A(sub_434_3_n79), .B(sub_434_3_carry_24_), .Z(N302)
         );
  XOR2_X1 sub_434_3_U4 ( .A(sub_434_3_n80), .B(sub_434_3_carry_23_), .Z(N301)
         );
  XOR2_X1 sub_434_3_U3 ( .A(sub_434_3_n81), .B(sub_434_3_carry_22_), .Z(N300)
         );
  XOR2_X1 sub_434_3_U2 ( .A(sub_434_3_n82), .B(sub_434_3_carry_21_), .Z(N299)
         );
  XOR2_X1 sub_434_3_U1 ( .A(sub_434_3_n83), .B(sub_434_3_n84), .Z(N298) );
  INV_X4 sub_434_b0_U80 ( .A(N227), .ZN(sub_434_b0_n70) );
  INV_X4 sub_434_b0_U79 ( .A(opa_r1[1]), .ZN(sub_434_b0_n69) );
  INV_X4 sub_434_b0_U78 ( .A(opa_r1[2]), .ZN(sub_434_b0_n68) );
  INV_X4 sub_434_b0_U77 ( .A(opa_r1[3]), .ZN(sub_434_b0_n67) );
  INV_X4 sub_434_b0_U76 ( .A(opa_r1[4]), .ZN(sub_434_b0_n66) );
  INV_X4 sub_434_b0_U75 ( .A(opa_r1[5]), .ZN(sub_434_b0_n65) );
  INV_X4 sub_434_b0_U74 ( .A(opa_r1[6]), .ZN(sub_434_b0_n64) );
  INV_X4 sub_434_b0_U73 ( .A(opa_r1[7]), .ZN(sub_434_b0_n63) );
  INV_X4 sub_434_b0_U72 ( .A(opa_r1[8]), .ZN(sub_434_b0_n62) );
  INV_X4 sub_434_b0_U71 ( .A(opa_r1[9]), .ZN(sub_434_b0_n61) );
  INV_X4 sub_434_b0_U70 ( .A(opa_r1[10]), .ZN(sub_434_b0_n60) );
  INV_X4 sub_434_b0_U69 ( .A(opa_r1[11]), .ZN(sub_434_b0_n59) );
  INV_X4 sub_434_b0_U68 ( .A(opa_r1[12]), .ZN(sub_434_b0_n58) );
  INV_X4 sub_434_b0_U67 ( .A(opa_r1[13]), .ZN(sub_434_b0_n57) );
  INV_X4 sub_434_b0_U66 ( .A(opa_r1[14]), .ZN(sub_434_b0_n56) );
  INV_X4 sub_434_b0_U65 ( .A(opa_r1[15]), .ZN(sub_434_b0_n55) );
  INV_X4 sub_434_b0_U64 ( .A(opa_r1[16]), .ZN(sub_434_b0_n54) );
  INV_X4 sub_434_b0_U63 ( .A(opa_r1[17]), .ZN(sub_434_b0_n53) );
  INV_X4 sub_434_b0_U62 ( .A(opa_r1[18]), .ZN(sub_434_b0_n52) );
  INV_X4 sub_434_b0_U61 ( .A(opa_r1[19]), .ZN(sub_434_b0_n51) );
  INV_X4 sub_434_b0_U60 ( .A(opa_r1[20]), .ZN(sub_434_b0_n50) );
  INV_X4 sub_434_b0_U59 ( .A(opa_r1[21]), .ZN(sub_434_b0_n49) );
  INV_X4 sub_434_b0_U58 ( .A(opa_r1[22]), .ZN(sub_434_b0_n48) );
  INV_X4 sub_434_b0_U57 ( .A(N224), .ZN(sub_434_b0_n47) );
  INV_X4 sub_434_b0_U56 ( .A(sub_434_b0_n46), .ZN(sub_434_b0_carry_3_) );
  NAND2_X2 sub_434_b0_U55 ( .A1(sub_434_b0_n68), .A2(sub_434_b0_n3), .ZN(
        sub_434_b0_n46) );
  INV_X4 sub_434_b0_U54 ( .A(sub_434_b0_n45), .ZN(sub_434_b0_carry_5_) );
  NAND2_X2 sub_434_b0_U53 ( .A1(sub_434_b0_n66), .A2(sub_434_b0_n2), .ZN(
        sub_434_b0_n45) );
  INV_X4 sub_434_b0_U52 ( .A(sub_434_b0_n44), .ZN(sub_434_b0_carry_8_) );
  NAND2_X2 sub_434_b0_U51 ( .A1(sub_434_b0_n63), .A2(sub_434_b0_n12), .ZN(
        sub_434_b0_n44) );
  INV_X4 sub_434_b0_U50 ( .A(sub_434_b0_n43), .ZN(sub_434_b0_carry_10_) );
  NAND2_X2 sub_434_b0_U49 ( .A1(sub_434_b0_n61), .A2(sub_434_b0_n11), .ZN(
        sub_434_b0_n43) );
  INV_X4 sub_434_b0_U48 ( .A(sub_434_b0_n42), .ZN(sub_434_b0_carry_12_) );
  NAND2_X2 sub_434_b0_U47 ( .A1(sub_434_b0_n59), .A2(sub_434_b0_n10), .ZN(
        sub_434_b0_n42) );
  INV_X4 sub_434_b0_U46 ( .A(sub_434_b0_n41), .ZN(sub_434_b0_carry_14_) );
  NAND2_X2 sub_434_b0_U45 ( .A1(sub_434_b0_n57), .A2(sub_434_b0_n9), .ZN(
        sub_434_b0_n41) );
  INV_X4 sub_434_b0_U44 ( .A(sub_434_b0_n40), .ZN(sub_434_b0_carry_16_) );
  NAND2_X2 sub_434_b0_U43 ( .A1(sub_434_b0_n55), .A2(sub_434_b0_n8), .ZN(
        sub_434_b0_n40) );
  INV_X4 sub_434_b0_U42 ( .A(sub_434_b0_n39), .ZN(sub_434_b0_carry_18_) );
  NAND2_X2 sub_434_b0_U41 ( .A1(sub_434_b0_n53), .A2(sub_434_b0_n7), .ZN(
        sub_434_b0_n39) );
  INV_X4 sub_434_b0_U40 ( .A(sub_434_b0_n38), .ZN(sub_434_b0_carry_20_) );
  NAND2_X2 sub_434_b0_U39 ( .A1(sub_434_b0_n51), .A2(sub_434_b0_n6), .ZN(
        sub_434_b0_n38) );
  INV_X4 sub_434_b0_U38 ( .A(sub_434_b0_n37), .ZN(sub_434_b0_carry_22_) );
  NAND2_X2 sub_434_b0_U37 ( .A1(sub_434_b0_n49), .A2(sub_434_b0_n5), .ZN(
        sub_434_b0_n37) );
  NAND2_X2 sub_434_b0_U36 ( .A1(sub_434_b0_n47), .A2(sub_434_b0_n4), .ZN(N251)
         );
  XOR2_X2 sub_434_b0_U35 ( .A(sub_434_b0_n69), .B(sub_434_b0_n70), .Z(N228) );
  XOR2_X2 sub_434_b0_U34 ( .A(sub_434_b0_n47), .B(sub_434_b0_n4), .Z(N250) );
  XOR2_X2 sub_434_b0_U33 ( .A(sub_434_b0_n48), .B(sub_434_b0_carry_22_), .Z(
        N249) );
  XOR2_X2 sub_434_b0_U32 ( .A(sub_434_b0_n49), .B(sub_434_b0_n5), .Z(N248) );
  XOR2_X2 sub_434_b0_U31 ( .A(sub_434_b0_n50), .B(sub_434_b0_carry_20_), .Z(
        N247) );
  XOR2_X2 sub_434_b0_U30 ( .A(sub_434_b0_n51), .B(sub_434_b0_n6), .Z(N246) );
  XOR2_X2 sub_434_b0_U29 ( .A(sub_434_b0_n52), .B(sub_434_b0_carry_18_), .Z(
        N245) );
  XOR2_X2 sub_434_b0_U28 ( .A(sub_434_b0_n53), .B(sub_434_b0_n7), .Z(N244) );
  XOR2_X2 sub_434_b0_U27 ( .A(sub_434_b0_n54), .B(sub_434_b0_carry_16_), .Z(
        N243) );
  XOR2_X2 sub_434_b0_U26 ( .A(sub_434_b0_n55), .B(sub_434_b0_n8), .Z(N242) );
  XOR2_X2 sub_434_b0_U25 ( .A(sub_434_b0_n56), .B(sub_434_b0_carry_14_), .Z(
        N241) );
  XOR2_X2 sub_434_b0_U24 ( .A(sub_434_b0_n57), .B(sub_434_b0_n9), .Z(N240) );
  XOR2_X2 sub_434_b0_U23 ( .A(sub_434_b0_n58), .B(sub_434_b0_carry_12_), .Z(
        N239) );
  XOR2_X2 sub_434_b0_U22 ( .A(sub_434_b0_n59), .B(sub_434_b0_n10), .Z(N238) );
  XOR2_X2 sub_434_b0_U21 ( .A(sub_434_b0_n60), .B(sub_434_b0_carry_10_), .Z(
        N237) );
  XOR2_X2 sub_434_b0_U20 ( .A(sub_434_b0_n61), .B(sub_434_b0_n11), .Z(N236) );
  XOR2_X2 sub_434_b0_U19 ( .A(sub_434_b0_n62), .B(sub_434_b0_carry_8_), .Z(
        N235) );
  XOR2_X2 sub_434_b0_U18 ( .A(sub_434_b0_n63), .B(sub_434_b0_n12), .Z(N234) );
  XOR2_X2 sub_434_b0_U17 ( .A(sub_434_b0_n64), .B(sub_434_b0_n1), .Z(N233) );
  XOR2_X2 sub_434_b0_U16 ( .A(sub_434_b0_n65), .B(sub_434_b0_carry_5_), .Z(
        N232) );
  XOR2_X2 sub_434_b0_U15 ( .A(sub_434_b0_n66), .B(sub_434_b0_n2), .Z(N231) );
  XOR2_X2 sub_434_b0_U14 ( .A(sub_434_b0_n67), .B(sub_434_b0_carry_3_), .Z(
        N230) );
  XOR2_X2 sub_434_b0_U13 ( .A(sub_434_b0_n68), .B(sub_434_b0_n3), .Z(N229) );
  AND2_X4 sub_434_b0_U12 ( .A1(sub_434_b0_n64), .A2(sub_434_b0_n1), .ZN(
        sub_434_b0_n12) );
  AND2_X4 sub_434_b0_U11 ( .A1(sub_434_b0_n62), .A2(sub_434_b0_carry_8_), .ZN(
        sub_434_b0_n11) );
  AND2_X4 sub_434_b0_U10 ( .A1(sub_434_b0_n60), .A2(sub_434_b0_carry_10_), 
        .ZN(sub_434_b0_n10) );
  AND2_X4 sub_434_b0_U9 ( .A1(sub_434_b0_n58), .A2(sub_434_b0_carry_12_), .ZN(
        sub_434_b0_n9) );
  AND2_X4 sub_434_b0_U8 ( .A1(sub_434_b0_n56), .A2(sub_434_b0_carry_14_), .ZN(
        sub_434_b0_n8) );
  AND2_X4 sub_434_b0_U7 ( .A1(sub_434_b0_n54), .A2(sub_434_b0_carry_16_), .ZN(
        sub_434_b0_n7) );
  AND2_X4 sub_434_b0_U6 ( .A1(sub_434_b0_n52), .A2(sub_434_b0_carry_18_), .ZN(
        sub_434_b0_n6) );
  AND2_X4 sub_434_b0_U5 ( .A1(sub_434_b0_n50), .A2(sub_434_b0_carry_20_), .ZN(
        sub_434_b0_n5) );
  AND2_X4 sub_434_b0_U4 ( .A1(sub_434_b0_n48), .A2(sub_434_b0_carry_22_), .ZN(
        sub_434_b0_n4) );
  AND2_X4 sub_434_b0_U3 ( .A1(sub_434_b0_n69), .A2(sub_434_b0_n70), .ZN(
        sub_434_b0_n3) );
  AND2_X4 sub_434_b0_U2 ( .A1(sub_434_b0_n67), .A2(sub_434_b0_carry_3_), .ZN(
        sub_434_b0_n2) );
  AND2_X4 sub_434_b0_U1 ( .A1(sub_434_b0_n65), .A2(sub_434_b0_carry_5_), .ZN(
        sub_434_b0_n1) );
  AND2_X1 sll_384_U49 ( .A1(fracta_mul[0]), .A2(sll_384_n4), .ZN(
        sll_384_ML_int_1__0_) );
  AND2_X1 sll_384_U48 ( .A1(sll_384_ML_int_1__0_), .A2(sll_384_n7), .ZN(
        sll_384_ML_int_2__0_) );
  AND2_X1 sll_384_U47 ( .A1(sll_384_ML_int_1__1_), .A2(sll_384_n7), .ZN(
        sll_384_ML_int_2__1_) );
  AND2_X1 sll_384_U46 ( .A1(sll_384_ML_int_2__0_), .A2(sll_384_n1), .ZN(
        sll_384_ML_int_3__0_) );
  AND2_X1 sll_384_U45 ( .A1(sll_384_ML_int_2__1_), .A2(sll_384_n1), .ZN(
        sll_384_ML_int_3__1_) );
  AND2_X1 sll_384_U44 ( .A1(sll_384_ML_int_2__2_), .A2(sll_384_n1), .ZN(
        sll_384_ML_int_3__2_) );
  AND2_X1 sll_384_U43 ( .A1(sll_384_ML_int_2__3_), .A2(sll_384_n1), .ZN(
        sll_384_ML_int_3__3_) );
  NAND2_X1 sll_384_U42 ( .A1(sll_384_ML_int_3__0_), .A2(sll_384_n2), .ZN(
        sll_384_n24) );
  NAND2_X1 sll_384_U41 ( .A1(sll_384_ML_int_3__1_), .A2(sll_384_n2), .ZN(
        sll_384_n23) );
  NAND2_X1 sll_384_U40 ( .A1(sll_384_ML_int_3__2_), .A2(sll_384_n2), .ZN(
        sll_384_n22) );
  NAND2_X1 sll_384_U39 ( .A1(sll_384_ML_int_3__3_), .A2(sll_384_n2), .ZN(
        sll_384_n21) );
  NAND2_X1 sll_384_U38 ( .A1(sll_384_ML_int_3__4_), .A2(sll_384_n2), .ZN(
        sll_384_n20) );
  NAND2_X1 sll_384_U37 ( .A1(sll_384_ML_int_3__5_), .A2(sll_384_n2), .ZN(
        sll_384_n19) );
  NAND2_X1 sll_384_U36 ( .A1(sll_384_ML_int_3__6_), .A2(sll_384_n2), .ZN(
        sll_384_n18) );
  NAND2_X1 sll_384_U35 ( .A1(sll_384_ML_int_3__7_), .A2(sll_384_n2), .ZN(
        sll_384_n17) );
  NOR2_X1 sll_384_U34 ( .A1(n2587), .A2(sll_384_n24), .ZN(N172) );
  AND2_X1 sll_384_U33 ( .A1(sll_384_ML_int_4__10_), .A2(sll_384_n16), .ZN(N182) );
  AND2_X1 sll_384_U32 ( .A1(sll_384_ML_int_4__11_), .A2(sll_384_n16), .ZN(N183) );
  AND2_X1 sll_384_U31 ( .A1(sll_384_ML_int_4__12_), .A2(sll_384_n16), .ZN(N184) );
  AND2_X1 sll_384_U30 ( .A1(sll_384_ML_int_4__13_), .A2(sll_384_n16), .ZN(N185) );
  AND2_X1 sll_384_U29 ( .A1(sll_384_ML_int_4__14_), .A2(sll_384_n16), .ZN(N186) );
  AND2_X1 sll_384_U28 ( .A1(sll_384_ML_int_4__15_), .A2(sll_384_n16), .ZN(N187) );
  NOR2_X1 sll_384_U27 ( .A1(n2587), .A2(sll_384_n23), .ZN(N173) );
  NOR2_X1 sll_384_U26 ( .A1(n2587), .A2(sll_384_n22), .ZN(N174) );
  NOR2_X1 sll_384_U25 ( .A1(n2587), .A2(sll_384_n21), .ZN(N175) );
  NOR2_X1 sll_384_U24 ( .A1(n2587), .A2(sll_384_n20), .ZN(N176) );
  NOR2_X1 sll_384_U23 ( .A1(n2587), .A2(sll_384_n19), .ZN(N177) );
  NOR2_X1 sll_384_U22 ( .A1(n2587), .A2(sll_384_n18), .ZN(N178) );
  NOR2_X1 sll_384_U21 ( .A1(n2587), .A2(sll_384_n17), .ZN(N179) );
  AND2_X1 sll_384_U20 ( .A1(sll_384_ML_int_4__8_), .A2(sll_384_n16), .ZN(N180)
         );
  AND2_X1 sll_384_U19 ( .A1(sll_384_ML_int_4__9_), .A2(sll_384_n16), .ZN(N181)
         );
  INV_X4 sll_384_U18 ( .A(n2587), .ZN(sll_384_n16) );
  INV_X4 sll_384_U17 ( .A(sll_384_n17), .ZN(sll_384_n15) );
  INV_X4 sll_384_U16 ( .A(sll_384_n21), .ZN(sll_384_n14) );
  INV_X4 sll_384_U15 ( .A(sll_384_n19), .ZN(sll_384_n13) );
  INV_X4 sll_384_U14 ( .A(sll_384_n23), .ZN(sll_384_n12) );
  INV_X4 sll_384_U13 ( .A(sll_384_n18), .ZN(sll_384_n11) );
  INV_X4 sll_384_U12 ( .A(sll_384_n22), .ZN(sll_384_n10) );
  INV_X4 sll_384_U11 ( .A(sll_384_n20), .ZN(sll_384_n9) );
  INV_X4 sll_384_U10 ( .A(sll_384_n24), .ZN(sll_384_n8) );
  INV_X4 sll_384_U9 ( .A(sll_384_n2), .ZN(sll_384_n3) );
  INV_X4 sll_384_U8 ( .A(n2597), .ZN(sll_384_n2) );
  INV_X4 sll_384_U7 ( .A(N107), .ZN(sll_384_n1) );
  INV_X4 sll_384_U6 ( .A(sll_384_n7), .ZN(sll_384_n6) );
  INV_X4 sll_384_U5 ( .A(N141), .ZN(sll_384_n7) );
  INV_X4 sll_384_U4 ( .A(sll_384_n4), .ZN(sll_384_n5) );
  INV_X4 sll_384_U3 ( .A(N170), .ZN(sll_384_n4) );
  MUX2_X2 sll_384_M1_0_1 ( .A(n2586), .B(fracta_mul[0]), .S(sll_384_n5), .Z(
        sll_384_ML_int_1__1_) );
  MUX2_X2 sll_384_M1_0_2 ( .A(fracta_mul[2]), .B(n2586), .S(sll_384_n5), .Z(
        sll_384_ML_int_1__2_) );
  MUX2_X2 sll_384_M1_0_3 ( .A(fracta_mul[3]), .B(fracta_mul[2]), .S(sll_384_n5), .Z(sll_384_ML_int_1__3_) );
  MUX2_X2 sll_384_M1_0_4 ( .A(fracta_mul[4]), .B(fracta_mul[3]), .S(sll_384_n5), .Z(sll_384_ML_int_1__4_) );
  MUX2_X2 sll_384_M1_0_5 ( .A(fracta_mul[5]), .B(fracta_mul[4]), .S(sll_384_n5), .Z(sll_384_ML_int_1__5_) );
  MUX2_X2 sll_384_M1_0_6 ( .A(fracta_mul[6]), .B(fracta_mul[5]), .S(sll_384_n5), .Z(sll_384_ML_int_1__6_) );
  MUX2_X2 sll_384_M1_0_7 ( .A(fracta_mul[7]), .B(fracta_mul[6]), .S(sll_384_n5), .Z(sll_384_ML_int_1__7_) );
  MUX2_X2 sll_384_M1_0_8 ( .A(fracta_mul[8]), .B(fracta_mul[7]), .S(sll_384_n5), .Z(sll_384_ML_int_1__8_) );
  MUX2_X2 sll_384_M1_0_9 ( .A(fracta_mul[9]), .B(fracta_mul[8]), .S(sll_384_n5), .Z(sll_384_ML_int_1__9_) );
  MUX2_X2 sll_384_M1_0_10 ( .A(fracta_mul[10]), .B(fracta_mul[9]), .S(
        sll_384_n5), .Z(sll_384_ML_int_1__10_) );
  MUX2_X2 sll_384_M1_0_11 ( .A(fracta_mul[11]), .B(fracta_mul[10]), .S(
        sll_384_n5), .Z(sll_384_ML_int_1__11_) );
  MUX2_X2 sll_384_M1_0_12 ( .A(fracta_mul[12]), .B(fracta_mul[11]), .S(
        sll_384_n5), .Z(sll_384_ML_int_1__12_) );
  MUX2_X2 sll_384_M1_0_13 ( .A(fracta_mul[13]), .B(fracta_mul[12]), .S(
        sll_384_n5), .Z(sll_384_ML_int_1__13_) );
  MUX2_X2 sll_384_M1_0_14 ( .A(fracta_mul[14]), .B(fracta_mul[13]), .S(N170), 
        .Z(sll_384_ML_int_1__14_) );
  MUX2_X2 sll_384_M1_0_15 ( .A(fracta_mul[15]), .B(fracta_mul[14]), .S(N170), 
        .Z(sll_384_ML_int_1__15_) );
  MUX2_X2 sll_384_M1_0_16 ( .A(fracta_mul[16]), .B(fracta_mul[15]), .S(
        sll_384_n5), .Z(sll_384_ML_int_1__16_) );
  MUX2_X2 sll_384_M1_0_17 ( .A(fracta_mul[17]), .B(fracta_mul[16]), .S(N170), 
        .Z(sll_384_ML_int_1__17_) );
  MUX2_X2 sll_384_M1_0_18 ( .A(fracta_mul[18]), .B(fracta_mul[17]), .S(N170), 
        .Z(sll_384_ML_int_1__18_) );
  MUX2_X2 sll_384_M1_0_19 ( .A(fracta_mul[19]), .B(fracta_mul[18]), .S(N170), 
        .Z(sll_384_ML_int_1__19_) );
  MUX2_X2 sll_384_M1_0_20 ( .A(fracta_mul[20]), .B(fracta_mul[19]), .S(N170), 
        .Z(sll_384_ML_int_1__20_) );
  MUX2_X2 sll_384_M1_0_21 ( .A(fracta_mul[21]), .B(fracta_mul[20]), .S(N170), 
        .Z(sll_384_ML_int_1__21_) );
  MUX2_X2 sll_384_M1_0_22 ( .A(fracta_mul[22]), .B(fracta_mul[21]), .S(N170), 
        .Z(sll_384_ML_int_1__22_) );
  MUX2_X2 sll_384_M1_0_23 ( .A(u2_N124), .B(fracta_mul[22]), .S(N170), .Z(
        sll_384_ML_int_1__23_) );
  MUX2_X2 sll_384_M1_1_2 ( .A(sll_384_ML_int_1__2_), .B(sll_384_ML_int_1__0_), 
        .S(sll_384_n6), .Z(sll_384_ML_int_2__2_) );
  MUX2_X2 sll_384_M1_1_3 ( .A(sll_384_ML_int_1__3_), .B(sll_384_ML_int_1__1_), 
        .S(sll_384_n6), .Z(sll_384_ML_int_2__3_) );
  MUX2_X2 sll_384_M1_1_4 ( .A(sll_384_ML_int_1__4_), .B(sll_384_ML_int_1__2_), 
        .S(sll_384_n6), .Z(sll_384_ML_int_2__4_) );
  MUX2_X2 sll_384_M1_1_5 ( .A(sll_384_ML_int_1__5_), .B(sll_384_ML_int_1__3_), 
        .S(sll_384_n6), .Z(sll_384_ML_int_2__5_) );
  MUX2_X2 sll_384_M1_1_6 ( .A(sll_384_ML_int_1__6_), .B(sll_384_ML_int_1__4_), 
        .S(sll_384_n6), .Z(sll_384_ML_int_2__6_) );
  MUX2_X2 sll_384_M1_1_7 ( .A(sll_384_ML_int_1__7_), .B(sll_384_ML_int_1__5_), 
        .S(sll_384_n6), .Z(sll_384_ML_int_2__7_) );
  MUX2_X2 sll_384_M1_1_8 ( .A(sll_384_ML_int_1__8_), .B(sll_384_ML_int_1__6_), 
        .S(sll_384_n6), .Z(sll_384_ML_int_2__8_) );
  MUX2_X2 sll_384_M1_1_9 ( .A(sll_384_ML_int_1__9_), .B(sll_384_ML_int_1__7_), 
        .S(sll_384_n6), .Z(sll_384_ML_int_2__9_) );
  MUX2_X2 sll_384_M1_1_10 ( .A(sll_384_ML_int_1__10_), .B(sll_384_ML_int_1__8_), .S(sll_384_n6), .Z(sll_384_ML_int_2__10_) );
  MUX2_X2 sll_384_M1_1_11 ( .A(sll_384_ML_int_1__11_), .B(sll_384_ML_int_1__9_), .S(sll_384_n6), .Z(sll_384_ML_int_2__11_) );
  MUX2_X2 sll_384_M1_1_12 ( .A(sll_384_ML_int_1__12_), .B(
        sll_384_ML_int_1__10_), .S(sll_384_n6), .Z(sll_384_ML_int_2__12_) );
  MUX2_X2 sll_384_M1_1_13 ( .A(sll_384_ML_int_1__13_), .B(
        sll_384_ML_int_1__11_), .S(sll_384_n6), .Z(sll_384_ML_int_2__13_) );
  MUX2_X2 sll_384_M1_1_14 ( .A(sll_384_ML_int_1__14_), .B(
        sll_384_ML_int_1__12_), .S(sll_384_n6), .Z(sll_384_ML_int_2__14_) );
  MUX2_X2 sll_384_M1_1_15 ( .A(sll_384_ML_int_1__15_), .B(
        sll_384_ML_int_1__13_), .S(sll_384_n6), .Z(sll_384_ML_int_2__15_) );
  MUX2_X2 sll_384_M1_1_16 ( .A(sll_384_ML_int_1__16_), .B(
        sll_384_ML_int_1__14_), .S(sll_384_n6), .Z(sll_384_ML_int_2__16_) );
  MUX2_X2 sll_384_M1_1_17 ( .A(sll_384_ML_int_1__17_), .B(
        sll_384_ML_int_1__15_), .S(sll_384_n6), .Z(sll_384_ML_int_2__17_) );
  MUX2_X2 sll_384_M1_1_18 ( .A(sll_384_ML_int_1__18_), .B(
        sll_384_ML_int_1__16_), .S(sll_384_n6), .Z(sll_384_ML_int_2__18_) );
  MUX2_X2 sll_384_M1_1_19 ( .A(sll_384_ML_int_1__19_), .B(
        sll_384_ML_int_1__17_), .S(sll_384_n6), .Z(sll_384_ML_int_2__19_) );
  MUX2_X2 sll_384_M1_1_20 ( .A(sll_384_ML_int_1__20_), .B(
        sll_384_ML_int_1__18_), .S(N141), .Z(sll_384_ML_int_2__20_) );
  MUX2_X2 sll_384_M1_1_21 ( .A(sll_384_ML_int_1__21_), .B(
        sll_384_ML_int_1__19_), .S(N141), .Z(sll_384_ML_int_2__21_) );
  MUX2_X2 sll_384_M1_1_22 ( .A(sll_384_ML_int_1__22_), .B(
        sll_384_ML_int_1__20_), .S(sll_384_n6), .Z(sll_384_ML_int_2__22_) );
  MUX2_X2 sll_384_M1_1_23 ( .A(sll_384_ML_int_1__23_), .B(
        sll_384_ML_int_1__21_), .S(N141), .Z(sll_384_ML_int_2__23_) );
  MUX2_X2 sll_384_M1_2_4 ( .A(sll_384_ML_int_2__4_), .B(sll_384_ML_int_2__0_), 
        .S(N107), .Z(sll_384_ML_int_3__4_) );
  MUX2_X2 sll_384_M1_2_5 ( .A(sll_384_ML_int_2__5_), .B(sll_384_ML_int_2__1_), 
        .S(N107), .Z(sll_384_ML_int_3__5_) );
  MUX2_X2 sll_384_M1_2_6 ( .A(sll_384_ML_int_2__6_), .B(sll_384_ML_int_2__2_), 
        .S(N107), .Z(sll_384_ML_int_3__6_) );
  MUX2_X2 sll_384_M1_2_7 ( .A(sll_384_ML_int_2__7_), .B(sll_384_ML_int_2__3_), 
        .S(N107), .Z(sll_384_ML_int_3__7_) );
  MUX2_X2 sll_384_M1_2_8 ( .A(sll_384_ML_int_2__8_), .B(sll_384_ML_int_2__4_), 
        .S(N107), .Z(sll_384_ML_int_3__8_) );
  MUX2_X2 sll_384_M1_2_9 ( .A(sll_384_ML_int_2__9_), .B(sll_384_ML_int_2__5_), 
        .S(N107), .Z(sll_384_ML_int_3__9_) );
  MUX2_X2 sll_384_M1_2_10 ( .A(sll_384_ML_int_2__10_), .B(sll_384_ML_int_2__6_), .S(N107), .Z(sll_384_ML_int_3__10_) );
  MUX2_X2 sll_384_M1_2_11 ( .A(sll_384_ML_int_2__11_), .B(sll_384_ML_int_2__7_), .S(N107), .Z(sll_384_ML_int_3__11_) );
  MUX2_X2 sll_384_M1_2_12 ( .A(sll_384_ML_int_2__12_), .B(sll_384_ML_int_2__8_), .S(N107), .Z(sll_384_ML_int_3__12_) );
  MUX2_X2 sll_384_M1_2_13 ( .A(sll_384_ML_int_2__13_), .B(sll_384_ML_int_2__9_), .S(N107), .Z(sll_384_ML_int_3__13_) );
  MUX2_X2 sll_384_M1_2_14 ( .A(sll_384_ML_int_2__14_), .B(
        sll_384_ML_int_2__10_), .S(N107), .Z(sll_384_ML_int_3__14_) );
  MUX2_X2 sll_384_M1_2_15 ( .A(sll_384_ML_int_2__15_), .B(
        sll_384_ML_int_2__11_), .S(N107), .Z(sll_384_ML_int_3__15_) );
  MUX2_X2 sll_384_M1_2_16 ( .A(sll_384_ML_int_2__16_), .B(
        sll_384_ML_int_2__12_), .S(N107), .Z(sll_384_ML_int_3__16_) );
  MUX2_X2 sll_384_M1_2_17 ( .A(sll_384_ML_int_2__17_), .B(
        sll_384_ML_int_2__13_), .S(N107), .Z(sll_384_ML_int_3__17_) );
  MUX2_X2 sll_384_M1_2_18 ( .A(sll_384_ML_int_2__18_), .B(
        sll_384_ML_int_2__14_), .S(N107), .Z(sll_384_ML_int_3__18_) );
  MUX2_X2 sll_384_M1_2_19 ( .A(sll_384_ML_int_2__19_), .B(
        sll_384_ML_int_2__15_), .S(N107), .Z(sll_384_ML_int_3__19_) );
  MUX2_X2 sll_384_M1_2_20 ( .A(sll_384_ML_int_2__20_), .B(
        sll_384_ML_int_2__16_), .S(N107), .Z(sll_384_ML_int_3__20_) );
  MUX2_X2 sll_384_M1_2_21 ( .A(sll_384_ML_int_2__21_), .B(
        sll_384_ML_int_2__17_), .S(N107), .Z(sll_384_ML_int_3__21_) );
  MUX2_X2 sll_384_M1_2_22 ( .A(sll_384_ML_int_2__22_), .B(
        sll_384_ML_int_2__18_), .S(N107), .Z(sll_384_ML_int_3__22_) );
  MUX2_X2 sll_384_M1_2_23 ( .A(sll_384_ML_int_2__23_), .B(
        sll_384_ML_int_2__19_), .S(N107), .Z(sll_384_ML_int_3__23_) );
  MUX2_X2 sll_384_M1_3_8 ( .A(sll_384_ML_int_3__8_), .B(sll_384_ML_int_3__0_), 
        .S(sll_384_n3), .Z(sll_384_ML_int_4__8_) );
  MUX2_X2 sll_384_M1_3_9 ( .A(sll_384_ML_int_3__9_), .B(sll_384_ML_int_3__1_), 
        .S(sll_384_n3), .Z(sll_384_ML_int_4__9_) );
  MUX2_X2 sll_384_M1_3_10 ( .A(sll_384_ML_int_3__10_), .B(sll_384_ML_int_3__2_), .S(sll_384_n3), .Z(sll_384_ML_int_4__10_) );
  MUX2_X2 sll_384_M1_3_11 ( .A(sll_384_ML_int_3__11_), .B(sll_384_ML_int_3__3_), .S(sll_384_n3), .Z(sll_384_ML_int_4__11_) );
  MUX2_X2 sll_384_M1_3_12 ( .A(sll_384_ML_int_3__12_), .B(sll_384_ML_int_3__4_), .S(sll_384_n3), .Z(sll_384_ML_int_4__12_) );
  MUX2_X2 sll_384_M1_3_13 ( .A(sll_384_ML_int_3__13_), .B(sll_384_ML_int_3__5_), .S(n2597), .Z(sll_384_ML_int_4__13_) );
  MUX2_X2 sll_384_M1_3_14 ( .A(sll_384_ML_int_3__14_), .B(sll_384_ML_int_3__6_), .S(n2597), .Z(sll_384_ML_int_4__14_) );
  MUX2_X2 sll_384_M1_3_15 ( .A(sll_384_ML_int_3__15_), .B(sll_384_ML_int_3__7_), .S(sll_384_n3), .Z(sll_384_ML_int_4__15_) );
  MUX2_X2 sll_384_M1_3_16 ( .A(sll_384_ML_int_3__16_), .B(sll_384_ML_int_3__8_), .S(sll_384_n3), .Z(sll_384_ML_int_4__16_) );
  MUX2_X2 sll_384_M1_3_17 ( .A(sll_384_ML_int_3__17_), .B(sll_384_ML_int_3__9_), .S(sll_384_n3), .Z(sll_384_ML_int_4__17_) );
  MUX2_X2 sll_384_M1_3_18 ( .A(sll_384_ML_int_3__18_), .B(
        sll_384_ML_int_3__10_), .S(sll_384_n3), .Z(sll_384_ML_int_4__18_) );
  MUX2_X2 sll_384_M1_3_19 ( .A(sll_384_ML_int_3__19_), .B(
        sll_384_ML_int_3__11_), .S(sll_384_n3), .Z(sll_384_ML_int_4__19_) );
  MUX2_X2 sll_384_M1_3_20 ( .A(sll_384_ML_int_3__20_), .B(
        sll_384_ML_int_3__12_), .S(sll_384_n3), .Z(sll_384_ML_int_4__20_) );
  MUX2_X2 sll_384_M1_3_21 ( .A(sll_384_ML_int_3__21_), .B(
        sll_384_ML_int_3__13_), .S(sll_384_n3), .Z(sll_384_ML_int_4__21_) );
  MUX2_X2 sll_384_M1_3_22 ( .A(sll_384_ML_int_3__22_), .B(
        sll_384_ML_int_3__14_), .S(sll_384_n3), .Z(sll_384_ML_int_4__22_) );
  MUX2_X2 sll_384_M1_3_23 ( .A(sll_384_ML_int_3__23_), .B(
        sll_384_ML_int_3__15_), .S(sll_384_n3), .Z(sll_384_ML_int_4__23_) );
  MUX2_X2 sll_384_M1_4_16 ( .A(sll_384_ML_int_4__16_), .B(sll_384_n8), .S(
        n2587), .Z(N188) );
  MUX2_X2 sll_384_M1_4_17 ( .A(sll_384_ML_int_4__17_), .B(sll_384_n12), .S(
        n2587), .Z(N189) );
  MUX2_X2 sll_384_M1_4_18 ( .A(sll_384_ML_int_4__18_), .B(sll_384_n10), .S(
        n2587), .Z(N190) );
  MUX2_X2 sll_384_M1_4_19 ( .A(sll_384_ML_int_4__19_), .B(sll_384_n14), .S(
        n2587), .Z(N191) );
  MUX2_X2 sll_384_M1_4_20 ( .A(sll_384_ML_int_4__20_), .B(sll_384_n9), .S(
        n2587), .Z(N192) );
  MUX2_X2 sll_384_M1_4_21 ( .A(sll_384_ML_int_4__21_), .B(sll_384_n13), .S(
        n2587), .Z(N193) );
  MUX2_X2 sll_384_M1_4_22 ( .A(sll_384_ML_int_4__22_), .B(sll_384_n11), .S(
        n2587), .Z(N194) );
  MUX2_X2 sll_384_M1_4_23 ( .A(sll_384_ML_int_4__23_), .B(sll_384_n15), .S(
        n2587), .Z(N195) );
  NAND2_X1 r473_U82 ( .A1(fracta_mul[20]), .A2(r473_n7), .ZN(r473_n37) );
  NAND2_X1 r473_U81 ( .A1(fracta_mul[19]), .A2(r473_n8), .ZN(r473_n36) );
  NAND2_X1 r473_U80 ( .A1(fracta_mul[18]), .A2(r473_n9), .ZN(r473_n41) );
  NAND2_X1 r473_U79 ( .A1(fracta_mul[17]), .A2(r473_n10), .ZN(r473_n39) );
  NAND2_X1 r473_U78 ( .A1(fracta_mul[16]), .A2(r473_n11), .ZN(r473_n40) );
  NAND2_X1 r473_U77 ( .A1(fracta_mul[15]), .A2(r473_n12), .ZN(r473_n43) );
  NAND2_X1 r473_U76 ( .A1(fracta_mul[14]), .A2(r473_n13), .ZN(r473_n45) );
  NAND2_X1 r473_U75 ( .A1(fracta_mul[13]), .A2(r473_n14), .ZN(r473_n44) );
  NAND2_X1 r473_U74 ( .A1(fracta_mul[12]), .A2(r473_n15), .ZN(r473_n48) );
  NAND2_X1 r473_U73 ( .A1(fracta_mul[11]), .A2(r473_n16), .ZN(r473_n46) );
  NAND2_X1 r473_U72 ( .A1(fracta_mul[10]), .A2(r473_n17), .ZN(r473_n47) );
  NAND2_X1 r473_U71 ( .A1(fracta_mul[9]), .A2(r473_n18), .ZN(r473_n50) );
  NAND2_X1 r473_U70 ( .A1(fracta_mul[8]), .A2(r473_n19), .ZN(r473_n52) );
  NAND2_X1 r473_U69 ( .A1(fracta_mul[7]), .A2(r473_n20), .ZN(r473_n51) );
  NAND2_X1 r473_U68 ( .A1(fracta_mul[6]), .A2(r473_n21), .ZN(r473_n56) );
  NAND2_X1 r473_U67 ( .A1(fracta_mul[5]), .A2(r473_n22), .ZN(r473_n58) );
  NAND2_X1 r473_U66 ( .A1(fracta_mul[4]), .A2(r473_n23), .ZN(r473_n57) );
  NAND2_X1 r473_U65 ( .A1(fracta_mul[3]), .A2(r473_n24), .ZN(r473_n54) );
  NOR2_X1 r473_U64 ( .A1(r473_n27), .A2(fracta_mul[0]), .ZN(r473_n80) );
  AOI21_X1 r473_U63 ( .B1(r473_n5), .B2(r473_n80), .A(u6_N1), .ZN(r473_n81) );
  OAI211_X1 r473_U62 ( .C1(r473_n80), .C2(r473_n5), .A(r473_n4), .B(r473_n53), 
        .ZN(r473_n79) );
  OAI221_X1 r473_U61 ( .B1(fracta_mul[2]), .B2(r473_n25), .C1(fracta_mul[3]), 
        .C2(r473_n24), .A(r473_n79), .ZN(r473_n78) );
  NAND3_X1 r473_U60 ( .A1(r473_n57), .A2(r473_n54), .A3(r473_n78), .ZN(
        r473_n77) );
  OAI221_X1 r473_U59 ( .B1(fracta_mul[4]), .B2(r473_n23), .C1(fracta_mul[5]), 
        .C2(r473_n22), .A(r473_n77), .ZN(r473_n76) );
  NAND3_X1 r473_U58 ( .A1(r473_n56), .A2(r473_n58), .A3(r473_n76), .ZN(
        r473_n75) );
  OAI221_X1 r473_U57 ( .B1(fracta_mul[6]), .B2(r473_n21), .C1(fracta_mul[7]), 
        .C2(r473_n20), .A(r473_n75), .ZN(r473_n74) );
  NAND3_X1 r473_U56 ( .A1(r473_n52), .A2(r473_n51), .A3(r473_n74), .ZN(
        r473_n73) );
  OAI221_X1 r473_U55 ( .B1(fracta_mul[8]), .B2(r473_n19), .C1(fracta_mul[9]), 
        .C2(r473_n18), .A(r473_n73), .ZN(r473_n72) );
  NAND3_X1 r473_U54 ( .A1(r473_n47), .A2(r473_n50), .A3(r473_n72), .ZN(
        r473_n71) );
  OAI221_X1 r473_U53 ( .B1(fracta_mul[10]), .B2(r473_n17), .C1(fracta_mul[11]), 
        .C2(r473_n16), .A(r473_n71), .ZN(r473_n70) );
  NAND3_X1 r473_U52 ( .A1(r473_n48), .A2(r473_n46), .A3(r473_n70), .ZN(
        r473_n69) );
  OAI221_X1 r473_U51 ( .B1(fracta_mul[12]), .B2(r473_n15), .C1(fracta_mul[13]), 
        .C2(r473_n14), .A(r473_n69), .ZN(r473_n68) );
  NAND3_X1 r473_U50 ( .A1(r473_n45), .A2(r473_n44), .A3(r473_n68), .ZN(
        r473_n67) );
  OAI221_X1 r473_U49 ( .B1(fracta_mul[14]), .B2(r473_n13), .C1(fracta_mul[15]), 
        .C2(r473_n12), .A(r473_n67), .ZN(r473_n66) );
  NAND3_X1 r473_U48 ( .A1(r473_n40), .A2(r473_n43), .A3(r473_n66), .ZN(
        r473_n65) );
  OAI221_X1 r473_U47 ( .B1(fracta_mul[16]), .B2(r473_n11), .C1(fracta_mul[17]), 
        .C2(r473_n10), .A(r473_n65), .ZN(r473_n64) );
  NAND3_X1 r473_U46 ( .A1(r473_n41), .A2(r473_n39), .A3(r473_n64), .ZN(
        r473_n63) );
  OAI221_X1 r473_U45 ( .B1(fracta_mul[18]), .B2(r473_n9), .C1(fracta_mul[19]), 
        .C2(r473_n8), .A(r473_n63), .ZN(r473_n62) );
  NAND3_X1 r473_U44 ( .A1(r473_n37), .A2(r473_n36), .A3(r473_n62), .ZN(
        r473_n61) );
  OAI221_X1 r473_U43 ( .B1(fracta_mul[20]), .B2(r473_n7), .C1(fracta_mul[21]), 
        .C2(r473_n6), .A(r473_n61), .ZN(r473_n60) );
  NAND2_X1 r473_U42 ( .A1(fracta_mul[21]), .A2(r473_n6), .ZN(r473_n35) );
  AND3_X1 r473_U41 ( .A1(r473_n56), .A2(r473_n57), .A3(r473_n58), .ZN(r473_n55) );
  NAND4_X1 r473_U40 ( .A1(r473_n53), .A2(r473_n28), .A3(r473_n54), .A4(
        r473_n55), .ZN(r473_n29) );
  AND3_X1 r473_U39 ( .A1(r473_n50), .A2(r473_n51), .A3(r473_n52), .ZN(r473_n49) );
  NAND4_X1 r473_U38 ( .A1(r473_n46), .A2(r473_n47), .A3(r473_n48), .A4(
        r473_n49), .ZN(r473_n30) );
  AND3_X1 r473_U37 ( .A1(r473_n43), .A2(r473_n44), .A3(r473_n45), .ZN(r473_n42) );
  NAND4_X1 r473_U36 ( .A1(r473_n39), .A2(r473_n40), .A3(r473_n41), .A4(
        r473_n42), .ZN(r473_n31) );
  AND2_X1 r473_U35 ( .A1(fracta_mul[0]), .A2(r473_n27), .ZN(r473_n38) );
  OAI22_X1 r473_U34 ( .A1(n2586), .A2(r473_n38), .B1(r473_n38), .B2(r473_n26), 
        .ZN(r473_n33) );
  AND3_X1 r473_U33 ( .A1(r473_n35), .A2(r473_n36), .A3(r473_n37), .ZN(r473_n34) );
  OAI211_X1 r473_U32 ( .C1(u6_N22), .C2(r473_n3), .A(r473_n33), .B(r473_n34), 
        .ZN(r473_n32) );
  NOR4_X1 r473_U31 ( .A1(r473_n29), .A2(r473_n30), .A3(r473_n31), .A4(r473_n32), .ZN(u1_N131) );
  INV_X4 r473_U30 ( .A(u6_N0), .ZN(r473_n27) );
  INV_X4 r473_U29 ( .A(u6_N1), .ZN(r473_n26) );
  INV_X4 r473_U28 ( .A(u6_N2), .ZN(r473_n25) );
  INV_X4 r473_U27 ( .A(u6_N3), .ZN(r473_n24) );
  INV_X4 r473_U26 ( .A(u6_N4), .ZN(r473_n23) );
  INV_X4 r473_U25 ( .A(u6_N5), .ZN(r473_n22) );
  INV_X4 r473_U24 ( .A(u6_N9), .ZN(r473_n18) );
  INV_X4 r473_U23 ( .A(n3049), .ZN(r473_n6) );
  INV_X4 r473_U22 ( .A(r473_n81), .ZN(r473_n4) );
  INV_X4 r473_U21 ( .A(fracta_mul[22]), .ZN(r473_n3) );
  INV_X4 r473_U20 ( .A(r473_n59), .ZN(r473_n2) );
  INV_X4 r473_U19 ( .A(r473_n28), .ZN(u1_N130) );
  OAI211_X2 r473_U18 ( .C1(u6_N22), .C2(r473_n3), .A(r473_n60), .B(r473_n35), 
        .ZN(r473_n59) );
  AOI21_X4 r473_U17 ( .B1(r473_n3), .B2(u6_N22), .A(r473_n2), .ZN(r473_n28) );
  INV_X1 r473_U16 ( .A(n2586), .ZN(r473_n5) );
  INV_X1 r473_U15 ( .A(n3040), .ZN(r473_n7) );
  INV_X1 r473_U14 ( .A(u6_N18), .ZN(r473_n9) );
  NAND2_X2 r473_U13 ( .A1(fracta_mul[2]), .A2(r473_n25), .ZN(r473_n53) );
  INV_X1 r473_U12 ( .A(u6_N17), .ZN(r473_n10) );
  INV_X1 r473_U11 ( .A(n2963), .ZN(r473_n11) );
  INV_X1 r473_U10 ( .A(u6_N13), .ZN(r473_n14) );
  INV_X1 r473_U9 ( .A(n2968), .ZN(r473_n8) );
  INV_X1 r473_U8 ( .A(n2986), .ZN(r473_n15) );
  INV_X1 r473_U7 ( .A(n2982), .ZN(r473_n16) );
  INV_X1 r473_U6 ( .A(n2672), .ZN(r473_n13) );
  INV_X2 r473_U5 ( .A(u6_N8), .ZN(r473_n19) );
  INV_X2 r473_U4 ( .A(u6_N10), .ZN(r473_n17) );
  INV_X1 r473_U3 ( .A(u6_N15), .ZN(r473_n12) );
  INV_X1 r473_U2 ( .A(u6_N7), .ZN(r473_n20) );
  INV_X1 r473_U1 ( .A(u6_N6), .ZN(r473_n21) );
  INV_X4 sub_1_root_sub_0_root_u4_add_496_U17 ( .A(div_opa_ldz_r2[1]), .ZN(
        sub_1_root_sub_0_root_u4_add_496_n9) );
  INV_X4 sub_1_root_sub_0_root_u4_add_496_U16 ( .A(div_opa_ldz_r2[2]), .ZN(
        sub_1_root_sub_0_root_u4_add_496_n8) );
  INV_X4 sub_1_root_sub_0_root_u4_add_496_U15 ( .A(div_opa_ldz_r2[3]), .ZN(
        sub_1_root_sub_0_root_u4_add_496_n7) );
  INV_X4 sub_1_root_sub_0_root_u4_add_496_U14 ( .A(div_opa_ldz_r2[4]), .ZN(
        sub_1_root_sub_0_root_u4_add_496_n6) );
  XNOR2_X2 sub_1_root_sub_0_root_u4_add_496_U13 ( .A(
        sub_1_root_sub_0_root_u4_add_496_n10), .B(net85905), .ZN(u4_ldz_dif_0_) );
  NAND2_X2 sub_1_root_sub_0_root_u4_add_496_U12 ( .A1(div_opa_ldz_r2[0]), .A2(
        sub_1_root_sub_0_root_u4_add_496_n5), .ZN(
        sub_1_root_sub_0_root_u4_add_496_carry_1_) );
  XNOR2_X2 sub_1_root_sub_0_root_u4_add_496_U11 ( .A(net85937), .B(
        sub_1_root_sub_0_root_u4_add_496_carry_7_), .ZN(u4_ldz_dif_7_) );
  INV_X4 sub_1_root_sub_0_root_u4_add_496_U10 ( .A(
        sub_1_root_sub_0_root_u4_add_496_carry_6_), .ZN(
        sub_1_root_sub_0_root_u4_add_496_n4) );
  INV_X4 sub_1_root_sub_0_root_u4_add_496_U9 ( .A(net85933), .ZN(
        sub_1_root_sub_0_root_u4_add_496_n3) );
  XNOR2_X2 sub_1_root_sub_0_root_u4_add_496_U8 ( .A(net85933), .B(
        sub_1_root_sub_0_root_u4_add_496_carry_6_), .ZN(u4_ldz_dif_6_) );
  NAND2_X2 sub_1_root_sub_0_root_u4_add_496_U7 ( .A1(
        sub_1_root_sub_0_root_u4_add_496_n3), .A2(
        sub_1_root_sub_0_root_u4_add_496_n4), .ZN(
        sub_1_root_sub_0_root_u4_add_496_carry_7_) );
  INV_X4 sub_1_root_sub_0_root_u4_add_496_U6 ( .A(
        sub_1_root_sub_0_root_u4_add_496_carry_5_), .ZN(
        sub_1_root_sub_0_root_u4_add_496_n2) );
  INV_X4 sub_1_root_sub_0_root_u4_add_496_U5 ( .A(net85929), .ZN(
        sub_1_root_sub_0_root_u4_add_496_n1) );
  XNOR2_X2 sub_1_root_sub_0_root_u4_add_496_U4 ( .A(net85929), .B(
        sub_1_root_sub_0_root_u4_add_496_carry_5_), .ZN(u4_ldz_dif_5_) );
  NAND2_X2 sub_1_root_sub_0_root_u4_add_496_U3 ( .A1(
        sub_1_root_sub_0_root_u4_add_496_n1), .A2(
        sub_1_root_sub_0_root_u4_add_496_n2), .ZN(
        sub_1_root_sub_0_root_u4_add_496_carry_6_) );
  INV_X2 sub_1_root_sub_0_root_u4_add_496_U2 ( .A(net85905), .ZN(
        sub_1_root_sub_0_root_u4_add_496_n5) );
  INV_X1 sub_1_root_sub_0_root_u4_add_496_U1 ( .A(div_opa_ldz_r2[0]), .ZN(
        sub_1_root_sub_0_root_u4_add_496_n10) );
  FA_X1 sub_1_root_sub_0_root_u4_add_496_U2_1 ( .A(n3091), .B(
        sub_1_root_sub_0_root_u4_add_496_n9), .CI(
        sub_1_root_sub_0_root_u4_add_496_carry_1_), .CO(
        sub_1_root_sub_0_root_u4_add_496_carry_2_), .S(u4_ldz_dif_1_) );
  FA_X1 sub_1_root_sub_0_root_u4_add_496_U2_2 ( .A(n3089), .B(
        sub_1_root_sub_0_root_u4_add_496_n8), .CI(
        sub_1_root_sub_0_root_u4_add_496_carry_2_), .CO(
        sub_1_root_sub_0_root_u4_add_496_carry_3_), .S(u4_ldz_dif_2_) );
  FA_X1 sub_1_root_sub_0_root_u4_add_496_U2_3 ( .A(n3088), .B(
        sub_1_root_sub_0_root_u4_add_496_n7), .CI(
        sub_1_root_sub_0_root_u4_add_496_carry_3_), .CO(
        sub_1_root_sub_0_root_u4_add_496_carry_4_), .S(u4_ldz_dif_3_) );
  FA_X1 sub_1_root_sub_0_root_u4_add_496_U2_4 ( .A(n3085), .B(
        sub_1_root_sub_0_root_u4_add_496_n6), .CI(
        sub_1_root_sub_0_root_u4_add_496_carry_4_), .CO(
        sub_1_root_sub_0_root_u4_add_496_carry_5_), .S(u4_ldz_dif_4_) );
  INV_X4 u5_mult_79_U3136 ( .A(fracta_mul[22]), .ZN(u5_mult_79_n1859) );
  INV_X4 u5_mult_79_U3135 ( .A(fracta_mul[21]), .ZN(u5_mult_79_n1857) );
  INV_X4 u5_mult_79_U3134 ( .A(fracta_mul[20]), .ZN(u5_mult_79_n1856) );
  NOR2_X4 u5_mult_79_U3133 ( .A1(u5_mult_79_n1818), .A2(u5_mult_79_n1773), 
        .ZN(u5_mult_79_ab_19__5_) );
  NOR2_X4 u5_mult_79_U3132 ( .A1(u5_mult_79_n1812), .A2(u5_mult_79_n1773), 
        .ZN(u5_mult_79_ab_19__7_) );
  NOR2_X4 u5_mult_79_U3131 ( .A1(u5_mult_79_n1794), .A2(u5_mult_79_n1773), 
        .ZN(u5_mult_79_ab_19__16_) );
  NOR2_X4 u5_mult_79_U3130 ( .A1(u5_mult_79_n1791), .A2(u5_mult_79_n1773), 
        .ZN(u5_mult_79_ab_19__17_) );
  NOR2_X4 u5_mult_79_U3129 ( .A1(u5_mult_79_n1788), .A2(u5_mult_79_n1773), 
        .ZN(u5_mult_79_ab_19__18_) );
  NOR2_X4 u5_mult_79_U3128 ( .A1(u5_mult_79_n1785), .A2(u5_mult_79_n1773), 
        .ZN(u5_mult_79_ab_19__19_) );
  NOR2_X4 u5_mult_79_U3127 ( .A1(u5_mult_79_n1783), .A2(u5_mult_79_n1773), 
        .ZN(u5_mult_79_ab_19__21_) );
  INV_X4 u5_mult_79_U3126 ( .A(fracta_mul[19]), .ZN(u5_mult_79_n1855) );
  NOR2_X4 u5_mult_79_U3125 ( .A1(u5_mult_79_n1815), .A2(u5_mult_79_n1770), 
        .ZN(u5_mult_79_ab_18__6_) );
  NOR2_X4 u5_mult_79_U3124 ( .A1(u5_mult_79_n1812), .A2(u5_mult_79_n1770), 
        .ZN(u5_mult_79_ab_18__7_) );
  NOR2_X4 u5_mult_79_U3123 ( .A1(u5_mult_79_n1809), .A2(u5_mult_79_n1770), 
        .ZN(u5_mult_79_ab_18__8_) );
  NOR2_X4 u5_mult_79_U3122 ( .A1(u5_mult_79_n1806), .A2(u5_mult_79_n1770), 
        .ZN(u5_mult_79_ab_18__9_) );
  NOR2_X4 u5_mult_79_U3121 ( .A1(u5_mult_79_n1801), .A2(u5_mult_79_n1771), 
        .ZN(u5_mult_79_ab_18__11_) );
  NOR2_X4 u5_mult_79_U3120 ( .A1(u5_mult_79_n1868), .A2(u5_mult_79_n1771), 
        .ZN(u5_mult_79_ab_18__13_) );
  NOR2_X4 u5_mult_79_U3119 ( .A1(u5_mult_79_n1867), .A2(u5_mult_79_n1771), 
        .ZN(u5_mult_79_ab_18__14_) );
  NOR2_X4 u5_mult_79_U3118 ( .A1(u5_mult_79_n1794), .A2(u5_mult_79_n1771), 
        .ZN(u5_mult_79_ab_18__16_) );
  NOR2_X4 u5_mult_79_U3117 ( .A1(u5_mult_79_n1788), .A2(u5_mult_79_n1771), 
        .ZN(u5_mult_79_ab_18__18_) );
  NOR2_X4 u5_mult_79_U3116 ( .A1(u5_mult_79_n1338), .A2(u5_mult_79_n1771), 
        .ZN(u5_mult_79_ab_18__20_) );
  NOR2_X4 u5_mult_79_U3115 ( .A1(u5_mult_79_n1783), .A2(u5_mult_79_n1771), 
        .ZN(u5_mult_79_ab_18__21_) );
  NOR2_X4 u5_mult_79_U3114 ( .A1(u5_mult_79_n1832), .A2(u5_mult_79_n1767), 
        .ZN(u5_mult_79_ab_17__23_) );
  NOR2_X4 u5_mult_79_U3113 ( .A1(u5_mult_79_n1781), .A2(u5_mult_79_n1771), 
        .ZN(u5_mult_79_ab_18__22_) );
  INV_X4 u5_mult_79_U3112 ( .A(fracta_mul[18]), .ZN(u5_mult_79_n1854) );
  NOR2_X4 u5_mult_79_U3111 ( .A1(u5_mult_79_n1826), .A2(u5_mult_79_n1767), 
        .ZN(u5_mult_79_ab_17__2_) );
  NOR2_X4 u5_mult_79_U3110 ( .A1(u5_mult_79_n1823), .A2(u5_mult_79_n1767), 
        .ZN(u5_mult_79_ab_17__3_) );
  NOR2_X4 u5_mult_79_U3109 ( .A1(u5_mult_79_n1809), .A2(u5_mult_79_n1767), 
        .ZN(u5_mult_79_ab_17__8_) );
  NOR2_X4 u5_mult_79_U3108 ( .A1(u5_mult_79_n1806), .A2(u5_mult_79_n1767), 
        .ZN(u5_mult_79_ab_17__9_) );
  NOR2_X4 u5_mult_79_U3107 ( .A1(u5_mult_79_n1803), .A2(u5_mult_79_n1767), 
        .ZN(u5_mult_79_ab_17__10_) );
  NOR2_X4 u5_mult_79_U3106 ( .A1(u5_mult_79_n1801), .A2(u5_mult_79_n1768), 
        .ZN(u5_mult_79_ab_17__11_) );
  NOR2_X4 u5_mult_79_U3105 ( .A1(u5_mult_79_n1796), .A2(u5_mult_79_n1768), 
        .ZN(u5_mult_79_ab_17__15_) );
  NOR2_X4 u5_mult_79_U3104 ( .A1(u5_mult_79_n1791), .A2(u5_mult_79_n1768), 
        .ZN(u5_mult_79_ab_17__17_) );
  NOR2_X4 u5_mult_79_U3103 ( .A1(u5_mult_79_n1785), .A2(u5_mult_79_n1768), 
        .ZN(u5_mult_79_ab_17__19_) );
  NOR2_X4 u5_mult_79_U3102 ( .A1(u5_mult_79_n1338), .A2(u5_mult_79_n1768), 
        .ZN(u5_mult_79_ab_17__20_) );
  INV_X4 u5_mult_79_U3101 ( .A(fracta_mul[17]), .ZN(u5_mult_79_n1853) );
  NOR2_X4 u5_mult_79_U3100 ( .A1(u5_mult_79_n1834), .A2(u5_mult_79_n1764), 
        .ZN(u5_mult_79_ab_16__0_) );
  NOR2_X4 u5_mult_79_U3099 ( .A1(u5_mult_79_n1823), .A2(u5_mult_79_n1764), 
        .ZN(u5_mult_79_ab_16__3_) );
  NOR2_X4 u5_mult_79_U3098 ( .A1(u5_mult_79_n1821), .A2(u5_mult_79_n1764), 
        .ZN(u5_mult_79_ab_16__4_) );
  NOR2_X4 u5_mult_79_U3097 ( .A1(u5_mult_79_n1812), .A2(u5_mult_79_n1764), 
        .ZN(u5_mult_79_ab_16__7_) );
  NOR2_X4 u5_mult_79_U3096 ( .A1(u5_mult_79_n1809), .A2(u5_mult_79_n1764), 
        .ZN(u5_mult_79_ab_16__8_) );
  NOR2_X4 u5_mult_79_U3095 ( .A1(u5_mult_79_n1803), .A2(u5_mult_79_n1764), 
        .ZN(u5_mult_79_ab_16__10_) );
  NOR2_X4 u5_mult_79_U3094 ( .A1(u5_mult_79_n1801), .A2(u5_mult_79_n1765), 
        .ZN(u5_mult_79_ab_16__11_) );
  NOR2_X4 u5_mult_79_U3093 ( .A1(u5_mult_79_n1868), .A2(u5_mult_79_n1765), 
        .ZN(u5_mult_79_ab_16__13_) );
  NOR2_X4 u5_mult_79_U3092 ( .A1(u5_mult_79_n1796), .A2(u5_mult_79_n1765), 
        .ZN(u5_mult_79_ab_16__15_) );
  NOR2_X4 u5_mult_79_U3091 ( .A1(u5_mult_79_n1791), .A2(u5_mult_79_n1765), 
        .ZN(u5_mult_79_ab_16__17_) );
  NOR2_X4 u5_mult_79_U3090 ( .A1(u5_mult_79_n1783), .A2(u5_mult_79_n1765), 
        .ZN(u5_mult_79_ab_16__21_) );
  INV_X4 u5_mult_79_U3089 ( .A(fracta_mul[16]), .ZN(u5_mult_79_n1852) );
  NOR2_X4 u5_mult_79_U3088 ( .A1(u5_mult_79_n1821), .A2(u5_mult_79_n1761), 
        .ZN(u5_mult_79_ab_15__4_) );
  NOR2_X4 u5_mult_79_U3087 ( .A1(u5_mult_79_n1818), .A2(u5_mult_79_n1761), 
        .ZN(u5_mult_79_ab_15__5_) );
  NOR2_X4 u5_mult_79_U3086 ( .A1(u5_mult_79_n1815), .A2(u5_mult_79_n1761), 
        .ZN(u5_mult_79_ab_15__6_) );
  NOR2_X4 u5_mult_79_U3085 ( .A1(u5_mult_79_n1812), .A2(u5_mult_79_n1761), 
        .ZN(u5_mult_79_ab_15__7_) );
  NOR2_X4 u5_mult_79_U3084 ( .A1(u5_mult_79_n1809), .A2(u5_mult_79_n1761), 
        .ZN(u5_mult_79_ab_15__8_) );
  NOR2_X4 u5_mult_79_U3083 ( .A1(u5_mult_79_n1806), .A2(u5_mult_79_n1761), 
        .ZN(u5_mult_79_ab_15__9_) );
  NOR2_X4 u5_mult_79_U3082 ( .A1(u5_mult_79_n1801), .A2(u5_mult_79_n1762), 
        .ZN(u5_mult_79_ab_15__11_) );
  NOR2_X4 u5_mult_79_U3081 ( .A1(u5_mult_79_n1799), .A2(u5_mult_79_n1762), 
        .ZN(u5_mult_79_ab_15__12_) );
  NOR2_X4 u5_mult_79_U3080 ( .A1(u5_mult_79_n1796), .A2(u5_mult_79_n1762), 
        .ZN(u5_mult_79_ab_15__15_) );
  NOR2_X4 u5_mult_79_U3079 ( .A1(u5_mult_79_n1794), .A2(u5_mult_79_n1762), 
        .ZN(u5_mult_79_ab_15__16_) );
  NOR2_X4 u5_mult_79_U3078 ( .A1(u5_mult_79_n1788), .A2(u5_mult_79_n1762), 
        .ZN(u5_mult_79_ab_15__18_) );
  NOR2_X4 u5_mult_79_U3077 ( .A1(u5_mult_79_n1785), .A2(u5_mult_79_n1762), 
        .ZN(u5_mult_79_ab_15__19_) );
  INV_X4 u5_mult_79_U3076 ( .A(fracta_mul[15]), .ZN(u5_mult_79_n1851) );
  NOR2_X4 u5_mult_79_U3075 ( .A1(u5_mult_79_n1828), .A2(u5_mult_79_n1758), 
        .ZN(u5_mult_79_ab_14__1_) );
  NOR2_X4 u5_mult_79_U3074 ( .A1(u5_mult_79_n1823), .A2(u5_mult_79_n1758), 
        .ZN(u5_mult_79_ab_14__3_) );
  NOR2_X4 u5_mult_79_U3073 ( .A1(u5_mult_79_n1821), .A2(u5_mult_79_n1758), 
        .ZN(u5_mult_79_ab_14__4_) );
  NOR2_X4 u5_mult_79_U3072 ( .A1(u5_mult_79_n1818), .A2(u5_mult_79_n1758), 
        .ZN(u5_mult_79_ab_14__5_) );
  NOR2_X4 u5_mult_79_U3071 ( .A1(u5_mult_79_n1815), .A2(u5_mult_79_n1758), 
        .ZN(u5_mult_79_ab_14__6_) );
  NOR2_X4 u5_mult_79_U3070 ( .A1(u5_mult_79_n1812), .A2(u5_mult_79_n1758), 
        .ZN(u5_mult_79_ab_14__7_) );
  NOR2_X4 u5_mult_79_U3069 ( .A1(u5_mult_79_n1809), .A2(u5_mult_79_n1758), 
        .ZN(u5_mult_79_ab_14__8_) );
  NOR2_X4 u5_mult_79_U3068 ( .A1(u5_mult_79_n1799), .A2(u5_mult_79_n1759), 
        .ZN(u5_mult_79_ab_14__12_) );
  NOR2_X4 u5_mult_79_U3067 ( .A1(u5_mult_79_n1794), .A2(u5_mult_79_n1759), 
        .ZN(u5_mult_79_ab_14__16_) );
  NOR2_X4 u5_mult_79_U3066 ( .A1(u5_mult_79_n1791), .A2(u5_mult_79_n1759), 
        .ZN(u5_mult_79_ab_14__17_) );
  NOR2_X4 u5_mult_79_U3065 ( .A1(u5_mult_79_n1338), .A2(u5_mult_79_n1759), 
        .ZN(u5_mult_79_ab_14__20_) );
  NOR2_X4 u5_mult_79_U3064 ( .A1(u5_mult_79_n1783), .A2(u5_mult_79_n1759), 
        .ZN(u5_mult_79_ab_14__21_) );
  NOR2_X4 u5_mult_79_U3063 ( .A1(u5_mult_79_n1832), .A2(u5_mult_79_n1755), 
        .ZN(u5_mult_79_ab_13__23_) );
  INV_X4 u5_mult_79_U3062 ( .A(fracta_mul[14]), .ZN(u5_mult_79_n1850) );
  NOR2_X4 u5_mult_79_U3061 ( .A1(u5_mult_79_n1818), .A2(u5_mult_79_n1755), 
        .ZN(u5_mult_79_ab_13__5_) );
  NOR2_X4 u5_mult_79_U3060 ( .A1(u5_mult_79_n1815), .A2(u5_mult_79_n1755), 
        .ZN(u5_mult_79_ab_13__6_) );
  NOR2_X4 u5_mult_79_U3059 ( .A1(u5_mult_79_n1809), .A2(u5_mult_79_n1755), 
        .ZN(u5_mult_79_ab_13__8_) );
  NOR2_X4 u5_mult_79_U3058 ( .A1(u5_mult_79_n1868), .A2(u5_mult_79_n1756), 
        .ZN(u5_mult_79_ab_13__13_) );
  NOR2_X4 u5_mult_79_U3057 ( .A1(u5_mult_79_n1788), .A2(u5_mult_79_n1756), 
        .ZN(u5_mult_79_ab_13__18_) );
  NOR2_X4 u5_mult_79_U3056 ( .A1(u5_mult_79_n1781), .A2(u5_mult_79_n1756), 
        .ZN(u5_mult_79_ab_13__22_) );
  INV_X4 u5_mult_79_U3055 ( .A(fracta_mul[13]), .ZN(u5_mult_79_n1849) );
  NOR2_X4 u5_mult_79_U3054 ( .A1(u5_mult_79_n1815), .A2(u5_mult_79_n1752), 
        .ZN(u5_mult_79_ab_12__6_) );
  NOR2_X4 u5_mult_79_U3053 ( .A1(u5_mult_79_n1809), .A2(u5_mult_79_n1752), 
        .ZN(u5_mult_79_ab_12__8_) );
  NOR2_X4 u5_mult_79_U3052 ( .A1(u5_mult_79_n1806), .A2(u5_mult_79_n1752), 
        .ZN(u5_mult_79_ab_12__9_) );
  NOR2_X4 u5_mult_79_U3051 ( .A1(u5_mult_79_n1801), .A2(u5_mult_79_n1753), 
        .ZN(u5_mult_79_ab_12__11_) );
  NOR2_X4 u5_mult_79_U3050 ( .A1(u5_mult_79_n1868), .A2(u5_mult_79_n1753), 
        .ZN(u5_mult_79_ab_12__13_) );
  NOR2_X4 u5_mult_79_U3049 ( .A1(u5_mult_79_n1796), .A2(u5_mult_79_n1753), 
        .ZN(u5_mult_79_ab_12__15_) );
  NOR2_X4 u5_mult_79_U3048 ( .A1(u5_mult_79_n1794), .A2(u5_mult_79_n1753), 
        .ZN(u5_mult_79_ab_12__16_) );
  NOR2_X4 u5_mult_79_U3047 ( .A1(u5_mult_79_n1338), .A2(u5_mult_79_n1753), 
        .ZN(u5_mult_79_ab_12__20_) );
  INV_X4 u5_mult_79_U3046 ( .A(fracta_mul[12]), .ZN(u5_mult_79_n1848) );
  NOR2_X4 u5_mult_79_U3045 ( .A1(u5_mult_79_n1815), .A2(u5_mult_79_n1749), 
        .ZN(u5_mult_79_ab_11__6_) );
  NOR2_X4 u5_mult_79_U3044 ( .A1(u5_mult_79_n1812), .A2(u5_mult_79_n1749), 
        .ZN(u5_mult_79_ab_11__7_) );
  NOR2_X4 u5_mult_79_U3043 ( .A1(u5_mult_79_n1809), .A2(u5_mult_79_n1749), 
        .ZN(u5_mult_79_ab_11__8_) );
  NOR2_X4 u5_mult_79_U3042 ( .A1(u5_mult_79_n1806), .A2(u5_mult_79_n1749), 
        .ZN(u5_mult_79_ab_11__9_) );
  NOR2_X4 u5_mult_79_U3041 ( .A1(u5_mult_79_n1803), .A2(u5_mult_79_n1749), 
        .ZN(u5_mult_79_ab_11__10_) );
  NOR2_X4 u5_mult_79_U3040 ( .A1(u5_mult_79_n1799), .A2(u5_mult_79_n1750), 
        .ZN(u5_mult_79_ab_11__12_) );
  NOR2_X4 u5_mult_79_U3039 ( .A1(u5_mult_79_n1868), .A2(u5_mult_79_n1750), 
        .ZN(u5_mult_79_ab_11__13_) );
  NOR2_X4 u5_mult_79_U3038 ( .A1(u5_mult_79_n1794), .A2(u5_mult_79_n1750), 
        .ZN(u5_mult_79_ab_11__16_) );
  NOR2_X4 u5_mult_79_U3037 ( .A1(u5_mult_79_n1791), .A2(u5_mult_79_n1750), 
        .ZN(u5_mult_79_ab_11__17_) );
  NOR2_X4 u5_mult_79_U3036 ( .A1(u5_mult_79_n1788), .A2(u5_mult_79_n1750), 
        .ZN(u5_mult_79_ab_11__18_) );
  NOR2_X4 u5_mult_79_U3035 ( .A1(u5_mult_79_n1785), .A2(u5_mult_79_n1750), 
        .ZN(u5_mult_79_ab_11__19_) );
  NOR2_X4 u5_mult_79_U3034 ( .A1(u5_mult_79_n1338), .A2(u5_mult_79_n1750), 
        .ZN(u5_mult_79_ab_11__20_) );
  NOR2_X4 u5_mult_79_U3033 ( .A1(u5_mult_79_n1781), .A2(u5_mult_79_n1750), 
        .ZN(u5_mult_79_ab_11__22_) );
  INV_X4 u5_mult_79_U3032 ( .A(fracta_mul[11]), .ZN(u5_mult_79_n1847) );
  NOR2_X4 u5_mult_79_U3031 ( .A1(u5_mult_79_n1820), .A2(u5_mult_79_n1746), 
        .ZN(u5_mult_79_ab_10__4_) );
  NOR2_X4 u5_mult_79_U3030 ( .A1(u5_mult_79_n1805), .A2(u5_mult_79_n1746), 
        .ZN(u5_mult_79_ab_10__9_) );
  NOR2_X4 u5_mult_79_U3029 ( .A1(u5_mult_79_n1800), .A2(u5_mult_79_n1747), 
        .ZN(u5_mult_79_ab_10__11_) );
  NOR2_X4 u5_mult_79_U3028 ( .A1(u5_mult_79_n1798), .A2(u5_mult_79_n1747), 
        .ZN(u5_mult_79_ab_10__12_) );
  NOR2_X4 u5_mult_79_U3027 ( .A1(u5_mult_79_n1796), .A2(u5_mult_79_n1747), 
        .ZN(u5_mult_79_ab_10__15_) );
  NOR2_X4 u5_mult_79_U3026 ( .A1(u5_mult_79_n1338), .A2(u5_mult_79_n1747), 
        .ZN(u5_mult_79_ab_10__20_) );
  INV_X4 u5_mult_79_U3025 ( .A(fracta_mul[10]), .ZN(u5_mult_79_n1846) );
  NOR2_X4 u5_mult_79_U3024 ( .A1(u5_mult_79_n1817), .A2(u5_mult_79_n1743), 
        .ZN(u5_mult_79_ab_9__5_) );
  NOR2_X4 u5_mult_79_U3023 ( .A1(u5_mult_79_n1811), .A2(u5_mult_79_n1743), 
        .ZN(u5_mult_79_ab_9__7_) );
  NOR2_X4 u5_mult_79_U3022 ( .A1(u5_mult_79_n1868), .A2(u5_mult_79_n1744), 
        .ZN(u5_mult_79_ab_9__13_) );
  NOR2_X4 u5_mult_79_U3021 ( .A1(u5_mult_79_n1796), .A2(u5_mult_79_n1744), 
        .ZN(u5_mult_79_ab_9__15_) );
  NOR2_X4 u5_mult_79_U3020 ( .A1(u5_mult_79_n1793), .A2(u5_mult_79_n1744), 
        .ZN(u5_mult_79_ab_9__16_) );
  NOR2_X4 u5_mult_79_U3019 ( .A1(u5_mult_79_n1790), .A2(u5_mult_79_n1744), 
        .ZN(u5_mult_79_ab_9__17_) );
  INV_X4 u5_mult_79_U3018 ( .A(fracta_mul[9]), .ZN(u5_mult_79_n1845) );
  NOR2_X4 u5_mult_79_U3017 ( .A1(u5_mult_79_n1825), .A2(u5_mult_79_n1740), 
        .ZN(u5_mult_79_ab_8__2_) );
  NOR2_X4 u5_mult_79_U3016 ( .A1(u5_mult_79_n1823), .A2(u5_mult_79_n1740), 
        .ZN(u5_mult_79_ab_8__3_) );
  NOR2_X4 u5_mult_79_U3015 ( .A1(u5_mult_79_n1820), .A2(u5_mult_79_n1740), 
        .ZN(u5_mult_79_ab_8__4_) );
  NOR2_X4 u5_mult_79_U3014 ( .A1(u5_mult_79_n1811), .A2(u5_mult_79_n1740), 
        .ZN(u5_mult_79_ab_8__7_) );
  NOR2_X4 u5_mult_79_U3013 ( .A1(u5_mult_79_n1808), .A2(u5_mult_79_n1740), 
        .ZN(u5_mult_79_ab_8__8_) );
  NOR2_X4 u5_mult_79_U3012 ( .A1(u5_mult_79_n1796), .A2(u5_mult_79_n1741), 
        .ZN(u5_mult_79_ab_8__15_) );
  NOR2_X4 u5_mult_79_U3011 ( .A1(u5_mult_79_n1793), .A2(u5_mult_79_n1741), 
        .ZN(u5_mult_79_ab_8__16_) );
  NOR2_X4 u5_mult_79_U3010 ( .A1(u5_mult_79_n1790), .A2(u5_mult_79_n1741), 
        .ZN(u5_mult_79_ab_8__17_) );
  NOR2_X4 u5_mult_79_U3009 ( .A1(u5_mult_79_n1787), .A2(u5_mult_79_n1741), 
        .ZN(u5_mult_79_ab_8__18_) );
  INV_X4 u5_mult_79_U3008 ( .A(fracta_mul[8]), .ZN(u5_mult_79_n1844) );
  NOR2_X4 u5_mult_79_U3007 ( .A1(u5_mult_79_n1825), .A2(u5_mult_79_n1737), 
        .ZN(u5_mult_79_ab_7__2_) );
  NOR2_X4 u5_mult_79_U3006 ( .A1(u5_mult_79_n1823), .A2(u5_mult_79_n1737), 
        .ZN(u5_mult_79_ab_7__3_) );
  NOR2_X4 u5_mult_79_U3005 ( .A1(u5_mult_79_n1820), .A2(u5_mult_79_n1737), 
        .ZN(u5_mult_79_ab_7__4_) );
  NOR2_X4 u5_mult_79_U3004 ( .A1(u5_mult_79_n1817), .A2(u5_mult_79_n1737), 
        .ZN(u5_mult_79_ab_7__5_) );
  NOR2_X4 u5_mult_79_U3003 ( .A1(u5_mult_79_n1808), .A2(u5_mult_79_n1737), 
        .ZN(u5_mult_79_ab_7__8_) );
  NOR2_X4 u5_mult_79_U3002 ( .A1(u5_mult_79_n1802), .A2(u5_mult_79_n1737), 
        .ZN(u5_mult_79_ab_7__10_) );
  NOR2_X4 u5_mult_79_U3001 ( .A1(u5_mult_79_n1800), .A2(u5_mult_79_n1738), 
        .ZN(u5_mult_79_ab_7__11_) );
  NOR2_X4 u5_mult_79_U3000 ( .A1(u5_mult_79_n1868), .A2(u5_mult_79_n1738), 
        .ZN(u5_mult_79_ab_7__13_) );
  NOR2_X4 u5_mult_79_U2999 ( .A1(u5_mult_79_n1793), .A2(u5_mult_79_n1738), 
        .ZN(u5_mult_79_ab_7__16_) );
  NOR2_X4 u5_mult_79_U2998 ( .A1(u5_mult_79_n1790), .A2(u5_mult_79_n1738), 
        .ZN(u5_mult_79_ab_7__17_) );
  NOR2_X4 u5_mult_79_U2997 ( .A1(u5_mult_79_n1787), .A2(u5_mult_79_n1738), 
        .ZN(u5_mult_79_ab_7__18_) );
  NOR2_X4 u5_mult_79_U2996 ( .A1(u5_mult_79_n1338), .A2(u5_mult_79_n1738), 
        .ZN(u5_mult_79_ab_7__20_) );
  INV_X4 u5_mult_79_U2995 ( .A(fracta_mul[7]), .ZN(u5_mult_79_n1843) );
  NOR2_X4 u5_mult_79_U2994 ( .A1(u5_mult_79_n1825), .A2(u5_mult_79_n1734), 
        .ZN(u5_mult_79_ab_6__2_) );
  NOR2_X4 u5_mult_79_U2993 ( .A1(u5_mult_79_n1823), .A2(u5_mult_79_n1734), 
        .ZN(u5_mult_79_ab_6__3_) );
  NOR2_X4 u5_mult_79_U2992 ( .A1(u5_mult_79_n1820), .A2(u5_mult_79_n1734), 
        .ZN(u5_mult_79_ab_6__4_) );
  NOR2_X4 u5_mult_79_U2991 ( .A1(u5_mult_79_n1814), .A2(u5_mult_79_n1734), 
        .ZN(u5_mult_79_ab_6__6_) );
  NOR2_X4 u5_mult_79_U2990 ( .A1(u5_mult_79_n1808), .A2(u5_mult_79_n1734), 
        .ZN(u5_mult_79_ab_6__8_) );
  NOR2_X4 u5_mult_79_U2989 ( .A1(u5_mult_79_n1805), .A2(u5_mult_79_n1734), 
        .ZN(u5_mult_79_ab_6__9_) );
  NOR2_X4 u5_mult_79_U2988 ( .A1(u5_mult_79_n1802), .A2(u5_mult_79_n1734), 
        .ZN(u5_mult_79_ab_6__10_) );
  NOR2_X4 u5_mult_79_U2987 ( .A1(u5_mult_79_n1800), .A2(u5_mult_79_n1735), 
        .ZN(u5_mult_79_ab_6__11_) );
  NOR2_X4 u5_mult_79_U2986 ( .A1(u5_mult_79_n1798), .A2(u5_mult_79_n1735), 
        .ZN(u5_mult_79_ab_6__12_) );
  NOR2_X4 u5_mult_79_U2985 ( .A1(u5_mult_79_n1796), .A2(u5_mult_79_n1735), 
        .ZN(u5_mult_79_ab_6__15_) );
  NOR2_X4 u5_mult_79_U2984 ( .A1(u5_mult_79_n1793), .A2(u5_mult_79_n1735), 
        .ZN(u5_mult_79_ab_6__16_) );
  NOR2_X4 u5_mult_79_U2983 ( .A1(u5_mult_79_n1790), .A2(u5_mult_79_n1735), 
        .ZN(u5_mult_79_ab_6__17_) );
  NOR2_X4 u5_mult_79_U2982 ( .A1(u5_mult_79_n1787), .A2(u5_mult_79_n1735), 
        .ZN(u5_mult_79_ab_6__18_) );
  INV_X4 u5_mult_79_U2981 ( .A(fracta_mul[6]), .ZN(u5_mult_79_n1842) );
  NOR2_X4 u5_mult_79_U2980 ( .A1(u5_mult_79_n1825), .A2(u5_mult_79_n1731), 
        .ZN(u5_mult_79_ab_5__2_) );
  NOR2_X4 u5_mult_79_U2979 ( .A1(u5_mult_79_n1811), .A2(u5_mult_79_n1731), 
        .ZN(u5_mult_79_ab_5__7_) );
  NOR2_X4 u5_mult_79_U2978 ( .A1(u5_mult_79_n1802), .A2(u5_mult_79_n1731), 
        .ZN(u5_mult_79_ab_5__10_) );
  NOR2_X4 u5_mult_79_U2977 ( .A1(u5_mult_79_n1800), .A2(u5_mult_79_n1732), 
        .ZN(u5_mult_79_ab_5__11_) );
  NOR2_X4 u5_mult_79_U2976 ( .A1(u5_mult_79_n1798), .A2(u5_mult_79_n1732), 
        .ZN(u5_mult_79_ab_5__12_) );
  NOR2_X4 u5_mult_79_U2975 ( .A1(u5_mult_79_n1868), .A2(u5_mult_79_n1732), 
        .ZN(u5_mult_79_ab_5__13_) );
  NOR2_X4 u5_mult_79_U2974 ( .A1(u5_mult_79_n1793), .A2(u5_mult_79_n1732), 
        .ZN(u5_mult_79_ab_5__16_) );
  NOR2_X4 u5_mult_79_U2973 ( .A1(u5_mult_79_n1790), .A2(u5_mult_79_n1732), 
        .ZN(u5_mult_79_ab_5__17_) );
  NOR2_X4 u5_mult_79_U2972 ( .A1(u5_mult_79_n1787), .A2(u5_mult_79_n1732), 
        .ZN(u5_mult_79_ab_5__18_) );
  INV_X4 u5_mult_79_U2971 ( .A(fracta_mul[5]), .ZN(u5_mult_79_n1841) );
  NOR2_X4 u5_mult_79_U2970 ( .A1(u5_mult_79_n1811), .A2(u5_mult_79_n1728), 
        .ZN(u5_mult_79_ab_4__7_) );
  NOR2_X4 u5_mult_79_U2969 ( .A1(u5_mult_79_n1800), .A2(u5_mult_79_n1729), 
        .ZN(u5_mult_79_ab_4__11_) );
  NOR2_X4 u5_mult_79_U2968 ( .A1(u5_mult_79_n1868), .A2(u5_mult_79_n1729), 
        .ZN(u5_mult_79_ab_4__13_) );
  NOR2_X4 u5_mult_79_U2967 ( .A1(u5_mult_79_n1867), .A2(u5_mult_79_n1729), 
        .ZN(u5_mult_79_ab_4__14_) );
  NOR2_X4 u5_mult_79_U2966 ( .A1(u5_mult_79_n1796), .A2(u5_mult_79_n1729), 
        .ZN(u5_mult_79_ab_4__15_) );
  NOR2_X4 u5_mult_79_U2965 ( .A1(u5_mult_79_n1790), .A2(u5_mult_79_n1729), 
        .ZN(u5_mult_79_ab_4__17_) );
  INV_X4 u5_mult_79_U2964 ( .A(fracta_mul[4]), .ZN(u5_mult_79_n1840) );
  NOR2_X4 u5_mult_79_U2963 ( .A1(u5_mult_79_n1808), .A2(u5_mult_79_n1725), 
        .ZN(u5_mult_79_ab_3__8_) );
  NOR2_X4 u5_mult_79_U2962 ( .A1(u5_mult_79_n1805), .A2(u5_mult_79_n1725), 
        .ZN(u5_mult_79_ab_3__9_) );
  NOR2_X4 u5_mult_79_U2961 ( .A1(u5_mult_79_n1802), .A2(u5_mult_79_n1725), 
        .ZN(u5_mult_79_ab_3__10_) );
  NOR2_X4 u5_mult_79_U2960 ( .A1(u5_mult_79_n1800), .A2(u5_mult_79_n1726), 
        .ZN(u5_mult_79_ab_3__11_) );
  NOR2_X4 u5_mult_79_U2959 ( .A1(u5_mult_79_n1798), .A2(u5_mult_79_n1726), 
        .ZN(u5_mult_79_ab_3__12_) );
  NOR2_X4 u5_mult_79_U2958 ( .A1(u5_mult_79_n1868), .A2(u5_mult_79_n1726), 
        .ZN(u5_mult_79_ab_3__13_) );
  NOR2_X4 u5_mult_79_U2957 ( .A1(u5_mult_79_n1796), .A2(u5_mult_79_n1726), 
        .ZN(u5_mult_79_ab_3__15_) );
  NOR2_X4 u5_mult_79_U2956 ( .A1(u5_mult_79_n1793), .A2(u5_mult_79_n1726), 
        .ZN(u5_mult_79_ab_3__16_) );
  NOR2_X4 u5_mult_79_U2955 ( .A1(u5_mult_79_n1790), .A2(u5_mult_79_n1726), 
        .ZN(u5_mult_79_ab_3__17_) );
  NOR2_X4 u5_mult_79_U2954 ( .A1(u5_mult_79_n1787), .A2(u5_mult_79_n1726), 
        .ZN(u5_mult_79_ab_3__18_) );
  NOR2_X4 u5_mult_79_U2953 ( .A1(u5_mult_79_n1338), .A2(u5_mult_79_n1726), 
        .ZN(u5_mult_79_ab_3__20_) );
  NOR2_X4 u5_mult_79_U2952 ( .A1(u5_mult_79_n1798), .A2(u5_mult_79_n1723), 
        .ZN(u5_mult_79_ab_2__12_) );
  NOR2_X4 u5_mult_79_U2951 ( .A1(u5_mult_79_n1796), .A2(u5_mult_79_n1723), 
        .ZN(u5_mult_79_ab_2__15_) );
  NOR2_X4 u5_mult_79_U2950 ( .A1(u5_mult_79_n1831), .A2(u5_mult_79_n1719), 
        .ZN(u5_mult_79_ab_1__23_) );
  NOR2_X4 u5_mult_79_U2949 ( .A1(u5_mult_79_n1835), .A2(u5_mult_79_n46), .ZN(
        u5_mult_79_ab_1__0_) );
  INV_X4 u5_mult_79_U2948 ( .A(u6_N0), .ZN(u5_mult_79_n1881) );
  INV_X4 u5_mult_79_U2947 ( .A(u6_N1), .ZN(u5_mult_79_n1878) );
  NOR2_X4 u5_mult_79_U2946 ( .A1(u5_mult_79_n1882), .A2(u5_mult_79_n1825), 
        .ZN(u5_mult_79_ab_0__2_) );
  NOR2_X4 u5_mult_79_U2945 ( .A1(u5_mult_79_n1825), .A2(u5_mult_79_n46), .ZN(
        u5_mult_79_ab_1__2_) );
  INV_X4 u5_mult_79_U2944 ( .A(u6_N2), .ZN(u5_mult_79_n1877) );
  INV_X4 u5_mult_79_U2943 ( .A(u6_N3), .ZN(u5_mult_79_n1876) );
  NOR2_X4 u5_mult_79_U2942 ( .A1(u5_mult_79_n1882), .A2(u5_mult_79_n1820), 
        .ZN(u5_mult_79_ab_0__4_) );
  NOR2_X4 u5_mult_79_U2941 ( .A1(u5_mult_79_n1820), .A2(u5_mult_79_n1719), 
        .ZN(u5_mult_79_ab_1__4_) );
  INV_X4 u5_mult_79_U2940 ( .A(u6_N4), .ZN(u5_mult_79_n1875) );
  NOR2_X4 u5_mult_79_U2939 ( .A1(u5_mult_79_n1882), .A2(u5_mult_79_n1817), 
        .ZN(u5_mult_79_ab_0__5_) );
  NOR2_X4 u5_mult_79_U2938 ( .A1(u5_mult_79_n1817), .A2(u5_mult_79_n1719), 
        .ZN(u5_mult_79_ab_1__5_) );
  NOR2_X4 u5_mult_79_U2937 ( .A1(u5_mult_79_n1882), .A2(u5_mult_79_n1814), 
        .ZN(u5_mult_79_ab_0__6_) );
  NOR2_X4 u5_mult_79_U2936 ( .A1(u5_mult_79_n1814), .A2(u5_mult_79_n1720), 
        .ZN(u5_mult_79_ab_1__6_) );
  NOR2_X4 u5_mult_79_U2935 ( .A1(u5_mult_79_n1882), .A2(u5_mult_79_n1811), 
        .ZN(u5_mult_79_ab_0__7_) );
  NOR2_X4 u5_mult_79_U2934 ( .A1(u5_mult_79_n1882), .A2(u5_mult_79_n1808), 
        .ZN(u5_mult_79_ab_0__8_) );
  NOR2_X4 u5_mult_79_U2933 ( .A1(u5_mult_79_n1808), .A2(u5_mult_79_n1719), 
        .ZN(u5_mult_79_ab_1__8_) );
  NOR2_X4 u5_mult_79_U2932 ( .A1(u5_mult_79_n1882), .A2(u5_mult_79_n1805), 
        .ZN(u5_mult_79_ab_0__9_) );
  NOR2_X4 u5_mult_79_U2931 ( .A1(u5_mult_79_n1805), .A2(u5_mult_79_n1719), 
        .ZN(u5_mult_79_ab_1__9_) );
  NOR2_X4 u5_mult_79_U2930 ( .A1(u5_mult_79_n1882), .A2(u5_mult_79_n1802), 
        .ZN(u5_mult_79_ab_0__10_) );
  NOR2_X4 u5_mult_79_U2929 ( .A1(u5_mult_79_n1802), .A2(u5_mult_79_n1720), 
        .ZN(u5_mult_79_ab_1__10_) );
  NOR2_X4 u5_mult_79_U2928 ( .A1(u5_mult_79_n1882), .A2(u5_mult_79_n1800), 
        .ZN(u5_mult_79_ab_0__11_) );
  NOR2_X4 u5_mult_79_U2927 ( .A1(u5_mult_79_n1800), .A2(u5_mult_79_n1719), 
        .ZN(u5_mult_79_ab_1__11_) );
  NOR2_X4 u5_mult_79_U2926 ( .A1(u5_mult_79_n1882), .A2(u5_mult_79_n1798), 
        .ZN(u5_mult_79_ab_0__12_) );
  NOR2_X4 u5_mult_79_U2925 ( .A1(u5_mult_79_n1798), .A2(u5_mult_79_n1720), 
        .ZN(u5_mult_79_ab_1__12_) );
  NOR2_X4 u5_mult_79_U2924 ( .A1(u5_mult_79_n1882), .A2(u5_mult_79_n1868), 
        .ZN(u5_mult_79_ab_0__13_) );
  NOR2_X4 u5_mult_79_U2923 ( .A1(u5_mult_79_n1868), .A2(u5_mult_79_n1720), 
        .ZN(u5_mult_79_ab_1__13_) );
  NOR2_X4 u5_mult_79_U2922 ( .A1(u5_mult_79_n1882), .A2(u5_mult_79_n1866), 
        .ZN(u5_mult_79_ab_0__15_) );
  NOR2_X4 u5_mult_79_U2921 ( .A1(u5_mult_79_n1866), .A2(u5_mult_79_n1719), 
        .ZN(u5_mult_79_ab_1__15_) );
  NOR2_X4 u5_mult_79_U2920 ( .A1(u5_mult_79_n1882), .A2(u5_mult_79_n1793), 
        .ZN(u5_mult_79_ab_0__16_) );
  NOR2_X4 u5_mult_79_U2919 ( .A1(u5_mult_79_n1790), .A2(u5_mult_79_n1720), 
        .ZN(u5_mult_79_ab_1__17_) );
  NOR2_X4 u5_mult_79_U2918 ( .A1(u5_mult_79_n1882), .A2(u5_mult_79_n1787), 
        .ZN(u5_mult_79_ab_0__18_) );
  NOR2_X4 u5_mult_79_U2917 ( .A1(u5_mult_79_n1787), .A2(u5_mult_79_n1720), 
        .ZN(u5_mult_79_ab_1__18_) );
  NOR2_X4 u5_mult_79_U2916 ( .A1(u5_mult_79_n1861), .A2(u5_mult_79_n1719), 
        .ZN(u5_mult_79_ab_1__20_) );
  NOR2_X4 u5_mult_79_U2915 ( .A1(u5_mult_79_n1882), .A2(u5_mult_79_n1780), 
        .ZN(u5_mult_79_ab_0__22_) );
  NOR2_X4 u5_mult_79_U2914 ( .A1(u5_mult_79_n1781), .A2(u5_mult_79_n1719), 
        .ZN(u5_mult_79_ab_1__22_) );
  INV_X32 u5_mult_79_U2913 ( .A(u5_mult_79_n1836), .ZN(u5_mult_79_n1835) );
  INV_X32 u5_mult_79_U2912 ( .A(u5_mult_79_n1836), .ZN(u5_mult_79_n1834) );
  INV_X32 u5_mult_79_U2911 ( .A(u5_mult_79_n1877), .ZN(u5_mult_79_n1827) );
  INV_X32 u5_mult_79_U2910 ( .A(u5_mult_79_n1827), .ZN(u5_mult_79_n1826) );
  INV_X32 u5_mult_79_U2909 ( .A(u5_mult_79_n1827), .ZN(u5_mult_79_n1825) );
  INV_X32 u5_mult_79_U2908 ( .A(u5_mult_79_n1875), .ZN(u5_mult_79_n1822) );
  INV_X32 u5_mult_79_U2907 ( .A(u5_mult_79_n1822), .ZN(u5_mult_79_n1821) );
  INV_X32 u5_mult_79_U2906 ( .A(u5_mult_79_n1822), .ZN(u5_mult_79_n1820) );
  INV_X32 u5_mult_79_U2905 ( .A(u5_mult_79_n1874), .ZN(u5_mult_79_n1819) );
  INV_X32 u5_mult_79_U2904 ( .A(u5_mult_79_n1819), .ZN(u5_mult_79_n1818) );
  INV_X32 u5_mult_79_U2903 ( .A(u5_mult_79_n1819), .ZN(u5_mult_79_n1817) );
  INV_X32 u5_mult_79_U2902 ( .A(u5_mult_79_n1816), .ZN(u5_mult_79_n1815) );
  INV_X32 u5_mult_79_U2901 ( .A(u5_mult_79_n1816), .ZN(u5_mult_79_n1814) );
  INV_X32 u5_mult_79_U2900 ( .A(u5_mult_79_n1813), .ZN(u5_mult_79_n1811) );
  INV_X32 u5_mult_79_U2899 ( .A(u5_mult_79_n1810), .ZN(u5_mult_79_n1809) );
  INV_X32 u5_mult_79_U2898 ( .A(u5_mult_79_n1810), .ZN(u5_mult_79_n1808) );
  INV_X32 u5_mult_79_U2897 ( .A(u5_mult_79_n1870), .ZN(u5_mult_79_n1807) );
  INV_X32 u5_mult_79_U2896 ( .A(u5_mult_79_n1807), .ZN(u5_mult_79_n1806) );
  INV_X32 u5_mult_79_U2895 ( .A(u5_mult_79_n1807), .ZN(u5_mult_79_n1805) );
  INV_X32 u5_mult_79_U2894 ( .A(u5_mult_79_n1804), .ZN(u5_mult_79_n1803) );
  INV_X32 u5_mult_79_U2893 ( .A(u5_mult_79_n1804), .ZN(u5_mult_79_n1802) );
  INV_X32 u5_mult_79_U2892 ( .A(n2982), .ZN(u5_mult_79_n1800) );
  INV_X32 u5_mult_79_U2891 ( .A(u5_mult_79_n1797), .ZN(u5_mult_79_n1796) );
  INV_X32 u5_mult_79_U2890 ( .A(u5_mult_79_n1795), .ZN(u5_mult_79_n1794) );
  INV_X32 u5_mult_79_U2889 ( .A(u5_mult_79_n1795), .ZN(u5_mult_79_n1793) );
  INV_X32 u5_mult_79_U2888 ( .A(u5_mult_79_n1792), .ZN(u5_mult_79_n1791) );
  INV_X32 u5_mult_79_U2887 ( .A(u5_mult_79_n1792), .ZN(u5_mult_79_n1790) );
  INV_X32 u5_mult_79_U2886 ( .A(u5_mult_79_n1789), .ZN(u5_mult_79_n1787) );
  INV_X32 u5_mult_79_U2885 ( .A(u5_mult_79_n1782), .ZN(u5_mult_79_n1781) );
  INV_X32 u5_mult_79_U2884 ( .A(u5_mult_79_n1782), .ZN(u5_mult_79_n1780) );
  INV_X32 u5_mult_79_U2883 ( .A(u5_mult_79_n1772), .ZN(u5_mult_79_n1770) );
  INV_X32 u5_mult_79_U2882 ( .A(u5_mult_79_n1769), .ZN(u5_mult_79_n1767) );
  INV_X32 u5_mult_79_U2881 ( .A(u5_mult_79_n1766), .ZN(u5_mult_79_n1765) );
  INV_X32 u5_mult_79_U2880 ( .A(u5_mult_79_n1766), .ZN(u5_mult_79_n1764) );
  INV_X32 u5_mult_79_U2879 ( .A(u5_mult_79_n1851), .ZN(u5_mult_79_n1763) );
  INV_X32 u5_mult_79_U2878 ( .A(u5_mult_79_n1763), .ZN(u5_mult_79_n1762) );
  INV_X32 u5_mult_79_U2877 ( .A(u5_mult_79_n1763), .ZN(u5_mult_79_n1761) );
  INV_X32 u5_mult_79_U2876 ( .A(u5_mult_79_n1757), .ZN(u5_mult_79_n1756) );
  INV_X32 u5_mult_79_U2875 ( .A(u5_mult_79_n1757), .ZN(u5_mult_79_n1755) );
  INV_X32 u5_mult_79_U2874 ( .A(u5_mult_79_n1754), .ZN(u5_mult_79_n1752) );
  INV_X32 u5_mult_79_U2873 ( .A(u5_mult_79_n1751), .ZN(u5_mult_79_n1749) );
  INV_X32 u5_mult_79_U2872 ( .A(u5_mult_79_n1748), .ZN(u5_mult_79_n1747) );
  INV_X32 u5_mult_79_U2871 ( .A(u5_mult_79_n1748), .ZN(u5_mult_79_n1746) );
  INV_X32 u5_mult_79_U2870 ( .A(u5_mult_79_n1845), .ZN(u5_mult_79_n1745) );
  INV_X32 u5_mult_79_U2869 ( .A(u5_mult_79_n1745), .ZN(u5_mult_79_n1744) );
  INV_X32 u5_mult_79_U2868 ( .A(u5_mult_79_n1745), .ZN(u5_mult_79_n1743) );
  INV_X32 u5_mult_79_U2867 ( .A(u5_mult_79_n1742), .ZN(u5_mult_79_n1741) );
  INV_X32 u5_mult_79_U2866 ( .A(u5_mult_79_n1742), .ZN(u5_mult_79_n1740) );
  INV_X32 u5_mult_79_U2865 ( .A(u5_mult_79_n1739), .ZN(u5_mult_79_n1738) );
  INV_X32 u5_mult_79_U2864 ( .A(u5_mult_79_n1739), .ZN(u5_mult_79_n1737) );
  INV_X32 u5_mult_79_U2863 ( .A(u5_mult_79_n1736), .ZN(u5_mult_79_n1735) );
  INV_X32 u5_mult_79_U2862 ( .A(u5_mult_79_n1736), .ZN(u5_mult_79_n1734) );
  INV_X32 u5_mult_79_U2861 ( .A(u5_mult_79_n1733), .ZN(u5_mult_79_n1732) );
  INV_X32 u5_mult_79_U2860 ( .A(u5_mult_79_n1733), .ZN(u5_mult_79_n1731) );
  INV_X32 u5_mult_79_U2859 ( .A(u5_mult_79_n1730), .ZN(u5_mult_79_n1729) );
  INV_X32 u5_mult_79_U2858 ( .A(u5_mult_79_n1730), .ZN(u5_mult_79_n1728) );
  INV_X32 u5_mult_79_U2857 ( .A(u5_mult_79_n1727), .ZN(u5_mult_79_n1726) );
  INV_X32 u5_mult_79_U2856 ( .A(u5_mult_79_n1727), .ZN(u5_mult_79_n1725) );
  INV_X32 u5_mult_79_U2855 ( .A(u5_mult_79_n1724), .ZN(u5_mult_79_n1723) );
  INV_X32 u5_mult_79_U2854 ( .A(u5_mult_79_n1724), .ZN(u5_mult_79_n1722) );
  INV_X32 u5_mult_79_U2853 ( .A(u5_mult_79_n1721), .ZN(u5_mult_79_n1720) );
  INV_X8 u5_mult_79_U2852 ( .A(n3050), .ZN(u5_mult_79_n1837) );
  INV_X16 u5_mult_79_U2851 ( .A(u5_mult_79_n1837), .ZN(u5_mult_79_n1721) );
  INV_X4 u5_mult_79_U2850 ( .A(u5_mult_79_n1717), .ZN(u5_mult_79_SUMB_1__22_)
         );
  XNOR2_X2 u5_mult_79_U2849 ( .A(u5_mult_79_n623), .B(u5_mult_79_ab_1__22_), 
        .ZN(u5_mult_79_n1717) );
  INV_X4 u5_mult_79_U2848 ( .A(u5_mult_79_n1716), .ZN(u5_mult_79_CARRYB_1__22_) );
  INV_X4 u5_mult_79_U2847 ( .A(u5_mult_79_n1715), .ZN(u5_mult_79_SUMB_1__21_)
         );
  XNOR2_X2 u5_mult_79_U2846 ( .A(u5_mult_79_ab_0__22_), .B(u5_mult_79_n1121), 
        .ZN(u5_mult_79_n1715) );
  INV_X4 u5_mult_79_U2845 ( .A(u5_mult_79_n1714), .ZN(u5_mult_79_CARRYB_1__21_) );
  INV_X4 u5_mult_79_U2844 ( .A(u5_mult_79_n1713), .ZN(u5_mult_79_SUMB_1__20_)
         );
  XNOR2_X2 u5_mult_79_U2843 ( .A(u5_mult_79_ab_1__20_), .B(
        u5_mult_79_ab_0__21_), .ZN(u5_mult_79_n1713) );
  INV_X4 u5_mult_79_U2842 ( .A(u5_mult_79_n1712), .ZN(u5_mult_79_CARRYB_1__20_) );
  NAND2_X2 u5_mult_79_U2841 ( .A1(u5_mult_79_ab_0__21_), .A2(
        u5_mult_79_ab_1__20_), .ZN(u5_mult_79_n1712) );
  INV_X4 u5_mult_79_U2840 ( .A(u5_mult_79_n1711), .ZN(u5_mult_79_SUMB_1__19_)
         );
  XNOR2_X2 u5_mult_79_U2839 ( .A(u5_mult_79_ab_1__19_), .B(
        u5_mult_79_ab_0__20_), .ZN(u5_mult_79_n1711) );
  INV_X4 u5_mult_79_U2838 ( .A(u5_mult_79_n1710), .ZN(u5_mult_79_CARRYB_1__19_) );
  INV_X4 u5_mult_79_U2837 ( .A(u5_mult_79_n1709), .ZN(u5_mult_79_SUMB_1__18_)
         );
  XNOR2_X2 u5_mult_79_U2836 ( .A(u5_mult_79_ab_1__18_), .B(
        u5_mult_79_ab_0__19_), .ZN(u5_mult_79_n1709) );
  INV_X4 u5_mult_79_U2835 ( .A(u5_mult_79_n1708), .ZN(u5_mult_79_CARRYB_1__18_) );
  XNOR2_X2 u5_mult_79_U2834 ( .A(u5_mult_79_ab_1__17_), .B(
        u5_mult_79_ab_0__18_), .ZN(u5_mult_79_n1707) );
  INV_X4 u5_mult_79_U2833 ( .A(u5_mult_79_n1706), .ZN(u5_mult_79_SUMB_1__16_)
         );
  XNOR2_X2 u5_mult_79_U2832 ( .A(u5_mult_79_ab_1__16_), .B(
        u5_mult_79_ab_0__17_), .ZN(u5_mult_79_n1706) );
  INV_X4 u5_mult_79_U2831 ( .A(u5_mult_79_n1705), .ZN(u5_mult_79_CARRYB_1__16_) );
  INV_X4 u5_mult_79_U2830 ( .A(u5_mult_79_n1704), .ZN(u5_mult_79_SUMB_1__15_)
         );
  XNOR2_X2 u5_mult_79_U2829 ( .A(u5_mult_79_ab_1__15_), .B(
        u5_mult_79_ab_0__16_), .ZN(u5_mult_79_n1704) );
  INV_X4 u5_mult_79_U2828 ( .A(u5_mult_79_n1703), .ZN(u5_mult_79_CARRYB_1__15_) );
  NAND2_X2 u5_mult_79_U2827 ( .A1(u5_mult_79_ab_0__16_), .A2(
        u5_mult_79_ab_1__15_), .ZN(u5_mult_79_n1703) );
  INV_X4 u5_mult_79_U2826 ( .A(u5_mult_79_n1702), .ZN(u5_mult_79_SUMB_1__14_)
         );
  XNOR2_X2 u5_mult_79_U2825 ( .A(u5_mult_79_ab_1__14_), .B(
        u5_mult_79_ab_0__15_), .ZN(u5_mult_79_n1702) );
  INV_X4 u5_mult_79_U2824 ( .A(u5_mult_79_n1701), .ZN(u5_mult_79_CARRYB_1__14_) );
  NAND2_X2 u5_mult_79_U2823 ( .A1(u5_mult_79_ab_0__15_), .A2(
        u5_mult_79_ab_1__14_), .ZN(u5_mult_79_n1701) );
  INV_X4 u5_mult_79_U2822 ( .A(u5_mult_79_n1700), .ZN(u5_mult_79_SUMB_1__13_)
         );
  XNOR2_X2 u5_mult_79_U2821 ( .A(u5_mult_79_ab_1__13_), .B(
        u5_mult_79_ab_0__14_), .ZN(u5_mult_79_n1700) );
  INV_X4 u5_mult_79_U2820 ( .A(u5_mult_79_n1699), .ZN(u5_mult_79_CARRYB_1__13_) );
  INV_X4 u5_mult_79_U2819 ( .A(u5_mult_79_n1698), .ZN(u5_mult_79_SUMB_1__12_)
         );
  XNOR2_X2 u5_mult_79_U2818 ( .A(u5_mult_79_ab_1__12_), .B(
        u5_mult_79_ab_0__13_), .ZN(u5_mult_79_n1698) );
  INV_X4 u5_mult_79_U2817 ( .A(u5_mult_79_n1697), .ZN(u5_mult_79_CARRYB_1__12_) );
  NAND2_X2 u5_mult_79_U2816 ( .A1(u5_mult_79_ab_0__13_), .A2(
        u5_mult_79_ab_1__12_), .ZN(u5_mult_79_n1697) );
  INV_X4 u5_mult_79_U2815 ( .A(u5_mult_79_n1696), .ZN(u5_mult_79_SUMB_1__11_)
         );
  XNOR2_X2 u5_mult_79_U2814 ( .A(u5_mult_79_ab_1__11_), .B(
        u5_mult_79_ab_0__12_), .ZN(u5_mult_79_n1696) );
  INV_X4 u5_mult_79_U2813 ( .A(u5_mult_79_n1695), .ZN(u5_mult_79_CARRYB_1__11_) );
  INV_X4 u5_mult_79_U2812 ( .A(u5_mult_79_n1694), .ZN(u5_mult_79_SUMB_1__10_)
         );
  XNOR2_X2 u5_mult_79_U2811 ( .A(u5_mult_79_ab_1__10_), .B(
        u5_mult_79_ab_0__11_), .ZN(u5_mult_79_n1694) );
  INV_X4 u5_mult_79_U2810 ( .A(u5_mult_79_n1693), .ZN(u5_mult_79_CARRYB_1__10_) );
  NAND2_X2 u5_mult_79_U2809 ( .A1(u5_mult_79_ab_0__11_), .A2(
        u5_mult_79_ab_1__10_), .ZN(u5_mult_79_n1693) );
  INV_X4 u5_mult_79_U2808 ( .A(u5_mult_79_n1692), .ZN(u5_mult_79_SUMB_1__9_)
         );
  XNOR2_X2 u5_mult_79_U2807 ( .A(u5_mult_79_ab_1__9_), .B(u5_mult_79_ab_0__10_), .ZN(u5_mult_79_n1692) );
  INV_X4 u5_mult_79_U2806 ( .A(u5_mult_79_n1691), .ZN(u5_mult_79_SUMB_1__8_)
         );
  XNOR2_X2 u5_mult_79_U2805 ( .A(u5_mult_79_ab_1__8_), .B(u5_mult_79_ab_0__9_), 
        .ZN(u5_mult_79_n1691) );
  INV_X4 u5_mult_79_U2804 ( .A(u5_mult_79_n1690), .ZN(u5_mult_79_CARRYB_1__8_)
         );
  NAND2_X2 u5_mult_79_U2803 ( .A1(u5_mult_79_ab_0__9_), .A2(
        u5_mult_79_ab_1__8_), .ZN(u5_mult_79_n1690) );
  INV_X4 u5_mult_79_U2802 ( .A(u5_mult_79_n1689), .ZN(u5_mult_79_SUMB_1__7_)
         );
  XNOR2_X2 u5_mult_79_U2801 ( .A(u5_mult_79_ab_1__7_), .B(u5_mult_79_ab_0__8_), 
        .ZN(u5_mult_79_n1689) );
  INV_X4 u5_mult_79_U2800 ( .A(u5_mult_79_n1688), .ZN(u5_mult_79_CARRYB_1__7_)
         );
  NAND2_X2 u5_mult_79_U2799 ( .A1(u5_mult_79_ab_0__8_), .A2(
        u5_mult_79_ab_1__7_), .ZN(u5_mult_79_n1688) );
  INV_X4 u5_mult_79_U2798 ( .A(u5_mult_79_n1687), .ZN(u5_mult_79_SUMB_1__6_)
         );
  XNOR2_X2 u5_mult_79_U2797 ( .A(u5_mult_79_ab_1__6_), .B(u5_mult_79_ab_0__7_), 
        .ZN(u5_mult_79_n1687) );
  INV_X4 u5_mult_79_U2796 ( .A(u5_mult_79_n1686), .ZN(u5_mult_79_CARRYB_1__6_)
         );
  NAND2_X2 u5_mult_79_U2795 ( .A1(u5_mult_79_ab_0__7_), .A2(
        u5_mult_79_ab_1__6_), .ZN(u5_mult_79_n1686) );
  INV_X4 u5_mult_79_U2794 ( .A(u5_mult_79_n1685), .ZN(u5_mult_79_SUMB_1__5_)
         );
  XNOR2_X2 u5_mult_79_U2793 ( .A(u5_mult_79_ab_1__5_), .B(u5_mult_79_ab_0__6_), 
        .ZN(u5_mult_79_n1685) );
  INV_X4 u5_mult_79_U2792 ( .A(u5_mult_79_n1684), .ZN(u5_mult_79_CARRYB_1__5_)
         );
  NAND2_X2 u5_mult_79_U2791 ( .A1(u5_mult_79_ab_0__6_), .A2(
        u5_mult_79_ab_1__5_), .ZN(u5_mult_79_n1684) );
  INV_X4 u5_mult_79_U2790 ( .A(u5_mult_79_n1683), .ZN(u5_mult_79_SUMB_1__4_)
         );
  XNOR2_X2 u5_mult_79_U2789 ( .A(u5_mult_79_ab_1__4_), .B(u5_mult_79_ab_0__5_), 
        .ZN(u5_mult_79_n1683) );
  INV_X4 u5_mult_79_U2788 ( .A(u5_mult_79_n1682), .ZN(u5_mult_79_CARRYB_1__4_)
         );
  NAND2_X2 u5_mult_79_U2787 ( .A1(u5_mult_79_ab_0__5_), .A2(
        u5_mult_79_ab_1__4_), .ZN(u5_mult_79_n1682) );
  INV_X4 u5_mult_79_U2786 ( .A(u5_mult_79_n1681), .ZN(u5_mult_79_SUMB_1__3_)
         );
  XNOR2_X2 u5_mult_79_U2785 ( .A(u5_mult_79_ab_1__3_), .B(u5_mult_79_ab_0__4_), 
        .ZN(u5_mult_79_n1681) );
  INV_X4 u5_mult_79_U2784 ( .A(u5_mult_79_n1680), .ZN(u5_mult_79_CARRYB_1__3_)
         );
  NAND2_X2 u5_mult_79_U2783 ( .A1(u5_mult_79_ab_0__4_), .A2(
        u5_mult_79_ab_1__3_), .ZN(u5_mult_79_n1680) );
  INV_X4 u5_mult_79_U2782 ( .A(u5_mult_79_n1679), .ZN(u5_mult_79_SUMB_1__2_)
         );
  XNOR2_X2 u5_mult_79_U2781 ( .A(u5_mult_79_ab_1__2_), .B(u5_mult_79_ab_0__3_), 
        .ZN(u5_mult_79_n1679) );
  INV_X4 u5_mult_79_U2780 ( .A(u5_mult_79_n1678), .ZN(u5_mult_79_CARRYB_1__2_)
         );
  NAND2_X2 u5_mult_79_U2779 ( .A1(u5_mult_79_ab_0__3_), .A2(
        u5_mult_79_ab_1__2_), .ZN(u5_mult_79_n1678) );
  INV_X4 u5_mult_79_U2778 ( .A(u5_mult_79_n1677), .ZN(u5_mult_79_SUMB_1__1_)
         );
  XNOR2_X2 u5_mult_79_U2777 ( .A(u5_mult_79_ab_1__1_), .B(u5_mult_79_ab_0__2_), 
        .ZN(u5_mult_79_n1677) );
  INV_X4 u5_mult_79_U2776 ( .A(u5_mult_79_n1676), .ZN(u5_mult_79_CARRYB_1__1_)
         );
  NAND2_X2 u5_mult_79_U2775 ( .A1(u5_mult_79_ab_0__2_), .A2(
        u5_mult_79_ab_1__1_), .ZN(u5_mult_79_n1676) );
  INV_X4 u5_mult_79_U2774 ( .A(u5_mult_79_n1675), .ZN(u5_mult_79_CARRYB_1__0_)
         );
  NAND2_X2 u5_mult_79_U2773 ( .A1(u5_mult_79_ab_0__1_), .A2(
        u5_mult_79_ab_1__0_), .ZN(u5_mult_79_n1675) );
  INV_X4 u5_mult_79_U2772 ( .A(u5_mult_79_n1674), .ZN(u5_mult_79_CLA_CARRY[45]) );
  NAND2_X2 u5_mult_79_U2771 ( .A1(u5_mult_79_SUMB_23__22_), .A2(
        u5_mult_79_CARRYB_23__21_), .ZN(u5_mult_79_n1674) );
  INV_X4 u5_mult_79_U2770 ( .A(u5_mult_79_n1673), .ZN(u5_mult_79_CLA_SUM[44])
         );
  XNOR2_X2 u5_mult_79_U2769 ( .A(u5_mult_79_CARRYB_23__20_), .B(
        u5_mult_79_SUMB_23__21_), .ZN(u5_mult_79_n1673) );
  INV_X4 u5_mult_79_U2768 ( .A(u5_mult_79_n1672), .ZN(u5_mult_79_CLA_CARRY[44]) );
  NAND2_X2 u5_mult_79_U2767 ( .A1(u5_mult_79_SUMB_23__21_), .A2(
        u5_mult_79_CARRYB_23__20_), .ZN(u5_mult_79_n1672) );
  INV_X4 u5_mult_79_U2766 ( .A(u5_mult_79_n1671), .ZN(u5_mult_79_CLA_SUM[43])
         );
  XNOR2_X2 u5_mult_79_U2765 ( .A(u5_mult_79_CARRYB_23__19_), .B(
        u5_mult_79_SUMB_23__20_), .ZN(u5_mult_79_n1671) );
  INV_X4 u5_mult_79_U2764 ( .A(u5_mult_79_n1670), .ZN(u5_mult_79_CLA_SUM[42])
         );
  XNOR2_X2 u5_mult_79_U2763 ( .A(u5_mult_79_CARRYB_23__18_), .B(
        u5_mult_79_SUMB_23__19_), .ZN(u5_mult_79_n1670) );
  INV_X4 u5_mult_79_U2762 ( .A(u5_mult_79_n1669), .ZN(u5_mult_79_CLA_SUM[41])
         );
  XNOR2_X2 u5_mult_79_U2761 ( .A(u5_mult_79_CARRYB_23__17_), .B(
        u5_mult_79_SUMB_23__18_), .ZN(u5_mult_79_n1669) );
  INV_X4 u5_mult_79_U2760 ( .A(u5_mult_79_n1668), .ZN(u5_mult_79_CLA_CARRY[41]) );
  NAND2_X2 u5_mult_79_U2759 ( .A1(u5_mult_79_SUMB_23__18_), .A2(
        u5_mult_79_CARRYB_23__17_), .ZN(u5_mult_79_n1668) );
  INV_X4 u5_mult_79_U2758 ( .A(u5_mult_79_n1667), .ZN(u5_mult_79_CLA_SUM[40])
         );
  XNOR2_X2 u5_mult_79_U2757 ( .A(u5_mult_79_CARRYB_23__16_), .B(
        u5_mult_79_SUMB_23__17_), .ZN(u5_mult_79_n1667) );
  XNOR2_X2 u5_mult_79_U2756 ( .A(u5_mult_79_SUMB_23__16_), .B(
        u5_mult_79_CARRYB_23__15_), .ZN(u5_mult_79_n1666) );
  INV_X4 u5_mult_79_U2755 ( .A(u5_mult_79_n1665), .ZN(u5_mult_79_CLA_SUM[38])
         );
  XNOR2_X2 u5_mult_79_U2754 ( .A(u5_mult_79_SUMB_23__15_), .B(
        u5_mult_79_CARRYB_23__14_), .ZN(u5_mult_79_n1665) );
  INV_X4 u5_mult_79_U2753 ( .A(u5_mult_79_n1664), .ZN(u5_mult_79_CLA_SUM[37])
         );
  XNOR2_X2 u5_mult_79_U2752 ( .A(u5_mult_79_SUMB_23__14_), .B(
        u5_mult_79_CARRYB_23__13_), .ZN(u5_mult_79_n1664) );
  INV_X4 u5_mult_79_U2751 ( .A(u5_mult_79_n1663), .ZN(u5_mult_79_CLA_CARRY[37]) );
  INV_X4 u5_mult_79_U2750 ( .A(u5_mult_79_n1662), .ZN(u5_mult_79_CLA_SUM[36])
         );
  XNOR2_X2 u5_mult_79_U2749 ( .A(u5_mult_79_CARRYB_23__12_), .B(
        u5_mult_79_SUMB_23__13_), .ZN(u5_mult_79_n1662) );
  INV_X4 u5_mult_79_U2748 ( .A(u5_mult_79_n1661), .ZN(u5_mult_79_CLA_CARRY[36]) );
  NAND2_X2 u5_mult_79_U2747 ( .A1(u5_mult_79_n393), .A2(
        u5_mult_79_CARRYB_23__12_), .ZN(u5_mult_79_n1661) );
  INV_X4 u5_mult_79_U2746 ( .A(u5_mult_79_n1660), .ZN(u5_mult_79_CLA_SUM[35])
         );
  XNOR2_X2 u5_mult_79_U2745 ( .A(u5_mult_79_CARRYB_23__11_), .B(
        u5_mult_79_SUMB_23__12_), .ZN(u5_mult_79_n1660) );
  XNOR2_X2 u5_mult_79_U2744 ( .A(u5_mult_79_SUMB_23__11_), .B(
        u5_mult_79_CARRYB_23__10_), .ZN(u5_mult_79_n1659) );
  INV_X4 u5_mult_79_U2743 ( .A(u5_mult_79_n1658), .ZN(u5_mult_79_CLA_CARRY[34]) );
  XNOR2_X2 u5_mult_79_U2742 ( .A(u5_mult_79_SUMB_23__10_), .B(
        u5_mult_79_CARRYB_23__9_), .ZN(u5_mult_79_n1657) );
  INV_X4 u5_mult_79_U2741 ( .A(u5_mult_79_n1656), .ZN(u5_mult_79_CLA_CARRY[33]) );
  INV_X4 u5_mult_79_U2740 ( .A(u5_mult_79_n1655), .ZN(u5_mult_79_CLA_SUM[32])
         );
  XNOR2_X2 u5_mult_79_U2739 ( .A(u5_mult_79_CARRYB_23__8_), .B(
        u5_mult_79_SUMB_23__9_), .ZN(u5_mult_79_n1655) );
  INV_X4 u5_mult_79_U2738 ( .A(u5_mult_79_n1653), .ZN(u5_mult_79_CLA_SUM[30])
         );
  XNOR2_X2 u5_mult_79_U2737 ( .A(u5_mult_79_SUMB_23__7_), .B(
        u5_mult_79_CARRYB_23__6_), .ZN(u5_mult_79_n1653) );
  INV_X4 u5_mult_79_U2736 ( .A(u5_mult_79_n1652), .ZN(u5_mult_79_CLA_SUM[29])
         );
  XNOR2_X2 u5_mult_79_U2735 ( .A(u5_mult_79_SUMB_23__6_), .B(
        u5_mult_79_CARRYB_23__5_), .ZN(u5_mult_79_n1652) );
  XNOR2_X2 u5_mult_79_U2734 ( .A(u5_mult_79_SUMB_23__5_), .B(
        u5_mult_79_CARRYB_23__4_), .ZN(u5_mult_79_n1651) );
  XNOR2_X2 u5_mult_79_U2733 ( .A(u5_mult_79_SUMB_23__4_), .B(
        u5_mult_79_CARRYB_23__3_), .ZN(u5_mult_79_n1650) );
  INV_X4 u5_mult_79_U2732 ( .A(u5_mult_79_n1649), .ZN(u5_mult_79_CLA_CARRY[27]) );
  INV_X4 u5_mult_79_U2731 ( .A(u5_mult_79_n1648), .ZN(u5_mult_79_CLA_CARRY[26]) );
  INV_X4 u5_mult_79_U2730 ( .A(u5_mult_79_n1647), .ZN(u5_mult_79_CLA_SUM[25])
         );
  INV_X32 u5_mult_79_U2729 ( .A(u5_mult_79_n1721), .ZN(u5_mult_79_n1719) );
  NOR2_X2 u5_mult_79_U2728 ( .A1(u5_mult_79_n1780), .A2(u5_mult_79_n1723), 
        .ZN(u5_mult_79_ab_2__22_) );
  NAND2_X1 u5_mult_79_U2727 ( .A1(u5_mult_79_ab_19__7_), .A2(
        u5_mult_79_CARRYB_18__7_), .ZN(u5_mult_79_n1642) );
  NAND2_X1 u5_mult_79_U2726 ( .A1(u5_mult_79_ab_18__8_), .A2(
        u5_mult_79_CARRYB_17__8_), .ZN(u5_mult_79_n1639) );
  NOR2_X1 u5_mult_79_U2725 ( .A1(u5_mult_79_n1823), .A2(u5_mult_79_n1778), 
        .ZN(u5_mult_79_ab_21__3_) );
  NOR2_X1 u5_mult_79_U2724 ( .A1(u5_mult_79_n1823), .A2(u5_mult_79_n1775), 
        .ZN(u5_mult_79_ab_20__3_) );
  NAND3_X2 u5_mult_79_U2723 ( .A1(u5_mult_79_n1632), .A2(u5_mult_79_n1633), 
        .A3(u5_mult_79_n1634), .ZN(u5_mult_79_CARRYB_20__3_) );
  NAND2_X2 u5_mult_79_U2722 ( .A1(u5_mult_79_ab_20__3_), .A2(
        u5_mult_79_SUMB_19__4_), .ZN(u5_mult_79_n1633) );
  NAND2_X1 u5_mult_79_U2721 ( .A1(u5_mult_79_CARRYB_3__19_), .A2(
        u5_mult_79_SUMB_3__20_), .ZN(u5_mult_79_n1631) );
  NAND2_X1 u5_mult_79_U2720 ( .A1(u5_mult_79_ab_4__19_), .A2(
        u5_mult_79_SUMB_3__20_), .ZN(u5_mult_79_n1630) );
  NAND2_X1 u5_mult_79_U2719 ( .A1(u5_mult_79_ab_4__19_), .A2(
        u5_mult_79_CARRYB_3__19_), .ZN(u5_mult_79_n1629) );
  NAND2_X2 u5_mult_79_U2718 ( .A1(u5_mult_79_ab_3__20_), .A2(
        u5_mult_79_SUMB_2__21_), .ZN(u5_mult_79_n1627) );
  XOR2_X2 u5_mult_79_U2717 ( .A(u5_mult_79_n1625), .B(u5_mult_79_n341), .Z(
        u5_mult_79_SUMB_3__20_) );
  NAND2_X2 u5_mult_79_U2716 ( .A1(u5_mult_79_CARRYB_1__21_), .A2(
        u5_mult_79_SUMB_1__22_), .ZN(u5_mult_79_n1622) );
  NOR2_X1 u5_mult_79_U2715 ( .A1(u5_mult_79_n1783), .A2(u5_mult_79_n1729), 
        .ZN(u5_mult_79_ab_4__21_) );
  NOR2_X1 u5_mult_79_U2714 ( .A1(u5_mult_79_n1806), .A2(u5_mult_79_n1764), 
        .ZN(u5_mult_79_ab_16__9_) );
  NAND3_X2 u5_mult_79_U2713 ( .A1(u5_mult_79_n1616), .A2(u5_mult_79_n1617), 
        .A3(u5_mult_79_n1618), .ZN(u5_mult_79_CARRYB_3__22_) );
  NAND2_X2 u5_mult_79_U2712 ( .A1(u5_mult_79_ab_2__23_), .A2(
        u5_mult_79_ab_3__22_), .ZN(u5_mult_79_n1618) );
  NAND2_X2 u5_mult_79_U2711 ( .A1(u5_mult_79_ab_17__8_), .A2(
        u5_mult_79_SUMB_16__9_), .ZN(u5_mult_79_n1611) );
  XOR2_X2 u5_mult_79_U2710 ( .A(u5_mult_79_n1609), .B(u5_mult_79_SUMB_16__9_), 
        .Z(u5_mult_79_SUMB_17__8_) );
  NAND3_X2 u5_mult_79_U2709 ( .A1(u5_mult_79_n1606), .A2(u5_mult_79_n1607), 
        .A3(u5_mult_79_n1608), .ZN(u5_mult_79_CARRYB_16__9_) );
  NAND2_X1 u5_mult_79_U2708 ( .A1(u5_mult_79_ab_16__9_), .A2(
        u5_mult_79_CARRYB_15__9_), .ZN(u5_mult_79_n1608) );
  NOR2_X2 u5_mult_79_U2707 ( .A1(u5_mult_79_n1783), .A2(u5_mult_79_n1726), 
        .ZN(u5_mult_79_ab_3__21_) );
  NAND2_X2 u5_mult_79_U2706 ( .A1(u5_mult_79_ab_18__7_), .A2(
        u5_mult_79_CARRYB_17__7_), .ZN(u5_mult_79_n1613) );
  NAND3_X2 u5_mult_79_U2705 ( .A1(u5_mult_79_n1597), .A2(u5_mult_79_n1598), 
        .A3(u5_mult_79_n1599), .ZN(u5_mult_79_CARRYB_19__5_) );
  NAND2_X2 u5_mult_79_U2704 ( .A1(u5_mult_79_ab_18__6_), .A2(
        u5_mult_79_SUMB_17__7_), .ZN(u5_mult_79_n1595) );
  NAND3_X4 u5_mult_79_U2703 ( .A1(u5_mult_79_n1591), .A2(u5_mult_79_n1592), 
        .A3(u5_mult_79_n1593), .ZN(u5_mult_79_CARRYB_17__7_) );
  NOR2_X1 u5_mult_79_U2702 ( .A1(u5_mult_79_n1821), .A2(u5_mult_79_n1773), 
        .ZN(u5_mult_79_ab_19__4_) );
  NOR2_X1 u5_mult_79_U2701 ( .A1(u5_mult_79_n1787), .A2(u5_mult_79_n1729), 
        .ZN(u5_mult_79_ab_4__18_) );
  NOR2_X1 u5_mult_79_U2700 ( .A1(u5_mult_79_n1815), .A2(u5_mult_79_n1764), 
        .ZN(u5_mult_79_ab_16__6_) );
  NAND3_X2 u5_mult_79_U2699 ( .A1(u5_mult_79_n1588), .A2(u5_mult_79_n1589), 
        .A3(u5_mult_79_n1590), .ZN(u5_mult_79_CARRYB_19__4_) );
  NAND3_X2 u5_mult_79_U2698 ( .A1(u5_mult_79_n1585), .A2(u5_mult_79_n1586), 
        .A3(u5_mult_79_n1587), .ZN(u5_mult_79_CARRYB_6__16_) );
  NAND2_X1 u5_mult_79_U2697 ( .A1(u5_mult_79_ab_6__16_), .A2(
        u5_mult_79_CARRYB_5__16_), .ZN(u5_mult_79_n1585) );
  NAND2_X2 u5_mult_79_U2696 ( .A1(u5_mult_79_CARRYB_4__17_), .A2(
        u5_mult_79_SUMB_4__18_), .ZN(u5_mult_79_n1584) );
  NAND2_X2 u5_mult_79_U2695 ( .A1(u5_mult_79_ab_5__17_), .A2(
        u5_mult_79_SUMB_4__18_), .ZN(u5_mult_79_n1583) );
  NAND2_X1 u5_mult_79_U2694 ( .A1(u5_mult_79_ab_5__17_), .A2(
        u5_mult_79_CARRYB_4__17_), .ZN(u5_mult_79_n1582) );
  NAND2_X1 u5_mult_79_U2693 ( .A1(u5_mult_79_ab_4__18_), .A2(
        u5_mult_79_CARRYB_3__18_), .ZN(u5_mult_79_n1581) );
  NOR2_X1 u5_mult_79_U2692 ( .A1(u5_mult_79_n1785), .A2(u5_mult_79_n1738), 
        .ZN(u5_mult_79_ab_7__19_) );
  NAND3_X2 u5_mult_79_U2691 ( .A1(u5_mult_79_n1572), .A2(u5_mult_79_n1573), 
        .A3(u5_mult_79_n1574), .ZN(u5_mult_79_CARRYB_7__19_) );
  NAND2_X1 u5_mult_79_U2690 ( .A1(u5_mult_79_ab_7__19_), .A2(
        u5_mult_79_CARRYB_6__19_), .ZN(u5_mult_79_n1573) );
  NAND2_X1 u5_mult_79_U2689 ( .A1(u5_mult_79_CARRYB_17__9_), .A2(
        u5_mult_79_SUMB_17__10_), .ZN(u5_mult_79_n1571) );
  NAND2_X1 u5_mult_79_U2688 ( .A1(u5_mult_79_ab_18__9_), .A2(
        u5_mult_79_CARRYB_17__9_), .ZN(u5_mult_79_n1569) );
  NAND2_X2 u5_mult_79_U2687 ( .A1(u5_mult_79_n350), .A2(
        u5_mult_79_SUMB_16__11_), .ZN(u5_mult_79_n1568) );
  NAND2_X2 u5_mult_79_U2686 ( .A1(u5_mult_79_SUMB_16__11_), .A2(
        u5_mult_79_ab_17__10_), .ZN(u5_mult_79_n1567) );
  NAND2_X1 u5_mult_79_U2685 ( .A1(u5_mult_79_ab_17__10_), .A2(
        u5_mult_79_CARRYB_16__10_), .ZN(u5_mult_79_n1566) );
  NAND3_X2 u5_mult_79_U2684 ( .A1(u5_mult_79_n1562), .A2(u5_mult_79_n1563), 
        .A3(u5_mult_79_n1564), .ZN(u5_mult_79_CARRYB_22__5_) );
  NAND2_X1 u5_mult_79_U2683 ( .A1(u5_mult_79_CARRYB_21__5_), .A2(
        u5_mult_79_SUMB_21__6_), .ZN(u5_mult_79_n1564) );
  NAND2_X1 u5_mult_79_U2682 ( .A1(u5_mult_79_ab_22__5_), .A2(
        u5_mult_79_SUMB_21__6_), .ZN(u5_mult_79_n1563) );
  NAND2_X1 u5_mult_79_U2681 ( .A1(u5_mult_79_ab_22__5_), .A2(
        u5_mult_79_CARRYB_21__5_), .ZN(u5_mult_79_n1562) );
  XOR2_X2 u5_mult_79_U2680 ( .A(u5_mult_79_n1558), .B(u5_mult_79_n381), .Z(
        u5_mult_79_SUMB_21__6_) );
  NAND2_X1 u5_mult_79_U2679 ( .A1(u5_mult_79_SUMB_23__4_), .A2(
        u5_mult_79_CARRYB_23__3_), .ZN(u5_mult_79_n1649) );
  NOR2_X1 u5_mult_79_U2678 ( .A1(u5_mult_79_n1867), .A2(u5_mult_79_n1759), 
        .ZN(u5_mult_79_ab_14__14_) );
  NOR2_X1 u5_mult_79_U2677 ( .A1(u5_mult_79_n1783), .A2(u5_mult_79_n1732), 
        .ZN(u5_mult_79_ab_5__21_) );
  NAND3_X2 u5_mult_79_U2676 ( .A1(u5_mult_79_n1556), .A2(u5_mult_79_n1555), 
        .A3(u5_mult_79_n1557), .ZN(u5_mult_79_CARRYB_14__14_) );
  NAND2_X1 u5_mult_79_U2675 ( .A1(u5_mult_79_ab_14__14_), .A2(
        u5_mult_79_CARRYB_13__14_), .ZN(u5_mult_79_n1557) );
  NAND2_X2 u5_mult_79_U2674 ( .A1(u5_mult_79_ab_14__14_), .A2(u5_mult_79_n472), 
        .ZN(u5_mult_79_n1556) );
  NAND2_X1 u5_mult_79_U2673 ( .A1(u5_mult_79_ab_17__11_), .A2(
        u5_mult_79_CARRYB_16__11_), .ZN(u5_mult_79_n1548) );
  NAND3_X4 u5_mult_79_U2672 ( .A1(u5_mult_79_n1546), .A2(u5_mult_79_n1545), 
        .A3(u5_mult_79_n1547), .ZN(u5_mult_79_CARRYB_16__12_) );
  NAND2_X2 u5_mult_79_U2671 ( .A1(u5_mult_79_n1134), .A2(
        u5_mult_79_CARRYB_15__12_), .ZN(u5_mult_79_n1547) );
  NAND2_X2 u5_mult_79_U2670 ( .A1(u5_mult_79_ab_16__12_), .A2(u5_mult_79_n1134), .ZN(u5_mult_79_n1546) );
  NAND2_X1 u5_mult_79_U2669 ( .A1(u5_mult_79_ab_16__12_), .A2(
        u5_mult_79_CARRYB_15__12_), .ZN(u5_mult_79_n1545) );
  XNOR2_X2 u5_mult_79_U2668 ( .A(u5_mult_79_CARRYB_3__19_), .B(
        u5_mult_79_ab_4__19_), .ZN(u5_mult_79_n1544) );
  XNOR2_X2 u5_mult_79_U2667 ( .A(u5_mult_79_n284), .B(u5_mult_79_ab_4__21_), 
        .ZN(u5_mult_79_n1543) );
  NOR2_X1 u5_mult_79_U2666 ( .A1(u5_mult_79_n1821), .A2(u5_mult_79_n1775), 
        .ZN(u5_mult_79_ab_20__4_) );
  NAND3_X2 u5_mult_79_U2665 ( .A1(u5_mult_79_n1540), .A2(u5_mult_79_n1541), 
        .A3(u5_mult_79_n1542), .ZN(u5_mult_79_CARRYB_20__4_) );
  NAND3_X2 u5_mult_79_U2664 ( .A1(u5_mult_79_n1537), .A2(u5_mult_79_n1538), 
        .A3(u5_mult_79_n1539), .ZN(u5_mult_79_CARRYB_6__15_) );
  NAND2_X2 u5_mult_79_U2663 ( .A1(u5_mult_79_CARRYB_4__16_), .A2(
        u5_mult_79_SUMB_4__17_), .ZN(u5_mult_79_n1536) );
  NAND2_X2 u5_mult_79_U2662 ( .A1(u5_mult_79_ab_5__16_), .A2(
        u5_mult_79_SUMB_4__17_), .ZN(u5_mult_79_n1535) );
  XOR2_X2 u5_mult_79_U2661 ( .A(u5_mult_79_n1533), .B(u5_mult_79_SUMB_4__17_), 
        .Z(u5_mult_79_SUMB_5__16_) );
  NAND3_X2 u5_mult_79_U2660 ( .A1(u5_mult_79_n1530), .A2(u5_mult_79_n1531), 
        .A3(u5_mult_79_n1532), .ZN(u5_mult_79_CARRYB_4__17_) );
  NAND2_X1 u5_mult_79_U2659 ( .A1(u5_mult_79_CARRYB_3__17_), .A2(
        u5_mult_79_SUMB_3__18_), .ZN(u5_mult_79_n1532) );
  NAND2_X1 u5_mult_79_U2658 ( .A1(u5_mult_79_ab_4__17_), .A2(
        u5_mult_79_SUMB_3__18_), .ZN(u5_mult_79_n1531) );
  NAND2_X1 u5_mult_79_U2657 ( .A1(u5_mult_79_ab_4__17_), .A2(
        u5_mult_79_CARRYB_3__17_), .ZN(u5_mult_79_n1530) );
  NAND2_X2 u5_mult_79_U2656 ( .A1(u5_mult_79_ab_3__18_), .A2(u5_mult_79_n423), 
        .ZN(u5_mult_79_n1528) );
  NAND2_X1 u5_mult_79_U2655 ( .A1(u5_mult_79_ab_3__18_), .A2(
        u5_mult_79_CARRYB_2__18_), .ZN(u5_mult_79_n1527) );
  NAND2_X2 u5_mult_79_U2654 ( .A1(u5_mult_79_CARRYB_16__7_), .A2(
        u5_mult_79_n354), .ZN(u5_mult_79_n1591) );
  XNOR2_X2 u5_mult_79_U2653 ( .A(u5_mult_79_CARRYB_13__14_), .B(
        u5_mult_79_n1526), .ZN(u5_mult_79_n1554) );
  INV_X8 u5_mult_79_U2652 ( .A(n3035), .ZN(u5_mult_79_n1863) );
  NOR2_X1 u5_mult_79_U2651 ( .A1(u5_mult_79_n1868), .A2(u5_mult_79_n1759), 
        .ZN(u5_mult_79_ab_14__13_) );
  CLKBUF_X2 u5_mult_79_U2650 ( .A(u5_mult_79_CARRYB_13__13_), .Z(
        u5_mult_79_n1524) );
  NAND3_X2 u5_mult_79_U2649 ( .A1(u5_mult_79_n1522), .A2(u5_mult_79_n1523), 
        .A3(u5_mult_79_n1521), .ZN(u5_mult_79_CARRYB_14__13_) );
  NAND2_X1 u5_mult_79_U2648 ( .A1(u5_mult_79_ab_18__11_), .A2(
        u5_mult_79_CARRYB_17__11_), .ZN(u5_mult_79_n1515) );
  NAND3_X4 u5_mult_79_U2647 ( .A1(u5_mult_79_n1613), .A2(u5_mult_79_n1614), 
        .A3(u5_mult_79_n1615), .ZN(u5_mult_79_CARRYB_18__7_) );
  NAND2_X2 u5_mult_79_U2646 ( .A1(u5_mult_79_ab_17__7_), .A2(
        u5_mult_79_CARRYB_16__7_), .ZN(u5_mult_79_n1593) );
  XNOR2_X2 u5_mult_79_U2645 ( .A(u5_mult_79_ab_18__7_), .B(
        u5_mult_79_CARRYB_17__7_), .ZN(u5_mult_79_n1513) );
  NAND3_X2 u5_mult_79_U2644 ( .A1(u5_mult_79_n1509), .A2(u5_mult_79_n1510), 
        .A3(u5_mult_79_n1511), .ZN(u5_mult_79_CARRYB_23__2_) );
  NAND2_X2 u5_mult_79_U2643 ( .A1(u5_mult_79_ab_23__2_), .A2(
        u5_mult_79_CARRYB_22__2_), .ZN(u5_mult_79_n1510) );
  NAND2_X1 u5_mult_79_U2642 ( .A1(u5_mult_79_ab_23__2_), .A2(
        u5_mult_79_SUMB_22__3_), .ZN(u5_mult_79_n1509) );
  NAND2_X2 u5_mult_79_U2641 ( .A1(u5_mult_79_ab_22__2_), .A2(u5_mult_79_n280), 
        .ZN(u5_mult_79_n1506) );
  NAND3_X2 u5_mult_79_U2640 ( .A1(u5_mult_79_n1501), .A2(u5_mult_79_n1502), 
        .A3(u5_mult_79_n1503), .ZN(u5_mult_79_CARRYB_16__4_) );
  NAND2_X2 u5_mult_79_U2639 ( .A1(u5_mult_79_n133), .A2(
        u5_mult_79_CARRYB_14__5_), .ZN(u5_mult_79_n1500) );
  NAND2_X1 u5_mult_79_U2638 ( .A1(u5_mult_79_ab_15__5_), .A2(
        u5_mult_79_CARRYB_14__5_), .ZN(u5_mult_79_n1498) );
  NAND3_X4 u5_mult_79_U2637 ( .A1(u5_mult_79_n1495), .A2(u5_mult_79_n1496), 
        .A3(u5_mult_79_n1497), .ZN(u5_mult_79_CARRYB_17__9_) );
  NAND2_X2 u5_mult_79_U2636 ( .A1(u5_mult_79_CARRYB_16__9_), .A2(
        u5_mult_79_SUMB_16__10_), .ZN(u5_mult_79_n1497) );
  NAND2_X2 u5_mult_79_U2635 ( .A1(u5_mult_79_ab_17__9_), .A2(
        u5_mult_79_SUMB_16__10_), .ZN(u5_mult_79_n1496) );
  NAND3_X2 u5_mult_79_U2634 ( .A1(u5_mult_79_n1492), .A2(u5_mult_79_n1493), 
        .A3(u5_mult_79_n1494), .ZN(u5_mult_79_CARRYB_16__10_) );
  NAND2_X1 u5_mult_79_U2633 ( .A1(u5_mult_79_CARRYB_15__10_), .A2(
        u5_mult_79_ab_16__10_), .ZN(u5_mult_79_n1492) );
  NAND2_X1 u5_mult_79_U2632 ( .A1(u5_mult_79_ab_15__11_), .A2(
        u5_mult_79_CARRYB_14__11_), .ZN(u5_mult_79_n1489) );
  NAND2_X1 u5_mult_79_U2631 ( .A1(u5_mult_79_ab_14__12_), .A2(
        u5_mult_79_CARRYB_13__12_), .ZN(u5_mult_79_n1486) );
  NOR2_X1 u5_mult_79_U2630 ( .A1(u5_mult_79_n1798), .A2(u5_mult_79_n1741), 
        .ZN(u5_mult_79_ab_8__12_) );
  NAND3_X2 u5_mult_79_U2629 ( .A1(u5_mult_79_n1485), .A2(u5_mult_79_n1484), 
        .A3(u5_mult_79_n1483), .ZN(u5_mult_79_CARRYB_8__12_) );
  NAND2_X2 u5_mult_79_U2628 ( .A1(u5_mult_79_ab_8__12_), .A2(
        u5_mult_79_SUMB_7__13_), .ZN(u5_mult_79_n1484) );
  NAND2_X1 u5_mult_79_U2627 ( .A1(u5_mult_79_ab_16__7_), .A2(
        u5_mult_79_CARRYB_15__7_), .ZN(u5_mult_79_n1480) );
  XNOR2_X2 u5_mult_79_U2626 ( .A(u5_mult_79_n1512), .B(u5_mult_79_n352), .ZN(
        u5_mult_79_SUMB_18__6_) );
  XNOR2_X2 u5_mult_79_U2625 ( .A(u5_mult_79_n1513), .B(u5_mult_79_n377), .ZN(
        u5_mult_79_SUMB_18__7_) );
  NAND2_X2 u5_mult_79_U2624 ( .A1(u5_mult_79_ab_20__4_), .A2(
        u5_mult_79_SUMB_19__5_), .ZN(u5_mult_79_n1541) );
  NOR2_X1 u5_mult_79_U2623 ( .A1(u5_mult_79_n1818), .A2(u5_mult_79_n1767), 
        .ZN(u5_mult_79_ab_17__5_) );
  NOR2_X1 u5_mult_79_U2622 ( .A1(u5_mult_79_n1818), .A2(u5_mult_79_n1764), 
        .ZN(u5_mult_79_ab_16__5_) );
  NAND2_X1 u5_mult_79_U2621 ( .A1(u5_mult_79_ab_17__5_), .A2(
        u5_mult_79_CARRYB_16__5_), .ZN(u5_mult_79_n1476) );
  NAND2_X2 u5_mult_79_U2620 ( .A1(u5_mult_79_ab_17__5_), .A2(
        u5_mult_79_SUMB_16__6_), .ZN(u5_mult_79_n1475) );
  NAND3_X2 u5_mult_79_U2619 ( .A1(u5_mult_79_n1471), .A2(u5_mult_79_n1472), 
        .A3(u5_mult_79_n1473), .ZN(u5_mult_79_CARRYB_16__5_) );
  NAND2_X1 u5_mult_79_U2618 ( .A1(u5_mult_79_ab_16__5_), .A2(
        u5_mult_79_CARRYB_15__5_), .ZN(u5_mult_79_n1473) );
  NAND2_X2 u5_mult_79_U2617 ( .A1(u5_mult_79_ab_16__5_), .A2(
        u5_mult_79_SUMB_15__6_), .ZN(u5_mult_79_n1472) );
  NAND2_X1 u5_mult_79_U2616 ( .A1(u5_mult_79_SUMB_15__6_), .A2(
        u5_mult_79_CARRYB_15__5_), .ZN(u5_mult_79_n1471) );
  NAND3_X2 u5_mult_79_U2615 ( .A1(u5_mult_79_n1470), .A2(u5_mult_79_n1469), 
        .A3(u5_mult_79_n1468), .ZN(u5_mult_79_CARRYB_13__8_) );
  NAND2_X1 u5_mult_79_U2614 ( .A1(u5_mult_79_ab_13__8_), .A2(
        u5_mult_79_CARRYB_12__8_), .ZN(u5_mult_79_n1468) );
  NAND2_X2 u5_mult_79_U2613 ( .A1(u5_mult_79_n103), .A2(
        u5_mult_79_SUMB_11__10_), .ZN(u5_mult_79_n1467) );
  NAND2_X2 u5_mult_79_U2612 ( .A1(u5_mult_79_ab_12__9_), .A2(
        u5_mult_79_SUMB_11__10_), .ZN(u5_mult_79_n1466) );
  NAND3_X2 u5_mult_79_U2611 ( .A1(u5_mult_79_n1462), .A2(u5_mult_79_n1463), 
        .A3(u5_mult_79_n1464), .ZN(u5_mult_79_CARRYB_11__10_) );
  NAND2_X1 u5_mult_79_U2610 ( .A1(u5_mult_79_ab_11__10_), .A2(
        u5_mult_79_CARRYB_10__10_), .ZN(u5_mult_79_n1462) );
  NAND3_X2 u5_mult_79_U2609 ( .A1(u5_mult_79_n1459), .A2(u5_mult_79_n1460), 
        .A3(u5_mult_79_n1461), .ZN(u5_mult_79_CARRYB_10__11_) );
  NAND2_X1 u5_mult_79_U2608 ( .A1(u5_mult_79_ab_10__11_), .A2(
        u5_mult_79_CARRYB_9__11_), .ZN(u5_mult_79_n1459) );
  NAND3_X2 u5_mult_79_U2607 ( .A1(u5_mult_79_n1455), .A2(u5_mult_79_n1456), 
        .A3(u5_mult_79_n1457), .ZN(u5_mult_79_CARRYB_23__9_) );
  NAND2_X1 u5_mult_79_U2606 ( .A1(u5_mult_79_CARRYB_22__9_), .A2(
        u5_mult_79_SUMB_22__10_), .ZN(u5_mult_79_n1457) );
  NAND2_X1 u5_mult_79_U2605 ( .A1(u5_mult_79_ab_23__9_), .A2(
        u5_mult_79_SUMB_22__10_), .ZN(u5_mult_79_n1456) );
  NAND2_X1 u5_mult_79_U2604 ( .A1(u5_mult_79_ab_23__9_), .A2(
        u5_mult_79_CARRYB_22__9_), .ZN(u5_mult_79_n1455) );
  XNOR2_X2 u5_mult_79_U2603 ( .A(u5_mult_79_n28), .B(u5_mult_79_ab_7__19_), 
        .ZN(u5_mult_79_n1451) );
  XNOR2_X2 u5_mult_79_U2602 ( .A(u5_mult_79_SUMB_23__3_), .B(u5_mult_79_n1450), 
        .ZN(u5_mult_79_n1449) );
  INV_X4 u5_mult_79_U2601 ( .A(u5_mult_79_CARRYB_23__2_), .ZN(u5_mult_79_n1450) );
  NAND2_X1 u5_mult_79_U2600 ( .A1(u5_mult_79_SUMB_23__3_), .A2(
        u5_mult_79_CARRYB_23__2_), .ZN(u5_mult_79_n1648) );
  NAND2_X2 u5_mult_79_U2599 ( .A1(u5_mult_79_CARRYB_16__8_), .A2(
        u5_mult_79_n127), .ZN(u5_mult_79_n1612) );
  NAND2_X2 u5_mult_79_U2598 ( .A1(u5_mult_79_ab_19__7_), .A2(
        u5_mult_79_SUMB_18__8_), .ZN(u5_mult_79_n1643) );
  NOR2_X1 u5_mult_79_U2597 ( .A1(u5_mult_79_n1831), .A2(u5_mult_79_n1737), 
        .ZN(u5_mult_79_ab_7__23_) );
  NOR2_X1 u5_mult_79_U2596 ( .A1(u5_mult_79_n1780), .A2(u5_mult_79_n1741), 
        .ZN(u5_mult_79_ab_8__22_) );
  NOR2_X1 u5_mult_79_U2595 ( .A1(u5_mult_79_n1801), .A2(u5_mult_79_n1773), 
        .ZN(u5_mult_79_ab_19__11_) );
  NOR2_X1 u5_mult_79_U2594 ( .A1(u5_mult_79_n1803), .A2(u5_mult_79_n1775), 
        .ZN(u5_mult_79_ab_20__10_) );
  NAND3_X2 u5_mult_79_U2593 ( .A1(u5_mult_79_n1446), .A2(u5_mult_79_n1447), 
        .A3(u5_mult_79_n1448), .ZN(u5_mult_79_CARRYB_8__22_) );
  NAND2_X2 u5_mult_79_U2592 ( .A1(u5_mult_79_ab_7__23_), .A2(
        u5_mult_79_ab_8__22_), .ZN(u5_mult_79_n1448) );
  NAND2_X2 u5_mult_79_U2591 ( .A1(u5_mult_79_ab_8__22_), .A2(
        u5_mult_79_CARRYB_7__22_), .ZN(u5_mult_79_n1446) );
  XOR2_X1 u5_mult_79_U2590 ( .A(u5_mult_79_CARRYB_7__22_), .B(u5_mult_79_n1445), .Z(u5_mult_79_SUMB_8__22_) );
  XOR2_X2 u5_mult_79_U2589 ( .A(u5_mult_79_ab_8__22_), .B(u5_mult_79_ab_7__23_), .Z(u5_mult_79_n1445) );
  NAND3_X2 u5_mult_79_U2588 ( .A1(u5_mult_79_n1442), .A2(u5_mult_79_n1443), 
        .A3(u5_mult_79_n1444), .ZN(u5_mult_79_CARRYB_19__11_) );
  NAND2_X1 u5_mult_79_U2587 ( .A1(u5_mult_79_ab_19__11_), .A2(
        u5_mult_79_CARRYB_18__11_), .ZN(u5_mult_79_n1444) );
  NAND2_X1 u5_mult_79_U2586 ( .A1(u5_mult_79_CARRYB_18__11_), .A2(
        u5_mult_79_SUMB_18__12_), .ZN(u5_mult_79_n1442) );
  NAND2_X2 u5_mult_79_U2585 ( .A1(u5_mult_79_ab_14__16_), .A2(u5_mult_79_n484), 
        .ZN(u5_mult_79_n1437) );
  NAND3_X2 u5_mult_79_U2584 ( .A1(u5_mult_79_n1433), .A2(u5_mult_79_n1434), 
        .A3(u5_mult_79_n1435), .ZN(u5_mult_79_CARRYB_22__8_) );
  NAND2_X1 u5_mult_79_U2583 ( .A1(u5_mult_79_ab_22__8_), .A2(
        u5_mult_79_CARRYB_21__8_), .ZN(u5_mult_79_n1433) );
  NAND3_X2 u5_mult_79_U2582 ( .A1(u5_mult_79_n1430), .A2(u5_mult_79_n1431), 
        .A3(u5_mult_79_n1432), .ZN(u5_mult_79_CARRYB_21__9_) );
  NAND2_X1 u5_mult_79_U2581 ( .A1(u5_mult_79_ab_20__10_), .A2(
        u5_mult_79_CARRYB_19__10_), .ZN(u5_mult_79_n1429) );
  NAND2_X1 u5_mult_79_U2580 ( .A1(u5_mult_79_ab_3__20_), .A2(u5_mult_79_n337), 
        .ZN(u5_mult_79_n1626) );
  XNOR2_X2 u5_mult_79_U2579 ( .A(u5_mult_79_CARRYB_13__13_), .B(
        u5_mult_79_ab_14__13_), .ZN(u5_mult_79_n1425) );
  NAND2_X2 u5_mult_79_U2578 ( .A1(u5_mult_79_ab_18__8_), .A2(
        u5_mult_79_SUMB_17__9_), .ZN(u5_mult_79_n1640) );
  NAND2_X2 u5_mult_79_U2577 ( .A1(u5_mult_79_SUMB_17__9_), .A2(
        u5_mult_79_CARRYB_17__8_), .ZN(u5_mult_79_n1641) );
  XNOR2_X2 u5_mult_79_U2576 ( .A(u5_mult_79_n1424), .B(
        u5_mult_79_CARRYB_18__7_), .ZN(u5_mult_79_n1638) );
  NAND2_X1 u5_mult_79_U2575 ( .A1(u5_mult_79_ab_7__13_), .A2(
        u5_mult_79_CARRYB_6__13_), .ZN(u5_mult_79_n1415) );
  NAND2_X1 u5_mult_79_U2574 ( .A1(u5_mult_79_ab_6__14_), .A2(
        u5_mult_79_CARRYB_5__14_), .ZN(u5_mult_79_n1412) );
  NAND3_X2 u5_mult_79_U2573 ( .A1(u5_mult_79_n1480), .A2(u5_mult_79_n1481), 
        .A3(u5_mult_79_n1482), .ZN(u5_mult_79_CARRYB_16__7_) );
  INV_X8 u5_mult_79_U2572 ( .A(n2967), .ZN(u5_mult_79_n1862) );
  INV_X16 u5_mult_79_U2571 ( .A(u5_mult_79_n1863), .ZN(u5_mult_79_n1789) );
  XNOR2_X2 u5_mult_79_U2570 ( .A(u5_mult_79_CARRYB_11__12_), .B(
        u5_mult_79_ab_12__12_), .ZN(u5_mult_79_n1411) );
  NOR2_X1 u5_mult_79_U2569 ( .A1(u5_mult_79_n1803), .A2(u5_mult_79_n1755), 
        .ZN(u5_mult_79_ab_13__10_) );
  NAND3_X2 u5_mult_79_U2568 ( .A1(u5_mult_79_n1405), .A2(u5_mult_79_n1406), 
        .A3(u5_mult_79_n1407), .ZN(u5_mult_79_CARRYB_12__11_) );
  NAND2_X1 u5_mult_79_U2567 ( .A1(u5_mult_79_ab_11__12_), .A2(
        u5_mult_79_CARRYB_10__12_), .ZN(u5_mult_79_n1402) );
  XOR2_X2 u5_mult_79_U2566 ( .A(u5_mult_79_n1401), .B(u5_mult_79_n307), .Z(
        u5_mult_79_SUMB_12__11_) );
  NAND2_X1 u5_mult_79_U2565 ( .A1(u5_mult_79_ab_7__16_), .A2(
        u5_mult_79_CARRYB_6__16_), .ZN(u5_mult_79_n1395) );
  NAND2_X1 u5_mult_79_U2564 ( .A1(u5_mult_79_ab_13__12_), .A2(
        u5_mult_79_SUMB_12__13_), .ZN(u5_mult_79_n1393) );
  NAND2_X1 u5_mult_79_U2563 ( .A1(u5_mult_79_ab_13__12_), .A2(
        u5_mult_79_CARRYB_12__12_), .ZN(u5_mult_79_n1392) );
  NAND3_X2 u5_mult_79_U2562 ( .A1(u5_mult_79_n1389), .A2(u5_mult_79_n1390), 
        .A3(u5_mult_79_n1391), .ZN(u5_mult_79_CARRYB_12__13_) );
  NAND2_X2 u5_mult_79_U2561 ( .A1(u5_mult_79_CARRYB_11__13_), .A2(
        u5_mult_79_n490), .ZN(u5_mult_79_n1391) );
  NAND2_X2 u5_mult_79_U2560 ( .A1(u5_mult_79_ab_12__13_), .A2(u5_mult_79_n490), 
        .ZN(u5_mult_79_n1390) );
  NAND2_X1 u5_mult_79_U2559 ( .A1(u5_mult_79_ab_12__13_), .A2(
        u5_mult_79_CARRYB_11__13_), .ZN(u5_mult_79_n1389) );
  NAND2_X2 u5_mult_79_U2558 ( .A1(u5_mult_79_ab_2__21_), .A2(
        u5_mult_79_CARRYB_1__21_), .ZN(u5_mult_79_n1624) );
  NAND2_X2 u5_mult_79_U2557 ( .A1(u5_mult_79_ab_2__21_), .A2(
        u5_mult_79_SUMB_1__22_), .ZN(u5_mult_79_n1623) );
  NOR2_X4 u5_mult_79_U2556 ( .A1(u5_mult_79_n1860), .A2(u5_mult_79_n1723), 
        .ZN(u5_mult_79_ab_2__21_) );
  INV_X8 u5_mult_79_U2555 ( .A(n3032), .ZN(u5_mult_79_n1864) );
  NAND2_X2 u5_mult_79_U2554 ( .A1(u5_mult_79_CARRYB_20__1_), .A2(
        u5_mult_79_ab_21__1_), .ZN(u5_mult_79_n1387) );
  NAND3_X2 u5_mult_79_U2553 ( .A1(u5_mult_79_n1383), .A2(u5_mult_79_n1384), 
        .A3(u5_mult_79_n1385), .ZN(u5_mult_79_CARRYB_20__1_) );
  NAND3_X2 u5_mult_79_U2552 ( .A1(u5_mult_79_n1380), .A2(u5_mult_79_n1381), 
        .A3(u5_mult_79_n1382), .ZN(u5_mult_79_CARRYB_4__15_) );
  NAND2_X1 u5_mult_79_U2551 ( .A1(u5_mult_79_CARRYB_3__15_), .A2(
        u5_mult_79_SUMB_3__16_), .ZN(u5_mult_79_n1382) );
  NAND2_X1 u5_mult_79_U2550 ( .A1(u5_mult_79_ab_4__15_), .A2(
        u5_mult_79_CARRYB_3__15_), .ZN(u5_mult_79_n1380) );
  NAND2_X1 u5_mult_79_U2549 ( .A1(u5_mult_79_ab_9__17_), .A2(
        u5_mult_79_CARRYB_8__17_), .ZN(u5_mult_79_n1373) );
  NAND2_X2 u5_mult_79_U2548 ( .A1(u5_mult_79_n1376), .A2(
        u5_mult_79_SUMB_7__19_), .ZN(u5_mult_79_n1372) );
  NAND2_X2 u5_mult_79_U2547 ( .A1(u5_mult_79_ab_8__18_), .A2(
        u5_mult_79_SUMB_7__19_), .ZN(u5_mult_79_n1371) );
  NAND2_X2 u5_mult_79_U2546 ( .A1(u5_mult_79_ab_8__18_), .A2(u5_mult_79_n1376), 
        .ZN(u5_mult_79_n1370) );
  XOR2_X2 u5_mult_79_U2545 ( .A(u5_mult_79_n1369), .B(u5_mult_79_SUMB_8__18_), 
        .Z(u5_mult_79_SUMB_9__17_) );
  XOR2_X2 u5_mult_79_U2544 ( .A(u5_mult_79_ab_9__17_), .B(
        u5_mult_79_CARRYB_8__17_), .Z(u5_mult_79_n1369) );
  XOR2_X2 u5_mult_79_U2543 ( .A(u5_mult_79_n1368), .B(u5_mult_79_SUMB_7__19_), 
        .Z(u5_mult_79_SUMB_8__18_) );
  NAND3_X4 u5_mult_79_U2542 ( .A1(u5_mult_79_n1367), .A2(u5_mult_79_n1366), 
        .A3(u5_mult_79_n1365), .ZN(u5_mult_79_CARRYB_16__11_) );
  NAND2_X2 u5_mult_79_U2541 ( .A1(u5_mult_79_ab_16__11_), .A2(
        u5_mult_79_SUMB_15__12_), .ZN(u5_mult_79_n1367) );
  NAND2_X2 u5_mult_79_U2540 ( .A1(u5_mult_79_n1268), .A2(
        u5_mult_79_SUMB_15__12_), .ZN(u5_mult_79_n1366) );
  NAND2_X1 u5_mult_79_U2539 ( .A1(u5_mult_79_CARRYB_15__11_), .A2(
        u5_mult_79_ab_16__11_), .ZN(u5_mult_79_n1365) );
  XNOR2_X2 u5_mult_79_U2538 ( .A(u5_mult_79_ab_15__15_), .B(
        u5_mult_79_CARRYB_14__15_), .ZN(u5_mult_79_n1361) );
  XNOR2_X2 u5_mult_79_U2537 ( .A(u5_mult_79_CARRYB_11__11_), .B(
        u5_mult_79_n1360), .ZN(u5_mult_79_n1401) );
  NOR2_X1 u5_mult_79_U2536 ( .A1(u5_mult_79_n1799), .A2(u5_mult_79_n1768), 
        .ZN(u5_mult_79_ab_17__12_) );
  NOR2_X1 u5_mult_79_U2535 ( .A1(u5_mult_79_n1805), .A2(u5_mult_79_n1859), 
        .ZN(u5_mult_79_ab_22__9_) );
  NAND3_X2 u5_mult_79_U2534 ( .A1(u5_mult_79_n1357), .A2(u5_mult_79_n1358), 
        .A3(u5_mult_79_n1359), .ZN(u5_mult_79_CARRYB_17__12_) );
  NAND2_X1 u5_mult_79_U2533 ( .A1(u5_mult_79_ab_17__12_), .A2(
        u5_mult_79_CARRYB_16__12_), .ZN(u5_mult_79_n1359) );
  NAND2_X2 u5_mult_79_U2532 ( .A1(u5_mult_79_ab_17__12_), .A2(
        u5_mult_79_SUMB_16__13_), .ZN(u5_mult_79_n1358) );
  NAND2_X1 u5_mult_79_U2531 ( .A1(u5_mult_79_SUMB_16__13_), .A2(
        u5_mult_79_CARRYB_16__12_), .ZN(u5_mult_79_n1357) );
  NAND2_X2 u5_mult_79_U2530 ( .A1(u5_mult_79_ab_22__9_), .A2(
        u5_mult_79_CARRYB_21__9_), .ZN(u5_mult_79_n1356) );
  NAND2_X2 u5_mult_79_U2529 ( .A1(u5_mult_79_ab_22__9_), .A2(
        u5_mult_79_SUMB_21__10_), .ZN(u5_mult_79_n1355) );
  NOR2_X1 u5_mult_79_U2528 ( .A1(u5_mult_79_n1785), .A2(u5_mult_79_n1726), 
        .ZN(u5_mult_79_ab_3__19_) );
  NOR2_X1 u5_mult_79_U2527 ( .A1(u5_mult_79_n1785), .A2(u5_mult_79_n1729), 
        .ZN(u5_mult_79_ab_4__19_) );
  NOR2_X1 u5_mult_79_U2526 ( .A1(u5_mult_79_n1785), .A2(u5_mult_79_n1732), 
        .ZN(u5_mult_79_ab_5__19_) );
  NOR2_X1 u5_mult_79_U2525 ( .A1(u5_mult_79_n1785), .A2(u5_mult_79_n1741), 
        .ZN(u5_mult_79_ab_8__19_) );
  NOR2_X1 u5_mult_79_U2524 ( .A1(u5_mult_79_n1785), .A2(u5_mult_79_n1744), 
        .ZN(u5_mult_79_ab_9__19_) );
  NOR2_X1 u5_mult_79_U2523 ( .A1(u5_mult_79_n1785), .A2(u5_mult_79_n1747), 
        .ZN(u5_mult_79_ab_10__19_) );
  NOR2_X1 u5_mult_79_U2522 ( .A1(u5_mult_79_n1785), .A2(u5_mult_79_n1859), 
        .ZN(u5_mult_79_ab_22__19_) );
  NOR2_X1 u5_mult_79_U2521 ( .A1(u5_mult_79_n1879), .A2(u5_mult_79_n1785), 
        .ZN(u5_mult_79_ab_23__19_) );
  NAND2_X2 u5_mult_79_U2520 ( .A1(u5_mult_79_ab_0__20_), .A2(
        u5_mult_79_ab_1__19_), .ZN(u5_mult_79_n1710) );
  NOR2_X4 u5_mult_79_U2519 ( .A1(u5_mult_79_n1882), .A2(u5_mult_79_n1862), 
        .ZN(u5_mult_79_ab_0__19_) );
  INV_X32 u5_mult_79_U2518 ( .A(u5_mult_79_n1786), .ZN(u5_mult_79_n1785) );
  INV_X8 u5_mult_79_U2517 ( .A(u5_mult_79_n1862), .ZN(u5_mult_79_n1786) );
  XNOR2_X2 u5_mult_79_U2516 ( .A(u5_mult_79_n337), .B(u5_mult_79_n1353), .ZN(
        u5_mult_79_n1625) );
  XNOR2_X2 u5_mult_79_U2515 ( .A(u5_mult_79_n1352), .B(
        u5_mult_79_CARRYB_21__2_), .ZN(u5_mult_79_n1504) );
  NAND3_X4 u5_mult_79_U2514 ( .A1(u5_mult_79_n1349), .A2(u5_mult_79_n1350), 
        .A3(u5_mult_79_n1351), .ZN(u5_mult_79_CARRYB_3__15_) );
  NAND2_X2 u5_mult_79_U2513 ( .A1(u5_mult_79_ab_3__15_), .A2(
        u5_mult_79_CARRYB_2__15_), .ZN(u5_mult_79_n1350) );
  NAND3_X2 u5_mult_79_U2512 ( .A1(u5_mult_79_n1346), .A2(u5_mult_79_n1347), 
        .A3(u5_mult_79_n1348), .ZN(u5_mult_79_CARRYB_2__15_) );
  NAND2_X1 u5_mult_79_U2511 ( .A1(u5_mult_79_CARRYB_1__15_), .A2(
        u5_mult_79_SUMB_1__16_), .ZN(u5_mult_79_n1348) );
  NAND2_X2 u5_mult_79_U2510 ( .A1(u5_mult_79_ab_2__15_), .A2(
        u5_mult_79_SUMB_1__16_), .ZN(u5_mult_79_n1347) );
  NAND2_X1 u5_mult_79_U2509 ( .A1(u5_mult_79_ab_2__15_), .A2(
        u5_mult_79_CARRYB_1__15_), .ZN(u5_mult_79_n1346) );
  NAND2_X1 u5_mult_79_U2508 ( .A1(u5_mult_79_ab_5__13_), .A2(
        u5_mult_79_CARRYB_4__13_), .ZN(u5_mult_79_n1343) );
  INV_X8 u5_mult_79_U2507 ( .A(n3039), .ZN(u5_mult_79_n1861) );
  NAND3_X4 u5_mult_79_U2506 ( .A1(u5_mult_79_n1568), .A2(u5_mult_79_n1567), 
        .A3(u5_mult_79_n1566), .ZN(u5_mult_79_CARRYB_17__10_) );
  NAND3_X2 u5_mult_79_U2505 ( .A1(u5_mult_79_n1332), .A2(u5_mult_79_n1333), 
        .A3(u5_mult_79_n1334), .ZN(u5_mult_79_CARRYB_15__14_) );
  NAND2_X2 u5_mult_79_U2504 ( .A1(u5_mult_79_ab_15__14_), .A2(u5_mult_79_n294), 
        .ZN(u5_mult_79_n1333) );
  NAND2_X1 u5_mult_79_U2503 ( .A1(u5_mult_79_ab_15__14_), .A2(
        u5_mult_79_CARRYB_14__14_), .ZN(u5_mult_79_n1332) );
  INV_X8 u5_mult_79_U2502 ( .A(n2942), .ZN(u5_mult_79_n1866) );
  AND2_X2 u5_mult_79_U2501 ( .A1(u5_mult_79_n1789), .A2(n3000), .ZN(
        u5_mult_79_ab_2__18_) );
  XNOR2_X2 u5_mult_79_U2500 ( .A(u5_mult_79_n1331), .B(u5_mult_79_SUMB_14__13_), .ZN(u5_mult_79_SUMB_15__12_) );
  XNOR2_X2 u5_mult_79_U2499 ( .A(u5_mult_79_SUMB_22__3_), .B(u5_mult_79_n1330), 
        .ZN(u5_mult_79_n1508) );
  NOR2_X2 u5_mult_79_U2498 ( .A1(u5_mult_79_n1806), .A2(u5_mult_79_n1758), 
        .ZN(u5_mult_79_ab_14__9_) );
  NOR2_X1 u5_mult_79_U2497 ( .A1(u5_mult_79_n1868), .A2(u5_mult_79_n1741), 
        .ZN(u5_mult_79_ab_8__13_) );
  NAND2_X1 u5_mult_79_U2496 ( .A1(u5_mult_79_ab_8__13_), .A2(u5_mult_79_n268), 
        .ZN(u5_mult_79_n1326) );
  NAND2_X2 u5_mult_79_U2495 ( .A1(u5_mult_79_n32), .A2(u5_mult_79_ab_8__13_), 
        .ZN(u5_mult_79_n1325) );
  NAND2_X2 u5_mult_79_U2494 ( .A1(u5_mult_79_CARRYB_14__9_), .A2(
        u5_mult_79_n463), .ZN(u5_mult_79_n1320) );
  NAND2_X2 u5_mult_79_U2493 ( .A1(u5_mult_79_n463), .A2(u5_mult_79_ab_15__9_), 
        .ZN(u5_mult_79_n1319) );
  NAND2_X2 u5_mult_79_U2492 ( .A1(u5_mult_79_ab_4__14_), .A2(
        u5_mult_79_CARRYB_3__14_), .ZN(u5_mult_79_n1340) );
  XNOR2_X2 u5_mult_79_U2491 ( .A(u5_mult_79_n1315), .B(u5_mult_79_SUMB_15__8_), 
        .ZN(u5_mult_79_SUMB_16__7_) );
  NAND2_X2 u5_mult_79_U2490 ( .A1(u5_mult_79_ab_16__8_), .A2(
        u5_mult_79_CARRYB_15__8_), .ZN(u5_mult_79_n1321) );
  NAND2_X2 u5_mult_79_U2489 ( .A1(u5_mult_79_CARRYB_15__8_), .A2(
        u5_mult_79_SUMB_15__9_), .ZN(u5_mult_79_n1323) );
  NOR2_X1 u5_mult_79_U2488 ( .A1(u5_mult_79_n1831), .A2(u5_mult_79_n1731), 
        .ZN(u5_mult_79_ab_5__23_) );
  NOR2_X1 u5_mult_79_U2487 ( .A1(u5_mult_79_n1780), .A2(u5_mult_79_n1735), 
        .ZN(u5_mult_79_ab_6__22_) );
  NAND3_X2 u5_mult_79_U2486 ( .A1(u5_mult_79_n1312), .A2(u5_mult_79_n1313), 
        .A3(u5_mult_79_n1314), .ZN(u5_mult_79_CARRYB_6__22_) );
  NAND2_X2 u5_mult_79_U2485 ( .A1(u5_mult_79_ab_5__23_), .A2(
        u5_mult_79_ab_6__22_), .ZN(u5_mult_79_n1314) );
  NAND2_X2 u5_mult_79_U2484 ( .A1(u5_mult_79_n498), .A2(u5_mult_79_ab_5__23_), 
        .ZN(u5_mult_79_n1313) );
  NAND2_X2 u5_mult_79_U2483 ( .A1(u5_mult_79_ab_6__22_), .A2(u5_mult_79_n498), 
        .ZN(u5_mult_79_n1312) );
  NAND2_X1 u5_mult_79_U2482 ( .A1(u5_mult_79_n213), .A2(
        u5_mult_79_SUMB_22__11_), .ZN(u5_mult_79_n1311) );
  NAND2_X1 u5_mult_79_U2481 ( .A1(u5_mult_79_ab_23__10_), .A2(
        u5_mult_79_SUMB_22__11_), .ZN(u5_mult_79_n1310) );
  NAND2_X1 u5_mult_79_U2480 ( .A1(u5_mult_79_ab_23__10_), .A2(u5_mult_79_n213), 
        .ZN(u5_mult_79_n1309) );
  NAND2_X1 u5_mult_79_U2479 ( .A1(u5_mult_79_ab_22__11_), .A2(
        u5_mult_79_SUMB_21__12_), .ZN(u5_mult_79_n1307) );
  XNOR2_X2 u5_mult_79_U2478 ( .A(u5_mult_79_ab_16__7_), .B(
        u5_mult_79_CARRYB_15__7_), .ZN(u5_mult_79_n1315) );
  XNOR2_X2 u5_mult_79_U2477 ( .A(u5_mult_79_ab_16__12_), .B(
        u5_mult_79_CARRYB_15__12_), .ZN(u5_mult_79_n1305) );
  NAND2_X2 u5_mult_79_U2476 ( .A1(u5_mult_79_ab_12__12_), .A2(
        u5_mult_79_SUMB_11__13_), .ZN(u5_mult_79_n1422) );
  NAND2_X2 u5_mult_79_U2475 ( .A1(u5_mult_79_CARRYB_11__12_), .A2(
        u5_mult_79_SUMB_11__13_), .ZN(u5_mult_79_n1423) );
  NAND2_X1 u5_mult_79_U2474 ( .A1(u5_mult_79_CARRYB_12__12_), .A2(
        u5_mult_79_SUMB_12__13_), .ZN(u5_mult_79_n1394) );
  XNOR2_X2 u5_mult_79_U2473 ( .A(u5_mult_79_ab_22__5_), .B(
        u5_mult_79_CARRYB_21__5_), .ZN(u5_mult_79_n1303) );
  NAND2_X2 u5_mult_79_U2472 ( .A1(u5_mult_79_ab_19__5_), .A2(
        u5_mult_79_SUMB_18__6_), .ZN(u5_mult_79_n1598) );
  XNOR2_X2 u5_mult_79_U2471 ( .A(u5_mult_79_n124), .B(u5_mult_79_n1302), .ZN(
        u5_mult_79_SUMB_17__7_) );
  XNOR2_X2 u5_mult_79_U2470 ( .A(u5_mult_79_CARRYB_21__9_), .B(
        u5_mult_79_ab_22__9_), .ZN(u5_mult_79_n1301) );
  XNOR2_X2 u5_mult_79_U2469 ( .A(u5_mult_79_n361), .B(u5_mult_79_n1301), .ZN(
        u5_mult_79_SUMB_22__9_) );
  XNOR2_X2 u5_mult_79_U2468 ( .A(u5_mult_79_n1300), .B(u5_mult_79_n321), .ZN(
        u5_mult_79_SUMB_20__3_) );
  XNOR2_X2 u5_mult_79_U2467 ( .A(u5_mult_79_ab_2__15_), .B(
        u5_mult_79_CARRYB_1__15_), .ZN(u5_mult_79_n1299) );
  XNOR2_X2 u5_mult_79_U2466 ( .A(u5_mult_79_n1299), .B(u5_mult_79_SUMB_1__16_), 
        .ZN(u5_mult_79_SUMB_2__15_) );
  NOR2_X1 u5_mult_79_U2465 ( .A1(u5_mult_79_n1793), .A2(u5_mult_79_n1729), 
        .ZN(u5_mult_79_ab_4__16_) );
  NOR2_X2 u5_mult_79_U2464 ( .A1(u5_mult_79_n1806), .A2(u5_mult_79_n1755), 
        .ZN(u5_mult_79_ab_13__9_) );
  NAND2_X2 u5_mult_79_U2463 ( .A1(u5_mult_79_ab_10__12_), .A2(
        u5_mult_79_SUMB_9__13_), .ZN(u5_mult_79_n1297) );
  NAND2_X1 u5_mult_79_U2462 ( .A1(u5_mult_79_ab_10__12_), .A2(
        u5_mult_79_CARRYB_9__12_), .ZN(u5_mult_79_n1296) );
  NAND2_X2 u5_mult_79_U2461 ( .A1(u5_mult_79_CARRYB_8__13_), .A2(
        u5_mult_79_SUMB_8__14_), .ZN(u5_mult_79_n1295) );
  NAND2_X2 u5_mult_79_U2460 ( .A1(u5_mult_79_ab_9__13_), .A2(
        u5_mult_79_SUMB_8__14_), .ZN(u5_mult_79_n1294) );
  NAND2_X1 u5_mult_79_U2459 ( .A1(u5_mult_79_ab_4__16_), .A2(u5_mult_79_n269), 
        .ZN(u5_mult_79_n1292) );
  NAND2_X2 u5_mult_79_U2458 ( .A1(u5_mult_79_ab_4__16_), .A2(
        u5_mult_79_SUMB_3__17_), .ZN(u5_mult_79_n1291) );
  NAND3_X4 u5_mult_79_U2457 ( .A1(u5_mult_79_n1284), .A2(u5_mult_79_n1285), 
        .A3(u5_mult_79_n1286), .ZN(u5_mult_79_CARRYB_14__8_) );
  NAND2_X2 u5_mult_79_U2456 ( .A1(u5_mult_79_SUMB_13__9_), .A2(
        u5_mult_79_CARRYB_13__8_), .ZN(u5_mult_79_n1286) );
  NAND2_X2 u5_mult_79_U2455 ( .A1(u5_mult_79_SUMB_13__9_), .A2(
        u5_mult_79_ab_14__8_), .ZN(u5_mult_79_n1285) );
  NAND2_X1 u5_mult_79_U2454 ( .A1(u5_mult_79_ab_14__8_), .A2(
        u5_mult_79_CARRYB_13__8_), .ZN(u5_mult_79_n1284) );
  NAND3_X4 u5_mult_79_U2453 ( .A1(u5_mult_79_n1281), .A2(u5_mult_79_n1282), 
        .A3(u5_mult_79_n1283), .ZN(u5_mult_79_CARRYB_13__9_) );
  NAND2_X2 u5_mult_79_U2452 ( .A1(u5_mult_79_ab_13__9_), .A2(
        u5_mult_79_CARRYB_12__9_), .ZN(u5_mult_79_n1283) );
  NAND2_X2 u5_mult_79_U2451 ( .A1(u5_mult_79_ab_13__9_), .A2(
        u5_mult_79_SUMB_12__10_), .ZN(u5_mult_79_n1282) );
  NAND2_X2 u5_mult_79_U2450 ( .A1(u5_mult_79_CARRYB_12__9_), .A2(
        u5_mult_79_SUMB_12__10_), .ZN(u5_mult_79_n1281) );
  NAND3_X2 u5_mult_79_U2449 ( .A1(u5_mult_79_n1278), .A2(u5_mult_79_n1279), 
        .A3(u5_mult_79_n1280), .ZN(u5_mult_79_CARRYB_8__17_) );
  NAND2_X2 u5_mult_79_U2448 ( .A1(u5_mult_79_SUMB_7__18_), .A2(
        u5_mult_79_ab_8__17_), .ZN(u5_mult_79_n1279) );
  NAND3_X2 u5_mult_79_U2447 ( .A1(u5_mult_79_n1275), .A2(u5_mult_79_n1276), 
        .A3(u5_mult_79_n1277), .ZN(u5_mult_79_CARRYB_7__18_) );
  NAND3_X2 u5_mult_79_U2446 ( .A1(u5_mult_79_n1272), .A2(u5_mult_79_n1273), 
        .A3(u5_mult_79_n1274), .ZN(u5_mult_79_CARRYB_10__15_) );
  NAND2_X1 u5_mult_79_U2445 ( .A1(u5_mult_79_ab_10__15_), .A2(
        u5_mult_79_CARRYB_9__15_), .ZN(u5_mult_79_n1272) );
  XNOR2_X2 u5_mult_79_U2444 ( .A(u5_mult_79_ab_12__13_), .B(
        u5_mult_79_CARRYB_11__13_), .ZN(u5_mult_79_n1267) );
  XNOR2_X2 u5_mult_79_U2443 ( .A(u5_mult_79_n1267), .B(u5_mult_79_n490), .ZN(
        u5_mult_79_SUMB_12__13_) );
  NAND3_X2 u5_mult_79_U2442 ( .A1(u5_mult_79_n1580), .A2(u5_mult_79_n1579), 
        .A3(u5_mult_79_n1581), .ZN(u5_mult_79_CARRYB_4__18_) );
  INV_X8 u5_mult_79_U2441 ( .A(n2962), .ZN(u5_mult_79_n1865) );
  XNOR2_X2 u5_mult_79_U2440 ( .A(u5_mult_79_n1266), .B(
        u5_mult_79_CARRYB_2__15_), .ZN(u5_mult_79_SUMB_3__15_) );
  NAND2_X2 u5_mult_79_U2439 ( .A1(u5_mult_79_ab_16__10_), .A2(
        u5_mult_79_SUMB_15__11_), .ZN(u5_mult_79_n1493) );
  XNOR2_X2 u5_mult_79_U2438 ( .A(u5_mult_79_ab_23__9_), .B(
        u5_mult_79_CARRYB_22__9_), .ZN(u5_mult_79_n1265) );
  XNOR2_X2 u5_mult_79_U2437 ( .A(u5_mult_79_n1265), .B(u5_mult_79_n110), .ZN(
        u5_mult_79_SUMB_23__9_) );
  XNOR2_X2 u5_mult_79_U2436 ( .A(u5_mult_79_CARRYB_3__20_), .B(
        u5_mult_79_ab_4__20_), .ZN(u5_mult_79_n1264) );
  XNOR2_X2 u5_mult_79_U2435 ( .A(u5_mult_79_CARRYB_22__10_), .B(
        u5_mult_79_ab_23__10_), .ZN(u5_mult_79_n1263) );
  XNOR2_X2 u5_mult_79_U2434 ( .A(u5_mult_79_n1263), .B(u5_mult_79_SUMB_22__11_), .ZN(u5_mult_79_SUMB_23__10_) );
  NOR2_X2 u5_mult_79_U2433 ( .A1(u5_mult_79_n1867), .A2(u5_mult_79_n1726), 
        .ZN(u5_mult_79_ab_3__14_) );
  NAND2_X1 u5_mult_79_U2432 ( .A1(u5_mult_79_ab_20__2_), .A2(
        u5_mult_79_SUMB_19__3_), .ZN(u5_mult_79_n1261) );
  NAND2_X1 u5_mult_79_U2431 ( .A1(u5_mult_79_CARRYB_19__2_), .A2(
        u5_mult_79_SUMB_19__3_), .ZN(u5_mult_79_n1260) );
  NAND3_X2 u5_mult_79_U2430 ( .A1(u5_mult_79_n1254), .A2(u5_mult_79_n1255), 
        .A3(u5_mult_79_n1256), .ZN(u5_mult_79_CARRYB_7__10_) );
  NAND2_X1 u5_mult_79_U2429 ( .A1(u5_mult_79_ab_7__10_), .A2(
        u5_mult_79_CARRYB_6__10_), .ZN(u5_mult_79_n1254) );
  NAND3_X2 u5_mult_79_U2428 ( .A1(u5_mult_79_n1253), .A2(u5_mult_79_n1252), 
        .A3(u5_mult_79_n1251), .ZN(u5_mult_79_CARRYB_6__11_) );
  NAND2_X2 u5_mult_79_U2427 ( .A1(u5_mult_79_n285), .A2(
        u5_mult_79_CARRYB_5__11_), .ZN(u5_mult_79_n1253) );
  NAND2_X2 u5_mult_79_U2426 ( .A1(u5_mult_79_SUMB_5__12_), .A2(
        u5_mult_79_ab_6__11_), .ZN(u5_mult_79_n1252) );
  NAND2_X1 u5_mult_79_U2425 ( .A1(u5_mult_79_ab_6__11_), .A2(
        u5_mult_79_CARRYB_5__11_), .ZN(u5_mult_79_n1251) );
  XOR2_X2 u5_mult_79_U2424 ( .A(u5_mult_79_n1250), .B(u5_mult_79_n285), .Z(
        u5_mult_79_SUMB_6__11_) );
  NAND3_X2 u5_mult_79_U2423 ( .A1(u5_mult_79_n1247), .A2(u5_mult_79_n1248), 
        .A3(u5_mult_79_n1249), .ZN(u5_mult_79_CARRYB_3__14_) );
  NAND2_X2 u5_mult_79_U2422 ( .A1(u5_mult_79_ab_3__14_), .A2(
        u5_mult_79_CARRYB_2__14_), .ZN(u5_mult_79_n1248) );
  XNOR2_X2 u5_mult_79_U2421 ( .A(u5_mult_79_n1246), .B(u5_mult_79_n300), .ZN(
        u5_mult_79_SUMB_19__10_) );
  NOR2_X1 u5_mult_79_U2420 ( .A1(u5_mult_79_n1814), .A2(u5_mult_79_n1859), 
        .ZN(u5_mult_79_ab_22__6_) );
  NAND3_X2 u5_mult_79_U2419 ( .A1(u5_mult_79_n1243), .A2(u5_mult_79_n1244), 
        .A3(u5_mult_79_n1245), .ZN(u5_mult_79_CARRYB_22__6_) );
  NAND2_X1 u5_mult_79_U2418 ( .A1(u5_mult_79_ab_22__6_), .A2(
        u5_mult_79_CARRYB_21__6_), .ZN(u5_mult_79_n1245) );
  NAND2_X2 u5_mult_79_U2417 ( .A1(u5_mult_79_ab_22__6_), .A2(
        u5_mult_79_SUMB_21__7_), .ZN(u5_mult_79_n1244) );
  NAND2_X2 u5_mult_79_U2416 ( .A1(u5_mult_79_ab_15__12_), .A2(
        u5_mult_79_CARRYB_14__12_), .ZN(u5_mult_79_n1241) );
  NAND3_X2 u5_mult_79_U2415 ( .A1(u5_mult_79_n1237), .A2(u5_mult_79_n1236), 
        .A3(u5_mult_79_n1238), .ZN(u5_mult_79_CARRYB_14__17_) );
  NAND2_X1 u5_mult_79_U2414 ( .A1(u5_mult_79_CARRYB_13__17_), .A2(
        u5_mult_79_SUMB_13__18_), .ZN(u5_mult_79_n1238) );
  NAND2_X1 u5_mult_79_U2413 ( .A1(u5_mult_79_ab_14__17_), .A2(
        u5_mult_79_SUMB_13__18_), .ZN(u5_mult_79_n1237) );
  NAND2_X1 u5_mult_79_U2412 ( .A1(u5_mult_79_ab_14__17_), .A2(
        u5_mult_79_CARRYB_13__17_), .ZN(u5_mult_79_n1236) );
  NAND2_X2 u5_mult_79_U2411 ( .A1(u5_mult_79_ab_13__18_), .A2(
        u5_mult_79_SUMB_12__19_), .ZN(u5_mult_79_n1234) );
  NAND2_X1 u5_mult_79_U2410 ( .A1(u5_mult_79_ab_13__18_), .A2(
        u5_mult_79_CARRYB_12__18_), .ZN(u5_mult_79_n1233) );
  XOR2_X2 u5_mult_79_U2409 ( .A(u5_mult_79_n1232), .B(u5_mult_79_n477), .Z(
        u5_mult_79_SUMB_13__18_) );
  NAND2_X2 u5_mult_79_U2408 ( .A1(u5_mult_79_ab_6__21_), .A2(u5_mult_79_n436), 
        .ZN(u5_mult_79_n1227) );
  NAND2_X1 u5_mult_79_U2407 ( .A1(u5_mult_79_ab_6__21_), .A2(
        u5_mult_79_CARRYB_5__21_), .ZN(u5_mult_79_n1226) );
  NAND3_X2 u5_mult_79_U2406 ( .A1(u5_mult_79_n1223), .A2(u5_mult_79_n1224), 
        .A3(u5_mult_79_n1225), .ZN(u5_mult_79_CARRYB_20__11_) );
  NAND2_X1 u5_mult_79_U2405 ( .A1(u5_mult_79_ab_20__11_), .A2(
        u5_mult_79_CARRYB_19__11_), .ZN(u5_mult_79_n1223) );
  NAND2_X2 u5_mult_79_U2404 ( .A1(u5_mult_79_SUMB_18__13_), .A2(
        u5_mult_79_CARRYB_18__12_), .ZN(u5_mult_79_n1222) );
  NAND2_X2 u5_mult_79_U2403 ( .A1(u5_mult_79_ab_19__12_), .A2(
        u5_mult_79_SUMB_18__13_), .ZN(u5_mult_79_n1221) );
  INV_X1 u5_mult_79_U2402 ( .A(u5_mult_79_SUMB_3__20_), .ZN(u5_mult_79_n1217)
         );
  NAND2_X2 u5_mult_79_U2401 ( .A1(u5_mult_79_n1216), .A2(u5_mult_79_n1217), 
        .ZN(u5_mult_79_n1219) );
  INV_X4 u5_mult_79_U2400 ( .A(u5_mult_79_n1525), .ZN(u5_mult_79_n1212) );
  NAND3_X4 u5_mult_79_U2399 ( .A1(u5_mult_79_n1209), .A2(u5_mult_79_n1210), 
        .A3(u5_mult_79_n1211), .ZN(u5_mult_79_CARRYB_9__15_) );
  NAND2_X2 u5_mult_79_U2398 ( .A1(u5_mult_79_ab_9__15_), .A2(
        u5_mult_79_SUMB_8__16_), .ZN(u5_mult_79_n1210) );
  NAND2_X1 u5_mult_79_U2397 ( .A1(u5_mult_79_ab_9__15_), .A2(
        u5_mult_79_CARRYB_8__15_), .ZN(u5_mult_79_n1209) );
  NAND2_X2 u5_mult_79_U2396 ( .A1(u5_mult_79_CARRYB_7__16_), .A2(
        u5_mult_79_n89), .ZN(u5_mult_79_n1208) );
  NAND2_X2 u5_mult_79_U2395 ( .A1(u5_mult_79_ab_8__16_), .A2(u5_mult_79_n89), 
        .ZN(u5_mult_79_n1207) );
  INV_X1 u5_mult_79_U2394 ( .A(u5_mult_79_ab_17__11_), .ZN(u5_mult_79_n1202)
         );
  NAND2_X2 u5_mult_79_U2393 ( .A1(u5_mult_79_ab_16__6_), .A2(
        u5_mult_79_SUMB_15__7_), .ZN(u5_mult_79_n1577) );
  NAND2_X2 u5_mult_79_U2392 ( .A1(u5_mult_79_ab_19__5_), .A2(
        u5_mult_79_CARRYB_18__5_), .ZN(u5_mult_79_n1597) );
  NAND2_X2 u5_mult_79_U2391 ( .A1(u5_mult_79_CARRYB_18__5_), .A2(
        u5_mult_79_SUMB_18__6_), .ZN(u5_mult_79_n1599) );
  NOR2_X1 u5_mult_79_U2390 ( .A1(u5_mult_79_n1818), .A2(u5_mult_79_n1770), 
        .ZN(u5_mult_79_ab_18__5_) );
  NAND3_X4 u5_mult_79_U2389 ( .A1(u5_mult_79_n1199), .A2(u5_mult_79_n1200), 
        .A3(u5_mult_79_n1201), .ZN(u5_mult_79_CARRYB_18__5_) );
  NAND2_X2 u5_mult_79_U2388 ( .A1(u5_mult_79_ab_18__5_), .A2(
        u5_mult_79_SUMB_17__6_), .ZN(u5_mult_79_n1200) );
  XOR2_X2 u5_mult_79_U2387 ( .A(u5_mult_79_n1198), .B(u5_mult_79_n491), .Z(
        u5_mult_79_SUMB_18__5_) );
  NAND3_X2 u5_mult_79_U2386 ( .A1(u5_mult_79_n1195), .A2(u5_mult_79_n1196), 
        .A3(u5_mult_79_n1197), .ZN(u5_mult_79_CARRYB_3__13_) );
  NAND2_X1 u5_mult_79_U2385 ( .A1(u5_mult_79_SUMB_2__14_), .A2(
        u5_mult_79_CARRYB_2__13_), .ZN(u5_mult_79_n1197) );
  NAND2_X1 u5_mult_79_U2384 ( .A1(u5_mult_79_ab_3__13_), .A2(
        u5_mult_79_SUMB_2__14_), .ZN(u5_mult_79_n1196) );
  NAND2_X1 u5_mult_79_U2383 ( .A1(u5_mult_79_ab_3__13_), .A2(
        u5_mult_79_CARRYB_2__13_), .ZN(u5_mult_79_n1195) );
  NAND3_X4 u5_mult_79_U2382 ( .A1(u5_mult_79_n1192), .A2(u5_mult_79_n1193), 
        .A3(u5_mult_79_n1194), .ZN(u5_mult_79_CARRYB_2__14_) );
  NAND2_X2 u5_mult_79_U2381 ( .A1(u5_mult_79_CARRYB_1__14_), .A2(
        u5_mult_79_SUMB_1__15_), .ZN(u5_mult_79_n1194) );
  NAND2_X2 u5_mult_79_U2380 ( .A1(u5_mult_79_ab_2__14_), .A2(
        u5_mult_79_SUMB_1__15_), .ZN(u5_mult_79_n1193) );
  NAND2_X2 u5_mult_79_U2379 ( .A1(u5_mult_79_ab_2__14_), .A2(
        u5_mult_79_CARRYB_1__14_), .ZN(u5_mult_79_n1192) );
  XOR2_X2 u5_mult_79_U2378 ( .A(u5_mult_79_n1191), .B(u5_mult_79_SUMB_1__15_), 
        .Z(u5_mult_79_SUMB_2__14_) );
  XOR2_X2 u5_mult_79_U2377 ( .A(u5_mult_79_ab_2__14_), .B(
        u5_mult_79_CARRYB_1__14_), .Z(u5_mult_79_n1191) );
  NAND3_X2 u5_mult_79_U2376 ( .A1(u5_mult_79_n1188), .A2(u5_mult_79_n1189), 
        .A3(u5_mult_79_n1190), .ZN(u5_mult_79_CARRYB_22__4_) );
  NAND2_X1 u5_mult_79_U2375 ( .A1(u5_mult_79_ab_22__4_), .A2(
        u5_mult_79_SUMB_21__5_), .ZN(u5_mult_79_n1190) );
  NAND2_X1 u5_mult_79_U2374 ( .A1(u5_mult_79_SUMB_21__5_), .A2(
        u5_mult_79_CARRYB_21__4_), .ZN(u5_mult_79_n1189) );
  NAND2_X1 u5_mult_79_U2373 ( .A1(u5_mult_79_ab_22__4_), .A2(
        u5_mult_79_CARRYB_21__4_), .ZN(u5_mult_79_n1188) );
  NAND2_X2 u5_mult_79_U2372 ( .A1(u5_mult_79_n457), .A2(u5_mult_79_n466), .ZN(
        u5_mult_79_n1187) );
  NAND2_X2 u5_mult_79_U2371 ( .A1(u5_mult_79_ab_21__5_), .A2(u5_mult_79_n466), 
        .ZN(u5_mult_79_n1186) );
  NAND2_X1 u5_mult_79_U2370 ( .A1(u5_mult_79_CARRYB_2__14_), .A2(
        u5_mult_79_SUMB_2__15_), .ZN(u5_mult_79_n1247) );
  NAND2_X2 u5_mult_79_U2369 ( .A1(u5_mult_79_n324), .A2(
        u5_mult_79_CARRYB_2__15_), .ZN(u5_mult_79_n1351) );
  NAND3_X2 u5_mult_79_U2368 ( .A1(u5_mult_79_n1260), .A2(u5_mult_79_n1261), 
        .A3(u5_mult_79_n1262), .ZN(u5_mult_79_CARRYB_20__2_) );
  NAND2_X2 u5_mult_79_U2367 ( .A1(u5_mult_79_ab_3__16_), .A2(
        u5_mult_79_CARRYB_2__16_), .ZN(u5_mult_79_n1377) );
  NOR2_X1 u5_mult_79_U2366 ( .A1(u5_mult_79_n1823), .A2(u5_mult_79_n1770), 
        .ZN(u5_mult_79_ab_18__3_) );
  NOR2_X1 u5_mult_79_U2365 ( .A1(u5_mult_79_n1828), .A2(u5_mult_79_n1859), 
        .ZN(u5_mult_79_ab_22__1_) );
  NAND2_X2 u5_mult_79_U2364 ( .A1(u5_mult_79_ab_2__16_), .A2(
        u5_mult_79_CARRYB_1__16_), .ZN(u5_mult_79_n1182) );
  NAND3_X2 u5_mult_79_U2363 ( .A1(u5_mult_79_n1178), .A2(u5_mult_79_n1179), 
        .A3(u5_mult_79_n1180), .ZN(u5_mult_79_CARRYB_18__3_) );
  NAND2_X1 u5_mult_79_U2362 ( .A1(u5_mult_79_SUMB_17__4_), .A2(
        u5_mult_79_ab_18__3_), .ZN(u5_mult_79_n1180) );
  NAND2_X2 u5_mult_79_U2361 ( .A1(u5_mult_79_ab_22__1_), .A2(
        u5_mult_79_SUMB_21__2_), .ZN(u5_mult_79_n1176) );
  NAND2_X2 u5_mult_79_U2360 ( .A1(u5_mult_79_ab_19__4_), .A2(
        u5_mult_79_SUMB_18__5_), .ZN(u5_mult_79_n1589) );
  NAND2_X2 u5_mult_79_U2359 ( .A1(u5_mult_79_n1130), .A2(
        u5_mult_79_SUMB_16__6_), .ZN(u5_mult_79_n1474) );
  NOR2_X2 u5_mult_79_U2358 ( .A1(u5_mult_79_n1834), .A2(u5_mult_79_n1829), 
        .ZN(u5_mult_79_ab_23__0_) );
  NAND2_X2 u5_mult_79_U2357 ( .A1(u5_mult_79_ab_23__0_), .A2(
        u5_mult_79_SUMB_22__1_), .ZN(u5_mult_79_n1174) );
  NAND3_X2 u5_mult_79_U2356 ( .A1(u5_mult_79_n1168), .A2(u5_mult_79_n1169), 
        .A3(u5_mult_79_n1170), .ZN(u5_mult_79_CARRYB_8__7_) );
  NAND2_X1 u5_mult_79_U2355 ( .A1(u5_mult_79_ab_8__7_), .A2(
        u5_mult_79_SUMB_7__8_), .ZN(u5_mult_79_n1169) );
  NAND3_X2 u5_mult_79_U2354 ( .A1(u5_mult_79_n1165), .A2(u5_mult_79_n1166), 
        .A3(u5_mult_79_n1167), .ZN(u5_mult_79_CARRYB_7__8_) );
  NAND2_X2 u5_mult_79_U2353 ( .A1(u5_mult_79_ab_7__8_), .A2(
        u5_mult_79_SUMB_6__9_), .ZN(u5_mult_79_n1166) );
  NAND2_X1 u5_mult_79_U2352 ( .A1(u5_mult_79_ab_7__8_), .A2(u5_mult_79_n10), 
        .ZN(u5_mult_79_n1165) );
  NAND3_X2 u5_mult_79_U2351 ( .A1(u5_mult_79_n1161), .A2(u5_mult_79_n1162), 
        .A3(u5_mult_79_n1163), .ZN(u5_mult_79_CARRYB_4__11_) );
  NAND2_X1 u5_mult_79_U2350 ( .A1(u5_mult_79_CARRYB_3__11_), .A2(
        u5_mult_79_SUMB_3__12_), .ZN(u5_mult_79_n1163) );
  NAND2_X1 u5_mult_79_U2349 ( .A1(u5_mult_79_ab_4__11_), .A2(
        u5_mult_79_SUMB_3__12_), .ZN(u5_mult_79_n1162) );
  NAND2_X1 u5_mult_79_U2348 ( .A1(u5_mult_79_ab_4__11_), .A2(
        u5_mult_79_CARRYB_3__11_), .ZN(u5_mult_79_n1161) );
  NAND2_X2 u5_mult_79_U2347 ( .A1(u5_mult_79_CARRYB_2__12_), .A2(
        u5_mult_79_SUMB_2__13_), .ZN(u5_mult_79_n1160) );
  NAND2_X2 u5_mult_79_U2346 ( .A1(u5_mult_79_ab_3__12_), .A2(
        u5_mult_79_SUMB_2__13_), .ZN(u5_mult_79_n1159) );
  NAND2_X1 u5_mult_79_U2345 ( .A1(u5_mult_79_ab_3__12_), .A2(
        u5_mult_79_CARRYB_2__12_), .ZN(u5_mult_79_n1158) );
  XOR2_X2 u5_mult_79_U2344 ( .A(u5_mult_79_n1157), .B(u5_mult_79_SUMB_3__12_), 
        .Z(u5_mult_79_SUMB_4__11_) );
  XOR2_X2 u5_mult_79_U2343 ( .A(u5_mult_79_ab_4__11_), .B(
        u5_mult_79_CARRYB_3__11_), .Z(u5_mult_79_n1157) );
  XOR2_X2 u5_mult_79_U2342 ( .A(u5_mult_79_n1156), .B(u5_mult_79_n326), .Z(
        u5_mult_79_SUMB_3__12_) );
  XOR2_X2 u5_mult_79_U2341 ( .A(u5_mult_79_ab_3__12_), .B(
        u5_mult_79_CARRYB_2__12_), .Z(u5_mult_79_n1156) );
  NAND2_X1 u5_mult_79_U2340 ( .A1(u5_mult_79_CARRYB_23__9_), .A2(
        u5_mult_79_SUMB_23__10_), .ZN(u5_mult_79_n1656) );
  NOR2_X1 u5_mult_79_U2339 ( .A1(u5_mult_79_n1829), .A2(u5_mult_79_n1798), 
        .ZN(u5_mult_79_ab_23__12_) );
  NAND3_X2 u5_mult_79_U2338 ( .A1(u5_mult_79_n1153), .A2(u5_mult_79_n1154), 
        .A3(u5_mult_79_n1155), .ZN(u5_mult_79_CARRYB_23__12_) );
  NAND2_X1 u5_mult_79_U2337 ( .A1(u5_mult_79_ab_23__12_), .A2(
        u5_mult_79_CARRYB_22__12_), .ZN(u5_mult_79_n1155) );
  NAND2_X1 u5_mult_79_U2336 ( .A1(u5_mult_79_ab_23__12_), .A2(
        u5_mult_79_SUMB_22__13_), .ZN(u5_mult_79_n1154) );
  NAND2_X1 u5_mult_79_U2335 ( .A1(u5_mult_79_CARRYB_22__12_), .A2(
        u5_mult_79_SUMB_22__13_), .ZN(u5_mult_79_n1153) );
  NAND2_X2 u5_mult_79_U2334 ( .A1(u5_mult_79_ab_5__20_), .A2(
        u5_mult_79_SUMB_4__21_), .ZN(u5_mult_79_n1151) );
  NAND3_X2 u5_mult_79_U2333 ( .A1(u5_mult_79_n1354), .A2(u5_mult_79_n1355), 
        .A3(u5_mult_79_n1356), .ZN(u5_mult_79_CARRYB_22__9_) );
  XNOR2_X2 u5_mult_79_U2332 ( .A(u5_mult_79_CARRYB_13__17_), .B(
        u5_mult_79_ab_14__17_), .ZN(u5_mult_79_n1148) );
  NAND2_X2 u5_mult_79_U2331 ( .A1(u5_mult_79_ab_11__20_), .A2(
        u5_mult_79_CARRYB_10__20_), .ZN(u5_mult_79_n1146) );
  NAND3_X2 u5_mult_79_U2330 ( .A1(u5_mult_79_n1142), .A2(u5_mult_79_n1143), 
        .A3(u5_mult_79_n1144), .ZN(u5_mult_79_CARRYB_10__20_) );
  NAND2_X2 u5_mult_79_U2329 ( .A1(u5_mult_79_ab_10__20_), .A2(
        u5_mult_79_SUMB_9__21_), .ZN(u5_mult_79_n1144) );
  NAND2_X1 u5_mult_79_U2328 ( .A1(u5_mult_79_SUMB_9__21_), .A2(
        u5_mult_79_CARRYB_9__20_), .ZN(u5_mult_79_n1143) );
  NAND2_X1 u5_mult_79_U2327 ( .A1(u5_mult_79_CARRYB_9__20_), .A2(
        u5_mult_79_ab_10__20_), .ZN(u5_mult_79_n1142) );
  NAND3_X2 u5_mult_79_U2326 ( .A1(u5_mult_79_n1139), .A2(u5_mult_79_n1140), 
        .A3(u5_mult_79_n1141), .ZN(u5_mult_79_CARRYB_18__14_) );
  NAND2_X2 u5_mult_79_U2325 ( .A1(u5_mult_79_CARRYB_16__15_), .A2(
        u5_mult_79_SUMB_16__16_), .ZN(u5_mult_79_n1138) );
  NAND2_X2 u5_mult_79_U2324 ( .A1(u5_mult_79_ab_17__15_), .A2(
        u5_mult_79_SUMB_16__16_), .ZN(u5_mult_79_n1137) );
  NAND2_X2 u5_mult_79_U2323 ( .A1(u5_mult_79_ab_17__11_), .A2(
        u5_mult_79_CARRYB_16__11_), .ZN(u5_mult_79_n1204) );
  XNOR2_X2 u5_mult_79_U2322 ( .A(u5_mult_79_CARRYB_21__4_), .B(
        u5_mult_79_ab_22__4_), .ZN(u5_mult_79_n1131) );
  XNOR2_X2 u5_mult_79_U2321 ( .A(u5_mult_79_n1131), .B(u5_mult_79_SUMB_21__5_), 
        .ZN(u5_mult_79_SUMB_22__4_) );
  NAND2_X1 u5_mult_79_U2320 ( .A1(u5_mult_79_ab_5__21_), .A2(
        u5_mult_79_CARRYB_4__21_), .ZN(u5_mult_79_n1553) );
  CLKBUF_X3 u5_mult_79_U2319 ( .A(u5_mult_79_CARRYB_16__5_), .Z(
        u5_mult_79_n1130) );
  NAND3_X2 u5_mult_79_U2318 ( .A1(u5_mult_79_n1127), .A2(u5_mult_79_n1128), 
        .A3(u5_mult_79_n1129), .ZN(u5_mult_79_CARRYB_7__11_) );
  NAND2_X1 u5_mult_79_U2317 ( .A1(u5_mult_79_CARRYB_6__11_), .A2(
        u5_mult_79_SUMB_6__12_), .ZN(u5_mult_79_n1129) );
  NAND2_X1 u5_mult_79_U2316 ( .A1(u5_mult_79_ab_7__11_), .A2(
        u5_mult_79_SUMB_6__12_), .ZN(u5_mult_79_n1128) );
  NAND2_X1 u5_mult_79_U2315 ( .A1(u5_mult_79_ab_7__11_), .A2(
        u5_mult_79_CARRYB_6__11_), .ZN(u5_mult_79_n1127) );
  NAND2_X2 u5_mult_79_U2314 ( .A1(u5_mult_79_SUMB_5__13_), .A2(
        u5_mult_79_CARRYB_5__12_), .ZN(u5_mult_79_n1126) );
  NAND2_X2 u5_mult_79_U2313 ( .A1(u5_mult_79_SUMB_5__13_), .A2(
        u5_mult_79_ab_6__12_), .ZN(u5_mult_79_n1125) );
  XOR2_X2 u5_mult_79_U2312 ( .A(u5_mult_79_n1123), .B(u5_mult_79_SUMB_6__12_), 
        .Z(u5_mult_79_SUMB_7__11_) );
  NAND2_X2 u5_mult_79_U2311 ( .A1(u5_mult_79_CARRYB_3__21_), .A2(
        u5_mult_79_n284), .ZN(u5_mult_79_n1619) );
  NAND2_X1 u5_mult_79_U2310 ( .A1(u5_mult_79_ab_5__16_), .A2(
        u5_mult_79_CARRYB_4__16_), .ZN(u5_mult_79_n1534) );
  XNOR2_X2 u5_mult_79_U2309 ( .A(u5_mult_79_ab_4__17_), .B(
        u5_mult_79_CARRYB_3__17_), .ZN(u5_mult_79_n1120) );
  XNOR2_X2 u5_mult_79_U2308 ( .A(u5_mult_79_n1120), .B(u5_mult_79_SUMB_3__18_), 
        .ZN(u5_mult_79_SUMB_4__17_) );
  NAND2_X2 u5_mult_79_U2307 ( .A1(u5_mult_79_ab_7__19_), .A2(
        u5_mult_79_SUMB_6__20_), .ZN(u5_mult_79_n1574) );
  XNOR2_X2 u5_mult_79_U2306 ( .A(u5_mult_79_n1118), .B(
        u5_mult_79_CARRYB_10__20_), .ZN(u5_mult_79_SUMB_11__20_) );
  NOR2_X1 u5_mult_79_U2305 ( .A1(u5_mult_79_n1818), .A2(u5_mult_79_n1752), 
        .ZN(u5_mult_79_ab_12__5_) );
  NOR2_X1 u5_mult_79_U2304 ( .A1(u5_mult_79_n1818), .A2(u5_mult_79_n1749), 
        .ZN(u5_mult_79_ab_11__5_) );
  NAND2_X2 u5_mult_79_U2303 ( .A1(u5_mult_79_n385), .A2(u5_mult_79_ab_12__5_), 
        .ZN(u5_mult_79_n1116) );
  NAND2_X1 u5_mult_79_U2302 ( .A1(u5_mult_79_ab_11__5_), .A2(
        u5_mult_79_CARRYB_10__5_), .ZN(u5_mult_79_n1114) );
  NAND3_X4 u5_mult_79_U2301 ( .A1(u5_mult_79_n1505), .A2(u5_mult_79_n1506), 
        .A3(u5_mult_79_n1507), .ZN(u5_mult_79_CARRYB_22__2_) );
  NAND3_X2 u5_mult_79_U2300 ( .A1(u5_mult_79_n1109), .A2(u5_mult_79_n1110), 
        .A3(u5_mult_79_n1111), .ZN(u5_mult_79_CARRYB_12__6_) );
  NAND2_X1 u5_mult_79_U2299 ( .A1(u5_mult_79_CARRYB_11__6_), .A2(
        u5_mult_79_ab_12__6_), .ZN(u5_mult_79_n1109) );
  NAND2_X2 u5_mult_79_U2298 ( .A1(u5_mult_79_ab_11__7_), .A2(
        u5_mult_79_SUMB_10__8_), .ZN(u5_mult_79_n1107) );
  NAND2_X1 u5_mult_79_U2297 ( .A1(u5_mult_79_ab_11__7_), .A2(
        u5_mult_79_CARRYB_10__7_), .ZN(u5_mult_79_n1106) );
  NOR2_X1 u5_mult_79_U2296 ( .A1(u5_mult_79_n1805), .A2(u5_mult_79_n1737), 
        .ZN(u5_mult_79_ab_7__9_) );
  NOR2_X1 u5_mult_79_U2295 ( .A1(u5_mult_79_n1812), .A2(u5_mult_79_n1752), 
        .ZN(u5_mult_79_ab_12__7_) );
  NAND3_X2 u5_mult_79_U2294 ( .A1(u5_mult_79_n1103), .A2(u5_mult_79_n1104), 
        .A3(u5_mult_79_n1105), .ZN(u5_mult_79_CARRYB_7__9_) );
  NAND2_X1 u5_mult_79_U2293 ( .A1(u5_mult_79_ab_7__9_), .A2(
        u5_mult_79_CARRYB_6__9_), .ZN(u5_mult_79_n1105) );
  NAND2_X2 u5_mult_79_U2292 ( .A1(u5_mult_79_ab_7__9_), .A2(
        u5_mult_79_SUMB_6__10_), .ZN(u5_mult_79_n1104) );
  NAND2_X1 u5_mult_79_U2291 ( .A1(u5_mult_79_CARRYB_6__9_), .A2(
        u5_mult_79_SUMB_6__10_), .ZN(u5_mult_79_n1103) );
  NAND3_X2 u5_mult_79_U2290 ( .A1(u5_mult_79_n1100), .A2(u5_mult_79_n1101), 
        .A3(u5_mult_79_n1102), .ZN(u5_mult_79_CARRYB_14__5_) );
  NAND2_X1 u5_mult_79_U2289 ( .A1(u5_mult_79_CARRYB_13__5_), .A2(
        u5_mult_79_SUMB_13__6_), .ZN(u5_mult_79_n1102) );
  NAND2_X1 u5_mult_79_U2288 ( .A1(u5_mult_79_ab_14__5_), .A2(
        u5_mult_79_SUMB_13__6_), .ZN(u5_mult_79_n1101) );
  NAND2_X1 u5_mult_79_U2287 ( .A1(u5_mult_79_ab_14__5_), .A2(
        u5_mult_79_CARRYB_13__5_), .ZN(u5_mult_79_n1100) );
  NAND3_X2 u5_mult_79_U2286 ( .A1(u5_mult_79_n1097), .A2(u5_mult_79_n1098), 
        .A3(u5_mult_79_n1099), .ZN(u5_mult_79_CARRYB_13__6_) );
  NAND2_X2 u5_mult_79_U2285 ( .A1(u5_mult_79_SUMB_12__7_), .A2(
        u5_mult_79_CARRYB_12__6_), .ZN(u5_mult_79_n1099) );
  NAND2_X2 u5_mult_79_U2284 ( .A1(u5_mult_79_ab_13__6_), .A2(
        u5_mult_79_SUMB_12__7_), .ZN(u5_mult_79_n1098) );
  NAND2_X1 u5_mult_79_U2283 ( .A1(u5_mult_79_ab_13__6_), .A2(
        u5_mult_79_CARRYB_12__6_), .ZN(u5_mult_79_n1097) );
  NAND3_X2 u5_mult_79_U2282 ( .A1(u5_mult_79_n1095), .A2(u5_mult_79_n1094), 
        .A3(u5_mult_79_n1096), .ZN(u5_mult_79_CARRYB_12__7_) );
  NAND2_X2 u5_mult_79_U2281 ( .A1(u5_mult_79_ab_11__13_), .A2(
        u5_mult_79_CARRYB_10__13_), .ZN(u5_mult_79_n1418) );
  NOR2_X2 u5_mult_79_U2280 ( .A1(u5_mult_79_n1868), .A2(u5_mult_79_n1747), 
        .ZN(u5_mult_79_ab_10__13_) );
  NOR2_X1 u5_mult_79_U2279 ( .A1(u5_mult_79_n1812), .A2(u5_mult_79_n1775), 
        .ZN(u5_mult_79_ab_20__7_) );
  NOR2_X1 u5_mult_79_U2278 ( .A1(u5_mult_79_n1801), .A2(u5_mult_79_n1756), 
        .ZN(u5_mult_79_ab_13__11_) );
  NAND3_X4 u5_mult_79_U2277 ( .A1(u5_mult_79_n1091), .A2(u5_mult_79_n1092), 
        .A3(u5_mult_79_n1093), .ZN(u5_mult_79_CARRYB_10__13_) );
  NAND2_X2 u5_mult_79_U2276 ( .A1(u5_mult_79_ab_10__13_), .A2(
        u5_mult_79_SUMB_9__14_), .ZN(u5_mult_79_n1092) );
  NAND2_X2 u5_mult_79_U2275 ( .A1(u5_mult_79_CARRYB_9__13_), .A2(
        u5_mult_79_SUMB_9__14_), .ZN(u5_mult_79_n1091) );
  NAND3_X2 u5_mult_79_U2274 ( .A1(u5_mult_79_n1088), .A2(u5_mult_79_n1089), 
        .A3(u5_mult_79_n1090), .ZN(u5_mult_79_CARRYB_20__7_) );
  NAND2_X1 u5_mult_79_U2273 ( .A1(u5_mult_79_ab_20__7_), .A2(
        u5_mult_79_CARRYB_19__7_), .ZN(u5_mult_79_n1090) );
  NAND2_X1 u5_mult_79_U2272 ( .A1(u5_mult_79_CARRYB_19__7_), .A2(
        u5_mult_79_SUMB_19__8_), .ZN(u5_mult_79_n1088) );
  NAND3_X2 u5_mult_79_U2271 ( .A1(u5_mult_79_n1085), .A2(u5_mult_79_n1086), 
        .A3(u5_mult_79_n1087), .ZN(u5_mult_79_CARRYB_13__11_) );
  NAND2_X1 u5_mult_79_U2270 ( .A1(u5_mult_79_ab_13__11_), .A2(
        u5_mult_79_CARRYB_12__11_), .ZN(u5_mult_79_n1087) );
  NAND2_X2 u5_mult_79_U2269 ( .A1(u5_mult_79_ab_13__11_), .A2(
        u5_mult_79_SUMB_12__12_), .ZN(u5_mult_79_n1086) );
  NAND2_X4 u5_mult_79_U2268 ( .A1(u5_mult_79_n623), .A2(u5_mult_79_ab_1__22_), 
        .ZN(u5_mult_79_n1716) );
  XNOR2_X2 u5_mult_79_U2267 ( .A(u5_mult_79_n1083), .B(u5_mult_79_n21), .ZN(
        u5_mult_79_SUMB_8__17_) );
  NOR2_X4 u5_mult_79_U2266 ( .A1(u5_mult_79_n1831), .A2(u5_mult_79_n1722), 
        .ZN(u5_mult_79_ab_2__23_) );
  NAND2_X2 u5_mult_79_U2265 ( .A1(u5_mult_79_ab_20__2_), .A2(
        u5_mult_79_CARRYB_19__2_), .ZN(u5_mult_79_n1262) );
  XOR2_X2 u5_mult_79_U2264 ( .A(u5_mult_79_ab_8__18_), .B(
        u5_mult_79_CARRYB_7__18_), .Z(u5_mult_79_n1368) );
  NAND3_X4 u5_mult_79_U2263 ( .A1(u5_mult_79_n1206), .A2(u5_mult_79_n1207), 
        .A3(u5_mult_79_n1208), .ZN(u5_mult_79_CARRYB_8__16_) );
  NOR2_X1 u5_mult_79_U2262 ( .A1(u5_mult_79_n1783), .A2(u5_mult_79_n1750), 
        .ZN(u5_mult_79_ab_11__21_) );
  NOR2_X1 u5_mult_79_U2261 ( .A1(u5_mult_79_n1783), .A2(u5_mult_79_n1753), 
        .ZN(u5_mult_79_ab_12__21_) );
  NAND3_X2 u5_mult_79_U2260 ( .A1(u5_mult_79_n1080), .A2(u5_mult_79_n1081), 
        .A3(u5_mult_79_n1082), .ZN(u5_mult_79_CARRYB_11__21_) );
  NAND2_X1 u5_mult_79_U2259 ( .A1(u5_mult_79_ab_11__21_), .A2(
        u5_mult_79_SUMB_10__22_), .ZN(u5_mult_79_n1082) );
  NAND3_X2 u5_mult_79_U2258 ( .A1(u5_mult_79_n1077), .A2(u5_mult_79_n1078), 
        .A3(u5_mult_79_n1079), .ZN(u5_mult_79_CARRYB_12__21_) );
  NAND3_X2 u5_mult_79_U2257 ( .A1(u5_mult_79_n1074), .A2(u5_mult_79_n1075), 
        .A3(u5_mult_79_n1076), .ZN(u5_mult_79_CARRYB_15__19_) );
  NAND2_X2 u5_mult_79_U2256 ( .A1(u5_mult_79_ab_15__19_), .A2(
        u5_mult_79_SUMB_14__20_), .ZN(u5_mult_79_n1075) );
  NAND2_X2 u5_mult_79_U2255 ( .A1(u5_mult_79_ab_14__20_), .A2(
        u5_mult_79_SUMB_13__21_), .ZN(u5_mult_79_n1072) );
  XOR2_X2 u5_mult_79_U2254 ( .A(u5_mult_79_n1070), .B(u5_mult_79_SUMB_14__20_), 
        .Z(u5_mult_79_SUMB_15__19_) );
  NAND3_X2 u5_mult_79_U2253 ( .A1(u5_mult_79_n1343), .A2(u5_mult_79_n1344), 
        .A3(u5_mult_79_n1345), .ZN(u5_mult_79_CARRYB_5__13_) );
  XNOR2_X2 u5_mult_79_U2252 ( .A(u5_mult_79_CARRYB_2__13_), .B(
        u5_mult_79_ab_3__13_), .ZN(u5_mult_79_n1068) );
  XNOR2_X2 u5_mult_79_U2251 ( .A(u5_mult_79_n1068), .B(u5_mult_79_SUMB_2__14_), 
        .ZN(u5_mult_79_SUMB_3__13_) );
  NOR2_X1 u5_mult_79_U2250 ( .A1(u5_mult_79_n1783), .A2(u5_mult_79_n1738), 
        .ZN(u5_mult_79_ab_7__21_) );
  NOR2_X2 u5_mult_79_U2249 ( .A1(u5_mult_79_n1785), .A2(u5_mult_79_n1756), 
        .ZN(u5_mult_79_ab_13__19_) );
  NAND2_X1 u5_mult_79_U2248 ( .A1(u5_mult_79_ab_7__21_), .A2(
        u5_mult_79_SUMB_6__22_), .ZN(u5_mult_79_n1067) );
  NAND2_X2 u5_mult_79_U2247 ( .A1(u5_mult_79_CARRYB_6__21_), .A2(
        u5_mult_79_ab_7__21_), .ZN(u5_mult_79_n1066) );
  XOR2_X2 u5_mult_79_U2246 ( .A(u5_mult_79_CARRYB_6__21_), .B(u5_mult_79_n1064), .Z(u5_mult_79_SUMB_7__21_) );
  NAND3_X2 u5_mult_79_U2245 ( .A1(u5_mult_79_n1061), .A2(u5_mult_79_n1062), 
        .A3(u5_mult_79_n1063), .ZN(u5_mult_79_CARRYB_13__19_) );
  NAND2_X1 u5_mult_79_U2244 ( .A1(u5_mult_79_ab_13__19_), .A2(
        u5_mult_79_SUMB_12__20_), .ZN(u5_mult_79_n1063) );
  NAND2_X2 u5_mult_79_U2243 ( .A1(u5_mult_79_ab_13__19_), .A2(
        u5_mult_79_CARRYB_12__19_), .ZN(u5_mult_79_n1062) );
  NAND3_X2 u5_mult_79_U2242 ( .A1(u5_mult_79_n1058), .A2(u5_mult_79_n1059), 
        .A3(u5_mult_79_n1060), .ZN(u5_mult_79_CARRYB_23__11_) );
  NAND2_X1 u5_mult_79_U2241 ( .A1(u5_mult_79_CARRYB_22__11_), .A2(
        u5_mult_79_SUMB_22__12_), .ZN(u5_mult_79_n1060) );
  NAND2_X1 u5_mult_79_U2240 ( .A1(u5_mult_79_ab_23__11_), .A2(
        u5_mult_79_SUMB_22__12_), .ZN(u5_mult_79_n1059) );
  NAND2_X1 u5_mult_79_U2239 ( .A1(u5_mult_79_ab_23__11_), .A2(
        u5_mult_79_CARRYB_22__11_), .ZN(u5_mult_79_n1058) );
  NAND3_X4 u5_mult_79_U2238 ( .A1(u5_mult_79_n1055), .A2(u5_mult_79_n1056), 
        .A3(u5_mult_79_n1057), .ZN(u5_mult_79_CARRYB_22__12_) );
  NAND2_X2 u5_mult_79_U2237 ( .A1(u5_mult_79_SUMB_21__13_), .A2(
        u5_mult_79_CARRYB_21__12_), .ZN(u5_mult_79_n1057) );
  NAND2_X2 u5_mult_79_U2236 ( .A1(u5_mult_79_SUMB_21__13_), .A2(
        u5_mult_79_ab_22__12_), .ZN(u5_mult_79_n1056) );
  NAND2_X2 u5_mult_79_U2235 ( .A1(u5_mult_79_CARRYB_21__1_), .A2(
        u5_mult_79_SUMB_21__2_), .ZN(u5_mult_79_n1175) );
  NAND2_X2 u5_mult_79_U2234 ( .A1(u5_mult_79_ab_15__11_), .A2(
        u5_mult_79_SUMB_14__12_), .ZN(u5_mult_79_n1490) );
  XNOR2_X2 u5_mult_79_U2233 ( .A(u5_mult_79_CARRYB_16__5_), .B(
        u5_mult_79_ab_17__5_), .ZN(u5_mult_79_n1053) );
  XNOR2_X2 u5_mult_79_U2232 ( .A(u5_mult_79_SUMB_16__6_), .B(u5_mult_79_n1053), 
        .ZN(u5_mult_79_SUMB_17__5_) );
  XNOR2_X1 u5_mult_79_U2231 ( .A(u5_mult_79_SUMB_23__2_), .B(
        u5_mult_79_CARRYB_23__1_), .ZN(u5_mult_79_n1647) );
  NAND3_X2 u5_mult_79_U2230 ( .A1(u5_mult_79_n1639), .A2(u5_mult_79_n1640), 
        .A3(u5_mult_79_n1641), .ZN(u5_mult_79_CARRYB_18__8_) );
  NAND2_X2 u5_mult_79_U2229 ( .A1(u5_mult_79_CARRYB_14__11_), .A2(
        u5_mult_79_SUMB_14__12_), .ZN(u5_mult_79_n1491) );
  XNOR2_X2 u5_mult_79_U2228 ( .A(u5_mult_79_SUMB_2__16_), .B(
        u5_mult_79_ab_3__15_), .ZN(u5_mult_79_n1266) );
  NAND2_X2 u5_mult_79_U2227 ( .A1(u5_mult_79_CARRYB_14__8_), .A2(
        u5_mult_79_SUMB_14__9_), .ZN(u5_mult_79_n1479) );
  NAND2_X2 u5_mult_79_U2226 ( .A1(u5_mult_79_CARRYB_17__5_), .A2(
        u5_mult_79_SUMB_17__6_), .ZN(u5_mult_79_n1199) );
  NAND2_X2 u5_mult_79_U2225 ( .A1(u5_mult_79_ab_4__21_), .A2(u5_mult_79_n284), 
        .ZN(u5_mult_79_n1621) );
  NOR2_X2 u5_mult_79_U2224 ( .A1(u5_mult_79_n1867), .A2(u5_mult_79_n1778), 
        .ZN(u5_mult_79_ab_21__14_) );
  NOR2_X2 u5_mult_79_U2223 ( .A1(u5_mult_79_n1867), .A2(u5_mult_79_n1776), 
        .ZN(u5_mult_79_ab_20__14_) );
  NOR2_X2 u5_mult_79_U2222 ( .A1(u5_mult_79_n1867), .A2(u5_mult_79_n1773), 
        .ZN(u5_mult_79_ab_19__14_) );
  NOR2_X2 u5_mult_79_U2221 ( .A1(u5_mult_79_n1867), .A2(u5_mult_79_n1768), 
        .ZN(u5_mult_79_ab_17__14_) );
  NOR2_X2 u5_mult_79_U2220 ( .A1(u5_mult_79_n1867), .A2(u5_mult_79_n1765), 
        .ZN(u5_mult_79_ab_16__14_) );
  NOR2_X2 u5_mult_79_U2219 ( .A1(u5_mult_79_n1867), .A2(u5_mult_79_n1756), 
        .ZN(u5_mult_79_ab_13__14_) );
  NOR2_X2 u5_mult_79_U2218 ( .A1(u5_mult_79_n1867), .A2(u5_mult_79_n1753), 
        .ZN(u5_mult_79_ab_12__14_) );
  NOR2_X2 u5_mult_79_U2217 ( .A1(u5_mult_79_n1867), .A2(u5_mult_79_n1750), 
        .ZN(u5_mult_79_ab_11__14_) );
  NOR2_X2 u5_mult_79_U2216 ( .A1(u5_mult_79_n1867), .A2(u5_mult_79_n1747), 
        .ZN(u5_mult_79_ab_10__14_) );
  NOR2_X2 u5_mult_79_U2215 ( .A1(u5_mult_79_n1867), .A2(u5_mult_79_n1732), 
        .ZN(u5_mult_79_ab_5__14_) );
  NOR2_X2 u5_mult_79_U2214 ( .A1(u5_mult_79_n1867), .A2(u5_mult_79_n1859), 
        .ZN(u5_mult_79_ab_22__14_) );
  NOR2_X2 u5_mult_79_U2213 ( .A1(u5_mult_79_n1879), .A2(u5_mult_79_n1867), 
        .ZN(u5_mult_79_ab_23__14_) );
  XNOR2_X2 u5_mult_79_U2212 ( .A(u5_mult_79_ab_15__11_), .B(
        u5_mult_79_CARRYB_14__11_), .ZN(u5_mult_79_n1052) );
  XNOR2_X2 u5_mult_79_U2211 ( .A(u5_mult_79_n1052), .B(u5_mult_79_SUMB_14__12_), .ZN(u5_mult_79_SUMB_15__11_) );
  NAND2_X2 u5_mult_79_U2210 ( .A1(u5_mult_79_ab_15__8_), .A2(
        u5_mult_79_SUMB_14__9_), .ZN(u5_mult_79_n1478) );
  NAND3_X4 u5_mult_79_U2209 ( .A1(u5_mult_79_n1477), .A2(u5_mult_79_n1478), 
        .A3(u5_mult_79_n1479), .ZN(u5_mult_79_CARRYB_15__8_) );
  XNOR2_X2 u5_mult_79_U2208 ( .A(u5_mult_79_ab_7__10_), .B(
        u5_mult_79_CARRYB_6__10_), .ZN(u5_mult_79_n1051) );
  XNOR2_X2 u5_mult_79_U2207 ( .A(u5_mult_79_n1051), .B(u5_mult_79_SUMB_6__11_), 
        .ZN(u5_mult_79_SUMB_7__10_) );
  XNOR2_X2 u5_mult_79_U2206 ( .A(u5_mult_79_n1508), .B(u5_mult_79_n1050), .ZN(
        u5_mult_79_SUMB_23__2_) );
  NAND2_X4 u5_mult_79_U2205 ( .A1(u5_mult_79_n1218), .A2(u5_mult_79_n1219), 
        .ZN(u5_mult_79_SUMB_4__19_) );
  INV_X4 u5_mult_79_U2204 ( .A(u5_mult_79_n1544), .ZN(u5_mult_79_n1216) );
  NAND2_X2 u5_mult_79_U2203 ( .A1(u5_mult_79_ab_8__17_), .A2(
        u5_mult_79_CARRYB_7__17_), .ZN(u5_mult_79_n1278) );
  NOR2_X4 u5_mult_79_U2202 ( .A1(u5_mult_79_n1793), .A2(u5_mult_79_n1723), 
        .ZN(u5_mult_79_ab_2__16_) );
  XNOR2_X2 u5_mult_79_U2201 ( .A(u5_mult_79_SUMB_15__6_), .B(u5_mult_79_n1132), 
        .ZN(u5_mult_79_SUMB_16__5_) );
  NOR2_X2 u5_mult_79_U2200 ( .A1(u5_mult_79_n1796), .A2(u5_mult_79_n1759), 
        .ZN(u5_mult_79_ab_14__15_) );
  NOR2_X1 u5_mult_79_U2199 ( .A1(u5_mult_79_n1803), .A2(u5_mult_79_n1857), 
        .ZN(u5_mult_79_ab_21__10_) );
  NAND2_X2 u5_mult_79_U2198 ( .A1(u5_mult_79_ab_19__12_), .A2(
        u5_mult_79_CARRYB_18__12_), .ZN(u5_mult_79_n1220) );
  NOR2_X2 u5_mult_79_U2197 ( .A1(u5_mult_79_n1799), .A2(u5_mult_79_n1771), 
        .ZN(u5_mult_79_ab_18__12_) );
  NOR2_X1 u5_mult_79_U2196 ( .A1(u5_mult_79_n1829), .A2(u5_mult_79_n1808), 
        .ZN(u5_mult_79_ab_23__8_) );
  NOR2_X1 u5_mult_79_U2195 ( .A1(u5_mult_79_n1796), .A2(u5_mult_79_n1750), 
        .ZN(u5_mult_79_ab_11__15_) );
  NAND3_X4 u5_mult_79_U2194 ( .A1(u5_mult_79_n1047), .A2(u5_mult_79_n1048), 
        .A3(u5_mult_79_n1049), .ZN(u5_mult_79_CARRYB_14__15_) );
  NAND2_X2 u5_mult_79_U2193 ( .A1(u5_mult_79_SUMB_13__16_), .A2(
        u5_mult_79_ab_14__15_), .ZN(u5_mult_79_n1048) );
  NAND2_X1 u5_mult_79_U2192 ( .A1(u5_mult_79_ab_21__10_), .A2(
        u5_mult_79_CARRYB_20__10_), .ZN(u5_mult_79_n1046) );
  NAND2_X2 u5_mult_79_U2191 ( .A1(u5_mult_79_ab_21__10_), .A2(
        u5_mult_79_SUMB_20__11_), .ZN(u5_mult_79_n1045) );
  NAND2_X1 u5_mult_79_U2190 ( .A1(u5_mult_79_ab_18__12_), .A2(
        u5_mult_79_CARRYB_17__12_), .ZN(u5_mult_79_n1043) );
  NAND3_X2 u5_mult_79_U2189 ( .A1(u5_mult_79_n1038), .A2(u5_mult_79_n1039), 
        .A3(u5_mult_79_n1040), .ZN(u5_mult_79_CARRYB_23__8_) );
  NAND2_X1 u5_mult_79_U2188 ( .A1(u5_mult_79_ab_23__8_), .A2(
        u5_mult_79_CARRYB_22__8_), .ZN(u5_mult_79_n1040) );
  NAND2_X1 u5_mult_79_U2187 ( .A1(u5_mult_79_ab_23__8_), .A2(
        u5_mult_79_SUMB_22__9_), .ZN(u5_mult_79_n1039) );
  NAND2_X1 u5_mult_79_U2186 ( .A1(u5_mult_79_CARRYB_22__8_), .A2(
        u5_mult_79_SUMB_22__9_), .ZN(u5_mult_79_n1038) );
  NAND3_X2 u5_mult_79_U2185 ( .A1(u5_mult_79_n1035), .A2(u5_mult_79_n1036), 
        .A3(u5_mult_79_n1037), .ZN(u5_mult_79_CARRYB_11__15_) );
  NAND2_X1 u5_mult_79_U2184 ( .A1(u5_mult_79_ab_11__15_), .A2(
        u5_mult_79_CARRYB_10__15_), .ZN(u5_mult_79_n1037) );
  NAND2_X2 u5_mult_79_U2183 ( .A1(u5_mult_79_ab_11__15_), .A2(
        u5_mult_79_SUMB_10__16_), .ZN(u5_mult_79_n1036) );
  NAND2_X1 u5_mult_79_U2182 ( .A1(u5_mult_79_CARRYB_10__15_), .A2(
        u5_mult_79_SUMB_10__16_), .ZN(u5_mult_79_n1035) );
  XOR2_X2 u5_mult_79_U2181 ( .A(u5_mult_79_SUMB_10__16_), .B(u5_mult_79_n1034), 
        .Z(u5_mult_79_SUMB_11__15_) );
  XNOR2_X2 u5_mult_79_U2180 ( .A(u5_mult_79_n1033), .B(
        u5_mult_79_CARRYB_6__11_), .ZN(u5_mult_79_n1123) );
  NAND2_X2 u5_mult_79_U2179 ( .A1(u5_mult_79_n1212), .A2(u5_mult_79_n1213), 
        .ZN(u5_mult_79_n1215) );
  XNOR2_X2 u5_mult_79_U2178 ( .A(u5_mult_79_CARRYB_10__15_), .B(
        u5_mult_79_n1032), .ZN(u5_mult_79_n1034) );
  NAND2_X4 u5_mult_79_U2177 ( .A1(u5_mult_79_ab_22__2_), .A2(
        u5_mult_79_CARRYB_21__2_), .ZN(u5_mult_79_n1505) );
  NOR2_X2 u5_mult_79_U2176 ( .A1(u5_mult_79_n1826), .A2(u5_mult_79_n1778), 
        .ZN(u5_mult_79_ab_21__2_) );
  NOR2_X1 u5_mult_79_U2175 ( .A1(u5_mult_79_n1826), .A2(u5_mult_79_n1773), 
        .ZN(u5_mult_79_ab_19__2_) );
  NOR2_X2 u5_mult_79_U2174 ( .A1(u5_mult_79_n1811), .A2(u5_mult_79_n1737), 
        .ZN(u5_mult_79_ab_7__7_) );
  NAND3_X4 u5_mult_79_U2173 ( .A1(u5_mult_79_n1028), .A2(u5_mult_79_n1029), 
        .A3(u5_mult_79_n1030), .ZN(u5_mult_79_CARRYB_21__2_) );
  NAND2_X2 u5_mult_79_U2172 ( .A1(u5_mult_79_SUMB_20__3_), .A2(
        u5_mult_79_ab_21__2_), .ZN(u5_mult_79_n1029) );
  NAND2_X2 u5_mult_79_U2171 ( .A1(u5_mult_79_SUMB_20__3_), .A2(
        u5_mult_79_CARRYB_20__2_), .ZN(u5_mult_79_n1028) );
  NAND3_X4 u5_mult_79_U2170 ( .A1(u5_mult_79_n1025), .A2(u5_mult_79_n1026), 
        .A3(u5_mult_79_n1027), .ZN(u5_mult_79_CARRYB_19__2_) );
  NAND2_X2 u5_mult_79_U2169 ( .A1(u5_mult_79_ab_19__2_), .A2(
        u5_mult_79_CARRYB_18__2_), .ZN(u5_mult_79_n1026) );
  NAND3_X2 u5_mult_79_U2168 ( .A1(u5_mult_79_n1022), .A2(u5_mult_79_n1023), 
        .A3(u5_mult_79_n1024), .ZN(u5_mult_79_CARRYB_10__4_) );
  NAND2_X1 u5_mult_79_U2167 ( .A1(u5_mult_79_CARRYB_9__4_), .A2(
        u5_mult_79_SUMB_9__5_), .ZN(u5_mult_79_n1024) );
  NAND2_X1 u5_mult_79_U2166 ( .A1(u5_mult_79_ab_10__4_), .A2(
        u5_mult_79_CARRYB_9__4_), .ZN(u5_mult_79_n1022) );
  NAND3_X2 u5_mult_79_U2165 ( .A1(u5_mult_79_n1019), .A2(u5_mult_79_n1020), 
        .A3(u5_mult_79_n1021), .ZN(u5_mult_79_CARRYB_9__5_) );
  NAND2_X2 u5_mult_79_U2164 ( .A1(u5_mult_79_ab_9__5_), .A2(
        u5_mult_79_SUMB_8__6_), .ZN(u5_mult_79_n1020) );
  NAND2_X1 u5_mult_79_U2163 ( .A1(u5_mult_79_ab_9__5_), .A2(
        u5_mult_79_CARRYB_8__5_), .ZN(u5_mult_79_n1019) );
  NAND2_X1 u5_mult_79_U2162 ( .A1(u5_mult_79_ab_7__7_), .A2(
        u5_mult_79_CARRYB_6__7_), .ZN(u5_mult_79_n1018) );
  NAND2_X2 u5_mult_79_U2161 ( .A1(u5_mult_79_CARRYB_15__9_), .A2(
        u5_mult_79_n448), .ZN(u5_mult_79_n1606) );
  XNOR2_X2 u5_mult_79_U2160 ( .A(u5_mult_79_ab_2__16_), .B(u5_mult_79_n1707), 
        .ZN(u5_mult_79_n1181) );
  NAND3_X2 u5_mult_79_U2159 ( .A1(u5_mult_79_n1145), .A2(u5_mult_79_n1146), 
        .A3(u5_mult_79_n1147), .ZN(u5_mult_79_CARRYB_11__20_) );
  XNOR2_X2 u5_mult_79_U2158 ( .A(u5_mult_79_n1014), .B(
        u5_mult_79_CARRYB_5__12_), .ZN(u5_mult_79_n1122) );
  XNOR2_X2 u5_mult_79_U2157 ( .A(u5_mult_79_CARRYB_6__19_), .B(
        u5_mult_79_n1451), .ZN(u5_mult_79_SUMB_7__19_) );
  NAND3_X2 u5_mult_79_U2156 ( .A1(u5_mult_79_n1491), .A2(u5_mult_79_n1490), 
        .A3(u5_mult_79_n1489), .ZN(u5_mult_79_CARRYB_15__11_) );
  BUF_X4 u5_mult_79_U2155 ( .A(u5_mult_79_CARRYB_7__18_), .Z(u5_mult_79_n1376)
         );
  NAND2_X1 u5_mult_79_U2154 ( .A1(u5_mult_79_CARRYB_15__10_), .A2(
        u5_mult_79_SUMB_15__11_), .ZN(u5_mult_79_n1494) );
  NOR2_X1 u5_mult_79_U2153 ( .A1(u5_mult_79_n1783), .A2(u5_mult_79_n1735), 
        .ZN(u5_mult_79_ab_6__21_) );
  NOR2_X1 u5_mult_79_U2152 ( .A1(u5_mult_79_n1783), .A2(u5_mult_79_n1741), 
        .ZN(u5_mult_79_ab_8__21_) );
  NOR2_X1 u5_mult_79_U2151 ( .A1(u5_mult_79_n1783), .A2(u5_mult_79_n1744), 
        .ZN(u5_mult_79_ab_9__21_) );
  NOR2_X1 u5_mult_79_U2150 ( .A1(u5_mult_79_n1783), .A2(u5_mult_79_n1747), 
        .ZN(u5_mult_79_ab_10__21_) );
  NOR2_X1 u5_mult_79_U2149 ( .A1(u5_mult_79_n1783), .A2(u5_mult_79_n1859), 
        .ZN(u5_mult_79_ab_22__21_) );
  NOR2_X1 u5_mult_79_U2148 ( .A1(u5_mult_79_n1829), .A2(u5_mult_79_n1783), 
        .ZN(u5_mult_79_ab_23__21_) );
  NOR2_X1 u5_mult_79_U2147 ( .A1(u5_mult_79_n1796), .A2(u5_mult_79_n1855), 
        .ZN(u5_mult_79_ab_19__15_) );
  NOR2_X1 u5_mult_79_U2146 ( .A1(u5_mult_79_n1796), .A2(u5_mult_79_n1771), 
        .ZN(u5_mult_79_ab_18__15_) );
  NAND3_X2 u5_mult_79_U2145 ( .A1(u5_mult_79_n1011), .A2(u5_mult_79_n1012), 
        .A3(u5_mult_79_n1013), .ZN(u5_mult_79_CARRYB_19__15_) );
  NAND2_X1 u5_mult_79_U2144 ( .A1(u5_mult_79_CARRYB_18__15_), .A2(
        u5_mult_79_ab_19__15_), .ZN(u5_mult_79_n1013) );
  NAND2_X2 u5_mult_79_U2143 ( .A1(u5_mult_79_ab_19__15_), .A2(
        u5_mult_79_SUMB_18__16_), .ZN(u5_mult_79_n1012) );
  XOR2_X2 u5_mult_79_U2142 ( .A(u5_mult_79_SUMB_18__16_), .B(u5_mult_79_n1010), 
        .Z(u5_mult_79_SUMB_19__15_) );
  NAND3_X2 u5_mult_79_U2141 ( .A1(u5_mult_79_n1007), .A2(u5_mult_79_n1008), 
        .A3(u5_mult_79_n1009), .ZN(u5_mult_79_CARRYB_18__15_) );
  NAND2_X1 u5_mult_79_U2140 ( .A1(u5_mult_79_ab_18__15_), .A2(
        u5_mult_79_CARRYB_17__15_), .ZN(u5_mult_79_n1009) );
  NAND2_X2 u5_mult_79_U2139 ( .A1(u5_mult_79_ab_18__15_), .A2(
        u5_mult_79_SUMB_17__16_), .ZN(u5_mult_79_n1008) );
  INV_X4 u5_mult_79_U2138 ( .A(n2986), .ZN(u5_mult_79_n1799) );
  CLKBUF_X3 u5_mult_79_U2137 ( .A(u5_mult_79_CARRYB_15__11_), .Z(
        u5_mult_79_n1268) );
  NOR2_X2 u5_mult_79_U2136 ( .A1(u5_mult_79_n1780), .A2(u5_mult_79_n1732), 
        .ZN(u5_mult_79_ab_5__22_) );
  NOR2_X1 u5_mult_79_U2135 ( .A1(u5_mult_79_n1780), .A2(u5_mult_79_n1729), 
        .ZN(u5_mult_79_ab_4__22_) );
  NOR2_X2 u5_mult_79_U2134 ( .A1(u5_mult_79_n1780), .A2(u5_mult_79_n1726), 
        .ZN(u5_mult_79_ab_3__22_) );
  NAND2_X2 u5_mult_79_U2133 ( .A1(u5_mult_79_n279), .A2(u5_mult_79_SUMB_3__17_), .ZN(u5_mult_79_n1290) );
  NAND3_X4 u5_mult_79_U2132 ( .A1(u5_mult_79_n1290), .A2(u5_mult_79_n1291), 
        .A3(u5_mult_79_n1292), .ZN(u5_mult_79_CARRYB_4__16_) );
  NOR2_X1 u5_mult_79_U2131 ( .A1(u5_mult_79_n1794), .A2(u5_mult_79_n1768), 
        .ZN(u5_mult_79_ab_17__16_) );
  NOR2_X1 u5_mult_79_U2130 ( .A1(u5_mult_79_n1794), .A2(u5_mult_79_n1765), 
        .ZN(u5_mult_79_ab_16__16_) );
  NAND2_X1 u5_mult_79_U2129 ( .A1(u5_mult_79_ab_17__16_), .A2(
        u5_mult_79_CARRYB_16__16_), .ZN(u5_mult_79_n1006) );
  NAND2_X2 u5_mult_79_U2128 ( .A1(u5_mult_79_ab_17__16_), .A2(
        u5_mult_79_SUMB_16__17_), .ZN(u5_mult_79_n1005) );
  NAND2_X1 u5_mult_79_U2127 ( .A1(u5_mult_79_ab_16__16_), .A2(
        u5_mult_79_CARRYB_15__16_), .ZN(u5_mult_79_n1003) );
  NAND2_X2 u5_mult_79_U2126 ( .A1(u5_mult_79_SUMB_14__7_), .A2(
        u5_mult_79_ab_15__6_), .ZN(u5_mult_79_n999) );
  NAND2_X2 u5_mult_79_U2125 ( .A1(u5_mult_79_n781), .A2(u5_mult_79_SUMB_13__8_), .ZN(u5_mult_79_n997) );
  NAND2_X2 u5_mult_79_U2124 ( .A1(u5_mult_79_ab_14__7_), .A2(
        u5_mult_79_SUMB_13__8_), .ZN(u5_mult_79_n996) );
  NAND2_X2 u5_mult_79_U2123 ( .A1(u5_mult_79_ab_14__7_), .A2(u5_mult_79_n781), 
        .ZN(u5_mult_79_n995) );
  NAND2_X1 u5_mult_79_U2122 ( .A1(u5_mult_79_ab_12__8_), .A2(
        u5_mult_79_CARRYB_11__8_), .ZN(u5_mult_79_n992) );
  NAND2_X2 u5_mult_79_U2121 ( .A1(u5_mult_79_CARRYB_10__9_), .A2(
        u5_mult_79_n433), .ZN(u5_mult_79_n991) );
  NOR2_X1 u5_mult_79_U2120 ( .A1(u5_mult_79_n1788), .A2(u5_mult_79_n1768), 
        .ZN(u5_mult_79_ab_17__18_) );
  NAND3_X2 u5_mult_79_U2119 ( .A1(u5_mult_79_n986), .A2(u5_mult_79_n987), .A3(
        u5_mult_79_n988), .ZN(u5_mult_79_CARRYB_17__18_) );
  NAND2_X1 u5_mult_79_U2118 ( .A1(u5_mult_79_ab_17__18_), .A2(
        u5_mult_79_SUMB_16__19_), .ZN(u5_mult_79_n988) );
  NAND2_X2 u5_mult_79_U2117 ( .A1(u5_mult_79_ab_17__18_), .A2(
        u5_mult_79_CARRYB_16__18_), .ZN(u5_mult_79_n987) );
  NAND2_X2 u5_mult_79_U2116 ( .A1(u5_mult_79_n373), .A2(
        u5_mult_79_CARRYB_16__18_), .ZN(u5_mult_79_n986) );
  NOR2_X2 u5_mult_79_U2115 ( .A1(u5_mult_79_n1791), .A2(u5_mult_79_n1753), 
        .ZN(u5_mult_79_ab_12__17_) );
  NOR2_X1 u5_mult_79_U2114 ( .A1(u5_mult_79_n1787), .A2(u5_mult_79_n1747), 
        .ZN(u5_mult_79_ab_10__18_) );
  NAND3_X2 u5_mult_79_U2113 ( .A1(u5_mult_79_n983), .A2(u5_mult_79_n984), .A3(
        u5_mult_79_n985), .ZN(u5_mult_79_CARRYB_12__17_) );
  NAND2_X1 u5_mult_79_U2112 ( .A1(u5_mult_79_ab_12__17_), .A2(
        u5_mult_79_CARRYB_11__17_), .ZN(u5_mult_79_n985) );
  NAND2_X1 u5_mult_79_U2111 ( .A1(u5_mult_79_CARRYB_11__17_), .A2(
        u5_mult_79_SUMB_11__18_), .ZN(u5_mult_79_n983) );
  XOR2_X2 u5_mult_79_U2110 ( .A(u5_mult_79_SUMB_11__18_), .B(u5_mult_79_n982), 
        .Z(u5_mult_79_SUMB_12__17_) );
  NAND3_X2 u5_mult_79_U2109 ( .A1(u5_mult_79_n979), .A2(u5_mult_79_n980), .A3(
        u5_mult_79_n981), .ZN(u5_mult_79_CARRYB_10__18_) );
  NAND2_X1 u5_mult_79_U2108 ( .A1(u5_mult_79_ab_10__18_), .A2(
        u5_mult_79_CARRYB_9__18_), .ZN(u5_mult_79_n981) );
  NAND2_X1 u5_mult_79_U2107 ( .A1(u5_mult_79_CARRYB_9__18_), .A2(
        u5_mult_79_SUMB_9__19_), .ZN(u5_mult_79_n979) );
  INV_X16 u5_mult_79_U2106 ( .A(u5_mult_79_n1784), .ZN(u5_mult_79_n1783) );
  INV_X32 u5_mult_79_U2105 ( .A(n3039), .ZN(u5_mult_79_n1338) );
  NOR2_X2 u5_mult_79_U2104 ( .A1(u5_mult_79_n1338), .A2(u5_mult_79_n1735), 
        .ZN(u5_mult_79_ab_6__20_) );
  NOR2_X4 u5_mult_79_U2103 ( .A1(u5_mult_79_n1338), .A2(u5_mult_79_n1732), 
        .ZN(u5_mult_79_ab_5__20_) );
  NOR2_X4 u5_mult_79_U2102 ( .A1(u5_mult_79_n1338), .A2(u5_mult_79_n1729), 
        .ZN(u5_mult_79_ab_4__20_) );
  XNOR2_X2 u5_mult_79_U2101 ( .A(u5_mult_79_CARRYB_9__12_), .B(
        u5_mult_79_ab_10__12_), .ZN(u5_mult_79_n978) );
  XNOR2_X2 u5_mult_79_U2100 ( .A(u5_mult_79_n978), .B(u5_mult_79_n311), .ZN(
        u5_mult_79_SUMB_10__12_) );
  NAND2_X2 u5_mult_79_U2099 ( .A1(u5_mult_79_CARRYB_15__4_), .A2(
        u5_mult_79_ab_16__4_), .ZN(u5_mult_79_n1501) );
  XNOR2_X2 u5_mult_79_U2098 ( .A(u5_mult_79_n1119), .B(u5_mult_79_SUMB_6__21_), 
        .ZN(u5_mult_79_SUMB_7__20_) );
  NAND3_X2 u5_mult_79_U2097 ( .A1(u5_mult_79_n1172), .A2(u5_mult_79_n1173), 
        .A3(u5_mult_79_n1174), .ZN(u5_mult_79_CARRYB_23__0_) );
  NAND2_X2 u5_mult_79_U2096 ( .A1(u5_mult_79_CARRYB_6__18_), .A2(
        u5_mult_79_SUMB_6__19_), .ZN(u5_mult_79_n1277) );
  NAND2_X2 u5_mult_79_U2095 ( .A1(u5_mult_79_ab_9__17_), .A2(
        u5_mult_79_SUMB_8__18_), .ZN(u5_mult_79_n1374) );
  XNOR2_X2 u5_mult_79_U2094 ( .A(u5_mult_79_CARRYB_11__6_), .B(
        u5_mult_79_ab_12__6_), .ZN(u5_mult_79_n977) );
  XNOR2_X2 u5_mult_79_U2093 ( .A(u5_mult_79_n977), .B(u5_mult_79_SUMB_11__7_), 
        .ZN(u5_mult_79_SUMB_12__6_) );
  XNOR2_X2 u5_mult_79_U2092 ( .A(u5_mult_79_ab_7__18_), .B(
        u5_mult_79_CARRYB_6__18_), .ZN(u5_mult_79_n976) );
  XNOR2_X2 u5_mult_79_U2091 ( .A(u5_mult_79_n976), .B(u5_mult_79_SUMB_6__19_), 
        .ZN(u5_mult_79_SUMB_7__18_) );
  NAND2_X2 u5_mult_79_U2090 ( .A1(u5_mult_79_ab_22__10_), .A2(
        u5_mult_79_SUMB_21__11_), .ZN(u5_mult_79_n1453) );
  NAND3_X2 u5_mult_79_U2089 ( .A1(u5_mult_79_n1603), .A2(u5_mult_79_n1604), 
        .A3(u5_mult_79_n1605), .ZN(u5_mult_79_CARRYB_4__20_) );
  NOR2_X1 u5_mult_79_U2088 ( .A1(u5_mult_79_n1867), .A2(u5_mult_79_n1741), 
        .ZN(u5_mult_79_ab_8__14_) );
  NOR2_X1 u5_mult_79_U2087 ( .A1(u5_mult_79_n1867), .A2(u5_mult_79_n1738), 
        .ZN(u5_mult_79_ab_7__14_) );
  NAND2_X2 u5_mult_79_U2086 ( .A1(u5_mult_79_ab_8__14_), .A2(
        u5_mult_79_SUMB_7__15_), .ZN(u5_mult_79_n974) );
  NAND2_X1 u5_mult_79_U2085 ( .A1(u5_mult_79_ab_7__14_), .A2(
        u5_mult_79_CARRYB_6__14_), .ZN(u5_mult_79_n972) );
  NAND2_X2 u5_mult_79_U2084 ( .A1(u5_mult_79_ab_7__14_), .A2(
        u5_mult_79_SUMB_6__15_), .ZN(u5_mult_79_n971) );
  NAND2_X2 u5_mult_79_U2083 ( .A1(u5_mult_79_CARRYB_20__3_), .A2(
        u5_mult_79_SUMB_20__4_), .ZN(u5_mult_79_n1635) );
  NOR2_X2 u5_mult_79_U2082 ( .A1(u5_mult_79_n1785), .A2(u5_mult_79_n1723), 
        .ZN(u5_mult_79_ab_2__19_) );
  NAND3_X2 u5_mult_79_U2081 ( .A1(u5_mult_79_n1534), .A2(u5_mult_79_n1535), 
        .A3(u5_mult_79_n1536), .ZN(u5_mult_79_CARRYB_5__16_) );
  XNOR2_X2 u5_mult_79_U2080 ( .A(u5_mult_79_n968), .B(u5_mult_79_CARRYB_4__16_), .ZN(u5_mult_79_n1533) );
  NAND2_X2 u5_mult_79_U2079 ( .A1(u5_mult_79_CARRYB_21__2_), .A2(
        u5_mult_79_n280), .ZN(u5_mult_79_n1507) );
  NAND2_X2 u5_mult_79_U2078 ( .A1(u5_mult_79_CARRYB_9__15_), .A2(
        u5_mult_79_SUMB_9__16_), .ZN(u5_mult_79_n1274) );
  XNOR2_X2 u5_mult_79_U2077 ( .A(u5_mult_79_ab_11__12_), .B(
        u5_mult_79_CARRYB_10__12_), .ZN(u5_mult_79_n967) );
  XNOR2_X2 u5_mult_79_U2076 ( .A(u5_mult_79_n967), .B(u5_mult_79_SUMB_10__13_), 
        .ZN(u5_mult_79_SUMB_11__12_) );
  XNOR2_X2 u5_mult_79_U2075 ( .A(u5_mult_79_CARRYB_11__8_), .B(
        u5_mult_79_ab_12__8_), .ZN(u5_mult_79_n966) );
  XNOR2_X2 u5_mult_79_U2074 ( .A(u5_mult_79_n966), .B(u5_mult_79_SUMB_11__9_), 
        .ZN(u5_mult_79_SUMB_12__8_) );
  NAND3_X4 u5_mult_79_U2073 ( .A1(u5_mult_79_n1465), .A2(u5_mult_79_n1466), 
        .A3(u5_mult_79_n1467), .ZN(u5_mult_79_CARRYB_12__9_) );
  INV_X8 u5_mult_79_U2072 ( .A(n2944), .ZN(u5_mult_79_n1869) );
  NAND2_X1 u5_mult_79_U2071 ( .A1(u5_mult_79_ab_22__7_), .A2(
        u5_mult_79_CARRYB_21__7_), .ZN(u5_mult_79_n962) );
  NAND3_X4 u5_mult_79_U2070 ( .A1(u5_mult_79_n959), .A2(u5_mult_79_n960), .A3(
        u5_mult_79_n961), .ZN(u5_mult_79_CARRYB_21__8_) );
  NAND2_X2 u5_mult_79_U2069 ( .A1(u5_mult_79_CARRYB_20__8_), .A2(
        u5_mult_79_SUMB_20__9_), .ZN(u5_mult_79_n961) );
  NAND2_X2 u5_mult_79_U2068 ( .A1(u5_mult_79_ab_21__8_), .A2(u5_mult_79_n367), 
        .ZN(u5_mult_79_n960) );
  XOR2_X2 u5_mult_79_U2067 ( .A(u5_mult_79_ab_21__8_), .B(
        u5_mult_79_CARRYB_20__8_), .Z(u5_mult_79_n958) );
  NAND2_X2 u5_mult_79_U2066 ( .A1(u5_mult_79_CARRYB_15__4_), .A2(
        u5_mult_79_SUMB_15__5_), .ZN(u5_mult_79_n1503) );
  XNOR2_X2 u5_mult_79_U2065 ( .A(u5_mult_79_CARRYB_13__9_), .B(
        u5_mult_79_ab_14__9_), .ZN(u5_mult_79_n957) );
  XNOR2_X2 u5_mult_79_U2064 ( .A(u5_mult_79_n286), .B(u5_mult_79_n957), .ZN(
        u5_mult_79_SUMB_14__9_) );
  NAND2_X1 u5_mult_79_U2063 ( .A1(u5_mult_79_CARRYB_21__11_), .A2(
        u5_mult_79_SUMB_21__12_), .ZN(u5_mult_79_n1308) );
  XNOR2_X2 u5_mult_79_U2062 ( .A(u5_mult_79_ab_22__7_), .B(
        u5_mult_79_CARRYB_21__7_), .ZN(u5_mult_79_n956) );
  XNOR2_X2 u5_mult_79_U2061 ( .A(u5_mult_79_n956), .B(u5_mult_79_SUMB_21__8_), 
        .ZN(u5_mult_79_SUMB_22__7_) );
  NAND3_X2 u5_mult_79_U2060 ( .A1(u5_mult_79_n954), .A2(u5_mult_79_n955), .A3(
        u5_mult_79_n953), .ZN(u5_mult_79_CARRYB_18__13_) );
  NAND2_X2 u5_mult_79_U2059 ( .A1(u5_mult_79_SUMB_17__14_), .A2(
        u5_mult_79_ab_18__13_), .ZN(u5_mult_79_n954) );
  NOR2_X1 u5_mult_79_U2058 ( .A1(u5_mult_79_n1834), .A2(u5_mult_79_n1758), 
        .ZN(u5_mult_79_ab_14__0_) );
  NOR2_X1 u5_mult_79_U2057 ( .A1(u5_mult_79_n1834), .A2(u5_mult_79_n1755), 
        .ZN(u5_mult_79_ab_13__0_) );
  NAND3_X2 u5_mult_79_U2056 ( .A1(u5_mult_79_n947), .A2(u5_mult_79_n948), .A3(
        u5_mult_79_n949), .ZN(u5_mult_79_CARRYB_14__0_) );
  NAND2_X1 u5_mult_79_U2055 ( .A1(u5_mult_79_ab_14__0_), .A2(
        u5_mult_79_CARRYB_13__0_), .ZN(u5_mult_79_n949) );
  NAND2_X2 u5_mult_79_U2054 ( .A1(u5_mult_79_ab_14__0_), .A2(
        u5_mult_79_SUMB_13__1_), .ZN(u5_mult_79_n948) );
  XOR2_X2 u5_mult_79_U2053 ( .A(u5_mult_79_SUMB_13__1_), .B(u5_mult_79_n946), 
        .Z(u5_N14) );
  XOR2_X2 u5_mult_79_U2052 ( .A(u5_mult_79_CARRYB_13__0_), .B(
        u5_mult_79_ab_14__0_), .Z(u5_mult_79_n946) );
  NAND3_X2 u5_mult_79_U2051 ( .A1(u5_mult_79_n943), .A2(u5_mult_79_n944), .A3(
        u5_mult_79_n945), .ZN(u5_mult_79_CARRYB_13__0_) );
  NAND2_X1 u5_mult_79_U2050 ( .A1(u5_mult_79_ab_13__0_), .A2(
        u5_mult_79_CARRYB_12__0_), .ZN(u5_mult_79_n945) );
  NAND2_X2 u5_mult_79_U2049 ( .A1(u5_mult_79_ab_13__0_), .A2(
        u5_mult_79_SUMB_12__1_), .ZN(u5_mult_79_n944) );
  NAND2_X1 u5_mult_79_U2048 ( .A1(u5_mult_79_CARRYB_12__0_), .A2(
        u5_mult_79_SUMB_12__1_), .ZN(u5_mult_79_n943) );
  XOR2_X2 u5_mult_79_U2047 ( .A(u5_mult_79_SUMB_12__1_), .B(u5_mult_79_n942), 
        .Z(u5_N13) );
  XOR2_X2 u5_mult_79_U2046 ( .A(u5_mult_79_CARRYB_12__0_), .B(
        u5_mult_79_ab_13__0_), .Z(u5_mult_79_n942) );
  NAND3_X2 u5_mult_79_U2045 ( .A1(u5_mult_79_n939), .A2(u5_mult_79_n940), .A3(
        u5_mult_79_n941), .ZN(u5_mult_79_CARRYB_17__0_) );
  NAND2_X2 u5_mult_79_U2044 ( .A1(u5_mult_79_CARRYB_16__0_), .A2(
        u5_mult_79_SUMB_16__1_), .ZN(u5_mult_79_n941) );
  NAND2_X2 u5_mult_79_U2043 ( .A1(u5_mult_79_ab_17__0_), .A2(
        u5_mult_79_CARRYB_16__0_), .ZN(u5_mult_79_n940) );
  NAND2_X2 u5_mult_79_U2042 ( .A1(u5_mult_79_ab_17__0_), .A2(
        u5_mult_79_SUMB_16__1_), .ZN(u5_mult_79_n939) );
  XOR2_X2 u5_mult_79_U2041 ( .A(u5_mult_79_n938), .B(u5_mult_79_CARRYB_16__0_), 
        .Z(u5_N17) );
  NAND3_X2 u5_mult_79_U2040 ( .A1(u5_mult_79_n935), .A2(u5_mult_79_n936), .A3(
        u5_mult_79_n937), .ZN(u5_mult_79_CARRYB_16__0_) );
  NAND2_X1 u5_mult_79_U2039 ( .A1(u5_mult_79_CARRYB_15__0_), .A2(
        u5_mult_79_SUMB_15__1_), .ZN(u5_mult_79_n937) );
  NAND2_X2 u5_mult_79_U2038 ( .A1(u5_mult_79_ab_16__0_), .A2(
        u5_mult_79_SUMB_15__1_), .ZN(u5_mult_79_n936) );
  NAND2_X1 u5_mult_79_U2037 ( .A1(u5_mult_79_ab_16__0_), .A2(
        u5_mult_79_CARRYB_15__0_), .ZN(u5_mult_79_n935) );
  XOR2_X2 u5_mult_79_U2036 ( .A(u5_mult_79_n934), .B(u5_mult_79_SUMB_15__1_), 
        .Z(u5_N16) );
  NOR2_X1 u5_mult_79_U2035 ( .A1(u5_mult_79_n1826), .A2(u5_mult_79_n1752), 
        .ZN(u5_mult_79_ab_12__2_) );
  NOR2_X1 u5_mult_79_U2034 ( .A1(u5_mult_79_n1826), .A2(u5_mult_79_n1749), 
        .ZN(u5_mult_79_ab_11__2_) );
  NOR2_X1 u5_mult_79_U2033 ( .A1(u5_mult_79_n1826), .A2(u5_mult_79_n1758), 
        .ZN(u5_mult_79_ab_14__2_) );
  NAND3_X2 u5_mult_79_U2032 ( .A1(u5_mult_79_n931), .A2(u5_mult_79_n932), .A3(
        u5_mult_79_n933), .ZN(u5_mult_79_CARRYB_12__2_) );
  NAND2_X2 u5_mult_79_U2031 ( .A1(u5_mult_79_ab_12__2_), .A2(
        u5_mult_79_SUMB_11__3_), .ZN(u5_mult_79_n932) );
  XOR2_X2 u5_mult_79_U2030 ( .A(u5_mult_79_SUMB_11__3_), .B(u5_mult_79_n930), 
        .Z(u5_mult_79_SUMB_12__2_) );
  XOR2_X2 u5_mult_79_U2029 ( .A(u5_mult_79_CARRYB_11__2_), .B(
        u5_mult_79_ab_12__2_), .Z(u5_mult_79_n930) );
  NAND3_X2 u5_mult_79_U2028 ( .A1(u5_mult_79_n927), .A2(u5_mult_79_n928), .A3(
        u5_mult_79_n929), .ZN(u5_mult_79_CARRYB_11__2_) );
  NAND2_X2 u5_mult_79_U2027 ( .A1(u5_mult_79_ab_11__2_), .A2(
        u5_mult_79_SUMB_10__3_), .ZN(u5_mult_79_n928) );
  NAND2_X1 u5_mult_79_U2026 ( .A1(u5_mult_79_CARRYB_10__2_), .A2(
        u5_mult_79_SUMB_10__3_), .ZN(u5_mult_79_n927) );
  NAND3_X2 u5_mult_79_U2025 ( .A1(u5_mult_79_n924), .A2(u5_mult_79_n925), .A3(
        u5_mult_79_n926), .ZN(u5_mult_79_CARRYB_14__2_) );
  NAND2_X2 u5_mult_79_U2024 ( .A1(u5_mult_79_SUMB_13__3_), .A2(
        u5_mult_79_ab_14__2_), .ZN(u5_mult_79_n925) );
  NOR2_X2 u5_mult_79_U2023 ( .A1(u5_mult_79_n1814), .A2(u5_mult_79_n1740), 
        .ZN(u5_mult_79_ab_8__6_) );
  NOR2_X1 u5_mult_79_U2022 ( .A1(u5_mult_79_n1814), .A2(u5_mult_79_n1737), 
        .ZN(u5_mult_79_ab_7__6_) );
  NOR2_X1 u5_mult_79_U2021 ( .A1(u5_mult_79_n1821), .A2(u5_mult_79_n1749), 
        .ZN(u5_mult_79_ab_11__4_) );
  NOR2_X2 u5_mult_79_U2020 ( .A1(u5_mult_79_n1817), .A2(u5_mult_79_n1746), 
        .ZN(u5_mult_79_ab_10__5_) );
  NAND2_X1 u5_mult_79_U2019 ( .A1(u5_mult_79_ab_8__6_), .A2(
        u5_mult_79_CARRYB_7__6_), .ZN(u5_mult_79_n923) );
  NAND3_X2 u5_mult_79_U2018 ( .A1(u5_mult_79_n918), .A2(u5_mult_79_n919), .A3(
        u5_mult_79_n920), .ZN(u5_mult_79_CARRYB_7__6_) );
  NAND2_X1 u5_mult_79_U2017 ( .A1(u5_mult_79_ab_7__6_), .A2(
        u5_mult_79_CARRYB_6__6_), .ZN(u5_mult_79_n920) );
  NAND2_X1 u5_mult_79_U2016 ( .A1(u5_mult_79_CARRYB_6__6_), .A2(
        u5_mult_79_SUMB_6__7_), .ZN(u5_mult_79_n918) );
  NAND3_X2 u5_mult_79_U2015 ( .A1(u5_mult_79_n915), .A2(u5_mult_79_n916), .A3(
        u5_mult_79_n917), .ZN(u5_mult_79_CARRYB_11__4_) );
  NAND2_X1 u5_mult_79_U2014 ( .A1(u5_mult_79_ab_11__4_), .A2(
        u5_mult_79_CARRYB_10__4_), .ZN(u5_mult_79_n917) );
  NAND2_X2 u5_mult_79_U2013 ( .A1(u5_mult_79_ab_11__4_), .A2(
        u5_mult_79_SUMB_10__5_), .ZN(u5_mult_79_n916) );
  NAND2_X1 u5_mult_79_U2012 ( .A1(u5_mult_79_SUMB_10__5_), .A2(
        u5_mult_79_CARRYB_10__4_), .ZN(u5_mult_79_n915) );
  NAND2_X1 u5_mult_79_U2011 ( .A1(u5_mult_79_ab_10__5_), .A2(
        u5_mult_79_CARRYB_9__5_), .ZN(u5_mult_79_n914) );
  NAND2_X2 u5_mult_79_U2010 ( .A1(u5_mult_79_SUMB_9__6_), .A2(
        u5_mult_79_ab_10__5_), .ZN(u5_mult_79_n913) );
  NAND2_X2 u5_mult_79_U2009 ( .A1(u5_mult_79_CARRYB_9__5_), .A2(
        u5_mult_79_SUMB_9__6_), .ZN(u5_mult_79_n912) );
  NAND2_X2 u5_mult_79_U2008 ( .A1(u5_mult_79_CARRYB_11__5_), .A2(
        u5_mult_79_n385), .ZN(u5_mult_79_n1115) );
  NAND2_X2 u5_mult_79_U2007 ( .A1(u5_mult_79_n783), .A2(u5_mult_79_SUMB_17__7_), .ZN(u5_mult_79_n1596) );
  XNOR2_X2 u5_mult_79_U2006 ( .A(u5_mult_79_n911), .B(u5_mult_79_CARRYB_2__14_), .ZN(u5_mult_79_SUMB_3__14_) );
  NAND2_X2 u5_mult_79_U2005 ( .A1(u5_mult_79_n376), .A2(u5_mult_79_n267), .ZN(
        u5_mult_79_n1243) );
  NAND3_X2 u5_mult_79_U2004 ( .A1(u5_mult_79_n1622), .A2(u5_mult_79_n1623), 
        .A3(u5_mult_79_n1624), .ZN(u5_mult_79_CARRYB_2__21_) );
  NAND2_X2 u5_mult_79_U2003 ( .A1(u5_mult_79_SUMB_15__9_), .A2(
        u5_mult_79_ab_16__8_), .ZN(u5_mult_79_n1322) );
  NAND3_X2 u5_mult_79_U2002 ( .A1(u5_mult_79_n1415), .A2(u5_mult_79_n1417), 
        .A3(u5_mult_79_n1416), .ZN(u5_mult_79_CARRYB_7__13_) );
  NAND2_X2 u5_mult_79_U2001 ( .A1(u5_mult_79_ab_15__8_), .A2(
        u5_mult_79_CARRYB_14__8_), .ZN(u5_mult_79_n1477) );
  XNOR2_X2 u5_mult_79_U2000 ( .A(u5_mult_79_SUMB_10__22_), .B(
        u5_mult_79_ab_11__21_), .ZN(u5_mult_79_n910) );
  XNOR2_X2 u5_mult_79_U1999 ( .A(u5_mult_79_SUMB_18__5_), .B(u5_mult_79_n909), 
        .ZN(u5_mult_79_SUMB_19__4_) );
  XNOR2_X2 u5_mult_79_U1998 ( .A(u5_mult_79_SUMB_10__3_), .B(u5_mult_79_n908), 
        .ZN(u5_mult_79_SUMB_11__2_) );
  XNOR2_X2 u5_mult_79_U1997 ( .A(u5_mult_79_ab_8__16_), .B(
        u5_mult_79_CARRYB_7__16_), .ZN(u5_mult_79_n906) );
  XNOR2_X2 u5_mult_79_U1996 ( .A(u5_mult_79_n906), .B(u5_mult_79_SUMB_7__17_), 
        .ZN(u5_mult_79_SUMB_8__16_) );
  NAND2_X2 u5_mult_79_U1995 ( .A1(u5_mult_79_ab_10__15_), .A2(
        u5_mult_79_SUMB_9__16_), .ZN(u5_mult_79_n1273) );
  XNOR2_X2 u5_mult_79_U1994 ( .A(u5_mult_79_ab_10__4_), .B(
        u5_mult_79_CARRYB_9__4_), .ZN(u5_mult_79_n905) );
  XNOR2_X2 u5_mult_79_U1993 ( .A(u5_mult_79_n905), .B(u5_mult_79_SUMB_9__5_), 
        .ZN(u5_mult_79_SUMB_10__4_) );
  XNOR2_X2 u5_mult_79_U1992 ( .A(u5_mult_79_n904), .B(u5_mult_79_n389), .ZN(
        u5_mult_79_SUMB_17__9_) );
  XNOR2_X2 u5_mult_79_U1991 ( .A(u5_mult_79_ab_7__16_), .B(
        u5_mult_79_CARRYB_6__16_), .ZN(u5_mult_79_n903) );
  XNOR2_X2 u5_mult_79_U1990 ( .A(u5_mult_79_SUMB_6__17_), .B(u5_mult_79_n903), 
        .ZN(u5_mult_79_SUMB_7__16_) );
  NAND2_X2 u5_mult_79_U1989 ( .A1(u5_mult_79_ab_9__13_), .A2(
        u5_mult_79_CARRYB_8__13_), .ZN(u5_mult_79_n1293) );
  NAND2_X2 u5_mult_79_U1988 ( .A1(u5_mult_79_CARRYB_18__7_), .A2(
        u5_mult_79_SUMB_18__8_), .ZN(u5_mult_79_n1644) );
  NAND3_X4 u5_mult_79_U1987 ( .A1(u5_mult_79_n1150), .A2(u5_mult_79_n1151), 
        .A3(u5_mult_79_n1152), .ZN(u5_mult_79_CARRYB_5__20_) );
  NAND3_X4 u5_mult_79_U1986 ( .A1(u5_mult_79_n897), .A2(u5_mult_79_n898), .A3(
        u5_mult_79_n899), .ZN(u5_mult_79_CARRYB_13__14_) );
  NAND2_X1 u5_mult_79_U1985 ( .A1(u5_mult_79_ab_13__14_), .A2(
        u5_mult_79_CARRYB_12__14_), .ZN(u5_mult_79_n899) );
  NAND2_X2 u5_mult_79_U1984 ( .A1(u5_mult_79_CARRYB_12__14_), .A2(
        u5_mult_79_SUMB_12__15_), .ZN(u5_mult_79_n897) );
  XNOR2_X2 u5_mult_79_U1983 ( .A(u5_mult_79_ab_10__15_), .B(
        u5_mult_79_CARRYB_9__15_), .ZN(u5_mult_79_n892) );
  XNOR2_X2 u5_mult_79_U1982 ( .A(u5_mult_79_n891), .B(u5_mult_79_SUMB_19__5_), 
        .ZN(u5_mult_79_SUMB_20__4_) );
  XNOR2_X2 u5_mult_79_U1981 ( .A(u5_mult_79_ab_6__16_), .B(
        u5_mult_79_CARRYB_5__16_), .ZN(u5_mult_79_n890) );
  XNOR2_X2 u5_mult_79_U1980 ( .A(u5_mult_79_n890), .B(u5_mult_79_n34), .ZN(
        u5_mult_79_SUMB_6__16_) );
  NAND3_X2 u5_mult_79_U1979 ( .A1(u5_mult_79_n1454), .A2(u5_mult_79_n1453), 
        .A3(u5_mult_79_n1452), .ZN(u5_mult_79_CARRYB_22__10_) );
  XNOR2_X2 u5_mult_79_U1978 ( .A(u5_mult_79_CARRYB_7__13_), .B(
        u5_mult_79_ab_8__13_), .ZN(u5_mult_79_n889) );
  XNOR2_X2 u5_mult_79_U1977 ( .A(u5_mult_79_SUMB_7__14_), .B(u5_mult_79_n889), 
        .ZN(u5_mult_79_SUMB_8__13_) );
  NOR2_X1 u5_mult_79_U1976 ( .A1(u5_mult_79_n1823), .A2(u5_mult_79_n1749), 
        .ZN(u5_mult_79_ab_11__3_) );
  NAND3_X2 u5_mult_79_U1975 ( .A1(u5_mult_79_n886), .A2(u5_mult_79_n887), .A3(
        u5_mult_79_n888), .ZN(u5_mult_79_CARRYB_11__3_) );
  NAND2_X1 u5_mult_79_U1974 ( .A1(u5_mult_79_ab_11__3_), .A2(
        u5_mult_79_SUMB_10__4_), .ZN(u5_mult_79_n888) );
  NAND3_X2 u5_mult_79_U1973 ( .A1(u5_mult_79_n883), .A2(u5_mult_79_n884), .A3(
        u5_mult_79_n885), .ZN(u5_mult_79_CARRYB_6__6_) );
  NAND2_X1 u5_mult_79_U1972 ( .A1(u5_mult_79_ab_6__6_), .A2(
        u5_mult_79_SUMB_5__7_), .ZN(u5_mult_79_n884) );
  NAND2_X1 u5_mult_79_U1971 ( .A1(u5_mult_79_CARRYB_4__7_), .A2(
        u5_mult_79_SUMB_4__8_), .ZN(u5_mult_79_n882) );
  NAND2_X1 u5_mult_79_U1970 ( .A1(u5_mult_79_ab_5__7_), .A2(
        u5_mult_79_SUMB_4__8_), .ZN(u5_mult_79_n881) );
  NAND2_X1 u5_mult_79_U1969 ( .A1(u5_mult_79_ab_5__7_), .A2(
        u5_mult_79_CARRYB_4__7_), .ZN(u5_mult_79_n880) );
  XOR2_X2 u5_mult_79_U1968 ( .A(u5_mult_79_n879), .B(u5_mult_79_SUMB_4__8_), 
        .Z(u5_mult_79_SUMB_5__7_) );
  XOR2_X2 u5_mult_79_U1967 ( .A(u5_mult_79_ab_5__7_), .B(
        u5_mult_79_CARRYB_4__7_), .Z(u5_mult_79_n879) );
  NAND2_X2 u5_mult_79_U1966 ( .A1(u5_mult_79_CARRYB_2__22_), .A2(
        u5_mult_79_ab_3__22_), .ZN(u5_mult_79_n1616) );
  NAND2_X2 u5_mult_79_U1965 ( .A1(u5_mult_79_CARRYB_2__22_), .A2(
        u5_mult_79_ab_2__23_), .ZN(u5_mult_79_n1617) );
  INV_X8 u5_mult_79_U1964 ( .A(u6_N23), .ZN(u5_mult_79_n1880) );
  XNOR2_X2 u5_mult_79_U1963 ( .A(u5_mult_79_ab_9__16_), .B(
        u5_mult_79_CARRYB_8__16_), .ZN(u5_mult_79_n878) );
  XNOR2_X2 u5_mult_79_U1962 ( .A(u5_mult_79_ab_20__1_), .B(
        u5_mult_79_CARRYB_19__1_), .ZN(u5_mult_79_n877) );
  XNOR2_X2 u5_mult_79_U1961 ( .A(u5_mult_79_ab_6__15_), .B(
        u5_mult_79_CARRYB_5__15_), .ZN(u5_mult_79_n1031) );
  XNOR2_X2 u5_mult_79_U1960 ( .A(u5_mult_79_ab_3__16_), .B(
        u5_mult_79_CARRYB_2__16_), .ZN(u5_mult_79_n876) );
  XNOR2_X2 u5_mult_79_U1959 ( .A(u5_mult_79_n876), .B(u5_mult_79_n488), .ZN(
        u5_mult_79_SUMB_3__16_) );
  NAND2_X4 u5_mult_79_U1958 ( .A1(u5_mult_79_n1202), .A2(u5_mult_79_n1203), 
        .ZN(u5_mult_79_n1205) );
  NAND2_X4 u5_mult_79_U1957 ( .A1(u5_mult_79_n1204), .A2(u5_mult_79_n1205), 
        .ZN(u5_mult_79_n1525) );
  NAND2_X2 u5_mult_79_U1956 ( .A1(u5_mult_79_ab_21__1_), .A2(
        u5_mult_79_SUMB_20__2_), .ZN(u5_mult_79_n1386) );
  NAND3_X4 u5_mult_79_U1955 ( .A1(u5_mult_79_n1402), .A2(u5_mult_79_n1403), 
        .A3(u5_mult_79_n1404), .ZN(u5_mult_79_CARRYB_11__12_) );
  NOR2_X1 u5_mult_79_U1954 ( .A1(u5_mult_79_n1821), .A2(u5_mult_79_n1755), 
        .ZN(u5_mult_79_ab_13__4_) );
  NAND3_X2 u5_mult_79_U1953 ( .A1(u5_mult_79_n873), .A2(u5_mult_79_n874), .A3(
        u5_mult_79_n875), .ZN(u5_mult_79_CARRYB_13__4_) );
  NAND2_X2 u5_mult_79_U1952 ( .A1(u5_mult_79_ab_13__4_), .A2(
        u5_mult_79_SUMB_12__5_), .ZN(u5_mult_79_n874) );
  NAND2_X1 u5_mult_79_U1951 ( .A1(u5_mult_79_n372), .A2(u5_mult_79_SUMB_12__5_), .ZN(u5_mult_79_n873) );
  CLKBUF_X2 u5_mult_79_U1950 ( .A(u5_mult_79_CARRYB_4__10_), .Z(
        u5_mult_79_n872) );
  NAND3_X2 u5_mult_79_U1949 ( .A1(u5_mult_79_n869), .A2(u5_mult_79_n870), .A3(
        u5_mult_79_n871), .ZN(u5_mult_79_CARRYB_6__9_) );
  NAND2_X2 u5_mult_79_U1948 ( .A1(u5_mult_79_ab_6__9_), .A2(
        u5_mult_79_SUMB_5__10_), .ZN(u5_mult_79_n870) );
  NAND2_X1 u5_mult_79_U1947 ( .A1(u5_mult_79_ab_6__9_), .A2(
        u5_mult_79_CARRYB_5__9_), .ZN(u5_mult_79_n869) );
  NAND3_X2 u5_mult_79_U1946 ( .A1(u5_mult_79_n866), .A2(u5_mult_79_n867), .A3(
        u5_mult_79_n868), .ZN(u5_mult_79_CARRYB_5__10_) );
  NAND2_X1 u5_mult_79_U1945 ( .A1(u5_mult_79_ab_5__10_), .A2(
        u5_mult_79_SUMB_4__11_), .ZN(u5_mult_79_n867) );
  XOR2_X2 u5_mult_79_U1944 ( .A(u5_mult_79_n865), .B(u5_mult_79_SUMB_4__11_), 
        .Z(u5_mult_79_SUMB_5__10_) );
  XOR2_X2 u5_mult_79_U1943 ( .A(u5_mult_79_ab_5__10_), .B(
        u5_mult_79_CARRYB_4__10_), .Z(u5_mult_79_n865) );
  NAND3_X2 u5_mult_79_U1942 ( .A1(u5_mult_79_n862), .A2(u5_mult_79_n863), .A3(
        u5_mult_79_n864), .ZN(u5_mult_79_CARRYB_17__2_) );
  NAND2_X1 u5_mult_79_U1941 ( .A1(u5_mult_79_ab_17__2_), .A2(
        u5_mult_79_SUMB_16__3_), .ZN(u5_mult_79_n863) );
  NAND2_X2 u5_mult_79_U1940 ( .A1(u5_mult_79_CARRYB_15__3_), .A2(
        u5_mult_79_SUMB_15__4_), .ZN(u5_mult_79_n861) );
  NAND2_X2 u5_mult_79_U1939 ( .A1(u5_mult_79_ab_16__3_), .A2(u5_mult_79_n312), 
        .ZN(u5_mult_79_n860) );
  NAND2_X2 u5_mult_79_U1938 ( .A1(u5_mult_79_CARRYB_15__3_), .A2(
        u5_mult_79_ab_16__3_), .ZN(u5_mult_79_n859) );
  XNOR2_X2 u5_mult_79_U1937 ( .A(u5_mult_79_SUMB_2__15_), .B(
        u5_mult_79_ab_3__14_), .ZN(u5_mult_79_n911) );
  NAND2_X2 u5_mult_79_U1936 ( .A1(u5_mult_79_n492), .A2(u5_mult_79_SUMB_19__2_), .ZN(u5_mult_79_n1385) );
  XNOR2_X2 u5_mult_79_U1935 ( .A(u5_mult_79_CARRYB_12__10_), .B(
        u5_mult_79_n858), .ZN(u5_mult_79_SUMB_13__10_) );
  NAND2_X2 u5_mult_79_U1934 ( .A1(u5_mult_79_ab_13__8_), .A2(
        u5_mult_79_SUMB_12__9_), .ZN(u5_mult_79_n1469) );
  NAND2_X2 u5_mult_79_U1933 ( .A1(u5_mult_79_ab_8__15_), .A2(
        u5_mult_79_CARRYB_7__15_), .ZN(u5_mult_79_n1398) );
  NOR2_X1 u5_mult_79_U1932 ( .A1(u5_mult_79_n1796), .A2(u5_mult_79_n1738), 
        .ZN(u5_mult_79_ab_7__15_) );
  NOR2_X1 u5_mult_79_U1931 ( .A1(u5_mult_79_n1867), .A2(u5_mult_79_n1744), 
        .ZN(u5_mult_79_ab_9__14_) );
  NAND2_X2 u5_mult_79_U1930 ( .A1(u5_mult_79_ab_7__15_), .A2(
        u5_mult_79_CARRYB_6__15_), .ZN(u5_mult_79_n856) );
  NAND3_X2 u5_mult_79_U1929 ( .A1(u5_mult_79_n852), .A2(u5_mult_79_n853), .A3(
        u5_mult_79_n854), .ZN(u5_mult_79_CARRYB_9__14_) );
  NAND2_X1 u5_mult_79_U1928 ( .A1(u5_mult_79_ab_9__14_), .A2(
        u5_mult_79_CARRYB_8__14_), .ZN(u5_mult_79_n854) );
  INV_X8 u5_mult_79_U1927 ( .A(u5_mult_79_CARRYB_16__11_), .ZN(
        u5_mult_79_n1203) );
  XNOR2_X2 u5_mult_79_U1926 ( .A(u5_mult_79_n848), .B(u5_mult_79_CARRYB_5__11_), .ZN(u5_mult_79_n1250) );
  XNOR2_X2 u5_mult_79_U1925 ( .A(u5_mult_79_CARRYB_3__16_), .B(
        u5_mult_79_ab_4__16_), .ZN(u5_mult_79_n847) );
  XNOR2_X2 u5_mult_79_U1924 ( .A(u5_mult_79_SUMB_3__17_), .B(u5_mult_79_n847), 
        .ZN(u5_mult_79_SUMB_4__16_) );
  XOR2_X2 u5_mult_79_U1923 ( .A(u5_mult_79_n105), .B(u5_mult_79_n1015), .Z(
        u5_mult_79_SUMB_7__7_) );
  NAND2_X2 u5_mult_79_U1922 ( .A1(u5_mult_79_ab_8__6_), .A2(
        u5_mult_79_SUMB_7__7_), .ZN(u5_mult_79_n922) );
  NAND2_X2 u5_mult_79_U1921 ( .A1(u5_mult_79_n282), .A2(
        u5_mult_79_CARRYB_4__21_), .ZN(u5_mult_79_n1551) );
  INV_X4 u5_mult_79_U1920 ( .A(u5_mult_79_CARRYB_14__12_), .ZN(
        u5_mult_79_n1240) );
  XNOR2_X2 u5_mult_79_U1919 ( .A(u5_mult_79_n846), .B(u5_mult_79_SUMB_16__3_), 
        .ZN(u5_mult_79_SUMB_17__2_) );
  NOR2_X1 u5_mult_79_U1918 ( .A1(u5_mult_79_n1808), .A2(u5_mult_79_n1743), 
        .ZN(u5_mult_79_ab_9__8_) );
  NAND2_X1 u5_mult_79_U1917 ( .A1(u5_mult_79_ab_9__8_), .A2(
        u5_mult_79_CARRYB_8__8_), .ZN(u5_mult_79_n845) );
  NAND2_X1 u5_mult_79_U1916 ( .A1(u5_mult_79_CARRYB_8__8_), .A2(
        u5_mult_79_SUMB_8__9_), .ZN(u5_mult_79_n843) );
  XOR2_X2 u5_mult_79_U1915 ( .A(u5_mult_79_SUMB_8__9_), .B(u5_mult_79_n842), 
        .Z(u5_mult_79_SUMB_9__8_) );
  XOR2_X2 u5_mult_79_U1914 ( .A(u5_mult_79_CARRYB_8__8_), .B(
        u5_mult_79_ab_9__8_), .Z(u5_mult_79_n842) );
  NAND3_X4 u5_mult_79_U1913 ( .A1(u5_mult_79_n839), .A2(u5_mult_79_n840), .A3(
        u5_mult_79_n841), .ZN(u5_mult_79_CARRYB_6__10_) );
  NAND2_X2 u5_mult_79_U1912 ( .A1(u5_mult_79_CARRYB_5__10_), .A2(
        u5_mult_79_SUMB_5__11_), .ZN(u5_mult_79_n841) );
  NAND2_X2 u5_mult_79_U1911 ( .A1(u5_mult_79_ab_6__10_), .A2(
        u5_mult_79_SUMB_5__11_), .ZN(u5_mult_79_n840) );
  NAND2_X1 u5_mult_79_U1910 ( .A1(u5_mult_79_ab_6__10_), .A2(
        u5_mult_79_CARRYB_5__10_), .ZN(u5_mult_79_n839) );
  NAND3_X4 u5_mult_79_U1909 ( .A1(u5_mult_79_n836), .A2(u5_mult_79_n837), .A3(
        u5_mult_79_n838), .ZN(u5_mult_79_CARRYB_5__11_) );
  NAND2_X2 u5_mult_79_U1908 ( .A1(u5_mult_79_CARRYB_4__11_), .A2(
        u5_mult_79_SUMB_4__12_), .ZN(u5_mult_79_n838) );
  NAND2_X2 u5_mult_79_U1907 ( .A1(u5_mult_79_ab_5__11_), .A2(
        u5_mult_79_SUMB_4__12_), .ZN(u5_mult_79_n837) );
  NAND2_X1 u5_mult_79_U1906 ( .A1(u5_mult_79_ab_5__11_), .A2(
        u5_mult_79_CARRYB_4__11_), .ZN(u5_mult_79_n836) );
  XOR2_X2 u5_mult_79_U1905 ( .A(u5_mult_79_n835), .B(u5_mult_79_SUMB_5__11_), 
        .Z(u5_mult_79_SUMB_6__10_) );
  XNOR2_X2 u5_mult_79_U1904 ( .A(u5_mult_79_n1181), .B(u5_mult_79_n1705), .ZN(
        u5_mult_79_SUMB_2__16_) );
  XNOR2_X2 u5_mult_79_U1903 ( .A(u5_mult_79_SUMB_16__19_), .B(
        u5_mult_79_ab_17__18_), .ZN(u5_mult_79_n834) );
  XNOR2_X2 u5_mult_79_U1902 ( .A(u5_mult_79_n126), .B(u5_mult_79_n834), .ZN(
        u5_mult_79_SUMB_17__18_) );
  NAND3_X2 u5_mult_79_U1901 ( .A1(u5_mult_79_n1017), .A2(u5_mult_79_n1016), 
        .A3(u5_mult_79_n1018), .ZN(u5_mult_79_CARRYB_7__7_) );
  NAND3_X4 u5_mult_79_U1900 ( .A1(u5_mult_79_n1486), .A2(u5_mult_79_n1487), 
        .A3(u5_mult_79_n1488), .ZN(u5_mult_79_CARRYB_14__12_) );
  INV_X1 u5_mult_79_U1899 ( .A(u5_mult_79_SUMB_13__18_), .ZN(u5_mult_79_n831)
         );
  INV_X2 u5_mult_79_U1898 ( .A(u5_mult_79_n1148), .ZN(u5_mult_79_n830) );
  NAND2_X1 u5_mult_79_U1897 ( .A1(u5_mult_79_n1148), .A2(
        u5_mult_79_SUMB_13__18_), .ZN(u5_mult_79_n832) );
  NAND2_X4 u5_mult_79_U1896 ( .A1(u5_mult_79_ab_14__12_), .A2(u5_mult_79_n1426), .ZN(u5_mult_79_n1487) );
  XNOR2_X2 u5_mult_79_U1895 ( .A(u5_mult_79_CARRYB_3__21_), .B(
        u5_mult_79_n1543), .ZN(u5_mult_79_SUMB_4__21_) );
  NAND2_X2 u5_mult_79_U1894 ( .A1(u5_mult_79_n969), .A2(u5_mult_79_SUMB_4__21_), .ZN(u5_mult_79_n1150) );
  XNOR2_X2 u5_mult_79_U1893 ( .A(u5_mult_79_n829), .B(u5_mult_79_n433), .ZN(
        u5_mult_79_SUMB_11__9_) );
  XNOR2_X2 u5_mult_79_U1892 ( .A(u5_mult_79_n828), .B(u5_mult_79_n476), .ZN(
        u5_mult_79_SUMB_14__15_) );
  XNOR2_X2 u5_mult_79_U1891 ( .A(u5_mult_79_SUMB_3__21_), .B(u5_mult_79_n1264), 
        .ZN(u5_mult_79_SUMB_4__20_) );
  NAND2_X2 u5_mult_79_U1890 ( .A1(u5_mult_79_ab_19__10_), .A2(
        u5_mult_79_CARRYB_18__10_), .ZN(u5_mult_79_n1518) );
  NAND2_X4 u5_mult_79_U1889 ( .A1(u5_mult_79_n1214), .A2(u5_mult_79_n1215), 
        .ZN(u5_mult_79_SUMB_17__11_) );
  NOR2_X2 u5_mult_79_U1888 ( .A1(u5_mult_79_n1803), .A2(u5_mult_79_n1770), 
        .ZN(u5_mult_79_ab_18__10_) );
  NAND3_X4 u5_mult_79_U1887 ( .A1(u5_mult_79_n825), .A2(u5_mult_79_n826), .A3(
        u5_mult_79_n827), .ZN(u5_mult_79_CARRYB_18__10_) );
  NAND2_X2 u5_mult_79_U1886 ( .A1(u5_mult_79_ab_18__10_), .A2(
        u5_mult_79_CARRYB_17__10_), .ZN(u5_mult_79_n827) );
  NAND2_X4 u5_mult_79_U1885 ( .A1(u5_mult_79_ab_18__10_), .A2(
        u5_mult_79_SUMB_17__11_), .ZN(u5_mult_79_n826) );
  NAND2_X1 u5_mult_79_U1884 ( .A1(u5_mult_79_ab_12__15_), .A2(
        u5_mult_79_CARRYB_11__15_), .ZN(u5_mult_79_n822) );
  NAND2_X1 u5_mult_79_U1883 ( .A1(u5_mult_79_ab_11__16_), .A2(
        u5_mult_79_CARRYB_10__16_), .ZN(u5_mult_79_n819) );
  NAND3_X4 u5_mult_79_U1882 ( .A1(u5_mult_79_n816), .A2(u5_mult_79_n817), .A3(
        u5_mult_79_n818), .ZN(u5_mult_79_CARRYB_21__7_) );
  NAND2_X2 u5_mult_79_U1881 ( .A1(u5_mult_79_CARRYB_20__7_), .A2(
        u5_mult_79_SUMB_20__8_), .ZN(u5_mult_79_n818) );
  NAND2_X2 u5_mult_79_U1880 ( .A1(u5_mult_79_ab_21__7_), .A2(
        u5_mult_79_SUMB_20__8_), .ZN(u5_mult_79_n817) );
  NAND3_X4 u5_mult_79_U1879 ( .A1(u5_mult_79_n813), .A2(u5_mult_79_n814), .A3(
        u5_mult_79_n815), .ZN(u5_mult_79_CARRYB_20__8_) );
  NAND2_X2 u5_mult_79_U1878 ( .A1(u5_mult_79_SUMB_19__9_), .A2(
        u5_mult_79_CARRYB_19__8_), .ZN(u5_mult_79_n815) );
  NAND2_X2 u5_mult_79_U1877 ( .A1(u5_mult_79_ab_20__8_), .A2(
        u5_mult_79_SUMB_19__9_), .ZN(u5_mult_79_n814) );
  NAND2_X1 u5_mult_79_U1876 ( .A1(u5_mult_79_ab_20__8_), .A2(
        u5_mult_79_CARRYB_19__8_), .ZN(u5_mult_79_n813) );
  XOR2_X2 u5_mult_79_U1875 ( .A(u5_mult_79_n812), .B(u5_mult_79_n374), .Z(
        u5_mult_79_SUMB_21__7_) );
  XNOR2_X2 u5_mult_79_U1874 ( .A(u5_mult_79_CARRYB_6__7_), .B(u5_mult_79_n811), 
        .ZN(u5_mult_79_n1015) );
  NAND2_X2 u5_mult_79_U1873 ( .A1(u5_mult_79_ab_20__1_), .A2(
        u5_mult_79_SUMB_19__2_), .ZN(u5_mult_79_n1384) );
  NOR2_X2 u5_mult_79_U1872 ( .A1(u5_mult_79_n1867), .A2(u5_mult_79_n1723), 
        .ZN(u5_mult_79_ab_2__14_) );
  XNOR2_X2 u5_mult_79_U1871 ( .A(u5_mult_79_ab_4__14_), .B(
        u5_mult_79_CARRYB_3__14_), .ZN(u5_mult_79_n809) );
  XNOR2_X2 u5_mult_79_U1870 ( .A(u5_mult_79_ab_11__9_), .B(
        u5_mult_79_CARRYB_10__9_), .ZN(u5_mult_79_n829) );
  XNOR2_X2 u5_mult_79_U1869 ( .A(u5_mult_79_SUMB_11__22_), .B(
        u5_mult_79_ab_12__21_), .ZN(u5_mult_79_n808) );
  XNOR2_X2 u5_mult_79_U1868 ( .A(u5_mult_79_n877), .B(u5_mult_79_SUMB_19__2_), 
        .ZN(u5_mult_79_SUMB_20__1_) );
  XNOR2_X2 u5_mult_79_U1867 ( .A(u5_mult_79_CARRYB_11__9_), .B(
        u5_mult_79_ab_12__9_), .ZN(u5_mult_79_n807) );
  XNOR2_X2 u5_mult_79_U1866 ( .A(u5_mult_79_n807), .B(u5_mult_79_n364), .ZN(
        u5_mult_79_SUMB_12__9_) );
  NAND3_X2 u5_mult_79_U1865 ( .A1(u5_mult_79_n1373), .A2(u5_mult_79_n1374), 
        .A3(u5_mult_79_n1375), .ZN(u5_mult_79_CARRYB_9__17_) );
  XNOR2_X2 u5_mult_79_U1864 ( .A(u5_mult_79_n806), .B(u5_mult_79_CARRYB_4__13_), .ZN(u5_mult_79_n1339) );
  NAND2_X2 u5_mult_79_U1863 ( .A1(u5_mult_79_CARRYB_13__16_), .A2(
        u5_mult_79_n484), .ZN(u5_mult_79_n1438) );
  NAND2_X2 u5_mult_79_U1862 ( .A1(u5_mult_79_n1544), .A2(
        u5_mult_79_SUMB_3__20_), .ZN(u5_mult_79_n1218) );
  NAND2_X2 u5_mult_79_U1861 ( .A1(u5_mult_79_SUMB_13__3_), .A2(
        u5_mult_79_CARRYB_13__2_), .ZN(u5_mult_79_n924) );
  XNOR2_X2 u5_mult_79_U1860 ( .A(u5_mult_79_n805), .B(u5_mult_79_SUMB_13__8_), 
        .ZN(u5_mult_79_SUMB_14__7_) );
  NOR2_X1 u5_mult_79_U1859 ( .A1(u5_mult_79_n1791), .A2(u5_mult_79_n1771), 
        .ZN(u5_mult_79_ab_18__17_) );
  NAND3_X2 u5_mult_79_U1858 ( .A1(u5_mult_79_n804), .A2(u5_mult_79_n803), .A3(
        u5_mult_79_n802), .ZN(u5_mult_79_CARRYB_18__17_) );
  NAND2_X1 u5_mult_79_U1857 ( .A1(u5_mult_79_ab_18__17_), .A2(
        u5_mult_79_CARRYB_17__17_), .ZN(u5_mult_79_n803) );
  NAND2_X1 u5_mult_79_U1856 ( .A1(u5_mult_79_n334), .A2(
        u5_mult_79_CARRYB_17__17_), .ZN(u5_mult_79_n802) );
  XOR2_X2 u5_mult_79_U1855 ( .A(u5_mult_79_CARRYB_17__17_), .B(u5_mult_79_n801), .Z(u5_mult_79_SUMB_18__17_) );
  NAND3_X4 u5_mult_79_U1854 ( .A1(u5_mult_79_n1610), .A2(u5_mult_79_n1611), 
        .A3(u5_mult_79_n1612), .ZN(u5_mult_79_CARRYB_17__8_) );
  NAND2_X2 u5_mult_79_U1853 ( .A1(u5_mult_79_CARRYB_7__6_), .A2(
        u5_mult_79_SUMB_7__7_), .ZN(u5_mult_79_n921) );
  NAND2_X1 u5_mult_79_U1852 ( .A1(u5_mult_79_CARRYB_7__7_), .A2(
        u5_mult_79_SUMB_7__8_), .ZN(u5_mult_79_n1170) );
  NAND2_X2 u5_mult_79_U1851 ( .A1(u5_mult_79_ab_7__18_), .A2(
        u5_mult_79_SUMB_6__19_), .ZN(u5_mult_79_n1276) );
  XNOR2_X2 u5_mult_79_U1850 ( .A(u5_mult_79_SUMB_6__22_), .B(u5_mult_79_n800), 
        .ZN(u5_mult_79_n1064) );
  NAND2_X1 u5_mult_79_U1849 ( .A1(u5_mult_79_SUMB_18__5_), .A2(
        u5_mult_79_CARRYB_18__4_), .ZN(u5_mult_79_n1588) );
  NAND3_X2 u5_mult_79_U1848 ( .A1(u5_mult_79_n1500), .A2(u5_mult_79_n1499), 
        .A3(u5_mult_79_n1498), .ZN(u5_mult_79_CARRYB_15__5_) );
  NAND3_X4 u5_mult_79_U1847 ( .A1(u5_mult_79_n973), .A2(u5_mult_79_n974), .A3(
        u5_mult_79_n975), .ZN(u5_mult_79_CARRYB_8__14_) );
  NAND3_X2 u5_mult_79_U1846 ( .A1(u5_mult_79_n1233), .A2(u5_mult_79_n1234), 
        .A3(u5_mult_79_n1235), .ZN(u5_mult_79_CARRYB_13__18_) );
  XNOR2_X2 u5_mult_79_U1845 ( .A(u5_mult_79_CARRYB_19__4_), .B(
        u5_mult_79_ab_20__4_), .ZN(u5_mult_79_n891) );
  NAND2_X2 u5_mult_79_U1844 ( .A1(u5_mult_79_ab_20__4_), .A2(
        u5_mult_79_CARRYB_19__4_), .ZN(u5_mult_79_n1542) );
  NAND2_X2 u5_mult_79_U1843 ( .A1(u5_mult_79_n268), .A2(u5_mult_79_n32), .ZN(
        u5_mult_79_n1324) );
  NAND2_X2 u5_mult_79_U1842 ( .A1(u5_mult_79_CARRYB_5__20_), .A2(
        u5_mult_79_SUMB_5__21_), .ZN(u5_mult_79_n900) );
  XNOR2_X2 u5_mult_79_U1841 ( .A(u5_mult_79_SUMB_17__18_), .B(u5_mult_79_n799), 
        .ZN(u5_mult_79_n801) );
  INV_X8 u5_mult_79_U1840 ( .A(fracta_mul[3]), .ZN(u5_mult_79_n1839) );
  NAND3_X4 u5_mult_79_U1839 ( .A1(u5_mult_79_n1474), .A2(u5_mult_79_n1475), 
        .A3(u5_mult_79_n1476), .ZN(u5_mult_79_CARRYB_17__5_) );
  XNOR2_X2 u5_mult_79_U1838 ( .A(u5_mult_79_CARRYB_15__5_), .B(
        u5_mult_79_ab_16__5_), .ZN(u5_mult_79_n1132) );
  INV_X8 u5_mult_79_U1837 ( .A(n2923), .ZN(u5_mult_79_n1870) );
  XNOR2_X2 u5_mult_79_U1836 ( .A(u5_mult_79_ab_3__22_), .B(
        u5_mult_79_ab_2__23_), .ZN(u5_mult_79_n797) );
  XNOR2_X1 u5_mult_79_U1835 ( .A(u5_mult_79_CARRYB_2__22_), .B(u5_mult_79_n797), .ZN(u5_mult_79_SUMB_3__22_) );
  NAND2_X2 u5_mult_79_U1834 ( .A1(u5_mult_79_CARRYB_5__14_), .A2(
        u5_mult_79_n496), .ZN(u5_mult_79_n1414) );
  NAND3_X2 u5_mult_79_U1833 ( .A1(u5_mult_79_n1559), .A2(u5_mult_79_n1560), 
        .A3(u5_mult_79_n1561), .ZN(u5_mult_79_CARRYB_21__6_) );
  XNOR2_X2 u5_mult_79_U1832 ( .A(u5_mult_79_ab_23__11_), .B(
        u5_mult_79_CARRYB_22__11_), .ZN(u5_mult_79_n796) );
  NAND3_X2 u5_mult_79_U1831 ( .A1(u5_mult_79_n912), .A2(u5_mult_79_n913), .A3(
        u5_mult_79_n914), .ZN(u5_mult_79_CARRYB_10__5_) );
  XNOR2_X2 u5_mult_79_U1830 ( .A(u5_mult_79_CARRYB_15__16_), .B(
        u5_mult_79_ab_16__16_), .ZN(u5_mult_79_n795) );
  XNOR2_X2 u5_mult_79_U1829 ( .A(u5_mult_79_n23), .B(u5_mult_79_n795), .ZN(
        u5_mult_79_SUMB_16__16_) );
  NAND3_X4 u5_mult_79_U1828 ( .A1(u5_mult_79_n1115), .A2(u5_mult_79_n1116), 
        .A3(u5_mult_79_n1117), .ZN(u5_mult_79_CARRYB_12__5_) );
  XNOR2_X2 u5_mult_79_U1827 ( .A(u5_mult_79_CARRYB_10__5_), .B(
        u5_mult_79_ab_11__5_), .ZN(u5_mult_79_n794) );
  XNOR2_X2 u5_mult_79_U1826 ( .A(u5_mult_79_n404), .B(u5_mult_79_n794), .ZN(
        u5_mult_79_SUMB_11__5_) );
  XNOR2_X2 u5_mult_79_U1825 ( .A(u5_mult_79_CARRYB_12__9_), .B(
        u5_mult_79_ab_13__9_), .ZN(u5_mult_79_n793) );
  XNOR2_X2 u5_mult_79_U1824 ( .A(u5_mult_79_n793), .B(u5_mult_79_SUMB_12__10_), 
        .ZN(u5_mult_79_SUMB_13__9_) );
  NAND2_X2 u5_mult_79_U1823 ( .A1(u5_mult_79_CARRYB_5__6_), .A2(
        u5_mult_79_SUMB_5__7_), .ZN(u5_mult_79_n885) );
  NAND2_X2 u5_mult_79_U1822 ( .A1(u5_mult_79_ab_6__6_), .A2(
        u5_mult_79_CARRYB_5__6_), .ZN(u5_mult_79_n883) );
  NOR2_X1 u5_mult_79_U1821 ( .A1(u5_mult_79_n1814), .A2(u5_mult_79_n1731), 
        .ZN(u5_mult_79_ab_5__6_) );
  NOR2_X1 u5_mult_79_U1820 ( .A1(u5_mult_79_n1828), .A2(u5_mult_79_n1764), 
        .ZN(u5_mult_79_ab_16__1_) );
  NAND3_X4 u5_mult_79_U1819 ( .A1(u5_mult_79_n790), .A2(u5_mult_79_n791), .A3(
        u5_mult_79_n792), .ZN(u5_mult_79_CARRYB_5__6_) );
  NAND2_X1 u5_mult_79_U1818 ( .A1(u5_mult_79_ab_5__6_), .A2(
        u5_mult_79_CARRYB_4__6_), .ZN(u5_mult_79_n792) );
  NAND2_X2 u5_mult_79_U1817 ( .A1(u5_mult_79_n262), .A2(u5_mult_79_n387), .ZN(
        u5_mult_79_n790) );
  XOR2_X2 u5_mult_79_U1816 ( .A(u5_mult_79_n387), .B(u5_mult_79_n789), .Z(
        u5_mult_79_SUMB_5__6_) );
  NAND3_X2 u5_mult_79_U1815 ( .A1(u5_mult_79_n786), .A2(u5_mult_79_n787), .A3(
        u5_mult_79_n788), .ZN(u5_mult_79_CARRYB_16__1_) );
  NAND2_X1 u5_mult_79_U1814 ( .A1(u5_mult_79_ab_16__1_), .A2(
        u5_mult_79_SUMB_15__2_), .ZN(u5_mult_79_n788) );
  NAND2_X1 u5_mult_79_U1813 ( .A1(u5_mult_79_ab_16__1_), .A2(
        u5_mult_79_CARRYB_15__1_), .ZN(u5_mult_79_n787) );
  NAND2_X1 u5_mult_79_U1812 ( .A1(u5_mult_79_SUMB_15__2_), .A2(
        u5_mult_79_CARRYB_15__1_), .ZN(u5_mult_79_n786) );
  XNOR2_X2 u5_mult_79_U1811 ( .A(u5_mult_79_CARRYB_2__21_), .B(
        u5_mult_79_ab_3__21_), .ZN(u5_mult_79_n785) );
  XNOR2_X2 u5_mult_79_U1810 ( .A(u5_mult_79_n401), .B(u5_mult_79_n785), .ZN(
        u5_mult_79_SUMB_3__21_) );
  XNOR2_X2 u5_mult_79_U1809 ( .A(u5_mult_79_ab_13__12_), .B(
        u5_mult_79_CARRYB_12__12_), .ZN(u5_mult_79_n784) );
  XNOR2_X2 u5_mult_79_U1808 ( .A(u5_mult_79_SUMB_12__13_), .B(u5_mult_79_n784), 
        .ZN(u5_mult_79_SUMB_13__12_) );
  NAND2_X2 u5_mult_79_U1807 ( .A1(u5_mult_79_SUMB_13__16_), .A2(
        u5_mult_79_n442), .ZN(u5_mult_79_n1047) );
  NAND2_X2 u5_mult_79_U1806 ( .A1(u5_mult_79_ab_7__18_), .A2(
        u5_mult_79_CARRYB_6__18_), .ZN(u5_mult_79_n1275) );
  INV_X4 u5_mult_79_U1805 ( .A(u5_mult_79_n782), .ZN(u5_mult_79_n783) );
  INV_X4 u5_mult_79_U1804 ( .A(u5_mult_79_n780), .ZN(u5_mult_79_n781) );
  XNOR2_X2 u5_mult_79_U1803 ( .A(u5_mult_79_n511), .B(u5_mult_79_n779), .ZN(
        u5_mult_79_SUMB_21__2_) );
  NAND2_X2 u5_mult_79_U1802 ( .A1(u5_mult_79_CARRYB_8__15_), .A2(
        u5_mult_79_SUMB_8__16_), .ZN(u5_mult_79_n1211) );
  NAND2_X4 u5_mult_79_U1801 ( .A1(u5_mult_79_ab_18__5_), .A2(
        u5_mult_79_CARRYB_17__5_), .ZN(u5_mult_79_n1201) );
  XNOR2_X2 u5_mult_79_U1800 ( .A(u5_mult_79_CARRYB_6__8_), .B(u5_mult_79_n777), 
        .ZN(u5_mult_79_n1164) );
  XNOR2_X2 u5_mult_79_U1799 ( .A(u5_mult_79_n776), .B(u5_mult_79_SUMB_14__7_), 
        .ZN(u5_mult_79_SUMB_15__6_) );
  NOR2_X1 u5_mult_79_U1798 ( .A1(u5_mult_79_n1832), .A2(u5_mult_79_n1761), 
        .ZN(u5_mult_79_ab_15__23_) );
  NOR2_X1 u5_mult_79_U1797 ( .A1(u5_mult_79_n1781), .A2(u5_mult_79_n1765), 
        .ZN(u5_mult_79_ab_16__22_) );
  NAND3_X2 u5_mult_79_U1796 ( .A1(u5_mult_79_n773), .A2(u5_mult_79_n774), .A3(
        u5_mult_79_n775), .ZN(u5_mult_79_CARRYB_16__22_) );
  NAND2_X2 u5_mult_79_U1795 ( .A1(u5_mult_79_ab_15__23_), .A2(
        u5_mult_79_ab_16__22_), .ZN(u5_mult_79_n775) );
  NAND2_X2 u5_mult_79_U1794 ( .A1(u5_mult_79_ab_15__23_), .A2(
        u5_mult_79_CARRYB_15__22_), .ZN(u5_mult_79_n774) );
  NAND2_X2 u5_mult_79_U1793 ( .A1(u5_mult_79_ab_16__22_), .A2(
        u5_mult_79_CARRYB_15__22_), .ZN(u5_mult_79_n773) );
  XOR2_X1 u5_mult_79_U1792 ( .A(u5_mult_79_CARRYB_15__22_), .B(u5_mult_79_n772), .Z(u5_mult_79_SUMB_16__22_) );
  XOR2_X2 u5_mult_79_U1791 ( .A(u5_mult_79_ab_16__22_), .B(
        u5_mult_79_ab_15__23_), .Z(u5_mult_79_n772) );
  NAND3_X2 u5_mult_79_U1790 ( .A1(u5_mult_79_n1596), .A2(u5_mult_79_n1595), 
        .A3(u5_mult_79_n1594), .ZN(u5_mult_79_CARRYB_18__6_) );
  NOR2_X1 u5_mult_79_U1789 ( .A1(u5_mult_79_n1831), .A2(u5_mult_79_n1749), 
        .ZN(u5_mult_79_ab_11__23_) );
  NOR2_X1 u5_mult_79_U1788 ( .A1(u5_mult_79_n1781), .A2(u5_mult_79_n1753), 
        .ZN(u5_mult_79_ab_12__22_) );
  NAND3_X2 u5_mult_79_U1787 ( .A1(u5_mult_79_n769), .A2(u5_mult_79_n770), .A3(
        u5_mult_79_n771), .ZN(u5_mult_79_CARRYB_12__22_) );
  NAND2_X2 u5_mult_79_U1786 ( .A1(u5_mult_79_ab_11__23_), .A2(
        u5_mult_79_ab_12__22_), .ZN(u5_mult_79_n771) );
  NAND2_X2 u5_mult_79_U1785 ( .A1(u5_mult_79_ab_11__23_), .A2(
        u5_mult_79_CARRYB_11__22_), .ZN(u5_mult_79_n770) );
  NAND2_X2 u5_mult_79_U1784 ( .A1(u5_mult_79_ab_12__22_), .A2(
        u5_mult_79_CARRYB_11__22_), .ZN(u5_mult_79_n769) );
  XOR2_X1 u5_mult_79_U1783 ( .A(u5_mult_79_CARRYB_11__22_), .B(u5_mult_79_n768), .Z(u5_mult_79_SUMB_12__22_) );
  XOR2_X2 u5_mult_79_U1782 ( .A(u5_mult_79_ab_12__22_), .B(
        u5_mult_79_ab_11__23_), .Z(u5_mult_79_n768) );
  NOR2_X1 u5_mult_79_U1781 ( .A1(u5_mult_79_n1868), .A2(u5_mult_79_n1773), 
        .ZN(u5_mult_79_ab_19__13_) );
  NAND3_X2 u5_mult_79_U1780 ( .A1(u5_mult_79_n765), .A2(u5_mult_79_n766), .A3(
        u5_mult_79_n767), .ZN(u5_mult_79_CARRYB_11__18_) );
  NAND2_X2 u5_mult_79_U1779 ( .A1(u5_mult_79_CARRYB_10__18_), .A2(
        u5_mult_79_SUMB_10__19_), .ZN(u5_mult_79_n767) );
  NAND2_X2 u5_mult_79_U1778 ( .A1(u5_mult_79_ab_11__18_), .A2(
        u5_mult_79_SUMB_10__19_), .ZN(u5_mult_79_n766) );
  NAND2_X1 u5_mult_79_U1777 ( .A1(u5_mult_79_ab_11__18_), .A2(
        u5_mult_79_CARRYB_10__18_), .ZN(u5_mult_79_n765) );
  NAND3_X2 u5_mult_79_U1776 ( .A1(u5_mult_79_n762), .A2(u5_mult_79_n763), .A3(
        u5_mult_79_n764), .ZN(u5_mult_79_CARRYB_10__19_) );
  NAND2_X1 u5_mult_79_U1775 ( .A1(u5_mult_79_CARRYB_9__19_), .A2(
        u5_mult_79_SUMB_9__20_), .ZN(u5_mult_79_n764) );
  NAND2_X1 u5_mult_79_U1774 ( .A1(u5_mult_79_ab_10__19_), .A2(
        u5_mult_79_SUMB_9__20_), .ZN(u5_mult_79_n763) );
  NAND2_X2 u5_mult_79_U1773 ( .A1(u5_mult_79_ab_19__13_), .A2(u5_mult_79_n440), 
        .ZN(u5_mult_79_n760) );
  NAND2_X1 u5_mult_79_U1772 ( .A1(u5_mult_79_SUMB_18__14_), .A2(
        u5_mult_79_n396), .ZN(u5_mult_79_n759) );
  NAND3_X4 u5_mult_79_U1771 ( .A1(u5_mult_79_n756), .A2(u5_mult_79_n757), .A3(
        u5_mult_79_n758), .ZN(u5_mult_79_CARRYB_16__15_) );
  NAND2_X2 u5_mult_79_U1770 ( .A1(u5_mult_79_SUMB_15__16_), .A2(
        u5_mult_79_ab_16__15_), .ZN(u5_mult_79_n758) );
  NAND2_X2 u5_mult_79_U1769 ( .A1(u5_mult_79_ab_15__16_), .A2(
        u5_mult_79_SUMB_14__17_), .ZN(u5_mult_79_n755) );
  NAND2_X2 u5_mult_79_U1768 ( .A1(u5_mult_79_ab_4__20_), .A2(
        u5_mult_79_CARRYB_3__20_), .ZN(u5_mult_79_n1605) );
  NAND2_X1 u5_mult_79_U1767 ( .A1(u5_mult_79_CARRYB_3__20_), .A2(
        u5_mult_79_SUMB_3__21_), .ZN(u5_mult_79_n1603) );
  XNOR2_X2 u5_mult_79_U1766 ( .A(u5_mult_79_CARRYB_11__17_), .B(
        u5_mult_79_n752), .ZN(u5_mult_79_n982) );
  NAND2_X1 u5_mult_79_U1765 ( .A1(u5_mult_79_CARRYB_8__17_), .A2(
        u5_mult_79_SUMB_8__18_), .ZN(u5_mult_79_n1375) );
  XNOR2_X2 u5_mult_79_U1764 ( .A(u5_mult_79_n751), .B(u5_mult_79_SUMB_12__9_), 
        .ZN(u5_mult_79_SUMB_13__8_) );
  INV_X4 u5_mult_79_U1763 ( .A(u5_mult_79_ab_18__5_), .ZN(u5_mult_79_n1054) );
  INV_X4 u5_mult_79_U1762 ( .A(u5_mult_79_n1054), .ZN(u5_mult_79_n748) );
  INV_X2 u5_mult_79_U1761 ( .A(u5_mult_79_CARRYB_17__5_), .ZN(u5_mult_79_n747)
         );
  NAND2_X1 u5_mult_79_U1760 ( .A1(u5_mult_79_CARRYB_17__5_), .A2(
        u5_mult_79_n1054), .ZN(u5_mult_79_n749) );
  NAND3_X2 u5_mult_79_U1759 ( .A1(u5_mult_79_n744), .A2(u5_mult_79_n745), .A3(
        u5_mult_79_n746), .ZN(u5_mult_79_CARRYB_5__19_) );
  NAND2_X1 u5_mult_79_U1758 ( .A1(u5_mult_79_SUMB_4__20_), .A2(
        u5_mult_79_ab_5__19_), .ZN(u5_mult_79_n746) );
  NAND2_X2 u5_mult_79_U1757 ( .A1(u5_mult_79_ab_5__19_), .A2(
        u5_mult_79_CARRYB_4__19_), .ZN(u5_mult_79_n745) );
  NAND3_X2 u5_mult_79_U1756 ( .A1(u5_mult_79_n741), .A2(u5_mult_79_n743), .A3(
        u5_mult_79_n742), .ZN(u5_mult_79_CARRYB_12__16_) );
  NAND2_X1 u5_mult_79_U1755 ( .A1(u5_mult_79_ab_12__16_), .A2(
        u5_mult_79_CARRYB_11__16_), .ZN(u5_mult_79_n741) );
  NAND3_X2 u5_mult_79_U1754 ( .A1(u5_mult_79_n738), .A2(u5_mult_79_n739), .A3(
        u5_mult_79_n740), .ZN(u5_mult_79_CARRYB_11__17_) );
  NAND2_X2 u5_mult_79_U1753 ( .A1(u5_mult_79_ab_11__17_), .A2(
        u5_mult_79_SUMB_10__18_), .ZN(u5_mult_79_n739) );
  NAND2_X1 u5_mult_79_U1752 ( .A1(u5_mult_79_ab_11__17_), .A2(
        u5_mult_79_CARRYB_10__17_), .ZN(u5_mult_79_n738) );
  XNOR2_X1 u5_mult_79_U1751 ( .A(u5_mult_79_ab_10__11_), .B(
        u5_mult_79_CARRYB_9__11_), .ZN(u5_mult_79_n737) );
  XNOR2_X2 u5_mult_79_U1750 ( .A(u5_mult_79_n737), .B(u5_mult_79_n450), .ZN(
        u5_mult_79_SUMB_10__11_) );
  NAND3_X4 u5_mult_79_U1749 ( .A1(u5_mult_79_n1289), .A2(u5_mult_79_n1288), 
        .A3(u5_mult_79_n1287), .ZN(u5_mult_79_CARRYB_15__7_) );
  NAND2_X1 u5_mult_79_U1748 ( .A1(u5_mult_79_ab_8__7_), .A2(
        u5_mult_79_CARRYB_7__7_), .ZN(u5_mult_79_n1168) );
  NAND2_X1 u5_mult_79_U1747 ( .A1(u5_mult_79_CARRYB_5__9_), .A2(
        u5_mult_79_SUMB_5__10_), .ZN(u5_mult_79_n871) );
  XNOR2_X2 u5_mult_79_U1746 ( .A(u5_mult_79_CARRYB_18__4_), .B(
        u5_mult_79_ab_19__4_), .ZN(u5_mult_79_n909) );
  NAND2_X2 u5_mult_79_U1745 ( .A1(u5_mult_79_CARRYB_16__11_), .A2(
        u5_mult_79_n454), .ZN(u5_mult_79_n1550) );
  XNOR2_X2 u5_mult_79_U1744 ( .A(u5_mult_79_n1304), .B(u5_mult_79_n258), .ZN(
        u5_mult_79_SUMB_21__1_) );
  NOR2_X1 u5_mult_79_U1743 ( .A1(u5_mult_79_n1806), .A2(u5_mult_79_n1773), 
        .ZN(u5_mult_79_ab_19__9_) );
  NAND2_X1 u5_mult_79_U1742 ( .A1(u5_mult_79_ab_19__9_), .A2(
        u5_mult_79_CARRYB_18__9_), .ZN(u5_mult_79_n736) );
  NAND2_X2 u5_mult_79_U1741 ( .A1(u5_mult_79_ab_19__9_), .A2(
        u5_mult_79_SUMB_18__10_), .ZN(u5_mult_79_n735) );
  NAND2_X1 u5_mult_79_U1740 ( .A1(u5_mult_79_CARRYB_18__9_), .A2(
        u5_mult_79_SUMB_18__10_), .ZN(u5_mult_79_n734) );
  NAND3_X4 u5_mult_79_U1739 ( .A1(u5_mult_79_n733), .A2(u5_mult_79_n732), .A3(
        u5_mult_79_n731), .ZN(u5_mult_79_CARRYB_6__17_) );
  NAND2_X2 u5_mult_79_U1738 ( .A1(u5_mult_79_CARRYB_5__17_), .A2(
        u5_mult_79_n128), .ZN(u5_mult_79_n733) );
  NAND2_X2 u5_mult_79_U1737 ( .A1(u5_mult_79_n128), .A2(u5_mult_79_ab_6__17_), 
        .ZN(u5_mult_79_n732) );
  NAND2_X1 u5_mult_79_U1736 ( .A1(u5_mult_79_ab_6__17_), .A2(
        u5_mult_79_CARRYB_5__17_), .ZN(u5_mult_79_n731) );
  NAND3_X2 u5_mult_79_U1735 ( .A1(u5_mult_79_n728), .A2(u5_mult_79_n729), .A3(
        u5_mult_79_n730), .ZN(u5_mult_79_CARRYB_5__18_) );
  NAND2_X1 u5_mult_79_U1734 ( .A1(u5_mult_79_CARRYB_4__18_), .A2(
        u5_mult_79_SUMB_4__19_), .ZN(u5_mult_79_n730) );
  NAND2_X1 u5_mult_79_U1733 ( .A1(u5_mult_79_ab_5__18_), .A2(
        u5_mult_79_SUMB_4__19_), .ZN(u5_mult_79_n729) );
  NAND2_X1 u5_mult_79_U1732 ( .A1(u5_mult_79_ab_5__18_), .A2(
        u5_mult_79_CARRYB_4__18_), .ZN(u5_mult_79_n728) );
  NAND3_X2 u5_mult_79_U1731 ( .A1(u5_mult_79_n725), .A2(u5_mult_79_n726), .A3(
        u5_mult_79_n727), .ZN(u5_mult_79_CARRYB_13__13_) );
  NAND2_X2 u5_mult_79_U1730 ( .A1(u5_mult_79_n356), .A2(
        u5_mult_79_SUMB_12__14_), .ZN(u5_mult_79_n727) );
  NAND2_X2 u5_mult_79_U1729 ( .A1(u5_mult_79_ab_13__13_), .A2(
        u5_mult_79_SUMB_12__14_), .ZN(u5_mult_79_n726) );
  NAND2_X1 u5_mult_79_U1728 ( .A1(u5_mult_79_ab_13__13_), .A2(
        u5_mult_79_CARRYB_12__13_), .ZN(u5_mult_79_n725) );
  NAND2_X2 u5_mult_79_U1727 ( .A1(u5_mult_79_ab_12__14_), .A2(
        u5_mult_79_SUMB_11__15_), .ZN(u5_mult_79_n723) );
  XOR2_X2 u5_mult_79_U1726 ( .A(u5_mult_79_ab_13__13_), .B(
        u5_mult_79_CARRYB_12__13_), .Z(u5_mult_79_n721) );
  XOR2_X2 u5_mult_79_U1725 ( .A(u5_mult_79_n720), .B(u5_mult_79_SUMB_11__15_), 
        .Z(u5_mult_79_SUMB_12__14_) );
  XOR2_X2 u5_mult_79_U1724 ( .A(u5_mult_79_ab_12__14_), .B(
        u5_mult_79_CARRYB_11__14_), .Z(u5_mult_79_n720) );
  NAND2_X2 u5_mult_79_U1723 ( .A1(u5_mult_79_SUMB_20__2_), .A2(
        u5_mult_79_CARRYB_20__1_), .ZN(u5_mult_79_n1388) );
  XNOR2_X2 u5_mult_79_U1722 ( .A(u5_mult_79_CARRYB_12__19_), .B(
        u5_mult_79_n719), .ZN(u5_mult_79_SUMB_13__19_) );
  NAND2_X2 u5_mult_79_U1721 ( .A1(u5_mult_79_ab_6__14_), .A2(u5_mult_79_n496), 
        .ZN(u5_mult_79_n1413) );
  NAND3_X2 u5_mult_79_U1720 ( .A1(u5_mult_79_n716), .A2(u5_mult_79_n717), .A3(
        u5_mult_79_n718), .ZN(u5_mult_79_CARRYB_3__11_) );
  NAND2_X1 u5_mult_79_U1719 ( .A1(u5_mult_79_ab_3__11_), .A2(
        u5_mult_79_SUMB_2__12_), .ZN(u5_mult_79_n718) );
  NAND2_X1 u5_mult_79_U1718 ( .A1(u5_mult_79_SUMB_2__12_), .A2(u5_mult_79_n288), .ZN(u5_mult_79_n717) );
  NAND2_X1 u5_mult_79_U1717 ( .A1(u5_mult_79_ab_3__11_), .A2(u5_mult_79_n288), 
        .ZN(u5_mult_79_n716) );
  NAND3_X4 u5_mult_79_U1716 ( .A1(u5_mult_79_n713), .A2(u5_mult_79_n714), .A3(
        u5_mult_79_n715), .ZN(u5_mult_79_CARRYB_2__12_) );
  NAND2_X2 u5_mult_79_U1715 ( .A1(u5_mult_79_CARRYB_1__12_), .A2(
        u5_mult_79_SUMB_1__13_), .ZN(u5_mult_79_n715) );
  NAND2_X2 u5_mult_79_U1714 ( .A1(u5_mult_79_ab_2__12_), .A2(
        u5_mult_79_SUMB_1__13_), .ZN(u5_mult_79_n714) );
  NAND2_X2 u5_mult_79_U1713 ( .A1(u5_mult_79_ab_2__12_), .A2(
        u5_mult_79_CARRYB_1__12_), .ZN(u5_mult_79_n713) );
  XOR2_X2 u5_mult_79_U1712 ( .A(u5_mult_79_n712), .B(u5_mult_79_SUMB_2__12_), 
        .Z(u5_mult_79_SUMB_3__11_) );
  XOR2_X2 u5_mult_79_U1711 ( .A(u5_mult_79_n711), .B(u5_mult_79_SUMB_1__13_), 
        .Z(u5_mult_79_SUMB_2__12_) );
  XOR2_X2 u5_mult_79_U1710 ( .A(u5_mult_79_ab_2__12_), .B(
        u5_mult_79_CARRYB_1__12_), .Z(u5_mult_79_n711) );
  NAND2_X1 u5_mult_79_U1709 ( .A1(u5_mult_79_ab_9__7_), .A2(
        u5_mult_79_CARRYB_8__7_), .ZN(u5_mult_79_n708) );
  NAND2_X2 u5_mult_79_U1708 ( .A1(u5_mult_79_CARRYB_7__8_), .A2(
        u5_mult_79_SUMB_7__9_), .ZN(u5_mult_79_n707) );
  NAND2_X2 u5_mult_79_U1707 ( .A1(u5_mult_79_ab_8__8_), .A2(
        u5_mult_79_SUMB_7__9_), .ZN(u5_mult_79_n706) );
  NAND2_X2 u5_mult_79_U1706 ( .A1(u5_mult_79_ab_8__8_), .A2(
        u5_mult_79_CARRYB_7__8_), .ZN(u5_mult_79_n705) );
  XNOR2_X2 u5_mult_79_U1705 ( .A(u5_mult_79_SUMB_12__20_), .B(
        u5_mult_79_ab_13__19_), .ZN(u5_mult_79_n719) );
  NAND2_X2 u5_mult_79_U1704 ( .A1(u5_mult_79_ab_0__22_), .A2(
        u5_mult_79_ab_1__21_), .ZN(u5_mult_79_n1714) );
  INV_X8 u5_mult_79_U1703 ( .A(u5_mult_79_n1866), .ZN(u5_mult_79_n1797) );
  NAND2_X4 u5_mult_79_U1702 ( .A1(u5_mult_79_ab_0__12_), .A2(
        u5_mult_79_ab_1__11_), .ZN(u5_mult_79_n1695) );
  XNOR2_X2 u5_mult_79_U1701 ( .A(u5_mult_79_ab_4__15_), .B(
        u5_mult_79_CARRYB_3__15_), .ZN(u5_mult_79_n778) );
  NAND3_X2 u5_mult_79_U1700 ( .A1(u5_mult_79_n1642), .A2(u5_mult_79_n1643), 
        .A3(u5_mult_79_n1644), .ZN(u5_mult_79_CARRYB_19__7_) );
  NAND2_X2 u5_mult_79_U1699 ( .A1(u5_mult_79_ab_11__9_), .A2(
        u5_mult_79_CARRYB_10__9_), .ZN(u5_mult_79_n989) );
  NAND2_X1 u5_mult_79_U1698 ( .A1(u5_mult_79_ab_7__6_), .A2(
        u5_mult_79_SUMB_6__7_), .ZN(u5_mult_79_n919) );
  NAND3_X1 u5_mult_79_U1697 ( .A1(u5_mult_79_n1603), .A2(u5_mult_79_n1604), 
        .A3(u5_mult_79_n1605), .ZN(u5_mult_79_n969) );
  NOR2_X2 u5_mult_79_U1696 ( .A1(u5_mult_79_n1798), .A2(u5_mult_79_n1738), 
        .ZN(u5_mult_79_ab_7__12_) );
  NAND3_X2 u5_mult_79_U1695 ( .A1(u5_mult_79_n702), .A2(u5_mult_79_n703), .A3(
        u5_mult_79_n704), .ZN(u5_mult_79_CARRYB_7__12_) );
  NAND2_X1 u5_mult_79_U1694 ( .A1(u5_mult_79_ab_7__12_), .A2(
        u5_mult_79_CARRYB_6__12_), .ZN(u5_mult_79_n704) );
  NAND2_X2 u5_mult_79_U1693 ( .A1(u5_mult_79_n9), .A2(u5_mult_79_SUMB_4__13_), 
        .ZN(u5_mult_79_n701) );
  NAND2_X2 u5_mult_79_U1692 ( .A1(u5_mult_79_ab_5__12_), .A2(
        u5_mult_79_SUMB_4__13_), .ZN(u5_mult_79_n700) );
  NAND2_X1 u5_mult_79_U1691 ( .A1(u5_mult_79_ab_5__12_), .A2(
        u5_mult_79_CARRYB_4__12_), .ZN(u5_mult_79_n699) );
  NAND3_X4 u5_mult_79_U1690 ( .A1(u5_mult_79_n696), .A2(u5_mult_79_n697), .A3(
        u5_mult_79_n698), .ZN(u5_mult_79_CARRYB_4__13_) );
  NAND2_X2 u5_mult_79_U1689 ( .A1(u5_mult_79_CARRYB_3__13_), .A2(
        u5_mult_79_SUMB_3__14_), .ZN(u5_mult_79_n698) );
  NAND2_X2 u5_mult_79_U1688 ( .A1(u5_mult_79_ab_4__13_), .A2(
        u5_mult_79_SUMB_3__14_), .ZN(u5_mult_79_n697) );
  NAND2_X1 u5_mult_79_U1687 ( .A1(u5_mult_79_ab_4__13_), .A2(
        u5_mult_79_CARRYB_3__13_), .ZN(u5_mult_79_n696) );
  NAND2_X1 u5_mult_79_U1686 ( .A1(u5_mult_79_SUMB_16__15_), .A2(
        u5_mult_79_CARRYB_16__14_), .ZN(u5_mult_79_n952) );
  NAND2_X1 u5_mult_79_U1685 ( .A1(u5_mult_79_ab_19__13_), .A2(u5_mult_79_n396), 
        .ZN(u5_mult_79_n761) );
  NAND3_X2 u5_mult_79_U1684 ( .A1(u5_mult_79_n563), .A2(u5_mult_79_n693), .A3(
        u5_mult_79_n694), .ZN(u5_mult_79_CARRYB_18__16_) );
  NAND2_X2 u5_mult_79_U1683 ( .A1(u5_mult_79_CARRYB_17__16_), .A2(
        u5_mult_79_SUMB_17__17_), .ZN(u5_mult_79_n694) );
  NAND3_X2 u5_mult_79_U1682 ( .A1(u5_mult_79_n690), .A2(u5_mult_79_n691), .A3(
        u5_mult_79_n692), .ZN(u5_mult_79_CARRYB_17__17_) );
  NAND2_X1 u5_mult_79_U1681 ( .A1(u5_mult_79_CARRYB_16__17_), .A2(
        u5_mult_79_SUMB_16__18_), .ZN(u5_mult_79_n692) );
  NAND2_X1 u5_mult_79_U1680 ( .A1(u5_mult_79_ab_17__17_), .A2(
        u5_mult_79_SUMB_16__18_), .ZN(u5_mult_79_n691) );
  NAND2_X1 u5_mult_79_U1679 ( .A1(u5_mult_79_ab_17__17_), .A2(
        u5_mult_79_CARRYB_16__17_), .ZN(u5_mult_79_n690) );
  XOR2_X2 u5_mult_79_U1678 ( .A(u5_mult_79_n689), .B(u5_mult_79_SUMB_16__18_), 
        .Z(u5_mult_79_SUMB_17__17_) );
  XNOR2_X2 u5_mult_79_U1677 ( .A(u5_mult_79_ab_8__7_), .B(
        u5_mult_79_CARRYB_7__7_), .ZN(u5_mult_79_n688) );
  XNOR2_X2 u5_mult_79_U1676 ( .A(u5_mult_79_CARRYB_6__14_), .B(
        u5_mult_79_ab_7__14_), .ZN(u5_mult_79_n687) );
  XNOR2_X2 u5_mult_79_U1675 ( .A(u5_mult_79_n30), .B(u5_mult_79_n687), .ZN(
        u5_mult_79_SUMB_7__14_) );
  NAND2_X2 u5_mult_79_U1674 ( .A1(u5_mult_79_ab_16__13_), .A2(
        u5_mult_79_SUMB_15__14_), .ZN(u5_mult_79_n1336) );
  NAND2_X2 u5_mult_79_U1673 ( .A1(u5_mult_79_n430), .A2(
        u5_mult_79_SUMB_15__14_), .ZN(u5_mult_79_n1337) );
  NAND2_X1 u5_mult_79_U1672 ( .A1(u5_mult_79_SUMB_6__8_), .A2(
        u5_mult_79_CARRYB_6__7_), .ZN(u5_mult_79_n1016) );
  XNOR2_X2 u5_mult_79_U1671 ( .A(u5_mult_79_CARRYB_10__4_), .B(
        u5_mult_79_ab_11__4_), .ZN(u5_mult_79_n686) );
  NOR2_X2 u5_mult_79_U1670 ( .A1(u5_mult_79_n1811), .A2(u5_mult_79_n1734), 
        .ZN(u5_mult_79_ab_6__7_) );
  NOR2_X1 u5_mult_79_U1669 ( .A1(u5_mult_79_n1828), .A2(u5_mult_79_n1767), 
        .ZN(u5_mult_79_ab_17__1_) );
  NAND3_X2 u5_mult_79_U1668 ( .A1(u5_mult_79_n683), .A2(u5_mult_79_n684), .A3(
        u5_mult_79_n685), .ZN(u5_mult_79_CARRYB_6__7_) );
  NAND2_X1 u5_mult_79_U1667 ( .A1(u5_mult_79_ab_6__7_), .A2(
        u5_mult_79_CARRYB_5__7_), .ZN(u5_mult_79_n685) );
  NAND2_X2 u5_mult_79_U1666 ( .A1(u5_mult_79_ab_6__7_), .A2(
        u5_mult_79_SUMB_5__8_), .ZN(u5_mult_79_n684) );
  NAND2_X2 u5_mult_79_U1665 ( .A1(u5_mult_79_CARRYB_5__7_), .A2(
        u5_mult_79_SUMB_5__8_), .ZN(u5_mult_79_n683) );
  XOR2_X2 u5_mult_79_U1664 ( .A(u5_mult_79_SUMB_5__8_), .B(u5_mult_79_n682), 
        .Z(u5_mult_79_SUMB_6__7_) );
  XOR2_X2 u5_mult_79_U1663 ( .A(u5_mult_79_CARRYB_5__7_), .B(
        u5_mult_79_ab_6__7_), .Z(u5_mult_79_n682) );
  NAND3_X2 u5_mult_79_U1662 ( .A1(u5_mult_79_n679), .A2(u5_mult_79_n680), .A3(
        u5_mult_79_n681), .ZN(u5_mult_79_CARRYB_17__1_) );
  NAND2_X1 u5_mult_79_U1661 ( .A1(u5_mult_79_ab_17__1_), .A2(
        u5_mult_79_CARRYB_16__1_), .ZN(u5_mult_79_n681) );
  NAND2_X1 u5_mult_79_U1660 ( .A1(u5_mult_79_ab_17__1_), .A2(
        u5_mult_79_SUMB_16__2_), .ZN(u5_mult_79_n680) );
  NAND2_X1 u5_mult_79_U1659 ( .A1(u5_mult_79_CARRYB_16__1_), .A2(
        u5_mult_79_SUMB_16__2_), .ZN(u5_mult_79_n679) );
  XOR2_X2 u5_mult_79_U1658 ( .A(u5_mult_79_n383), .B(u5_mult_79_n678), .Z(
        u5_mult_79_SUMB_17__1_) );
  XOR2_X2 u5_mult_79_U1657 ( .A(u5_mult_79_CARRYB_16__1_), .B(
        u5_mult_79_ab_17__1_), .Z(u5_mult_79_n678) );
  NAND2_X1 u5_mult_79_U1656 ( .A1(u5_mult_79_ab_14__4_), .A2(
        u5_mult_79_CARRYB_13__4_), .ZN(u5_mult_79_n675) );
  NAND2_X2 u5_mult_79_U1655 ( .A1(u5_mult_79_SUMB_12__6_), .A2(
        u5_mult_79_CARRYB_12__5_), .ZN(u5_mult_79_n674) );
  NAND2_X2 u5_mult_79_U1654 ( .A1(u5_mult_79_SUMB_12__6_), .A2(
        u5_mult_79_ab_13__5_), .ZN(u5_mult_79_n673) );
  NAND2_X1 u5_mult_79_U1653 ( .A1(u5_mult_79_ab_13__5_), .A2(
        u5_mult_79_CARRYB_12__5_), .ZN(u5_mult_79_n672) );
  XNOR2_X2 u5_mult_79_U1652 ( .A(u5_mult_79_ab_16__8_), .B(
        u5_mult_79_CARRYB_15__8_), .ZN(u5_mult_79_n671) );
  INV_X1 u5_mult_79_U1651 ( .A(u5_mult_79_n1707), .ZN(u5_mult_79_SUMB_1__17_)
         );
  NAND3_X2 u5_mult_79_U1650 ( .A1(u5_mult_79_n970), .A2(u5_mult_79_n971), .A3(
        u5_mult_79_n972), .ZN(u5_mult_79_CARRYB_7__14_) );
  NAND2_X2 u5_mult_79_U1649 ( .A1(u5_mult_79_CARRYB_6__14_), .A2(
        u5_mult_79_SUMB_6__15_), .ZN(u5_mult_79_n970) );
  NAND3_X4 u5_mult_79_U1648 ( .A1(u5_mult_79_n1340), .A2(u5_mult_79_n1341), 
        .A3(u5_mult_79_n1342), .ZN(u5_mult_79_CARRYB_4__14_) );
  XNOR2_X2 u5_mult_79_U1647 ( .A(u5_mult_79_CARRYB_20__6_), .B(u5_mult_79_n670), .ZN(u5_mult_79_n1558) );
  XNOR2_X2 u5_mult_79_U1646 ( .A(u5_mult_79_n442), .B(u5_mult_79_ab_14__15_), 
        .ZN(u5_mult_79_n828) );
  NAND2_X2 u5_mult_79_U1645 ( .A1(u5_mult_79_ab_4__20_), .A2(
        u5_mult_79_SUMB_3__21_), .ZN(u5_mult_79_n1604) );
  XNOR2_X2 u5_mult_79_U1644 ( .A(u5_mult_79_CARRYB_21__6_), .B(
        u5_mult_79_ab_22__6_), .ZN(u5_mult_79_n669) );
  XNOR2_X2 u5_mult_79_U1643 ( .A(u5_mult_79_n376), .B(u5_mult_79_n669), .ZN(
        u5_mult_79_SUMB_22__6_) );
  XNOR2_X2 u5_mult_79_U1642 ( .A(u5_mult_79_CARRYB_4__6_), .B(u5_mult_79_n668), 
        .ZN(u5_mult_79_n789) );
  NOR2_X1 u5_mult_79_U1641 ( .A1(u5_mult_79_n1817), .A2(u5_mult_79_n1731), 
        .ZN(u5_mult_79_ab_5__5_) );
  NAND3_X2 u5_mult_79_U1640 ( .A1(u5_mult_79_n665), .A2(u5_mult_79_n666), .A3(
        u5_mult_79_n667), .ZN(u5_mult_79_CARRYB_14__1_) );
  NAND2_X1 u5_mult_79_U1639 ( .A1(u5_mult_79_SUMB_13__2_), .A2(
        u5_mult_79_CARRYB_13__1_), .ZN(u5_mult_79_n667) );
  NAND2_X2 u5_mult_79_U1638 ( .A1(u5_mult_79_ab_14__1_), .A2(
        u5_mult_79_CARRYB_13__1_), .ZN(u5_mult_79_n666) );
  NAND2_X1 u5_mult_79_U1637 ( .A1(u5_mult_79_ab_14__1_), .A2(
        u5_mult_79_SUMB_13__2_), .ZN(u5_mult_79_n665) );
  XOR2_X1 u5_mult_79_U1636 ( .A(u5_mult_79_ab_14__1_), .B(
        u5_mult_79_SUMB_13__2_), .Z(u5_mult_79_n664) );
  NAND3_X2 u5_mult_79_U1635 ( .A1(u5_mult_79_n661), .A2(u5_mult_79_n662), .A3(
        u5_mult_79_n663), .ZN(u5_mult_79_CARRYB_13__1_) );
  NAND2_X2 u5_mult_79_U1634 ( .A1(u5_mult_79_ab_13__1_), .A2(
        u5_mult_79_SUMB_12__2_), .ZN(u5_mult_79_n663) );
  NAND2_X1 u5_mult_79_U1633 ( .A1(u5_mult_79_CARRYB_12__1_), .A2(
        u5_mult_79_SUMB_12__2_), .ZN(u5_mult_79_n662) );
  NAND2_X1 u5_mult_79_U1632 ( .A1(u5_mult_79_CARRYB_12__1_), .A2(
        u5_mult_79_ab_13__1_), .ZN(u5_mult_79_n661) );
  NAND3_X4 u5_mult_79_U1631 ( .A1(u5_mult_79_n658), .A2(u5_mult_79_n659), .A3(
        u5_mult_79_n660), .ZN(u5_mult_79_CARRYB_19__0_) );
  NAND2_X2 u5_mult_79_U1630 ( .A1(u5_mult_79_ab_19__0_), .A2(u5_mult_79_n250), 
        .ZN(u5_mult_79_n660) );
  NAND2_X2 u5_mult_79_U1629 ( .A1(u5_mult_79_ab_19__0_), .A2(
        u5_mult_79_CARRYB_18__0_), .ZN(u5_mult_79_n659) );
  NAND2_X2 u5_mult_79_U1628 ( .A1(u5_mult_79_n250), .A2(
        u5_mult_79_CARRYB_18__0_), .ZN(u5_mult_79_n658) );
  NAND3_X2 u5_mult_79_U1627 ( .A1(u5_mult_79_n654), .A2(u5_mult_79_n655), .A3(
        u5_mult_79_n656), .ZN(u5_mult_79_CARRYB_21__0_) );
  NAND2_X2 u5_mult_79_U1626 ( .A1(u5_mult_79_SUMB_20__1_), .A2(
        u5_mult_79_CARRYB_20__0_), .ZN(u5_mult_79_n656) );
  NAND2_X2 u5_mult_79_U1625 ( .A1(u5_mult_79_ab_21__0_), .A2(
        u5_mult_79_CARRYB_20__0_), .ZN(u5_mult_79_n655) );
  NAND2_X2 u5_mult_79_U1624 ( .A1(u5_mult_79_SUMB_20__1_), .A2(
        u5_mult_79_ab_21__0_), .ZN(u5_mult_79_n654) );
  NAND3_X2 u5_mult_79_U1623 ( .A1(u5_mult_79_n650), .A2(u5_mult_79_n651), .A3(
        u5_mult_79_n652), .ZN(u5_mult_79_CARRYB_20__0_) );
  NAND2_X1 u5_mult_79_U1622 ( .A1(u5_mult_79_CARRYB_19__0_), .A2(
        u5_mult_79_SUMB_19__1_), .ZN(u5_mult_79_n652) );
  NAND2_X2 u5_mult_79_U1621 ( .A1(u5_mult_79_ab_20__0_), .A2(
        u5_mult_79_CARRYB_19__0_), .ZN(u5_mult_79_n650) );
  XOR2_X1 u5_mult_79_U1620 ( .A(u5_mult_79_n649), .B(u5_mult_79_n343), .Z(
        u5_N20) );
  XOR2_X2 u5_mult_79_U1619 ( .A(u5_mult_79_ab_20__0_), .B(
        u5_mult_79_CARRYB_19__0_), .Z(u5_mult_79_n649) );
  NAND3_X2 u5_mult_79_U1618 ( .A1(u5_mult_79_n646), .A2(u5_mult_79_n647), .A3(
        u5_mult_79_n648), .ZN(u5_mult_79_CARRYB_7__3_) );
  NAND2_X1 u5_mult_79_U1617 ( .A1(u5_mult_79_CARRYB_6__3_), .A2(
        u5_mult_79_SUMB_6__4_), .ZN(u5_mult_79_n648) );
  NAND2_X1 u5_mult_79_U1616 ( .A1(u5_mult_79_ab_7__3_), .A2(
        u5_mult_79_SUMB_6__4_), .ZN(u5_mult_79_n647) );
  NAND2_X1 u5_mult_79_U1615 ( .A1(u5_mult_79_ab_7__3_), .A2(
        u5_mult_79_CARRYB_6__3_), .ZN(u5_mult_79_n646) );
  NAND3_X4 u5_mult_79_U1614 ( .A1(u5_mult_79_n643), .A2(u5_mult_79_n644), .A3(
        u5_mult_79_n645), .ZN(u5_mult_79_CARRYB_6__4_) );
  NAND2_X2 u5_mult_79_U1613 ( .A1(u5_mult_79_CARRYB_5__4_), .A2(
        u5_mult_79_SUMB_5__5_), .ZN(u5_mult_79_n645) );
  NAND2_X2 u5_mult_79_U1612 ( .A1(u5_mult_79_ab_6__4_), .A2(
        u5_mult_79_SUMB_5__5_), .ZN(u5_mult_79_n644) );
  NAND2_X2 u5_mult_79_U1611 ( .A1(u5_mult_79_ab_6__4_), .A2(
        u5_mult_79_CARRYB_5__4_), .ZN(u5_mult_79_n643) );
  XOR2_X2 u5_mult_79_U1610 ( .A(u5_mult_79_n642), .B(u5_mult_79_SUMB_6__4_), 
        .Z(u5_mult_79_SUMB_7__3_) );
  XOR2_X2 u5_mult_79_U1609 ( .A(u5_mult_79_ab_7__3_), .B(
        u5_mult_79_CARRYB_6__3_), .Z(u5_mult_79_n642) );
  XOR2_X2 u5_mult_79_U1608 ( .A(u5_mult_79_n641), .B(u5_mult_79_SUMB_5__5_), 
        .Z(u5_mult_79_SUMB_6__4_) );
  XOR2_X2 u5_mult_79_U1607 ( .A(u5_mult_79_ab_6__4_), .B(
        u5_mult_79_CARRYB_5__4_), .Z(u5_mult_79_n641) );
  NAND3_X2 u5_mult_79_U1606 ( .A1(u5_mult_79_n638), .A2(u5_mult_79_n639), .A3(
        u5_mult_79_n640), .ZN(u5_mult_79_CARRYB_5__5_) );
  NAND2_X1 u5_mult_79_U1605 ( .A1(u5_mult_79_ab_5__5_), .A2(
        u5_mult_79_CARRYB_4__5_), .ZN(u5_mult_79_n640) );
  NAND2_X2 u5_mult_79_U1604 ( .A1(u5_mult_79_ab_5__5_), .A2(
        u5_mult_79_SUMB_4__6_), .ZN(u5_mult_79_n639) );
  NAND2_X1 u5_mult_79_U1603 ( .A1(u5_mult_79_CARRYB_4__5_), .A2(
        u5_mult_79_SUMB_4__6_), .ZN(u5_mult_79_n638) );
  NAND2_X1 u5_mult_79_U1602 ( .A1(u5_mult_79_CARRYB_14__16_), .A2(
        u5_mult_79_ab_15__16_), .ZN(u5_mult_79_n753) );
  XNOR2_X2 u5_mult_79_U1601 ( .A(u5_mult_79_n1303), .B(u5_mult_79_n413), .ZN(
        u5_mult_79_SUMB_22__5_) );
  XNOR2_X2 u5_mult_79_U1600 ( .A(u5_mult_79_n1411), .B(u5_mult_79_n325), .ZN(
        u5_mult_79_SUMB_12__12_) );
  NAND2_X2 u5_mult_79_U1599 ( .A1(u5_mult_79_n23), .A2(u5_mult_79_ab_16__16_), 
        .ZN(u5_mult_79_n1002) );
  XNOR2_X2 u5_mult_79_U1598 ( .A(u5_mult_79_SUMB_12__11_), .B(
        u5_mult_79_ab_13__10_), .ZN(u5_mult_79_n858) );
  NAND2_X2 u5_mult_79_U1597 ( .A1(u5_mult_79_ab_3__21_), .A2(
        u5_mult_79_CARRYB_2__21_), .ZN(u5_mult_79_n1602) );
  NAND3_X2 u5_mult_79_U1596 ( .A1(u5_mult_79_n1626), .A2(u5_mult_79_n1627), 
        .A3(u5_mult_79_n1628), .ZN(u5_mult_79_CARRYB_3__20_) );
  NAND3_X4 u5_mult_79_U1595 ( .A1(u5_mult_79_n1001), .A2(u5_mult_79_n1002), 
        .A3(u5_mult_79_n1003), .ZN(u5_mult_79_CARRYB_16__16_) );
  XNOR2_X2 u5_mult_79_U1594 ( .A(u5_mult_79_ab_5__17_), .B(
        u5_mult_79_CARRYB_4__17_), .ZN(u5_mult_79_n637) );
  XNOR2_X2 u5_mult_79_U1593 ( .A(u5_mult_79_SUMB_4__18_), .B(u5_mult_79_n637), 
        .ZN(u5_mult_79_SUMB_5__17_) );
  NAND2_X2 u5_mult_79_U1592 ( .A1(u5_mult_79_n28), .A2(
        u5_mult_79_CARRYB_6__19_), .ZN(u5_mult_79_n1572) );
  NOR2_X2 u5_mult_79_U1591 ( .A1(u5_mult_79_n1785), .A2(u5_mult_79_n1735), 
        .ZN(u5_mult_79_ab_6__19_) );
  NAND3_X2 u5_mult_79_U1590 ( .A1(u5_mult_79_n634), .A2(u5_mult_79_n635), .A3(
        u5_mult_79_n636), .ZN(u5_mult_79_CARRYB_6__19_) );
  NAND2_X1 u5_mult_79_U1589 ( .A1(u5_mult_79_ab_6__19_), .A2(
        u5_mult_79_CARRYB_5__19_), .ZN(u5_mult_79_n636) );
  NAND2_X2 u5_mult_79_U1588 ( .A1(u5_mult_79_ab_6__19_), .A2(
        u5_mult_79_SUMB_5__20_), .ZN(u5_mult_79_n635) );
  NAND2_X2 u5_mult_79_U1587 ( .A1(u5_mult_79_SUMB_15__16_), .A2(
        u5_mult_79_CARRYB_15__15_), .ZN(u5_mult_79_n757) );
  NAND2_X2 u5_mult_79_U1586 ( .A1(u5_mult_79_ab_17__15_), .A2(
        u5_mult_79_CARRYB_16__15_), .ZN(u5_mult_79_n1136) );
  NAND3_X4 u5_mult_79_U1585 ( .A1(u5_mult_79_n1136), .A2(u5_mult_79_n1137), 
        .A3(u5_mult_79_n1138), .ZN(u5_mult_79_CARRYB_17__15_) );
  XNOR2_X2 u5_mult_79_U1584 ( .A(u5_mult_79_n633), .B(u5_mult_79_SUMB_17__14_), 
        .ZN(u5_mult_79_SUMB_18__13_) );
  NAND2_X2 u5_mult_79_U1583 ( .A1(u5_mult_79_ab_17__11_), .A2(u5_mult_79_n454), 
        .ZN(u5_mult_79_n1549) );
  NAND2_X2 u5_mult_79_U1582 ( .A1(u5_mult_79_n23), .A2(
        u5_mult_79_CARRYB_15__16_), .ZN(u5_mult_79_n1001) );
  XNOR2_X2 u5_mult_79_U1581 ( .A(u5_mult_79_n1031), .B(u5_mult_79_n407), .ZN(
        u5_mult_79_SUMB_6__15_) );
  XOR2_X2 u5_mult_79_U1580 ( .A(u5_mult_79_n1638), .B(u5_mult_79_SUMB_18__8_), 
        .Z(u5_mult_79_SUMB_19__7_) );
  NAND2_X2 u5_mult_79_U1579 ( .A1(u5_mult_79_ab_14__15_), .A2(u5_mult_79_n442), 
        .ZN(u5_mult_79_n1049) );
  NAND3_X2 u5_mult_79_U1578 ( .A1(u5_mult_79_n822), .A2(u5_mult_79_n823), .A3(
        u5_mult_79_n824), .ZN(u5_mult_79_CARRYB_12__15_) );
  XNOR2_X2 u5_mult_79_U1577 ( .A(u5_mult_79_CARRYB_12__11_), .B(
        u5_mult_79_n632), .ZN(u5_mult_79_n1084) );
  NAND2_X2 u5_mult_79_U1576 ( .A1(u5_mult_79_n1524), .A2(
        u5_mult_79_SUMB_13__14_), .ZN(u5_mult_79_n1521) );
  XNOR2_X2 u5_mult_79_U1575 ( .A(u5_mult_79_CARRYB_16__16_), .B(
        u5_mult_79_ab_17__16_), .ZN(u5_mult_79_n631) );
  XNOR2_X2 u5_mult_79_U1574 ( .A(u5_mult_79_n631), .B(u5_mult_79_SUMB_16__17_), 
        .ZN(u5_mult_79_SUMB_17__16_) );
  NAND2_X1 u5_mult_79_U1573 ( .A1(u5_mult_79_ab_8__12_), .A2(
        u5_mult_79_CARRYB_7__12_), .ZN(u5_mult_79_n1485) );
  NAND2_X1 u5_mult_79_U1572 ( .A1(u5_mult_79_SUMB_7__13_), .A2(
        u5_mult_79_CARRYB_7__12_), .ZN(u5_mult_79_n1483) );
  NAND2_X2 u5_mult_79_U1571 ( .A1(u5_mult_79_n322), .A2(
        u5_mult_79_CARRYB_12__10_), .ZN(u5_mult_79_n1408) );
  NOR2_X1 u5_mult_79_U1570 ( .A1(u5_mult_79_n1803), .A2(u5_mult_79_n1752), 
        .ZN(u5_mult_79_ab_12__10_) );
  NAND3_X4 u5_mult_79_U1569 ( .A1(u5_mult_79_n628), .A2(u5_mult_79_n629), .A3(
        u5_mult_79_n630), .ZN(u5_mult_79_CARRYB_12__10_) );
  NAND2_X1 u5_mult_79_U1568 ( .A1(u5_mult_79_ab_12__10_), .A2(
        u5_mult_79_CARRYB_11__10_), .ZN(u5_mult_79_n630) );
  NAND2_X2 u5_mult_79_U1567 ( .A1(u5_mult_79_ab_12__10_), .A2(
        u5_mult_79_SUMB_11__11_), .ZN(u5_mult_79_n629) );
  NAND2_X2 u5_mult_79_U1566 ( .A1(u5_mult_79_CARRYB_11__10_), .A2(
        u5_mult_79_SUMB_11__11_), .ZN(u5_mult_79_n628) );
  NAND2_X2 u5_mult_79_U1565 ( .A1(u5_mult_79_CARRYB_7__14_), .A2(
        u5_mult_79_SUMB_7__15_), .ZN(u5_mult_79_n973) );
  XNOR2_X2 u5_mult_79_U1564 ( .A(u5_mult_79_n892), .B(u5_mult_79_SUMB_9__16_), 
        .ZN(u5_mult_79_SUMB_10__15_) );
  NAND2_X2 u5_mult_79_U1563 ( .A1(u5_mult_79_ab_14__13_), .A2(u5_mult_79_n1524), .ZN(u5_mult_79_n1523) );
  NAND3_X2 u5_mult_79_U1562 ( .A1(u5_mult_79_n1071), .A2(u5_mult_79_n1072), 
        .A3(u5_mult_79_n1073), .ZN(u5_mult_79_CARRYB_14__20_) );
  NAND3_X2 u5_mult_79_U1561 ( .A1(u5_mult_79_n1515), .A2(u5_mult_79_n1516), 
        .A3(u5_mult_79_n1517), .ZN(u5_mult_79_CARRYB_18__11_) );
  XNOR2_X2 u5_mult_79_U1560 ( .A(u5_mult_79_n627), .B(u5_mult_79_CARRYB_14__9_), .ZN(u5_mult_79_n1317) );
  NAND3_X2 u5_mult_79_U1559 ( .A1(u5_mult_79_n1527), .A2(u5_mult_79_n1528), 
        .A3(u5_mult_79_n1529), .ZN(u5_mult_79_CARRYB_3__18_) );
  NAND2_X2 u5_mult_79_U1558 ( .A1(u5_mult_79_CARRYB_2__18_), .A2(
        u5_mult_79_n422), .ZN(u5_mult_79_n1529) );
  INV_X2 u5_mult_79_U1557 ( .A(u5_mult_79_ab_7__20_), .ZN(u5_mult_79_n624) );
  NAND2_X2 u5_mult_79_U1556 ( .A1(u5_mult_79_CARRYB_10__12_), .A2(
        u5_mult_79_SUMB_10__13_), .ZN(u5_mult_79_n1404) );
  NAND3_X4 u5_mult_79_U1555 ( .A1(u5_mult_79_n1412), .A2(u5_mult_79_n1413), 
        .A3(u5_mult_79_n1414), .ZN(u5_mult_79_CARRYB_6__14_) );
  NAND2_X2 u5_mult_79_U1554 ( .A1(u5_mult_79_n850), .A2(u5_mult_79_n851), .ZN(
        u5_mult_79_n1135) );
  INV_X2 u5_mult_79_U1553 ( .A(u5_mult_79_n1554), .ZN(u5_mult_79_n893) );
  NAND3_X2 u5_mult_79_U1552 ( .A1(u5_mult_79_n675), .A2(u5_mult_79_n676), .A3(
        u5_mult_79_n677), .ZN(u5_mult_79_CARRYB_14__4_) );
  NAND2_X2 u5_mult_79_U1551 ( .A1(u5_mult_79_ab_5__20_), .A2(u5_mult_79_n969), 
        .ZN(u5_mult_79_n1152) );
  NAND2_X2 u5_mult_79_U1550 ( .A1(u5_mult_79_ab_15__15_), .A2(
        u5_mult_79_SUMB_14__16_), .ZN(u5_mult_79_n1440) );
  NAND2_X2 u5_mult_79_U1549 ( .A1(u5_mult_79_CARRYB_14__15_), .A2(
        u5_mult_79_SUMB_14__16_), .ZN(u5_mult_79_n1441) );
  XNOR2_X2 u5_mult_79_U1548 ( .A(u5_mult_79_ab_6__21_), .B(
        u5_mult_79_CARRYB_5__21_), .ZN(u5_mult_79_n621) );
  XNOR2_X2 u5_mult_79_U1547 ( .A(u5_mult_79_n621), .B(u5_mult_79_n436), .ZN(
        u5_mult_79_SUMB_6__21_) );
  NAND3_X4 u5_mult_79_U1546 ( .A1(u5_mult_79_n1548), .A2(u5_mult_79_n1549), 
        .A3(u5_mult_79_n1550), .ZN(u5_mult_79_CARRYB_17__11_) );
  XNOR2_X2 u5_mult_79_U1545 ( .A(u5_mult_79_CARRYB_16__12_), .B(
        u5_mult_79_ab_17__12_), .ZN(u5_mult_79_n620) );
  XNOR2_X2 u5_mult_79_U1544 ( .A(u5_mult_79_SUMB_16__13_), .B(u5_mult_79_n620), 
        .ZN(u5_mult_79_SUMB_17__12_) );
  NAND2_X2 u5_mult_79_U1543 ( .A1(u5_mult_79_CARRYB_14__19_), .A2(
        u5_mult_79_SUMB_14__20_), .ZN(u5_mult_79_n1076) );
  NAND3_X2 u5_mult_79_U1542 ( .A1(u5_mult_79_n753), .A2(u5_mult_79_n754), .A3(
        u5_mult_79_n755), .ZN(u5_mult_79_CARRYB_15__16_) );
  NAND2_X2 u5_mult_79_U1541 ( .A1(u5_mult_79_n166), .A2(
        u5_mult_79_SUMB_14__17_), .ZN(u5_mult_79_n754) );
  XNOR2_X2 u5_mult_79_U1540 ( .A(u5_mult_79_CARRYB_4__21_), .B(
        u5_mult_79_ab_5__21_), .ZN(u5_mult_79_n618) );
  XNOR2_X2 u5_mult_79_U1539 ( .A(u5_mult_79_n282), .B(u5_mult_79_n618), .ZN(
        u5_mult_79_SUMB_5__21_) );
  NAND3_X4 u5_mult_79_U1538 ( .A1(u5_mult_79_n1439), .A2(u5_mult_79_n1440), 
        .A3(u5_mult_79_n1441), .ZN(u5_mult_79_CARRYB_15__15_) );
  NAND2_X4 u5_mult_79_U1537 ( .A1(u5_mult_79_CARRYB_15__15_), .A2(
        u5_mult_79_ab_16__15_), .ZN(u5_mult_79_n756) );
  NAND2_X1 u5_mult_79_U1536 ( .A1(u5_mult_79_ab_9__16_), .A2(
        u5_mult_79_SUMB_8__17_), .ZN(u5_mult_79_n1270) );
  NAND2_X1 u5_mult_79_U1535 ( .A1(u5_mult_79_ab_9__16_), .A2(
        u5_mult_79_CARRYB_8__16_), .ZN(u5_mult_79_n1269) );
  INV_X4 u5_mult_79_U1534 ( .A(u5_mult_79_n616), .ZN(u5_mult_79_n617) );
  NAND2_X2 u5_mult_79_U1533 ( .A1(u5_mult_79_n1270), .A2(u5_mult_79_n1271), 
        .ZN(u5_mult_79_n616) );
  NAND3_X4 u5_mult_79_U1532 ( .A1(u5_mult_79_n613), .A2(u5_mult_79_n614), .A3(
        u5_mult_79_n615), .ZN(u5_mult_79_CARRYB_7__17_) );
  NAND2_X2 u5_mult_79_U1531 ( .A1(u5_mult_79_ab_7__17_), .A2(
        u5_mult_79_SUMB_6__18_), .ZN(u5_mult_79_n614) );
  NAND3_X4 u5_mult_79_U1530 ( .A1(u5_mult_79_n612), .A2(u5_mult_79_n611), .A3(
        u5_mult_79_n610), .ZN(u5_mult_79_CARRYB_6__18_) );
  NAND2_X1 u5_mult_79_U1529 ( .A1(u5_mult_79_ab_6__18_), .A2(
        u5_mult_79_CARRYB_5__18_), .ZN(u5_mult_79_n610) );
  INV_X1 u5_mult_79_U1528 ( .A(u5_mult_79_CARRYB_7__17_), .ZN(u5_mult_79_n607)
         );
  INV_X1 u5_mult_79_U1527 ( .A(u5_mult_79_ab_8__17_), .ZN(u5_mult_79_n606) );
  NAND2_X2 u5_mult_79_U1526 ( .A1(u5_mult_79_n608), .A2(u5_mult_79_n609), .ZN(
        u5_mult_79_n1083) );
  NAND2_X2 u5_mult_79_U1525 ( .A1(u5_mult_79_n606), .A2(u5_mult_79_n607), .ZN(
        u5_mult_79_n609) );
  NAND2_X1 u5_mult_79_U1524 ( .A1(u5_mult_79_ab_8__17_), .A2(
        u5_mult_79_CARRYB_7__17_), .ZN(u5_mult_79_n608) );
  NAND3_X2 u5_mult_79_U1523 ( .A1(u5_mult_79_n603), .A2(u5_mult_79_n604), .A3(
        u5_mult_79_n605), .ZN(u5_mult_79_CARRYB_8__21_) );
  NAND2_X2 u5_mult_79_U1522 ( .A1(u5_mult_79_ab_8__21_), .A2(
        u5_mult_79_SUMB_7__22_), .ZN(u5_mult_79_n604) );
  NAND2_X2 u5_mult_79_U1521 ( .A1(u5_mult_79_CARRYB_20__14_), .A2(
        u5_mult_79_SUMB_20__15_), .ZN(u5_mult_79_n602) );
  NAND2_X2 u5_mult_79_U1520 ( .A1(u5_mult_79_ab_21__14_), .A2(
        u5_mult_79_SUMB_20__15_), .ZN(u5_mult_79_n601) );
  NAND2_X1 u5_mult_79_U1519 ( .A1(u5_mult_79_ab_21__14_), .A2(
        u5_mult_79_CARRYB_20__14_), .ZN(u5_mult_79_n600) );
  NAND3_X2 u5_mult_79_U1518 ( .A1(u5_mult_79_n597), .A2(u5_mult_79_n598), .A3(
        u5_mult_79_n599), .ZN(u5_mult_79_CARRYB_20__15_) );
  NAND2_X2 u5_mult_79_U1517 ( .A1(u5_mult_79_ab_20__15_), .A2(
        u5_mult_79_SUMB_19__16_), .ZN(u5_mult_79_n598) );
  NAND2_X1 u5_mult_79_U1516 ( .A1(u5_mult_79_ab_20__15_), .A2(
        u5_mult_79_CARRYB_19__15_), .ZN(u5_mult_79_n597) );
  XOR2_X2 u5_mult_79_U1515 ( .A(u5_mult_79_n596), .B(u5_mult_79_SUMB_20__15_), 
        .Z(u5_mult_79_SUMB_21__14_) );
  XOR2_X2 u5_mult_79_U1514 ( .A(u5_mult_79_CARRYB_20__14_), .B(
        u5_mult_79_ab_21__14_), .Z(u5_mult_79_n596) );
  NAND2_X2 u5_mult_79_U1513 ( .A1(u5_mult_79_ab_3__14_), .A2(
        u5_mult_79_SUMB_2__15_), .ZN(u5_mult_79_n1249) );
  NAND2_X1 u5_mult_79_U1512 ( .A1(u5_mult_79_SUMB_5__20_), .A2(
        u5_mult_79_CARRYB_5__19_), .ZN(u5_mult_79_n634) );
  NAND2_X2 u5_mult_79_U1511 ( .A1(u5_mult_79_CARRYB_8__7_), .A2(
        u5_mult_79_SUMB_8__8_), .ZN(u5_mult_79_n710) );
  NAND2_X4 u5_mult_79_U1510 ( .A1(u5_mult_79_n749), .A2(u5_mult_79_n750), .ZN(
        u5_mult_79_n1198) );
  XOR2_X2 u5_mult_79_U1509 ( .A(u5_mult_79_n275), .B(u5_mult_79_n1575), .Z(
        u5_mult_79_SUMB_16__6_) );
  XNOR2_X2 u5_mult_79_U1508 ( .A(u5_mult_79_CARRYB_8__14_), .B(
        u5_mult_79_ab_9__14_), .ZN(u5_mult_79_n594) );
  XNOR2_X2 u5_mult_79_U1507 ( .A(u5_mult_79_n29), .B(u5_mult_79_n594), .ZN(
        u5_mult_79_SUMB_9__14_) );
  NAND2_X2 u5_mult_79_U1506 ( .A1(u5_mult_79_SUMB_14__8_), .A2(
        u5_mult_79_ab_15__7_), .ZN(u5_mult_79_n1289) );
  NAND3_X4 u5_mult_79_U1505 ( .A1(u5_mult_79_n1629), .A2(u5_mult_79_n1630), 
        .A3(u5_mult_79_n1631), .ZN(u5_mult_79_CARRYB_4__19_) );
  NAND2_X2 u5_mult_79_U1504 ( .A1(u5_mult_79_CARRYB_4__19_), .A2(
        u5_mult_79_SUMB_4__20_), .ZN(u5_mult_79_n744) );
  NAND2_X2 u5_mult_79_U1503 ( .A1(u5_mult_79_ab_15__19_), .A2(
        u5_mult_79_CARRYB_14__19_), .ZN(u5_mult_79_n1074) );
  NAND2_X2 u5_mult_79_U1502 ( .A1(u5_mult_79_ab_5__10_), .A2(u5_mult_79_n872), 
        .ZN(u5_mult_79_n866) );
  NAND2_X2 u5_mult_79_U1501 ( .A1(u5_mult_79_n872), .A2(u5_mult_79_SUMB_4__11_), .ZN(u5_mult_79_n868) );
  NAND3_X2 u5_mult_79_U1500 ( .A1(u5_mult_79_n591), .A2(u5_mult_79_n592), .A3(
        u5_mult_79_n593), .ZN(u5_mult_79_CARRYB_3__17_) );
  NAND2_X1 u5_mult_79_U1499 ( .A1(u5_mult_79_ab_3__17_), .A2(u5_mult_79_n266), 
        .ZN(u5_mult_79_n591) );
  NAND3_X4 u5_mult_79_U1498 ( .A1(u5_mult_79_n588), .A2(u5_mult_79_n589), .A3(
        u5_mult_79_n590), .ZN(u5_mult_79_CARRYB_2__18_) );
  NAND2_X2 u5_mult_79_U1497 ( .A1(u5_mult_79_CARRYB_1__18_), .A2(
        u5_mult_79_SUMB_1__19_), .ZN(u5_mult_79_n590) );
  NAND2_X2 u5_mult_79_U1496 ( .A1(u5_mult_79_ab_2__18_), .A2(
        u5_mult_79_SUMB_1__19_), .ZN(u5_mult_79_n589) );
  NAND2_X2 u5_mult_79_U1495 ( .A1(u5_mult_79_ab_2__18_), .A2(
        u5_mult_79_CARRYB_1__18_), .ZN(u5_mult_79_n588) );
  XOR2_X2 u5_mult_79_U1494 ( .A(u5_mult_79_CARRYB_2__17_), .B(
        u5_mult_79_ab_3__17_), .Z(u5_mult_79_n587) );
  XOR2_X2 u5_mult_79_U1493 ( .A(u5_mult_79_n586), .B(u5_mult_79_SUMB_1__19_), 
        .Z(u5_mult_79_SUMB_2__18_) );
  XOR2_X2 u5_mult_79_U1492 ( .A(u5_mult_79_ab_2__18_), .B(
        u5_mult_79_CARRYB_1__18_), .Z(u5_mult_79_n586) );
  NAND2_X2 u5_mult_79_U1491 ( .A1(u5_mult_79_CARRYB_21__3_), .A2(
        u5_mult_79_SUMB_21__4_), .ZN(u5_mult_79_n585) );
  NAND2_X2 u5_mult_79_U1490 ( .A1(u5_mult_79_ab_22__3_), .A2(
        u5_mult_79_SUMB_21__4_), .ZN(u5_mult_79_n584) );
  NAND3_X2 u5_mult_79_U1489 ( .A1(u5_mult_79_n580), .A2(u5_mult_79_n581), .A3(
        u5_mult_79_n582), .ZN(u5_mult_79_CARRYB_21__4_) );
  NAND2_X2 u5_mult_79_U1488 ( .A1(u5_mult_79_ab_21__4_), .A2(u5_mult_79_n420), 
        .ZN(u5_mult_79_n582) );
  NAND2_X2 u5_mult_79_U1487 ( .A1(u5_mult_79_n111), .A2(u5_mult_79_n420), .ZN(
        u5_mult_79_n581) );
  NAND2_X1 u5_mult_79_U1486 ( .A1(u5_mult_79_n111), .A2(u5_mult_79_ab_21__4_), 
        .ZN(u5_mult_79_n580) );
  NAND2_X1 u5_mult_79_U1485 ( .A1(u5_mult_79_CARRYB_19__3_), .A2(
        u5_mult_79_SUMB_19__4_), .ZN(u5_mult_79_n1632) );
  XNOR2_X2 u5_mult_79_U1484 ( .A(u5_mult_79_CARRYB_18__13_), .B(
        u5_mult_79_ab_19__13_), .ZN(u5_mult_79_n579) );
  XNOR2_X2 u5_mult_79_U1483 ( .A(u5_mult_79_n440), .B(u5_mult_79_n579), .ZN(
        u5_mult_79_SUMB_19__13_) );
  NAND3_X2 u5_mult_79_U1482 ( .A1(u5_mult_79_n1379), .A2(u5_mult_79_n1378), 
        .A3(u5_mult_79_n1377), .ZN(u5_mult_79_CARRYB_3__16_) );
  XNOR2_X2 u5_mult_79_U1481 ( .A(u5_mult_79_n577), .B(u5_mult_79_n437), .ZN(
        u5_mult_79_SUMB_19__12_) );
  NAND2_X2 u5_mult_79_U1480 ( .A1(u5_mult_79_ab_21__2_), .A2(
        u5_mult_79_CARRYB_20__2_), .ZN(u5_mult_79_n1030) );
  NAND2_X2 u5_mult_79_U1479 ( .A1(u5_mult_79_ab_6__12_), .A2(
        u5_mult_79_CARRYB_5__12_), .ZN(u5_mult_79_n1124) );
  NAND3_X4 u5_mult_79_U1478 ( .A1(u5_mult_79_n1124), .A2(u5_mult_79_n1125), 
        .A3(u5_mult_79_n1126), .ZN(u5_mult_79_CARRYB_6__12_) );
  XOR2_X2 u5_mult_79_U1477 ( .A(u5_mult_79_CARRYB_12__18_), .B(
        u5_mult_79_ab_13__18_), .Z(u5_mult_79_n1232) );
  NAND2_X2 u5_mult_79_U1476 ( .A1(u5_mult_79_CARRYB_16__16_), .A2(
        u5_mult_79_SUMB_16__17_), .ZN(u5_mult_79_n1004) );
  NAND2_X2 u5_mult_79_U1475 ( .A1(u5_mult_79_CARRYB_5__21_), .A2(
        u5_mult_79_n436), .ZN(u5_mult_79_n1228) );
  NAND3_X4 u5_mult_79_U1474 ( .A1(u5_mult_79_n1226), .A2(u5_mult_79_n1227), 
        .A3(u5_mult_79_n1228), .ZN(u5_mult_79_CARRYB_6__21_) );
  NAND2_X2 u5_mult_79_U1473 ( .A1(u5_mult_79_SUMB_18__3_), .A2(
        u5_mult_79_CARRYB_18__2_), .ZN(u5_mult_79_n1025) );
  INV_X8 u5_mult_79_U1472 ( .A(n2921), .ZN(u5_mult_79_n1871) );
  NAND2_X2 u5_mult_79_U1471 ( .A1(u5_mult_79_ab_18__16_), .A2(
        u5_mult_79_SUMB_17__17_), .ZN(u5_mult_79_n693) );
  NAND2_X1 u5_mult_79_U1470 ( .A1(u5_mult_79_CARRYB_22__0_), .A2(
        u5_mult_79_ab_23__0_), .ZN(u5_mult_79_n1173) );
  NAND2_X1 u5_mult_79_U1469 ( .A1(u5_mult_79_CARRYB_22__0_), .A2(
        u5_mult_79_n253), .ZN(u5_mult_79_n1172) );
  NAND2_X2 u5_mult_79_U1468 ( .A1(u5_mult_79_n4), .A2(u5_mult_79_ab_11__20_), 
        .ZN(u5_mult_79_n1145) );
  NAND2_X2 u5_mult_79_U1467 ( .A1(u5_mult_79_n4), .A2(
        u5_mult_79_CARRYB_10__20_), .ZN(u5_mult_79_n1147) );
  NAND2_X1 u5_mult_79_U1466 ( .A1(u5_mult_79_CARRYB_17__15_), .A2(
        u5_mult_79_SUMB_17__16_), .ZN(u5_mult_79_n1007) );
  XNOR2_X2 u5_mult_79_U1465 ( .A(u5_mult_79_CARRYB_18__15_), .B(
        u5_mult_79_n575), .ZN(u5_mult_79_n1010) );
  NAND2_X1 u5_mult_79_U1464 ( .A1(u5_mult_79_CARRYB_3__18_), .A2(
        u5_mult_79_SUMB_3__19_), .ZN(u5_mult_79_n1579) );
  NAND2_X2 u5_mult_79_U1463 ( .A1(u5_mult_79_ab_9__7_), .A2(
        u5_mult_79_SUMB_8__8_), .ZN(u5_mult_79_n709) );
  NAND2_X2 u5_mult_79_U1462 ( .A1(u5_mult_79_ab_16__4_), .A2(
        u5_mult_79_SUMB_15__5_), .ZN(u5_mult_79_n1502) );
  XOR2_X2 u5_mult_79_U1461 ( .A(u5_mult_79_ab_15__19_), .B(
        u5_mult_79_CARRYB_14__19_), .Z(u5_mult_79_n1070) );
  NOR2_X1 u5_mult_79_U1460 ( .A1(u5_mult_79_n1785), .A2(u5_mult_79_n1759), 
        .ZN(u5_mult_79_ab_14__19_) );
  NAND3_X4 u5_mult_79_U1459 ( .A1(u5_mult_79_n572), .A2(u5_mult_79_n573), .A3(
        u5_mult_79_n574), .ZN(u5_mult_79_CARRYB_16__17_) );
  NAND2_X2 u5_mult_79_U1458 ( .A1(u5_mult_79_n130), .A2(
        u5_mult_79_SUMB_15__18_), .ZN(u5_mult_79_n574) );
  NAND2_X2 u5_mult_79_U1457 ( .A1(u5_mult_79_ab_16__17_), .A2(
        u5_mult_79_SUMB_15__18_), .ZN(u5_mult_79_n573) );
  NAND3_X2 u5_mult_79_U1456 ( .A1(u5_mult_79_n569), .A2(u5_mult_79_n570), .A3(
        u5_mult_79_n571), .ZN(u5_mult_79_CARRYB_15__18_) );
  NAND2_X1 u5_mult_79_U1455 ( .A1(u5_mult_79_ab_15__18_), .A2(
        u5_mult_79_SUMB_14__19_), .ZN(u5_mult_79_n571) );
  NAND2_X1 u5_mult_79_U1454 ( .A1(u5_mult_79_CARRYB_14__18_), .A2(
        u5_mult_79_SUMB_14__19_), .ZN(u5_mult_79_n570) );
  NAND2_X1 u5_mult_79_U1453 ( .A1(u5_mult_79_CARRYB_14__18_), .A2(
        u5_mult_79_ab_15__18_), .ZN(u5_mult_79_n569) );
  XOR2_X2 u5_mult_79_U1452 ( .A(u5_mult_79_n568), .B(u5_mult_79_SUMB_14__19_), 
        .Z(u5_mult_79_SUMB_15__18_) );
  XOR2_X2 u5_mult_79_U1451 ( .A(u5_mult_79_CARRYB_14__18_), .B(
        u5_mult_79_ab_15__18_), .Z(u5_mult_79_n568) );
  NAND3_X2 u5_mult_79_U1450 ( .A1(u5_mult_79_n565), .A2(u5_mult_79_n566), .A3(
        u5_mult_79_n567), .ZN(u5_mult_79_CARRYB_14__19_) );
  NAND2_X1 u5_mult_79_U1449 ( .A1(u5_mult_79_ab_14__19_), .A2(
        u5_mult_79_CARRYB_13__19_), .ZN(u5_mult_79_n567) );
  NAND2_X2 u5_mult_79_U1448 ( .A1(u5_mult_79_ab_14__19_), .A2(
        u5_mult_79_SUMB_13__20_), .ZN(u5_mult_79_n566) );
  NAND2_X2 u5_mult_79_U1447 ( .A1(u5_mult_79_CARRYB_13__19_), .A2(
        u5_mult_79_SUMB_13__20_), .ZN(u5_mult_79_n565) );
  INV_X4 u5_mult_79_U1446 ( .A(u5_mult_79_CARRYB_17__16_), .ZN(u5_mult_79_n562) );
  INV_X1 u5_mult_79_U1445 ( .A(u5_mult_79_ab_18__16_), .ZN(u5_mult_79_n561) );
  NAND2_X2 u5_mult_79_U1444 ( .A1(u5_mult_79_n563), .A2(u5_mult_79_n564), .ZN(
        u5_mult_79_n619) );
  NAND2_X2 u5_mult_79_U1443 ( .A1(u5_mult_79_n561), .A2(u5_mult_79_n562), .ZN(
        u5_mult_79_n564) );
  NAND3_X4 u5_mult_79_U1442 ( .A1(u5_mult_79_n1388), .A2(u5_mult_79_n1387), 
        .A3(u5_mult_79_n1386), .ZN(u5_mult_79_CARRYB_21__1_) );
  INV_X4 u5_mult_79_U1441 ( .A(u5_mult_79_CARRYB_17__9_), .ZN(u5_mult_79_n558)
         );
  NAND2_X2 u5_mult_79_U1440 ( .A1(u5_mult_79_n1514), .A2(
        u5_mult_79_CARRYB_17__9_), .ZN(u5_mult_79_n559) );
  NOR2_X1 u5_mult_79_U1439 ( .A1(u5_mult_79_n1785), .A2(u5_mult_79_n1776), 
        .ZN(u5_mult_79_ab_20__19_) );
  NAND3_X2 u5_mult_79_U1438 ( .A1(u5_mult_79_n555), .A2(u5_mult_79_n556), .A3(
        u5_mult_79_n557), .ZN(u5_mult_79_CARRYB_22__17_) );
  NAND2_X1 u5_mult_79_U1437 ( .A1(u5_mult_79_CARRYB_21__17_), .A2(
        u5_mult_79_SUMB_21__18_), .ZN(u5_mult_79_n557) );
  NAND2_X1 u5_mult_79_U1436 ( .A1(u5_mult_79_ab_22__17_), .A2(
        u5_mult_79_SUMB_21__18_), .ZN(u5_mult_79_n556) );
  NAND2_X1 u5_mult_79_U1435 ( .A1(u5_mult_79_ab_22__17_), .A2(
        u5_mult_79_CARRYB_21__17_), .ZN(u5_mult_79_n555) );
  NAND3_X2 u5_mult_79_U1434 ( .A1(u5_mult_79_n552), .A2(u5_mult_79_n553), .A3(
        u5_mult_79_n554), .ZN(u5_mult_79_CARRYB_21__18_) );
  NAND2_X1 u5_mult_79_U1433 ( .A1(u5_mult_79_ab_21__18_), .A2(
        u5_mult_79_SUMB_20__19_), .ZN(u5_mult_79_n554) );
  NAND2_X1 u5_mult_79_U1432 ( .A1(u5_mult_79_CARRYB_20__18_), .A2(
        u5_mult_79_SUMB_20__19_), .ZN(u5_mult_79_n553) );
  NAND2_X1 u5_mult_79_U1431 ( .A1(u5_mult_79_CARRYB_20__18_), .A2(
        u5_mult_79_ab_21__18_), .ZN(u5_mult_79_n552) );
  XOR2_X2 u5_mult_79_U1430 ( .A(u5_mult_79_n551), .B(u5_mult_79_SUMB_21__18_), 
        .Z(u5_mult_79_SUMB_22__17_) );
  XOR2_X2 u5_mult_79_U1429 ( .A(u5_mult_79_ab_22__17_), .B(
        u5_mult_79_CARRYB_21__17_), .Z(u5_mult_79_n551) );
  XOR2_X2 u5_mult_79_U1428 ( .A(u5_mult_79_n550), .B(u5_mult_79_SUMB_20__19_), 
        .Z(u5_mult_79_SUMB_21__18_) );
  XOR2_X2 u5_mult_79_U1427 ( .A(u5_mult_79_CARRYB_20__18_), .B(
        u5_mult_79_ab_21__18_), .Z(u5_mult_79_n550) );
  NAND3_X2 u5_mult_79_U1426 ( .A1(u5_mult_79_n547), .A2(u5_mult_79_n548), .A3(
        u5_mult_79_n549), .ZN(u5_mult_79_CARRYB_20__19_) );
  NAND2_X1 u5_mult_79_U1425 ( .A1(u5_mult_79_ab_20__19_), .A2(
        u5_mult_79_CARRYB_19__19_), .ZN(u5_mult_79_n549) );
  NAND2_X2 u5_mult_79_U1424 ( .A1(u5_mult_79_ab_20__19_), .A2(
        u5_mult_79_SUMB_19__20_), .ZN(u5_mult_79_n548) );
  NAND2_X1 u5_mult_79_U1423 ( .A1(u5_mult_79_CARRYB_19__19_), .A2(
        u5_mult_79_SUMB_19__20_), .ZN(u5_mult_79_n547) );
  XOR2_X2 u5_mult_79_U1422 ( .A(u5_mult_79_SUMB_19__20_), .B(u5_mult_79_n546), 
        .Z(u5_mult_79_SUMB_20__19_) );
  XOR2_X2 u5_mult_79_U1421 ( .A(u5_mult_79_CARRYB_19__19_), .B(
        u5_mult_79_ab_20__19_), .Z(u5_mult_79_n546) );
  XNOR2_X2 u5_mult_79_U1420 ( .A(u5_mult_79_CARRYB_4__12_), .B(u5_mult_79_n545), .ZN(u5_mult_79_n695) );
  NAND2_X2 u5_mult_79_U1419 ( .A1(u5_mult_79_ab_20__1_), .A2(u5_mult_79_n492), 
        .ZN(u5_mult_79_n1383) );
  NAND2_X2 u5_mult_79_U1418 ( .A1(u5_mult_79_ab_14__4_), .A2(
        u5_mult_79_SUMB_13__5_), .ZN(u5_mult_79_n676) );
  NAND3_X2 u5_mult_79_U1417 ( .A1(u5_mult_79_n1392), .A2(u5_mult_79_n1393), 
        .A3(u5_mult_79_n1394), .ZN(u5_mult_79_CARRYB_13__12_) );
  XNOR2_X2 u5_mult_79_U1416 ( .A(u5_mult_79_n544), .B(u5_mult_79_n121), .ZN(
        u5_mult_79_SUMB_16__3_) );
  NAND2_X2 u5_mult_79_U1415 ( .A1(u5_mult_79_SUMB_14__8_), .A2(
        u5_mult_79_CARRYB_14__7_), .ZN(u5_mult_79_n1288) );
  NAND2_X2 u5_mult_79_U1414 ( .A1(u5_mult_79_CARRYB_15__7_), .A2(
        u5_mult_79_SUMB_15__8_), .ZN(u5_mult_79_n1482) );
  XNOR2_X2 u5_mult_79_U1413 ( .A(u5_mult_79_CARRYB_20__7_), .B(u5_mult_79_n543), .ZN(u5_mult_79_n812) );
  XNOR2_X2 u5_mult_79_U1412 ( .A(u5_mult_79_n27), .B(u5_mult_79_ab_7__13_), 
        .ZN(u5_mult_79_n542) );
  NOR2_X1 u5_mult_79_U1411 ( .A1(u5_mult_79_n1831), .A2(u5_mult_79_n1743), 
        .ZN(u5_mult_79_ab_9__23_) );
  NOR2_X1 u5_mult_79_U1410 ( .A1(u5_mult_79_n1780), .A2(u5_mult_79_n1747), 
        .ZN(u5_mult_79_ab_10__22_) );
  INV_X4 u5_mult_79_U1409 ( .A(u5_mult_79_n1880), .ZN(u5_mult_79_n1833) );
  NAND3_X2 u5_mult_79_U1408 ( .A1(u5_mult_79_n539), .A2(u5_mult_79_n540), .A3(
        u5_mult_79_n541), .ZN(u5_mult_79_CARRYB_10__22_) );
  NAND2_X2 u5_mult_79_U1407 ( .A1(u5_mult_79_ab_9__23_), .A2(
        u5_mult_79_ab_10__22_), .ZN(u5_mult_79_n541) );
  NAND2_X2 u5_mult_79_U1406 ( .A1(u5_mult_79_n212), .A2(u5_mult_79_ab_9__23_), 
        .ZN(u5_mult_79_n540) );
  NAND2_X2 u5_mult_79_U1405 ( .A1(u5_mult_79_ab_10__22_), .A2(u5_mult_79_n212), 
        .ZN(u5_mult_79_n539) );
  XOR2_X1 u5_mult_79_U1404 ( .A(u5_mult_79_n212), .B(u5_mult_79_n538), .Z(
        u5_mult_79_SUMB_10__22_) );
  XOR2_X2 u5_mult_79_U1403 ( .A(u5_mult_79_ab_10__22_), .B(
        u5_mult_79_ab_9__23_), .Z(u5_mult_79_n538) );
  NAND3_X4 u5_mult_79_U1402 ( .A1(u5_mult_79_n535), .A2(u5_mult_79_n536), .A3(
        u5_mult_79_n537), .ZN(u5_mult_79_CARRYB_18__18_) );
  NAND2_X2 u5_mult_79_U1401 ( .A1(u5_mult_79_CARRYB_17__18_), .A2(
        u5_mult_79_SUMB_17__19_), .ZN(u5_mult_79_n537) );
  NAND2_X2 u5_mult_79_U1400 ( .A1(u5_mult_79_ab_18__18_), .A2(
        u5_mult_79_SUMB_17__19_), .ZN(u5_mult_79_n536) );
  NAND2_X1 u5_mult_79_U1399 ( .A1(u5_mult_79_ab_18__18_), .A2(
        u5_mult_79_CARRYB_17__18_), .ZN(u5_mult_79_n535) );
  NAND2_X2 u5_mult_79_U1398 ( .A1(u5_mult_79_CARRYB_16__19_), .A2(
        u5_mult_79_SUMB_16__20_), .ZN(u5_mult_79_n534) );
  NAND2_X2 u5_mult_79_U1397 ( .A1(u5_mult_79_ab_17__19_), .A2(
        u5_mult_79_SUMB_16__20_), .ZN(u5_mult_79_n533) );
  NAND2_X1 u5_mult_79_U1396 ( .A1(u5_mult_79_ab_17__19_), .A2(
        u5_mult_79_CARRYB_16__19_), .ZN(u5_mult_79_n532) );
  XOR2_X2 u5_mult_79_U1395 ( .A(u5_mult_79_n531), .B(u5_mult_79_SUMB_17__19_), 
        .Z(u5_mult_79_SUMB_18__18_) );
  XOR2_X2 u5_mult_79_U1394 ( .A(u5_mult_79_ab_18__18_), .B(
        u5_mult_79_CARRYB_17__18_), .Z(u5_mult_79_n531) );
  XOR2_X2 u5_mult_79_U1393 ( .A(u5_mult_79_n530), .B(u5_mult_79_n106), .Z(
        u5_mult_79_SUMB_17__19_) );
  XOR2_X2 u5_mult_79_U1392 ( .A(u5_mult_79_ab_17__19_), .B(
        u5_mult_79_CARRYB_16__19_), .Z(u5_mult_79_n530) );
  NAND3_X4 u5_mult_79_U1391 ( .A1(u5_mult_79_n527), .A2(u5_mult_79_n528), .A3(
        u5_mult_79_n529), .ZN(u5_mult_79_CARRYB_22__14_) );
  NAND2_X2 u5_mult_79_U1390 ( .A1(u5_mult_79_CARRYB_21__14_), .A2(
        u5_mult_79_SUMB_21__15_), .ZN(u5_mult_79_n529) );
  NAND2_X2 u5_mult_79_U1389 ( .A1(u5_mult_79_ab_22__14_), .A2(
        u5_mult_79_SUMB_21__15_), .ZN(u5_mult_79_n528) );
  NAND2_X1 u5_mult_79_U1388 ( .A1(u5_mult_79_ab_22__14_), .A2(
        u5_mult_79_CARRYB_21__14_), .ZN(u5_mult_79_n527) );
  NAND3_X2 u5_mult_79_U1387 ( .A1(u5_mult_79_n524), .A2(u5_mult_79_n525), .A3(
        u5_mult_79_n526), .ZN(u5_mult_79_CARRYB_21__15_) );
  NAND2_X2 u5_mult_79_U1386 ( .A1(u5_mult_79_CARRYB_20__15_), .A2(
        u5_mult_79_SUMB_20__16_), .ZN(u5_mult_79_n526) );
  NAND2_X2 u5_mult_79_U1385 ( .A1(u5_mult_79_ab_21__15_), .A2(
        u5_mult_79_SUMB_20__16_), .ZN(u5_mult_79_n525) );
  NAND2_X1 u5_mult_79_U1384 ( .A1(u5_mult_79_ab_21__15_), .A2(
        u5_mult_79_CARRYB_20__15_), .ZN(u5_mult_79_n524) );
  XOR2_X2 u5_mult_79_U1383 ( .A(u5_mult_79_n523), .B(u5_mult_79_SUMB_21__15_), 
        .Z(u5_mult_79_SUMB_22__14_) );
  XOR2_X2 u5_mult_79_U1382 ( .A(u5_mult_79_ab_22__14_), .B(
        u5_mult_79_CARRYB_21__14_), .Z(u5_mult_79_n523) );
  NAND2_X1 u5_mult_79_U1381 ( .A1(u5_mult_79_CARRYB_8__16_), .A2(
        u5_mult_79_SUMB_8__17_), .ZN(u5_mult_79_n1271) );
  NAND2_X1 u5_mult_79_U1380 ( .A1(u5_mult_79_SUMB_20__11_), .A2(
        u5_mult_79_CARRYB_20__10_), .ZN(u5_mult_79_n1044) );
  XNOR2_X1 u5_mult_79_U1379 ( .A(u5_mult_79_n375), .B(u5_mult_79_ab_16__4_), 
        .ZN(u5_mult_79_n521) );
  XNOR2_X2 u5_mult_79_U1378 ( .A(u5_mult_79_n521), .B(u5_mult_79_n351), .ZN(
        u5_mult_79_SUMB_16__4_) );
  NAND2_X2 u5_mult_79_U1377 ( .A1(u5_mult_79_ab_7__13_), .A2(
        u5_mult_79_SUMB_6__14_), .ZN(u5_mult_79_n1416) );
  XNOR2_X2 u5_mult_79_U1376 ( .A(u5_mult_79_CARRYB_20__2_), .B(
        u5_mult_79_ab_21__2_), .ZN(u5_mult_79_n779) );
  NAND2_X2 u5_mult_79_U1375 ( .A1(u5_mult_79_ab_17__8_), .A2(u5_mult_79_n518), 
        .ZN(u5_mult_79_n520) );
  NAND2_X2 u5_mult_79_U1374 ( .A1(u5_mult_79_n1458), .A2(
        u5_mult_79_CARRYB_16__8_), .ZN(u5_mult_79_n519) );
  NAND2_X1 u5_mult_79_U1373 ( .A1(u5_mult_79_CARRYB_11__14_), .A2(
        u5_mult_79_SUMB_11__15_), .ZN(u5_mult_79_n724) );
  NAND2_X1 u5_mult_79_U1372 ( .A1(u5_mult_79_ab_12__14_), .A2(
        u5_mult_79_CARRYB_11__14_), .ZN(u5_mult_79_n722) );
  NAND2_X1 u5_mult_79_U1371 ( .A1(u5_mult_79_CARRYB_20__9_), .A2(
        u5_mult_79_SUMB_20__10_), .ZN(u5_mult_79_n1432) );
  NAND2_X1 u5_mult_79_U1370 ( .A1(u5_mult_79_ab_21__9_), .A2(
        u5_mult_79_SUMB_20__10_), .ZN(u5_mult_79_n1431) );
  XNOR2_X2 u5_mult_79_U1369 ( .A(u5_mult_79_n517), .B(u5_mult_79_n119), .ZN(
        u5_mult_79_SUMB_22__3_) );
  XNOR2_X2 u5_mult_79_U1368 ( .A(u5_mult_79_ab_21__1_), .B(
        u5_mult_79_SUMB_20__2_), .ZN(u5_mult_79_n1304) );
  NAND2_X2 u5_mult_79_U1367 ( .A1(u5_mult_79_ab_12__16_), .A2(
        u5_mult_79_SUMB_11__17_), .ZN(u5_mult_79_n742) );
  XNOR2_X2 u5_mult_79_U1366 ( .A(u5_mult_79_ab_13__8_), .B(
        u5_mult_79_CARRYB_12__8_), .ZN(u5_mult_79_n751) );
  XNOR2_X2 u5_mult_79_U1365 ( .A(u5_mult_79_n516), .B(u5_mult_79_n368), .ZN(
        u5_mult_79_SUMB_20__8_) );
  NAND3_X2 u5_mult_79_U1364 ( .A1(u5_mult_79_n995), .A2(u5_mult_79_n996), .A3(
        u5_mult_79_n997), .ZN(u5_mult_79_CARRYB_14__7_) );
  NAND2_X2 u5_mult_79_U1363 ( .A1(u5_mult_79_CARRYB_13__14_), .A2(
        u5_mult_79_n472), .ZN(u5_mult_79_n1555) );
  NAND2_X2 u5_mult_79_U1362 ( .A1(u5_mult_79_ab_3__15_), .A2(u5_mult_79_n324), 
        .ZN(u5_mult_79_n1349) );
  XNOR2_X2 u5_mult_79_U1361 ( .A(u5_mult_79_n515), .B(u5_mult_79_n485), .ZN(
        u5_mult_79_SUMB_17__15_) );
  NAND2_X1 u5_mult_79_U1360 ( .A1(u5_mult_79_SUMB_5__19_), .A2(
        u5_mult_79_CARRYB_5__18_), .ZN(u5_mult_79_n612) );
  NAND2_X2 u5_mult_79_U1359 ( .A1(u5_mult_79_ab_14__13_), .A2(
        u5_mult_79_SUMB_13__14_), .ZN(u5_mult_79_n1522) );
  XNOR2_X2 u5_mult_79_U1358 ( .A(u5_mult_79_ab_22__10_), .B(
        u5_mult_79_CARRYB_21__10_), .ZN(u5_mult_79_n514) );
  XNOR2_X2 u5_mult_79_U1357 ( .A(u5_mult_79_n514), .B(u5_mult_79_n494), .ZN(
        u5_mult_79_SUMB_22__10_) );
  XNOR2_X2 u5_mult_79_U1356 ( .A(u5_mult_79_n513), .B(u5_mult_79_n347), .ZN(
        u5_mult_79_SUMB_15__7_) );
  NAND2_X2 u5_mult_79_U1355 ( .A1(u5_mult_79_ab_22__3_), .A2(
        u5_mult_79_CARRYB_21__3_), .ZN(u5_mult_79_n583) );
  NAND3_X2 u5_mult_79_U1354 ( .A1(u5_mult_79_n1569), .A2(u5_mult_79_n1570), 
        .A3(u5_mult_79_n1571), .ZN(u5_mult_79_CARRYB_18__9_) );
  NAND2_X2 u5_mult_79_U1353 ( .A1(u5_mult_79_ab_22__7_), .A2(
        u5_mult_79_SUMB_21__8_), .ZN(u5_mult_79_n963) );
  NAND2_X2 u5_mult_79_U1352 ( .A1(u5_mult_79_CARRYB_21__7_), .A2(
        u5_mult_79_SUMB_21__8_), .ZN(u5_mult_79_n964) );
  NAND2_X1 u5_mult_79_U1351 ( .A1(u5_mult_79_ab_6__15_), .A2(
        u5_mult_79_CARRYB_5__15_), .ZN(u5_mult_79_n1537) );
  NOR2_X2 u5_mult_79_U1350 ( .A1(u5_mult_79_n1831), .A2(u5_mult_79_n1725), 
        .ZN(u5_mult_79_ab_3__23_) );
  NOR2_X2 u5_mult_79_U1349 ( .A1(u5_mult_79_n1831), .A2(u5_mult_79_n1740), 
        .ZN(u5_mult_79_ab_8__23_) );
  NOR2_X2 u5_mult_79_U1348 ( .A1(u5_mult_79_n1831), .A2(u5_mult_79_n1746), 
        .ZN(u5_mult_79_ab_10__23_) );
  INV_X4 u5_mult_79_U1347 ( .A(u5_mult_79_CARRYB_22__2_), .ZN(u5_mult_79_n1050) );
  XNOR2_X2 u5_mult_79_U1346 ( .A(u5_mult_79_n595), .B(u5_mult_79_n12), .ZN(
        u5_mult_79_SUMB_8__12_) );
  XNOR2_X2 u5_mult_79_U1345 ( .A(u5_mult_79_n576), .B(u5_mult_79_n320), .ZN(
        u5_mult_79_SUMB_12__16_) );
  NAND2_X2 u5_mult_79_U1344 ( .A1(u5_mult_79_ab_19__2_), .A2(
        u5_mult_79_SUMB_18__3_), .ZN(u5_mult_79_n1027) );
  NAND3_X2 u5_mult_79_U1343 ( .A1(u5_mult_79_n1185), .A2(u5_mult_79_n1186), 
        .A3(u5_mult_79_n1187), .ZN(u5_mult_79_CARRYB_21__5_) );
  XNOR2_X2 u5_mult_79_U1342 ( .A(u5_mult_79_ab_17__15_), .B(
        u5_mult_79_CARRYB_16__15_), .ZN(u5_mult_79_n515) );
  NAND2_X4 u5_mult_79_U1341 ( .A1(u5_mult_79_n617), .A2(u5_mult_79_n1269), 
        .ZN(u5_mult_79_CARRYB_9__16_) );
  XNOR2_X2 u5_mult_79_U1340 ( .A(u5_mult_79_CARRYB_19__2_), .B(
        u5_mult_79_ab_20__2_), .ZN(u5_mult_79_n512) );
  XNOR2_X2 u5_mult_79_U1339 ( .A(u5_mult_79_n512), .B(u5_mult_79_n109), .ZN(
        u5_mult_79_SUMB_20__2_) );
  NAND3_X4 u5_mult_79_U1338 ( .A1(u5_mult_79_n1175), .A2(u5_mult_79_n1176), 
        .A3(u5_mult_79_n1177), .ZN(u5_mult_79_CARRYB_22__1_) );
  NOR2_X1 u5_mult_79_U1337 ( .A1(u5_mult_79_n1829), .A2(u5_mult_79_n1828), 
        .ZN(u5_mult_79_ab_23__1_) );
  CLKBUF_X3 u5_mult_79_U1336 ( .A(u5_mult_79_SUMB_20__3_), .Z(u5_mult_79_n511)
         );
  NAND3_X2 u5_mult_79_U1335 ( .A1(u5_mult_79_n508), .A2(u5_mult_79_n509), .A3(
        u5_mult_79_n510), .ZN(u5_mult_79_CARRYB_23__1_) );
  NAND2_X2 u5_mult_79_U1334 ( .A1(u5_mult_79_ab_23__1_), .A2(
        u5_mult_79_SUMB_22__2_), .ZN(u5_mult_79_n509) );
  NAND2_X2 u5_mult_79_U1333 ( .A1(u5_mult_79_ab_10__9_), .A2(
        u5_mult_79_SUMB_9__10_), .ZN(u5_mult_79_n504) );
  NAND2_X1 u5_mult_79_U1332 ( .A1(u5_mult_79_CARRYB_9__9_), .A2(
        u5_mult_79_ab_10__9_), .ZN(u5_mult_79_n502) );
  XNOR2_X2 u5_mult_79_U1331 ( .A(u5_mult_79_ab_18__8_), .B(
        u5_mult_79_CARRYB_17__8_), .ZN(u5_mult_79_n501) );
  XNOR2_X2 u5_mult_79_U1330 ( .A(u5_mult_79_SUMB_17__9_), .B(u5_mult_79_n501), 
        .ZN(u5_mult_79_SUMB_18__8_) );
  XNOR2_X2 u5_mult_79_U1329 ( .A(u5_mult_79_CARRYB_3__18_), .B(
        u5_mult_79_ab_4__18_), .ZN(u5_mult_79_n500) );
  XNOR2_X2 u5_mult_79_U1328 ( .A(u5_mult_79_SUMB_3__19_), .B(u5_mult_79_n500), 
        .ZN(u5_mult_79_SUMB_4__18_) );
  NAND2_X2 u5_mult_79_U1327 ( .A1(u5_mult_79_ab_11__12_), .A2(
        u5_mult_79_SUMB_10__13_), .ZN(u5_mult_79_n1403) );
  XOR2_X2 u5_mult_79_U1326 ( .A(u5_mult_79_n587), .B(u5_mult_79_SUMB_2__18_), 
        .Z(u5_mult_79_SUMB_3__17_) );
  NAND2_X4 u5_mult_79_U1325 ( .A1(u5_mult_79_CARRYB_17__10_), .A2(
        u5_mult_79_SUMB_17__11_), .ZN(u5_mult_79_n825) );
  NAND2_X2 u5_mult_79_U1324 ( .A1(u5_mult_79_n849), .A2(u5_mult_79_ab_18__14_), 
        .ZN(u5_mult_79_n851) );
  INV_X4 u5_mult_79_U1323 ( .A(u5_mult_79_n497), .ZN(u5_mult_79_n498) );
  INV_X4 u5_mult_79_U1322 ( .A(u5_mult_79_n495), .ZN(u5_mult_79_n496) );
  INV_X2 u5_mult_79_U1321 ( .A(u5_mult_79_SUMB_5__15_), .ZN(u5_mult_79_n495)
         );
  INV_X1 u5_mult_79_U1320 ( .A(u5_mult_79_n367), .ZN(u5_mult_79_n493) );
  CLKBUF_X2 u5_mult_79_U1319 ( .A(u5_mult_79_CARRYB_19__1_), .Z(
        u5_mult_79_n492) );
  CLKBUF_X3 u5_mult_79_U1318 ( .A(u5_mult_79_SUMB_17__6_), .Z(u5_mult_79_n491)
         );
  INV_X2 u5_mult_79_U1317 ( .A(u5_mult_79_SUMB_11__14_), .ZN(u5_mult_79_n489)
         );
  INV_X8 u5_mult_79_U1316 ( .A(u5_mult_79_n487), .ZN(u5_mult_79_n488) );
  INV_X2 u5_mult_79_U1315 ( .A(u5_mult_79_SUMB_2__17_), .ZN(u5_mult_79_n487)
         );
  XNOR2_X2 u5_mult_79_U1314 ( .A(u5_mult_79_ab_6__18_), .B(
        u5_mult_79_CARRYB_5__18_), .ZN(u5_mult_79_n486) );
  INV_X4 u5_mult_79_U1313 ( .A(u5_mult_79_n483), .ZN(u5_mult_79_n484) );
  INV_X2 u5_mult_79_U1312 ( .A(u5_mult_79_SUMB_13__17_), .ZN(u5_mult_79_n483)
         );
  XNOR2_X2 u5_mult_79_U1311 ( .A(u5_mult_79_n481), .B(u5_mult_79_SUMB_14__17_), 
        .ZN(u5_mult_79_SUMB_15__16_) );
  XNOR2_X2 u5_mult_79_U1310 ( .A(u5_mult_79_CARRYB_1__21_), .B(
        u5_mult_79_ab_2__21_), .ZN(u5_mult_79_n480) );
  XNOR2_X2 u5_mult_79_U1309 ( .A(u5_mult_79_SUMB_1__22_), .B(u5_mult_79_n480), 
        .ZN(u5_mult_79_SUMB_2__21_) );
  XNOR2_X2 u5_mult_79_U1308 ( .A(u5_mult_79_n479), .B(u5_mult_79_SUMB_15__11_), 
        .ZN(u5_mult_79_SUMB_16__10_) );
  XNOR2_X2 u5_mult_79_U1307 ( .A(u5_mult_79_n688), .B(u5_mult_79_SUMB_7__8_), 
        .ZN(u5_mult_79_SUMB_8__7_) );
  NAND2_X1 u5_mult_79_U1306 ( .A1(u5_mult_79_n304), .A2(u5_mult_79_SUMB_20__7_), .ZN(u5_mult_79_n1561) );
  CLKBUF_X2 u5_mult_79_U1305 ( .A(u5_mult_79_SUMB_12__19_), .Z(u5_mult_79_n477) );
  XNOR2_X2 u5_mult_79_U1304 ( .A(u5_mult_79_CARRYB_20__3_), .B(
        u5_mult_79_ab_21__3_), .ZN(u5_mult_79_n475) );
  XNOR2_X1 u5_mult_79_U1303 ( .A(u5_mult_79_CARRYB_11__7_), .B(
        u5_mult_79_ab_12__7_), .ZN(u5_mult_79_n473) );
  XNOR2_X2 u5_mult_79_U1302 ( .A(u5_mult_79_n473), .B(u5_mult_79_n316), .ZN(
        u5_mult_79_SUMB_12__7_) );
  INV_X4 u5_mult_79_U1301 ( .A(u5_mult_79_n471), .ZN(u5_mult_79_n472) );
  INV_X2 u5_mult_79_U1300 ( .A(u5_mult_79_SUMB_13__15_), .ZN(u5_mult_79_n471)
         );
  XNOR2_X2 u5_mult_79_U1299 ( .A(u5_mult_79_ab_12__15_), .B(
        u5_mult_79_CARRYB_11__15_), .ZN(u5_mult_79_n470) );
  XNOR2_X2 u5_mult_79_U1298 ( .A(u5_mult_79_n470), .B(u5_mult_79_n302), .ZN(
        u5_mult_79_SUMB_12__15_) );
  XNOR2_X2 u5_mult_79_U1297 ( .A(u5_mult_79_n958), .B(u5_mult_79_n493), .ZN(
        u5_mult_79_SUMB_21__8_) );
  XNOR2_X1 u5_mult_79_U1296 ( .A(u5_mult_79_ab_6__9_), .B(
        u5_mult_79_CARRYB_5__9_), .ZN(u5_mult_79_n468) );
  XNOR2_X2 u5_mult_79_U1295 ( .A(u5_mult_79_n468), .B(u5_mult_79_SUMB_5__10_), 
        .ZN(u5_mult_79_SUMB_6__9_) );
  XNOR2_X2 u5_mult_79_U1294 ( .A(u5_mult_79_n467), .B(u5_mult_79_SUMB_10__11_), 
        .ZN(u5_mult_79_SUMB_11__10_) );
  INV_X4 u5_mult_79_U1293 ( .A(u5_mult_79_n465), .ZN(u5_mult_79_n466) );
  INV_X2 u5_mult_79_U1292 ( .A(u5_mult_79_SUMB_20__6_), .ZN(u5_mult_79_n465)
         );
  XNOR2_X2 u5_mult_79_U1291 ( .A(u5_mult_79_ab_6__14_), .B(
        u5_mult_79_CARRYB_5__14_), .ZN(u5_mult_79_n464) );
  XNOR2_X2 u5_mult_79_U1290 ( .A(u5_mult_79_n464), .B(u5_mult_79_n496), .ZN(
        u5_mult_79_SUMB_6__14_) );
  XNOR2_X2 u5_mult_79_U1289 ( .A(u5_mult_79_n461), .B(u5_mult_79_n426), .ZN(
        u5_mult_79_SUMB_15__14_) );
  XNOR2_X2 u5_mult_79_U1288 ( .A(u5_mult_79_n385), .B(u5_mult_79_n460), .ZN(
        u5_mult_79_SUMB_12__5_) );
  XNOR2_X2 u5_mult_79_U1287 ( .A(u5_mult_79_CARRYB_6__9_), .B(
        u5_mult_79_ab_7__9_), .ZN(u5_mult_79_n459) );
  XNOR2_X2 u5_mult_79_U1286 ( .A(u5_mult_79_SUMB_6__10_), .B(u5_mult_79_n459), 
        .ZN(u5_mult_79_SUMB_7__9_) );
  XNOR2_X2 u5_mult_79_U1285 ( .A(u5_mult_79_n878), .B(u5_mult_79_n318), .ZN(
        u5_mult_79_SUMB_9__16_) );
  XNOR2_X2 u5_mult_79_U1284 ( .A(u5_mult_79_CARRYB_15__9_), .B(
        u5_mult_79_ab_16__9_), .ZN(u5_mult_79_n458) );
  XNOR2_X2 u5_mult_79_U1283 ( .A(u5_mult_79_n448), .B(u5_mult_79_n458), .ZN(
        u5_mult_79_SUMB_16__9_) );
  XNOR2_X2 u5_mult_79_U1282 ( .A(u5_mult_79_ab_15__5_), .B(
        u5_mult_79_CARRYB_14__5_), .ZN(u5_mult_79_n456) );
  NAND3_X2 u5_mult_79_U1281 ( .A1(u5_mult_79_n952), .A2(u5_mult_79_n951), .A3(
        u5_mult_79_n950), .ZN(u5_mult_79_CARRYB_17__14_) );
  XNOR2_X2 u5_mult_79_U1280 ( .A(u5_mult_79_ab_15__8_), .B(
        u5_mult_79_CARRYB_14__8_), .ZN(u5_mult_79_n455) );
  XNOR2_X2 u5_mult_79_U1279 ( .A(u5_mult_79_n455), .B(u5_mult_79_n125), .ZN(
        u5_mult_79_SUMB_15__8_) );
  XNOR2_X2 u5_mult_79_U1278 ( .A(u5_mult_79_CARRYB_20__4_), .B(
        u5_mult_79_ab_21__4_), .ZN(u5_mult_79_n453) );
  XNOR2_X2 u5_mult_79_U1277 ( .A(u5_mult_79_n453), .B(u5_mult_79_n420), .ZN(
        u5_mult_79_SUMB_21__4_) );
  XNOR2_X2 u5_mult_79_U1276 ( .A(u5_mult_79_SUMB_20__11_), .B(u5_mult_79_n452), 
        .ZN(u5_mult_79_SUMB_21__10_) );
  XNOR2_X2 u5_mult_79_U1275 ( .A(u5_mult_79_n45), .B(u5_mult_79_n451), .ZN(
        u5_mult_79_SUMB_11__13_) );
  XNOR2_X2 u5_mult_79_U1274 ( .A(u5_mult_79_n542), .B(u5_mult_79_n427), .ZN(
        u5_mult_79_SUMB_7__13_) );
  NAND3_X2 u5_mult_79_U1273 ( .A1(u5_mult_79_n1106), .A2(u5_mult_79_n1107), 
        .A3(u5_mult_79_n1108), .ZN(u5_mult_79_CARRYB_11__7_) );
  INV_X2 u5_mult_79_U1272 ( .A(u5_mult_79_n449), .ZN(u5_mult_79_n450) );
  XNOR2_X2 u5_mult_79_U1271 ( .A(u5_mult_79_SUMB_13__14_), .B(u5_mult_79_n1425), .ZN(u5_mult_79_SUMB_14__13_) );
  NAND2_X1 u5_mult_79_U1270 ( .A1(u5_mult_79_CARRYB_14__12_), .A2(
        u5_mult_79_SUMB_14__13_), .ZN(u5_mult_79_n1364) );
  INV_X8 u5_mult_79_U1269 ( .A(u5_mult_79_n447), .ZN(u5_mult_79_n448) );
  XNOR2_X2 u5_mult_79_U1268 ( .A(u5_mult_79_CARRYB_16__14_), .B(
        u5_mult_79_ab_17__14_), .ZN(u5_mult_79_n446) );
  XNOR2_X2 u5_mult_79_U1267 ( .A(u5_mult_79_n446), .B(u5_mult_79_SUMB_16__15_), 
        .ZN(u5_mult_79_SUMB_17__14_) );
  XNOR2_X2 u5_mult_79_U1266 ( .A(u5_mult_79_ab_18__11_), .B(
        u5_mult_79_CARRYB_17__11_), .ZN(u5_mult_79_n445) );
  XNOR2_X2 u5_mult_79_U1265 ( .A(u5_mult_79_SUMB_17__12_), .B(u5_mult_79_n445), 
        .ZN(u5_mult_79_SUMB_18__11_) );
  XNOR2_X2 u5_mult_79_U1264 ( .A(u5_mult_79_CARRYB_17__10_), .B(
        u5_mult_79_ab_18__10_), .ZN(u5_mult_79_n444) );
  XNOR2_X2 u5_mult_79_U1263 ( .A(u5_mult_79_SUMB_17__11_), .B(u5_mult_79_n444), 
        .ZN(u5_mult_79_SUMB_18__10_) );
  XNOR2_X1 u5_mult_79_U1262 ( .A(u5_mult_79_CARRYB_18__9_), .B(
        u5_mult_79_ab_19__9_), .ZN(u5_mult_79_n443) );
  XNOR2_X2 u5_mult_79_U1261 ( .A(u5_mult_79_SUMB_18__10_), .B(u5_mult_79_n443), 
        .ZN(u5_mult_79_SUMB_19__9_) );
  XOR2_X1 u5_mult_79_U1260 ( .A(u5_mult_79_n1135), .B(u5_mult_79_n421), .Z(
        u5_mult_79_SUMB_18__14_) );
  XOR2_X2 u5_mult_79_U1259 ( .A(u5_mult_79_n1135), .B(u5_mult_79_n421), .Z(
        u5_mult_79_n440) );
  XNOR2_X2 u5_mult_79_U1258 ( .A(u5_mult_79_CARRYB_19__7_), .B(
        u5_mult_79_ab_20__7_), .ZN(u5_mult_79_n438) );
  NAND3_X2 u5_mult_79_U1257 ( .A1(u5_mult_79_n900), .A2(u5_mult_79_n901), .A3(
        u5_mult_79_n902), .ZN(u5_mult_79_CARRYB_6__20_) );
  XNOR2_X1 u5_mult_79_U1256 ( .A(u5_mult_79_SUMB_19__8_), .B(u5_mult_79_n438), 
        .ZN(u5_mult_79_SUMB_20__7_) );
  NAND2_X1 u5_mult_79_U1255 ( .A1(u5_mult_79_SUMB_19__8_), .A2(
        u5_mult_79_ab_20__7_), .ZN(u5_mult_79_n1089) );
  NAND3_X2 u5_mult_79_U1254 ( .A1(u5_mult_79_n859), .A2(u5_mult_79_n860), .A3(
        u5_mult_79_n861), .ZN(u5_mult_79_CARRYB_16__3_) );
  INV_X4 u5_mult_79_U1253 ( .A(u5_mult_79_CARRYB_15__13_), .ZN(u5_mult_79_n429) );
  XNOR2_X2 u5_mult_79_U1252 ( .A(u5_mult_79_CARRYB_11__10_), .B(
        u5_mult_79_ab_12__10_), .ZN(u5_mult_79_n428) );
  XNOR2_X2 u5_mult_79_U1251 ( .A(u5_mult_79_SUMB_11__11_), .B(u5_mult_79_n428), 
        .ZN(u5_mult_79_SUMB_12__10_) );
  NAND2_X2 u5_mult_79_U1250 ( .A1(u5_mult_79_ab_6__15_), .A2(
        u5_mult_79_SUMB_5__16_), .ZN(u5_mult_79_n1538) );
  CLKBUF_X2 u5_mult_79_U1249 ( .A(u5_mult_79_SUMB_6__14_), .Z(u5_mult_79_n427)
         );
  XNOR2_X2 u5_mult_79_U1248 ( .A(u5_mult_79_CARRYB_11__5_), .B(
        u5_mult_79_ab_12__5_), .ZN(u5_mult_79_n460) );
  CLKBUF_X3 u5_mult_79_U1247 ( .A(u5_mult_79_n294), .Z(u5_mult_79_n426) );
  NAND2_X2 u5_mult_79_U1246 ( .A1(u5_mult_79_ab_12__5_), .A2(
        u5_mult_79_CARRYB_11__5_), .ZN(u5_mult_79_n1117) );
  XNOR2_X2 u5_mult_79_U1245 ( .A(u5_mult_79_ab_6__17_), .B(
        u5_mult_79_CARRYB_5__17_), .ZN(u5_mult_79_n425) );
  XNOR2_X2 u5_mult_79_U1244 ( .A(u5_mult_79_n425), .B(u5_mult_79_n305), .ZN(
        u5_mult_79_SUMB_6__17_) );
  XNOR2_X2 u5_mult_79_U1243 ( .A(u5_mult_79_ab_9__13_), .B(
        u5_mult_79_CARRYB_8__13_), .ZN(u5_mult_79_n424) );
  XNOR2_X2 u5_mult_79_U1242 ( .A(u5_mult_79_n424), .B(u5_mult_79_n24), .ZN(
        u5_mult_79_SUMB_9__13_) );
  XNOR2_X2 u5_mult_79_U1241 ( .A(u5_mult_79_ab_22__3_), .B(
        u5_mult_79_CARRYB_21__3_), .ZN(u5_mult_79_n517) );
  INV_X2 u5_mult_79_U1240 ( .A(u5_mult_79_n454), .ZN(u5_mult_79_n1213) );
  FA_X1 u5_mult_79_U1239 ( .A(u5_mult_79_ab_2__19_), .B(
        u5_mult_79_CARRYB_1__19_), .CI(u5_mult_79_SUMB_1__20_), .S(
        u5_mult_79_n423) );
  FA_X1 u5_mult_79_U1238 ( .A(u5_mult_79_SUMB_1__20_), .B(
        u5_mult_79_CARRYB_1__19_), .CI(u5_mult_79_ab_2__19_), .S(
        u5_mult_79_n422) );
  BUF_X8 u5_mult_79_U1237 ( .A(u5_mult_79_SUMB_17__15_), .Z(u5_mult_79_n421)
         );
  INV_X4 u5_mult_79_U1236 ( .A(u5_mult_79_n419), .ZN(u5_mult_79_n420) );
  INV_X2 u5_mult_79_U1235 ( .A(u5_mult_79_SUMB_20__5_), .ZN(u5_mult_79_n419)
         );
  XNOR2_X2 u5_mult_79_U1234 ( .A(u5_mult_79_ab_14__8_), .B(
        u5_mult_79_CARRYB_13__8_), .ZN(u5_mult_79_n418) );
  XNOR2_X2 u5_mult_79_U1233 ( .A(u5_mult_79_n418), .B(u5_mult_79_SUMB_13__9_), 
        .ZN(u5_mult_79_SUMB_14__8_) );
  XNOR2_X2 u5_mult_79_U1232 ( .A(u5_mult_79_n431), .B(u5_mult_79_n113), .ZN(
        u5_mult_79_SUMB_13__5_) );
  CLKBUF_X3 u5_mult_79_U1231 ( .A(u5_mult_79_SUMB_13__5_), .Z(u5_mult_79_n417)
         );
  XNOR2_X2 u5_mult_79_U1230 ( .A(u5_mult_79_ab_23__12_), .B(
        u5_mult_79_CARRYB_22__12_), .ZN(u5_mult_79_n416) );
  XNOR2_X2 u5_mult_79_U1229 ( .A(u5_mult_79_SUMB_22__13_), .B(u5_mult_79_n416), 
        .ZN(u5_mult_79_SUMB_23__12_) );
  INV_X2 u5_mult_79_U1228 ( .A(u5_mult_79_n412), .ZN(u5_mult_79_n413) );
  INV_X1 u5_mult_79_U1227 ( .A(u5_mult_79_SUMB_21__6_), .ZN(u5_mult_79_n412)
         );
  NAND2_X1 u5_mult_79_U1226 ( .A1(u5_mult_79_n1504), .A2(u5_mult_79_n474), 
        .ZN(u5_mult_79_n1258) );
  BUF_X8 u5_mult_79_U1225 ( .A(u5_mult_79_SUMB_21__2_), .Z(u5_mult_79_n411) );
  NAND2_X1 u5_mult_79_U1224 ( .A1(u5_mult_79_ab_21__5_), .A2(
        u5_mult_79_CARRYB_20__5_), .ZN(u5_mult_79_n1185) );
  XNOR2_X2 u5_mult_79_U1223 ( .A(u5_mult_79_n8), .B(u5_mult_79_n410), .ZN(
        u5_mult_79_SUMB_10__13_) );
  XNOR2_X2 u5_mult_79_U1222 ( .A(u5_mult_79_ab_22__12_), .B(
        u5_mult_79_CARRYB_21__12_), .ZN(u5_mult_79_n409) );
  XNOR2_X2 u5_mult_79_U1221 ( .A(u5_mult_79_n409), .B(u5_mult_79_n499), .ZN(
        u5_mult_79_SUMB_22__12_) );
  XNOR2_X2 u5_mult_79_U1220 ( .A(u5_mult_79_ab_21__9_), .B(
        u5_mult_79_CARRYB_20__9_), .ZN(u5_mult_79_n408) );
  XNOR2_X2 u5_mult_79_U1219 ( .A(u5_mult_79_n408), .B(u5_mult_79_SUMB_20__10_), 
        .ZN(u5_mult_79_SUMB_21__9_) );
  CLKBUF_X2 u5_mult_79_U1218 ( .A(u5_mult_79_SUMB_5__16_), .Z(u5_mult_79_n407)
         );
  NAND2_X2 u5_mult_79_U1217 ( .A1(u5_mult_79_n401), .A2(
        u5_mult_79_CARRYB_2__21_), .ZN(u5_mult_79_n1600) );
  INV_X4 u5_mult_79_U1216 ( .A(u5_mult_79_n405), .ZN(u5_mult_79_n406) );
  INV_X4 u5_mult_79_U1215 ( .A(u5_mult_79_n403), .ZN(u5_mult_79_n404) );
  INV_X2 u5_mult_79_U1214 ( .A(u5_mult_79_SUMB_10__6_), .ZN(u5_mult_79_n403)
         );
  NAND2_X1 u5_mult_79_U1213 ( .A1(u5_mult_79_SUMB_6__8_), .A2(
        u5_mult_79_ab_7__7_), .ZN(u5_mult_79_n1017) );
  XNOR2_X2 u5_mult_79_U1212 ( .A(u5_mult_79_SUMB_7__7_), .B(u5_mult_79_n402), 
        .ZN(u5_mult_79_SUMB_8__6_) );
  NAND2_X1 u5_mult_79_U1211 ( .A1(u5_mult_79_ab_15__15_), .A2(
        u5_mult_79_CARRYB_14__15_), .ZN(u5_mult_79_n1439) );
  BUF_X4 u5_mult_79_U1210 ( .A(u5_mult_79_SUMB_13__16_), .Z(u5_mult_79_n476)
         );
  NAND2_X2 u5_mult_79_U1209 ( .A1(u5_mult_79_CARRYB_17__7_), .A2(
        u5_mult_79_SUMB_17__8_), .ZN(u5_mult_79_n1615) );
  NAND2_X2 u5_mult_79_U1208 ( .A1(u5_mult_79_ab_18__7_), .A2(
        u5_mult_79_SUMB_17__8_), .ZN(u5_mult_79_n1614) );
  INV_X4 u5_mult_79_U1207 ( .A(u5_mult_79_n400), .ZN(u5_mult_79_n401) );
  INV_X2 u5_mult_79_U1206 ( .A(u5_mult_79_SUMB_2__22_), .ZN(u5_mult_79_n400)
         );
  XNOR2_X2 u5_mult_79_U1205 ( .A(u5_mult_79_n415), .B(u5_mult_79_n399), .ZN(
        u5_mult_79_SUMB_18__3_) );
  XNOR2_X2 u5_mult_79_U1204 ( .A(u5_mult_79_n398), .B(u5_mult_79_n482), .ZN(
        u5_mult_79_SUMB_7__17_) );
  XNOR2_X2 u5_mult_79_U1203 ( .A(u5_mult_79_n406), .B(u5_mult_79_ab_11__8_), 
        .ZN(u5_mult_79_n397) );
  NAND2_X1 u5_mult_79_U1202 ( .A1(u5_mult_79_ab_9__8_), .A2(
        u5_mult_79_SUMB_8__9_), .ZN(u5_mult_79_n844) );
  NAND3_X2 u5_mult_79_U1201 ( .A1(u5_mult_79_n759), .A2(u5_mult_79_n760), .A3(
        u5_mult_79_n761), .ZN(u5_mult_79_CARRYB_19__13_) );
  XNOR2_X2 u5_mult_79_U1200 ( .A(u5_mult_79_ab_17__9_), .B(
        u5_mult_79_CARRYB_16__9_), .ZN(u5_mult_79_n904) );
  XNOR2_X2 u5_mult_79_U1199 ( .A(u5_mult_79_n441), .B(u5_mult_79_n394), .ZN(
        u5_mult_79_SUMB_18__12_) );
  INV_X2 u5_mult_79_U1198 ( .A(u5_mult_79_n392), .ZN(u5_mult_79_n393) );
  XNOR2_X2 u5_mult_79_U1197 ( .A(u5_mult_79_SUMB_10__5_), .B(u5_mult_79_n686), 
        .ZN(u5_mult_79_SUMB_11__4_) );
  XNOR2_X2 u5_mult_79_U1196 ( .A(u5_mult_79_ab_8__8_), .B(
        u5_mult_79_CARRYB_7__8_), .ZN(u5_mult_79_n391) );
  XNOR2_X2 u5_mult_79_U1195 ( .A(u5_mult_79_n391), .B(u5_mult_79_SUMB_7__9_), 
        .ZN(u5_mult_79_SUMB_8__8_) );
  XNOR2_X2 u5_mult_79_U1194 ( .A(u5_mult_79_CARRYB_12__14_), .B(
        u5_mult_79_ab_13__14_), .ZN(u5_mult_79_n390) );
  XNOR2_X2 u5_mult_79_U1193 ( .A(u5_mult_79_SUMB_12__15_), .B(u5_mult_79_n390), 
        .ZN(u5_mult_79_SUMB_13__14_) );
  XNOR2_X2 u5_mult_79_U1192 ( .A(u5_mult_79_CARRYB_9__5_), .B(
        u5_mult_79_ab_10__5_), .ZN(u5_mult_79_n388) );
  XNOR2_X2 u5_mult_79_U1191 ( .A(u5_mult_79_n115), .B(u5_mult_79_n388), .ZN(
        u5_mult_79_SUMB_10__5_) );
  XNOR2_X2 u5_mult_79_U1190 ( .A(u5_mult_79_ab_19__12_), .B(
        u5_mult_79_CARRYB_18__12_), .ZN(u5_mult_79_n577) );
  NAND2_X1 u5_mult_79_U1189 ( .A1(u5_mult_79_CARRYB_9__9_), .A2(
        u5_mult_79_SUMB_9__10_), .ZN(u5_mult_79_n503) );
  XNOR2_X2 u5_mult_79_U1188 ( .A(u5_mult_79_n456), .B(u5_mult_79_n133), .ZN(
        u5_mult_79_SUMB_15__5_) );
  INV_X4 u5_mult_79_U1187 ( .A(u5_mult_79_n386), .ZN(u5_mult_79_n387) );
  INV_X2 u5_mult_79_U1186 ( .A(u5_mult_79_SUMB_4__7_), .ZN(u5_mult_79_n386) );
  INV_X4 u5_mult_79_U1185 ( .A(u5_mult_79_n384), .ZN(u5_mult_79_n385) );
  INV_X2 u5_mult_79_U1184 ( .A(u5_mult_79_SUMB_11__6_), .ZN(u5_mult_79_n384)
         );
  NAND2_X1 u5_mult_79_U1183 ( .A1(u5_mult_79_SUMB_6__9_), .A2(u5_mult_79_n10), 
        .ZN(u5_mult_79_n1167) );
  CLKBUF_X2 u5_mult_79_U1182 ( .A(u5_mult_79_SUMB_16__2_), .Z(u5_mult_79_n383)
         );
  XNOR2_X2 u5_mult_79_U1181 ( .A(u5_mult_79_n382), .B(u5_mult_79_SUMB_10__18_), 
        .ZN(u5_mult_79_SUMB_11__17_) );
  INV_X4 u5_mult_79_U1180 ( .A(u5_mult_79_n380), .ZN(u5_mult_79_n381) );
  XNOR2_X2 u5_mult_79_U1179 ( .A(u5_mult_79_n379), .B(u5_mult_79_n395), .ZN(
        u5_mult_79_SUMB_6__20_) );
  XNOR2_X2 u5_mult_79_U1178 ( .A(u5_mult_79_CARRYB_7__14_), .B(
        u5_mult_79_ab_8__14_), .ZN(u5_mult_79_n378) );
  XNOR2_X2 u5_mult_79_U1177 ( .A(u5_mult_79_SUMB_7__15_), .B(u5_mult_79_n378), 
        .ZN(u5_mult_79_SUMB_8__14_) );
  NAND2_X4 u5_mult_79_U1176 ( .A1(u5_mult_79_n519), .A2(u5_mult_79_n520), .ZN(
        u5_mult_79_n1609) );
  XOR2_X2 u5_mult_79_U1175 ( .A(u5_mult_79_n127), .B(u5_mult_79_n1609), .Z(
        u5_mult_79_n377) );
  XOR2_X2 u5_mult_79_U1174 ( .A(u5_mult_79_n812), .B(u5_mult_79_n374), .Z(
        u5_mult_79_n376) );
  FA_X1 u5_mult_79_U1173 ( .A(u5_mult_79_CARRYB_14__4_), .B(
        u5_mult_79_ab_15__4_), .CI(u5_mult_79_SUMB_14__5_), .CO(
        u5_mult_79_n375), .S(u5_mult_79_n312) );
  CLKBUF_X2 u5_mult_79_U1172 ( .A(u5_mult_79_CARRYB_12__4_), .Z(
        u5_mult_79_n372) );
  XNOR2_X2 u5_mult_79_U1171 ( .A(u5_mult_79_CARRYB_10__16_), .B(
        u5_mult_79_ab_11__16_), .ZN(u5_mult_79_n371) );
  XNOR2_X1 u5_mult_79_U1170 ( .A(u5_mult_79_n371), .B(u5_mult_79_SUMB_10__17_), 
        .ZN(u5_mult_79_SUMB_11__16_) );
  XNOR2_X1 u5_mult_79_U1169 ( .A(u5_mult_79_CARRYB_13__19_), .B(
        u5_mult_79_ab_14__19_), .ZN(u5_mult_79_n370) );
  XNOR2_X2 u5_mult_79_U1168 ( .A(u5_mult_79_SUMB_13__20_), .B(u5_mult_79_n370), 
        .ZN(u5_mult_79_SUMB_14__19_) );
  XNOR2_X2 u5_mult_79_U1167 ( .A(u5_mult_79_n369), .B(
        u5_mult_79_CARRYB_16__17_), .ZN(u5_mult_79_n689) );
  INV_X4 u5_mult_79_U1166 ( .A(u5_mult_79_SUMB_20__7_), .ZN(u5_mult_79_n380)
         );
  NAND2_X2 u5_mult_79_U1165 ( .A1(u5_mult_79_n366), .A2(u5_mult_79_ab_14__20_), 
        .ZN(u5_mult_79_n1071) );
  XNOR2_X2 u5_mult_79_U1164 ( .A(u5_mult_79_n366), .B(u5_mult_79_n434), .ZN(
        u5_mult_79_n1069) );
  CLKBUF_X3 u5_mult_79_U1163 ( .A(u5_mult_79_SUMB_19__9_), .Z(u5_mult_79_n368)
         );
  INV_X4 u5_mult_79_U1162 ( .A(u5_mult_79_SUMB_14__10_), .ZN(u5_mult_79_n462)
         );
  INV_X8 u5_mult_79_U1161 ( .A(u5_mult_79_n462), .ZN(u5_mult_79_n463) );
  XNOR2_X2 u5_mult_79_U1160 ( .A(u5_mult_79_n1317), .B(u5_mult_79_n462), .ZN(
        u5_mult_79_SUMB_15__9_) );
  XNOR2_X2 u5_mult_79_U1159 ( .A(u5_mult_79_ab_5__18_), .B(
        u5_mult_79_CARRYB_4__18_), .ZN(u5_mult_79_n578) );
  NAND2_X1 u5_mult_79_U1158 ( .A1(u5_mult_79_n337), .A2(u5_mult_79_SUMB_2__21_), .ZN(u5_mult_79_n1628) );
  INV_X4 u5_mult_79_U1157 ( .A(u5_mult_79_n365), .ZN(u5_mult_79_n366) );
  INV_X2 u5_mult_79_U1156 ( .A(u5_mult_79_CARRYB_13__20_), .ZN(u5_mult_79_n365) );
  NAND2_X1 u5_mult_79_U1155 ( .A1(u5_mult_79_SUMB_23__14_), .A2(
        u5_mult_79_CARRYB_23__13_), .ZN(u5_mult_79_n1663) );
  XNOR2_X2 u5_mult_79_U1154 ( .A(u5_mult_79_n357), .B(u5_mult_79_n809), .ZN(
        u5_mult_79_SUMB_4__14_) );
  NAND2_X2 u5_mult_79_U1153 ( .A1(u5_mult_79_n406), .A2(u5_mult_79_SUMB_10__9_), .ZN(u5_mult_79_n507) );
  NAND2_X2 u5_mult_79_U1152 ( .A1(u5_mult_79_ab_11__8_), .A2(u5_mult_79_n295), 
        .ZN(u5_mult_79_n506) );
  INV_X2 u5_mult_79_U1151 ( .A(u5_mult_79_n360), .ZN(u5_mult_79_n361) );
  INV_X1 u5_mult_79_U1150 ( .A(u5_mult_79_SUMB_21__10_), .ZN(u5_mult_79_n360)
         );
  XNOR2_X2 u5_mult_79_U1149 ( .A(u5_mult_79_n411), .B(u5_mult_79_n359), .ZN(
        u5_mult_79_SUMB_22__1_) );
  XNOR2_X2 u5_mult_79_U1148 ( .A(u5_mult_79_n397), .B(u5_mult_79_n296), .ZN(
        u5_mult_79_SUMB_11__8_) );
  NAND2_X2 u5_mult_79_U1147 ( .A1(u5_mult_79_ab_21__8_), .A2(
        u5_mult_79_CARRYB_20__8_), .ZN(u5_mult_79_n959) );
  CLKBUF_X3 u5_mult_79_U1146 ( .A(u5_mult_79_CARRYB_12__13_), .Z(
        u5_mult_79_n356) );
  XNOR2_X2 u5_mult_79_U1145 ( .A(u5_mult_79_ab_12__16_), .B(
        u5_mult_79_CARRYB_11__16_), .ZN(u5_mult_79_n576) );
  NAND3_X2 u5_mult_79_U1144 ( .A1(u5_mult_79_n672), .A2(u5_mult_79_n673), .A3(
        u5_mult_79_n674), .ZN(u5_mult_79_CARRYB_13__5_) );
  XNOR2_X2 u5_mult_79_U1143 ( .A(u5_mult_79_n355), .B(u5_mult_79_SUMB_3__14_), 
        .ZN(u5_mult_79_SUMB_4__13_) );
  XNOR2_X2 u5_mult_79_U1142 ( .A(u5_mult_79_n20), .B(u5_mult_79_n671), .ZN(
        u5_mult_79_n354) );
  XNOR2_X2 u5_mult_79_U1141 ( .A(u5_mult_79_SUMB_22__2_), .B(u5_mult_79_n353), 
        .ZN(u5_mult_79_SUMB_23__1_) );
  XNOR2_X2 u5_mult_79_U1140 ( .A(u5_mult_79_CARRYB_15__10_), .B(
        u5_mult_79_ab_16__10_), .ZN(u5_mult_79_n479) );
  XNOR2_X2 u5_mult_79_U1139 ( .A(u5_mult_79_n619), .B(u5_mult_79_n297), .ZN(
        u5_mult_79_SUMB_18__16_) );
  CLKBUF_X3 u5_mult_79_U1138 ( .A(u5_mult_79_SUMB_15__5_), .Z(u5_mult_79_n351)
         );
  NAND2_X2 u5_mult_79_U1137 ( .A1(u5_mult_79_ab_6__18_), .A2(
        u5_mult_79_SUMB_5__19_), .ZN(u5_mult_79_n611) );
  INV_X2 u5_mult_79_U1136 ( .A(u5_mult_79_n349), .ZN(u5_mult_79_n350) );
  INV_X1 u5_mult_79_U1135 ( .A(u5_mult_79_CARRYB_16__10_), .ZN(u5_mult_79_n349) );
  XNOR2_X2 u5_mult_79_U1134 ( .A(u5_mult_79_n348), .B(u5_mult_79_CARRYB_6__15_), .ZN(u5_mult_79_SUMB_7__15_) );
  XNOR2_X1 u5_mult_79_U1133 ( .A(u5_mult_79_CARRYB_15__3_), .B(
        u5_mult_79_ab_16__3_), .ZN(u5_mult_79_n544) );
  XNOR2_X2 u5_mult_79_U1132 ( .A(u5_mult_79_n346), .B(u5_mult_79_n308), .ZN(
        u5_mult_79_SUMB_10__9_) );
  XNOR2_X2 u5_mult_79_U1131 ( .A(u5_mult_79_ab_3__18_), .B(
        u5_mult_79_CARRYB_2__18_), .ZN(u5_mult_79_n345) );
  XNOR2_X2 u5_mult_79_U1130 ( .A(u5_mult_79_n345), .B(u5_mult_79_SUMB_2__19_), 
        .ZN(u5_mult_79_SUMB_3__18_) );
  XNOR2_X2 u5_mult_79_U1129 ( .A(u5_mult_79_n344), .B(u5_mult_79_SUMB_12__7_), 
        .ZN(u5_mult_79_SUMB_13__6_) );
  INV_X4 u5_mult_79_U1128 ( .A(u5_mult_79_n342), .ZN(u5_mult_79_n343) );
  INV_X2 u5_mult_79_U1127 ( .A(u5_mult_79_SUMB_19__1_), .ZN(u5_mult_79_n342)
         );
  CLKBUF_X2 u5_mult_79_U1126 ( .A(u5_mult_79_SUMB_2__21_), .Z(u5_mult_79_n341)
         );
  XNOR2_X2 u5_mult_79_U1125 ( .A(u5_mult_79_CARRYB_7__12_), .B(
        u5_mult_79_ab_8__12_), .ZN(u5_mult_79_n595) );
  XNOR2_X2 u5_mult_79_U1124 ( .A(u5_mult_79_CARRYB_15__11_), .B(
        u5_mult_79_n1316), .ZN(u5_mult_79_n340) );
  XOR2_X2 u5_mult_79_U1123 ( .A(u5_mult_79_n340), .B(u5_mult_79_SUMB_15__12_), 
        .Z(u5_mult_79_SUMB_16__11_) );
  XNOR2_X2 u5_mult_79_U1122 ( .A(u5_mult_79_CARRYB_9__9_), .B(
        u5_mult_79_ab_10__9_), .ZN(u5_mult_79_n346) );
  INV_X2 u5_mult_79_U1121 ( .A(u5_mult_79_n338), .ZN(u5_mult_79_n339) );
  INV_X1 u5_mult_79_U1120 ( .A(u5_mult_79_CARRYB_22__0_), .ZN(u5_mult_79_n338)
         );
  INV_X4 u5_mult_79_U1119 ( .A(u5_mult_79_n336), .ZN(u5_mult_79_n337) );
  INV_X2 u5_mult_79_U1118 ( .A(u5_mult_79_CARRYB_2__20_), .ZN(u5_mult_79_n336)
         );
  NAND2_X2 u5_mult_79_U1117 ( .A1(u5_mult_79_ab_12__8_), .A2(u5_mult_79_n116), 
        .ZN(u5_mult_79_n993) );
  NAND2_X2 u5_mult_79_U1116 ( .A1(u5_mult_79_n48), .A2(u5_mult_79_n116), .ZN(
        u5_mult_79_n994) );
  NAND3_X4 u5_mult_79_U1115 ( .A1(u5_mult_79_n992), .A2(u5_mult_79_n993), .A3(
        u5_mult_79_n994), .ZN(u5_mult_79_CARRYB_12__8_) );
  CLKBUF_X3 u5_mult_79_U1114 ( .A(u5_mult_79_SUMB_16__19_), .Z(u5_mult_79_n373) );
  CLKBUF_X2 u5_mult_79_U1113 ( .A(u5_mult_79_SUMB_17__18_), .Z(u5_mult_79_n334) );
  XNOR2_X2 u5_mult_79_U1112 ( .A(u5_mult_79_ab_10__19_), .B(
        u5_mult_79_CARRYB_9__19_), .ZN(u5_mult_79_n332) );
  XNOR2_X2 u5_mult_79_U1111 ( .A(u5_mult_79_n332), .B(u5_mult_79_n323), .ZN(
        u5_mult_79_SUMB_10__19_) );
  XNOR2_X2 u5_mult_79_U1110 ( .A(u5_mult_79_n330), .B(u5_mult_79_SUMB_15__18_), 
        .ZN(u5_mult_79_SUMB_16__17_) );
  XNOR2_X2 u5_mult_79_U1109 ( .A(u5_mult_79_CARRYB_21__1_), .B(
        u5_mult_79_ab_22__1_), .ZN(u5_mult_79_n359) );
  XOR2_X2 u5_mult_79_U1108 ( .A(u5_mult_79_n798), .B(u5_mult_79_CARRYB_13__16_), .Z(u5_mult_79_n329) );
  XNOR2_X2 u5_mult_79_U1107 ( .A(u5_mult_79_n329), .B(u5_mult_79_n484), .ZN(
        u5_mult_79_SUMB_14__16_) );
  XNOR2_X2 u5_mult_79_U1106 ( .A(u5_mult_79_CARRYB_18__11_), .B(
        u5_mult_79_ab_19__11_), .ZN(u5_mult_79_n328) );
  XNOR2_X2 u5_mult_79_U1105 ( .A(u5_mult_79_SUMB_18__12_), .B(u5_mult_79_n328), 
        .ZN(u5_mult_79_SUMB_19__11_) );
  NAND2_X1 u5_mult_79_U1104 ( .A1(u5_mult_79_ab_19__4_), .A2(
        u5_mult_79_CARRYB_18__4_), .ZN(u5_mult_79_n1590) );
  XNOR2_X2 u5_mult_79_U1103 ( .A(u5_mult_79_CARRYB_9__18_), .B(
        u5_mult_79_ab_10__18_), .ZN(u5_mult_79_n327) );
  XNOR2_X2 u5_mult_79_U1102 ( .A(u5_mult_79_SUMB_9__19_), .B(u5_mult_79_n327), 
        .ZN(u5_mult_79_SUMB_10__18_) );
  INV_X4 u5_mult_79_U1101 ( .A(u5_mult_79_n363), .ZN(u5_mult_79_n364) );
  CLKBUF_X3 u5_mult_79_U1100 ( .A(u5_mult_79_SUMB_2__13_), .Z(u5_mult_79_n326)
         );
  XNOR2_X2 u5_mult_79_U1099 ( .A(u5_mult_79_n1705), .B(u5_mult_79_n1181), .ZN(
        u5_mult_79_n324) );
  CLKBUF_X2 u5_mult_79_U1098 ( .A(u5_mult_79_SUMB_9__20_), .Z(u5_mult_79_n323)
         );
  XOR2_X2 u5_mult_79_U1097 ( .A(u5_mult_79_n1401), .B(u5_mult_79_n307), .Z(
        u5_mult_79_n322) );
  BUF_X8 u5_mult_79_U1096 ( .A(u5_mult_79_SUMB_19__4_), .Z(u5_mult_79_n321) );
  CLKBUF_X2 u5_mult_79_U1095 ( .A(u5_mult_79_SUMB_11__17_), .Z(u5_mult_79_n320) );
  NAND2_X2 u5_mult_79_U1094 ( .A1(u5_mult_79_ab_18__9_), .A2(u5_mult_79_n558), 
        .ZN(u5_mult_79_n560) );
  XNOR2_X2 u5_mult_79_U1093 ( .A(u5_mult_79_CARRYB_4__19_), .B(u5_mult_79_n319), .ZN(u5_mult_79_SUMB_5__19_) );
  INV_X2 u5_mult_79_U1092 ( .A(u5_mult_79_n317), .ZN(u5_mult_79_n318) );
  INV_X1 u5_mult_79_U1091 ( .A(u5_mult_79_SUMB_8__17_), .ZN(u5_mult_79_n317)
         );
  XNOR2_X2 u5_mult_79_U1090 ( .A(u5_mult_79_ab_11__10_), .B(
        u5_mult_79_CARRYB_10__10_), .ZN(u5_mult_79_n467) );
  NAND2_X2 u5_mult_79_U1089 ( .A1(u5_mult_79_ab_22__12_), .A2(
        u5_mult_79_CARRYB_21__12_), .ZN(u5_mult_79_n1055) );
  NAND2_X4 u5_mult_79_U1088 ( .A1(u5_mult_79_ab_20__0_), .A2(u5_mult_79_n343), 
        .ZN(u5_mult_79_n651) );
  BUF_X8 u5_mult_79_U1087 ( .A(u5_mult_79_SUMB_11__8_), .Z(u5_mult_79_n316) );
  BUF_X8 u5_mult_79_U1086 ( .A(u5_mult_79_SUMB_20__4_), .Z(u5_mult_79_n315) );
  CLKBUF_X3 u5_mult_79_U1085 ( .A(u5_mult_79_SUMB_4__21_), .Z(u5_mult_79_n314)
         );
  XNOR2_X1 u5_mult_79_U1084 ( .A(u5_mult_79_ab_17__10_), .B(
        u5_mult_79_CARRYB_16__10_), .ZN(u5_mult_79_n313) );
  XNOR2_X2 u5_mult_79_U1083 ( .A(u5_mult_79_n313), .B(u5_mult_79_n335), .ZN(
        u5_mult_79_SUMB_17__10_) );
  INV_X2 u5_mult_79_U1082 ( .A(u5_mult_79_n310), .ZN(u5_mult_79_n311) );
  XNOR2_X2 u5_mult_79_U1081 ( .A(u5_mult_79_CARRYB_5__19_), .B(
        u5_mult_79_ab_6__19_), .ZN(u5_mult_79_n309) );
  XNOR2_X2 u5_mult_79_U1080 ( .A(u5_mult_79_SUMB_5__20_), .B(u5_mult_79_n309), 
        .ZN(u5_mult_79_SUMB_6__19_) );
  XNOR2_X2 u5_mult_79_U1079 ( .A(u5_mult_79_n486), .B(u5_mult_79_SUMB_5__19_), 
        .ZN(u5_mult_79_SUMB_6__18_) );
  CLKBUF_X3 u5_mult_79_U1078 ( .A(u5_mult_79_SUMB_6__18_), .Z(u5_mult_79_n482)
         );
  NAND2_X2 u5_mult_79_U1077 ( .A1(u5_mult_79_ab_7__20_), .A2(
        u5_mult_79_CARRYB_6__20_), .ZN(u5_mult_79_n1229) );
  CLKBUF_X3 u5_mult_79_U1076 ( .A(u5_mult_79_SUMB_11__12_), .Z(u5_mult_79_n307) );
  INV_X1 u5_mult_79_U1075 ( .A(u5_mult_79_CARRYB_18__2_), .ZN(u5_mult_79_n306)
         );
  XNOR2_X2 u5_mult_79_U1074 ( .A(u5_mult_79_n578), .B(u5_mult_79_SUMB_4__19_), 
        .ZN(u5_mult_79_n305) );
  CLKBUF_X2 u5_mult_79_U1073 ( .A(u5_mult_79_CARRYB_20__6_), .Z(
        u5_mult_79_n304) );
  NAND2_X2 u5_mult_79_U1072 ( .A1(u5_mult_79_ab_17__9_), .A2(
        u5_mult_79_CARRYB_16__9_), .ZN(u5_mult_79_n1495) );
  CLKBUF_X3 u5_mult_79_U1071 ( .A(u5_mult_79_SUMB_7__22_), .Z(u5_mult_79_n303)
         );
  INV_X2 u5_mult_79_U1070 ( .A(u5_mult_79_SUMB_9__13_), .ZN(u5_mult_79_n310)
         );
  CLKBUF_X3 u5_mult_79_U1069 ( .A(u5_mult_79_SUMB_11__16_), .Z(u5_mult_79_n302) );
  XNOR2_X2 u5_mult_79_U1068 ( .A(u5_mult_79_CARRYB_4__20_), .B(
        u5_mult_79_ab_5__20_), .ZN(u5_mult_79_n301) );
  XNOR2_X2 u5_mult_79_U1067 ( .A(u5_mult_79_n314), .B(u5_mult_79_n301), .ZN(
        u5_mult_79_SUMB_5__20_) );
  XOR2_X2 u5_mult_79_U1066 ( .A(u5_mult_79_n362), .B(u5_mult_79_CARRYB_10__18_), .Z(u5_mult_79_n299) );
  XNOR2_X2 u5_mult_79_U1065 ( .A(u5_mult_79_n299), .B(u5_mult_79_SUMB_10__19_), 
        .ZN(u5_mult_79_SUMB_11__18_) );
  CLKBUF_X3 u5_mult_79_U1064 ( .A(u5_mult_79_CARRYB_20__5_), .Z(
        u5_mult_79_n457) );
  XOR2_X2 u5_mult_79_U1063 ( .A(u5_mult_79_CARRYB_20__5_), .B(u5_mult_79_n522), 
        .Z(u5_mult_79_n298) );
  XNOR2_X2 u5_mult_79_U1062 ( .A(u5_mult_79_n298), .B(u5_mult_79_n466), .ZN(
        u5_mult_79_SUMB_21__5_) );
  NAND2_X2 u5_mult_79_U1061 ( .A1(u5_mult_79_CARRYB_6__17_), .A2(
        u5_mult_79_SUMB_6__18_), .ZN(u5_mult_79_n615) );
  NAND2_X4 u5_mult_79_U1060 ( .A1(u5_mult_79_n286), .A2(
        u5_mult_79_CARRYB_13__9_), .ZN(u5_mult_79_n1327) );
  NAND2_X4 u5_mult_79_U1059 ( .A1(u5_mult_79_SUMB_13__10_), .A2(
        u5_mult_79_ab_14__9_), .ZN(u5_mult_79_n1328) );
  BUF_X8 u5_mult_79_U1058 ( .A(u5_mult_79_SUMB_17__17_), .Z(u5_mult_79_n297)
         );
  NAND3_X2 u5_mult_79_U1057 ( .A1(u5_mult_79_n880), .A2(u5_mult_79_n881), .A3(
        u5_mult_79_n882), .ZN(u5_mult_79_CARRYB_5__7_) );
  CLKBUF_X3 u5_mult_79_U1056 ( .A(u5_mult_79_SUMB_5__21_), .Z(u5_mult_79_n395)
         );
  XNOR2_X1 u5_mult_79_U1055 ( .A(u5_mult_79_n346), .B(u5_mult_79_n308), .ZN(
        u5_mult_79_n296) );
  XNOR2_X2 u5_mult_79_U1054 ( .A(u5_mult_79_n346), .B(u5_mult_79_n308), .ZN(
        u5_mult_79_n295) );
  XNOR2_X2 u5_mult_79_U1053 ( .A(u5_mult_79_n292), .B(u5_mult_79_n476), .ZN(
        u5_mult_79_n294) );
  NAND3_X2 u5_mult_79_U1052 ( .A1(u5_mult_79_n1422), .A2(u5_mult_79_n1423), 
        .A3(u5_mult_79_n1421), .ZN(u5_mult_79_CARRYB_12__12_) );
  XOR2_X2 u5_mult_79_U1051 ( .A(u5_mult_79_ab_14__12_), .B(
        u5_mult_79_CARRYB_13__12_), .Z(u5_mult_79_n293) );
  XNOR2_X2 u5_mult_79_U1050 ( .A(u5_mult_79_n293), .B(u5_mult_79_n228), .ZN(
        u5_mult_79_SUMB_14__12_) );
  INV_X4 u5_mult_79_U1049 ( .A(u5_mult_79_CARRYB_5__22_), .ZN(u5_mult_79_n497)
         );
  XNOR2_X2 u5_mult_79_U1048 ( .A(u5_mult_79_n497), .B(u5_mult_79_n241), .ZN(
        u5_mult_79_SUMB_6__22_) );
  XNOR2_X2 u5_mult_79_U1047 ( .A(u5_mult_79_n442), .B(u5_mult_79_ab_14__15_), 
        .ZN(u5_mult_79_n292) );
  INV_X2 u5_mult_79_U1046 ( .A(u5_mult_79_n290), .ZN(u5_mult_79_n291) );
  INV_X1 u5_mult_79_U1045 ( .A(u5_mult_79_SUMB_7__16_), .ZN(u5_mult_79_n290)
         );
  INV_X4 u5_mult_79_U1044 ( .A(u5_mult_79_n289), .ZN(u5_mult_79_SUMB_7__8_) );
  XNOR2_X2 u5_mult_79_U1043 ( .A(u5_mult_79_n1164), .B(u5_mult_79_SUMB_6__9_), 
        .ZN(u5_mult_79_n289) );
  XNOR2_X2 u5_mult_79_U1042 ( .A(u5_mult_79_CARRYB_5__20_), .B(
        u5_mult_79_ab_6__20_), .ZN(u5_mult_79_n379) );
  INV_X2 u5_mult_79_U1041 ( .A(u5_mult_79_CARRYB_2__11_), .ZN(u5_mult_79_n287)
         );
  XNOR2_X2 u5_mult_79_U1040 ( .A(u5_mult_79_CARRYB_12__10_), .B(
        u5_mult_79_n858), .ZN(u5_mult_79_n286) );
  XOR2_X2 u5_mult_79_U1039 ( .A(u5_mult_79_n695), .B(u5_mult_79_SUMB_4__13_), 
        .Z(u5_mult_79_n285) );
  INV_X4 u5_mult_79_U1038 ( .A(u5_mult_79_SUMB_3__22_), .ZN(u5_mult_79_n283)
         );
  INV_X4 u5_mult_79_U1037 ( .A(u5_mult_79_n281), .ZN(u5_mult_79_n282) );
  INV_X2 u5_mult_79_U1036 ( .A(u5_mult_79_SUMB_4__22_), .ZN(u5_mult_79_n281)
         );
  NAND3_X2 u5_mult_79_U1035 ( .A1(u5_mult_79_n1309), .A2(u5_mult_79_n1310), 
        .A3(u5_mult_79_n1311), .ZN(u5_mult_79_CARRYB_23__10_) );
  XNOR2_X2 u5_mult_79_U1034 ( .A(u5_mult_79_n315), .B(u5_mult_79_n475), .ZN(
        u5_mult_79_n280) );
  INV_X2 u5_mult_79_U1033 ( .A(u5_mult_79_n278), .ZN(u5_mult_79_n279) );
  INV_X1 u5_mult_79_U1032 ( .A(u5_mult_79_n269), .ZN(u5_mult_79_n278) );
  INV_X4 u5_mult_79_U1031 ( .A(u5_mult_79_n276), .ZN(u5_mult_79_n277) );
  INV_X2 u5_mult_79_U1030 ( .A(u5_mult_79_CARRYB_14__6_), .ZN(u5_mult_79_n276)
         );
  INV_X2 u5_mult_79_U1029 ( .A(u5_mult_79_n274), .ZN(u5_mult_79_n275) );
  INV_X1 u5_mult_79_U1028 ( .A(u5_mult_79_SUMB_15__7_), .ZN(u5_mult_79_n274)
         );
  NAND3_X2 u5_mult_79_U1027 ( .A1(u5_mult_79_n1041), .A2(u5_mult_79_n1042), 
        .A3(u5_mult_79_n1043), .ZN(u5_mult_79_CARRYB_18__12_) );
  CLKBUF_X2 u5_mult_79_U1026 ( .A(u5_mult_79_SUMB_12__5_), .Z(u5_mult_79_n273)
         );
  XNOR2_X2 u5_mult_79_U1025 ( .A(u5_mult_79_SUMB_18__11_), .B(u5_mult_79_n1246), .ZN(u5_mult_79_n333) );
  NAND2_X2 u5_mult_79_U1024 ( .A1(u5_mult_79_ab_7__17_), .A2(
        u5_mult_79_CARRYB_6__17_), .ZN(u5_mult_79_n613) );
  NAND2_X1 u5_mult_79_U1023 ( .A1(u5_mult_79_ab_4__18_), .A2(
        u5_mult_79_SUMB_3__19_), .ZN(u5_mult_79_n1580) );
  NAND2_X2 u5_mult_79_U1022 ( .A1(u5_mult_79_SUMB_10__17_), .A2(
        u5_mult_79_CARRYB_10__16_), .ZN(u5_mult_79_n821) );
  NAND3_X4 u5_mult_79_U1021 ( .A1(u5_mult_79_n1600), .A2(u5_mult_79_n1601), 
        .A3(u5_mult_79_n1602), .ZN(u5_mult_79_CARRYB_3__21_) );
  NAND2_X2 u5_mult_79_U1020 ( .A1(u5_mult_79_ab_21__6_), .A2(u5_mult_79_n304), 
        .ZN(u5_mult_79_n1559) );
  NAND2_X2 u5_mult_79_U1019 ( .A1(u5_mult_79_n354), .A2(u5_mult_79_ab_17__7_), 
        .ZN(u5_mult_79_n1592) );
  XNOR2_X2 u5_mult_79_U1018 ( .A(u5_mult_79_CARRYB_17__15_), .B(
        u5_mult_79_ab_18__15_), .ZN(u5_mult_79_n272) );
  NAND2_X1 u5_mult_79_U1017 ( .A1(u5_mult_79_ab_12__17_), .A2(
        u5_mult_79_SUMB_11__18_), .ZN(u5_mult_79_n984) );
  NAND2_X2 u5_mult_79_U1016 ( .A1(u5_mult_79_ab_10__18_), .A2(
        u5_mult_79_SUMB_9__19_), .ZN(u5_mult_79_n980) );
  XNOR2_X2 u5_mult_79_U1015 ( .A(u5_mult_79_CARRYB_6__12_), .B(
        u5_mult_79_ab_7__12_), .ZN(u5_mult_79_n271) );
  XNOR2_X2 u5_mult_79_U1014 ( .A(u5_mult_79_SUMB_6__13_), .B(u5_mult_79_n271), 
        .ZN(u5_mult_79_SUMB_7__12_) );
  INV_X2 u5_mult_79_U1013 ( .A(u5_mult_79_n287), .ZN(u5_mult_79_n288) );
  XNOR2_X2 u5_mult_79_U1012 ( .A(u5_mult_79_CARRYB_5__10_), .B(u5_mult_79_n270), .ZN(u5_mult_79_n835) );
  XNOR2_X2 u5_mult_79_U1011 ( .A(u5_mult_79_n287), .B(u5_mult_79_ab_3__11_), 
        .ZN(u5_mult_79_n712) );
  NAND2_X4 u5_mult_79_U1010 ( .A1(u5_mult_79_ab_3__16_), .A2(u5_mult_79_n488), 
        .ZN(u5_mult_79_n1378) );
  NOR2_X4 u5_mult_79_U1009 ( .A1(u5_mult_79_n1880), .A2(u5_mult_79_n1882), 
        .ZN(u5_mult_79_n623) );
  NAND3_X2 u5_mult_79_U1008 ( .A1(u5_mult_79_n1379), .A2(u5_mult_79_n1378), 
        .A3(u5_mult_79_n1377), .ZN(u5_mult_79_n269) );
  NAND2_X2 u5_mult_79_U1007 ( .A1(u5_mult_79_CARRYB_10__5_), .A2(
        u5_mult_79_n404), .ZN(u5_mult_79_n1112) );
  NAND3_X4 u5_mult_79_U1006 ( .A1(u5_mult_79_n1112), .A2(u5_mult_79_n1113), 
        .A3(u5_mult_79_n1114), .ZN(u5_mult_79_CARRYB_11__5_) );
  INV_X16 u5_mult_79_U1005 ( .A(n2969), .ZN(u5_mult_79_n1867) );
  NAND3_X2 u5_mult_79_U1004 ( .A1(u5_mult_79_n1415), .A2(u5_mult_79_n1417), 
        .A3(u5_mult_79_n1416), .ZN(u5_mult_79_n268) );
  CLKBUF_X3 u5_mult_79_U1003 ( .A(u5_mult_79_CARRYB_21__6_), .Z(
        u5_mult_79_n267) );
  CLKBUF_X2 u5_mult_79_U1002 ( .A(u5_mult_79_CARRYB_2__17_), .Z(
        u5_mult_79_n266) );
  NAND2_X4 u5_mult_79_U1001 ( .A1(u5_mult_79_n387), .A2(u5_mult_79_ab_5__6_), 
        .ZN(u5_mult_79_n791) );
  NAND2_X2 u5_mult_79_U1000 ( .A1(u5_mult_79_ab_6__16_), .A2(
        u5_mult_79_SUMB_5__17_), .ZN(u5_mult_79_n1586) );
  NAND2_X2 u5_mult_79_U999 ( .A1(u5_mult_79_SUMB_5__17_), .A2(
        u5_mult_79_CARRYB_5__16_), .ZN(u5_mult_79_n1587) );
  NAND2_X2 u5_mult_79_U998 ( .A1(u5_mult_79_ab_16__7_), .A2(
        u5_mult_79_SUMB_15__8_), .ZN(u5_mult_79_n1481) );
  NAND2_X2 u5_mult_79_U997 ( .A1(u5_mult_79_ab_0__17_), .A2(
        u5_mult_79_ab_1__16_), .ZN(u5_mult_79_n1705) );
  NAND2_X4 u5_mult_79_U996 ( .A1(u5_mult_79_ab_22__1_), .A2(
        u5_mult_79_CARRYB_21__1_), .ZN(u5_mult_79_n1177) );
  XNOR2_X1 u5_mult_79_U995 ( .A(u5_mult_79_CARRYB_6__6_), .B(
        u5_mult_79_ab_7__6_), .ZN(u5_mult_79_n907) );
  XNOR2_X2 u5_mult_79_U994 ( .A(u5_mult_79_SUMB_6__7_), .B(u5_mult_79_n907), 
        .ZN(u5_mult_79_SUMB_7__6_) );
  XNOR2_X2 u5_mult_79_U993 ( .A(u5_mult_79_ab_9__15_), .B(
        u5_mult_79_CARRYB_8__15_), .ZN(u5_mult_79_n264) );
  XNOR2_X2 u5_mult_79_U992 ( .A(u5_mult_79_n264), .B(u5_mult_79_SUMB_8__16_), 
        .ZN(u5_mult_79_SUMB_9__15_) );
  NAND2_X2 u5_mult_79_U991 ( .A1(u5_mult_79_SUMB_3__15_), .A2(
        u5_mult_79_CARRYB_3__14_), .ZN(u5_mult_79_n1342) );
  INV_X4 u5_mult_79_U990 ( .A(u5_mult_79_n1657), .ZN(u5_mult_79_CLA_SUM[33])
         );
  XNOR2_X2 u5_mult_79_U989 ( .A(u5_mult_79_n303), .B(u5_mult_79_n263), .ZN(
        u5_mult_79_SUMB_8__21_) );
  NAND3_X4 u5_mult_79_U988 ( .A1(u5_mult_79_n1324), .A2(u5_mult_79_n1325), 
        .A3(u5_mult_79_n1326), .ZN(u5_mult_79_CARRYB_8__13_) );
  NAND2_X1 u5_mult_79_U987 ( .A1(u5_mult_79_CARRYB_13__4_), .A2(
        u5_mult_79_SUMB_13__5_), .ZN(u5_mult_79_n677) );
  XNOR2_X2 u5_mult_79_U986 ( .A(u5_mult_79_ab_13__5_), .B(
        u5_mult_79_CARRYB_12__5_), .ZN(u5_mult_79_n431) );
  XOR2_X2 u5_mult_79_U985 ( .A(u5_mult_79_n340), .B(u5_mult_79_n14), .Z(
        u5_mult_79_n335) );
  NAND2_X2 u5_mult_79_U984 ( .A1(u5_mult_79_CARRYB_10__3_), .A2(
        u5_mult_79_ab_11__3_), .ZN(u5_mult_79_n887) );
  NAND2_X2 u5_mult_79_U983 ( .A1(u5_mult_79_CARRYB_10__3_), .A2(
        u5_mult_79_SUMB_10__4_), .ZN(u5_mult_79_n886) );
  INV_X8 u5_mult_79_U982 ( .A(n2769), .ZN(u5_mult_79_n1872) );
  BUF_X4 u5_mult_79_U981 ( .A(u5_mult_79_CARRYB_4__6_), .Z(u5_mult_79_n262) );
  XNOR2_X1 u5_mult_79_U980 ( .A(u5_mult_79_ab_5__11_), .B(
        u5_mult_79_CARRYB_4__11_), .ZN(u5_mult_79_n261) );
  XNOR2_X2 u5_mult_79_U979 ( .A(u5_mult_79_n261), .B(u5_mult_79_SUMB_4__12_), 
        .ZN(u5_mult_79_SUMB_5__11_) );
  XNOR2_X2 u5_mult_79_U978 ( .A(u5_mult_79_CARRYB_14__7_), .B(
        u5_mult_79_ab_15__7_), .ZN(u5_mult_79_n513) );
  INV_X16 u5_mult_79_U977 ( .A(u5_mult_79_n1865), .ZN(u5_mult_79_n1795) );
  NAND2_X2 u5_mult_79_U976 ( .A1(u5_mult_79_ab_14__2_), .A2(
        u5_mult_79_CARRYB_13__2_), .ZN(u5_mult_79_n926) );
  NAND2_X2 u5_mult_79_U975 ( .A1(u5_mult_79_CARRYB_11__2_), .A2(
        u5_mult_79_SUMB_11__3_), .ZN(u5_mult_79_n931) );
  NAND3_X2 u5_mult_79_U974 ( .A1(u5_mult_79_n1298), .A2(u5_mult_79_n1297), 
        .A3(u5_mult_79_n1296), .ZN(u5_mult_79_CARRYB_10__12_) );
  NAND3_X2 u5_mult_79_U973 ( .A1(u5_mult_79_n855), .A2(u5_mult_79_n856), .A3(
        u5_mult_79_n857), .ZN(u5_mult_79_CARRYB_7__15_) );
  NAND2_X1 u5_mult_79_U972 ( .A1(u5_mult_79_CARRYB_5__15_), .A2(
        u5_mult_79_SUMB_5__16_), .ZN(u5_mult_79_n1539) );
  NAND2_X2 u5_mult_79_U971 ( .A1(u5_mult_79_ab_6__20_), .A2(
        u5_mult_79_CARRYB_5__20_), .ZN(u5_mult_79_n902) );
  NAND2_X2 u5_mult_79_U970 ( .A1(u5_mult_79_SUMB_5__21_), .A2(
        u5_mult_79_ab_6__20_), .ZN(u5_mult_79_n901) );
  XNOR2_X2 u5_mult_79_U969 ( .A(u5_mult_79_n260), .B(u5_mult_79_SUMB_21__9_), 
        .ZN(u5_mult_79_SUMB_22__8_) );
  NAND2_X1 u5_mult_79_U968 ( .A1(u5_mult_79_CARRYB_8__5_), .A2(
        u5_mult_79_SUMB_8__6_), .ZN(u5_mult_79_n1021) );
  NAND2_X2 u5_mult_79_U967 ( .A1(u5_mult_79_ab_12__7_), .A2(
        u5_mult_79_CARRYB_11__7_), .ZN(u5_mult_79_n1096) );
  NOR2_X2 u5_mult_79_U966 ( .A1(u5_mult_79_n1882), .A2(u5_mult_79_n1867), .ZN(
        u5_mult_79_ab_0__14_) );
  NAND2_X2 u5_mult_79_U965 ( .A1(u5_mult_79_ab_0__14_), .A2(
        u5_mult_79_ab_1__13_), .ZN(u5_mult_79_n1699) );
  NAND3_X2 u5_mult_79_U964 ( .A1(u5_mult_79_n583), .A2(u5_mult_79_n584), .A3(
        u5_mult_79_n585), .ZN(u5_mult_79_CARRYB_22__3_) );
  NAND2_X2 u5_mult_79_U963 ( .A1(u5_mult_79_n381), .A2(u5_mult_79_ab_21__6_), 
        .ZN(u5_mult_79_n1560) );
  NAND2_X2 u5_mult_79_U962 ( .A1(u5_mult_79_SUMB_3__15_), .A2(
        u5_mult_79_ab_4__14_), .ZN(u5_mult_79_n1341) );
  NAND2_X2 u5_mult_79_U961 ( .A1(u5_mult_79_ab_13__4_), .A2(u5_mult_79_n372), 
        .ZN(u5_mult_79_n875) );
  NAND2_X1 u5_mult_79_U960 ( .A1(u5_mult_79_ab_10__4_), .A2(
        u5_mult_79_SUMB_9__5_), .ZN(u5_mult_79_n1023) );
  XNOR2_X2 u5_mult_79_U959 ( .A(u5_mult_79_n415), .B(u5_mult_79_n399), .ZN(
        u5_mult_79_n259) );
  NAND2_X2 u5_mult_79_U958 ( .A1(u5_mult_79_CARRYB_23__1_), .A2(
        u5_mult_79_SUMB_23__2_), .ZN(u5_mult_79_n1646) );
  CLKBUF_X2 u5_mult_79_U957 ( .A(u5_mult_79_CARRYB_20__1_), .Z(u5_mult_79_n258) );
  INV_X4 u5_mult_79_U956 ( .A(u5_mult_79_n1504), .ZN(u5_mult_79_n1257) );
  XNOR2_X2 u5_mult_79_U955 ( .A(u5_mult_79_n277), .B(u5_mult_79_ab_15__6_), 
        .ZN(u5_mult_79_n776) );
  XNOR2_X2 u5_mult_79_U954 ( .A(u5_mult_79_SUMB_17__4_), .B(
        u5_mult_79_ab_18__3_), .ZN(u5_mult_79_n399) );
  CLKBUF_X3 u5_mult_79_U953 ( .A(u5_mult_79_CARRYB_17__3_), .Z(u5_mult_79_n415) );
  XNOR2_X2 u5_mult_79_U952 ( .A(u5_mult_79_CARRYB_8__5_), .B(
        u5_mult_79_ab_9__5_), .ZN(u5_mult_79_n257) );
  XNOR2_X2 u5_mult_79_U951 ( .A(u5_mult_79_n257), .B(u5_mult_79_SUMB_8__6_), 
        .ZN(u5_mult_79_SUMB_9__5_) );
  XNOR2_X2 u5_mult_79_U950 ( .A(u5_mult_79_n273), .B(u5_mult_79_n256), .ZN(
        u5_mult_79_SUMB_13__4_) );
  XNOR2_X2 u5_mult_79_U949 ( .A(u5_mult_79_ab_6__6_), .B(
        u5_mult_79_CARRYB_5__6_), .ZN(u5_mult_79_n255) );
  XNOR2_X1 u5_mult_79_U948 ( .A(u5_mult_79_n255), .B(u5_mult_79_SUMB_5__7_), 
        .ZN(u5_mult_79_SUMB_6__6_) );
  XNOR2_X2 u5_mult_79_U947 ( .A(u5_mult_79_ab_4__13_), .B(
        u5_mult_79_CARRYB_3__13_), .ZN(u5_mult_79_n355) );
  NAND2_X2 u5_mult_79_U946 ( .A1(u5_mult_79_CARRYB_23__0_), .A2(
        u5_mult_79_SUMB_23__1_), .ZN(u5_mult_79_n1645) );
  INV_X4 u5_mult_79_U945 ( .A(u5_mult_79_n1645), .ZN(u5_mult_79_CLA_CARRY[24])
         );
  NAND3_X4 u5_mult_79_U944 ( .A1(u5_mult_79_n505), .A2(u5_mult_79_n506), .A3(
        u5_mult_79_n507), .ZN(u5_mult_79_CARRYB_11__8_) );
  NAND2_X2 u5_mult_79_U943 ( .A1(u5_mult_79_ab_11__8_), .A2(u5_mult_79_n406), 
        .ZN(u5_mult_79_n505) );
  NAND2_X1 u5_mult_79_U942 ( .A1(u5_mult_79_SUMB_17__4_), .A2(
        u5_mult_79_CARRYB_17__3_), .ZN(u5_mult_79_n1178) );
  XOR2_X2 u5_mult_79_U941 ( .A(u5_mult_79_n1171), .B(u5_mult_79_n339), .Z(
        u5_N23) );
  INV_X8 u5_mult_79_U940 ( .A(n2523), .ZN(u5_mult_79_n1873) );
  NAND2_X2 u5_mult_79_U939 ( .A1(u5_mult_79_ab_23__1_), .A2(
        u5_mult_79_CARRYB_22__1_), .ZN(u5_mult_79_n510) );
  XNOR2_X2 u5_mult_79_U938 ( .A(u5_mult_79_CARRYB_22__1_), .B(
        u5_mult_79_ab_23__1_), .ZN(u5_mult_79_n353) );
  XNOR2_X2 u5_mult_79_U937 ( .A(u5_mult_79_n253), .B(u5_mult_79_n254), .ZN(
        u5_mult_79_n1171) );
  XNOR2_X2 u5_mult_79_U936 ( .A(u5_mult_79_n359), .B(u5_mult_79_n411), .ZN(
        u5_mult_79_n253) );
  XNOR2_X2 u5_mult_79_U935 ( .A(u5_mult_79_ab_13__6_), .B(
        u5_mult_79_CARRYB_12__6_), .ZN(u5_mult_79_n344) );
  INV_X1 u5_mult_79_U934 ( .A(u5_mult_79_CARRYB_18__0_), .ZN(u5_mult_79_n252)
         );
  XNOR2_X1 u5_mult_79_U933 ( .A(u5_mult_79_CARRYB_13__2_), .B(
        u5_mult_79_ab_14__2_), .ZN(u5_mult_79_n251) );
  XNOR2_X1 u5_mult_79_U932 ( .A(u5_mult_79_SUMB_15__2_), .B(
        u5_mult_79_ab_16__1_), .ZN(u5_mult_79_n248) );
  XNOR2_X2 u5_mult_79_U931 ( .A(u5_mult_79_n248), .B(u5_mult_79_CARRYB_15__1_), 
        .ZN(u5_mult_79_SUMB_16__1_) );
  XOR2_X2 u5_mult_79_U930 ( .A(u5_mult_79_n664), .B(u5_mult_79_CARRYB_13__1_), 
        .Z(u5_mult_79_SUMB_14__1_) );
  NAND2_X2 u5_mult_79_U929 ( .A1(u5_mult_79_CARRYB_13__0_), .A2(
        u5_mult_79_SUMB_13__1_), .ZN(u5_mult_79_n947) );
  XNOR2_X2 u5_mult_79_U928 ( .A(u5_mult_79_n247), .B(u5_mult_79_SUMB_16__1_), 
        .ZN(u5_mult_79_n938) );
  XOR2_X1 u5_mult_79_U927 ( .A(u5_mult_79_ab_1__0_), .B(u5_mult_79_ab_0__1_), 
        .Z(u5_N1) );
  INV_X4 u5_mult_79_U926 ( .A(u5_mult_79_ab_18__14_), .ZN(u5_mult_79_n965) );
  INV_X4 u5_mult_79_U925 ( .A(u5_mult_79_ab_17__8_), .ZN(u5_mult_79_n1458) );
  INV_X4 u5_mult_79_U924 ( .A(u5_mult_79_ab_18__9_), .ZN(u5_mult_79_n1514) );
  INV_X16 u5_mult_79_U923 ( .A(u5_mult_79_n1774), .ZN(u5_mult_79_n1773) );
  INV_X4 u5_mult_79_U922 ( .A(u5_mult_79_n1855), .ZN(u5_mult_79_n1774) );
  INV_X8 u5_mult_79_U921 ( .A(u5_mult_79_n1779), .ZN(u5_mult_79_n1778) );
  INV_X4 u5_mult_79_U920 ( .A(u5_mult_79_n1857), .ZN(u5_mult_79_n1779) );
  AND2_X2 u5_mult_79_U919 ( .A1(u5_mult_79_ab_23__23_), .A2(
        u5_mult_79_CARRYB_23__22_), .ZN(u5_mult_79_n245) );
  AND2_X4 u5_mult_79_U918 ( .A1(u5_mult_79_SUMB_23__20_), .A2(
        u5_mult_79_CARRYB_23__19_), .ZN(u5_mult_79_n244) );
  XOR2_X2 u5_mult_79_U917 ( .A(u5_mult_79_CARRYB_23__22_), .B(
        u5_mult_79_ab_23__23_), .Z(u5_mult_79_n243) );
  XOR2_X2 u5_mult_79_U916 ( .A(u5_mult_79_CARRYB_23__21_), .B(
        u5_mult_79_SUMB_23__22_), .Z(u5_mult_79_n242) );
  XOR2_X1 u5_mult_79_U915 ( .A(u5_mult_79_ab_6__22_), .B(u5_mult_79_ab_5__23_), 
        .Z(u5_mult_79_n241) );
  INV_X4 u5_mult_79_U914 ( .A(u5_mult_79_n478), .ZN(u5_mult_79_n442) );
  INV_X2 u5_mult_79_U913 ( .A(u5_mult_79_CARRYB_13__15_), .ZN(u5_mult_79_n478)
         );
  AND2_X2 u5_mult_79_U912 ( .A1(u5_mult_79_ab_0__10_), .A2(u5_mult_79_ab_1__9_), .ZN(u5_mult_79_n240) );
  AND2_X2 u5_mult_79_U911 ( .A1(u5_mult_79_ab_0__18_), .A2(
        u5_mult_79_ab_1__17_), .ZN(u5_mult_79_n239) );
  AND2_X2 u5_mult_79_U910 ( .A1(u5_mult_79_SUMB_23__5_), .A2(
        u5_mult_79_CARRYB_23__4_), .ZN(u5_mult_79_n238) );
  AND2_X4 u5_mult_79_U909 ( .A1(u5_mult_79_SUMB_23__15_), .A2(
        u5_mult_79_CARRYB_23__14_), .ZN(u5_mult_79_n237) );
  AND2_X4 u5_mult_79_U908 ( .A1(u5_mult_79_SUMB_23__17_), .A2(
        u5_mult_79_CARRYB_23__16_), .ZN(u5_mult_79_n236) );
  AND2_X4 u5_mult_79_U907 ( .A1(u5_mult_79_SUMB_23__19_), .A2(
        u5_mult_79_CARRYB_23__18_), .ZN(u5_mult_79_n235) );
  AND2_X4 u5_mult_79_U906 ( .A1(u5_mult_79_SUMB_23__7_), .A2(
        u5_mult_79_CARRYB_23__6_), .ZN(u5_mult_79_n232) );
  AND2_X4 u5_mult_79_U905 ( .A1(u5_mult_79_SUMB_23__16_), .A2(
        u5_mult_79_CARRYB_23__15_), .ZN(u5_mult_79_n231) );
  AND2_X4 u5_mult_79_U904 ( .A1(u5_mult_79_SUMB_23__9_), .A2(
        u5_mult_79_CARRYB_23__8_), .ZN(u5_mult_79_n230) );
  AND2_X2 u5_mult_79_U903 ( .A1(u5_mult_79_SUMB_23__12_), .A2(
        u5_mult_79_CARRYB_23__11_), .ZN(u5_mult_79_n229) );
  XNOR2_X2 u5_mult_79_U902 ( .A(u5_mult_79_n721), .B(u5_mult_79_SUMB_12__14_), 
        .ZN(u5_mult_79_n228) );
  INV_X1 u5_mult_79_U901 ( .A(u2_N124), .ZN(u5_mult_79_n1879) );
  INV_X4 u5_mult_79_U900 ( .A(u5_mult_79_n1830), .ZN(u5_mult_79_n1829) );
  INV_X4 u5_mult_79_U899 ( .A(u5_mult_79_n1879), .ZN(u5_mult_79_n1830) );
  INV_X16 u5_mult_79_U898 ( .A(u6_N1), .ZN(u5_mult_79_n1828) );
  INV_X16 u5_mult_79_U897 ( .A(u5_mult_79_n1824), .ZN(u5_mult_79_n1823) );
  INV_X4 u5_mult_79_U896 ( .A(u5_mult_79_n1876), .ZN(u5_mult_79_n1824) );
  NOR2_X1 u5_mult_79_U895 ( .A1(u5_mult_79_n1882), .A2(u5_mult_79_n1834), .ZN(
        u5_N0) );
  NOR2_X2 u5_mult_79_U894 ( .A1(u5_mult_79_n1835), .A2(u5_mult_79_n1722), .ZN(
        u5_mult_79_ab_2__0_) );
  NOR2_X2 u5_mult_79_U893 ( .A1(u5_mult_79_n1835), .A2(u5_mult_79_n1734), .ZN(
        u5_mult_79_ab_6__0_) );
  NOR2_X2 u5_mult_79_U892 ( .A1(u5_mult_79_n1835), .A2(u5_mult_79_n1746), .ZN(
        u5_mult_79_ab_10__0_) );
  NOR2_X2 u5_mult_79_U891 ( .A1(u5_mult_79_n1834), .A2(u5_mult_79_n1761), .ZN(
        u5_mult_79_ab_15__0_) );
  NOR2_X1 u5_mult_79_U890 ( .A1(u5_mult_79_n1834), .A2(u5_mult_79_n1770), .ZN(
        u5_mult_79_ab_18__0_) );
  NOR2_X1 u5_mult_79_U889 ( .A1(u5_mult_79_n1834), .A2(u5_mult_79_n1859), .ZN(
        u5_mult_79_ab_22__0_) );
  NOR2_X1 u5_mult_79_U888 ( .A1(u5_mult_79_n1828), .A2(u5_mult_79_n1722), .ZN(
        u5_mult_79_ab_2__1_) );
  NOR2_X1 u5_mult_79_U887 ( .A1(u5_mult_79_n1828), .A2(u5_mult_79_n1734), .ZN(
        u5_mult_79_ab_6__1_) );
  NOR2_X1 u5_mult_79_U886 ( .A1(u5_mult_79_n1828), .A2(u5_mult_79_n1746), .ZN(
        u5_mult_79_ab_10__1_) );
  INV_X4 u5_mult_79_U885 ( .A(u5_mult_79_ab_23__0_), .ZN(u5_mult_79_n254) );
  NOR2_X1 u5_mult_79_U884 ( .A1(u5_mult_79_n1832), .A2(u5_mult_79_n1829), .ZN(
        u5_mult_79_ab_23__23_) );
  NOR2_X1 u5_mult_79_U883 ( .A1(u5_mult_79_n1879), .A2(u5_mult_79_n1780), .ZN(
        u5_mult_79_ab_23__22_) );
  NOR2_X1 u5_mult_79_U882 ( .A1(u5_mult_79_n1832), .A2(u5_mult_79_n1859), .ZN(
        u5_mult_79_ab_22__23_) );
  NOR2_X1 u5_mult_79_U881 ( .A1(u5_mult_79_n1834), .A2(u5_mult_79_n1775), .ZN(
        u5_mult_79_ab_20__0_) );
  INV_X8 u5_mult_79_U880 ( .A(u5_mult_79_n1839), .ZN(u5_mult_79_n1727) );
  NOR2_X2 u5_mult_79_U879 ( .A1(u5_mult_79_n1825), .A2(u5_mult_79_n1722), .ZN(
        u5_mult_79_ab_2__2_) );
  INV_X8 u5_mult_79_U878 ( .A(u5_mult_79_n1840), .ZN(u5_mult_79_n1730) );
  INV_X8 u5_mult_79_U877 ( .A(u5_mult_79_n1841), .ZN(u5_mult_79_n1733) );
  INV_X8 u5_mult_79_U876 ( .A(u5_mult_79_n1843), .ZN(u5_mult_79_n1739) );
  INV_X8 u5_mult_79_U875 ( .A(u5_mult_79_n1844), .ZN(u5_mult_79_n1742) );
  INV_X4 u5_mult_79_U874 ( .A(u5_mult_79_n1847), .ZN(u5_mult_79_n1751) );
  NOR2_X2 u5_mult_79_U873 ( .A1(u5_mult_79_n1825), .A2(u5_mult_79_n1746), .ZN(
        u5_mult_79_ab_10__2_) );
  INV_X4 u5_mult_79_U872 ( .A(u5_mult_79_n1848), .ZN(u5_mult_79_n1754) );
  NOR2_X1 u5_mult_79_U871 ( .A1(u5_mult_79_n1823), .A2(u5_mult_79_n1746), .ZN(
        u5_mult_79_ab_10__3_) );
  NOR2_X2 u5_mult_79_U870 ( .A1(u5_mult_79_n1828), .A2(u5_mult_79_n1755), .ZN(
        u5_mult_79_ab_13__1_) );
  NOR2_X1 u5_mult_79_U869 ( .A1(u5_mult_79_n1828), .A2(u5_mult_79_n1770), .ZN(
        u5_mult_79_ab_18__1_) );
  NOR2_X1 u5_mult_79_U868 ( .A1(u5_mult_79_n1828), .A2(u5_mult_79_n1775), .ZN(
        u5_mult_79_ab_20__1_) );
  INV_X4 u5_mult_79_U867 ( .A(u5_mult_79_ab_23__2_), .ZN(u5_mult_79_n1330) );
  INV_X4 u5_mult_79_U866 ( .A(u5_mult_79_n1650), .ZN(u5_mult_79_n1718) );
  INV_X4 u5_mult_79_U865 ( .A(u5_mult_79_n1659), .ZN(u5_mult_79_CLA_SUM[34])
         );
  INV_X8 u5_mult_79_U864 ( .A(u5_mult_79_n1777), .ZN(u5_mult_79_n1775) );
  NOR2_X1 u5_mult_79_U863 ( .A1(u5_mult_79_n1823), .A2(u5_mult_79_n1722), .ZN(
        u5_mult_79_ab_2__3_) );
  INV_X4 u5_mult_79_U862 ( .A(u5_mult_79_n1849), .ZN(u5_mult_79_n1757) );
  INV_X4 u5_mult_79_U861 ( .A(u5_mult_79_n1850), .ZN(u5_mult_79_n1760) );
  INV_X8 u5_mult_79_U860 ( .A(u5_mult_79_n1852), .ZN(u5_mult_79_n1766) );
  INV_X4 u5_mult_79_U859 ( .A(u5_mult_79_n1853), .ZN(u5_mult_79_n1769) );
  INV_X4 u5_mult_79_U858 ( .A(u5_mult_79_ab_19__2_), .ZN(u5_mult_79_n810) );
  NOR2_X1 u5_mult_79_U857 ( .A1(u5_mult_79_n1826), .A2(u5_mult_79_n1775), .ZN(
        u5_mult_79_ab_20__2_) );
  INV_X4 u5_mult_79_U856 ( .A(u5_mult_79_ab_22__2_), .ZN(u5_mult_79_n1352) );
  NOR2_X1 u5_mult_79_U855 ( .A1(u5_mult_79_n1829), .A2(u5_mult_79_n1817), .ZN(
        u5_mult_79_ab_23__5_) );
  NOR2_X1 u5_mult_79_U854 ( .A1(u5_mult_79_n1829), .A2(u5_mult_79_n1814), .ZN(
        u5_mult_79_ab_23__6_) );
  NAND3_X2 u5_mult_79_U853 ( .A1(u5_mult_79_n962), .A2(u5_mult_79_n963), .A3(
        u5_mult_79_n964), .ZN(u5_mult_79_CARRYB_22__7_) );
  NOR2_X1 u5_mult_79_U852 ( .A1(u5_mult_79_n1829), .A2(u5_mult_79_n1811), .ZN(
        u5_mult_79_ab_23__7_) );
  NOR2_X1 u5_mult_79_U851 ( .A1(u5_mult_79_n1829), .A2(u5_mult_79_n1796), .ZN(
        u5_mult_79_ab_23__15_) );
  NOR2_X1 u5_mult_79_U850 ( .A1(u5_mult_79_n1829), .A2(u5_mult_79_n1793), .ZN(
        u5_mult_79_ab_23__16_) );
  NOR2_X1 u5_mult_79_U849 ( .A1(u5_mult_79_n1879), .A2(u5_mult_79_n1787), .ZN(
        u5_mult_79_ab_23__18_) );
  NOR2_X1 u5_mult_79_U848 ( .A1(u5_mult_79_n1829), .A2(u5_mult_79_n1790), .ZN(
        u5_mult_79_ab_23__17_) );
  NOR2_X1 u5_mult_79_U847 ( .A1(u5_mult_79_n1829), .A2(u5_mult_79_n1338), .ZN(
        u5_mult_79_ab_23__20_) );
  INV_X4 u5_mult_79_U846 ( .A(u5_mult_79_n1856), .ZN(u5_mult_79_n1777) );
  NOR2_X1 u5_mult_79_U845 ( .A1(u5_mult_79_n1823), .A2(u5_mult_79_n1859), .ZN(
        u5_mult_79_ab_22__3_) );
  NOR2_X1 u5_mult_79_U844 ( .A1(u5_mult_79_n1829), .A2(u5_mult_79_n1805), .ZN(
        u5_mult_79_ab_23__9_) );
  NOR2_X1 u5_mult_79_U843 ( .A1(u5_mult_79_n1829), .A2(u5_mult_79_n1802), .ZN(
        u5_mult_79_ab_23__10_) );
  NOR2_X1 u5_mult_79_U842 ( .A1(u5_mult_79_n1829), .A2(u5_mult_79_n1800), .ZN(
        u5_mult_79_ab_23__11_) );
  NOR2_X2 u5_mult_79_U841 ( .A1(u5_mult_79_n1817), .A2(u5_mult_79_n1722), .ZN(
        u5_mult_79_ab_2__5_) );
  NOR2_X2 u5_mult_79_U840 ( .A1(u5_mult_79_n1814), .A2(u5_mult_79_n1746), .ZN(
        u5_mult_79_ab_10__6_) );
  NOR2_X1 u5_mult_79_U839 ( .A1(u5_mult_79_n1821), .A2(u5_mult_79_n1778), .ZN(
        u5_mult_79_ab_21__4_) );
  NOR2_X2 u5_mult_79_U838 ( .A1(u5_mult_79_n1818), .A2(u5_mult_79_n1778), .ZN(
        u5_mult_79_ab_21__5_) );
  NOR2_X1 u5_mult_79_U837 ( .A1(u5_mult_79_n1820), .A2(u5_mult_79_n1859), .ZN(
        u5_mult_79_ab_22__4_) );
  NOR2_X1 u5_mult_79_U836 ( .A1(u5_mult_79_n1809), .A2(u5_mult_79_n1778), .ZN(
        u5_mult_79_ab_21__8_) );
  NOR2_X1 u5_mult_79_U835 ( .A1(u5_mult_79_n1806), .A2(u5_mult_79_n1778), .ZN(
        u5_mult_79_ab_21__9_) );
  INV_X4 u5_mult_79_U834 ( .A(u5_mult_79_ab_21__10_), .ZN(u5_mult_79_n622) );
  NOR2_X1 u5_mult_79_U833 ( .A1(u5_mult_79_n1802), .A2(u5_mult_79_n1859), .ZN(
        u5_mult_79_ab_22__10_) );
  NAND3_X2 u5_mult_79_U832 ( .A1(u5_mult_79_n1044), .A2(u5_mult_79_n1045), 
        .A3(u5_mult_79_n1046), .ZN(u5_mult_79_CARRYB_21__10_) );
  NOR2_X1 u5_mult_79_U831 ( .A1(u5_mult_79_n1800), .A2(u5_mult_79_n1859), .ZN(
        u5_mult_79_ab_22__11_) );
  NOR2_X1 u5_mult_79_U830 ( .A1(u5_mult_79_n1798), .A2(u5_mult_79_n1859), .ZN(
        u5_mult_79_ab_22__12_) );
  NOR2_X1 u5_mult_79_U829 ( .A1(u5_mult_79_n1796), .A2(u5_mult_79_n1778), .ZN(
        u5_mult_79_ab_21__15_) );
  NOR2_X1 u5_mult_79_U828 ( .A1(u5_mult_79_n1788), .A2(u5_mult_79_n1778), .ZN(
        u5_mult_79_ab_21__18_) );
  INV_X16 u5_mult_79_U827 ( .A(n2986), .ZN(u5_mult_79_n1798) );
  NOR2_X1 u5_mult_79_U826 ( .A1(u5_mult_79_n1781), .A2(u5_mult_79_n1773), .ZN(
        u5_mult_79_ab_19__22_) );
  NOR2_X1 u5_mult_79_U825 ( .A1(u5_mult_79_n1832), .A2(u5_mult_79_n1770), .ZN(
        u5_mult_79_ab_18__23_) );
  NOR2_X2 u5_mult_79_U824 ( .A1(u5_mult_79_n1814), .A2(u5_mult_79_n1722), .ZN(
        u5_mult_79_ab_2__6_) );
  NOR2_X1 u5_mult_79_U823 ( .A1(u5_mult_79_n1815), .A2(u5_mult_79_n1773), .ZN(
        u5_mult_79_ab_19__6_) );
  NOR2_X2 u5_mult_79_U822 ( .A1(u5_mult_79_n1815), .A2(u5_mult_79_n1778), .ZN(
        u5_mult_79_ab_21__6_) );
  NOR2_X1 u5_mult_79_U821 ( .A1(u5_mult_79_n1812), .A2(u5_mult_79_n1778), .ZN(
        u5_mult_79_ab_21__7_) );
  NOR2_X1 u5_mult_79_U820 ( .A1(u5_mult_79_n1809), .A2(u5_mult_79_n1773), .ZN(
        u5_mult_79_ab_19__8_) );
  NOR2_X1 u5_mult_79_U819 ( .A1(u5_mult_79_n1809), .A2(u5_mult_79_n1775), .ZN(
        u5_mult_79_ab_20__8_) );
  NOR2_X1 u5_mult_79_U818 ( .A1(u5_mult_79_n1806), .A2(u5_mult_79_n1775), .ZN(
        u5_mult_79_ab_20__9_) );
  NOR2_X2 u5_mult_79_U817 ( .A1(u5_mult_79_n1801), .A2(u5_mult_79_n1776), .ZN(
        u5_mult_79_ab_20__11_) );
  INV_X16 u5_mult_79_U816 ( .A(n2982), .ZN(u5_mult_79_n1801) );
  NOR2_X1 u5_mult_79_U815 ( .A1(u5_mult_79_n1796), .A2(u5_mult_79_n1776), .ZN(
        u5_mult_79_ab_20__15_) );
  INV_X2 u5_mult_79_U814 ( .A(u5_mult_79_ab_19__15_), .ZN(u5_mult_79_n575) );
  NOR2_X2 u5_mult_79_U813 ( .A1(u5_mult_79_n1811), .A2(u5_mult_79_n1722), .ZN(
        u5_mult_79_ab_2__7_) );
  NOR2_X2 u5_mult_79_U812 ( .A1(u5_mult_79_n1808), .A2(u5_mult_79_n1722), .ZN(
        u5_mult_79_ab_2__8_) );
  INV_X4 u5_mult_79_U811 ( .A(u5_mult_79_ab_19__7_), .ZN(u5_mult_79_n1424) );
  INV_X2 u5_mult_79_U810 ( .A(u5_mult_79_ab_18__17_), .ZN(u5_mult_79_n799) );
  NOR2_X2 u5_mult_79_U809 ( .A1(u5_mult_79_n1799), .A2(u5_mult_79_n1773), .ZN(
        u5_mult_79_ab_19__12_) );
  NOR2_X2 u5_mult_79_U808 ( .A1(u5_mult_79_n1805), .A2(u5_mult_79_n1722), .ZN(
        u5_mult_79_ab_2__9_) );
  NOR2_X2 u5_mult_79_U807 ( .A1(u5_mult_79_n1802), .A2(u5_mult_79_n1722), .ZN(
        u5_mult_79_ab_2__10_) );
  NOR2_X2 u5_mult_79_U806 ( .A1(u5_mult_79_n1800), .A2(u5_mult_79_n1723), .ZN(
        u5_mult_79_ab_2__11_) );
  NAND2_X2 u5_mult_79_U805 ( .A1(u5_mult_79_CARRYB_14__7_), .A2(
        u5_mult_79_ab_15__7_), .ZN(u5_mult_79_n1287) );
  INV_X4 u5_mult_79_U804 ( .A(u5_mult_79_ab_15__9_), .ZN(u5_mult_79_n627) );
  INV_X4 u5_mult_79_U803 ( .A(u5_mult_79_ab_15__12_), .ZN(u5_mult_79_n1239) );
  NAND2_X1 u5_mult_79_U802 ( .A1(u5_mult_79_ab_15__12_), .A2(
        u5_mult_79_SUMB_14__13_), .ZN(u5_mult_79_n1363) );
  INV_X4 u5_mult_79_U801 ( .A(u5_mult_79_n429), .ZN(u5_mult_79_n430) );
  NAND3_X2 u5_mult_79_U800 ( .A1(u5_mult_79_n502), .A2(u5_mult_79_n503), .A3(
        u5_mult_79_n504), .ZN(u5_mult_79_CARRYB_10__9_) );
  NOR2_X2 u5_mult_79_U799 ( .A1(u5_mult_79_n1867), .A2(u5_mult_79_n1762), .ZN(
        u5_mult_79_ab_15__14_) );
  NOR2_X2 u5_mult_79_U798 ( .A1(u5_mult_79_n1868), .A2(u5_mult_79_n1723), .ZN(
        u5_mult_79_ab_2__13_) );
  NOR2_X2 u5_mult_79_U797 ( .A1(u5_mult_79_n1802), .A2(u5_mult_79_n1746), .ZN(
        u5_mult_79_ab_10__10_) );
  NOR2_X2 u5_mult_79_U796 ( .A1(u5_mult_79_n1790), .A2(u5_mult_79_n1747), .ZN(
        u5_mult_79_ab_10__17_) );
  NOR2_X2 u5_mult_79_U795 ( .A1(u5_mult_79_n1793), .A2(u5_mult_79_n1747), .ZN(
        u5_mult_79_ab_10__16_) );
  NOR2_X2 u5_mult_79_U794 ( .A1(u5_mult_79_n1867), .A2(u5_mult_79_n1735), .ZN(
        u5_mult_79_ab_6__14_) );
  NOR2_X2 u5_mult_79_U793 ( .A1(u5_mult_79_n1790), .A2(u5_mult_79_n1723), .ZN(
        u5_mult_79_ab_2__17_) );
  NOR2_X2 u5_mult_79_U792 ( .A1(u5_mult_79_n1338), .A2(u5_mult_79_n1723), .ZN(
        u5_mult_79_ab_2__20_) );
  NOR2_X2 u5_mult_79_U791 ( .A1(u5_mult_79_n1835), .A2(u5_mult_79_n1725), .ZN(
        u5_mult_79_ab_3__0_) );
  NOR2_X2 u5_mult_79_U790 ( .A1(u5_mult_79_n1835), .A2(u5_mult_79_n1737), .ZN(
        u5_mult_79_ab_7__0_) );
  NOR2_X2 u5_mult_79_U789 ( .A1(u5_mult_79_n1835), .A2(u5_mult_79_n1749), .ZN(
        u5_mult_79_ab_11__0_) );
  INV_X4 u5_mult_79_U788 ( .A(u5_mult_79_ab_17__0_), .ZN(u5_mult_79_n247) );
  NOR2_X2 u5_mult_79_U787 ( .A1(u5_mult_79_n1882), .A2(u5_mult_79_n1828), .ZN(
        u5_mult_79_ab_0__1_) );
  NOR2_X1 u5_mult_79_U786 ( .A1(u5_mult_79_n1828), .A2(u5_mult_79_n1725), .ZN(
        u5_mult_79_ab_3__1_) );
  NOR2_X1 u5_mult_79_U785 ( .A1(u5_mult_79_n1828), .A2(u5_mult_79_n1737), .ZN(
        u5_mult_79_ab_7__1_) );
  NOR2_X1 u5_mult_79_U784 ( .A1(u5_mult_79_n1828), .A2(u5_mult_79_n1749), .ZN(
        u5_mult_79_ab_11__1_) );
  NOR2_X1 u5_mult_79_U783 ( .A1(u5_mult_79_n1834), .A2(u5_mult_79_n1778), .ZN(
        u5_mult_79_ab_21__0_) );
  NOR2_X2 u5_mult_79_U782 ( .A1(u5_mult_79_n1878), .A2(u5_mult_79_n1719), .ZN(
        u5_mult_79_ab_1__1_) );
  NOR2_X2 u5_mult_79_U781 ( .A1(u5_mult_79_n1825), .A2(u5_mult_79_n1725), .ZN(
        u5_mult_79_ab_3__2_) );
  INV_X8 u5_mult_79_U780 ( .A(u5_mult_79_n1842), .ZN(u5_mult_79_n1736) );
  INV_X8 u5_mult_79_U779 ( .A(u5_mult_79_n1846), .ZN(u5_mult_79_n1748) );
  INV_X16 u5_mult_79_U778 ( .A(u5_mult_79_n1760), .ZN(u5_mult_79_n1758) );
  NOR2_X2 u5_mult_79_U777 ( .A1(u5_mult_79_n1826), .A2(u5_mult_79_n1755), .ZN(
        u5_mult_79_ab_13__2_) );
  NOR2_X1 u5_mult_79_U776 ( .A1(u5_mult_79_n1823), .A2(u5_mult_79_n1755), .ZN(
        u5_mult_79_ab_13__3_) );
  INV_X4 u5_mult_79_U775 ( .A(u5_mult_79_n1854), .ZN(u5_mult_79_n1772) );
  NOR2_X1 u5_mult_79_U774 ( .A1(u5_mult_79_n1828), .A2(u5_mult_79_n1778), .ZN(
        u5_mult_79_ab_21__1_) );
  INV_X4 u5_mult_79_U773 ( .A(u5_mult_79_n1666), .ZN(u5_mult_79_CLA_SUM[39])
         );
  NOR2_X1 u5_mult_79_U772 ( .A1(u5_mult_79_n1859), .A2(u5_mult_79_n1780), .ZN(
        u5_mult_79_ab_22__22_) );
  NOR2_X1 u5_mult_79_U771 ( .A1(u5_mult_79_n1832), .A2(u5_mult_79_n1778), .ZN(
        u5_mult_79_ab_21__23_) );
  NOR2_X2 u5_mult_79_U770 ( .A1(u5_mult_79_n1882), .A2(u5_mult_79_n1876), .ZN(
        u5_mult_79_ab_0__3_) );
  NOR2_X2 u5_mult_79_U769 ( .A1(u5_mult_79_n1820), .A2(u5_mult_79_n1743), .ZN(
        u5_mult_79_ab_9__4_) );
  NOR2_X1 u5_mult_79_U768 ( .A1(u5_mult_79_n1829), .A2(u5_mult_79_n1825), .ZN(
        u5_mult_79_ab_23__2_) );
  NOR2_X1 u5_mult_79_U767 ( .A1(u5_mult_79_n1829), .A2(u5_mult_79_n1823), .ZN(
        u5_mult_79_ab_23__3_) );
  NOR2_X1 u5_mult_79_U766 ( .A1(u5_mult_79_n1829), .A2(u5_mult_79_n1820), .ZN(
        u5_mult_79_ab_23__4_) );
  NOR2_X1 u5_mult_79_U765 ( .A1(u5_mult_79_n1829), .A2(u5_mult_79_n1868), .ZN(
        u5_mult_79_ab_23__13_) );
  NOR2_X2 u5_mult_79_U764 ( .A1(u5_mult_79_n1876), .A2(u5_mult_79_n1720), .ZN(
        u5_mult_79_ab_1__3_) );
  NOR2_X2 u5_mult_79_U763 ( .A1(u5_mult_79_n1820), .A2(u5_mult_79_n1722), .ZN(
        u5_mult_79_ab_2__4_) );
  NOR2_X1 u5_mult_79_U762 ( .A1(u5_mult_79_n1825), .A2(u5_mult_79_n1859), .ZN(
        u5_mult_79_ab_22__2_) );
  INV_X4 u5_mult_79_U761 ( .A(u5_mult_79_ab_22__11_), .ZN(u5_mult_79_n469) );
  NAND3_X2 u5_mult_79_U760 ( .A1(u5_mult_79_n1307), .A2(u5_mult_79_n1308), 
        .A3(u5_mult_79_n1306), .ZN(u5_mult_79_CARRYB_22__11_) );
  CLKBUF_X3 u5_mult_79_U759 ( .A(u5_mult_79_SUMB_21__13_), .Z(u5_mult_79_n499)
         );
  NOR2_X1 u5_mult_79_U758 ( .A1(u5_mult_79_n1790), .A2(u5_mult_79_n1859), .ZN(
        u5_mult_79_ab_22__17_) );
  NOR2_X1 u5_mult_79_U757 ( .A1(u5_mult_79_n1787), .A2(u5_mult_79_n1859), .ZN(
        u5_mult_79_ab_22__18_) );
  NOR2_X1 u5_mult_79_U756 ( .A1(u5_mult_79_n1338), .A2(u5_mult_79_n1859), .ZN(
        u5_mult_79_ab_22__20_) );
  NOR2_X2 u5_mult_79_U755 ( .A1(u5_mult_79_n1817), .A2(u5_mult_79_n1725), .ZN(
        u5_mult_79_ab_3__5_) );
  NOR2_X2 u5_mult_79_U754 ( .A1(u5_mult_79_n1814), .A2(u5_mult_79_n1728), .ZN(
        u5_mult_79_ab_4__6_) );
  NAND3_X2 u5_mult_79_U753 ( .A1(u5_mult_79_n921), .A2(u5_mult_79_n922), .A3(
        u5_mult_79_n923), .ZN(u5_mult_79_CARRYB_8__6_) );
  NOR2_X2 u5_mult_79_U752 ( .A1(u5_mult_79_n1814), .A2(u5_mult_79_n1743), .ZN(
        u5_mult_79_ab_9__6_) );
  INV_X4 u5_mult_79_U751 ( .A(u5_mult_79_ab_21__7_), .ZN(u5_mult_79_n543) );
  NOR2_X1 u5_mult_79_U750 ( .A1(u5_mult_79_n1811), .A2(u5_mult_79_n1859), .ZN(
        u5_mult_79_ab_22__7_) );
  INV_X16 u5_mult_79_U749 ( .A(u5_mult_79_n1777), .ZN(u5_mult_79_n1776) );
  INV_X2 u5_mult_79_U748 ( .A(u5_mult_79_ab_9__7_), .ZN(u5_mult_79_n265) );
  NAND2_X2 u5_mult_79_U747 ( .A1(u5_mult_79_n747), .A2(u5_mult_79_n748), .ZN(
        u5_mult_79_n750) );
  NOR2_X1 u5_mult_79_U746 ( .A1(u5_mult_79_n1815), .A2(u5_mult_79_n1775), .ZN(
        u5_mult_79_ab_20__6_) );
  INV_X8 u5_mult_79_U745 ( .A(u5_mult_79_n1871), .ZN(u5_mult_79_n1810) );
  INV_X4 u5_mult_79_U744 ( .A(u5_mult_79_ab_20__11_), .ZN(u5_mult_79_n1149) );
  INV_X8 u5_mult_79_U743 ( .A(u5_mult_79_n1869), .ZN(u5_mult_79_n1804) );
  INV_X4 u5_mult_79_U742 ( .A(u5_mult_79_ab_17__17_), .ZN(u5_mult_79_n369) );
  NAND3_X2 u5_mult_79_U741 ( .A1(u5_mult_79_n1004), .A2(u5_mult_79_n1005), 
        .A3(u5_mult_79_n1006), .ZN(u5_mult_79_CARRYB_17__16_) );
  NOR2_X1 u5_mult_79_U740 ( .A1(u5_mult_79_n1832), .A2(u5_mult_79_n1764), .ZN(
        u5_mult_79_ab_16__23_) );
  NOR2_X2 u5_mult_79_U739 ( .A1(u5_mult_79_n1781), .A2(u5_mult_79_n1768), .ZN(
        u5_mult_79_ab_17__22_) );
  INV_X4 u5_mult_79_U738 ( .A(u5_mult_79_ab_16__11_), .ZN(u5_mult_79_n1316) );
  NAND2_X2 u5_mult_79_U737 ( .A1(u5_mult_79_n1239), .A2(u5_mult_79_n1240), 
        .ZN(u5_mult_79_n1242) );
  NOR2_X2 u5_mult_79_U736 ( .A1(u5_mult_79_n1785), .A2(u5_mult_79_n1765), .ZN(
        u5_mult_79_ab_16__19_) );
  NOR2_X1 u5_mult_79_U735 ( .A1(u5_mult_79_n1338), .A2(u5_mult_79_n1765), .ZN(
        u5_mult_79_ab_16__20_) );
  NOR2_X1 u5_mult_79_U734 ( .A1(u5_mult_79_n1783), .A2(u5_mult_79_n1768), .ZN(
        u5_mult_79_ab_17__21_) );
  NOR2_X2 u5_mult_79_U733 ( .A1(u5_mult_79_n1799), .A2(u5_mult_79_n1765), .ZN(
        u5_mult_79_ab_16__12_) );
  NOR2_X1 u5_mult_79_U732 ( .A1(u5_mult_79_n1798), .A2(u5_mult_79_n1729), .ZN(
        u5_mult_79_ab_4__12_) );
  INV_X4 u5_mult_79_U731 ( .A(u5_mult_79_ab_7__11_), .ZN(u5_mult_79_n1033) );
  NAND2_X2 u5_mult_79_U730 ( .A1(u5_mult_79_ab_14__9_), .A2(
        u5_mult_79_CARRYB_13__9_), .ZN(u5_mult_79_n1329) );
  NOR2_X2 u5_mult_79_U729 ( .A1(u5_mult_79_n1791), .A2(u5_mult_79_n1756), .ZN(
        u5_mult_79_ab_13__17_) );
  INV_X4 u5_mult_79_U728 ( .A(u5_mult_79_ab_5__13_), .ZN(u5_mult_79_n806) );
  INV_X16 u5_mult_79_U727 ( .A(u5_mult_79_n1751), .ZN(u5_mult_79_n1750) );
  INV_X16 u5_mult_79_U726 ( .A(u5_mult_79_n1760), .ZN(u5_mult_79_n1759) );
  INV_X2 u5_mult_79_U725 ( .A(u5_mult_79_ab_13__11_), .ZN(u5_mult_79_n632) );
  NOR2_X2 u5_mult_79_U724 ( .A1(u5_mult_79_n1799), .A2(u5_mult_79_n1756), .ZN(
        u5_mult_79_ab_13__12_) );
  NAND2_X2 u5_mult_79_U723 ( .A1(u5_mult_79_SUMB_12__15_), .A2(
        u5_mult_79_ab_13__14_), .ZN(u5_mult_79_n898) );
  NOR2_X2 u5_mult_79_U722 ( .A1(u5_mult_79_n1800), .A2(u5_mult_79_n1744), .ZN(
        u5_mult_79_ab_9__11_) );
  NOR2_X1 u5_mult_79_U721 ( .A1(u5_mult_79_n1798), .A2(u5_mult_79_n1744), .ZN(
        u5_mult_79_ab_9__12_) );
  INV_X4 u5_mult_79_U720 ( .A(u5_mult_79_n489), .ZN(u5_mult_79_n490) );
  NOR2_X2 u5_mult_79_U719 ( .A1(u5_mult_79_n1799), .A2(u5_mult_79_n1753), .ZN(
        u5_mult_79_ab_12__12_) );
  NOR2_X1 u5_mult_79_U718 ( .A1(u5_mult_79_n1796), .A2(u5_mult_79_n1756), .ZN(
        u5_mult_79_ab_13__15_) );
  NOR2_X2 u5_mult_79_U717 ( .A1(u5_mult_79_n1780), .A2(u5_mult_79_n1744), .ZN(
        u5_mult_79_ab_9__22_) );
  NAND3_X2 u5_mult_79_U716 ( .A1(u5_mult_79_n1370), .A2(u5_mult_79_n1371), 
        .A3(u5_mult_79_n1372), .ZN(u5_mult_79_CARRYB_8__18_) );
  NOR2_X2 u5_mult_79_U715 ( .A1(u5_mult_79_n1787), .A2(u5_mult_79_n1744), .ZN(
        u5_mult_79_ab_9__18_) );
  NOR2_X1 u5_mult_79_U714 ( .A1(u5_mult_79_n1338), .A2(u5_mult_79_n1741), .ZN(
        u5_mult_79_ab_8__20_) );
  INV_X4 u5_mult_79_U713 ( .A(u5_mult_79_n283), .ZN(u5_mult_79_n284) );
  INV_X4 u5_mult_79_U712 ( .A(u5_mult_79_ab_3__20_), .ZN(u5_mult_79_n1353) );
  NOR2_X2 u5_mult_79_U711 ( .A1(u5_mult_79_n1835), .A2(u5_mult_79_n1728), .ZN(
        u5_mult_79_ab_4__0_) );
  NOR2_X2 u5_mult_79_U710 ( .A1(u5_mult_79_n1835), .A2(u5_mult_79_n1740), .ZN(
        u5_mult_79_ab_8__0_) );
  NOR2_X2 u5_mult_79_U709 ( .A1(u5_mult_79_n1834), .A2(u5_mult_79_n1752), .ZN(
        u5_mult_79_ab_12__0_) );
  NOR2_X1 u5_mult_79_U708 ( .A1(u5_mult_79_n1828), .A2(u5_mult_79_n1728), .ZN(
        u5_mult_79_ab_4__1_) );
  NOR2_X1 u5_mult_79_U707 ( .A1(u5_mult_79_n1828), .A2(u5_mult_79_n1740), .ZN(
        u5_mult_79_ab_8__1_) );
  NOR2_X1 u5_mult_79_U706 ( .A1(u5_mult_79_n1828), .A2(u5_mult_79_n1752), .ZN(
        u5_mult_79_ab_12__1_) );
  NOR2_X1 u5_mult_79_U705 ( .A1(u5_mult_79_n1828), .A2(u5_mult_79_n1761), .ZN(
        u5_mult_79_ab_15__1_) );
  NOR2_X1 u5_mult_79_U704 ( .A1(u5_mult_79_n1834), .A2(u5_mult_79_n1767), .ZN(
        u5_mult_79_ab_17__0_) );
  INV_X8 u5_mult_79_U703 ( .A(n3000), .ZN(u5_mult_79_n1838) );
  INV_X16 u5_mult_79_U702 ( .A(u5_mult_79_n1838), .ZN(u5_mult_79_n1724) );
  NOR2_X2 u5_mult_79_U701 ( .A1(u5_mult_79_n1826), .A2(u5_mult_79_n1761), .ZN(
        u5_mult_79_ab_15__2_) );
  NOR2_X1 u5_mult_79_U700 ( .A1(u5_mult_79_n1828), .A2(u5_mult_79_n1773), .ZN(
        u5_mult_79_ab_19__1_) );
  NOR2_X1 u5_mult_79_U699 ( .A1(u5_mult_79_n1823), .A2(u5_mult_79_n1725), .ZN(
        u5_mult_79_ab_3__3_) );
  NOR2_X1 u5_mult_79_U698 ( .A1(u5_mult_79_n1823), .A2(u5_mult_79_n1761), .ZN(
        u5_mult_79_ab_15__3_) );
  NOR2_X1 u5_mult_79_U697 ( .A1(u5_mult_79_n1780), .A2(u5_mult_79_n1778), .ZN(
        u5_mult_79_ab_21__22_) );
  NOR2_X1 u5_mult_79_U696 ( .A1(u5_mult_79_n1832), .A2(u5_mult_79_n1775), .ZN(
        u5_mult_79_ab_20__23_) );
  NOR2_X2 u5_mult_79_U695 ( .A1(u5_mult_79_n1820), .A2(u5_mult_79_n1725), .ZN(
        u5_mult_79_ab_3__4_) );
  NOR2_X2 u5_mult_79_U694 ( .A1(u5_mult_79_n1821), .A2(u5_mult_79_n1770), .ZN(
        u5_mult_79_ab_18__4_) );
  NOR2_X1 u5_mult_79_U693 ( .A1(u5_mult_79_n1796), .A2(u5_mult_79_n1859), .ZN(
        u5_mult_79_ab_22__15_) );
  NAND3_X2 u5_mult_79_U692 ( .A1(u5_mult_79_n600), .A2(u5_mult_79_n601), .A3(
        u5_mult_79_n602), .ZN(u5_mult_79_CARRYB_21__14_) );
  NOR2_X1 u5_mult_79_U691 ( .A1(u5_mult_79_n1868), .A2(u5_mult_79_n1859), .ZN(
        u5_mult_79_ab_22__13_) );
  NOR2_X1 u5_mult_79_U690 ( .A1(u5_mult_79_n1793), .A2(u5_mult_79_n1859), .ZN(
        u5_mult_79_ab_22__16_) );
  NOR2_X2 u5_mult_79_U689 ( .A1(u5_mult_79_n1817), .A2(u5_mult_79_n1728), .ZN(
        u5_mult_79_ab_4__5_) );
  NAND2_X2 u5_mult_79_U688 ( .A1(u5_mult_79_ab_11__5_), .A2(u5_mult_79_n404), 
        .ZN(u5_mult_79_n1113) );
  NOR2_X1 u5_mult_79_U687 ( .A1(u5_mult_79_n1818), .A2(u5_mult_79_n1775), .ZN(
        u5_mult_79_ab_20__5_) );
  INV_X4 u5_mult_79_U686 ( .A(u5_mult_79_ab_21__6_), .ZN(u5_mult_79_n670) );
  NOR2_X1 u5_mult_79_U685 ( .A1(u5_mult_79_n1817), .A2(u5_mult_79_n1859), .ZN(
        u5_mult_79_ab_22__5_) );
  INV_X8 u5_mult_79_U684 ( .A(u5_mult_79_n1872), .ZN(u5_mult_79_n1813) );
  NOR2_X1 u5_mult_79_U683 ( .A1(u5_mult_79_n1801), .A2(u5_mult_79_n1778), .ZN(
        u5_mult_79_ab_21__11_) );
  NOR2_X1 u5_mult_79_U682 ( .A1(u5_mult_79_n1799), .A2(u5_mult_79_n1778), .ZN(
        u5_mult_79_ab_21__12_) );
  NOR2_X1 u5_mult_79_U681 ( .A1(u5_mult_79_n1338), .A2(u5_mult_79_n1778), .ZN(
        u5_mult_79_ab_21__20_) );
  NOR2_X1 u5_mult_79_U680 ( .A1(u5_mult_79_n1785), .A2(u5_mult_79_n1778), .ZN(
        u5_mult_79_ab_21__19_) );
  NOR2_X1 u5_mult_79_U679 ( .A1(u5_mult_79_n1783), .A2(u5_mult_79_n1778), .ZN(
        u5_mult_79_ab_21__21_) );
  INV_X2 u5_mult_79_U678 ( .A(u5_mult_79_ab_5__6_), .ZN(u5_mult_79_n668) );
  NOR2_X2 u5_mult_79_U677 ( .A1(u5_mult_79_n1808), .A2(u5_mult_79_n1731), .ZN(
        u5_mult_79_ab_5__8_) );
  INV_X16 u5_mult_79_U676 ( .A(u5_mult_79_n1772), .ZN(u5_mult_79_n1771) );
  NOR2_X2 u5_mult_79_U675 ( .A1(u5_mult_79_n1805), .A2(u5_mult_79_n1731), .ZN(
        u5_mult_79_ab_5__9_) );
  INV_X4 u5_mult_79_U674 ( .A(u5_mult_79_ab_6__10_), .ZN(u5_mult_79_n270) );
  NOR2_X2 u5_mult_79_U673 ( .A1(u5_mult_79_n1788), .A2(u5_mult_79_n1765), .ZN(
        u5_mult_79_ab_16__18_) );
  INV_X16 u5_mult_79_U672 ( .A(u5_mult_79_n1769), .ZN(u5_mult_79_n1768) );
  INV_X4 u5_mult_79_U671 ( .A(u5_mult_79_ab_6__11_), .ZN(u5_mult_79_n848) );
  NOR2_X2 u5_mult_79_U670 ( .A1(u5_mult_79_n1803), .A2(u5_mult_79_n1761), .ZN(
        u5_mult_79_ab_15__10_) );
  NOR2_X2 u5_mult_79_U669 ( .A1(u5_mult_79_n1791), .A2(u5_mult_79_n1762), .ZN(
        u5_mult_79_ab_15__17_) );
  NOR2_X2 u5_mult_79_U668 ( .A1(u5_mult_79_n1338), .A2(u5_mult_79_n1762), .ZN(
        u5_mult_79_ab_15__20_) );
  NOR2_X1 u5_mult_79_U667 ( .A1(u5_mult_79_n1783), .A2(u5_mult_79_n1762), .ZN(
        u5_mult_79_ab_15__21_) );
  NOR2_X2 u5_mult_79_U666 ( .A1(u5_mult_79_n1781), .A2(u5_mult_79_n1762), .ZN(
        u5_mult_79_ab_15__22_) );
  NOR2_X1 u5_mult_79_U665 ( .A1(u5_mult_79_n1832), .A2(u5_mult_79_n1758), .ZN(
        u5_mult_79_ab_14__23_) );
  INV_X4 u5_mult_79_U664 ( .A(u5_mult_79_ab_6__12_), .ZN(u5_mult_79_n1014) );
  INV_X4 u5_mult_79_U663 ( .A(u5_mult_79_n228), .ZN(u5_mult_79_n1426) );
  NOR2_X2 u5_mult_79_U662 ( .A1(u5_mult_79_n1868), .A2(u5_mult_79_n1762), .ZN(
        u5_mult_79_ab_15__13_) );
  INV_X4 u5_mult_79_U661 ( .A(u5_mult_79_ab_14__16_), .ZN(u5_mult_79_n798) );
  NAND3_X2 u5_mult_79_U660 ( .A1(u5_mult_79_n1436), .A2(u5_mult_79_n1437), 
        .A3(u5_mult_79_n1438), .ZN(u5_mult_79_CARRYB_14__16_) );
  INV_X2 u5_mult_79_U659 ( .A(u5_mult_79_ab_11__15_), .ZN(u5_mult_79_n1032) );
  INV_X16 u5_mult_79_U658 ( .A(u5_mult_79_n1754), .ZN(u5_mult_79_n1753) );
  NOR2_X2 u5_mult_79_U657 ( .A1(u5_mult_79_n1868), .A2(u5_mult_79_n1735), .ZN(
        u5_mult_79_ab_6__13_) );
  NOR2_X2 u5_mult_79_U656 ( .A1(u5_mult_79_n1338), .A2(u5_mult_79_n1744), .ZN(
        u5_mult_79_ab_9__20_) );
  INV_X4 u5_mult_79_U655 ( .A(u5_mult_79_ab_5__16_), .ZN(u5_mult_79_n968) );
  NOR2_X1 u5_mult_79_U654 ( .A1(u5_mult_79_n1796), .A2(u5_mult_79_n1732), .ZN(
        u5_mult_79_ab_5__15_) );
  NOR2_X2 u5_mult_79_U653 ( .A1(u5_mult_79_n1835), .A2(u5_mult_79_n1731), .ZN(
        u5_mult_79_ab_5__0_) );
  NOR2_X2 u5_mult_79_U652 ( .A1(u5_mult_79_n1835), .A2(u5_mult_79_n1743), .ZN(
        u5_mult_79_ab_9__0_) );
  NOR2_X1 u5_mult_79_U651 ( .A1(u5_mult_79_n1828), .A2(u5_mult_79_n1731), .ZN(
        u5_mult_79_ab_5__1_) );
  NOR2_X1 u5_mult_79_U650 ( .A1(u5_mult_79_n1828), .A2(u5_mult_79_n1743), .ZN(
        u5_mult_79_ab_9__1_) );
  NOR2_X2 u5_mult_79_U649 ( .A1(u5_mult_79_n1825), .A2(u5_mult_79_n1743), .ZN(
        u5_mult_79_ab_9__2_) );
  NOR2_X2 u5_mult_79_U648 ( .A1(u5_mult_79_n1826), .A2(u5_mult_79_n1764), .ZN(
        u5_mult_79_ab_16__2_) );
  NOR2_X1 u5_mult_79_U647 ( .A1(u5_mult_79_n1823), .A2(u5_mult_79_n1728), .ZN(
        u5_mult_79_ab_4__3_) );
  NOR2_X1 u5_mult_79_U646 ( .A1(u5_mult_79_n1823), .A2(u5_mult_79_n1743), .ZN(
        u5_mult_79_ab_9__3_) );
  NOR2_X2 u5_mult_79_U645 ( .A1(u5_mult_79_n1821), .A2(u5_mult_79_n1752), .ZN(
        u5_mult_79_ab_12__4_) );
  NOR2_X1 u5_mult_79_U644 ( .A1(u5_mult_79_n1823), .A2(u5_mult_79_n1773), .ZN(
        u5_mult_79_ab_19__3_) );
  INV_X8 u5_mult_79_U643 ( .A(n3003), .ZN(u5_mult_79_n1858) );
  INV_X16 u5_mult_79_U642 ( .A(u5_mult_79_n1858), .ZN(u5_mult_79_n1782) );
  NOR2_X2 u5_mult_79_U641 ( .A1(u5_mult_79_n1820), .A2(u5_mult_79_n1728), .ZN(
        u5_mult_79_ab_4__4_) );
  NOR2_X2 u5_mult_79_U640 ( .A1(u5_mult_79_n1817), .A2(u5_mult_79_n1740), .ZN(
        u5_mult_79_ab_8__5_) );
  INV_X4 u5_mult_79_U639 ( .A(u5_mult_79_ab_21__5_), .ZN(u5_mult_79_n522) );
  NOR2_X1 u5_mult_79_U638 ( .A1(u5_mult_79_n1791), .A2(u5_mult_79_n1778), .ZN(
        u5_mult_79_ab_21__17_) );
  NOR2_X1 u5_mult_79_U637 ( .A1(u5_mult_79_n1868), .A2(u5_mult_79_n1778), .ZN(
        u5_mult_79_ab_21__13_) );
  NOR2_X1 u5_mult_79_U636 ( .A1(u5_mult_79_n1794), .A2(u5_mult_79_n1778), .ZN(
        u5_mult_79_ab_21__16_) );
  NOR2_X2 u5_mult_79_U635 ( .A1(u5_mult_79_n1814), .A2(u5_mult_79_n1725), .ZN(
        u5_mult_79_ab_3__6_) );
  NOR2_X2 u5_mult_79_U634 ( .A1(u5_mult_79_n1811), .A2(u5_mult_79_n1725), .ZN(
        u5_mult_79_ab_3__7_) );
  INV_X4 u5_mult_79_U633 ( .A(u5_mult_79_ab_7__8_), .ZN(u5_mult_79_n777) );
  NOR2_X1 u5_mult_79_U632 ( .A1(u5_mult_79_n1799), .A2(u5_mult_79_n1776), .ZN(
        u5_mult_79_ab_20__12_) );
  NOR2_X1 u5_mult_79_U631 ( .A1(u5_mult_79_n1338), .A2(u5_mult_79_n1773), .ZN(
        u5_mult_79_ab_19__20_) );
  INV_X4 u5_mult_79_U630 ( .A(u5_mult_79_ab_7__7_), .ZN(u5_mult_79_n811) );
  NOR2_X2 u5_mult_79_U629 ( .A1(u5_mult_79_n1805), .A2(u5_mult_79_n1740), .ZN(
        u5_mult_79_ab_8__9_) );
  NAND3_X2 u5_mult_79_U628 ( .A1(u5_mult_79_n705), .A2(u5_mult_79_n706), .A3(
        u5_mult_79_n707), .ZN(u5_mult_79_CARRYB_8__8_) );
  NOR2_X2 u5_mult_79_U627 ( .A1(u5_mult_79_n1812), .A2(u5_mult_79_n1755), .ZN(
        u5_mult_79_ab_13__7_) );
  NOR2_X2 u5_mult_79_U626 ( .A1(u5_mult_79_n1802), .A2(u5_mult_79_n1740), .ZN(
        u5_mult_79_ab_8__10_) );
  INV_X4 u5_mult_79_U625 ( .A(u5_mult_79_ab_14__20_), .ZN(u5_mult_79_n434) );
  NOR2_X1 u5_mult_79_U624 ( .A1(u5_mult_79_n1801), .A2(u5_mult_79_n1759), .ZN(
        u5_mult_79_ab_14__11_) );
  NOR2_X1 u5_mult_79_U623 ( .A1(u5_mult_79_n1803), .A2(u5_mult_79_n1758), .ZN(
        u5_mult_79_ab_14__10_) );
  NOR2_X2 u5_mult_79_U622 ( .A1(u5_mult_79_n1788), .A2(u5_mult_79_n1759), .ZN(
        u5_mult_79_ab_14__18_) );
  NOR2_X2 u5_mult_79_U621 ( .A1(u5_mult_79_n1800), .A2(u5_mult_79_n1741), .ZN(
        u5_mult_79_ab_8__11_) );
  NAND3_X2 u5_mult_79_U620 ( .A1(u5_mult_79_n722), .A2(u5_mult_79_n723), .A3(
        u5_mult_79_n724), .ZN(u5_mult_79_CARRYB_12__14_) );
  INV_X4 u5_mult_79_U619 ( .A(u5_mult_79_ab_11__18_), .ZN(u5_mult_79_n362) );
  INV_X4 u5_mult_79_U618 ( .A(u5_mult_79_ab_12__17_), .ZN(u5_mult_79_n752) );
  INV_X2 u5_mult_79_U617 ( .A(u5_mult_79_ab_7__21_), .ZN(u5_mult_79_n800) );
  INV_X4 u5_mult_79_U616 ( .A(u5_mult_79_n1881), .ZN(u5_mult_79_n1836) );
  NOR2_X2 u5_mult_79_U615 ( .A1(u5_mult_79_n1825), .A2(u5_mult_79_n1728), .ZN(
        u5_mult_79_ab_4__2_) );
  NOR2_X1 u5_mult_79_U614 ( .A1(u5_mult_79_n1823), .A2(u5_mult_79_n1731), .ZN(
        u5_mult_79_ab_5__3_) );
  NOR2_X1 u5_mult_79_U613 ( .A1(u5_mult_79_n1823), .A2(u5_mult_79_n1752), .ZN(
        u5_mult_79_ab_12__3_) );
  NOR2_X1 u5_mult_79_U612 ( .A1(u5_mult_79_n1826), .A2(u5_mult_79_n1770), .ZN(
        u5_mult_79_ab_18__2_) );
  NOR2_X2 u5_mult_79_U611 ( .A1(u5_mult_79_n1820), .A2(u5_mult_79_n1731), .ZN(
        u5_mult_79_ab_5__4_) );
  NOR2_X1 u5_mult_79_U610 ( .A1(u5_mult_79_n1832), .A2(u5_mult_79_n1773), .ZN(
        u5_mult_79_ab_19__23_) );
  NOR2_X1 u5_mult_79_U609 ( .A1(u5_mult_79_n1781), .A2(u5_mult_79_n1776), .ZN(
        u5_mult_79_ab_20__22_) );
  NOR2_X2 u5_mult_79_U608 ( .A1(u5_mult_79_n1817), .A2(u5_mult_79_n1734), .ZN(
        u5_mult_79_ab_6__5_) );
  NOR2_X2 u5_mult_79_U607 ( .A1(u5_mult_79_n1821), .A2(u5_mult_79_n1767), .ZN(
        u5_mult_79_ab_17__4_) );
  INV_X8 u5_mult_79_U606 ( .A(u5_mult_79_n1873), .ZN(u5_mult_79_n1816) );
  NOR2_X1 u5_mult_79_U605 ( .A1(u5_mult_79_n1794), .A2(u5_mult_79_n1776), .ZN(
        u5_mult_79_ab_20__16_) );
  NOR2_X1 u5_mult_79_U604 ( .A1(u5_mult_79_n1791), .A2(u5_mult_79_n1776), .ZN(
        u5_mult_79_ab_20__17_) );
  NOR2_X1 u5_mult_79_U603 ( .A1(u5_mult_79_n1788), .A2(u5_mult_79_n1776), .ZN(
        u5_mult_79_ab_20__18_) );
  NOR2_X1 u5_mult_79_U602 ( .A1(u5_mult_79_n1868), .A2(u5_mult_79_n1776), .ZN(
        u5_mult_79_ab_20__13_) );
  NOR2_X1 u5_mult_79_U601 ( .A1(u5_mult_79_n1783), .A2(u5_mult_79_n1776), .ZN(
        u5_mult_79_ab_20__21_) );
  NOR2_X1 u5_mult_79_U600 ( .A1(u5_mult_79_n1338), .A2(u5_mult_79_n1776), .ZN(
        u5_mult_79_ab_20__20_) );
  NOR2_X2 u5_mult_79_U599 ( .A1(u5_mult_79_n1808), .A2(u5_mult_79_n1728), .ZN(
        u5_mult_79_ab_4__8_) );
  NOR2_X2 u5_mult_79_U598 ( .A1(u5_mult_79_n1805), .A2(u5_mult_79_n1728), .ZN(
        u5_mult_79_ab_4__9_) );
  NAND3_X2 u5_mult_79_U597 ( .A1(u5_mult_79_n708), .A2(u5_mult_79_n709), .A3(
        u5_mult_79_n710), .ZN(u5_mult_79_CARRYB_9__7_) );
  NOR2_X2 u5_mult_79_U596 ( .A1(u5_mult_79_n1811), .A2(u5_mult_79_n1746), .ZN(
        u5_mult_79_ab_10__7_) );
  INV_X16 u5_mult_79_U595 ( .A(u5_mult_79_n1813), .ZN(u5_mult_79_n1812) );
  NOR2_X2 u5_mult_79_U594 ( .A1(u5_mult_79_n1805), .A2(u5_mult_79_n1743), .ZN(
        u5_mult_79_ab_9__9_) );
  NOR2_X2 u5_mult_79_U593 ( .A1(u5_mult_79_n1802), .A2(u5_mult_79_n1728), .ZN(
        u5_mult_79_ab_4__10_) );
  NOR2_X2 u5_mult_79_U592 ( .A1(u5_mult_79_n1802), .A2(u5_mult_79_n1743), .ZN(
        u5_mult_79_ab_9__10_) );
  NOR2_X1 u5_mult_79_U591 ( .A1(u5_mult_79_n1783), .A2(u5_mult_79_n1756), .ZN(
        u5_mult_79_ab_13__21_) );
  NOR2_X1 u5_mult_79_U590 ( .A1(u5_mult_79_n1338), .A2(u5_mult_79_n1756), .ZN(
        u5_mult_79_ab_13__20_) );
  NOR2_X1 u5_mult_79_U589 ( .A1(u5_mult_79_n1781), .A2(u5_mult_79_n1759), .ZN(
        u5_mult_79_ab_14__22_) );
  INV_X4 u5_mult_79_U588 ( .A(u5_mult_79_ab_5__12_), .ZN(u5_mult_79_n545) );
  NOR2_X1 u5_mult_79_U587 ( .A1(u5_mult_79_n1785), .A2(u5_mult_79_n1753), .ZN(
        u5_mult_79_ab_12__19_) );
  NOR2_X1 u5_mult_79_U586 ( .A1(u5_mult_79_n1788), .A2(u5_mult_79_n1753), .ZN(
        u5_mult_79_ab_12__18_) );
  INV_X4 u5_mult_79_U585 ( .A(u5_mult_79_ab_12__11_), .ZN(u5_mult_79_n1360) );
  INV_X2 u5_mult_79_U584 ( .A(u5_mult_79_ab_14__14_), .ZN(u5_mult_79_n1526) );
  XNOR2_X2 u5_mult_79_U583 ( .A(u5_mult_79_n166), .B(u5_mult_79_ab_15__16_), 
        .ZN(u5_mult_79_n481) );
  NAND2_X2 u5_mult_79_U582 ( .A1(u5_mult_79_ab_10__19_), .A2(
        u5_mult_79_CARRYB_9__19_), .ZN(u5_mult_79_n762) );
  NAND2_X2 u5_mult_79_U581 ( .A1(u5_mult_79_ab_18__13_), .A2(
        u5_mult_79_CARRYB_17__13_), .ZN(u5_mult_79_n953) );
  NAND2_X2 u5_mult_79_U580 ( .A1(u5_mult_79_SUMB_17__14_), .A2(
        u5_mult_79_CARRYB_17__13_), .ZN(u5_mult_79_n955) );
  NAND3_X4 u5_mult_79_U579 ( .A1(u5_mult_79_n1337), .A2(u5_mult_79_n1336), 
        .A3(u5_mult_79_n1335), .ZN(u5_mult_79_CARRYB_16__13_) );
  NOR2_X1 u5_mult_79_U578 ( .A1(u5_mult_79_n1868), .A2(u5_mult_79_n1768), .ZN(
        u5_mult_79_ab_17__13_) );
  NAND2_X2 u5_mult_79_U577 ( .A1(u5_mult_79_ab_14__16_), .A2(
        u5_mult_79_CARRYB_13__16_), .ZN(u5_mult_79_n1436) );
  NOR2_X1 u5_mult_79_U576 ( .A1(u5_mult_79_n1794), .A2(u5_mult_79_n1756), .ZN(
        u5_mult_79_ab_13__16_) );
  INV_X8 u5_mult_79_U575 ( .A(u5_mult_79_n1833), .ZN(u5_mult_79_n1831) );
  INV_X4 u5_mult_79_U574 ( .A(u5_mult_79_n1833), .ZN(u5_mult_79_n1832) );
  NAND2_X1 u5_mult_79_U573 ( .A1(u5_mult_79_ab_9__19_), .A2(
        u5_mult_79_CARRYB_8__19_), .ZN(u5_mult_79_n227) );
  NAND2_X2 u5_mult_79_U572 ( .A1(u5_mult_79_ab_9__19_), .A2(
        u5_mult_79_SUMB_8__20_), .ZN(u5_mult_79_n226) );
  XOR2_X2 u5_mult_79_U571 ( .A(u5_mult_79_SUMB_8__20_), .B(u5_mult_79_n224), 
        .Z(u5_mult_79_SUMB_9__19_) );
  XOR2_X2 u5_mult_79_U570 ( .A(u5_mult_79_CARRYB_8__19_), .B(
        u5_mult_79_ab_9__19_), .Z(u5_mult_79_n224) );
  NAND3_X4 u5_mult_79_U569 ( .A1(u5_mult_79_n221), .A2(u5_mult_79_n222), .A3(
        u5_mult_79_n223), .ZN(u5_mult_79_CARRYB_17__13_) );
  NAND2_X1 u5_mult_79_U568 ( .A1(u5_mult_79_ab_17__13_), .A2(
        u5_mult_79_CARRYB_16__13_), .ZN(u5_mult_79_n223) );
  NAND2_X2 u5_mult_79_U567 ( .A1(u5_mult_79_ab_17__13_), .A2(u5_mult_79_n40), 
        .ZN(u5_mult_79_n222) );
  NAND2_X2 u5_mult_79_U566 ( .A1(u5_mult_79_CARRYB_16__13_), .A2(
        u5_mult_79_n40), .ZN(u5_mult_79_n221) );
  NAND3_X2 u5_mult_79_U565 ( .A1(u5_mult_79_n218), .A2(u5_mult_79_n219), .A3(
        u5_mult_79_n220), .ZN(u5_mult_79_CARRYB_13__16_) );
  NAND2_X1 u5_mult_79_U564 ( .A1(u5_mult_79_ab_13__16_), .A2(
        u5_mult_79_CARRYB_12__16_), .ZN(u5_mult_79_n220) );
  NAND2_X2 u5_mult_79_U563 ( .A1(u5_mult_79_ab_13__16_), .A2(
        u5_mult_79_SUMB_12__17_), .ZN(u5_mult_79_n219) );
  NAND2_X1 u5_mult_79_U562 ( .A1(u5_mult_79_CARRYB_12__16_), .A2(
        u5_mult_79_SUMB_12__17_), .ZN(u5_mult_79_n218) );
  XOR2_X2 u5_mult_79_U561 ( .A(u5_mult_79_n38), .B(u5_mult_79_n217), .Z(
        u5_mult_79_SUMB_13__16_) );
  XOR2_X2 u5_mult_79_U560 ( .A(u5_mult_79_CARRYB_12__16_), .B(
        u5_mult_79_ab_13__16_), .Z(u5_mult_79_n217) );
  NAND3_X2 u5_mult_79_U559 ( .A1(u5_mult_79_n214), .A2(u5_mult_79_n215), .A3(
        u5_mult_79_n216), .ZN(u5_mult_79_CARRYB_21__11_) );
  NAND2_X1 u5_mult_79_U558 ( .A1(u5_mult_79_ab_21__11_), .A2(
        u5_mult_79_CARRYB_20__11_), .ZN(u5_mult_79_n216) );
  NAND2_X2 u5_mult_79_U557 ( .A1(u5_mult_79_ab_21__11_), .A2(
        u5_mult_79_SUMB_20__12_), .ZN(u5_mult_79_n215) );
  NAND2_X1 u5_mult_79_U556 ( .A1(u5_mult_79_SUMB_20__12_), .A2(
        u5_mult_79_CARRYB_20__11_), .ZN(u5_mult_79_n214) );
  NAND2_X2 u5_mult_79_U555 ( .A1(u5_mult_79_SUMB_1__17_), .A2(
        u5_mult_79_ab_2__16_), .ZN(u5_mult_79_n1184) );
  NAND2_X1 u5_mult_79_U554 ( .A1(u5_mult_79_SUMB_1__17_), .A2(
        u5_mult_79_CARRYB_1__16_), .ZN(u5_mult_79_n1183) );
  CLKBUF_X3 u5_mult_79_U553 ( .A(u5_mult_79_CARRYB_10__21_), .Z(
        u5_mult_79_n439) );
  NAND3_X2 u5_mult_79_U552 ( .A1(u5_mult_79_n991), .A2(u5_mult_79_n990), .A3(
        u5_mult_79_n989), .ZN(u5_mult_79_CARRYB_11__9_) );
  INV_X4 u5_mult_79_U551 ( .A(u5_mult_79_n211), .ZN(u5_mult_79_n212) );
  INV_X2 u5_mult_79_U550 ( .A(u5_mult_79_CARRYB_9__22_), .ZN(u5_mult_79_n211)
         );
  NAND2_X2 u5_mult_79_U549 ( .A1(u5_mult_79_ab_12__21_), .A2(
        u5_mult_79_CARRYB_11__21_), .ZN(u5_mult_79_n1078) );
  NAND3_X4 u5_mult_79_U548 ( .A1(u5_mult_79_n532), .A2(u5_mult_79_n533), .A3(
        u5_mult_79_n534), .ZN(u5_mult_79_CARRYB_17__19_) );
  NOR2_X1 u5_mult_79_U547 ( .A1(u5_mult_79_n1785), .A2(u5_mult_79_n1771), .ZN(
        u5_mult_79_ab_18__19_) );
  NOR2_X1 u5_mult_79_U546 ( .A1(u5_mult_79_n1831), .A2(u5_mult_79_n1734), .ZN(
        u5_mult_79_ab_6__23_) );
  NOR2_X1 u5_mult_79_U545 ( .A1(u5_mult_79_n1780), .A2(u5_mult_79_n1738), .ZN(
        u5_mult_79_ab_7__22_) );
  NAND3_X2 u5_mult_79_U544 ( .A1(u5_mult_79_n208), .A2(u5_mult_79_n209), .A3(
        u5_mult_79_n210), .ZN(u5_mult_79_CARRYB_18__19_) );
  NAND2_X1 u5_mult_79_U543 ( .A1(u5_mult_79_ab_18__19_), .A2(
        u5_mult_79_CARRYB_17__19_), .ZN(u5_mult_79_n210) );
  NAND2_X1 u5_mult_79_U542 ( .A1(u5_mult_79_ab_18__19_), .A2(
        u5_mult_79_SUMB_17__20_), .ZN(u5_mult_79_n209) );
  NAND2_X1 u5_mult_79_U541 ( .A1(u5_mult_79_CARRYB_17__19_), .A2(
        u5_mult_79_SUMB_17__20_), .ZN(u5_mult_79_n208) );
  NAND3_X2 u5_mult_79_U540 ( .A1(u5_mult_79_n205), .A2(u5_mult_79_n206), .A3(
        u5_mult_79_n207), .ZN(u5_mult_79_CARRYB_7__22_) );
  NAND2_X2 u5_mult_79_U539 ( .A1(u5_mult_79_ab_7__22_), .A2(
        u5_mult_79_ab_6__23_), .ZN(u5_mult_79_n207) );
  NAND2_X2 u5_mult_79_U538 ( .A1(u5_mult_79_ab_7__22_), .A2(
        u5_mult_79_CARRYB_6__22_), .ZN(u5_mult_79_n206) );
  NAND2_X2 u5_mult_79_U537 ( .A1(u5_mult_79_ab_6__23_), .A2(
        u5_mult_79_CARRYB_6__22_), .ZN(u5_mult_79_n205) );
  XOR2_X2 u5_mult_79_U536 ( .A(u5_mult_79_CARRYB_6__22_), .B(u5_mult_79_n204), 
        .Z(u5_mult_79_SUMB_7__22_) );
  XOR2_X2 u5_mult_79_U535 ( .A(u5_mult_79_ab_6__23_), .B(u5_mult_79_ab_7__22_), 
        .Z(u5_mult_79_n204) );
  XNOR2_X2 u5_mult_79_U534 ( .A(u5_mult_79_CARRYB_14__14_), .B(
        u5_mult_79_ab_15__14_), .ZN(u5_mult_79_n461) );
  NAND2_X2 u5_mult_79_U533 ( .A1(u5_mult_79_SUMB_10__17_), .A2(
        u5_mult_79_ab_11__16_), .ZN(u5_mult_79_n820) );
  NAND3_X4 u5_mult_79_U532 ( .A1(u5_mult_79_n1182), .A2(u5_mult_79_n1183), 
        .A3(u5_mult_79_n1184), .ZN(u5_mult_79_CARRYB_2__16_) );
  NAND2_X2 u5_mult_79_U531 ( .A1(u5_mult_79_n27), .A2(u5_mult_79_SUMB_6__14_), 
        .ZN(u5_mult_79_n1417) );
  NAND2_X2 u5_mult_79_U530 ( .A1(u5_mult_79_ab_16__17_), .A2(u5_mult_79_n130), 
        .ZN(u5_mult_79_n572) );
  NAND3_X4 u5_mult_79_U529 ( .A1(u5_mult_79_n819), .A2(u5_mult_79_n820), .A3(
        u5_mult_79_n821), .ZN(u5_mult_79_CARRYB_11__16_) );
  NAND2_X2 u5_mult_79_U528 ( .A1(u5_mult_79_n893), .A2(u5_mult_79_n472), .ZN(
        u5_mult_79_n896) );
  NAND3_X4 u5_mult_79_U527 ( .A1(u5_mult_79_n1518), .A2(u5_mult_79_n1519), 
        .A3(u5_mult_79_n1520), .ZN(u5_mult_79_CARRYB_19__10_) );
  NAND2_X2 u5_mult_79_U526 ( .A1(u5_mult_79_SUMB_11__22_), .A2(
        u5_mult_79_CARRYB_11__21_), .ZN(u5_mult_79_n1077) );
  NAND2_X1 u5_mult_79_U525 ( .A1(u5_mult_79_ab_12__21_), .A2(
        u5_mult_79_SUMB_11__22_), .ZN(u5_mult_79_n1079) );
  NAND2_X2 u5_mult_79_U524 ( .A1(u5_mult_79_SUMB_6__22_), .A2(
        u5_mult_79_CARRYB_6__21_), .ZN(u5_mult_79_n1065) );
  NAND2_X2 u5_mult_79_U523 ( .A1(u5_mult_79_ab_12__7_), .A2(
        u5_mult_79_SUMB_11__8_), .ZN(u5_mult_79_n1095) );
  NAND2_X2 u5_mult_79_U522 ( .A1(u5_mult_79_CARRYB_15__6_), .A2(
        u5_mult_79_SUMB_15__7_), .ZN(u5_mult_79_n1576) );
  NAND2_X2 u5_mult_79_U521 ( .A1(u5_mult_79_CARRYB_17__14_), .A2(
        u5_mult_79_SUMB_17__15_), .ZN(u5_mult_79_n1141) );
  NAND2_X1 u5_mult_79_U520 ( .A1(u5_mult_79_SUMB_23__11_), .A2(
        u5_mult_79_CARRYB_23__10_), .ZN(u5_mult_79_n1658) );
  INV_X4 u5_mult_79_U519 ( .A(u5_mult_79_n1789), .ZN(u5_mult_79_n1788) );
  XNOR2_X1 u5_mult_79_U518 ( .A(u5_mult_79_n783), .B(u5_mult_79_ab_18__6_), 
        .ZN(u5_mult_79_n1512) );
  NAND2_X2 u5_mult_79_U517 ( .A1(u5_mult_79_SUMB_17__12_), .A2(
        u5_mult_79_CARRYB_17__11_), .ZN(u5_mult_79_n1517) );
  NAND2_X2 u5_mult_79_U516 ( .A1(u5_mult_79_SUMB_6__17_), .A2(
        u5_mult_79_ab_7__16_), .ZN(u5_mult_79_n1396) );
  NAND2_X2 u5_mult_79_U515 ( .A1(u5_mult_79_CARRYB_6__16_), .A2(
        u5_mult_79_SUMB_6__17_), .ZN(u5_mult_79_n1397) );
  NAND2_X2 u5_mult_79_U514 ( .A1(u5_mult_79_CARRYB_10__13_), .A2(
        u5_mult_79_n45), .ZN(u5_mult_79_n1420) );
  NAND2_X2 u5_mult_79_U513 ( .A1(u5_mult_79_ab_21__7_), .A2(
        u5_mult_79_CARRYB_20__7_), .ZN(u5_mult_79_n816) );
  NAND3_X2 u5_mult_79_U512 ( .A1(u5_mult_79_n201), .A2(u5_mult_79_n202), .A3(
        u5_mult_79_n203), .ZN(u5_mult_79_CARRYB_21__13_) );
  NAND2_X1 u5_mult_79_U511 ( .A1(u5_mult_79_ab_21__13_), .A2(
        u5_mult_79_SUMB_20__14_), .ZN(u5_mult_79_n203) );
  NAND2_X1 u5_mult_79_U510 ( .A1(u5_mult_79_CARRYB_20__13_), .A2(
        u5_mult_79_SUMB_20__14_), .ZN(u5_mult_79_n202) );
  NAND2_X1 u5_mult_79_U509 ( .A1(u5_mult_79_CARRYB_20__13_), .A2(
        u5_mult_79_ab_21__13_), .ZN(u5_mult_79_n201) );
  NAND3_X4 u5_mult_79_U508 ( .A1(u5_mult_79_n198), .A2(u5_mult_79_n199), .A3(
        u5_mult_79_n200), .ZN(u5_mult_79_CARRYB_20__14_) );
  NAND2_X2 u5_mult_79_U507 ( .A1(u5_mult_79_ab_20__14_), .A2(
        u5_mult_79_SUMB_19__15_), .ZN(u5_mult_79_n200) );
  NAND2_X2 u5_mult_79_U506 ( .A1(u5_mult_79_CARRYB_19__14_), .A2(
        u5_mult_79_SUMB_19__15_), .ZN(u5_mult_79_n199) );
  NAND2_X1 u5_mult_79_U505 ( .A1(u5_mult_79_CARRYB_19__14_), .A2(
        u5_mult_79_ab_20__14_), .ZN(u5_mult_79_n198) );
  XOR2_X2 u5_mult_79_U504 ( .A(u5_mult_79_n197), .B(u5_mult_79_SUMB_20__14_), 
        .Z(u5_mult_79_SUMB_21__13_) );
  XOR2_X2 u5_mult_79_U503 ( .A(u5_mult_79_CARRYB_20__13_), .B(
        u5_mult_79_ab_21__13_), .Z(u5_mult_79_n197) );
  XOR2_X2 u5_mult_79_U502 ( .A(u5_mult_79_n196), .B(u5_mult_79_n17), .Z(
        u5_mult_79_SUMB_20__14_) );
  XOR2_X2 u5_mult_79_U501 ( .A(u5_mult_79_CARRYB_19__14_), .B(
        u5_mult_79_ab_20__14_), .Z(u5_mult_79_n196) );
  INV_X4 u5_mult_79_U500 ( .A(u5_mult_79_SUMB_11__10_), .ZN(u5_mult_79_n363)
         );
  NAND3_X4 u5_mult_79_U499 ( .A1(u5_mult_79_n699), .A2(u5_mult_79_n700), .A3(
        u5_mult_79_n701), .ZN(u5_mult_79_CARRYB_5__12_) );
  INV_X8 u5_mult_79_U498 ( .A(u5_mult_79_n432), .ZN(u5_mult_79_n433) );
  CLKBUF_X3 u5_mult_79_U497 ( .A(u5_mult_79_SUMB_14__8_), .Z(u5_mult_79_n347)
         );
  BUF_X8 u5_mult_79_U496 ( .A(u5_mult_79_SUMB_17__7_), .Z(u5_mult_79_n352) );
  NOR2_X4 u5_mult_79_U495 ( .A1(u5_mult_79_n1812), .A2(u5_mult_79_n1767), .ZN(
        u5_mult_79_ab_17__7_) );
  NAND3_X2 u5_mult_79_U494 ( .A1(u5_mult_79_n1480), .A2(u5_mult_79_n1481), 
        .A3(u5_mult_79_n1482), .ZN(u5_mult_79_n195) );
  INV_X1 u5_mult_79_U493 ( .A(u5_mult_79_ab_17__7_), .ZN(u5_mult_79_n192) );
  INV_X4 u5_mult_79_U492 ( .A(u5_mult_79_n195), .ZN(u5_mult_79_n191) );
  NAND2_X4 u5_mult_79_U491 ( .A1(u5_mult_79_n193), .A2(u5_mult_79_n194), .ZN(
        u5_mult_79_n1302) );
  NAND2_X4 u5_mult_79_U490 ( .A1(u5_mult_79_n191), .A2(u5_mult_79_n192), .ZN(
        u5_mult_79_n194) );
  NAND2_X2 u5_mult_79_U489 ( .A1(u5_mult_79_n195), .A2(u5_mult_79_ab_17__7_), 
        .ZN(u5_mult_79_n193) );
  NAND3_X4 u5_mult_79_U488 ( .A1(u5_mult_79_n1395), .A2(u5_mult_79_n1396), 
        .A3(u5_mult_79_n1397), .ZN(u5_mult_79_CARRYB_7__16_) );
  XNOR2_X2 u5_mult_79_U487 ( .A(u5_mult_79_CARRYB_17__12_), .B(
        u5_mult_79_ab_18__12_), .ZN(u5_mult_79_n394) );
  NAND2_X4 u5_mult_79_U486 ( .A1(u5_mult_79_n895), .A2(u5_mult_79_n896), .ZN(
        u5_mult_79_SUMB_14__14_) );
  XNOR2_X2 u5_mult_79_U485 ( .A(u5_mult_79_ab_7__17_), .B(
        u5_mult_79_CARRYB_6__17_), .ZN(u5_mult_79_n398) );
  NAND2_X2 u5_mult_79_U484 ( .A1(u5_mult_79_ab_15__12_), .A2(
        u5_mult_79_CARRYB_14__12_), .ZN(u5_mult_79_n1362) );
  NAND3_X2 u5_mult_79_U483 ( .A1(u5_mult_79_n1362), .A2(u5_mult_79_n1364), 
        .A3(u5_mult_79_n1363), .ZN(u5_mult_79_CARRYB_15__12_) );
  XNOR2_X1 u5_mult_79_U482 ( .A(u5_mult_79_n1339), .B(u5_mult_79_SUMB_4__14_), 
        .ZN(u5_mult_79_n190) );
  XNOR2_X2 u5_mult_79_U481 ( .A(u5_mult_79_n1122), .B(u5_mult_79_n190), .ZN(
        u5_mult_79_SUMB_6__12_) );
  XNOR2_X2 u5_mult_79_U480 ( .A(u5_mult_79_SUMB_17__16_), .B(u5_mult_79_n272), 
        .ZN(u5_mult_79_SUMB_18__15_) );
  NAND2_X2 u5_mult_79_U479 ( .A1(u5_mult_79_ab_12__6_), .A2(
        u5_mult_79_SUMB_11__7_), .ZN(u5_mult_79_n1110) );
  CLKBUF_X2 u5_mult_79_U478 ( .A(u5_mult_79_SUMB_10__8_), .Z(u5_mult_79_n358)
         );
  INV_X8 u5_mult_79_U477 ( .A(u5_mult_79_n1133), .ZN(u5_mult_79_n1134) );
  INV_X8 u5_mult_79_U476 ( .A(n2526), .ZN(u5_mult_79_n1860) );
  INV_X4 u5_mult_79_U475 ( .A(u5_mult_79_n1860), .ZN(u5_mult_79_n1784) );
  NAND2_X2 u5_mult_79_U474 ( .A1(u5_mult_79_CARRYB_11__6_), .A2(
        u5_mult_79_SUMB_11__7_), .ZN(u5_mult_79_n1111) );
  CLKBUF_X3 u5_mult_79_U473 ( .A(u5_mult_79_SUMB_16__10_), .Z(u5_mult_79_n389)
         );
  NAND2_X2 u5_mult_79_U472 ( .A1(u5_mult_79_ab_12__11_), .A2(
        u5_mult_79_CARRYB_11__11_), .ZN(u5_mult_79_n1405) );
  NOR2_X2 u5_mult_79_U471 ( .A1(u5_mult_79_n1801), .A2(u5_mult_79_n1750), .ZN(
        u5_mult_79_ab_11__11_) );
  NAND2_X4 u5_mult_79_U470 ( .A1(u5_mult_79_n559), .A2(u5_mult_79_n560), .ZN(
        u5_mult_79_n1565) );
  NAND3_X4 u5_mult_79_U469 ( .A1(u5_mult_79_n187), .A2(u5_mult_79_n188), .A3(
        u5_mult_79_n189), .ZN(u5_mult_79_CARRYB_11__11_) );
  NAND2_X2 u5_mult_79_U468 ( .A1(u5_mult_79_ab_11__11_), .A2(
        u5_mult_79_SUMB_10__12_), .ZN(u5_mult_79_n188) );
  NAND2_X2 u5_mult_79_U467 ( .A1(u5_mult_79_CARRYB_10__11_), .A2(
        u5_mult_79_SUMB_10__12_), .ZN(u5_mult_79_n187) );
  NAND3_X2 u5_mult_79_U466 ( .A1(u5_mult_79_n184), .A2(u5_mult_79_n185), .A3(
        u5_mult_79_n186), .ZN(u5_mult_79_CARRYB_14__10_) );
  NAND2_X1 u5_mult_79_U465 ( .A1(u5_mult_79_ab_14__10_), .A2(
        u5_mult_79_CARRYB_13__10_), .ZN(u5_mult_79_n186) );
  NAND2_X1 u5_mult_79_U464 ( .A1(u5_mult_79_ab_14__10_), .A2(
        u5_mult_79_SUMB_13__11_), .ZN(u5_mult_79_n185) );
  NAND2_X1 u5_mult_79_U463 ( .A1(u5_mult_79_CARRYB_13__10_), .A2(
        u5_mult_79_SUMB_13__11_), .ZN(u5_mult_79_n184) );
  INV_X1 u5_mult_79_U462 ( .A(u5_mult_79_SUMB_17__10_), .ZN(u5_mult_79_n180)
         );
  INV_X4 u5_mult_79_U461 ( .A(u5_mult_79_n1565), .ZN(u5_mult_79_n179) );
  NAND2_X2 u5_mult_79_U460 ( .A1(u5_mult_79_n181), .A2(u5_mult_79_n182), .ZN(
        u5_mult_79_SUMB_18__9_) );
  NAND2_X2 u5_mult_79_U459 ( .A1(u5_mult_79_n1565), .A2(u5_mult_79_n180), .ZN(
        u5_mult_79_n181) );
  XNOR2_X2 u5_mult_79_U458 ( .A(u5_mult_79_ab_16__17_), .B(u5_mult_79_n130), 
        .ZN(u5_mult_79_n330) );
  INV_X32 u5_mult_79_U457 ( .A(u5_mult_79_ab_14__7_), .ZN(u5_mult_79_n178) );
  XNOR2_X2 u5_mult_79_U456 ( .A(u5_mult_79_n178), .B(u5_mult_79_n780), .ZN(
        u5_mult_79_n805) );
  NAND2_X1 u5_mult_79_U455 ( .A1(u5_mult_79_ab_21__9_), .A2(
        u5_mult_79_CARRYB_20__9_), .ZN(u5_mult_79_n1430) );
  NAND2_X2 u5_mult_79_U454 ( .A1(u5_mult_79_CARRYB_6__10_), .A2(
        u5_mult_79_SUMB_6__11_), .ZN(u5_mult_79_n1256) );
  NAND2_X2 u5_mult_79_U453 ( .A1(u5_mult_79_ab_7__10_), .A2(
        u5_mult_79_SUMB_6__11_), .ZN(u5_mult_79_n1255) );
  CLKBUF_X3 u5_mult_79_U452 ( .A(u5_mult_79_SUMB_17__13_), .Z(u5_mult_79_n441)
         );
  CLKBUF_X3 u5_mult_79_U451 ( .A(u5_mult_79_SUMB_21__11_), .Z(u5_mult_79_n494)
         );
  NAND2_X1 u5_mult_79_U450 ( .A1(u5_mult_79_ab_17__14_), .A2(
        u5_mult_79_CARRYB_16__14_), .ZN(u5_mult_79_n950) );
  NAND2_X1 u5_mult_79_U449 ( .A1(u5_mult_79_CARRYB_10__17_), .A2(
        u5_mult_79_SUMB_10__18_), .ZN(u5_mult_79_n740) );
  NAND2_X2 u5_mult_79_U448 ( .A1(u5_mult_79_CARRYB_10__7_), .A2(
        u5_mult_79_SUMB_10__8_), .ZN(u5_mult_79_n1108) );
  NAND2_X2 u5_mult_79_U447 ( .A1(u5_mult_79_ab_18__14_), .A2(
        u5_mult_79_SUMB_17__15_), .ZN(u5_mult_79_n1140) );
  NOR2_X4 u5_mult_79_U446 ( .A1(u5_mult_79_n1867), .A2(u5_mult_79_n1719), .ZN(
        u5_mult_79_ab_1__14_) );
  NAND2_X2 u5_mult_79_U445 ( .A1(u5_mult_79_CARRYB_12__8_), .A2(
        u5_mult_79_SUMB_12__9_), .ZN(u5_mult_79_n1470) );
  NAND2_X1 u5_mult_79_U444 ( .A1(u5_mult_79_ab_17__14_), .A2(
        u5_mult_79_SUMB_16__15_), .ZN(u5_mult_79_n951) );
  NAND2_X2 u5_mult_79_U443 ( .A1(u5_mult_79_ab_18__14_), .A2(
        u5_mult_79_CARRYB_17__14_), .ZN(u5_mult_79_n1139) );
  INV_X2 u5_mult_79_U442 ( .A(u5_mult_79_CARRYB_17__14_), .ZN(u5_mult_79_n849)
         );
  NAND2_X1 u5_mult_79_U441 ( .A1(u5_mult_79_n965), .A2(
        u5_mult_79_CARRYB_17__14_), .ZN(u5_mult_79_n850) );
  NAND2_X2 u5_mult_79_U440 ( .A1(u5_mult_79_ab_11__13_), .A2(u5_mult_79_n45), 
        .ZN(u5_mult_79_n1419) );
  NAND2_X2 u5_mult_79_U439 ( .A1(u5_mult_79_CARRYB_12__11_), .A2(
        u5_mult_79_SUMB_12__12_), .ZN(u5_mult_79_n1085) );
  CLKBUF_X3 u5_mult_79_U438 ( .A(u5_mult_79_SUMB_11__13_), .Z(u5_mult_79_n325)
         );
  XNOR2_X2 u5_mult_79_U437 ( .A(u5_mult_79_CARRYB_20__11_), .B(
        u5_mult_79_ab_21__11_), .ZN(u5_mult_79_n177) );
  XNOR2_X2 u5_mult_79_U436 ( .A(u5_mult_79_SUMB_20__12_), .B(u5_mult_79_n177), 
        .ZN(u5_mult_79_SUMB_21__11_) );
  NAND2_X2 u5_mult_79_U435 ( .A1(u5_mult_79_ab_9__14_), .A2(
        u5_mult_79_SUMB_8__15_), .ZN(u5_mult_79_n853) );
  NAND2_X2 u5_mult_79_U434 ( .A1(u5_mult_79_CARRYB_13__12_), .A2(
        u5_mult_79_n1426), .ZN(u5_mult_79_n1488) );
  NAND2_X1 u5_mult_79_U433 ( .A1(u5_mult_79_ab_18__9_), .A2(
        u5_mult_79_SUMB_17__10_), .ZN(u5_mult_79_n1570) );
  NAND2_X2 u5_mult_79_U432 ( .A1(u5_mult_79_n179), .A2(u5_mult_79_SUMB_17__10_), .ZN(u5_mult_79_n182) );
  NAND3_X2 u5_mult_79_U431 ( .A1(u5_mult_79_n174), .A2(u5_mult_79_n175), .A3(
        u5_mult_79_n176), .ZN(u5_mult_79_CARRYB_10__10_) );
  NAND2_X1 u5_mult_79_U430 ( .A1(u5_mult_79_ab_10__10_), .A2(
        u5_mult_79_SUMB_9__11_), .ZN(u5_mult_79_n176) );
  NAND2_X1 u5_mult_79_U429 ( .A1(u5_mult_79_CARRYB_9__10_), .A2(
        u5_mult_79_SUMB_9__11_), .ZN(u5_mult_79_n175) );
  NAND2_X1 u5_mult_79_U428 ( .A1(u5_mult_79_CARRYB_9__10_), .A2(
        u5_mult_79_ab_10__10_), .ZN(u5_mult_79_n174) );
  NAND3_X4 u5_mult_79_U427 ( .A1(u5_mult_79_n171), .A2(u5_mult_79_n172), .A3(
        u5_mult_79_n173), .ZN(u5_mult_79_CARRYB_9__11_) );
  NAND2_X2 u5_mult_79_U426 ( .A1(u5_mult_79_SUMB_8__12_), .A2(
        u5_mult_79_CARRYB_8__11_), .ZN(u5_mult_79_n173) );
  NAND2_X2 u5_mult_79_U425 ( .A1(u5_mult_79_ab_9__11_), .A2(
        u5_mult_79_SUMB_8__12_), .ZN(u5_mult_79_n172) );
  NAND2_X2 u5_mult_79_U424 ( .A1(u5_mult_79_ab_9__11_), .A2(
        u5_mult_79_CARRYB_8__11_), .ZN(u5_mult_79_n171) );
  NAND2_X1 u5_mult_79_U423 ( .A1(u5_mult_79_CARRYB_21__9_), .A2(
        u5_mult_79_SUMB_21__10_), .ZN(u5_mult_79_n1354) );
  NAND2_X2 u5_mult_79_U422 ( .A1(u5_mult_79_CARRYB_18__10_), .A2(
        u5_mult_79_SUMB_18__11_), .ZN(u5_mult_79_n1520) );
  NAND2_X2 u5_mult_79_U421 ( .A1(u5_mult_79_ab_22__8_), .A2(
        u5_mult_79_SUMB_21__9_), .ZN(u5_mult_79_n1434) );
  NAND2_X2 u5_mult_79_U420 ( .A1(u5_mult_79_SUMB_21__9_), .A2(
        u5_mult_79_CARRYB_21__8_), .ZN(u5_mult_79_n1435) );
  BUF_X8 u5_mult_79_U419 ( .A(u5_mult_79_SUMB_16__16_), .Z(u5_mult_79_n485) );
  NAND2_X4 u5_mult_79_U418 ( .A1(u5_mult_79_n832), .A2(u5_mult_79_n833), .ZN(
        u5_mult_79_SUMB_14__17_) );
  NAND2_X4 u5_mult_79_U417 ( .A1(u5_mult_79_n830), .A2(u5_mult_79_n831), .ZN(
        u5_mult_79_n833) );
  NAND3_X4 u5_mult_79_U416 ( .A1(u5_mult_79_n1576), .A2(u5_mult_79_n1577), 
        .A3(u5_mult_79_n1578), .ZN(u5_mult_79_CARRYB_16__6_) );
  XNOR2_X2 u5_mult_79_U415 ( .A(u5_mult_79_SUMB_6__16_), .B(
        u5_mult_79_ab_7__15_), .ZN(u5_mult_79_n348) );
  NAND2_X2 u5_mult_79_U414 ( .A1(u5_mult_79_SUMB_19__11_), .A2(
        u5_mult_79_CARRYB_19__10_), .ZN(u5_mult_79_n1427) );
  NAND2_X2 u5_mult_79_U413 ( .A1(u5_mult_79_SUMB_17__12_), .A2(
        u5_mult_79_ab_18__11_), .ZN(u5_mult_79_n1516) );
  NAND2_X2 u5_mult_79_U412 ( .A1(u5_mult_79_CARRYB_7__15_), .A2(
        u5_mult_79_SUMB_7__16_), .ZN(u5_mult_79_n1400) );
  NAND3_X2 u5_mult_79_U411 ( .A1(u5_mult_79_n168), .A2(u5_mult_79_n169), .A3(
        u5_mult_79_n170), .ZN(u5_mult_79_CARRYB_8__20_) );
  NAND2_X2 u5_mult_79_U410 ( .A1(u5_mult_79_ab_8__20_), .A2(
        u5_mult_79_CARRYB_7__20_), .ZN(u5_mult_79_n169) );
  NAND2_X1 u5_mult_79_U409 ( .A1(u5_mult_79_SUMB_7__21_), .A2(
        u5_mult_79_CARRYB_7__20_), .ZN(u5_mult_79_n168) );
  XOR2_X2 u5_mult_79_U408 ( .A(u5_mult_79_n36), .B(u5_mult_79_n167), .Z(
        u5_mult_79_SUMB_8__20_) );
  XOR2_X2 u5_mult_79_U407 ( .A(u5_mult_79_SUMB_7__21_), .B(
        u5_mult_79_ab_8__20_), .Z(u5_mult_79_n167) );
  NAND3_X2 u5_mult_79_U406 ( .A1(u5_mult_79_n1436), .A2(u5_mult_79_n1437), 
        .A3(u5_mult_79_n1438), .ZN(u5_mult_79_n166) );
  INV_X4 u5_mult_79_U405 ( .A(u5_mult_79_SUMB_22__12_), .ZN(u5_mult_79_n163)
         );
  INV_X4 u5_mult_79_U404 ( .A(u5_mult_79_n796), .ZN(u5_mult_79_n162) );
  NAND2_X2 u5_mult_79_U403 ( .A1(u5_mult_79_n164), .A2(u5_mult_79_n165), .ZN(
        u5_mult_79_SUMB_23__11_) );
  NAND2_X4 u5_mult_79_U402 ( .A1(u5_mult_79_n162), .A2(u5_mult_79_n163), .ZN(
        u5_mult_79_n165) );
  NAND2_X1 u5_mult_79_U401 ( .A1(u5_mult_79_n796), .A2(u5_mult_79_SUMB_22__12_), .ZN(u5_mult_79_n164) );
  NAND3_X4 u5_mult_79_U400 ( .A1(u5_mult_79_n159), .A2(u5_mult_79_n160), .A3(
        u5_mult_79_n161), .ZN(u5_mult_79_CARRYB_21__12_) );
  NAND2_X2 u5_mult_79_U399 ( .A1(u5_mult_79_CARRYB_20__12_), .A2(
        u5_mult_79_SUMB_20__13_), .ZN(u5_mult_79_n161) );
  NAND2_X2 u5_mult_79_U398 ( .A1(u5_mult_79_ab_21__12_), .A2(
        u5_mult_79_SUMB_20__13_), .ZN(u5_mult_79_n160) );
  NAND2_X1 u5_mult_79_U397 ( .A1(u5_mult_79_ab_21__12_), .A2(
        u5_mult_79_CARRYB_20__12_), .ZN(u5_mult_79_n159) );
  NAND3_X4 u5_mult_79_U396 ( .A1(u5_mult_79_n156), .A2(u5_mult_79_n157), .A3(
        u5_mult_79_n158), .ZN(u5_mult_79_CARRYB_20__13_) );
  NAND2_X2 u5_mult_79_U395 ( .A1(u5_mult_79_CARRYB_19__13_), .A2(
        u5_mult_79_SUMB_19__14_), .ZN(u5_mult_79_n158) );
  NAND2_X2 u5_mult_79_U394 ( .A1(u5_mult_79_ab_20__13_), .A2(
        u5_mult_79_SUMB_19__14_), .ZN(u5_mult_79_n157) );
  NAND2_X1 u5_mult_79_U393 ( .A1(u5_mult_79_ab_20__13_), .A2(
        u5_mult_79_CARRYB_19__13_), .ZN(u5_mult_79_n156) );
  XOR2_X2 u5_mult_79_U392 ( .A(u5_mult_79_n155), .B(u5_mult_79_SUMB_20__13_), 
        .Z(u5_mult_79_SUMB_21__12_) );
  XOR2_X2 u5_mult_79_U391 ( .A(u5_mult_79_ab_21__12_), .B(
        u5_mult_79_CARRYB_20__12_), .Z(u5_mult_79_n155) );
  XNOR2_X2 u5_mult_79_U390 ( .A(u5_mult_79_CARRYB_23__7_), .B(
        u5_mult_79_SUMB_23__8_), .ZN(u5_mult_79_n1654) );
  NAND2_X4 u5_mult_79_U389 ( .A1(u5_mult_79_n433), .A2(u5_mult_79_ab_11__9_), 
        .ZN(u5_mult_79_n990) );
  INV_X4 u5_mult_79_U388 ( .A(u5_mult_79_SUMB_10__10_), .ZN(u5_mult_79_n432)
         );
  XOR2_X2 u5_mult_79_U387 ( .A(u5_mult_79_n695), .B(u5_mult_79_SUMB_4__13_), 
        .Z(u5_mult_79_SUMB_5__12_) );
  NAND2_X4 u5_mult_79_U386 ( .A1(u5_mult_79_ab_16__6_), .A2(
        u5_mult_79_CARRYB_15__6_), .ZN(u5_mult_79_n1578) );
  NAND3_X2 u5_mult_79_U385 ( .A1(u5_mult_79_n1160), .A2(u5_mult_79_n1159), 
        .A3(u5_mult_79_n1158), .ZN(u5_mult_79_CARRYB_3__12_) );
  NAND3_X4 u5_mult_79_U384 ( .A1(u5_mult_79_n1427), .A2(u5_mult_79_n1428), 
        .A3(u5_mult_79_n1429), .ZN(u5_mult_79_CARRYB_20__10_) );
  NOR2_X4 u5_mult_79_U383 ( .A1(u5_mult_79_n1815), .A2(u5_mult_79_n1767), .ZN(
        u5_mult_79_ab_17__6_) );
  INV_X4 u5_mult_79_U382 ( .A(u5_mult_79_n778), .ZN(u5_mult_79_n151) );
  NAND2_X4 u5_mult_79_U381 ( .A1(u5_mult_79_n153), .A2(u5_mult_79_n154), .ZN(
        u5_mult_79_SUMB_4__15_) );
  NAND2_X4 u5_mult_79_U380 ( .A1(u5_mult_79_n151), .A2(u5_mult_79_n152), .ZN(
        u5_mult_79_n154) );
  NAND2_X2 u5_mult_79_U379 ( .A1(u5_mult_79_n778), .A2(u5_mult_79_SUMB_3__16_), 
        .ZN(u5_mult_79_n153) );
  NAND2_X1 u5_mult_79_U378 ( .A1(u5_mult_79_ab_17__6_), .A2(
        u5_mult_79_CARRYB_16__6_), .ZN(u5_mult_79_n150) );
  NAND2_X2 u5_mult_79_U377 ( .A1(u5_mult_79_ab_17__6_), .A2(
        u5_mult_79_SUMB_16__7_), .ZN(u5_mult_79_n149) );
  NAND2_X2 u5_mult_79_U376 ( .A1(u5_mult_79_CARRYB_16__6_), .A2(
        u5_mult_79_SUMB_16__7_), .ZN(u5_mult_79_n148) );
  XOR2_X2 u5_mult_79_U375 ( .A(u5_mult_79_n122), .B(u5_mult_79_n147), .Z(
        u5_mult_79_SUMB_17__6_) );
  XOR2_X2 u5_mult_79_U374 ( .A(u5_mult_79_CARRYB_16__6_), .B(
        u5_mult_79_ab_17__6_), .Z(u5_mult_79_n147) );
  XNOR2_X2 u5_mult_79_U373 ( .A(u5_mult_79_CARRYB_19__8_), .B(
        u5_mult_79_ab_20__8_), .ZN(u5_mult_79_n516) );
  NOR2_X4 u5_mult_79_U372 ( .A1(u5_mult_79_n1860), .A2(u5_mult_79_n1719), .ZN(
        u5_mult_79_n1121) );
  NAND2_X2 u5_mult_79_U371 ( .A1(u5_mult_79_CARRYB_18__15_), .A2(
        u5_mult_79_SUMB_18__16_), .ZN(u5_mult_79_n1011) );
  NAND2_X1 u5_mult_79_U370 ( .A1(u5_mult_79_CARRYB_19__15_), .A2(
        u5_mult_79_SUMB_19__16_), .ZN(u5_mult_79_n599) );
  INV_X2 u5_mult_79_U369 ( .A(u5_mult_79_SUMB_23__13_), .ZN(u5_mult_79_n392)
         );
  NOR2_X4 u5_mult_79_U368 ( .A1(u5_mult_79_n1882), .A2(u5_mult_79_n1860), .ZN(
        u5_mult_79_ab_0__21_) );
  NAND2_X4 u5_mult_79_U367 ( .A1(u5_mult_79_ab_16__9_), .A2(u5_mult_79_n448), 
        .ZN(u5_mult_79_n1607) );
  NAND2_X2 u5_mult_79_U366 ( .A1(u5_mult_79_ab_13__10_), .A2(
        u5_mult_79_CARRYB_12__10_), .ZN(u5_mult_79_n1409) );
  NAND3_X4 u5_mult_79_U365 ( .A1(u5_mult_79_n1408), .A2(u5_mult_79_n1410), 
        .A3(u5_mult_79_n1409), .ZN(u5_mult_79_CARRYB_13__10_) );
  NAND2_X4 u5_mult_79_U364 ( .A1(u5_mult_79_SUMB_7__18_), .A2(
        u5_mult_79_CARRYB_7__17_), .ZN(u5_mult_79_n1280) );
  XNOR2_X2 u5_mult_79_U363 ( .A(u5_mult_79_SUMB_4__20_), .B(
        u5_mult_79_ab_5__19_), .ZN(u5_mult_79_n319) );
  INV_X8 u5_mult_79_U362 ( .A(u5_mult_79_n1654), .ZN(u5_mult_79_CLA_SUM[31])
         );
  NAND2_X2 u5_mult_79_U361 ( .A1(u5_mult_79_ab_8__14_), .A2(
        u5_mult_79_CARRYB_7__14_), .ZN(u5_mult_79_n975) );
  NAND2_X1 u5_mult_79_U360 ( .A1(u5_mult_79_CARRYB_17__12_), .A2(
        u5_mult_79_SUMB_17__13_), .ZN(u5_mult_79_n1041) );
  NAND3_X2 u5_mult_79_U359 ( .A1(u5_mult_79_n144), .A2(u5_mult_79_n145), .A3(
        u5_mult_79_n146), .ZN(u5_mult_79_CARRYB_17__21_) );
  NAND2_X2 u5_mult_79_U358 ( .A1(u5_mult_79_ab_17__21_), .A2(
        u5_mult_79_SUMB_16__22_), .ZN(u5_mult_79_n146) );
  NAND2_X2 u5_mult_79_U357 ( .A1(u5_mult_79_ab_17__21_), .A2(
        u5_mult_79_CARRYB_16__21_), .ZN(u5_mult_79_n145) );
  NAND2_X2 u5_mult_79_U356 ( .A1(u5_mult_79_SUMB_16__22_), .A2(
        u5_mult_79_CARRYB_16__21_), .ZN(u5_mult_79_n144) );
  XOR2_X1 u5_mult_79_U355 ( .A(u5_mult_79_CARRYB_16__21_), .B(u5_mult_79_n143), 
        .Z(u5_mult_79_SUMB_17__21_) );
  XOR2_X2 u5_mult_79_U354 ( .A(u5_mult_79_SUMB_16__22_), .B(
        u5_mult_79_ab_17__21_), .Z(u5_mult_79_n143) );
  NAND3_X2 u5_mult_79_U353 ( .A1(u5_mult_79_n140), .A2(u5_mult_79_n141), .A3(
        u5_mult_79_n142), .ZN(u5_mult_79_CARRYB_21__17_) );
  NAND2_X1 u5_mult_79_U352 ( .A1(u5_mult_79_CARRYB_20__17_), .A2(
        u5_mult_79_SUMB_20__18_), .ZN(u5_mult_79_n142) );
  NAND2_X1 u5_mult_79_U351 ( .A1(u5_mult_79_ab_21__17_), .A2(
        u5_mult_79_SUMB_20__18_), .ZN(u5_mult_79_n141) );
  NAND2_X1 u5_mult_79_U350 ( .A1(u5_mult_79_ab_21__17_), .A2(
        u5_mult_79_CARRYB_20__17_), .ZN(u5_mult_79_n140) );
  NAND3_X4 u5_mult_79_U349 ( .A1(u5_mult_79_n137), .A2(u5_mult_79_n138), .A3(
        u5_mult_79_n139), .ZN(u5_mult_79_CARRYB_20__18_) );
  NAND2_X1 u5_mult_79_U348 ( .A1(u5_mult_79_CARRYB_19__18_), .A2(
        u5_mult_79_SUMB_19__19_), .ZN(u5_mult_79_n139) );
  NAND2_X1 u5_mult_79_U347 ( .A1(u5_mult_79_ab_20__18_), .A2(
        u5_mult_79_SUMB_19__19_), .ZN(u5_mult_79_n138) );
  NAND2_X1 u5_mult_79_U346 ( .A1(u5_mult_79_ab_20__18_), .A2(
        u5_mult_79_CARRYB_19__18_), .ZN(u5_mult_79_n137) );
  XOR2_X2 u5_mult_79_U345 ( .A(u5_mult_79_n136), .B(u5_mult_79_SUMB_20__18_), 
        .Z(u5_mult_79_SUMB_21__17_) );
  XOR2_X2 u5_mult_79_U344 ( .A(u5_mult_79_ab_21__17_), .B(
        u5_mult_79_CARRYB_20__17_), .Z(u5_mult_79_n136) );
  XOR2_X2 u5_mult_79_U343 ( .A(u5_mult_79_n135), .B(u5_mult_79_SUMB_19__19_), 
        .Z(u5_mult_79_SUMB_20__18_) );
  XOR2_X2 u5_mult_79_U342 ( .A(u5_mult_79_ab_20__18_), .B(
        u5_mult_79_CARRYB_19__18_), .Z(u5_mult_79_n135) );
  CLKBUF_X3 u5_mult_79_U341 ( .A(u5_mult_79_SUMB_3__15_), .Z(u5_mult_79_n357)
         );
  XNOR2_X2 u5_mult_79_U340 ( .A(u5_mult_79_ab_20__15_), .B(
        u5_mult_79_CARRYB_19__15_), .ZN(u5_mult_79_n134) );
  XNOR2_X2 u5_mult_79_U339 ( .A(u5_mult_79_n134), .B(u5_mult_79_SUMB_19__16_), 
        .ZN(u5_mult_79_SUMB_20__15_) );
  INV_X4 u5_mult_79_U338 ( .A(u5_mult_79_n132), .ZN(u5_mult_79_n133) );
  INV_X2 u5_mult_79_U337 ( .A(u5_mult_79_SUMB_14__6_), .ZN(u5_mult_79_n132) );
  XNOR2_X2 u5_mult_79_U336 ( .A(u5_mult_79_ab_8__15_), .B(
        u5_mult_79_CARRYB_7__15_), .ZN(u5_mult_79_n131) );
  XNOR2_X2 u5_mult_79_U335 ( .A(u5_mult_79_n131), .B(u5_mult_79_n291), .ZN(
        u5_mult_79_SUMB_8__15_) );
  INV_X4 u5_mult_79_U334 ( .A(u5_mult_79_n129), .ZN(u5_mult_79_n130) );
  INV_X2 u5_mult_79_U333 ( .A(u5_mult_79_CARRYB_15__17_), .ZN(u5_mult_79_n129)
         );
  XNOR2_X2 u5_mult_79_U332 ( .A(u5_mult_79_n578), .B(u5_mult_79_SUMB_4__19_), 
        .ZN(u5_mult_79_n128) );
  NAND2_X2 u5_mult_79_U331 ( .A1(u5_mult_79_ab_19__10_), .A2(u5_mult_79_n300), 
        .ZN(u5_mult_79_n1519) );
  XNOR2_X2 u5_mult_79_U330 ( .A(u5_mult_79_n439), .B(u5_mult_79_n910), .ZN(
        u5_mult_79_SUMB_11__21_) );
  NAND2_X1 u5_mult_79_U329 ( .A1(u5_mult_79_SUMB_6__21_), .A2(
        u5_mult_79_CARRYB_6__20_), .ZN(u5_mult_79_n1231) );
  XNOR2_X2 u5_mult_79_U328 ( .A(u5_mult_79_ab_11__13_), .B(
        u5_mult_79_CARRYB_10__13_), .ZN(u5_mult_79_n451) );
  XNOR2_X2 u5_mult_79_U327 ( .A(u5_mult_79_n458), .B(u5_mult_79_n448), .ZN(
        u5_mult_79_n127) );
  NAND3_X4 u5_mult_79_U326 ( .A1(u5_mult_79_n1635), .A2(u5_mult_79_n1636), 
        .A3(u5_mult_79_n1637), .ZN(u5_mult_79_CARRYB_21__3_) );
  XOR2_X2 u5_mult_79_U325 ( .A(u5_mult_79_CARRYB_13__10_), .B(
        u5_mult_79_ab_14__10_), .Z(u5_mult_79_n183) );
  XNOR2_X2 u5_mult_79_U324 ( .A(u5_mult_79_CARRYB_10__17_), .B(
        u5_mult_79_ab_11__17_), .ZN(u5_mult_79_n382) );
  NAND2_X1 u5_mult_79_U323 ( .A1(u5_mult_79_SUMB_6__21_), .A2(
        u5_mult_79_ab_7__20_), .ZN(u5_mult_79_n1230) );
  CLKBUF_X2 u5_mult_79_U322 ( .A(u5_mult_79_CARRYB_16__18_), .Z(
        u5_mult_79_n126) );
  CLKBUF_X2 u5_mult_79_U321 ( .A(u5_mult_79_SUMB_14__9_), .Z(u5_mult_79_n125)
         );
  NAND2_X1 u5_mult_79_U320 ( .A1(u5_mult_79_CARRYB_17__3_), .A2(
        u5_mult_79_ab_18__3_), .ZN(u5_mult_79_n1179) );
  CLKBUF_X2 u5_mult_79_U319 ( .A(u5_mult_79_n354), .Z(u5_mult_79_n124) );
  XNOR2_X2 u5_mult_79_U318 ( .A(u5_mult_79_ab_16__13_), .B(u5_mult_79_n430), 
        .ZN(u5_mult_79_n123) );
  XNOR2_X2 u5_mult_79_U317 ( .A(u5_mult_79_n123), .B(u5_mult_79_n37), .ZN(
        u5_mult_79_SUMB_16__13_) );
  NAND2_X1 u5_mult_79_U316 ( .A1(u5_mult_79_CARRYB_19__4_), .A2(
        u5_mult_79_SUMB_19__5_), .ZN(u5_mult_79_n1540) );
  NAND2_X2 u5_mult_79_U315 ( .A1(u5_mult_79_ab_18__6_), .A2(u5_mult_79_n783), 
        .ZN(u5_mult_79_n1594) );
  NAND3_X2 u5_mult_79_U314 ( .A1(u5_mult_79_n1320), .A2(u5_mult_79_n1319), 
        .A3(u5_mult_79_n1318), .ZN(u5_mult_79_CARRYB_15__9_) );
  XOR2_X2 u5_mult_79_U313 ( .A(u5_mult_79_SUMB_13__11_), .B(u5_mult_79_n183), 
        .Z(u5_mult_79_SUMB_14__10_) );
  CLKBUF_X3 u5_mult_79_U312 ( .A(u5_mult_79_SUMB_16__7_), .Z(u5_mult_79_n122)
         );
  CLKBUF_X2 u5_mult_79_U311 ( .A(u5_mult_79_n312), .Z(u5_mult_79_n121) );
  XNOR2_X2 u5_mult_79_U310 ( .A(u5_mult_79_n120), .B(u5_mult_79_SUMB_13__6_), 
        .ZN(u5_mult_79_SUMB_14__5_) );
  NAND2_X2 u5_mult_79_U309 ( .A1(u5_mult_79_ab_16__13_), .A2(u5_mult_79_n430), 
        .ZN(u5_mult_79_n1335) );
  NAND2_X2 u5_mult_79_U308 ( .A1(u5_mult_79_ab_4__21_), .A2(
        u5_mult_79_CARRYB_3__21_), .ZN(u5_mult_79_n1620) );
  NAND3_X2 u5_mult_79_U307 ( .A1(u5_mult_79_n1619), .A2(u5_mult_79_n1620), 
        .A3(u5_mult_79_n1621), .ZN(u5_mult_79_CARRYB_4__21_) );
  NAND2_X4 u5_mult_79_U306 ( .A1(u5_mult_79_ab_3__21_), .A2(u5_mult_79_n401), 
        .ZN(u5_mult_79_n1601) );
  CLKBUF_X3 u5_mult_79_U305 ( .A(u5_mult_79_SUMB_21__4_), .Z(u5_mult_79_n119)
         );
  XNOR2_X2 u5_mult_79_U304 ( .A(u5_mult_79_ab_19__5_), .B(
        u5_mult_79_CARRYB_18__5_), .ZN(u5_mult_79_n118) );
  XNOR2_X2 u5_mult_79_U303 ( .A(u5_mult_79_n118), .B(u5_mult_79_SUMB_18__6_), 
        .ZN(u5_mult_79_SUMB_19__5_) );
  NAND2_X2 u5_mult_79_U302 ( .A1(u5_mult_79_ab_12__9_), .A2(u5_mult_79_n103), 
        .ZN(u5_mult_79_n1465) );
  NAND2_X2 u5_mult_79_U301 ( .A1(u5_mult_79_ab_11__11_), .A2(
        u5_mult_79_CARRYB_10__11_), .ZN(u5_mult_79_n189) );
  NAND3_X4 u5_mult_79_U300 ( .A1(u5_mult_79_n1551), .A2(u5_mult_79_n1553), 
        .A3(u5_mult_79_n1552), .ZN(u5_mult_79_CARRYB_5__21_) );
  NOR2_X1 u5_mult_79_U299 ( .A1(u5_mult_79_n1831), .A2(u5_mult_79_n1752), .ZN(
        u5_mult_79_ab_12__23_) );
  XNOR2_X2 u5_mult_79_U298 ( .A(u5_mult_79_CARRYB_10__11_), .B(
        u5_mult_79_ab_11__11_), .ZN(u5_mult_79_n117) );
  XNOR2_X2 u5_mult_79_U297 ( .A(u5_mult_79_n35), .B(u5_mult_79_n117), .ZN(
        u5_mult_79_SUMB_11__11_) );
  XNOR2_X2 u5_mult_79_U296 ( .A(u5_mult_79_n829), .B(u5_mult_79_n433), .ZN(
        u5_mult_79_n116) );
  NAND2_X2 u5_mult_79_U295 ( .A1(u5_mult_79_ab_11__10_), .A2(
        u5_mult_79_SUMB_10__11_), .ZN(u5_mult_79_n1463) );
  NAND2_X1 u5_mult_79_U294 ( .A1(u5_mult_79_ab_10__11_), .A2(
        u5_mult_79_SUMB_9__12_), .ZN(u5_mult_79_n1460) );
  NAND2_X1 u5_mult_79_U293 ( .A1(u5_mult_79_CARRYB_9__11_), .A2(
        u5_mult_79_SUMB_9__12_), .ZN(u5_mult_79_n1461) );
  INV_X2 u5_mult_79_U292 ( .A(u5_mult_79_SUMB_9__12_), .ZN(u5_mult_79_n449) );
  XNOR2_X2 u5_mult_79_U291 ( .A(u5_mult_79_CARRYB_9__13_), .B(
        u5_mult_79_ab_10__13_), .ZN(u5_mult_79_n410) );
  INV_X2 u5_mult_79_U290 ( .A(u5_mult_79_n114), .ZN(u5_mult_79_n115) );
  INV_X4 u5_mult_79_U289 ( .A(u5_mult_79_n112), .ZN(u5_mult_79_n113) );
  INV_X4 u5_mult_79_U288 ( .A(u5_mult_79_SUMB_12__6_), .ZN(u5_mult_79_n112) );
  NAND3_X2 u5_mult_79_U287 ( .A1(u5_mult_79_n1540), .A2(u5_mult_79_n1541), 
        .A3(u5_mult_79_n1542), .ZN(u5_mult_79_n111) );
  XNOR2_X2 u5_mult_79_U286 ( .A(u5_mult_79_n514), .B(u5_mult_79_n494), .ZN(
        u5_mult_79_n110) );
  NAND2_X2 u5_mult_79_U285 ( .A1(u5_mult_79_ab_0__19_), .A2(
        u5_mult_79_ab_1__18_), .ZN(u5_mult_79_n1708) );
  XNOR2_X2 u5_mult_79_U284 ( .A(u5_mult_79_CARRYB_17__19_), .B(
        u5_mult_79_ab_18__19_), .ZN(u5_mult_79_n107) );
  XNOR2_X2 u5_mult_79_U283 ( .A(u5_mult_79_SUMB_17__20_), .B(u5_mult_79_n107), 
        .ZN(u5_mult_79_SUMB_18__19_) );
  CLKBUF_X2 u5_mult_79_U282 ( .A(u5_mult_79_SUMB_16__20_), .Z(u5_mult_79_n106)
         );
  INV_X2 u5_mult_79_U281 ( .A(u5_mult_79_n104), .ZN(u5_mult_79_n105) );
  INV_X2 u5_mult_79_U280 ( .A(u5_mult_79_SUMB_6__8_), .ZN(u5_mult_79_n104) );
  NAND2_X2 u5_mult_79_U279 ( .A1(u5_mult_79_ab_18__16_), .A2(
        u5_mult_79_CARRYB_17__16_), .ZN(u5_mult_79_n563) );
  NAND3_X2 u5_mult_79_U278 ( .A1(u5_mult_79_n991), .A2(u5_mult_79_n990), .A3(
        u5_mult_79_n989), .ZN(u5_mult_79_n103) );
  NAND3_X4 u5_mult_79_U277 ( .A1(u5_mult_79_n1327), .A2(u5_mult_79_n1328), 
        .A3(u5_mult_79_n1329), .ZN(u5_mult_79_CARRYB_14__9_) );
  NAND2_X2 u5_mult_79_U276 ( .A1(u5_mult_79_ab_15__9_), .A2(
        u5_mult_79_CARRYB_14__9_), .ZN(u5_mult_79_n1318) );
  XNOR2_X2 u5_mult_79_U275 ( .A(u5_mult_79_ab_9__11_), .B(
        u5_mult_79_CARRYB_8__11_), .ZN(u5_mult_79_n102) );
  XNOR2_X2 u5_mult_79_U274 ( .A(u5_mult_79_n102), .B(u5_mult_79_SUMB_8__12_), 
        .ZN(u5_mult_79_SUMB_9__11_) );
  NOR2_X2 u5_mult_79_U273 ( .A1(u5_mult_79_n1882), .A2(u5_mult_79_n1861), .ZN(
        u5_mult_79_ab_0__20_) );
  NOR2_X2 u5_mult_79_U272 ( .A1(u5_mult_79_n1882), .A2(u5_mult_79_n1790), .ZN(
        u5_mult_79_ab_0__17_) );
  NOR2_X2 u5_mult_79_U271 ( .A1(u5_mult_79_n1811), .A2(u5_mult_79_n1720), .ZN(
        u5_mult_79_ab_1__7_) );
  NOR2_X2 u5_mult_79_U270 ( .A1(u5_mult_79_n1793), .A2(u5_mult_79_n1720), .ZN(
        u5_mult_79_ab_1__16_) );
  NOR2_X2 u5_mult_79_U269 ( .A1(u5_mult_79_n1862), .A2(u5_mult_79_n1720), .ZN(
        u5_mult_79_ab_1__19_) );
  NOR2_X2 u5_mult_79_U268 ( .A1(u5_mult_79_n1860), .A2(u5_mult_79_n1720), .ZN(
        u5_mult_79_ab_1__21_) );
  INV_X4 u5_mult_79_U267 ( .A(u5_mult_79_CARRYB_13__7_), .ZN(u5_mult_79_n780)
         );
  NAND2_X4 u5_mult_79_U266 ( .A1(u5_mult_79_n133), .A2(u5_mult_79_ab_15__5_), 
        .ZN(u5_mult_79_n1499) );
  XNOR2_X2 u5_mult_79_U265 ( .A(u5_mult_79_CARRYB_9__10_), .B(
        u5_mult_79_ab_10__10_), .ZN(u5_mult_79_n101) );
  XNOR2_X2 u5_mult_79_U264 ( .A(u5_mult_79_n101), .B(u5_mult_79_SUMB_9__11_), 
        .ZN(u5_mult_79_SUMB_10__10_) );
  INV_X32 u5_mult_79_U263 ( .A(n3030), .ZN(u5_mult_79_n1882) );
  NAND3_X2 u5_mult_79_U262 ( .A1(u5_mult_79_n148), .A2(u5_mult_79_n149), .A3(
        u5_mult_79_n150), .ZN(u5_mult_79_CARRYB_17__6_) );
  INV_X4 u5_mult_79_U261 ( .A(u5_mult_79_CARRYB_17__6_), .ZN(u5_mult_79_n782)
         );
  XNOR2_X2 u5_mult_79_U260 ( .A(u5_mult_79_CARRYB_7__6_), .B(
        u5_mult_79_ab_8__6_), .ZN(u5_mult_79_n402) );
  XNOR2_X2 u5_mult_79_U259 ( .A(u5_mult_79_ab_14__4_), .B(
        u5_mult_79_CARRYB_13__4_), .ZN(u5_mult_79_n100) );
  XNOR2_X2 u5_mult_79_U258 ( .A(u5_mult_79_n100), .B(u5_mult_79_n417), .ZN(
        u5_mult_79_SUMB_14__4_) );
  CLKBUF_X2 u5_mult_79_U257 ( .A(u5_mult_79_SUMB_13__3_), .Z(u5_mult_79_n99)
         );
  XOR2_X2 u5_mult_79_U256 ( .A(u5_mult_79_n265), .B(u5_mult_79_CARRYB_8__7_), 
        .Z(u5_mult_79_n98) );
  XNOR2_X2 u5_mult_79_U255 ( .A(u5_mult_79_n98), .B(u5_mult_79_SUMB_8__8_), 
        .ZN(u5_mult_79_SUMB_9__7_) );
  XOR2_X2 u5_mult_79_U254 ( .A(u5_mult_79_CARRYB_23__0_), .B(
        u5_mult_79_SUMB_23__1_), .Z(u5_N24) );
  XNOR2_X2 u5_mult_79_U253 ( .A(u5_mult_79_n259), .B(u5_mult_79_n810), .ZN(
        u5_mult_79_n96) );
  XNOR2_X2 u5_mult_79_U252 ( .A(u5_mult_79_n306), .B(u5_mult_79_n96), .ZN(
        u5_mult_79_SUMB_19__2_) );
  CLKBUF_X3 u5_mult_79_U251 ( .A(u5_mult_79_CARRYB_16__2_), .Z(u5_mult_79_n331) );
  NAND2_X2 u5_mult_79_U250 ( .A1(u5_mult_79_ab_17__2_), .A2(u5_mult_79_n331), 
        .ZN(u5_mult_79_n862) );
  NAND2_X2 u5_mult_79_U249 ( .A1(u5_mult_79_n331), .A2(u5_mult_79_SUMB_16__3_), 
        .ZN(u5_mult_79_n864) );
  XNOR2_X2 u5_mult_79_U248 ( .A(u5_mult_79_ab_14__5_), .B(
        u5_mult_79_CARRYB_13__5_), .ZN(u5_mult_79_n120) );
  XNOR2_X2 u5_mult_79_U247 ( .A(u5_mult_79_CARRYB_4__5_), .B(
        u5_mult_79_ab_5__5_), .ZN(u5_mult_79_n95) );
  XNOR2_X2 u5_mult_79_U246 ( .A(u5_mult_79_n95), .B(u5_mult_79_SUMB_4__6_), 
        .ZN(u5_mult_79_SUMB_5__5_) );
  INV_X32 u5_mult_79_U245 ( .A(n3005), .ZN(u5_mult_79_n1868) );
  CLKBUF_X3 u5_mult_79_U244 ( .A(u5_mult_79_SUMB_19__3_), .Z(u5_mult_79_n109)
         );
  INV_X32 u5_mult_79_U243 ( .A(u5_mult_79_ab_21__0_), .ZN(u5_mult_79_n94) );
  XNOR2_X2 u5_mult_79_U242 ( .A(u5_mult_79_SUMB_20__1_), .B(u5_mult_79_n94), 
        .ZN(u5_mult_79_n653) );
  AND3_X4 u5_mult_79_U241 ( .A1(u5_mult_79_n650), .A2(u5_mult_79_n651), .A3(
        u5_mult_79_n652), .ZN(u5_mult_79_n93) );
  XNOR2_X2 u5_mult_79_U240 ( .A(u5_mult_79_n653), .B(u5_mult_79_n93), .ZN(
        u5_N21) );
  XNOR2_X2 u5_mult_79_U239 ( .A(u5_mult_79_n99), .B(u5_mult_79_n251), .ZN(
        u5_mult_79_SUMB_14__2_) );
  INV_X8 u5_mult_79_U238 ( .A(u6_N5), .ZN(u5_mult_79_n1874) );
  XNOR2_X2 u5_mult_79_U237 ( .A(u5_mult_79_n657), .B(u5_mult_79_n252), .ZN(
        u5_N19) );
  INV_X8 u5_mult_79_U236 ( .A(u5_mult_79_n249), .ZN(u5_mult_79_n250) );
  NOR2_X1 u5_mult_79_U235 ( .A1(u5_mult_79_n1834), .A2(u5_mult_79_n1773), .ZN(
        u5_mult_79_ab_19__0_) );
  INV_X4 u5_mult_79_U234 ( .A(u5_mult_79_SUMB_18__1_), .ZN(u5_mult_79_n249) );
  XNOR2_X2 u5_mult_79_U233 ( .A(u5_mult_79_n249), .B(u5_mult_79_ab_19__0_), 
        .ZN(u5_mult_79_n657) );
  XNOR2_X2 u5_mult_79_U232 ( .A(u5_mult_79_SUMB_10__4_), .B(
        u5_mult_79_ab_11__3_), .ZN(u5_mult_79_n92) );
  XNOR2_X2 u5_mult_79_U231 ( .A(u5_mult_79_n414), .B(u5_mult_79_n92), .ZN(
        u5_mult_79_SUMB_11__3_) );
  XNOR2_X1 u5_mult_79_U230 ( .A(u5_mult_79_CARRYB_10__2_), .B(
        u5_mult_79_ab_11__2_), .ZN(u5_mult_79_n908) );
  XNOR2_X1 u5_mult_79_U229 ( .A(u5_mult_79_CARRYB_12__1_), .B(
        u5_mult_79_ab_13__1_), .ZN(u5_mult_79_n91) );
  XNOR2_X2 u5_mult_79_U228 ( .A(u5_mult_79_n91), .B(u5_mult_79_SUMB_12__2_), 
        .ZN(u5_mult_79_SUMB_13__1_) );
  NAND2_X2 u5_mult_79_U227 ( .A1(u5_mult_79_ab_12__2_), .A2(
        u5_mult_79_CARRYB_11__2_), .ZN(u5_mult_79_n933) );
  NAND2_X2 u5_mult_79_U226 ( .A1(u5_mult_79_ab_11__2_), .A2(
        u5_mult_79_CARRYB_10__2_), .ZN(u5_mult_79_n929) );
  BUF_X4 u5_mult_79_U225 ( .A(u5_mult_79_CARRYB_10__3_), .Z(u5_mult_79_n414)
         );
  INV_X32 u5_mult_79_U224 ( .A(u5_mult_79_ab_16__0_), .ZN(u5_mult_79_n90) );
  XNOR2_X2 u5_mult_79_U223 ( .A(u5_mult_79_n90), .B(u5_mult_79_CARRYB_15__0_), 
        .ZN(u5_mult_79_n934) );
  AND2_X2 u5_mult_79_U222 ( .A1(u5_mult_79_SUMB_23__8_), .A2(
        u5_mult_79_CARRYB_23__7_), .ZN(u5_mult_79_n234) );
  NOR2_X1 u5_mult_79_U221 ( .A1(u5_mult_79_n1831), .A2(u5_mult_79_n1728), .ZN(
        u5_mult_79_ab_4__23_) );
  INV_X2 u5_mult_79_U220 ( .A(u5_mult_79_SUMB_5__22_), .ZN(u5_mult_79_n435) );
  INV_X4 u5_mult_79_U219 ( .A(u5_mult_79_n472), .ZN(u5_mult_79_n894) );
  NAND2_X4 u5_mult_79_U218 ( .A1(u5_mult_79_n1554), .A2(u5_mult_79_n894), .ZN(
        u5_mult_79_n895) );
  XNOR2_X2 u5_mult_79_U217 ( .A(u5_mult_79_n1361), .B(u5_mult_79_SUMB_14__16_), 
        .ZN(u5_mult_79_SUMB_15__15_) );
  NAND2_X2 u5_mult_79_U216 ( .A1(u5_mult_79_ab_3__17_), .A2(
        u5_mult_79_SUMB_2__18_), .ZN(u5_mult_79_n592) );
  NAND2_X2 u5_mult_79_U215 ( .A1(u5_mult_79_SUMB_2__18_), .A2(u5_mult_79_n266), 
        .ZN(u5_mult_79_n593) );
  NAND2_X4 u5_mult_79_U214 ( .A1(u5_mult_79_n366), .A2(u5_mult_79_SUMB_13__21_), .ZN(u5_mult_79_n1073) );
  NAND2_X2 u5_mult_79_U213 ( .A1(u5_mult_79_ab_18__17_), .A2(u5_mult_79_n334), 
        .ZN(u5_mult_79_n804) );
  NAND2_X4 u5_mult_79_U212 ( .A1(u5_mult_79_n282), .A2(u5_mult_79_ab_5__21_), 
        .ZN(u5_mult_79_n1552) );
  XNOR2_X2 u5_mult_79_U211 ( .A(u5_mult_79_CARRYB_7__21_), .B(
        u5_mult_79_ab_8__21_), .ZN(u5_mult_79_n263) );
  NAND2_X2 u5_mult_79_U210 ( .A1(u5_mult_79_ab_10__13_), .A2(
        u5_mult_79_CARRYB_9__13_), .ZN(u5_mult_79_n1093) );
  NAND2_X1 u5_mult_79_U209 ( .A1(u5_mult_79_ab_12__15_), .A2(
        u5_mult_79_SUMB_11__16_), .ZN(u5_mult_79_n823) );
  NAND2_X1 u5_mult_79_U208 ( .A1(u5_mult_79_CARRYB_11__15_), .A2(
        u5_mult_79_SUMB_11__16_), .ZN(u5_mult_79_n824) );
  NAND2_X2 u5_mult_79_U207 ( .A1(u5_mult_79_ab_8__15_), .A2(
        u5_mult_79_SUMB_7__16_), .ZN(u5_mult_79_n1399) );
  XNOR2_X2 u5_mult_79_U206 ( .A(u5_mult_79_n398), .B(u5_mult_79_n482), .ZN(
        u5_mult_79_n89) );
  NAND2_X2 u5_mult_79_U205 ( .A1(u5_mult_79_ab_12__12_), .A2(
        u5_mult_79_CARRYB_11__12_), .ZN(u5_mult_79_n1421) );
  NAND2_X4 u5_mult_79_U204 ( .A1(u5_mult_79_CARRYB_2__16_), .A2(
        u5_mult_79_n488), .ZN(u5_mult_79_n1379) );
  NAND2_X2 u5_mult_79_U203 ( .A1(u5_mult_79_SUMB_7__22_), .A2(
        u5_mult_79_CARRYB_7__21_), .ZN(u5_mult_79_n603) );
  NAND3_X4 u5_mult_79_U202 ( .A1(u5_mult_79_n1065), .A2(u5_mult_79_n1066), 
        .A3(u5_mult_79_n1067), .ZN(u5_mult_79_CARRYB_7__21_) );
  NAND2_X4 u5_mult_79_U201 ( .A1(u5_mult_79_ab_8__21_), .A2(
        u5_mult_79_CARRYB_7__21_), .ZN(u5_mult_79_n605) );
  BUF_X8 u5_mult_79_U200 ( .A(u5_mult_79_SUMB_18__13_), .Z(u5_mult_79_n437) );
  XNOR2_X2 u5_mult_79_U199 ( .A(u5_mult_79_CARRYB_22__8_), .B(
        u5_mult_79_ab_23__8_), .ZN(u5_mult_79_n88) );
  XNOR2_X2 u5_mult_79_U198 ( .A(u5_mult_79_SUMB_22__9_), .B(u5_mult_79_n88), 
        .ZN(u5_mult_79_SUMB_23__8_) );
  NAND2_X2 u5_mult_79_U197 ( .A1(u5_mult_79_n277), .A2(u5_mult_79_SUMB_14__7_), 
        .ZN(u5_mult_79_n1000) );
  NAND2_X2 u5_mult_79_U196 ( .A1(u5_mult_79_ab_7__23_), .A2(
        u5_mult_79_CARRYB_7__22_), .ZN(u5_mult_79_n1447) );
  NAND2_X2 u5_mult_79_U195 ( .A1(u5_mult_79_CARRYB_14__14_), .A2(
        u5_mult_79_SUMB_14__15_), .ZN(u5_mult_79_n1334) );
  NAND2_X1 u5_mult_79_U194 ( .A1(u5_mult_79_ab_22__10_), .A2(
        u5_mult_79_CARRYB_21__10_), .ZN(u5_mult_79_n1452) );
  NAND2_X1 u5_mult_79_U193 ( .A1(u5_mult_79_CARRYB_21__10_), .A2(
        u5_mult_79_SUMB_21__11_), .ZN(u5_mult_79_n1454) );
  XOR2_X2 u5_mult_79_U192 ( .A(u5_mult_79_CARRYB_15__6_), .B(
        u5_mult_79_ab_16__6_), .Z(u5_mult_79_n1575) );
  NAND2_X4 u5_mult_79_U191 ( .A1(u5_mult_79_n277), .A2(u5_mult_79_ab_15__6_), 
        .ZN(u5_mult_79_n998) );
  NAND2_X1 u5_mult_79_U190 ( .A1(u5_mult_79_ab_22__11_), .A2(
        u5_mult_79_CARRYB_21__11_), .ZN(u5_mult_79_n1306) );
  NAND2_X1 u5_mult_79_U189 ( .A1(u5_mult_79_SUMB_17__13_), .A2(
        u5_mult_79_ab_18__12_), .ZN(u5_mult_79_n1042) );
  NAND3_X1 u5_mult_79_U188 ( .A1(u5_mult_79_n1454), .A2(u5_mult_79_n1453), 
        .A3(u5_mult_79_n1452), .ZN(u5_mult_79_n213) );
  NAND2_X1 u5_mult_79_U187 ( .A1(u5_mult_79_SUMB_11__17_), .A2(
        u5_mult_79_CARRYB_11__16_), .ZN(u5_mult_79_n743) );
  INV_X4 u5_mult_79_U186 ( .A(u5_mult_79_SUMB_15__13_), .ZN(u5_mult_79_n1133)
         );
  NAND2_X4 u5_mult_79_U185 ( .A1(u5_mult_79_ab_20__10_), .A2(
        u5_mult_79_SUMB_19__11_), .ZN(u5_mult_79_n1428) );
  XOR2_X2 u5_mult_79_U184 ( .A(u5_mult_79_SUMB_12__12_), .B(u5_mult_79_n1084), 
        .Z(u5_mult_79_SUMB_13__11_) );
  NAND3_X4 u5_mult_79_U183 ( .A1(u5_mult_79_n1398), .A2(u5_mult_79_n1399), 
        .A3(u5_mult_79_n1400), .ZN(u5_mult_79_CARRYB_8__15_) );
  NAND2_X2 u5_mult_79_U182 ( .A1(u5_mult_79_CARRYB_4__13_), .A2(
        u5_mult_79_SUMB_4__14_), .ZN(u5_mult_79_n1345) );
  NAND2_X1 u5_mult_79_U181 ( .A1(u5_mult_79_ab_5__13_), .A2(
        u5_mult_79_SUMB_4__14_), .ZN(u5_mult_79_n1344) );
  XOR2_X1 u5_mult_79_U180 ( .A(u5_mult_79_n1339), .B(u5_mult_79_SUMB_4__14_), 
        .Z(u5_mult_79_SUMB_5__13_) );
  CLKBUF_X3 u5_mult_79_U179 ( .A(u5_mult_79_SUMB_9__10_), .Z(u5_mult_79_n308)
         );
  INV_X1 u5_mult_79_U178 ( .A(u5_mult_79_n280), .ZN(u5_mult_79_n474) );
  NAND2_X2 u5_mult_79_U177 ( .A1(u5_mult_79_ab_8__20_), .A2(
        u5_mult_79_SUMB_7__21_), .ZN(u5_mult_79_n170) );
  XNOR2_X2 u5_mult_79_U176 ( .A(u5_mult_79_n4), .B(u5_mult_79_ab_11__20_), 
        .ZN(u5_mult_79_n1118) );
  XNOR2_X2 u5_mult_79_U175 ( .A(u5_mult_79_CARRYB_11__21_), .B(u5_mult_79_n808), .ZN(u5_mult_79_SUMB_12__21_) );
  NAND2_X1 u5_mult_79_U174 ( .A1(u5_mult_79_CARRYB_11__11_), .A2(
        u5_mult_79_SUMB_11__12_), .ZN(u5_mult_79_n1407) );
  NAND2_X1 u5_mult_79_U173 ( .A1(u5_mult_79_ab_12__11_), .A2(
        u5_mult_79_SUMB_11__12_), .ZN(u5_mult_79_n1406) );
  NAND3_X4 u5_mult_79_U172 ( .A1(u5_mult_79_n225), .A2(u5_mult_79_n226), .A3(
        u5_mult_79_n227), .ZN(u5_mult_79_CARRYB_9__19_) );
  NAND2_X2 u5_mult_79_U171 ( .A1(u5_mult_79_CARRYB_8__19_), .A2(
        u5_mult_79_SUMB_8__20_), .ZN(u5_mult_79_n225) );
  INV_X4 u5_mult_79_U170 ( .A(u5_mult_79_n435), .ZN(u5_mult_79_n436) );
  NAND3_X4 u5_mult_79_U169 ( .A1(u5_mult_79_n1418), .A2(u5_mult_79_n1419), 
        .A3(u5_mult_79_n1420), .ZN(u5_mult_79_CARRYB_11__13_) );
  INV_X4 u5_mult_79_U168 ( .A(u5_mult_79_ab_18__13_), .ZN(u5_mult_79_n85) );
  INV_X8 u5_mult_79_U167 ( .A(u5_mult_79_CARRYB_17__13_), .ZN(u5_mult_79_n84)
         );
  NAND2_X4 u5_mult_79_U166 ( .A1(u5_mult_79_n84), .A2(u5_mult_79_n85), .ZN(
        u5_mult_79_n87) );
  NAND2_X2 u5_mult_79_U165 ( .A1(u5_mult_79_CARRYB_17__13_), .A2(
        u5_mult_79_ab_18__13_), .ZN(u5_mult_79_n86) );
  NAND3_X2 u5_mult_79_U164 ( .A1(u5_mult_79_n1220), .A2(u5_mult_79_n1221), 
        .A3(u5_mult_79_n1222), .ZN(u5_mult_79_CARRYB_19__12_) );
  INV_X32 u5_mult_79_U163 ( .A(u5_mult_79_n622), .ZN(u5_mult_79_n83) );
  XNOR2_X2 u5_mult_79_U162 ( .A(u5_mult_79_CARRYB_20__10_), .B(u5_mult_79_n83), 
        .ZN(u5_mult_79_n452) );
  NAND2_X2 u5_mult_79_U161 ( .A1(u5_mult_79_CARRYB_11__7_), .A2(
        u5_mult_79_SUMB_11__8_), .ZN(u5_mult_79_n1094) );
  NAND2_X1 u5_mult_79_U160 ( .A1(u5_mult_79_CARRYB_10__21_), .A2(
        u5_mult_79_SUMB_10__22_), .ZN(u5_mult_79_n1080) );
  NAND2_X1 u5_mult_79_U159 ( .A1(u5_mult_79_CARRYB_10__21_), .A2(
        u5_mult_79_ab_11__21_), .ZN(u5_mult_79_n1081) );
  NAND3_X2 u5_mult_79_U158 ( .A1(u5_mult_79_n80), .A2(u5_mult_79_n81), .A3(
        u5_mult_79_n82), .ZN(u5_mult_79_CARRYB_13__21_) );
  NAND2_X1 u5_mult_79_U157 ( .A1(u5_mult_79_ab_13__21_), .A2(
        u5_mult_79_SUMB_12__22_), .ZN(u5_mult_79_n82) );
  NAND2_X2 u5_mult_79_U156 ( .A1(u5_mult_79_ab_13__21_), .A2(
        u5_mult_79_CARRYB_12__21_), .ZN(u5_mult_79_n81) );
  NAND2_X1 u5_mult_79_U155 ( .A1(u5_mult_79_SUMB_12__22_), .A2(
        u5_mult_79_CARRYB_12__21_), .ZN(u5_mult_79_n80) );
  XOR2_X2 u5_mult_79_U154 ( .A(u5_mult_79_CARRYB_12__21_), .B(u5_mult_79_n79), 
        .Z(u5_mult_79_SUMB_13__21_) );
  XOR2_X2 u5_mult_79_U153 ( .A(u5_mult_79_SUMB_12__22_), .B(
        u5_mult_79_ab_13__21_), .Z(u5_mult_79_n79) );
  NAND2_X2 u5_mult_79_U152 ( .A1(u5_mult_79_ab_4__15_), .A2(
        u5_mult_79_SUMB_3__16_), .ZN(u5_mult_79_n1381) );
  INV_X4 u5_mult_79_U151 ( .A(u5_mult_79_SUMB_3__16_), .ZN(u5_mult_79_n152) );
  XNOR2_X2 u5_mult_79_U150 ( .A(u5_mult_79_SUMB_19__11_), .B(u5_mult_79_n108), 
        .ZN(u5_mult_79_SUMB_20__10_) );
  XNOR2_X1 u5_mult_79_U149 ( .A(u5_mult_79_CARRYB_19__10_), .B(
        u5_mult_79_ab_20__10_), .ZN(u5_mult_79_n108) );
  NAND3_X4 u5_mult_79_U148 ( .A1(u5_mult_79_n1293), .A2(u5_mult_79_n1294), 
        .A3(u5_mult_79_n1295), .ZN(u5_mult_79_CARRYB_9__13_) );
  CLKBUF_X3 u5_mult_79_U147 ( .A(u5_mult_79_CARRYB_18__13_), .Z(
        u5_mult_79_n396) );
  NAND2_X2 u5_mult_79_U146 ( .A1(u5_mult_79_CARRYB_10__10_), .A2(
        u5_mult_79_SUMB_10__11_), .ZN(u5_mult_79_n1464) );
  NAND2_X2 u5_mult_79_U145 ( .A1(u5_mult_79_CARRYB_22__1_), .A2(
        u5_mult_79_SUMB_22__2_), .ZN(u5_mult_79_n508) );
  NAND2_X4 u5_mult_79_U144 ( .A1(u5_mult_79_n1258), .A2(u5_mult_79_n1259), 
        .ZN(u5_mult_79_SUMB_22__2_) );
  NAND2_X2 u5_mult_79_U143 ( .A1(u5_mult_79_SUMB_22__3_), .A2(
        u5_mult_79_CARRYB_22__2_), .ZN(u5_mult_79_n1511) );
  INV_X2 u5_mult_79_U142 ( .A(u5_mult_79_SUMB_15__10_), .ZN(u5_mult_79_n447)
         );
  INV_X4 u5_mult_79_U141 ( .A(u5_mult_79_CARRYB_10__8_), .ZN(u5_mult_79_n405)
         );
  NAND3_X4 u5_mult_79_U140 ( .A1(u5_mult_79_n843), .A2(u5_mult_79_n844), .A3(
        u5_mult_79_n845), .ZN(u5_mult_79_CARRYB_9__8_) );
  NOR2_X4 u5_mult_79_U139 ( .A1(u5_mult_79_n1808), .A2(u5_mult_79_n1746), .ZN(
        u5_mult_79_ab_10__8_) );
  NAND3_X4 u5_mult_79_U138 ( .A1(u5_mult_79_n76), .A2(u5_mult_79_n77), .A3(
        u5_mult_79_n78), .ZN(u5_mult_79_CARRYB_10__8_) );
  NAND2_X4 u5_mult_79_U137 ( .A1(u5_mult_79_ab_10__8_), .A2(
        u5_mult_79_CARRYB_9__8_), .ZN(u5_mult_79_n78) );
  NAND2_X2 u5_mult_79_U136 ( .A1(u5_mult_79_ab_10__8_), .A2(u5_mult_79_n42), 
        .ZN(u5_mult_79_n77) );
  NAND2_X2 u5_mult_79_U135 ( .A1(u5_mult_79_CARRYB_9__8_), .A2(u5_mult_79_n42), 
        .ZN(u5_mult_79_n76) );
  XOR2_X2 u5_mult_79_U134 ( .A(u5_mult_79_n42), .B(u5_mult_79_n75), .Z(
        u5_mult_79_SUMB_10__8_) );
  XOR2_X2 u5_mult_79_U133 ( .A(u5_mult_79_CARRYB_9__8_), .B(
        u5_mult_79_ab_10__8_), .Z(u5_mult_79_n75) );
  NAND2_X2 u5_mult_79_U132 ( .A1(u5_mult_79_SUMB_12__20_), .A2(
        u5_mult_79_CARRYB_12__19_), .ZN(u5_mult_79_n1061) );
  NAND2_X2 u5_mult_79_U131 ( .A1(u5_mult_79_CARRYB_19__11_), .A2(
        u5_mult_79_SUMB_19__12_), .ZN(u5_mult_79_n1225) );
  NAND2_X4 u5_mult_79_U130 ( .A1(u5_mult_79_ab_21__3_), .A2(
        u5_mult_79_CARRYB_20__3_), .ZN(u5_mult_79_n1637) );
  INV_X4 u5_mult_79_U129 ( .A(u5_mult_79_CARRYB_16__8_), .ZN(u5_mult_79_n518)
         );
  NAND2_X2 u5_mult_79_U128 ( .A1(u5_mult_79_CARRYB_9__12_), .A2(
        u5_mult_79_SUMB_9__13_), .ZN(u5_mult_79_n1298) );
  NAND2_X4 u5_mult_79_U127 ( .A1(u5_mult_79_ab_13__10_), .A2(u5_mult_79_n322), 
        .ZN(u5_mult_79_n1410) );
  NAND2_X2 u5_mult_79_U126 ( .A1(u5_mult_79_ab_19__11_), .A2(
        u5_mult_79_SUMB_18__12_), .ZN(u5_mult_79_n1443) );
  XNOR2_X2 u5_mult_79_U125 ( .A(u5_mult_79_n74), .B(u5_mult_79_SUMB_9__21_), 
        .ZN(u5_mult_79_SUMB_10__20_) );
  NAND2_X2 u5_mult_79_U124 ( .A1(u5_mult_79_ab_8__16_), .A2(
        u5_mult_79_CARRYB_7__16_), .ZN(u5_mult_79_n1206) );
  INV_X16 u5_mult_79_U123 ( .A(u5_mult_79_n1864), .ZN(u5_mult_79_n1792) );
  NAND2_X1 u5_mult_79_U122 ( .A1(u5_mult_79_ab_7__15_), .A2(
        u5_mult_79_SUMB_6__16_), .ZN(u5_mult_79_n857) );
  NAND2_X1 u5_mult_79_U121 ( .A1(u5_mult_79_SUMB_6__16_), .A2(
        u5_mult_79_CARRYB_6__15_), .ZN(u5_mult_79_n855) );
  NAND2_X2 u5_mult_79_U120 ( .A1(u5_mult_79_n1525), .A2(u5_mult_79_n454), .ZN(
        u5_mult_79_n1214) );
  NOR2_X2 u5_mult_79_U119 ( .A1(u5_mult_79_n1803), .A2(u5_mult_79_n1773), .ZN(
        u5_mult_79_ab_19__10_) );
  NAND3_X2 u5_mult_79_U118 ( .A1(u5_mult_79_n734), .A2(u5_mult_79_n735), .A3(
        u5_mult_79_n736), .ZN(u5_mult_79_CARRYB_19__9_) );
  NOR2_X4 u5_mult_79_U117 ( .A1(u5_mult_79_n1808), .A2(u5_mult_79_n1859), .ZN(
        u5_mult_79_ab_22__8_) );
  INV_X2 u5_mult_79_U116 ( .A(u5_mult_79_n1305), .ZN(u5_mult_79_n71) );
  INV_X2 u5_mult_79_U115 ( .A(u5_mult_79_n1134), .ZN(u5_mult_79_n70) );
  NAND2_X4 u5_mult_79_U114 ( .A1(u5_mult_79_n72), .A2(u5_mult_79_n73), .ZN(
        u5_mult_79_n454) );
  NAND2_X4 u5_mult_79_U113 ( .A1(u5_mult_79_n70), .A2(u5_mult_79_n71), .ZN(
        u5_mult_79_n73) );
  NAND2_X1 u5_mult_79_U112 ( .A1(u5_mult_79_n1134), .A2(u5_mult_79_n1305), 
        .ZN(u5_mult_79_n72) );
  INV_X2 u5_mult_79_U111 ( .A(u5_mult_79_CARRYB_18__10_), .ZN(u5_mult_79_n67)
         );
  INV_X4 u5_mult_79_U110 ( .A(u5_mult_79_ab_19__10_), .ZN(u5_mult_79_n66) );
  NAND2_X4 u5_mult_79_U109 ( .A1(u5_mult_79_n68), .A2(u5_mult_79_n69), .ZN(
        u5_mult_79_n1246) );
  NAND2_X2 u5_mult_79_U108 ( .A1(u5_mult_79_n66), .A2(u5_mult_79_n67), .ZN(
        u5_mult_79_n69) );
  NAND2_X2 u5_mult_79_U107 ( .A1(u5_mult_79_ab_19__10_), .A2(
        u5_mult_79_CARRYB_18__10_), .ZN(u5_mult_79_n68) );
  XOR2_X2 u5_mult_79_U106 ( .A(u5_mult_79_SUMB_19__10_), .B(u5_mult_79_n65), 
        .Z(u5_mult_79_n367) );
  XOR2_X2 u5_mult_79_U105 ( .A(u5_mult_79_CARRYB_19__9_), .B(
        u5_mult_79_ab_20__9_), .Z(u5_mult_79_n65) );
  INV_X4 u5_mult_79_U104 ( .A(u5_mult_79_CARRYB_21__8_), .ZN(u5_mult_79_n62)
         );
  INV_X16 u5_mult_79_U103 ( .A(u5_mult_79_ab_22__8_), .ZN(u5_mult_79_n61) );
  NAND2_X4 u5_mult_79_U102 ( .A1(u5_mult_79_n63), .A2(u5_mult_79_n64), .ZN(
        u5_mult_79_n260) );
  NAND2_X4 u5_mult_79_U101 ( .A1(u5_mult_79_n61), .A2(u5_mult_79_n62), .ZN(
        u5_mult_79_n64) );
  NAND2_X1 u5_mult_79_U100 ( .A1(u5_mult_79_ab_22__8_), .A2(
        u5_mult_79_CARRYB_21__8_), .ZN(u5_mult_79_n63) );
  NAND2_X1 u5_mult_79_U99 ( .A1(u5_mult_79_CARRYB_8__14_), .A2(
        u5_mult_79_SUMB_8__15_), .ZN(u5_mult_79_n852) );
  INV_X8 u5_mult_79_U98 ( .A(u5_mult_79_n1651), .ZN(u5_mult_79_CLA_SUM[28]) );
  XNOR2_X2 u5_mult_79_U97 ( .A(u5_mult_79_CARRYB_9__20_), .B(
        u5_mult_79_ab_10__20_), .ZN(u5_mult_79_n74) );
  INV_X1 u5_mult_79_U96 ( .A(u5_mult_79_SUMB_13__21_), .ZN(u5_mult_79_n58) );
  INV_X4 u5_mult_79_U95 ( .A(u5_mult_79_n1069), .ZN(u5_mult_79_n57) );
  NAND2_X4 u5_mult_79_U94 ( .A1(u5_mult_79_n59), .A2(u5_mult_79_n60), .ZN(
        u5_mult_79_SUMB_14__20_) );
  NAND2_X2 u5_mult_79_U93 ( .A1(u5_mult_79_n57), .A2(u5_mult_79_SUMB_13__21_), 
        .ZN(u5_mult_79_n60) );
  NAND2_X2 u5_mult_79_U92 ( .A1(u5_mult_79_n1069), .A2(u5_mult_79_n58), .ZN(
        u5_mult_79_n59) );
  NAND3_X4 u5_mult_79_U91 ( .A1(u5_mult_79_n54), .A2(u5_mult_79_n55), .A3(
        u5_mult_79_n56), .ZN(u5_mult_79_CARRYB_20__16_) );
  NAND2_X2 u5_mult_79_U90 ( .A1(u5_mult_79_ab_20__16_), .A2(
        u5_mult_79_SUMB_19__17_), .ZN(u5_mult_79_n56) );
  NAND2_X2 u5_mult_79_U89 ( .A1(u5_mult_79_CARRYB_19__16_), .A2(
        u5_mult_79_SUMB_19__17_), .ZN(u5_mult_79_n55) );
  NAND2_X2 u5_mult_79_U88 ( .A1(u5_mult_79_CARRYB_19__16_), .A2(
        u5_mult_79_ab_20__16_), .ZN(u5_mult_79_n54) );
  NAND3_X2 u5_mult_79_U87 ( .A1(u5_mult_79_n51), .A2(u5_mult_79_n52), .A3(
        u5_mult_79_n53), .ZN(u5_mult_79_CARRYB_19__17_) );
  NAND2_X2 u5_mult_79_U86 ( .A1(u5_mult_79_ab_19__17_), .A2(
        u5_mult_79_SUMB_18__18_), .ZN(u5_mult_79_n53) );
  NAND2_X1 u5_mult_79_U85 ( .A1(u5_mult_79_CARRYB_18__17_), .A2(
        u5_mult_79_SUMB_18__18_), .ZN(u5_mult_79_n52) );
  NAND2_X1 u5_mult_79_U84 ( .A1(u5_mult_79_CARRYB_18__17_), .A2(
        u5_mult_79_ab_19__17_), .ZN(u5_mult_79_n51) );
  XOR2_X2 u5_mult_79_U83 ( .A(u5_mult_79_n50), .B(u5_mult_79_SUMB_19__17_), 
        .Z(u5_mult_79_SUMB_20__16_) );
  XOR2_X2 u5_mult_79_U82 ( .A(u5_mult_79_CARRYB_19__16_), .B(
        u5_mult_79_ab_20__16_), .Z(u5_mult_79_n50) );
  XOR2_X2 u5_mult_79_U81 ( .A(u5_mult_79_n49), .B(u5_mult_79_SUMB_18__18_), 
        .Z(u5_mult_79_SUMB_19__17_) );
  XOR2_X2 u5_mult_79_U80 ( .A(u5_mult_79_CARRYB_18__17_), .B(
        u5_mult_79_ab_19__17_), .Z(u5_mult_79_n49) );
  NAND2_X2 u5_mult_79_U79 ( .A1(u5_mult_79_ab_20__11_), .A2(
        u5_mult_79_SUMB_19__12_), .ZN(u5_mult_79_n1224) );
  NAND2_X4 u5_mult_79_U78 ( .A1(u5_mult_79_ab_21__3_), .A2(
        u5_mult_79_SUMB_20__4_), .ZN(u5_mult_79_n1636) );
  NAND3_X2 u5_mult_79_U77 ( .A1(u5_mult_79_n1000), .A2(u5_mult_79_n999), .A3(
        u5_mult_79_n998), .ZN(u5_mult_79_CARRYB_15__6_) );
  NAND2_X2 u5_mult_79_U76 ( .A1(u5_mult_79_n1257), .A2(u5_mult_79_n280), .ZN(
        u5_mult_79_n1259) );
  INV_X8 u5_mult_79_U75 ( .A(u5_mult_79_n1646), .ZN(u5_mult_79_CLA_CARRY[25])
         );
  INV_X2 u5_mult_79_U74 ( .A(u5_mult_79_n47), .ZN(u5_mult_79_n48) );
  INV_X1 u5_mult_79_U73 ( .A(u5_mult_79_CARRYB_11__8_), .ZN(u5_mult_79_n47) );
  INV_X4 u5_mult_79_U72 ( .A(u5_mult_79_CARRYB_6__20_), .ZN(u5_mult_79_n625)
         );
  NAND2_X4 u5_mult_79_U71 ( .A1(u5_mult_79_n625), .A2(u5_mult_79_n624), .ZN(
        u5_mult_79_n626) );
  NAND2_X4 u5_mult_79_U70 ( .A1(u5_mult_79_n1229), .A2(u5_mult_79_n626), .ZN(
        u5_mult_79_n1119) );
  NAND3_X1 u5_mult_79_U69 ( .A1(u5_mult_79_n1229), .A2(u5_mult_79_n1230), .A3(
        u5_mult_79_n1231), .ZN(u5_mult_79_CARRYB_7__20_) );
  BUF_X4 u5_mult_79_U68 ( .A(u5_mult_79_n1720), .Z(u5_mult_79_n46) );
  INV_X4 u5_mult_79_U67 ( .A(u5_mult_79_n44), .ZN(u5_mult_79_n45) );
  INV_X2 u5_mult_79_U66 ( .A(u5_mult_79_SUMB_10__14_), .ZN(u5_mult_79_n44) );
  XOR2_X2 u5_mult_79_U65 ( .A(u5_mult_79_n469), .B(u5_mult_79_CARRYB_21__11_), 
        .Z(u5_mult_79_n43) );
  XNOR2_X2 u5_mult_79_U64 ( .A(u5_mult_79_SUMB_21__12_), .B(u5_mult_79_n43), 
        .ZN(u5_mult_79_SUMB_22__11_) );
  INV_X8 u5_mult_79_U63 ( .A(u5_mult_79_n41), .ZN(u5_mult_79_n42) );
  INV_X4 u5_mult_79_U62 ( .A(u5_mult_79_SUMB_9__9_), .ZN(u5_mult_79_n41) );
  INV_X4 u5_mult_79_U61 ( .A(u5_mult_79_n39), .ZN(u5_mult_79_n40) );
  INV_X2 u5_mult_79_U60 ( .A(u5_mult_79_SUMB_16__14_), .ZN(u5_mult_79_n39) );
  CLKBUF_X3 u5_mult_79_U59 ( .A(u5_mult_79_SUMB_12__17_), .Z(u5_mult_79_n38)
         );
  CLKBUF_X3 u5_mult_79_U58 ( .A(u5_mult_79_SUMB_15__14_), .Z(u5_mult_79_n37)
         );
  NAND3_X2 u5_mult_79_U57 ( .A1(u5_mult_79_n1582), .A2(u5_mult_79_n1583), .A3(
        u5_mult_79_n1584), .ZN(u5_mult_79_CARRYB_5__17_) );
  CLKBUF_X3 u5_mult_79_U56 ( .A(u5_mult_79_CARRYB_7__20_), .Z(u5_mult_79_n36)
         );
  XNOR2_X1 u5_mult_79_U55 ( .A(u5_mult_79_n445), .B(u5_mult_79_SUMB_17__12_), 
        .ZN(u5_mult_79_n300) );
  NAND2_X1 u5_mult_79_U54 ( .A1(u5_mult_79_CARRYB_6__12_), .A2(
        u5_mult_79_SUMB_6__13_), .ZN(u5_mult_79_n702) );
  NAND2_X1 u5_mult_79_U53 ( .A1(u5_mult_79_ab_7__12_), .A2(
        u5_mult_79_SUMB_6__13_), .ZN(u5_mult_79_n703) );
  CLKBUF_X3 u5_mult_79_U52 ( .A(u5_mult_79_SUMB_10__12_), .Z(u5_mult_79_n35)
         );
  INV_X4 u5_mult_79_U51 ( .A(u5_mult_79_n33), .ZN(u5_mult_79_n34) );
  INV_X2 u5_mult_79_U50 ( .A(u5_mult_79_SUMB_5__17_), .ZN(u5_mult_79_n33) );
  XNOR2_X2 u5_mult_79_U49 ( .A(u5_mult_79_CARRYB_12__4_), .B(
        u5_mult_79_ab_13__4_), .ZN(u5_mult_79_n256) );
  XNOR2_X2 u5_mult_79_U48 ( .A(u5_mult_79_n30), .B(u5_mult_79_n687), .ZN(
        u5_mult_79_n32) );
  XNOR2_X1 u5_mult_79_U47 ( .A(u5_mult_79_ab_20__13_), .B(
        u5_mult_79_CARRYB_19__13_), .ZN(u5_mult_79_n31) );
  XNOR2_X2 u5_mult_79_U46 ( .A(u5_mult_79_n31), .B(u5_mult_79_n5), .ZN(
        u5_mult_79_SUMB_20__13_) );
  CLKBUF_X3 u5_mult_79_U45 ( .A(u5_mult_79_SUMB_6__15_), .Z(u5_mult_79_n30) );
  CLKBUF_X3 u5_mult_79_U44 ( .A(u5_mult_79_SUMB_8__15_), .Z(u5_mult_79_n29) );
  XNOR2_X2 u5_mult_79_U43 ( .A(u5_mult_79_n379), .B(u5_mult_79_n395), .ZN(
        u5_mult_79_n28) );
  INV_X4 u5_mult_79_U42 ( .A(u5_mult_79_n26), .ZN(u5_mult_79_n27) );
  INV_X2 u5_mult_79_U41 ( .A(u5_mult_79_CARRYB_6__13_), .ZN(u5_mult_79_n26) );
  XNOR2_X2 u5_mult_79_U40 ( .A(u5_mult_79_ab_11__7_), .B(
        u5_mult_79_CARRYB_10__7_), .ZN(u5_mult_79_n25) );
  XNOR2_X2 u5_mult_79_U39 ( .A(u5_mult_79_n25), .B(u5_mult_79_n358), .ZN(
        u5_mult_79_SUMB_11__7_) );
  CLKBUF_X2 u5_mult_79_U38 ( .A(u5_mult_79_SUMB_8__14_), .Z(u5_mult_79_n24) );
  INV_X4 u5_mult_79_U37 ( .A(u5_mult_79_n22), .ZN(u5_mult_79_n23) );
  INV_X2 u5_mult_79_U36 ( .A(u5_mult_79_SUMB_15__17_), .ZN(u5_mult_79_n22) );
  CLKBUF_X2 u5_mult_79_U35 ( .A(u5_mult_79_SUMB_7__18_), .Z(u5_mult_79_n21) );
  INV_X4 u5_mult_79_U34 ( .A(u5_mult_79_n19), .ZN(u5_mult_79_n20) );
  INV_X2 u5_mult_79_U33 ( .A(u5_mult_79_SUMB_15__9_), .ZN(u5_mult_79_n19) );
  XNOR2_X2 u5_mult_79_U32 ( .A(u5_mult_79_CARRYB_16__2_), .B(
        u5_mult_79_ab_17__2_), .ZN(u5_mult_79_n846) );
  XNOR2_X2 u5_mult_79_U31 ( .A(u5_mult_79_ab_21__15_), .B(
        u5_mult_79_CARRYB_20__15_), .ZN(u5_mult_79_n18) );
  XNOR2_X2 u5_mult_79_U30 ( .A(u5_mult_79_n18), .B(u5_mult_79_SUMB_20__16_), 
        .ZN(u5_mult_79_SUMB_21__15_) );
  CLKBUF_X2 u5_mult_79_U29 ( .A(u5_mult_79_SUMB_19__15_), .Z(u5_mult_79_n17)
         );
  INV_X4 u5_mult_79_U28 ( .A(u5_mult_79_SUMB_19__12_), .ZN(u5_mult_79_n16) );
  XNOR2_X2 u5_mult_79_U27 ( .A(u5_mult_79_n1149), .B(u5_mult_79_CARRYB_19__11_), .ZN(u5_mult_79_n15) );
  XNOR2_X2 u5_mult_79_U26 ( .A(u5_mult_79_n15), .B(u5_mult_79_n16), .ZN(
        u5_mult_79_SUMB_20__11_) );
  BUF_X8 u5_mult_79_U25 ( .A(u5_mult_79_SUMB_20__8_), .Z(u5_mult_79_n374) );
  AND2_X2 u5_mult_79_U24 ( .A1(u5_mult_79_SUMB_23__6_), .A2(
        u5_mult_79_CARRYB_23__5_), .ZN(u5_mult_79_n233) );
  NAND2_X4 u5_mult_79_U23 ( .A1(u5_mult_79_n1241), .A2(u5_mult_79_n1242), .ZN(
        u5_mult_79_n1331) );
  XNOR2_X2 u5_mult_79_U22 ( .A(u5_mult_79_n1331), .B(u5_mult_79_SUMB_14__13_), 
        .ZN(u5_mult_79_n14) );
  XNOR2_X1 u5_mult_79_U21 ( .A(u5_mult_79_CARRYB_19__3_), .B(
        u5_mult_79_ab_20__3_), .ZN(u5_mult_79_n1300) );
  NAND2_X1 u5_mult_79_U20 ( .A1(u5_mult_79_CARRYB_19__3_), .A2(
        u5_mult_79_ab_20__3_), .ZN(u5_mult_79_n1634) );
  XNOR2_X2 u5_mult_79_U19 ( .A(u5_mult_79_CARRYB_15__15_), .B(
        u5_mult_79_ab_16__15_), .ZN(u5_mult_79_n13) );
  XNOR2_X2 u5_mult_79_U18 ( .A(u5_mult_79_n13), .B(u5_mult_79_SUMB_15__16_), 
        .ZN(u5_mult_79_SUMB_16__15_) );
  INV_X2 u5_mult_79_U17 ( .A(u5_mult_79_n11), .ZN(u5_mult_79_n12) );
  INV_X1 u5_mult_79_U16 ( .A(u5_mult_79_SUMB_7__13_), .ZN(u5_mult_79_n11) );
  CLKBUF_X2 u5_mult_79_U15 ( .A(u5_mult_79_CARRYB_6__8_), .Z(u5_mult_79_n10)
         );
  NAND3_X4 u5_mult_79_U14 ( .A1(u5_mult_79_n1323), .A2(u5_mult_79_n1322), .A3(
        u5_mult_79_n1321), .ZN(u5_mult_79_CARRYB_16__8_) );
  NAND2_X2 u5_mult_79_U13 ( .A1(u5_mult_79_ab_17__8_), .A2(
        u5_mult_79_CARRYB_16__8_), .ZN(u5_mult_79_n1610) );
  CLKBUF_X2 u5_mult_79_U12 ( .A(u5_mult_79_CARRYB_4__12_), .Z(u5_mult_79_n9)
         );
  INV_X2 u5_mult_79_U11 ( .A(u5_mult_79_n7), .ZN(u5_mult_79_n8) );
  INV_X1 u5_mult_79_U10 ( .A(u5_mult_79_SUMB_9__14_), .ZN(u5_mult_79_n7) );
  INV_X1 u5_mult_79_U9 ( .A(u5_mult_79_SUMB_9__6_), .ZN(u5_mult_79_n114) );
  NAND2_X4 u5_mult_79_U8 ( .A1(u5_mult_79_n86), .A2(u5_mult_79_n87), .ZN(
        u5_mult_79_n633) );
  XNOR2_X2 u5_mult_79_U7 ( .A(u5_mult_79_CARRYB_16__13_), .B(
        u5_mult_79_ab_17__13_), .ZN(u5_mult_79_n6) );
  XNOR2_X2 u5_mult_79_U6 ( .A(u5_mult_79_n40), .B(u5_mult_79_n6), .ZN(
        u5_mult_79_SUMB_17__13_) );
  NAND2_X1 u5_mult_79_U5 ( .A1(u5_mult_79_CARRYB_12__18_), .A2(
        u5_mult_79_SUMB_12__19_), .ZN(u5_mult_79_n1235) );
  CLKBUF_X2 u5_mult_79_U4 ( .A(u5_mult_79_SUMB_19__14_), .Z(u5_mult_79_n5) );
  INV_X4 u5_mult_79_U3 ( .A(u5_mult_79_n3), .ZN(u5_mult_79_n4) );
  INV_X2 u5_mult_79_U2 ( .A(u5_mult_79_SUMB_10__21_), .ZN(u5_mult_79_n3) );
  FA_X1 u5_mult_79_S3_2_22 ( .A(u5_mult_79_ab_2__22_), .B(
        u5_mult_79_CARRYB_1__22_), .CI(u5_mult_79_ab_1__23_), .CO(
        u5_mult_79_CARRYB_2__22_), .S(u5_mult_79_SUMB_2__22_) );
  FA_X1 u5_mult_79_S2_2_20 ( .A(u5_mult_79_ab_2__20_), .B(
        u5_mult_79_CARRYB_1__20_), .CI(u5_mult_79_SUMB_1__21_), .CO(
        u5_mult_79_CARRYB_2__20_), .S(u5_mult_79_SUMB_2__20_) );
  FA_X1 u5_mult_79_S2_2_19 ( .A(u5_mult_79_ab_2__19_), .B(
        u5_mult_79_CARRYB_1__19_), .CI(u5_mult_79_SUMB_1__20_), .CO(
        u5_mult_79_CARRYB_2__19_), .S(u5_mult_79_SUMB_2__19_) );
  FA_X1 u5_mult_79_S2_2_17 ( .A(u5_mult_79_n239), .B(u5_mult_79_ab_2__17_), 
        .CI(u5_mult_79_SUMB_1__18_), .CO(u5_mult_79_CARRYB_2__17_), .S(
        u5_mult_79_SUMB_2__17_) );
  FA_X1 u5_mult_79_S2_2_13 ( .A(u5_mult_79_ab_2__13_), .B(
        u5_mult_79_CARRYB_1__13_), .CI(u5_mult_79_SUMB_1__14_), .CO(
        u5_mult_79_CARRYB_2__13_), .S(u5_mult_79_SUMB_2__13_) );
  FA_X1 u5_mult_79_S2_2_11 ( .A(u5_mult_79_ab_2__11_), .B(
        u5_mult_79_CARRYB_1__11_), .CI(u5_mult_79_SUMB_1__12_), .CO(
        u5_mult_79_CARRYB_2__11_), .S(u5_mult_79_SUMB_2__11_) );
  FA_X1 u5_mult_79_S2_2_10 ( .A(u5_mult_79_ab_2__10_), .B(
        u5_mult_79_CARRYB_1__10_), .CI(u5_mult_79_SUMB_1__11_), .CO(
        u5_mult_79_CARRYB_2__10_), .S(u5_mult_79_SUMB_2__10_) );
  FA_X1 u5_mult_79_S2_2_9 ( .A(u5_mult_79_ab_2__9_), .B(u5_mult_79_n240), .CI(
        u5_mult_79_SUMB_1__10_), .CO(u5_mult_79_CARRYB_2__9_), .S(
        u5_mult_79_SUMB_2__9_) );
  FA_X1 u5_mult_79_S2_2_8 ( .A(u5_mult_79_ab_2__8_), .B(
        u5_mult_79_CARRYB_1__8_), .CI(u5_mult_79_SUMB_1__9_), .CO(
        u5_mult_79_CARRYB_2__8_), .S(u5_mult_79_SUMB_2__8_) );
  FA_X1 u5_mult_79_S2_2_7 ( .A(u5_mult_79_ab_2__7_), .B(
        u5_mult_79_CARRYB_1__7_), .CI(u5_mult_79_SUMB_1__8_), .CO(
        u5_mult_79_CARRYB_2__7_), .S(u5_mult_79_SUMB_2__7_) );
  FA_X1 u5_mult_79_S2_2_6 ( .A(u5_mult_79_ab_2__6_), .B(
        u5_mult_79_CARRYB_1__6_), .CI(u5_mult_79_SUMB_1__7_), .CO(
        u5_mult_79_CARRYB_2__6_), .S(u5_mult_79_SUMB_2__6_) );
  FA_X1 u5_mult_79_S2_2_5 ( .A(u5_mult_79_ab_2__5_), .B(
        u5_mult_79_CARRYB_1__5_), .CI(u5_mult_79_SUMB_1__6_), .CO(
        u5_mult_79_CARRYB_2__5_), .S(u5_mult_79_SUMB_2__5_) );
  FA_X1 u5_mult_79_S2_2_4 ( .A(u5_mult_79_ab_2__4_), .B(
        u5_mult_79_CARRYB_1__4_), .CI(u5_mult_79_SUMB_1__5_), .CO(
        u5_mult_79_CARRYB_2__4_), .S(u5_mult_79_SUMB_2__4_) );
  FA_X1 u5_mult_79_S2_2_3 ( .A(u5_mult_79_ab_2__3_), .B(
        u5_mult_79_CARRYB_1__3_), .CI(u5_mult_79_SUMB_1__4_), .CO(
        u5_mult_79_CARRYB_2__3_), .S(u5_mult_79_SUMB_2__3_) );
  FA_X1 u5_mult_79_S2_2_2 ( .A(u5_mult_79_ab_2__2_), .B(
        u5_mult_79_CARRYB_1__2_), .CI(u5_mult_79_SUMB_1__3_), .CO(
        u5_mult_79_CARRYB_2__2_), .S(u5_mult_79_SUMB_2__2_) );
  FA_X1 u5_mult_79_S2_2_1 ( .A(u5_mult_79_ab_2__1_), .B(
        u5_mult_79_CARRYB_1__1_), .CI(u5_mult_79_SUMB_1__2_), .CO(
        u5_mult_79_CARRYB_2__1_), .S(u5_mult_79_SUMB_2__1_) );
  FA_X1 u5_mult_79_S1_2_0 ( .A(u5_mult_79_ab_2__0_), .B(
        u5_mult_79_CARRYB_1__0_), .CI(u5_mult_79_SUMB_1__1_), .CO(
        u5_mult_79_CARRYB_2__0_), .S(u5_N2) );
  FA_X1 u5_mult_79_S2_3_19 ( .A(u5_mult_79_ab_3__19_), .B(
        u5_mult_79_CARRYB_2__19_), .CI(u5_mult_79_SUMB_2__20_), .CO(
        u5_mult_79_CARRYB_3__19_), .S(u5_mult_79_SUMB_3__19_) );
  FA_X1 u5_mult_79_S2_3_10 ( .A(u5_mult_79_CARRYB_2__10_), .B(
        u5_mult_79_ab_3__10_), .CI(u5_mult_79_SUMB_2__11_), .CO(
        u5_mult_79_CARRYB_3__10_), .S(u5_mult_79_SUMB_3__10_) );
  FA_X1 u5_mult_79_S2_3_9 ( .A(u5_mult_79_ab_3__9_), .B(
        u5_mult_79_CARRYB_2__9_), .CI(u5_mult_79_SUMB_2__10_), .CO(
        u5_mult_79_CARRYB_3__9_), .S(u5_mult_79_SUMB_3__9_) );
  FA_X1 u5_mult_79_S2_3_8 ( .A(u5_mult_79_ab_3__8_), .B(
        u5_mult_79_CARRYB_2__8_), .CI(u5_mult_79_SUMB_2__9_), .CO(
        u5_mult_79_CARRYB_3__8_), .S(u5_mult_79_SUMB_3__8_) );
  FA_X1 u5_mult_79_S2_3_7 ( .A(u5_mult_79_ab_3__7_), .B(
        u5_mult_79_CARRYB_2__7_), .CI(u5_mult_79_SUMB_2__8_), .CO(
        u5_mult_79_CARRYB_3__7_), .S(u5_mult_79_SUMB_3__7_) );
  FA_X1 u5_mult_79_S2_3_6 ( .A(u5_mult_79_ab_3__6_), .B(
        u5_mult_79_CARRYB_2__6_), .CI(u5_mult_79_SUMB_2__7_), .CO(
        u5_mult_79_CARRYB_3__6_), .S(u5_mult_79_SUMB_3__6_) );
  FA_X1 u5_mult_79_S2_3_5 ( .A(u5_mult_79_ab_3__5_), .B(
        u5_mult_79_CARRYB_2__5_), .CI(u5_mult_79_SUMB_2__6_), .CO(
        u5_mult_79_CARRYB_3__5_), .S(u5_mult_79_SUMB_3__5_) );
  FA_X1 u5_mult_79_S2_3_4 ( .A(u5_mult_79_ab_3__4_), .B(
        u5_mult_79_CARRYB_2__4_), .CI(u5_mult_79_SUMB_2__5_), .CO(
        u5_mult_79_CARRYB_3__4_), .S(u5_mult_79_SUMB_3__4_) );
  FA_X1 u5_mult_79_S2_3_3 ( .A(u5_mult_79_ab_3__3_), .B(
        u5_mult_79_CARRYB_2__3_), .CI(u5_mult_79_SUMB_2__4_), .CO(
        u5_mult_79_CARRYB_3__3_), .S(u5_mult_79_SUMB_3__3_) );
  FA_X1 u5_mult_79_S2_3_2 ( .A(u5_mult_79_ab_3__2_), .B(
        u5_mult_79_CARRYB_2__2_), .CI(u5_mult_79_SUMB_2__3_), .CO(
        u5_mult_79_CARRYB_3__2_), .S(u5_mult_79_SUMB_3__2_) );
  FA_X1 u5_mult_79_S2_3_1 ( .A(u5_mult_79_ab_3__1_), .B(
        u5_mult_79_CARRYB_2__1_), .CI(u5_mult_79_SUMB_2__2_), .CO(
        u5_mult_79_CARRYB_3__1_), .S(u5_mult_79_SUMB_3__1_) );
  FA_X1 u5_mult_79_S1_3_0 ( .A(u5_mult_79_ab_3__0_), .B(
        u5_mult_79_CARRYB_2__0_), .CI(u5_mult_79_SUMB_2__1_), .CO(
        u5_mult_79_CARRYB_3__0_), .S(u5_N3) );
  FA_X1 u5_mult_79_S3_4_22 ( .A(u5_mult_79_ab_4__22_), .B(u5_mult_79_ab_3__23_), .CI(u5_mult_79_CARRYB_3__22_), .CO(u5_mult_79_CARRYB_4__22_), .S(
        u5_mult_79_SUMB_4__22_) );
  FA_X1 u5_mult_79_S2_4_12 ( .A(u5_mult_79_CARRYB_3__12_), .B(
        u5_mult_79_ab_4__12_), .CI(u5_mult_79_SUMB_3__13_), .CO(
        u5_mult_79_CARRYB_4__12_), .S(u5_mult_79_SUMB_4__12_) );
  FA_X1 u5_mult_79_S2_4_10 ( .A(u5_mult_79_CARRYB_3__10_), .B(
        u5_mult_79_ab_4__10_), .CI(u5_mult_79_SUMB_3__11_), .CO(
        u5_mult_79_CARRYB_4__10_), .S(u5_mult_79_SUMB_4__10_) );
  FA_X1 u5_mult_79_S2_4_9 ( .A(u5_mult_79_ab_4__9_), .B(
        u5_mult_79_CARRYB_3__9_), .CI(u5_mult_79_SUMB_3__10_), .CO(
        u5_mult_79_CARRYB_4__9_), .S(u5_mult_79_SUMB_4__9_) );
  FA_X1 u5_mult_79_S2_4_8 ( .A(u5_mult_79_ab_4__8_), .B(
        u5_mult_79_CARRYB_3__8_), .CI(u5_mult_79_SUMB_3__9_), .CO(
        u5_mult_79_CARRYB_4__8_), .S(u5_mult_79_SUMB_4__8_) );
  FA_X1 u5_mult_79_S2_4_7 ( .A(u5_mult_79_ab_4__7_), .B(
        u5_mult_79_CARRYB_3__7_), .CI(u5_mult_79_SUMB_3__8_), .CO(
        u5_mult_79_CARRYB_4__7_), .S(u5_mult_79_SUMB_4__7_) );
  FA_X1 u5_mult_79_S2_4_6 ( .A(u5_mult_79_CARRYB_3__6_), .B(
        u5_mult_79_ab_4__6_), .CI(u5_mult_79_SUMB_3__7_), .CO(
        u5_mult_79_CARRYB_4__6_), .S(u5_mult_79_SUMB_4__6_) );
  FA_X1 u5_mult_79_S2_4_5 ( .A(u5_mult_79_ab_4__5_), .B(
        u5_mult_79_CARRYB_3__5_), .CI(u5_mult_79_SUMB_3__6_), .CO(
        u5_mult_79_CARRYB_4__5_), .S(u5_mult_79_SUMB_4__5_) );
  FA_X1 u5_mult_79_S2_4_4 ( .A(u5_mult_79_ab_4__4_), .B(
        u5_mult_79_CARRYB_3__4_), .CI(u5_mult_79_SUMB_3__5_), .CO(
        u5_mult_79_CARRYB_4__4_), .S(u5_mult_79_SUMB_4__4_) );
  FA_X1 u5_mult_79_S2_4_3 ( .A(u5_mult_79_ab_4__3_), .B(
        u5_mult_79_CARRYB_3__3_), .CI(u5_mult_79_SUMB_3__4_), .CO(
        u5_mult_79_CARRYB_4__3_), .S(u5_mult_79_SUMB_4__3_) );
  FA_X1 u5_mult_79_S2_4_2 ( .A(u5_mult_79_ab_4__2_), .B(
        u5_mult_79_CARRYB_3__2_), .CI(u5_mult_79_SUMB_3__3_), .CO(
        u5_mult_79_CARRYB_4__2_), .S(u5_mult_79_SUMB_4__2_) );
  FA_X1 u5_mult_79_S2_4_1 ( .A(u5_mult_79_ab_4__1_), .B(
        u5_mult_79_CARRYB_3__1_), .CI(u5_mult_79_SUMB_3__2_), .CO(
        u5_mult_79_CARRYB_4__1_), .S(u5_mult_79_SUMB_4__1_) );
  FA_X1 u5_mult_79_S1_4_0 ( .A(u5_mult_79_ab_4__0_), .B(
        u5_mult_79_CARRYB_3__0_), .CI(u5_mult_79_SUMB_3__1_), .CO(
        u5_mult_79_CARRYB_4__0_), .S(u5_N4) );
  FA_X1 u5_mult_79_S3_5_22 ( .A(u5_mult_79_ab_5__22_), .B(u5_mult_79_ab_4__23_), .CI(u5_mult_79_CARRYB_4__22_), .CO(u5_mult_79_CARRYB_5__22_), .S(
        u5_mult_79_SUMB_5__22_) );
  FA_X1 u5_mult_79_S2_5_15 ( .A(u5_mult_79_ab_5__15_), .B(
        u5_mult_79_CARRYB_4__15_), .CI(u5_mult_79_SUMB_4__16_), .CO(
        u5_mult_79_CARRYB_5__15_), .S(u5_mult_79_SUMB_5__15_) );
  FA_X1 u5_mult_79_S2_5_14 ( .A(u5_mult_79_CARRYB_4__14_), .B(
        u5_mult_79_ab_5__14_), .CI(u5_mult_79_SUMB_4__15_), .CO(
        u5_mult_79_CARRYB_5__14_), .S(u5_mult_79_SUMB_5__14_) );
  FA_X1 u5_mult_79_S2_5_9 ( .A(u5_mult_79_CARRYB_4__9_), .B(
        u5_mult_79_ab_5__9_), .CI(u5_mult_79_SUMB_4__10_), .CO(
        u5_mult_79_CARRYB_5__9_), .S(u5_mult_79_SUMB_5__9_) );
  FA_X1 u5_mult_79_S2_5_8 ( .A(u5_mult_79_ab_5__8_), .B(
        u5_mult_79_CARRYB_4__8_), .CI(u5_mult_79_SUMB_4__9_), .CO(
        u5_mult_79_CARRYB_5__8_), .S(u5_mult_79_SUMB_5__8_) );
  FA_X1 u5_mult_79_S2_5_4 ( .A(u5_mult_79_ab_5__4_), .B(
        u5_mult_79_CARRYB_4__4_), .CI(u5_mult_79_SUMB_4__5_), .CO(
        u5_mult_79_CARRYB_5__4_), .S(u5_mult_79_SUMB_5__4_) );
  FA_X1 u5_mult_79_S2_5_3 ( .A(u5_mult_79_ab_5__3_), .B(
        u5_mult_79_CARRYB_4__3_), .CI(u5_mult_79_SUMB_4__4_), .CO(
        u5_mult_79_CARRYB_5__3_), .S(u5_mult_79_SUMB_5__3_) );
  FA_X1 u5_mult_79_S2_5_2 ( .A(u5_mult_79_ab_5__2_), .B(
        u5_mult_79_CARRYB_4__2_), .CI(u5_mult_79_SUMB_4__3_), .CO(
        u5_mult_79_CARRYB_5__2_), .S(u5_mult_79_SUMB_5__2_) );
  FA_X1 u5_mult_79_S2_5_1 ( .A(u5_mult_79_ab_5__1_), .B(
        u5_mult_79_CARRYB_4__1_), .CI(u5_mult_79_SUMB_4__2_), .CO(
        u5_mult_79_CARRYB_5__1_), .S(u5_mult_79_SUMB_5__1_) );
  FA_X1 u5_mult_79_S1_5_0 ( .A(u5_mult_79_ab_5__0_), .B(
        u5_mult_79_CARRYB_4__0_), .CI(u5_mult_79_SUMB_4__1_), .CO(
        u5_mult_79_CARRYB_5__0_), .S(u5_N5) );
  FA_X1 u5_mult_79_S2_6_13 ( .A(u5_mult_79_ab_6__13_), .B(
        u5_mult_79_CARRYB_5__13_), .CI(u5_mult_79_SUMB_5__14_), .CO(
        u5_mult_79_CARRYB_6__13_), .S(u5_mult_79_SUMB_6__13_) );
  FA_X1 u5_mult_79_S2_6_8 ( .A(u5_mult_79_CARRYB_5__8_), .B(
        u5_mult_79_ab_6__8_), .CI(u5_mult_79_SUMB_5__9_), .CO(
        u5_mult_79_CARRYB_6__8_), .S(u5_mult_79_SUMB_6__8_) );
  FA_X1 u5_mult_79_S2_6_5 ( .A(u5_mult_79_ab_6__5_), .B(
        u5_mult_79_CARRYB_5__5_), .CI(u5_mult_79_SUMB_5__6_), .CO(
        u5_mult_79_CARRYB_6__5_), .S(u5_mult_79_SUMB_6__5_) );
  FA_X1 u5_mult_79_S2_6_3 ( .A(u5_mult_79_ab_6__3_), .B(
        u5_mult_79_CARRYB_5__3_), .CI(u5_mult_79_SUMB_5__4_), .CO(
        u5_mult_79_CARRYB_6__3_), .S(u5_mult_79_SUMB_6__3_) );
  FA_X1 u5_mult_79_S2_6_2 ( .A(u5_mult_79_ab_6__2_), .B(
        u5_mult_79_CARRYB_5__2_), .CI(u5_mult_79_SUMB_5__3_), .CO(
        u5_mult_79_CARRYB_6__2_), .S(u5_mult_79_SUMB_6__2_) );
  FA_X1 u5_mult_79_S2_6_1 ( .A(u5_mult_79_ab_6__1_), .B(
        u5_mult_79_CARRYB_5__1_), .CI(u5_mult_79_SUMB_5__2_), .CO(
        u5_mult_79_CARRYB_6__1_), .S(u5_mult_79_SUMB_6__1_) );
  FA_X1 u5_mult_79_S1_6_0 ( .A(u5_mult_79_ab_6__0_), .B(
        u5_mult_79_CARRYB_5__0_), .CI(u5_mult_79_SUMB_5__1_), .CO(
        u5_mult_79_CARRYB_6__0_), .S(u5_N6) );
  FA_X1 u5_mult_79_S2_7_5 ( .A(u5_mult_79_CARRYB_6__5_), .B(
        u5_mult_79_ab_7__5_), .CI(u5_mult_79_SUMB_6__6_), .CO(
        u5_mult_79_CARRYB_7__5_), .S(u5_mult_79_SUMB_7__5_) );
  FA_X1 u5_mult_79_S2_7_4 ( .A(u5_mult_79_ab_7__4_), .B(
        u5_mult_79_CARRYB_6__4_), .CI(u5_mult_79_SUMB_6__5_), .CO(
        u5_mult_79_CARRYB_7__4_), .S(u5_mult_79_SUMB_7__4_) );
  FA_X1 u5_mult_79_S2_7_2 ( .A(u5_mult_79_ab_7__2_), .B(
        u5_mult_79_CARRYB_6__2_), .CI(u5_mult_79_SUMB_6__3_), .CO(
        u5_mult_79_CARRYB_7__2_), .S(u5_mult_79_SUMB_7__2_) );
  FA_X1 u5_mult_79_S2_7_1 ( .A(u5_mult_79_ab_7__1_), .B(
        u5_mult_79_CARRYB_6__1_), .CI(u5_mult_79_SUMB_6__2_), .CO(
        u5_mult_79_CARRYB_7__1_), .S(u5_mult_79_SUMB_7__1_) );
  FA_X1 u5_mult_79_S1_7_0 ( .A(u5_mult_79_ab_7__0_), .B(
        u5_mult_79_CARRYB_6__0_), .CI(u5_mult_79_SUMB_6__1_), .CO(
        u5_mult_79_CARRYB_7__0_), .S(u5_N7) );
  FA_X1 u5_mult_79_S2_8_19 ( .A(u5_mult_79_CARRYB_7__19_), .B(
        u5_mult_79_ab_8__19_), .CI(u5_mult_79_SUMB_7__20_), .CO(
        u5_mult_79_CARRYB_8__19_), .S(u5_mult_79_SUMB_8__19_) );
  FA_X1 u5_mult_79_S2_8_11 ( .A(u5_mult_79_ab_8__11_), .B(
        u5_mult_79_CARRYB_7__11_), .CI(u5_mult_79_SUMB_7__12_), .CO(
        u5_mult_79_CARRYB_8__11_), .S(u5_mult_79_SUMB_8__11_) );
  FA_X1 u5_mult_79_S2_8_10 ( .A(u5_mult_79_CARRYB_7__10_), .B(
        u5_mult_79_ab_8__10_), .CI(u5_mult_79_SUMB_7__11_), .CO(
        u5_mult_79_CARRYB_8__10_), .S(u5_mult_79_SUMB_8__10_) );
  FA_X1 u5_mult_79_S2_8_9 ( .A(u5_mult_79_ab_8__9_), .B(
        u5_mult_79_CARRYB_7__9_), .CI(u5_mult_79_SUMB_7__10_), .CO(
        u5_mult_79_CARRYB_8__9_), .S(u5_mult_79_SUMB_8__9_) );
  FA_X1 u5_mult_79_S2_8_5 ( .A(u5_mult_79_CARRYB_7__5_), .B(
        u5_mult_79_ab_8__5_), .CI(u5_mult_79_SUMB_7__6_), .CO(
        u5_mult_79_CARRYB_8__5_), .S(u5_mult_79_SUMB_8__5_) );
  FA_X1 u5_mult_79_S2_8_4 ( .A(u5_mult_79_ab_8__4_), .B(
        u5_mult_79_CARRYB_7__4_), .CI(u5_mult_79_SUMB_7__5_), .CO(
        u5_mult_79_CARRYB_8__4_), .S(u5_mult_79_SUMB_8__4_) );
  FA_X1 u5_mult_79_S2_8_3 ( .A(u5_mult_79_ab_8__3_), .B(
        u5_mult_79_CARRYB_7__3_), .CI(u5_mult_79_SUMB_7__4_), .CO(
        u5_mult_79_CARRYB_8__3_), .S(u5_mult_79_SUMB_8__3_) );
  FA_X1 u5_mult_79_S2_8_2 ( .A(u5_mult_79_ab_8__2_), .B(
        u5_mult_79_CARRYB_7__2_), .CI(u5_mult_79_SUMB_7__3_), .CO(
        u5_mult_79_CARRYB_8__2_), .S(u5_mult_79_SUMB_8__2_) );
  FA_X1 u5_mult_79_S2_8_1 ( .A(u5_mult_79_ab_8__1_), .B(
        u5_mult_79_CARRYB_7__1_), .CI(u5_mult_79_SUMB_7__2_), .CO(
        u5_mult_79_CARRYB_8__1_), .S(u5_mult_79_SUMB_8__1_) );
  FA_X1 u5_mult_79_S1_8_0 ( .A(u5_mult_79_ab_8__0_), .B(
        u5_mult_79_CARRYB_7__0_), .CI(u5_mult_79_SUMB_7__1_), .CO(
        u5_mult_79_CARRYB_8__0_), .S(u5_N8) );
  FA_X1 u5_mult_79_S3_9_22 ( .A(u5_mult_79_ab_9__22_), .B(u5_mult_79_ab_8__23_), .CI(u5_mult_79_CARRYB_8__22_), .CO(u5_mult_79_CARRYB_9__22_), .S(
        u5_mult_79_SUMB_9__22_) );
  FA_X1 u5_mult_79_S2_9_21 ( .A(u5_mult_79_CARRYB_8__21_), .B(
        u5_mult_79_ab_9__21_), .CI(u5_mult_79_SUMB_8__22_), .CO(
        u5_mult_79_CARRYB_9__21_), .S(u5_mult_79_SUMB_9__21_) );
  FA_X1 u5_mult_79_S2_9_20 ( .A(u5_mult_79_CARRYB_8__20_), .B(
        u5_mult_79_ab_9__20_), .CI(u5_mult_79_SUMB_8__21_), .CO(
        u5_mult_79_CARRYB_9__20_), .S(u5_mult_79_SUMB_9__20_) );
  FA_X1 u5_mult_79_S2_9_18 ( .A(u5_mult_79_CARRYB_8__18_), .B(
        u5_mult_79_ab_9__18_), .CI(u5_mult_79_SUMB_8__19_), .CO(
        u5_mult_79_CARRYB_9__18_), .S(u5_mult_79_SUMB_9__18_) );
  FA_X1 u5_mult_79_S2_9_12 ( .A(u5_mult_79_CARRYB_8__12_), .B(
        u5_mult_79_ab_9__12_), .CI(u5_mult_79_SUMB_8__13_), .CO(
        u5_mult_79_CARRYB_9__12_), .S(u5_mult_79_SUMB_9__12_) );
  FA_X1 u5_mult_79_S2_9_10 ( .A(u5_mult_79_ab_9__10_), .B(
        u5_mult_79_CARRYB_8__10_), .CI(u5_mult_79_SUMB_8__11_), .CO(
        u5_mult_79_CARRYB_9__10_), .S(u5_mult_79_SUMB_9__10_) );
  FA_X1 u5_mult_79_S2_9_9 ( .A(u5_mult_79_CARRYB_8__9_), .B(
        u5_mult_79_ab_9__9_), .CI(u5_mult_79_SUMB_8__10_), .CO(
        u5_mult_79_CARRYB_9__9_), .S(u5_mult_79_SUMB_9__9_) );
  FA_X1 u5_mult_79_S2_9_6 ( .A(u5_mult_79_ab_9__6_), .B(
        u5_mult_79_CARRYB_8__6_), .CI(u5_mult_79_SUMB_8__7_), .CO(
        u5_mult_79_CARRYB_9__6_), .S(u5_mult_79_SUMB_9__6_) );
  FA_X1 u5_mult_79_S2_9_4 ( .A(u5_mult_79_CARRYB_8__4_), .B(
        u5_mult_79_ab_9__4_), .CI(u5_mult_79_SUMB_8__5_), .CO(
        u5_mult_79_CARRYB_9__4_), .S(u5_mult_79_SUMB_9__4_) );
  FA_X1 u5_mult_79_S2_9_3 ( .A(u5_mult_79_CARRYB_8__3_), .B(
        u5_mult_79_ab_9__3_), .CI(u5_mult_79_SUMB_8__4_), .CO(
        u5_mult_79_CARRYB_9__3_), .S(u5_mult_79_SUMB_9__3_) );
  FA_X1 u5_mult_79_S2_9_2 ( .A(u5_mult_79_ab_9__2_), .B(
        u5_mult_79_CARRYB_8__2_), .CI(u5_mult_79_SUMB_8__3_), .CO(
        u5_mult_79_CARRYB_9__2_), .S(u5_mult_79_SUMB_9__2_) );
  FA_X1 u5_mult_79_S2_9_1 ( .A(u5_mult_79_ab_9__1_), .B(
        u5_mult_79_CARRYB_8__1_), .CI(u5_mult_79_SUMB_8__2_), .CO(
        u5_mult_79_CARRYB_9__1_), .S(u5_mult_79_SUMB_9__1_) );
  FA_X1 u5_mult_79_S1_9_0 ( .A(u5_mult_79_ab_9__0_), .B(
        u5_mult_79_CARRYB_8__0_), .CI(u5_mult_79_SUMB_8__1_), .CO(
        u5_mult_79_CARRYB_9__0_), .S(u5_N9) );
  FA_X1 u5_mult_79_S2_10_21 ( .A(u5_mult_79_CARRYB_9__21_), .B(
        u5_mult_79_ab_10__21_), .CI(u5_mult_79_SUMB_9__22_), .CO(
        u5_mult_79_CARRYB_10__21_), .S(u5_mult_79_SUMB_10__21_) );
  FA_X1 u5_mult_79_S2_10_17 ( .A(u5_mult_79_ab_10__17_), .B(
        u5_mult_79_CARRYB_9__17_), .CI(u5_mult_79_SUMB_9__18_), .CO(
        u5_mult_79_CARRYB_10__17_), .S(u5_mult_79_SUMB_10__17_) );
  FA_X1 u5_mult_79_S2_10_16 ( .A(u5_mult_79_ab_10__16_), .B(
        u5_mult_79_CARRYB_9__16_), .CI(u5_mult_79_SUMB_9__17_), .CO(
        u5_mult_79_CARRYB_10__16_), .S(u5_mult_79_SUMB_10__16_) );
  FA_X1 u5_mult_79_S2_10_14 ( .A(u5_mult_79_ab_10__14_), .B(
        u5_mult_79_CARRYB_9__14_), .CI(u5_mult_79_SUMB_9__15_), .CO(
        u5_mult_79_CARRYB_10__14_), .S(u5_mult_79_SUMB_10__14_) );
  FA_X1 u5_mult_79_S2_10_7 ( .A(u5_mult_79_ab_10__7_), .B(
        u5_mult_79_CARRYB_9__7_), .CI(u5_mult_79_SUMB_9__8_), .CO(
        u5_mult_79_CARRYB_10__7_), .S(u5_mult_79_SUMB_10__7_) );
  FA_X1 u5_mult_79_S2_10_6 ( .A(u5_mult_79_ab_10__6_), .B(
        u5_mult_79_CARRYB_9__6_), .CI(u5_mult_79_SUMB_9__7_), .CO(
        u5_mult_79_CARRYB_10__6_), .S(u5_mult_79_SUMB_10__6_) );
  FA_X1 u5_mult_79_S2_10_3 ( .A(u5_mult_79_CARRYB_9__3_), .B(
        u5_mult_79_ab_10__3_), .CI(u5_mult_79_SUMB_9__4_), .CO(
        u5_mult_79_CARRYB_10__3_), .S(u5_mult_79_SUMB_10__3_) );
  FA_X1 u5_mult_79_S2_10_2 ( .A(u5_mult_79_ab_10__2_), .B(
        u5_mult_79_CARRYB_9__2_), .CI(u5_mult_79_SUMB_9__3_), .CO(
        u5_mult_79_CARRYB_10__2_), .S(u5_mult_79_SUMB_10__2_) );
  FA_X1 u5_mult_79_S2_10_1 ( .A(u5_mult_79_ab_10__1_), .B(
        u5_mult_79_CARRYB_9__1_), .CI(u5_mult_79_SUMB_9__2_), .CO(
        u5_mult_79_CARRYB_10__1_), .S(u5_mult_79_SUMB_10__1_) );
  FA_X1 u5_mult_79_S1_10_0 ( .A(u5_mult_79_ab_10__0_), .B(
        u5_mult_79_CARRYB_9__0_), .CI(u5_mult_79_SUMB_9__1_), .CO(
        u5_mult_79_CARRYB_10__0_), .S(u5_N10) );
  FA_X1 u5_mult_79_S3_11_22 ( .A(u5_mult_79_ab_11__22_), .B(
        u5_mult_79_CARRYB_10__22_), .CI(u5_mult_79_ab_10__23_), .CO(
        u5_mult_79_CARRYB_11__22_), .S(u5_mult_79_SUMB_11__22_) );
  FA_X1 u5_mult_79_S2_11_19 ( .A(u5_mult_79_CARRYB_10__19_), .B(
        u5_mult_79_ab_11__19_), .CI(u5_mult_79_SUMB_10__20_), .CO(
        u5_mult_79_CARRYB_11__19_), .S(u5_mult_79_SUMB_11__19_) );
  FA_X1 u5_mult_79_S2_11_14 ( .A(u5_mult_79_ab_11__14_), .B(
        u5_mult_79_CARRYB_10__14_), .CI(u5_mult_79_SUMB_10__15_), .CO(
        u5_mult_79_CARRYB_11__14_), .S(u5_mult_79_SUMB_11__14_) );
  FA_X1 u5_mult_79_S2_11_6 ( .A(u5_mult_79_CARRYB_10__6_), .B(
        u5_mult_79_ab_11__6_), .CI(u5_mult_79_SUMB_10__7_), .CO(
        u5_mult_79_CARRYB_11__6_), .S(u5_mult_79_SUMB_11__6_) );
  FA_X1 u5_mult_79_S2_11_1 ( .A(u5_mult_79_ab_11__1_), .B(
        u5_mult_79_CARRYB_10__1_), .CI(u5_mult_79_SUMB_10__2_), .CO(
        u5_mult_79_CARRYB_11__1_), .S(u5_mult_79_SUMB_11__1_) );
  FA_X1 u5_mult_79_S1_11_0 ( .A(u5_mult_79_ab_11__0_), .B(
        u5_mult_79_CARRYB_10__0_), .CI(u5_mult_79_SUMB_10__1_), .CO(
        u5_mult_79_CARRYB_11__0_), .S(u5_N11) );
  FA_X1 u5_mult_79_S2_12_20 ( .A(u5_mult_79_CARRYB_11__20_), .B(
        u5_mult_79_ab_12__20_), .CI(u5_mult_79_SUMB_11__21_), .CO(
        u5_mult_79_CARRYB_12__20_), .S(u5_mult_79_SUMB_12__20_) );
  FA_X1 u5_mult_79_S2_12_19 ( .A(u5_mult_79_ab_12__19_), .B(
        u5_mult_79_CARRYB_11__19_), .CI(u5_mult_79_SUMB_11__20_), .CO(
        u5_mult_79_CARRYB_12__19_), .S(u5_mult_79_SUMB_12__19_) );
  FA_X1 u5_mult_79_S2_12_18 ( .A(u5_mult_79_ab_12__18_), .B(
        u5_mult_79_CARRYB_11__18_), .CI(u5_mult_79_SUMB_11__19_), .CO(
        u5_mult_79_CARRYB_12__18_), .S(u5_mult_79_SUMB_12__18_) );
  FA_X1 u5_mult_79_S2_12_4 ( .A(u5_mult_79_ab_12__4_), .B(
        u5_mult_79_CARRYB_11__4_), .CI(u5_mult_79_SUMB_11__5_), .CO(
        u5_mult_79_CARRYB_12__4_), .S(u5_mult_79_SUMB_12__4_) );
  FA_X1 u5_mult_79_S2_12_3 ( .A(u5_mult_79_CARRYB_11__3_), .B(
        u5_mult_79_ab_12__3_), .CI(u5_mult_79_SUMB_11__4_), .CO(
        u5_mult_79_CARRYB_12__3_), .S(u5_mult_79_SUMB_12__3_) );
  FA_X1 u5_mult_79_S2_12_1 ( .A(u5_mult_79_ab_12__1_), .B(
        u5_mult_79_CARRYB_11__1_), .CI(u5_mult_79_SUMB_11__2_), .CO(
        u5_mult_79_CARRYB_12__1_), .S(u5_mult_79_SUMB_12__1_) );
  FA_X1 u5_mult_79_S1_12_0 ( .A(u5_mult_79_ab_12__0_), .B(
        u5_mult_79_CARRYB_11__0_), .CI(u5_mult_79_SUMB_11__1_), .CO(
        u5_mult_79_CARRYB_12__0_), .S(u5_N12) );
  FA_X1 u5_mult_79_S3_13_22 ( .A(u5_mult_79_ab_13__22_), .B(
        u5_mult_79_CARRYB_12__22_), .CI(u5_mult_79_ab_12__23_), .CO(
        u5_mult_79_CARRYB_13__22_), .S(u5_mult_79_SUMB_13__22_) );
  FA_X1 u5_mult_79_S2_13_20 ( .A(u5_mult_79_CARRYB_12__20_), .B(
        u5_mult_79_ab_13__20_), .CI(u5_mult_79_SUMB_12__21_), .CO(
        u5_mult_79_CARRYB_13__20_), .S(u5_mult_79_SUMB_13__20_) );
  FA_X1 u5_mult_79_S2_13_17 ( .A(u5_mult_79_ab_13__17_), .B(
        u5_mult_79_CARRYB_12__17_), .CI(u5_mult_79_SUMB_12__18_), .CO(
        u5_mult_79_CARRYB_13__17_), .S(u5_mult_79_SUMB_13__17_) );
  FA_X1 u5_mult_79_S2_13_15 ( .A(u5_mult_79_ab_13__15_), .B(
        u5_mult_79_CARRYB_12__15_), .CI(u5_mult_79_SUMB_12__16_), .CO(
        u5_mult_79_CARRYB_13__15_), .S(u5_mult_79_SUMB_13__15_) );
  FA_X1 u5_mult_79_S2_13_7 ( .A(u5_mult_79_CARRYB_12__7_), .B(
        u5_mult_79_ab_13__7_), .CI(u5_mult_79_SUMB_12__8_), .CO(
        u5_mult_79_CARRYB_13__7_), .S(u5_mult_79_SUMB_13__7_) );
  FA_X1 u5_mult_79_S2_13_3 ( .A(u5_mult_79_CARRYB_12__3_), .B(
        u5_mult_79_ab_13__3_), .CI(u5_mult_79_SUMB_12__4_), .CO(
        u5_mult_79_CARRYB_13__3_), .S(u5_mult_79_SUMB_13__3_) );
  FA_X1 u5_mult_79_S2_13_2 ( .A(u5_mult_79_ab_13__2_), .B(
        u5_mult_79_CARRYB_12__2_), .CI(u5_mult_79_SUMB_12__3_), .CO(
        u5_mult_79_CARRYB_13__2_), .S(u5_mult_79_SUMB_13__2_) );
  FA_X1 u5_mult_79_S3_14_22 ( .A(u5_mult_79_ab_14__22_), .B(
        u5_mult_79_CARRYB_13__22_), .CI(u5_mult_79_ab_13__23_), .CO(
        u5_mult_79_CARRYB_14__22_), .S(u5_mult_79_SUMB_14__22_) );
  FA_X1 u5_mult_79_S2_14_21 ( .A(u5_mult_79_ab_14__21_), .B(
        u5_mult_79_CARRYB_13__21_), .CI(u5_mult_79_SUMB_13__22_), .CO(
        u5_mult_79_CARRYB_14__21_), .S(u5_mult_79_SUMB_14__21_) );
  FA_X1 u5_mult_79_S2_14_18 ( .A(u5_mult_79_CARRYB_13__18_), .B(
        u5_mult_79_ab_14__18_), .CI(u5_mult_79_SUMB_13__19_), .CO(
        u5_mult_79_CARRYB_14__18_), .S(u5_mult_79_SUMB_14__18_) );
  FA_X1 u5_mult_79_S2_14_11 ( .A(u5_mult_79_ab_14__11_), .B(
        u5_mult_79_CARRYB_13__11_), .CI(u5_mult_79_SUMB_13__12_), .CO(
        u5_mult_79_CARRYB_14__11_), .S(u5_mult_79_SUMB_14__11_) );
  FA_X1 u5_mult_79_S2_14_6 ( .A(u5_mult_79_CARRYB_13__6_), .B(
        u5_mult_79_ab_14__6_), .CI(u5_mult_79_SUMB_13__7_), .CO(
        u5_mult_79_CARRYB_14__6_), .S(u5_mult_79_SUMB_14__6_) );
  FA_X1 u5_mult_79_S2_14_3 ( .A(u5_mult_79_SUMB_13__4_), .B(
        u5_mult_79_ab_14__3_), .CI(u5_mult_79_CARRYB_13__3_), .CO(
        u5_mult_79_CARRYB_14__3_), .S(u5_mult_79_SUMB_14__3_) );
  FA_X1 u5_mult_79_S3_15_22 ( .A(u5_mult_79_ab_15__22_), .B(
        u5_mult_79_CARRYB_14__22_), .CI(u5_mult_79_ab_14__23_), .CO(
        u5_mult_79_CARRYB_15__22_), .S(u5_mult_79_SUMB_15__22_) );
  FA_X1 u5_mult_79_S2_15_21 ( .A(u5_mult_79_ab_15__21_), .B(
        u5_mult_79_CARRYB_14__21_), .CI(u5_mult_79_SUMB_14__22_), .CO(
        u5_mult_79_CARRYB_15__21_), .S(u5_mult_79_SUMB_15__21_) );
  FA_X1 u5_mult_79_S2_15_20 ( .A(u5_mult_79_ab_15__20_), .B(
        u5_mult_79_CARRYB_14__20_), .CI(u5_mult_79_SUMB_14__21_), .CO(
        u5_mult_79_CARRYB_15__20_), .S(u5_mult_79_SUMB_15__20_) );
  FA_X1 u5_mult_79_S2_15_17 ( .A(u5_mult_79_CARRYB_14__17_), .B(
        u5_mult_79_ab_15__17_), .CI(u5_mult_79_SUMB_14__18_), .CO(
        u5_mult_79_CARRYB_15__17_), .S(u5_mult_79_SUMB_15__17_) );
  FA_X1 u5_mult_79_S2_15_13 ( .A(u5_mult_79_ab_15__13_), .B(
        u5_mult_79_CARRYB_14__13_), .CI(u5_mult_79_SUMB_14__14_), .CO(
        u5_mult_79_CARRYB_15__13_), .S(u5_mult_79_SUMB_15__13_) );
  FA_X1 u5_mult_79_S2_15_10 ( .A(u5_mult_79_CARRYB_14__10_), .B(
        u5_mult_79_ab_15__10_), .CI(u5_mult_79_SUMB_14__11_), .CO(
        u5_mult_79_CARRYB_15__10_), .S(u5_mult_79_SUMB_15__10_) );
  FA_X1 u5_mult_79_S2_15_4 ( .A(u5_mult_79_CARRYB_14__4_), .B(
        u5_mult_79_ab_15__4_), .CI(u5_mult_79_SUMB_14__5_), .CO(
        u5_mult_79_CARRYB_15__4_), .S(u5_mult_79_SUMB_15__4_) );
  FA_X1 u5_mult_79_S2_15_3 ( .A(u5_mult_79_SUMB_14__4_), .B(
        u5_mult_79_ab_15__3_), .CI(u5_mult_79_CARRYB_14__3_), .CO(
        u5_mult_79_CARRYB_15__3_), .S(u5_mult_79_SUMB_15__3_) );
  FA_X1 u5_mult_79_S2_15_2 ( .A(u5_mult_79_ab_15__2_), .B(
        u5_mult_79_CARRYB_14__2_), .CI(u5_mult_79_SUMB_14__3_), .CO(
        u5_mult_79_CARRYB_15__2_), .S(u5_mult_79_SUMB_15__2_) );
  FA_X1 u5_mult_79_S2_15_1 ( .A(u5_mult_79_CARRYB_14__1_), .B(
        u5_mult_79_ab_15__1_), .CI(u5_mult_79_SUMB_14__2_), .CO(
        u5_mult_79_CARRYB_15__1_), .S(u5_mult_79_SUMB_15__1_) );
  FA_X1 u5_mult_79_S1_15_0 ( .A(u5_mult_79_ab_15__0_), .B(
        u5_mult_79_CARRYB_14__0_), .CI(u5_mult_79_SUMB_14__1_), .CO(
        u5_mult_79_CARRYB_15__0_), .S(u5_N15) );
  FA_X1 u5_mult_79_S2_16_21 ( .A(u5_mult_79_ab_16__21_), .B(
        u5_mult_79_CARRYB_15__21_), .CI(u5_mult_79_SUMB_15__22_), .CO(
        u5_mult_79_CARRYB_16__21_), .S(u5_mult_79_SUMB_16__21_) );
  FA_X1 u5_mult_79_S2_16_20 ( .A(u5_mult_79_ab_16__20_), .B(
        u5_mult_79_CARRYB_15__20_), .CI(u5_mult_79_SUMB_15__21_), .CO(
        u5_mult_79_CARRYB_16__20_), .S(u5_mult_79_SUMB_16__20_) );
  FA_X1 u5_mult_79_S2_16_19 ( .A(u5_mult_79_CARRYB_15__19_), .B(
        u5_mult_79_ab_16__19_), .CI(u5_mult_79_SUMB_15__20_), .CO(
        u5_mult_79_CARRYB_16__19_), .S(u5_mult_79_SUMB_16__19_) );
  FA_X1 u5_mult_79_S2_16_18 ( .A(u5_mult_79_ab_16__18_), .B(
        u5_mult_79_CARRYB_15__18_), .CI(u5_mult_79_SUMB_15__19_), .CO(
        u5_mult_79_CARRYB_16__18_), .S(u5_mult_79_SUMB_16__18_) );
  FA_X1 u5_mult_79_S2_16_14 ( .A(u5_mult_79_ab_16__14_), .B(
        u5_mult_79_CARRYB_15__14_), .CI(u5_mult_79_SUMB_15__15_), .CO(
        u5_mult_79_CARRYB_16__14_), .S(u5_mult_79_SUMB_16__14_) );
  FA_X1 u5_mult_79_S2_16_2 ( .A(u5_mult_79_CARRYB_15__2_), .B(
        u5_mult_79_ab_16__2_), .CI(u5_mult_79_SUMB_15__3_), .CO(
        u5_mult_79_CARRYB_16__2_), .S(u5_mult_79_SUMB_16__2_) );
  FA_X1 u5_mult_79_S3_17_22 ( .A(u5_mult_79_ab_17__22_), .B(
        u5_mult_79_CARRYB_16__22_), .CI(u5_mult_79_ab_16__23_), .CO(
        u5_mult_79_CARRYB_17__22_), .S(u5_mult_79_SUMB_17__22_) );
  FA_X1 u5_mult_79_S2_17_20 ( .A(u5_mult_79_CARRYB_16__20_), .B(
        u5_mult_79_ab_17__20_), .CI(u5_mult_79_SUMB_16__21_), .CO(
        u5_mult_79_CARRYB_17__20_), .S(u5_mult_79_SUMB_17__20_) );
  FA_X1 u5_mult_79_S2_17_4 ( .A(u5_mult_79_ab_17__4_), .B(
        u5_mult_79_CARRYB_16__4_), .CI(u5_mult_79_SUMB_16__5_), .CO(
        u5_mult_79_CARRYB_17__4_), .S(u5_mult_79_SUMB_17__4_) );
  FA_X1 u5_mult_79_S2_17_3 ( .A(u5_mult_79_CARRYB_16__3_), .B(
        u5_mult_79_ab_17__3_), .CI(u5_mult_79_SUMB_16__4_), .CO(
        u5_mult_79_CARRYB_17__3_), .S(u5_mult_79_SUMB_17__3_) );
  FA_X1 u5_mult_79_S3_18_22 ( .A(u5_mult_79_ab_18__22_), .B(
        u5_mult_79_CARRYB_17__22_), .CI(u5_mult_79_ab_17__23_), .CO(
        u5_mult_79_CARRYB_18__22_), .S(u5_mult_79_SUMB_18__22_) );
  FA_X1 u5_mult_79_S2_18_21 ( .A(u5_mult_79_ab_18__21_), .B(
        u5_mult_79_CARRYB_17__21_), .CI(u5_mult_79_SUMB_17__22_), .CO(
        u5_mult_79_CARRYB_18__21_), .S(u5_mult_79_SUMB_18__21_) );
  FA_X1 u5_mult_79_S2_18_20 ( .A(u5_mult_79_CARRYB_17__20_), .B(
        u5_mult_79_ab_18__20_), .CI(u5_mult_79_SUMB_17__21_), .CO(
        u5_mult_79_CARRYB_18__20_), .S(u5_mult_79_SUMB_18__20_) );
  FA_X1 u5_mult_79_S2_18_4 ( .A(u5_mult_79_SUMB_17__5_), .B(
        u5_mult_79_ab_18__4_), .CI(u5_mult_79_CARRYB_17__4_), .CO(
        u5_mult_79_CARRYB_18__4_), .S(u5_mult_79_SUMB_18__4_) );
  FA_X1 u5_mult_79_S2_18_2 ( .A(u5_mult_79_CARRYB_17__2_), .B(
        u5_mult_79_ab_18__2_), .CI(u5_mult_79_SUMB_17__3_), .CO(
        u5_mult_79_CARRYB_18__2_), .S(u5_mult_79_SUMB_18__2_) );
  FA_X1 u5_mult_79_S2_18_1 ( .A(u5_mult_79_SUMB_17__2_), .B(
        u5_mult_79_ab_18__1_), .CI(u5_mult_79_CARRYB_17__1_), .CO(
        u5_mult_79_CARRYB_18__1_), .S(u5_mult_79_SUMB_18__1_) );
  FA_X1 u5_mult_79_S1_18_0 ( .A(u5_mult_79_ab_18__0_), .B(
        u5_mult_79_CARRYB_17__0_), .CI(u5_mult_79_SUMB_17__1_), .CO(
        u5_mult_79_CARRYB_18__0_), .S(u5_N18) );
  FA_X1 u5_mult_79_S3_19_22 ( .A(u5_mult_79_ab_19__22_), .B(
        u5_mult_79_CARRYB_18__22_), .CI(u5_mult_79_ab_18__23_), .CO(
        u5_mult_79_CARRYB_19__22_), .S(u5_mult_79_SUMB_19__22_) );
  FA_X1 u5_mult_79_S2_19_21 ( .A(u5_mult_79_ab_19__21_), .B(
        u5_mult_79_CARRYB_18__21_), .CI(u5_mult_79_SUMB_18__22_), .CO(
        u5_mult_79_CARRYB_19__21_), .S(u5_mult_79_SUMB_19__21_) );
  FA_X1 u5_mult_79_S2_19_20 ( .A(u5_mult_79_ab_19__20_), .B(
        u5_mult_79_SUMB_18__21_), .CI(u5_mult_79_CARRYB_18__20_), .CO(
        u5_mult_79_CARRYB_19__20_), .S(u5_mult_79_SUMB_19__20_) );
  FA_X1 u5_mult_79_S2_19_19 ( .A(u5_mult_79_ab_19__19_), .B(
        u5_mult_79_CARRYB_18__19_), .CI(u5_mult_79_SUMB_18__20_), .CO(
        u5_mult_79_CARRYB_19__19_), .S(u5_mult_79_SUMB_19__19_) );
  FA_X1 u5_mult_79_S2_19_18 ( .A(u5_mult_79_ab_19__18_), .B(
        u5_mult_79_CARRYB_18__18_), .CI(u5_mult_79_SUMB_18__19_), .CO(
        u5_mult_79_CARRYB_19__18_), .S(u5_mult_79_SUMB_19__18_) );
  FA_X1 u5_mult_79_S2_19_16 ( .A(u5_mult_79_ab_19__16_), .B(
        u5_mult_79_CARRYB_18__16_), .CI(u5_mult_79_SUMB_18__17_), .CO(
        u5_mult_79_CARRYB_19__16_), .S(u5_mult_79_SUMB_19__16_) );
  FA_X1 u5_mult_79_S2_19_14 ( .A(u5_mult_79_ab_19__14_), .B(
        u5_mult_79_CARRYB_18__14_), .CI(u5_mult_79_SUMB_18__15_), .CO(
        u5_mult_79_CARRYB_19__14_), .S(u5_mult_79_SUMB_19__14_) );
  FA_X1 u5_mult_79_S2_19_8 ( .A(u5_mult_79_CARRYB_18__8_), .B(
        u5_mult_79_ab_19__8_), .CI(u5_mult_79_SUMB_18__9_), .CO(
        u5_mult_79_CARRYB_19__8_), .S(u5_mult_79_SUMB_19__8_) );
  FA_X1 u5_mult_79_S2_19_6 ( .A(u5_mult_79_CARRYB_18__6_), .B(
        u5_mult_79_ab_19__6_), .CI(u5_mult_79_SUMB_18__7_), .CO(
        u5_mult_79_CARRYB_19__6_), .S(u5_mult_79_SUMB_19__6_) );
  FA_X1 u5_mult_79_S2_19_3 ( .A(u5_mult_79_CARRYB_18__3_), .B(
        u5_mult_79_ab_19__3_), .CI(u5_mult_79_SUMB_18__4_), .CO(
        u5_mult_79_CARRYB_19__3_), .S(u5_mult_79_SUMB_19__3_) );
  FA_X1 u5_mult_79_S2_19_1 ( .A(u5_mult_79_CARRYB_18__1_), .B(
        u5_mult_79_ab_19__1_), .CI(u5_mult_79_SUMB_18__2_), .CO(
        u5_mult_79_CARRYB_19__1_), .S(u5_mult_79_SUMB_19__1_) );
  FA_X1 u5_mult_79_S3_20_22 ( .A(u5_mult_79_ab_20__22_), .B(
        u5_mult_79_CARRYB_19__22_), .CI(u5_mult_79_ab_19__23_), .CO(
        u5_mult_79_CARRYB_20__22_), .S(u5_mult_79_SUMB_20__22_) );
  FA_X1 u5_mult_79_S2_20_21 ( .A(u5_mult_79_ab_20__21_), .B(
        u5_mult_79_CARRYB_19__21_), .CI(u5_mult_79_SUMB_19__22_), .CO(
        u5_mult_79_CARRYB_20__21_), .S(u5_mult_79_SUMB_20__21_) );
  FA_X1 u5_mult_79_S2_20_20 ( .A(u5_mult_79_ab_20__20_), .B(
        u5_mult_79_CARRYB_19__20_), .CI(u5_mult_79_SUMB_19__21_), .CO(
        u5_mult_79_CARRYB_20__20_), .S(u5_mult_79_SUMB_20__20_) );
  FA_X1 u5_mult_79_S2_20_17 ( .A(u5_mult_79_CARRYB_19__17_), .B(
        u5_mult_79_ab_20__17_), .CI(u5_mult_79_SUMB_19__18_), .CO(
        u5_mult_79_CARRYB_20__17_), .S(u5_mult_79_SUMB_20__17_) );
  FA_X1 u5_mult_79_S2_20_12 ( .A(u5_mult_79_ab_20__12_), .B(
        u5_mult_79_CARRYB_19__12_), .CI(u5_mult_79_SUMB_19__13_), .CO(
        u5_mult_79_CARRYB_20__12_), .S(u5_mult_79_SUMB_20__12_) );
  FA_X1 u5_mult_79_S2_20_9 ( .A(u5_mult_79_CARRYB_19__9_), .B(
        u5_mult_79_ab_20__9_), .CI(u5_mult_79_n333), .CO(
        u5_mult_79_CARRYB_20__9_), .S(u5_mult_79_SUMB_20__9_) );
  FA_X1 u5_mult_79_S2_20_6 ( .A(u5_mult_79_CARRYB_19__6_), .B(
        u5_mult_79_ab_20__6_), .CI(u5_mult_79_SUMB_19__7_), .CO(
        u5_mult_79_CARRYB_20__6_), .S(u5_mult_79_SUMB_20__6_) );
  FA_X1 u5_mult_79_S2_20_5 ( .A(u5_mult_79_CARRYB_19__5_), .B(
        u5_mult_79_ab_20__5_), .CI(u5_mult_79_SUMB_19__6_), .CO(
        u5_mult_79_CARRYB_20__5_), .S(u5_mult_79_SUMB_20__5_) );
  FA_X1 u5_mult_79_S3_21_22 ( .A(u5_mult_79_ab_21__22_), .B(
        u5_mult_79_CARRYB_20__22_), .CI(u5_mult_79_ab_20__23_), .CO(
        u5_mult_79_CARRYB_21__22_), .S(u5_mult_79_SUMB_21__22_) );
  FA_X1 u5_mult_79_S2_21_21 ( .A(u5_mult_79_ab_21__21_), .B(
        u5_mult_79_CARRYB_20__21_), .CI(u5_mult_79_SUMB_20__22_), .CO(
        u5_mult_79_CARRYB_21__21_), .S(u5_mult_79_SUMB_21__21_) );
  FA_X1 u5_mult_79_S2_21_20 ( .A(u5_mult_79_ab_21__20_), .B(
        u5_mult_79_CARRYB_20__20_), .CI(u5_mult_79_SUMB_20__21_), .CO(
        u5_mult_79_CARRYB_21__20_), .S(u5_mult_79_SUMB_21__20_) );
  FA_X1 u5_mult_79_S2_21_19 ( .A(u5_mult_79_ab_21__19_), .B(
        u5_mult_79_CARRYB_20__19_), .CI(u5_mult_79_SUMB_20__20_), .CO(
        u5_mult_79_CARRYB_21__19_), .S(u5_mult_79_SUMB_21__19_) );
  FA_X1 u5_mult_79_S2_21_16 ( .A(u5_mult_79_CARRYB_20__16_), .B(
        u5_mult_79_ab_21__16_), .CI(u5_mult_79_SUMB_20__17_), .CO(
        u5_mult_79_CARRYB_21__16_), .S(u5_mult_79_SUMB_21__16_) );
  FA_X1 u5_mult_79_S3_22_22 ( .A(u5_mult_79_ab_22__22_), .B(
        u5_mult_79_CARRYB_21__22_), .CI(u5_mult_79_ab_21__23_), .CO(
        u5_mult_79_CARRYB_22__22_), .S(u5_mult_79_SUMB_22__22_) );
  FA_X1 u5_mult_79_S2_22_21 ( .A(u5_mult_79_ab_22__21_), .B(
        u5_mult_79_CARRYB_21__21_), .CI(u5_mult_79_SUMB_21__22_), .CO(
        u5_mult_79_CARRYB_22__21_), .S(u5_mult_79_SUMB_22__21_) );
  FA_X1 u5_mult_79_S2_22_20 ( .A(u5_mult_79_ab_22__20_), .B(
        u5_mult_79_CARRYB_21__20_), .CI(u5_mult_79_SUMB_21__21_), .CO(
        u5_mult_79_CARRYB_22__20_), .S(u5_mult_79_SUMB_22__20_) );
  FA_X1 u5_mult_79_S2_22_19 ( .A(u5_mult_79_ab_22__19_), .B(
        u5_mult_79_CARRYB_21__19_), .CI(u5_mult_79_SUMB_21__20_), .CO(
        u5_mult_79_CARRYB_22__19_), .S(u5_mult_79_SUMB_22__19_) );
  FA_X1 u5_mult_79_S2_22_18 ( .A(u5_mult_79_ab_22__18_), .B(
        u5_mult_79_CARRYB_21__18_), .CI(u5_mult_79_SUMB_21__19_), .CO(
        u5_mult_79_CARRYB_22__18_), .S(u5_mult_79_SUMB_22__18_) );
  FA_X1 u5_mult_79_S2_22_16 ( .A(u5_mult_79_ab_22__16_), .B(
        u5_mult_79_CARRYB_21__16_), .CI(u5_mult_79_SUMB_21__17_), .CO(
        u5_mult_79_CARRYB_22__16_), .S(u5_mult_79_SUMB_22__16_) );
  FA_X1 u5_mult_79_S2_22_15 ( .A(u5_mult_79_CARRYB_21__15_), .B(
        u5_mult_79_ab_22__15_), .CI(u5_mult_79_SUMB_21__16_), .CO(
        u5_mult_79_CARRYB_22__15_), .S(u5_mult_79_SUMB_22__15_) );
  FA_X1 u5_mult_79_S2_22_13 ( .A(u5_mult_79_ab_22__13_), .B(
        u5_mult_79_CARRYB_21__13_), .CI(u5_mult_79_SUMB_21__14_), .CO(
        u5_mult_79_CARRYB_22__13_), .S(u5_mult_79_SUMB_22__13_) );
  FA_X1 u5_mult_79_S1_22_0 ( .A(u5_mult_79_CARRYB_21__0_), .B(
        u5_mult_79_ab_22__0_), .CI(u5_mult_79_SUMB_21__1_), .CO(
        u5_mult_79_CARRYB_22__0_), .S(u5_N22) );
  FA_X1 u5_mult_79_S5_22 ( .A(u5_mult_79_ab_23__22_), .B(
        u5_mult_79_CARRYB_22__22_), .CI(u5_mult_79_ab_22__23_), .CO(
        u5_mult_79_CARRYB_23__22_), .S(u5_mult_79_SUMB_23__22_) );
  FA_X1 u5_mult_79_S4_21 ( .A(u5_mult_79_ab_23__21_), .B(
        u5_mult_79_CARRYB_22__21_), .CI(u5_mult_79_SUMB_22__22_), .CO(
        u5_mult_79_CARRYB_23__21_), .S(u5_mult_79_SUMB_23__21_) );
  FA_X1 u5_mult_79_S4_20 ( .A(u5_mult_79_ab_23__20_), .B(
        u5_mult_79_CARRYB_22__20_), .CI(u5_mult_79_SUMB_22__21_), .CO(
        u5_mult_79_CARRYB_23__20_), .S(u5_mult_79_SUMB_23__20_) );
  FA_X1 u5_mult_79_S4_19 ( .A(u5_mult_79_ab_23__19_), .B(
        u5_mult_79_CARRYB_22__19_), .CI(u5_mult_79_SUMB_22__20_), .CO(
        u5_mult_79_CARRYB_23__19_), .S(u5_mult_79_SUMB_23__19_) );
  FA_X1 u5_mult_79_S4_18 ( .A(u5_mult_79_ab_23__18_), .B(
        u5_mult_79_CARRYB_22__18_), .CI(u5_mult_79_SUMB_22__19_), .CO(
        u5_mult_79_CARRYB_23__18_), .S(u5_mult_79_SUMB_23__18_) );
  FA_X1 u5_mult_79_S4_17 ( .A(u5_mult_79_ab_23__17_), .B(
        u5_mult_79_CARRYB_22__17_), .CI(u5_mult_79_SUMB_22__18_), .CO(
        u5_mult_79_CARRYB_23__17_), .S(u5_mult_79_SUMB_23__17_) );
  FA_X1 u5_mult_79_S4_16 ( .A(u5_mult_79_CARRYB_22__16_), .B(
        u5_mult_79_ab_23__16_), .CI(u5_mult_79_SUMB_22__17_), .CO(
        u5_mult_79_CARRYB_23__16_), .S(u5_mult_79_SUMB_23__16_) );
  FA_X1 u5_mult_79_S4_15 ( .A(u5_mult_79_CARRYB_22__15_), .B(
        u5_mult_79_ab_23__15_), .CI(u5_mult_79_SUMB_22__16_), .CO(
        u5_mult_79_CARRYB_23__15_), .S(u5_mult_79_SUMB_23__15_) );
  FA_X1 u5_mult_79_S4_14 ( .A(u5_mult_79_ab_23__14_), .B(
        u5_mult_79_CARRYB_22__14_), .CI(u5_mult_79_SUMB_22__15_), .CO(
        u5_mult_79_CARRYB_23__14_), .S(u5_mult_79_SUMB_23__14_) );
  FA_X1 u5_mult_79_S4_13 ( .A(u5_mult_79_CARRYB_22__13_), .B(
        u5_mult_79_ab_23__13_), .CI(u5_mult_79_SUMB_22__14_), .CO(
        u5_mult_79_CARRYB_23__13_), .S(u5_mult_79_SUMB_23__13_) );
  FA_X1 u5_mult_79_S4_7 ( .A(u5_mult_79_ab_23__7_), .B(
        u5_mult_79_CARRYB_22__7_), .CI(u5_mult_79_SUMB_22__8_), .CO(
        u5_mult_79_CARRYB_23__7_), .S(u5_mult_79_SUMB_23__7_) );
  FA_X1 u5_mult_79_S4_6 ( .A(u5_mult_79_CARRYB_22__6_), .B(
        u5_mult_79_ab_23__6_), .CI(u5_mult_79_SUMB_22__7_), .CO(
        u5_mult_79_CARRYB_23__6_), .S(u5_mult_79_SUMB_23__6_) );
  FA_X1 u5_mult_79_S4_5 ( .A(u5_mult_79_ab_23__5_), .B(
        u5_mult_79_CARRYB_22__5_), .CI(u5_mult_79_SUMB_22__6_), .CO(
        u5_mult_79_CARRYB_23__5_), .S(u5_mult_79_SUMB_23__5_) );
  FA_X1 u5_mult_79_S4_4 ( .A(u5_mult_79_ab_23__4_), .B(
        u5_mult_79_CARRYB_22__4_), .CI(u5_mult_79_SUMB_22__5_), .CO(
        u5_mult_79_CARRYB_23__4_), .S(u5_mult_79_SUMB_23__4_) );
  FA_X1 u5_mult_79_S4_3 ( .A(u5_mult_79_CARRYB_22__3_), .B(
        u5_mult_79_ab_23__3_), .CI(u5_mult_79_SUMB_22__4_), .CO(
        u5_mult_79_CARRYB_23__3_), .S(u5_mult_79_SUMB_23__3_) );
  INV_X4 u5_mult_79_FS_1_U309 ( .A(u5_mult_79_CLA_CARRY[24]), .ZN(
        u5_mult_79_FS_1_n284) );
  XNOR2_X2 u5_mult_79_FS_1_U308 ( .A(u5_mult_79_FS_1_n282), .B(
        u5_mult_79_FS_1_n56), .ZN(u5_N26) );
  XNOR2_X2 u5_mult_79_FS_1_U307 ( .A(u5_mult_79_FS_1_n280), .B(
        u5_mult_79_FS_1_n281), .ZN(u5_N27) );
  INV_X4 u5_mult_79_FS_1_U306 ( .A(u5_mult_79_FS_1_n279), .ZN(
        u5_mult_79_FS_1_n270) );
  NOR2_X4 u5_mult_79_FS_1_U305 ( .A1(u5_mult_79_CLA_SUM[28]), .A2(
        u5_mult_79_CLA_CARRY[27]), .ZN(u5_mult_79_FS_1_n261) );
  INV_X4 u5_mult_79_FS_1_U304 ( .A(u5_mult_79_FS_1_n278), .ZN(
        u5_mult_79_FS_1_n271) );
  XNOR2_X2 u5_mult_79_FS_1_U303 ( .A(u5_mult_79_FS_1_n269), .B(
        u5_mult_79_FS_1_n271), .ZN(u5_N28) );
  INV_X4 u5_mult_79_FS_1_U302 ( .A(u5_mult_79_n238), .ZN(u5_mult_79_FS_1_n267)
         );
  INV_X4 u5_mult_79_FS_1_U301 ( .A(u5_mult_79_FS_1_n253), .ZN(
        u5_mult_79_FS_1_n197) );
  XNOR2_X2 u5_mult_79_FS_1_U300 ( .A(u5_mult_79_FS_1_n264), .B(
        u5_mult_79_FS_1_n265), .ZN(u5_N29) );
  INV_X4 u5_mult_79_FS_1_U299 ( .A(u5_mult_79_n233), .ZN(u5_mult_79_FS_1_n262)
         );
  INV_X4 u5_mult_79_FS_1_U298 ( .A(u5_mult_79_CLA_SUM[30]), .ZN(
        u5_mult_79_FS_1_n263) );
  NAND2_X2 u5_mult_79_FS_1_U297 ( .A1(u5_mult_79_n233), .A2(
        u5_mult_79_CLA_SUM[30]), .ZN(u5_mult_79_FS_1_n220) );
  NOR2_X4 u5_mult_79_FS_1_U296 ( .A1(u5_mult_79_FS_1_n254), .A2(
        u5_mult_79_FS_1_n261), .ZN(u5_mult_79_FS_1_n213) );
  NOR2_X4 u5_mult_79_FS_1_U295 ( .A1(u5_mult_79_n1718), .A2(
        u5_mult_79_CLA_CARRY[26]), .ZN(u5_mult_79_FS_1_n259) );
  NOR2_X4 u5_mult_79_FS_1_U294 ( .A1(u5_mult_79_CLA_SUM[28]), .A2(
        u5_mult_79_CLA_CARRY[27]), .ZN(u5_mult_79_FS_1_n258) );
  INV_X4 u5_mult_79_FS_1_U293 ( .A(u5_mult_79_FS_1_n258), .ZN(
        u5_mult_79_FS_1_n257) );
  NAND2_X2 u5_mult_79_FS_1_U292 ( .A1(u5_mult_79_FS_1_n252), .A2(
        u5_mult_79_FS_1_n253), .ZN(u5_mult_79_FS_1_n241) );
  XNOR2_X2 u5_mult_79_FS_1_U291 ( .A(u5_mult_79_FS_1_n249), .B(
        u5_mult_79_FS_1_n248), .ZN(u5_N30) );
  INV_X4 u5_mult_79_FS_1_U290 ( .A(u5_mult_79_n232), .ZN(u5_mult_79_FS_1_n246)
         );
  INV_X4 u5_mult_79_FS_1_U289 ( .A(u5_mult_79_CLA_SUM[31]), .ZN(
        u5_mult_79_FS_1_n247) );
  INV_X4 u5_mult_79_FS_1_U288 ( .A(u5_mult_79_n234), .ZN(u5_mult_79_FS_1_n238)
         );
  INV_X4 u5_mult_79_FS_1_U287 ( .A(u5_mult_79_CLA_SUM[32]), .ZN(
        u5_mult_79_FS_1_n239) );
  NAND2_X2 u5_mult_79_FS_1_U286 ( .A1(u5_mult_79_n234), .A2(
        u5_mult_79_CLA_SUM[32]), .ZN(u5_mult_79_FS_1_n202) );
  XNOR2_X2 u5_mult_79_FS_1_U285 ( .A(u5_mult_79_FS_1_n235), .B(
        u5_mult_79_FS_1_n234), .ZN(u5_N32) );
  INV_X4 u5_mult_79_FS_1_U284 ( .A(u5_mult_79_n230), .ZN(u5_mult_79_FS_1_n232)
         );
  INV_X4 u5_mult_79_FS_1_U283 ( .A(u5_mult_79_FS_1_n231), .ZN(
        u5_mult_79_FS_1_n223) );
  INV_X4 u5_mult_79_FS_1_U282 ( .A(u5_mult_79_FS_1_n202), .ZN(
        u5_mult_79_FS_1_n227) );
  XNOR2_X2 u5_mult_79_FS_1_U281 ( .A(u5_mult_79_FS_1_n224), .B(
        u5_mult_79_FS_1_n223), .ZN(u5_N33) );
  NAND2_X2 u5_mult_79_FS_1_U280 ( .A1(u5_mult_79_CLA_CARRY[33]), .A2(
        u5_mult_79_CLA_SUM[34]), .ZN(u5_mult_79_FS_1_n222) );
  INV_X4 u5_mult_79_FS_1_U279 ( .A(u5_mult_79_FS_1_n222), .ZN(
        u5_mult_79_FS_1_n189) );
  NOR2_X4 u5_mult_79_FS_1_U278 ( .A1(u5_mult_79_CLA_SUM[34]), .A2(
        u5_mult_79_CLA_CARRY[33]), .ZN(u5_mult_79_FS_1_n181) );
  INV_X4 u5_mult_79_FS_1_U277 ( .A(u5_mult_79_FS_1_n221), .ZN(
        u5_mult_79_FS_1_n190) );
  INV_X4 u5_mult_79_FS_1_U276 ( .A(u5_mult_79_FS_1_n220), .ZN(
        u5_mult_79_FS_1_n216) );
  INV_X4 u5_mult_79_FS_1_U275 ( .A(u5_mult_79_FS_1_n199), .ZN(
        u5_mult_79_FS_1_n219) );
  NOR2_X4 u5_mult_79_FS_1_U274 ( .A1(u5_mult_79_FS_1_n219), .A2(
        u5_mult_79_FS_1_n204), .ZN(u5_mult_79_FS_1_n218) );
  NAND3_X4 u5_mult_79_FS_1_U273 ( .A1(u5_mult_79_FS_1_n218), .A2(
        u5_mult_79_FS_1_n210), .A3(u5_mult_79_FS_1_n8), .ZN(
        u5_mult_79_FS_1_n217) );
  NAND2_X2 u5_mult_79_FS_1_U272 ( .A1(u5_mult_79_FS_1_n204), .A2(
        u5_mult_79_FS_1_n201), .ZN(u5_mult_79_FS_1_n198) );
  NAND3_X2 u5_mult_79_FS_1_U271 ( .A1(u5_mult_79_FS_1_n201), .A2(
        u5_mult_79_FS_1_n202), .A3(u5_mult_79_FS_1_n203), .ZN(
        u5_mult_79_FS_1_n200) );
  INV_X4 u5_mult_79_FS_1_U270 ( .A(u5_mult_79_FS_1_n53), .ZN(
        u5_mult_79_FS_1_n194) );
  NOR3_X4 u5_mult_79_FS_1_U269 ( .A1(u5_mult_79_FS_1_n61), .A2(
        u5_mult_79_FS_1_n194), .A3(u5_mult_79_FS_1_n195), .ZN(
        u5_mult_79_FS_1_n193) );
  NAND3_X4 u5_mult_79_FS_1_U268 ( .A1(u5_mult_79_FS_1_n191), .A2(
        u5_mult_79_FS_1_n192), .A3(u5_mult_79_FS_1_n193), .ZN(
        u5_mult_79_FS_1_n173) );
  NAND2_X2 u5_mult_79_FS_1_U267 ( .A1(u5_mult_79_CLA_CARRY[34]), .A2(
        u5_mult_79_CLA_SUM[35]), .ZN(u5_mult_79_FS_1_n183) );
  INV_X4 u5_mult_79_FS_1_U266 ( .A(u5_mult_79_CLA_CARRY[34]), .ZN(
        u5_mult_79_FS_1_n186) );
  XNOR2_X2 u5_mult_79_FS_1_U265 ( .A(u5_mult_79_FS_1_n185), .B(
        u5_mult_79_FS_1_n14), .ZN(u5_N35) );
  NAND3_X4 u5_mult_79_FS_1_U264 ( .A1(u5_mult_79_CLA_SUM[34]), .A2(
        u5_mult_79_CLA_CARRY[33]), .A3(u5_mult_79_FS_1_n182), .ZN(
        u5_mult_79_FS_1_n184) );
  NAND2_X2 u5_mult_79_FS_1_U263 ( .A1(u5_mult_79_FS_1_n173), .A2(
        u5_mult_79_FS_1_n172), .ZN(u5_mult_79_FS_1_n179) );
  NAND2_X2 u5_mult_79_FS_1_U262 ( .A1(u5_mult_79_FS_1_n178), .A2(
        u5_mult_79_FS_1_n179), .ZN(u5_mult_79_FS_1_n174) );
  NAND2_X2 u5_mult_79_FS_1_U261 ( .A1(u5_mult_79_n229), .A2(
        u5_mult_79_CLA_SUM[36]), .ZN(u5_mult_79_FS_1_n156) );
  INV_X4 u5_mult_79_FS_1_U260 ( .A(u5_mult_79_n229), .ZN(u5_mult_79_FS_1_n176)
         );
  INV_X4 u5_mult_79_FS_1_U259 ( .A(u5_mult_79_CLA_SUM[36]), .ZN(
        u5_mult_79_FS_1_n177) );
  XNOR2_X2 u5_mult_79_FS_1_U258 ( .A(u5_mult_79_FS_1_n174), .B(
        u5_mult_79_FS_1_n175), .ZN(u5_N36) );
  NAND2_X2 u5_mult_79_FS_1_U257 ( .A1(u5_mult_79_FS_1_n172), .A2(
        u5_mult_79_FS_1_n171), .ZN(u5_mult_79_FS_1_n161) );
  OAI211_X2 u5_mult_79_FS_1_U256 ( .C1(u5_mult_79_FS_1_n169), .C2(
        u5_mult_79_FS_1_n161), .A(u5_mult_79_FS_1_n10), .B(
        u5_mult_79_FS_1_n156), .ZN(u5_mult_79_FS_1_n165) );
  NAND2_X2 u5_mult_79_FS_1_U255 ( .A1(u5_mult_79_CLA_CARRY[36]), .A2(
        u5_mult_79_CLA_SUM[37]), .ZN(u5_mult_79_FS_1_n159) );
  INV_X4 u5_mult_79_FS_1_U254 ( .A(u5_mult_79_CLA_CARRY[36]), .ZN(
        u5_mult_79_FS_1_n167) );
  INV_X4 u5_mult_79_FS_1_U253 ( .A(u5_mult_79_CLA_SUM[37]), .ZN(
        u5_mult_79_FS_1_n168) );
  XNOR2_X2 u5_mult_79_FS_1_U252 ( .A(u5_mult_79_FS_1_n165), .B(
        u5_mult_79_FS_1_n166), .ZN(u5_N37) );
  NOR2_X4 u5_mult_79_FS_1_U251 ( .A1(u5_mult_79_CLA_SUM[38]), .A2(
        u5_mult_79_CLA_CARRY[37]), .ZN(u5_mult_79_FS_1_n135) );
  NOR2_X4 u5_mult_79_FS_1_U250 ( .A1(u5_mult_79_FS_1_n108), .A2(
        u5_mult_79_FS_1_n60), .ZN(u5_mult_79_FS_1_n164) );
  INV_X4 u5_mult_79_FS_1_U249 ( .A(u5_mult_79_FS_1_n161), .ZN(
        u5_mult_79_FS_1_n160) );
  INV_X4 u5_mult_79_FS_1_U248 ( .A(u5_mult_79_FS_1_n159), .ZN(
        u5_mult_79_FS_1_n97) );
  INV_X4 u5_mult_79_FS_1_U247 ( .A(u5_mult_79_FS_1_n158), .ZN(
        u5_mult_79_FS_1_n157) );
  AOI21_X4 u5_mult_79_FS_1_U246 ( .B1(u5_mult_79_FS_1_n155), .B2(
        u5_mult_79_FS_1_n156), .A(u5_mult_79_FS_1_n157), .ZN(
        u5_mult_79_FS_1_n98) );
  OAI21_X4 u5_mult_79_FS_1_U245 ( .B1(u5_mult_79_FS_1_n153), .B2(
        u5_mult_79_FS_1_n51), .A(u5_mult_79_FS_1_n154), .ZN(
        u5_mult_79_FS_1_n117) );
  XNOR2_X2 u5_mult_79_FS_1_U244 ( .A(u5_mult_79_FS_1_n152), .B(
        u5_mult_79_FS_1_n151), .ZN(u5_N38) );
  INV_X4 u5_mult_79_FS_1_U243 ( .A(u5_mult_79_n237), .ZN(u5_mult_79_FS_1_n148)
         );
  NAND2_X2 u5_mult_79_FS_1_U242 ( .A1(u5_mult_79_n237), .A2(
        u5_mult_79_CLA_SUM[39]), .ZN(u5_mult_79_FS_1_n144) );
  INV_X4 u5_mult_79_FS_1_U241 ( .A(u5_mult_79_FS_1_n144), .ZN(
        u5_mult_79_FS_1_n129) );
  XNOR2_X2 u5_mult_79_FS_1_U240 ( .A(u5_mult_79_FS_1_n145), .B(
        u5_mult_79_FS_1_n146), .ZN(u5_N39) );
  NAND2_X2 u5_mult_79_FS_1_U239 ( .A1(u5_mult_79_CLA_CARRY[37]), .A2(
        u5_mult_79_CLA_SUM[38]), .ZN(u5_mult_79_FS_1_n134) );
  INV_X4 u5_mult_79_FS_1_U238 ( .A(u5_mult_79_n231), .ZN(u5_mult_79_FS_1_n140)
         );
  INV_X4 u5_mult_79_FS_1_U237 ( .A(u5_mult_79_CLA_SUM[40]), .ZN(
        u5_mult_79_FS_1_n141) );
  NAND2_X2 u5_mult_79_FS_1_U236 ( .A1(u5_mult_79_FS_1_n140), .A2(
        u5_mult_79_FS_1_n141), .ZN(u5_mult_79_FS_1_n139) );
  INV_X4 u5_mult_79_FS_1_U235 ( .A(u5_mult_79_FS_1_n139), .ZN(
        u5_mult_79_FS_1_n132) );
  NAND2_X2 u5_mult_79_FS_1_U234 ( .A1(u5_mult_79_n231), .A2(
        u5_mult_79_CLA_SUM[40]), .ZN(u5_mult_79_FS_1_n120) );
  INV_X4 u5_mult_79_FS_1_U233 ( .A(u5_mult_79_FS_1_n120), .ZN(
        u5_mult_79_FS_1_n138) );
  NOR2_X4 u5_mult_79_FS_1_U232 ( .A1(u5_mult_79_FS_1_n132), .A2(
        u5_mult_79_FS_1_n138), .ZN(u5_mult_79_FS_1_n137) );
  XNOR2_X2 u5_mult_79_FS_1_U231 ( .A(u5_mult_79_FS_1_n136), .B(
        u5_mult_79_FS_1_n137), .ZN(u5_N40) );
  NOR3_X4 u5_mult_79_FS_1_U230 ( .A1(u5_mult_79_FS_1_n135), .A2(
        u5_mult_79_FS_1_n132), .A3(u5_mult_79_FS_1_n133), .ZN(
        u5_mult_79_FS_1_n122) );
  INV_X4 u5_mult_79_FS_1_U229 ( .A(u5_mult_79_FS_1_n134), .ZN(
        u5_mult_79_FS_1_n130) );
  INV_X4 u5_mult_79_FS_1_U228 ( .A(u5_mult_79_n236), .ZN(u5_mult_79_FS_1_n126)
         );
  INV_X4 u5_mult_79_FS_1_U227 ( .A(u5_mult_79_CLA_SUM[41]), .ZN(
        u5_mult_79_FS_1_n127) );
  NAND2_X2 u5_mult_79_FS_1_U226 ( .A1(u5_mult_79_FS_1_n126), .A2(
        u5_mult_79_FS_1_n127), .ZN(u5_mult_79_FS_1_n118) );
  NAND2_X2 u5_mult_79_FS_1_U225 ( .A1(u5_mult_79_n236), .A2(
        u5_mult_79_CLA_SUM[41]), .ZN(u5_mult_79_FS_1_n119) );
  INV_X4 u5_mult_79_FS_1_U224 ( .A(u5_mult_79_FS_1_n119), .ZN(
        u5_mult_79_FS_1_n125) );
  NOR2_X4 u5_mult_79_FS_1_U223 ( .A1(u5_mult_79_FS_1_n26), .A2(
        u5_mult_79_FS_1_n125), .ZN(u5_mult_79_FS_1_n124) );
  XNOR2_X2 u5_mult_79_FS_1_U222 ( .A(u5_mult_79_FS_1_n123), .B(
        u5_mult_79_FS_1_n124), .ZN(u5_N41) );
  INV_X4 u5_mult_79_FS_1_U221 ( .A(u5_mult_79_CLA_CARRY[41]), .ZN(
        u5_mult_79_FS_1_n115) );
  INV_X4 u5_mult_79_FS_1_U220 ( .A(u5_mult_79_CLA_SUM[42]), .ZN(
        u5_mult_79_FS_1_n116) );
  NAND2_X2 u5_mult_79_FS_1_U219 ( .A1(u5_mult_79_CLA_CARRY[41]), .A2(
        u5_mult_79_CLA_SUM[42]), .ZN(u5_mult_79_FS_1_n114) );
  INV_X4 u5_mult_79_FS_1_U218 ( .A(u5_mult_79_FS_1_n114), .ZN(
        u5_mult_79_FS_1_n99) );
  NOR2_X4 u5_mult_79_FS_1_U217 ( .A1(u5_mult_79_FS_1_n113), .A2(
        u5_mult_79_FS_1_n99), .ZN(u5_mult_79_FS_1_n112) );
  XNOR2_X2 u5_mult_79_FS_1_U216 ( .A(u5_mult_79_FS_1_n111), .B(
        u5_mult_79_FS_1_n112), .ZN(u5_N42) );
  NAND2_X2 u5_mult_79_FS_1_U215 ( .A1(u5_mult_79_n235), .A2(
        u5_mult_79_CLA_SUM[43]), .ZN(u5_mult_79_FS_1_n90) );
  INV_X4 u5_mult_79_FS_1_U214 ( .A(u5_mult_79_n235), .ZN(u5_mult_79_FS_1_n109)
         );
  INV_X4 u5_mult_79_FS_1_U213 ( .A(u5_mult_79_CLA_SUM[43]), .ZN(
        u5_mult_79_FS_1_n110) );
  NAND2_X2 u5_mult_79_FS_1_U212 ( .A1(u5_mult_79_FS_1_n109), .A2(
        u5_mult_79_FS_1_n110), .ZN(u5_mult_79_FS_1_n84) );
  NAND2_X2 u5_mult_79_FS_1_U211 ( .A1(u5_mult_79_FS_1_n90), .A2(
        u5_mult_79_FS_1_n84), .ZN(u5_mult_79_FS_1_n91) );
  NOR2_X4 u5_mult_79_FS_1_U210 ( .A1(u5_mult_79_FS_1_n103), .A2(
        u5_mult_79_FS_1_n104), .ZN(u5_mult_79_FS_1_n92) );
  INV_X4 u5_mult_79_FS_1_U209 ( .A(u5_mult_79_FS_1_n51), .ZN(
        u5_mult_79_FS_1_n101) );
  OAI21_X4 u5_mult_79_FS_1_U208 ( .B1(u5_mult_79_FS_1_n25), .B2(
        u5_mult_79_FS_1_n99), .A(u5_mult_79_FS_1_n100), .ZN(
        u5_mult_79_FS_1_n42) );
  INV_X4 u5_mult_79_FS_1_U207 ( .A(u5_mult_79_FS_1_n42), .ZN(
        u5_mult_79_FS_1_n95) );
  OAI21_X4 u5_mult_79_FS_1_U206 ( .B1(u5_mult_79_FS_1_n97), .B2(
        u5_mult_79_FS_1_n98), .A(u5_mult_79_FS_1_n22), .ZN(u5_mult_79_FS_1_n38) );
  NOR2_X4 u5_mult_79_FS_1_U205 ( .A1(u5_mult_79_FS_1_n95), .A2(
        u5_mult_79_FS_1_n96), .ZN(u5_mult_79_FS_1_n94) );
  OAI21_X4 u5_mult_79_FS_1_U204 ( .B1(u5_mult_79_FS_1_n92), .B2(
        u5_mult_79_FS_1_n93), .A(u5_mult_79_FS_1_n94), .ZN(u5_mult_79_FS_1_n68) );
  INV_X4 u5_mult_79_FS_1_U203 ( .A(u5_mult_79_FS_1_n90), .ZN(
        u5_mult_79_FS_1_n79) );
  INV_X4 u5_mult_79_FS_1_U202 ( .A(u5_mult_79_n244), .ZN(u5_mult_79_FS_1_n88)
         );
  INV_X4 u5_mult_79_FS_1_U201 ( .A(u5_mult_79_CLA_SUM[44]), .ZN(
        u5_mult_79_FS_1_n89) );
  NAND2_X2 u5_mult_79_FS_1_U200 ( .A1(u5_mult_79_FS_1_n88), .A2(
        u5_mult_79_FS_1_n89), .ZN(u5_mult_79_FS_1_n81) );
  INV_X4 u5_mult_79_FS_1_U199 ( .A(u5_mult_79_FS_1_n81), .ZN(
        u5_mult_79_FS_1_n82) );
  NAND2_X2 u5_mult_79_FS_1_U198 ( .A1(u5_mult_79_n244), .A2(
        u5_mult_79_CLA_SUM[44]), .ZN(u5_mult_79_FS_1_n87) );
  INV_X4 u5_mult_79_FS_1_U197 ( .A(u5_mult_79_FS_1_n87), .ZN(
        u5_mult_79_FS_1_n80) );
  NOR2_X4 u5_mult_79_FS_1_U196 ( .A1(u5_mult_79_FS_1_n82), .A2(
        u5_mult_79_FS_1_n80), .ZN(u5_mult_79_FS_1_n86) );
  XNOR2_X2 u5_mult_79_FS_1_U195 ( .A(u5_mult_79_FS_1_n85), .B(
        u5_mult_79_FS_1_n86), .ZN(u5_N44) );
  INV_X4 u5_mult_79_FS_1_U194 ( .A(u5_mult_79_FS_1_n84), .ZN(
        u5_mult_79_FS_1_n83) );
  NOR2_X4 u5_mult_79_FS_1_U193 ( .A1(u5_mult_79_FS_1_n82), .A2(
        u5_mult_79_FS_1_n83), .ZN(u5_mult_79_FS_1_n72) );
  OAI21_X4 u5_mult_79_FS_1_U192 ( .B1(u5_mult_79_FS_1_n79), .B2(
        u5_mult_79_FS_1_n80), .A(u5_mult_79_FS_1_n81), .ZN(u5_mult_79_FS_1_n78) );
  INV_X4 u5_mult_79_FS_1_U191 ( .A(u5_mult_79_FS_1_n78), .ZN(
        u5_mult_79_FS_1_n70) );
  INV_X4 u5_mult_79_FS_1_U190 ( .A(u5_mult_79_CLA_CARRY[44]), .ZN(
        u5_mult_79_FS_1_n76) );
  INV_X4 u5_mult_79_FS_1_U189 ( .A(u5_mult_79_n242), .ZN(u5_mult_79_FS_1_n77)
         );
  NAND2_X2 u5_mult_79_FS_1_U188 ( .A1(u5_mult_79_FS_1_n76), .A2(
        u5_mult_79_FS_1_n77), .ZN(u5_mult_79_FS_1_n71) );
  INV_X4 u5_mult_79_FS_1_U187 ( .A(u5_mult_79_FS_1_n71), .ZN(
        u5_mult_79_FS_1_n75) );
  NOR2_X4 u5_mult_79_FS_1_U186 ( .A1(u5_mult_79_FS_1_n75), .A2(
        u5_mult_79_FS_1_n11), .ZN(u5_mult_79_FS_1_n74) );
  XNOR2_X2 u5_mult_79_FS_1_U185 ( .A(u5_mult_79_FS_1_n73), .B(
        u5_mult_79_FS_1_n74), .ZN(u5_N45) );
  NAND2_X2 u5_mult_79_FS_1_U184 ( .A1(u5_mult_79_FS_1_n72), .A2(
        u5_mult_79_FS_1_n71), .ZN(u5_mult_79_FS_1_n52) );
  INV_X4 u5_mult_79_FS_1_U183 ( .A(u5_mult_79_FS_1_n52), .ZN(
        u5_mult_79_FS_1_n40) );
  OAI21_X4 u5_mult_79_FS_1_U182 ( .B1(u5_mult_79_FS_1_n11), .B2(
        u5_mult_79_FS_1_n70), .A(u5_mult_79_FS_1_n71), .ZN(u5_mult_79_FS_1_n69) );
  INV_X4 u5_mult_79_FS_1_U181 ( .A(u5_mult_79_FS_1_n69), .ZN(
        u5_mult_79_FS_1_n45) );
  INV_X4 u5_mult_79_FS_1_U180 ( .A(u5_mult_79_CLA_CARRY[45]), .ZN(
        u5_mult_79_FS_1_n66) );
  INV_X4 u5_mult_79_FS_1_U179 ( .A(u5_mult_79_n243), .ZN(u5_mult_79_FS_1_n67)
         );
  NAND2_X2 u5_mult_79_FS_1_U178 ( .A1(u5_mult_79_FS_1_n66), .A2(
        u5_mult_79_FS_1_n67), .ZN(u5_mult_79_FS_1_n41) );
  INV_X4 u5_mult_79_FS_1_U177 ( .A(u5_mult_79_FS_1_n41), .ZN(
        u5_mult_79_FS_1_n64) );
  NAND2_X2 u5_mult_79_FS_1_U176 ( .A1(u5_mult_79_CLA_CARRY[45]), .A2(
        u5_mult_79_n243), .ZN(u5_mult_79_FS_1_n65) );
  INV_X4 u5_mult_79_FS_1_U175 ( .A(u5_mult_79_FS_1_n65), .ZN(
        u5_mult_79_FS_1_n46) );
  NOR2_X4 u5_mult_79_FS_1_U174 ( .A1(u5_mult_79_FS_1_n64), .A2(
        u5_mult_79_FS_1_n46), .ZN(u5_mult_79_FS_1_n63) );
  XNOR2_X2 u5_mult_79_FS_1_U173 ( .A(u5_mult_79_FS_1_n62), .B(
        u5_mult_79_FS_1_n63), .ZN(u5_N46) );
  NAND2_X2 u5_mult_79_FS_1_U172 ( .A1(u5_mult_79_FS_1_n21), .A2(
        u5_mult_79_FS_1_n41), .ZN(u5_mult_79_FS_1_n50) );
  NAND2_X2 u5_mult_79_FS_1_U171 ( .A1(u5_mult_79_FS_1_n40), .A2(
        u5_mult_79_FS_1_n41), .ZN(u5_mult_79_FS_1_n43) );
  AOI21_X4 u5_mult_79_FS_1_U170 ( .B1(u5_mult_79_FS_1_n45), .B2(
        u5_mult_79_FS_1_n41), .A(u5_mult_79_FS_1_n46), .ZN(u5_mult_79_FS_1_n44) );
  NAND2_X2 u5_mult_79_FS_1_U169 ( .A1(u5_mult_79_FS_1_n40), .A2(
        u5_mult_79_FS_1_n41), .ZN(u5_mult_79_FS_1_n39) );
  XNOR2_X2 u5_mult_79_FS_1_U168 ( .A(u5_mult_79_FS_1_n33), .B(
        u5_mult_79_FS_1_n32), .ZN(u5_N47) );
  NAND2_X1 u5_mult_79_FS_1_U167 ( .A1(u5_mult_79_FS_1_n4), .A2(
        u5_mult_79_CLA_CARRY[25]), .ZN(u5_mult_79_FS_1_n276) );
  NAND2_X1 u5_mult_79_FS_1_U166 ( .A1(u5_mult_79_CLA_CARRY[27]), .A2(
        u5_mult_79_CLA_SUM[28]), .ZN(u5_mult_79_FS_1_n279) );
  NOR2_X1 u5_mult_79_FS_1_U165 ( .A1(u5_mult_79_FS_1_n61), .A2(
        u5_mult_79_FS_1_n2), .ZN(u5_mult_79_FS_1_n59) );
  OAI21_X1 u5_mult_79_FS_1_U164 ( .B1(u5_mult_79_FS_1_n274), .B2(
        u5_mult_79_FS_1_n260), .A(u5_mult_79_FS_1_n213), .ZN(
        u5_mult_79_FS_1_n250) );
  NOR2_X1 u5_mult_79_FS_1_U163 ( .A1(u5_mult_79_FS_1_n270), .A2(
        u5_mult_79_FS_1_n258), .ZN(u5_mult_79_FS_1_n278) );
  NAND2_X1 u5_mult_79_FS_1_U162 ( .A1(u5_mult_79_FS_1_n244), .A2(
        u5_mult_79_FS_1_n215), .ZN(u5_mult_79_FS_1_n243) );
  NOR2_X2 u5_mult_79_FS_1_U161 ( .A1(u5_mult_79_FS_1_n108), .A2(
        u5_mult_79_FS_1_n2), .ZN(u5_mult_79_FS_1_n191) );
  NOR2_X1 u5_mult_79_FS_1_U160 ( .A1(u5_mult_79_FS_1_n1), .A2(
        u5_mult_79_FS_1_n276), .ZN(u5_mult_79_FS_1_n275) );
  OAI21_X1 u5_mult_79_FS_1_U159 ( .B1(u5_mult_79_FS_1_n1), .B2(
        u5_mult_79_FS_1_n250), .A(u5_mult_79_FS_1_n251), .ZN(
        u5_mult_79_FS_1_n249) );
  NAND2_X4 u5_mult_79_FS_1_U158 ( .A1(u5_mult_79_n1718), .A2(
        u5_mult_79_CLA_CARRY[26]), .ZN(u5_mult_79_FS_1_n215) );
  NAND3_X2 u5_mult_79_FS_1_U157 ( .A1(u5_mult_79_FS_1_n228), .A2(
        u5_mult_79_FS_1_n229), .A3(u5_mult_79_FS_1_n220), .ZN(
        u5_mult_79_FS_1_n237) );
  INV_X4 u5_mult_79_FS_1_U156 ( .A(u5_mult_79_n245), .ZN(u5_mult_79_FS_1_n32)
         );
  NOR2_X4 u5_mult_79_FS_1_U155 ( .A1(u5_mult_79_FS_1_n162), .A2(
        u5_mult_79_FS_1_n163), .ZN(u5_mult_79_FS_1_n153) );
  NAND2_X1 u5_mult_79_FS_1_U154 ( .A1(u5_mult_79_FS_1_n242), .A2(
        u5_mult_79_FS_1_n215), .ZN(u5_mult_79_FS_1_n281) );
  INV_X8 u5_mult_79_FS_1_U153 ( .A(u5_mult_79_FS_1_n24), .ZN(
        u5_mult_79_FS_1_n56) );
  NAND2_X4 u5_mult_79_FS_1_U152 ( .A1(u5_mult_79_FS_1_n239), .A2(
        u5_mult_79_FS_1_n238), .ZN(u5_mult_79_FS_1_n211) );
  NAND2_X4 u5_mult_79_FS_1_U151 ( .A1(u5_mult_79_FS_1_n262), .A2(
        u5_mult_79_FS_1_n263), .ZN(u5_mult_79_FS_1_n209) );
  INV_X8 u5_mult_79_FS_1_U150 ( .A(u5_mult_79_FS_1_n266), .ZN(
        u5_mult_79_FS_1_n254) );
  NAND2_X4 u5_mult_79_FS_1_U149 ( .A1(u5_mult_79_FS_1_n232), .A2(
        u5_mult_79_FS_1_n233), .ZN(u5_mult_79_FS_1_n199) );
  NAND2_X4 u5_mult_79_FS_1_U148 ( .A1(u5_mult_79_FS_1_n216), .A2(
        u5_mult_79_FS_1_n55), .ZN(u5_mult_79_FS_1_n58) );
  INV_X8 u5_mult_79_FS_1_U147 ( .A(u5_mult_79_FS_1_n58), .ZN(
        u5_mult_79_FS_1_n108) );
  NAND2_X4 u5_mult_79_FS_1_U146 ( .A1(u5_mult_79_FS_1_n246), .A2(
        u5_mult_79_FS_1_n247), .ZN(u5_mult_79_FS_1_n210) );
  NAND2_X4 u5_mult_79_FS_1_U145 ( .A1(u5_mult_79_FS_1_n267), .A2(
        u5_mult_79_FS_1_n268), .ZN(u5_mult_79_FS_1_n266) );
  INV_X16 u5_mult_79_FS_1_U144 ( .A(u5_mult_79_FS_1_n217), .ZN(
        u5_mult_79_FS_1_n55) );
  NAND2_X4 u5_mult_79_FS_1_U143 ( .A1(u5_mult_79_FS_1_n55), .A2(
        u5_mult_79_FS_1_n6), .ZN(u5_mult_79_FS_1_n54) );
  INV_X8 u5_mult_79_FS_1_U142 ( .A(u5_mult_79_FS_1_n211), .ZN(
        u5_mult_79_FS_1_n204) );
  NAND2_X1 u5_mult_79_FS_1_U141 ( .A1(u5_mult_79_FS_1_n58), .A2(
        u5_mult_79_FS_1_n59), .ZN(u5_mult_79_FS_1_n47) );
  NAND2_X4 u5_mult_79_FS_1_U140 ( .A1(u5_mult_79_FS_1_n197), .A2(
        u5_mult_79_FS_1_n55), .ZN(u5_mult_79_FS_1_n106) );
  NAND2_X1 u5_mult_79_FS_1_U139 ( .A1(u5_mult_79_FS_1_n211), .A2(
        u5_mult_79_FS_1_n199), .ZN(u5_mult_79_FS_1_n207) );
  NAND3_X2 u5_mult_79_FS_1_U138 ( .A1(u5_mult_79_FS_1_n198), .A2(
        u5_mult_79_FS_1_n199), .A3(u5_mult_79_FS_1_n200), .ZN(
        u5_mult_79_FS_1_n53) );
  NAND2_X1 u5_mult_79_FS_1_U137 ( .A1(u5_mult_79_FS_1_n201), .A2(
        u5_mult_79_FS_1_n199), .ZN(u5_mult_79_FS_1_n231) );
  NAND2_X2 u5_mult_79_FS_1_U136 ( .A1(u5_mult_79_n230), .A2(
        u5_mult_79_CLA_SUM[33]), .ZN(u5_mult_79_FS_1_n201) );
  NAND2_X4 u5_mult_79_FS_1_U135 ( .A1(u5_mult_79_FS_1_n186), .A2(
        u5_mult_79_FS_1_n187), .ZN(u5_mult_79_FS_1_n182) );
  NAND2_X4 u5_mult_79_FS_1_U134 ( .A1(u5_mult_79_FS_1_n170), .A2(
        u5_mult_79_FS_1_n171), .ZN(u5_mult_79_FS_1_n155) );
  NAND2_X1 u5_mult_79_FS_1_U133 ( .A1(u5_mult_79_FS_1_n211), .A2(
        u5_mult_79_FS_1_n202), .ZN(u5_mult_79_FS_1_n234) );
  NAND2_X4 u5_mult_79_FS_1_U132 ( .A1(u5_mult_79_FS_1_n105), .A2(
        u5_mult_79_FS_1_n23), .ZN(u5_mult_79_FS_1_n104) );
  NAND2_X4 u5_mult_79_FS_1_U131 ( .A1(u5_mult_79_FS_1_n183), .A2(
        u5_mult_79_FS_1_n184), .ZN(u5_mult_79_FS_1_n170) );
  INV_X2 u5_mult_79_FS_1_U130 ( .A(u5_mult_79_FS_1_n210), .ZN(
        u5_mult_79_FS_1_n230) );
  NAND2_X1 u5_mult_79_FS_1_U129 ( .A1(u5_mult_79_FS_1_n203), .A2(
        u5_mult_79_FS_1_n210), .ZN(u5_mult_79_FS_1_n240) );
  NOR2_X1 u5_mult_79_FS_1_U128 ( .A1(u5_mult_79_FS_1_n38), .A2(
        u5_mult_79_FS_1_n39), .ZN(u5_mult_79_FS_1_n37) );
  AOI21_X4 u5_mult_79_FS_1_U127 ( .B1(u5_mult_79_FS_1_n40), .B2(
        u5_mult_79_FS_1_n68), .A(u5_mult_79_FS_1_n45), .ZN(u5_mult_79_FS_1_n62) );
  AOI21_X4 u5_mult_79_FS_1_U126 ( .B1(u5_mult_79_FS_1_n72), .B2(
        u5_mult_79_FS_1_n68), .A(u5_mult_79_FS_1_n70), .ZN(u5_mult_79_FS_1_n73) );
  AOI21_X4 u5_mult_79_FS_1_U125 ( .B1(u5_mult_79_FS_1_n84), .B2(
        u5_mult_79_FS_1_n68), .A(u5_mult_79_FS_1_n79), .ZN(u5_mult_79_FS_1_n85) );
  NOR2_X1 u5_mult_79_FS_1_U124 ( .A1(u5_mult_79_FS_1_n97), .A2(
        u5_mult_79_FS_1_n98), .ZN(u5_mult_79_FS_1_n154) );
  INV_X2 u5_mult_79_FS_1_U123 ( .A(u5_mult_79_FS_1_n181), .ZN(
        u5_mult_79_FS_1_n188) );
  NOR2_X1 u5_mult_79_FS_1_U122 ( .A1(u5_mult_79_FS_1_n189), .A2(
        u5_mult_79_FS_1_n181), .ZN(u5_mult_79_FS_1_n221) );
  INV_X4 u5_mult_79_FS_1_U121 ( .A(u5_mult_79_FS_1_n28), .ZN(
        u5_mult_79_FS_1_n29) );
  NOR2_X4 u5_mult_79_FS_1_U120 ( .A1(u5_mult_79_FS_1_n206), .A2(
        u5_mult_79_FS_1_n29), .ZN(u5_mult_79_FS_1_n60) );
  NOR2_X2 u5_mult_79_FS_1_U119 ( .A1(u5_mult_79_FS_1_n207), .A2(
        u5_mult_79_FS_1_n208), .ZN(u5_mult_79_FS_1_n28) );
  INV_X4 u5_mult_79_FS_1_U118 ( .A(u5_mult_79_FS_1_n105), .ZN(
        u5_mult_79_FS_1_n205) );
  NAND2_X4 u5_mult_79_FS_1_U117 ( .A1(u5_mult_79_FS_1_n160), .A2(
        u5_mult_79_FS_1_n158), .ZN(u5_mult_79_FS_1_n51) );
  NAND3_X1 u5_mult_79_FS_1_U116 ( .A1(u5_mult_79_FS_1_n23), .A2(
        u5_mult_79_FS_1_n105), .A3(u5_mult_79_FS_1_n54), .ZN(
        u5_mult_79_FS_1_n48) );
  NAND2_X4 u5_mult_79_FS_1_U115 ( .A1(u5_mult_79_FS_1_n148), .A2(
        u5_mult_79_FS_1_n149), .ZN(u5_mult_79_FS_1_n147) );
  NAND2_X1 u5_mult_79_FS_1_U114 ( .A1(u5_mult_79_n238), .A2(
        u5_mult_79_FS_1_n16), .ZN(u5_mult_79_FS_1_n253) );
  NAND2_X2 u5_mult_79_FS_1_U113 ( .A1(u5_mult_79_CLA_CARRY[25]), .A2(
        u5_mult_79_n1449), .ZN(u5_mult_79_FS_1_n214) );
  NOR2_X1 u5_mult_79_FS_1_U112 ( .A1(u5_mult_79_FS_1_n254), .A2(
        u5_mult_79_FS_1_n197), .ZN(u5_mult_79_FS_1_n265) );
  INV_X2 u5_mult_79_FS_1_U111 ( .A(u5_mult_79_FS_1_n173), .ZN(
        u5_mult_79_FS_1_n169) );
  AOI21_X2 u5_mult_79_FS_1_U110 ( .B1(u5_mult_79_FS_1_n173), .B2(
        u5_mult_79_FS_1_n188), .A(u5_mult_79_FS_1_n189), .ZN(
        u5_mult_79_FS_1_n185) );
  INV_X8 u5_mult_79_FS_1_U109 ( .A(u5_mult_79_CLA_SUM[39]), .ZN(
        u5_mult_79_FS_1_n149) );
  NAND2_X4 u5_mult_79_FS_1_U108 ( .A1(u5_mult_79_FS_1_n122), .A2(
        u5_mult_79_FS_1_n118), .ZN(u5_mult_79_FS_1_n121) );
  NOR2_X1 u5_mult_79_FS_1_U107 ( .A1(u5_mult_79_FS_1_n133), .A2(
        u5_mult_79_FS_1_n135), .ZN(u5_mult_79_FS_1_n142) );
  NOR2_X1 u5_mult_79_FS_1_U106 ( .A1(u5_mult_79_FS_1_n13), .A2(
        u5_mult_79_FS_1_n135), .ZN(u5_mult_79_FS_1_n151) );
  AOI21_X2 u5_mult_79_FS_1_U105 ( .B1(u5_mult_79_FS_1_n122), .B2(
        u5_mult_79_FS_1_n117), .A(u5_mult_79_FS_1_n128), .ZN(
        u5_mult_79_FS_1_n123) );
  OAI21_X1 u5_mult_79_FS_1_U104 ( .B1(u5_mult_79_FS_1_n133), .B2(
        u5_mult_79_FS_1_n134), .A(u5_mult_79_FS_1_n144), .ZN(
        u5_mult_79_FS_1_n143) );
  NOR2_X4 u5_mult_79_FS_1_U103 ( .A1(u5_mult_79_FS_1_n254), .A2(
        u5_mult_79_FS_1_n255), .ZN(u5_mult_79_FS_1_n196) );
  AOI21_X2 u5_mult_79_FS_1_U102 ( .B1(u5_mult_79_FS_1_n142), .B2(
        u5_mult_79_FS_1_n117), .A(u5_mult_79_FS_1_n143), .ZN(
        u5_mult_79_FS_1_n136) );
  AOI21_X2 u5_mult_79_FS_1_U101 ( .B1(u5_mult_79_FS_1_n150), .B2(
        u5_mult_79_FS_1_n117), .A(u5_mult_79_FS_1_n13), .ZN(
        u5_mult_79_FS_1_n145) );
  AOI21_X2 u5_mult_79_FS_1_U100 ( .B1(u5_mult_79_FS_1_n102), .B2(
        u5_mult_79_FS_1_n117), .A(u5_mult_79_FS_1_n20), .ZN(
        u5_mult_79_FS_1_n111) );
  NAND2_X1 u5_mult_79_FS_1_U99 ( .A1(u5_mult_79_FS_1_n17), .A2(
        u5_mult_79_FS_1_n120), .ZN(u5_mult_79_FS_1_n128) );
  NAND2_X4 u5_mult_79_FS_1_U98 ( .A1(u5_mult_79_FS_1_n176), .A2(
        u5_mult_79_FS_1_n177), .ZN(u5_mult_79_FS_1_n171) );
  AND2_X4 u5_mult_79_FS_1_U97 ( .A1(u5_mult_79_FS_1_n119), .A2(
        u5_mult_79_FS_1_n120), .ZN(u5_mult_79_FS_1_n27) );
  AOI21_X4 u5_mult_79_FS_1_U96 ( .B1(u5_mult_79_FS_1_n17), .B2(
        u5_mult_79_FS_1_n27), .A(u5_mult_79_FS_1_n26), .ZN(u5_mult_79_FS_1_n25) );
  NAND2_X2 u5_mult_79_FS_1_U95 ( .A1(u5_mult_79_FS_1_n34), .A2(
        u5_mult_79_FS_1_n35), .ZN(u5_mult_79_FS_1_n33) );
  INV_X2 u5_mult_79_FS_1_U94 ( .A(u5_mult_79_FS_1_n170), .ZN(
        u5_mult_79_FS_1_n178) );
  OAI21_X2 u5_mult_79_FS_1_U93 ( .B1(u5_mult_79_FS_1_n7), .B2(
        u5_mult_79_FS_1_n241), .A(u5_mult_79_FS_1_n209), .ZN(
        u5_mult_79_FS_1_n229) );
  NAND2_X1 u5_mult_79_FS_1_U92 ( .A1(u5_mult_79_FS_1_n209), .A2(
        u5_mult_79_FS_1_n220), .ZN(u5_mult_79_FS_1_n248) );
  OAI21_X2 u5_mult_79_FS_1_U91 ( .B1(u5_mult_79_FS_1_n47), .B2(
        u5_mult_79_FS_1_n48), .A(u5_mult_79_FS_1_n49), .ZN(u5_mult_79_FS_1_n34) );
  NOR2_X4 u5_mult_79_FS_1_U90 ( .A1(u5_mult_79_FS_1_n180), .A2(
        u5_mult_79_FS_1_n181), .ZN(u5_mult_79_FS_1_n172) );
  INV_X4 u5_mult_79_FS_1_U89 ( .A(u5_mult_79_FS_1_n30), .ZN(
        u5_mult_79_FS_1_n31) );
  INV_X1 u5_mult_79_FS_1_U88 ( .A(u5_mult_79_FS_1_n182), .ZN(
        u5_mult_79_FS_1_n180) );
  NAND2_X4 u5_mult_79_FS_1_U87 ( .A1(u5_mult_79_FS_1_n106), .A2(
        u5_mult_79_FS_1_n54), .ZN(u5_mult_79_FS_1_n30) );
  NAND2_X1 u5_mult_79_FS_1_U86 ( .A1(u5_mult_79_FS_1_n156), .A2(
        u5_mult_79_FS_1_n171), .ZN(u5_mult_79_FS_1_n175) );
  INV_X8 u5_mult_79_FS_1_U85 ( .A(u5_mult_79_FS_1_n245), .ZN(
        u5_mult_79_FS_1_n57) );
  INV_X8 u5_mult_79_FS_1_U84 ( .A(u5_mult_79_FS_1_n147), .ZN(
        u5_mult_79_FS_1_n133) );
  NAND2_X2 u5_mult_79_FS_1_U83 ( .A1(u5_mult_79_FS_1_n214), .A2(
        u5_mult_79_FS_1_n215), .ZN(u5_mult_79_FS_1_n212) );
  INV_X8 u5_mult_79_FS_1_U82 ( .A(u5_mult_79_FS_1_n194), .ZN(
        u5_mult_79_FS_1_n23) );
  INV_X8 u5_mult_79_FS_1_U81 ( .A(u5_mult_79_FS_1_n100), .ZN(
        u5_mult_79_FS_1_n113) );
  NAND2_X4 u5_mult_79_FS_1_U80 ( .A1(u5_mult_79_FS_1_n115), .A2(
        u5_mult_79_FS_1_n116), .ZN(u5_mult_79_FS_1_n100) );
  NOR2_X4 u5_mult_79_FS_1_U79 ( .A1(u5_mult_79_FS_1_n121), .A2(
        u5_mult_79_FS_1_n113), .ZN(u5_mult_79_FS_1_n22) );
  NOR2_X2 u5_mult_79_FS_1_U78 ( .A1(u5_mult_79_FS_1_n121), .A2(
        u5_mult_79_FS_1_n113), .ZN(u5_mult_79_FS_1_n21) );
  BUF_X8 u5_mult_79_FS_1_U77 ( .A(u5_mult_79_FS_1_n25), .Z(u5_mult_79_FS_1_n20) );
  OAI21_X1 u5_mult_79_FS_1_U76 ( .B1(u5_mult_79_FS_1_n25), .B2(
        u5_mult_79_FS_1_n99), .A(u5_mult_79_FS_1_n100), .ZN(
        u5_mult_79_FS_1_n19) );
  BUF_X16 u5_mult_79_FS_1_U75 ( .A(u5_mult_79_CLA_SUM[38]), .Z(
        u5_mult_79_FS_1_n18) );
  INV_X1 u5_mult_79_FS_1_U74 ( .A(u5_mult_79_FS_1_n135), .ZN(
        u5_mult_79_FS_1_n150) );
  OAI21_X2 u5_mult_79_FS_1_U73 ( .B1(u5_mult_79_FS_1_n19), .B2(
        u5_mult_79_FS_1_n43), .A(u5_mult_79_FS_1_n44), .ZN(u5_mult_79_FS_1_n36) );
  NOR2_X2 u5_mult_79_FS_1_U72 ( .A1(u5_mult_79_FS_1_n37), .A2(
        u5_mult_79_FS_1_n36), .ZN(u5_mult_79_FS_1_n35) );
  NOR2_X2 u5_mult_79_FS_1_U71 ( .A1(u5_mult_79_FS_1_n204), .A2(
        u5_mult_79_FS_1_n230), .ZN(u5_mult_79_FS_1_n225) );
  INV_X8 u5_mult_79_FS_1_U70 ( .A(u5_mult_79_CLA_SUM[29]), .ZN(
        u5_mult_79_FS_1_n268) );
  INV_X1 u5_mult_79_FS_1_U69 ( .A(u5_mult_79_FS_1_n268), .ZN(
        u5_mult_79_FS_1_n16) );
  XNOR2_X2 u5_mult_79_FS_1_U68 ( .A(u5_mult_79_FS_1_n173), .B(
        u5_mult_79_FS_1_n190), .ZN(u5_N34) );
  INV_X2 u5_mult_79_FS_1_U67 ( .A(u5_mult_79_FS_1_n237), .ZN(
        u5_mult_79_FS_1_n236) );
  XNOR2_X2 u5_mult_79_FS_1_U66 ( .A(u5_mult_79_FS_1_n237), .B(
        u5_mult_79_FS_1_n240), .ZN(u5_N31) );
  NAND3_X2 u5_mult_79_FS_1_U65 ( .A1(u5_mult_79_FS_1_n56), .A2(
        u5_mult_79_FS_1_n8), .A3(u5_mult_79_FS_1_n57), .ZN(
        u5_mult_79_FS_1_n228) );
  AOI21_X2 u5_mult_79_FS_1_U64 ( .B1(u5_mult_79_FS_1_n269), .B2(
        u5_mult_79_FS_1_n257), .A(u5_mult_79_FS_1_n270), .ZN(
        u5_mult_79_FS_1_n264) );
  NAND2_X2 u5_mult_79_FS_1_U63 ( .A1(u5_mult_79_CLA_SUM[28]), .A2(
        u5_mult_79_CLA_CARRY[27]), .ZN(u5_mult_79_FS_1_n255) );
  NOR2_X2 u5_mult_79_FS_1_U62 ( .A1(u5_mult_79_FS_1_n275), .A2(
        u5_mult_79_FS_1_n274), .ZN(u5_mult_79_FS_1_n273) );
  INV_X2 u5_mult_79_FS_1_U61 ( .A(u5_mult_79_FS_1_n277), .ZN(
        u5_mult_79_FS_1_n283) );
  NAND3_X2 u5_mult_79_FS_1_U60 ( .A1(u5_mult_79_FS_1_n256), .A2(
        u5_mult_79_FS_1_n242), .A3(u5_mult_79_FS_1_n257), .ZN(
        u5_mult_79_FS_1_n245) );
  AND2_X2 u5_mult_79_FS_1_U59 ( .A1(u5_mult_79_FS_1_n284), .A2(
        u5_mult_79_FS_1_n285), .ZN(u5_mult_79_FS_1_n15) );
  AND2_X2 u5_mult_79_FS_1_U58 ( .A1(u5_mult_79_FS_1_n183), .A2(
        u5_mult_79_FS_1_n182), .ZN(u5_mult_79_FS_1_n14) );
  INV_X4 u5_mult_79_FS_1_U57 ( .A(u5_mult_79_FS_1_n215), .ZN(
        u5_mult_79_FS_1_n274) );
  INV_X2 u5_mult_79_FS_1_U56 ( .A(u5_mult_79_FS_1_n118), .ZN(
        u5_mult_79_FS_1_n26) );
  AND2_X2 u5_mult_79_FS_1_U55 ( .A1(u5_mult_79_CLA_CARRY[37]), .A2(
        u5_mult_79_FS_1_n18), .ZN(u5_mult_79_FS_1_n13) );
  AND2_X4 u5_mult_79_FS_1_U54 ( .A1(u5_mult_79_CLA_CARRY[44]), .A2(
        u5_mult_79_n242), .ZN(u5_mult_79_FS_1_n11) );
  NOR2_X2 u5_mult_79_FS_1_U53 ( .A1(u5_mult_79_FS_1_n133), .A2(
        u5_mult_79_FS_1_n129), .ZN(u5_mult_79_FS_1_n146) );
  INV_X4 u5_mult_79_FS_1_U52 ( .A(u5_mult_79_FS_1_n205), .ZN(
        u5_mult_79_FS_1_n192) );
  NOR2_X2 u5_mult_79_FS_1_U51 ( .A1(u5_mult_79_FS_1_n132), .A2(
        u5_mult_79_FS_1_n133), .ZN(u5_mult_79_FS_1_n131) );
  NAND2_X1 u5_mult_79_FS_1_U50 ( .A1(u5_mult_79_FS_1_n159), .A2(
        u5_mult_79_FS_1_n158), .ZN(u5_mult_79_FS_1_n166) );
  OR2_X1 u5_mult_79_FS_1_U49 ( .A1(u5_mult_79_FS_1_n277), .A2(
        u5_mult_79_FS_1_n259), .ZN(u5_mult_79_FS_1_n12) );
  INV_X8 u5_mult_79_FS_1_U48 ( .A(u5_mult_79_CLA_SUM[35]), .ZN(
        u5_mult_79_FS_1_n187) );
  NOR3_X2 u5_mult_79_FS_1_U47 ( .A1(u5_mult_79_FS_1_n50), .A2(
        u5_mult_79_FS_1_n51), .A3(u5_mult_79_FS_1_n52), .ZN(
        u5_mult_79_FS_1_n49) );
  INV_X2 u5_mult_79_FS_1_U46 ( .A(u5_mult_79_FS_1_n9), .ZN(u5_mult_79_FS_1_n10) );
  INV_X1 u5_mult_79_FS_1_U45 ( .A(u5_mult_79_FS_1_n155), .ZN(
        u5_mult_79_FS_1_n9) );
  INV_X8 u5_mult_79_FS_1_U44 ( .A(u5_mult_79_CLA_SUM[33]), .ZN(
        u5_mult_79_FS_1_n233) );
  NAND2_X4 u5_mult_79_FS_1_U43 ( .A1(u5_mult_79_FS_1_n21), .A2(
        u5_mult_79_FS_1_n101), .ZN(u5_mult_79_FS_1_n93) );
  NAND2_X4 u5_mult_79_FS_1_U42 ( .A1(u5_mult_79_FS_1_n167), .A2(
        u5_mult_79_FS_1_n168), .ZN(u5_mult_79_FS_1_n158) );
  INV_X1 u5_mult_79_FS_1_U41 ( .A(u5_mult_79_FS_1_n117), .ZN(
        u5_mult_79_FS_1_n152) );
  NAND2_X2 u5_mult_79_FS_1_U40 ( .A1(u5_mult_79_FS_1_n209), .A2(
        u5_mult_79_FS_1_n210), .ZN(u5_mult_79_FS_1_n208) );
  NAND2_X4 u5_mult_79_FS_1_U39 ( .A1(u5_mult_79_FS_1_n164), .A2(
        u5_mult_79_FS_1_n105), .ZN(u5_mult_79_FS_1_n162) );
  NAND3_X2 u5_mult_79_FS_1_U38 ( .A1(u5_mult_79_FS_1_n54), .A2(
        u5_mult_79_FS_1_n106), .A3(u5_mult_79_FS_1_n53), .ZN(
        u5_mult_79_FS_1_n163) );
  NAND2_X4 u5_mult_79_FS_1_U37 ( .A1(u5_mult_79_n232), .A2(
        u5_mult_79_CLA_SUM[31]), .ZN(u5_mult_79_FS_1_n203) );
  NAND2_X4 u5_mult_79_FS_1_U36 ( .A1(u5_mult_79_FS_1_n107), .A2(
        u5_mult_79_FS_1_n31), .ZN(u5_mult_79_FS_1_n103) );
  NAND2_X4 u5_mult_79_FS_1_U35 ( .A1(u5_mult_79_FS_1_n262), .A2(
        u5_mult_79_FS_1_n263), .ZN(u5_mult_79_FS_1_n8) );
  INV_X4 u5_mult_79_FS_1_U34 ( .A(u5_mult_79_FS_1_n106), .ZN(
        u5_mult_79_FS_1_n61) );
  AOI21_X2 u5_mult_79_FS_1_U33 ( .B1(u5_mult_79_FS_1_n225), .B2(
        u5_mult_79_FS_1_n226), .A(u5_mult_79_FS_1_n227), .ZN(
        u5_mult_79_FS_1_n224) );
  OAI21_X4 u5_mult_79_FS_1_U32 ( .B1(u5_mult_79_FS_1_n129), .B2(
        u5_mult_79_FS_1_n130), .A(u5_mult_79_FS_1_n131), .ZN(
        u5_mult_79_FS_1_n17) );
  AND3_X4 u5_mult_79_FS_1_U31 ( .A1(u5_mult_79_FS_1_n243), .A2(
        u5_mult_79_FS_1_n242), .A3(u5_mult_79_FS_1_n213), .ZN(
        u5_mult_79_FS_1_n7) );
  OAI21_X2 u5_mult_79_FS_1_U30 ( .B1(u5_mult_79_FS_1_n236), .B2(
        u5_mult_79_FS_1_n230), .A(u5_mult_79_FS_1_n203), .ZN(
        u5_mult_79_FS_1_n235) );
  INV_X8 u5_mult_79_FS_1_U29 ( .A(u5_mult_79_FS_1_n196), .ZN(
        u5_mult_79_FS_1_n252) );
  INV_X4 u5_mult_79_FS_1_U28 ( .A(u5_mult_79_FS_1_n252), .ZN(
        u5_mult_79_FS_1_n6) );
  OAI21_X4 u5_mult_79_FS_1_U27 ( .B1(u5_mult_79_FS_1_n272), .B2(
        u5_mult_79_FS_1_n12), .A(u5_mult_79_FS_1_n273), .ZN(
        u5_mult_79_FS_1_n269) );
  OAI21_X2 u5_mult_79_FS_1_U26 ( .B1(u5_mult_79_FS_1_n272), .B2(
        u5_mult_79_FS_1_n5), .A(u5_mult_79_FS_1_n276), .ZN(
        u5_mult_79_FS_1_n280) );
  NAND2_X1 u5_mult_79_FS_1_U25 ( .A1(u5_mult_79_FS_1_n276), .A2(
        u5_mult_79_FS_1_n283), .ZN(u5_mult_79_FS_1_n282) );
  NOR2_X4 u5_mult_79_FS_1_U24 ( .A1(u5_mult_79_n1449), .A2(
        u5_mult_79_CLA_CARRY[25]), .ZN(u5_mult_79_FS_1_n277) );
  INV_X2 u5_mult_79_FS_1_U23 ( .A(u5_mult_79_FS_1_n283), .ZN(
        u5_mult_79_FS_1_n5) );
  NAND3_X4 u5_mult_79_FS_1_U22 ( .A1(u5_mult_79_FS_1_n55), .A2(
        u5_mult_79_FS_1_n56), .A3(u5_mult_79_FS_1_n57), .ZN(
        u5_mult_79_FS_1_n105) );
  INV_X8 u5_mult_79_FS_1_U21 ( .A(u5_mult_79_FS_1_n56), .ZN(
        u5_mult_79_FS_1_n272) );
  NAND2_X4 u5_mult_79_FS_1_U20 ( .A1(u5_mult_79_CLA_CARRY[24]), .A2(
        u5_mult_79_CLA_SUM[25]), .ZN(u5_mult_79_FS_1_n24) );
  INV_X1 u5_mult_79_FS_1_U19 ( .A(u5_mult_79_CLA_SUM[25]), .ZN(
        u5_mult_79_FS_1_n285) );
  NOR2_X2 u5_mult_79_FS_1_U18 ( .A1(u5_mult_79_FS_1_n15), .A2(
        u5_mult_79_FS_1_n56), .ZN(u5_N25) );
  NOR2_X4 u5_mult_79_FS_1_U17 ( .A1(u5_mult_79_FS_1_n2), .A2(
        u5_mult_79_FS_1_n108), .ZN(u5_mult_79_FS_1_n107) );
  XNOR2_X2 u5_mult_79_FS_1_U16 ( .A(u5_mult_79_FS_1_n68), .B(
        u5_mult_79_FS_1_n91), .ZN(u5_N43) );
  INV_X4 u5_mult_79_FS_1_U15 ( .A(u5_mult_79_FS_1_n38), .ZN(
        u5_mult_79_FS_1_n96) );
  NOR2_X4 u5_mult_79_FS_1_U14 ( .A1(u5_mult_79_FS_1_n277), .A2(
        u5_mult_79_FS_1_n254), .ZN(u5_mult_79_FS_1_n256) );
  INV_X8 u5_mult_79_FS_1_U13 ( .A(u5_mult_79_FS_1_n259), .ZN(
        u5_mult_79_FS_1_n242) );
  INV_X4 u5_mult_79_FS_1_U12 ( .A(u5_mult_79_FS_1_n54), .ZN(
        u5_mult_79_FS_1_n195) );
  INV_X2 u5_mult_79_FS_1_U11 ( .A(u5_mult_79_FS_1_n121), .ZN(
        u5_mult_79_FS_1_n102) );
  NAND4_X2 u5_mult_79_FS_1_U10 ( .A1(u5_mult_79_FS_1_n220), .A2(
        u5_mult_79_FS_1_n203), .A3(u5_mult_79_FS_1_n228), .A4(
        u5_mult_79_FS_1_n229), .ZN(u5_mult_79_FS_1_n226) );
  NAND2_X1 u5_mult_79_FS_1_U9 ( .A1(u5_mult_79_CLA_CARRY[25]), .A2(
        u5_mult_79_n1449), .ZN(u5_mult_79_FS_1_n244) );
  INV_X2 u5_mult_79_FS_1_U8 ( .A(u5_mult_79_FS_1_n3), .ZN(u5_mult_79_FS_1_n4)
         );
  INV_X1 u5_mult_79_FS_1_U7 ( .A(u5_mult_79_n1449), .ZN(u5_mult_79_FS_1_n3) );
  NAND3_X4 u5_mult_79_FS_1_U6 ( .A1(u5_mult_79_FS_1_n213), .A2(
        u5_mult_79_FS_1_n242), .A3(u5_mult_79_FS_1_n212), .ZN(
        u5_mult_79_FS_1_n206) );
  NOR2_X4 u5_mult_79_FS_1_U5 ( .A1(u5_mult_79_FS_1_n206), .A2(
        u5_mult_79_FS_1_n29), .ZN(u5_mult_79_FS_1_n2) );
  AOI21_X1 u5_mult_79_FS_1_U4 ( .B1(u5_mult_79_FS_1_n56), .B2(
        u5_mult_79_FS_1_n57), .A(u5_mult_79_FS_1_n241), .ZN(
        u5_mult_79_FS_1_n251) );
  INV_X1 u5_mult_79_FS_1_U3 ( .A(u5_mult_79_FS_1_n242), .ZN(u5_mult_79_FS_1_n1) );
  INV_X1 u5_mult_79_FS_1_U2 ( .A(u5_mult_79_FS_1_n244), .ZN(
        u5_mult_79_FS_1_n260) );
  INV_X4 u4_add_395_U91 ( .A(u4_fract_out_0_), .ZN(u4_fract_out_pl1_0_) );
  NAND4_X2 u4_add_395_U90 ( .A1(u4_fract_out_3_), .A2(u4_fract_out_2_), .A3(
        u4_fract_out_1_), .A4(u4_fract_out_0_), .ZN(u4_add_395_n25) );
  INV_X4 u4_add_395_U89 ( .A(u4_add_395_n25), .ZN(u4_add_395_n21) );
  NAND2_X2 u4_add_395_U88 ( .A1(u4_fract_out_7_), .A2(u4_fract_out_6_), .ZN(
        u4_add_395_n67) );
  NAND2_X2 u4_add_395_U87 ( .A1(u4_fract_out_4_), .A2(u4_fract_out_5_), .ZN(
        u4_add_395_n68) );
  NAND2_X2 u4_add_395_U86 ( .A1(u4_add_395_n21), .A2(u4_add_395_n66), .ZN(
        u4_add_395_n13) );
  INV_X4 u4_add_395_U85 ( .A(u4_add_395_n13), .ZN(u4_add_395_n15) );
  XNOR2_X2 u4_add_395_U84 ( .A(u4_add_395_n3), .B(u4_add_395_n65), .ZN(
        u4_fract_out_pl1_10_) );
  XNOR2_X2 u4_add_395_U83 ( .A(u4_fract_out_11_), .B(u4_add_395_n64), .ZN(
        u4_fract_out_pl1_11_) );
  NAND2_X2 u4_add_395_U82 ( .A1(u4_add_395_n1), .A2(u4_add_395_n15), .ZN(
        u4_add_395_n63) );
  INV_X4 u4_add_395_U81 ( .A(u4_add_395_n63), .ZN(u4_add_395_n60) );
  INV_X4 u4_add_395_U80 ( .A(u4_fract_out_12_), .ZN(u4_add_395_n62) );
  XNOR2_X2 u4_add_395_U79 ( .A(u4_add_395_n60), .B(u4_add_395_n62), .ZN(
        u4_fract_out_pl1_12_) );
  NAND2_X2 u4_add_395_U78 ( .A1(u4_add_395_n60), .A2(u4_fract_out_12_), .ZN(
        u4_add_395_n61) );
  XNOR2_X2 u4_add_395_U77 ( .A(u4_add_395_n10), .B(u4_add_395_n61), .ZN(
        u4_fract_out_pl1_13_) );
  INV_X4 u4_add_395_U76 ( .A(u4_add_395_n59), .ZN(u4_add_395_n57) );
  XNOR2_X2 u4_add_395_U75 ( .A(u4_add_395_n57), .B(u4_add_395_n58), .ZN(
        u4_fract_out_pl1_14_) );
  NAND2_X2 u4_add_395_U74 ( .A1(u4_add_395_n57), .A2(u4_fract_out_14_), .ZN(
        u4_add_395_n56) );
  NAND2_X2 u4_add_395_U73 ( .A1(u4_fract_out_12_), .A2(u4_fract_out_13_), .ZN(
        u4_add_395_n54) );
  NAND3_X4 u4_add_395_U72 ( .A1(u4_add_395_n1), .A2(u4_add_395_n53), .A3(
        u4_add_395_n15), .ZN(u4_add_395_n42) );
  INV_X4 u4_add_395_U71 ( .A(u4_add_395_n42), .ZN(u4_add_395_n49) );
  XNOR2_X2 u4_add_395_U70 ( .A(u4_fract_out_17_), .B(u4_add_395_n52), .ZN(
        u4_fract_out_pl1_17_) );
  INV_X4 u4_add_395_U69 ( .A(u4_fract_out_17_), .ZN(u4_add_395_n51) );
  NAND2_X2 u4_add_395_U68 ( .A1(u4_add_395_n48), .A2(u4_add_395_n49), .ZN(
        u4_add_395_n47) );
  INV_X4 u4_add_395_U67 ( .A(u4_add_395_n47), .ZN(u4_add_395_n45) );
  INV_X4 u4_add_395_U66 ( .A(u4_fract_out_18_), .ZN(u4_add_395_n46) );
  XNOR2_X2 u4_add_395_U65 ( .A(u4_add_395_n45), .B(u4_add_395_n46), .ZN(
        u4_fract_out_pl1_18_) );
  NAND2_X2 u4_add_395_U64 ( .A1(u4_add_395_n45), .A2(u4_fract_out_18_), .ZN(
        u4_add_395_n44) );
  NOR2_X4 u4_add_395_U63 ( .A1(u4_add_395_n42), .A2(u4_add_395_n43), .ZN(
        u4_add_395_n39) );
  NAND3_X4 u4_add_395_U62 ( .A1(u4_fract_out_12_), .A2(u4_fract_out_13_), .A3(
        u4_fract_out_14_), .ZN(u4_add_395_n34) );
  NAND3_X4 u4_add_395_U61 ( .A1(u4_fract_out_8_), .A2(u4_fract_out_6_), .A3(
        u4_fract_out_7_), .ZN(u4_add_395_n32) );
  NAND3_X4 u4_add_395_U60 ( .A1(u4_fract_out_3_), .A2(u4_fract_out_5_), .A3(
        u4_fract_out_4_), .ZN(u4_add_395_n31) );
  NAND2_X2 u4_add_395_U59 ( .A1(u4_fract_out_1_), .A2(u4_fract_out_0_), .ZN(
        u4_add_395_n29) );
  XNOR2_X2 u4_add_395_U58 ( .A(u4_fract_out_2_), .B(u4_add_395_n29), .ZN(
        u4_fract_out_pl1_2_) );
  INV_X4 u4_add_395_U57 ( .A(u4_fract_out_2_), .ZN(u4_add_395_n28) );
  INV_X4 u4_add_395_U56 ( .A(u4_fract_out_3_), .ZN(u4_add_395_n27) );
  XNOR2_X2 u4_add_395_U55 ( .A(u4_add_395_n26), .B(u4_add_395_n27), .ZN(
        u4_fract_out_pl1_3_) );
  INV_X4 u4_add_395_U54 ( .A(u4_fract_out_4_), .ZN(u4_add_395_n23) );
  XNOR2_X2 u4_add_395_U53 ( .A(u4_add_395_n21), .B(u4_add_395_n23), .ZN(
        u4_fract_out_pl1_4_) );
  INV_X4 u4_add_395_U52 ( .A(u4_fract_out_5_), .ZN(u4_add_395_n22) );
  XNOR2_X2 u4_add_395_U51 ( .A(u4_add_395_n24), .B(u4_add_395_n22), .ZN(
        u4_fract_out_pl1_5_) );
  NOR2_X4 u4_add_395_U50 ( .A1(u4_add_395_n22), .A2(u4_add_395_n23), .ZN(
        u4_add_395_n20) );
  NAND2_X2 u4_add_395_U49 ( .A1(u4_add_395_n20), .A2(u4_add_395_n21), .ZN(
        u4_add_395_n19) );
  INV_X4 u4_add_395_U48 ( .A(u4_add_395_n19), .ZN(u4_add_395_n17) );
  INV_X4 u4_add_395_U47 ( .A(u4_fract_out_6_), .ZN(u4_add_395_n18) );
  XNOR2_X2 u4_add_395_U46 ( .A(u4_add_395_n17), .B(u4_add_395_n18), .ZN(
        u4_fract_out_pl1_6_) );
  NAND2_X2 u4_add_395_U45 ( .A1(u4_add_395_n17), .A2(u4_fract_out_6_), .ZN(
        u4_add_395_n16) );
  XNOR2_X2 u4_add_395_U44 ( .A(u4_fract_out_7_), .B(u4_add_395_n16), .ZN(
        u4_fract_out_pl1_7_) );
  INV_X4 u4_add_395_U43 ( .A(u4_fract_out_8_), .ZN(u4_add_395_n14) );
  XNOR2_X2 u4_add_395_U42 ( .A(u4_add_395_n15), .B(u4_add_395_n14), .ZN(
        u4_fract_out_pl1_8_) );
  XNOR2_X2 u4_add_395_U41 ( .A(u4_add_395_n11), .B(u4_add_395_n12), .ZN(
        u4_fract_out_pl1_9_) );
  XNOR2_X1 u4_add_395_U40 ( .A(n3017), .B(u4_add_395_n38), .ZN(
        u4_fract_out_pl1_22_) );
  NAND3_X2 u4_add_395_U39 ( .A1(u4_add_395_n10), .A2(u4_fract_out_12_), .A3(
        u4_add_395_n60), .ZN(u4_add_395_n59) );
  INV_X2 u4_add_395_U38 ( .A(u4_fract_out_14_), .ZN(u4_add_395_n58) );
  NAND4_X1 u4_add_395_U37 ( .A1(u4_fract_out_19_), .A2(u4_fract_out_17_), .A3(
        u4_fract_out_18_), .A4(u4_fract_out_16_), .ZN(u4_add_395_n43) );
  CLKBUF_X3 u4_add_395_U36 ( .A(u4_fract_out_13_), .Z(u4_add_395_n10) );
  NAND2_X1 u4_add_395_U35 ( .A1(u4_add_395_n3), .A2(u4_fract_out_10_), .ZN(
        u4_add_395_n64) );
  NAND2_X1 u4_add_395_U34 ( .A1(u4_fract_out_15_), .A2(u4_fract_out_14_), .ZN(
        u4_add_395_n55) );
  XNOR2_X1 u4_add_395_U33 ( .A(u4_fract_out_15_), .B(u4_add_395_n56), .ZN(
        u4_fract_out_pl1_15_) );
  NAND2_X1 u4_add_395_U32 ( .A1(u4_add_395_n49), .A2(u4_fract_out_16_), .ZN(
        u4_add_395_n52) );
  XNOR2_X1 u4_add_395_U31 ( .A(u4_fract_out_16_), .B(u4_add_395_n42), .ZN(
        u4_fract_out_pl1_16_) );
  INV_X1 u4_add_395_U30 ( .A(u4_fract_out_16_), .ZN(u4_add_395_n50) );
  XNOR2_X1 u4_add_395_U29 ( .A(u4_fract_out_19_), .B(u4_add_395_n44), .ZN(
        u4_fract_out_pl1_19_) );
  INV_X1 u4_add_395_U28 ( .A(u4_fract_out_10_), .ZN(u4_add_395_n65) );
  NAND3_X2 u4_add_395_U27 ( .A1(u4_fract_out_15_), .A2(u4_fract_out_17_), .A3(
        u4_fract_out_16_), .ZN(u4_add_395_n35) );
  OR2_X4 u4_add_395_U26 ( .A1(u4_add_395_n34), .A2(u4_add_395_n35), .ZN(
        u4_add_395_n8) );
  OR2_X4 u4_add_395_U25 ( .A1(u4_add_395_n36), .A2(u4_add_395_n37), .ZN(
        u4_add_395_n7) );
  XNOR2_X1 u4_add_395_U24 ( .A(u4_fract_out_21_), .B(u4_add_395_n40), .ZN(
        u4_fract_out_pl1_21_) );
  NOR2_X2 u4_add_395_U23 ( .A1(u4_add_395_n54), .A2(u4_add_395_n55), .ZN(
        u4_add_395_n53) );
  NOR2_X2 u4_add_395_U22 ( .A1(u4_add_395_n50), .A2(u4_add_395_n51), .ZN(
        u4_add_395_n48) );
  NOR2_X4 u4_add_395_U21 ( .A1(u4_add_395_n30), .A2(u4_add_395_n31), .ZN(
        u4_add_395_n5) );
  XOR2_X1 u4_add_395_U20 ( .A(u4_fract_out_1_), .B(u4_fract_out_0_), .Z(
        u4_fract_out_pl1_1_) );
  NOR2_X1 u4_add_395_U19 ( .A1(u4_add_395_n13), .A2(u4_add_395_n14), .ZN(
        u4_add_395_n11) );
  NOR2_X1 u4_add_395_U18 ( .A1(u4_add_395_n25), .A2(u4_add_395_n23), .ZN(
        u4_add_395_n24) );
  NOR2_X1 u4_add_395_U17 ( .A1(u4_add_395_n28), .A2(u4_add_395_n29), .ZN(
        u4_add_395_n26) );
  NOR2_X2 u4_add_395_U16 ( .A1(u4_add_395_n67), .A2(u4_add_395_n68), .ZN(
        u4_add_395_n66) );
  INV_X4 u4_add_395_U15 ( .A(u4_add_395_n5), .ZN(u4_add_395_n9) );
  INV_X1 u4_add_395_U14 ( .A(u4_fract_out_9_), .ZN(u4_add_395_n12) );
  NAND2_X1 u4_add_395_U13 ( .A1(u4_add_395_n39), .A2(u4_fract_out_20_), .ZN(
        u4_add_395_n40) );
  NAND3_X1 u4_add_395_U12 ( .A1(u4_fract_out_21_), .A2(u4_fract_out_20_), .A3(
        u4_add_395_n39), .ZN(u4_add_395_n38) );
  INV_X1 u4_add_395_U11 ( .A(u4_fract_out_20_), .ZN(u4_add_395_n41) );
  XNOR2_X1 u4_add_395_U10 ( .A(u4_add_395_n39), .B(u4_add_395_n41), .ZN(
        u4_fract_out_pl1_20_) );
  OR2_X4 u4_add_395_U9 ( .A1(u4_add_395_n32), .A2(u4_add_395_n33), .ZN(
        u4_add_395_n2) );
  NAND3_X2 u4_add_395_U8 ( .A1(u4_fract_out_18_), .A2(u4_fract_out_19_), .A3(
        u4_fract_out_20_), .ZN(u4_add_395_n36) );
  NAND3_X2 u4_add_395_U7 ( .A1(u4_fract_out_2_), .A2(u4_fract_out_0_), .A3(
        u4_fract_out_1_), .ZN(u4_add_395_n30) );
  NOR4_X4 u4_add_395_U6 ( .A1(u4_add_395_n7), .A2(u4_add_395_n8), .A3(
        u4_add_395_n2), .A4(u4_add_395_n9), .ZN(u4_fract_out_pl1_23_) );
  AND3_X2 u4_add_395_U5 ( .A1(u4_fract_out_8_), .A2(u4_fract_out_9_), .A3(
        u4_add_395_n15), .ZN(u4_add_395_n3) );
  AND4_X4 u4_add_395_U4 ( .A1(u4_fract_out_11_), .A2(u4_fract_out_10_), .A3(
        u4_fract_out_9_), .A4(u4_fract_out_8_), .ZN(u4_add_395_n1) );
  NAND3_X4 u4_add_395_U3 ( .A1(u4_fract_out_9_), .A2(u4_fract_out_11_), .A3(
        u4_fract_out_10_), .ZN(u4_add_395_n33) );
  NAND2_X2 u4_add_395_U2 ( .A1(n3017), .A2(u4_fract_out_21_), .ZN(
        u4_add_395_n37) );
  NAND2_X2 u4_sub_495_U80 ( .A1(u4_exp_in_pl1_0_), .A2(u4_sub_495_n35), .ZN(
        u4_sub_495_n29) );
  INV_X4 u4_sub_495_U79 ( .A(u4_exp_in_pl1_0_), .ZN(u4_sub_495_n34) );
  NAND2_X2 u4_sub_495_U78 ( .A1(u4_ldz_all_0_), .A2(u4_sub_495_n34), .ZN(
        u4_sub_495_n30) );
  NAND2_X2 u4_sub_495_U77 ( .A1(u4_sub_495_n29), .A2(u4_sub_495_n30), .ZN(
        u4_div_exp2_0_) );
  NOR2_X4 u4_sub_495_U76 ( .A1(u4_sub_495_n22), .A2(u4_sub_495_n32), .ZN(
        u4_sub_495_n31) );
  INV_X4 u4_sub_495_U75 ( .A(u4_sub_495_n31), .ZN(u4_sub_495_n27) );
  INV_X4 u4_sub_495_U74 ( .A(u4_sub_495_n30), .ZN(u4_sub_495_n28) );
  XNOR2_X2 u4_sub_495_U73 ( .A(u4_sub_495_n27), .B(u4_sub_495_n24), .ZN(
        u4_div_exp2_1_) );
  INV_X4 u4_sub_495_U72 ( .A(u4_exp_in_pl1_1_), .ZN(u4_sub_495_n26) );
  XNOR2_X2 u4_sub_495_U71 ( .A(u4_sub_495_net32054), .B(u4_sub_495_net32055), 
        .ZN(u4_div_exp2_2_) );
  XNOR2_X2 u4_sub_495_U70 ( .A(u4_sub_495_net32044), .B(u4_sub_495_net32045), 
        .ZN(u4_div_exp2_3_) );
  XNOR2_X2 u4_sub_495_U69 ( .A(u4_sub_495_net32028), .B(u4_sub_495_net94054), 
        .ZN(u4_div_exp2_5_) );
  NAND2_X2 u4_sub_495_U68 ( .A1(u4_sub_495_n28), .A2(u4_sub_495_n29), .ZN(
        u4_sub_495_n24) );
  INV_X1 u4_sub_495_U67 ( .A(u4_sub_495_net95073), .ZN(u4_sub_495_net32045) );
  NAND2_X4 u4_sub_495_U66 ( .A1(u4_exp_in_pl1_1_), .A2(u4_sub_495_n33), .ZN(
        u4_sub_495_net32050) );
  XNOR2_X2 u4_sub_495_U65 ( .A(u4_sub_495_net91261), .B(u4_sub_495_n23), .ZN(
        u4_div_exp2_4_) );
  INV_X2 u4_sub_495_U64 ( .A(u4_ldz_all_0_), .ZN(u4_sub_495_n35) );
  INV_X4 u4_sub_495_U63 ( .A(u4_ldz_all_1_), .ZN(u4_sub_495_n33) );
  NOR2_X2 u4_sub_495_U62 ( .A1(u4_exp_in_pl1_1_), .A2(u4_sub_495_n33), .ZN(
        u4_sub_495_n32) );
  AND2_X2 u4_sub_495_U61 ( .A1(u4_exp_in_pl1_1_), .A2(u4_sub_495_n33), .ZN(
        u4_sub_495_n22) );
  NAND2_X4 u4_sub_495_U60 ( .A1(u4_sub_495_n24), .A2(u4_sub_495_n25), .ZN(
        u4_sub_495_net32051) );
  INV_X4 u4_sub_495_U59 ( .A(u4_exp_in_pl1_5_), .ZN(u4_sub_495_n20) );
  NAND2_X4 u4_sub_495_U58 ( .A1(u4_ldz_all_5_), .A2(u4_sub_495_n20), .ZN(
        u4_sub_495_net32027) );
  INV_X4 u4_sub_495_U57 ( .A(u4_ldz_all_5_), .ZN(u4_sub_495_n21) );
  NAND2_X4 u4_sub_495_U56 ( .A1(u4_sub_495_n21), .A2(u4_exp_in_pl1_5_), .ZN(
        u4_sub_495_net32025) );
  NAND2_X1 u4_sub_495_U55 ( .A1(u4_sub_495_net32051), .A2(u4_sub_495_net32050), 
        .ZN(u4_sub_495_net32055) );
  INV_X4 u4_sub_495_U54 ( .A(u4_exp_in_pl1_3_), .ZN(u4_sub_495_net32052) );
  NAND2_X2 u4_sub_495_U53 ( .A1(u4_ldz_all_3_), .A2(u4_sub_495_net32052), .ZN(
        u4_sub_495_net32043) );
  NAND2_X4 u4_sub_495_U52 ( .A1(u4_sub_495_net32050), .A2(u4_sub_495_net32051), 
        .ZN(u4_sub_495_net32047) );
  INV_X4 u4_sub_495_U51 ( .A(u4_ldz_all_3_), .ZN(u4_sub_495_n19) );
  NAND2_X4 u4_sub_495_U50 ( .A1(u4_exp_in_pl1_3_), .A2(u4_sub_495_n19), .ZN(
        u4_sub_495_net32042) );
  INV_X4 u4_sub_495_U49 ( .A(u4_exp_in_pl1_4_), .ZN(u4_sub_495_n17) );
  INV_X4 u4_sub_495_U48 ( .A(n2924), .ZN(u4_sub_495_n18) );
  NAND2_X4 u4_sub_495_U47 ( .A1(u4_sub_495_n18), .A2(u4_exp_in_pl1_4_), .ZN(
        u4_sub_495_net32031) );
  NAND2_X1 u4_sub_495_U46 ( .A1(u4_sub_495_net32042), .A2(u4_sub_495_net32043), 
        .ZN(u4_sub_495_net32044) );
  INV_X4 u4_sub_495_U45 ( .A(u4_sub_495_net32036), .ZN(u4_sub_495_net32029) );
  INV_X2 u4_sub_495_U44 ( .A(u4_sub_495_net32031), .ZN(u4_sub_495_net32035) );
  INV_X4 u4_sub_495_U43 ( .A(u4_exp_in_pl1_6_), .ZN(u4_sub_495_n12) );
  INV_X4 u4_sub_495_U42 ( .A(u4_sub_495_net32015), .ZN(u4_sub_495_net32019) );
  NAND2_X2 u4_sub_495_U41 ( .A1(u4_ldz_all_6_), .A2(u4_sub_495_n12), .ZN(
        u4_sub_495_net32015) );
  INV_X4 u4_sub_495_U40 ( .A(u4_sub_495_net32043), .ZN(u4_sub_495_net32040) );
  AOI21_X1 u4_sub_495_U39 ( .B1(u4_sub_495_net32047), .B2(u4_sub_495_net32046), 
        .A(u4_sub_495_net32048), .ZN(u4_sub_495_net95073) );
  AOI21_X4 u4_sub_495_U38 ( .B1(u4_sub_495_net32047), .B2(u4_sub_495_net32046), 
        .A(u4_sub_495_net32048), .ZN(u4_sub_495_n16) );
  OAI21_X4 u4_sub_495_U37 ( .B1(u4_sub_495_net32040), .B2(u4_sub_495_n16), .A(
        u4_sub_495_net32042), .ZN(u4_sub_495_net32039) );
  OAI21_X2 u4_sub_495_U36 ( .B1(u4_sub_495_net32030), .B2(u4_sub_495_net32029), 
        .A(u4_sub_495_net32031), .ZN(u4_sub_495_net94054) );
  INV_X8 u4_sub_495_U35 ( .A(u4_sub_495_net32039), .ZN(u4_sub_495_net32030) );
  OAI21_X4 u4_sub_495_U34 ( .B1(u4_sub_495_net32030), .B2(u4_sub_495_net32029), 
        .A(u4_sub_495_net32031), .ZN(u4_sub_495_n15) );
  INV_X4 u4_sub_495_U33 ( .A(u4_sub_495_net32027), .ZN(u4_sub_495_n14) );
  OAI21_X4 u4_sub_495_U32 ( .B1(u4_sub_495_net32024), .B2(u4_sub_495_n14), .A(
        u4_sub_495_net32025), .ZN(u4_sub_495_n11) );
  INV_X4 u4_sub_495_U31 ( .A(u4_ldz_all_6_), .ZN(u4_sub_495_n13) );
  NAND2_X2 u4_sub_495_U30 ( .A1(u4_exp_in_pl1_6_), .A2(u4_sub_495_n13), .ZN(
        u4_sub_495_net32021) );
  NOR2_X4 u4_sub_495_U29 ( .A1(u4_sub_495_net32016), .A2(u4_sub_495_net32019), 
        .ZN(u4_sub_495_net32018) );
  INV_X4 u4_sub_495_U28 ( .A(u4_sub_495_net32021), .ZN(u4_sub_495_net32016) );
  AOI21_X4 u4_sub_495_U27 ( .B1(u4_sub_495_n11), .B2(u4_sub_495_net32015), .A(
        u4_sub_495_net32016), .ZN(u4_sub_495_net32012) );
  NAND2_X2 u4_sub_495_U26 ( .A1(u4_sub_495_n9), .A2(u4_ldz_all_2_), .ZN(
        u4_sub_495_net32046) );
  INV_X4 u4_sub_495_U25 ( .A(u4_exp_in_pl1_2_), .ZN(u4_sub_495_n9) );
  NAND2_X1 u4_sub_495_U24 ( .A1(u4_sub_495_net32049), .A2(u4_sub_495_net32046), 
        .ZN(u4_sub_495_net32054) );
  INV_X8 u4_sub_495_U23 ( .A(u4_sub_495_net32049), .ZN(u4_sub_495_net32048) );
  NAND2_X4 u4_sub_495_U22 ( .A1(u4_sub_495_n10), .A2(u4_exp_in_pl1_2_), .ZN(
        u4_sub_495_net32049) );
  NOR2_X2 u4_sub_495_U21 ( .A1(u4_sub_495_net32035), .A2(u4_sub_495_net32029), 
        .ZN(u4_sub_495_n23) );
  INV_X4 u4_sub_495_U20 ( .A(u4_sub_495_n11), .ZN(u4_sub_495_net32017) );
  INV_X1 u4_sub_495_U19 ( .A(u4_exp_in_pl1_7_), .ZN(u4_sub_495_net32013) );
  INV_X4 u4_sub_495_U18 ( .A(u4_sub_495_net32013), .ZN(u4_sub_495_n6) );
  INV_X4 u4_sub_495_U17 ( .A(u4_sub_495_net32012), .ZN(u4_sub_495_n5) );
  NAND2_X4 u4_sub_495_U16 ( .A1(u4_sub_495_n7), .A2(u4_sub_495_n8), .ZN(
        u4_div_exp2_7_) );
  NAND2_X4 u4_sub_495_U15 ( .A1(u4_sub_495_n5), .A2(u4_sub_495_n6), .ZN(
        u4_sub_495_n8) );
  NAND2_X2 u4_sub_495_U14 ( .A1(u4_sub_495_net32013), .A2(u4_sub_495_net32012), 
        .ZN(u4_sub_495_n7) );
  NAND2_X4 u4_sub_495_U13 ( .A1(u4_ldz_all_1_), .A2(u4_sub_495_n26), .ZN(
        u4_sub_495_n25) );
  INV_X8 u4_sub_495_U12 ( .A(u4_ldz_all_2_), .ZN(u4_sub_495_n10) );
  BUF_X4 u4_sub_495_U11 ( .A(u4_sub_495_net32030), .Z(u4_sub_495_net91261) );
  NAND2_X4 u4_sub_495_U10 ( .A1(u4_sub_495_net32025), .A2(u4_sub_495_net32027), 
        .ZN(u4_sub_495_net32028) );
  INV_X4 u4_sub_495_U9 ( .A(u4_sub_495_net32018), .ZN(u4_sub_495_n2) );
  INV_X4 u4_sub_495_U8 ( .A(u4_sub_495_net32017), .ZN(u4_sub_495_n1) );
  NAND2_X4 u4_sub_495_U7 ( .A1(u4_sub_495_n3), .A2(u4_sub_495_n4), .ZN(
        u4_div_exp2_6_) );
  NAND2_X4 u4_sub_495_U6 ( .A1(u4_sub_495_n1), .A2(u4_sub_495_n2), .ZN(
        u4_sub_495_n4) );
  NAND2_X2 u4_sub_495_U5 ( .A1(u4_sub_495_net32017), .A2(u4_sub_495_net32018), 
        .ZN(u4_sub_495_n3) );
  NAND2_X2 u4_sub_495_U4 ( .A1(n2924), .A2(u4_sub_495_n17), .ZN(
        u4_sub_495_net32036) );
  INV_X8 u4_sub_495_U3 ( .A(u4_sub_495_n15), .ZN(u4_sub_495_net32024) );
  INV_X4 u4_add_463_U22 ( .A(n4756), .ZN(u4_exp_out_pl1_0_) );
  XNOR2_X2 u4_add_463_U21 ( .A(u4_exp_out_2_), .B(u4_add_463_n13), .ZN(
        u4_exp_out_pl1_2_) );
  INV_X4 u4_add_463_U20 ( .A(u4_exp_out_2_), .ZN(u4_add_463_n14) );
  XNOR2_X2 u4_add_463_U19 ( .A(u4_add_463_n11), .B(u4_add_463_n12), .ZN(
        u4_exp_out_pl1_3_) );
  INV_X4 u4_add_463_U18 ( .A(u4_add_463_n5), .ZN(u4_add_463_n9) );
  XNOR2_X2 u4_add_463_U17 ( .A(u4_add_463_n1), .B(u4_add_463_n10), .ZN(
        u4_exp_out_pl1_4_) );
  NAND2_X2 u4_add_463_U16 ( .A1(n4756), .A2(u4_add_463_n4), .ZN(u4_add_463_n3)
         );
  XNOR2_X1 u4_add_463_U15 ( .A(net95138), .B(u4_add_463_n3), .ZN(
        u4_exp_out_pl1_7_) );
  NAND3_X1 u4_add_463_U14 ( .A1(n2476), .A2(net94896), .A3(u4_exp_out_4_), 
        .ZN(u4_add_463_n6) );
  XNOR2_X1 u4_add_463_U13 ( .A(n2476), .B(u4_add_463_n7), .ZN(
        u4_exp_out_pl1_6_) );
  NAND3_X1 u4_add_463_U12 ( .A1(u4_add_463_n9), .A2(u4_exp_out_4_), .A3(n4756), 
        .ZN(u4_add_463_n8) );
  NAND3_X1 u4_add_463_U11 ( .A1(net94896), .A2(u4_exp_out_4_), .A3(
        u4_add_463_n1), .ZN(u4_add_463_n7) );
  NAND3_X1 u4_add_463_U10 ( .A1(u4_exp_out_2_), .A2(net94566), .A3(net94948), 
        .ZN(u4_add_463_n5) );
  INV_X1 u4_add_463_U9 ( .A(net94566), .ZN(u4_add_463_n12) );
  NAND2_X1 u4_add_463_U8 ( .A1(net94948), .A2(n4756), .ZN(u4_add_463_n13) );
  XNOR2_X1 u4_add_463_U7 ( .A(net94896), .B(u4_add_463_n8), .ZN(
        u4_exp_out_pl1_5_) );
  NOR2_X1 u4_add_463_U6 ( .A1(u4_add_463_n5), .A2(u4_add_463_n6), .ZN(
        u4_add_463_n4) );
  INV_X1 u4_add_463_U5 ( .A(u4_exp_out_4_), .ZN(u4_add_463_n10) );
  XOR2_X1 u4_add_463_U4 ( .A(net94948), .B(n4756), .Z(u4_exp_out_pl1_1_) );
  NOR2_X2 u4_add_463_U3 ( .A1(u4_add_463_n13), .A2(u4_add_463_n14), .ZN(
        u4_add_463_n11) );
  AND2_X2 u4_add_463_U2 ( .A1(u4_add_463_n9), .A2(n4756), .ZN(u4_add_463_n1)
         );
  NOR2_X4 u4_add_493_U82 ( .A1(u4_add_493_n1), .A2(u4_add_493_n72), .ZN(
        u4_div_exp1_0_) );
  INV_X4 u4_add_493_U81 ( .A(u4_exp_in_mi1_1_), .ZN(u4_add_493_n71) );
  NAND2_X2 u4_add_493_U80 ( .A1(u4_add_493_n70), .A2(u4_add_493_n71), .ZN(
        u4_add_493_n67) );
  NAND2_X2 u4_add_493_U79 ( .A1(u4_add_493_n67), .A2(u4_add_493_n55), .ZN(
        u4_add_493_n69) );
  XNOR2_X2 u4_add_493_U78 ( .A(u4_add_493_n69), .B(u4_add_493_n1), .ZN(
        u4_div_exp1_1_) );
  INV_X4 u4_add_493_U77 ( .A(u4_add_493_n53), .ZN(u4_add_493_n68) );
  NAND2_X2 u4_add_493_U76 ( .A1(u4_add_493_n59), .A2(u4_add_493_n68), .ZN(
        u4_add_493_n63) );
  INV_X4 u4_add_493_U75 ( .A(u4_add_493_n67), .ZN(u4_add_493_n65) );
  NOR2_X4 u4_add_493_U74 ( .A1(u4_add_493_n65), .A2(u4_add_493_n66), .ZN(
        u4_add_493_n45) );
  INV_X4 u4_add_493_U73 ( .A(u4_add_493_n45), .ZN(u4_add_493_n64) );
  XNOR2_X2 u4_add_493_U72 ( .A(u4_add_493_n63), .B(u4_add_493_n60), .ZN(
        u4_div_exp1_2_) );
  INV_X4 u4_add_493_U71 ( .A(n2656), .ZN(u4_add_493_n62) );
  NAND2_X2 u4_add_493_U70 ( .A1(u4_add_493_n61), .A2(u4_add_493_n62), .ZN(
        u4_add_493_n54) );
  NAND2_X2 u4_add_493_U69 ( .A1(u4_add_493_n54), .A2(u4_add_493_n40), .ZN(
        u4_add_493_n56) );
  INV_X4 u4_add_493_U68 ( .A(u4_add_493_n60), .ZN(u4_add_493_n58) );
  OAI21_X4 u4_add_493_U67 ( .B1(u4_add_493_n53), .B2(u4_add_493_n58), .A(
        u4_add_493_n59), .ZN(u4_add_493_n57) );
  XNOR2_X2 u4_add_493_U66 ( .A(u4_add_493_n56), .B(u4_add_493_n57), .ZN(
        u4_div_exp1_3_) );
  INV_X4 u4_add_493_U65 ( .A(u4_add_493_n24), .ZN(u4_add_493_n38) );
  INV_X4 u4_add_493_U64 ( .A(u4_add_493_n55), .ZN(u4_add_493_n44) );
  INV_X4 u4_add_493_U63 ( .A(u4_add_493_n54), .ZN(u4_add_493_n51) );
  INV_X4 u4_add_493_U62 ( .A(u4_add_493_n43), .ZN(u4_add_493_n47) );
  INV_X4 u4_add_493_U61 ( .A(u4_exp_in_mi1_2_), .ZN(u4_add_493_n52) );
  NOR3_X4 u4_add_493_U60 ( .A1(u4_add_493_n50), .A2(u4_add_493_n51), .A3(
        u4_add_493_n52), .ZN(u4_add_493_n41) );
  NOR2_X4 u4_add_493_U59 ( .A1(u4_add_493_n41), .A2(u4_add_493_n49), .ZN(
        u4_add_493_n48) );
  OAI21_X4 u4_add_493_U58 ( .B1(u4_add_493_n46), .B2(u4_add_493_n47), .A(
        u4_add_493_n48), .ZN(u4_add_493_n25) );
  XNOR2_X2 u4_add_493_U57 ( .A(u4_add_493_n2), .B(u4_add_493_n25), .ZN(
        u4_div_exp1_4_) );
  NAND2_X2 u4_add_493_U56 ( .A1(u4_add_493_n42), .A2(u4_add_493_n43), .ZN(
        u4_add_493_n35) );
  NAND2_X2 u4_add_493_U55 ( .A1(u4_add_493_n41), .A2(u4_add_493_n42), .ZN(
        u4_add_493_n36) );
  OAI211_X2 u4_add_493_U54 ( .C1(u4_add_493_n34), .C2(u4_add_493_n35), .A(
        u4_add_493_n36), .B(u4_add_493_n37), .ZN(u4_add_493_n30) );
  INV_X4 u4_add_493_U53 ( .A(u4_fi_ldz_2a_5_), .ZN(u4_add_493_n32) );
  INV_X4 u4_add_493_U52 ( .A(u4_exp_in_mi1_5_), .ZN(u4_add_493_n33) );
  NAND2_X2 u4_add_493_U51 ( .A1(u4_add_493_n32), .A2(u4_add_493_n33), .ZN(
        u4_add_493_n28) );
  NAND2_X2 u4_add_493_U50 ( .A1(u4_fi_ldz_2a_5_), .A2(u4_exp_in_mi1_5_), .ZN(
        u4_add_493_n22) );
  NAND2_X2 u4_add_493_U49 ( .A1(u4_add_493_n28), .A2(u4_add_493_n22), .ZN(
        u4_add_493_n31) );
  XNOR2_X2 u4_add_493_U48 ( .A(u4_add_493_n30), .B(u4_add_493_n31), .ZN(
        u4_div_exp1_5_) );
  INV_X4 u4_add_493_U47 ( .A(u4_fi_ldz_2a_6_), .ZN(u4_add_493_n15) );
  INV_X4 u4_add_493_U46 ( .A(u4_exp_in_mi1_6_), .ZN(u4_add_493_n29) );
  NAND2_X2 u4_add_493_U45 ( .A1(u4_add_493_n15), .A2(u4_add_493_n29), .ZN(
        u4_add_493_n14) );
  NAND2_X2 u4_add_493_U44 ( .A1(u4_fi_ldz_2a_6_), .A2(u4_exp_in_mi1_6_), .ZN(
        u4_add_493_n12) );
  NAND2_X2 u4_add_493_U43 ( .A1(u4_add_493_n14), .A2(u4_add_493_n12), .ZN(
        u4_add_493_n17) );
  INV_X4 u4_add_493_U42 ( .A(u4_add_493_n28), .ZN(u4_add_493_n27) );
  INV_X4 u4_add_493_U41 ( .A(u4_add_493_n25), .ZN(u4_add_493_n23) );
  NAND2_X2 u4_add_493_U40 ( .A1(u4_add_493_n23), .A2(u4_add_493_n24), .ZN(
        u4_add_493_n20) );
  INV_X4 u4_add_493_U39 ( .A(u4_add_493_n22), .ZN(u4_add_493_n21) );
  AOI21_X4 u4_add_493_U38 ( .B1(u4_add_493_n19), .B2(u4_add_493_n20), .A(
        u4_add_493_n21), .ZN(u4_add_493_n18) );
  INV_X4 u4_add_493_U37 ( .A(u4_add_493_n18), .ZN(u4_add_493_n13) );
  XNOR2_X2 u4_add_493_U36 ( .A(u4_add_493_n17), .B(u4_add_493_n13), .ZN(
        u4_div_exp1_6_) );
  NAND2_X2 u4_add_493_U35 ( .A1(u4_exp_in_mi1_7_), .A2(u4_fi_ldz_2a_6_), .ZN(
        u4_add_493_n7) );
  INV_X4 u4_add_493_U34 ( .A(u4_exp_in_mi1_7_), .ZN(u4_add_493_n16) );
  NAND2_X2 u4_add_493_U33 ( .A1(u4_add_493_n15), .A2(u4_add_493_n16), .ZN(
        u4_add_493_n9) );
  NAND2_X2 u4_add_493_U32 ( .A1(u4_add_493_n7), .A2(u4_add_493_n9), .ZN(
        u4_add_493_n10) );
  INV_X4 u4_add_493_U31 ( .A(u4_add_493_n14), .ZN(u4_add_493_n11) );
  OAI21_X4 u4_add_493_U30 ( .B1(u4_add_493_n11), .B2(u4_add_493_n18), .A(
        u4_add_493_n12), .ZN(u4_add_493_n8) );
  XNOR2_X2 u4_add_493_U29 ( .A(u4_add_493_n10), .B(u4_add_493_n8), .ZN(
        u4_div_exp1_7_) );
  INV_X4 u4_add_493_U28 ( .A(u4_add_493_n9), .ZN(u4_add_493_n5) );
  INV_X4 u4_add_493_U27 ( .A(u4_add_493_n8), .ZN(u4_add_493_n6) );
  OAI21_X4 u4_add_493_U26 ( .B1(u4_add_493_n5), .B2(u4_add_493_n6), .A(
        u4_add_493_n7), .ZN(u4_add_493_n4) );
  XNOR2_X2 u4_add_493_U25 ( .A(u4_add_493_n3), .B(u4_add_493_n4), .ZN(
        u4_div_exp1_8_) );
  NAND2_X1 u4_add_493_U24 ( .A1(net22501), .A2(n4757), .ZN(u4_add_493_n66) );
  NOR2_X1 u4_add_493_U23 ( .A1(net22501), .A2(n4757), .ZN(u4_add_493_n72) );
  INV_X4 u4_add_493_U22 ( .A(net86044), .ZN(u4_add_493_n3) );
  NOR2_X4 u4_add_493_U21 ( .A1(u4_add_493_n45), .A2(u4_add_493_n44), .ZN(
        u4_add_493_n46) );
  NAND2_X2 u4_add_493_U20 ( .A1(u4_add_493_n64), .A2(u4_add_493_n55), .ZN(
        u4_add_493_n60) );
  NAND2_X1 u4_add_493_U19 ( .A1(net33106), .A2(u4_exp_in_mi1_1_), .ZN(
        u4_add_493_n55) );
  NAND2_X1 u4_add_493_U18 ( .A1(u4_fi_ldz_2a_3_), .A2(n2656), .ZN(
        u4_add_493_n40) );
  INV_X1 u4_add_493_U17 ( .A(net33106), .ZN(u4_add_493_n70) );
  INV_X1 u4_add_493_U16 ( .A(u4_fi_ldz_2a_3_), .ZN(u4_add_493_n61) );
  NOR2_X2 u4_add_493_U15 ( .A1(u4_add_493_n26), .A2(u4_add_493_n40), .ZN(
        u4_add_493_n39) );
  INV_X2 u4_add_493_U14 ( .A(u4_add_493_n26), .ZN(u4_add_493_n42) );
  NOR2_X2 u4_add_493_U13 ( .A1(u4_exp_in_mi1_4_), .A2(u4_fi_ldz_2a_4_), .ZN(
        u4_add_493_n26) );
  NOR2_X2 u4_add_493_U12 ( .A1(u4_add_493_n44), .A2(u4_add_493_n45), .ZN(
        u4_add_493_n34) );
  INV_X2 u4_add_493_U11 ( .A(u4_add_493_n40), .ZN(u4_add_493_n49) );
  NAND2_X1 u4_add_493_U10 ( .A1(u4_fi_ldz_2a_4_), .A2(u4_exp_in_mi1_4_), .ZN(
        u4_add_493_n24) );
  OR2_X2 u4_add_493_U9 ( .A1(u4_add_493_n26), .A2(u4_add_493_n38), .ZN(
        u4_add_493_n2) );
  AND2_X2 u4_add_493_U8 ( .A1(n4757), .A2(net22501), .ZN(u4_add_493_n1) );
  NOR2_X2 u4_add_493_U7 ( .A1(u4_add_493_n26), .A2(u4_add_493_n27), .ZN(
        u4_add_493_n19) );
  NOR2_X2 u4_add_493_U6 ( .A1(u4_add_493_n38), .A2(u4_add_493_n39), .ZN(
        u4_add_493_n37) );
  NOR2_X2 u4_add_493_U5 ( .A1(u4_add_493_n51), .A2(u4_add_493_n53), .ZN(
        u4_add_493_n43) );
  NOR2_X1 u4_add_493_U4 ( .A1(u4_exp_in_mi1_2_), .A2(net23043), .ZN(
        u4_add_493_n53) );
  INV_X1 u4_add_493_U3 ( .A(net23043), .ZN(u4_add_493_n50) );
  NAND2_X1 u4_add_493_U2 ( .A1(net23043), .A2(u4_exp_in_mi1_2_), .ZN(
        u4_add_493_n59) );
  INV_X4 add_0_root_sub_0_root_u4_add_496_U75 ( .A(u4_ldz_dif_1_), .ZN(
        add_0_root_sub_0_root_u4_add_496_n65) );
  NAND2_X2 add_0_root_sub_0_root_u4_add_496_U74 ( .A1(
        add_0_root_sub_0_root_u4_add_496_n64), .A2(
        add_0_root_sub_0_root_u4_add_496_n65), .ZN(
        add_0_root_sub_0_root_u4_add_496_n59) );
  NAND2_X2 add_0_root_sub_0_root_u4_add_496_U73 ( .A1(
        add_0_root_sub_0_root_u4_add_496_n59), .A2(
        add_0_root_sub_0_root_u4_add_496_n46), .ZN(
        add_0_root_sub_0_root_u4_add_496_n61) );
  XNOR2_X2 add_0_root_sub_0_root_u4_add_496_U72 ( .A(
        add_0_root_sub_0_root_u4_add_496_n61), .B(
        add_0_root_sub_0_root_u4_add_496_n62), .ZN(u4_div_exp3[1]) );
  INV_X4 add_0_root_sub_0_root_u4_add_496_U71 ( .A(
        add_0_root_sub_0_root_u4_add_496_n44), .ZN(
        add_0_root_sub_0_root_u4_add_496_n60) );
  NAND2_X2 add_0_root_sub_0_root_u4_add_496_U70 ( .A1(
        add_0_root_sub_0_root_u4_add_496_n51), .A2(
        add_0_root_sub_0_root_u4_add_496_n60), .ZN(
        add_0_root_sub_0_root_u4_add_496_n55) );
  INV_X4 add_0_root_sub_0_root_u4_add_496_U69 ( .A(
        add_0_root_sub_0_root_u4_add_496_n59), .ZN(
        add_0_root_sub_0_root_u4_add_496_n57) );
  XNOR2_X2 add_0_root_sub_0_root_u4_add_496_U68 ( .A(
        add_0_root_sub_0_root_u4_add_496_n55), .B(
        add_0_root_sub_0_root_u4_add_496_n52), .ZN(u4_div_exp3[2]) );
  INV_X4 add_0_root_sub_0_root_u4_add_496_U67 ( .A(u4_ldz_dif_3_), .ZN(
        add_0_root_sub_0_root_u4_add_496_n54) );
  NAND2_X2 add_0_root_sub_0_root_u4_add_496_U66 ( .A1(
        add_0_root_sub_0_root_u4_add_496_n53), .A2(
        add_0_root_sub_0_root_u4_add_496_n54), .ZN(
        add_0_root_sub_0_root_u4_add_496_n45) );
  NAND2_X2 add_0_root_sub_0_root_u4_add_496_U65 ( .A1(
        add_0_root_sub_0_root_u4_add_496_n45), .A2(
        add_0_root_sub_0_root_u4_add_496_n30), .ZN(
        add_0_root_sub_0_root_u4_add_496_n48) );
  INV_X4 add_0_root_sub_0_root_u4_add_496_U64 ( .A(
        add_0_root_sub_0_root_u4_add_496_n52), .ZN(
        add_0_root_sub_0_root_u4_add_496_n50) );
  XNOR2_X2 add_0_root_sub_0_root_u4_add_496_U63 ( .A(
        add_0_root_sub_0_root_u4_add_496_n48), .B(
        add_0_root_sub_0_root_u4_add_496_n49), .ZN(u4_div_exp3[3]) );
  INV_X4 add_0_root_sub_0_root_u4_add_496_U62 ( .A(
        add_0_root_sub_0_root_u4_add_496_n14), .ZN(
        add_0_root_sub_0_root_u4_add_496_n28) );
  INV_X4 add_0_root_sub_0_root_u4_add_496_U61 ( .A(
        add_0_root_sub_0_root_u4_add_496_n47), .ZN(
        add_0_root_sub_0_root_u4_add_496_n36) );
  INV_X4 add_0_root_sub_0_root_u4_add_496_U60 ( .A(
        add_0_root_sub_0_root_u4_add_496_n46), .ZN(
        add_0_root_sub_0_root_u4_add_496_n33) );
  INV_X4 add_0_root_sub_0_root_u4_add_496_U59 ( .A(
        add_0_root_sub_0_root_u4_add_496_n45), .ZN(
        add_0_root_sub_0_root_u4_add_496_n42) );
  INV_X4 add_0_root_sub_0_root_u4_add_496_U58 ( .A(
        add_0_root_sub_0_root_u4_add_496_n31), .ZN(
        add_0_root_sub_0_root_u4_add_496_n38) );
  INV_X4 add_0_root_sub_0_root_u4_add_496_U57 ( .A(u4_ldz_dif_2_), .ZN(
        add_0_root_sub_0_root_u4_add_496_n43) );
  NOR3_X4 add_0_root_sub_0_root_u4_add_496_U56 ( .A1(
        add_0_root_sub_0_root_u4_add_496_n41), .A2(
        add_0_root_sub_0_root_u4_add_496_n42), .A3(
        add_0_root_sub_0_root_u4_add_496_n43), .ZN(
        add_0_root_sub_0_root_u4_add_496_n26) );
  NOR2_X4 add_0_root_sub_0_root_u4_add_496_U55 ( .A1(
        add_0_root_sub_0_root_u4_add_496_n26), .A2(
        add_0_root_sub_0_root_u4_add_496_n40), .ZN(
        add_0_root_sub_0_root_u4_add_496_n39) );
  OAI21_X4 add_0_root_sub_0_root_u4_add_496_U54 ( .B1(
        add_0_root_sub_0_root_u4_add_496_n37), .B2(
        add_0_root_sub_0_root_u4_add_496_n38), .A(
        add_0_root_sub_0_root_u4_add_496_n39), .ZN(
        add_0_root_sub_0_root_u4_add_496_n15) );
  XNOR2_X2 add_0_root_sub_0_root_u4_add_496_U53 ( .A(
        add_0_root_sub_0_root_u4_add_496_n36), .B(
        add_0_root_sub_0_root_u4_add_496_n15), .ZN(u4_div_exp3[4]) );
  INV_X4 add_0_root_sub_0_root_u4_add_496_U52 ( .A(u4_fi_ldz_2a_5_), .ZN(
        add_0_root_sub_0_root_u4_add_496_n34) );
  INV_X4 add_0_root_sub_0_root_u4_add_496_U51 ( .A(u4_ldz_dif_5_), .ZN(
        add_0_root_sub_0_root_u4_add_496_n35) );
  NAND2_X2 add_0_root_sub_0_root_u4_add_496_U50 ( .A1(
        add_0_root_sub_0_root_u4_add_496_n34), .A2(
        add_0_root_sub_0_root_u4_add_496_n35), .ZN(
        add_0_root_sub_0_root_u4_add_496_n18) );
  NAND2_X2 add_0_root_sub_0_root_u4_add_496_U49 ( .A1(u4_fi_ldz_2a_5_), .A2(
        u4_ldz_dif_5_), .ZN(add_0_root_sub_0_root_u4_add_496_n12) );
  NAND2_X2 add_0_root_sub_0_root_u4_add_496_U48 ( .A1(
        add_0_root_sub_0_root_u4_add_496_n18), .A2(
        add_0_root_sub_0_root_u4_add_496_n12), .ZN(
        add_0_root_sub_0_root_u4_add_496_n21) );
  INV_X4 add_0_root_sub_0_root_u4_add_496_U47 ( .A(
        add_0_root_sub_0_root_u4_add_496_n16), .ZN(
        add_0_root_sub_0_root_u4_add_496_n27) );
  NAND2_X2 add_0_root_sub_0_root_u4_add_496_U46 ( .A1(
        add_0_root_sub_0_root_u4_add_496_n26), .A2(
        add_0_root_sub_0_root_u4_add_496_n27), .ZN(
        add_0_root_sub_0_root_u4_add_496_n25) );
  OAI211_X2 add_0_root_sub_0_root_u4_add_496_U45 ( .C1(
        add_0_root_sub_0_root_u4_add_496_n37), .C2(
        add_0_root_sub_0_root_u4_add_496_n23), .A(
        add_0_root_sub_0_root_u4_add_496_n24), .B(
        add_0_root_sub_0_root_u4_add_496_n25), .ZN(
        add_0_root_sub_0_root_u4_add_496_n22) );
  XNOR2_X2 add_0_root_sub_0_root_u4_add_496_U44 ( .A(
        add_0_root_sub_0_root_u4_add_496_n21), .B(
        add_0_root_sub_0_root_u4_add_496_n22), .ZN(u4_div_exp3[5]) );
  INV_X4 add_0_root_sub_0_root_u4_add_496_U43 ( .A(u4_fi_ldz_2a_6_), .ZN(
        add_0_root_sub_0_root_u4_add_496_n19) );
  INV_X4 add_0_root_sub_0_root_u4_add_496_U42 ( .A(u4_ldz_dif_6_), .ZN(
        add_0_root_sub_0_root_u4_add_496_n20) );
  NAND2_X2 add_0_root_sub_0_root_u4_add_496_U41 ( .A1(
        add_0_root_sub_0_root_u4_add_496_n19), .A2(
        add_0_root_sub_0_root_u4_add_496_n20), .ZN(
        add_0_root_sub_0_root_u4_add_496_n6) );
  NAND2_X2 add_0_root_sub_0_root_u4_add_496_U40 ( .A1(u4_fi_ldz_2a_6_), .A2(
        u4_ldz_dif_6_), .ZN(add_0_root_sub_0_root_u4_add_496_n5) );
  NAND2_X2 add_0_root_sub_0_root_u4_add_496_U39 ( .A1(
        add_0_root_sub_0_root_u4_add_496_n6), .A2(
        add_0_root_sub_0_root_u4_add_496_n5), .ZN(
        add_0_root_sub_0_root_u4_add_496_n7) );
  INV_X4 add_0_root_sub_0_root_u4_add_496_U38 ( .A(
        add_0_root_sub_0_root_u4_add_496_n18), .ZN(
        add_0_root_sub_0_root_u4_add_496_n17) );
  INV_X4 add_0_root_sub_0_root_u4_add_496_U37 ( .A(
        add_0_root_sub_0_root_u4_add_496_n15), .ZN(
        add_0_root_sub_0_root_u4_add_496_n13) );
  NAND2_X2 add_0_root_sub_0_root_u4_add_496_U36 ( .A1(
        add_0_root_sub_0_root_u4_add_496_n13), .A2(
        add_0_root_sub_0_root_u4_add_496_n14), .ZN(
        add_0_root_sub_0_root_u4_add_496_n10) );
  INV_X4 add_0_root_sub_0_root_u4_add_496_U35 ( .A(
        add_0_root_sub_0_root_u4_add_496_n12), .ZN(
        add_0_root_sub_0_root_u4_add_496_n11) );
  AOI21_X4 add_0_root_sub_0_root_u4_add_496_U34 ( .B1(
        add_0_root_sub_0_root_u4_add_496_n9), .B2(
        add_0_root_sub_0_root_u4_add_496_n10), .A(
        add_0_root_sub_0_root_u4_add_496_n11), .ZN(
        add_0_root_sub_0_root_u4_add_496_n4) );
  INV_X4 add_0_root_sub_0_root_u4_add_496_U33 ( .A(
        add_0_root_sub_0_root_u4_add_496_n4), .ZN(
        add_0_root_sub_0_root_u4_add_496_n8) );
  XNOR2_X2 add_0_root_sub_0_root_u4_add_496_U32 ( .A(
        add_0_root_sub_0_root_u4_add_496_n7), .B(
        add_0_root_sub_0_root_u4_add_496_n8), .ZN(u4_div_exp3[6]) );
  XNOR2_X2 add_0_root_sub_0_root_u4_add_496_U31 ( .A(u4_fi_ldz_2a_6_), .B(
        u4_ldz_dif_7_), .ZN(add_0_root_sub_0_root_u4_add_496_n1) );
  INV_X4 add_0_root_sub_0_root_u4_add_496_U30 ( .A(
        add_0_root_sub_0_root_u4_add_496_n6), .ZN(
        add_0_root_sub_0_root_u4_add_496_n3) );
  XNOR2_X2 add_0_root_sub_0_root_u4_add_496_U29 ( .A(
        add_0_root_sub_0_root_u4_add_496_n1), .B(
        add_0_root_sub_0_root_u4_add_496_n2), .ZN(u4_div_exp3[7]) );
  NAND2_X1 add_0_root_sub_0_root_u4_add_496_U28 ( .A1(u4_ldz_dif_0_), .A2(
        n4757), .ZN(add_0_root_sub_0_root_u4_add_496_n58) );
  NAND2_X1 add_0_root_sub_0_root_u4_add_496_U27 ( .A1(n4757), .A2(
        u4_ldz_dif_0_), .ZN(add_0_root_sub_0_root_u4_add_496_n63) );
  OAI21_X1 add_0_root_sub_0_root_u4_add_496_U26 ( .B1(u4_ldz_dif_0_), .B2(
        n4757), .A(add_0_root_sub_0_root_u4_add_496_n63), .ZN(
        add_0_root_sub_0_root_u4_add_496_n66) );
  NAND2_X1 add_0_root_sub_0_root_u4_add_496_U25 ( .A1(u4_fi_ldz_2a_3_), .A2(
        u4_ldz_dif_3_), .ZN(add_0_root_sub_0_root_u4_add_496_n30) );
  NAND2_X1 add_0_root_sub_0_root_u4_add_496_U24 ( .A1(net33106), .A2(
        u4_ldz_dif_1_), .ZN(add_0_root_sub_0_root_u4_add_496_n46) );
  INV_X4 add_0_root_sub_0_root_u4_add_496_U23 ( .A(
        add_0_root_sub_0_root_u4_add_496_n66), .ZN(u4_div_exp3[0]) );
  INV_X4 add_0_root_sub_0_root_u4_add_496_U22 ( .A(
        add_0_root_sub_0_root_u4_add_496_n63), .ZN(
        add_0_root_sub_0_root_u4_add_496_n62) );
  NAND2_X2 add_0_root_sub_0_root_u4_add_496_U21 ( .A1(
        add_0_root_sub_0_root_u4_add_496_n56), .A2(
        add_0_root_sub_0_root_u4_add_496_n46), .ZN(
        add_0_root_sub_0_root_u4_add_496_n52) );
  INV_X1 add_0_root_sub_0_root_u4_add_496_U20 ( .A(net33106), .ZN(
        add_0_root_sub_0_root_u4_add_496_n64) );
  INV_X1 add_0_root_sub_0_root_u4_add_496_U19 ( .A(u4_fi_ldz_2a_3_), .ZN(
        add_0_root_sub_0_root_u4_add_496_n53) );
  NOR2_X2 add_0_root_sub_0_root_u4_add_496_U18 ( .A1(u4_ldz_dif_4_), .A2(
        u4_fi_ldz_2a_4_), .ZN(add_0_root_sub_0_root_u4_add_496_n16) );
  NAND2_X1 add_0_root_sub_0_root_u4_add_496_U17 ( .A1(u4_fi_ldz_2a_4_), .A2(
        u4_ldz_dif_4_), .ZN(add_0_root_sub_0_root_u4_add_496_n14) );
  OAI21_X1 add_0_root_sub_0_root_u4_add_496_U16 ( .B1(u4_ldz_dif_4_), .B2(
        u4_fi_ldz_2a_4_), .A(add_0_root_sub_0_root_u4_add_496_n31), .ZN(
        add_0_root_sub_0_root_u4_add_496_n23) );
  INV_X2 add_0_root_sub_0_root_u4_add_496_U15 ( .A(
        add_0_root_sub_0_root_u4_add_496_n32), .ZN(
        add_0_root_sub_0_root_u4_add_496_n56) );
  INV_X2 add_0_root_sub_0_root_u4_add_496_U14 ( .A(
        add_0_root_sub_0_root_u4_add_496_n30), .ZN(
        add_0_root_sub_0_root_u4_add_496_n40) );
  NOR2_X2 add_0_root_sub_0_root_u4_add_496_U13 ( .A1(
        add_0_root_sub_0_root_u4_add_496_n16), .A2(
        add_0_root_sub_0_root_u4_add_496_n30), .ZN(
        add_0_root_sub_0_root_u4_add_496_n29) );
  OAI21_X2 add_0_root_sub_0_root_u4_add_496_U12 ( .B1(
        add_0_root_sub_0_root_u4_add_496_n3), .B2(
        add_0_root_sub_0_root_u4_add_496_n4), .A(
        add_0_root_sub_0_root_u4_add_496_n5), .ZN(
        add_0_root_sub_0_root_u4_add_496_n2) );
  OAI21_X2 add_0_root_sub_0_root_u4_add_496_U11 ( .B1(
        add_0_root_sub_0_root_u4_add_496_n44), .B2(
        add_0_root_sub_0_root_u4_add_496_n50), .A(
        add_0_root_sub_0_root_u4_add_496_n51), .ZN(
        add_0_root_sub_0_root_u4_add_496_n49) );
  NOR2_X2 add_0_root_sub_0_root_u4_add_496_U10 ( .A1(
        add_0_root_sub_0_root_u4_add_496_n57), .A2(
        add_0_root_sub_0_root_u4_add_496_n58), .ZN(
        add_0_root_sub_0_root_u4_add_496_n32) );
  NOR2_X2 add_0_root_sub_0_root_u4_add_496_U9 ( .A1(
        add_0_root_sub_0_root_u4_add_496_n28), .A2(
        add_0_root_sub_0_root_u4_add_496_n29), .ZN(
        add_0_root_sub_0_root_u4_add_496_n24) );
  NOR2_X2 add_0_root_sub_0_root_u4_add_496_U8 ( .A1(
        add_0_root_sub_0_root_u4_add_496_n42), .A2(
        add_0_root_sub_0_root_u4_add_496_n44), .ZN(
        add_0_root_sub_0_root_u4_add_496_n31) );
  NOR2_X2 add_0_root_sub_0_root_u4_add_496_U7 ( .A1(
        add_0_root_sub_0_root_u4_add_496_n16), .A2(
        add_0_root_sub_0_root_u4_add_496_n17), .ZN(
        add_0_root_sub_0_root_u4_add_496_n9) );
  NOR2_X2 add_0_root_sub_0_root_u4_add_496_U6 ( .A1(
        add_0_root_sub_0_root_u4_add_496_n16), .A2(
        add_0_root_sub_0_root_u4_add_496_n28), .ZN(
        add_0_root_sub_0_root_u4_add_496_n47) );
  NOR2_X4 add_0_root_sub_0_root_u4_add_496_U5 ( .A1(
        add_0_root_sub_0_root_u4_add_496_n32), .A2(
        add_0_root_sub_0_root_u4_add_496_n33), .ZN(
        add_0_root_sub_0_root_u4_add_496_n37) );
  NOR2_X1 add_0_root_sub_0_root_u4_add_496_U4 ( .A1(u4_ldz_dif_2_), .A2(
        net23043), .ZN(add_0_root_sub_0_root_u4_add_496_n44) );
  INV_X1 add_0_root_sub_0_root_u4_add_496_U3 ( .A(net23043), .ZN(
        add_0_root_sub_0_root_u4_add_496_n41) );
  NAND2_X1 add_0_root_sub_0_root_u4_add_496_U2 ( .A1(net23043), .A2(
        u4_ldz_dif_2_), .ZN(add_0_root_sub_0_root_u4_add_496_n51) );
  INV_X4 u4_add_465_U22 ( .A(net85905), .ZN(u4_exp_in_pl1_0_) );
  XNOR2_X2 u4_add_465_U21 ( .A(n3089), .B(u4_add_465_n10), .ZN(
        u4_exp_in_pl1_2_) );
  XNOR2_X2 u4_add_465_U20 ( .A(n3088), .B(u4_add_465_n12), .ZN(
        u4_exp_in_pl1_3_) );
  NAND2_X2 u4_add_465_U19 ( .A1(n3088), .A2(n3089), .ZN(u4_add_465_n11) );
  INV_X4 u4_add_465_U18 ( .A(n3085), .ZN(u4_add_465_n9) );
  XNOR2_X2 u4_add_465_U17 ( .A(u4_add_465_n7), .B(u4_add_465_n9), .ZN(
        u4_exp_in_pl1_4_) );
  NAND2_X2 u4_add_465_U16 ( .A1(n3085), .A2(u4_add_465_n7), .ZN(u4_add_465_n8)
         );
  XNOR2_X2 u4_add_465_U15 ( .A(exp_r[5]), .B(u4_add_465_n8), .ZN(
        u4_exp_in_pl1_5_) );
  NAND3_X4 u4_add_465_U14 ( .A1(exp_r[5]), .A2(n3085), .A3(u4_add_465_n7), 
        .ZN(u4_add_465_n3) );
  XNOR2_X2 u4_add_465_U13 ( .A(net85933), .B(u4_add_465_n3), .ZN(
        u4_exp_in_pl1_6_) );
  INV_X4 u4_add_465_U12 ( .A(net85933), .ZN(u4_add_465_n6) );
  NOR2_X4 u4_add_465_U11 ( .A1(u4_add_465_n3), .A2(u4_add_465_n6), .ZN(
        u4_add_465_n4) );
  INV_X4 u4_add_465_U10 ( .A(net85937), .ZN(u4_add_465_n5) );
  XNOR2_X2 u4_add_465_U9 ( .A(u4_add_465_n4), .B(u4_add_465_n5), .ZN(
        u4_exp_in_pl1_7_) );
  INV_X4 u4_add_465_U8 ( .A(u4_add_465_n3), .ZN(u4_add_465_n2) );
  INV_X4 u4_add_465_U7 ( .A(u4_add_465_n1), .ZN(u4_exp_in_pl1_8_) );
  NAND3_X1 u4_add_465_U6 ( .A1(n3089), .A2(net85905), .A3(n3091), .ZN(
        u4_add_465_n12) );
  NAND2_X1 u4_add_465_U5 ( .A1(n3091), .A2(net85905), .ZN(u4_add_465_n10) );
  XOR2_X2 u4_add_465_U4 ( .A(n3091), .B(net85905), .Z(u4_exp_in_pl1_1_) );
  NAND3_X2 u4_add_465_U3 ( .A1(net85933), .A2(net85937), .A3(u4_add_465_n2), 
        .ZN(u4_add_465_n1) );
  NOR2_X2 u4_add_465_U2 ( .A1(u4_add_465_n10), .A2(u4_add_465_n11), .ZN(
        u4_add_465_n7) );
  INV_X4 sub_1_root_u1_sub_130_aco_U109 ( .A(u1_exp_small[0]), .ZN(
        sub_1_root_u1_sub_130_aco_n69) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U108 ( .A1(n5316), .A2(
        sub_1_root_u1_sub_130_aco_n69), .ZN(sub_1_root_u1_sub_130_aco_n99) );
  INV_X4 sub_1_root_u1_sub_130_aco_U107 ( .A(sub_1_root_u1_sub_130_aco_n99), 
        .ZN(sub_1_root_u1_sub_130_aco_n96) );
  NOR2_X4 sub_1_root_u1_sub_130_aco_U106 ( .A1(sub_1_root_u1_sub_130_aco_n96), 
        .A2(sub_1_root_u1_sub_130_aco_n98), .ZN(sub_1_root_u1_sub_130_aco_n97)
         );
  XNOR2_X2 sub_1_root_u1_sub_130_aco_U105 ( .A(n5317), .B(
        sub_1_root_u1_sub_130_aco_n97), .ZN(u1_exp_diff2[0]) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U104 ( .A1(u1_exp_small[0]), .A2(
        sub_1_root_u1_sub_130_aco_n52), .ZN(sub_1_root_u1_sub_130_aco_n95) );
  AOI21_X4 sub_1_root_u1_sub_130_aco_U103 ( .B1(sub_1_root_u1_sub_130_aco_n95), 
        .B2(sub_1_root_u1_sub_130_aco_n53), .A(sub_1_root_u1_sub_130_aco_n96), 
        .ZN(sub_1_root_u1_sub_130_aco_n91) );
  INV_X4 sub_1_root_u1_sub_130_aco_U102 ( .A(n5315), .ZN(
        sub_1_root_u1_sub_130_aco_n94) );
  INV_X4 sub_1_root_u1_sub_130_aco_U101 ( .A(u1_exp_small[1]), .ZN(
        sub_1_root_u1_sub_130_aco_n93) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U100 ( .A1(n5315), .A2(
        sub_1_root_u1_sub_130_aco_n93), .ZN(sub_1_root_u1_sub_130_aco_n10) );
  INV_X4 sub_1_root_u1_sub_130_aco_U99 ( .A(sub_1_root_u1_sub_130_aco_n10), 
        .ZN(sub_1_root_u1_sub_130_aco_n38) );
  XNOR2_X2 sub_1_root_u1_sub_130_aco_U98 ( .A(sub_1_root_u1_sub_130_aco_n91), 
        .B(sub_1_root_u1_sub_130_aco_n92), .ZN(u1_exp_diff2[1]) );
  INV_X4 sub_1_root_u1_sub_130_aco_U97 ( .A(n5314), .ZN(
        sub_1_root_u1_sub_130_aco_n90) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U96 ( .A1(u1_exp_small[2]), .A2(
        sub_1_root_u1_sub_130_aco_n90), .ZN(sub_1_root_u1_sub_130_aco_n71) );
  INV_X4 sub_1_root_u1_sub_130_aco_U95 ( .A(u1_exp_small[2]), .ZN(
        sub_1_root_u1_sub_130_aco_n89) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U94 ( .A1(n5314), .A2(
        sub_1_root_u1_sub_130_aco_n89), .ZN(sub_1_root_u1_sub_130_aco_n66) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U93 ( .A1(sub_1_root_u1_sub_130_aco_n71), 
        .A2(sub_1_root_u1_sub_130_aco_n66), .ZN(sub_1_root_u1_sub_130_aco_n83)
         );
  INV_X4 sub_1_root_u1_sub_130_aco_U92 ( .A(n5317), .ZN(
        sub_1_root_u1_sub_130_aco_n53) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U91 ( .A1(u1_exp_small[0]), .A2(
        sub_1_root_u1_sub_130_aco_n52), .ZN(sub_1_root_u1_sub_130_aco_n87) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U90 ( .A1(sub_1_root_u1_sub_130_aco_n85), 
        .A2(sub_1_root_u1_sub_130_aco_n86), .ZN(sub_1_root_u1_sub_130_aco_n84)
         );
  XNOR2_X2 sub_1_root_u1_sub_130_aco_U89 ( .A(sub_1_root_u1_sub_130_aco_n83), 
        .B(sub_1_root_u1_sub_130_aco_n84), .ZN(u1_exp_diff2[2]) );
  NOR2_X4 sub_1_root_u1_sub_130_aco_U88 ( .A1(sub_1_root_u1_sub_130_aco_n80), 
        .A2(sub_1_root_u1_sub_130_aco_n81), .ZN(sub_1_root_u1_sub_130_aco_n78)
         );
  INV_X4 sub_1_root_u1_sub_130_aco_U87 ( .A(sub_1_root_u1_sub_130_aco_n71), 
        .ZN(sub_1_root_u1_sub_130_aco_n79) );
  AOI211_X4 sub_1_root_u1_sub_130_aco_U86 ( .C1(sub_1_root_u1_sub_130_aco_n77), 
        .C2(sub_1_root_u1_sub_130_aco_n78), .A(sub_1_root_u1_sub_130_aco_n79), 
        .B(sub_1_root_u1_sub_130_aco_n70), .ZN(sub_1_root_u1_sub_130_aco_n75)
         );
  INV_X4 sub_1_root_u1_sub_130_aco_U85 ( .A(sub_1_root_u1_sub_130_aco_n66), 
        .ZN(sub_1_root_u1_sub_130_aco_n76) );
  NOR2_X4 sub_1_root_u1_sub_130_aco_U84 ( .A1(sub_1_root_u1_sub_130_aco_n75), 
        .A2(sub_1_root_u1_sub_130_aco_n76), .ZN(sub_1_root_u1_sub_130_aco_n73)
         );
  INV_X4 sub_1_root_u1_sub_130_aco_U83 ( .A(n5313), .ZN(
        sub_1_root_u1_sub_130_aco_n64) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U82 ( .A1(u1_exp_small[3]), .A2(
        sub_1_root_u1_sub_130_aco_n64), .ZN(sub_1_root_u1_sub_130_aco_n72) );
  INV_X4 sub_1_root_u1_sub_130_aco_U81 ( .A(u1_exp_small[3]), .ZN(
        sub_1_root_u1_sub_130_aco_n74) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U80 ( .A1(n5313), .A2(
        sub_1_root_u1_sub_130_aco_n74), .ZN(sub_1_root_u1_sub_130_aco_n65) );
  XNOR2_X2 sub_1_root_u1_sub_130_aco_U79 ( .A(sub_1_root_u1_sub_130_aco_n73), 
        .B(sub_1_root_u1_sub_130_aco_n1), .ZN(u1_exp_diff2[3]) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U78 ( .A1(sub_1_root_u1_sub_130_aco_n71), 
        .A2(sub_1_root_u1_sub_130_aco_n72), .ZN(sub_1_root_u1_sub_130_aco_n13)
         );
  NOR2_X4 sub_1_root_u1_sub_130_aco_U77 ( .A1(sub_1_root_u1_sub_130_aco_n70), 
        .A2(sub_1_root_u1_sub_130_aco_n13), .ZN(sub_1_root_u1_sub_130_aco_n61)
         );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U76 ( .A1(n5316), .A2(
        sub_1_root_u1_sub_130_aco_n69), .ZN(sub_1_root_u1_sub_130_aco_n67) );
  NAND3_X2 sub_1_root_u1_sub_130_aco_U75 ( .A1(sub_1_root_u1_sub_130_aco_n67), 
        .A2(sub_1_root_u1_sub_130_aco_n10), .A3(sub_1_root_u1_sub_130_aco_n68), 
        .ZN(sub_1_root_u1_sub_130_aco_n62) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U74 ( .A1(sub_1_root_u1_sub_130_aco_n65), 
        .A2(sub_1_root_u1_sub_130_aco_n66), .ZN(sub_1_root_u1_sub_130_aco_n17)
         );
  INV_X4 sub_1_root_u1_sub_130_aco_U73 ( .A(sub_1_root_u1_sub_130_aco_n17), 
        .ZN(sub_1_root_u1_sub_130_aco_n33) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U72 ( .A1(u1_exp_small[3]), .A2(
        sub_1_root_u1_sub_130_aco_n64), .ZN(sub_1_root_u1_sub_130_aco_n16) );
  INV_X4 sub_1_root_u1_sub_130_aco_U71 ( .A(sub_1_root_u1_sub_130_aco_n16), 
        .ZN(sub_1_root_u1_sub_130_aco_n34) );
  NOR2_X4 sub_1_root_u1_sub_130_aco_U70 ( .A1(sub_1_root_u1_sub_130_aco_n33), 
        .A2(sub_1_root_u1_sub_130_aco_n34), .ZN(sub_1_root_u1_sub_130_aco_n63)
         );
  AOI21_X4 sub_1_root_u1_sub_130_aco_U69 ( .B1(sub_1_root_u1_sub_130_aco_n61), 
        .B2(sub_1_root_u1_sub_130_aco_n62), .A(sub_1_root_u1_sub_130_aco_n63), 
        .ZN(sub_1_root_u1_sub_130_aco_n57) );
  INV_X4 sub_1_root_u1_sub_130_aco_U68 ( .A(n5312), .ZN(
        sub_1_root_u1_sub_130_aco_n60) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U67 ( .A1(u1_exp_small[4]), .A2(
        sub_1_root_u1_sub_130_aco_n60), .ZN(sub_1_root_u1_sub_130_aco_n36) );
  INV_X4 sub_1_root_u1_sub_130_aco_U66 ( .A(sub_1_root_u1_sub_130_aco_n36), 
        .ZN(sub_1_root_u1_sub_130_aco_n49) );
  INV_X4 sub_1_root_u1_sub_130_aco_U65 ( .A(u1_exp_small[4]), .ZN(
        sub_1_root_u1_sub_130_aco_n59) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U64 ( .A1(n5312), .A2(
        sub_1_root_u1_sub_130_aco_n59), .ZN(sub_1_root_u1_sub_130_aco_n24) );
  INV_X4 sub_1_root_u1_sub_130_aco_U63 ( .A(sub_1_root_u1_sub_130_aco_n24), 
        .ZN(sub_1_root_u1_sub_130_aco_n47) );
  XNOR2_X2 sub_1_root_u1_sub_130_aco_U62 ( .A(sub_1_root_u1_sub_130_aco_n57), 
        .B(sub_1_root_u1_sub_130_aco_n58), .ZN(u1_exp_diff2[4]) );
  INV_X4 sub_1_root_u1_sub_130_aco_U61 ( .A(u1_exp_small[5]), .ZN(
        sub_1_root_u1_sub_130_aco_n56) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U60 ( .A1(n5311), .A2(
        sub_1_root_u1_sub_130_aco_n56), .ZN(sub_1_root_u1_sub_130_aco_n21) );
  INV_X4 sub_1_root_u1_sub_130_aco_U59 ( .A(n5311), .ZN(
        sub_1_root_u1_sub_130_aco_n55) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U58 ( .A1(u1_exp_small[5]), .A2(
        sub_1_root_u1_sub_130_aco_n55), .ZN(sub_1_root_u1_sub_130_aco_n32) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U57 ( .A1(sub_1_root_u1_sub_130_aco_n21), 
        .A2(sub_1_root_u1_sub_130_aco_n32), .ZN(sub_1_root_u1_sub_130_aco_n42)
         );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U56 ( .A1(u1_exp_small[0]), .A2(
        sub_1_root_u1_sub_130_aco_n52), .ZN(sub_1_root_u1_sub_130_aco_n54) );
  NAND3_X2 sub_1_root_u1_sub_130_aco_U55 ( .A1(sub_1_root_u1_sub_130_aco_n51), 
        .A2(sub_1_root_u1_sub_130_aco_n53), .A3(sub_1_root_u1_sub_130_aco_n54), 
        .ZN(sub_1_root_u1_sub_130_aco_n11) );
  INV_X4 sub_1_root_u1_sub_130_aco_U54 ( .A(sub_1_root_u1_sub_130_aco_n11), 
        .ZN(sub_1_root_u1_sub_130_aco_n37) );
  INV_X4 sub_1_root_u1_sub_130_aco_U53 ( .A(sub_1_root_u1_sub_130_aco_n12), 
        .ZN(sub_1_root_u1_sub_130_aco_n39) );
  NOR3_X4 sub_1_root_u1_sub_130_aco_U52 ( .A1(sub_1_root_u1_sub_130_aco_n37), 
        .A2(sub_1_root_u1_sub_130_aco_n38), .A3(sub_1_root_u1_sub_130_aco_n39), 
        .ZN(sub_1_root_u1_sub_130_aco_n44) );
  INV_X4 sub_1_root_u1_sub_130_aco_U51 ( .A(sub_1_root_u1_sub_130_aco_n13), 
        .ZN(sub_1_root_u1_sub_130_aco_n35) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U50 ( .A1(sub_1_root_u1_sub_130_aco_n35), 
        .A2(sub_1_root_u1_sub_130_aco_n36), .ZN(sub_1_root_u1_sub_130_aco_n45)
         );
  NOR3_X4 sub_1_root_u1_sub_130_aco_U49 ( .A1(sub_1_root_u1_sub_130_aco_n33), 
        .A2(sub_1_root_u1_sub_130_aco_n49), .A3(sub_1_root_u1_sub_130_aco_n34), 
        .ZN(sub_1_root_u1_sub_130_aco_n48) );
  NOR2_X4 sub_1_root_u1_sub_130_aco_U48 ( .A1(sub_1_root_u1_sub_130_aco_n47), 
        .A2(sub_1_root_u1_sub_130_aco_n48), .ZN(sub_1_root_u1_sub_130_aco_n46)
         );
  OAI21_X4 sub_1_root_u1_sub_130_aco_U47 ( .B1(sub_1_root_u1_sub_130_aco_n44), 
        .B2(sub_1_root_u1_sub_130_aco_n45), .A(sub_1_root_u1_sub_130_aco_n46), 
        .ZN(sub_1_root_u1_sub_130_aco_n43) );
  XNOR2_X2 sub_1_root_u1_sub_130_aco_U46 ( .A(sub_1_root_u1_sub_130_aco_n42), 
        .B(sub_1_root_u1_sub_130_aco_n43), .ZN(u1_exp_diff2[5]) );
  INV_X4 sub_1_root_u1_sub_130_aco_U45 ( .A(u1_exp_small[6]), .ZN(
        sub_1_root_u1_sub_130_aco_n41) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U44 ( .A1(n5310), .A2(
        sub_1_root_u1_sub_130_aco_n41), .ZN(sub_1_root_u1_sub_130_aco_n22) );
  INV_X4 sub_1_root_u1_sub_130_aco_U43 ( .A(n5310), .ZN(
        sub_1_root_u1_sub_130_aco_n40) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U42 ( .A1(u1_exp_small[6]), .A2(
        sub_1_root_u1_sub_130_aco_n40), .ZN(sub_1_root_u1_sub_130_aco_n8) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U41 ( .A1(sub_1_root_u1_sub_130_aco_n22), 
        .A2(sub_1_root_u1_sub_130_aco_n8), .ZN(sub_1_root_u1_sub_130_aco_n25)
         );
  NOR3_X4 sub_1_root_u1_sub_130_aco_U40 ( .A1(sub_1_root_u1_sub_130_aco_n37), 
        .A2(sub_1_root_u1_sub_130_aco_n38), .A3(sub_1_root_u1_sub_130_aco_n39), 
        .ZN(sub_1_root_u1_sub_130_aco_n27) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U39 ( .A1(sub_1_root_u1_sub_130_aco_n36), 
        .A2(sub_1_root_u1_sub_130_aco_n32), .ZN(sub_1_root_u1_sub_130_aco_n14)
         );
  INV_X4 sub_1_root_u1_sub_130_aco_U38 ( .A(sub_1_root_u1_sub_130_aco_n14), 
        .ZN(sub_1_root_u1_sub_130_aco_n15) );
  NAND2_X2 sub_1_root_u1_sub_130_aco_U37 ( .A1(sub_1_root_u1_sub_130_aco_n15), 
        .A2(sub_1_root_u1_sub_130_aco_n35), .ZN(sub_1_root_u1_sub_130_aco_n28)
         );
  NOR2_X4 sub_1_root_u1_sub_130_aco_U36 ( .A1(sub_1_root_u1_sub_130_aco_n33), 
        .A2(sub_1_root_u1_sub_130_aco_n34), .ZN(sub_1_root_u1_sub_130_aco_n30)
         );
  INV_X4 sub_1_root_u1_sub_130_aco_U35 ( .A(sub_1_root_u1_sub_130_aco_n32), 
        .ZN(sub_1_root_u1_sub_130_aco_n23) );
  AOI21_X4 sub_1_root_u1_sub_130_aco_U34 ( .B1(sub_1_root_u1_sub_130_aco_n24), 
        .B2(sub_1_root_u1_sub_130_aco_n21), .A(sub_1_root_u1_sub_130_aco_n23), 
        .ZN(sub_1_root_u1_sub_130_aco_n31) );
  AOI21_X4 sub_1_root_u1_sub_130_aco_U33 ( .B1(sub_1_root_u1_sub_130_aco_n30), 
        .B2(sub_1_root_u1_sub_130_aco_n15), .A(sub_1_root_u1_sub_130_aco_n31), 
        .ZN(sub_1_root_u1_sub_130_aco_n29) );
  XNOR2_X2 sub_1_root_u1_sub_130_aco_U32 ( .A(sub_1_root_u1_sub_130_aco_n25), 
        .B(sub_1_root_u1_sub_130_aco_n26), .ZN(u1_exp_diff2[6]) );
  INV_X4 sub_1_root_u1_sub_130_aco_U31 ( .A(sub_1_root_u1_sub_130_aco_n8), 
        .ZN(sub_1_root_u1_sub_130_aco_n20) );
  NAND4_X2 sub_1_root_u1_sub_130_aco_U30 ( .A1(sub_1_root_u1_sub_130_aco_n15), 
        .A2(sub_1_root_u1_sub_130_aco_n16), .A3(sub_1_root_u1_sub_130_aco_n17), 
        .A4(sub_1_root_u1_sub_130_aco_n8), .ZN(sub_1_root_u1_sub_130_aco_n5)
         );
  NAND3_X4 sub_1_root_u1_sub_130_aco_U29 ( .A1(sub_1_root_u1_sub_130_aco_n7), 
        .A2(sub_1_root_u1_sub_130_aco_n8), .A3(sub_1_root_u1_sub_130_aco_n9), 
        .ZN(sub_1_root_u1_sub_130_aco_n6) );
  XNOR2_X2 sub_1_root_u1_sub_130_aco_U28 ( .A(sub_1_root_u1_sub_130_aco_n2), 
        .B(sub_1_root_u1_sub_130_aco_n3), .ZN(u1_exp_diff2[7]) );
  NAND2_X4 sub_1_root_u1_sub_130_aco_U27 ( .A1(u1_exp_small[1]), .A2(
        sub_1_root_u1_sub_130_aco_n94), .ZN(sub_1_root_u1_sub_130_aco_n51) );
  NAND2_X4 sub_1_root_u1_sub_130_aco_U26 ( .A1(sub_1_root_u1_sub_130_aco_n50), 
        .A2(sub_1_root_u1_sub_130_aco_n51), .ZN(sub_1_root_u1_sub_130_aco_n12)
         );
  NAND3_X1 sub_1_root_u1_sub_130_aco_U25 ( .A1(sub_1_root_u1_sub_130_aco_n51), 
        .A2(sub_1_root_u1_sub_130_aco_n53), .A3(sub_1_root_u1_sub_130_aco_n87), 
        .ZN(sub_1_root_u1_sub_130_aco_n86) );
  AOI21_X2 sub_1_root_u1_sub_130_aco_U24 ( .B1(sub_1_root_u1_sub_130_aco_n88), 
        .B2(sub_1_root_u1_sub_130_aco_n51), .A(sub_1_root_u1_sub_130_aco_n38), 
        .ZN(sub_1_root_u1_sub_130_aco_n85) );
  INV_X8 sub_1_root_u1_sub_130_aco_U23 ( .A(sub_1_root_u1_sub_130_aco_n51), 
        .ZN(sub_1_root_u1_sub_130_aco_n70) );
  XOR2_X1 sub_1_root_u1_sub_130_aco_U22 ( .A(u1_exp_small[7]), .B(n5309), .Z(
        sub_1_root_u1_sub_130_aco_n2) );
  AND2_X2 sub_1_root_u1_sub_130_aco_U21 ( .A1(sub_1_root_u1_sub_130_aco_n72), 
        .A2(sub_1_root_u1_sub_130_aco_n65), .ZN(sub_1_root_u1_sub_130_aco_n1)
         );
  OAI21_X1 sub_1_root_u1_sub_130_aco_U20 ( .B1(n5316), .B2(
        sub_1_root_u1_sub_130_aco_n69), .A(sub_1_root_u1_sub_130_aco_n53), 
        .ZN(sub_1_root_u1_sub_130_aco_n68) );
  OAI21_X2 sub_1_root_u1_sub_130_aco_U19 ( .B1(sub_1_root_u1_sub_130_aco_n27), 
        .B2(sub_1_root_u1_sub_130_aco_n28), .A(sub_1_root_u1_sub_130_aco_n29), 
        .ZN(sub_1_root_u1_sub_130_aco_n26) );
  NOR2_X2 sub_1_root_u1_sub_130_aco_U18 ( .A1(sub_1_root_u1_sub_130_aco_n18), 
        .A2(sub_1_root_u1_sub_130_aco_n19), .ZN(sub_1_root_u1_sub_130_aco_n4)
         );
  NAND3_X2 sub_1_root_u1_sub_130_aco_U17 ( .A1(sub_1_root_u1_sub_130_aco_n4), 
        .A2(sub_1_root_u1_sub_130_aco_n5), .A3(sub_1_root_u1_sub_130_aco_n6), 
        .ZN(sub_1_root_u1_sub_130_aco_n3) );
  NOR2_X2 sub_1_root_u1_sub_130_aco_U16 ( .A1(sub_1_root_u1_sub_130_aco_n38), 
        .A2(sub_1_root_u1_sub_130_aco_n82), .ZN(sub_1_root_u1_sub_130_aco_n77)
         );
  NOR2_X1 sub_1_root_u1_sub_130_aco_U15 ( .A1(u1_exp_small[0]), .A2(
        sub_1_root_u1_sub_130_aco_n52), .ZN(sub_1_root_u1_sub_130_aco_n88) );
  NOR2_X2 sub_1_root_u1_sub_130_aco_U14 ( .A1(sub_1_root_u1_sub_130_aco_n49), 
        .A2(sub_1_root_u1_sub_130_aco_n47), .ZN(sub_1_root_u1_sub_130_aco_n58)
         );
  NOR3_X2 sub_1_root_u1_sub_130_aco_U13 ( .A1(sub_1_root_u1_sub_130_aco_n23), 
        .A2(sub_1_root_u1_sub_130_aco_n24), .A3(sub_1_root_u1_sub_130_aco_n20), 
        .ZN(sub_1_root_u1_sub_130_aco_n18) );
  OAI21_X2 sub_1_root_u1_sub_130_aco_U12 ( .B1(sub_1_root_u1_sub_130_aco_n20), 
        .B2(sub_1_root_u1_sub_130_aco_n21), .A(sub_1_root_u1_sub_130_aco_n22), 
        .ZN(sub_1_root_u1_sub_130_aco_n19) );
  NOR2_X2 sub_1_root_u1_sub_130_aco_U11 ( .A1(sub_1_root_u1_sub_130_aco_n13), 
        .A2(sub_1_root_u1_sub_130_aco_n14), .ZN(sub_1_root_u1_sub_130_aco_n7)
         );
  NAND3_X2 sub_1_root_u1_sub_130_aco_U10 ( .A1(sub_1_root_u1_sub_130_aco_n10), 
        .A2(sub_1_root_u1_sub_130_aco_n11), .A3(sub_1_root_u1_sub_130_aco_n12), 
        .ZN(sub_1_root_u1_sub_130_aco_n9) );
  NOR2_X1 sub_1_root_u1_sub_130_aco_U9 ( .A1(u1_exp_small[0]), .A2(
        sub_1_root_u1_sub_130_aco_n52), .ZN(sub_1_root_u1_sub_130_aco_n82) );
  NOR2_X1 sub_1_root_u1_sub_130_aco_U8 ( .A1(n5317), .A2(u1_exp_small[0]), 
        .ZN(sub_1_root_u1_sub_130_aco_n81) );
  NOR2_X1 sub_1_root_u1_sub_130_aco_U7 ( .A1(n5317), .A2(
        sub_1_root_u1_sub_130_aco_n52), .ZN(sub_1_root_u1_sub_130_aco_n80) );
  NOR2_X2 sub_1_root_u1_sub_130_aco_U6 ( .A1(n5316), .A2(
        sub_1_root_u1_sub_130_aco_n69), .ZN(sub_1_root_u1_sub_130_aco_n98) );
  NOR2_X2 sub_1_root_u1_sub_130_aco_U5 ( .A1(sub_1_root_u1_sub_130_aco_n70), 
        .A2(sub_1_root_u1_sub_130_aco_n38), .ZN(sub_1_root_u1_sub_130_aco_n92)
         );
  INV_X8 sub_1_root_u1_sub_130_aco_U4 ( .A(n5316), .ZN(
        sub_1_root_u1_sub_130_aco_n52) );
  NOR2_X2 sub_1_root_u1_sub_130_aco_U3 ( .A1(u1_exp_small[0]), .A2(
        sub_1_root_u1_sub_130_aco_n52), .ZN(sub_1_root_u1_sub_130_aco_n50) );
  NOR2_X4 u4_sub_469_U72 ( .A1(u4_sub_469_n59), .A2(u4_sub_469_n60), .ZN(
        u4_sub_469_n55) );
  INV_X4 u4_sub_469_U71 ( .A(u4_exp_in_pl1_1_), .ZN(u4_sub_469_n58) );
  XNOR2_X2 u4_sub_469_U70 ( .A(u4_sub_469_n55), .B(u4_sub_469_n56), .ZN(
        u4_exp_next_mi_1_) );
  AOI21_X4 u4_sub_469_U69 ( .B1(u4_sub_469_n51), .B2(u4_sub_469_n52), .A(
        u4_sub_469_n11), .ZN(u4_sub_469_n45) );
  INV_X4 u4_sub_469_U68 ( .A(u4_exp_in_pl1_2_), .ZN(u4_sub_469_n49) );
  OAI21_X4 u4_sub_469_U67 ( .B1(u4_sub_469_n9), .B2(u4_sub_469_n45), .A(
        u4_sub_469_n46), .ZN(u4_sub_469_n44) );
  INV_X4 u4_sub_469_U66 ( .A(u4_exp_in_pl1_3_), .ZN(u4_sub_469_n42) );
  NOR2_X4 u4_sub_469_U65 ( .A1(u4_sub_469_n40), .A2(u4_sub_469_n36), .ZN(
        u4_sub_469_n39) );
  OAI21_X4 u4_sub_469_U64 ( .B1(u4_sub_469_n37), .B2(u4_sub_469_n36), .A(
        u4_sub_469_n38), .ZN(u4_sub_469_n35) );
  INV_X4 u4_sub_469_U63 ( .A(u4_exp_in_pl1_4_), .ZN(u4_sub_469_n33) );
  NAND2_X2 u4_sub_469_U62 ( .A1(u4_fi_ldz_mi1_4_), .A2(u4_sub_469_n33), .ZN(
        u4_sub_469_n32) );
  INV_X4 u4_sub_469_U61 ( .A(u4_fi_ldz_mi1_5_), .ZN(u4_sub_469_n27) );
  INV_X4 u4_sub_469_U60 ( .A(u4_exp_in_pl1_5_), .ZN(u4_sub_469_n26) );
  NAND2_X2 u4_sub_469_U59 ( .A1(u4_fi_ldz_mi1_5_), .A2(u4_sub_469_n26), .ZN(
        u4_sub_469_n25) );
  INV_X4 u4_sub_469_U58 ( .A(u4_sub_469_n25), .ZN(u4_sub_469_n22) );
  NOR2_X4 u4_sub_469_U57 ( .A1(u4_sub_469_n2), .A2(u4_sub_469_n22), .ZN(
        u4_sub_469_n24) );
  XNOR2_X2 u4_sub_469_U56 ( .A(u4_sub_469_n23), .B(u4_sub_469_n24), .ZN(
        u4_exp_next_mi_5_) );
  XNOR2_X2 u4_sub_469_U55 ( .A(u4_sub_469_n6), .B(u4_sub_469_n21), .ZN(
        u4_exp_next_mi_6_) );
  INV_X4 u4_sub_469_U54 ( .A(u4_sub_469_n17), .ZN(u4_sub_469_n19) );
  XNOR2_X2 u4_sub_469_U53 ( .A(u4_sub_469_n20), .B(u4_sub_469_n19), .ZN(
        u4_exp_next_mi_7_) );
  INV_X4 u4_sub_469_U52 ( .A(u4_sub_469_n18), .ZN(u4_sub_469_n17) );
  XNOR2_X2 u4_sub_469_U51 ( .A(u4_sub_469_n14), .B(u4_sub_469_n15), .ZN(
        u4_exp_next_mi_8_) );
  INV_X8 u4_sub_469_U50 ( .A(u4_sub_469_n44), .ZN(u4_sub_469_n37) );
  NAND2_X4 u4_sub_469_U49 ( .A1(u4_sub_469_n50), .A2(u4_exp_in_pl1_2_), .ZN(
        u4_sub_469_n46) );
  INV_X2 u4_sub_469_U48 ( .A(u4_sub_469_n53), .ZN(u4_sub_469_n60) );
  INV_X1 u4_sub_469_U47 ( .A(u4_sub_469_n54), .ZN(u4_sub_469_n59) );
  INV_X4 u4_sub_469_U46 ( .A(u4_exp_in_pl1_8_), .ZN(u4_sub_469_n15) );
  NOR2_X4 u4_sub_469_U45 ( .A1(u4_sub_469_n61), .A2(u4_exp_in_pl1_0_), .ZN(
        u4_sub_469_n54) );
  INV_X4 u4_sub_469_U44 ( .A(u4_exp_in_pl1_6_), .ZN(u4_sub_469_n21) );
  INV_X4 u4_sub_469_U43 ( .A(u4_exp_in_pl1_7_), .ZN(u4_sub_469_n18) );
  NAND2_X4 u4_sub_469_U42 ( .A1(u4_sub_469_n6), .A2(u4_sub_469_n21), .ZN(
        u4_sub_469_n16) );
  INV_X4 u4_sub_469_U41 ( .A(u4_fi_ldz_mi1_3_), .ZN(u4_sub_469_n43) );
  NAND2_X4 u4_sub_469_U40 ( .A1(u4_sub_469_n43), .A2(u4_exp_in_pl1_3_), .ZN(
        u4_sub_469_n38) );
  NAND2_X4 u4_sub_469_U39 ( .A1(u4_exp_in_pl1_4_), .A2(u4_sub_469_n34), .ZN(
        u4_sub_469_n30) );
  INV_X2 u4_sub_469_U38 ( .A(u4_sub_469_n51), .ZN(u4_sub_469_n57) );
  INV_X4 u4_sub_469_U37 ( .A(u4_fi_ldz_mi1_4_), .ZN(u4_sub_469_n34) );
  NAND2_X4 u4_sub_469_U36 ( .A1(u4_sub_469_n12), .A2(u4_sub_469_n13), .ZN(
        u4_exp_next_mi_4_) );
  NAND2_X2 u4_sub_469_U35 ( .A1(u4_sub_469_n42), .A2(u4_fi_ldz_mi1_3_), .ZN(
        u4_sub_469_n41) );
  NOR2_X4 u4_sub_469_U34 ( .A1(u4_sub_469_n50), .A2(u4_sub_469_n10), .ZN(
        u4_sub_469_n9) );
  NAND2_X4 u4_sub_469_U33 ( .A1(u4_fi_ldz_mi1_1_), .A2(u4_sub_469_n58), .ZN(
        u4_sub_469_n51) );
  NOR2_X4 u4_sub_469_U32 ( .A1(u4_fi_ldz_mi1_1_), .A2(u4_sub_469_n58), .ZN(
        u4_sub_469_n11) );
  INV_X8 u4_sub_469_U31 ( .A(n4757), .ZN(u4_sub_469_n61) );
  NAND2_X4 u4_sub_469_U30 ( .A1(u4_exp_in_pl1_0_), .A2(u4_sub_469_n61), .ZN(
        u4_sub_469_n53) );
  NOR2_X4 u4_sub_469_U29 ( .A1(u4_sub_469_n16), .A2(u4_sub_469_n17), .ZN(
        u4_sub_469_n14) );
  INV_X4 u4_sub_469_U28 ( .A(u4_sub_469_n8), .ZN(u4_sub_469_n31) );
  NAND2_X4 u4_sub_469_U27 ( .A1(u4_sub_469_n30), .A2(u4_sub_469_n32), .ZN(
        u4_sub_469_n8) );
  NAND2_X2 u4_sub_469_U26 ( .A1(u4_sub_469_n8), .A2(u4_sub_469_n35), .ZN(
        u4_sub_469_n13) );
  NOR2_X1 u4_sub_469_U25 ( .A1(u4_exp_in_pl1_0_), .A2(u4_sub_469_n61), .ZN(
        u4_sub_469_n62) );
  NAND2_X2 u4_sub_469_U24 ( .A1(u4_sub_469_n31), .A2(u4_sub_469_n1), .ZN(
        u4_sub_469_n12) );
  NOR2_X2 u4_sub_469_U23 ( .A1(u4_sub_469_n48), .A2(u4_sub_469_n9), .ZN(
        u4_sub_469_n47) );
  XNOR2_X2 u4_sub_469_U22 ( .A(u4_sub_469_n47), .B(u4_sub_469_n5), .ZN(
        u4_exp_next_mi_2_) );
  AOI21_X4 u4_sub_469_U21 ( .B1(u4_sub_469_n4), .B2(u4_sub_469_n25), .A(
        u4_sub_469_n2), .ZN(u4_sub_469_n6) );
  INV_X4 u4_sub_469_U20 ( .A(u4_sub_469_n32), .ZN(u4_sub_469_n29) );
  OAI21_X4 u4_sub_469_U19 ( .B1(u4_sub_469_n1), .B2(u4_sub_469_n29), .A(
        u4_sub_469_n30), .ZN(u4_sub_469_n4) );
  OR2_X4 u4_sub_469_U18 ( .A1(u4_sub_469_n60), .A2(u4_sub_469_n62), .ZN(
        u4_exp_next_mi_0_) );
  AND2_X2 u4_sub_469_U17 ( .A1(u4_exp_in_pl1_5_), .A2(u4_sub_469_n27), .ZN(
        u4_sub_469_n2) );
  INV_X4 u4_sub_469_U16 ( .A(u4_sub_469_n49), .ZN(u4_sub_469_n10) );
  NAND2_X2 u4_sub_469_U15 ( .A1(u4_sub_469_n53), .A2(u4_sub_469_n54), .ZN(
        u4_sub_469_n52) );
  INV_X8 u4_sub_469_U14 ( .A(u4_sub_469_n38), .ZN(u4_sub_469_n40) );
  INV_X4 u4_sub_469_U13 ( .A(u4_sub_469_n28), .ZN(u4_sub_469_n23) );
  NOR2_X4 u4_sub_469_U12 ( .A1(u4_sub_469_n57), .A2(u4_sub_469_n7), .ZN(
        u4_sub_469_n56) );
  INV_X2 u4_sub_469_U11 ( .A(u4_sub_469_n46), .ZN(u4_sub_469_n48) );
  INV_X4 u4_sub_469_U10 ( .A(u4_sub_469_n16), .ZN(u4_sub_469_n20) );
  INV_X8 u4_sub_469_U9 ( .A(u4_sub_469_n41), .ZN(u4_sub_469_n36) );
  NOR2_X2 u4_sub_469_U8 ( .A1(u4_fi_ldz_mi1_1_), .A2(u4_sub_469_n58), .ZN(
        u4_sub_469_n7) );
  CLKBUF_X2 u4_sub_469_U7 ( .A(u4_sub_469_n45), .Z(u4_sub_469_n5) );
  OAI21_X2 u4_sub_469_U6 ( .B1(u4_sub_469_n1), .B2(u4_sub_469_n29), .A(
        u4_sub_469_n30), .ZN(u4_sub_469_n28) );
  XNOR2_X2 u4_sub_469_U5 ( .A(u4_sub_469_n37), .B(u4_sub_469_n39), .ZN(
        u4_exp_next_mi_3_) );
  INV_X8 u4_sub_469_U4 ( .A(u4_sub_469_n35), .ZN(u4_sub_469_n1) );
  INV_X8 u4_sub_469_U3 ( .A(u4_fi_ldz_mi1_2_), .ZN(u4_sub_469_n50) );
endmodule

