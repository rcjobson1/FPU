`define BIT_SIZE 31
`define EXP_SIZE 7
`define EXP_BIAS 127

module multiplication(clk, opa, opb, product);




endmodule // multiplication
